`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
sSWLwNpLqLeR2hab8l6ZJrl3sNn3hpv8u3Ogl2NahcAavs5u5oCkrsBNdhU4mx2b
6gLDr2sgn5BIfcshaIQTpXJjxcL7DZD67Pp5BYEC+wCC7Gh1ygdTLxC5Fk0i2Ugr
nTrmZoLPXA/1ztg5Nm7iVq84SeL2GjiacPfDgwYwzEs=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2022880), data_block
8OyoJidNwRGiKrQ1gFoBSkohj6EEQOLPeXCLZskovXVoq9ot3VyWABkMYO8HBUce
s/ZYnC0SQLQ8qunZfZf8kRms2oNAgYXYT/kuocKUj7PzN9op4SUuYJ34EaaB2x2U
k4Pq0O1nqDkCYwnKguEJDeyJq5xK/6AT6911e0/Wwwx/gV0DT82/tkQyN18I+jn/
lZpRpCsK8TMBNxu5/XmZlScj89hd2u2G8HWdPkflZ+kr3hW7L9D4wPBS66tGbLGl
BAqyVk3dxdanIb1hHjy7StiQpQe2+eT9MccBM/ObEfXVQVaDSJcY1deURnZ74U4M
k30TP+LYM8gj2zTOqmeswbKvezaeUrrYaKydUAt35xZPcvgM8KKCFiilmhzC2+Qo
CSR2MD9KTNlf9gLbGfPmV7o47beVIvXwgunuJhNfqoojLZA6t05A/xIgHi8jADqz
hcGSvn7VW3iW5BajJ6gY4ofCfGMu8ALVfFLP/lebI+w2k5MmCqqpHpvXyQw+wQvl
MkakgFMuppmI0UOJc8TIxooQm8RuFUD/GZ1yRPN5Gm54m25+ieYzjlI+CT0o2GOI
H+8LPEsat4K2fTOBlKvRCtTXFyEhw7yhbhzl8ypXpgzDWN8GJ2rApZBQ3UWayhI9
UeUceb4NHxo3m7hCqOCZbP2xI5D9Cd5f8hS4dBMP70P2zkBRjgOnh7QaV4bnBpma
wu108vjiWtmK0I7nVvJ9cQ7WnZaxTPLUaPKCthq2uabdqxssW9ieVQfN7/Q1gh6a
mwZuJGuOGHaHf5LCcEvroLeeCTNPnu+AoXuvr2UcoH5VVksTlF2zmKwH40tgGvuX
a1uWJJPlZfI9P4216C++XTjvPli5STPsUZjNcu3uSwsUKUik2PfGxpH2w+bUPOdC
4Uw5odRWTBEo3RXFu4rnRgTKAfQEXp+Nk7wQEWXPShQknpnGAh2pAUhCc9MAkkUO
IiOsfFIyFHvi9KZ4/yV24c0tcjUEn0ZiogFCbVorqzGSSliRecCvx+pXb4gPxEN4
zAklBLJoy6mzFImuPEJhUIahTiTUfLCLV5kkZO66QI5sq5IKKlVOrlVNluRhh80q
Nmc58iOTwyVXjc1GDm8GouXNBlEbyWnw8JiZm2KoiC/Kb9aux7MazCcKG8IpH0VH
My4Uf1SJBehJo0GKOYl07O7W8vt5m94L8e1CSFPeeYsx1YlD8vp25H41vigZR+i9
ud7ADwO+wEbznb5c+zMc+aA97EV7h9dYFp2X/PE4tk+XWxdKWwQEKfXa58W8pvj4
FySugyLiuu1qqa13BvAeYwjWRr4lT9ErknPpJnWfwyY91uQmNWtafl4m1mPm7HSH
R7G3PNZrHHGXF2sXf+B1tODJ5vwvH+ehC8aUvgNgUJLIiiqNNeIzifkBS56hZI28
5iL88k2VGCEj2JQhix7ebkqFroVBZEUMTUOPHFlBCbyxzFwUyuN9AN8TdcWyFtMY
sHyYvI6hNYslNEa5Yd4ahFB/tlaseAFyHSDkg8y57zWiW0zPpuotmB4DYz/eTmKv
xUpy+fz8xMWLa+aDkpxTqZy/jqZEWS6GVUR5X6PlmAsP44I23oT8u8zq+nOIo5Uz
nwricJev0W3tmjBO0XqkhOhF6seBEj/QI0Bw76fLzI/0T06FtXVUufS8Ikmj2XSP
lPTEtQgqpw7O1FO7gJ7P8vX/ArWF7WWRu2IEA0yIQ30wQWuPOmfjKGlQXGgHDmJ4
KgrK2Hp0KaTzmCo7PsuqE3cTrxwuQ/h+jsx1LUdDLZLDHXJ6LrQsVRdHeYoGm7rP
exA/AbQzRAUHF3HuzsnRCpkuqw+9KKHPr8zj1PGpbgm3UdnEn9E81l8uU4Lem0lR
kXUI434RBo9lk0/6FdKcBL2OlHrnc9GWBj6bcppuD1GKFwuzQt9A9AR7KP3kKiZB
x5+fW2IJ6/6FehKWlwSGQaAsl656cDmxSQ0dG7T644+f31RGeqnkYhMH16PmYHTS
3be7zdEL9SzE1MEKSTvFjeQ+YgaO2GvyYi1xNXLXtL0HRAfjdiV14cuWJZAivlyT
RHZmQHvkO9mG18vjJZ7g0cObWvcwwCLWocSLDhLFFIofaO6K+/M7+C3Ui01vZA6m
Z+SsLnmNNE14F0BI7wwr9FpZhCW5H3ATpYHWETTfBoC4BCxGD4XtV9V/YiJGQKn7
kmKZnzMjDr2FlIi2v7DwUwQdva6wReRv96CmJ6Dtr649kaGUUf8ubUvFVdUAbT+q
xAd0jYoSnV22B2AJmsS7zW/WGDkfdkD5SU6wz1f0fsAlxEeIHrKeP0FC7YddBN7A
7bzGuU9wrPtnc3HdKOsEErS1g5xLW2f5Yu+59HGIsFjiFe/VANQ1EyQdiEfRX9Jj
XeJjrlKxxszz/6grQ3RCKJLj8oNCqUe0/aQALUNitA6wjWqkE6mNEhdb7iLr4lCQ
GrYDDsF3xu3d3v+tZNsGNJ8Nr5gb9QiBGECdc5XJMIRUb32z3YqNShCLJEZj9Pht
hq/ac607hqX2pOS0J2LiO6xkWu7ChgF7XekMb1KaeCbAWLF+WyPZgZdPYi8LB7Qw
cLauH34BlDptu9tC61m5SQCWluda4CmYNDatxu+dHPIqSlM33qXcgPyj8A3Wguzn
tcjGQA1dQlWr6+/5c1zrLpK8sxUcNzd7Wa9HCSZoh8UGwaHq0/oOTe0L5aMX8qHy
h3ZfYf6IfbRV333lccQwuCnzZIAbrp3kn9b8DCRokuj2tge8X1U3J8zUtCLfaR5O
fV8fncqR0CxPRgtwSjxbjlmINKz/oL8FwNGBRCfCbtegg9NeogqHNZKPu41VVryL
GUzJ0nUW3R3Kgttpxd0w2R/sS1iyeCu3Sq8lb+OugyvXNcF35bCQrByJm5xySBku
yiyB/SxbmS7dbxjr4/F7LLQk+mytJT39IK7MGL7Oer3S/ACR5FsU0ZD933BMh/Xc
mPSKeQV9fsZakZwn6sRQVITtVq6ZpV8dQfDOV5GrFh8HUsExhrWC2Eq0xsfzJBna
29dVEkn5oP4Qm1+w1UX8EHzF9Ux8ldXG9seQLQIDTDZdtPKeK0Y87bxlXQb8jKWM
iVEryetq6vupyWL8GWBpNvcOx9hGPHptCndsnX5coZYgJwRdgGj+qRLEmXe4Z0sa
nNB16QBbCqO/sb6lN1X1awIkoD7kPeZpWc4b42epONK/q8UP+vQSo0ODc4JB0E1v
1x9uTL1P0O71Qhk3UOgC5CVmcPBl2/L8FGzDL2O5o33T1kMVrZWJjWHVius2Dj3z
nqSXd/mdjBQm+iV87sFeiC6yGwHmjUhsiEoU4vRUuwLWBlIQeKLrZEmcfhCfVJct
HioCTI+payYhtIFAGgsgmRufA7+D2QQAcJIFw6iv2rwCigECRnswih3pRFHwXLAL
H/FIc6hLCNHh6j2CyAEMTvqlS5AIpgMqBU7Aui8gBWSVK6p3WKoQHfz/jYWGACfw
P+gNmsHpSuj0MwxQumJKFm5l+j7uhdJgvaDgNmFdZCRuiN7BZ7NJDKnk7UzZQuXG
9hjiuymwTit2gNjpQNfCa+vtHfCz0UFqiAp+WglUKG+ZAKNU4rvWiNqo+MqrGhL3
ojcw95akGyNBS9ujuR7QlUzaR5pxEt9NeMM86oD6bsdBsa+M1LvRr2Zvxyyuih4a
LBz0xusggVMTJwc018p3sz2N82HgOdNdvEjAughLuG8/NiWLP4HuOAk/qwl70kz3
O1eOXJcW3eAksP4CEcgcwWHIk6ly3UHK9NizfIkkoSuSj5G2KCJpdNurxNOSpiD2
oFEULIcGVSom5T8JLO/Rkn9R0envXfUoPmShola/6lR2LPoe3hanSoiu6QLU0WdF
au/uiibXyIaopYuRfyZs4cexWF9VawIpyAXQuRxmxhTYM0scG2yWBqga2pKp3YNB
IMNIxTsLz7MSOObr3jvyiXNsDNFkSyTa6SgUBId42jX5Gdg59VbuIXGmueafSG4a
5PTnwjVvZY7Buv9rxBuz/aCVu3ip50pnqXHTKz4S8hQwtVS7c6UwObA/+QxR07iE
LBtBR6HnMhRzh8rsMD7dl3px+AcKzpp4J7SeOXRks81vY8GGb7tCU3yAjbByl+mz
dld/7tshgd6UoRoVLFTWa0IdMxgedwRK5tKvvju/MMQyzbkUx7FD0NdcC1abttaI
78oys5PBztmqbzrPPXutTg6gGEjP4b3FlXHltIWsM8lQLRxkyA642bWbqS5AVQoQ
eaohrqHxbmAPMf7C36zdaRr+QqKfQSMMe+q++fEQIO7HTNL1Zb4Bfktkn0xTO5sk
LV39tRacXsjSUKG9E4uHN0xa0zosfugCVJ9sWJ/tfMwLA7x5X7b1LTjK9IYWY7md
6fDea+ZBhiREKydZ5WKr9OFZN+AqrkHfiMHyQ8UrtD7D8J2c7uXsUz8KeA3sh1Je
r5/0BfJwiEIRHBfHN7eHptlW6uti3L6fC50EvnIHC3FT6v+k9xTSO8P/8x0YlanE
8RqvlpSQKVG3Oe1ipmJa4P+Wi0DDB7t7f6YK8LcZxwIo/fXGDbKCiCr576DUPCnF
bN7SHW3JLb8/JDzm52yuzGe+PoWgUNNDsSkwhgFnErrei9WmQB886XNISWBJYZPr
dMr/Pvs56nUmLE/1OI7oXjDtkVWsB9Wn/gDUkWIgWfVJv+Me3eD9N+BLdd7Hn5oc
Eb4r3HtK9Hyw9cSgOKpiP1ZjFafIpmxDdfWG9zaKu7RN40t+4filyQcnGMp9YEQQ
trPG7BKQsMILANJm0ib9lyiiIyCF34+jUmwdwEW0EclnNZDQKgIaTl91wQp6Izxj
I/U+Y3OtT6BC7VMVe54mn/QsTB+EgyUWCftzHFUMUaRydO8n38du1sIiDy1H58nk
fl8UQNawsAmYKTsuCtEZVw1uOtwjCP6AMlqb6hjXxSB/Cr9K4Ly3vn0hb8OzNe9G
2GKU+lZUdnPFZxbcZ+yTmdVHupODPoltd5d7YyjT3lmo9CjUjVY3wgHAoYw2ENg7
Xft6NfrNwgsp4DmZyj23wM7RcEDvlaVbuqkDGRWxy/GJ0Xeg9f1wsmKO2WZHLmPa
z0Kr83OLmtYs9LYDHFuFAsXBslI9LrvF0T+MxUDoF8AyUo5eFHFUOVMghc/CGath
hCEnBJXY9y8mKSqj/pxuQbt4FzULj8sj4vrp5C+lWaWKkqkBuJ5LH5DJHEA2AtXv
Tz7bFYnJE8E/1288+AHBrYM+vjXXoyiEnY6Oo3/3WFi8uJfR+gyF4P5L6vTkMnu8
yuG2qzHBG2fuESl9pgNhHUBx1n0rX40HMAxuVhTVEom540A7iNypqsHHLAQvzZTV
XFoIAawyr6FeY+GxzaTAau0RGt5SAFHUtrL7g903ZVFfa4hgWcV2CuBdfO/qPcOh
jZ9bYUsljLIn1K30P8P9gORU7m6ALkDU8fTD5I1xda06hyx6qBltJ8AoZh0AoKfS
rAwMXD3M8/dE7GTXwzkSbyVCjTx6HUm4p/BEizqNcDR7MVO54vylLzWTZsJOb1LU
O3fgbWKAmAESjbupI7gkSbAiGlg7Uh8LadoWinoIP2JKWuUf8qlmZ4boqhpYcWG4
5wM46JnPFgMIzj8p0deC25jgMFsGceaHaneKxH34pe4cy8o/swP+W0AGzCCkDp4J
hegWyQmU5AQot0jiqdRuHyJvAs5jjTKtyBSCt6ZWLsKW+t/ATCd3x+jpsOrXcxr4
P3CxCSQQQdwgJbA49jOTZkRfucAA0oCbjveLgRNBDaCedHGSEHf6y8Hi1Do/QfP4
soSSZW6ogKszkE7ge/krG7sznxvonKyTP2ecaieSmn8+DyXiyZfm3iMlhwb3Qwew
hzyLAdoidKcjsPGvoCpR93dTU6nAp+6tP4YoX1vCWEqbRpA84O0U+/FRPvYIZyhr
masPVM0/RdshtflXf6Yd62sHrMCZEemyhzGylB4C1YF1pXjFHW9Mc8us9+g+bbf3
s8afIz5ocMcnFyVlFw7NfskVQjyHwT6LQfuVE5R5nKj5rx3/DjSIrnxiqi+pfSWB
ZLvu972yiEprzNpXu33y8BgbNM7OwLwR8sCMT4rNbb8AGsyJB3D+7pBk80230Vrl
3FPT68aiGrWQBFvogravB4jHP4xr/VDNCUQ4bANgaqqIpwCtClbXLkfYZJRXZAkh
h7i9AvFNtqDd9VDv0mLuGXw6wWBSDh+QJ9EQxOgDDglLEsJdgWQUwtaGA+5nOluR
GBb0ohkq4eWPk0NW11ofgDs/2qStTBj26dYJ1BGLa79IZRaVcOLnuasAZWKr3zv5
M9KgUSlB69lfEL8WVDxdSofqB+APsh8gk2vSfbhiI0mBHOJpSlzJ5IhzVgITQm0l
PWbS8MYmKQz3uGMWe5fSMmreRPQnyBwpkLt75HRUS4vwUScvi+Mq5CoPGssfYYR/
g9sESkWNN/k7rt8PqgTeUIJT0flBf+1ItPruZM0Uzf+/MNttkCZ2zmjdRY9Q1YuY
JjyzrOBVg/x0LZMy7kRWEfw+3vRxxJmiZuZ/cLGWjQv5xSkJyFMFtxtl5fRV7dpH
ggL9XqrKSzWFkgXdPgcw/lw5GKkopySlRdOBzhFVszNIHHVt9lHVrxvDZHQCYLrx
JqGtmyDX8lcV5Hl3ihhhxUULet6TSatTOtY2ju6kFYmOgtPG8LtFv0qKzj4GYKXj
muXablAd/Wo9VWNfM4wEDxbZBn8FDWy7+U0Qx9wmN8kTzQ2ZD5R6KdMivITu5VsT
J7rnteDKV9RrMcukjEwzWqv62lcliUX5R8C2VBQ7bQydYqtuwh7KUU7/s3QOpKmJ
DwoqMqzRiSVw8GZLaFAYYsFCcGqKihZg55NX4dap+bzAMInnKR9Qz7FrmoaEpMCO
pks8Im6E3ZyN7Z77Pmhwj72eqm2yVixM/KRV4xbiT+K70zAO1Hz8a5uVwv89It6F
1fG31QJ898zB5UyDua+CMM8pHC0XHGDQQCVw+qClinkMheD8nUbw6yCIrabB7F2E
C+Pfa7U8/hDB4i5rLbCjxKKuZwQkuJUuqhezZ6VqHiH0Qn1g2BQDaaBwl9IV5Crw
xaK7/MDmZ6NcBcbwlAwdEp0gvh7B8LRciErIZSt5ZXhvpe+ANRPlHKcJmiWMvQNM
7u6hFea9WXe7Kee5otvupAq7iiRzgHKBSKtl/rNoCbvM2q0lJ/NjuWJBy4ucaS+L
OmNIv/Q6ctqrDB3TuLUlrhXgb1shApaBAuETXHSAx6/qlTjDNpYFqImKxjE4U7eH
7cB3isr6pn128Igc61hhWzQCjXdJrca5lzf6rNT6oFBqHoktwtA6z1WX1AD4tpFb
r2CdFtSr9+Gh/ExN36zVzksW9WhSGhLbjpMY35iHKVQ7TQSO6PQI1w8GYIIE2Mr8
/FBioOA4g3+cUZvquVwbxhZy0IWAZCy3vmBCHMZWjfUYuq3+LodJlDgRNjnlS8Ml
8bozGJKAJgj/sqAiNdaVHqcOG1KWOJOSZ1p4Dhb5+5NAGde4316BAUjgBxcIaEMD
VScXZy6gMfdoY+6zEcOG60zI6lo8UbwtbyQcljpD77r4rCqdEggcSv593nKTAqjY
wGDEOfy8jrDfsSOOyOnejjC9ZmhwCk8z/WgcooGmOBL5JXwIhqs16QeF8++hxQdb
FiKIZuPMKJ4s34aAlhC5VfAOdngJtVoQAd5kpdX7BSM/7QuVDI89rIge9IJSJXGW
DrXAwFFA2hkqD5qLW1BiUlHHvK+xceeNzeU7d+eI0DmqNDxCwGwAx5CPlwbcs5v8
6WyacJ80FvfrlltA/ImkKeiqnlFgxmZfUvxuoQwjRbHAQFaJ9VOn54IOhcg/zaIL
dNd57SwfhA/zfmCKfUhxe1ueT03OM4KvRw7csXQWzn+OVYtXuc5j/HmPfgJtfOCN
XovkLim5dv2r7hHMQTvAWGXnZsVigU1mFkkdnXiXo+JxRpaT9SK2mDJeq8F4WAwp
0wWY3QR1eiZxTgcZrmUEMK9VGebmWZQDDoPuH8lW+c/HRM6wWT+5lK7MGMHa3CPZ
eHj+co2fVtoQl8lTYz9kHAOWNGhbLihSmuuG/iObSS/Y1shi4PSIVDJv1d5UAy7Y
AX77c57he6yENtKsu9B0Xe+lW7zbztbhRVMuRAzg9PvCnSnIgThGtL+3LLeO2tDN
aOy0oEb4lpiZz9DMvJl/uvqWvN9IN3jR/QMrW3MWI98JJpot1Zwu7/28lS+/Q4s+
B2IzHtslHEb+M+RlsLgSh9t48rX3bCX9DxM/VwW/hRjhwJqeTozbEHdsUQx0CFrP
NFgvPXpcfQDqCQZ6o2fpR/vJSxiSojnl9LXTuRrLrX+OlnH+0nff3C8ts9oDwn4K
DvOPrjcG1Hq5RYPekd8uT8v5NdA6XCKGThSPGTf/veB/C034yVH0vt515i+0ySiJ
k7ThOK08lWnsAgTc6qRRMx53yau1YDcle7gESQU8+oYzQNCRRIOJKoQvFa57K9As
aBXitDXb+vK56uzlZ2jonCthtVdZQiw70w16t+q1DpR0yJRwRb4C+3AcQ4Zs2Eyb
RjtnMEkamEQsCrFLP6f513SnWZ9NVLbgdCoSnsSBZ/zxh/f2Bx9fiWt8qAnbdITg
NEkMuLJMvUgBWvGsO16vapQb9VST3GiVtsgd27Ys1z0diKb9nb5sZl9abV97Q1ot
sfzuoQpzeA8plLcRr7hNqHLHdADLTY99bMvXtTWH3KCBlib0DmmIasjgdV0qI0El
/XQnMhJVUxwQge+9B4NoViu7aOLmYvh9LQJNFMWngpO3GCqWT+i4gNHaQnpkpQnS
hLjjkZz0vWVeRPBgYJRsJhmGo+S43e5LNXJsDLyF0EzCNR/gAb1lJLS6DODPI5U3
rhyP1TOEMw7BE56rpliH18QVVcMOJEMdfg6IVv90LxujjY587dA6VH1dtPtLN3Wq
09N/+8hrHhgHppM9003WDbHIPiOmEkOPSHBXHoO0Fqv+Z1PftXEPi6lNC5ri6WSi
cNGR0iqOP1qkeG6v1d4/MmAPf11Gxf4w0tN22pArbma+9WMHvpHU+3HAtAgSKP1B
jlByXAHWO1Yi2CjvXo/QnVTbJS44d7MCycE9N4ploe4vws30yi/W2GDFOpkeGKrl
FAtd6/VO2mmt8cTxLS4B6aHHSE7eBy5sRim8Btw8yMGsctvJNpH7nK5EHixfedk1
KhglncBSl6JBEKC7btH7KJ5GYJ9q2nu0rcyiRGwoffP+WGza5fmMZt9d1cOo4gl8
qlKSsMUdZ54prJc4au7pkVEPG7KLEugVtuNUGXB+FaF4uXdfDQVgh2XcPUEsAad4
6geJ7+02QNUtBjpx6CrvKhaLl3IjyemvAz8hL0JxkPC7BGq7G2gcf/7gi4dugGpe
UvGUZlvASWra+AGblZnwtkiy+Y086tU/aH0cmDRQrczt5yQQ/OlBMDlKBct03AAW
5k4RliZB1dhslVvH7PABKyWEQpfLfT10uEcUZO4VZQwvqfZm9JgQ0gsMb2fVt/K+
yvkgdGvDlE5dSPOAcERJdWop4D3rEzsoeZ7c+w6QbNWcCWPtS9ndvQZ/QiytMhN9
0GsWQgk35jEmTZjxeka+ODcOBoztsLQ13/bz8hHebnxSavgy0QTS1IjNkqhbOPof
MOLaCMIINcYQAjW6f/PMuN2Vt8pYT6kBTEWAWemKysep1SxKYePQkp9Y8nsU9qSc
YDGcAj8mLDeP4s8eICeFQOmfrWw3U/2iZaLC+ZYc+W2sl+Rptdn6xSJZKiEV90Pd
PJd0rPH8mmqdRYmmK4kkMEYN50UVFUIocEmiK0tJyrxO1/+C+OPiYvYsKTTkVqPD
YDaEBkZ+Ggh6Y5VL/9I8eu+2b+ia1fRqvBefzQjIUvA/FN4maLHtlkIwgvwiCkTE
sMoeXX9wt4OucuNsnFiKkTtZOPf/zRmy4zW1zdoGFCF1w3i9nKmOGUCcndmvgOfZ
vFqLIjpg0gxifvZgOGklxCzFj5j6Au+Jaum0oc7QuyCqfeXXEzARW9AaULlTX3ro
vPVcC1xw5z2n4YJqdb4xYT2vQZHZY8CiGWrOqkRhJCqbsn4JuBVto/+oVOBDN66a
7l9Du3ZlWWVuCeIuPKzxsXqOTiY3ouHSHIpo9rwt2ihPie4Ikyx7sexRiUTMsqzL
1EqIwFsiyncCxPdSlaKemnF5RG1DQiQOw+keXP+cFB46nmwN10xzbwasz62WOTJT
p3FBMQEdkiqvJp8oMfgIICC3ybhHmoeqtFis4gFoczSau429tU1HEGzu8l1wGSJY
wAxBHN5KHklP2BtPNblE99u7YyxGkQqFWd4YDOznGARzK69SVrucI+XOXR/tBfTo
eMENEr2jTphu19hGA+/oBUu7/YVKNPgYwQXqL2NUZvZE1NVZHob+r1MAZrxK1Evp
i6WdP+wJIwsRCZT8AfmsZiYLEhN5vF9W8P+YvsJkiwJNTTjXsDwO1/Mw6sal8hkH
wjftDHoTUaFOtogwPVGdo6+/6BWla9odDxMcdXIGnNun/Q7gIKY2NJjhPDxLxs4E
tGtD1z6CPv7L/wj9tTOMnKq9PpiZT2CZEiLn8dDIIz1bNqxdzwobRSEW740JBDIh
YIkO3XyE6kzY+T7zRAnH759goviMmJbbtr32Hk0v03aJlSvRtqpGP4je93f9auaY
vlaMgDorH82OiQisp77GipN9c/n+DHzdB0TT41G7Uvs2c74B7JAUfpDpBA4ggSJL
/J3cU0yK0lLIZYxGb/0Yf/Svntrt0tgmKeIIWxCMYCJRBNzGKmCmPXVGIH2R6Xx/
B7JDuVJ0cXc5Ujnar8bOWEU11RbaId2vlJYCKiZxIXuqLoYhDpKv7kIPywTtDipK
2hZOvN+thPgPMmMK4FERsHVjZZ1ZqVvluO1yd3OtmqZREMb/lF4Eu8W51NgBPWmj
R+jvdeoFl4NN16Gcb7JXEgWJXdMQlRLsUHa34VtmzrxvOMOg93ThAnDqtStlR5LV
mH6UDRWfznwD8CAOVCFISYXQfSYHpsXzrl+FSPhPHAwqulOJfUJFbN7cCciQaT6N
cfbkI7UaULNgy9hUQG5cF3nm/iWbVMaFk/BGnYfG30yOZOLmlZjIoqWD5PeXBSpR
DCtc+42AA/KY4adHAQV8VHF+9BIcgaQz+0YkC2ezFjEd++uFggX2WwwSZjDIN/Uj
lMdRMCSCTSAaheLvx0tknQyBNDzbVen8YbqZIdEWxfWODSz+s+Ls/Cg9Xcb1Don4
+VJJBo4/Y03rGJc57Vrtv1lwCyPCkogU/UCPHAeh4Fe/Xc220WAyCIpRy/9WgvOD
BwEqiCBM4c7FojhHxT/fxzFVXHtErlmS+FYwyk2GFoc5+BsuEB3hjJroH3E4BdE/
4698G07RnfRqw++CuYDzXnPHZmjakVMccb+yF1s/ezqcY5f+2E7iY9eLf8LSsidy
6gEszE8ws89uUdxDXHIyc3YqAsabgBtzIAmSxc+y6C+gwytDLccZpSpLMY3/KYCB
O82VsiWe5WXFFDYeuCwi/YM9vX7oBq5HwyEDZVjnqHF2dy529nm2eRwbezna/dXa
HpMwwL2tLTHl3nkHSG88GDbPPl6FHSB55sRdtxZNuvW4ftDN+1YfsP6LN8zIJaqZ
wXA8DZA5V3xvFMScbDEhcLJBV1uOiA1LYGoJ1i6TjyvJEYTqqu5k+/sDtDZXwE4K
1ryqLxzjlji3gyxUVIrxtcZhmn8mjbv510aa9RLRcPLn+x28lyzSOovn9lF9P0ct
p0BzaCIlC9P8imXoBs17Sglbe8e6UjsQ6UClKAfYXkeEiAucqdMZLpgsYT2RilK8
osT8slVobttI3X9tDlatu3h0prl88yXXKFROGJpPJ+RUm5YbMCLzFq1tJP11550e
7MzBUhyactbrMksW1Fyuo4XD7uSI4VyivNWLU/8Am5ZPsY3Vep9I8M66bYk3zLPR
Gvsio3gxFT2ybpyCHlqKA+R/mmW5mSw3nV1QFczw3OUd5RZ2uOhGQDgDpnUCDPWn
txq6TOG5udCQPsuE9kSCk/N8WUz03h+N1NoF22P80o5mN9Eh95l7HFGPSpTm8h6Q
7t+I7hzoI/IrRJ7mJ3q1VYDe0VXLoKqug2CV4uxjnMhRqeNt0ZlrbeAaQ/AH+xDl
lF6JHyb7M8IE+lNx6PIgL5hX/ITz0kGRgDlH8GbLTYxCN5HbCcZbO80ZS3CisPei
Rp8xhNinuFpX+5xBr0AG/X8fRIZc6vBYYsWlNJIPQFqjWRbt+YFjVzfz9Sc04vsJ
IoCfsv7Nx+a5pa1FmzeUHa5d97FyH3a6BdrCoY7mEu2UGnPdoxAh4+hUMxR6mdUA
JfTwEDVj93aucbS3fuHAiERsSKX3yC6n+1wZXwBxryu1iJsb9Goo8L0HQM3wA+Q2
nrCcy1uvtizTegGQoCJScQNemoJzE7vT7rk6Wu1OwtFYQypD2di1OCFq29QZRHd0
/QHqNq53bw6a7CItvqcSFSxXHFwvgbBb5zSQLzId41MtMeqky6xMDTAp8cztBUpx
aygJA+BDkf1VjALONQFYXLRRHIupqPOIlL1KCz3KCrhf1wgPqvoZlm3RBtE2+76t
urePfv1wMYeTjkXydyYF1xouXavGCyvH7kFp8V+NQ7teXLCzo6h+rjFTNKI9mEbF
IvorZCbOxjq4nlzbK2K6cBs9jUrTroUSMT6D6B8JRIzq9ZH+UXpx0N+U66dRCwgi
jsWuTXw0CBCrc2tAyHpGN3V12lNpVJ6lZPEi85LAL489KwkrpEbADx7knT0Pf2Ew
MVEa81a/dXu6ToHT7+EwYyAQRpZiuv0Ytdk8m8xxr6Qb8c3kRVD1jv9YBuIxi0Lb
zK3io09ZTnPTND3gMf9V1VUVxAp4mm6A9GCCc36wZKOd0BKCPFNKFKzgo8IzhGig
tEYxS5YRYEprhoWQTEDcXOsjDyiaMjUFfHrKtu9yK6EtH6Lk3NIjYUxer/8Bclll
4/hHRnaIUkUBIdYKDDC/5buprNqO6TdPZA0yWpyNTV34DkfG+8aD4sfDX882eHBd
Znb/SXZAagjS/0o4c32l9uf8LG9rL34aPk0YEOapADrau+iWso1dZsbiNIc13RPu
nIIrgj0FbQpwm2qZe3FnxHKlsSw7vvr3eABKaSh2Tpbzq6QG+abbRZjW5dqlQtw9
EqDI5pMGJik/Us/t6FLj3QiuS0MIAEu+oef04mHKUhtNB9YsgAO+Zi6S3dvHnj4R
6NXfjdDXx+vE1QE1fy+FStmLhtDFLJ0s/YGXfQKxEOzdV96NV8GpqniDwTMntLpL
2MYnwlj3/18l41f86mnL6+sJpyTcepY0/muE4dcriben21wZHiaOGMXgxTQwZCIk
owCTRYBYd45Kcfugf7EhedsX4BJ7yOuLtNLTsBn1QisJwb/hhVBjVzYcTHia/Dum
iDoT2egZwej6oEvLe9HT75qZoBaHISI4HtLFPFcBleFv/GvFzCVsOcOrq5MWRtFr
9Fy7kLyXDW6vi6iAMFa3dnL+fBQEBtbZmYwiayAFfFAuuhVoWkc+x87yzaH+/5jr
NQfK9GEFkvZcn4bPRSKoMfZ/BTKd6KhrPXqpJhNjB5hbPeoxeJShR3BQswnQ5AL/
8+H2yKvQhjVf+iR22JBJU6KbpFlDDZ2fWH3LucZZOGsaz8IkzmORmWcmIIdK9ENs
HZ1F8Kp7hiPMO9r8ZBQOC8CSRPaSz+IEWtXrtO6MB4eL9e2e7L5SEuRGUljhEf2B
hcAXuqBMlY/AL50a8CuTobny9L5xtf9DH2fBQqM12TlgLygxS+aO0RNECHRpcJ6w
Cnr34c+ivtODlHVnfqAe4x5T2omGgSVvAAakwM74MAvL3Rzq2Jc4eELR7gGSrb1l
/y13QRQp928enCq3LArRoZX8l9pOY1CWQXupoOx0kE0Fyx9bm693PbWJsOnt/DxM
86iPb0GAHX7+DHypcIWi46wWFxYY7QQhsiNq4s++X9juIsPbVXPxas8jQPnArvOV
go6S2wAk49olgHJttrbEEYG3Hzy+BuShGPuKAZlmfaMuEck2AlVLJYVi2At9NB80
oJmZunIM+K9KV6/GdCW6T18oQf0Od9bQmQAjIE3QG52foBGqvZUPFkYrKSw/vX2z
4TDPX1R+Cygm5BLUePAIe3tBazpHF85pBRRWeYMzULBRz9eIJ43Cb/pQW8tQn3Np
L1vJg24rZmLdmHXt5eucQu/v+5DNPA792JPQhQfsZconXSoFTa2BLSsWE0sDVipL
I6iEZOG6q7x/p72zIPnVx6YoGnaEOefct1OEIpHv/wObQOhw+KZxJ5Lw6wPc7IEV
kf335iOktRQFUIQGehgUxkCe4OUGfoP/ToKvC5t+hYI+nkTfzRPi8cdj7HGFa6e8
EHFq6FmFXTgGM+vBH4GUM6oI98J8l9FC7EajTInem3F/YK5273uPCD2LHAaBjtwm
gv/ZNB8Lsf9ykwYVu1WbXf6ObPjlE2InU2eAdSfjQLEbM4VZCmQb0UOHF7ofa63H
wV8QKh6Hg7BmDW9ffzsXS/pkdWryemOaBwYLz1zPAPu2gcMWYB0JSsdFAiogZ2p2
SSxrgwtDw3jr0dV1wrndqiWv460Bp3QvvXqrh9ulft2FPhVfH4NixR1/VAk+FOhl
GiQAw0bjQhBQ0WAUzndGZvnjeKiexTbi7RjGmaugQYQmP77ki4ZJS1ER7u+yKOHt
WFCogJBi6ZKeYfAXvCpAVNc1MtWeO07cGJHD4bQ3EaVpghYy7BUyp0QMHLrroZHQ
KfIs6qLLaUHDw7d3ymisjwX+p46bpJ7yUMWHw9EycA3LghR51dQSCXzY+qLA2ICO
MvDoYYhiDFy4HZ81RA0P7SYeO9QRZZtI7PtY7TJ85K01croYi7QkcgxokM0WBf/q
a8mrYHSOWHkAR4Z06I7pEbG/79B1ujHhU4QaQmHWGgJEE3bcnsKhSi3fBumPaXn3
yz47Qb1WsfU8n1EFGSbu4aH6kR8jZHZIwOLScAkwmRvNlUufrzhtQCGNPxgRHSuX
rWKC04DJnKzEq058wTsTI69nfOuj/C8SBLHmiJVkzwakI/z48ms5A+uPDpCi+I2N
832QMhhT03oVynDgFddUf3UqV9NSjD3+RtbPK0h9qxTUabjdUpZbotuNL6yymH2O
fTFXCbHoHJHRFVu3HKLP4xbc1B8anN0VrY7KdIpyZt8I/n4mZp7AiP+c1+sWJD7g
wsAKm97tut48CFXcIefTy1qibu1FxZZNKQKV0nxBjaWzwBcsS/afGMRNasRyJBOX
Bpzb04422SLhhSnRRPeVCIhYEw2LBrK+/l8tLoOd8ZhxY1QUL5DrJIHG+sS8fo1G
oYiZqMJL6hp7z7KYERB7DmKab0sypsToEO3Li32f0tZRb9rZVOY/unh44rCh0HOh
7wlhbHJimCjJVNOnHmZVJ31Z1Cy5GBCp7BTXzDieIJAIxk+n/zIqvc+R5LCkpRuM
eJ8T5IYStzhw05rFQ7lFWwICqWkoJQFPT827wH3xZnit6oopuIAmugyXGNGDqXfN
TGyTOiEGofUtC949xbUdTC0IpI6Wta6BKD74KpU0VCGJXYn9TRxUK2kN+79Qid4R
KgvX6ybroRZ7P6slDnVEBXfjajPqy3LD/1Ck2C5IBB6oLgUj/eXFM/8b6AeyP4oC
v71Pgi13cIZNs8Wnm8msgzPQ/ZUa+3fdzlwdGFrulG6iPU0Qrv8nlzV3O1sqPkJ0
G41FryYROQNzZnwU9Vf+iWNHwlderdvqyVd/vBS83xBeZVgkylHy70rinomM9Eac
yLWnFn1khba2hDJ9bGJYaNMYcsyR4gdTjN/68kHhWLukTOGnZPEJ8l18euOoPk8P
lT+Ity9+RHWqacYSvrkKXiNSSNYW7WBm6enYTMssdsB8x7+aBQT4d5PCLSDgaT/y
AT+JcFb3Prp8h5wetem98Tlq1Db4fGyb3KdWmZDdHshIzUIFn2eD6xYnIRbIZE4l
qQFle+Jzzpvjcv7p9+97YyiBBGsbkqrFf0I1KPsR04Nd5hrELO6DsCQPvGb6vI3c
hxfXJvc+U9j/TiPD67iPyRhfJ/b1FLxZWDh5X2pwPDyVFtRdsFgAPOn0v4G1Lbs1
AWjdxouoo33UMd0jEQn9JgByLEh+3G6McdnhWbFooq0/xvYLKWg8WakAegOO0R6j
+XDSZ9NItAhsQOFo9F+AJAT6FJOZ+//Tre5Ix/SV0ViIIMPr2DndBUVLVAXD1Ejc
xSbgjRcfYw7yKYVj+ekCUMp3oKkvEvvad0B32+2VAMmyvR28HKjAGyqlQgCDr1J3
O+MEPnNFiFfNGXarSGheJ+5NcHnOyk77pn5SUDsoK37nRLsaKORLxt4CRBS4FwJP
w+SPkpwmU2FxfTRycXRIVMFk+qMdaivM69nDucZvh5I6+C8InIe7nJx6CYHtzsur
Sh8n7B3rqpkuqRhkPiUJnBCveySnXtwqacmXpw6230IWWvZBlvx4lpxIzIe4JGzP
G3/oJ9V5Druca0CnkfWMO/u33mN0HtQ92HRA040Or/Isq/ZzOCipIZmmoz7N8Yrv
3D31W9N4GCNmaXurjzyXW5JhWk+nJud3G4bS3lo+UXcVR4ZsxrLIWyY/cGGpjExu
vbgL0B9lRpqWOnyr6ZqD472whiejlf+XgJ0SP8SAT8vx4gJMF/qZB0zd2LCQPuxy
cZ2ENZm+D9tzpPI+QCIehe3mLtIsFnNuzkBQTKexH5krTkidph999qCcvIJkCc8G
I0juT3pKp9vlB+UZgfDdTBx9/iJsqL9CUPDZK8AO19X4b3CmmE01Bip3ArDH8PPc
80ZGCxhJGYaWcIHeZTmrb98QAo2QK+nka2Xs+tm/hLmgWecItrDycijwT3094Wym
NvVuWV610Z4bZgy1ovRxZfG9/i7QQdqygFJfRdQEYRsTsw3wso2qzNRE1OsDpqOT
Iq2zM51NCC6r6W7VMFrevITGbvpmYncOUx7e/DVTB95hmbUA/UakacKhGwPujgHS
qHHtn1IWS1UN5Agb4e1co1muVMbPVyGi5VhA5Fq1bz7jFkfX0otT9EM0qxbGzRia
c2h6jITtm3JW6bNUV3jRNnsn+eVWSQ3HxCZs3Pbp5n3goReZXvetNgxaT2Q2d2ks
MHSvGLJ/zxPE9M8XN2wsAj6xPYbprdJFw5TCUQLqiwDPimdhUS94DZ9w3i6nrwx8
y+bDGhgS+AiOFmxiLZ9Gx3HL1zrfSlLiPxAcyZz5DnEMfG2/xOqqIXCDdtWpHipo
uM6CGp8qBpPfERsmQZT+0BIBsfh4v2/EbUJlf7wAB0nIpAZbGJROdQiknvxvUD2w
xpurnTQMMaHWTy3Mf76mB0nVnGFxLLjzOtegtL+wj57HAeu7b1OB7FJ16rGELYqC
HZhhaqnVaps6GhkZieEoNIY7egLxmbjQDSjoEH7B8wmTfpbbYWjRX2p+rkwl8nVk
TJ5bTmM3JYKdVnkL7tGISre9+CxJD/jtMk44Fx7BJQ+jneVxxbL8Vymu+x6OVc/l
vCgl5En/uZD1jPfcTvjtskB/2KjCGMpHlQOvEcXu/xRBzo4DAf9pHgoD/z25Yk6j
nEKlHzaHGpE/zb6gmObLNH/5pv7b8eawxgtOcYo/rAFq/EbhLRuXRQG37oDhsuzt
0r29sq08LG6kUuk2+8BvL+NzW5/msbIBxRWJB14adi0cpqIUrTRNVbrmBpxMB+pA
cQzcICod/g0ESFMo4NTiOAnxJ2IVzshDRWQADk+yLfnHHdk0hwCtKOXHiKbN0d+Y
fGtNfUI75BzHm1G37uJExINJjFG/b9+3x5jbB79U/CugV4uXPySZeMXfTGs2CocY
4QyPsYK0SzRoNQZXqByCdpDI2xFykZ4tuvk/R4Ic2y1OzLlH/4HQGCDHBR2qGYJE
AppWmgH+ZvMdBLJNS3GH04JyfkEAgCNSbg5Rdz8ZwHeXkY7SV3wrIMN29VvOLgxi
zcsaEkV6FZRNQi8NZ8WAxSRhGj9opNriULqKU5FdzWfG16HnSzHUB0QHsY0uWmyi
jZfgUufLFBA3BNRPPVYGFcqa8ltw5p7iPUQyyuWwxuqjZgyZXxuOYHmX7mX2ADA7
8RIs56qrY1pEN1ZrzOyUxfy+dBrAJYgkWwtrLS3VrAR101qwlRyUBxEmbtVNQ6SX
HSznQcH0CYszOL1dBeBQXnEqwb0eqJaBMot+timCyebzSb76X7SlaZ0M6ENEf023
pTWeLvY7SXtWvGX2NRflD92vv31PVwy/Q0TzY911I0UQBiG1zxq/2EkDct0ZzlQO
xSn+Dew/9plwv6vDAFFTlZzgNKsb6eCpSd0VCN6gypKjEzNhvlehJohyz5Ki1nYS
0vfczT/VH576ghjpXRUZsHnux9ldaSy+VDioTKjPlCWXeq2pa4sY8QJt9uxBecVY
wY67GKlMEnECNW4EbN1qe011tNwkdGnENSN3p7KpnlV1DCO9rlVsuaZbMXyYeCYw
xyMHGVCa2WM9yk4w4HOfLilqd3ejR03BEeH+o2iqFN9wjUI5m/QeGz6gQKRCAz/c
Db7RYGXT5+g4qXIkyrYoQ/TQ43B2EITivFVqvQR8e9IP669RCkB4kEAiVcZmz65h
VKfwL3bN3aSUZqi+ZkjB0UiObuJrpumhtfTUp1zP6vWNqXy5SJu7ZFpaLlmi64vr
xdbJfcMgzOoyARcLtTNkVg7mHrQddOw5a0G3KbkhIZ2HN3lhGdqALQLghrF0ilNk
hPS3+nVCg6LnPHZ/0bag86vKqIO8uiU5mSAz9/12zvHlNaLNrLgywiLcRpUVEk7d
KTgpBmKbJ4SP/rJ5cWfAU+82vCQdEHBLjHTvlKG37hsSLDC423A7G2ZBxmMB9tiw
xjM64RK+sAWPey/uvQENmkzJcSsYCu8DOqlRBxSM1clcCSeOjrFtJm71EGUCoegN
6C+n9b19dHJFaZrrLcHKpIctA6FFVarUvIgh0blKJAim1GYS7ldMQA7Nwc7YB+gD
RijgqHzKrjtkcFZ2eGT567Wj30dQ54yVKwLwHC53ej+nwYdzfZXwsn9lsuEQsvVs
nrIsrZdVLFJZdm2AD/VoF0rNemK/cENtQDaS393T04LZUins7XPWD286o3iDBTja
eTXAxs/Qi2J1TrWgExMGBdlQ/LXtJDWGL8CbnOb63mCHmDHBNGtQ8Skusv72mDBb
AQcEPqkc/DcJ+NZKb4pFK10OjFCDVvlMbCncdMqthDfSJtfMiw0Qm204CJFoYj8T
X/QG0a1UbMqo/mldDY6cXA69d5AzWlPKcqV1JKhodeuPM80nk+DjobjcbLhb5e9w
ZlBfNvhJLfThVyEoLILEDYOC3xvwe+tLz8WiAg1AGQl4CZG45o7Qg+AbZw1HxLpF
ArH+cWksqe9xarvO0KbLh4T3txN/gvXGTV8c3tsZXmx6OyoeppXdh7fzYGE0z8gT
2KYocw4bZ+voZfRicXxJKOHjsRyx/L4dSrkvKzGlyYxRc2V7exlh5NpLuJDlgN6G
iTUCUOq2UNiyjtIzHqdtotV/XtACpfrQZkFWkJKTV19TFbjUo04A4GOagYsPHnyQ
dSAEysAQfp+m77EVBB4XS+CI4KNJhXXu3wehahPrGdtOOjKvcLmhoNCTXNcoDcP4
W3RdMsOgz7sp/Hef/L4e2Zr251VjL+MhfYo2+QHzrzkn/toO5/1gVZnN/9aO1Sw/
zFN/pl1VCZXEnK15vg+L8ZM/6bCF8sfOzdRC8EUlO12jIUeZPBrURLfElM1t3Pgt
nVQNln48w7TPxpbVZTqyvNFKIguqG9A3dDhNvOa3FkZjGVrsyFLKv1f32maYU1WQ
EeDtVjs8CAkxKNPTCywLveSfQpv817j2hUf54R61jCJDS6IxrRSgsGJjWsb5XM9K
MJVyyv1DWYBp9T6QU10gtjzj63iYow6jYjfyIT98j9zksc1YAV+t8DndNhpaG+Bd
mXPJmd46oTSgjGAYElsucDz+gc8oDTT19Z8lDX0sL0EO9HzuxvzMDISTlD2mKUZO
Oiftv8bCgo+3suUGIQKA/LhTbqokGsvJ0zNFsRW5fqYg235OAwBx8GGLuetpynY5
CRxwoWShuKD9lQjjyZmyfNBLZ7GDP+BkjizXoDEg/a/cEiThR9nvdUez6Iu7rIfe
l2sRhASjq/RBXEg8nTcwpwHt3STUrYtT/O6B97b3FtnJu0/q46j+Q8v1Phj+XAHV
maPimzUnJjwVzBG/2SmHnSnRZ7gl/9KPI+LWpzM3v2nFh0qAoBmXEPXcLJ5JcxpI
JOYNjXUotsStbIozFes5OtjsKTcKofBuHqqoc6MSgnH4YhXpy4Jqu84C3sdzvEIz
C697XMJud0mN3jmWv21snjAMd9BPF5X9CnBY4UCjwKOhug7cb4gfJeF7HblXgMXO
wxRrsmJ3/e2kIJzav1RJUMWuqY7QNtuuwvD8/BzLszk2q7btG5O0bvbKZH9BO6z8
qcLyOnUCDaZDG2Ua5NL/JmVV+JXD1PF64svt3Vg5zx97ZFLjkpIcpR43VnuqiG0o
KxW8mHl2ypMfz4FV8Vrmox8jVaccXDfaumw14FZA3/8jPt+JVMYFikGWjvnwY42P
BPui/y85T6WFJdv+OoLyqE+zndeNXSykeacij+KD0EfOFfuZBNRxuqBIu/19wFkB
9xwGNJLpvmDN0xfgsou0tgb1S++F6jUECtJtO1km1AzkEIWPC+lvmnuxj16xPPg1
GSDsk2P2fXNe6vYa2xVTu6QJuAjMjQ9aru7OdM0hDtThg0jhE2RNAsmUx0HddTGW
8K7m1C/i8tHuzfVtfs3i26IIUrIqvwcAQYZnSZhS3VEIrkJG8KB5+Rrni5pzH1rx
6fMTmfXmQSuLV6ayKlhqjGY8t70xCFpIPixzLYr/mzgPheWU7QQY5fPPN5JxQK82
7FEU0Vt1RehUdXE48dpHDSaWlT6EX2XchHK9bgkOtDS8Zp8Mz/dkXZ8Zp/aFMHd8
HSosQp9rW9Y7xf3YJdwPlgqxZfGsgWCDsVT1qlUIoBY4uUfHbzsqLGGs55kt1DX6
6/gOe2O2WxW0TgGKTkIPdadycZgNLqqbR8JiGsgzWN9oZ0CIkzwd0YT9dyLPCvUb
j85bxNSSmXbE9Dinj9Sah5fYqFfv3W8FpLoqpQQ9/UfJ9BToUFqPKadKwwVa63u0
R16WF6tW3FIzWGcZb+G6y4TRIXeG6aitsvjH8PnSzoI+8NrJPAWCvhgZKvEE2ng4
W9AJbTrbdoHK2njR2qCmWNiLQtK+xpOa2R0Bm3XPLORAunifNvv8DUurcPdvln/w
csyBMJubG7JwiXzO3OKxnKnbvmITFvUZd6FBCx6ZOv5PEqt7NJ2bqiDU1Y+50aMT
6G5KXHNwpGkAyuNYvMhQTHRQ6PlaWWNJ59nFK7YCZ4yCsvPUo7H2Q3FwjuF1aKoE
AB1xn+n9IbqrxPzUll/2r/havHYJ51Yhij+jv776+1NQEreYgJi12E4QkdWoVnln
pwxlmngnPKSVTgZ+z1jp5Bl50t2VHcXwnmU2ssA1NuPmCqH7pjFV5qY9VaamCeOS
7lFGcUi7RfbgZjrPf8st+rS6xXoaOySD7WuTbjHJHexLs2nfY1zwORJ2jk4tP8ZN
WqLy5CJ3EZs0zLLM+95R9UeLBuUiJpS33yUX3OCd4U6VnW2CCmumXHPtemrwdpWp
bAvCH3V8iewj9b6sDQobJvk0Q11t6RDK0Azp1nmoBFM+PBdIG97HUUTr/ufh4smV
6tCC3t+O1rSIxN6k8iGRep5KvTHxZys7m75xoDS+o6a8eJ0Opjd5UqEB9isXq64A
dFRk3JABhY71W0vkBPT/BemL0s4dlCEfBmsU/7joNqXa+mui4U3Dv6tBqSjKa/Zb
SBUgDuFvJxw5y+819xrUD6M4vV70oDDBpY6Y20DpNUzkfIifLQJUtzQ1Hu3fM41X
o77f/YlvcBOwaFhNgYHM+4X+5D5fKezZ/GaXCzTu5Na/8IBmi8K4EAS8yQ+SokVi
FDS2dxEfu8FMGEZhx6QQXJYos0vewriE8iG+n4oH2djEipAMVX+C5hEb0ZBAHBOe
SYd29GwGreYX7cLYxmJ7vxImp0+C9FXQy2t7/ycMdmsDJshXUyPp/ez5fKSWJW4y
cIU8EPlID0mVwqJe5nI9xtu0KX5ZAb9griNKzkt+uafE8lfgxKCwcuMTUWsvDVqM
5SVjr73YdgcAEkab2wXSPC6rldoFsYrRk9xWj52+XqbQIfuhz909FEn//dY3I3+h
ZHTtdevv7Is9vsL0N+34gqisSW026ZpXgKMIEqnCqL6uWCYssLKT7PTBeUanPAW9
YZFc36lv76P9wHVAUbFc1pODN0sK/5K/W9fwW8uG11mrOJHHbvg6cjqgvHiDWd3P
rXmLR5GkNdkDylpZVFEsZWzq2l4fS660lDjwGT2ehlsCcCWLZoXUV4V43YlhFq2E
EpyriH7JPIulG89sF7NysrN+U5LqbP4z+r9Ouz2YkAnBLcI0axcNWn/GMFxL5suv
VfvmMCnSi7VVGJpnKmSG2b54+0L4m/pVc9oysJXxPNSnid/nL1t/XUhLJr1uG1gV
AfxfTwg3ODOZ/W2B80D3B9rZ6gsl+6T7rn61zoIkL0/JCM9z76CiBi7s4KdxpxKT
e8tdkz3sm02rBoEzaMbn/DLP2COQlV505quPg+tj5Hq5eMDyHv/T+hVTL1CFapmQ
NHbhHfTVM4+uLCr2QV7buc2+LyWETelZShP1Pxd35LXWc2Y9qwoe9t6wigDlthOA
DJ24Yhy6jE3tm7isP9GKeepTJTNxXcjIk0iZYlN7qepezhVeTdczbRF4nVYiJSVN
jRHRIm5QuM3X9oZVo5SxrMASAco0BpnQWavEAmnF32/ckAafRkOVpSzJqSqFKub8
9ZluYT/Jjt25Lf9nKGVAw6dJOAv4GGXNfN52Keza0sd5elYSMzFJ2KdkC7LrQfeQ
Gg/R0jWiaXlolP0P0bUzuWZKSYbUFkR075e1jns8XjnZLOhEbzB4QOd7kzYrmM8J
AHtDOCe/19UQ4eW++QFB5+U8seRbE6M88M8YaovUn4WwBV4KBbbGzpDnFEwxT/XK
rNB6hIJ9rsGpDBEeURPMgtsfLsa92PpRfC7zhZMBwtqXK5McCrb8EvgkOSUF2+sa
n4gMuO2Xjw22zJLnYnJwCXdtoB0IDLnZmEbDYbUXjrLMuS8WGIt6s7lGp6uqjAIp
GkC2bzCTc8T8Lc16FcurGBUDyRegiOH/RGqRKJwDWx/Dv7D2AvbhdaqrR3WkgW1x
ZmOpHItZcBKrqox15/lwQuzQ7WXRx1PlVNITwbO+HgQsa79qs5SKurDjdVREygdC
FHjjt2BovOhUOzxSus/06llPT1IsagrT19/cVCnKyVDQHm4JIa6iv/xeTV0P833D
w9gACvt1oOllUG4ZBHtMoGc2nIS6ZtxcxBWAZTuMKjw4Q98N50DDcW1ch0mpyi+/
KSwFUvNEcXn0pP1d1EyA/XrepHpNp8kGq1HswLfQudJ4kVM90jkZUI+bMGWVqzOB
FH1/YK36aMC+IENyDZCQhuYRie5UqHq8l/TGiGJ57k8QXlmwvv/9xeHxLg49E1iY
kkbN46hm5jl5pRXl/UqgPk3rHJ56G/8k8uyvthnMH2nseRSp7Yyp0DayJKVwLljt
jeKOVZTghPEbr0FQGemazMXE0RKgMZz10ksaSyF9GHZp8MYQAwoc8pOrKqVtoaTJ
CDluUKim1D/sX6RauTUsfaOZa7f1xc+0COHsJaV5dhY/biyoXWypdxXfF3mG0WG9
RIVBLGhmWwyI24JXR070YCBKdZPFh97jBqtF8hpjXpLaz9oCu64T1Ow3hpHtd3Vs
nj5Y1PlM3IR6wjGJb9LYOdCgiU0aqt3UsvSgPSZ9E1JC8YNqHNAaB6WGGOdf8fvK
KcC2nvb9g9pInElwhetCgvj09/YVFIj4ggxADntKx3SO5N8okTBwMkdeH4H5ihAv
mtkV6YE0v7jfmDVUZ2ZGHnYRmzn19IRzdQoHFYasNIqBvGlYQOSRAF9kup+bO9Us
ZSXcznlHuhNCgTAWuuA11f1PtViNH20k5SxNXN1IaaQeOoDwjedrYyO2v9Y1pZR9
KJVAJPtyrgxmAPpQbCZltD7OPZRP3hBh8esMqzt7Tk03GTAgPYqh6+vHkChkf72w
Zh1s3x+1dOtZrutKNEU6ifC21pt0TbYLzJaOulSx89DFHUhaY5b+VxvcZ4Llicds
omlfYuV+rrkJNqLRC7pecBMBEvmsgU/h7FUk3jX6kWGCDrIygNTgz7BlFqiLKWSB
yeaOYjImbynnMwhHfJ+nm1WQobIn9UF7PpUTcqpbGpgVTLF5dEDfjMeAnBpOGryM
bPaJhSqLstUT4vdfYJrL31KFDWNGXkgJxMhdYafbGSFggXrkpRSJLU05HF0xpRsG
UvXMjh2wKwqf949VHPqh+lTXhg+s6oA117E1WbGjda9hTmyqM43XdmCE5buBcL3H
1wqB36UqIuKP1uNqOSicx5SKEKoH/Lqs/O1mdI+9ZXG9iGQkQYCBBGNvkW9ZWExh
je1xvx1QeTYKJVfHcK49jvX+Qz65f/9HvOQvMhCmaTGnrvFYBdfFa0TcmA/lquG3
Sf316Jd2R9yJvQswGhfsD/oEx0SATQisjnrBFr3mWLQyNu3+tpgMOh6Zr+neDEFD
+DGOhVg91oQdCKVpC3mz6F90T17eviW9WPF1My0ogOptrBEVRGWkEshLBr8p3RHv
WAu8zXtok5RNH6ETHK7AvPO6RcBOpbFNz0vGhUowWLXUUZ1X56VKZABtfanKZV/Z
7nG1s4IdI4ChJAGzBfMeHhtSPXO8BFzo5jaSoPHOoY/+z8Ja+tneHHZLz1ypMJWH
uEXQozxDIUVKgUIQIfsf3mOMN+S8uaDJKHj0W8A3GPhKrLToy8UnTw4EDqu4vRR0
Z6zbDw2m/DTyio6WxFbqv/vD4cU7GV409uueQInhOOINujt+Y0ddfOLAGn8sXv7j
MMc6dJ9ToZYI6voXmGPvrr1cEKawVMoBgiec2Qlln+rrk00BuQskW2GqqH5yabUE
7WlRcoOMf2YHlZdDRmxJHuzAPaA6+y3Pj8405CpH1EwnlkziMjD87XiM5VdpmRYo
XLloV+K91hljc1k7HTbJKLoVbFcuunYKOKWTwXJBpYbLTfFjwtWNuPexrF6npTFW
WL1WCWYUa2Aqi7uWOnq4K7lZ1ATLet6BOhqyWqhKJb0VU0eVCPmiaTSArU/rsXVH
wnzkpuCFfzPrrX0qLn927LyiiYtS3HpcU5XXR01RWnbObT4/f7JfZrgwE9CP39Ph
SoBapefM4bUf/FVpjwBlRtII6pQVDftlASPnWfKxZVsbHIv0NWY2Bi9y4/sEUdAf
0ySKSFDRIyZ/t8KM03UJKBp7K6tkQigAMXKUPuLgchcNiQqczN+MCQ47D953JZbY
9cZWzfLlXxpmLlUeacSwWtvB4wynpLKLZKEM+DoK9hI1odx7eEL80kxLGmzCLv2B
XB+ziBPFb6xzqxnTmsdti7Y39PglE5eypnjkasqtTqYEcGuLseQ5HRGtlo5id4po
4fcndfJ4vbba2e0LtitB20mbmkuJHsIKupEOW+/Z4g/4U0J69bLJicrXG8uhgc0e
gY/uVfZMavjOFMQa94pS/WOOLXRjuiwfbru3UPrr5wO7p2nCsTmNoygMYf0L0FC7
54zztXc3+Z+RoY6byemAZ2G9Q3lFzjWgUGhOb6Y7vuq5ceTbmL6ZuoP9jDxosyUk
eDSS+uVBMhTDmwvD60/abhyYqtohvO0mWYktDdUGDEV5CSbWFeEvegJ5jI5ZZ55h
Sur2VNwaET131M4+P6WlSdkevEi0YphiWtBZL9y1J3sNf+8WNBL7n+e8FBn8qn9G
pSoBQ8yMldZVhGiXVy8fF//B8vy25Hd1SBeZz5gugKZ2kaW9VJkjTYwCMuJ1T4ov
GI7QeG7I8DkQyRQbC2LMBj8GrI//QguqT8VOUW58naFz4p4vddiasrBIgE1x1ZOY
L4r47LkvDbrkBbNqmAl8Fgk60/lVwAYeDEK0udSrxRcUXWzeVvO52xXw/8FgNycF
pmVnUYsq8Rt9289nztxhpf/2RCgF/Wkv17QAwJ8ZQIdrv1qEAFUN/KzBMUI6Xtay
yf6wPOjCQovUuhyLMruZrYLiH3sgzUlAQqOKvRoP7pJqXCEZ3BWxuov2mrd/ury4
1DwIYGgiTuc/vEdMwlcBVf3ZO/eBBwMp6evnm0WNJ3qLAw+ICaBpC6aH8fmF0yCH
nmv8N+mhElQPtHxcAdlUJQkw6urJDugF2RW54cBzHRdMqyf8mRXAKyXEsDNC/Quh
owxUE8L9TcN4Kba/VzSNDTa8utJ/OasMFCXIjHJWmVD0OfLWsFkKnAVg+9SJYzWL
uFBI+/ZAQfaRzr3OtDKJ3MpOSFTbPJ9Dy9biynnD+HveSlWopbLzXmB/3odPdSNL
y9TqFwGK5GPoXlYs1l5AqZqeyWynLYYATDFQ4/0ezC4l33Jz3a4kSeuTlGQXKrfh
VhJ5sz9rUoh53z2FFvlbynOCH7IpVTZVdOIPxyRBK0L4I1Svl1RGqZyasAEgCNLU
oJMO5dtjs0UZjroxBQHECWLpFYaR/BLGpd6m/DTy++PijUKG5wvj6hAS+72JmHEL
v9KvDxT9+c1YshmCzdYgGQYusPn3IKCQI1nSIpwQ0XJZCnftAZn80xn3OuNstnHY
Pw85KCnDiQbLUGJ2Nd/+qpKU/fHjR1+KbWPxS6WsvZ12+ch5kA+BRvVWV3EtqfXW
BYXli7D+5PjX3fGP6PEWPLXDpbVNC2mnEDiF78thMrhW12kFFVgzOXzkmu7e5c44
zYmuGcxmrHT5Yu2GiCWnpHdko83ef/4SdCRtQw+1rpJY5Cz0OBp89eFiWH826nQR
uVCuFYozgz9cW2H3P1LPxuY0N+CkvEOrGlVsXyWQSiW8b/QW+CRYUHCG6g6RvIwd
Fa9VDzHfFR6RDEvqYXvYSBCIUAjgTO0bCQeiw5YbJUD8N6cccZbH67RwKomUP1hP
oZKXchxxw2Ons8rkJNF+FsT7fl4Xm13nTNHaujOQ3D0nGLv4lUdXDgFdRvnSZq2K
pUgAjGk4KrF6TJL+k79BACAt7W88GfWBuh0fM/9en5yFSKzjRbl2HrbnnrzpA4qc
DsspSnotoiEHyAMu2//dFGHcH8Y/6yIQQ2PJ8AhwZT8y1IUIMiSGLveQEX48NA/1
pgj1CCt4tbivtr4+UzAonJUv4fUOzpFBja07thk60zJq30WY7hlGGlCh1QoUdNHK
tJFfhaFy2GxhK18exlh/x2OLAPAy4oT1OtpdqwsL9h60nvRPO1e2/be7u520iQ4R
QVT2VgcT8q1FChL6NSiCFULbSH/a5JpW7FcQ6km4fe+3PnQ2I85t3EnE671FWo0/
14aqkZ8vYCnQNP+hz5Gi0Ox+554o+Kl3wR/Wxnc1KKyKhmRLzyUpq/fHr5D7pcOE
IJGXUStH+CW56STwTVTap9ojAji6wr5VwZWAv4WG3nQDFMXzSI6dv1ATdzrAN9nA
nB4Zf519nwM9ufMmpzre0/rxwOUlhpAnal5TCJuIf5YwlD7jAPW8MX1z+YFgDeyu
hAE7g2HzJAWosIMJMrVexm1v1oee3PZr5oNlg4aGhh00bKIln9/+Nyfbxdvi6xxf
Dr32ay+Kng/11baR/1lVoJpIBgeO9MXJLiMgRxAun79jhAs1c7SBbQULGty5cZVZ
n3Pix+h4OACGU3EKqFQY8SI9j1DH34gnqWZ/jA9v7QQl04McBPFN4tLz2RCvGvTG
ifHKit+RTOJ1l4AM1EfD43o49vfKwWBKQj76TJqwicSIu29husx1PBmz1YwNluAi
yiHTufyBOR9Cdpo01sg7c162+Xi+TkmXZxRFh9FojKbzFeQz+D7GkqLeMT9uIWmH
3XN6N37npP3FdeOtnirWwk/SOygTj5+qNhXFuyQoL+71p6xtZVxaD304+f8jBw48
81pvLL9VVGm/dmDSgWU51znVJuEVaNKIVJaPrywMgauJTahi/UvJ89HLJ90sai1h
gbl794rcEi9e0K/D2JbcjCz5FC/vnBiecklPjBhJ8HhjI9hQZ60YQpU2TVsP1Bzo
a7yemvOY32bt85UdYukePQNyNZX+hMZL7BHyPwXY/5yR9y0uPkcOE8a9HiOcnOnn
CPtAgOu9gAa8dJRV8igSFHKqDrhzwpbPhGOOcSNU9flAYE3FteYr/XAs+Ipaf+Jq
ZXPDMktpamT8HzntwE4FWntq4CYmU/XJNLtkfCVtPnygKHVLfF3kTTATq2mCtzhF
2XzzOWPC/UCsviff4osfkL3ldEDuB0WynxxkPg1YyBxVobwlcQm9KSojLBXfomnH
veqoNxkTBdFp5xzJNx1Gti8ZOFWtykEsSLJ6GP3hwylU5zy3eNznQXuWMokCTwfY
DMVl8WT2zmmAPWwnltvzqSZupidp13ErnNKnJX7jNYK7cBD/rNay+NXo+p2srQS9
B56gNdN8zxMxZ2sLXBuj2D95vs9953hh+glKZb6JJUhTaN7qT9UiXAepEPWDYeEw
UROgHlkDF8199jZJzZB8+ntLUh7UkeqmIyGKrz4ERfPLWovdoBU/yv4Zr4r27D+1
6vnbkHJh3o0tJKlnTLYSOH91xdMEPKwJ18unzFXBer4vKFuq1fmVUlo92g405alJ
CPemstmd0k3mDNCCAHR5H3b7xh97Vumw+vSPu9yP57zxJquASLylJpvosZmh7ZTg
DgsCKigTKqkHJ5ref7RFou49NNfmFA9QueQEqdK0MLnIhS2pKfWt921MowQ/a3o1
OOXDO6xhx6NgW3ArRZmf2h/dYbConLqNsxjv2oO7IozQas6w66+TEJYj2cDxcH9v
IHHh9QGKypcSlkGNlY4d2msmA1KQ6HtWjDWR/WKnx5ur+xlrggPJA0DjBEtnfNzr
ID6wLgZDfsuVaBqDb5LhON0rV6hJTchydYrmtJQr5AZWW7RHMQZDqYA9IM1PHi7h
hDdDxtsGhzGu++mRJ1Mxrm302OQVe2l/tnJx7UxCmWrCq9JtxrHArwgnBzgyY1CT
9cv5JEHdBTivNfoyzF7x/oj/gK4L/zR9qgLb0tAyPcKBc3bKdus4dIriSZ1PCx7i
dg0ZsxFql0tnJH48af8gNjzXQtp0NKv1IQOMmIZwW5RVau/KnBaW5c1hEuvrcPt3
4L932/TdxnZDkspZmkBftIlDi88EPKhgLjfVoIYdJnXUVgR/ndz+r4j0U1uC58/s
OY1tV//qz3BR45XC7iAmq4lCbfIYeOBLlykb5ZKzuNJnw+6GxAY3btunMiwFXZ9p
l2oS4JeO+nMvMd4H9xQDb11OdHz6tjkpddRwUtGFt5HiTm2n72KwDKanyaSQxZ1g
DA3nIFoEaxMdWKzCwuKics9pYnc69AcnsGnWkIXoO2jEq07pHP6NFOlJfnbyK/vL
n2WZLBOBO/b2chXoJMIbTpRYjB9+KClF0JgoIB7THtC7de3lJ6r57P0P5v8D7T+N
f5K5EIh8Llk9b5sHF/Wooja8LW3DVDdeZltDczsN1HjS7dh8t2b/I1f8pVmsK5Vm
Nz43Ryz7bqF054ZntR+spM7LPStoKrdhCD3uj8s9vZakzLcSejkKiDXJXTVCpKd5
AwV9dyZhLDjrusCiuL4m9Ok14yVqDVliQHs38qtuPNImD1uLQnRdac0LCPtSLz/z
sV5f0gouoqlUY6f4UnVVMAMBCObcDnNA4HTIDO5O+fU2dU7ka7JfkirBXZNjWvOb
Vw7LRXlEiAhcUZj+4Us5WJVmyQ9zCvj+U8YK2c9bKbCmzqe4RHO7ePd5ibnos1C3
9JyVfvPSBpDJrw7ReKLjuLPS02KTfTDYTo32DruYU4ppFOz3c/PWXa4wTsQ5pvze
GLcjk+KJHdSoKKH0NuVUKuPNNsh/APqw8vVyBHznfYdYxVWHetNqTcoWUk3N5um5
kLGxDiIPo/rYZb2TgzMtb0kFkKfzYWYDi7rU9wnAqoPTldDdnapY+VKnQcAHWmoY
ReRBiTFdYcyWUeAGcKWmWAiJPsQHWDwVvZk5g2eRjy7NHI8pG5CLuwYvFDruarCU
N2T0Fym6j5tc7iK8xep/9hzuOAQhrEBYKwyjwMqWNECzfSlnwWr9KieMwlrPJgd4
1Ddfm/e6fmvD46B1yHgub+cFTPwKeT/2WdMmiE3K49Af2h+roNNfcO0OE/NNMkrC
EVIIPqEGzT4d9yuWrU1+OdNw8g9SOxa20u0PgXsZSIp+ho1MQwBvurl8Zp4mmkZh
cxSd7MCDuMbH7aC1YlkEnlJ2qdd+FzEskpLUjoPRN9J68H3VwfvBVkULPDDMGO0K
SWbx0stUxQ3n+4fz3I9GRX92lIztPVptsOoongJZrRywUb8YLR4XBCmuA8TVCvDy
sB+9h9tt9LA0rQDcKqEahn4NlVTbP8EXYEitmz7jhpo1y7A1bo4tI0gHFj/9HdOg
cNj8yhTIv3Q/KPx8wE3pFFPV8fZvXoVjKfi4VnO4K1WlG+JLpxzGRsiUl4uG7vnH
ZsBym5UJ9hich75Et8PABd6EVYX3EiUWWlzXUuXrvGwrOFrt5k1Tnv+xvl0jcB/T
OFWxX2f1NpdrBGGf4VVnXsUYACEZZHSOSY5lIzCuovj4dri6TCK09y38OB2hOofJ
MgSmw0rveIoXI5DOCAtGhipvyv8xAul16rdtrkKLL9qNewijR+S+0FdbkiCS0KNN
lg6H2bwYQNkCssOKjMK6qtI5lKnxk+P0zmIy5KlAufBSjTNGP5mzCAWa9BSpQb0/
Z0rt60Gz1ErLy/JfCom7tr2faXV3VrY2/OMZ4re8tjrg7IvbAZ46VroW59SgzL3D
dS7Yt9v1OIkYG8kb70mBd5UCPyAdWbgO83Pi0FnfQ+BQhEyDghPbG+uK2Y4zlZc+
M+PEvVw1YWXlULvuOM32kpRiN76M9rEgZ9YJe8kA+nulpH4jmY6mEWFHFCPHN3s+
X3LIFJJoGeNwEfmOuz/B7jM09k5zMtEI4AQku+BrdfqWSPZAKVtS7OU4DGN5Wm9C
85nYY56wBle4+/r1OruZ4WntIEEjFBFpmDipaVc78NCYqzWthi3ubsmNfIPlYWPg
Nwtadm4KtXQDuCEytamAdhbVmnbrw4RKFcFHVH6cwXHCGZZHdGpKSboVNcNnGxZ6
3I/CdvtfiSiIenveGdzZ7hXDTRNLHeAognFf8mGRmfj/4HChw5+qLZ0UM8dZcrE0
0/UPZY7QrvHMDX1z3JkYXspJn1KbfBGup/pYuaxS5URUa5nybKhUn7pik249zPOh
gtkVMGVHpgk8QFF8TGN7NJADq6CI2qrlHYAZ8B6dpG96YIaMXDTl9H40FOFvMtZ9
Fa7bdO11eWNloB428qvC0S+u2yxZGe2gJ4cRTR+IcZW/0iNp3Ku5IxeRl0mj9FDw
9dLVSqbk64vLQ+M0DUXbRLSfqixzVys3bWndX87Ne1qyXbt3AKVBalnBavX1QjPs
4gW0fDu847EcRjMdWLSnH8hmOoatytWSAwk12EFn+OwcDfjwL1p/yjIl+Z+p2NvM
4HOADyyaPbt3CX+FjYK/pXuRpXloasJ+0oxqHZLqH6igO/pMVv/LEzUZ7FQmqQNG
iipOeZW2JH3ifZEaWilhxmLxwh1I0gPqnhI2kpzPKxNibWVUDmjOdYFfrqaxR+32
Dfr+3St27DnbzHV9Ecam4n4MVqozPYx4NCFJZT8JEYZoEEh36BXHwSbeHqtM740W
+m+tamcA2W/BAREkITq1ECxjiBX6FRUvTqtp+O7+Lbg842ThRm2pVZkcoM+DK7pG
cKZsCY82tKKCrTEcVb764NMrZgvpXZr8le/ivlM5GIETRvwlcBCWV6nzGZLARtfY
A2evwhYc25OijgoOVKPSJVKNyb5oWjmVVOcBIT9BK85CBk97vv1Mvb+3eaCXEYX9
gOXdXSH3L8ePaNRqtFTyIUjuUgx5EPxdCqijkSQT33D3RmytktZUSx75XyIRHS4W
NwM17y03Xv3hVPoUOjFB+niZ3mTgZeC+MSUgNweA4LyXnjdq1VvOdKDi0kooj/We
yYErmAhimwMFo/iK06WqfMf9kghCinr23d3dyEo3GqAkvFMLjJczo6cNBwbUIb3A
LBFbUYMc/UBPz3xG10hhJChyGETyl1P1A5kpJ4aB3FrwEr0s0WP94/xIE3g+o3gN
DDqJh/PAG7uble4SJ5dBxUyhumcElbx4Ry1idL8RCQCppM1aPbC/rtmt4oMNoKSK
JnY719puxkPEWfYrX8BID1eeUYSVOBC8G0Jnjb1WdBYwIv2e1wCDEJmWLpJiij/J
nGpwDx2oKSEIL5R0mDdVGlZJcuNvWUGKn7ZpUOQ+ERG4CKqy/axW1Fq+BB+i+x/G
KjAfMRFkydmuvy27868LSb47osZj6Cgu+zK2ZAOkgpxjLzZ3Lz8cfaZbqLbDguhl
wAlZh7Cr4XeI/+p2C2QtbegZ3gI4ekbN2JyORiH+HJzkL7VEDZT0Gr742p2iH3mf
VzH+MespaDo4OlmXH95A7XEHKoYAQixG2bdscZbXVRrWzUEi/+MVwkNoSpOZGSCI
4yPUAFJ3ZFMhPr4u8zpmyhdrZ7eJ0uRCKTusYlGljM6gpGi6O14+FgWBm4dfqKUb
PBEmz9LhFVlaGWLsPbECZHMkYaTKMVj90NbuCr1Lj6GYO/2J0Rxn4godtyxTjFD4
bcN8Xa6bgJCf9cfnDZTkF+WyUyHpAkOOSYYQfj8EeCMphUEEl9tTXlRia9YpDQCK
JuqpTaqW4XjE8UqUtuhzXxTF8oH5wKYnQe+Ih57GUbQudMiBPrwdiVXWsBTl0p87
h4/roggL/gcy76Fjzbk2XYNyC4o0Zl9yGVNnxaegdIdu07tT7xC3dr+w0ghpAEfb
MFj8J1517/UFcVa/y6rk7rN4k2oWwAMuBarCSeiCH7G4EQEAuzJNalxjavs+wr/D
KZjuEjrJUTUQ6DU8JdS87LA/pxfKETY7ktmARh0zLttpBdd/EhbJw75rvZMiqCYZ
kQD/sTXQLR1CWVgTMEjgT4J53sfCD0F0f8m5IyJ/eU1/xlsBbNnarXb723Jz0ovW
lgnUj6jry3wVbtH8JQMbUJeJO7J2e5TdPIIa+7rgXs4KRum5ufvOlOU9Kkhc7rPZ
PdMEO07/5T4wsUitnpL++mX18ysW/tswA6cLWTA7Nbmigmq16gaqx5/VnyTfBTUJ
a9EGFPhGqzI19YDIZ7zfAemWvrgTiXkucvqkFeEkBK48YnksRtwuA4afB8iFAmSN
WiFOqWigl3o95MzrYHQNwdfbfXcBAt9sZ/omGZ68R/ySwsuvpFN3qRDDvbJIJdFO
nLIFoWCyzeq2HqcSK7grjerNQWMl3MuZZfmlreyfJ7jlsywO1gK0m8JXT+asPZX4
0YNDnhsmRFC/fEjpM/6WQKs7CYFS7swET2fA9E60mplcE/nY2Vz8drx46Z7HwlA1
SgvS55btG9sK6v3+7MHVU6E7y03IFgtgwnL9x/tSozosAaA0yQgYBut/tOw7N5i9
VBUDwyNVh1eLCFOmTCMSHJtPbmWjQ1HxJKvxFinHXBmDraMo64CYp1Y3XJgQgzPq
hf7AeE6csbhwq/r17bWtIsZG5tJ6bsz5QzEqyhMlzg54HzJjhO6WfUfaKA2/Uzqv
UwOdMkBKAmrJK0k7QbOTOS07PzELT8BL76VjIUblms2zG9QU1iR8yJZxBz+pbKQW
D1+g4Xowi7csxPcOp066gcwCeGlxgdm5kJENMnSAHHRcbDTCwE2Woa+7zOzwmwGV
Ay0NU5n94tXZV8NMoMY37L3NyoKwDw6sAW4+O1alAa/I0dZbSAJ50n3LG9q4U2VW
S8wMdNMgWWxargT9ZumL7pItfCivcKqP7hry9nSxSkynfUY/8LINizuiPH8HZk32
EHb5uCpRwMyKmPZODO8y51hg/owIb+CX+hMRJMmjhDQwHwaLJ75qsArVPKU5TiOs
Va4mpk8E07ej6waFOVBR3ZUAmtdPuWLRe7K7RMRSVDJVyBGE1/veCLq1INREJ/Gs
SS4v46DW+YU6sX6xKzR7FkDAwSHhpC1vdWszqwoiulfj3oi7xC89mRzzIbnetJLz
+rF8CgM6GfxKyGWiomtePU8ny/6HlFiXum8kR3QMkmA8S5aZovATCKSqSmtFOI/U
nb376JCs9Ul6O2+xXBBRCx+3b47Cf+MhL8pTcTPSRTktUwuXfQJ1Du5Cavt6mgXX
1TUSE/pM7kgmPAoCwKa/J8r0vmUDPqxlco21OWBZryFwnFg7bpjOum6kAw3edVtP
t4dJ1KsW58HeLSIIhJJwD6HNY+A085YZgioA5Zv8MNxfBf2vQMUKwViZdDfEGCQ5
3huDYyeI0E57uorq4fSLdHV+lof48wvHzyWIPvQ9ZVsYxsWyZkDHE4MaLbZzpuxY
b/XRHJ1gLOpzKe6ZZTKSNkcTXLVFbDVYZIfkHwpnttnj39BGL6imUhbX5drbpFIv
WiCGz6XYy1LnEVtdLBT4hkfRyJH8HxGSvDiwFSNN98rAp6umY2Ezs+86JxCT2nUR
ySxL/OhOQ73zRsvTsnzmdbjgx2ISaga7AlE3fw8Wiq8c9M/9Z97YndPgsi4ayEBx
1g8jZIvaC/oSwI1sT3vrFAHs5fLQNWA5hrA4Ejxl68BXDfWHOWEJwIxY8NjKn5H4
kXv4/pcoFdDDH8JBMrCW3Zv42udfrpXmPg7eLwkfgWOuNygoAkPPUNYc81aseZc+
zqhlSs0quroFxFvhofnmTmrUphgiw6CEQ78uOocsjyemrTFntUZWCqLTj8UviWvK
SK/lBp8R8pQr1lOQY0DKAo/e71NrMDhpINmlRMXCqirlQiD54HkF1mWDWt1Js8am
uiVmqHWzc/A4VH493UoVeGrHOLh/j59RbMNDEAethEHVnfRxRUuRLdeUClgXuj4k
X2+BhOAcHuIGtmBX1tjUY+IU3dbLis2c65edQn6nH5gJMHyJV6lDJO5gCAGmlWtk
nhzkfJz765wZopyXFBCE6rKBE5o5jaBR4A5K//meEg2xELoIFbsPHFqFUTQIi029
KjVCHk9zuWIEFqBRvrBDMRtwc4scwTUqtuI1V73PHSrsCH+iUG3qP/QY/Qtacw7e
qDFlfyXvDRJE8iDSqIcd+RJjcWzIPRchj4+Qv227xIKUUtbC6xG5AtX6ae3G4XEi
ZLXCNsaJmEOeNHyPVi4xXJDefjJ5iJ7ZpouGgoDluMVKsfIZ3341nOCaIB67+UT1
s4+I8J/Wo8v5aWg+S6leP3Bw5l7BSqGX2IyKxLbqZjM3oa0WIDkceB4ZAzTQ73AL
z34t3faAH9kyZx7SvB7xKhTudWTRsM6okfH2A3NjmN9JpbfSeisYTbLZeA0J7Bhl
Xme1mCLPzYKSCXLrm6/jiK3ueIivniRF6vpekVQTJjxHuSy3LL3uRCaWUugf6ccx
9C54luGwxXQFPS6N2/x2skTy5jS76m3f/lZZrI08DLQw7lKATzESLW7NR36mURzE
HIzDbjtGrnxMw2GnnvloQbUYQKyDMXuaRYZhYDPXQlHULLDwHwMnCFMiOui/bZbO
9309Fgj5KsPYxY+EyXxsXVoqZEc/TCi5IJrjByH0QUPb/mdJVYmIHDLhHqKGa+fm
qSp0VtCt2QhARd7TnrpfX/iPissoLCJ2+a/hybxX3ZdbOdVnR4NLRFxiUaOi6lRO
tBiIk9AymMJesfT5HJkFw+8kOeZg0Ddse11O1A6xg7fb8xnV5gGNeTpwRUdlgP/+
my5AXgKM9Re83GMQyqFO+k1pyB+vG7fIKppMgsYm8SMWAseY0GByKi9Fu/aIejaC
hLpvhCAp10qYhxseXm1AYtJMWGd9OFMWB7Bd9sXFBt4POf8YDSfiP9zU31lLb6lQ
qlB/MD4CtC0546S+r0006MC9p+PPVO6ejs5Nuanxecum6INAuHxdHq2SUjjMfbF7
KYv3kfoPD3l9TfD0M3TNVS65oAMl6+tfmPNoGdb+gAN9m65MjZluM7Nw3S4bLZU4
SFaBWMLzsUx6cnXQEFSz8dFRcPjFLQne+KswIEdLlRLAu+q8RgXmjvpgkdcz2pSP
SxVEV9iw6cnxw1qvtPwyHCrK66VyVChTzFjamELPItQA6W7bsTMHWsOojgI4W/EH
lqQJ7queHksqLlo+cjat0xvLFb7B+ydB6k20q7oHGxDFNyekLfLFzKABd0gHJWOP
PMuy3cdqWDS7rHGege2htTjWdWGzm1v/mLvV+HYWc8rOzP/E3N/WZzZgWbWbsuZC
SKgLtYDRRiS766S9WYvR2iEXeDgGdDychmDOHaXac3/1dR8kNh3ezIo/M+b/hCLw
mSkyRJMmkLQrEuGevskJ6K0gFKeG+Qv195d5JUuj3zRzhfpMzKGZUOqu+ag2aE6t
WiEB+2xzOh7rWWM78jHkEN3J6WJkptuvv4+L/Er8+My0qPInKme9mEU4y4S4dhW4
aZm1vI7zn1yhHd9jMjrSZpjPM0tNefFwyswm7Ty1ywYRdxEFi8Pkzyj9cF4dq6M6
QuGLPUCbUutA7F07Af9ksqOxZqZXT74kpPIeP2viRiPtEyQnbkID9jH59Y1hTiwV
pjIGEkLdrTxd42qkKGqnnd2gFXpsqanwgJt0tCWPfqcgKmR97+qiUN7BJDgTm+tp
J9EMac5ptVtFIPABH1unN94ceK66OE9upmQVbp7VwxLmdT/iZ/mXU9E72TnNk7QO
8czFPLubFo3dBe5eqJ//paOyRKXz/cXnjmeicg3vH2XPkPnrd4DQgR8u5H6QRvSS
8EYdIwTTijRmuvTBaE3K7p/nU3yKHAIZYg0ODoYCmzriCiAKpkSmPY0FoyF/bA9F
9Ly2PUtaJtqpdXGvwFieWPcFSMFT0GpkKn1FedJzryOQy5Gpln2uLU+RfCaexBdT
XRTUCQDjaLErrSh++cFxyE5rfkg7+ttrKP8904SIYniHYe/OE9nbqPJiIuGUB6Hd
cenKX+18kov/zE+HT59Lg6EPaifTjJA2DO9iDYKzOjXgyH07f+xedKJs+JvR/wmL
1V0KGpgYp6g8CTHQFOt1+0HFurOpqqSM/m8fdI0P3qViNNrn4On9RoVcdhXFvhp7
775x5S+1Gzhu31PDBQtTNPPNVDO3OAz36Jermo5sR3O4YIwMkO5s3kY7DiBpVgeP
9+9/+GSBQMeAX8Hqzgr3q0tAJ08z1w8nvCSEUyQxwE7hCIdS09hojSRSSevmihR7
y2rCV+QRNE7p5+tvr7SMw+7mvMOHHICd8x7ivvVlugpxqhEgi35tEkGCitzfmfIt
qYpAR3VslnXTsiOQ/rn23QVDs0WoE2wokrD5xAGkIjtF6uJkJ4uT1vx+hw8aYR67
pbZYKGflLt8w/+ccuWvz1bmLZjHjPZHC4j9u4B7tr/ZIkYdzHRdQyUklEjhbSc5O
NDrEyoHkf1DnEbIkc+P5f0Vjj8DF22DkT6qJ/hAHtdXRfVOmftvf1y99tX1K+aBE
rcms+tFPREeUq0Yp1eepo0uVa01U1T5HIe6L2fVhqfYhXWYNLWhqX+5LdB6tXoDn
O3j5GEij3BVigxd2TC1cWjeb1V1fjFmlaqGwEliWDpFTc8tP5lONBLMX+PizO5hh
EbcPW0jqXI7TR3TcolOTefBUJlzrZouV2tIjolInizIEvFlDrTGJYnES7Erx7ids
MuuPBCka4IsOV8XVr9pXn+YAbYPkPj/i43GOTBllcPGy/suSHruED1GXIQ7rpazF
gvjOSIM14o2x3WbedyufwVzyCqMsZ8mXDTy/Oya3j3oSK+EKmp3Qpm6v7zrR4as7
JQ6HUufRaEXBEXAa7Th3VxxzjkmWXvW0pqHnGf+JpvqkYNlR6VRPj8kfULSZWmJy
rF4Um68pmz7mSBIgzWpie0uGpd2jlPyQptk9cCZ7ItZCZZ7FQS5fk/5vWnMvDe+W
tZJzEDNi7np/kQ6zEzKMD/wq1oS3F3FjV35aWksVOF2Ztl0w+mKoy3JPr+auOsZ9
3BJ0mwz+mWUviffhrhhoRge6efembC0FzAWNlMBChhQynwtsLCoWOIs3Y8weUDJz
QVdmkM5Nb6CUaQb68zS2W6H7QbzgqZ8mZO2/BQ7TEIT0Q2DsvT5LO8Zx/9q15JKB
AzSWIy5uQQHiP3yw4YxhfgZjbPH9eylI7lO3x8U2zf9Q8oSFlcRmyLXNHV+UrhxR
es44IrN7atvyXoO2W8okKjmhorrJO4T0bLl5b9xHb1nHw8dtvG7zEMb7jVCHtY8J
o8z1LV4bVOZWE3zFc1oo6a0EAJksvGXinrm+/mY2ZcLW0g9edVHG9MrhVol4Ouh9
WLXU5+Q+HDMnWhpKkIIopNSC33UU1pqK2ydeUWk9i7NrYmJ15kn34SH0HFKdOlsV
Fr5uRwpDVzdq33Bz2AX7nyEgscachDJgiJ1+YMpnH3bAPhGsUuk5CMGWsa7edl+X
hW8hEAFYj6IUN7jDUcnD4NydiZGIPhKTfr4ofk5TdQBUl67CEckSyCuKYM5M9LlB
JynG1CZsK4brf5j1xyNKepvXICAa4GikAwaxBImhzCdbim3Vcf2nGMRugWBKWemp
Z4/v38gPgGp7NvSxlV+O4rpta6AbgR+b6+woikgI+/B7TRrEeNjPqRKE0TiIDrKz
7J2xoxJxObIr190v3rUUsc1iU9jAqBsnBB1ILXvFS7kLSGEI9DIJBaYWwkaytBAS
aW9kgmQkHcP5VO09/gOigGr3OWisem/ZPjf1w2mGjVsYxI1pcwndOVFsehaD21Th
cCugjrIILIEmrIeIawianPJ7bNPwXV5rBARQ4VrFaqiSRauZJTZ152FoUusFe6KC
AFOs/pSdKTlkFB+aSPbFfk9uqfkYDA0ip7pZyB80bQv9hYrowNoGbgmSJMqkyINf
GActfLlDuc2yAOXO10ALibY04GZZIlhP73yyZG7Su3BAOMxvQFlUQkVYWP94SQG1
lqfcS/pBPXidDjm1z6Et5cwRt7GdvnOVs+0FksvgpT5LYEN6A6lSpVegsKmrKzRk
CsZF0UVlSmkpLM0nH7hVhBCgowcHHbWZi+0YNVWZEsCWUrG6Bc9fD1ZXfPdd8XkL
YEWtT7S8hWy/M7BYaU1Vl4mwz5rSSvYUI6fDFuLL389O93DVQSMIfEUWzuSzsfIy
+jTI70euNyCEEAYHQvGxdEf9kVz8bJTFZ9IBtDNsiuujeIKfqlwhBjK03DPASjhg
pqwl4XUD+nk8BPdvstOKDrlUbkkMg1tZIqj8CNh7lMIJ2Obf+NmNbShzAFvUHPmx
NbxYRmCH9s+2srjJYPeYXDCOaX5bT2zMdb8uJJFDra7RofIWYl2R27ByaGafSGq0
ajfN/CJt+IuJy4yydsacJHYhbcImtxsIlvSeuqE3qbhDJJXHaFo5I/6ff+wX8B/T
LquakTJq9Pdf8CkIR4ps5h0mhckbz6sptlBJOH5uAQg4tdvrT78AqbCT0xg85Vuh
j3JePrIV4o/WYvS0Npa9RSmHBK0OeL0aun+Tkw4hwyiY66aNnqTgtZQfsfaTG/LW
KzdSl6cn8ykP17lJu89MiYjiSUNTDWlEZ7BWsFbvLYPlkXOyrJDxr3P6uP7SFMqb
2z234NbuqXcNleahWvO9Gqfx1c0MqlMg4O1c5AXKYSMwsRUENVJkeXFFGZSHXlry
9NL/vPZ6mJZSYdACCuPkwSwn5RLNBLLEM1jiNpliCNHixGGW3Ic3RVqiesC8LSGx
q3S89aJsFtv1fKdrHamXqDYdDXQGtFtoSYbShLFDpGiuPmjHzfTEFvn/QrRWIdus
TxeX3xtGNyHEiu+pMgE1G293KXkoih7Ma32gCWHLeYBx4ugjBgmpSXl4/B/a8/TG
WdAmW67mu5GcCEfQTK8HeMXpghaMgIEhgYyzypzvxwwbF0fNjSTwlmhnweAhzKtM
9cFe9i/1eF3Hmtr/h6LWPAqEyKVKe511T/EQGuNY19aMMUUK5c0YUB7gG3yZiTgZ
K3rai2Q1aSMzI1GyBfN3TB+KNY+ZMhw7vlSLHVPDG9UhA48rDDsqMUJOHV/5j0NW
kYi8uzOJEEN+yR5z9zvgU4OjZHdRUldT6MNNKkje/SKk0GpQ2IziD5SpidaP2zWl
29d7/x6x/Azyl6I1R0v1Sm00rBUxnlF69b4J6F8sWEuUSuHle9hAFv+Hk0gnVJht
5lazkmsv9kqenVFdpL3xGa3F++wMVyNxMuQW9KGpu5HvfjUdOpQCM15hmu7ww7ps
AcueC8AgRIPuTH9sMycmP/RRc+dQtQVb2X+nm7DLpVABbLrS9di27v3rKfKSU4JA
nOqv8Kf+KftwXGrGgdFFP07gOqBHUco8tn2pznjF5lprDlt4hPwzPkZn+YC0J7bO
+wxTtvIoP1T7COQEccVADkRymYANqtFloThthypWrJWAmQ+VlOJmA1PrEak3U39t
WOfHSW700Mg54ADxquTwqiatt7hBGgqKtuaJNjXfMjL2LBdbquJeSnQSCHQEz8/3
AaUVwgUx90PAZ/sWC8Kd9hc/iwmwoc+8WoTejkwt8AeRe8c/Wzb1Z6sXzuuzcEdu
NUxT/pfPTLDpwiWBEIj+AOY92yNKyCxVLUrMoLq2vn7zbZdrujQV0sD1lqa5KbQO
wn8Nd7/vK4l6lu4IaCIQbuHSSqX9vMhx44YHOmbc5FgVQpC3HJ9rofrpbTfOuaWb
App6/4OqBPt89FamjkZxFA/0QqOAKogC5zZva5RrEDIbBIAO8c4U5r5asDawNYp0
5fiaFudZJABVuiBaLHKDLS48a6k47kodaAwyBX8IQsCaMl6DxOViSnRKc2N/4RXd
sTAjL5TJAgiiHUrqgzYzuvkMoLCn57y00sybS7rhMrxDTpzW/EIPp4Eq7MaNXacz
eXBHsWOMl2kver5H5xydsYouV8A0OeWPNHZZVKTdNqrSxEnbHrAtvAe0t03cRHmc
DzZuIkeJlFMwiRjqmZq/nPdSU3QpnJnB2ndH0BlRKZHBnf1VtTtR2no7T4QAzAAP
HQg5ylPWcnJcYkMOHhyLy0e9Sr2uXGKLUvC2GQJ3luQbAnSyO/PhZ7SyiN7mZvQO
+JfhRWsg2tCjgzPGDllPnowAFL8jpXCqciUnLJ1eSF75dhA/8Nae30wQ1RLW3AVe
1p3L7/T9Ie3ryXdmMYtKR1LIyqcCv0yy4lVt0o64WXfzCSiy2AG736FjXmYaJo/4
F2EghQksugCgttWhnDQekhDNHM3xmYiyyoPX5ZmgkOJ8Q84kLN6T9XmxTi/5i1sm
kg4SnsVnH/TAuwkFvkM86aQiR/yM8HtJ7IDjCak7GrRIpuk2nlZ4QqruoNK3jO7l
esRO/+88f8XyyP6SGFHw6ldyjUiH85LFpNgvMFAVMK637AYV449YoLgjzj4+Ybop
aKQGxonJgLIcK5pKG7Z8jai/gPAapQ46YiYk6twL60Qg4vjVAmleNV5y3JKu1wnN
XYtZRmD2IM0EIjSAQrC97WpnIDxOX/F70Rlf08kLtkfYzppXubfFmIfPxa8SiEbd
QU+u8Rm5NgLQ0cXy4gb/7KAd6tgQQzekV2KZioubF4ie/o41i2U4AldGp9t7CTQe
EBMxdpL98vcvR97qKoPGYlH2aiEPs2NFLKPnBwJB8yIkzPVkYIt2o0piJzbSW93l
UzU/kjgyh9pO9msoqSaiL4jm/c/OW/qsehh9htztaTYfJY/PEb7Xk4cv5L2Ih0OV
qurqjMhjKajhpi2jxHmo53GkULhIaO/vj3suwpDacZgWKv2ad8eLfbqsXjX5x8pp
+iP0Trm/n+CZeWOhB/tCWF9gBhakuBJqEYzQcWXVx3ch3IlLfypkYtvVWaBx8asA
aRVYuIEZ9tApKY6xQ8AaWRkp+pyNPjMthxeAGp1qwOM54BAAr88iPjaE6/uO//Qa
j/nbkTIId2HjkQt3ZOVKuT3DFjhrKEZLaGDFAeU4nmo/vBK/p13qQMEAqygESbzt
ZBD08ln0Azrk0eDoB+onIcXLIz+S6m6kpywIuK9V7eAbYeF7ql4v9sMpgaU+KyvG
sfiZ/l1eRG2ryLVNvolg28qk6J4ySY72PfdjTN9wsGoIdkTiZHBeni2er4RdZmqV
PabUrcbTYMsPTOsJUHGJ9DGBKAYpS41tNi3lxrCGS9K1s5L14Upx59TEH4rzcW6X
htYmbo14ViavQs7X5UBKd2A3dBv+jrxPrPSQpy1OTPwlpMB4EWl5FYKZLg80tIDK
Q31HGiIL0yvJtzq8FKAHfP/kpzBi6AGImusRsPlb8qfsPPEW3vxQKZKqdP6sonSG
MebFcmrwIjqKQgbyVHxLe2vo9A2b1xoorSFAFEi+xzLa/D99UfsSnHSRsSDuxz5E
oHn1MY63qzQ8eNCAPHD8+td6wfy3n7VEfZpOUIBlVhHd1OIT2qM3tBLp3FFXGDWn
iNql+JrxWZsWcCZqAxTBVkYICfETVvR4rIFNbTT5xEgt8bDAAVbGP9LrxCTnXHZQ
B5mC+SHcYBpXmn8GfOeX7pjb0sxSWFfftXFJrzlWeAVl4fWgxkcQPJf+I+8niS3V
DM6I0rqQPy2d1yJa58kmTfmSN7hT7yLwqWMULLDENDYbpo9B/+T78qEQQlIP7JxW
Zj5Fl601sbR/W1R1nmEj++GqaRKrhmyIXyogkNMpcSor0wlSQ5nKR9KabS2Z+Vh7
4ctyRp93be6sgIpp7CUE5Ojn+UdnttzZUsVICknqnsdMc7XsQXFECYOTDIqELXjw
QEjLHbRrcgmWNupSInFNvVCGNPmpFjVCmURzcUssFYJThttpar9pwz9qPrkacuW5
eZ36FqhVdaT0Tk/4LSPb+jntd51DmMq1QWVe08PCjwJexm4DTQjB8Pc/yPstk/oL
S057jI4E5IK1pLoi3+jKrw05AsioOQKm2HQXC+D2KS9ULz0ImQ2bxrP9VtDHqc3y
9C4Uu8vJwpfWMt+CXGMVh+TMytjF4qM3aLpi4gXNsp10731aIJTnAsMaZ1Z6h+PV
PYm3+KKbkkfIrCLqEHYrM9KWSLlwtsKvCPxgdZfrRhbMnTS5+Pr/yvRlni83O8z9
6n+71MWYPCbGS3uIOqt5GpXL0VQo+THoezB8xKYOppyAzryZkavN1hjXxxlP5yYL
cEDqD74LTMxYNcAVfNTPa4hx+JdWThU/P7BCTLPUqefEQyey/VYH75upj86IyIQA
Dt23fqZC/QTcocBM3GA/PoStK6DPevxIHgBhTdxvk6lRJ0Ynacz8KfSWP17gKAoE
7cLD3j9jfGBowIwOxcc9F3p1vP+yiizmznasqT+5BJYxvtucvfbDwhqAQXli3Izs
o7sNc0jIWdCyB1fW0WgeLPrL71h6l75Z1LEKKAHAp8jhX0zZ7zbn/a0Wwi+MZD+7
qev8Vsg+/uPA/P4fOS54IdPYsGYMpLzIwURxtfTUtxouyjKw/1l3Ccr9mnLxz7OV
7xLOHJ7rc0UFoK9GTQvJAkXNypMGAUoWxcXCUJyZp1rfgJIdwNJbLKH68LYhA/ds
OYVtj46klnYbXFvs4ld5Bsf3ZrcYb8yli4HE/u72bZSPtEdj5TMFWJP64KIrMw90
lDyCg6AwUBgEpzwD01lNlwlBN6xmveSXyYgv1/Q0tVJYTotPAW7IXo/tArz9THuR
mTfgRSb7JQGWgKMMSqc/W+HrbDsZvhJD0GfQM6iWDX18XIJZj2BQtNXuFLxa9yNg
U2pMwQqDiFa9v8GIfOkjhtt4XDs8yvIQWowhbD1d8fTTSsK90lvZzF/jMFGkGTOf
Kzql8CpUJU6ZbeY/Tu66UcL7w85zMwiS8DyZr3NVcT0TZSkoaJsvA+z5xhEytJmM
Pqda1ajbe5c0yv+M0U2vNNVOS/G7coX2GIccuI3W2+YgLg9lxEmRaUK/vJyax4jr
NpfDfTZhdYzpmsoECbcbhkAXCpuwqgM1u2SB8fIsyZZT47CsX31bXc7wHCOrLRNv
bFxohVeNtCBNEerDqaQl1rflyuFRBhkcRwcjOTNlWdGoyYX6OhV6ntXx4K2kg5uy
cKijQsrhhOPVV88L7E+SubBmEEVGNawpEJjfyNR7OULRcSaTzcBl7MkmThRDhaMX
2ZsexiBlRlPL49Qx9d8EKATaD7Ju8EwSi3OysCalUYSc4LZwxz4zugquSkd4Q52f
WeA18v9bbDA9nEnlxv64Xh0y1BjB9JQwLVTxjYgmSrM8eRAn6iuZ0Ni8ON6C2QOO
TGWMaKe0TcyZywa/nmpGMNi3K0cTKsuftw201Mehqfe53Cttu/O9pxxgcEIsI8YP
UNzix4h9OYsBKobxvPQt3oCEF9utWMWFMICOxSFbL5Mn+q8EPCnd5gFMrm04gekN
YN70PWBLYASqcgjp1lkFf5k7SaRvscW17quDGdsXkrV0FRpEidO1hKuoj5LYfFh7
Hei82Mivz29XJQe+c5HyL9uYMLV8QUJGdH1AXd+82KsW4OJazEHx/2Pc4aqXepaC
TVGwWWHrN0bD0RnR93hoob2tznJftYCeT0G4jTfcKdkf68dsivGkgFTyK2oOCj63
YU5qg6UP/L9DmKw13sqJnxqJ1pkhe3GBH2/84ijCaJ+Nvp0PpPj/wqiJ0NwBMHRv
+SvvD+3AAr7Di1rKv+Ab6cT4jgLGfNPLoIqx4Dr1VmR8cMb7TLpucek4kqKWl754
8S+ZpaDRHOqNJF5PtpoZq5JGEY1LT+79UTtPZrthBRrUYsmkgnnUwkpFDvwGI0EL
JPn/nI2fBUEZfV70JsYN0Vq1Qh+kwHfnAuNPogWo18N27c3YqLJelJ4/mQ3/0x/6
ZlcYZQAsJSPjouXBZdDjDeDa90y0PHcIY7+/4e/WAbmbR+JHA6XuJU6fT/eoLNCY
fUqKapxLrrBJj0K5SepeAEP82GqZ3+qNzi+5QrmMnTdVsSZDRYfgPeoADnHlmK2d
/NIQ3yyGew98ZChscZpt/Ui2EYTa8Uwfdoe9Xu1B3RlvMSCz/sWfIiTyg29R8xkH
PgobA9WqRHThjSJMR46Va+VXD+dPhLASDceVZkvxIE/KmdlrK3+VWjcDqn0dJ2/Z
Ps2c14Q9l+3Zed3FrzjvaxvW0pAOrLJXrugFcyo8h1Fn/TRpJpH5CTCxZ4E69lWW
LHG3wQ9il7XvGZvGQPYgmftkjFpo1DQ13yZpaWF+a5iEjsksuWRAdghEsfDXq56W
Nh92V+kSHQAeZ1pl5mnRJ6eSeZtLtehIUlxDPZQmBOrsvkEdZijdGzBw9G5Ons8+
YQBiyuhc4CKk/QThxFsN711ID6yQhYCC5CSj/S0XyB/Zg7jXg3OAKxr+6B9HwQR6
wgEjkrFD9YoCsivi/fKWWjmg+Vfl/t4jP14+hvDmywEIsKdHkciP2r5+sK6vosP9
LKkeOBb+j2TXr/h45kaRZYGM8MDPpdtDTVWwugjrgbPNJ4eU3t/3aeRvCLvRpiIa
TjDtLBM9Qy1AMvmERxYYGPe32XAF+NXyNV8XmJ25Wt7Xp1GOMpgt3e36TmPAIOT3
nZcUZRYNTnG6deUdIM9h9S1LEmMhE/vGrLCszxATgxay+QPc6ttEGhlNQcBuV0yl
DVVmw3dH7tzHVmN50iWa6O4uZByFs6cHk/S1S6OXTqYDwvc6RXZgg+m7n12vO4dF
JXV1q6vIj0FZS6r2+a2re0D9wPjzjT9DnwhEI1I8ClJqg6GemDakTubnDRGxo5Nm
/jJ6Xby+ykFhM62TxEum9kuBqvq9fIw34y+yt6XORpJIFt9ePiCDa95FN9DQW3MZ
sNDOPPdMWa97M08u0Cy+sxgXWcH4QmIDItDHChgX6vZB5KXuiH+PxWMacgg/q4wo
miMfpLeS3QRZtOWGOa/pffwC46EGlJO7u4Mzc4oiPV3CaaOROa55Ka/+svUGwoFe
Fz6tBNXhAryRKfcqU1PqT2LTV4g8Bnr/AeEMp9rhHR8f2/8l8Jw2bY3ihR++h/VI
WGqrJV3ZdHp4ChcUEuZ/JvvbVyG+xrOfomCtMEh4TrGElPSSuK+RLN07a9WD1U2o
JWUJrduhhOXRSPxCgB7Px/5R1xuvkszwo3TPLm+ji4szShogHCm8fjsyBmP2ViXy
riQUmOOeUEcqhXCJ64VZZTX6SKpKJ2nWJAZwjzbIg1sNey7XoFeRXltHRKt/P9Xw
hN4GbO0ZLP4h61eTy4I+zNlocz1nmDlWAsgYqg3tgJjLE28jWgMgoI2Tiq9/n4nR
nCYNmbyvJl7c9Xe1J8z7NqiazHwdiKYt3TiMiGc07GfHeRfXWin3ad95kkx9yvpz
2vvX5ICHLvRyxuUWErUvAVf4gc6wl/MQirV2/tgTpO4dKPb1I2FSxiHufPUIezCf
QGro13eM4Gys9NOzxqnqYeoqOsza/GmWuDRLOn80sTzHFVrjc23BUirg9taNvoKx
puB8AM0WDXKuEzBtIcCOqmuNui4u108FkbRkZjweeGVlem6fKg7Lhd7k78BXyNj8
Hok11MVb8G2+rqXQm3RWKDhRcU3v2mw02Z0ZGOM36OEmHJ48ghes0EoeQJ0QKz2p
a2mf7htdRQkkdO5Ap344aciv6CzSCDoztJanbSbD1hgsYQUTqducKfVAXgS65JFc
ny7TaznQRGSaDTwSMFMQKN3Zb7YlwOklI4/XCne+mIaRXgiloGMQKcllkUTqwrSl
zAA+oXPVtecR8pkjcKEWs40l1fkKPWPfwW38uDNH959CTKjf585RLk/KmHY8qlA0
+KAwcVErnIU91cw2EKQlbo3n4SGjp2FD2NiVIqR/0XyeDzV2TlKUsT8i/7sBhZrx
TcsD3xpKe6t4MZl1A/0cfrOv7rOWR1RUlFeV0njrpf13I+LizWlKBFzwcwgiybWC
c3zXqx/TZIubKmwEFr45W1dPTi2kesAYFcW2h/48sEDG3f98XbJ4iT06wJzZqqau
2QPGRaScbknmTrwL7Kh89iIdTHMOVjV9wMbio56BDRF4LOiQ133q58M1MW0AwyTe
8CgvYMu/AzWc3AysRrYNuQD9/QBYcb+IQSuVAvqw/ICywBMMFeo5UzoviDqomf96
YvqyuG8/1nGoOR8FSNoVtqxisoyScmKIlfQsm9m9eaf/0CIVJEYimW05mYwjfE07
EPsBZhWJ2vSce/Y0NFKzkCxcsB2T/TajlDwAGBF4soVwofa6vAbAN0oEQyi/ibO5
2UaukOjUmLvkBouDxjPJ7cJdcffXwjCsXwI1FbBs9cTb7zixIasMSCOsB4C5F/5S
MojotSulzPMH/rbvt5CEpWE4GZuTpyUrRDi/R7wlhnXdycig/SfFe9LfuY7JJCfi
9MCXScHLVhWMArQNCXXEznpnLlb92RM5Y8X1Sd8KjjM6Mgt9q8Tco9zeiTYpwjDy
hpJmsodjiyNS7j4caodseEzIfIdbMlXdMT1Ynl3QO5scP2AiAe8/pcjcX92KNI60
VdY34qTDj8dx1jC7RGtOwaPAtUfTYYX1cTFN+CO70wqizjLkGEIdpr4+qwHsXp5K
q1EHS0ufvZVSeu5JLkSNu8Nbgc113fktsCNUO1h+DC+CvKwH94W2okkEMuULKeKX
MDJLptr0VgoITTqKsE/YYyFo30Ee5eAqH/OhaSuBLYzllyXmiQUl44gXYQbzKLxf
zYjUvdQnJbIB7NELayw83XGgn2zQD6fca3gyzNAAY8hbpRXS+bwlJ3O0uNyq/BP1
XJSByAwt7LNTn3gaNm3t3pdWQBL/TpMhvSFszjKoFE0rQsx/NfWvhnFmacBwkWci
TPf2LBhkVc2DBdYHnKwW45aLgLitBWKHvQy4NYlL9tjl3Mqzy8g4wrln+oN4f74V
oYyvxmp4BkFXyngXReDDKbSDjecmD0nNsaVqeRFqxH4xcgiP6uWd/bsk7TyODKbx
64G+H6hznIcTe+IVlz+xdxPoHNKw/3G9sjII+ZZYCFJfcOHudBrbv4XrlKVvkyq7
xgvB8eGznX8+LBq3P2Osuiso6OWhK5p4zIJzrsVDbYCmnyLejwi9xGXMRuq+cP/j
Mwi/wNeQB6wahQOrZLqYNdjHOFgXgg0Sn8M19AhW7g8vqHXGr0/3y0c27zbTtQ3O
24A7/fKVqQyFIxM9HowQ1+6fNN4HkagkBfh6DUSx9n8BN+RFdrgPNcwrYkP22kbb
0O4K/EiiWDChlSFlqYNfRORk27ysFhWeLp5FOOGm0OdDtVEv0/PaxaTELVFOzIfJ
vuzpZ/7Scr7q4gJCGOj4vGaL4SDK+osn0ymr4FIsTQFUfTDA8DqpD6URdCw25hi9
IdjRhwtMgBU88I6QBSMjLwSCy8oMgjf19IC16qF84xzmVEBt85t0l+SBmrRdnRSj
gXJLGX1mznc634003j8bp2UBAhz6I5U1l4zgkXoD6qE5+eHzq2X5gZZ+dJ8gR95A
gJ3+cZ5a0ZKVhbwfFJ7MXC+q/dkVZHj041mK5y1e+Se9Xzt7BDVmbSD9INGMhI/S
fsey3tltCMOZ94HoYt8iupNDqRv4iDF2Xwkry2BBe3xHWWZ188X3RAND6eoNGkBx
lohTHI6E/IKddQ1DarbM/aRS8rzNBVyc/L2gx8T8QU8Uwzy773OeTdDyhDEzaCcb
QKJ2F4RJBUli/rx8RU/Yfdy1yFu+qy2B8Jq90mLFMJ/Gubt5wyg2acC+v737wCfJ
WrqDyOdovO1HNZ6ZmigoMx0NAuSPxLvrHwiUeW8H7MbUJ6i023GJyxr9pT+jTNlV
ZPGDItazbmpkMaYFny1V6y29QB4Xe30NR8/+yqViunXrzE5Qy2XXvCKqsWV6Yh8Q
AKyj5Ca0a0IK66WuUGWTZujYL6SRR82NuptAyENk0uL/Q76ZsdO7VDT24Dmza3lr
mpZfd8wYZFQv3RUldAGPiaNdfa2dZHvFEcaHamhAke/rQV+E6D/ebGlPU0nhbaIu
gjbUWA47oV3l8Un0NfC+KR6Y/B4GfcvdbEsIn1YFML5qNTmVThvsYkQVBQF8DXj/
ER8EFQc1HlpaNLxvSnsLR0Fjk4d5eWxRF8osZ/O7Wi53nUQhAM7CQFA5sz8fQixm
d19f5sgxZCE/1gJ9bUM+SXSFhNUSgVSFdPYjoGDAK/iS3T22ppwNd8KfhhVwu2F3
SG7VKzIdFl6d4x7pMy7GsG2qhRUd6FC8Bu8LYNFUHbrqDUrk8WddJ9bKVZWfP46j
0KS8lfe/coYGqAC9h9FslLISF5z2SFvjB1Jhj9g2NFGWBz4AJff8U9LkJI5z+XWZ
w192K2rJJAPuKtVfkK4Ecsj7Y7IPT/A96Rt24T4r0iMsF+KLpU2/4HJH9H2GoOTc
B+GJUR1mAv/zV8FcZCo0kTMVQQdTB6WGsHEX9q/LbCgu8vfyxAB6xdnbLW6jwC8O
GUjW+a51OFVrnjTysLmyiLk64w2DGSWdUoXOKorwHZ8GgElSRsyn8I98qv7LU6tL
QKYZOv+72jiTvmpIGQ5ZG/ZsRsVfCjNVVR+8G5Y6tBYK1QiWgAdugqNou5OmXaJa
jDne6cmD/oaoq8q6Ji/ItNURWVDasXz0v2Br/0a26LEdJjrKqD1eXAQ3B1MZa/vg
C5mDHkklODsXuBlSXrSEzQ7+oV0ehXlCTw4zmSK3EBlcHxDwcCorkeeacvlPXp3d
3Vhtx6EACbuuWBl/e2llg/DfnYoqVF0UcRq6C95xqkQeXeS1Ld84RtpAsJ9Uxsyp
MBzAZPOXbAiGbJkYGyplysbJTBAXysdoLnNI0bbyg0IXn0pfvOyDP01Yjv7jKLfJ
H3geYoatH0TSrZfdOZCZRe+X9HVRH5dEKAA9+72jiMDzLaN4LyA9A8jSVA7+g96Z
BFgjaXQ50z5RWeFn8duB0WTZIP3XYSxubUPx+CkU6Vob621SWauqjDwmhskxEfv6
7xyZ4YrJYNYr0QbRm6+SgVzOT6+0s0PDkHs9pGpiySuaBCFEuoD1smIDGKpVdOV3
mOV2y5SvxbuhUFoZ/fMmCfizmV2YVb4tKNmxKqRfrqh3LLgkf4GhnyrN8EnaZN3p
U87eAsr8NXc1CU/CNEBxbXRxwtFv6p4jnIZN62IeafNNwPl64xQH/UgRCqLwRXS9
fNMZ8/lpq7rXP8hEOvbu7PEuDGCwDlmVORrgRcD1z6V6fEnohrUx/vPxHfDq4IJf
lF5/m/1WaZ0ya5lTeRiHh0k5CpFTZWCI58xK8CYFbN0B1cPF/8LkuNCXJHgaTA6q
bRgejeXZLGPNftt+ae5z+WK6fSVlFwL4znT3HbxWQL9GjfKnwq1RHVh7ykr3XNVw
x5K3MW6wx97RJ6HDdPY6HYv7Q/WGp/QPDjuPnpS33JxVvnqwR21HlTEJBOu2sPGZ
bA8cgEWqEBOqy83MO/ts8EHKjd0zcrNe4BpPz96Osim1Q75Tz2y0Wtk2v/27YpJe
900THpOnK4G9z32yH3AAf7tnSxoGZO7CGjTTrudSoCdto6uILhFF8D+EJcTBOUdE
baHTwawNAKW621YkXGMgaI3pIXhEPg4Ed1ABi3bGcaQjvz+LaoVJrpB/d9K1l0TR
ecluia89hIE1uDMGcsQpffGJhjw8rcfOaW5GsOOco/GpxUpMLWVJ0kgF3S8+wg+A
6b1Dr9MMzbN9Zc5kQv4VvhmZPflR9ciz4mOP3qXOBU0yUvf+iWTK9aYde6qFYUSu
z6MI38XVL7zExcTkx0sJLpxA1iiOzuFyPWA2LUw56uGXG6GofTdi1vNRKGCWvd8U
nIL9565gmX8Ptdl23uGSFeFZCjCPop1d+0MRkc0EoPoDqTK0yV2Pnjk1WjTuX63P
mR2PGBIk066f93GWIRNCSva8OsxRAUaOp8liIiee3q035VMEzLP6iVh5C++FzceH
Pxaq2U/cgnBZQwTd75erPnQraRBclzg3DZZRKQ5JnrU80gpucGVAl/J5uNfHOr2k
UmTD9HcSgk2EpXL6l4WcqYXIt0QnKFflMd1MzdoQKQExYIX3yFGPH5WZx33XLwNk
fo6FIHMR8q5xCdLl6pu8wjYb44c1yYIF6RVc19n4mzjh4lLZz/1DjwyguQOsiQ/a
jyJ5FFusGIU0LNyuVV3C+aaL39maFpix8+JxuGHGKMCEW0cSBJD8j6GfGVjydlRb
qu8QRlxdywxLpNetK4RfJbXESr8SO/uSuJaJine93gi8ksIRkBBJ2/N3U9PT5YLA
AL91vwlPY8i3UGM2GHJ5HgCPCCupMY0kXOrx52YvWzF7KdGpY3WQ4dloc4sCxPMO
w/pUBmvOsiXn03bs/q28a120NOhAwBTcIlZB7TCJcOGwyl5v3rFvn6GO/p6u7Uiv
ErHQH0OuYVrD/OZAGnernGr86nlnpzUteP3HLy3gLQBT6IS98phh6q2VZ+FTZpj8
gkssMx8305+6AY2/28qDN6ZFx2ik8q5jcHRba+G7d31TZTEYG6YuhhWeIwWHveZw
cr+KTYUAcCtozx/N0IMb4LB5KccNKGtaZMeryulBI+RL8YBfrg/wFMqlN5X+BR+H
AI6SWWXm6GHxNCrLu8DN1PrKkzrr7vuguFKjwtmLaNqvSouTw0eXBCJ1Lzeu/2ex
m75RoqAtxsu3QBOFRi7hXQMbSxzOWiv4sxzqHUGuNHFv+ImYrE5fARq20M69/lrU
oWblVHJJlJVa8b4WI8S9N0yQzRAO/tFmGmyemSxjGTI3VVt7pmZCCR4LmujSqSlY
ubNbkCePMpA4afF7SdNCkl/mpz/B9Na/7oxa+BUMaPb9tb9ty6uUj3pUh0SQfcLW
WNJycESZqNXp5Hu24bQa3IsI+txdZORpBzSb/PcGgfWmOqF4E7ZNS/FHKIqYG7Zr
fHmMiby/bc/m/oAm9oG8jCTydh8f1Zc8bFqtvUQWh5W0Zttz4vXZySFYWneSk0wi
2xuqIfv9Ijv/8AqiEEe3l8t08epUy1LeUKY9a9Y+cHGrqSXw/sCae66ly8n6QvDb
sgrfsYsViUpDbXvx9b9w0VYRqCKpOP2pJ6/8vSX6msI6Xa2IwncpnRV2IfwT05tH
YHLZiCPFseGaNXnDGruO7wrXSdj6LKZMILGvMZq9XnQUt0jLVbyQwQKH0QuVfAVo
GHIJkj6vOQpfMcZJSiKK3TmWwwG3Y6ZUddvcmDxB/BWlyq5nemjNIZ1F2smB/1Ii
b4zFbQz3TouHeqWDmEKtYHhEE1wbkJ+TUJCSkVBTGIV2wR13r9fGSc9TkDaqND3p
RN3QKq6PRRLjEVcBhZ2eOxVG8SY7w9nlMxc3ZjWcl/hf5IEaLAAiCf115/fcbQrL
UP8Ru+DF5nWcCszz8utlg546VBtzT7HIUe8fA85b8yLOgYr7ezy1MS/BVqQ2treH
XMM5OSZjjc18Ahqak1LnL97eY5zPGCyyP5wmRyrUOsu8a8EmECwjf5vNzJQWnN0R
G+2nieaY4xHRwPs2+1To4Y62J4/Jdz57eCTxLqghaNskfEVjk1ZlpXfLy6Le0V5q
zwX10PiADwA0q6KH0z7sO8ueosiqmcTzjEL4HmId1os9G8JtFmeCs12S1Qbj32aK
1d7nnvstz1aTlB1kXKusNOzFDKecvrGDsDHT0K8yRV0GUVsxvXbDczVy7TwJQXwQ
3TygUaoGTz9stSt0ql+T7nbXUldvQzp28BRr9CD7WOhjA2HLGvYDaxLFNHnXMoD0
LVq7F7GrFnN2bynx1ss+lusN8B0Pcg4D4+kVOQHOxALQdCIxkfpqMXJbhZlhdxMj
5FL1KL/GQ8sCwwzk89SoeR89LpnsNE18U93QZK/O6p1rsSWJwC1TuwjuWM5J8TSD
DIsihPFeUQVYg9TRX6tRAWkC/IR6093Tcq2IN+Er6y4OFagt+zqG96//ZnZxvAs0
ku53hUs95nlNeEaUWbfCH9GsIJgU0OwFdtNXKaWDtOQY0b/rBWNOQP/PJx4oNyOa
qmYa1m6EcvyR+CeE6H2u8aYWEVBscmqCdzkYK+skeGXxEYYwfgwEVJEEhLK8V1A9
Xwtd/cqmlsNaKATCArk6319mZSNP9KuQ1QADJGBeFhDWPY+c4Z5gAMM25ga/RXUT
GiSjC2zHrHFtKnHzRNtMC5Ruhm/oXtAgLfQp6SopgbUHPi2RqF/YtSujrTMaMoUF
pFuyVJ7+zIJaFPR65uDr5NJK7gLJCEkJk1AEvXEXIZu/iw31DqeCNdxXX2tBwvDc
M1wePui91v/noCTkQAcD3hq4zuoZMhvHv3c6dIKfOKu3xGzn3fusUr7wJ99NFvi5
gSYHL+qFQ+1Nk3Ueo+eBb2pYjkpx3ggt39otOHMfdgNwPK+OyUH4ugTJg0JKsOWM
jGKZRhvh7uUnjNoWf6BoD5YkeYOBATlIewE2X2cUCEP0FH5cTzZkN58jglHR9Yip
qdMGx5zoRiIJ8qJP1T9FQ6527TnIvrMZQqKTdAlkKGDnpXz1kJXEiC2qG9DnqfZx
cVDDfAeaAi2k4y+FZmx6m3FjyGYlqjNP0kFpsBhzfT0g8latVwVjAk1gTB2A9Lhm
c4geJkldB8H1a6wOy/7wqs5yP2ZRyYksAHDLyiWwjE2ChmaNw+WQABGBxr8iVDGp
UAfKT1DxM/Fx0AonrXKyRe3NHFo/w59/QU/e8fwP2/XQhq4qoGgdHu/XOnmvtEWb
qUnPfg0h9nKrkT2pWHbbzY8TTW14HqtlbpOniJdsK8eW/p7itB5Y4LN8d2vaYprS
jk2aA2hru7ww6mVnTW4CDQ3FAP38b+1uXDhDWb5rc/UDIIfO6swdGp6g5OSXya/9
L+T+AsyjdgCNMX7eeBvpL7YampFv4zVy/ub3u7x0Syeu0uqfSLhxvFpNG2oaY2/e
+1lRiQccaVQgtlHL3Nmw6kjpapVuj73KITXWeZF0BO01kEBf+39vG50KVWLlWPM0
2dyMyOwaDTeHlCGotLaSXa//otZMk+DEYfZ4FLafPgrLDWdtODYfToZ7l+2d0y3J
XQcG2lxFsxy2uG33NoUaud8ezs2nAOgv6Jw2pf06WdgPSKnkl1te0NvufTmz7zCI
amfNFDu3xPeSgdGm//s6ssfbnftj1yHi+OcuIBx522CKSwkvisvkHi50INrclmTG
Ro9FUPdpiN9iPA+mPsmyxJAxoI2hYCi8oM1DSVLCQ3yc3v37Ww35QUVC/MXATvlc
gGgV00ThHMAaeXWLJ9NRwp376JJLYvNgaGmrbUWtZ8fxQc/l1Ekp45DNqzdvVTni
s8U9rnnOhlqEkRjEy6VoHHzfCMNa8QXwwAazAurBJJmAzH69OcxIc7FERyIZh3ar
GTSq7JsVDCboWYE6HVLxqjf3h2L2dSF7QAYVn0a/w35gLlhJwOXxmOu5SRjSlgSF
OufZwYyXUdLhoDOjXJG9JUEVSjr0e6sQ2mb7RdBX4JRDy6EdVMKelRj4wI1TUQ54
z50Cj7VSD4alApEMcRH7B1vJBf36fFrTD8U7LOCXKcX9eSMRBH9W7JPTdZruMIdI
P8g+BJsP4E5mzu6/pAQwR54Lk+wQEOUDCUzE29j9B1V2wb5+Qn0pju5usHXoJJQT
TX+NY13Vn3hiEGy9Uoy2/Heb0Z+0d5lPL0mm+P1mscOUE5nOnmRRc6VxWQvTkc2H
3Oktqmj1lmK/U97Dp7XaAFnjP/7kEUukP0zDcjbKqdwTF/BRUX4NVBDr+im9UB/s
IBjWdEtxyJhW5HoMutka1ULxvfFQBwJbuc56Oi8zfnQpHHreN2nDl4FVv4oe8gyD
y5NaSjlQbs4dh1nfeJ8iFDUFICJf8xp35HtR/3hJcIkW/9r20syhhbqAccad4A9/
NE+bHfumBNBMKqYjHuJnE1N+Oz0rEciPEipCp13YtoHgY0GzPOaNUmkwzUTWVk5a
XFn7SuxOhXgoqbNUwqX5ql4EtIHEKKwvVjluB871oHleFh5dWI119d89h7XLkKOl
zdAyDJFT42wUcFtkPzwA6cQeNpB1My8gZM9gGDOTbyG5lgCiR8HCcmJiM52+HMfi
76QeDFTb9T+AvWydye7C1oFg29j6MQSAllxOgv1NF6n1aYnifq2wwvM+Yko6SDxb
dmGTO/B4gUycDI4g04Ck8wQb4x9dkLhqX6j9UBuIlQfppZAt5IXR7FI7aR3dbKWi
8pFD8I/PN379sy9PK3m0JDImBJOt71OrnIl5wu5NPribvDzNTgg3dG+dkd91/AF2
SxgDbHKWcJfeaVD3WwoZUHl+Ams+OippWjVhWcyRaKeSCJgRMbzqw3XevJZcO7hU
B41F4ls2sEyRWeOnEowmVDmyOKUFAv8dIklod7BaFNU/ptf+5JE+22q8jrruIj6h
S29mAhsfryV3rxH3gUqaW2nKMzrkqKCOcHsRLQbyx1mcLoC4JlanjdRufyCh27k2
Kk+eDDnn7962XheXXN9axADQMYMXrvUtlcRitVZ/JnzPxvIIL9f5Gk6Z7Dy/25xn
yEwn44wJjsi/LQLnyh0vRIJMRiwL+kNfyFkccFkmEZ3TGxSUlEFfESDlwZrbKR2Z
Wqypfw+bVAfd/18NrafQQaVcrYdCAQbnbMBI3yFx4g07+PoaWsJidrj55x4B+57L
yozVmb8R45MoRU0yp8WPfC36nCkNQK3sqymOdmoKRVFjqR0C/H//+n27yjFWP/JK
MuFs8XvcetPT47NeANMtLaCjV6m6K2IWD4ga/6fDDRP8FzF4UJ0YoMu9gkc9Nwk5
YO6ep1t3x4AnrXv4IiBlUPvgfNLpV2PWhfjwry/6khU5huEeEWqbOKTbEfj+TY4P
XwVGcN2Od1H6mYXAq1xWWc3l/UtHTTItRGWCjSFn7rC0UpkXZrnjg9yOLBgNuPb1
zgqy1n2E+uSDYxgOOQN9d9SBLCTGMM0lR8StqhJs0kLqGLyK8GBXq0i6legsF2AW
6kBUfvlAS0AgwH3HiGE+QRvsTqzmcOJevQpIF5WkRdegtDiLQgixB0Df2+BjqKrQ
zbbZ9OcWAYPaPYuk1fVp0bA/kACaoQMBWii6+YvLxWe6x4Plk2ug4VR0XDLvr+zJ
ETG+n3VCe7FdZSPL5hMHRiblxOWRNV66QHdqexomdK5BR2k9oA9SKRvFfZyna4os
i07VXxgPPEs8aXT8PFYPPqeU4GC2IJcQrS5byQMYhWtSiFkbODMYYxF9VTNBwiuf
KhZCc/czsBAWIcLxtdBtXTeb7xYLp/6MGJJQIJZdxn0VchhS0yAdgLbnHTAhPJzI
fgBiRtjRCB6BtkceBzXP9bJ6hiJ1INgf7N2JR3ikdLJ6BjICXYLpFSkbq6I3PHB3
X2TKg2wClK+3OiXJz/tqSbCCgPbvwAPJQZjrzOGjPqvrNParcpq2QgSSxfEU2fln
9c/kdTHFjSTFAyPBOYBJySrCElQjxDCc6EN9k6XHYVW5cKZcHogLCmki7qjN15UB
KDyB9JKQoCLeIZeaePQSDnOhwt74gFn5nGXoSS0xS2xbIp5oDHEReQz2zJ/wgIGX
2JKFIKCMigv0aNaT8aUhuoywnrBJb3IB4A3J1dtT01hVPqEt1Ud6W9RpJsOhfZum
/IY5fAallMWlMvA0j/Jo4CKpf8PsKUv4h1+/viEI0WguieGomLlmYap+AiS7i791
/CYRsRjEes/WODNkyU3di5HuF+Xn7RLGx3VL73zz7NIyWnAFcxWKz8a6LtvjFoQD
WirHLJ/cNQr/wlmW21yViCi4dUVdIQHOFzvZEwBItWipk5tzm7yehWVdXs5Cc2Gw
DFw22Fn6noSXUpv5OP/OrovQOxMpGgdPwxzoC05Y/RzHDpVglNII5cdZKST0EiKd
N9Bqy0T7ZP1HZs7USU2Bc8lY90mtNnFGqKPALWPRLYeX+lPJKnJaYrcgia1dNQN4
9q/ldlgNuaI947GjSe195hf6j81qVZfEl2enm1A6+OrbvywgM9ECnCrAf0GQnH10
1CfZ+nawpOaeAYUU/ienpt0joe2Cu1jwe459JCThpLvzM11gITlh+/3nvIWU3XJt
jmdJozVx5ckHEAhp07lJyX6NH7ViIHDgVU9E3n3Oy4Hc4V2zqFodqUHMLA8TxVVQ
BR4omKZkkNmKUQsIjNE/FHNIfHMPBVAsuLKTGkvuemx2xOfiXpWEAYw+WVYZQCCV
D4Tvu9aO20X41cbhMbLvtq5p5WI15ridg2TG2GS5WLZ15Psm1tFApvflZD5ppirI
1xiHwnw7G2W+VAJeLiU3fvvSyvBPIEysss1LuXRPbgbYTaRKnxwLw42WkCBegaG7
dr8FyDNSKwvlQYd9tHvudiVuhRJelRaQvfI+NZRHfVlHNpwc/0hNG3JZxYxPHpfR
jztFVMcRhA0bhKSp7YduDVqtrh2DaHJ/HNnkbyaf6pAMOeIIJObWN4MT4bi6ncHK
ctFogSXuscnEkORukcg8XUEEGUIYYb30ZnTJR4GYcdIVuLqoXskr0AnqCis1YtDW
6DtHyJehraGSXm1RqlKiRmWmSevQ4Nuo7b8xxDeS/Xzl23HPCqOCg14EWOwSNigG
UhIJg29sSOXoqgBJiVWyG1YhatYh5sagXvbki+7tX++eJuaMODwI1GwEXbF4Vn6s
og3lKzpU1un2Wx0Aa6jSOEQTbx1VjudcLtGgSasH7imVtC1Dy+6HVS1gpviZunGd
SlGbWQzgOtdEW9SNLZuzlXk4/W21gcbfquBfxl/95XwdzXouxkA3yetCjpVD+J1K
sjuokTzKcjzOPZVh084O/W03+lfWt22/FY6n3sWX0e1NxozQa0zzC/DX2jSI5S91
gW8u3VY+VgHOtcsqzV1xvDJytlz4z6jZ6iPfhNM4MvpoADInraJZxxc7mqiyi1iu
tCA9EtJRPpeLg1NYOt6+vbBdzthxLyEzwTgJniqQh+wo0TYxfNqAnhyWMRXJoip9
ca1uHfwp/s7lB+QrD4x9e3H5etGnw35222b+OzNTFWmzeTDATM3GFFSWvMl3JlpS
61+VM2WwtLI5CBRsKhaKafoMZPImbqe8w3onjeyCGcldY37D5es0xqm6TPtWw6be
JMqtEk+EW7DVNgdxQUPahOIBwv0f6VD1TlTXiJB9y8Zcn2Ac5xDNgVYLTugWRCBm
HzUHNTJt9t/IVk3/kRiW9BqtdFdaK18kclK7I4Q576kOYrVWXHa+v8gp3HwYjEKV
G0xJ3byJecgluN2h/du8faZtO7whd58fMhLvEpHjXviDcscmzwXeEvZGkSOq9kSL
9IP3Olj1F14NxeXP78CtPls3oQ3YEKBS0QiA40wIdHgJCFTMAz/Gh8iARdN9KKvS
5C0Y52HdDCUXlbqWtiB6OLkCM2035kgTL4kTNKXmt+vzismgK5+otwrIaRyW6huS
eahFKvx34SwrwHvUe79pmoNtK+GJKCoS2SYBvPfrOv3V60jozIGWyvd3dPDCSzfL
2NRiTEC5Z4mB5ph6eP2dO9XKdLXqVm5cFhELopL0s2NQp42R3iUsB3jknsRx9lAt
K+IjmWwXIDx52dqC2lXC2IISEyhVhdyOHHyt2/49Ppupe4UtJeLcPHYBPj2gxsu1
uPS9tRnKpFuuaibnc7o5Gcs9ifZjYHvaGpAY9HZ8nt/YJWMMZ+uT1T7IudaAOivu
ZR9A7esbL+nWJCaMrT0PVoqpyXRH0hMPz0usY0GbOKRKV+W0hMXzBDLrCfSlO9OZ
QH4INXRc4KpNqAlbhx2DJG0YeszrJXnXxZhOecQoKqe83VhJxB7YPN1rRVczP8oq
kX2lO02Qeh75PLD2UYPlXwkEE4cfJ4WiQSuyygpbUo2QGwBMhhi9k9PPvyb4Mdzd
RXLkoj/SMrpuMfCRBu+ks/ylKUMunx4qkfhL+6PYmiyKIIMoNGuWnG3IQs/mDxNF
C3zlSH+nwEiayIL+8qKPapkizwKR1S+n33V7OgtqzMpocSUmKVBeXmrZ+QsynSfg
OwZQRiu/YiF/lcqUropvRoE996fEIwhxxLYXonqq0Sv1Uqmy9heCHvSTBYQdfQ1y
+01MZlUspRxYnGBfsbNPHvRHiUP9Oa/cDe/X3W/FuXB6b8HYZU/bkduyjswjLuLa
P2osOabTnFkEONpxqsm+iH2mkOBO9rkpnm3M+eDzGKwEuIOTtDO9nu8bcO8g/8x3
8zr2dpJ7zrQpGXjM7At4FWUsc5LFgz3Q5zt4E4av4TgzHoxEXgslKKKXQ8huHzG5
br8KHjk7i7qV3pFecCbExziAYRK9Q49KfhLOr6vEsviYLIccrMTT42HEaOD/S7R8
k7ya+3jwNupOaDFYoTmAS9Kik2VpP34nnQBGUptjgtR2Zo86chjaazbbLfgJRXJ5
5qwOKsMZRhKMFToHotGR+a7iKYugm6uiDh5FNPCE6Rf9kuRSsU9B/ObEXFkftX3Q
5GjCsQpGXauEDP9Fprk6Mc8qdUeTOTPiPLTwP+VcVZWcQw9etIQmBIOh660LN0hG
Nh1Y6aaD/4NXrXzsUN7fKisv8LSr2xsDKJIruZNYVyFnU32vLEBwtN3MBmQj8dkQ
dokhMsd7gT+OH28VIcV9rLisg8mUz/2LDynguAS7Z/mPJlCUNDzXBoRXQL34Hcpu
3K9yXiSwaqA89vLtefkpOEM8nQEWnvgecbVvDBRw+bARQ1JzZrWK6nPI4ibuV7Rg
3NsZqVBSwr5/QgQ7tyPEtIkanspqtXW7Nc6aEFRWVJHIMiuVlNeaB2gpw4DXsdUR
QF6LSl56CLEZ3hWXEPGSVK8gs7CP8T9vuMQQBwrRNrHylq9QqhukZcK0uxME/B7Q
9/qmzno/gWphKUk4XIfiwhYJyT4092DIkpILiyNxdMh7QAznbiDPsGNElUZDBSGc
G9EGirxPBjMorNpSAtDMxfH1swNFwud9otJa1sdDO9mNLi4rLDrpxo6BKB5ILgMI
0Gi8COdqFbIqfqWUs5N2Fe+bSfLc9SzSLSwPxvWwDfjRz50FEvCEIMDV/hN+azD4
9YU3A99UZvwoDuZow8G1pzDpwgSMzvQzxXFHVxnBKCa2wHQchbpXOBsMQJA7NQ60
f8Ne3c1IIgxFNAQerCaNXdsRmsl3v6c/8HlTg6yG8XB87UJ0c22eoi0lEczcyLNF
QzW/6BGPnch+Uk5hreiE6W1YA5LNg0KnpetGcvBFutn5544SuHYiJycZn0PByQlv
a5vcWuJxjlQSfx3WZ4pVVVXoXfvoWPMR/+yOrAV3Ee87Ft/gk5yHc7498FRuiw+9
oONfiIFZpYPzTYs+i8G1YvBfDorWAXKbyTFXbArap8ekN4T36oQ6x8vvtfzVlNgQ
V1/YIAzfJdxsqUqTaHElq8dwDy6ymxUVH5tvNyvHthAWZE48jH82NVisl2pWQy4A
dB4t+5kVvaTY3dUAwNXAGZ4mJyOzL6xtFUhqimG0Xs9bx4b6y016TGUsddfEs8IA
1EdTMjEAOhnevHygRer0UoM0Rpxa+rPLO+mjY0F1q8ZlSoZgfuIfg+Hj5gH92hmE
/a9j0Us+bZjySBYF1UOwTSPtg9i+2AM7jqBvL9oyLrWZfQz3PwvUq8Ha6PN+l1uq
zPIXU7tmStTAjM7vurD4TLgN5EHwZmNZYwkqaGundttAYsvjgMALtRp1QwMKhE+K
8e43+UsXQmk5PRb1+LK1TI5mLSrZApqejyfsNZ4fgmHxetDswS7WfywoNR95xTL6
FpqN6dGyZPQSumuyvtHCzvvjnQSsy8MyvJfb0ph/cS4sIx8hrRv0NFU2/f3A0t3A
Y+Puywbcra4+GCbbqw0UUD1g+APPhL5Hn6jUKzJUMukhSZY5fZdk1+M8iZD9Y2s+
kEkcn68fxAV9590DoyFVxfPjV5nbC8Wzt1nyLlPkeZO98EUlmpj21/owI4xJtsL9
dPz6C+vjsxOp40d0LoB4FbdPY8qHWd4x9034DAFfbIGCzsWcxeNgsxwWifvF2aIe
jieGHW7F6iPobHJZEgsoeMgUsvoghybJ7jPyQ26mvTL88SUuCtQyojBODthSjpo0
YVVsuUmBfoLWsdAKtBONmN/GeoO6KZDminIql0lhSHOXcL6Fh/Slr16HXnb9uNz4
Ze8TKnoWbtGrL1OH5LI2dfYeT/vbUjR0uHBxNwg4wVZjYEclrC7dISJ3+WwR8v8l
Vv42XhEm9GLcciWSJlLxOFwrvFMWBzYl1qgZ2TgkQdiaRkl5b+FZDnlvm5jLw3TO
TqEsC+6J+8WYi5Y4LY0po7bjYxMSq+e/HZw6bvTYWCDykGD8iE66FIRlDfD1HqM5
nm+hjB/UC1CBFiXueT7Bsx4u8UvpLgTC1hBOnHJbapGgECuIO05wDvUt+DVSVuM5
TOzR2off/kVZwzWOl3UVPlJ4eQj25NeccmLcTePuwe0buD/0he8VgjMQF49acp/A
gecCr9C4R1wXard1blTbG4TyhW1yDCP/JamGRRW5UeoLyh4KUXKj5xMvGYJXN3Ie
01zsapaijSOECTEdkN+7+BHEux7lCZLtizs91DbBCU+WObxOOuFEYw85x2mL7IEo
s/ontEuwdMu/MWRB4POndsyn957FH9K5OzPjKMw6IuhiWzswPT6moo+vXWUsAvVx
p4zJJUBf4o3GWMXQfgLQe0WY+ZkA0vwWYTjIjWQOnQnky0b5YIB1IoYrn/5Ok7mr
yo0u/gpoU4OhyZUGI47IseY7v36n4esyQuyJ72Y1CpVz00nWoZ8L8xZ6po+Qzk4G
OHa9930LRvT+PoyiCAhwKxX8eF5joj6hu4OzJlu5TmEwItqaPB6W06JQOHHIRAy3
RlvOKVI4gpOUudv6HF42GbANOwIYvFKpSZvEtTeBm+nCZS+p+nde/mOyIuudPQYj
/Cp4oDFf6qwXDaE5ts0s+aTVxJ0gtJSw0myg+ECnhvwHroIs8zz7fa5TLEYgEPLA
DwrFHycFwh1A1rjYMbWbEwO+zRzjfZNIZAvpSyR/8IvRooBWE4y9yGyqPYVZki7S
/Fq75EbDbl8ozl/+kJNMSBz8b+XidF4ZLb2ZYhIu+tsjdI+gBzMPEydA0MLElGWF
mkYQYrlVZikkVfQoBG/eZYdrmmCCAsLDfVZaSWMvx5f0wxYV7yb+JkbI2wl50tQP
n/3ev6+ArO7vTqQTvW/rdfrnCS+LHGV1FLE3vOEh2K4cA5FImmsA7kVf+Lz9MgP2
dUNvY14Pd/OC30liuJa6QwkAjL6R353JPQ3GePR1NOcSDFYrRWckvKyoYC6spRji
EOEq+BzR/b7t6JxcTuYa0vyLw9yTCLXPBwU7bcCW2EkFIv3D3Jy3zBmb9aObWg69
Pr1BFWeemig7klhOTLURuyPkAZX39qEURq8icMPQUNDOfW+Ya/HL80vuBDUgpb/p
b5QGxW3TJdIw2Z3f8hbHK0A1sNN0BtrYHO62jCSf2r8mLgzrIsvHMeYoYptTk4Z5
vLYxlWif/TfxEHahtxU2dJAd9TtaYMg0T+t2sJ73V6yj4wdXT/IrXy50SyRPfWI4
HLAYXBwUzksb8yDynMKu4h5SbFYH9hYz8bESCm8J8QccgzZKf56CQcSU2j21/K7h
yOEjgH71uBC6QL8hocTO5NWGK6Qd0LEB3KsnRw3WBHXr7UomWTHFIJvSUIR1zrae
ctDBR2H9Kxew7WgoYGrUHAnbo8XPEjognlgnDnkJ6zK3eSNI7xwoO74rhX3q4Jab
CcTNhvUWJmUc1mEwf2HlOn2ii8MB2SVXTmyBOkUm7nma/WjLuoXV3UT5UFEHMpfP
kYfzaRgalHWTxklacJpHzynmDNAFFdXa48iEVBax6KZf4nAH3OCQ6T7ZpSnP9fMF
eIfUrtmcG3nsgY6uSnpxHmsrSFtcQJSPu8bYbEHL7OwPBEvtwPcRf6J4SUo5BkOh
g4slabmxW2icRAlcP5MnCPnnLh6PqK99yQsXIDpfUnZ5PxG7lavMsOyum7YEjKmc
Nr3BcAVwU0zkIdsCppD9c+5TQaktXJpvegG5taS/9vyx0xEtBJ02sxa8yhBtZAF2
rQhu2BRlNSzEDR+jtJ13ldx2rCTBPuw3yw6oYL2uhpZYkOTTUh+CHh+HGj/r9pCc
iMmvViq4jhBcBgZVntHGwEIoUAkZQ2/O/VvxamjwMihL/VDPujynLshWPBuSA9FZ
x9GxOCNHF6bS5QxzlfkA0mRO/ZaDKnx6kHUENOKf6rEa1t8LFvtWdfyjXdTzeh3y
eh/OOKLn0tVo8pdLv/wATXXV/xwtjbN3BEum3zL1c+sK0evbus+4897L3aIrYzDR
wn+3ujORnkqWN8ORCzQ9yhdi1XSrqHCsV76UF8RMwu/5ZL6JpFSlFV1+HtzUBZBp
jJyl/pDL7ZycF/4lr9ZcS8gYwRuZGK0rW7pDYU5k0MvDbrSLLBPNmhHWFv8pXtLj
DXJiql0ZnGt72Nu2tf79L3gX2XbcdxR5EHqzk+ibrJ0xlez2EcafTJ4S04EIWaUm
uW8IZmhwvMyUyAequ0wUitaZUqHd8C5POje7APT0kh5+G2V32t67oqyCtTkTkJl+
s7BU3FZy6A9tyAo0o+FKCYa33HzmEmf9f0yZj/y+6DPRvMrG/C3W4yXzrWOl+4bU
boNGmphGHifJV8LlRTCm3dPsdgZNHHh+USwwwyycnT+aM3D9k8V4Ki8Mb1Qc0am5
cM+sY0zMrOyTCi25aAA/wYZD3KGLkdUypexUabl2NndmYAHbGyIelT57BkDd/yBr
1xZsTo6NDpS04JxkI4PM0a6Sqr2VSCv6EnRo3Z9c/EioYrmFPs+Tu7V1FY0BPviH
98v63lbtmGyHzK7+CTB1jVsjVqgDm6me9d+zoakbB99N85OTP8/8TTMJboe+dphz
mOFBO/YjMAbmb5itvgpEALi5O3otyn+B5E3zPPdhQwIjtTNhFM/jkmVo5Gzas88I
O2oLri2MpuzsI3jompNxhzlB8/rH2mz0uhTuSAcEt518CwYwwlKdKTdOPtr5aMJY
BaFn9E/1P23lc9EXT79ZCCfpOzW/QCrs+HIdIcEoiroYYAwswf3aIZAC7Yr5Omws
Tp9wRg1qIkRG5JgxUrc6mcxS7N/sPi0OET8lDEWkF47ioGpSbmqQNsQzSHe1kEzB
d5TKkKSQWWIT8zcBCcKVtjji5Rn1sNTsIKV3hEWuHNJNcFFKyDjV8vhmTfpkd4S/
nz9tpIZfBtr7MkT854EjvAc4MJ+LNFXF8+cY5TWUJeaAHkPeA0dtj/I+J6v+Jbka
vexcBz2/JjzVZsZAhx1wqhOs0xP67PZCP5DeQ2hIZaARA+nlS/PlABewizedJ7er
/4YaQN4CZtJ4FccgKOpbKmhE3mkyS+1mgEr7fVfeKBOFzdCW+udjZvTiuqc7v3+1
UnRn7ii+krhgxs1Zu7ZfrZOkItZzkm7eD5jqFbzNa/DhBUYtpqNefjdX+AkxWOaV
Kqek/sF0B66wrxTy61s67o/ZiDYJQeVCsBmuTBDKmIlyD/yVEnNPuM4sO4Er/D74
jsm0Lf5pkqtEY2YiDQNDZMPKJfzN9hms/tuggUJ7DzyUaHpq928lRbDfYAGlm7PW
GPECKz5s6jBdYf7rUt9mFS4L7utvgJO4AGE1Ij3/FJEyuNJzKFEj05v21hUXJCkH
5dBmF5SP8UiE3P33WS+LG4EcoQuJ5mID5mVr04ny7FLnpHQf2XxJRIcBLU+fq8Z9
W+oUgPeeqwomI0F0tHdJUEou3Q3keHEiJhsoLIeduQ49cPoqXyWxDlcST48q+3NA
hrgYFNi07ZaBulVFnsGithdZabYU3ryu/B+Odvk6Ry/+/IXOOq0OVDrV+WAU/sPD
trscVyXGF+J1lE3uUXioq1XC2joDYufME+b03xsq9SbANsqQgn5D2RClJynFoaoB
iSiEO9XTejNc3CwI5cEg8+YxQi2i+443e5Pt3vtWpX5bvBWxq3nvqKMCJ4De4Qb4
5a7yvPl/Rf8ORbWsVNr1SnLhSFX9vWLvJfWvUE+zlJeaYL4KXLzddvsY2B7233F5
AO1Gk1HXAG7WadU1M2SI/4WUXAn03T3kJLA/8mSVH+W+Kwh89B2oKTP1wk0XEmVA
Syq7ejZF8GJaRkBbN459mGm3w07txRecfYWhhH+qoPm79HXhWwfq+2B2TDkU0MQJ
x1avPWWaHZwB0DVdPSfiJljTIzg3GApVqlMnDwtD+nw/fBNpjBSHSG6PkV+2xy99
nH5653zt5Rmy2Cv37quo8MCIc6tW3/ktIkjVEXv8QgIgIb51ayiGYCiRGB6OLcvS
St2DhSulLTS36tKZS16ReAc4u+QKCvsMSwhDBXm+GcxZmXLNFPAzWQ/n91MjnMcR
QZdgclcWPl7T2x9z3f3KYOluYVP4ShBa2iWZwL7X/NCBlEUBP1fKd3Q3EDKfn60D
Q/ilkejUYUxGZ9sMdiUzUMcCvYz5zNfByHKCY53ySE/6Ph7iJC57Py7hqgfO7OWH
NsthgW72mhPXjK71G0o0VDNv1Vx/zCTqDn6F0pATI8+Gu5EWgv+1qFMfLmVuEoYR
WKWC8kBzujL5+GG1s+bGxTPsYbw+zk7v30e3ikQOhKCitKdUu5brQMArF2mg/q0V
6doOCABqTBLRa2PpSGS7WnKGNs38rKkpUM/hznxpUUmVa6rWVqbYbDWj+l3pY1K2
dxgsVu848ObQLXtj02IAG60HwIjbvehO1UW1PqMI9j59tIuG0v4m0srVznstKwUo
MYBBsJiM1w9th4t8JU3TyAKRTRJ06dG8rTVhDOxZ92MwNpNweiNswlZUYRdI+pZ0
FcjQ1RQHNcS+Obedj5lu2ONOW6W3WYeyPYaVr7ztb+Ka8Lm07ZUXW1PxBxtdQAyw
KcCYSbKYDKawT3XfmjmLcJW5TQwTYkzwt1D9D+wcl4JayB4T7mQK1xH7+bUtkTAg
nTwAa1mVIb16suO0y/6dUTYXDBBHAGjfyYNoUdRe42qw/xCWXbc7rtP4Lishy7mz
sEbeM11lhvC3LqJGvcTjrkmKLDDS/M49aJ2ggrO5bozzqG48FTQ5IF8nCeBptLl7
x8XWX/HagwodHLcT5vYSQF5HfQV3Yoe6SwuSYqK5m8yME6thcx4RfVGerZ7jwDK4
05dwROqXq92i/JYjQrUAXeAEBKNRrEiNIbNDWO+WMi/W6o0loaHCbGCCaoWnBoDo
sx9P7RvD2d0m5XVo30oFoI264JFM+VU+iL1dFA3Y+QhOt7U5lg8WZWy2sNyWN+mu
t2pUzMbytYSsc0kmPDeUbSo2fckPcSHTr6lRh93rvVxeMS+R3RND+ikO5bhkOd4v
id3Q9v0PAHPMUwkQiF8IMRAVWA/F3gksiO0E276ZpwPBNppwWTsMS8O7bnIy5X0r
sJqQ0KlRfyjTeFJ4jdN7oxlsp3I9mI135QIklQ+ZZfolOlvNALuicaA+23Yd47u2
SHpoScMyHHIqBAp04KiirthentUykikxLXgJp3rzhRIXlmiZLINvhRT4WYObbYcp
8iRFLeUflM/zMoPvfjiQW+D89nkdDWYZuii5mN+OG9nQENZGJWj1w2DlKrsY/krS
70d7/hyy/d7qDImjyUUnuHIG2YFGYlKJGeihuS++Xqgli/eWfZCumsVJ5LoC8hP7
MKosN33r5Ewni+ehSCQzkahho9UlKtn83CpznhAeIOy0JapRtkZR+e49otG+i326
qLfRoBr49seiV3q/aRZAInFDwECTnsqhIEtbGa+UeBMDZIvDl5Qiy02D51hyqDPb
VMAUYzC2/QcJ2XSJG5K0SAVxiQLRMGi1LvLJ4Ivuf65gkCUfiHbd9PerFx2t5rTV
ZNIl4qiTg30FoiR/lWWggdJwB86fSeXlJZ/r9Zf1jMJf/IFXZmGxKJ1THIeNf1D5
qg3xBznVq4BcbvK1uO3S9M/bMKZqK22YsHNOSQvKX2HSfADEPVNl/L5xpz0gwfep
takZpMauOfDdrcMzD9OeLJO0+x8t3HWDG4I5F7sqQEVQ6lSDgkc4TR/TzxU8Q0zN
iePOPqnhDFieTIzfXQb5Zi/PmKO7TSVwhQ4F4bAf1xTSz/nLUR4DE+boO1TYol4Z
iQxLwQfbN5oJbILLUF2t8JnT9fCUHJgnWyxUkHI3K57C3D41ECPfxG4HcIkjJqgd
KFGuuDtQ2jgOHu/7F4N3CcOUmmWoHbHoqbB3DLdIDsFfjAzWJhRvA+OX35C9aOkk
PIJwokJFSJd16fyTincci3GBSfco7UnuOppsByVpedgW1Zo90ULLtXa8ehSxPz75
zQPqiGjMkUCRHuwAXenE8Tv2rEx1bjiLHzR4Z2wOlmjlOPtxOAmTFwyZlVX8ock/
K1JvBwmNPbIbFk0r1urdxKGgLfosTSNlB3MEffWZy4KTr7rsg4Q70pDuE7DpgmxN
DReWzlAhYC9xjLxkPrEU/KqFFKfFoW4EKPcQJVBfttGnCjYDMtK0p+dceur7Ppja
3JaoObrIzcAZy/ElBwfdv1kvIE9VH40NWJj+B2maIP7gfyrwy3XEXl/9Rgit0+WV
PXUX2ydwr9dEHuQWTL2qfxGdDwXxTGZmKactvRX9JFxBq6XhPuIJKAEC1wL84XO1
CkVkh2Td1DFzgIWcVhlYX/XTwx5TqBaYyuGBUha3ePVGkKChK7aSfbT0Zsheufvi
W9d6786MFriQjtAHiBEdYzwNNxXoL3Ldnv+pOWen9s5D8/DuTGGOkmwqqFWfuvme
EFdCN2m5zQ/cYoy2b0VtJO2HToiQfTGvLqI08IeD+qBPbBIrpa1adCtMR/V1LZOR
1vPVhN9fXeMpXjMPNdjydNPs00LnKz83/MFxbgsjFMpvgstoM18PvYo+1ZR3CnTG
+gNUOAQyl5OIqIbCUwejp/GnIt1zcfb+bb0L/+jE6/XJ2sax0btutCKFQdOtbGIk
r6ShqinZWXfC8vZ+K4S6s6mv7y/4avUiHQUvOndvqv0bu+hU9b5OqUfvkZo/hIja
WK+LBiZkOI46g4jZ/AxP/4px9nCJBdsQC41ACaeO39EWyDNt7p1nCw9kwep9HUjA
Grpz2vyw9EWAtqrft3yTLh/I+pNg6hubtlfscWbMGQBZdcZMGqlp0lN4wlERLXV4
XItMIyGLTHitThy9AN7mBOPRAr5F46Y2VV83kdP2FCWJnGwLJlpI99NRE0DXxtFB
N1POfLbbdkoUKKH8wBgoO/aCH8lqEFx7tObRujEyT4cMtGlzdjDY9uB5KYvKTOUD
cXJm69Bx+REKeOg4OXqhsw/8xhVbcdldzj9bK8zrGo6dP9+fA71AJT55JlYXZw7R
fgMyddjeKJlsDWItMHqywM4L8AYNuuuDmdLwh36sIbvGLyo16nay91sn9Mvi8hVt
tvSiYc5ZTWhRqte7YYTqYlqzmdO7f3itWigLeA8X35UFLsa66l9OqIwdVIkeLGsP
OUd3nkfhRnPWZTreFCbyF6ms77aQaDPfkuVfB4bczyr3lurpOVf/flaTa3AX6dyq
rAOWiliJiJk78w7+ye4muHwZpPCWeMsyqeMZNXaTsf+fW3mLQttkqb0LaC5fiCmU
Zd0uM64Tm2fmReohCeXpbzQRilCQEWSdTZXgVJzf5SiLGvl3C2mnjSdM643Sc+C0
+VDPhiQts81O1jaji5s2lkL0VHo6kJJdCfEYshHo6kmywBUkR1VSmLTe+a05UyUh
ZrT4s3LIxcs4ldb0vqFnUAMA6xNGt20qHb1L8GDAkOiEtY7MXQc3fAJ/QGoNqHB7
gsc9kWbXhlij6UlP8uyEJFZfMz4kU+voO41uqXPS/+nSC50BaBP0QeF5WJP/Rq3M
jEfqKDjV6pTgJb5dG7Ps5ajQa9P3H2oZRkUtlAeJK6XEOs5n36QFero/d6yKdzzM
7mj/BaNZCACcKGRSnYP1J5hUYiVCtY5oipOsZN7gKpB2oQfBBJdHG7DIV5WCdY5g
gkG2Gj7XaTR+/GJ935oMK6rp3TePA0NxEf9Fm8vZrXO5yipAixxVp+tX93gSHfJz
OLJeLWGf+ug9j8epkHJ6JFKWUU4F3Bmwp7KTPLy0SPZfatAJjz2Dlq6iS3DGBW0l
hSCeIcbGW4X6hM3O/Rh/r2wyzYzBSGMibgOnfSr/KDojVfpkAZgxWjoBsKyTiHUi
21kZaDp8xTw+bUFsvrG8GxR/pWSfwrGIkY2oIV8gfyT0ZQgtPvld1Uai1bSc/Z0K
tJxKLi6Y+hASPGU48Dqv+M7lbNQfNI0QlQ7IHvbA3bla13ECozXIPfuCgRdot+rv
3hJcNkbhv1GCVwwFfAW1lTDoqTVJBvg6K83OQQiTcWBiQb4UC19ywFBMBW8VvH49
SDPe7FjQKbBgSRN4WoIDWD9//nu6nETjCUbMBn8gI+LKVKgI5JeYKLxeN66ERHOS
S4Um0BzhprFndLml5pC5WXcQU6sxlnyva0OA7NAOMgH10E4LmGBAvClFNSZM+ixv
AOxcUGWqQo1IAOLa/rUN+9aZq1L2kRLndWe1UZzT9s3ARh8sLdIiOa5P+5TzPxRw
24ok2TBQZ5QvhqMy/WfdnJhtS1f1PXowSiy0CCy3Zp3fZuEwge9XR78E/03IXuBO
EGJNRkrxJyDzR1VOX1yVXLz3KfBXbeWWrdCdigNV1yE4un5yS4eXF6DMRhyt8VB9
ySJT2j3y1mUBCUm4Iygi7cXu0j5fLaySE0JKg+rRxKdrpSB+vIfIhhnF5xcJOX5c
JbaLyT1N2iga7nWJ0S1GG88bEU1GukT0cyvRkuGmZH4OLrpeM5wwQEo7IGQozFqF
aVG+6plrix8tsxkEoNJkAWTNKwxnBifdSQVTQir0gK7pTLwnVm135eingiDqCNqP
3AWI2Lq2Yb8/hROfUX3Ow8t3DtMqIumxAxLt0/4toPyiSmu2/ziFQ8T3B36zVuJE
B2ba44UNxChy5IOose7SMXPrPGOEGkegyu6ms7ucqIG8SJ0MpOI9Hl3VWxmakAvw
k2RLF297lyd/VKZ24/RnCOGW1Eg053I1+kYgNc6fUeODyqtMr7XgcYPLh4ip4R5G
3avRGD4X6sB83IKzWEMgCW26R4z/CTkWYQSXT8KApVG2s6Sp3XT+iF1WhYTX/JkV
hzntpCUwqv/ch5TKZ/7ErUqGU5QCnYaOWUmEX1fepJbWRpnXvnKBKwiK6lEj3vtF
4A9sAEWpJNUvj+/NdvmoMiIZti+DqOVTjCix/sEsH+WmmwnSJJnLZJVF1msgOFDI
hBrKrE1V3tfya92oehgiLjYEOu7YXZ00PXuRjuFbL5RdVA4h6Zhtx9p0iqsFGM8d
24JY3KYbg0N0iGfsAM8gNKKdtIVPKWUjois7LOfomM9hvFg7ljd8JOGP+YbsJRTg
RpMV6tihRi/0DpQwkwTbEnk5+a8GdbayCW8HDz1NeZVJFVM97q7UEK8Ew9KEgUI2
Q44HNYfX5oUmlg37UN5fg2R/QE12lOJ898brB+LfA5KR+uuJ709Q/IZWRZ4KKo+C
ZVn6CwMnreFjCCpB/9sEFHSFxyK93qIkryEjdzIcKvuu78ZNj5MgWWo+ZE3z81Yo
twhfeFo8jMec9Zgnfax4wb5cOVTv/TFh5zaAxFmNqNEs30cdrIY9ouSKZdeI56wF
jmPRT6PHFMizlbj5ZaRdo+fQwwCLI1VFlWZmoog/UDvL3NnsiOuFba2H7VEnH21x
F24J22O1SDELpqcZMFWPH2h7VDPtWROXPCVA03HfNvI2XCyT1DhJ0RiIVND2Sxka
C5Z34/XcX09jhwHNDkqT74jZbF58eVjEmTLq/kEgVYyTEkDHNzgsW7SMMtb+eB8Y
EArIvZjHwt5e58iBlbOjMOH767mdSiJfzpIwDCTWRwAyJb+F0+9GRSodRszhrozi
y71xj46+SpO++xHNYFHjPq8hZUS0n6P1RFD16oucAqIu3QmE5FUsTiafP1srCDZA
1lrJHe0EQ/NmyjYBiK3fT+ijI+C0iz+fwSMPOXEj0JlYNbvDaiLSixyC/VOwYD2R
vQ3XXx+FAp3Toy0pRHZpITRFQgEg+IfUs7h2fJWXIZJB2xfM3JbBVXyLlz6s+Qhg
T1M4htE6FPjQXuOVWemhKTLJZ3c00uoMVTSVKeluxZDGqzcmq2pzBDywtX6RV2tf
CM42rswmlQrMtrxYKoJroDDhkPDzlijcDzcTiOxdnJj0uIFw3ttZhtW4W6IDf/EG
P8dRV2Dbj1ANHAW7rqnEaeOjUSTIj72AWTi3vMLdddOqZ5EhMvgHeROZo2UDkeEW
hmKgO7eTTxrJY8JGV+mBbAnzvka1eeYuiRkG8NwVZ2gxDzmj1MBhCEKGDIoE5Qz1
9XaXA2knlw1CHKleMnLQ1LPhpQiYvvXdq0MPmtwPV0FRpUNLx/fx/3+OkUXx4S6v
V6vf+cUQIZIBdprZ8JiH0l8cHG8h34by/JgaO+D7V9pWINr9Lfgk8Tn6DYaEhC0y
p58XPEEDt4UXazVJ1ZAb2r1rficQYXLNswbGmTKfIVjVJQrLTcutDERsm7+Tsoqa
8dOSMT23wxqawGv2Xn4kSazDpgYk8TkWpXEdxDsgDRjKfwWuiBkIc1oLnXEKAGKN
TlipRltdlr+9kw24pRb6bluSKTJEx8QR36sUBq4sFjGxgWHlQyj9rq0IVXFRnbPo
1vewNcH75oJtYAK04nYob+4mS2yllXVzPQAS+OyBMfG0/Xu951aBZ+qQfTK5H3jh
/NrKNiusyVey2CiHAfZ3yRmdzprMrqB6DaOs4SCiwVyi7WMXnES2FaCmKGl2RvEL
S/G02wMjBg4I2rXQg89QVcJk4nWFj7hKuYPbfcJ2H+3QlAEhE2H+LJmxrXwvJI3A
pv6bBm2lpky9OWZA/+QNHDl5WaIPycT72E5cRGMPFSQUjbMl7i9IBk9miWqkErXY
FIpIacqvZpsTI5s+6+IEpUQD7a9ZcEWsgh+3DMTQQrNAzGd7cOgQ5yOywYrurq/n
OoLCbML+hSAErwOZvfV0ToiLHFkojxnLlh3PLvb8KTXmme76owR9jltYeEHHASjy
hOiJu2Z1N+OCd1tmc7PBWT4SI+nUCmVtfOUKSdzD86htUo9gCqD0xf/nTNuY8doG
nPsfrEToknGM8oomIpLud8cNyqFunEora8MxXa4aLGvoq6ZZro1CIygbh1RkB5Zs
MSbB9lBSueDyUJLMO4FmQxnu1Wt/F7zM222A1JKkJMFeD6qU7pNZLy0UX5URBD97
qjE0Og+EUUgVLFpUCRWMgsUCU/JcOqEsWt00uqfDjUo4m31anP4KqHXYwXj4ZiRU
aCA+yFE59lB7Knx5oHYpxp1F0c3q3YwioidwnvzDSgQthTSSR1Zl3uEIJBJ4FmrK
W+n4hlPtqPqSqmsb9EWx3IjfOF8ygiQwdXmjVmJ82pPX1lS6fWbSpttOSHh0xIv/
IbIG2JRlge+qX973IR7yaEWzV1ju1kZU2U2S3+fj//VEhUuF3efsCG7Azx5oaxPc
opU+uUcC0QUMoIXr5eE30KnR/bFc1NrgSlqmvFOoZeJWbgLb4V8ccZgxbL2BwpDk
TI92Vj216K97ITAlgA18nXMBzgboXCAg/iXDzZuBc++nxW/hUnTLP4i7ob0bJeGB
ZmtrNFPwpJ5OIJQDwKRxmJ25w5MKNzZFcZooIhgbTYl01S63jN9xNhC9AfHAA2w8
zbPJt3v/ib8c1XACet8yOOplJdM6hOgbTSiiNw8xDdtJvbdcVew0I2Yze3uQ8g/1
QoctbU27QX3EDOTQSd8dp3C2hIkeMJy2W6fLZR/d0jFEwRDp93SCPiqyA/CKqyxb
13pEc/EmcL8Q+mUaVMyWtomYuWFrZCOwQ7cyJuCtrdDnPziKa/lKKPkEB+pdikR0
xc+O7eyQ5+PaZGfaNLPTUTJO82TUd+l8pLj46URnorpfKDTyJxfDeXpfcWza8qN2
S08UlSlebx5cwI7+hCvpxoVd0uu/HFwmqo4JXVZ95IhW7PlP8pyQ7bK29Jf1VUBF
DfDEwdx0NnjEa9u5eIeccLj6XXmfv6KKsa0gYGkrcgF2RT2flWkJY1JikazPsakO
CSSS1ycyBNbePrzbfmR5R0f+6lIZBbTPJHP+swFYMd6QZdQph13PKw9gCEri1osx
tw+8Ft79mZdqNZM7xLNsjIRB+frYm+1oWIggGfq5eY5AZ94As+imU8F6ZlgW/rCU
Rr/qNVdth5C+Q54PRc8vT6SrJMIpLMz0eWdlw1aWobi+oYvX8pTidQ37baLn3YBL
rfzsm20LadXVvhEhGmMm9EHVQamUhU+BESOvJPOrmKVyV5molZjqHgGBNGU66rNe
w9uw8a6PXgDYr4lWJkD2gwj+BmBe81EIDEb2OpET1IPNGbZR2I3QsX6hQvBkNR3n
e544rA6kVrLr0P7zsQwDVpI7JHjyvSmjlJXfpPtoAfG+0ynDv5CG6XqxylsFhRoi
wrlE9gI/jVUM+IlVfc93IMp4INf9MfsmYvo3ZU6hddQ18Ub+ackixv8LGdvdsuB+
fkN34QUb+qKq++AUSDTkZgUBVUBk1BozLTIRmqt3h9CKaADeLkocNRaq6ntpGKFA
Mkuc5EfodBvqgusw2u8NGMafcP816Su2gbADaaglIJvp6vmwVy7Dpx4ZM1mMM+cz
T4PXPhjIK99nCRhTPK0fzIo1imkl3r2r55BFAvMNwFptMlrqmnbp1vE1jlr4jXS8
up7atpX3jEWq95df3VUF8k+0nE/bTvVuRDwSsoK5wY4S2lmZNdhcnZwgqjioWYm9
a2qrlAiN0r0yoFU87ytcpetgTrGyobZI33WzvH7XqHdrbHy4lf56dKgC5FwwyfkU
KXDhB265WLXXTtuP2NkarWMwsdCARyEP9iU9zKcyceQ2CU/I8cTvjZsLXEXLG1WL
1LCL6VA6LgGXmtPwidoAoUEsFm4EPSntTxTyOcV2mP7jekDqMn72CGRo7YsEagbO
MgcnNHvgAvvlWDT3ltxSOMjqrJnKkv20vhgPUdzAahmhTZNhgmDhkeESbcE+TlAL
ZHaW3UZwn46MUkXVwbe0typvZiUp/qdwzXJ2sAg4lGE3pjGIvRsiNHIYjJcz2jF/
rIexFp9k7dHUFHu7yVurGhpAimUFnq4WY1BcGpDeytqysBCQ5r9uMYsgBCk1ypG0
6809hRImXzR1KRgYHzK0Vw9nOpibmeJvbZIv0HpQsJ3lPuZa6QZzytCCfzKPJaKA
Gkhs5QKYYp+0nCquXbco0bSRI9YBf0kdVhyA4PDNkA4JA5rUPprB4MvAO17Zdlf/
iXGRJej5BF0tJZxP/on2eYUWdJ1in2PMRWFgcBzV2ZGWg1vupPvlxO920M7dunEU
siWUt0BfHYVhhEuBqSTP1g4tqWK6pFRm0K2bwalvoTapRuLJPfU+SOTe4woAAuaO
TWVfZhH+TCJzYRS9mO5Px7YkFf5Lia8EDW5Bcgfup4fS+biOl+eRXDQyhVoIjfck
jREy+SBUlbf2/8l6/+X/GiOy+iTQOyPFe0R/+tlotXzhIm76M/MLkCSVyHDa1ifO
Q7e8FvZ5YfU7rMf3zqdt/yrUB1weZSzXQe/uQA3HCzvnYlaucK7aTYgdbUZvoUCD
C4Y1DT5XWnI7D8Nm8+ktrODNqDYkK7duk/Qk13mo3veeZqoc0rDcjpiK1FgW2Ztk
VIE9WAhHTc8zyvy9i/vRNlsfKprIclIpmbgyz+BVEAScwm2R3q6US3dh3K7zFTuH
/Ik6Mi2tEm0LVsN5xTz3plotp/6RK3m+W3qd5TFKR4oW4AwrVpjZ8TVaStCv5+Uo
8aHNE2O5lqqWLfi/ZXwPvplgmtNk4sBnGiH5A7KI08ubbNW4dPpUZC1a9zSpOIOI
Zf/RneDAmJ/D7VRwhJFbTabtDYi3l/cEbr8ICk2OK1xL5aDOSNnz/vG3mUweyamy
0GaV8r11HpXGZPwXV8qDMk+QxR/Z4AwFMuwg01gr+CIRQhJlFdwK+ssVJPtR29hS
9akIcUnGVWrUfVQH1P4Z2W80zJgzA5Fu2190n6TFpLkWMJVML1CkiQDq/XTz+gLc
v9lFbk7nGeGFcw3wCz3ntj30rHlV7YacqTYyaUVjv53CdHOGEOv2NPyhJgv3oyvw
wCh8cobzTm1P9zib5+oVZgdUqn3YF2Jo1j469eXLAfeemo53fk02TYlFztrki65d
NsVRh/9L0r6IZgUbCRmPhGLAR0sWSvXO2klZbnI+0AjdxoS8X6UYeyfgE+RMfobR
w8M4N7k6RN9UsxCeUZfiZbDSpyKZmZnkzLA93jIGghOGI9ag51Zql1zkG8cTsW4h
BdaIOTwv2boB6HsV/NfUo1lZMCYzjqTjKC8gis4gUT4XN/KWzfcHgPB/8PiWfh7J
8hlwT8gG6cqvKe1FlWfkjMxcRAvrH+SrZJTbgL6D1noAKEICowG968VJijBGvx4M
6TQw8WE20wTDndjf+qKd48f3LeJBwXf0dSAdrkdVycP0KsuSdR5Lo+QbzknmrAQa
ITglHYv6RYIPLSpa/SxB7Po3+dH7S5hxIozS7bfNo+jLR+/2p9ao0fqgDAxElzMo
uPxvwmJX2eflXnk+WtViTetuhsdKmNUwGsyKqpkzYYJZlprkzvhjKvvGDN9C6oyN
iPgwI5tK/OaEuh1tgTR3HkbCOm9lTccHl0xDLTWJrZJz2V/5rJO1dH8fB3o0ymiX
+a79WJRxjnxIWr1ysGlqF8ABQXqs2HjUjo6QHMADS1WynPA1HbSSHCfsCLcvaTPB
siQs5W8Lxtp6yQfxImnl3rFuiz/ptQGsJEREWMud3CoMPsJdY9eyAfZXA3/aoCOK
lNc9M2n/6yeukPVAXApTTYhUKafSu9//YnWXD92FMt0gMT3uETqIvHGgEFCmRLvB
oHf8mtK6XtUeSF0CAay57r3Y1bWz+x7E2GmDSYsJbRCwVKR4jOz5RXNdFSqh6v/e
BBFp9SgMug7GeN2aSr3vwVVnV+aPTAw5pMEDvNxqIS+Ft4U0SL6kWAesXCDfacqz
4wPM2LFWdYHYYMOf0IT3dpC17VyXrRvhRFfExQ2u/k8VbqVc+Z2Lz8QP4JLOFZSW
FqKMlxNuh8FsoBJQGpcxklYkbBubIknmknzAB9c6I90HnMWVOMCSgqS4bvVHq02k
Mdezf9lDN5dvPhc4L7e1Iwml6vuNtFY7ASAx7+wn89Irdu7legar2G6Uv3yb3Hgz
5NxQiQ+9VcWpQbboounaUBE50CbqITDlZxKCjq0KJYx4ZsiWi0MCvzDkBrg6I+y7
8DqXxaAGhNxIlO1T9zcfVw8VqFUDrCaJamWJB0DkRSQboYLsEeP7P5aBNIoBb5pp
MU/Wx+pbIJatosRp3To/Sd0KX5T0xmuTEB21bjDY8J+DlHfLrPUWv78SJrr0latn
GRqsbHYExV3XD96Ltb0r5QIH41bN9VVr9grFMPuGWlsCEDrNQxOo47IX7Npl++gx
GWrIKsetUGXIDGsnJlQUr9t6VYy8JmMh3f11WawvKV+9HdhdBsKNM7uD7VBiW7i2
VW8EK4WXiFzBRCZI2oTBQMOHU0n575yr0y4XVoyqIgsAuiq+mk0e3UUS3HkT4WeO
pVpoHsnH/VLB30DQF+OYPc8tjF2recUA3C7iemkiooQGektQw9uK319XwCenNQvQ
uwoDCCniK0Xbl+fl/+82Hf62HkhgHGJncdyTDEFEmVUKNDdrez9girGsCZ9ijdJT
GSjpTJrzS357bB1u++syY4s0Xs+vfc9N2aA70jzttA89BO+F7dNzRS/CWRcjUtln
+K0dINIuvu9wu5M9hUO1U1ToT4DWCx9qLYuz/9FqtCbf7KrNNIFQCqQFII8qSbj0
cc5kWmnMPv6nCphuKq66IQ6GkZ9imuTN3b5/gVP+kjqDAF1t74836v61CNrqeowm
cGfLK1fbHZnQKSb9RrkDsxk5yuQmeiX5eggZm1S3VonMbPu9HyOzwnRwel2IRVl+
Ru4+fuCEcKkzRvFiO7ZTCiw6WHicM4D3uHwf05xavJbsueczaoPqiLF2KZabpWeS
eKyi9ikBPItKSGnOzITBiFFsXkX1d8S4CE4v0RPF6Ym21Y1wCvN6B6qOlIpQup7v
8gy7QvTFTGh73OuMT5nsowuAdCYV/+qlI1l0RjqfBCoP0pTV8CmZzuiIisP/GMx+
C7JYTCnFo0XyaeP85Qnv4xWjmPKmYoAzXtHp1U53CKzsDWKww0zpjEeVnNqbiKVB
gQf7uYs0jkaNk/qt2DvvhDmNQMPMlxrC1hCPH3F6zbmVvizR7CYXDc7RqFHgkeH2
IGTA1cFFEQw+xyTV5cZ+9uka5jj9P6/IRUyPB/+l8V4mxO/eIFDNlUhTfCbnmnLt
ZrMH1VRTF3oZvOTPaBPAleikCg0FP1hhJV1JW0FQtJBE6ChNK6umGf9MPCJXavZq
9s2JlbXWctQMmC2CskZ63BaLMEMVXGWQjmmrVCEopiogi412YWoUzIbzLtzV3cyl
Se2dM801s9GmMe2jEiHeY8hhvDHAppJmC/2LvLn+fHSocmlqzpCl9v19BneBwv6C
5IvRSfktFypgBAOKpy2q1/eSpn4YzH+vAEN7YPf/2Io5bVznEcy7uAj5RGcLloAS
L1ytNLPC9WKr63o0XesVCviDjStDrV1OuVyP4KYrEbVANIK7unXlmCYlqwHJTRZU
jw3k+Q+scwBUNZOHdxQ+L1GFHlqbQaG8ty0zkK7+Sr1L20FUWhCpMAErXKZWgzVT
dnKeyiSOVEk1nFnDjqcuO7KaYwGeFg122OzFm3BB9ibYvz9KmxMina0w+2tqmBYO
8GJH7XOw06QFpzeRX+ATkcq7+MqKDsf875BhIPaBdKcme2w9YbIl8W1UHDR6yMpH
QtB/vSaKQFVZqnkaXBGA/0vyud+IXHafi+yl2s0X6U6dYV1vR3S/Edy7OsZtHfI2
vQF1tXRjb6gKgLgCesVvwSU7kyz+hUT424SScF1rSwGnnPrvQ4WrIWwcdRXclWWb
Z9dhuCKh4zv5MrcQK7fXK+2jEvlyLcKW5cHp4u0N6BDMeDMZxA0yRrHTwEqch0CK
YCHhpVbislQCnamEM8avHfvjQsWI2jHnpFDEl8FT+Om5wBmVRSaFoME2uMRiKkKG
5uaF2LJKGqNZnm+0OgNqFumdaomI7aV4Cx10laHazJy9Avj11XbBXrwk0ENNub8u
6tIhimHx5v+nWZouEGAdfGV/yAh/4caREw1HMLajORudmZZjU4Hk2tDpuCxV8d3t
z3YY4Ufvuy/weO5wghJxNuR/W/zsZKBPzynDW1dQO5ojCefKqxOYxwqXB7n7i8kS
keFvvtRnUB71UQQlVF/GhDTKSR4QudYEcLdYy0jI/vDG+ah3WDDVVPg4SH1916Xl
6awlLV91/NjerEjhgeu96UFrx6zcmnWHZ6W1G90s46cq8T2wMWGUB4pQvKzkjYfW
olC7P1jD2IQj6ejfVvB6Ig1t0wqYiQWdc9nmFmZhIxD7dGlK6RMDrey7vTZK8WMS
Cq4+bVNy8arUs1SSBXCH79e28sHKAg7cXUZaVfUGJPIYd4DFQk8nTG5YYpJa4OCW
XDDutTbHn5QfOLfReMUFKvv/pwPUXcQKAv2u/rQjh9G2tlXrLeFmjNlh+QRB3ken
Q5ncnch6MwyWzLBOluE5wjIaNT/NCpAC1rS3wZGY6Kx6wQBxTpqabokO/pFHdIx9
x/2IPTndP51Mx4I6c8rJEA99iFdxqA1zzVIi8esCCNKQ0sOTppUpwxOsTbS6NnoU
1gHG8e+t8GFCxYazVQHuedgi/eSWSh74eG8JNrw62e+Q/8iHTcFAZMRM9gPAArgC
tNYRumJP+n8uwEgh0TuWy5lstNl8efaNWuoCuLxPppV0cBJarJJIyhLPIoVEOVi9
9HQW6M0IPJAVDTaznx5QnUu9EWCeHUcHyEBBwkWKmvoxw0WPbZKcjuvq7uvI9t7m
ErckauCVr0LWOAPvzcAB26a8jDFWD6u++wSPojtIBTMmhk8CQF9pAnSA0CxsUgdG
dvQtoyMXGSMkUIz3g0iJvs1Nhr+cQV7Qi+LtKqPklVUXvH1xACATwE0nZUmHXkYS
jjCxzMuLsIVjJ6akhNMytA8w1QAgOMExjOOnZlJW2kTcFgJCo/UFCGbgt17tEHZd
HfVFXoANmuZUpR7kWHkF+o8ZfNHGiDWnpEhpoK7gZqHdflhMMwRFgs0KB6DizVX8
UeRuW2NLH2Gpz3ttn9CmvgiOh2mlvc+JR6YwYKFW7rZ97+x70xXnYgtNQbrcHc9h
SM3E61pwAAgcyXNAcZyr7eYPzZPCu2B+DZgw/0KovwiIvTCrD0Anssd+OdhOPlYk
1lb3w0pu0m1/GVwz/wQ+fSbMh6Y92y4GYgs5KNCKgTjtF51so20dHmnTICCM88AF
aZfbU2vqljVjxWw2cQOgnLGKoI5iqdFRMD2f3xVaQN0euUWn69msxTM2Fa5XzzI8
W71JdQ8jwQ9tcSo5UAA/cBnnUynKxEiYzqXtKNw8hPqYcKBN9XDz6xNIbV29WolH
H3zDzTdGOGXroBbiRjhB6etwKxNE6YRdwX+jM3ULwL8oEq/jKtH2dziWezfumuQ3
pR+yWWmlFgvU6YGP4EUjRqIz7kMTo9tet2bFhwFfc6pTF2DTbypd8Eabi1RMjh8G
hNqvtPxMCQkoBA2INAWHt/cQn26apXG9Pz17vYRvl13OIzrCgrwx/1PKcAJKCwB2
eYv3Tl+g+t0OxOdkV+mK/r0Xfjzs5ihXM4xO9M0RJE5VSGcxGBI+ilLBBFZrJs+9
yKV5IAwx7jieBhwQBiL+1S3xGi2cACMZ2JcyqR0fWBzu1zT3fE/YZ54ZMrE/+lV+
excVbuPHsYHoNtrsCC/UwSDJCdBuxCsPxISMs1TzmfFZMz49pdA9SoS3zpZKjixS
fVV4wEinAo9e6ZFM2q5nOx5S9lWFGW3fES/Hi5mcTebnoMzy0LJJD09B8B0M0nTs
sV9VNsJ/dOKJbKI8co5VfmOcmidy+K6wcbPWnYPmX28ewSjdtB6COez/yJ412V1J
6Sn0i77weG1LVVehHJw0fe9DOs/l8ltT4rULiVRjb2MCIiV8ueaJgqLMyf96PbtK
AfmorfFJdw8SIbdkKEy7V1EuzhxkcermLRQVX166cb7eBCv8g+xWEKwwvC/E4FlY
E02zLYGFEp9ntdO29j995T2JIXbjEO0S1oQQJI8cvPjuE8DNDo9g0sx6kL5LeURe
+30Eb73g9qUGUjBkUeNL9ABAcvHI4jKZqFx8/wrRWhYJXz/u7laKLh8910MM6zws
HdEIhwA/HVfYuzGwAi6/3nd8P2eKKhLcpq9xgPtIQxQ464hB//bpizhcU3Am+OnP
bGCcmCiVSAoGnuOyvP2R2VyS3lC5rnigTRqa8K75qCy+xfI5zFte4ZjKE9fofzV7
uQ8Xwgz7JVKjg0kk/aMQE2+diR1ulKvw7Ji6MayosWIdUMqUBrQk8e9VKpRXM4uS
zrWQM8XqejChnL9e/sgrZyoK9m0I9KGj/QFlv07DWb4AJNLXEhTDfhEcnLo++STU
RHhkL1xDAiRmhrdGRinp3qe1uE0kgHMWlD1/C8Sh+QE7TDGJBX2t9iIUdXtQpDp0
F+7WpyIU3UEeL4ZcdwORW2i6lM2yVJSYo0/De+l5AxLtWB64BA+nTGwl0LjEyucw
SGlYKNHqh0jYqE2+t9oZUVutvoUSOJw+X2pNxmaNT84FxKj1aJStY6HIIlNiRgx2
SSfsNOZGlIoL4ivVAvY8KCmjrKND2+AyC7sXXXfi6xOGqySs8XjEMOv+Lnj2wvG/
Z/MY3oMT/+8vYSlr2DAk8Fst17JtCfZiYTm1gowgNc0twK3naB/XPVNYw2c0Gi5P
p0YwfoOPikYRVOOmz/qTykjrgkEnwR2bib395FC50jAoNcnKaEV9HKPhrxVW4FD+
esPY/Z6KPlVpyqadK19xEPNZZ4yY7om5wbBfeYCMrIYk/yDv6wAYKmMbtan6m6Y2
rYeOf8smwadXJauFW5jQXlFmnkDx2I4ppNbHOi/Cr+vxoFhG+HxnYiIS0jYEKSEk
/24flc9abA3nPTOyXvPlCfG9N5aoRnS2lpURwF95vGuArWhvQO80Vm8SokDSadDK
RX/8wtlwYdqinGJ8EDUhTk1BLuRVTsI+Vps3EHokdrnF4vikRv82f7tkEQWv8Bqi
crZ7N33MT+mZHY914cvPkWQlBTYCjRed9ODw+l9q2VOxkWEq76ulMuiRk9TY1HWs
lWK4dxw5dfoCRqhpNX6VoMyQJaGIbY7gdCSR2tvXcHYRQA0jZp82C9simrhEK31j
iieV/Ov5t5ymhI9jvxooTLIa2zeWncs7psGPkwbom/pvbSCk3Y+e3pwoBHmBqQQW
wQaDXT3KxxAyNQAulygMvEFZdFF+KaOFvi+TmMfTC8U8QPH/Pw0O3urH8vlPO5LJ
Tv7+XrbUZWhFwwrtYKwuPiYajgIT3h6Lkb5HfcRAEBaSPkvM3tUx6BL0sTZWAHcn
ra57O7n9LKzcm1cfH57bjRTIbvDp9tFEsYVVvvknJIZhiBL+hXb7xAsTBZoLhSS/
NJoZhzpyjVQwP1oQ3faq/C0Bar0lZGBfrzfRk4SzkEMSo7sTdUGX0JIlzZIfFMKw
AdUNEA3j2nXM0bjGYhFhCpMJ5bhWsWzihV0m686arCgDtrRkuxcgl/AYUzmlpzck
S8lfZgcA00o2jxQ4FTIHXITL0aSc1q/2J9lGUgtwyyOnH8RRCuXl7MzsHfQC17Tu
/60KAF13wY+KmmOY8cbBfzTemlgKnm75r1Go841PBboeBPRgzRXaK7G8Iu2Rdg7x
6xJGFiTpxZr80GAVSU1xvjEiViGtyhyp6+kV7DVQjwwXYHhuGl2B5oPf/djN+6dK
NSq56Zg8VcUgFj17b9yCDUXvzZE0Pa9v4+4OS5Hjbkq7jpa2BCVg4Q6qdcOwyKEa
unskrxuETxoamo4iA4v55hgVRSerNYxwD2pCflDbmnvi0SeZdz8EP2TtzJllGktm
e3+Z1OEaft5ROk1QKYd2vHOA3Dsffe624bzZ9n6b5D6XBgbZHGQGiqVEnvnr3N5Z
IhGMjSwetafw5XgDPTmY1Cwb876cGANVileStDiJfOwkBasbqCb5vVv7dO2FGHp8
YkgBkAj6FttfTsLWSUQzxem84eMgM4YWj7/JFtwLpXEMcJys5V6e44S+GFGGxptP
p3OWO1K3x4Y1jQQCcP6AnT6ien9y+TsrcaGPvKpjGCMzTD5R4vAHxpvu33hbq98w
wHFdFfPfjQ6URO3iYqvnFNiE/Cp25MjAD0rJtz/J4R8BEu6oRbby8pABOLKJk67k
GxRQ5f6g0n9extLA34B4e5UbTpLCJD+nFDhljWnuwxZUm2tapghEem4BRZzAFQPO
XCzaspkpIdgjmQp1IaBIZASEqPnF8zWyyhGQ/IbajdZEf+u5844mKijab6oUTV8E
wGE01ucdNPCOlULhaMGEiP4W/hSmF+SeaN0AqhjCYQinYs6yrb6kQG+uDE6NFZvS
3BVq3oNWYlTsocqmxbO/WeVYVC4E5xW02SeJnSVwVq1iadYwyyNVmtpRy/wVzoLK
8TZpmtUU84xlidchIPE1LwpdHBKQib30fwyNXxDi5Cd42NoyREEWEVYH0GjbzMQn
FjSvf/LKupZcvtKNqqWJ3FAz2ZFUUtG6O96MW2Dk2kK3n5zk0xS7wChVIX0TFqV+
9FL52EBZuBsHLx6sryoy3ucqX4lQUinGexUANtZ/L7DnOl4qLYmRpoQp7PWOtiK8
TYP8iXnAHBpIyITgYJgNI3PHGUXU2i1C5kxPekX6TFRITosiL7h63lwb0XG1rYm3
X11iuH8DZAMxw3GeQq/9V0K3khunKHFEaRdGyGjR5AHHFkaLq9otWPecgEeATOjr
AZLQr7rRxuo/eJ5ReLdWZgbtnfwLeJGUPlZFrCgSq2p9irKvnt+6hUeoKKqj9laa
LOJk3JuqRoXQturjl0q4DC5jbLZ5nxCvH7N+R+xv9zQEb6u8xic6oi5+G6R8WVzY
bZ7MmtOSai8O2zauQXCQ3xQUWCJZxVpm86q3OoqLj9JP9PyX1yclfIWO6FpvBwzm
cOCW/nc8WkO19y2ATyyQO3mSUOJTMknVSG3JHJ5yC04CLs4WmgXof0XkPeeyPEH8
949UjBAWr8uIqaKAAFd99FiE01TuXvQBX2Q3izO3R4wsOGd7Q1OSvIcPGIWlsaIs
unKnEldHaPYzl9x5ILKgWJvON00VwsswD4fHYPbYAr1Kep/NNSlOtkioKuWTq/3+
s7wC/Xj3txYyAhNl5G351X6ZlcGoNO/nwLV+OJeSQlcreYIO+1lFZ5nvjbvtu3Ni
BDFRsY6xAm0/eZC+MVpzWyfcxQTq59tes73gGVjs/vIrer+2zQOvjNprxQVNP4XP
BSdUsJ1fkHgKok78MaSGgT9nWmOcfgAYBLnQNKL2ZorJkA5yhiTa7UazkmO8Hmbz
jvx22iQZo5FQs6bnImxXkTGiFZ7ShfvuS0HgXvHWiRhJ05NKpxo/6/3KDH3DOfno
uMnnRcdsBK09FrmYAIs2+VUYeVrHxuksuExcpNyFCX+2sD8gEIE/cAoIZRCb9M62
Pr/PssJ9APCKArd3+8ybb3MliqYLY2NM05uW47yyQAAN+8Pgze+Fcy4ACVHOdgnH
avK2eV460vbi7cQN938Til9cTkdX9Q1E7FNpZ0xbUyMltnPRp0/oDfp7GFVYZAqt
fZFpZidTos64p9gUBD9BTOGul5AaHvQ0oRD6QjQ75TFC1VEkzmVMJNW+DyNrScFM
dtWd5v9nelZZLyLjaZEQc7cbkWdMgE9Tkx6x08cP6AWK4E4Q2WXdATOyrF6Fp1oj
/+ckKe7QvTLEQr2IZ3QWXlNywlUATbTTcDZYmhy5jIPHn7WiJwkjOhgTH9axWSsn
D5uGYrjDDwVH8JZQ9Usyj7o7qio+A3J+nUTw2MnT/k2F+UJYRnZstGX38+sMm+9Y
q+OFD8NhDFlpuS7ovMhM2PhSexTCW0WfEgg1nAy2LgB8ghUHvVsxeQdTGgOnMI67
bq+asfQhOm5ma4iQ7tmNyK91oytI4IM0v/S4ifoz3uGXnB5xipNRmmQ1KyB7meyq
dBOb8eknl7oOjEbvYfOrEgd0yVFsJ9WD6Rs12kZU4NlKCmBbpFM9sy/6O5b+/o0U
wX+TrFZntO/K0Rc/lyivM4B2z6kIDrNWTzdgzoDdhzW0QXIE4toOrMTZeJr6cczg
2u2o2Iw8axOk3eqlzpTzeg8R4KfOMVGfCgnTd2s6p1BRVdo4R7KD4hkq5OmgASH5
OZK0OaBwUOYVYzRTkNfwx/CoU6x2+v7dDChUQ4GsOAriO6Mh+8aTd/v38BvpzMOs
yhZ3doWsoU13JmOqfb2Ggvmpq7QV33SmV7oK1Td3aDCmGlXCGz7c6wiz7DC1a/3W
D8J57kDyYFjTugNC7SU0+IKpO9F+8pIoLmVottE1M2R5AQM82Z1hDLc1mK/skzNQ
qyTZPllUBw2ACuYWM/P5kzD98IDpeFvI3SNHDeobjefTqZEd4iqHEe1hMby1imiL
FDPnrZfaoo8F9Ln0MHOC8ER7/ZJFq87hKEJQIsE9fXy8GJMFcL8zyALgaH8RAFRE
4in9CxRrKlaF7lBBPARrbxxDGlFD59YEDZsZBDYnngkzC5bwtHtfmGiEIbLnmdz+
G/91k2wh3V1DlGECDTRmvrCDqfeYzFMwHAgdi7VG731jBiqCUSV9GkF2Wz2wdBSj
Hps28y5c2Vkbgt6sCmACIsHEPvvHucu1T74nniRBXstgeJN///z8NH6YTJPj1H3C
Xb4tW1JGNk8y/XCKoywFmHpcxRflY4S02QHix+eFXT6NxI5J7a/Kau9/lopRoTPp
BkVBE9wg1y5/DJEbAQDD74TYmc+gLk3fnxq+oVOY3Ps79kCRC4FFUex2fMf+9CCs
jIFE9/vpW5BMbf15n4ot/QSpkbQgat3EzB24Es78AQn7r6LtdtqmIFyIRtiwnpUK
5PJ2uf0Q8c2qbvKY0hNKiysAGaQQngofkdrAsrrgnYCQQs1pUKmrhgtKSqoVeCEX
h/gcNQwu7C1e5yMJEQnunIIkq2SOEk75DUq9pgZC6b7TAR0eHxXhWYt54HUM04dw
X9ORwz+9xWHxXswPnqJDbVMHJw0SDR0KUCqIdG4q1rknZ3tVwL/T2xcqT/hS/cGF
fXmjuuGK3cSG8w4yCqJWdV/cfTlSJn7vs3MFO1RCMsxeoDieRe2/m7oKhC3KREgw
ieZR4XeShz/HXSYjZbSW87W1k1HjQI43wz1u7pBRH6rHqkfTCflvK7ttUIzKjzWP
FW1XPycFhBPboyFrGMaFsil0MFOsDqxkUElJc2q8w/TQi1jBMEfMMwLS+dNRb2Zj
R1Sik1HIrVVtzjIRLdSI3vIPUj4L3Dvq1zv6sjQEmYrJ2lsHFtXpCC02VbMyy7iU
2D85Rf6ZZkl4oAZG0pSp626vHBywMBDWUE6Wiw4UvG1fsYAj6MspKD2v1GTqWerG
P5Sclr4OwWNcUnMezJ2x9y2S5grgHws1ZEB0nzcYlMHhltCl0DzrQDXgPwcjyOWD
lPZqAVPOu8LBqq4pv4F8LzUBY3FeUUlsRcLDUp9LD3CzW1YIo7sWFweOQG47QIhQ
Qg/DGPqu711lVVMo/+Uhmh7/PB900zhiJJ37CNCmSx9nct1KL1V1f/0YA6mojEtr
9SRqI+EZUQYwHLfmuY0yuduLvC7HxQi6dDassL7o/GcdkgrRASVyEXA52S8STz/Q
XG+quLgxG1L6vPLj1CwNHyOIDjEV7wJCctvT25kiqjzLAHZJQnZ6CbUBrENA3+qp
eHHCktd5ZW2u4E0edxIkFIcvCZzGZgjKBMPf+h34oXG2f84HV+ENWeSmpGSOZlYF
jxoGtCLJOKawzRvMHDJvQbz/o+gryv7Y9BLZUkVvQl56IEDnzzbmlWdv+r6pLi9h
e0fQcf8eB6ZnAkqM2L2iJAkBOmCu7nO+AzPvxgXiZDioOiztjPTjBxXu+fr2P8yA
INdjcy8jVRR0JbHlmll0kbn3LGlOM5V70BCPFFUnkhQXA90IPAyNuwe2M3yZWCVN
2j95c7CaOMpEdDwy1HH4d8F+gDINclqn26pg7I9jv61nfKyBASmDfPAA4z1M10Rv
BraTC6t4TOr871l0KekABy7Et8ri0TvUJCXLmh28yPccTfxnd4bFizkzJ0lTxjkK
UhCvTrCwyvn8zJwPY6Qi0Q+NVZin7QpeSMO+DztpLiiRFDQmPycKTWc42u7AVNfj
Dk+M6/ge/PhWhQDU5RvVy3B4bN0jE1uPZQqVvhWI/OjtS1Kr9Geum8r9P9nHUTgL
2GFBw1xWL3PAazYUn1/d0DwUYu7i3iorIEUeexmeAqr+Z9VnK/ZOVhav/2DcTsAn
y5SbfZA5AIqvJLwNd2rUaRcTQv9d8wjUueKDXXNQyfehCwr4iXApNkJ1z9B73jQy
ybsbz+rxoxN2BEH0CtIZ9cgzQ2j1mM2NQt+bpWcXaHXiWNZpzLjdbLRixOEA5emZ
3n5ZDylqq32QI469vZP9sBJ5D+8z3VdSzPby2CWZs6xVX6qHGlzn9k3nIXUMSdSn
nCxlNmYDGaUUBx79fVolNVmKA8vnnfQc8mj7aG7/xTWi0uXK/L+jJNwQHbpI1cUC
Q72lqpxqp0LWrmPxo4VwLsBD+WApzAqZJEfzxP2/aw8ofN8TNs3mhJkNizjX+Tqq
vpiPEmAaqZP1giV2SdIGaDihHgW8YpjstAbtXPvDw7olJ3+x0Pl3Z646wq0AHfjM
KEyuGeW3k3ELH3gx/t68kngmv6jDcIVVX5xX8SVF+VXkfEpBkwF5HEDHxsUuZ7KD
wo3bZOQoxqXxPHJRBopyt8vFXjkpIfY8qq7t9b6CfCacfLEqoKouhzm/7C6bPYK8
dJ/URihbxv9+Aci7vvF9rNbRacaCBMkuGTVK1TaUNGSKsEfaM2ciOYOdWDPJgtjd
pS5d2YH+RxCNpBYoCOIUieB2EMZG+QfHH+jCRMmXCa/EoLfNNM+bIm7q8LBqt0B6
5zczlAXj9uPznBuGG5SpQhi6J7mFMn4ctCmbjx5Py38318abmAZnoGNrzWdANlmW
F5EesMvxy2gV0fVmuFG7282E2nRY0rs8vSlZ7U7HPo2CcLE+Ikk14rjWlY8OHVzo
cR3cA9RsU690Xd78U/3V/Y+FVq+GiVQC21M9Fg1OeVZxygYrxRqJYcvX/R0SjA24
xnBIsRobXEAL/dt8pqkaNCTQE+pVyiQtgz1nEbepC3OqR4qL7MTw0Q/jujvepPaU
PV76Y5SDvHQfpZc4diR7ikvBsyv4Zi5/g3HtGBJrZkZkRf4meIp+6w8/r+mra37o
xiXei91CSW8DvFbRLp9Yv1NWSorOd2fe91/NVwWC9CobpdFaQkPdrirYtWezPkqp
rfmNH1Tde7BamPfdw2tFWHMiSoqeOk4bU235icGOQAZH4fTOGy2KEBeC7jHxjpio
+GtUxXvVdfZaVWTuA+n1eOrD1sMTr5n83ZWlJEpQOKSkv1T/zhoC22r75+ybJY00
KFJBQSKFcBF7aPXrjs5p6+CpBGaOxkBDugH0iOoAfNc2SuHM14FpVv9EyXLTPaid
Z1W3S1GQN2P3jj3Fz6+W2m6Lc1fH5BmlSoWXFDMdFxh2zh+Cfyg+lr6pfBxnGC0i
T3ayYZqCqkQLjW1YR33U/iFfoQoFEUe1PaF8IJC7b+nmraP4toH1AWgmbNTCcVKt
IunTGwTI5RSEedMuL1uhqTPyvhKJeDLIojHK/nUlJ3ObgRisW9jPES3id+TQyKDw
x+R8oi8zX+Bx5U0JN8/W5zqNtXzsR8doA8VjDAsT9NkN28W9LoITa8aksWRaO8OE
mUX4szA5Wc2AF3xrZcPhcA8NO3kSIj9d/Mb6U8EJ99adKOQi7USWAeY70ZHwpLsJ
mBrMxhu19It6yusADxZIG+ZPUTaVQ0Bdy2y+3N3Sb5jwluUtgidO6xOANiIKU/aB
ieKtIXBlsKka7alGEYeSSGgCfijHJv2Q9D3k6HoOpgeQTuYcVfuo7aqcZ3P0As+G
aOv/poL/PLk4PAei8YhglhjBZbUP+p5zfcKH6el8IG7Hp4Dh7e36ayv9Wh1VwPyd
voXVhjWeWacMFfBWDvgAqGhbe0mAh+C+eiSQcPUEMkhLhdYbxOeOTkywZBxAbQZr
anZNJSuCjYHsciKm9Xfk30gidX7Ow8r+31gBu16GMDQ55I5bMMFgzS0BNl5ML2jg
yy33V/yGSRTZl+Nx4LGs7uCNEuHc6FZL/kdxpKEU2+gRBFdp9wmCIARRV4bOXeM5
BUWdVi99B1tiisTtQUNLPjpgoaVGRs6XKntG0aq57bxPTp8Qvw+++FvzeBq18MT6
cG/vQU/00nEEzsxfkI/ZEwnKCYh2wYEIY4JfpwZskMNw4lB/cz5+kVk6sP5aFFZf
aH5xmIdDw0J6lkULW2OvMi4Ybcy4HnltnVSf/aBPYobUFDnbj3S2I1k10BQYqLjM
Y88jHVO7m9iVCAqwqJ/iim2T3d3Zq0vO44NlRLNVycX4GzyT5PRzZ0LCqwNt1f0X
2qa2ZILmCB2dx0yzDZEolpsHGZex8Sm5C92CTpHwQF3hEbB/JzNBcoJH8eqL+Qw2
vXw7tDeCgmKHmQG2cl2iF2bJGwfYgT0DqeCms+yk8AyBx7QZEopTbAViXqXIT1Lg
GCfdIIRT3bLqGBDFEUlM8g2kwldWwdmFUgmD8TeDTSS0ZwDuplcH//Ov5dSzG8Um
3HvQMqAUmqNS+nsIA8rDtnHVmewDGbRsUBEiuTjsd99ngJ34Igd2CgM8omt/CcsI
rtBG5RPCd2HWESs9iq7WS5b5STBgIFN25UyTBw2cYN+GP15WZfuErKyVku1sAsoa
rwxUfOkYr4FztEgv1UWoe7S6pkAPROTUa/lhEqMgXIHUv76ISfZdadBn8QqDcfdA
0tlhmEPb5i7Wm90VFuWVAldgyj6w+slWy4ya36sCfngLJoOkMFY7so51/n1wlrvc
uzzI3HvzHz9z/Y1IIYxcUK+M4s4epX2saaTIUgPnzy9xUd4t9nCLSUCQnyDuLqNc
qULYUo/PMNAH75+8ts3tC4KUdcTf1ltd3OqwBb8wqHJq0kLleMpUo6lmnaopEwxj
uGW1tI0VHqCr9pAuSpsNoWC6sh/LIBLq8xde1FjuFB7Px/ZkvsaMQEWdLtNZ40Nq
nBobeRm/4wtmynK0CK9I1jpX8T1reyIPWgb+BhLACkE6Ei/GUqfsSPKyqH7cfCJd
8Nc1VcYvUWeLh2AdMX4CZxJX3NW/O/dbuUSMyhg1xY3RQN5wkLqLQ7MtslqBUtOW
jdAvYB7Jkdcq4PRmPTb9lflTc+EyYmUSZMN0w0XDKVX0Gf4Qf0Le3HSvQsfrarN3
q3tPMDsDy7nvrGMdivOGq2IJtR+RIf4sntOsMgzkFYJNBZwmIZXdWwzpHc9aTeu4
fF46NhKGXQrEuydn7neYtZxQbHKlPX1ktWPIhVz/UWvZGKCJa3BKZye33IT71K6E
0KzuGaQlQSdI2/srvzPTeaMzvtzqPrEUlhEqneSC0NtTZ+w/4xou8T4r1GoWzvmd
xrl8n2+ovHv8kkxeq0m5dn4gFMWdoG6AM21cuAFehit3Pgj4UbTL9bHjPka3g4fA
AQ0ZY9+0ODcNigTCtVaPAr2gLKHHnB1mveudsMj4qna3x4CdIdyDcoeTtXknY8Lz
E1Tlm1jjxbX1L6yZ5nZ8Weo44z68RedBLA6g17VwiuBOnKVqJUOaiVqKhwOTuSNa
bl1aUzW9z0227efCaI2Zx1aiNgn9AHlyOdP5HlIgdIhKzhdQZYZW5hAn+9wtP8k2
h4CW4MxHGc4jFoCppfi4l07/L0+dpLyzh6/w8vDwcnttTP6wIlwa9HWOa3ympxK5
DpoLYuqFOjDkFsIvqjDT6icFDs37jcxTInUKBhBLNtP98yzCgpS3rnyidpCVUAd9
astQ1pZvdoIbjlEJ6a+7XRzPSZRtp5c9Ybwhf4eyYl/VHZZGYvnXlodexho4nfcs
7PSwaqJwomic3OsIselHKzxMXG4k8JwiJUL+H+ZWxeMjAe9GHGHxmpLhEZqCKzCm
zxG8BPLeLO9DkCnjW/mnUtl/lCD70JYnLPRL+Ljh+WIedN1vHcxjnIijHOI0g7p/
0TRbAnHP69h/d/CCmpfOXJ4t9e/LK0HeJsa3eofLmYOj3roMk32EQy3bPAsxjDYW
QJqKjuXSUwxJ4tbPHh62mI0c+6NN1OY4bfqcTbYVflReIT3wxTed3CuH9SqViefY
V1kZgfqmCuMZuspeIbe/BSL3uuGCS1NA9bJ9a8qY9soau37ZdWBSyhJ8RYCbNKMn
RSZKpCft1X97jajf3nAK46lLv/3+FzCEkpttoirPK8KrQ0iNpRyLmwfMgtl7BJiV
K3cGLGyx6JxGRjqwBPOQxCtjo0sJUFgcZ/CD213GiSZdnXUfdfiqTgWxXvMWtpZu
zetL4D/1LCWhIfBg66MHKGhZCVEMHFaAlgAnVm4fXufXfBxDxE29NQIVCGaea52h
3mm4wNxwZw4+fRDfs9j2DL3Iv+jYhmuT+wiYHdCbQbdUYhcJgEtw4i5/W5a+E/fH
E+YsRCUGC1UM/r4fDxp0FMpucCTfTLnEUgKRR+5FeGJcUtg1NF411Ox4acUS0r/j
FI/Pe7xNZkuB5DiSu91+71unCMQvikD5zTnXAJndo+yJ+qMOTriHLSEQZcXbXrhY
6OejAuX++GSd2/1O+1OZaJrNnj9z+ZEQiwdk/c6K5wEqtxQFMmARht9BMdUoasHw
8hUhpGNbtNSTXTtleuvxTvIdq/QQ/pFDZ6nk5Oazb0FvakW0hFdRV9nadoSYxD7I
rpqGZlgpOgnx7D3Y1weGaMqIWu7jVWvNf1ez3+edVkPNKqRK00qmTlQMCtbhT6on
D40rUNV8XMPw1ELZS0y57B6NAypLYuF1/LRQ6xy4CTfcBWa/N+ZBZCGNfvjQFA00
uF1LF04Urwd1RM5Zcj5p/he1uxqVBQNBL4a3NFqJax3VQxgruhRBvCkLoSF1Z35n
2rgEvUJuKEcRG8zBwZ3zpeuSuLbP1tmxICm5g/i8eQO9YAafmLSl/5bwmjcqtFUp
pecdOY63V+dVvWWtwzweC1z8y9/ngm4S+5suKKBAq/QXoTjCGnA5a82VaV7+Nea9
pkq3C4Zc5wJ+0uFv+h0FpC19IYVcQ8RsZP6Kce8qX4qxExFV0cLkFRIXE4N86fEz
pk3RzKaUBo0OhFwIMFYL34Wr6KybwDeSX0NE6sPpki9eJ+DfyeWMmU5MvStgOYEy
xe1gvNvCKvLbfKdVlK3hTRIrMYEH/Y1Fr6qxZ8Uz/9vAADGX/4LdL4YUO220J5fJ
0mSLapFa2dNbbq7GIdHA+qhmkaPQhvnw9yPBbe7E8hZb4kZ6z75//I9uaQRQMub0
4tfGd8j4QGq0aJpUHRigf4sb88wAQx8yJ7flIzgo1ScYxfwb631WlDIYMFfwRxRC
ZtZ+s7SrDcyOMlHGULoJfG6l54k12mCednuO29f7cXUBNMAd4IhhqJGVCyrgkxBf
CJLw9Wix2nVT6k3jzOX/IJYGRDFLST55tPasX6GuSR6J7OfWQfIjRlX9FQjouzXn
ERc49n6RCVzIrR5MKDPIrsHSmaDLrLAiMNRWvgyElwj2eXKsLI99bAMjE6XPuWJu
z3OYNpqf+1RuM6ou22UjrMzLHFrkeoY8wzROlG94arLa+9rS48TTReRncSlme69w
WPRGQhhLYKtkIxqrs4M/N/INfK2MiwSksk9FgSHQ0f8vTgtqHmEdmO1TEigbOGSk
0EPeRLunoRF5scFcXk0RuY6FVB+XZuJzBWixpOne7HMahzxvmDfycLLUhvuQ0FQM
LOPpaDi8eiyoYc1FYUVo6GXnxI1Ou7o82msQQR1AGk8zR28gFoytmYuGOhtC63m8
QzT37bYFgKKiYw/x3DgBnQy8kw+om0Nq2dyeu0+Yt28/HNqqcyoQUqf0vKqdTxmz
BFBIsTuiJM9sbmVj6ZVz9BjFQKj74m6j0me2a+U20IyRgb9Y3ho1veZkWcG+DNjG
L2Cu8MmIyL+hARWOOKEZxDHSduKino24rjWK0dcIOWfZgv4HdcIFve3tIKNdQqqZ
RrFxeYP4MM12iutcfjx3NTZdC0jhwmORNdOK3zn1OiCSvXUQG4t8fjNE3VUdYPrY
uyxltRUwgigbUXLWM2qk6gwrM3yn1/eqUboTMLln7DLx+ShKYocvf8AiImonI8ry
1RNyJ3Ss/dp5vQK0W/nYDz60Hsba+qPD5iHZ4nmQICD4CSDfw4BoOMdD0DRgHU2N
ZO5amBY421XL53vOM3wycCwSk9mSJA1ctYEiLA8WNCwlSa/iZ5MoF+LWhYQwKXkn
RQVSitJt6HeonqfuzMpfa7kx7DnZwDd6sdBOoGEOmSJU8NJvF5nRzw8jxHtKfQuS
myVmEdAYfv6mPa9MkkT/7mwfiaHBjv6046o4Op5dQhnsvTX928kHfDc7f+NXtrAC
WtTBgJgN1XdPz7XzHkotA7qSJ1RQSdoWcITIELVS6KaOVMZZhAdWW7Mu9eliwJUT
EN6ZUqJErOhc5kXKDzQmiXQTgOcN1fk9MO0w41zqUbTAIa7PBV4+ryQSTHigamm5
0+s7zEi2U1FZINAZamyz9vycM4t5crLDOSMiSsyj/PaEg3dxdp78vBJ5mAe5EL4K
uGXSM/eCdbS15MV7AUmyQux2pY5f5RtkK3V0hYmxlpvqpwICnC5pRu1uFgj1SfXm
2e/DYp02AUJnVWXUbVVxUnEPUBUbhpVsQhF5jB9pIU6WjFyHo2CjMYIuM0On3EuE
MTYfhqQu4padKGderepfqCCc7OoaZ8HdXubLCRDRCoABoloCAv7M0Q1XP3kwi6Ta
gdc8+apgmxZdqY/Wq2ayxxIxWL2hv0WHgCGG+f5CKxHGes2PrP82UYKKCji6RL2i
J7jzT2ceoJcYW3K8BCiSvnFHHtG2eDGKEyy5aP3YTTdnhhwdWVraAhsOMLY0BvDE
c1yJSaYiSEnYgwBJTWhMcH5wUuWp/r6g2s7vMuqFrdPkhy34RPIUjj8maAPeDmcS
NEkNfCV4Ljzu9UPc1Lnfql5R1NzQnmqb7S5h0Ej3nFNVkTq4cIbCD3XvjwP1o/jU
eiuz/1YLwEBIYw9uT5A6tD4mKSCPqTCSRXOiO7hA5WQaBaVNfspB9NoLIk2Ry9uC
MX0aWZ+Vhi6kMhh2taiCmesh8vh0b1FCp++bny4GUjgB5AnUeU1jRr9aEN+Xe4V8
bZoPhM5HSq7LTmCby2raAYd2kBiU7qnk2xC5xxXYKoJ3y1xOCPx1njoUWmP/1xmw
gNMS0obzbkROCqTlOXg8WNnmZ3zFc+PHmNeH6GvLwATC2wGEdJgEXtCJwOsRGEB0
U84s8ZdWN6210YpTPRWxin4CtaQG1JjPds9gXaiDhPOwaCTYOzilLLAlVcJ/Sjjn
fsjs/s5XzNMHT+5CnBoGpQ0uaE0DIEP9c3oXID6tyJ2+5QpkDe6ktyXY6GKSLOfd
yKcYCRZA/jgvmO/RUHXE1nuKis8Nj4stxrFLVeNvrOrQlCUZMI+poxFdSm/Zlw9R
gAgHVldlFK6Sd2iHnQ9nrdmOrEnkVK/Kkwe4OMqmwgpBR4YjrI0qwrf9B7phraa+
jusVO/sJDhpVyZO1pPH4vGb2gQUsdZsw1KEAFEpvw0rfYQoz5Ald0TCcqVPiGjAx
yMrCtHYcOkcTUU4lgHJjtBCoZlM722hb/oY/zHqRJn1wKh5/CNqzJSVZ9SMrP2iB
KqUzX8weATK9u7afB4RPmsFeb8Xyr9eVuty4uevd0XB6VH5ZKsGT8veoHK8mWro2
r5/rtneDVKJCtvNMn/Y6Fy2XublUJbTEwibZkvnhEKQH9YSyaA6GK5X+MpSYm8/B
aHgcfaBOQ2b7pUXLPuAD0acdIfkHtGQQdBUIa+QJCLUFfC8gfAr6yZbw7nU3fsxy
DMnHdm1M7gT6NJFwqvynPhsEq1FDF5BQ5gD2oOf9oD5slaVUQZdZvv8Y0LZkaN8H
vTBBmAfyUcJf0vXGOYS57fFzhycop3s7cd4gRdU/xEQL8+hDY99PDDcp/hoJGiYV
pjnsVde3gkJyL8dGPecjVRcyXWgY//nXxrS9rKudTUcRCGRUZkTGx+ioAw8Yim/j
mPcfDQfGpkwCNc3i7WHTgQ6l+h+IbspM7vIbcXKIc27Ye34gFxtjQM9AUAxVlgTi
AKOoTjtOmWYub0XBUYI1Bk2Yywx1gVXUFF9bqyYrXpuHdQ7wXm5nC9eXDiFJsGTt
vTtHGdSSeeAu72nXP/lK7Pq2+j0ws+V2WGSNgN7QBd85A5Yb4gy7kQSKT0jCeYYi
+PAZSWRHci4bmXtwXGOqQZGPyMxTYNfKpB6ImF4cQIt8MAWeEnWO2kgVyLbHYCQP
1gC2oIYoEb8E7b9z/lU0wOt4AiHNnttY4kK2X7oGPLXoIN5tv2WInPP7J0w/c5ec
mVa7ur5l6N4sT++blOWUqB65s6ynRSUNI2ryZbPHqTGuXJCilIZFjXOUGw1h4ap7
Kx/nQl9z9eOq6h/K2GkMJfJEWwihTxo58fOrS129kAgD4Ffv/GMiRRaHMu7JBdOn
Jc6nfasVIy11akLd72MiLYLlrDw0h1LsvQB1Vsg4D13txbdFVfFDzFHaEzg/2rNR
H1ASx/OFkzEGxCZqp9OH1LdRvNPNMi/swKK/pF8vXNrnos0CghXipwzbhEDlQ9Lu
0ebGLGV1CmpKhSH8U40OuS0XFxkVXFGjyK9gXJc5iB5Me+7+N7h+AVmXRmhgs2qK
oYUURyiYjoLkTQkYIhmbWM87LbQpGva23uKbb9EKjmuWjYB9y+Kyjs4anpV4d2zg
mpl62B13uy8qmopMg4WEubR7wcsByPqFaYTt+S3Bo09KvYPEt90fKmzGkJ8EoeBs
nI44YdccxItd1cH7itKdysvVDWqwUaZeawXfPdwCeXxkpCxUFOy+8UXXJHaWEa8i
3VVXwbyYc5AL8bNQWxNfIQ9Fm3B+Ar9TE/tF5RweFHNoOkzmHrnlbrbYqkol2U4p
7oIRDw+5+9yi/s3u2EOf92ZBCTlGa3UZs3bQwIrYX2ImLU1VuWmNLfI+wNsxFmTd
RafssNFYDGHHL5LyVFCrF1OJLp9MJQRqSoTxdJnTh56RQUJJNn98w//l69uKVHnb
tUi8I6wWLucLt7aCsb04hwr2WBJ2WrClqmFLhZ1Rx7ze7PspAbUHsOX0Q+fA/MnF
bR/Q1UKNJUXCpZdGzgXoQhVVzaTGjd0VusVecOEZYdrj+Hhz/FAvDqSmzSsbkKoX
ruAxU8s/kVF6+C5TH3rffIgwLjJIHpRCEQISdEXVPFl+vrTYi8iCYZrriLj2pWhZ
i15wff7wKW8eWDw3nWA5cqqAftbNlzNT+/X/3ieZa8v1451YGWu7VpwRf37SjsRI
aIX9pF/dWGgqbQh2cfHw6ascp1EYbIayEE8+Sr913+x0o0shqSwBgTPzGojlkw2A
zVSRv7nr3m8qIMhgmJ1Ikl5dfAuMqETukHfEYW+pskScetuaAbLbPl67HIlhKcXo
FdmaMAGog55i9phFFJKs1Z0SXwqibWw1v4T/HCiJ793lEzV4NXwnmfM+6/Po+CUV
2WcsROa0HWrTmRa81m5AIvoKW3/R7JXjycsVzEolYSj3tfvw9A7I3flh7gEBWjcZ
Px7ebznb5ZMSbGJ5bDy1sVOlMruAbUy2jG9RcudoN4tMTo7TvKabKboGC7iO3Qqy
ER0KTa8RDg5T1SWRXtQVBE7BawNigWqGwLwfrnh1T0aMAGcbi2BbQv4i8WRzCTJU
NEryqz0l+Sgh9vmKVALVzUVl6807UjbOR6yMxDyb4BzcSOGU3tufmV6KhmUF3lex
/XIsPfZtsfD/2JqD9R2fyug0fh4J0Lei5Vu+QE9yrwcaLunGYbwm/H86UQjozjl+
QmT9KE9OJIrML2GRqEVXkSmMd41gCHiLdRceARa36mvbf8sJHwAPc//kC4fleweJ
kOplZYKTuk1DIY9yD5Ix2EEXwRPcEAR+7iH0el/OkjXgXPQ+5p+y9hTev7fgW/rT
KY0pAsAhkitg6bBHjcLjSzMG3HyFOv8Rx9LTV2Ck65U0Xi8cERAoDEghYou5aa7/
AcKC0FI0y7ny33nfFH6Uy77HQNUjnrQJtby0DYNxcBTt+k9Mre9UZCXwsPWllOI2
jwcO5XaPOwZwp6/zMxoy9nrC1OMopznoEEEiELz3Be40WHmjgUi2iy+6anJPdaZ/
lAU7yeQqJYOk8AYib6nswT/G8h7M4DbC6zrEtZdEv+abjaUDefA/ajSPqF/GUs87
KRaRMyvDQz5Bokg+UFWG0rBiTgYhyxOp1/fzvkHCNR3Bu7niWwOnkO9Wn5tuOYau
7Tfk6pkF8N/nx4PHrGYo69iJLF1ohATgwloTS2ThQGq8z8QtQWHXpmcnANdyGGuN
cfHcTcn+GO9JWUUeREyd13g3aFm2p8t9ce1Yj345AR3Zl/mZQA9jz3m5EODCgpFB
B1/QzUBKqE/BGV8J9IU4PhIF/lWuYGL8FprjwXqdVFKKO5huctTs6pQRA46v02RO
9vfHc8JS97DwgEBtMyxlmDqsK96+Q6GmaWhXKtQjl+UCOximTBEPYMKoNsoQ6lcz
g2h9m2uR4sIUGI8IsM7N0cR8NHvAsHJwlzY02CxsFqeH3ggOfzm8ajTIoh8hKkil
L68bjeEQP9sGVZP8804wyvg/BRklWbtPOg6Ya+sCdAe6ZnORHHKu6+W1Y71yQU2s
G1wXgLnuwiLEGKtRhq9pvyvuF/iyVgsr08JxnOtMrXzRFONDWNr5Q6TRnXdsAM09
5xbqJ92GFlODDvmTThvfRTGMgxoaYXPzcn71T9u5x5BH8GeOMT/hj7SExS7FPEyx
In/01aIgsVMcoK8T5RVr/TNYIaSrErIA017Nc1dIH5RlhbtPKSRpxQqzJOEkgb0U
mJB8/XutJgFdd5xevG59L1NZcR8EvpmUUPYBRT1AhMWMOyLKO+C874UpKlh728oz
ohrWPw/olC8Qvx51K7I5RwubfVsxqVOulUkMUk9BlhpCuZ5aCJSc70xntpqMaHpr
VTot9we/Kt4Fp4XjNXHmORg7IjRv5mBH9TyBGPxa6g4jzMB/gFan1tprHnSHdd03
mvyWT4MGt4UYXgNiOvT623wJIbAzd1R9iVuRY1r68xjVl07duH2ZcG1kjTMO0z7x
T7w9SiSuimChO/h9R1aSBcldtKVV2yXs0aGusitNxW97Jki8RatfFVQsaJ6Eco1v
B0VL9FwSwf+rh7+ETiXe/IDu/sI7LocR4Lfcd1yAXRjpABGMB2AYsZp+F59ZNmPg
TppGp9rXznM+O281x3ZaHpa6KAhgAopZDJDdrpTD5KwCxqrJNyGXuTO5hNGSbMG+
yylBP6RNDXf3x+fXsrMFUa7KS09CHqkChCBTjQElP82pMYfaJJ5VG/5x6Mnt3iDy
o3gHlBPexnRWT1sVVuR54e0OuQWgJakxEHXGG0by2KtFi6XoJKnj9RHhF81/U6ds
syIRK7KQceu/5glTZ8pgB8+I3O5987IZuTB9CzSIV1UwcL3+XIsukkj9iwkySneO
BNk+WlFM4fA10QOCGQLlYqbOby3GwBlNL9ots4rZwGcUFEL5oIR+fRBolqsf8iz9
WwRTgYF+QIRfjSR7JKFhKkYdKfvzfI2zp3qg31KFbcY8x3/fVShxC7nmzmNLNE80
NjEc5l1EBhcoov1L6SFbfjPx2TObQoHciga8i7dEUO5aKdvgnO3k6o0/YCmKB2wd
9dLYBAtZZYWJaRC9lZVXhMinQeSedwvVLMeTQ2VugP3AjmNLDJwzGvocWrDRA/AU
mRC3c/8jIGiRycaNpo79LaTVq4VTeS60tr7N1852FofLd6pShEpzkJnAz83PP+6g
2DSrMTil617XEcn1hb2sEet6NTpqS4qIfZgHyT0fTCww4Tt5Mo6IaMVEFesKiBmX
qXqtOWqsbtIQWEdyJ5/mBvBQ1xBG0yWRyqz3Jm3YEgBFlSlbXwFv0OKW2/TeL/+h
ZpnUv0MlNObVpTG/GZ6vNq32fHmb5bDGCgqn1MoWeP3GXTRG5zY3OG8q+q8r+QEe
go3o5Rtg1z0WZtTWz5MBfGSjdzvypfeul0DUZr5AiAyX5gFxzFHoAKFxJT0r05Zh
cRV8HWcFC02nbGGV7JpTRJxivBItgDsB/5o0ui67onKTPEpNPk+MoOb4l0LDW4gE
FMWWdF3cuOKWwkyhzfIIEVXmRLSR0E63dAUnQaW1mH+PzU5vX75S7l6GQH3Uaqzb
TqAfbKSZtEFHfV3+BKYPWDazZmfGIjKl2XtcZd8mlsVL6KCXGK1G1V2QC7yH3r9W
er4pBR5BdeNAHDgieXzIzZK8xoNEafpcB++9+QYr5tiI3eOH+sufa+kPPx55J1HK
T2sjLFgKnp49tBhXAsKoQerN1CyNdLPxYVLLNBY4yhaWYyuabPu39UpIdorTQOii
RguEu+6k8ft10eXEIiTDHRFPKWzsHa4+iw/R5H2cpUdaYotaKLcrakqVr/KVec29
uUeP6f0PiJo/76SvZa4otcFWB/E2SYim7xna9VWX1vIyJ31+xG/TJ62p2+49dOq9
KK99wYJXx+AICxwHH2d9Ye/h0UDuTixQsJVi5AU5fLdKlkuD8tndZLmN/OsRmqc0
X+yKgEQjZnaSIRs3Gpmli0e/5NXmYG1OCZeRc+xG0PRzov4iQEJhXldY1UtdlaZt
huJevNQfstB/Of3rBv50IONp0WCDA48ABSwBGR0Hn7ab0FTXiepAm5p6cPQ5d53w
GFlaDfy/Ba90ANTh3nKQS8QM5jOkUHcVS/uTA1pBvqlkWjC74QuPxbQKj3iU0aG3
D/l1o2GGdnW+kr1KGTin2xg8gBZYUFLfLYCfmZANiDCmUtOGlLgCzq/y1zQZwXqE
jLFi96Ckij0sG5fXXdb97emVgARb4RUMHfxU5gUxgiiV3u47Mu3Cfur4nfhjVCeD
yvaAzezQEcKc1w4A6RgjrBXwOk9sqWL8eTDAu+mm0kgeJuyHLd84sZnWb35W5C+3
guTyrkZOgKzfa76DoeuPsbcFt0nDbuz5qiYtvk9S6VAQiYgzNfnC2mVMMRC3sSNG
g82R9utZgzTC1sBpNho4uXvbrdg1LDNKF/ANJtWJrA1nNE+0JTzkXPgHrLJIfC7p
5aH+MPG2yeyElVyyd7T+FflYC0MVHBchvmXNWl+Cs+Jh4ChjsorkvwE+ujlN8J39
M40xT9esWIus8/0ZD3C7HTAQDIBVDjuAK/R8g0HXDbDZrsp9UzOru8PcB1pOzOZl
5e21rsFTGAxtgp0fzbjAHN8w+aA9GO74wzB+X1C/ILfqh7ckHUcJj5SyJAJYcjv7
DE6bSqqBdIVf5nZuUE4HUpzqUMyjEjDZbVJZhH7ri+LQIrktaTEQOZeeBG6pIaDB
4qSimfo+2NVaZzFE3Jz9LmDnKojxolTCkVa1PVfwwzqbb9J+y6735vG8Ob6OrB3N
lUJTnHGcFnhi+sgLuIu1ao7xFZ4+ZzZY5ScNxwg/jcNvux47cYjEjhLNfGJVyMwg
QpDhKruFhiSO+ksT6zs3s/f1ZSRVcWfiTss0S7s2NDS5qTHDT9DwfI/Y1nHhZ0k6
54rqwqzsmCJRvi2A5J6SpzlIMrjOmZq6g7Qlc1LtrR3H+IEVHOkTyiJzyERA03c+
UiAJCkFc/lT/2RuJnHUpRhbvO84ySlBdR2BG7acgvzFoKI/9oZFDw3DYGW/Bsf0m
Vuu5/AF1S2YrXATMpP3hyg+5JXu1dhlRlmHgcVPX1XLGDxSO874WmFlx3EjDm2pK
qgQMz5dYW1thaMw90/t7ipJ39Xupj25I78arm8WAcGqjTAOdkcQrS6u9rqR6BhOc
yUKCSePVAgBx31WECEhXMwko72GwoBNMQkpTsTDWyhsiXeO5Jhzw3g0G+3aZZOKF
QRoJwsxjrj5mXJ6M7lxQwMnpTCPwekw8pCn5OtW5UbUhzWOaEnK5FTBkjWcy2xVp
3XP4YZL94IzViP84GaS+9Ph5TP87eCzjEZd8rL2Rn5CGacfirxYJsJddjR2aegnQ
yIgGTeTPxtAX2UKzMstMscTH0VoDr7HEgb6vpIBacJxQz5/GHBNNRTpgGlRokpVp
hO/9VFBxpDd/Y3yroZ0MSRt7F8Ph2eLXNkkHoIM6SAyWrhgWoYoAk/jl1liyieHy
+Xl8iZy8QjQPTFiBoAmE6KOk0kYaDYwOQgLXX0xwVO8y8LMWLH/2w/OGXq37DCsi
CmeNSVeQ8xQiMnWJUKCWAH3Xu0MGB7s7VpoaMnp9HPBrlH/iVsGKvk2P2sYkPGIh
hZUuaL9NlD4nT2q5UHU8osWzbLMoRwl+PhDx3SkMsk0wGKf8fMfb2PHXOCfxZbnd
wgG5gh2iz0Z/itwMm3EEyXXNDxH3isx00qZMMgUQaiihjs797KVfv9HBYKVPUjbO
Sil0jPBYKuO/o4BEhCF0jM2cxFm9jrAoqnVnTpsaIoZtlT39zfN+RQDTB6FaxUKE
3rsSwgdMnve+ix0/7RWF19MsDtUYKtqHqtToC89OBR7tnMG8+RCyVJhTP0PVAxR3
APPcyVM8NDak4nbdHSsbDUUTcf8MFDlyU/ZYVgVWJpSrO623BTcz34YXslIJXE1T
m1Aas5uPykNXOuBvNB7EhDhEXimKu2qzB3Qld8NSYBhNGMNMK+hBTfHOIWPfwwB5
tiI1ovTH324vEef5FuSyRyeRygQc0aEYGjpTZ45BvHUTJvAo7pRfeeSzVh/OYE9j
wgA1eH6PWpVPOKdUjvzeQOQoJWwPk8mfHQh/BXf8vWKOYs0jsBQyo2hJwDw8/Ugc
aqUf7KPDZ0DqXwaXEC929v9nClvmOBglRnOWbIHFge93NRY+4f7ZxKeNyjVdE5iu
ktU0X57ZYv1Ide5YnyZvELjt2Kpso45tlYZm+Da1gv5oh84YjSNjEHjmAux5gwQi
9eYN6IurYF1QvrD3DGE3qcNjVHft6ajBANZdkS260tcBxyZ/NdXeQlLvZDmtbokR
0Fo+EkzmsqMt5l3uxCBROYownqxrGUpaXP2Efnb01t410Q3wh61Xg9lVyCvQwCNK
61HBazCvO+aJ2nzHaKa5ASoWbLFxewxWELvj2An5UeXyBdxrisKG5egZMa698+EX
jagcHkEcebS014AlqLSO+inIxwHun9ZWArHfWZp7re3DUhpfSsPhhYeftJI4RR3L
N+NKoBg4xylwxR+RSoQKIRnaLTCt3JYA7jBlNIq8wmD5GDC9p8K6jPhiuLATAnqb
nZvM128GdiE0YHDy5fnfLiAauN4cTuwIktIKUJl37HuHiAxh0Roa2PpuNV5UatnS
2TgnHtE3RCQq1dxACA/Yt47hOt8xiH8FF9S9NtY2nDIGPIqpPhCk04tnkGmaTZjt
jqrRYCq6tcsVB7JJzorYrKmsPd8KCVEzjc05/yF43Q1FT7zpGtS5gyWblE+vfqTe
+SsV3JAv2i46F+zzvVPTkOZmDFASmi9ySw8lrZKRVvElHAy1+xkX+tf/X/pS8sNQ
eHEMPt31UoBtaa8IZK689PQ1irvEbVQphwf6Tdu+hcLI+QRvFB5ErD1nDhHzvBDL
wjZtJ2M0eTIfWHcyJuyc0ykBgriiR7beLjHZZbkGFb+SwqLVfHd+oPfC6nGnN2/5
CJxBIsavkpVDcmGei9XibksMe6EoNpWsW/gwNsL0j99wzMRhdRM3zId/HjWIiY9C
Ts1MyI/KZ+NOMiqvZL4JArk8HvunDGuwGcHYWcLRZ1lLEnSM6TJOJcSH25/6pRS4
RVhP9vCOUAB1eoBbjYuMkIk5uYs8JbRh/MyUmJ6ektdqNMs8I7OELQdKDbOg5pwQ
qAnHypieI718yjwsGJm1uzKjwVV6k1Ti7XS/yZ6aTJsrSWyag4FcQW7ADq8ptWMu
Zmuh2ONTX9Tm/hfa1OX0iTBXGWf8pFTx/achzeD9yzZtnVDcRU4hXTNl6vOT2TLR
8Q7HWSzBMRKsDkqJz6gOmKjFqLGNLL6/0cGnZok1VFKs6fT3LPtWQ9wHcX2f3oT4
g6w+i4iMDKkxjZ8NRkXvGuoYHk+Ci5YA8WeVSQQTsnxPd8ACOcmVnC6Cs2y/nURt
/4SxPabgwWncvpMDmoZE1DJHNwXig1kDtMuQN4qbwNjuF9WjBQeYykQavaIDKOXr
ikZkKstIUFDCqXfahQJg/j/85ZMlCQucKciRhmfXdHGFqZ34pbZ7tQ7I7QH0QuHi
VRxlFdUmyH1SwUrXAI/nCSSTNxm9fR/kshkCAItTr6fI0+8CS2IP96PSVrqFsHau
BpJyvaE4PiN1MUqE7UcygBxEkQOTYTU0gJLVqPJWYca8V6HUVHUpq3zJsj3Bi/os
fY/+PTlyDkxSbDVcbnQqM56HIQell6crwdvfn+W1ibNDIc76fOEfSMR9o+TDrTw4
FkP59pGrXnnJSqLIidlhwXusem00YsXEy+XFerQUwaTHPTVRBWaC0RucUlTyjfx9
/UwuRsbLdh/57nqxz6HwnkrUK4q6ddi7B2GUhUUsvEqwTAaPowUwhSH8j9pNc5Jn
3uw7+MmnrHCrkLwu3npGp8hh/8kpoMv0JNeIRus5AE/id2I7RdPAh2VUHSUFSRX6
Sbfd0cR3ceiFm4R3Yzqie3xEoImLrBOaY/nSSSWZXerbXE2mdqngL6eBmC9a78WC
dfSyfKM6jM4Bn027Uwqb2qWEGr7qzj2YubaxQ6qc3/nLhf9GPDeXRlqr8OI9PCVO
y9WVA9P/WibdVo1/HkymaPt8XJdTySkrGDWmtYhcW2oT3rYBRpOFMDpq4Xbqt5te
/vGkM7XDxC0DgF4FrVW1OB/zBECbYeDBE65ESLTuF6xZujVXOEUJDHhT6id2xRwP
yVTdaBpnsGidl2VHm0f/s5m5kgDWFpU7ZJFsRnjh8v+2ifP1erLYmEdhsjsPTab8
3Cxuk1trG/Z0/KIHr4CSZUFHuwKXBRQpGYWvoXTCVxdrPybc6/A9G7EFlkwlFjNb
4ZvBw8pn3r+qwb35c+3KplKHNWmymsb4utvZmkPcOrtvYY9m+sqZjYXgAwYnOUyr
vwCVg1C578fNqFU7eBl4CbgM/yyegiHLSU1yrLCnmjoLwCu+tQ6xpMZDt8dL81IX
JGgsNVP11UoeN3n/sSXay7CFgZ+J4V7wjXp5LHynWW2HgMlyZsWOZPfUK9973h3n
eni1vjOIZ0wgm2jafzko1Q9G9yV9MalCBVEtlOJO4S3qZwpBMlxNGgJUO4MSx41B
5ePRmQBjqxUiKyB+4AY1eIDFMC8YXgbbpqv+eiuHx+E4eLryNHOz5y0GVf+eLHTN
wbj87uGLZ3KarzsHEUpz9uurKxv+qHGg/5/JmiizUnn9BtTZIrOU1uu9p8Cua+ew
W5Vs+tuF2akj5lM+EF7Gx6rEQrRhQ1I/cErOCN4oM/brs7UKHfj1joCXw4rLvzwy
X+5k7XIKXPzsyYloJ0bRS0t1Px6nHBotljOAPrWu/Zdyd/7qJvYi850RpO5mED6C
Kut2CBdYu0N1TJ/Z6mqb110rkNi3hJKQOUpU72JlR7FT/XIrMEjh3myJciy+MXJ1
rNSFFSebFaj9Vu/s8+f1YJPrTf8YfvnlD/Z/BcqmtYdeBfrC09fTsh08EBs3y7vc
+3uWn20TZaS1/niu5Yd6Cj9QSMJOcHJnyQi9QAoHKjNH697ffVXwqns59hUrggXa
dAg4XYkl7TBzjpITdUbWU2RHlSJEuDPdNMMS3W8dGGWEJlgMhOLkP2IcvdF9b1iU
EuF5SQdR5ZfQPpqB71Bq4G2pYvuNpq26Gh+B8M+OP4DIk4G7JoJucmDBiG5XFgd9
EPZwwxem5Pii+M/xXcAtmoDquy1Soha0HSWVz90UR507BjmC9zBSRgVxyDLanJmO
5KjONGCoO3Li0XdjTmWVwoeZ/1GQT3LZk06GAqi5ycR6Zt1/tdxUdH4W4z8aZdKT
5kCrg2+pEScV8Yy02iECty2vkDviOTcQb4IOgzslXixPnKgLELrRrE7DVykBzUyB
IduXQJc4swDr5ibRxDZNvelZrD8A61p3S4BDi7pAi5+7NEYDw8cEdXTIfCzOe1jP
2W6j4IBXLDql9Q34pS1CdctDb0s4iUX6SvmrUrvOAo6MZXETOpqMsfvrG1Yk7dlX
SlldbgorxXdbAEYSKFp1xF4MtWr0+QI3JVqS15cJys5mdRx7DIerB+r78hfJt+Je
gd4/WnqNxjcXohkjvwYJifxysMdoXAvfAc6S9fdMm0qTVdTeVf65cskuTRJrLqGV
f2Zwgk4LTreqtoyJpoSQz/OTSL5iHcnYsJO6MGCEwiNhvxJ9laL8taB553fa3Ury
S3FS/+4j7AnFrPLx0uOg1N/sMOO2LyPniE6TCsAQ75bpv45DjlB33elFnvcwbxR/
zf2skWVO+7oQsDq84g+RewDMTOFZ4olhoKU1pbaeiXKPPihI/fb5eN566q8ecDRy
IBz8YWc2PIIu+TWzjzeaDZGdmhl+4ZCjyC0MAPl+YQ/PYSiE9oL1f7SPCGHVW4tv
wX3JTIEvj7HKdkdETwNjiF+Aqi8R5XX++ZhFXh0OYvseO096eAsYCIJa12sGy2es
2DtLdKOW9jGbt0vniHIG4UShQdw1UdelgqNjk8fTGdgxv2JB4dRMLbdMpYnRs/sB
5TzPnDRW9n3fTLx9jYcngaZ0Ble1muJk1WBhDT2feMrH3YflF1sySgbrb5pDo1rS
KBfQP4rz6gHFx+MAd7N76kGzTyHcJOqv87RLrecL2GW+c9qaWsNEs6efbMnDxcAP
1Y5ws8QSu1NG0GHBOBfQHRyXK9d1FvuOf+4iJq3iircSMCKUpRCqz94olbg9Hudj
hArCDL+eNejaGazwZ7eAVD9MT/HuIzw49zj2/EHfmJraGdOowZ3YQggj3Z734/6d
ZAEYGdUyHdD2D6g7f6F+lPGWxL4PM6AVwjC6sX+dkXvpJSRLRSqu2RircxxWPqsc
FWNEtDCHIpWNaK9KLrRhjq5Ci7dJG+JYllFp+8wYt4kihy9TLqJCELbdk1Z0InMW
UiI0aifhxLcy/gBgY7YvJR/AkiMwbZMCByo+SlWawxY+GGRQVp2T9iINrQU9Jp8Y
mJkTys2yCYuafPiTwCMgyQ/ndIwqMyGdMYXekAMUzdP+1sTG93i3LzdCYdI353sf
J3Q1iXR8LrQqJL0HIQJKrS4LLwBmp7D9+3GQ41+fNcCS2BfzRnGZdtBumxfaz0e1
UZhRia1A9JcDLq3zXl/zmcor0UaRvUHbnemKzFDwjk6K83ZnhwaVpXbauxd6PQx1
tWmsMP2YrjLoxFMywCr0bgSN+WV6+wq5po+bJm6WIWdKa/vTG70Y3zAZRRDnPScO
p1joo2jF+gGgf9w88N2S6oGlbFUs+Z4cNpzkAVF5L/3KqeZef8bmTxAGyNFrO3TR
nXOURwy9wUF97M9O9YHC516ec88g+D06q2HFkdtP36xHgnuEhVWDguM0uu5yMI/m
1ZiE7DhuS2FdENhpnD5FUukiQUBBwwa2FCt5fUhZ1IvqGli1u0UqlMRTe5oWljW8
/1LsgUN83Icq/cuRqlWUMwkiQXEIJyhSYKkq3UVjk7ZvqHMCBa7EafVNwXISyPJg
kTb8gYAIfcfB3vjpCizKAvQ5nt6mQwe7s9YUEwbC0Zku88vuQrzfgsUIeIwmqQxM
W3Z1J7KlhTdVHNciEj/SowrVgdFWlVSRZbMCRBbX+ys+dTNKN4I2qeprvyvAfQB1
WcNhew1LWxsS3SO9u6LzHkTI/47U0cC+UTzUWKzQB/fJTfDigem4CRUN7zy9EJrU
55ggdlEDc19mgvlzqOuK23+WBpS/kRHECNGdcQL2GQDYsFfgh1IUUET8TaQ3r4oL
cSObquwSk187LJSIZQ/Wb0Us/pLbpRjW8ON5BKDXxAOfegxejdtvwwrGms2APQQA
XebDH5bOouroEmZqblqIJLOIsHHvcmYLfmnZ8SOeBEeD7lWFBR/WTBslUFErJWFE
iD0wIEF0n1v4u0kgSTsdREAd+WpbEZSEWzgpSbZ0TFROz7YKvE/4rHWob9BwmekS
Lfts0uAyCcGMMeABpgEtXz9l2CjRF0GA0wb7qZjgg28xYY24JFs3B0r9JhNWfC+h
Rv7reN1UniFdyUuH92ZcBcF8S4XCb+UluHVDA4nGdb783L/Zlwjh2KO3vnSRDrD5
Ux2YsqGSBMg7zIs0XWwMEtZfkYv89l8fR9C6ddEK5m+i8KV3t2LMinJu4CkoUnJG
4QfwbhF6xUar7vw/WVcxpHGhDADZ/E/84LP/D4uDitCYnXqJLeOgtFewEP8T88ft
9Ax9WNUYm0JBxERhLhl9s8a6imWd9dhDI+rPl1Kz9VxrdYADXa0BC2Mh13vZmkce
SGdIo2wnB5A78LeH5/UQscIJ7wIas/hpEfS4/grxF1yEXZGFJPMHfRuf4A7CIsIi
48elijQrtkQcqghv6dC+i9yQIi0gLF+FgFGmaCrcjEHRP9dL29f6JEOE3Zq5bXUo
/5z9M+3r65q5pE40ucJleIrTcX9cFy3y0wBLEqg4w4qgVhAHND52cttkM9SWSs4E
sNe9TC/Seaoz+p/RuhPk0S+d6l8bKGIw9GV0ytmMocvAqCbQIAaM+SRi688/zNxo
/w1LkXjVxscEZ8j74wgsoLtws5Wg2CQyyOW/2pyZMKEf+YtON7twJ65X0OpWRjXe
hWB/UXl00OaXm7HMjdCXGHMWJv0GSQxkd0pHPnMSeoFZb1qYRIZ9MItMF8ZfJ8mc
1ykSlXXF0r8dzab2Uk/rQqgwCwiqW/4nfNIyLAGgbG8U7jPAiD6JLYyfKzOhrDYu
m0jxXzEW6o0L/YnTswpTFm+I8xu2o+wOg89e5Ta8AbafDz2o6Q5FPbvc2vi9wMjF
+UgblZ0Hxb1onHcWg+lcLWQeFI2s7uok1jrQawn1M0XBxvJJv5zzU4Pql5LBHR/Y
8UDWBx0ngftAZ/ONCF6gj5mYceTFMmvxzaE65viwzEtK3ROo7kIaYAlD19VJZBgI
8qrrQJM3eT3kNSPcefrB9S4sjH6CCL3+dFOUPg8cdclUkQgRL8TWmGXZYDU8t1cl
eDVeXsBW0B8zMvHTz4j2thm+dfRhbf1EpA61x5kmpcvTALx/44PLaue7fhN4cl7M
WV8qI+JF9/XnoC3TDHBzWsLG/Uzbx6no+JnND4ioCaZDnQUDArYoB4BuCyQ5Rtt7
z/ElcrmIEEyZJcY6+Exlarkci0YQAGP6miUc8NlvkaNr2HP3UVfX1ZlP3RzCX40t
gR4t55GG1ISB7kEo1953OoC8FM54dxvqFfWFBiWsVb/GpnSmK0QrQYJ9Il6tycyl
9Q7T1b4f1ibnfVihhfJLCXfoXZW2uLdWaiK34xPTDNmFpWAMuojF14jX9LlBkiMb
8spaoF5mmMIqKPqU92+t0ZGraoNgGwVbelLlhCfxMrCRiSSP8ldoB2LQvXwVZWs3
ZvmXJLPUKaQYQA+IyRFNDqmEphjAcTltSvC89uzzYGLQRsUTBGcrtWf61xUal0BZ
8RFT0C7AqqALHdWfq3EWF9uGw9BJEeM+LCABiUqKBMgJRWvk+83LYWo5NThAVqUM
QVN+Us27HBf31bP1Epoj0XXKNnWm8hoYjgbgiQHQRUupX9FS3EkkOgrLj+xqwocQ
juOUQuj35jGn0d3frG45pXoGf4XL//uG5KetZEJL0Km+aLr8QcqmT2mSYQTH3JkR
ZNYZbs5qQFPgxE5TZ8QI93jcvP7gWU5SRkaUU8pO8i7nGwTuMXAOl/QY1DCeYtJD
jR2GtIv3FG5Oi3W9zQv/4bclMD2Ku4Qs9gJ7DCmHU9cUs1K3V6PEOaGkowcTqci8
+RsUd5rVhj8kt9D9J/KVzgM8vmhBxZrpIfiHeevDPCbJGzBkaq1+QTXmiTDgRR0s
eb4W7lr+a7X+wtsvekxzcyXcWdzV1cXgyDch2ogI1a0j8TK18ATf1doJY7esgjpi
KsMcB4xT6Nr9HR5X671vZ5FECTt5VtrJPYGrY3AnGi7QsxCdk/c9f0cYdrKPwxYB
uCGsN4CfEP3/munCV3GHknliyR/91H0gRsRi9oLwjyVbyVZIH1ajSTKUHOrDIMol
7l1iPaViduZOG8WZo6UAqYPjYfeOfdwijJrFGtFZEBK59ZbGsVB4+nQXt2BOJp9q
hYJm47zh83uGN/i933VaqwcCaBG2Ay8coRc9/VNqZSEhHWUoe21FrL2BvwcxWkVv
2Fwqy+ZBrAY48cD5g7CUOp1/3746EACZAPQQj7+QP/3m7xiyrkhuPiUzyevTxSGi
E0RK+X2oOR9VUD7o099+ofMjYKc+y8kUT3i1RZ6CWE/GSCcpiFtcfoPpiZnFJECy
tAAS9k3K39XUFsN0d8h1if4lwBnZ1sb9fUK0gpQCEmdAgsI9S3kXQ5hRvghFokvO
22tg3xJd45kupUf9Lrba+NpcvVOpFvISb7DjbVDhTwTO4rhMw/LcrSi85vMjYxLP
4voCtOZkJRj8aiaeSrIF84S2Th6DlH6ZUm3AEMGP6FnTe0+NZtW8AMLDDKYQgDYc
Um27vcSB74FkUY7sTGT9r5L+zJSzZJv9tD7sJa5ucnSlBPDHQ2LAEeI7AfxfRpzz
HHKUsMAVIRxNmvOvefrwRvgBetrZMpqplo7/3Faw+G81mZTRS3XSiIFNRcGAEFrF
VbR1asezPWOGMv3U8ochstiAoJpigxlaZ6a2TQcZLbjewa2Gs+N+zYs7MR3Hzbgo
aIVouY0Wl7LEA+gA7x3iLsCoHmleQgDWAGF1NE7JzSULHRISkjvuJ/QM8TmmTSP9
2Vs+8WddrdDK3JtA2P+qxfl6gCrjGzi7A1iH/ZlpnQCeMovgPOvLEjAesB1vRGpa
apjNfwd5V3Q808GzibycMJAgpwsPEhUp2crv/kNBei207meMj2eSU2eBjwfkS+lE
rGuIbCgZvdKSCTl8gqIo/7bVBGRlGjYuEAThGk4P/6Kou715o3pWwSi38pV18IKt
jkquLQ9HIRZaGoxgWzahbYwZ6jdSiYwIobqC/Mal/XAMQHi4Oz+sPQncn+hKag2v
2nNLEuF5hhkWPdIe0I/lHoyyUzxr9BrD158BXVjAe3Nh8a4WfDhR3bCt9nbINDWo
rkJJXW6uw5b16CBPi+LYnfBY2ctEscym13t3cwoLr0DZxazAPu/OJl5MBTPbaPK2
p5U/BTbMw3nJvso6rou1XTQuoqt597vIPg4R/pZSzL+2iEIJpZSGToamaqPrxG4K
iI+e3QjHzB0BhS//SGVE0hrlrM4YSMymYMLOH6IZ4R6l6b2yzRQtH9Jg5cZVHErm
A3lFycZdcr2aCDtg/C8/+pEM+ala2tkeIfNllGPeWyNaJbJKGgallUBmmpysRhp6
aOQUmm2o9iI79SGK2dZvukVMRvxt/2J1e3aRWexPvm6nzPTChpoMLodaJQ1eYgoE
ztzLV8RcoMd52o0y26TAJiR9yqV7R4xAOhY1d+aqrFC75ue6cBy94a5rxBVcC4JK
DsT5bzONOVzMK4ho0IANHlRyN6OSAJLGsO9dQxFPDAAZei8/m0iT0epjh7omd7Oj
EVPXciGZmobxoAQKSsL4IDqhd18YWKBOjyc3YXndI94qjwlxjJjD6vaHp8bI9DO1
jQCsslj2p0GYp2AAAMEgzbk/zwqgSE7sCfM4B0hgyatR7pXaDtuLNXu8st5i6AJP
jH93h11QxppUpcT2mt4kSZmugF1fnpkvwQG63HdJ+stl6VoMtEfVO/IzYB6WeXUw
RAar98wJLKRlFdVKSfB/ocXe8BhcSadY65lpxu6a8h3gKwZ+1LGjFzFxP/4fR9WQ
EDomlGzLvgcP3cb7ujGT4QVtNOymwknh7Xy/cxMKhGepmZNWOsCge5tFzJg52taa
si4I7yXFDQ89OgTEP682qGM/uCcaISI4fLcFdRtp1nIyulQfLKqvd2bAhQokXU6m
5LUldTUUNbT3xAAUjZ/Qjb5ycMOadCYDfnD9Rgsr5rb3cGjy3FqI9y9uxRKpvG2Q
co3QL+JolNAl+cG7HLk2ouvAndt2koERAEr+XCcqh6Aw+vkbkMlkBAJbR1INS8SF
WOXaC61vzz9FWT+f3fGl3x/gSoJ8dJxLnA7bkQy+4F+L7c0pmz3bC1aJJuBmLRJB
IA+hsXCiO4WJX2MH6QNa97laPpiF2TiTvXFoyB2kA8qfJBSYCEb0FXKeuuZ5j8n9
PyXADk0mLMz78Ov2b6S+qfsqTqj//I++7fAy/XI792QhgFhiZzk6ewB/wp8PKlVn
6YFiWyViO6pz+z240eSJ++0i3DwwOEIBl5BYiV3wzRlMvteg0MyDzV9BRTYUkFh2
vOA9Mcgc1MeEWakjbZCaB9eXi2na4rVpB9VlgxoZxRGkNBM1QsFYLlR906MYAM+8
rQ/mr3hJ5OON7EzdBAmWKVGp6aM8W3GySJRbKf7XbGizfC6y2Egt0Nqf2JMBoAgz
oocdGszQCDdqCiPa/3OB/KBmsIFs5geuVvAioNdQ1iIm5CP3UjAoBiKA5Pax6XJN
b99op3i+UjbR92CCwVx1wS7mektNpw4u/Z8eU/BvfDwd1+fnPSDeJK9qboG1Yi9P
8GTivDHXsgHf8Ed9ckzyj6b4L4cKlHscEfCcalTh+v/GSUJdcEqYVM3pEFaPtPpn
ibqJnVfAtEwJk8nY492jZt2zDrQetrZKD7OsTY6DwqNRuD369+vdSqofBg0rLE8g
uByfTuWcQKtbQy21R9/Ulgbu9ElbBnnAV4/h28R3VMBexz7Yvtw4TZiYhu5tZUuK
qTjqhFjYeMVwVXf7pRvEMdODqmX7WWEmkt1u9MBbHOUNAkBNWbmBY2AQlQR9CXuY
ltDm4tLJ3AyWsZA/weVzcLkTHAzqSmTFHgNleQ8XAr6Yjrmnq6aWvpqE/wlx4EtX
9QmxrEWC9+avN5OcH4Ij8Yq0lzEvwzvxFT92GBfWzW4iUB8SKjik7uSGVvZJA/lI
VSJeijnlJo3sZwA3fYqqBW8UvB/dZDBBQTyJz3OJ8lmZ6sPv4oE4AKMqAbedIfQu
yUDGMY9pEhcZpchRCAqH5BzmVb34BEwXtvhrXr8x6bSebOC0NWQOvQYFJA2dYvKS
P/khJgLyTEdz0SGn8viXZvocyKmMNG7a4aiqOgFDqrPA7RgRd5nqyL8T3qSKWgNp
JEgTpEDIqdj4bz/psr5b1uO3QbJ3kEaM6cMegp//yXI6ccn7k2L7UqQeGSHxGUrb
SL6b8ppHj6XyhQQ2RiJFeTuYCU+NzDOecFqKAGTlaL3vhs0M3Rg0YU/QM+gybSlD
BZaso0uHa6NI5sRAZvSX8tN993v/gfQh6z/QK5Zk24WK86RjmJ1FDTp1SOEtlebI
i8f8O27CMJACrEfqGhplQse/rwv0eQtl6LEHjYUfu434DZ5I19/jUTayglAYo+Z0
LjAQulHJnWib9NGJxA13bC3Fkn/rDsSAqssNrJt9WTrzhPwXciehlyBtd3oLy8qA
QL+PAe4yqXCRyMpGrer+XwDpUjzToLXvggfTht0qgK3RmO/eCO7tvVYv+ouXCWUo
SvO0qE1TZo7dBl0o7W6vR3RU5zuL/22N5FD0XdVmcfgVbfDKwjR4Ms6qTlduEmvV
wcHtz/hZInAxTLsFKRO55jRy0WGFUjFFng3R3BDhy0XPvlCL7gk/3kMqWs/PClP5
Tc1Q2h5bAFW5zxV/WKaB4+ONWogixdOmGHLrwYGybW8aoLlPz6poh0ACtG4hx+h2
R6MyIz0Vddc+puDTJot2CyR6OHP9hd/tckhbFIyvvxm6gI3n5bTeI39ejuqAIOdg
7IPAHg7VysamRFVDQy4JExsJTzTuTw3qpUajusaUEBYnx6MWavrgspWNJ7UubtYv
IkEU48BrfgvCrq0Cr3qeU0yDpk4iELOZqTvlJF/zVZ5I/550qhc+7L3W/mKs2ijp
tZgj32XDKrB4qhlMLWcsEUmdLPpa8PF2saxNxrggwxbW6DyYqtyrQj9Z0k4qY5TQ
MvdVl7awbr6ofsuojt1IiNXNnCW5i7z3IbljWEhqCMRenUHj+ih6CEJ7H4NX84fe
SK8qZRBGGaygL/AWmvyORpXPab7YCgUZpi5jNn3PCrjY7Akg7JRXM4oLVb1gSRXy
QN++dX7xMR7el30+LyunjO0DHwOv8Oo2OdoZlF4yKR0w8fcyFHPXOwIrA3x1Jnt8
TKEyT1Kz9eHwP4YSe3uiMyR9s2RnTk08DAusj2M6cAsJ8yu1QgCPVtdbCs/faAAd
vYIb2W3x+cRVLtQcAsqveGyYB2Ce90WVJAor8y3SMpr9pPGouy4DM5Zx1KMR2Edf
u9yZCUjp5jdJv5MSeCqndDomhIMKpvp/XL73WNqHIEpSIuMrBhXX05pAx3MbQ2hg
5tcOHB4tYWnKcV98659i8kq2wzGatYPi7wpwweMsvfQbdzeEmBv98gCWTXKO28lW
UKDrL/AaQxVMvtQi4gpzdei4PEp/CYxxnAEM5U4t/VAiq1q7CZgiXelqURUznxmZ
x4EvZxmEiUbFHR+PcRiEg4fKta7ut0LaAtqM3rLEuPMnyHQ86/QUyBpzMvW3K5ao
vze51nAjUgJlnRM27PfgLyAmYidbs6McwMTCCc+bTSeQETwRChLGqEaLZBMM9gup
1F/uePdWGprZomLTcdJIE2+PQ5KFZ+QcLPUnhRApvUBjR6SfNmb/5VD9DYMU9iSk
NKqSP+lQHfXVeLDvznL3DNGRO2gptmJ8AH3ddLLto16MLttvkHff/hQCWOXCiEq+
agBzFFJ2ttj8Y8rW+t33IQE46NgNilTPkfDJMSKl0muS1cSv/OdGMG2PMeUr8i1B
A7yE+/bcInW2ytAOz9xvBy1p0Gmlnvx4JzZq4Pxf+D4vGA+POcajLdHlzM3dwCrd
I5NNbt6KmWfkUyVSuloafSvOWeas+RSojPsH1kk8yCkCVZi8Eaz9cDoAbrbdhXSx
LMOrEYGZOW8zRAKJhENi/58sPzetz0GBEvxyKxoN5H7RisvOgbaDjaXJJTrl8EVs
gSVaviqZZRTUcq8J5kTJ/3PLwCpogWZL7kGqB1U2i/Yv14vC/dr/iehuqUgvhW+U
TFYYltH02LCd0/o8ybFnxZVVahAhFhG1LDPVX4XrxHztLXEeN3LBAsZ1z9EOtLS6
yEEK0T6ycz/v9oCljZCpsOeHYYBnW+BeIpzdvNTlH5mab2NGq3kWv29Q30VmY2YU
SHe1G6AiKIcPr0uBBendZNMYt0MTcLZlsq/6zFtcVrwDdjPnGv0c/klx86xDcdQ7
r8iEzhsN8FWQ62/jjHdjTER1hLqIvw3hd/7VKQYQTa+V4yv+4fjHnvgIz6CxawQi
psc1i4LGvpJT96woIZkI2gpV9rKJtJyaMJsVB+hsM2XCnSuMo5idbfgZG7Lv9U5o
TzgJOeqTmAcRX6lWVwz2vaszfo3Dn/p1au1aMKJPKl1YQnUIILjqrUy6GoxcM40R
o2p8BhON0a9H+RlI3Xzeh5p43E/e0+t0FbpHFKKB8LLaBV8tRK74vD80+5s1pUSv
KgJNdLsCAi1e8CRPeMAlDkJhWyftH2W255dGgwOCCCEM4sOV1csgy+vjGI7i2OTe
qPMpriQvGRL/cNWeqxi6d9GsPM3ZfVUbfw0yoR7wegtQfXEzBNuOZfIwtzHU2GiK
7P2l+s2EyfKadpuVk7OmRbFqUoQq68fndLtsgTf/gm1y6g+/sBnHQD5xiq0KzMRu
c0gQIF8wHFiaUai1e+N8cWWvInLfZDhl1ElECUG1F65TVOzF1lAYHB9pKD99WUWp
Hhprm4tqGJtgWaRMMj1uXQixy7GgRGRdN/2EOExmf3BF+8wmY3xN/+tk/wb5iyQw
DNFCulQvdQDYzMgQT58uIv0P/VQz0moAurquQsEcUwMbh1/AobK8zS9oZaIPpq9S
DbF5zmjFiNnlLhc0F+TX/LRib7SAU5zm9Im+4h7um1GBt31rzk2Hw5l9Iimc9J6Q
A13q5wHqkHRgzhkFjlS7H8KYK92ekKA+mqiSUmUr1GvW3Q0pryp9knuskk5kVb4o
6qeM3Ga9+IPOe/tf1//wrXFX2lywPwAWsvVt4/ouqu2E5RLEn2H6p+5ZWfjoiaeA
wROrE8+4104tDLqOCCf4RWml3J0XEuf4z9+tVDv7UsHUtQYK4MB5tIKuEzwvOBLY
TMRPQpt3p/C27I2PDJ12yc2V3peJudBhh+odvHknjCwON0dwbVZky8gIVwWSw9Nq
1ifjAqAqz+wDIZCnBj/nGiqPMJ7iqq1KCH+8+ygXswL/DQbiNx5ppsJmpvj4c4xp
ngxZpjojcNweF8tX8uKwWzjaO0tYwUQnRoAUATFyDNYrM2lj3kTYNNsfQe0fAgMy
Ya1HrVOfeG4WX8qI6WWv8EEwz5/88+b1cSnF2Z+HRi1d2xWUWvorgnySfsc4BMeI
3rGAwVgQXAs98xj7krvwvYOxY3qdwPKhVpt77j45RtydVQR70cA4ToSRxfbasuef
Sa5TC0Ko0bJuJeTNNEvXX7Y7RAwxLGhHDmryKILzmOHl24HB/eH+IOTdDH4sQ3gr
qgY5+ohBWaY/SWNh69yq4eMa6e3CV14YfiSC+ufv39PhKrbccQ6wdB7wc4B1eYBw
aFax8c2ba0XHEKbIOhkZ/h3XoAr0gseaW/YSZrYMeX+BkPW0FpBiKabMiwNnkayL
zUjpzMyR8TAykRmROfKIo0X0niuFRElhwhXNfDG7rufgzRINz/OBb1QYwpZecyD9
Rg3HqwgkFJ5RDFTbV52f/UzrAfydU/LWzAo0x2wB2rvMMQYNDSDHLH0hDjnq+ksd
Uvip2EQbURRgQOpc5LDzIAoUj2Sh7a/0XQHSNYrtsCIvSvlMKW9JpHMjryLNo5ak
JWWyna4CY7QNJbGA1mW2709iMk/BRr1TT278Z3aK3gF5lGrpYJhe+0yK+auvQ7EV
EXWqocoGzXfV+iqB0LhDfXGR2ikTQAVWyb7nEPBG/dBQEn6LRYsXOinkM1C9M+6i
gOKq3QxzKYOLCWOvwg5EIyqf5H/NzJvtZb3EEDAiBDCAq0ZiXSCOsCmmBIfsjkER
r6T5om0LHF9Nl7y92d99jMI4oWEAQlBB+OL+qTV0UzCsKNBxQ8AM02ftKVKh123t
OGr43xfP8QaajCusnAoCrTh5UgSASRz8NPoa41KcJo8mVRMCBIAyCGWSCViN+gGb
nIWhr/9tiZyPbb7ejpkhVIq2V0vD/UXGmiyKoNL+/cjKs5zesMzbPaiMTgjeDPhC
f3LQ7yxD7WO20oQvbBRc6snnvy3Xox/LyETYVvWEnhs4IoZS/+iMfnsdy2wBBn7J
INp3lXs6D6PZ0Ry87Gu/vnmVbXWpE+mbxf9vSMsZ2JiXFJaxnmVTfhHs13hNrH7A
g87LI4EQ4XFsSfdJADbq/gJ8c47y8/T6qp2ncG3hDUOTJr9PQSleX3J1r8W6dw/L
YoZ3wWPItAIPEB8W67cLv3CYp936WPpJFHu10SJbS/6eJeY372Oah7t/LCV1l7ca
Q72RA+noNcCLHg/RpusIVjmv/czwp0T01fQj25Q9KIjlfyv/U8edQnruum661pIA
r8P88wYV6Yf/GG3zluArAriTunKBF7HjOO2oEn35cZ9kb+uykvCOXGt+Tgt+ujce
JRsql6LkpAQTRb8MlweESYNe6fTAOVEpEdyX7ZwUZVio3tgHfs/X6T3KOPY6DAuQ
0FO1FvKlW+SkLebWH+krQiB69G2sR5K5dZI9wkVuklvpgFBl4KvICSkylB3kqKNy
nmFBUqwKoQpsePTAMixd83Ecrb6L5w9wfPru3Mtcav6/ucvQPT3JOKgS7PPD2NEK
QjHjCp1cWBtudZLCLJQqa0Ln13DE3pIPeR1LtuVAh1RHuwfdV3ykQg8cKYjp8fP/
GrhcUhY6lC7GXxcSYuPiimWwvtrPfs3410wTfFfAoDs6ZzyzWrEZ6fGRvwh5H6Tp
SJaA9O6My3BcmIkV0jJfrQIeGafq2v7Qpjo0x1cIWJ3ZTx+QteYmSEkVr9AT7bnm
AJL14q1r1pOGKrhZa5M49+sB/slJLlhpvEvCmTbY8diiMoYLt16tMaclvxJAM+Mc
AAonRLEZsTVZeJyrne/UytFXx1GLn45v9oPnKXxyXjy9bHcMsta7r4tiex7UFWEu
TwM+jTizA8aT7Y2uBANUGTL//5KdQcAHeoQht5wplyON8h62+/yjiU7pLMzXHUrh
Yj72NPOyEM08Cv33QjWzGzfrl/Oe1GViI+4itFHIOybaa9IrKOxw0jg374bh3SM8
TAxkFP0fKDvRSaTxN2TstkpYXTl0hLfOiDvLDP8B0ZksCx7TXG5jkkVU5HJfG2dD
+jfCl7au6TdDMrGRVdoh1MBt7v94nFSv+pcZKHdtjvbUCGBoLrS9bkv2pczPd7Gd
OKiIMdtPjbWHc0ByMr6ijA1OF3S4rgMFDKl4fiRh2iDTJNhp/h+cxvPnKTuz2+wp
N5MjgtzrarkN0g0FtiNjJueGyTWLM8sN9wGmCS37IDDCBaEs5SrDB4PFZ6bvN2X1
XDcPFh6PxD5tXqLKO3Q272cb0MLzEKZr2oYBDu09q7AceE4sAArH7WpYIts2eQ50
guy7QAyzlR8gtnpx1qkdGqwXrTIQZZjR2xMKA7VOqobNzRPqAVIMDL3t89O6Vq8r
qLfuf5jwC5PzJf0p1xAW7kPYKR2uQ3Dk/lFcUk0eoRBAqZ0LHHyhLQnWtahfP0fn
Cdvb5ulAErfaR8IO6cfLFT6+EWbLlw3Sp2O6gREw73ka6rp3obnH6N8YbFQnTunv
d9hl22Lu72OFq/mYuWs7yBBfSSx1mn751evIKqemloZ1mBYmKaDqv0MIH4DN5AFH
IrUI7hfYbjDuOampmjIVodB5eOE4SW471ryiaUE/qQtK7XwigCyQ3fjwDG+92hgL
c48RuNHQn1tGkcUXB+Gdu0W0o4qx+UZz3KWpOHARLgYtWy584K4ar2VnM4dARsXe
NH/miwEMbdgGUMn9XeQPG243Vy2jGgPF7Tcx7crjDsosnwbsU7il5AQm1JatfLUS
cs/xWyRf7y/5/Y7kZJrBTA9TUiZD7cBioDNo2aeam9QSgZhOEI8WiBz2zfsaI6K0
hcuDgDyNVI699rb5Mytc19xBf5cBGIg2beWAa+C92SQ+/kjzVoymHHc7yGebmvxL
K2Pmompg4KVTsI8qwp/hVe/4jOjvE+pAFj7IUroRNs4RgVvMu7ro/kE8jSh+fSYR
Ewwp+iOrmEe+0HlDQpR6dVQrILwg1vvo6IQzhblwA37gDtZGCnHUKpQ923afcJby
vjsYhItikTxiuo8crQ5zApjAmUHiO10gMxjD+SCvr1WfYYKOcbySBb1MWudAn+zQ
5lvfpRsFntF6i6wRhrKqAe1Sycg6p7hfrq7eO+g1OMSbU8ak8F6pVcw1c0DKd/68
y358QwlwJYLL1JiLzSqdvEeSsqEqMKq0RkCC8bne9+5exSxOg5B5FkD9C2UXBy99
wWJ+uZ2N54bgWBtgNuJ7+ZkXBiKGJmoeawU4PfTRNFee3YOzWN3eOivc9SL/lVXI
t+2CPGFzMP8gDWgMuLxnsTgQGJvAf/2/goFWMngAckv56LQMNxlh7VFXmvmypZqC
D7WkummH2/9xYbExthxuzycPbKP+tPzHt3fQy6nmBGWCSsJAOfe+eX549mzI6Nky
DqWaEm3XcdpRZaugTPj90zo+rGwtXC1/lL5EjaMC79Q8Pl5G454BCQFdcpBAMpmZ
0q//0v6D8F3wDze+kx92hr6xgWo8A75p4omaHD/ReBmW6Ez/JVNx+wr3fqVhRxnC
zj1cZREmE7cd9irz0lZGZVqZD0cDuvjMm4o+dNxZwvUiKxacviSyj7dcY3FN522o
CRyy2IFV6E90sWbA5WOSwnxtP3qInmxRbJg0JzixCBfK2LiRc7q+3fy3/DGpUn0H
wDL0dF868Auohfgie2TleczCG06/F+/OlIxcPNVnlGGeM70pHW1N8vVHm2oYqG9q
vCl4Av/XraNyTrI7zDT+hxLY+5Kw38Kw48bTGg1Nak6y6LgDe6GkPzYEhG2NBKlv
+k+kAfvpjVdDL7VZlCbmkPwe4hwofCc+HvtMw8WEGOmWYP/QBcUi3rfPW8luk5sL
1RGHw8qbRz5c0oc1iFV6TWGElMwBkPAmemdX9iW/pI7723ab2oys8HvUrAsf5OF3
LkXVz+khqzaX7TY8no3nzxgeL/AhcHIt1VY1SP1iLdEmSPJjLV/UbDmfhkd6EaOn
281fpi1Y6JQHvjJqbIxU54avPMcLb6iTyGu2C8QEEORVmdK13DOguWAa+99NXtT1
vtG3deoXMDQnDjtII+59QJ8oBGdfnqfXEogtWg7JftsHJyGgxy0L1fMw1CrzazMY
GbFUnOgEyyItMpjceJ0iVjOvCxRV5HjxEIaTGzxUALdAdnzvF6sLuhp9cuH0tL6H
DV5wWlanJEMAm+PuW8zV/0oxUJ/W92XH8TvndUYOXUHhCdEYEcjutgJ8KrcW36bp
Stc13feW+GRJjldTHUMYCh5iKpj3vjLDOOHrBX+5qlDnR6QDRwWNcvx9+ae5ICpk
5YaHBYkqXSfra0OSqC2D94EXSSqPicIlXbiB4JHhPYMICrs/tQPaBzJv2zeMyWzt
7h3wZzMFJw9orUv7zVa3dKwRv41p8yLeB3z4tyMkPgpKmflZRXFCDpvH/vZiEA9l
uF3kmu2xsYZnHBwAzHNEzH98hhPhLasenEO6s+tz8ZH8AZn8xVnrHqll0cXkXPGZ
qOA7X1CUV18tduSRL7iK3lg+KzF417En0p6FQAI4DC9SfsuzEWisshheK+kiWHV6
XCjGTJakUaIzBdEfatZdIwGeCzKDuc0Gw/SD4cQPbgGJz5lLp54PEw0ffRVaSnqz
tWx94IRq2+VSQUeQ2qotIvoTmVXmtssu8QWOpSmqRRnAOMYPPaXHzuLlQkRrJplz
Rk6KIHS/mHn1FeoMdHjWR6sRDjJLpyb5uCiOj/hWzvoJyzc6ZsLoEriUE06OcAtv
jWEo5Fh7uDtMhDPBsP2bz0iU3e/wSjuZvQo4MxAB8V5kBBSgfinNXgJNyGo7jEC/
f+xJnFL9VzBF4PklLokKhX0VeD2nn8tm6c2ZzV/zqTdPbJjM1TsqzinMU7NPPHW6
gFPDBbWeni7C7BsweXrPu9rdaqtKSr+sxquDVaUDGtb/HaBi+48idxoXhDPtTAjT
6ZIOpVzDtkey7yi2hKtxf3nEgUmkiwj0CS93hToCUWs0L1PX+iSlpTN+PzjkBO9I
jLZfKmyKDBmPPwr8Gw/HV8N16miDQzzzYrp3r0hui9Dv99YNOmDCyrGo1TFNF3oj
m8zitI99M21v5guBa0fQWxSWy/rYaNoAjuwZFJLQgbjOnQ0NS3TDQLCX2RnS1Q/D
qrw7w70Ajm5xJ+XFTBJGiZ1jRc1BGtnvpsHema87wmdKplCGgE5pYkGrN8epHF4k
f2WZqlP0lNRUJjoLmu5+xIwMYWWk1hcUUY8PMPLi3QnZWUvzTHIMA/D7r5V9Pd2I
FT7/qWkfPua1LxTDLYBXgLVyr34b+PvwGA9km53SLvZG+gkWig6o77hZ1DIbFHWs
9sZsCiWBpWIUGuy6HuG4GJ3dkuBAnbkBUG0C5zcHOpsO4HHupRe3FD0XwTQygOhn
jrtLnIxXmnBJbVUaAZoIQWOxeet5vzQTNnwyTgfAYNldnTp14Jz2lqnwVgZZgTD9
jmMiuj99tkgXKttG7X9yChYANuxrAAypBk6BwLPZm+u8XUSjgUYCDUMi/mi543xa
5HnEgTM763TVARjbaiRBJ1KuyJFw+oOfSboiX90MWO83TCk/rHLI9/fGVjg34623
l+RhK3UtYqG1kgwCmwUgxx6IOSD7oHMCPgL/MbT6KOMzZNVm3gQqkhNt5s2eURfr
k8U6o5R9nljEFxK2ZS9SxMZ+SsuLgN1wAGwD40hiyX3K3l+VvLeoRnS92DGlpnnb
CRwMCliV1FRmqfEL0fQeKkzNeBA089fL2SgbW2pxlXk6OUgXB6kfCfXiBy5++yWN
REBqfRGEDAGFjMB4/MxSNNZ4pNdd4LOE/4neltbso9rLdH1Py6NLXrX96+XruFV8
IQGF8lNntjrFvoW2TTWxSPD+5Ct7Lpux1gYH/dVfWx8hG7HcPcDkHoortgnpvxrD
hQexGcBtIXtfCLuG1SI2Yc4wisANDyAObZKiqnq3goxRqp0ydPuCpcmh1g7ZxuJ3
LtzeXavaPntlcS3RvKcHvmguvmdekseuLzjfeNni8fihH5Ayuxr6bfqbKSh553g3
h75hZUZi5Pvj4/Iq7b467u8fk5icHxrxKe60faL73RtFteRRf5rwHQi/y19YHi+6
4cGSfj7CsOuqsw1Fh8eKOvFFwAx3bxWl1tI1/bjO9+tmWGyLUGGmcJUaT72WGRNR
L+yacRRWV1v4kK1DrGqZO86h++jbUE/YY+Sl4dIepC876Yvo3MnYjwaIV5ss/P2c
JQY0QaRYwfpehLTO2bQtJH2MjHolpeVjpH5W8Q6klP6k0UxtrAyj2rVRvR0Ubu29
NjvxcMvaBdrLb1uSpcoSwwapHgByqykPv+yI6wZ+SkE3VN/6F8HuppAIiID89Ii5
2tD9tRYa0uwHPkLc+57C3Vi700Sur9cuio9YOrRk/nlhUbJxbaawgYu+SR6UgsPE
nQi2ixpchhuAappFI0O9tMcse6C17arx9py+R3TPqyWXC4+6WIPXIR+VDBn7Q3W6
VvaN47QDwgfo2ZIk4QMqvjVFfVHbuGCb8W3U1xqmeIuEFm+APnPr5a+Y1oM73Gwv
nZEzZBQYcDh11XojACOOBwMzegkFGDAwh86kmksXl638lmVxAhnaN8vcXub+uBra
iPsbnPPEsHCV+i7Wf5TWPuviCs9wnhq7eF2b7bPlIoTUW2sXsSQxNC4SKH13r/q3
tTUfBwwI/8wcsRKsZ6M1KnXYHXZhjjvqHnFe8jBYZiJChVyDIEltdSqFqLEwkihA
0zDj96UD/AmwQ3kRaLHMeRf4I063ruuZYur1zTpt2mXR3/Z2/HIcFKmZlPPtxV1z
2qU69NeYAuTiS4iS5csooDNddheBxaubZOjVFTHBYplX8YkPzUKGK78kN15vnDW7
5GHtFdsvttqArj9WGBOICkrj1Q8JcnxxL0o13BiDRJJEStFgHo7xrh9WT8mKPkxq
mFZPQMrdFzdZoW6R3TM6VmCg8dHk5VwQoejPMP4ICkS4sa4WMpPqEwu5V+/QwDUq
QYVRLFHHGf33vtGaLmp5oVUCdZFjzIWjE2AGd5DudhoceJVyo9N4/14Bpc1WaInU
v2DCbN8IBkEaXM9FdcsNZnMr0xKWeX0SjnEdrVISWDqd49TVB9AgZ1USXdbHZg6L
55Ribcx03f5cRCPtmfQ8E/UYF+NFhFl9D8UcNKKy4obtL7qX0N41oVDS/TW5RvxY
6ccdBlTe2S/H+ZZPdooC2M+2an2RMthTrr52zpZExM40Ldw8/2sqOQvUEQVx4fvh
1nlVIzkSixDLFKdAWmqsQSQjOtl8j/MVcWIRAnmftCm8JtYru2nfLIDyBWE740Lk
s0nX3IglcCFzpj4AEYMzfeeqCIuGraqJi+Oo9KDxu5SV4fguhPGGzquWOxjGliFc
cyuBJnqQbfgmwN7uOLo88Mm+JcjmEXwUEKFf2WEaPcHTpYlw6VL216WVQdAPFBN3
G1q4Ed1GA8WgUfFTfi/mEuFVhC6EHJuKzuCTUYl9ycQZPzI82NchwUGcvn+v9Mwz
EKxRD+u4udugoMnfYeMevTlkEpYN7ihBVGviDNrfcQLW3WFyisvAfO73kIhqHsrE
P2hdXhM8KYQBQyxCRTVfvDiw/ZH+pSiqoU8pboVyXmwO0rvkY+Cw/p3sq90r6n9j
0rMxykwnRCKlY9tICOS1PMEXVTVzwWNPwmuhHzOAphl6LKLYpSpmdxKi9ttXy+jg
LTHvudp6mrly0FR5+hrCywwL00DkO5O8jTU1Z4BAj6VJi06ldtWdOFxxkmYmE+8x
NVKvIdWYveZ+Es6HCGw2kaxqVEXhL8V6PYyc5TdavAefncSOyNEx3OGmyEOq3FKH
LtpEf/F8Q+dcN5qWzHag1jhHOxxEgq/suUJPXBvfhn/mpNoj61IGGqCOdy1OI6sx
qETF1k6RUhWTuk/75lN+2NxYdTvUaCSPaMcJDezJg5qv2wzOZzgCcOiFX7p3kIiT
sUcGy/oDDqG5YRFXSLA/GLoOkyre2iqVw1FTOIzOj6j16x7ml2WzBAld8c+PjFG7
9wExfWj+tIOxAPSK3y9fMzsZRNHi+UeG8bTbDNuz7W+5oRHivuIL34HxGO+XJ5/R
35ory3E6q9uj4cL8NNvhUEP6UJ36wwpKSZKqF3XJmyqLkmgUyP1bIop/D8daR9O1
em05KUdTXBdmxWutuXtyc0vmHgys75jdTh2Np81q0dvqE7mnZoM5xIlE75wFaxDq
mr5s022Q/KyGxfmiXzpTqtZSZmSpGQ/qCufKs16noymxHIE0lIc5xzVvqstRhcyN
REOBbZeEIFXOCnDbAE5JIz17ONc7G81P7GuD7NXJszem4tCgztZZ8FlDLzegz5HC
lhtZDf+zHFFkznrN2Cb244sRpr3eW5YI3ZmK+Dt7oghz3aOVDOxij61mFVExSS0G
lP9n6Cx2ijpMFp/PejrdEd4WBNGAN0ErkYK461anbgx8SFwSSeTjTFuXVMzcQOQT
DVLJaIVfXgdU0U3wEUFlchSnRNI9W+HnzJ6GqpzOASduFBNrT6aodAHHhIk+mw88
RFYP3yDOBcA+Zce1p9En89wlVUwyBsfOcevWHSsIiy1kSuv/xGVxlsefQc0r9FpE
ZeoegRV4sc7qsP325/QWJePxWDUbe0yLM+3Kg6sK23WB4NtHYd/W5+kDd7in1aHv
DPlYIyaoS4SSNd6mJFFeItXnNlaY05omfV17EKfIXKR99qPQb75byFa8o3aLiMl6
ogMvr11SGJptuY2NJHqmSHPJGD9hRtNhc4aROc/t5I4LM+LaEnd7X9mOimYDQmhI
xvPulSwkqSn/hAUCgeLEsqsYXgADf8qsusqjGZapshD17ofNtkQFzuzgU1w0UDp+
QdKM/AQtL3/EhSiO8x53+bwmJ2rmbKFYxwS/b3jV8zZX2vonTzm3WkeRwxfoYZW2
Tr5Nr3PW+iWyIG0TzAEVSlrhr47fChrarObzUupNTpq+y7lbvOP1BtwfMot+LlpM
Ac7/VkX1eZKLu/cRaS0RVAJ0YPFEgZ6GoLXdYTGkNLcbpDLEpj6sxYPcR2eEDmsR
o5ioR/0wE4QZQwMFKLcqLbxLxnFUKsy+Lf/UGqRsfd3L/ABp8carxAdqspQtgwGL
xW81Y+7LTZKbLYavacSf4CEdlupELSMJG0qsZlsEEESo0fwxK6FoV4e7CTUJd9an
7aogtq5jqci0jAGmM8UUm4TcyU3cTcAtxDFlBPsgnRNKUMrxJcIe0fdzE/DbAHVm
NH3v+btjZXuR1M/pAYUIXUiAhg15jLkMOA+EflMZcK4PWJNtOXI2UasThpj03bXz
d7hvAbnVhRJx10vtre0najoQGzvoyuO8OcXhoLeUgf74ezFq9setiXar8gQ3sNST
zYFHZLkLGRS5rYA8I2gCDtDHXXsOGZlZ6z08wC1Z8u0q2TJnD3ljlMsBx0Nd2FjO
kNtpgvAlilZv0pwR7q9h41jhcJuEWElE2N3wSWuKp1bqZj1zvB3I3RFg78j0ejEm
Ht17UuG0Ymu+AY8RaVqwB7DA8RPE8OMdTw1sv/xe6L0Y9rNK/gAslK2ebNHBHDGy
4lf+LgiL26+6XXvX0NI3szEA2PouWYWkv5BIjkts3XWLM7a25/qQ53c/WIzleQMH
EnxkQTJUkAXDAaNSqdotEtK2j+HhpSSurtGK3OEU3Z8lr7h+MH6zbYpPBAKrsfrT
eXaBvu3XIQ+ORX10Sn7H5dlU5QPAa1wkFI/hxTZ1+iCiKjuxrO8YlhOm0rMrBkS4
WJXEkqYwTAjtxzzg+mwncwiZBVwqPVnFdjAOndHubTe7CyzM/ex1cs+sEDXq+TB6
Wp3K6JPQObKnkLBdTJiQX1MEbmSFdI2VhRhykVxew8kFeeRZId1+d40FzgJ5eZJ7
Ka+jzOVON8O1tItOuzP9UCOS2F10D7sUVSKgJ38iMX+tMkOaB2iLLDoxZiH/s3fj
RYkRnOCHZ5EPqcYqzH3I512bpXJ0LngWEVFbtjJgu66FBoCfvqY/mNzV57wIhjWX
H7jedRxf/AXKfVBzaFabqMcpMWQVQmTsujlULIsEPcBIYQOKpJF25NfjK3jPKQ4E
qD/5RjSphNFru0icHCNpT9yeg47XkdkHx638TqpRN2UROm/LxNF0zasF/0REeBE6
7OusNbbl4FkzlCq/EPhcIJsQXN1uBpNZZnAqh/bkROSgBMizHb5ZDud6m/QJHGaL
PCreFfFn70+DgIOYzssa4DQdcPJFPk5AZIJ+JwohSoLBTyZhWMrwAjxB7RmQV/rX
CovKTksii05mjWVq3RPZfWEyXt/4AI5LlbDatW3RWi/tWyZovBQbsuHET9EFY4Hl
b8x9QypOnDxAJBaQkMGPXk0hQMHn3Lj5SnNvb6qeLnVU1SBl96AbOKPPctNJbqhs
MgsoSa7tycyGS4dokwQPsDOxwoeQpETfmxff/20h/dEKSM65zBStFcByXL5uJf7F
1NgS0l9H200CS6CajCrFawmHbSsoWJVgb1TKyWmCQ3vDOUcfa9zfkGo7BRaxmTkl
KDMEeyPxT1snB6EVy/eStW+mxklLFFRsYa2a9l9RjKyqRBUpqVfjxl1HAOhcCVPw
cpYTzNw9SJiUDIdRk6K9qxYh5gj7o/5UFBHYCmmuYbGzLQA1bzI9VkMhIRstisEr
vRfIM3+mZaIpEqaN01BWZGJQ174TGDeh8JYNrTM9cVi1kW5TJCN2VHSn0HVK3KZx
rwDrntMb9ik7kbjynnFmhxOmSc//SUj71VB+i6ITFU3x4wvItSyoIr1v1hNTDPnS
Nf4lGCpAEW5hseAQs3uLaLDzPsjJxc886daYouA7tqJyGCQwsFVHp8nYYWkS/6e5
ypbmU41vHuknitjOUAXOewc4t1UD3OZxiL2lHn4FKzW0rKfhbESajf8cBmgsP8xU
Obcs/w7b3iphYsVArZvmkMmVShXAuD9neJSyS+/kNn4jIx4D3JbXmYFkCiOcl+Ey
Cf0xd7rOE0NoC5cygvPIXuSfq/022T1f8/QkeFpVUK7+WCAHI1OTX/jEouLcUAGL
LJu/owpGukFhnkmDPbLWBmLktiDB6ZbJ3R1I+9U6pRbOQrDk8ZE3yOt3X7mmXVRX
qCAiC6sG38G/3hdq/NEXZhpWMEvCkFTxBiJdSXgwQvZim8q4LUZckRY6Gs9op9Sk
zITq5IMS+8tZJ/ZHdVhQ+LB5K/uPMHISQ6AhsqKAq6W18ChetPWATsgRQUEKXnv1
LmK7dDwHpdMDIPYcVEogXtMcha7To/BguZEJDkOL7xOWICC15Mxlpd5IC4TohQEU
J38pLUMdj1Na/DD5IWGkQzPPqimt3vFBXSW1Rj4CDnDpqaiF/Z99NFC2ji2ol9p9
ipuiO1t1lnTzndhKtTJzGGXXIUOCBThOGKw/bclEYSssPa3sR7J4zipFkYuUDyQg
s2lblc34gUYGe9SxCX92msoTP4FGM0L7tRFpnxJjb3Nem/JDhAkSiEKs3g3CcVMx
AL7XRpyZmdPDi0ux69P76fxXr05CIk0y5Iw9WtLrTsnPoRl9o8wf+jVUoAnLyua3
nN946S+6+7MF2LYWEif1XuHaLZA5C26x+Dv0pGo5IAzCH9X6yn74vTUGDKZxbktU
Qz1qPvPbpLpl6VZACnKo/+16y8TVxWlculnHeM21mavM1T0u4pdqqvhIfEh6An5L
dzDEl2qy3ST2RrCYMbsKA/9C3nJHQt34dj6N3pLqG4foZ38+rL+x+gY5MZ4ceIaZ
2XiyyzaRWcQm6jhwwV+umYEGHDnnbRJ+SqsxffD0YrRUKCESCh8K0IRiWiLCTQHX
zArZkR9XYrWs8oHXTjhVx++m7CAYNw8m/gtZ0DYUBnGHWoj0Ul2ZtGw7kHb6rfpr
EnS3WglBHR2OYb4D232EjcKCOKx+ecA1YKm6L3J9Cf3dm7PtPlh7CvvKtdlLP8Tz
c/7lwMz2Wf7T4OEKNmCA6LbNAYX64BeCGQ5JiKmgU7uFuo7om2uh9i4bhrzcOc2Z
ViBAGp888++A+w+0t5ftZ98DHif+KBW+vdE9wNe2EF+gJTsdVSMu7nRMMG/fcfEK
e/fRsVGIomXLXDyf+m2bJBcQOzjVTq93+4XfdWnfbrfrUceMIFOC6+Cs/lLY6Z8B
Ib66UknRBASWpB0/Pu1x0OyMIT1hVUDHk0Oh0WvtNPCSbBzdi0EXHzYbo/0lB4x0
zVeTafKEkSXYdvnC8bMst/RqeHc8kaoUC4zgJ3oc2KT4iz2WNPrIO4Be78ra3NPx
7fJcCtVFP/nMKI7eJJB93pasE8gNmqf4S/tnA2u/Wbe3f+blgpUpD2zMTDvUC929
SMuM3x5D4R8XsiK8e6MOMpCk/bwZs5bIDTzDkAQOtihQ9ZYVZmMiFx8btfpslql1
HTNdV8evSU6KzBDar3EPfAVPt2noIG4ajNriNsPlV1Au0QWqmToYP4SJXElMeMxK
MtuA0Pvq7Ylz57XBdz9G9li3m9i/LfNnjLCj+7rXAzP+vWTiSNjE/M8MtaNm+WBG
QfCCxs/c7Z7pyzkuxe+On7jhGB38+JHzY0HEG8p5NFhcywAQ6Ujp9xFaq2rc+6bW
TD/uAA+WifEoMNIWnv/wIfJNZCWHIKU2+uJ9nK35pu5djLD7QD+lgG4mMD2xTgCs
PVkRGSC65GuzdeRPqo8I9FxJ04Gqp1F8cSm/rAgC19T4yTWy9tcY+wGkLz2cWtSG
PV5fTU5ox/fcU/s//Jq00ttHbs43L3bqinUonn6bV7dinotNlrzfaA85qIhCUFtX
5f1lbLcPlASrIfw6LFQm4Hsi5SxOYO+zUStaTVUgRQpT8yP61ohn9po5+qf1hEB8
UcG7aat6I1W96AHYQbzueSCLzTDhzAkKLGR+Or7wZmdoTzgbILoTITilajsHlPf9
cNPtgvSTbZuRCPNb8OisNBcMurG66qZKi25zhEzQzO4kexTJNMtXMrtvL3WnBYc8
zas154sohKw7TzrUWjEQtwAKU2NXm36qvakNZwLk0QZ1Fdzc5lDhhfEzwfvnOPMO
UDisRy8ULyCJGQ7I1OpC1Ca0FKfI4TJ2INeGZeUxlh8ChrpOwVN281uHZeY4apaB
6Om4TA/nxqJv3rW+lEpK08NnDOgEG0TLezhkVrfsPdGrOY5CIjLeOQg17MmTFbqU
nhFmVRmt5i1YmkPo+uyiSvX7omC6wdiMvid1js5Jr2ItPhCBXfGb4uZf2u3aGvW0
bpFbqUZVB7aq3s6oW4fsvTyFLJ9xx/aHtRjuQWbGpgfZO4QbufwqBsV3gglUu4Bx
GP7qxlIrZiYJnfflpEoOatOLGAnmrvwbkOSj4/gfqYtC4t06liI4Ih0AHjMblNOm
sO+pLFoSqC0UikuEV6DqWSRSPqHppBpt/zuPw1YFM0rFltePWmjV3e+WvWll6DI4
I/jXmGdpBKLcEzBGZoIRaFzawQgkrCbOBoVQolFchhZZnXddAlhKVIeIkR8P7bUy
bvkiWRyacw3VynylFbMC5XxoqlvcusvdNvIjBVZmV+HoL0RPfgvJUKUn4sVRkfUv
b+a7SPKHjqKx0++FRzpTv9+Fjk8pcmd7XsEcp9N+aZUHdQmp9xXshngHTgmYUgxy
7ej07KVcdOXvJP6ddaUYx2k04yaJPE7/IDSevRpy4zihkqkZx+5A7mFs3eMvLGLO
XWaywzpXricg0K1owxGfLQY4s6YbjSNuHPR+YK4Az8yhrkNRlyjUNKfhz59OqCyM
h2i0gCU7Srqw1tGyJKxUmRIhn1Zha+VsjxZWpCqOpsMcovphBvJvlKkHCQ8WR3v2
pQN2cbLN2nU3VnRyU0WOD3ZAwMrd3rbmdanlPHkaZO+ADzCXfWBTIWnNJFPT9LFY
xXd8yuUSayqP0OZjfxszlDVorgIWOfaaIvEiFDPH4zTCWrFtvmwqBrP3+AANSwrI
UlwEUBGOYaznRZaz6ezrIKRb/ieTznxdsIWTHCgtsUapjhy5OJzZlxXi0ib2WPA5
+2Zn4sy3J8QH2/LO3PRGmvhCez7vsdH3KiEx5cI5kJGI0zb6/k+8X68OdzS6snE1
B3hvmp0QmFY/Ow2wRgxfSQqx1kbwbd3D4ik2e/DD4O1p+bnO0KSslvadm9mP/KzH
9ci+OAtXpVmtk92irRjoa6WdHYLCSWgLs6scVHK7mjEqgJtaPNT9YCuqQTLf+K7y
ClOrShPYCde4dvmL1uCh7Ky1BnwdJkgSrI3BXfCZ9xRuqNudQ9T/pS2dEGcERmnO
hxi4IKal2QP3xs3+SBHF3eSMHbKEuf73LbQDD35FMnfZfmvRm2OEzV+97LjRTrPd
3dCD6yZLRd3SSaNaUSragWLZxmZfWIm8gM3VBmxkk1ylCzSwLflwJwYmOpywV4T9
AWDX/zlq6AFw4B1uIQ97TWTfWrqrDKjB1naIpzMYVhaenqG+eHKg5y6aCM7GHfgT
2UxfCAb9b+/qV/SlLlmi6ZOI1Seid8lnd5zW6EhH8zzklwMRBJ1XaAKdAQY3dZ/c
9noRh+uu4ecEPn5rsL/qCZyeVsydU6z5Usq59jCS+fXNWkivxEbdvXQdg9IpDN7D
41xIMtl1bQc4qXs1dXJjimGm0b2eEb2ci9LzB8IzN18m3A6aoy8hSw0cXGWsOQso
O1kbSeEratkK3l2IPI2QqZPIfphmMP9XjJrP39JiOcsLYZUh3cgxCdcr1HeoGzc2
/Og4KAw0YS5J3O/fOZtClI598458F7Iy6/6sktufrecFSxdnVNs4YqgN6rs5/ydv
qc/8taHcGm0IugobrsYL1Il7SFy5k8DzewovaEX1i1h4+9Ktf19MlIYKe510mrQO
4DWtpvq9ngU51GwLYowcdQZ9YKwFKSMqmeJuOBo4ZGZHOmICIf1TKkWmsaEAUg2Z
JgaEK/1uTyeqnDT4ETiTJ65R/aulfvx+v/9MHfnmECoSmNHTJ0rQhLm/WNKHWJoU
vrhRrFtt52IEsC+vBhwtnoqcY790eh8dyj2MW8u+L0sQouZKbUW7H+1mxkNZ1qxw
O8hQ7hqpdtCi1i1Zp8z1N/sOoxnBIfKLo2v9mSI3LWtF5OzbTDGsdXL1DYrqUpmu
3CZK4Rs4iMZ82Xmx61Sh9o/ZuVbWz/RGUljbOk4EjHHQIWr5ytG9rRllkXNYP0rs
/duC7ci5gwtsza+a50FeY2m9+ybzonTnK0ziY3TEO8vHwbaQ0kIEABihc4YBV+3N
6n/rlrLNWn4c2PpGMBKcsyG6cqV8m+LGFGm7FacNxxDS7DBnM1lPSxjo50y5yLwF
BLz82Ie8ZsuRCkLc53b2Atz0oAblMmeL46YKD+PCwXmWdkFYxWimoXFN/+HOIEPl
g0j2fmWdjKits607Otw1C7nJUkle5uxAmZpbVrsgbQftkpG75F884hTxLFWAfP/T
2Xo6Y/F+0Mo5xIKDXL377X0Ep00jsnmA4LtL2KPolGM7xTiPrZLkkhavMYpnFYrM
MGrVAbZGnRSAV/0iYAuV9dfBCb8B0D5BoX9MWNau0kIyfwFMGyESZBbrnGRyfJsn
YqCkixqtaP5f27BkKInAgRJLySg6+QBrU6HeVwsoqYpWiX88v3ApcbyjPAXbzX6D
frEsWcHI807ufo6m2ciy9sI4+4kMepAHyk9VUWrKl7Wq8lNBtHXhdtovm9cqCoNb
CgLrWEMn/mqQowl1M6PyPiyG2u+2ajc1xkesOtMkzWEKEDfQATseZg3vh6YgrCgD
ilTDIHtUaGdNJGOWMoJJn+ldbZLMtKgr/y0GKJVK79wL833v9VE1jdl5ZiD9AVHg
Pur7wZc3OUw1PbfqdVkem8YYrE2/DhrYY22QsggTv9SKRRkLO+lKxS+xWXraTWFZ
hkXFrmMv+YlQrFcSxSiu/xXDPB0ZzGrun/d0CXzZvOsP7mxcKN/Ze13CmfkCwhUT
hm/DTwLEYejPeZOw+DT1slG8LkyUpEIkQfgQ9hB8Qffo9PUJtoDHsYwRUEwsrxir
VrlgbMCb8c9XzlLtc8yrE1HwP8hVW/h2BwEHsvzlbYeKxnWYCrbDQs2Qo2w6wqLx
0FuGdzAAipRa0YWn4bQY3OuWS7HxP799oxS1sN8y2gHWVHyfHTkytyvTafdoGdX3
XgTFDyBTDQUVOYxjjDz0yOsZH14doBANigfKHamlWPQWB5KPwSHTdMJgAdJpUgKn
yWmhwjj4FY/9Sq/F0DtPj8L/fJ5RyNsjaIDwyjRPOK35D38uuipziyec+t03D/9c
lOUovrlZs6HXYR9uMASmEYQ6cbrS41FITk11Y2EO9Bssr3H7NBs9iOwbl/83OE1X
TiAY9hPoS9ujuJlmKA/K2CcOtLpX06Tt6s2stF76H865sT22xMsNzIUbzpEwVEV9
sMEUTDAoJzrasD4/Cj1skHIVMPg8BSFBry1h9vc0Ob00K3tlssdkmEM10Nni+86c
6PmfMIevxa5ZKnCBCROVa9q5C0ef34MVdbjx7Z3h6bSnspf03yucZGyJZOYRcDaI
+P1nS+6lFjXuUppSMY16SRjJgyfTnFAFzBfs3HSSN1GzDudeTGIu8GDWnRtxb8lH
dwAxU0dKPST+VvIc8Ipy60CYk4A/WbUzUGHz1qSWt5KLlMYcSLrpnXo34g6M68xx
RcMnvm0AnHd38OPkRgqQ7jiZLjm6HUJdxj38WGrsMHxV8yQJMJ4r4XcZAgcgS41m
G29OBY4wgQXhVD/UHBdldw7Kg0cIX+sbvWH78kjFEOPSk/7EA6ibI7Wb4Jb5fir1
u7qa2H/lcMOXMg18FI6iqlpW/ZFB19bVOQXI827yFx3XWB2e8hpdRoGekbdYnte9
TCGelIHOUNxbNem9Ugazax1/l08d9EaNNfB1uAgwXcdVXaplSltONUvcbI7x71q6
i9fw6whL8c29Eaf+m2ZWzCIWH7QSKcVw76m2bmW2MHXFSPhh7ZjVSAycY6gJf7BM
qLtcSiViTsg+EKR7vPcJMccpB6U0Xgy7Nqvg6vcsXLeQiQzTpFLsSdnViJhYmm1O
WYJRdrPRlcm/PwoWM2JipOHYDjwOaL501gOleJhm1z0TgNwbhX0HBbU3As0XZ83A
MHsixodJ/e/XZeErdV7jx4ICAdewfynYQZFhovQnOfZYvET7Dz89u0uS7z6iacTn
ElnhnXufni6j/Rk8Xg9zeemHcdJkVxaq/yFo+AbzdNkFu0t0DVSZVjUFrZ9nykZG
GcK5bvrRo7cxBeiEgw2lCUyMcEX9uuTgUYZbAT3FkU5pY3BoTJtNLUqotz8bJpme
xqGyqkvIY5ks3Zwp1PPgijr2OgAJlqXK8bATxfPU53b3GG7Jjf7GuXcvSTIfYz0s
Izs1OBZPMcAV3OKEJgquNslW5cOHxzCzHRCrGKEbM96Z7RuiXyBAjvWjIjKQb2Z9
y88udwbTolHSoMaZ2KXkvg6kiyRGYl5s4Y5ceHhxuN1WMth8p4w/emF2q+DOOMw4
Y/BnLwng2NSZKHJffZ9icBMUdP3+/xId4U421Lpt4mYXecaS67bU8IK4HNtD2tAq
tN7gJhINhdxtMlNWlNiMs1tcEmhuCbAwF3UI/2iK8H73eyfs5q3ncaKl8VOyTv4H
bYgkaMrMsD8/Xly5PxMExJ3002BpxPKOx42M6u9Flsik3cnk2rI5JTD13RxnW57g
NtHRSODgZzWRG0s2IYX+L5F/TMpMxTrR8znMZksHAV8lM4S8L64B4D8V2ZvT5XHq
OJmuAR/Wlz7hvBDurMU6hNfGXoNr7uqja0AsbjjfADamfNFMu4s3UU9CNNBa+k6q
/IGiUC7zyjjyq2w8hSvTEZF9QLRAPFrN/t4a33LYdCRji+KTRyZL7hZEJJHydHxS
PvRMpzIZI0fBzAUAhu86T46OwuGkV8GdDr5X5NoTNe4wRXje1K3cUsUsIGzhOHpc
piXhWlJoE8XVKXY8FmkSBlvkHyNLQZmJ0Tc6gSyOL2EIPrpuTrzQjvxB/EtMKxDx
TJCpFcEJKQl0lfJN7FyAqnG3T4wUPZh67NSxIEcjSJ/klAsp1QWRy+8u/IQxkYQ/
2f73fLCe37v/7aX5zUB65/tnwXS9xdDuCR5o5pi44lswpVPsj+4ihCt+dJ2WXp4W
r0ffXROWE2GEqLwrjERJdtHAXflW473OBk3UOWS86AHMdPj0WeQGY19Tp7vTkLd7
nr2z+HA45oQWno+eDU16/Y2s4HZCWEpgofvo4oFKteaDNM4Vt9vzAxVZa1GJ6Vea
Yqg5uanIzo7+4OC3dHNIhqUZcew+8zIt/ve9/mXW14FT6nt8YmzKfT5GhL+6W89C
C6SDLEIdx8DQ8aP99HK0Y4j5Lh+kA3wgVPnGoxFsa0s7FNF56Wiwxs2LTtGpg0Hm
Ql4JS44u7lNxKpwM17i+obZ0ZQLKw5k5x/hU8ZcP/KNLZV111DyfF23UJkx0SnpT
YzTuhyOP8gL2BjFAh0jV766l8KaAf9ocOg6+Clo4I2cUo6qzS377nuDkeCEsIu5j
JNWrEkH2FH8x0r+3LXWAGgIWW8T7ZfzcXAUIXiV2OHxIrUSAbWRLT5+Ez8vk8KN5
mvB807YZ3NxFTHDb137HyoAEwiKwzVWH0f/RkM6Sw36nkvtVqIbIVcXRBMepJYM+
2v3xlfu9qNE73mejN+8ICHvwoTauXQOb00T1idwtYiR9goF8xY45Uyuce4yqtjS1
JiWIbsnXAqO2DvTjMAbRNtjwYYP4qTsOYXS8oDFmL0yqhoVskSWWGfM+1ZcVcfEH
VdRS5WqgHvcUZisY1QNUmtjHbeTAA8VapN6lEF0XQbH8AHkqxxXfyBX5/BCzPn25
8QhmVMJW4gQcZVyZKClJ1a4+uQAuuuJ6MhTYGAdJPe6MB+MLoFQIzKWPmXMDQA5b
Qz5+Svet795vfX0gnE5c+MU3Cjvt5M42LQoEJnuQrqz6ze7G40ED0qo1OzT22a3G
px6e1HuYMXEReGuY+0yuuxvKwIa1KuwN7XfGybWYk6lv9ie3SrlTDD+grjM+pCkn
JXQekbxAc8SnL4Kg9V4hmY0rhmSyhR1Yusjn5BD5RuA0c0/jYeww+j4yjKw8/KU9
fVNPsWeeXwnN51plby9neh6b8rCobP2rDZj04M9VhfxESP6SDo3Vtu8iZhDr3EXs
O0sYCD8qIS6ghAnYf3z+PxzvdtpQwzck0IEJfkB6G8BzlXcyZHnMzodlL71AM1sE
Fu2+qyWUTQBaLIkf34zUwUcsfzc7ZsvF4MygLJDRTwB+EbmlctVYOHXPtepSXCu5
LdXua9sAd6VOwTKTWsLU5Fc31+leX2S9YbMymtS9wzlP7U8GNR8fv/bT58TMTrGr
ZCEGp4kwwFNLCwzvPMQSHQZCl/EIbObhTq/TJDhE9ArYhvMxMqlTIPPGIFsVzpFd
z2R01fxKnDCKT0Zl3FgSNDZyYeuBdN6QD4XnJPX/hf+AI6oFeckDpfWSJ80G0KJW
aO4iPsyC19hxbzBYxh+nTGb49IfxwGDaJe6/NrWo2Mm5UrR/MMjRGGxgjZAH01sF
uxFyGbNEXEh+a6HHq1r58A2OISNOIo4N9ma5RARF6XEVovrzgEPFIA/bum22C905
OIRXwkVGPRx5g6wGFUofUqrr36a2Bq3qYIZm106C+UcVj4hYKZ/BS6RBaqm1bHmy
DaoplViqlJgVfwHDJzqPE+QVe0BZZBeux6xbwMa+0OMV6JRv4EQIPx9OoUrEvjce
l5vwLZ6aRK9faznM/3lNzX+OaXqcclyItJc3ktr7KQem57EEtdFu7/2ME+Bpa2ti
Y8HMu1pYn6UOjxGuwfGaidxBoZUQi3orucCASG5HI9dg+slbmwkFxQ9Ukb8gOieF
VT0LRVqvisKIva/rd4V0LPZd9AWi0hfNmFTrSIwMD/hLKEHkE40AZ60B9vv0soRq
vIlrocJQxL4uPVfS5/UDPD5nBjhmIDhtKdEyxHIurNtXikHZCDcfSZS/gKRWjr9x
EXkChiHL8zWXtkfnD1KrhUPaEE9MMwImulYEUJ1Uj2DWCZHP32/tQ2jAd7CtAc8T
vg36uULmP2C6ufkUkL/N0DgdW+HG7UlFoynitjNF3ynLUEuva36lQtHkR67nyhDP
W6z/jnG04kFIDk1llfHG/s7F0TzgQVqcmo6fvpiLkEvzA0HiSRwq3fA9QzKIi8OP
Zl8ObjY6VRkJL6fyOMspmDId5ae/yX000SWndVMeOndfvZ6u+XuC2AddTYjWHCIW
3oEFPTwCv/kYbqEMMZ5QV/DnbovM6Cj8fxeKaEsjsPBGcgGbabt79Z8CyRG2/07n
xJ+/RXcxAre1EbTSakW7r0FSqZHIuYpBrb36gHxuTjONVZhjSwkV0MTzCnAH6seB
9HeYp2Ahl0ljQcvqIlfrFy+w/jC1umntDiiEsIgPpuLu5AyQHZWT0qw34liVfVLx
LbdWJwHv2Nm+o6VJsrJIq8/3w6dcGjPVHoDDTIE2IYCyCi8ANjJGdnlu2RgwPlUJ
oxm0Bn+DbAOLhO+WfBtBHHoBmuxwtqHgSxHzM5GA/X0SXmNzaXr2+xK28WwVIP8f
d/yyayexKQbUPhHiizkzjXdjmeHfozEGf88uSJUn3wqWQcFesWhVf2usyxYuJslS
jUhBbuQiOQG6Uoduubf8T/p7l7UioccRtuVvV39thdpWsjH9zhESyuIpvz1lrQir
zkxTdX+z7DoOh75nNjHlgrKzBA/ged3FU9BSfflwP8tROmjFfWp44k07Cti5a41y
9xF0trhye2vaKImsJA4zspKKQRLPsvCo9JONObhyk46wcrKqPUbIcGxVyONzfwL9
PO5bktuFmDX2DoaY7KbM4i+6QIw5YdqLcIrMAq+8e7gNT0kxPf6y9PppWb69/xos
5LGVCiz5GnipFYb3FGAUrlw5/o7pWjXFfSr48TEJRCgObYLAQnXsn2OfT1MG7Up3
fjvEgn2RmKOOhZBr8j3X9xfIaIdxrqltoz77faVmprSrTM/G4ghmIcmGseW/3nOP
yWdOdj8qYavX8ZZDUtvHonkyfxuWRwZ//roMFMZSMopfpcZ69zbNR1XafUyXXena
zIlpMxahEX6CeiObgtWv4io7Q4RBnB2nJDqsm9OLAoKf+c1m5IwtEHNfIn9mzCsZ
3Vy3cLDpacv0yG77FD40acDx3Fm793THE5vtu7sxWTaA4ZVm8ntkkkmUlQSSHuoc
hhamX5H3ynuwPaMHESDKhVXa4PVxbNy07NQA0k8PcKEK4kAQKmuva1ETy/0Uh94M
fSyV8I/1q2EuAfXC3RsGPvOFB6ixyVMLNCfzl0+Ioh/UVqQe+cAkeqAcshttYJB+
0z0n0aCpHIUtwZR8Pe2Pfa7MsbhxPiHhcaVZAYjnH9UxXpeZMWPy96FGHbX5cxvt
Mrye1aBuQVvABM0hE4T7Wyp9kDkAe3fmNJuA4m+915QI8IX3SysT46C+UeFzrqft
+BKDCSXJCzyDYnDjG9SJ4kgpBNEbJpHLm+Xo26INCkahZ1jV6uZauSKx15j+/9sN
lNVzTCLUu5L44xMLC/N+xCvpvJlK7knar7cY3xSHo27FMjBMqoXz+jgMlfISU2Qj
GfarIABo8h3PI+KPoZGmjHrz73kjkCpiCL4pt0SzQxs1gxM02q/p5onDwC1D1ke7
bzf/Ztxhz1YZgCIa7kASlbPFCXqbYU+M6V2bEVPiI4FuvfYbdpcLmmzavtmlFwTd
r2V3R8y87/iKiznZSE7h7KmlVltL/jzQWlT+xXrzXfxmo9hGAQmBjlPge0YloaL0
qM20et2Cb6pONW9IsF1/kaGqGaYGP49/Jir2Jf5l39C2cwmghG24K8DLB/XE/YS6
B5J19g/8N6AEvhQQXQ0hZc+naIhu+CDVeHXQFQpPzXvKbs6m/ZWTDQ43ejk0eUh6
a0OqRtDzUoLSRUF9RJpVK7hL55osxTWwrqaz+Sz/edUXbRMlznCXBP7UsvXUhl/0
8h1b1/dZFjYhNcE5udn9JF/Yd37wx0h3ji3iIKcXuQARx2ybquOBwrDwtYLAgvv1
puN6ZjJ0wQH+iR5P5KrqUm2F+DTQSulwArc1o8tLkCXStJDlagPLlHmf0oxavTxv
VtIij1mD/raUXrPHW0bWod02JejGGmTqxrqKK0gP1kyYEBXEAOLj//HVK/t9aKU5
r66nz1d27WGnlMlVIPvHkBGTWJOPDZwQnrCiOk3eUUx3ftW55r0qbKNdp+NiM0Ar
3TD/aWP6tbhpHJQBaMlJA6lV5X9eJQD9WxFaFSES78yYYvzgM0nCl5tdxTxh6NGU
Fu/UmX35JPpeLxB2dHrsVfy2rvSG7u5CclYtmWwUpXVmx7iKFy2mlqe5kKE8wHQa
5uCBiWhie8NyiDtHyNt94FFZ2djms6Pf2A/QMpiV/S9ATEnGQ0nyM2lYE+7CmMwA
YEvmv2kT5SRRGyMWoZ5/+lH1N6CcXax4k2gEYV1UqLgREszsW216vPax70qJ/miB
503h/slSMOoO+U3xfjX6wpEnXzTc1rCPJ+Wp+e3AbkqsFM2QCWGjGEOqDcZbymRj
Kvtl7jSaXJzYNETJ/XFi+l8e/xtiB80MSWGSG2crGIzeL2EwPYzTaN4dlZtXW8KD
Xhmtmm3oytISS4dVV7Ef49sLkEhmlOKyGqI6lGgMnd2QqXGZmgLNld5ucT47S+p2
LTYDVCB/5cEjATFohgs9URHFa+IbDPTHXaSmE28wdPfqSddMWB7Z2ypfK1Ia1WXd
K2mJgh6GzIguq9Cs8YseFyP/+GFlgBvLLD4BolkWIj9bA+N2ISWKP59cd963ZmrI
5d7bYA2Hpi5ef+PrJ4bjxqGgkpRJGp3S2f4XTBoYlKgqco0tNnP2K9JasEbqdEfH
KlCrKTmtnW56q4qEF92kDjkqTDHSQwlJgHRCrOqole3Tkyj8O0OnrCwgF57VwDNb
oZIkCKConC7TRtAQ2W5qpIua3y6GH837c3b46a9vDqrtyWtPdR1vDqtM7wp8R9Qe
AAdR4QFXKpwoNyn0zBYBGK0fa2SuPhzLHjJUoorIA8vLpRocOSZbE0hSWqD95UUa
Buf593qFpBd2r0ODmlYZV2WWBfmgm3k8p9cg1vtZfRMmIhaIhMrBbWmyHjCc03zC
znnEeRUKiPmMNnZQ6Z0CPm3ViBa2Wsm2Fo8TBGwP5hPeJysUs0ZMmD/qrlHK+xxF
oIHnrMA5V/t1chdboc4x1ipvJi3zi1gRW4Pr0YWMWRBjLc3iJY6NfGD8v+vaoL9V
SpOt6UOKRkLEunV7pYrfyE96ULTg4hlsVN0IW9+UM8XAnxfNjTsWL4bu6gclgfqo
hMALg5plj50/3EsIGXmj/4V6hpLO3T4AeGxsfxy5F5XMEkxA52SxhAIHhnkwfBoL
xtZ2qXML48fA91OOT867bmTivMAvUujV4Pl9vEHx2MO+qYb6OMjO91V05lpAhUnw
VaNLlX3HjFJsLWDG+GnOABhq5Q7LwPKb1CvZUcj3zKorodJsaeoL0JND6GZQcXb0
GcS+QiR4NhgO1/xTGWu8hVB7A+WuxlHijC3Q4wUOIeFY5N1tSJLFuGnred4rMyZK
Sfxun8/gTTCQNdNkQp3mNyRRXm3kBTzsiE7aFwm5I3UUA4bJTCIQHuN7yasEVD+d
tjfDAIBP2f4VVPRUvt2cM2SUml2cv9mjCQ045b+lSjqrxtiOz+VW10ZTCrnctXNW
7wvPnshmEFtZf0T/qtoxAnC5HXW3rLBAbbkBiYCnj8sSV316zq6Mo7vj45fK6e45
qd6BHmsXbeDHqljqP8/qqmew5FQExm7JtIbbpp6lTgF4ei9LSdisVISBa2dyYPvL
xsohCe6a9pwV4VPAAlDySAMulaKDvFU4iDFEi1V0lrhg9ducdoKyEu4HxuBnuoX4
nLPGbzr7/fvWjv77EyNpFXOfh+yB6mUt7ThrsEhbeZyqZ/k8eBFSfcS6oxG6errX
+1lxByZ70jrgGs0cdtD3qYty6aN1Wcep3h5GqcbI5dMT5ThQo9YSwX4fqlNdkcX0
ylPiRsD6PxwrIaIc0qwUwFYSzPX5Q/YjgxB4NJBegU3uvDkr2HFnJsCctdky1uLn
Sptiei/c78djeSMWJKRWi49N5VabSMTdJQAKaNUgnXwAXX8+TERsRdiAQidrt/wC
WiD7PbXBzh7rsmV52pRAivLm81PA+Ocjktyf7k4BnDOKcDg8prKWWHbYTspoGFMe
4qD4ASrzYleQiHIMCrX1NQ1EcDwDAieDNpRHPLh5xw6HSaKIf0WBHzoGwongayCo
wljj4X3XeKkIJ7p6IwEH3WAam2ux7UQ122hcofKaEod14e4PrTJZ1o3FP00jmFF5
1Cq/9weK5e+HCWeh4+4ygWijialJY0ySR46TKcLdY9/MNjyDN93xR3dpu9bCltgI
d7sO6Z07s7nc64vWZi9NGPoH+3PVfCrzPt1pB89dzV5qOcJcWKtVTb3NRAVqOnye
YPApU6FKCi0Mi/hEgNU00iEvciVFMZqvBcZ2gs7svSlFIpPdEfdqD1Lqs+7R78nl
fvTza9DHFgC29WfSD/rf8aGgbWhPPkYlNwDYeUM0eJD6kCkE8v8qBBAQJigPqbM6
RjU2K3GQhR0i/sd0u+p1l2pa0ozXJnGFbH7EodddwZ7ptoap0y2prMTzbqTF/n92
Z9XwsKAxyzcPVcOTZAxIbnZIGx5TfsKGtxgYbO1hmtOHViRn6v4YIH/WpPIguJly
d4W0PtQhWpFQLV9xpZ2JLrOS91UV/IF/NNF+54X4vgS/7kn7RPk6jn5DH0VdkNga
xrOOp0fdB3hJr2n9sBJGhPuRflm7TaPKY3uLkF/TBnz582uQ5rDNQwlEqombXl/T
LuJvl2rQAbnMWjWoo637lLkCblzIjDvsIF9rfAWyvaZDFleS/tRG+OcIAVqXFUCn
GorFcaQqZh4rPFSXvoD5Eoji2OrJvbRD9Fq013hsgOX4NNfdrVXORvjhmL/zYN0N
Ao0tBq2TCO33tbATGv1ulJZye+4vN6ViVA7s6uKH8r+7lrm/QMe6fmUvykoLHrq1
ZlxzZD1vnuFIGwTjBx4GycTZQtYpEN24eNaB0bY8uSPt/LJlci5ueU0ODW8VZfy0
gVbQy8fEtzlvCuZUPZkxbPO7TNRH/4JXc/CVhMYbtX06zSolevTujCP4C2Da4D+F
uDV1q5FDGiHXJc2SQP7a2n7rljK4T/F974X3VxODaf/NsGiAdILQ3T826Y2uRg9Y
qbyso+oM6qrqTjYvMUS3uL8gWXf5tV+qRmRNZc6nBxTct8AaSLebW4u++AJ10tmo
nN+1WtmLuw6ijQsubqBqrilRK/AAjLI+nd8FLSZGaSB1ynrZkqtyQtfpr6QsPNnG
lh253lHLJlJU2t2YPl+1UNReVVKdSo0qWHkmZ0Zxd1Z1jVSJosweMuBp5dN4rlaC
KEplJ2wGfWuqFC0g2JwpM4jna8HVlNUswbfaVIoAhlvUnm0QAEQ6tHMX0LEEl4EK
ncDLDsD9cCfHdvAqzaX5q34glKFR9yLQRliauv8NFTJ6mvXEwfKAZn+Rr0DoaAjz
2dwdv6BRvtIWIUSAlFqck7JqLmBlymP5BFKsCEkbvBnjEDERt6W3+QmH0Q/0jsVQ
87r6Tkb6i4PPJlmtWrRSWNmO/f8K3vxBysKUGVmfTBayaMFkB6A7yJw3VvFhGCfB
lvDlX4AZN2+IelRS5rg49wDsrcNUKStVIk1oDCOGsSzDU5TPYcWVjouHbyOB+6hr
dY9yZ4XcgHSSfSEAhgAbMmjlLhJ183aohaJyCgvcIMWZEol2vEci8atZEIr06n20
tQMusLTa9xbz4AsKCywJRclCyYFM0sUtWxI/4wczFJSOhzJbpQPIPol4hXWLPwuN
ok8FbLSvYGXubvLXMsJVfM/XOeaySnfqRpkMZFN/lLnYVmT+CgH0TbLkHDMHljmY
MCiYyX8jxu9U8WuJxnKmZIUtGsdmFJJ3QOHUg9O/nmKWOW9gNQdmNgik8ZRkR9Iw
TJID/fFdUMDqy1UFm4cSrxnGvFL0JQHzKx/y+HFXSWh8pD3/NrmexVSyEJT4xugI
CxFKcBCgy2hn5KTL66Kt91aRXL/IHPvLpMGlLHGcAY3jAMvfYgjz7nEUUg8GuJGw
O2xi3uXnBVSZrCboBieuYc9vwsFB9LZgfKC+eH9IJZDlni0h0gm8ng2wjiQGDceh
w9+19LbAGl7gY6GwnlYpprt0fQOAc3tiZDbolJK9D/6BXhns4FjH8K5ez+j3jK6x
g+RtH9alA9rikpaCHJ3/dtxClE6FErdRBSsYKdiwlqZHJ590rVMB0+G0UQBnhEx1
ReJZE99CpxsFDrNV+mY/opQiUmT2n2+jWRA1JjZG3XLdppVlhKUPTQ4aTjDadKud
AE+2u4YK/JLxE0A32pTrzDdiyqK0yIDQyDSd6UZMutgapE5NQb0+LHLimLpWDoHB
yyI2EEqJURVfUlYshYJgNBLethgyaC1UQczCdiObD9mdC0zi2NIBHssgtjtoFikz
UybKCfyspClDOL109FThZ4lamm5hcnHnQThf0tkocF1tRgKFV9cTkHKn1G7HFh5I
C7WhkQK0JdDm4SUSRAFpB7QeUMBerxt4Lubif7tRIE7DJjwZdwcWXIvVhP/KG9/N
jpA6+KJd4EFzocGUgW7YP2yolG8vAi9FPg833IEY3N1C7SnCwXU0Iyk8F/+W8KPd
PVE6T17TQUj1lAaPeF5KovC1OFsAX2KmZQKyVH6RUp/F83kotUYXtPsYLNJQtoIs
+qc3C3zRIT4rfH9n7AzpqG/QvC7heaG298QXSMp4DPttRnKzLk3I0+2G/rXyMiVa
dWss3Q0qun4ZXz0ArJfmCzmoeXLpUF9963n2ZpP2GkZ0Ib6q+wUmgfTPvv8ldrqB
VqmvDMG/fp0UDAZCRGWOzVKmznhwnsIRa8Bq9BLOpml/0ag3vlK3yaL78EFCBRtl
+0wtVQppVv6BO6wkz3Scgg6nvaYCaTa3k0fpC3rytqpE6X3+9bIBEwsqd1Oyfl+S
zj/FzamPskBV/TyR3JdXETXrZtkDFAaTFTbKy0StoFWyva7BlBXnWjuwZwQqmY8x
XFmh0hcRm4ob5MjbxiEozJVa1BW09wQdgPVWbZv6iZnUhvAyvlDSPMTAeb1eHzfq
MuE/bGWpL8nsUhwJwij2OEs8ZtqaXjdjYLBwvWmH351U1Ts5ZWp8k41WzPS04CEf
KSyLj0eYqFScliXwvtzr4Wi4tkelV8s8v6U94CFP1ezH3UU73dslmSmZ1g1iR4JI
8KLJwmHk7XeRXxYCiCZPKogCOYtJwwDHbUjhFVY6o3XXDlpLv/Ny3RJsv01ELRaw
DQq0sNtpwgADupr9sgd0P29pAJzOIp4Y1thKMmsE6Uj2ICOe+DH7xuEEVv3B3+dO
Vg7+7C4KnYWUU7boD3R+rKKFjaEifnMe19ayL2A5lKe8qBKgw9DAHg2TrXEwlliX
W/r1QiyINRUP6JsDObLjmno2SolD68Fpf0Ct9vJXXlygyI79b3IjV2Ot8RVnsqnM
RT4Jjog2Xo/yP3AQV2UeIU8BzGRcROkxzt2BkyOB1Frz8h1eYK3xghBsofdz8a9p
ArS31Bvu0d3eLxpYqfG3b8pelNOi6hMS57Pak2ERMApQ1vryh4TI2h+PqIX87Tsp
I5fbWMVvURDC0+5YgkHKuQLwRbabzZ5Jte24yJZsA7/yMZyKR7JnrOye3jkHyCdQ
98syw8saj3xc0LGB1VxYALoS54H9hQUN9T+hsdS0UsgDb/Z27X147d/DRRbgjsLO
J0lDbTV23BTbuUV4N3Xy62FgCF+DRr4MS+ydmyseA9hD6ADTJe2D6ythnDOvtEg3
o3FiEKdJvfrEBCXwrUe3H1QJJNMPnihwfWmncDOr15ZV5AYANmp/LuzV6u2Y/1JY
EMTV7/qWAXA7PDHblHMzO7luc4Zt4lbWYOlsTUTco+wf8lYeVaLSq6KUnoPpGo9A
sNgJ2Igv3wi2XZBy4Lo2ySC1kcO5rAqSVKVeFR1zwy0ppe3ALeLYIHDWJapjvsW4
4ftoHBKHjE6Yh07rbR08o0zyT+IC0ASiTx7CSgNc5A/ZKah7bZeEEmTgo5seGhZL
Jm6ZZy53DHm+nHQZBN7P188vLxsY5EPnq9VNT4a15JJaUGhgB50rSrxQaHEhCJmg
mdbTguTOUMGlWk97onyVTSTgNWfIT+rYq7Sd8u6UCXyU/13XWGwQ2WJSp7YeN4cO
S6LOadebfXr21cy5tfWzbHaeoBmpMAJrvl69izMODmRFpZzgE6WKHoESCeW3xd3m
yCBSzUjbzKtKdpQXay3KqkeyYDL7XUVP0aMwEAV8/llDEFPLuupVtUROvnfk7bJk
NP6bj8Kysypw9wTFD2PIoJofq8yv59oAHb4MRqU+MnOcbTbmL3wLjFqR7biBEglI
9aSZA009kOcKNvkXF6JR29OQ4TZNPR1icIugLWsUmSYWHZgLhvJcTa2tpRS5Pmly
zBrA28LVrsbOhXqIQwjOuLFEZxKGPhDwseqigS78t23kLfXgetlD3CwaNrb364Ob
jS1jRTiXjkBFtv8Uo79P6sg/WYm8BROGaY47aw8mOMDnQ9gOgkZT2CzCmMItAvby
NRZNIIyhBZBKBW5g+53fTngYPcYlol6abJ+yZpKmfoXSI33qI9jcugp6pWeXeezd
Iw38DDE7NXWKb+1jgrVKe2KFjOYusrXe6QlCL6Bj+nkCUG260imjAoNBoOw0Tq9E
F/SE1w/CMQXTW5hRRjELwYk6cn2WQttdRMHKPmRTgUduVKQhntVIP3dUg9f8YOeB
mOCzcBUOp4ySUFo5BVgBLYBlbUAMtsX4SKJPoDJCZIZJuEdIvpuLzewuZmUfcWzu
pGEI2bapFvuIN96J/mThw3gc4yzFDvQAHp8rKe1wQe9ERdYwLjScO2fv8Y4jACT3
VM55/G+yV1j1ooOCuwykl7lNBqYbk2ceeaj7dXwioT4qNjkl9im0iwOc7RZoAyxT
Ico4xRWLs9VNwxdNyCSX/i4KlTecxFnFbng5lucLYjGUnqgJkDpZolFVaFVjmnRu
iy0njYO6JinNSga5O8T0t41EVJRNw0+5wxWI9siLVnHoJLri629ylMNCi4qv5sBI
qUc+mXmivqezKRbpevg+a81Xy+HWhyllsad6mjZOnNFFwMrl3+9OnHlW+iLhY2hm
MM1AmmWshbVSpty0y08r+k75btMxiofBW/iwizc23JTemmK2baKF+PcPIPnZSZr7
6PC+krzU886z3UOeBBUmSveqBDxchrbBCFvNQB+U9qE/MxFZpq1IjY94HERSDO5l
QfBqSgfaCYAemXu21fLCQCAIUWICFCGMCrWmbOV3IpL1E+BIHoSTRBbDn1j8o2op
bKMnxna7EVSWjMoBDJBZ47O5lHiiC68mE0Jwk2qoUw0hCf/Tbz3+tZ319XuA8tWu
tfbsvr7hDsMLJSJcHti8Yh6iarkdTPy/7y+D6NgPasSHfBrFuT7RQKFGs4OkRoxq
X01pkKrwi1pVALortTGMlQ3vlxyAYn0HMg7NoC0+qb3ktzKMUnnt6cqloS6vVLZa
NIhBfH8bLr41UaZkPGDXHbPDcxZ8uQiWMTU1xoYGaXfmuOzw1hocm1ZGGaQI4eaQ
nOk1T4QbHykQHM9zQptsJAjTcxtt1uY8Xrq8PqgLbEX9uXzbJt9BXMLWSx87avtJ
s/CY+nnot76OFLyOWsDXRKmI12PvaGVT9iBt4DtCnZBlwnliHGUWnFXMKGMZtkQ7
T9ffPyK+j9nLqrbWuxk+0b93xc/qG3W7wtShX8EmkjBkSXf1aDs4Q88dyQ36BDUS
md1XipYSFgfykNafA3Vb+f78pFbz/kShHvcH5c8/v+cfcezHah9zelHGhLF1J8kD
hHCsF9TOCr2LZrg0GTzWsAZ0RdD4K5CN/nEjkC+E17r1Mj28u6UWOvadMtBGYQyK
G49gr7g8U/5NhQeWIK2rVfAa8jPelSbjB9wyP/HUqdqJD1jiGNuFBNQhbwr4SMNM
VoPs7Pqj6lEyC0wtC5FSdbWilALmOtavvN40oMd8gx6i/SLE/fkETxloGdDHh2+y
WMPcUGKcG7MFJHT2Av7NSiZQ7p5w3GeANlizSwwfYsJMhwmoRt1cwIgmiW7F+BPP
03ZVP7fHu6m3aZigOITauhZ7ZsauYAYBJJGRuZLkJJyjzLdiJliqezdJAUv7fvB7
hDRTiIgJAoUw0ir46y3ldxC4P8Y949CK9Mn+qCbY57qYSZjR9HjBYVgRkPHwJJew
vnRLWi6CRXxsgpGMZ7BufIo+DvjSpYCrI1nX2WA2z0Tiz+vxvu7f9Nuy467GdyLp
tDMlhC2U+Nvw3lKq6DRh5tKuH3dXjUR3yxuY3OCFBQ3ydApKXGSltAYhjzSRXrhz
eH+ufjY8VpUIlf7+0yQ4DUlq/GHXJCjcw82vnLkMP5gck2+ejN+UVszFzfWNnvim
d5V7VS0vSGmfcDR7nmuArrbsEGbQEajJzWdupwDykmDhgyXd1bf6LF37is2X50UW
wqTtOKrpUyLLnL6hK6UZVTTtSPOFQeok5hS8jH54KnhB3u38JITwjsih6/c9t3w0
/P03B8m5eIgPHMVo5jwBrss8HLk8Iy09qHlIZnEiWtLme+LfazSTssU++hsW3PpQ
9F40FW1DqSurl0MWpSO2LUyrmjMd/9O4J+iTHvXk7+fZ8qBUpOROeqBpyIJH1czL
umxO/zloUDnFziR+0DGlvXKvXCbYU40JkoJ82ofApXgOsEbXxvdMXjsz1SjBZ1QT
nBAdx0kSkm87CTg4YT1BrsUsKj75c690Z3Y3w9xeOyYXj0QFuj7A5gfAlsv114IO
C4uTJqABK4s1/KyPwXvawfIdp61lisudtsq1CB4h0Wm3mQ21KUIknM897LLme2we
NvrsvX8eM+Nw5m17Th169d+t3C6RPXbyi0WolEM4g2n+Q8eRFw0BPzwnFXS+6kK6
GWhte6GlULH0bBBp0BxfjBU1GCgErFKgar7Ehon31d6YKnJy2xgBJQTfF+4Hs6KF
vpkpnqj+LDfKhOgTWbb+7Op5y/mVZIrBvsfJntb00N74RPHPrmRBBjgxCSYetuTh
awqyWj/6+9O13+0ScokDgx1nsCmVVS1TN8OZmVvKZNhSgn7cdq48PP50GrLJ2h4L
gsIxmNOkrpAXsvNX9pRvkl4j/Yt+fbM6iSYv0nVVbkBFlMaoV/8mYy9Cz3CCbO7t
+CfEWUn2KfbVWaonJqY1R9keT9GQERv4O9AsxS92nky81pXT20VXQeH2ipiTD2rK
Cfk2rcR253GeTpsKs+pWt9jbDUXcn3JMnUhjlr26z6LR2vpnUetexqSQgoLgV3tj
jY4QSBLMZ0GfVcpCs3+EOTx1mAOOXHjpWd11Jw3oT/W202/4vy6DPyPsHd9N9zbs
9YUS06OlA4Ivnyu/35YYzUkDrG8uBEaJ1QAnNowrU/qUGecs32s2ABUtT3MPk6p9
EVIAzGtJhs9NRXskKdf+m3ENEsmGWrOzQPaDo0WO8vD5wgjHuoPN8uRhsNzugL1b
FEVS/BsU6w7yHOtvnmN3c6mCnygxpt5HOPwZR5fCdYIBFiURrt9mLwNx0Y1Xyugo
zvDiESpL3BSzdHmZPx0FHFTTqzjk7iZW3BxM1foa23vPgr+DGjInidj8ogEn3KX6
2ZqpAdRok5ObRdCuBu06U2U9ES4rMCBDiUjGSYHSytA6/xMJ0oNVwMnQo+a5VgTO
HE3oIkZYQo+uNw072vwk5PIBp9nk2cW1uwSOgochrZ7/hiY8f+WQj4CeZPPAa5Mb
RZEGbgIYPNzuD8JOgMUBIuyb/3EeVk1rDMCz1QZBFeTER6T58CJ6n7vy2V8uS7wY
QXhiTJNOmKp40zcLPLyD4Bpea3zR7y1YxJNatzcQfrVYLJ/5c3UkjD5j+Ly0VRgh
vhY9h+FIoXJAGbxBcJsz2OSXDH83LARRVqdI0cJrBoafwbLH7kmqHXjRxb8bj3MF
0xJtrtDT7NRajIdBO2G7WnxXfV/tnZs4CK/r9ssikjlOspsE5+3J7Ym7r9TsQ3fb
kar9KHTWWkHy4p0fuIbf1py5XP3e8JxmcRN2zl0n0BDZltA8e3WcsXYhJ7y2/hlZ
8AT5+JBvp1ld5fc9cIaeQbSNUryOjqoFS8DpfNNnHisyPLTYy7ip72dl2vRKVIEN
Uk9/AgORdO94RkfPtlMuWXQMJjmn0++H4vWs8HDa1rflpaMkaX+mQtcEIfLJCLds
IENf+AdBjgsrlHrCgKSRuLagNhcDCb0/TucfC87t1NNzl9/jM+8IgDTQYK11l28S
9JXnWC0PXFpWBz9OsD4r6UCVtxdCrXd98coDpj/XYtV1jQzvP8NM3FqmgKimNsgL
odU7sbz0VmUvj0sIb3GzXz8stce0brlbrrbSMR9EfbHKa7Xy6Fq1m3QUNfz6h2rH
Fvdw5Xx/piuHKjosUcfnlVsj60RyquBGhwRVa1AnqB4eVPM2CwrgX30BRgcK5Xl2
1ohCQK1oA4IrSWZ5dA9iZ0ovco6wmM0xR26ax7q39jwdE0ZwkHN6uFOW+K7X4Liu
9sXF2bF2xjJdaWOjMJKSgGpCGvEKhAaS15IEMcsghMuHib8snfD3FmNWuyzv/8wT
8kw50FEzE6ESc9XmGLU45Iz4yQdIgpR/TLJH4ty4y+N/XMDT56wY7J0q/HK0CaD1
n7m3ahX5nB06RE3PhEsxvTEZY3EJlDMfIrV1k+0t1sih9xA0cqFIUjVeByzUPfIy
jzoTfzEpoP1DxZWmSJRSKwLvH5QhtI8mYaKz9rR5QoOxVGerht3WUwxHwsdr0PU1
EKvNsAhDLlvuoKWRGPVZmstZr7JTYspfA6d1BlhH+lpSStlSpdVufR/RX9PdaFW/
mN39LA2/t1n3+wNLmeGkBBicw1/H54EozYWcI/p1axxeTEEAsa+48ie0vVBM02X6
CxxGXOOxRbNBo2H2S4hZbCHDEkj66K2+7tZABmT34okJ6zQdU2nJL9n4wzRxe9jS
SO7X2LxlLjtC4UEpKGyj0moRTZzbnI0DTz9PfZsnxT+9My2QjtFwF/Mt9Tc9jP5Z
yeRBDayFVPWry56fBZLQPZg5ZNrVIITdi90GiXvOv6yKj4e9xz/lRtbMldmbt+tA
Y4NF/wTACmLGxhxM2L/iMi/GcGiANl3EyckPy+pF5plqDRPmA4z9CCb2WYtpkUB7
xhQgfXUUgoA9y+edg8dk6hAPaeEtrrc6agQYFtNy5DKdQLde34Bx4h3TzycOfsY7
JKXF52vJRGd9j+S9+vEbZHjYivVYz/Aii60kaOgfQcVc4EoQZzvOQeNeg2eLTRqS
UvQPzJ45oNN8773J47ZGRjlduLS2SdYeYpGmjgleLXBSmZVopQ1PUofICbnUpckX
CQMiG/zhu6mbcYsgHV7oKImccTIn5FA75Iw2FH/sdKa0KhUM0ulJ6o+DnrwnmIPt
+Qg3yO6AMKpyUyQZBn6zHRlN+cLir3cQG2svGASUYdSWuqQ2s9VR2txUiHcgyaz5
Lbiv0a09W814XiP8sUgBjjCXrL5/SblYgF+e3VqPRSnp8nrIrmOnmgrLiVtOIbP2
7TnOVxGBr3v9Pk26us1fbd9MG5L0Y1tNueJXUriz4GvHTuJwoysvvSqOy7SF75uG
gwn9QDFF/NKhE+KW3A6dDp19b5ti7+EgJ62Q7zT4l2LD8rwj47bu+ktIVESgUes+
1OqqyygFNyx8ApfbCNB8JrVri1mvDNBPIdg/wSIovGV1RmQuppCo5BM1WFOsDbZr
UW1dAwspEqiKWzxPIhmZorySHv0tsKG/+Afxda275pjybEVEpOwnMCMrKz8cnONZ
tWxEah3jGAEiOXLHhSYoHcrisnAhayZMzL30y7KoQ4a9GrzfD7+n3jAzuRvZqqp1
mKapcqws37m2IrYOe9tSbxr0i6HMxAvmVovEjrhsZFmeaE4p1VRToToVhO6SD9ZM
gz+DkiG0WZWfTwkJ66kMjZQrx0uKIN5YF3j4RXz6fQ0FVaBWYEQSqSUPEy/M+s2x
bCWzrxZ9ukUQLg/uREHRsxV/RDJlcYDltQlIPkZw9LJ3dIDKZzAOqeMPKEZqvbub
GLPsynvrmPBaTD/pkY73s1iRtlpW9rD8VfCDufzuhPin101+rAWbFDyxriXSWnZo
ZOJ/iqg6gPVGkunKgBLDGQMurMrFMvdemEMO9+rcHxOvnKNcbffP/rVpAcSk0wgH
XlAAdRw+cUk2P97fb2Zcvexjtk7J4kmmFX2zyej1Xuw3tiHTGvIddKjKO9VVhkFn
L/rwN7PuOTXcQX5l0mPyam+SHudgshv4uGwLx8TVB4w0n6Iz+D4RC6btjHnvAs4O
m4X4FnIufEeEdq+LzFIkF2YIpz4mcQkKMeTtb/6jBAkOhiC8FJZOJS+yx3jNlJHc
ngK8LXVzKeB6hxC3i55Mwz2IeLZvO6ScfbL8pKX3IPN0ruTR8y8NbA+AxOyENnil
7yL7rflUyXxDICWjjyY4KkUVzsgtJQ8QRZhZwyapIWMM0V265tX9jWXM7u4rJeLg
8b56tEN2CSyT4bTo9gNRmEGQxa3taG1/MJYY3sGq2j2cZqRFTQvQ9N2sTZ1SD76H
03L5KzDQTUvyx+DF791nTx/kZN2rcUCLbP9sGoM4riSGnA9QDiSewxRjiJrt0c0W
E635jETmeB8b9L7OAMYTmajj+IRLzqCG0wq5cMqWv9umeIrEVebm+c/88Xq3XQdI
467DB3XffiY85vU0z1ONINUPEGsvrwNZb0+zRcsd0tzOMPFGBu6bMS4kexEbrX/b
IQLklAjd/PBEQVUhADRsHn2aDxK/yL8HPjpL+b7aLHFe9FXyF+HV19pL0Aq2Do9t
tg6sKtD/vL6so0HsrBi6hfwSvZMfTfgQC1xaDt+DfiSWApccbFs8kr3y3Q2Hkxuf
D7otSBvLFkqxLTYhx4KSQ8TSXf0FEJwHzx1VRkYmLVkMHfF35F0bxXhG/Qpn/cxq
ijWBUiQZtVDjF8Rbe2PLW+1/4Ni3YTfLvuikzlIIhQAgpIYsC1Jwm4Rr8212liTj
dR7gKorN0ONPPZewClNlkikoZBpJNjXT44beasw/MVtwXSfDF7XVg/OTAk9qyEk/
AwObdF69ONiwm732k9mCns2ULjVdTNZxr5W4Cszulm02fp8JG5kwX1NnCOGPfJWp
cGohxfMt7CVO2qiqCB/XZoX4uSqbN+UcuZYIlHsOIAr9FZYyNNireYQOJDsZ31T9
fqNwE9YmjP5owRM+Z3skno1KaZOi1EXp7l8qT6DTvIIqIlwm73LYvbbr15tz6gr9
1GnWe5s5bw7z/YxsshZhwmqkeLrUi+x9wZ0ZSbllSb/Bxn9j4wLNVS2SlaIL6p1W
5sRTHNzKK//f9wmNmC8F4q7gaN3trMJn2erwRecjYcmyjrDTmcdqchwGihCIWd1P
m3GErgtnn9PvKvanv2ThhOwMby+YJGqKDrYkuBw7Gh9iecXE6y/9Ejkk1IgHkZKJ
y/3qGfzeOBnlYeBwqmOFyAMtAr3tuKxTmzLm1MX44VB8l175lSu0ocllry53D3Wm
9nCyjaDFc5PmapSn/QmydJrjlVACx7aJ/PASgdVORr+bDri3SqTCvi8dVwCPyYew
eRPxeOOdWtEs4coQ25miUx1JeuPoyN1vgldmBWz7jMvxQ5uFHBtszgDpJ1Iic74+
XTac3hjT/3mU/VZUMeWBufcRiZ8y4WMgzSclB6eRlwwPKzukpsgR38DuiB/n9Yer
295fkOAqYzDGkAuqnmZ4QcEVX63j4OIaso6Ji5/0UhJPTctypHt+ZDBq4ADEGpyb
k3riPbAFu0Ay3Oh5+tvltrMjiApHc/XUbZn8GYGGZH4mQo3uHe8IQNMfUOMN/tGI
EkAdGE0NxfVut3u0sSYiCr3b7y2oGz6Bl1pyXer9KUp1u4whxm2454sWE/Z0jnTs
Yhe+2b/IsFG9gSNU8OedVBjDZ5Cdl5UARCuqRZgGde5XtqcSaMea/2Oxi1yELYWz
QP6sgv448rYxtsm8TQ3+kn6DKkUZmjqmQWaGvVGbRkPtnBLuqsHN1IZM9Dg7gSCN
F1vBO4jQEADWW5rqCLG8YzPn8dLJ34dwLhbvgOihejmYX3/L0r+vxz+jPehKMccW
HUd8sNE/Vyk5U40c+HNQJXjDixJ80cqyvqrknsrP76NufMQzGlNu+wejqwSHDjgQ
DCfnrXWUCg5CDfiKd6H6zp05NsCpNwh6CHaMDO1OI95ygLPvkUoI1KqIuCBk+n06
mNgklJfmzLF6qUh1S77oY3yjx5fAl/pwaWaZFJ+kAgjjjJzA5smvHdfOA/mHgsKD
tpaGNF78R+O0Iso7uIC7pQAevGC3H0O6u/9LF92qW38E+OBG7MKVOqHwkYtPMOJt
xSqiiWbKNLF3crKqtlFtZHQcmATk90vBqwEPfhR+JZUu0zIQmx90HPDtCn42LsLC
MD2B0aNTBNOMdDzPIBsuw/Go+X/2hiE/yDZTmZy99EfzMSF6YgXjFjK/wuiAN0td
ddeGdyV3ZovBEo0mhHgpUbDT5/uNwL/1XGpiFG/ExgvW7jH21rCcgb1RA60XOQRf
zVybgce/2xTneYGvHHyoK+y46GI1pDtgVBIHpH8a0eG35ODzzTgf/m80wK3xznoN
Bpf9zDFL6EJzccgawzrjnRRQzokBE770oDFQxrkma9K1fbl/BZXt6fXArhqQZvun
DZNkm+nL+szL2vo8CBjgNG+uB49Z6CnP48wvdXKEUavkBUsrqFeNeLkYdhb7syMg
DvSEk+PSV/sX0wpX/eL1LAN2AEAGfbZ3VlAxyWGeQsYG3OlghkYrWgNxL7OEGGcQ
fVkNT8BqxvoPcecVUePrI85qlDqGDtZnvuCiPTKv3rUiotJkkVs+Sl7Fpom0wjI2
Ch4plTIRhD3MfBQ+ki2xwf8TWB3KfPnLnCjgpLeykgrO0hKBVPKYGUcXwjQv3DWw
nPWTg40xPjzXwy76QrQOC75oo0FuG5ty82IuaUTJUCen3NzY66DhUbyamcLTCQvj
MvgvuM/8Yc95cX0hzbG4AReCg9szU/B5HaVED6wI4CXN2ItJqIolYoWG01wdUfj2
6E6mNUadcNLJ6JlXAKaJ5csENL5k+vkAOAeE9WYp+YCR3UNDhRnuAVTtBAnajXh/
7eatpY0B5ykn1beFsxkg0jyYYFFiJGr8kDbqQrvisXuQ1i1qKwE67IhCw/QmNPbl
pCmRw2tDTrt1WZvCdEhSH+O/mQapmtTrzv8IOciZtdatabwOgccq7trLXieNP7VQ
yfxIqPlh9IGADoZR7IQBhJpMFkICZa1bXT6P4NpIrzqL2CWuPvTpcZu27rHH7yCG
lqmkfLqjl3bYA6aEk6fZgKjF+LDRHzHY0/t8WFdOPIKhvnAvgj8pEeNkQ9aucXOD
VfrvNyFpHhIdj0fhRkr7lfJ679d0epni4HESYUXBFthHye15WznQpNGmqmrBEO4m
FUnrFUVYbmU6coZZ7MbNo2doblHdlrgqC/b3zcgKorLDC2/NpJa1//PJp9knv/q1
CukjIFl8KNDJ2rzxh4FWnOKEd24EzTbWNQVg//qmxZl20clygxGDrPnmZb3EaLJZ
gHClx1y2VLM3VTB9r2jr6JaEXpCS8UfOHBPTs8fOjx+dWHBoJJOD6ntWTD2ICu7C
Ji98HVPS7Rp8FNIdqYIsJBFoF71/cPoaIZEdU/QT7AWNmDSEEz5K37sW2kI263RC
UFCBQau6aUwQroHTANGK8pUAtW7FWto7IFdpzySQTDfv+eQaONxy1ZYmLhxdqE7Q
fgD1pmCFcQFKq4mFwjSXCFWgJKbbQx9bLmk4Alpom7qhOkpKc/3f++JiWlzsRjcC
x5+8bpCp4Q27igVkLhx/BQkd2+fWAIPall7Vo5YLh/031bcq4OZfyDdS6jtH64Z8
Soq1l09cDDSlew5Tv8bSUlXxWVnCO0pCrUFlt62eEXN/RmE9J4JQnDTQ00LL20Xl
LJMCbbn88m4qEbSY6kS/W9/+muTwQbxWgYFd5SXnWurjzmvBIA4ci7DDy644YXer
nZl3AU7YBzN427O2MUkqxLM8dKlONK4lzsyNLluzjxB8ivbMTRJNL0VV4/CJSxav
g8AeP6y2T7ajCQ1Stmg+N/R/YqJosvfDuzTNkXYSSt+Qj+nHoz67v0PzedmAntDm
oEe9n2Cgv7z+JmZVUjuj77+F8YZK9MKOq2kE1ZecawH03alODxA3+Vc/E9QHq0gd
dsptXUt/X2oKufOGdIMiS6ZU0/ig88F1D+Qp6sJUKDuczjZgMD1/kj4Ug3kOH8Ou
U/50NX+VQPhiyjKSKBJ38z/vBJxjmfx95sItO/zFvpVPilFlqm/sJGPgk9cgO/Sn
VjWVUjIW0/mOQ1gN5Xp7SHFmSYlMBspezmxRNPtR9H5E9tmAcRkyWPxkVc4y4ai5
onNtZd+1D+5fbDsL8WekibvWNwgQRsLpnJDVNlstvAmCJIDh9vm/7kPyODEudrJT
xBtws0gwK5JAp7RA84S2on7xyMmAONrSDhvAF3wS6EbvNpo6oB8BDj8+uKlhsr1L
yMkwQkjp7EVSjgTuhOP7jtp4F2LFmEGWLNRg1vLBzpJ/4vnw0Iz4Wi2t0K3GSxeV
C9Mjl6pdlio1gwaicZ8yyzOyNaAkWDCwkdbxEg7yjSecb4E5VJ8a8hWVEuuipXhz
Kcvy/dMO+uv1s6izVbkjpneK6CgByXC0VlYQuRu8/hr4rWIFwxp4/aDK4cFxgjWF
MyqFm8N2XYgEkIXok4qaWxM+4wdeqdRxo//PngaVKP6z4At6VQ+YYFjBP4HwQRS3
EGN+E7+h/WPSc1vFLjKAHG0ufMyEfiEgZoPTuxgWmBiGjiYbKH9Z+9LjCHxWpUp5
S0TBKzuXvW5MdWH1Pc+4vVmE8ENNYxuq3g/nlGDBejcqwQxE8n6905Bwzjn8u3m0
nydhMMAyvDDkKZBNiDrOfHqeV398fSkdLxnr5DY3IxzKYsJQz0VRjQBa+yUq61lT
rh6r1oD7g/pLlXzujMRldA36EvY6OE80blZIpxEm0pCVMk0t1azq4Uk04E/P+PwL
sGeRvaQa7vkS38brxjPf+ay2yangD46WRuQOtYBzq1Pt0WiDiRfz8VwQB/51sCmW
uUYPTGIXVqOx7zBkGBGN7qI4WSjQmzIyyBq1ddZAx730UXtNDsR0dIPzzCV2Ydk8
6YhJk//swwV2pBJvGDLm9ntzaUzbZ0dHCe3jQF5nJ3/7DfAHwkRf+AeVVqc/Pc+8
ufSpWJB8YSr8bFqG5kFeetZsJDgkqIg32WNSPcfSLEkE3AXY0VZYgHDCiQzHe8Ja
DDmN5ZUq/6he3zuT/zwMvmzCwWbLQb/1yxeeIRLw011E6lYEmFV6iay/TQc3YVh0
o9J9TuBkOeTyamPA9S1wFW23Uy3J53Ph8uUEuX3OcmC6xdHcVWkzD0f+JetK3xdn
5LmPqiU0M+P8pUw6XAfYhqJbkSQLtALY1q/LtJat9vJNBfykmvSt0+o/ZzA57oR+
X5kRHIHGdBsKN904lZ8vW4BJUPCRnKMb4jLJu7TimhYqJpYiWAoTHgJ0m9djFxMc
aSXa6/1Oqm1WEM1bG8qTAkPciV/IZK69DZROkPCw3qE+ZY5MS5+WJCK7g4tnM4wb
XCAuVd9540cqAm4YjFmQDHBikLzhTviSlTL/K4A2LldKuNbXtQRNn6+i5jGrI8Lm
re+OwvG5a1ENNVNiGr6qv7eT8GEcUKJUI6m36Jtq6kwZbn0jGeWMR7XTKfSgxMMa
GPLVhcLfkOqBY+NMOg5bX+0escZA+xsV3jUTBZyOUJqKc5R0taLLmTipwjlXgq/k
CRI9YMyhKOdM0gN/tcehJoPxWNcn9j81ko8d2FecoZHLtYktR17XvHH8IgBAk8Q2
8K4UwR4Xafk4027WKQNxBj0eLD2FZO3G1sJjhZI1eYiTt8zytgSyQ4SiAqKyvqrd
0RAKm0eBuJHUdysUGNeZNRMTCnno2Im5sV2QsaPy1+Wh9y6fbhCA8vj1hoYGYAI1
QA+1s5rmoZzbCt8Yk7QAYwzxINxFckhNaFNgGg9xoAEuR8CX4HiFP6RmRmOvp94i
OeGzWYNgP9OltrdIFRPtrcEeV0aAW/S9ylU67fMPM/rIAIKlpts7qD9Eo1WwRUOu
DI+61oEZMYIt0uolub2U9rB1NK4oi60DPlovx5RTCXHEltlq//Bt2bAZgsYKH16r
Ng5bBu/Pu+PNcP/IR3s9JgWcP4wPhcAfHkITuFztoMBbnPd2jVtVuVKsR0QgJTEz
3tSnuMnnLVRndhToNKhoSca7lvBWDFqctGdp9pbEUuNF/RjXHSK5GcuPFvaMlSA0
cBqlg7mnYWvy0t4SgTUk4ZVeqt9/hr+W94q6FitWK9htJmSJX+DpWIQfzS0GJMK/
+MKmjX2KlpU1iEKtdshP+S2k0mK19K6Y/1FQG42uYsuH7K7WjMcepk7x4pauZYAB
XzZwBc6EXIA/sR0MQDNvWid4MGbMBAhLgz744Zx75g777rxH9lp/nR+EzW8JSTYx
e1XOhJcYknENKh6wlUifixWVuDP9mqAfsUYdlnlNc57jZvNuXnq76p20ZzVGHOBe
YLm1J7CihnYmtq2zxbWlHOm5L4xQmsQ5Lgy6rvrZAkhVNL9HGywa79j+K23RZLgo
KTSy2o36gLZmuxkLV0FAesmej2dmztsJaUzrp7/mpIwgj5a3UTmuApajUsYj2Wav
fdAmHZyk50+P4zr8EhK/CiNOxim8vOFDiBUiNAwZhJvZNFKGIvs1IVE8nlIxzYK5
/v3zRU/497sTozbJYwBjkK8IMNb2lOFGP5+sJIZz20ODmS34MGtANTl+8SRGdGHG
ard8PKgsreyJmdx5D95ZYug3b+BUUB2RTDnzdE29OZFB5YdZ0qgjvbUQ0YCNWbCa
TxLRiDnIddCusuyIQgmg5dScCSIAYJr7dEN0YzlwPSIjiwx0BmPMTdKmwjeJE0fF
KGl+S4GDB6fKITPsk13xJSdQA7QWD709uQUGOQrk9csQYXGO3VLdVcz5eUbpxq8o
O2YdcnEePgM5mZSDZFeenKJF4pLbTw16Q3wetUt/PdBZiTH5MqYCsj8q+dYtzPul
RzqHcmQtwVO9nS234TjRUKW2nMwYEZBn+bd2+ig2G8ZH4ns7LRr4sPtWnB+xoYbT
HrPkcg4MH6zbSQNIWcXsZVfUMx1SP0rxRsPyRTsQ2BZN//3tSE43M/5fJudALXx3
xOTa92Ck7rMAz/KInly9yUgD7brvGiJzO9ngIi9PuQ7tkQJkhoKuZOCaSdW8aQuJ
nQqDTjVWVkBOh10Po0EWMT6YwaQpbsW0oy7A6LBSI/qnMgAdTJaSFgLKnDf47BaE
mAq8HgfY7OqHVm95s9zNeJEjOue+5xZqnuj5KEoRIWYJzXF881gNRb498UzSqZa7
5xqm424VQXMDenwGpuTs7x6cfKFyWl3QzyOxBrrX7d0wRe4lLYV6szsQdgCrx4PH
Vz5egwdp0uHF/sfL2k8UCKsAAn6AOrBsxehr1W4b0fDQhniPpPOlZXvrujs5RA6B
5qzjF8ahWErWdSPVS7Bv9Rd5JIu5FAauPjOwwNzzujuN6iHZ5Hl5ysWOvugPXiv5
k0zQSQ/P6YmlPWK7WK4al9g75q+49USucCcddp31HeyHKH7FoiFrfuK+TFRlp1aL
Ghxu9UTctRNuxE2slEOm6b+I+EZfLSOO1xMkS4GZ0SfPtdhWaO9oUpeo3TpDNBmu
0vSpHDMYLIltV3zLqJKcjclLIYGTtrfFZ+Y8zhiRciHm1wHjshkuIVtC7m+VtsHX
YwQahzPcpKPpgKoUFBluFkPzDBZY8xiSeBtHHMjuQNcHHlnc9mfsrtgwr14et2Xo
1y3YL4dVLvOjEyhUwdz+oYVbu2mlzWXxBhfmS50pBNWytsdeOm1yLqLUFdRedEK2
X5KnPiMk0r78gpMzaf3GTXAoFNnvrP0wJTdSgdL10BTHhSy6GMJoiqpMc+NR38qL
QAoHPgb2RHE9thcWVJ0XEWQetc1Z1d7WCiyDyTiB0JcBeG+U7Mm1VDAdOz4aJtVO
aTtCOSnhYuw1E1OUtUDZ7kiMWQbXi05CcwQNiaeeg3S6LAgSNRH2J8xlQL75TpeD
ZPg/EEzr+zqJ6yRU68qYBOx0PSfKj/PDRE0R+pZPIWlUG74ZWd92WOtBjtJJvr/M
EhyWPTrtgTzH1EWLxp+YVV/LGpkZs0j+uiovYsiMHZWTSMP7CljgsgP+XpQyCVfK
Fa7f/CEC43sr5TFy3cMsmUQbKjxO0lgpXLbQ6qgq/8obI8N2MLKE0RR6A4Cc1yQU
qgj6wycilDuwZW+Gd+dztn+LSpF+bJ5TeLvEpHE4g89yVEMiDw9/NzfQQa71CGId
a2BL/760AcHcVWhzOGS/H2fJtatVdnZfyV2aPqLL0c6FXsnXfcUoQuO0Ll/hjQ2v
kvELnpcSvYr21Se3yi8Y2kY77J5BcY96xe9W7p2t4nYw39K54axJ3T0xACT4yO6j
Ad4r5/S5i1iZEp05K4Qpl3NZTnPYIpsK9OI7At06TEPyyy/T8U+/Y/wdymZDR37U
FLMDowK1enZ/RdkZPjrePaopH2GNBfMvR36CBkaynaXhtT78rEoinLAsJcl3ceIt
ilvZ8XDXEupD4vQwY5tpL69tjAyIIeSDzSMdkPHEcPiExu+SSUZb00xFd/cbtOAB
OTUUP2LJQ8uBIQ5sSm89Z5GzeU7eu1CpfjYxnSk64l5zSlnAyiNNCwJ2eOeuIJkl
j82TgSIO5IUuCw3G5S5cBJTGLsiTrGoK0T21gi1Vaz8ZWNpLrQIT9s81zL2RGsnr
lpayCBo7VSyYMxyEruS5w9PTbC1eMjko1HMBScf3hnbI24ZI/ziDVMZ95G9ZdBzF
NH7Kj/bAe5+inusfrc5Vo3vxePyMgQtsY3Zi/KuVMcATWYYikwa7mSJ5cKNYIXXi
3ZR9nMLpTh+emu5pbKEnlkMUMC/c2s2YSqiV4TyEXiGCTJeWngZ9NDQtBilPUW3f
2u9vU+RPsnOtnlpuO+BuYRcExuNOqOJgLO2icpCOb9vxFU4M9MzV4w1/ZGmMqiMH
t5/pG+hlEFrLgdU4H0o4z8DeBezbAvcieTQzC3Gh85XfK9XCDGhDE6QdUJXJ7vaw
bekETs7yWRoVQ2HQ7Aq4NTI8nAe6f6NcdqvWF1nTolkeS6IG116l48wPQeEXbSq+
i+MLjTYs0DjGoyhwxAjlGpuEbRBkeACT8f498eigRyaQFr8apJ66+PDLdhYrQ3ql
TKaHaj34ItsNDg2PnI3Lxl3a2dqdelLsdS6pD9wS0/zgGZaTyAF/tq2WC8AkTgLJ
2rMwOYx1AV3m8iV6b8eDZ+wpDvSWlBxsbdN46TPfEUWMnZJkB9ITggVtI6ZxGpby
pzzksKgNQ2hTkDFORgJHPOuMST10uLn+gnUQaSzEHKUI4g+iZyx5vug3w5Im+lnB
BwPWCDXLkTic8ZR2dozmPayILn6Bkm+DsmXAfAqyH3FKWr7D9/wYsJFB3jQiFfaw
nTOXT5jpEEfRfsQUieJostJtuGxUcFG6xZFVcb7oyJhQIkPHlD8sLLTF64S0v4Xz
kkDUwWGeNrUOap3Un59KlB/IqHuR69yNrHlmemKfCYVTIWChENgnZPASgHR9UVim
NTlBt6ZUtYrp42Qxcf373Xshayy0GsMDhW5HaMQP0rlHsrdZKUqTVzaTtetvCWqH
tSCwtC6KpdHqYOv/aHRT9Yf/5pnMELcRzk/iUDx7wVa+Bh31synhzIdPalmHfu8G
KFQlGlQ+6xqki0hQcrDWN/8zGwoyhVaqFZjMD/wEWHPnt9sJ2Y/nupthgl8cX12E
xbdfdyFfX0okoYHWbcCfr/YF+Dh/jqFpTYNkubvTzeeKQMWdLtfm8iJy+GvCDOuK
HZwqJNogzAb1eJWqKcFQJXgA7T20GByPutQbNCU5T8CuW1TZuCE2pbCpgJ2zOn5W
v/aPtuayL04KCN5hvAAm5yQZ9bveC013jl/MRFNH1TjlqdiTet8+60HCfUHpkr+D
uTtZJWcJBiKoX9nFYaIUGBqfyVu1evyYi/ava7Qq6gP0719WFHrKAkawlBuZ+ss+
CFyFI3DA6qsjrxfOeWc8NDC/ob1R99Y5P1AGDPYPIj4I+Hx/9uwGlgV+SF69ikhW
oNKh4pObQc7cWZ4RThivR2DIIqWZAeOPWhSuqXu5qQrELqCXpnXMDL1MkFeytsQJ
s7AA6BxWtxHoF0F0XRkbD+VYBHxG7WrDpLQgBZVO+IfzDn9ReqUzze8uM2259MhO
7caYD6lQYtNHMznwUq4PgZ2LUPG9uTGBZQPTh4OO0NJtc5qhiLjl6fGRGZOK8pnn
soUHOfJ1H8AAbSWXEnb9gJdYg33C7FtCGLhA4cSSZ7u/QX0rlRW5ptbb2NP7Zk81
vGkXm8KiHk51GK0t8JyoMxfXviA3xnBPnf0MAGQXgUp9YufKVv/JLpOfSKTF3bU6
3a4dAJ8DD4NiUzH7HKTymd1pYxZMSLw8Ygz1PoI1NjEoGcCN1G6J24ImJ9SBSvws
kEOasSn0S4XZYwzNXaJezRBwwuJBX+5MJNIlil5LefMUqv2DNA2quopb1ppJdqp0
b3sdCnCV+aZStycEs7xQB5SLEDCXU1OAp/uYAceTw5KPHrqjcQ5iBB4mV2iDHEvO
muxcKQ9QJLMM3lghNhoxqzuaWGIDjsSlOSO2HAJ0kcu2KBramPbP6MaRSVYx4U3Y
mXairvszfkNYSuUPzMrS36Ux89ojomEdX9w/oRDkmh0oGlxcSW455mZxhAxwYzqf
S4xzl4a4IM1+ctQN+QBP/Vqijmg+ggtrqNof/Ry7q3vOj/rFa2UPJ7xK9P/XLF5g
wgSgbWplpFEWcZjKhNZEn43OHx5a9u8d/aIeg/m0ZG2yDc/y/OOhq6vzZV5AdJHE
EuGt4kq1M7eb4npwLS+jsJyJRWpYnq0zkz4aO/toMl0mS59REbxWHicHHy4/8aff
h7hboh6zNvwyX3zuS+89MwuH1Fr92SnaPNP/ydLmKdtp6Gb3Go/dp1M7EOj9qP8w
bVisYSAjrYAb04EClVUPjuPu1zj087hDci2Fqy94XuvkY0svZtjT/KsuPPWiTmru
Zgh2mx6kDyFnwA8C2zmN9mgWimsDi7FyQ4vy/bmx4wmDRUu5fxW0QHioJduPRktr
02Xxu82dxM7Q0M9hVfrWLv75VgahjtEvvQpgFkHpFXFmRsA7s/vkDbjMrZ9Hg5HN
6gZlS8qKrZRO6purzXgw62FqFORyC0hFj9N+VCZPyqCSc9rPhAuAfTcGADKQ2LKT
7JYx57K/juPpCJOIUdPvAzG/KhyRdl1W5loUn+tLAl8ngSyJ/xC0HHX3IVm6PYAv
cr98y6x0/tCBJZTpqqs8dr2IqfsPRYf7DfIo/rYl8BTPgouHyb4xVcrzZmmCKdCj
UIHXunJxS2WZvFUSrmJYqKcONA5L0vAt1iiH/O3ImEuFfnj3rhUC7QrnTTNDbcZt
uTK1YwZeGx19unxPn3k4JTYIjqooL7F4E5XuQ47cU34egJtc+mSPbhy+/WEt+svh
BcPCvOpGqE92jk/aGAYm9GoNxGmNCGpNx77qAKM9k5IazTLi9RKJ4PFxk6vzRYfl
fz3hSn4Jeftg1Yl8c3c/Y05fk6AJHYjHiOP0LcypzjKa59KdULtHKY3bEDLTzbSO
Vp2TTu193LR0DtUlk0Y5M+TLXPwGvgxaS/qI6GXQeMT/dKJ6yWLIbrDJi1iR5mqx
yC8/9iLH51zyRkPp17muQI/Q0S4MBIs3uyMeKKr2Lt4RCuO2D4LvXE+KuGfBKWyz
Q6l+FfSHz8Y4CmlXLqoUbzloDJRmxZ7vccX357clw+WJ1SWyTniRaaKRNKcFdOV7
8vh0wLNJ6/jMnkHG7RqHe3PZJDYpC3cduzjBkTmhURL67aW9UBRwjvnsynsubErS
aQcxXtqrfOb+PNDaIZiVxaBVV+x2MmqAEDns4YcHqmiwdWR16UuBqfJi6Urk2sKC
nCJ8CF2XdJ1vdA65tVB82gOG402O8JHFLT2kW1/fB1dxmH6wH1MENb8xmTms2oY/
IijIzzpzAYOYTO4teas3rsPAle/cQC4NFk63Un2fJfY6jrdctiEIo/fSBDgqLQTZ
bSCw7mjqBDBO0AXrJTz5MOVO/i00ntvLi/3S3BWkBVQjIPZj2vVHn8W8/CkBsp0x
sno+2FON4up32JOh2Yd4eOYMhlBIcoirg3RsNRe5W5eAvNvhvgFcKQbyPUpkXhYi
QeZAbuTElUJ2vSGFwtWJHuRuAknMwB9x7z2P5jIFMk4JpVIKWNrdCf+Wz96rGcDM
ImCdf/5qFU/tXAqLMg3Gz0WBzj3uCDA8yy3AylzlgQNdgAkFKAlAMoXuHb1a1dzw
dzcm9toUTmU4ERj+vD7/xTEKuA574pDKhjnEWjYveGKvMvHI4/GXzIHY+ELMkv8J
BJ4PB3amYtm41Z72jGtrhqHCCYCGfdKrVvLpKtQnoUgxD+qnPn9j0aE0lr3MmTsU
n59N0KJ8YNYVywusUGSmh7TmYe2EjO9Os7Si975bmVidFY3s5tAU4duf1L/VY20Z
NstkY4k5JbTzmWyIiWBetLO6inC9PmuESsfrQJ0KGWDK1bgURbvJEgKXKy4AzCVJ
PRl8NJ1yn9hjmq8sJ5uSfrgPaNoeLZ11AmW5bf23RZfnDOoG9P89kWIYJMniksSy
kCaDKYjlz09ptPMn3J4GrAKCJNe37nyJd6pfOgJ1SAMVEf8D01WjrI4XXluwGIVC
1YEtI++7ksuCaaTYI1PiJRhwfAxkSMsc87B6Et/nE+yRZkK853kINftlOQK0ZWsU
vIrOmhyHCZRFxq1JP9zmeopUtO1KCTrt1q1M5KWn1dxxs2UHF0EolSRf1uXf587Z
xyBuzDXF8RpStvayvAI6x2vFieR0HNuba3gqYuu6uGgAYyZmz+PzabWrI5qQYHfx
DgHuJg+pfo35iXriIOtcdyYyjRa+LRT5K1BP6k4LmBWY5Z5A8KE2rwEI6hkv/ZtL
mIK+FhYIGVRys90GKYqgnZ5/Z6QYR2CU7rWRHwo04xSh94t12ULGU/K7N6mhIYO5
KKhh05gRqFtsJn/RrXVQ9uApjalrgzzc9ra6QXlcLNi/YtYFgGCKECpza/1ZdjqG
T/BbmvgTCMcHa6NiBMxsNBDaRV5BSFYzCaCmfunCFy7PE48mIuOyvqht6aPcFNFy
FctPx7PI8MS2TrgUMFSij/62CUvPKBzJuhBBoGvBMutJWIJRsmv1ufZn9yAhJvZD
V4RKCD5xf/hzzw9uCzXE5PWH3vFlI+sTz54oKNckUP6bPL86u/g75aHsihBUH6sG
LdW8b8NrlNGEHD7iYBH5Eikszq1DDYWU+Nu7Nl6DAxnBezNAeM3fqWDuN6NI5/M9
bVOMJtvSmlZuD4kyzySCQJxgiDOtq1UsKrWW2C3EhWo7t8odiSLUEMjcGVTnHN9J
QmBLH8Fwc3nx/9A90txXkgxUYzR+baNyLm+P0hdMqAMK7DBtNOkxB8sQ9yAAPtAH
2rvJip8E4M4hYkUNk4eN7WtavVnU5Q2MiDH8n8Tlqc3e0Qym1JtrIOLETLcCePnt
/LHGS2ygTGIxMvdpdhn0p2Y5ICiENgfqeJhC27j0ditPxLVEpLZHluGHMXLVeQx8
EgF8aIIJetOuTkYf5KefDzLGuvi5Uz9jVGfVvlJoPD+dWaN1bjoT88SB+o5chxrU
dmnZJC33W+O5Xnt2EsSf2zi66woev7WYDFzpL3P0hSAGSpmdwJqdKTJLu/GEaoui
jRUUx7VjcHU8aZR+XEublEO/W20pTqPpSqlZ4fSOFWs1Ss3QjCIxI1nFYkQ+yKoh
74zhHipTVZ+9lddS+qY7+dfnP0xJRRg+cxv6AzjG4VTYUrYbE/C5mQ6KcA5lv0dJ
oPmjnCKSz78YE9ToKuoT1heJdM58JamNHcDok7+CCMaKKAfKdWWr02rRzyH7tHmX
f4pZl2whSSEwps8ZRpL0/fGdC7Y4Gt8DkfPSEmReXUQg96f7DSewXTokcEdVvIqn
tDdNxkvigTNUk00fWaMAQUKRbjc13uySJrAbhD2KxP6Fq9RN7Xl7J3MD62CdPCi1
ORarNnDVBnYj2K7bPZU8Xc46TZjVebaCMWMlvKJpYmlk/G9CSqIrGWxjG4N3Qq7i
jWze7gjqQ2Y3U0SrHpvP8QjHF6E5c5vwDgsoPOYQ4lZZbtbCnUiF2+/O7jiJeMCO
uhLkogioeW2+E+skveyHVFdQqgg+r9EItCfCRRWHZBS2NYcRpjBYZFnmLmnsEF1V
r8CgDaW8gt/muiB7f5g0S+LZXESn6cyf78RYQsQqj1L6BYR3PEp9KKo2XvcN+GyL
xStIbFRiP78LjqdprOMch9Wo2eEG4mS0YZTYwLlyKYXVpK1HjZnbl25r4rihztjy
oOKpq1DwsYKusyn4Ch3GjaO4Wz9CFOU4gXiQMS/HxF+z9usLyO4Ou8TNkYaoq/vM
3QrR6bx4z2r/7/OSvxNww11sXiwsdlTdl5/+QHgJyMgA9bbeLw5lSMWi+y/8xeLb
meao8lPgEwW9vIXIo7rvOw8X6OsWqCpHsZ5lSK9ZMLHv0eykfGi62oD90Dys+uEy
mO/cIOm1x8AncITLzwX3JqKxqXALTtZW3ceiKTtprYgjOHDZGTnhly+uZTtQ8p6d
fOUxKyuToonGrSSQku/Gw5bkDDQknnpCo2n6K4k+2dQ8aYun+sx5g67SL0b7MREt
dfr90fuhYOhRjTWklDntJU9LCca9alKIeoOFO3XAdbxTtH6zpMZPXOTbbiVbHbR4
CtB7g6EVMV7SJDqLx1aODn+wlZQXyMXjWg+Hi0i56M7mnqC27FNcK7+wbyKcZ90a
svGmejLLugi2aIEfjImaAO6Hl2eVItVpIhwmtnK+CBiVEzoervPMZkm0NPxWL5rJ
tiQp68jAXz2rEUQAJxWL2lcAOT5HojxtPievgHtTtWNiPpx8i9SAgjBUDMmz3m3u
BnofwKEukZZ97IAd+HkBXJz9VPmni85QeoqUTc3n91UcCzsft4Pg6KRkfe8Xk+Oi
wCf6U3ExGljEVrherrwW+RgK7VeazHZGRWByuyvMNO8pXENrt1Fe1VDZmU+2Jm+3
LTD7su/LGhT6mq6GlxRQhe2QiwsJCr3wfISRRDO/kidHM9IwNw7KLmnUpVHouUE7
4ANg8W3BUhGpRg05LsVe2x4wLh3gKAKzxU93fCD1RSK1gvwyzGGlee3aw56ZKsNi
8aZvj2E16cwahVptgVP5418pboS5XTmnmaxGreawr0GOWT37DJyFGq0RL8rj06F3
C6IfJsdMyquHDGH4W8GMc8qiBflmTAWTueqI0W6rFsn9lEL8g6MFdoBnKjkFxU0T
e7e+oOG6BL4Xwfhqnezg2X5FKkpaljtEttgIG5/lvaW/R6yV6WBmOzjQ1OSUh3Dy
wfId8nwKzIo0HJSFs5EFwIZK9tnyvtgtLNLxseoroLHzRmR3iO9whB4dSoZgMUSz
C6WDUSvFzIWvHBSz62bs+lViVYrL8xeTCafr8KETn1MtI5aYE4EsuavwxItwfplA
dqXrj2jC1PTGcTXLDPEAQ5Q0cfAOlZUUPiD62HJqw2dHgipuFXzh4srmCXgyEeYr
R854XOi4nrcnmbM90ZuYB49PF2fPdqDkr/TqiWI3ixymX6Hd39PZcumc0mhdpsVA
klyXmlQF77KvFW2KgS/D/KYglVCI/1S/6Mdm3oFgcI4nAemsHV5BiFqP8xMPpVZg
BDs0izuorHrj8Yt5FbMbKrzuZk1jwze8jpyD2AOzvdpT0va5SlCpv1/SZB/9Vybc
DQAO+aUNvO6YNDuwDErLRxTxMqO+qwJonNKqAbNB6upkxhevN+4i1zI6aLhDCl/j
KvV35ckpX7UsieCnMx8mt+o91MMelG9mEbXSSml+xWqvqf1Xv9tVhos+lIJ7MOZ7
bf8GA7IOfcAn8Cn4uLpU8o3vf3EvQ3+Dy0Ze62yasMJmnEfDifjIYWouxDufMfQD
5vvkH9ydR6Gr50Jduak0Yz5UnkAfHKaDnl8HJ4LKQTZhv8uCA0aFX7rEj4X/0LwQ
k1DI5b17pP5P2mdnxZUeVTJCeiQnjC64KEHLZ5kAmb3bO2JrHY4zYRp7RPksuIIy
26Zl09hyNZr7zP1EQ6bE6HbVaUCZvy6PlCNF1pbaYK/Xi0Aozvf2X6jnFYQF3MiD
ojgkCZe9AqzCSa14bEgbbZmaZyIAIMXp/FezsmZhqbUZ7zHxsm6hQPWSNCu9F2VT
0Op1cTRwBYAb4F7TzTf67oo0ab52QBtnIdV2PsrPxspJYKlUSsdSOaqTRkRykz1a
7r0bnf0Ounu8if4H3b6DF2EYxPzVlqTEuLYedXq86poPb42mLDzXX49oQpIsB/0f
gCo5X5NZM5y7VmUiu3jqpTkWtMqDMhEJAMdQLglvPk98eNcr3Caen8tuzdDOYR8N
cwBmta0LWc73aE3Mr8pUzW3EK3BoNHJNAjMgyCPfsIC2bB06ZY9c4jOtkJT23tv2
E/9rwwYLu2EHpcBVs4lfQ1N3Qj7bkPk9Sdtas7gCxWzBvyv3+7GlVtsVxkgVdS+S
bAJ9KhqsqcSVE6OwyXQL/ccAgpKALeB+srTiEmNgU3CfVzwZt1dno0s3T7/ZHp4u
MmAm8IKUTY+/JlvXRqFFg1qCYy31nHeh93+sqruBKmcIdHqF8xtBGvDprtOjgR8H
SpztI1T1VKJZOon/wn0ZaqbGyY6P5fnpqHsRFBQam8ixL9mAFkO8F8/QtFK4JG9d
zUUI93Vb/hWg6dUl1i2dZC22GLLuxF+5NrZBLrquvkycHevUDUVcu+rET/FGgER6
igewMHCo+f7eqmHKyQosZ8D/8oQLyusA4Ik8xgwVi4fTHEvEMoKtb+qlrRP37iaG
NDvtzEm68AIyP+dT7BkAiJcw6/4/jWetYHCb2Mc8JblIaxFBojM8n3wusNXY5Bum
wRi7u7f0tcy6hfr/Q+Y8cF8wZ0IHeLFLHtW+mDbVtPhccLtdELMOu5KIJ8wJddHc
axvcAWbXlXuw21DmmzTxng8thKbW5yMxpnjUmJ8itQ2dT4YDUFxG86ftGRS6XHnZ
XczPOCXHk3sIVhQoK3i/GAsLdse+DrvFJM6BcB2EDrtGgxk+tk00oZsa/jWNUKRE
l40JWzmnTtW8nIhcfhjPiI7671+OONqtMu62rz7Fzs1m3GMUcTHkGuDtwntm29/6
uwmalPYmK+T9cU6lUzPO5S70lOus2Ym0B4Y+L9VQNwIOeJCDMAVZ7HIsygEXe4gK
KyAPBe0zH9e4KAJdGPL7fpoTGLMaQTS+UGYzks+H7j+Lt8VJEDRHXBtEn6CDwjkw
AonE0B+kIJvvXvYXHI8DJVDs+S4PhvPQlavjPt45FZBBREB2m+3f4u210gbmdLk6
wmRwhsC1RIqKHGzY1GBAbABFV9ZCvN4YnQlWzDEbqlqdPyAMbK1/hfggK9Sr95eg
HBVsPVCjpO5r39dX6PhxDkDs6T/mguzFowksG5pxX6Xen7kyHiC/x9dl7pdgnX3G
F+0gKkFdfjJwhRFwHkjQZv7yqs/CPRFPul8zvMV3xAXcyNecEnaVEKNmk69fhojC
IaICLEBLNbzrp4LXVLIakT5LQVAfZvdpfJQHdbNQhRW9M9pNOzfgT5xOZBqqZ1zX
8lNvY+lmMkb4LOCbSoEiPOVngnxDKApLYXVNlOkqd0bwK9AgtNlXa62YAFgYdFW2
B/kDQJYCCanIotsE2XdsmfUp9E6btzcKrphg0avyR5cFZeg1vOuV3H3sUkR97GdS
eUW8sF2qNjmjakX3vMjaO69a8PvvNhkSp7t3xzql4leftYMIQAHy/0iA6cTK/YQh
MBJJaGPpTnDmKToSWuQMiqA23jcLfLsZCGyIb0DRrdnJ3PFirr4uZ/abLNlwagh4
4zAhX+PH+hn+OpPKlYN+J/WDy+atIQWwQ5N5e60xRjp+qlmTTi0AF8frosnL0aDN
/y/DwBPVFYrXeaR3IWEyvwqB24DMrz0ixefRIin5gagNrdMwacy8yUgNc8dA+FJl
IFxfVFsT0wi3DkrMyYx5aq7WEQh47/z9m3mvFKljWLi1WRFIYWEzNL9tGEdm3fA+
LcahslJCQ5Ou2PVi+lOq0T+bwQG2RSvqn7aQKlo9VR7HElYWqaKvf+380g6E3tKu
nh3AqscpCvYmHDvZ9z7w2W38Eja8X/dKSYms9nsD2tHHRpr5Y66hpQjFvyITCOZV
gZpb9hUEuwwOfm92dFhd0q/0zT3QPnVl/spqHkY2CU+hnOaZ03IbdzjifDJIkVEs
ytFzBgXKA/LVcWZihc+iljDqNPXNUOsOL1foOKznSR465cH6xlsUFF1grrvSRv6O
8/yGEW1c5Ten0KokNjr/E+hkM2rBDmUN+osCwddQaYYfDBqQ8pUpCqxVsnZ9+wu5
1rNNiZvVQKMgkLRSS3ZvwdbxppSbHHWWYdtj8jzsDbsiLY3IJe0bJYuoBLZxC9uc
fvEz5gqMoCJer8RPT7Yy5rOByXwna06JHgwAEHvJFcDY9LnaBRPjLv1hFu59Vse2
qw7NCQ4SZfiKlm4a5zCep0NtNpimOSykzWQWsHTBTDI8G7LNbi/INsSWKeuPuMBH
eWtq40VOwLqaCRxSVq8t1dF5OBY62HKi2g2ngtACvLhLH0g2gN2fojY26Vzfh/Ex
0VHmN9usR8LSNlrDuMcMxGfii7tQHM7mHY5s4K+z28+2Ns6kSOix3Dyqe/T0pl2T
ZLhQZS7x+NRxM0CEBSaC5yR2bO12YuLVXqY5aVhdvPwnOD3iaGn0DYW+gLyzePc/
Z7qzY1QG+DwPWfTwlfANNKo33gAUq6PgYMsqHcwRacht/JrWb4vMJDBpu4Q5uCQ6
AQQW0IiyJe1tVjpl4f2c2wIvGI3M8825tVf7HMGg63OZ22mHa1K33o2XSkny84q7
60w3WvkQsH5GDkL6xXf8cKD8pZgc3wqgtbmI67KV2XZwravBMSgKPiQYVNDtNSLd
Te8ggTtEbKkBFvXx67rgvIYh96L1LLu9ABn045Oj+4YLLV1ees+RpUKwKq1YJRvI
bSrQG/fyMQ9fi9aMsnNGujqVVTE1z7V4LNnhmTA+oqiQMT08DIGyOTgVv3zagebv
lvN+88NN8LXDsq3ePWhh2sri7tWUqYHYhr9q/8Wuhj5OaV20Ghwm4NnnLPL0iMQt
ROHiEzputl6Jmg1o4V1/5Hj8x+W2XjKk+QRstoEvf5NUyGlWLL7XWX1DFA+HdPhu
jzrqJNHKaZpa3fYSDEI6pRvsxRUNVjieakTgQzOCmy6LUVo7ua1jRk7bSMy0gxdX
oHYWjU1pwNzNBWn7PANM5LgxTkc+WvQ9pcFg1l90IPZ9CgoWM8yIzLcGnmWLctAp
k/mu8aQqwYEQOo2FVL9LaGg9PN2VIWKlIWbUFczKrZns8xg/Wvoz9CprpALCnfDl
60JbbKrIhSKY3OiRyL7z0+owqr4yd6Wlzq1GXB8LKMjSyNaSejXY8xcHcodkvs6x
lsEGWRrAIyemcjYAmZ33GoCGkHNsR+u62hi2BZuFsRqUApvNANtjGgaPgbISKJah
nhf66v6WOsWIqP1XBg8yFpxTc/ZEUU7X3W2BrFYTWQd13CruKkztMHA8/2VWFnMM
1HqrLekmin7B2Ppoa0yhiR9nZ2h2KowO0pAmdpBNxK0D+AKcMs3tARC33SNdT1oB
j2N1/++UaCR5isAZusL3Dt1rue5CHBWdVanTfjr99qOHDxrQ01mzQCNfMqNsO1mj
wvVq8tEiPv9I6pC+XgFt94PEM7VAGCmqlXN+Nw5CaVlbxfpSkI/f9i8RAjwpdJrC
oEWdUniQG92389BBFtdJ89gb4IO0cLMyNs+Xsvqt9BgnVg/Ahk869u2F1XXe4Rlg
GFNvR013np3N4NtTe/s/2t3YGfMyRFfsfjFytKbKHhGC7LApDi0jfiH+2h6/2Rdz
EPgmQGwXimyv6E3ikVWMyv8Xce6CjtS+pFacvW84KycoixvAEp9jfBiFALT4SxHw
bkDGOXtHI45ya19jVJ3KPkyVzTuHx10RHn58emxy8sX48x7X2dohOPMEq1EYVyeA
S+K7BLReJS8j/YV37o/TDZAXElxc3k0CXz8J2MFJ/HawslhbpRT2/1RSVnkpPpQU
vxucAcxOqChchA9k/+ICvAVqNKwJkmQky397Oi/f+2gQqyVrlmsIvk25Ae1ky6fy
CH5RWraxCr+QkzIar1ptPX7+Va1TEh/ISlwlLXgIMpLLuOzFmw9RhF8ubHWR5KXD
n1DCkS/jO3nmYvPFxz991l3XaH9gFlmsz8wTKTRwvyePt8CS4lGxxi6qTce2Ih4S
fi2IzasoGoMp8Yko0LIl+HmPwo60XojwDNDCvXzrZMopYUPD97bZuxcequhGOUJt
K2yoKhSoIZrTIv6jFpanXSgruS6WNGqwLRK/rv8YVA36NI4KmIKYKx5fNKJy1o3N
vno8Ao9m3TDKiYioUikhVa42hqRZ3kEQXpPemEB0bLDSMTWQGn6K266tHLTYJNgU
w3zc+QqH5s8A0r9OVe6A43/J5nB7JQ9eboDHN4o9GN01VT0IGUVuwugsTAvduObN
ghtXUPhfsM6KrSGJ888yEtdOaeLN790OZ/OQnm9h/MeNoMcNa88f/XtLYG/koQlH
fBtdA8qKCbA+HumErETG4ePTM4FHrMqgWLRUh1dIt2ccZK/biMOoWIX5Kg4IBusw
Zi8Agouoi0GRuHhYdPrkR97UZrBIUyEKqq0elrP8y07E9u9STDh9cF/O0V+xu/Vf
XyRPLnoHNEkyVnrDWKC7yhtdfQxCg+/nN6pRCEcdRXrQy1HvvLU57zj1PJDbsrR1
ID+2I2CcbYoIP+sp7EyvGpQDOLaRkJPugO5zdx98fibEYE6iZCWw8rVHk/5Yo5WH
U12oDVz4T+6Tbacc6jOq/1EfyWbLoRmz4t9GvWD44yuiFEIdk+0edZTcFJi0iTs4
UlVMxk9boohlM0zPrQbISOdhQs8L3iFSyW1E6uE0H8n55FqQ5MOcrMSrlGYN2Etq
roQ2/HKyn50TpdyIc5qQbw+47yVeDPVvHiaEQqVacBzqH/7SoQjP5K3xqNw9ufZQ
zd4Vnk0tVNqkpASHWaRFRgFuq9aZ7V62CGszhEdkl2i1EEwi298TjOYNaasYHRRL
qJlhalJf6/1sHWFebtHlOMtmL9V/ZBD0GeRmaXJUZzq7bdhMdObuDIVnqpSYF7bj
6l7ATncFjeGGI2jlIhIFGU6qnM20vIqj5LGBY7+TEwjDk2PUhYlSMOwllfYs7Xpc
N0KDFCAZa5F/1RNt0VmTC+BxsxTHFdUn+jNSEF9hpx7kcHhpjpqJNyRuchaQcVk5
NgYJXnryzvcXoLnA+NFFvmWnV7PKSPglDCqIwhrSOSXHJVjvi3AwzF1R4JQzzg4r
bgBpTU1cJ9Gnjn+jYAZrtVpsYEieAnreDlsCq6Qms7GIFqkcg8x83shBjf9zh1Vh
rebT33PvsWHqCxjGL0MJ0V+BjSZjep6vaByUDrt4Pi+gp9h4TF+Sk5O2FbWTcA7O
atdFOH0UVL7sE6wuaJCuWzUqM9UBGRRaitTs16cVF9xnKxeCUlbvP+1+cXWXnZ+N
K7I6dl9EUI9kEd+Y9X/jvkphkxPfTEVMa7w7sSZ6fuGt5U1WSn3t4KiIp7CUee6T
mINCNulymfnrwGe/BafuwG8kAXUd50ZpwXAB9Y5bYxY97xS1wdy0+OOPxHhMhlxC
uapN+I6kJrp/jdZKaxK5zJk7CP0G0DNrhDKpvSNdJ1xBTi63PoEHBIlfcsluxv6+
yeb48ksyg2f4aJ3S//L46T93NvxJGWB3Zlohjhn5428YuWJHaexFb9j11ivd5LdZ
gyrP01arKJTvOsrm+R4Ur4O3Fx4HsYVjtHMSS84+vOXpgfy3x68lRwv+ZI3AvBKH
XzPAt8JIvOmv2c7fgzLOl5dHLR35Muy65WIyf5vaPNlmlP+6M8v3OWhJiLHBIHK0
BBXYlzDL9EOIeN0kIDd4cPJb1jiB5Fv7KPbka44VFatF/Tx3P3qFASl9cqYUhcuf
KwlaaVbDcg80fAeBF9qEd4nITsAdVHTABJrwxW1fvSJHI52+yVVXv06onnhOyqCl
2toHkxEGDpInC9NA1DOVeWeDMtyN5CPx1Bp4Pvqg5qAaCm44NeQxq53bufcLE54P
pQMBN1V8RYX56Z40xq6s9H7Dklveg47JzkZJQ5WgMrsRzOCiutuGUJ5dNmKvanUj
tNJuBrqaz/tYL8x5SuMbBwxb+Pl54yDBrTZ5l/oqe+J6ge3WLxDX832ndeObgDtn
CjHBYG78nnV7/8niK2a3vsNd3A9nfe5K0YEr70qyr9PAcEI6vA1vuiS+tL7AF7Gd
I1B7roo3RAPBXcysKjrGxHotJUax7o4WaqmPdxzFpbnFxXySvasfxzGvfOFGWpHr
07kA+FM7vB1g++R3L0OcleO+LAtGFC0vL4dYoZCd6GrX1B0xSY448X8q1UiN4WQB
ikbjLy+rnxh5mNy3fFz+Hb0VxEDQ7NXWPEm1R3TchvS/CPiRq23z7luawUibkJDI
9JnnvYJmzJemm5Wrvtc1+ID8KmSGhmXWorybMgJLApsCkVK/FU2A016BiY58Xs78
oEP9ifWccPM1h97hcM4FvkcnQ/kkEbOSORsKDkcIY1MyqKZUU8Z8hYN+1Drl/LgJ
A6B4MenksEjVJhyBAh5BXwPp8RnvZtyoPp95S0ltkdWFp4CKEJafCjeScHhvvqHc
F9woH0NQKaS2yuLqSHh6SsdmKswd3NI5MNIwKEoRHGs59U2CRWai2QM1PiBRsvyo
CKQv88YdRy6vV/a2dWaEIUDy/H0bUpjzXo3wHDjrZhRS6397cU1lzIysa2GyQyfw
PrIIFUn2gQfVMwwRlcxdSZXLbk5KM28xUXIPyP52XLB3tYKqxgz3vnAEk/7af3Nz
DmrBjkv8Pt5/S4CQTQhJsWIy6n690JxyytqqxHdTm1TMSVXqdcNAKe3a00lwQ11P
KgFGKyp1GH3qxXdku/MQepevwaAPP3T8BGUUWVmaFiXPaAtqBf+xQebzW1sC33Il
nTqUOGQ6QTZwcVpmrK8tKwgy7l4LhXRi4ciMeSY6+eU4Pdg6+hscKUG8GoXwkgLy
cXPSC+pTquAoxOtTaObgCBF/8Rm0uwYfXUgDKW5Kw7jWqGqpKf99ig8BAILV9Hc2
177YoS9mZXGkn6gAfIb159HbEtu8xZVFOiaEpv1DLHVwjIFO9VTwiW6SxuJTJvMm
6DUXZIeWfBWOkICFFCbns0P7ki2jxrYBbhhKvcW7Hu81TI3Hz05E2cTwSPi7OyFu
dc0JmVeoFNdoUxMgyvz5OBRM8BgHHBIXSwTdIIDCgR62qcwwBPJfaeCC5OMG8gT+
M0uXzds8FnExYl2hBYD6Y3LOChA2zlMOcwk3OrGIVG/EEzfGGOU943m7kYMCrUqf
TifEQgi7MbB79Za7IqRmpBqpxZFIgrAoaGv36SK2emFuBIx2hGGMt5CGTmOtrsFf
tUmUOIFicKsMFWrdyKZutT5wO7Zs3+WcduyF9vzOHKS7POvO31y9g6ja+DTo8b2C
Z87pUVPI5KCESOLkUubwVEHSNRgXdteCvpGQZ4RJ4+l1GF4GrN/K+Q4t5nljFWPA
g8fZw8eyuh5q5exj5oaEP7nxh9knmJFokb86HGlTsfnFISJ222nGpXFcUsp3PqQo
LwWTf8cnpYxryrQliVD7lVY8VxTUzBGlSk3Z9zqQSUxejPrSZWyxJNLzFFq4MF0u
FxoZz+KMLVWr+y4yCaFtzBw+uhpJkCEJEaZ81i6njI+XMuX99NRFBu1P8LnejHgZ
abnSXG3dBPd/NB6Tf9ZcT/YrTZXdenkp7V6qhSclNQxm5OQrNgxd7GWB563VQduR
21iGom7QbqdadYhrfx5ycdwfrM+uDtDBGIksP+LQz8R7+2N3AoHXlIX2z5v6zRUO
7mLXhuPWrp7eOPUtl+9WpKam+TBOxQZXYazC0QmdNsaN+upz3SKxFEGD/1tb2IOP
COVmFxcYVSJTeduTuaQmenJlq/DRraaouTEsc/E/rzhNZ8veuIW5/ybBf/F/seYv
DpiVSNe4yYtIKaQgA68c8XfOmLHdl8uCxBlXHKZVe1QV8jduoYt82sUq8A23CafA
i4cuNPtQUA85ZNl/gnEu2965qPZyeWcM/hsXxI/asNEsIgr4wwmX80LpO1CiObNk
QymFiUeG6rM3NHknP28u+wyXAnrYcmu4LZhnYWF1H/D1dZr9SxMTljG9zn+Xu4rg
jlgTCxwfhkMiLbBlZyPMp27Zl8cnmAnKZBx3NM6qRGu05+7VsDXNs7VLtRfoO/Ni
iolOpEzFjdhtoAGydvzkR/cWbfD5V6Y85gyxYl783q0bbzUlwTOU9tVs7c9DFP/G
o14nNKJ6n7Gcz4Yz1Bge4eRLKCgsqjmDu+WT4S7d1MkgihkK9CPzohKyK80vNP76
s2/Kvrbj0MS2eo7jJMjR6Ttq4U4DrC3i/qdCCDmwj6fgCampB+uNOpQIafMnwikk
9/E1/CF2a7YNKz+yVILTWigCYEnQvKFOhM5YTaYOfIQrxoLzOtgQYvd2fbv6muDf
d999bgkA996BhNq5btIqeMWuyrPrZZnxQfCe/Rne272D9sqo6nxNcX0oOh6Zhagn
PmdiAGfCysVmNFR3na7ORo8Z/a3BHv9bW8rfsDS+nALIdEpLunWd88J7F4QvZBFD
PLXCi1JSqTr5/MtgjeulZOF3psaehaurYgdOVEc2oGmlzpripm0HZeOpS5epaeNZ
Pj4JVbhA6HWYv0e0R57a2rnTptePTxxRYlQ0z+oBNwz/8EZNZWnWR0DHjW0SKJqV
KAZg9sluypk5ALYWfjtbJAptoGgAH+RPM19gqseNkws29MsNVn4djP72tDGH+hcN
elKHvg0dxUaMIKXAovU74hZE6KP3WjQTgHkZP3JTGgBqPRdBVNQka8azieg4mb/c
ZYrdvu6VILL2JuQ56rDBEemQEnnyFMiEhL4PvYCg8sWsFH+ekTN+SKApk8jRm7A5
23HQ7rjiLc6xZadstoD0bY91mFig0D1ZRfLNqjYWNGhDmvDujv+xvVVFaEF7BmY8
n9QnZo6qvbu8y1FxanWXQO2qpv/13QR2c3I1Y2P7rGoA3BoCtZZHm2o86I0NOHnC
PhenHOnaSArOTGd+Pv6UVGm4XPoKSng+E2pL3u0o8cxIJ5bhe9/MHWG79Mh+1fhF
QZszANFvLLx69LZKZ8/ccnkg3k9QK+xj8fvDVBNxlpLMJiAad1xpqa9GecYaoop6
bzBDZCwS3YcziNvZ1h5FrhAdRcjmR1HDHWG/dbJYVsDWq465qhFDxOkQk7r2FRB2
2fW8W6xvrI+le1IPgRqS8Zff/WevPijVLIXprvqQmhUP3nLbnJZHwK2Qp2dcYDmT
oBo5ZlwFYJZDHv8w04h9BOu5y8dEVflwyE8IeU/ei3fXW4G6rxxLQRzhtgKRc3Q3
vidyFl5Y6g5TdZ8/RnwwAqimQBIcpnCEN7TBPxw+1kxinhYX/sxhqK100ADnO7Iz
RVIeRC4tiFqvut39VusORswpdHBpfADvZlzklGWgjBBEgCVYrpB+zCLq7kIbR6li
LREmtrH63C1b8NSBN8zGoySu5/rH2E2XiIr117PlIOC6PpZZBktNWoF0PSSEXeDA
Ag+YbohjGbPTIbUnXAHz9W9v0h//A1l1KtNwWcDDD3VlG3SIE1ptDZU00gW9EI8S
mfZ+vLVEBUtlK2E0n/zhb3+kvCXNIVIdwple7BPbjDUgjzCqrPo6kGof4h/mVHbI
EXLd4eUve+OrCW1u/DyTHUXQJPXxtPmTwPkw4ux7hAKld+ZudicaNzWpLfNV2snk
6pqk8q86c49gDZcU1xj4lNFYUuSASE9sWJePjCTdEVAT0OOYjmBFrWXKgn9Us8Sr
QE4KXwQZ0COQx9qUCawKPOZvfUaITqjXe9QDKt1VyaPVKguTCTw4FMBvv72PXmtu
EzRo+46Lb7PQYsI51k+In9+q+riY/w5Ndi6Kfj/2ziUAZDpX9HLte0loUBSZV2WP
6s6iCUXOKW+dFxB6kEP944EHvEBhI9yaK49vVuSIJgBuvcuE0Wo2w8gWsgfo53rn
SBoDwGkytCZ+ffV0Q2tgU9Y6DC7erhn7Y8UfjXUhhRPqbfEqz5U3Fn4gNpiudJYu
dLMgWzAYIyKoaLgNLldGDUdjI/ls20p9YSpGNQ0FbuUVtHfso7UUx4dNk7Y7UTHl
b6phlp1P8Li//uGnIjDjgs9G4UbAOvAbF8ea54ivfbWINrSdRFuw3KtixyGIUOcD
6XQgC/Y/wr74IBYCGr/NFBjD4J3Lm83DifsJL02uuw0mNEvpprIW8VNv1Z7Wfpf2
D+Sc9kgQ//XBfHG8OqEY7XDoFOZP+bikD4l/2rxpUkYBfoZv5Esw8Hi3zkEOBdMj
7TNkQABomHGbY30eV48jsO5nT9CgwIU3u8L2YuvPTQ1HM1U9z9D1ZLmgof5K+jp4
JNz3s3Uo3f0FC4jsJN3Rxi5GTdM7+nNH+4fL1vGar8NH9GgOoMQxPqD/NcBmCFlf
RMvRxuFC9nIH7UFnuvtaL2/l+jozyv2Ea52CpqJCeLb09fDDeuepNNphTN87A/ST
4KPlRuQ/JP1Anbs8m+5ro/bMjuT57+04QnnbxN93cTPH7r3IlpsCZiKIfrN0fQWV
F3vYrtCeRtp/yXXBQggZZj52MHFKuAqUwBeFFNboQQTVKBRXxRZZY1RmVtNoGio7
v4oVAlRNrHfPBb8o6/5zr+BzVOxUw6PNEOtSgPOyZ2Yyt6RZvDXJwvQQJWOF+u4J
jILp/4Nav/uCxcQ8p0SJ22Ud6BuGKyd3+NwplhHo4AK+vyIJWzVPS6zt0vqw9y9o
RoonGuvGZABp7fjjBERZEef2jzJFn33hb0cL70xNdWSv4ZOadVQpYURLy5ZIsZO2
s9/1WcbBXNX3hix50kM/A5NC2ce3HmQ0Oz5ot6GQIjszzUnkxvYALW22MtJOobv6
LZ55cmK9Zeoaqyb2GVnrRNVJ9qzVSw3pnA/yw5xMVNexTTF1FvTWzkmqHrkCxiUC
YlxHF00ga4Ww3MD3OwwGj0OP3mbHoz7W0tklFSomo5BDAzkOwenn7bQTjZcRTwpE
UYMxK2ysb3TdCwS9NPREoPXTQhirFKsAkGaG53+Qtvhy+1JzWJtHS0pSSjCPxXaL
EE32hA4xyF7FV9L1zpkALBGqi98BlVrvuSjXdf34+ti8Y2rMCTQajXKkMqMbdeiR
7OWtvrxwGfbJbM16bblPlgOaI9B61S7JwIb7JZjOySAN9L3Osm0ytRHSaNbm9zhX
SCJrfdKYLWGET6dJLQ3y12UOL9e2vQgYwIisMV3jCt7MZWLZMajpPu1KzMgzctT9
4nLM1ZBNo3nBE2YqI4xBkIK1B/w80Ks40cK7Ix7dKxgsbpqXmrfT+dc0RXqiJwM8
mMH6tCFUxW+04QkfG8SSyGlIfX1lHMxY6qKL827fJf/gq7xSr9603PmFRA9vW/4b
K1G0bdmgQF9bn9xEkxzyupUAbuiXwu9lkbmXuYP3T5iedKg7T4EuJYNRgba7n0SH
yM9nidwgOW5gblGewGAMtCqLRI2B8eu94o/tYDPGsYKsH2ep29txddNBkGny2hbu
5EoAOlB5A4fGbmY3hdAfR0+PGoZi/CzMfDKqee/kCSYQXawv/CywN1U/1jeaulvq
vOWEtPmFQBFeaj6h3ttiaO4GtW+t/cwQFIfZXtr+j1kO/KxoLXKK/nxk3uVXkzqM
e85J2y1vG6cYLDUN+C0MUubS5mTbqVkGLrT8uRo2QfXEQvI3sudVzq0qug2TfSB8
G4Ky5PXhzJQuy+tvhYIh7pmzV7qccRK7ETkdTzZ06b4bSaS/h8f9pKuzZSQDzku/
ENfUslj0v4RjvKCW9NKk1P3M4fUUAzuGGj9vhHjefdphCmZqL14erozm9mCVZMsk
5OUxjgCjM5jAWe7mgMvM2aqRtfYHlOhYE+zm4SBKUTbhZJ9dl72xNO2RGNrDgb6d
lPgYD+Ih6jc6LlWAmDWkdRJNpI/RWVHT7JCv7UuLFvYrdcLlKaPAOMB2kRG+bBVb
s+LHl8RFbNxxjReGzXVojjim2Nb6XSAvbqPJd519oRoiobHslTj5NFTw0ON5t5/1
L5zmhcqWbo/5nZDPymTMcpiO7zFXAWSMMntawIL8jFxv+ntITW6B9Jj7m4s1qBSd
mHtP2ztLGL3TATK+GHfhyKox5A0qrqQrUMzlaxGIbJZojrEZsp3IYziHmKvnvAOk
fbXtRZFnXjeumxltnnAf8dnZ8m07yaPF5XvDB4s3pw9uEdNYmE5Al9JuoQy6VNyD
xzbMXthqWQVabxSh2iELE1FnAX13MlB9sP8buFDTNF6ac2t5N1oS+fHx8NBta9WZ
lKsNF0c0NUrHS6PYoPSrSxsBr48CkIbtH+BbyqSMHdtAjdRFhYIQ1hyuDfd8+OQJ
LOx7bsjTTQpr5/aMU2XXHeZxOkAcw/WXv1aSDOa75i5Rhn1X0mbKK+H5VryiJZ1G
7Gbh3gjj2GD8Qnbw2kKL+iCY31SDQ6zl9xJGGguSnrEzrX8ZQb1C1ZgAkY36LgYi
mTmiRjbTOAm99vbJIlY8f7V+NcgNdkGPVCgDUkEqWAhxiXrbfoGKA5dWLyiXkqdA
7DLp0ae3e7bzHC7AzYvLTkPI2KSBSW4E4C+wQTTju4PSiRii1FzdvKkjmJtdJiy4
ajLfRkh/yrlN9QFGsyB+ya8sKYuag4NEsm4HozmCqisNzJixLAJxGjH2yV346lX3
9ez9gM7jAAgBhfyVhgMsMxn6YsQZV2rdWo2/Xoq30eWAZzM8CmVo8KVePORN6Gmp
mHZ1sV/HRRzeye+oxToEQCKI1VcBCLP6kfA04GM5UJjVJnQ5dazdRY0Vowfvirh+
Z4ZcNNH+y4N+QwfS26ThUtlp668KVrMxrBganHTZyCtezQGotPR1Yvk3TX2OvXGC
W+sV40XR8B3zz3zHzklu6CtYobNDRLF105uXm9AeKLrEruTtUYSYRbntWt0OCeEc
19JtqcRsYj18+2IPWNJ7v6TB3OmUjSTpoZ43HcScyQZKmT9X4RPXyh5X+NiPfgfP
a++f3Y/C80pBCWf15AoNUJ669c7pDO3FdNnVquchysZ23/cyeJjVQe+U8xfeBJ5/
vUjDhPZrAxvD4alOdXRC2JwIN3XS5i3aFxQrTqWfdhsSRMAzcCl5GpBriio84dmM
ooGoI3y76aXfkZNMvVR3OmpbwFBgYXzk8HaO7g6ul5Go4qm8ztYmziu4VG7LvjFb
AviH6HpO7ZCXodbq99bcABpxKXe87BHChjNdxkwVAjzraaOU6P5d0naXxSXAQ5fE
mzarfVrqUcy8BNAthd6f6MkA5h55JryFNXcMWlFmL5plmBrxuE8YeG5Vo69LNhKt
FVFXmzz0Je09WGdAtqE46qsaHhCj1Iu7cPulx2aO8AKS3PXYGaHcWHNmGSdPund3
Yp71FXOeQsVZgUO8/7aVX0U3sSA9HCX/HuYenpTKbqcmg8gdX39igNDL0VTGoGqZ
QDxo723Ncbsl1pUR4lBUDuK/A93YnMEjtCq7TcOuc3BhLDDeyuJ9OfCp1ONWEC12
tk21CmNjRs1Hq2GZI/vWhMq8ZRbDkcm7kffp7KBAWWPtzB6mu1QsuvXAWcdQLcfB
gXCTN8wTshPQfRiG1gTrb3aqkcZSpndkT1H1OH6SnYYTazYJBjIWDacBEVmsR8e9
ZLC0bG2NBPuRHxB/gJ8e1Wd391rpKIGDCflT2H0oZL4kO8sAjHgOxBIxuxtqLRLL
bGnfg02ZG29u602O3OiPNtIoTsfMLZqWXoKCq2tee2/MSuhHPsxUuakOpEkZ9dgn
2mGp0v7v/Zr/ypXI6mkcAuGksBqxH8T4AMB8qD1Lz/Yqhz5UCbZKXcagqk3d/wRr
yLNK85Hp+KGP6AAN6qgM7GhTysrDXjjRqqZGYGHSOcZoj0VEQcLfO3aLFlnRg1oW
n/LRIu73htUfVe8bFc3q5eVLKi6H8cYA0VKcW2LLOGklL1cuu0H3xk0cEXnPDPMr
nlIQJ6k/j3I5r4lHqcUsF12jC2jJiVxg5rTYwtZGS3dTVMWwqIW2v0WSsXT23sxQ
5YEt1RSOEm58LeBGMZYfb9MY2Rdaw+RYQ5SZBYukr+y7wptaFyRGtbK/iyxHc6HC
kZmMyD8suLSxxMkgTI6RkcaL0Vtxigb0icD32jz/kh6LMpMfBYyjWBMdidvwX2KV
ALIXjUC7lSQ0hGTT9faGeQJuiHXV0nPjtX4Fq3nLJgz/TWnL+MQbfFNyQLVIhXXM
2XjU16D4pweae1nKGI9LhQdOjUEqf9irNQWa8tvtrSg/1jYfx1IyrqyGNEK/lqLY
9obG+SnjubMzDXiw58V6b7dSLzAjStZIAy3m0DH7Yrf8jpD84l1se2dOn9H51X0E
h+yuhQtB8pcIkPIUKMUNnYomII00LYgN7/GUYwVCaB4wL0kN4tegGbR+jxaKWYYF
+LTj6Ex/cMYMEvj4MjJkrboWAzlcDaa+tYunybv1RJcA1q6H4n01qPgMDOHwKUEg
2e2fp+PqKKlbfw0213yx8RcGUK3CFUFApICMvxqWEbyxXAqGF1SuSaILd74bVNUR
B7njqqIfmxDyxFH7wrUXRwjX9BWIqe46cGwLHB0XWfRNhNDOeIKK820lAMTO1ii3
bGVjqj355HYSIOi/dljw1r5g8v7er6hRAqEFkdAHQ4d0iUGGLDg5qlO43UHTxrDX
6lJnxOW3HuZQSJ05r07Q/xPmgy7icoutLTfpvsXtxxt3KVJe9m8ElZU+rzgp0QAl
4NHXv6mgVdIgXyUggBCimAS0al2NYlQJXILwPmEuc4XVzjOYB/lmlzCVlIOOWY7R
AMolK5WHyaWbu3mlUTuFUq49qpfgUJ1oFxaS6Q5Tiq0PRIWOSmvD+teuxUhcO+0m
ofp0d8I4Nad0dM5HgUlmIUbbmxRiS5noUSYbakmP/ixvrUfOzFy/77tYmQSTuksP
CQPjl1euPtTYlfIxNGtM0hINi5dtT9Dw64G1y8KmMvzsMf4kony24OKKJFFgM3Pj
Zt71Mp8VE5VV3rdE1SJu2BJQ4yNzpyHWAX7a9v92CGkQx8Zpl2cvHGd6ai9C+SBp
gtAWyG8JZaip/KMNbIF9x9TSZpHa4BZTPScX3E5OaEp/B2zlt/f6QlEeO3z8gBZv
BYtxAFLwhuSZQzgraiZuXdPa2KanYOAQmlIYbUg60j4wwkHBCSdSZ1U+VuV98cBW
F3ax8lRGFeYMRybpzP8IjRhI7iYjYarB9CXSpko5W3eEx2B9Vnf05JKM1gXT91KY
awllxoLUcuZrGpLObvCowkhQ5pp/yNYiwcCBpTGPMlgvwMZLqsK8ASW2obnfA2Ui
/tJid5NZwxah5C9RUk0v69NVbKhWHDHpUJovVl4GxwDp5frnUafc8Qit+8z51ku5
XYExlF03lnheURB8uDXUrNChb6brxgaFOS0jJMNIpr1Oi6IT0ESIEgMhT3SyAaMz
pnefAPl8JkPXrXCocngTYZfO8n5yiwz7eBHF2ZzSFjW3mbTOPsgUWSOmrUfEsHaE
HtW5N+O1ro+mSv2FSF8IHoEVl6q8u8hmEoUGUK+W5MFEopc/LPyavcIfhZjeRleH
9OzOWrOWCsn5peHJuXmSo1ZqxbOggyF9MyYMT5tyCFihBr92bCItPWRIvBEwojY2
MGT8398/+ncyoQWBLCkDOzVpIGJlCRGqJwmk2MVVQTeae+vtHQBethhFUBYL21x+
1FVueGWd4dGxGX6e7JAhVlQQkSZ4nGSJuUc9BEMaJEkD3gpdWKlVG//5o3XE1TBr
1fqjjs9Ha3HhML94LdIVOTqcRCD2KaTn+GeH8bXYcivJiGN36CTROz8BRC2+AsIZ
Zbx538sK3GQtIkZVUQNHX5WNHmY1RCrUu7S+txwwRdAxRPC80/LJAhTo+UKHdn+G
92FWK8nvpvddo3EYB2a7ym805bEPnKsvqZvtIhbswpcBVvmoKsOA9csgTkBOUJ/N
EGsTgwZ9dx+fHXJhvxWkjP+vKuZ9ZksUKsX/OJFsI/Xb8NK96/5Zrd7mWKSNaOs4
molwCb30RFuIcp1V3sDHeeJtgRpz/PRbyWkdpGlI58Dv/5j6VA6qBXEGxRZFIhm8
TPJDS6N+yj0xij/k/jSwMXwgrmJnBYYYhOylVpseW5m9KjJQDg1P6xsfnLQbkXg2
wIhqrmR+iuILuwe9YNAT98yKPPQglSQITuwK4sOcFxmydD4L7lT5AdfZYm1072QQ
oYB6CDi8sYOMu5KGzs7O6qzl09kFkSyUjsQ+S0+paCEBzwyumPw1Oj5Z7lMxigPj
1E3/W0xN1LesGs8cs43RbNYORZSu4mqWsXYWNkFv9hbffKIYuvLPiYtKrcF3jlrZ
+l+GPVRbiwsKhMehhcOWQghAYSQB0JHoozfQP58dFQ4U6EBxV6JYUVri5v1X8Yf5
8B82T5d7E9bxaFybTEsb7rQ8lCpxzeIgsbHFZtrktmL81lCeoTjFIX/5FkkIyAwM
ot8XwHgSfvReJ1t5NUM5jwja0NI5/auT8lENiGmihWTEI40lhajDbmUymv0LBuoz
Ai2IgnyvF895doKgmajaP6tsPqUIqe7imsql5ZwWyR5RpeeaQWww/GMUzNoM0wdu
ypBKmwKoMBci7UfXUuKIc/ZCtFNxq+zj+EsD7kR6rFcvxePAgV1YLA/Dqdjp2+V2
PluFPPjLE8SKIO/LeW+BiAfwBsblNLin4iplVjnjwmHR8HAm1+TMXySefDxoFXnV
mGT4FTw9s4SXBsAZZzOJpYvINPXO/jTU8/fMxQaF25P8Wmv7RDradRPqRo4kX7CY
zlvHFeGTbqk+6Hsdk4hTYojinUJGMCKW0MKIv0DzYAnk5OCYKxIOmFJnlSxwzG4b
VI5NZRnclLCxb78wpNrFG/EkIaMG+HdrkBJeFgYRt9GI+69O+IDGFj+mRXLitlv2
UUcRSrnFhn9oJddoIzq8DuFMSTzlCwZUV2dDOHlS+cyKFYCCkmlW78vOitVCwHHV
RpezE59XbQiR8gxoDgxI3b8dW/RzFUrH5ycmKbcf8GgRuRh6nhgFcA08Ag/ulDu+
7LKSDGWA5l1yMzcwrXk2PEEWzYCKbeQ7ssi7Fc8iI+5apjydtmZ4c40r/BkACfnb
HmUT4/YfbMp9A+4dQAcHiRZIFt3hxi4eZDQjaUFaijOwzEyIBaIjIAysHnt6vNwM
1sJHAvzsz/yQleL+OWAb14yKH6I6mGAx4y3txkFP1kbXUvhRqX0juLho/8NE2ymO
CJRDpfJt1KDsEmihlZ01kc31SgpQ7Qy8pke0zxCJl//fn9vDnFSnz72yofSSwV0N
BkPABY39kGePFv/J1ntaH+lRvmzIifLoS/oHfOAMI8QaQhlQqSZce/1UwgoC6RjN
9iz8yQTL4Vih8idrpiZeX+x1X4yCm5e8UWcC6cCF6lUXm7LH3/je/L59H81zxuD+
LB1uB+jtMRS9YGBwd8oXAjhNISAwt0RMdnFIlAXIUk7d4P4HAPfI0+AmEPQvfePl
+5qX1QACJ91gm+neiEIKdsBIriMAyBLddvEqDnWRQh8MPAIWWCUYlJ/Whz1qQkST
FFNP3jVh/V2ZIGVfKSEtUHhzhItPqS3FOby/pvjXcto20X+Mk2fjQy58TvLPLJoL
8uxwgpQ8uCN1ykZge9zzZGLmWFBRm2jy5Icw4hSp+UI5e4sJXnZCpuhVosDdkMeF
taUmWfa9b1Puc63bL/i3ByNs6t7tr0i31QOaoG/GeJ/448whRE+jjsTo7cZv9Xnu
DqrWaysj3MBlqOpySPHmTKoBUduxvb5EXXClfx43hw5qxWExjxhf/MtWE//mV/bN
/O98nf1IdRFHXp8kt9bhLWdLiRI4E7ZZmPF9CpNBDZDAkWTb4iYF/ThKVNldiy6I
9kzSW5242Yb6j+FkB+8vnZf9qEh1o0valcfmrJWOKVhAvM4l0hfQymVUZeX6pfSW
O9BLqZP/csP6ATtC445iaj+HA8t3OGpMI0Dsc3BOwVbieY5rkENflq/KT1D5Y9ns
4nX84mMsEYHcvDxKFkSkwpueuIVbeBAve8m/OsaspfEHBELWav/G+wPTJXoUVmNV
/t6a5zHID4pQd/KYHSZ/ofoWX24YIZVwDt8xXx5OltslFgbkLd2Nqy+1XAdsLc7s
dBbNoOPsiPRI/QvHSJotHNAyZA+Kv+8tuXceV16NK0+az9K3eQfAnVH7pZX7REmf
XWPvJKRyeuu6ZeGmTJTUSHZQHTTsGweXjLOXbqQm5tkcaNl5NrwwLNm2+t8Zcvia
bIfT4kwknHZKENEjtmA6c95g0xG7raOz8mrO77Yce6VTpvz2Cv6Jmrq3fkGLH5LK
SfPDkQSBov3hvr3g1vc1KO01GmrPNKLI9ZE0AC+4a/NCnZA7XeFui1/qAeYYn9xY
IdIf/L5zfvH4Ay8oqCcAogU79/5rjKooRffYrq63o21oF6p/so3vVa4ZcZoJdPjr
C7XV84s76mdRL0iwyC+iQML+AX48iERbpaWgZLEBN9Dczhb+f7XqRfwfL0OzXXHd
EmKG7tvXqntvGVcGEeu8M57nGskxEdOxlxhNz7Rke/kFe08te3qeOok7biZ1A+m7
KBHwwjxPJEwBzqlHhHe6P0vF1UW4l0zmY9BLeJaytpii13DJdEMYqihiLufE8GeF
0MOKg4ZxiDwfnjA+a/uVtAfTZCQod29MSrXiWcVMZMJr6cvJQm6s+3lYICL9S+ds
NXN75DkHVfvEwRVK4E+c/Qzvktf6dW4EmHKJfxQyVytVGhz3RcSxofyYFH/FkbYL
Rh0FjBfzfQi5xIItkovNq/GnQrZUetiHCDE5KmBp9JeZeHUrvvz48nWg4q1ElJN/
IaWX+Vm6qVnC8kxY3Gy0hL5V3Ay1v+CRP48LkKZRB/OmdP8mQzMQihoLbLZCgmdu
hAikRSFFyM0oYy9cO0vp9BhtcIBV06+C0orZh/8Nd0dawM0aWgAhKIwLAZaOVRmJ
pZyDlst/xNfxdRuGCcIzOosdOB/l1+bHi3rxg+VAatZVhjSFusKNHao8sLUMKiH1
PrvhNRW+LClWN58yJngm1TDGOYF1eup4YWnUq3O/mJrM3LjlXkAoFt9uDzJ12fKF
rGUkNjKwGDECXKJIL0fl0PDOOTv+hyFPhM5yFkKdNRDceJ6oEES9IbdfslxLeK4s
T10ryTctOaz7wLGeL5s0m5zzSXNvoTuTiP4hBI8ThLQF+0vPtOM3ik1adCqo+f8Z
q7zaUIBepMQ+RE7wOu0eRpliiJuZfGkX1ZTelOwVUMfo1dkM5q6MFxbDdj3G1QL/
3h44xjDk58+oaFCQXk0XFSUkBjw0xU7V9lLYbcViFu5F0j/v3M5V5v2XQbJAtmr8
tdO0fKAqcOEKa1lIdlCGzxPSCVBBdAjZfoIv/QekYNLmMwkDpLTS8iKEHoQzJL8c
5n446ltoOHFoViWQUc1YSHps5QpPZCCzzGK3ltM9P6G4tvNv3Ru3wsTp9ngTbODd
fffyx2Uwq3x9/Tu+y0xQojmeemdDOsgBzPP5n8EL0D9d7U4wOCBg0W69qMENU+PV
SG5Xf3QsZc63Fmk8mKoYsZU7EbGMMBF5tO3yT1trDm6ru1ESWqd7fE2gn4tlL2ik
VfcXLSxeKII0KgYk871NPZpVNTgU6wG8CYEs839/VCR7cacFTBq8sA30eqUb80Jm
6W9clameckDe3fPUAIqIeG76aQflbGK4u2ezJwwQpYt6pMemAA9lOxOpwlY97oa8
xqiFhkvcAojlP9yczLuL+wteMOe/dYDDZy8tl+bq8WSPaaF6O9/7WbY8Mvb+XXOk
W/qWhPn8f/u+Iif84j7Tm7KAScHFFroR/wYmMXHT9hsDc/QG7CyjzgK28aTPxef+
NgH4BtF6BpydNSfSDAQ22D/5iXR04U1QtTgprRDkhK20Tg0R8uNINFte2ngnIdv5
uyJPhNQMN7UCpO7eMR1Cr10soEMate2Z9x1uSn4m8ifmWtpp1mPV+mlqdIVtxuHQ
oqjdeFrxdAOH1OGnjRem1b0sLTMxFnV2UBQEtqu7ixWGamzqtqPiN2Hb3ks0MS2d
TuxS7n7TEIQCoZ1kuAeZ6cJqopCYKdFpPHudTK75MtJ6eviiJq1SSdRr6XM8+6Hp
XS+fTJBlI3d/5TrrNYohKN2XfvUowZNorTZYf8CsuKLoh35d2e2o+nJFHQ6Z26vY
3sqmCyGRofhMbodaMyyKmP8Bvr32SJY+IYQwiGp2Dw+CE3Q2ajMypCCo2EVCtDKv
6/JCKoB7tPn5cig9elvMHS2hRX61JY5C8xfMp6k2F+fUNbQWjUghMuHRPxhozz12
gcvUpcoj4LHptPQexbYth1Xg6OuFwAlC/Qa+O/a6qdS/Wamr27zlYTJacb2TAFYv
akM20lEB7YQnvdfuTBHw9DcJyHDZ2i2gaNzi03xSWyz/Wkl0ZovxyjzQtXKVt4TS
8mrJmu9jXhtHNv7CIaCcrjqu0oY+h8zkKtVoVR/wQE5+wGfEohj+XgDM1B5YPDWm
v7E9bzK5rnbWaECytvp/xnsY4jnSuQpC8IDS76a+ip5fz+vHRyyy/UwLT95nNYdi
GU+36X80uTHjpVtZUoma/zEWNlQWa9okdw2CaclYb06cFRIbsd/TAdRc26kqrcb1
JaHBb2RnCd/oijphYngvvx0ZJwgH2Q6BfHI/foP7Ygi56oxrrzoC0rlxZJ+gh6JH
xMIMtWmASBHuVVWvb3KkynUNyx2NS+eFaqM7MjrXkUdj1GXpMRNEnvO/Pl/Z8qPw
zzcIQKzbqVyR+BWQRASsZ9XCBeFOje+/bkTPi0GkTdU3aSFUOaH8+7x8WjPLYvx+
kMZlH4YKaPEFleFBWPikhUEt72khPgGmSaqp1l4M4nzME0BPikEh/zOD4YsaTFdy
q8mPhmvGrff/qXhzS9aKanhM7oJa9LSjFzWZ9oy6yva5V0dnzZJBS0pdMG032Ywu
XyOMGVrKpHXlOBZ6RpBQmr77MhWeYpIC4NUzaNb05fQsemQrdmKgbE1PxBWfrIXd
1LDhe1f+3dZ1LJBQxziE2mPMJxQU2jlFZFME5s/gMjpPb5U6BVgCblTd/hn0Vw8A
3XLvIGZRUyQMwdQ/sSfrUFlgi8EUNtmZ1l4KljT5vzE4jmg8Wfz/G2Cg0oTeJiJt
uaFurxS0imfYVyQdf+odFSU9QyqBb15BNbushf2ZJfmj3+izTaivQbHrMTZKmkwt
LEx5jzHwt0mahfvobm4UtMAZi6LBh87rspE7R/XrgdD9sJZDYEWyjirY9zbbuIxJ
PK/xjK9WiZI4mp9o2RPO062zwGUU9msQsoCT1rf01qllw0OosvMRzfXzxJo/fRGw
466SC4HNrRrCqJAnFXQl8GSxWb3UUNuP0gHNKX1XeGsHP1fD0E40Ccl0ou8JCkYu
NTkx+kxFEWl4AEqufCkr5xazjrn1EIjs70bVO5PB/X7le3Rk2GgqcWNEm16ITrAH
cGQlzigDCxo8x3aMyiIkns9HEStd/PXytuCH3JKWYjsXQq9gmlNIjY4Gc5CcyYO+
xbgQitz+mvtnsgfmzVl0jpuZL8ALQWqrSqr0UaVHvdwP+1SuGM6e+yhf4mZF4Ydf
5eHUXcIXt99ZxcXf+0zHGYZ1NDow3Z9F4TH4btNJfvyRwRqY8KaUkaZa0WLNOqeN
8Mipfc3qbz77w9fEHM9NC7JydGfExBZjHYnqxfxo90ycleoX6GfXmBFM6rpX+AOP
gzGmn/jTlT+OoPUSsaGLZZuJkuImmAc9ubFlKznTFNgcfbhQAzmvDWWt1R0qHdtr
AzWpiM96tstpcpoKhxrnF8zxT3wAyqRAV5PX0xm476GnBQYMA9I9up/EssCmbxtm
J6oPbkdVrpALKl3QbEKqMbPnYvFF5EGDG5Y7uuJqk9Z+iXX5o0wd+F2w9tFTwvG3
v8GWtLIpV9X2ZX4HPv9tNIz8r25NFsCwVMkUfQLL8lk1A/Zu7MRyfzoijfHb2jyZ
vhTtSK1PGHgWBnWbV6FpWMpwnRrRs9teEov48kC8tO9rMNPTCyafDrymtOY0u4iF
pUL5rk4s7mcckCRsWwh8nywoYlWCG8ce1ovI9+mSO9X+q9xkhYl1uuDqnEfZ2sz5
bx3ULlwPaJ8xmmRbC+C5u3FBi71qDRZgC+Fe/MTH/ktBV+p4DTKAKmFkZp5RwjIt
UE6cJNn9PKs0kVOVxqV5mGVtzdG/WA8q9JFWNpIAPZQbwQxU/sf8g2ixdeiRcu4p
eU2Xz+fzLP050kQ0r/j+FQ9tMxaGvnaewrcm4srHM4Rr7jCwwiscloL8Zqb2mUT/
ClLi6/sk4Qp5IylOyhjq8D5zTfWryiUVR5LtonFfdYx5Tx5x0uAN1mWYrJzWO+0r
/RHiGlAMYseFWl1TQDT/4dySNv9aEbvhl4Uaz7LwQCqOniu8zoi7TiQNDndep45a
GRiutJkcrndNtzPXvATaTYOn4CzHnEJT5AO9BFpET8I6+LjJKWCpp4G5zAWmOlW5
VesXJgI1LKhoFMdULOu7wbIKpdNpUOllyCX17hFy1XngS4iIApUXiHSFqqNZ7v2U
MViLcursKMAUFvT00UYr2BF1fDo5JZIBjjfTgrN5CjuBT5BSvwWwjiwSq8Nwcijb
Ri+pr+QQ4JlSNKtpsdMwxHYtmTAecB93erAzdZDMSmIHtpbPj8xlWFOQaDeiiOHS
3M8UIa7/jEXHtzyGNItPhip24cbV5CR4Qp/QZ6YsOWQ+oV4GgLy9+C+egUBoh1Ol
w04A3mIE7gDVTHcAxG9oEST6hMtgkSKhZBb9QaNtQBG2+7txy36HtfbxEQRBbS+6
y2udCR/KLwh5/wfnCEtIpM0bjDXSa/IaBdPGLcfIV+ZfXuEpi4OZHFVufhS/np7p
tqGpjqQtPEasJDONdCS4xTr+fub8H7Dyn4HN8/uEiuZGAy27IhSs8nnOis70hsNf
MKKDIAKOMp1RH1sAPB2Vya3W6V73Hz8WoV4jY6axQS1/D9F4aOMCmqM8LTqc0lx6
GG4uxpEqR7vDQQoMChUcDZy2NjfF0ptylVMz/QRbXtDKOTsx8lwpmVunE+gdN1+x
LkDl1DLJawaY96kiuKTe1DBLLLI8+WYkvnbl3u2EA9c7kmOstYMv+uIy3o6Q9i/W
8cJedwVfbLau4Z160r3fA/i5cxFRbWGbAHHYf31ZwqmcHpJVQNMmUNKo1oGFH1EJ
3Zs5XgtWPPLD2KwuusKVqoxnaz5yJjo5AKpdgC1zbn+wwD2Ljf84tyJiAh0ZgPcD
NEeN72hRthT+7lxbNXFwwLeadwvffbluHSN01F+p1JNzJNs+W6V7mB0NJxqNIIl4
E/b5sU5/Uqy82AOuEwOmUM+CJshGYz28yiYd36SLybuBpaFf42AlP2qoJBrJ13bX
tsFlzzRQy2N9lxE9CqNYCnV+5N/SGELqNdHb05NGMf1N7sF2VrTee3PYSBVWOQsR
FGpW+U/ghWt35ZY05+mdSfVf5F3pbSoq3S/CYo1chNU3Ofx0qg/E/9mkuJcuaQKU
Z83GlDfi1lnzP92fqDx/0R7LHOh5qwKpZZTE8ED7o0f9S3Ob8/eVAuoyZ46z5ANd
p0fCtD50MSvqwyYkYm+cpLy6aT5/3bLwYDmp2MTeRlVz4Zspl8aTlUKS4O9p3ZI3
52IpzresOx1sJ2bLmDFSJU6iatP/qBitxp3SkLeyzd4+VWFPNAFKAp1XtzCyWs+A
10po8FR3GA2PmNJh2tuDt5J8ebsPPsjvMMmK0zUjNgMX5/zMcAtyY0qyl+Y/G8SG
Z7mGmZVujpE8Z4yksa3GCfAiYgsturHfZTeYqNewwsu1i48x0f3eUe1DsQaEja0x
TpWsDWRAHVZyLoMQkwl1LOSSkhwjQKET1JRZ2Y0vcaQL3uEmkqC2AOLxnNb1ST1n
i0cMXFx9wFSstLE5K3t4rOKuBJeSUVedrE3PxFFR2nmkypOdvzz2BfHe7tmtLt5i
sULFL/L/sx1EfAZqgcBwiL32jOuE/9B1i6ZX1QiN4jguZjFOgoGma8caHSZv5tLr
aDl5m95h+HUkc9lSm0o8U7CZwH60UbrayCwX79HNEKDaw7NJBAAuMQvAAGtSwbCr
ZQUpRzSjBgNnNaa7HcDf3Jcd3EpNAF+nvf+lpKHVjYHnfeJ+Rej/y7rhuwzRoQVm
7QRUgOK0PPBONXK7zxFfTLBxGqymNbFZvP3aQU2unZfr1+z2DDY69HP3UpcFramz
IYvllUnim2eDo9fGdd1S8hMXJqef3/m0YklX6Tr/9ep9KE4BCh1enIcdmQodAPPk
ZdD2A1sPb2DRDAq88xSVPrp+/tR+6lmmVa7W6Z3M7P0RMIJIAjFQnFzSHdGH65yR
izBk6fpnUfXwPG0AzL2BnHX8eNoo412Juec264gl+tVom9k1ScypxkAjRhpZGIFd
JxhMGJDKwAsKfIqmtLHUL4aPyR2M0VYc+3Cr2ZP/atYJMw3VFuayhUhS9WwYGP2a
Y+ZDqS8KlL4bFdc5/lwF47VK123AjaENfq6U74VflJcvSDS34BE+w6RHzl6cHjbR
d6TMev4yMRheQCn2JLb0zFDXjGgAkktuutNt6Gb8jq/SwV0wN+KSy0Z9dRxKGCbE
WpfqrxgEUObREvt+n3PZBTbnDZu2VV6EGexZthkQSg8WKGPvv1bDQaf+5vTLiZ0Y
vCWJ0G3QFbc+3WkPiQJ3D4p++hXJNC+BSudyIWs+cEqi5MbAoMkG6mO2GqlVw7Bx
/WK9R1LobVM9NheArH9FGFJI+fQpiqgwTdyQZZl5OwU3DJ+0u5fFwk2nNr9quDZK
aUBtLzXUNaFKR7BWVBS1wpciKtgp6Jpcb5/H3z2zZS149RUNLtl6bYGVZT+X96ky
rOek5m0LiqAzKndxWe6xKgDtu4OSFlYBw1KHkEIflY2EgX95Ai0ONFgpR2vr7k/z
c5BsKwgsesauJoHH1hUp1Qp8bPSYgQx/SqqOVfG1tGVGekikujIzPqI8l7V4vn3F
iC62kMXAJSHmcMAGz5NxQ+2jlnWPyofuQgWuDt3zCOhNc9kwIwOoUbGecSRYzi73
e/UtkG58Mvyeb/mKeoSOMKGt8GXj8f+N4nY5TSZzO+hHCoCd0GKR+hogtVXZnCLw
FkcxTHB6KFEY1UgurdDYnkaAZ8Ib9ztSvtI9OhI2+0i/9aK3LSuKL5jo6N2P7BHE
WHk2Sb9v7/mZO/OFhUlHqeRd67vzCG7myz4pxx/362nRABJHaxJWfi99kLArS/gO
TxFzPs5hgMblcySQ+sM0SOaGI1d/DBI6Qv31oWmBpSC32atzkcbF3EMPd9URxv6s
zYfFeRmB7+NL0LlBh2ykTJ2b+bBkq5AMVHbujP9em+FIrtNlINH/lWmMuaCtn379
R3Uoynh/EvnjXFS/tbEUT27R403C+1jlO9+6wCUC4o4wP5u5afGhQUgBE+wlchvD
OgxLr4rPa4QSf28uzo4+RNZxnywBkRdQsaLV8DzeaIt/kMSpcNenU0pUtqGY+SRk
/7aXWArlY76aKEGsLCtySe9Ulw3w7PvjpqpKSZM6kKw4KCDoecLWthLfXCmbaA46
0JMIjfOzM3Ft3wcnOR6XoHSWuUxpZinile0XmKxnJM3rYiS/NuJbujoI5WN7WYdz
un3w5CpUjQyssMavKJRybYi8K5Nn6DYPk6oWxV2glCB5FGW7KIADUeAo56fJHjy+
Uwpa5nNZfNX+UUNkxlmcVjTMH+3VFcMST7paMiTmdoO11Z08xg+7gkF982+ZdYNs
xh00ADUCEluYhTiMWWCgFLTazNSoD7X04dYyuLC8nJafTbc3gn/yjRy2IqaztqYz
MoiT9iyxuamDOHKoTlwbJnPOK3VFMex8x1TpcYfmGzlrXt/TMVtJG4wwMW80Hlor
mF2KhTuRa1IiO3Yrs3SgZH2GbJcevRWtukJWTIeSv9sZ3CenTAQmPQXwX+3U0YQP
e7nMxQQYwjR0cnReOt4JHSsiyPn1JOuJ60iBsu0tj+geHF3FP82sfiHSv/32kSF7
wFbD+Sg4YwCOapTfBc8NsGcv0bJcs19sm3aWIVIOB4iRQb1OQQjxjuTrmpUYejxA
7uK7J2nWe5OKFfpAwCKZlWYy530+CkdGXqru+31Q5syI+nVPVABh8VoZqLPgDLDo
rJJqVZmf4tsgilRMGR5fw2NeQFRjC1pRUiy0e+H1eHG19j3Y4WSvNHQd6yC8KOEx
s5ag6msHif8mvhTxIJNoS2aJnzKh6Eym5M6BTdyIu+eoQJ/lgtTF/mFLDoJbdjmz
YrVP7wpud+3JsTZzDidXzMKcNV06OAAOVSvtE3qYLUA6y7Y+ne/sa7Ob7iWEG4Ho
uOqm08/UIGD4PJ5/pxMbBRrlJiXJ8KjadjQmkJhPm/lLw49qVqPellmD2vWW8F09
WKLhOwEV+Yrft1230pmfHrwqmnVWxKVKHQbzc6PITaSWtYQv+6vMFD2QVYvw0XcZ
p5qsW1EnFnNFCK0n3zGFxNiyjdsubNIyEG6DwSpPQOGUzoRWe++DKU6Wrbsm0Ar/
s2cRIjbISqpPVFwvPSYC2Z6zE3pnVU3t5CjyPQGIeStUjzaUolueMbtqmV2nbs4A
Z4EcD1FeS7cBgoI1fKwj/WF4ZJjjCLiNFGvii9yVwdIUhYR3zvy27qMIqzNyz6+j
oj8DB83ANsWayo9ruaMlHy/hRmMg58/OLG9MdyWT1XWwKpmR+JczfjE+W0eGgjFt
JSom1hnAVd98GjWOAz57nq/9Xm9/eASqJ7Wg8uC5NSZT2BEuqgD0xPftTw8LEuui
WPA4ySEeFKVL9FYREaJTnZMuDLPEaTOUuEKm8SGtwHK3ZKIN9Ldsq2R27J5jXe2U
cpJiLBe0sITJcSrvA6SE/dQspcZ1LXMG46UxJXjGlEPKWCklBwHnHHNA8/TF0a9C
T/7ayJkzfglNSKrdW8dHVafskCMCRHDrXCjMZrUNlCaLpgH3e2QuQz2EaMoV9USq
HZJww+RMH7daZMn1p6SGybJYIwj8aNUky3SfsaPg6Nmlkq+eX1ZzQzW+ZO1o7qym
GXZvInkuCXEvaMeKnmRryqKJqmaIRJGOgZRJ2H+rI8MLadqGNBQpGRguVZtEf7cK
aWnL3SYCli1ZInyfemuE/6PSqDWT4t0xMfoE5X6l+T4T2Uc0SQTeQfT0hjf4P1EY
YCNomuzNdoxFqiWz6EeY95T5tDJ+3cdhlglavjrz+twVMrsIWs4obJBNP47+22yp
rg4+TXQS+cFm5MHHpBbmIQbE4sTSYpq5rYPaZXRAjOGHGBOY6JqAwxMHEBwrMy4+
M5lIWvtK8QYgHbyeT2yQfc+Co8h07hEXvS2KHJ04ttCdTHQu2DxGKxKRa2friKiU
daY+YeoDT0GNxkMHTzaeqIzgDZjPDouQkat9nx1p0qd8TJN0vtuHeyJ5PCLxn5Oe
Nc6hw0mCmYzCoLBkhhd0A2rQIwNP3O4/hZ2UoY3dN3Z15Smm6TcsOovatGLF1nU5
zdJa1+niiXIxb3dRRphocEtJQ3BOJhpmR4PAylLfWzuMp+cdDLpgUifoFx4CN3k2
ZwodkUnEJQ4Tj5WYO0o/Swdg75UBjpqTV7ZagNGzhuDfBmlLokUmmE3vR90PldzA
8aXniGquBRsM7cupphq8r91I+qJrKVatD4ZJbcouN8K62UMn9newOLbtYIcIdhbT
RQ/04bQMV8gf3Z1uWBBHzHNHHTLm0+6AyRYj2tv0DJigvnA9OHFMSKU+iGcrj33g
GgjHfICG9HQxtmzNYkvIc9rafKwTgqp4RrvQfdvu9qFhFAe3/1pIRMCShYKEBpXE
rvfv2LNwJWcVJopwFns0Iw1Y8xlN39yxz1ro5imF/+k5wmsk8O/9fdm2V6rI3sNY
Ppj9a7ua7GwTkT+QtXDhvqN2e9WnFNQ6fuBNdRd/I+EAGGIAHQFjity4hYTeADRK
dZpVmXCqNfFHxRy2fliyC05g28XGjdV9WimFwDUvZ3pweMmBM8vyQ0EmmQGBOUKI
6TabsfVUf4atoM3PVo/+uzm3YKr9fO9cmiGL6clZVuE9rZDgSfoVKE/YsD7+k8Q3
z2JwOUQrNVFd/kWmAN7j/8CQeGbti1yGjS+w7S9l/L2NZOkrAyME50Tn9IKCxKbi
vm/RSqb8W3aw+gMhT/dKRv1wvBqeaR6lP/4ieNLAtLNx6mOvFqS3WYgP5P3UzRUC
X5mA+n6g6UqzwJWyyQ7/NWuJVY868NJSdsYvwZh6urIcUOsEFmmjpsdiK3xtyZ8G
hyav4hqRvqEx32Be3KK/A1NOxErttYsWDFYjDV/gOJrrAw42mH8Y8949yoU0t9bM
FLKPz/nSUWrSSBAUDkpJhOPXLvp8GRCPUhUIBRjtjUANhBo3ZBokAA534KL7tFxq
9/aF4cs3gRSTjj/rN4JMQV1P2o3SDuiTX1+S4AdXlPeYg5fnTg8IJ6da8rL7FDfm
2NYgDmdX18+B1hdl5O3xDH7Xwj/ywzovLr3CAME8XN5bF86zRxckxsK2c2fsL9Co
qn1bRim9EX6nDPX1439bnEw4QhprCrDrhRz0ylXmE6pAkrU+LoUK7AWu+o8UoooJ
Dxa28Pmym9TEh6TUhaS1Z0JwJnTv7ObQd/bqQUyiAM0csbB0FUOY/Z9/xcs4W9dr
iCSfhe+T9fEFe9Jdv4eZIloHx+5CZckNRRDZUlDKhu23U2ayxvbBSXFR9FclqVy6
EkAgPORlA1o7bWsGPGWcGu2yyPrrrlA73+Acelje5COBggmB8a3ZQe0CCJHIAiic
CsPXZapsj0aSCo3ToKNnu7bhh5JV6zeI5Zp9UWlBFRu6YsErznTLChJ096PEn6I7
Nl5OFE25seugQDi0OrEh27BEIVtOW5gtX0qud/EMcRowMWVmDFX6d5poNCvOyRtV
9XTbe16BHqxtXfXNrju8CoCmh8jOZYkmNomIE0IV83sFaMDGxfyLNuFxpWXs0HAV
yKVNLuGZ3a59DsxDaJymDwkbM+jD08gbxTQUvGZPueu+cRXk7SF6WwtgIN8ZoukC
aE3QjwSQNjqJCqrvIM147rfmQEtEJK9fLLPSqnf8CyAGmHBbruhDXUahmDSZcaZb
PRDuZPGed3YuECcs+8llldq7HwoZbVKEE33OMrtdX5uXakox9d6Qljft4oScEkMS
F1ED/cEBW2VE9ZgxdgpRkwhdIHzd8LQeVDjyuzRW6pU6yVAMcFBcI99yqggeDtie
4OkKHXFoChm1K4JXN4/MCC3HQ1FZV12CBmfkePGfiYbPePwxcxMGzjpygZatJmMA
HvylRP7pW0gYWqB8gTG9D8qGgbrtIiPaDlujJozuU+4C36iSjP70gz+hHUqu2bhV
f4eICpPRQb9rq3ZyDN+DaErb6TKAIwYJX15TJC+2SiGqJIDAZ6EQXu21amnUy9PP
iXe4J6ioEfd9kqhd3wsCYIShdiBTv1x0jJuzSokP04x2DhlVAECnW0a7wg97gJZI
3IfHmPI6FJURx0qrArvED/MGNY/2D6rH7WBbrWB0RXJuyR0agBFJGdTJucBgwEzZ
+DDYUZUHxFWKyflVLkXtVpm5aYSFdA27AG0zqjSh0psjh0o+yCRRmkGWe00mfAPm
lo0D3zHYi4TiD0HIRIUl4/ELTRtGee54cn+RQ0avlpsYhREeLHp63nbkwYDiayuM
2ReC4/noBS27q8hiW/ESIEhb94Y1sX+aul4F+swK5pxxlCAfS9t8je5MnFb6RPIl
PAQV+nfEHqd27QYC0pcT6Qt4FvAn9ezdOWI98A1OJcr8sim7rU7TpqSuWoeV+mUi
xZmxkVlbblX8i+Z6DCebt+G4L0Vk+eNXhnX/edQQVeyymjZObIM9qeGipyUei/Fp
ctHLHdRYNEk7k7oGWmqfk4RVgEQdhpyWsM+bAisvCneDGToZmM0ZCtNCsO0l9gfm
P+jvNx6xi8g8b2/rhgR+NpG/O+1PZZfYT3ybOohkB6wiqTLOT70WvEiwBbMwh6sd
l9ALVX82YJpXpayVQ3IokGm2AfsOpyrHrnsnTRRp6dbjCp0M2ppvfVcEdUq+tl+4
dZLtpyA3AchhaJVdzaMLxME2sWSsM+1WQtuvKJxo27fT79JQqf6ZwBqW/SXfNGMz
eo5/0gL3oT8G+0tXpraMRsQ3+/DHoA/jTJRrAl8p+F7Kf3G9kV01dWkL01elfjST
Fj7b1VrWnbX8ZDkpXhtr+bVfxYkGrMboPer1VdcyPXU8Z1Km0F/Y1B/6CF7cVs5E
1CMKdTCLgFNwNyZ02R9MZnsBPvv6uHsvJukn6Xk9K0VlHxyylUPZDZIHmrIoCqMJ
9gJTBEPyNZzF0MgEtO4aKykptiD04z+MhC71lRE3wESyM9NLnMxqlFwT0QrTkOvL
XQdiNkAKx4fCFHd+UOE/lya13ACjKp56JFTXx5FKmg3m9dz2gjcvIuhmYHBzE/zP
Mps9Co1RXSS1/I2b2XvYQ29FO4VdOWzgYNOypP030vtm7Vyts9e88d/8FO8JqrX7
PESqv3214qGt5n6o9Y3Sv8qCiqljrWJwjVMJ3v6A0mpuVZc9/X6ja+5oDk8IRBBX
jRlzeuRB19Hk95zB28nAZ8eKAVY73cvezre+dV20SBcBOX3AFYo+YPikq11h18TK
1MPZCM3TkpKEjsfi+2ZMvwedQ9VXQ1q+iMhfuyuAMIinrAGIjIPRhpLb3wQ4lLJq
mx1vep8i9GOC3e6bshpODYG5WlWf1KCNb7PgTGuo5AlOD6kzUrW7JIXIaGQN1l8v
t7t3hWJGCZseSbl7Lao/2xm2NsbVDIEJP4bB3jpE+6SgjmK/z1KDIt41wymaN99c
K43Jp1WK1TSjTzUHJR0kvGQVa27zYz5KEsd7CGCS3ovnBLypCS7H86QRVAwCoy/J
6uovv6lCzY2DAvpXtehDabY36ToVh+YvK+0/9Q2ehNMy0dDurdKkErrwbgfBHQVF
+G9GTOlTfFUUo5Tk7U49UDaqGpFblQhY3po/SlnMXjOMJKzysgFhdfg6fEjOaSA9
8p662t4RU/43GSPPKDw1fjNvq3GY4EiaJbMaiL3ya1rh2tU7NL1FDz5dUtU0/tE3
6HDFAT7qKPqIu+b4TZZY6ZJkSN772BDy3jQrGA0mmO3/DKXsRtQUoTwfjqd14etx
tejGjDmj1RMLOeIv9LwR2o/I438OdHdIzzIDG2lbwI8ao7sKTXe/xhC4R7s98ELH
BENolxFI8O03YPdcJ/U17O/fQKUr2qoG65p3VEZxuGM/nNxPmfAGhhk3mz2wiwSj
tSD1pmbj7zcEEEn+r2kvMRrRhllk29m3YmLiEtlr8eNpfG4+uKZ/Auc5jUqAB9rw
CN9vKQDUo5HfvUlbYRz6gl8Db8obCWz/IKbf7NYAzB3L+++2XRZyZw5LFRxBUvgR
2du/cY9Al1TNmbLSkwqRJR42JODbsbFB59z9nFacifHN1pj7huf3cQZrG92oTC/W
xGNDqVhLui1TeBJoKmyfZcw72i5b2ktU6X8unRx9Wzg4h18JB6G8+qRkg4ejxpud
q05K7ktY7DNyZLE8/3ESpzA0YAuFkyU5Hog1Ifbt7dLv2EBizBvxGEu0YzzkfgMD
JfGwNsu9aEmXxzCFmGcTOJNpuKJKJoSUWj58lsTQ5zy8IHl33jzZDaxI9vSjNTCC
gjPo6Sht4OW6R3dHsn0wo9K5bXCUeceseIbDbfa3YLUmiLlKkHjFLa6wQJh2m8TE
cOGsBtzvcqpJhG5ceyHw6dgoS/F+oi7aA6/asBvl+D4ndL2bRdYt2mGc6bkFtX+f
xvBmVP69rLYtPcwqXftUEeVRrgd+yM1pS9z1Uf0zzYrh+8fyyhR3JQL9er5X+vmm
fCUS3eLq8AKAcPBC7fKGiA3GEOa7Zuq4FuGRX2NsQNIsi88LOkC1Rp9ziw+igGoL
wxycMqGVLqsdYr17NQcgHFmE16v7gVkAnDZKKHP58M9vy3yoPQc/nxmOXbXqmQ9Q
2DLJa3rXa7tCJovBJx4MGmj50QhspivCoGYXs7OexZcmvmeZduLB0bhJmqnh8W5W
tjWt4Xfa/Oyzf3/SC79030LEvXuLHBVAKYNEuBawkjny9teSw1VDdbBKGWWKLY4W
JsNoq/9XzrXrPuLcfij9hni0FRtt8Vx23beFdZovyS7i90siLqmXnFr+ao8BFJgg
DO+zkylupWCTs6uXgeIFYMBYW6Ngs9/rpvhPX4rpTf2ATxWZjzFTCB9zWjls/82L
suOtHls1hqbHvlmrEdlilIkaKsiGt+6iR0y1DpYyVd1qla4b91NJiVXBFgQozPIc
Scd+AcWLbSD02H/sTofjtrYhNK1p8PvK5V7uatrvorwHAbTwWgmtPgxPIeF4G9HJ
fatLEKXWTd+L1VXibOo9vJn+RCvQTD9uwlu+dIM0vJ3qnJcaT6dVY0Gu8i9RApMN
R1kDBGLe5tzPS5i6KyTUy4lH0HKTCgEyVVuFfSfxr+kxGnkZeqLC/vpD3VrTHuSj
KWHvBwnO5jXTPbCa3lUpJof9ZLYXx7E3ZBhtmAP4nQJbEHXps1SERhxTM+hWyHe4
RyJRS+WLo63WJli9LH2dsNgJxObXCZx/5eq+O4wDUuIq3pnJwquG7EX8uChvvnVw
vb6rEUrLh4MkrCG5hcu6nlXFKKhSbgJZ6G1DTKg6N4zzOy+eCoKshVWjKkC6Il8v
QI2tj4uQkclnxpymAu+rRiNQtOf+0FoRmkamrpL8DZxUv1Ljd9/jBslJBDrliU/e
w4NnNCzPyGWZ+KN/vT9kTd4YU1mqhy9a2ObsPxN3OjmbxgXupaAKd/MWVLO0GEPJ
9lZcSBPVMVvcJjCHIoIBWOPK9iDn6YD0+iWAfrXXmePG5FkUhFmYSUnJzL6adNe3
dzvd31iyTbvFa6MFsQ0wE9weYkC6gus/U6JYcpLnezl0RceImtnhgQLCFy10/m+8
FjVWx+UvLosLYQC5Da/pu+gcTpWEdYYPix/2IycPNz6kVu84FAVRpC52FU+V652F
GBlaRo6TZ6W3u4py2VWodgjoqNfLPzUXwfVYe/KuUcb5475sYCP1Ueu6v8gsYRyL
kzHV9u3vhn9ejmS3SzcOueZrRXuX51+8vuHMegLN98fImCxuQJmTniBkUSzPrZl9
ZnBPvhvNptGIl34TT8RKzNO3hMBlHf42+2EQ2B6zFIinBj+bTKywgLD0OXkCcJC8
KPO8hK29xgzYA0yyF0lFoZh5FSipS1G1aPyPPBTAJuR/59GX7DqEuFZzSX7p33WB
RgMDoYy8Nk4GBpwKyYRhc2Nt/wAiC4bb4+SyIsxmIOhNw4iaG7BK9ZtcOWZ+KSgW
vAIhPmG04hmaF30zJe3mXSBjvrOricnP1g2jx3BxTAAqHFMshar4LoRkiHcczDhM
Es7Hz9YkrG4kB0F/FGJ5EbJNbMt2PTTZdwPnpsZTH0YiHHheit6RS5b9Bf3tNy2M
0hvVwesvd27o6bZgxf96EYWjvhILiK99qQgbfx+4sNmdmJ6cG0EUdN5KsFDGSVdt
rM8nOulutmVWf7ImtcevMldhedCWLOfD1yzK0A07lBT0Hhy/tbrPIGP5yKWpnaZm
32KOFvYwUv+33fWj8P4vg3HTz2hjsYzpzWtSScsmR4zczw5hVGqwyuX4Xg7fW++h
E678oqVTVgVOt9FdXMje9U8fFQUqyCMTNYouBsABs7sq6bm7hrBf+nmtCxe3uSdb
CQCwEqdL5VqV+T9hxNPSlBN8W1e2fTQe/zv//WbOpTSI+4uvA2X6R3LCyDk2uzv8
fnkFQRIbC0SaeEpDtvTDUJE1eQzt29L8SaSl5DAniRS9pMO6DDoJtsDqc2Ed7klS
cBS7L0sGnCxi3mvIpcw5i4u4G1U5gfJSGZDoQ7kGn7abEaP8xPE0Sz12Erc1wIXR
uNEoN8pCuBldbKdKK3P54BP1TMRcycXA9tuO0X+3RtNgBLDW6NyzQU3vka0Ssrdk
0yMx1NCqaiG7t1C5Bu/JxovpIk63N6fW2z/TMJY0ovWe4vSQkOm+1pHzEkqCmUu0
a0/KRcg2Zw0Gd8Tmd851p1f3wGCpsDRc5ThJD6vGnEmHMTstQ/0hlgggA/KY1lAx
gYCk5HGhzFjFlbupB/Fajk9/dYQKNy700D5zgdvga2ePhlYv74ZtXnMCmrqrpBsA
JyMTnJ0w4CEv9Xsl1StrTn2OsxY7aQwNAD1TomCa6jD4d5mxZ3XnDrcbzEH2mazT
j+V5EmmHd/MpnyB1g2AE7SNUwYVDmWtnsqJU6TQNiRz0ZNWP7qfjvp/574M1C620
W1EeYx0qw7hfSMjufOf8iyGl6aIqN2BrFlOjr7TbHhDVlhssVZNeD8jVOUmWSpLj
ga1KDu7hdD38OUauj2/Rexn4heh7CuWnAsA418u63sqVz7+vnU+mZTcPTxQl+Pj9
kIFS23WSR/NjXzl2+Fde8qAX+GvzShXL6+wqN3vC1CYlz3UCUk4B8bQEGCE+uJSB
9WoWHgx6U/1x5eHC7X46ko3D+3J1wrDgd5gcM7s/tdJHtnz9bryKqyi9J51y4S/f
QZQxRWj1h4LSr+0ruPjfgS1JyUJQK0XD4oYoCLiTDKeb2odYdzjovImLp2h7NzSQ
q5xWfuIL4HJ7IjBnmXuM2uHbOYufVB4r8I8eFq/rM9kMNVjWkjtw6mGs2kr/HIhT
MKSoPPxXCgn55Q60jLp6nI3tniM3DeYM3hXgn9Zjufy25Px8DDRNRubHBP/mYJRS
/PrKP33hkExnWsNBJO/FkMaQDQD3Ny57DOTQthYDlcSg+/0fld6CXtGsCdctIySx
yFDqzzCmDQ78IqLgZcxTm95y6BhwhRkD4CGYRHMV7itMoW++CKACAeFDacRb7yQb
Zzlp9F7QrbT2t37vktVUWMtghs5us7E48u/XJ/bSyy1lONGZFWrWjlSGdnjGtsme
n/HndM4HxC/MPm+4ghikRsJvXQNFCWVr8FmvjkjMhZ9S13gVSzFQJSa16FyY2bgk
RoY/KFLkf938gNh0D/aKjHdej4vCe3+ZdYFrmU6kQeIskVhSWivfzvoJ6Us6BT16
0lZItPe8b7/UGvBaaAQbz6AgtuIadJJlqEWBUdYiCQrdoci6d0Rkt6AmGadQzXt7
RzyG/ScYDnT3RYZWzyua/mfNstpomaYPfDPss8+bh/GiCVyT8okoSRGTOZqGHbgi
ejYPhtOkJ3zxrf3Uxo7U0Hj7mVb3yK64eieqAAj8Bm7GTIa1dVm06ogK+wz9N7xz
TsBDQn4NAxFN3FkvAs6X/jjbqTTrdQOezUTSvC95qo1+yXdkwHYovjIZT2bap8/P
v4JoHuMP9MpPrennkW1uBEfjH0OQDTn8avmt99fl7JL+fBpFdx0AAn4G6GwpCCfV
28p8lH/XOJjqvGshupeuWJp2fpGBXkiHDYwJsYOnVC4flpfzmRPG6ttsUNaaDWE2
CeBwsNVMw6wY34v7dRlww9zWMrFBrn/ABwFfqId5tmac9fRV3RJS4DlSORh3sDFh
hAz/U1HioRacY+rLw422rjyqAYy1abRthq9/yNt7qGkCv1uDHAdQsp/Q3RCFe5Dw
B0S5Iy2bsp3E+G3nNIyTzb8hWaAwzBjHOv/Ox6c/9SuDJSeDTKJCj0NQikeo62/L
/l712w1qBAy17pVe76CEUMTOymQAQM0aT7Nyb4kKOT+o0/nK1d7cwNlnxvx02NC3
L+ttViNrJ9V3zwN3G3hyLkuWMtcBiyjrQ1/KqISDy98Ivv58kuzcN4bHdHxidIUB
oY2O+6fz2NHtOqjzAzfQaklhzNMLtcMXwDuuntxmVVtZzE2c1tqoVX/G/ia34hIi
vFDwd0wtKfZYl5qTFLWqIzI7icuSiyMU/X/MArMKTVTbK+DDcMbpRV9y9zrVvhtY
/KRFxD6BKJQS0UFgLo3etR4Me3PqJmUXRR6H6+DCYPfvQX6XxypYeyBEIn84bw6s
ZxobiIbf8VvLbg9ZRfWdGjj4ZbBTVuvBoCGyVuFap5TdYM+ZyA5q50/2pmmTEKv3
m9JENqtQ9SUA0l+CyWHQ+dVZHTERATOLcprv3asGUsZDJ2rX3RKjchzUZECMs74c
XMoXZLFZtOJ3q6njDDDnQaFvpmCSoPpmj8eLUpSvvHDqXEArz/jsBAVn3hPQWBEO
WCqcUl1/LN4pKJWNs0/e9zp6+LtuWuQ5B/URKXttPymeE+VKy00xJ+oHzUo8Nf/c
fhk+ceA+j6K3RoOGynfsLov/dTcaWbBpcB2+iEEdtULobSDlJ3+xNYG6ktvbsqAu
jeHs9MRTuvT/L7hdJhJ2EKYGHEr06rvHWDEpKoAJCMRM7/h+kjlzjC8tFDcUITjt
m+u6nFkH7meJt06nmaw68YrydUmj0OvXKZp0n0BTD0ecVIcnhdvP2meVCfLZDZ6/
WNPiN/8xYuaNBkUm44bDjVEHWu6oFO3e2hUXUVF756xYb7nvm6REJX0jLgfiC69o
dl76iEqY/yMc1jgiCNbGGy5N1FSC5Si52qVYAsQ9+yLTWe2N1ARXyD43SYgrhPHK
9as+HZXZ5ycOcDk+WWRYXNGIrQ3dNgYvvifG2DGXNx2CPbRLm/VUEpg+UfZdJD2r
WiV4qA/2srZ7PqNb9QIfXgoOF3+mRs1X0+Juy08/oaNuJO5ZtmPm6l28buf5Ux0e
sM+dl1GeT1TtmUNJ7cRrpeUzb1I9OAYpG3//irlsDOHF8MkwVmhbL2QToe24UcmX
1k0jwAZwMUHFh1VvaxiJxU4LmHvGfk5F6QjI/SLZB3Mes6zoZTuK4BPnNmi2KM9d
tisS7c2DNfTLXClnF88VEiLJzrTtNjJ8ZbzDN21Rz8cbX8GII7GgK0IoC7L7Iy6Q
aprXh5N5ointpbHS/5qibAf85EEcJrXQ5HRSDcc0fBWjjEJEPMGMNBjSUvgMvA1Y
6L4GFjzVUcVfo+atsxNVHtfrdGsmhtYUTNqDGL4iMHpJ/0Uhuo0bl2Y1gwpxtkHa
fMoiCtNllyMa+ghWX5vL8CeQtyHSEOsRVP+z20QeOEwRo4saPrQaSei8fxipb4oa
E18wtenh0DPurSwcfhYX32O85JgOgzCusEI9weKXIKE0kGUcH0pKUFpLisgJc3DN
/jzRKvH3W7rpbqB9mfzTLMTcz6L2L9wHth5/fkqSEVKGi/rCVR3CyRQUxABmjXMI
fwziCBg0OzTn6myyy+pXpw/5d3xNIgMITpCugsSlj6Wi6J5JBGz5P89DAXnbJTTq
En+rqnNEZc0hmvm+R4XB8kj0kzAZL93dMpEi2r1d1TFsRyBLGfXA1kLuotQ5THmz
vJoYK9/qMkUsbE3l60ZR0T2tj4Et6kLewi6+Vgz6Ym6KgkA8QJZmWnqz+jGvOP1/
EoIj5HDMclxZMkpJNIJiNDVJwGNjQDDYCwKejxvBw/Fdj17i5UKO1RRc5YUp566N
X+pWtxy0TPVyqd9iRL3LRz/J23m7ZVf/uJozomJrrHyM6YM8RvNPgftLVfxwiALz
cfF7p0AWbpfiMH6xaICd63XD/u9k+dGDcA/lWtK3Ub5xkTy5yejna1TxHISgKeay
ARzDueJx5aN6KxtuDAVksufGGOygRy06A4XSLtXaBJc8nspA1ewyIGnCxhqyZUoo
ahlMB9rU+N2rGU45ymWWwz8Pu+Rcx2A1n9uGt5ewUDeRxv4qR+bF0kM4jHx7iTly
HVbSeDdAfWIvdVR+4xJ37zasUA7I4+9USIlKb/F/sa8fyPP2lZsZa65G/BSceIQf
JrVeGs9FHbN+x7v7jXinb/cVuxv+vmvruTYJq5iW1nh0s8YmbPD3ikCIOQ8o3c4D
K9UJUyUWL8hXd0qsytMjAeb5aiYhYViacou9FRYWudAO1e8cg9XIwoxU1lyVIBpa
VJMUOg0TcjjjTQG0XqyUrYWQPBaFztSVozOnmtslgnSAYdCgGepTbyXje6qoisMy
kl4ii8OtQupomloYqlGwJF4otrS4PQhptu6lnckqdduPom+KvQEYsrXImjwqA2Cq
/6wi00E+vbD6JycyHLPtyD24NxZfpYJjKFnL/bCaY2JX3BTvZ+uFP8J6yRnNY4cl
eBJKFuihata+MmVIZNK/Rc2PYTgynvDD0VhTCXy6HuTwCefhJGqSl8XhO2smFe2b
8JT/06kHq6wo9yiy47Q1IYN1GjwLyxQCX4u/Av8n7sQJNrRuT0CqG2Kmc6UPxP5Z
yQlLRZHfBvKgKQtznPJE3wWtk85oyv+STBHBRHNsBo+aqAV2yw+h0AJ5HTqjWBzD
khYTzcnP9u7TyaPgFh+F7jo2YP2Ba4LeoIxgOjGKURUgLHiNWEDP4T9kTg3d34fQ
l6OGOpiLNHsgoUYPlbV/99j0FlsSUwuYqVc8pFGyI5tC6G+ElMP8Q/vIk2XElLvM
28koD5pBofghptvH+rtw23VFW5Ia3RdCNxEkLysIaDlF15fm17N2msZ6CGDyHG6B
jd+3KVXFrqEqrp9WiPs47lhNy8EumCpb3HvGxL3cmO+8KGYha9YFIrpt3RxedGFU
fnTXCice6AE+S9LB8gyA12G56GTy/onCcRm4BuL27/CgiOzibvqc6IUBbtIgjrXU
bEpm7vpt8JNbn0kWfYSYZ29DaE0oGzbRvxcD7MWlt6LrKbgpbOzGmqxomdOFGeyW
b7qC8qb4VpPd7sqb4I/WGoudIwTxjvs4pYmMGsaRHyPIx+cML1dDoOJzbygEsBhO
QMEcmlwd8SkPxW/cJkmxFYFYl5EyCaANZQHxyeQjpQ1NxpJG8dzWzcZQ76Epsouq
TtcOuOxcM0SIxrsdgsMVkVjPFyQ+aawacLmkeFq6FpfVcUwk7GJFgNL9G5RAC5P+
Quis7ObUORFa3vXA6aQlZN3WnG77MvgfqTrS9yf5s/h/3OKMK1POPM/TNp/ZID6f
HEkvNDMMPBRkiYX2bqm+/JwBBsL6J1vLkOgWeMQmBteb0ATI2/eH1mMjgSN1s6BM
TBAvvzrX4z2qYXMpbHYEkhupwsRYY6RfbxRNAOSkxUvXCbr4HgLT+D2t2FkWNx8O
J/BwZfRnLSB70JI/PlEgr46kBl+MRonrfyxZdWhGCRpNH62PuFyZBOPDoV3aR1Rv
kCc2cpEqFOLCUGiugIqOhGxdxyhah24pyhuBQVPFpuOD0Mpb0ZTkMmRs37k/YX54
xk5rpQN+zLto1ZQSCTF4a1MS1WhyEG7CYPnIFWrVm/6nbU2pb1bY7QNwnt8OTm6e
VemNMon2UMBVi4wk+7+lOPhTCnx0bMNLpI6zbrwnLhn0UZ9nCRl22JQrao0f82fp
pKPx+ZaOLEIUcnztLjBeYtJ7XAiBZK3sn9TESWnBGTD02E8zio5dMzKvfaTWRUYH
bOM+JlWr3jbTS1vHsIfx2Q5+XyFNe1RJmZaIw/d3pvBtv7t7vmO9XYy1JUrOkz4n
PKbLt37jawLyX7T/npXTiCDH5r/uDZwbf2rMPRV0y4sa/wca/TbBLH/E/QxhS/Su
91jIWqa3+HYBfJ5RVd2kUHYTBn7gKtv/0//XMyNfNL13ERIILTevs/vAwVF70AyD
Q12BvrfzeLv8lHuG0LbQ63llqTDnd+JlKU1toD5ZwD8xbe3CIVRgjARJId2S5jL/
qsonBkY2TAM+rks4BhpiV4EPIZfAYnS3hACuvnkNhzJ6Y6bpQ+IrkDqSuX3+RvNF
lIB8EJgXjc207Ne5KhJEZscAFJb//zn1XvH9ktxMOsyvR0HWIxG0iNNVq1V8NOpK
85nG3B/98P1/mdA5n+67gUMhz/HXGzZH6P6rbsF6dGLJiArzgWt4UUscKh918fXQ
c8Jd0JMnxBPcVWwxnZuUUAj8g1jpLJaGWdkEZFKINpcvByFpu+5w1GEdZnUU9o1d
D2BZnvwnLssZ5V/3MPVhIOsc2E41YgXjh025EMbNb7TEX9Olx+ezxY2jLg0NU8dC
6Cz6/Mgov+ecpO5EpueVCSkTV6CpGf78OH8vHBqwNdYv7Ut6vu/2dwrKHNcrDsAS
g47gCcN2/vze0q3ZGC388ijMWH7h5GgKNH0ElQCXUAMLAVmHJs0iw8g5pBnMTfei
vGTTLM2imvx2+F0xIRhTqZTbZinTAwzAuEFLN8+FteDaC+980Wd/chmdamOjP5LT
cVfaZh7F+APeNcwFkPTK9aptbVfvDVWWGvFLCe3rlLab3D3r/gpOBDMBLbAgceMJ
5McPCW8Iao9deizAwsj/zOxYWK5yXjU4o7OiHVhVHt5jHueecbozS6mcLlOvBc15
qDY7bxDKSuEGQEGdgXbDpUTHwmihKtop3aak7qFjNZ7tVFos0UOMT2IPi6jOJLPo
ZhyAawapX74BiG3udjKebHFtDwgnmArTwWsgHwZQyWFLkX9q/HvaVl6Ypzzxt2mw
OF2LycEj9FChEclNh17VUAtBGdEoglbFDoMXEx+Yvdp6U0G/UhFwum5tjVEgfW+8
GFfoNDuPT7eUEAfMpu/r2bc7BkJFoURxFYpW9aEqTYRbjZgkXJd5huB1Rz3fPUOx
vDj3WAcFM+hrixRyHw3Peqa4Uf+NNq6kDTo/R1wEO3vM1y0r8CLuFSPvc8UusTux
3X/XQGIA9I+GmSomk0QHPbu8j3iAZ4r2NUX6PhUYfs80tnHTKD5OLbKaUjsHnN8k
Gxsk90Rwe1WseXR3Uu2PAdaVHZOGOquFYk78rEKgz2Qjgv0xJCj0kKoMxcv6CNkq
C0LBzc+KxoYCi3Mv/5Asdz/zz3g9y/Ct7fHFxVuz/sSNWiFh47NZ0NeWPqmHfa8d
n8S9D207voeQWy1X3xVP2pQ++P41r/CTWAW+N8F7KcutXL9bBV+h93elVxFqmw7y
Z2q0uakWVoZA40u5LO0oMceUNJXN0ewuCi1ZRYtuGET9oNdJ/nrmLHeKlT/Px1yT
doi4CEKSMTrVuROraEHnf5GXmH0UGZ63X6qsj6sypWyBJHaYz40NTOJHRtyFIpxs
EXSlIvGvsnYZwlpem5Na0I7/47d335CCyQ1K2SPeAi05d4zyLulMnCETNSXnqBWx
7QVDEkL+t3mPMNYF5tU41YS6MlYKUOd4bP2CVawXYIzggz8I3dUxHHJ0YwiTLdok
1Ybiuh+k6X19oA2PEM64tXesKlr2n8pFVvh3++U0/+SQyRGgw4s3NORHhSoNgzb4
m659zLv45xXupqkvY1/AcmOf0nJrGVN4+qB2Y3tmI+/eSa5SNbuAaicF+lY7Hz4q
yPjTTAlrqneGKixTLO5wXMinysD6VJmTT2SF2MWVZktNzj2ImoiwZIxPCoz9XU9a
0Ul9kaMWLXtqaVVZOwHyHjsRK1x2KfyTyOGqlfquk1DZXwd27fs5RNEkebVIqK0Z
S4VP6pSgl4Pj4JhJXVcZtRubjBlmVHZjm0jbXFow5VUnHs+PmZNzTb7vqo+JFIsM
51/wHx09lC1kjCrx+V+duyfMimUkY5Av2Qkv2m/H8e9k3QUtPE7HGm+fgWdJaJy4
zpbn5Q+/rOT5+yZkguX0w0pD3Zy6TvC7OX7lON5aBF/u4TmRGkd/N/U/pqPxJzuN
itHr9lDE0bEB3bkl3bG47vOrjjinGgMGIIvh5n9S/Xzxy0Lh607syTbR2fdt7eSD
bKb9mWkGBJOVw5ei9yA8HQCpzfuxBDqX+Gi3W7bMvTRVXeGALjW/bMjkFBaL8zyv
1uyCcN9VlItMsIXoFE5SuEbObaaWEqZjcBdNrhDgK3FX4Ub7VbdCMiz13K3NCfe1
AAahJLJI1u8vJpQKH11qUMLtW1YjUNmDfvhRPM43b4Fx9iliSGxOVehs79lvieVH
yZifi2GDEg3AwP/Bv+bkQXwAkyQ9+zoaJqKs7pEocjuhqBh2G8y2HnnEuCsi5m2i
EN2+27L+jthbQdazVUjBycQLoOcWRyNdNGgRJFeLxxRKBZTM5YZv8YaV9l7eRQPN
Y4z/bzjRZGd6NfDu5N7SGZtFlV3ge7GOqGjl3QwOQ9TDM6MHHRHL35vy1agbRTPy
AU57WnUl5+akDVx68DRPWx0+Z2MLlcz5OwIiYE+Y7fPlwrmqj2zE0OX5ArsdXZX9
hMKSpHpoRiO3SQh79VinKYPfjt9i1xbh9wFIGwGeM/OIbFSGHEoeKOjATwaW4bMm
PQGsrwi6LWRkKgqryAPJoaEn6ZdFS1OEdUGohFEZlWdChCGJo5yrr0NFPUP8cXGU
SbBYpFup5HO9mdC4SAow4aoURFlFYwS7KBJ8yexqGN74VP2myBFeCLgoXzYj+Ydd
Si1wtX34jS+Rv13eSjrenIxdvEboFqjJq4eTG8ttei3X4mZSWTlUHQWsb28bSvQp
MT3aKfr1akP7WHt25dyCxf+hrq1aWdKQRDpsgd6etcELAkIZSmNF8VWRpiyT/1yS
Vf9oE8uH2ZYQAMWUW5msL1ZDwZLQlQJWTwymaZoDfcJiKKIQWvICiESYSrnhXrte
KYfS6kd9dyqdmU0iJRE2aEDHh+zhR9t2mU7EaHIQ7VSj/++kzo9XTEo8QHSniu6C
llD3EQ8qmLQz4J2Oq23ZDsBPX9gUu2UVHd2+pyKD+x00XbLXesFTrJ8mZRKPSN7a
jlmIy43/jXCB9XxcWfo2ucuiS5vCL/UlA0IZRc8CT+h+jh0YAOdNhi2r56B+lnA0
2GBRFSyfi9MmJfomBdG94vSEzp+7hLc8DjLtUqI4mlNGR3QNBwTxF7WibfP4asJL
Gjy5BL4UUtonlPsn/v7kjrfYuroUlYHszbam2IJAgYyI8s392YwZLhhhDDLwcalU
VJsfVvH7NIdHdTWAcSvyDywBztkX1pLirpRe5CfCgP17xI3xLsN2UOHwQNqFBX4g
XLF+sgOXtfUwqYzXsS+nKMGbZZFJI3TNqs7XUu6cT/4r1EOBLWxdqyApV5lv1o+w
DXeNKTA4dyF3of0ak0jq7Xjz8FTNtp6afaEduu3XV5E7IkELEngwotDqoaLHyoBb
DJz6wFB9LoxNYObqrbLN5TssDMGYDb1vuLCQh5VQaddydwPJGXhFfVSumhbVFR7M
N5QiMGYF00SQheJQhSHOs2fveFIYCw0Un/kDeTOhx2uMp6dzjoC9vBpwq23lJwiJ
9KoY8EBwJLX5/nnQCFPySCPCRVFoH7M4encCmUgh8NWNtdH0zNEbRfaC4CUOYcNV
c+BkWcEm5GW4DdUi0anXJ7/qk+yZO15mOF6F/W/yPF3a3Jl35NDUpCFOeS6RuMHh
wXPUEttX443sXkiF0jXe8ufoIMrr6xCTdOIUQ6uNn47nziD69T3G5lYhPUvbjzEN
IVxUveJINdPqXdxBnuvgir76otJfeiZ9HFusArkCCL/vAkPCUSz/yXV47FW7yW4p
8N1jY81ir99gV3s89gtKvA9nKgdF9wNK7f1pFjdOTxOQ81vSMquNahnbl6pU07+m
rRwPPF3nLKUSpZ4L3pj5Jd/BOh+CKa3w+75CqLQmv05NLSVil9bCRc+a0LY0cQ0q
mFp45fJ1enVUIQD8z782cJAaGQGhciBRxFESNdjqg7NbPyBlHMSr/MaTxJYlCXgr
Qx0cuN/BHeAKtl2wWCia6t43koxKAFpSqu/u1OPNpJVIikdMDwcn0+wZHZvJcllT
CM3G9iH1V5ssLWzykCphceusj1Yjm1BPXv+WphYDQktwb1mn0Jt7RxvVquVuaOtG
ahf9S4U8Ivu1SLhSp9uGhuiFNh5kuwlcv+bG0chfkQxjYSTibECF1w4NaAtnOMiI
rufc1Cdh0e9InulHOSBTWdznHMUIVuxZQOLxKw3DVcF481b/X3Kzo4ZLjoZrGB9k
agez84fWOEgpbll25OATyU4FahoBCIMCLle5zV+FEwKBLeaCrQvF1Wn0WbFy9ZjZ
J/nOc8bvO8/VGh3tuQrrRZWPJ3AJQmIsP1fRiHM9azn36un/aqXB2OdzlyBsO5wY
56kjPZdSCmS43f7MX61atnM9LoaMqYkSDMaEWZZloSmge4bKrY8SQw8LCkRORzx4
qRnah/eIS+PPXVYHCkjpPAn7JGShkiz8hAcpOllCx5yxISnCB0HpM263L/vXBycy
MBWK4A7XAb645JdeV1LuX9VacoYz6GKBgvDWPjb2pNjke93++pUtlNzY2eEgIx5l
tRzMf++kb5HeOdpMzLJl3+cBHJ90x2zojQjYxhcd2m1XLTfbzXFQx6qEVmsomD3u
T3Coi2EWMnW0m/vNQNO2oFAdM7ieACR08W6oChpQJnnud9tBge/Or47t62XQl/HL
FZZ864ifixJbpUXfq1YhQA8NqECrbWpAw5dvSrl1qsE+DkYQFyD2vd3R0rcqJwnF
NS11yHqJUCDjW5PY6nel8OD2vJPfMUMDyB0MmcfELCJHia9dW5AKot9m4rb4a84R
L2434N7UirQxXWMmBo2mJiIGxb/7dJ7YMLoYBeshx1vFpa1N/rIX+0PoFDMi0NMU
sIfZYos51slxPk/DuBCfq4g+KKZO2EhN3l3XYUR9v/nzpMqp47mnMrzpNiAvpeZ4
7kSkrZ0EaWL/jY1ii3PraTqOg+flWY/9NJtYotvzPOE+gsShBpORO3+CwUiVY+5J
6r9mKDuFNMXpMaT1eT3vuBdoIUlDfHgZIoSiUys7Y/4drTz3GxZlPg7YQAEQ4TeB
ysgA7fK/qvBwN7FsCA5+34nqYhfnTqRntCFh7LQVLwah3szmj0/rquaeC55HK/bC
JiJn2cMbV4GiuGV4sr3wIAJuY8YnD+4RuZwd+hIqVKr5ZdXOJJNME2PWdTdzq2SA
kDkvCahWzLsT12NbMFsd5L38bCPOio4nRnePjSrbIBL9ssX4KTXACAMEcHlKWNxW
pxl4F6SimeHx1gE83LCTx1LwQs/ub3IbKH7HSKXWmCaGy9hVrhKuHni5yNmOJ9Ge
AkPWzKVE6PrbkVUYm8iKRyGJifPvNK0Hn4mES4TnY1HOVOcf4QY1Ry4uY/FS23p4
IUJz0MsNf6JpddjQtU4gH4M2LvC4sJeISiZqnyijq95l9yncXNZHdUcJQEDR8XPW
zSnQf2ExtLR7JDThXhLbNIkji7p+NdN9vu1QF89Ge54iyD29VwuNhRInfnaopolo
J5qHUBjU7KCDuOuZCbFfftoWu9UMzMSm6OE7/iEBUcXKKp4jlumzVX4lfYW50/tw
xP3y/L7bzr53hw1DQK6bzuEnFPzDd7CPYI+JJPylcOMNzXv8H80RTN6QxdnqZ+Zf
11FrnHvoWCRGnH/ZYMFVCWzEIsuXN/r9myilrCA2vVcMQqQzzrlqv7YM7krToO+X
BIPCOZAMldYuFYJe7eeId8Ld4yQdowDtmF781ehY0ilQwoxobB3oDIvZvcy26Jyb
2+/lHB/lwbFOnIbH2TxTQUjMXr38G+4vrKjjukYFZy00Ht9kpb51+Uouou9QCPpK
YKLeDTGGKKDAxrcgKvboriai6jvrn0zDdaaI+RdX5uWFxvOawEevZmtEmk+5uvCO
fMdXDWnhcFnby5TY/bL6UlqQ/1gQ/+CKMqvPMDhEjjbnwaX6fsFdpx7q8sF/jzid
JtpFYz9YFDvxWv//BUciAaaVPzRW6onL/xEuO6wxvWqfiqlOKNqsP0GmiZkTmAwT
FsIjQu/eLue8ApaTBy9aTtWAGoDxyrt9y3yHxpVRuG9fWR3RsjBB1XZ0aoWPJJ0s
Yqpgp9ufbZ22jRE7C1ADDLRaikTc/xtLdyogMzfs25Y8K0HqDXXyIkC8W9c0+4Cx
YQvZD4w0RdmA+0x9HzlxDpKcD73bcg3XGw8ri/7Anl8/9f19ThmLeAadfdyAPScA
mkmXMfiodgGW5zJmEIJVnmQhRmdlZ7BqGVND611iguL0JOd1MNytdtnsjqhBZ6SQ
f0pByaYQjRqPwShVbkOm4MTe5FAWCWVu9l93FYkaC2p8ViCcjJw4N2fCXcXEMfhj
1w+PKT9t/4oU5SeZtk9c0Qh0cyYGGB0Hh4a0sfuyGkyJLHvjMG9VS0Pp+xbXOZOl
wkTt6fBzod8YVXVMUhIIOOZCDfvdxSCTUvtzszjpBP/LQAyG0Uq2AwU0xYrjDmyg
giBsVsP0JceexFecYiL6FkTdUN65A/iWKSXac5oWaOEywjOCifiNUf0NL/4qNd92
FWE6mNiHQJLY4OwhQW4Wj8CemLnoiNHCM4JfNwUaKjvT3KFccF7eiBVCxBLrBnn/
a/ptTpjFO3ITh5FXUcOV27nfJ6a0U3VEzL0QsUtWhSGm2zjOa0Dhcd3d3rqyTsNY
mc606nzwBhyHjyMAlZmGSdUGp6rneeOyGeV6pb0LSh6Wz2UttpO7cUY7gDkzOECs
A8nf3nBSCH+N5frKinSkUZLPpd+HHC72ThLLO+OfNE7RsGF1ePisungKlnSgCtJs
K1bFiq4kHNRUYvi77o1NGPlqc3ODvH28wFoHZgVHAn5+DQ6xvdQvdNaQpglO+cId
OLCWYUjwe3gRJcvUwdYWj/8FPyFlz6y355FeexRMW3JgbIcrIvINHIkehs5/L3o6
NfqdOGUI0Y49WQseLDMfmP3YX5E5hBSz/dtjCfAw5XZr6mn/vYfUouthByddL/1H
bH1CXs/cA9lrglnFrEK8i5TbmKPEJVsqO2KLLc300D9Q6u3o5JTWjKGol0S7lHp3
V5Hk4M4oT1e6WVa5G8NEwnB+RTz7IoUxYKPtC3EBHfB1gDfO/gsRFgg3Eo3TB3kf
jBQEPtJrupTbUJ5e/XT/f1QeVp9ipZ9CkBXbaZmJbTqXkpLyfm0SS3jTMRmcCmcA
vp0Ub1MCgHzgSwwxUX/78Xd1KmnXS6jB48rdWQE/z2pIX72IG9ExL/0RixzBKtyR
dWz1Yqj50NoGpFGJGe35zc68Lev3DjLUgr8zLhqBs6JwMB35TGcQg7EITf6Ymvrq
ZoKqRY7EORaip3/wu2J5LDkIrf5TwecN+HDV1CVHvm3KaWna9hbkV5qLMwwIDpzo
zbW4/utPX6O52b97isySEJC11Wynuh7Vve/2T2zPySQcW2fK/Mdi07vcw/DeaZxS
rYOBvBf6wjZP6QiNSq6zIY7YPbQIXeHTF6CLXd+UsKwtZmT2x6dQsco8MlBAjXR+
G0cyDD2pw+2L5mBAofZO89vHpd0vQWjdN/okt00XGeuUdfTbSfR/DQhLKlXtmSFo
pUDkq7x50k6N4A9OaMCkIf1GJPMvUL2iiYeXg2djmIFotj/GpCZuW7gEnnFbN1AP
11rM3yJAvKhnQNouJIa4P+1Jl8E1IXMjg9qFAPySwiJ4IZQSuJ2OwzA5h/fsqZHS
P102oEanEYUOr/K+HfLMjp4fOP2/ojki+kb+3YpAsqKfkknmEVwBarpMgZRBDb6x
qtCESUh2k45PwkWHJXPMy1eUMwaLl9vkcYG/7/UzHz6E9K5dIVQK346G9ps0iruu
lw9p+IwiMvZprqOO4zO2mMB9gTODXzN9eRgjd0AC62yL1O5HxxtwN4gDHa1WELi6
WM4eHGQc/rIV71+uHn+X7JOHOLcHP8koWfgvGYzoklfqS+rl/2OVFUCwczwoX69Z
Vkqy7pjNEHdFAuOTWWQ1XRixGkZE702LKNHM/iJYzklpaQLfY8UlT/LhyudhydPx
5dEli6FPTzJ3NZTsDGW6WKsPIfin9gxe8II+N7OmspXeiICdLXR+1tnjoRL4LB1J
l/vdD6j09kzhxtF8quElCf1MdpySHxz12TiS5nDVotnOowzGEUPanQoeauaGYLPo
ruhKIE4HZQp30pkMuqXqh5WfNkgu9c3zacN4CdwroGIyxV7rn69nkSmvr+G8SqQF
x9ImNx0GQWJBfuPwBIaHkJH3512CNP7ykObzBD85neNw0LwxkoomKzHmcDnUpYA9
oGqBUTdNTzX5gOS5yu0BtSkYHERm4hjUKlkWYfRIIKMUNU9qyqZbgSCqiNJlQUhF
+Y2QgFrRhyK7iYAYHx0I8+uOOIVMlodF2HJz1BA0BmFV6wzsGUOKlj47EQc1LJBw
0xCQ3JmZqgldXr03GDzdmnl5OahRz7m5e/3PARHptT+Vx0hrs8Xhw1XT7NeZdtMq
VR+fyP+wTpEiceEvaYL8a0SbgjSL9OzC8Q0BCTBMHxv2PUhf92knRFeSqp3fHQ5/
Zhm0GXYXLLiLzg1PYHg+giDN1M+LeAiHAdxZJ1Ihxooxl9niWqDTX8SNjrp+RNEB
pdIZFcj5zk/8hh4/a5Chky7mRxS2+na4E30fmbNdhY/IojQxEmuZ9GV6+9gDkgE+
ppeBJz0GNVDMvpGPs4H4pBn9MOTr0XINO1TJ0FvxCwrDHvodjuxCrEa/HIbMAnBG
0m9WoR4b6bh7GpJ0qzg81I50WfA5idkTLkKN+BDnfBMYDwoM0XBqJpSpc0Iakc+T
7KS+jw3vAisM5NwZxopSfzh0DwkkK/212sHEyOV+0HpoYmXKsdtgAeanLKHp6X1Q
kRICPJsgde4zfyR6YPRRBKpofh2WJffj4FqmNPPrZorNMRWvr+63DTvkaAObvUtg
mnC0bmQrDXW7tU/CQyw0cMAJ0Yw/8ROC0a0ItItLZ/zQi0rlSb8HdMlbOhUkOFNf
GZsrp+qZhgB5pqiywCyHLmnjRVcbYSF2rbiJqTDsBVc/NjECxHATf2/2RJcRMiQo
q/817PLt0MHDTTyn7HSR68KiHZs6uv3WElwyfhfVbf+n/aDvNB1gEPgY/zUwFJL4
qR292txwv9AM3cp/vnc+H+/EVXSJXzPptf6JarIJlAw+ivGNpSv9tXShbMPOUGZN
PdPkbaex+3ah3QGmeHGRoyOsyw8tAvQ8TDKPVUp3FtSD70F+YZkC3qjnHsiIuRRG
psBSsyIeDZIOMCvlXLrZHEpsAw83qCy6NcmPFeug/qjjkr7EiqOv28lMaBz8v1/4
9nxnRn1wV0TWT27yiGeG23pIc90t8prDQMLixgXOzkQIgtrR+gt7Oad8tORifT6p
UjM+t8m1yQapy5o4qBODDl1jlD8YydU7TOxSIxDl8bcHC793aYWCrYja8t6d/vqm
SNGvpym3oXB4rUPaYOHC/kP+eyBtTckLN7Zhgvx2rrBAQU3m7/viv9Cm7Fqnk8DI
aP62xLPZ3+Yw40m0VXuJQT3SAN4Wfjq7A1t/7VpRLuIyYv6XqPbqUbE2NFgmnaq9
tCv+q+x5NsMPthF3oNSfCSctJna+JsXa4Ip2jHGdLTPYpjGjhT0v+NQd837L6RmU
3iRekzgmTk1Jw8xxhj+ueuBNmNmCOHq0KdRkFhQsAjhtZrK5o45Y1ce4QI6Va0RK
fHT/bAT1hJ6+PapYpuiezlAM6mzzR8ta6NY7CWFaR8qICFnjqCMK5EGwk5/a0BIo
X8JcuLn/zJxILaXy6v57wQqqc+I0UuhBj4ptuV3YZ01gzVMuCHUQRT7HnH/9Xh0K
KVExdr9Gb0TaOV9mU4aythf/XB1E7Bau7EQ93pR4bkzfJXU0WgayiMtDcx074Sxw
2HzLSr8GsZmHk1ZfJIBYv1TBZk/QZOoQPQqFegCQduQwO9VKS41LXcVNzEohVHHi
fOPTdgAgZxbdT7IeY72yDm3uKSO5VQPAbhMIO9Owp7xPRKC9ave5r5rRRo8V7YZ/
+Y1ywegJTndQr5zcj2ee31+lss4FgBqVDTOELrECCXyDPjK9xks1DD18PBiXXFXg
jViWZobWQ2xC7kVe4RNnua/C28BQAUGVTswTbDnQlDZJTmrYoSUZ+MM4UNMgkD3s
gh2eWcq0CvwBc5TjokGJS7TYwG0EosEj1crjmI1vULkNkeD/4cF+hf7GqAQBCUCC
tJqmclIKIWfDsypaWRgJYSEOazzQvWmYt3WB+dCfLAhmdq9bH3mOA3YseRmALY3L
PRseSUmlPtQA+oDcbBZIejvyFcQX1jUZdGry3I7uWlSxp5BV8bPZiQ7IxhkI32zP
XHDWrnkVFrbjAEJwxoox334/TAiSVP48oIoX18Ivoi3dlp6YVY7cSO6ua82G5wRC
BBJ39UNq9ziYfFNYH6Z0p/SXiu2AJ4SZDjZGZcZYxKx1A2NP2Go8NHBJK82WXxxm
2P3OJgpwhUd1UBcM0Nfm0XIZ0EkywztqBhs8B6fcS5bP0AfJQwN4+NU0EIRnDiC/
Xno+Cj90gKzZPkpB5q2Xoo9LJlEhTpM1CmcLDOeIgp3VAHPX4CQzldKF8Rcq6x9u
M/5JZdo6Ekte3Dh9HBlCKRWAHsnmQhrj0SMjZYsiRHvanr9oLQqaTSnZZTTFMzom
VbGME6SozOX3tvFIw2GUrXpqw8Y1i3AXicKDZN4VfiSZQwl/MHkOtRijzVr1fKPB
ObR3LxHjq/w2RHu01mLuWisGq/JtPIZsStNvySA0YB7tZ1oSf1cqIDm5Ih2ij57n
WpRg2XafQ0Gsva9T+KhlPqouP/3uZ/B+l/KrfQ/aWdLvIDI2qHtOxPxzGEszGmh2
AlGfXe9KmOvCU9OJuw3hxqrurnV1H6QHKGIX08QQdBi7Zc8GUQLAEWhdpmK29vBr
ciztulP+5PBD83LDznHltVsMl4jyrFqP7PZlL7I+/us3re4Gbdle4wfX98CuhGrv
WbX+7jFJG2Ao9dOl81XW3dYS0DJ84H/zbjBtLu/w+lWGlgQiWT79SYgt9sHmgrYs
jtk09il8HTElBckIV2aGOePKIgxJsRWrmhXNuxAxIGLjit+S8lZhSctpJ4rnuUOB
LwFDD2W6+xhVsSGPE3KWRwExFyrubNCq4xYk8FcQpT16pI+iJGJo7+gmjAkj4VQl
k7c9F5ycV1Qlk8ARaC1EIduddshiMKMd4BwuXGx/bnp87SxmZbmV/C4NbI0UmHZX
m90qvGu3pEl4J7Qx2LO7m+ffuUz/EzkMf7VPPw9NvFHADfh2abac5HY2pplnCJA+
v3lbLdANw6p89/O379PN9X0F219RJyYmwdF94PAfEx7YDa7SeyMRTjQlVpKnUS1F
Ucwd4SQUSt/0fi4796+DELJvzDLs1TvhK3tW6HVDL6YtIJhgKmzSc74h+T1NU7YK
ada45NGypEcOQX41l7jnevlEQV+xlb+YrpvEeGYtjUKLy0+wEShS02dZALWzttVr
aaXYuYJkXKlpD7SaV8gM9oC1f5+1H/tWcy9eTIfHGafhaumlnIjMNQlhmV15ydyY
PTaN7Jdu3tCMLT+5+wf3Y9NQyCf4odHtu36wf9gJtah3WblTAWCzIbYUPwnrxjoN
/YOqStlUesosBoXiTq4bmKKV5yvMj3qwwjWg3jIKLmsegFsbFbWMzN25YHOG/cbj
7ijEy3e2aJ7otkmiEUCTbCE9FYESjSWapwXNo0Y8ro1T59KYl9Omvtc0Oij9i+Ch
WKjHNmedtHT2gedAMUbYYcDhITjWnN6PyR7KxDn5L1ECBfjqqw/vFMUglgnuGsg3
sOe++tfR4STbGOhhuGTVWskzs+Vb+8VAUskLkU8WgdydcgmIIRD3ls2uxc0vRgTv
bjwkQL89aF0Dnz858t9m26LQNGPqX+3vcHvlQYE/kql/VHRnTl5eFOD5hbfX4VzS
gQ9l5uzlhXe+8rQ/nNbr/Gfu1E22eoCt5Ht3AwqvhwXYI2pVBuwCCmfME5JGM6rR
JMo6nagEdDRgc5nuplx6NmDiSy7oSMB5SfeDwabdDRfUgyu0SWOWZrJ13QfdLNXt
moTTGHiEUaeYSnTd7IE1l4L86CQe9Tw3AvMTTbXjKXC473UV/XJhkNd9o/QZFny8
74qFgUCW514bln/ayL4jZ7i7gX5IXQM7a7kg++yXW5MLw+1VG6rzRAPSnSWalaYl
agWpmBjYOuT+8XG9Rx8G5ACYuXBNpW++Ux+bN9t1/yqmT38BbvpDUIvU14lphaQg
9SQo5pt3RGAPh8VBUE+FyjV+vjiJ7WAPYWh514p/m9FqAwKRjch5WPXRlfzUoiww
VGoNBPjCJdoBcVvxG8zkO+gIsRtC+pHA+LxeIE7AA5N8IUqZfWhUQUNchxvHqcbc
J31Lf4+xelAi3GiS8gJ5766DS1OFD6AQh0NoFIRZZFxNzy3Fc6uqABmowK6Pdk+n
O4R4MCqXAp9gz1jC2YahaSossyYce8s5qMBg9wEwXew+yXHHmbRmdhgO2h0w4lDH
LvJtnpDU2HOvfen74B6xu/8rLnJCae4jY0tw+FAAFOKGJJVVfrVNMcFgz1Ml83Ev
TOLa96o8QByLbV1Y/LaSIRcoFB2TWCYUnRk/yOEcGskcDgcTyJlWcM7wKuFkTA38
tKrpZkTaQdhEna4wUeMFMca526XjnJqvndFOpZut3X98a8NUEy0TLqkh4MPnnexP
ZLdNEwyaAlRi2MzO8NEvYHS1FXz0WAGfqWt18h2sAUA+MwdApR0sCNXQdZD65wNF
dXEN2ZBPhsQ9XtmeUMCSXe2df5RdaS0zh5xYS7nUEpy5fArqLEYwOLcUEv/7ZSiE
0EDBr0AEYPOr6KQqkfv1jk7CmA2AEpwtTJ75yziTkjYaRKDL4iwUdJNB7dDsx/zA
0NzqXc2SJOXOVt7yTFEaIyYdmN8GlGN3n6BJ0jSSZ7nZ3cP72MhhUFALMmPxppoo
m96NW+3Aon5AEpri2gUM8KYk/b5jiT5hUQnMt+RMX6BFLkqvXSOrxoOsc8UpGMG+
FAvJq8qHMQkvFfzGHaJww7YWABiEGJO6CFbNL4Z1sOZejJ9pKnqZ4DlxQw5pr3Lz
v+fPmTtFN1TC2jJY02wYLraSj20owQChTq0x1f0Kmz52cyfOLwsWl5NAtNlHcSCB
KlhWF+5SkbgB0ucSvhk2dvCZXsTIFlysE6edd/vvTUNLczVjrYH98t1oirJ110zn
lUlQQOf2Nr+OtCR+LrNMDoYx6BzqVx8O9p9a+cOBuZMa5NRx6mnp0CoK15pfa60k
p/Qy31rpKsXRxqmjAw3/P54FdZ8DtAZDIAPhmjBBBJt2Yzqqg873N7tW8VDf/kbx
FOGmePEPwxh0MS/9XqRjPqp8vvwfOBh6UaAx7rlU0fdU21mpH3xgEm5otCrWpZm2
ttTrL/vs8yMycYxHrTc5pHa755rJrl4+bYxz5EpwSuV1uhnaZN9rI2yY9iYptkX/
T3xBeWy4ACdvCFbEIWVoRMVMqqbsN4cNIpI4x1VdmEBVs8mtO2fstB4O1iZrlNMj
I2nVGymuCFAHYxvX5JZE6KDTLN5kUcks2g/al324xH9hLbW5h93A6fbcR+YVG4bQ
VLbr6wuCRiNz193iJhy6I1Pngl/0iFRGd4rEeT53MWJwhZWQ9XC7cJrxrizF+tf3
+Lf5WE+JL++svIMIhM0zGiKaPwplSzZ/DVGyzNLlL9/Q91A4Jnwn/ByCC0BhU93r
JLUPcoWgxjBmysDTBuSQPp4XlWY+cofF4woO1M3UWv34eXuzd4iytbQdrWgxD5FB
MwgJzCiR5BbW1HkbKd32E7MQ73Tmn1I0solXt54s/y29xzQFJex6QUrpjY2Te9VD
7C030OC2lbIrCQhbbXGiMye0R5ZnYdcD4xBjYT2glQHFcS3MiN7/ootIrwQTJPt7
awsRiWJST039TllIMcg2D5dgf8+v4dkFi2AbHd+1mO1QlShrpQs5YR4ZN7FTWEFG
qmmignMdTRr1t1Oac+34BpxdH3kwYvSYmz71/j8HGWD57Epa9465T1zsaBcjgFiw
9ELTN/mtx+ZJXpRAxG80DeSSRIoFU3gHJGnHCgOpIJzyKT9sXgbeHZ2+ouRMiB4o
0bicxl/Nkk41aC0FVn+Jcy+zz5qxbFGXwxgqBWWvRvIT7TI8dVN3XEjt13azsUCU
52lIFVPnJjcvZc8sm5+WKurWAIvaeSiQCr3tVB+rPX/OEL5vTgtyzJB/d25Wc4lc
KYJBeGohIW/dEPDLaUc2kd9yhe9lPjVFE9x9EjSgkzjOMf18mp1J8PQ5xMF0b3ku
UkszdliFUzOpaLJ6dOUD3MrL1/LjDwnnjyIo2oaCj1gYVIAywmlc330NsS16FJY9
q2km8Ij/dAFlESpAtee7Lnky98bw8oKb0Z1eDHIO92tIxcOf/e5ALTN/XYZUrNGw
GC9jdhbtH/J9aPIolFvtk0wUyRj+eA9lf5IeyToIP+qEfVx8KgAifMOxnlNj9YiF
k1zlv+f8Z4qP96Rm/8KOB1eBTf3bEXW3Gw797c8qHajNoZwA2ZtVBYQHdE3Qri2E
rWQywbagYIeTSJzIaqQEMdfgXL3pnO5WtKssD3q/TNCpiAKfBZCd8RO26SWHqbeL
T/FZvho3I5NGqztrpU3yo37OAgL9MRxLrWR5Cv+36M08gy/x41LOsJgfywLr05us
KRByRAI3NVRiOMsZAjxQT9dN1pbp6YnrDfG4U+2i/zQpJXBFs0tazLu+FuB9Gg4P
44/URIxcfVoELPdJYCDjQRaym2qnwFqNdPhi6Dr/Aah0IsakUpfeK2ifDpPJijCV
aXq31TR36Tc8aKcCSN84MgEjUwV6dfx3eJ/E5BGtwf4nH3dc3EOXlfCu6hxwm1Gq
HVcyzyIdBr73g7ftijkYgu1prxl4aOT3i6JEBI5ZiKTVIjPrCMOld33CckceFxv3
FLcuN2nyni7Y+2490u0rFDKiKVCQwdhIAW5gv1Zm4Wmm/WBcGnTia+HokHlodox+
IDsaN1DSF0tjpVub6cGZ7ha5yUGDHo1GS+fnP8qbZvmSTs0QRbq/CsM4TyxkNn5l
y2h3ooJAuJuEf3XnUEJJlk2+oeGVXNvO6tj7hJ03RCm/pZXtBpb8aA6R31mAvVRP
BFafg+K/EqpGxL/umQEp92Bm8vlTtwGXykx1WC88n2vhLUc0DyyJYd1TPzGuGB75
fSx0xapBDS42RC+gWqCMpQaucBlUVVQT272uZgRrrCC6/95Ui82aXv99/QKx3v1n
54M0N1Iq9pbegZ0e8hGbZme/RapdG04ebNeWsD6bXFyzw+SvMFGY6zoq7SL60XWM
2G0yFlYNCAYX4Cbongg0ju0t5x2tgFVBxzrEjY8r71enZOLEp1xXuyUHIjQ3SnYj
Lc0sqkuZhgElgB28Amh1W4OYM88dmL5HuKA8kWUAiaLFHzt2Zt2W+hsON0n/0aNi
q00rR2nieI/l6r0QGvh+mDrVni96uRSzWlUqBwAQUsy5ycWrw0kMCtPD+Ywsr5wI
txq1jMa+8hysn1xdXJQnXfhPPmv4JpcyRKfYu1BDF3Z4ZeePiZ27NHtT9sotRvFb
s2yze0RWik6nXInoaxS9hZvJDWLjbsLvbPaxP6fs+tMMFI/b+AnQAEAzdmDDCnly
wCDAUHOa4Ur1SGOzf2UvzdfK9BzNIxVDOJ9uVgXJkxOMZExboU2z78xdAZmJieDz
sOFO7rmXm7BcFYP4jTUMVLG3viXGI3weGBr7S2dRyhLH7GM5oF5mfFmnhNcb4N4E
fPjr63EVWI7qCO8QvmvvDVibpFNHWVe/1fI9X1r/9D0vMx3ZIAqBH6ztYuMMpSzc
2OH6S9LBlusYOU/iSz4p39Pago/oUOSwPTDEJnbsns+Phnz2/rrR45eHyIxrH+a9
+LA71ms11ShXtCD9aLBpVvtPlHlG5WpAZ8bHzj/UoJncqj6GJHFrvJa8MYBlmR8s
xgMNPeBgAvOM4QUbw9cNXcJ0GbNuswu1QjxgYDtJXm25QEUDdpDJN4Bhnu32Lxx4
XvtOvdMRmnrihhZfPx4ltWUkavVNlKeAc9Pn5pVtGnIEGcGi+5fSJCYI96NDWZU6
Cyw8ArQeB+rsCuERLf21P1UaS8uEV76DpeHVWzCsG8vVZhXNoqBNDKxRsOweotwZ
EsGqVvXDXAlsjh8kZp1tuDTz2D30eeCMI/ZokY+38AFcqEag9G4+k72CP2ZL8OIA
H5XYUsnEm6dhpC0S0rbWdXnWZ8Yb4Aj8E6T5hFuSJPLUXWh10FUe9EJle/guKkvt
7dEkN/NEsDRwZQk9i3Rl3DCANyPfyZJ70F4m3hh979y/6lOU6sEui8jzMZrB47Va
mbYxK4UMvLZUfcbNdsbd1u+++5/kgIzDou1ON8d0p0yDm2do05fXNLBf4LSrsXzI
Ff0770oTHFZdCrhssc+RY0edeJSg1wI/N5xDKKE+hJPVQgb43o62fdlaPIolDleX
7BFkPwQA3+ww2EksaTpswIL2NrOhIToGRmEpZrmGk9ziP0IKWkeJJ6hnktyBdrRo
S5mJCo1SLbov7aypCg1zVZiCRaxkpeRHxNvAHIRJUxmlB735+hwkuIsrFzDfogzY
6ymejQtEIdvq8hU9FIBYHKfSnEeKvkYgsatwgPbgdOScIuW5qa7/3KxheF6SpcDR
Avr9AM676yHSwTGxen4oJo0QBdNDTJx1Gtu2G/sJPOeRicU47WggwMuNfEGWreNL
4Z66PR+jTlO9O2H0qC5XMA94nakpvLZGH3Upl+YkEYA3woPXa73qWQNIXrtrM9m9
5DE5+B4q7c9D0z1OqO1aEWW65tku8KiPtEFyTOuFLv+C3K4Nyumt976PXVnnc26R
/3Ka0IfPwFsHixLmZYkj9toVSkOndAkB6OjKB4+E6UtoUaVjf2Bk5cqExOHNRI90
GLF5d5tBRZH3YspHDkiHnbrw2huRdONFv/wwY1dQ+3q7NQ6BxltNlVRqnHiRCWNg
dsPS4064bUcoD8xtajpsRXMYp0I+5A0fOldXlLcj+/Ct3/K9aTWHiWLvbgv2ry6o
w3joyUvQoHLs+Eqxb4lJGIECuzBnSDSBCdjndM+o6OMAmwbKG9rnstnjcBhr8I9K
pJzVV2zDX4EXmtCTtTG6AwUZAcYfaEWCv3Sd/Zi8iWjVIpBJzGnmdboqh+Vzq9XO
7MLDuCJR3Tf08TRgQ7fS3kiglHX3BXz+R0Fsd0v6Ej3N47PYphKk+w00zQzzi7wT
kcEO7IiwLfbRsLURo1P9zJ+5sKJl8nN72ZQwYhsb/jgZRtmhQqBdoxZ8sNaDaO/r
TGbOo4obW+8Q51nWnf/3m++D9mHgDcEyjbZpKe4c8huvAK/fTlPfktTcZku40aoe
0grE6zdyB5wQhyfvurX9v3YCaStViChEeBWkVei4L/QyE9nquiwx+yiVQ9/lElzq
U516iqRcJJZLITBMjhDXr8OvDn9jeanqzte7bOfqMv2C30+NalHdw/0Fd+mBGR3/
ZEjUYUVMvxw4GSM4uDlzAFx31WwXw6xCIHjPFJ0szE+Gxq6/z9+ROd2gtiP5/NlX
nbt0R1FEWl+FzzC00YE6QUH4qZvRTr4k+2iNjMZARJ1TjxnTUNOqbG6l4CkBf4WL
8IEbKIllIKbwfoU6U4sSh9NsnZvTc0anPdkR5bCkDtVFnf7iWDqCV60AH8z1kByT
cLjrxJuhvDlXWiaV28GyEoOErRT+APxhM8HZx4bwfWCFtdLgm80Ox1TBHpcTsGS0
bse3gw9c99houiCNnibSVqwXu1Yolq7uM53X2ru3MTDnDm62hSu+cr1AkVYH5num
Ir3ehlEe+fI8k8IFE5MrrAsTZtZWmYrvdqj5Ztqz0iB/34NpoBcQ95yITKdbhQN9
8BZn8H13pgrUnR39u2XqEnGxTYd/tLbLXcZJmpyiM80IGPVbHDgcYE8O5RdXABbe
TT/sEPOT+Fmz0cc+rdrchLO8LkGVl05LWLpMd4AqP+2Xmik3y8yojzslttyUoTgp
9+4HaTbC3Yl8u7v1kTsMQOejx7Ogl/qZeJifbv0O+SBhII3PhurfKRnlYgM0qKKT
lxlIWRj+WgcASADBDcyPwPoTg6SM9DcOG18yRLyQwt7zfbIXXpFmxqEBZ2ur9+tX
zTPegkUTKGyZgJbv+D2OUCtzJi1uCzuJU6cMD8w/USchSCsc5ESXWaThIU8CYMTI
HpgkDNOzUHwWHf+2/lUCVJGrcVF1bGJYI6NI7/R15yo+o7B6u7XVxP4xwdzKgCVR
hM5qaxd5T4TkRlCiJwPUzX5eecgLWgqo133mOt4R8eCS3uuhllMKmEbiMvG8iFJO
eA30J6uaxf5ZSFBJ8CLza3DCS3tBfFULboArIYIl4e7oLttCZPXa4+jtCxLzEg86
ygDrV/0P/fFGHnZw5sww8TUNyfIZsp/zTDQWWuic2deI4OZymZcUWmjeWjgCPpqC
nHQdjJsk2vwJy5pSDyuOKBDFrSCm69cA9dZEeSEYqLWU0wfP8kFAMDYnFjwdG8SS
Dir/w5QH6bk3SWMrx6LHRWGUiXiTJi8pg4rkv7DXa+6Kq8IzXhwmpXclLS53zTSA
gU01HZO5UukALKNCt9VjiQxcv4IDBj+oDZBHJjhJzdmL1K6NyaA32v7nb9v+7qm2
ApsdDQ61hgURavDFj17UYYSWieLxEdK0fhJrAVHBqHpLix6AoaAP8xIcdXD2AGuC
dD1Ks4zhATYvNcLlUau7A+seSljERuqo2cnctBArD9/507A/J+KYFAtFK0JaVUEl
W7WKmHm5PO6imW0ZpMrafoond0Ja0ACHVIaPP/8EYmqmAkJQygGodxCq1eeVfD8H
KUZN6zQlGFgJAJ1HmUWwU+H9c8PMWUoUPNmXXTRAeZ3ki91T7bPI8X8rLbBDTuJK
mWbEuGKeUw2+x29xWTD+Oz1jW/uJW80XrtD/kRwciL64dkIcHVxpNUela2pZL4fE
BnTFguDjA9OwrJ5AaG0EDQ9h4bRwiN50i8KG9XD1ee4QedrPOlEGcd583sV72Kq/
J924h/MoHYDcMhLTcK22MiIMCH/B8AG3UGeowPPt2Jgi5rN4zMsom1Gt9HXovrUp
nj8Z96BQDU4GXYBmhsu+nsgLXd3bbm6BAfxnEjKT81GVQaHHGBVC972SFFscu8qm
3JwyGwCcBQio9ADTSI0cTaUK7VmDkPV6FAg+iFzwRliWlYofVezsmuQQ3s0ikOyV
nInb8u19gYbEB5ngpsbjxRJ7xN9K6fIFHm0nLVzX5P9DQmfkRVZDCZ9ORGgM7uWw
vZELgR2dq1mrl9LIHOkT+lRFVgHqVVuOvR6uH2OPlj+4kIervt+yypLQ31lbJwSA
gHIAU9aZg9sDdSvUTA2EUa4fy1VmFdyveaBXJpVEDCQkgfge9mNhx4y0N5/sZfer
mjzTE0DangK8rCP4Xx5ws08qBxEDczUdOQXmu+Fg57HR7Z1StkeEZC5aZYA3e67R
gFVB5KeSfdKyG6cS8s7Qhxz/olUHsGuv1OelZyKrZXPj68bQTXMzh5xsd73EwAHh
Blau0/5/83GebYB66NwWjd+clOtTex4fKXDw04A2bQicG2PgpZoixHcwOhCD98wn
sZbe9AART39VTaAE/ANkgXXVO0MGviUC1G3Q5dN2GawKiATWl3DDVIKtmitb63ua
CzixS9BKfJ4bk/Jua4YIzB7Xjhnjqu5jskh6h+Er+/Nm1hIhkmp4SECvixp6cGfd
HHaMqAdaytS8rLGtTkLc3QDLxEDDAcWdMITNlKTzN2j+A1WfoH16vDmlvOLL0ILK
2o1PaNplz3PDS/5JUIgMAiiZefnWHBlxFmwnI+ivTBm0KOwbb8Q2ZJnMeP38FEpL
6pG6MMVeq0Bew3Qq0jr9YZ905o4+0KYQ9zO061/ztRyKaCS7lZcYsualdFGVjcpS
we/d0c2G8HBMasmp7Q7r4dVhx/9xEqvmwDepKfvyHfvMhFlvbIHkuVFu/FQlAwvT
rR8MOIi313XFVAFfGfYpihyzQBWjQgVxkl69OxbUMi88Ssgq64kacbzyoBo6D1m+
xj0N+IjZo8nVprzSL+uSmv5j7gEEL5CJgbS/q8ibB782gs3qs86saPqhXcjSlNBb
cn5uQqxvoc5vas0fcOoQmbwntlBNI7iZhJHzc/yHV8/G1QN+tTXzhgN7RClezOlj
KvQsSIeGbXdwyzk1+QXtTrNhmK3qQ9AcxMLoleFhfb08E5dkDyR5cOIUOsUYSXTk
3bYgRhqm0wo4YJKbyYvrb5KZ5Oe/fOqTZriSajWQRm/yMik1ZJRThYglR0UAafgO
qrNxxmOElN4rWIZL9AUavxeN5oCc7gd+By5Pgj9pRsP77rjvc1kHLTH1z3FVCXol
rtYsswgShfMzc28YsUCYAT5X8H5gC4gJgaBaEtZ1g5PSjv+qLTxEVt/vkMq4gjfb
+9ZlifNjUOgxcJnIFaxva3nvih59/tFCW50Zr5pOnX0UEqQO3VWl8r9nKpBqxzsY
pslHSGR7+sqdHO3ADK3eJE9cPsjs5ffnn3BDuflgX2deoM+VX6e7E+bT1eNdBrAY
8lG+u9XiM8+JvlXFhxCYS19I95jxRIJIjBMFXHpi0i2eadtnnnMTDR6Jyb0vNkTK
m2d7cWfYoAuIpUB82Tu45v5GlSoImzLXZuVN+A09tseK4s/uGAu6B5ztB/B+hZpH
mVFeivIW6AP5NGdyrHKN9YyVb7e5YTL9qNYaNHOaMTx1dISCi6ph8bap8hFFUgj9
EL+IjU32AhYSjaPzsTSrvCgqtp3aj8AU9F8DeQSk7uJ27qCpP5NE670wcv+owqwg
CVT8nxbe9D86WQM95Hm/zjZ6bnzd4xepTFP9QNiA1u6J8//cBLExmItsQLtiT6M8
2GuHe00Nwjz3ZFlq+nw42a5/ot2zTBPnKpi9iDeJ+03+O/p/9l5CNVf+jY8vNVeF
TIFFdUPVhXVFruUijlbfi5fP5QmZipC0/KPBdH6AO6VwvUkY+xNGV9EXHX3Odwhq
JCfgy7m7N+vJZ0PwLd27OKRCLxkHZQ0ub5nTut5nyVV6Yf5Jo9WG/n8iFVQc4HwL
J7MRNWtFv3W43m/cG50zhm/M+AnB5RhI9E6jAqu4vtKRQiTGzDS9BQzDBTKl+VH+
N7JMb68EA8bHqzzfB02d3lHS9V/2gk9fxjZx/RFOMY4v6qwkE+r2JLFRoTZpkG04
3PE6yH9W5docv+2dFU2BO6f0IUp/uNC99ni5PbbW3i+OJoCwssZfs9chXpQQQKoF
SxHU10Bh7nXg40XRujd/UDKvEYWlvdj7ZIJ4F8u+2P0d5BuqqvsPOz3Fp4+iQ/GP
urq/Guiy1yZq9+JIbsQ1FrJcRaBpfOo8ycQOt3cA4+1PfyL0+gXEKrm7Fm/GCmTd
vE9S1iqa7yM/v1uaoXWr3/rUHzCyfLyoQhcJV0q5H4jWz8SJ2V7GmrAwMdte2Pv6
07FiFz33sW93yVkTpDsja0MJN0oZNVpGLLy8MCWMXklqK02KaxcDMiWZgc9xn+tY
hK92cPEJZ39ofs/oYaU1Axmwhqk8dkSo7CS7AvAzshE2qhBuk1/UFkoVK8YhxpPr
HsMTGYnkiXatXmPX6KuUt4zjcv+siPEHxMtTIGolNcR6IRP78gerORGDLtIxDtyI
jy8wShZq+BkCC7TmT5ehx4VsmO4ObK0qH1mrWv+otT25JhD6pXJPEU874dPQYun8
ISdP+HaH9cNqpCy0IkL1r0iqF+03opvlQAAE9NdwrWHPBJWvh5C4NC5PBes4TIch
uY4cLwpsWllVC2UWBRwZCv9r1fetZhVRRGYA6zweu9J0nWGCc/HojvI03OxvjFw9
HOO8CPaBUyKD/9olEXQQZzSil//+QvXfE2dSsAdCaTm4whHsYp22ze9yoNl4ffRK
2Cb90ibjiYyIfokhBW1Fx3I/Az/5NYQ9nBxMW0fmbQSSxJXyfZSoVRHNLR4T9MGi
DnnEzpNKQpBdAWG0zpM1IzjCSw+dmFFRSqCAQrIffqsWxKVGpLXtN3IIVT1ZwgVX
wGxEovCvsb+SrgkjvMkkdMXt4UXvvdIQ50PtJ8MzeIlZ8g1xTAezlWN+WzRH4LmW
AagdlGq/12bYpUa4+bkr70xGA9niAt++jwfyuXsjQLvnS0t2AjNmQwVQorZyyqqE
edTx21zGCnRn7OX4sdy5Lu+DsQ2cMV6Jyf/T9YhWXdvr00DuGNRVXAhd7NLFMBe2
JIkVWKgBX0Hdg0MBLPWX9VPKrmtshZQXNRuND78gOkQcr//x2lpNIJCcW/kFTtcT
30gaHYKZkD8moJGV8Em+LjBAGR+JVJyGajXa0EpGRfd6VpGpIDfH/Rsud3cjy6ck
EtdKWrq19Bn12CQxzJO5oiH/tNESlc8culfD0SRYcEp3xfkNU/1m+o3a9WvrbZyR
tUJLqSngN0gD5JJidd7k91N8yv3ul3h9MoZJgpn9CCZ88cx4w5R2hCLDFzMaHUl3
fLVHlc8dblA11uLeIKshGw+XU0cF/jnxMz/huFqRb8wK32I0J31bRp2e3VMWy23E
vKipbhHnGENffh0K10l8GrDO/JiXrhrxtyV7l5b3ayPVKWJCxat4pUsuB09liUu9
iTLxSRGbMRVOnsQiZhI4jWyMQVVl7O//BwspIz17QErmZe9NS04O5dw94lmxBIcl
ctgZLtV5IaYpmoUJWCtefySdGgs3FkbArpmhYLTK04db6r+gwUJqbMWYw39eLBqs
YqAuO2PmvDFDeYyqsTk/kV5izeM1Y00kj2VyGzdUT6lfW9mucOrgh5aUjFNDdZpS
bB8HhMWqTF5G14zA+y/kHTVf79GGErGnKID9qPOtCulhkvX85KJ4Qxis6m0zaep8
AeFJaK+nNgHd1gbTjaWigdJL2gxq4648UT9RC4bj7A7a9xvzluzsPnPVLgy5T6NX
VPbSA3+F/j4Wh8w6o6aY8HFAFGlvOH3TMU+k15He73V8+kF49HTpUhIcY7+BHjiV
RVaSjMT/yP8S3+6Q79nthmjdD6zrkcxGVDvNbMBCi5DlnBN/PVRGSyAu1TAOJPFD
oceZJKjEWgiMBvwqJUgKOeEhp/+7rg3cv/9rjP/e2cgTMeLs2y56yKUotbGhnOjR
kZk3TsIKrsGlVxq0gaupkq1dNM4cAAXEn3J3rBB6F8W8ENX2apIOGPEmN1fd/ZGH
M/jOz3tsXKXBuJATzGKs9ynsYzfaAhvPc8+EFvYCzU53qFW4cv0qZ7u3+O/uSO6y
koUj1v92GtoHV663ccKjli28zl3ZiI9R1auHR/R8xK3nLaal4I5VTc3XnQOGE+jL
1lqn5llKUM3C+11BFxseDn6c/Tm7bi6i8b5isvrWAp/1Crr3aYSBea+DEfozU8zF
Zam27yMFl3ZMgwEHM+2utZ1nW+ddj2H4LiMktAuP11aYYAui5RAw9UkdkT8BbdgR
YNKsbAmhJGmtQI2/uL/SeCrTjhH40ReF5pPG5M5679s89z1KVkUrI5013T9GTUvC
KM6lpe9lwCAx+Gxk+eeviAFYjiimOb9NAFQAi69c+8H5G3UsTjLiqeZgMKrGGGtb
+q3AXRzrkvzfKkl+/2EWr3xZfq8MC+osRoEbTmg1pEXVQKDRF1PRg+W7GuLp76ts
rzPOveq3rZFsW1EpT93qjIx3iJJlNzw1uUcUCzSRN1vdR9+qMg3/bxOlbAT34bzd
vxSAtg6PBXMg+jcMxRRR2Ptwmab0lMjOpb84C3NZtNa3bf8uJN3VwbV+tnVblP6q
Ipm6YrYKrCht6p0D/lb/W+C21n6CNTBfM0vlZNobzlpdIU11f/xQ0j1a56QcYDlO
FE5p61WLjQySr4L8GUp9WZBtu8xw24zmS2YFYPLOmX6XFRxiuK/M+ctHPXpuA4u+
P2lvkMllGHPczFWLtsm4AZ0ZwTuYwj3InMVAhc48R66xwWUC+5btoyvCyRUni4mL
OgDh1e5ixyccXrsb0voSTAgyH4ZmlHFsGd9to2V8dIyNWxVXWG3sDRnyIRmCMe7e
W0LkJc6zFqDXawLiol7D7rOiJNejvfoIij51a0NcG7ofUr0lSoT+uEP2ImsVedel
qU5ToNFLc/BWQ2jKkJ3mZHRwzqh3JehH2vA91c7JP9r16as4MKvZPDY6O5l3/jXT
yVIDaQrhsB2gNbx9akra3UH0uxvGAjLmL+VM+xpLaX+rFyG0RB7pT5SO4VRltkkw
GXEXoJGtC//+nmzkMJBm1dkBOGvHv61f2F6MGlEL0edPyjTFwlmB7kNjJ6MlQ8Ym
+A1oYMnx4hYRBgHuM0zooXAR8RMAebikg2iodzyIYJeo11OnIDpHGsjCU2M3KbaA
bgCJNtAMGdbtovy1hRE1+HBIB3nFbziFgo3XsP78MrBT1pRPqmWdbMcAjMZABpyb
U8tiU8+z4mYkDyvi2JSlgEZ95C8Hi+9hQ9o15fILzpXSb6p0OS4os7RnVU7dYFYr
G/c7GR6yutj5AVnqqfmWB2o8L2to7V3qpE5/oTN3l5hBKWzeVqSCSdbz2sBJm3rO
mgJROnMTNFkYTOKjezlrux3Ak0wvUOwLsvwJUDE5ErxIZwMC/r0B92VQQoK3xMII
QwpdaGhQLuKN4jUKlfR+yxfDqdWxkrUtOqwUT6SsYRYgvKVV3KnebYmoaciPmKV5
yWKquFOP1M8rj8W3NyBrVzQL82VLJeHE+RP82VoRrtGQS3W56QmTwnVq2L0GYj/v
uy7ldAwjmb1ONuc3pLjKGGJ+17SawRQuZU01ySejOmvwY4msdxlR54TeeU+MuECq
AnySfv6r79zKlCdPskDOB3hsbnJjhf+ZFlMai6eDGbsqw5TwiWGSZooX2rrm0Q5R
UMRtnTdwWoKXYOA6G6NYWMJdWRBXoXu5VQqOnC99cm0XjP5VddjPm9UIaZymU5o6
XuAwsVueSRj6s0f0wVK6YzEtMIY75c9OjTUup/ZsLVdgnJVgce/IwQNGWegDbr/n
7bi25wvXp5ik2WaT6LLhpFhH1BH/YX5FLW4KeQ52LTAPwl5ZHf4IP6PuTH/hLRhu
lo23Ho3gK9ITUyB4azN1nVGL//V9Wa2tG7WvX/uwHgRhDfVRcchh/gFDaET0bXZX
/NOHLmEhbiuHcUq+7Hz8WXS/FvxBkvW1s+v5kUGtwfsKaf6aXKwkb/1z2lerz1IH
uGoBlpVYcI4D4Nc3v4ApsfxDO1VjUrBD2984LINsHr+Be1FRhnIzIG3cmGYD9q27
NuItRbmvjXlhJMcAqjp583RyE1x4t+3muCOMqDJr10qnrk+Ujwv+1eeIrsp/5ser
Hkn7Wcf64GJnKW/dLaxwVvyezkGGpLmiZsPVVRzQD41+KsPMYVYK3cyEmzk+E8br
0l8RRTJ64kzVC5bgOo4LrJL12zlTplp5Yki1ogd4kpsbgA0Lm53VWnw66CUhQk00
ny1QF5wxakEGppZ/pgMujDCDnS/ffDdOM815cAM43HjzLqWCHi+kbB6EMDiYronT
0xjZTVpgaLCotuN7LDGtzzIl9rcdwQPCQvqmI1H7usYSYq1lgWYno8IB+d4/kS/p
M29x4ozYrTgCIljxNfI6Hs1Piog859EkL1SSCut/Y9BCScUKZsdEcUIwHXkK33IT
GVIUOBC9GPVBAPPByzeZPo621cxX2Yp6X0AjKH8hd61kowr+RH/2t0KgJby3vDjN
Lis9w4bhEQVtZSd2AbOHauO7YktPyrSYI5ZgqLLeAjfBzpopfnrSb5Rkd9Ufouiv
AOaiLiaaFqANO84IbE8qWcLJ9DzabPltFaKlDkqAWAeuUwFzELO4Sct5QJkWGSyM
zT4+LxN6Zg+PtHgNMeQ/Kat3Umkv10Uca+aAVUN0OkRYiY6uM3HgWFmJcD+OpFr9
ahG7yFnAvCLciOftjFhPq98AeWXfzUcrEWo2y9BsOtxmEgl34+ZwBjqtx0tiNwGt
2Wz0MVMPH+oOEh0Ex9sDPq0ThdOPH/nF0RtmvHsONutwBILeVZ2RY/Ne0yLFq3iN
HEmeWuPAE4YzUeikZUP6WaL9vBCWL7L5Pp3IEIVSZltoWj9qVhbCPZ0WX3uOB4lV
Biahxf683ukPLFlI+sUTrf4Dj6xmbTj6nP1/Uzrvcztq3xtKU1kgESpITPjD7vW1
8jeNB3WUqg7PxCu/YXF6VMfF65MjD7erwqGN9yZmPsTT2UCL7uKFaHUNncai2FnM
cAz2BWCOZYtHtuoNWFdq85RfJHlqavfkWXrBDgD496nBYh2udt1grl8e215c1hyk
ktCof5UQOnjNhRVQ8FQw7IG2pC3YsFdWwMM7vhoOJMRQQTvGec5Ac+8crCORvoQ2
Vk/P51c22dD55hbuHFk3+H58JRZsqG58mZt6ojcEhhNw2dZZK7Yx1dvgNkEgTYsY
/q71jYro8kKaTrV4sX72e4NZFbPQMgrOPnMChitobjTweqRiVdUmFzEBPnvSCVae
6jtNjHjR6gAlcY8VinXbnoQJjWP/toTjh2ccpWrPO5SqBHg/YHD7a865l2yjJCIj
XRgm35Iflwl3Tye03cc7457oV9TC0n1O18REkmFH/V2WQmCdDElaG0LIK8tTjSUk
ZbwLdjAema4xtLxfFBBUXCV2MtsYcFIxPKGZltl87/p1O/kQjrYCST4TYNMMs+0k
Ip2o5td1xDEaF0/2VyV0gsVWX26pGLvmjmRwmpJKhrj7FXisDkkl/hih7CvcyZsB
vFU+mAnTUxIr+79pbnXL78ltVVN0u4HRY1c1/X75xpFgbKrFMe6rMM92yfB4hH7N
EiE8yHgW/xL60wPnzYYftAObna67tZs+Pf2cQ8NpakKkerCMKpX9maP6PI1OxSrq
DRWvlFamNpaAml0i1n1HRrBJey+8imw3uGOAtG4L1ZxAM9QVZ5MLQR+86E28i0LB
ILmRVtRerIWo72wZJSG2Vdu2N1XtV3LCQqmqExNWV0PTtJMBacDOaC+sBIWbPtVs
N2fLvDWRzsrSQERYtP2vFYFfn+4k1EuyOH3GBiGw4ffsllvNwi/PRa6XjqNItgNU
k2wYZMmX7utd5bfhELpaXH6kNlSuq4rwBe0K4Ir5fN0VO1ZtyI3A6qxE01P5M4Ig
fp1bZ/7pUJYI3JB/vxTa17hi0aFJqeYC63/N4IyMb8S85+B4CbbZHrgPAIVOOty0
DHbAh8Z3nOT5SfhS/9w5AUwZK4qNP8wt8/2iqtYHbf79l6gswiEwcfEWeS/B0kbS
oaLD0g9tCrzyWFVUcrlaywXc91XzrI4POWMei6xofR3ifnfFiRcehsEr+paKAbL2
Z/O0JIgmU/XY5rsM1IC18Wlzaa/gZjOKtP02Qh5vlMm8K6QaJ9SFHVSP3hjcPTLX
SRZl+6RvWg4Go3aq2cXQMI1YFBtF+rxiCWi3pqROErPtt4QTadFYmsonmwHfC42v
frAHLCOwMhXHhp4aKsj4wfUuTOkCb7G+9CzKZMBtIbq9LoH6Rhw35c8nLz8hqCZn
SvXARwIsb8D15DStXOB6bAsl7Eoc1/ixh5fG+W4HInyTle11f/vehRF4Hds08B5+
TsPik7lGfgFJdKQ0ls8D9g9+ve1XXNo+POcFqygapYLjuSLq7DERQrtJSkKUyr0n
CSCZ6o0s3l3GCJlTJr1pw8DhgYD3uNgSMbZNYlwtJWIpT37wL7H+ZO7vMlohCqZS
vkZmhxL1GJCRZwNxJCdRtUB9mzg9jk+nPzC3G8w+ZtcuBIhDGw7WDp3gt957sCQv
+//0xUksvd04JEMNW68igUUi6s554vUmq8GfzALjxlA58+oFrLCHta/yst4Kq3Yd
gj7CAwn8ytYtDMOgFUURbWqqHz45y/5vwZOTsIKGySSqbdmlHetXC7T3mwfZHTvr
OmaR7rGy8uLXlnLLA4c6qJIMbx8PIQIr7PwoS75hmhpvfR3daNZmTQaM0EQcwE6I
vTylhc8/F/Llr9PCQKidpO3P/VmBkTyU4b065CHfuiMMdafNyG+TwmTRVH8DMdY9
Qd5nCqkzXfbMhiJT/avLCXKHA/ruF1wOglZFjGGqEpKbTyOvkAGeaxKz4nw9kQIw
Aeo3lmvVr9seV0lkStq1Lm5QjCrdtdEBJ0gJrsWwlE1avTvTreaiJDjG/HHDcwyi
UgBsWDDOxEBNrYKroQBfoV4GOnPEOVy6utOAX7S2Z4kA4frDF9clx5IbzFr09e6M
QdByze7jjeJSvfNte64y7xTqiHg/EY2RjeOG2nf06C4pruerdlcRIpz2pl9GEpHr
fCLFEHLDJVIpsVKS4r8OEDRIGU511X37NobwSkDg2d7NuyuPFs9JRD6l2lXACODw
JPZL2Axm7v8xZP7EoxKTIjbl+gfOcKGDHHwUo1RSQliImApHNZ9qxWD11cD+XToi
bf2vxc+BOVDgMDz0naHniT2TlEUr3y/RgKrWKAwl8TUDWmT1z27YBXy2KeLn/5AA
VX9OYGnn/KzlbnSjsQe7CNLSNtipjKn6izpOE9f0XhNwg+tzsxzy2RoOyFo/XqOO
RMgiRjDlRupQBmxpSX+EcOr/I7pW9QzTCvfgKCASVBbdCpGM0+RqAO1AstsIE10g
1Ym8aHYUjCqoaAER2ZoA9OO6NPYHIWLQt8IbM9AnTKmKPii6/6O4PxP+fOvn+qj7
o9TvwbnDjoU14guT7gV9V74XNT0WCnolshXajBC8Doryh/cY+EHkorzPHPMZZJci
SS29y0Fn+/mlFqMuqv3mppT5ANMCu7iBdxAP1vTAn4GZsyJKj8ovVSU/hNBX4M3E
bnj8601TIwxrV+QWR9+VdAhUizQu8449AzYgsyDeYEOE04L75KwDreHefSOjzfhr
oXthjUCzfF8HhT5c+B1O4eM/32BEgW52AyQ6g0FtB0FZhPXy0gRXoJc5lowOY4QC
+oi7zT2KmemssazUHz7R1rSvrnTzdDdITMPlHzYBDMIAi+gvAFx6Fqon9zKXDjv0
2y7/5Q68upNKMyzTeEHkdwIPqrFFr9HxZZbTljiWmIyQrXdbL4EPipudxaayUymG
PGMkIzzATz2UQTtQOx05WTEAJtGsGaeNv20tpmeyrIn+7b4KtKVmfpHKWClG0eOu
75e9y7DftmbtFwraPMWGWHtEGTlHyioH9+I9wxajxbehjOVvJWnJNZacP7CLHhoR
bfqs2Pd+gCCQNeVzLRQc+6eJloCDPUs1l4LDKInXXp8NF43dTXgrmbVXz9/nadId
+Pohkt1dZvRiYNx2KYDDAhgxtwV9mhX0o0w34/CH6Xb1RPtcaLXHQg/HiiNXDuBZ
Gkd300wg+c/bxGR4IKSf+4dyaBJvXE7FO0YacCJebpktOsgHqj6ekmJLPwyo2bkz
kzFvfrlbyIESEug+Op3zOi3drMxAIw4MHugVHvfwtVm961LQLMD8HmmxUq/Aq5MR
OnBWIIJuwGcfi6qbClvNoWApCfpqVyVjVrxDBpt9zroKWKFFNJk06OffaMxpJTQ2
McbutTwUsYBh5X2/HlNYVXHI7u00G2Ertd1VXcVybxZ6TJ6/l5de4BxQ8oAvYWiM
tfNYFW+KLvsyai4wAbb3tmoU57m88gE3iB1NWpcJaO+gZFB2OdWq3FPtNtFq3vF5
Wx3451V5XxLXok68zG5fht8nJf8qZ/sGvNYII5Wz8LVy+d6SsJoJ9SEtDAf/Lq+R
fxzmKj2Uu/GuAEw6G77LqouNxO+6Oq2dtZTOKQ5OD8RBrRa+ApUxoogMiOt032Kj
qbAad0iCy7PouwTHngXgMLvA84APSOm8D+kbRbijuIB2Enezph4R4TubGnUxKpdO
JxjOY1Tb8jdSEcTXqGl+Q4LeLSmlbeFSGUffT140vuhEBnWPotVa0PSAolQh0+v7
JbWpubhOPzx1RCVEwaJMPP8SuFZ5IX2Va1Whx1gCwDyERIqyJVqyRz3MVNkrA22r
Atudk4TQyDdji5ductZgNlZ6LFKFE+aYzBh3nUBGZ9ShOADNteKev/jojpZW+9A6
pfeT1+weJ/g2CsmBYYpLHdT3kwp5rdKgVBN+tLZN+aCRPLaAVUgQW0gmvqsQTp7O
ljwzuqSF0O7M/+aSwJg6XOrMXm9p/wDMJw4oUxLj/yD5YxHPoPVE3eEx+Fa6hPB8
ESrVaX+boeNKaOWvthh2dmhkI9/43CbENGuP8DSSbDZ/c0fhDy9OKTAosTLZYMIE
UtksRy/mnGJJHR3G2gbkYi6/DKcp5l6oi3K766m0fG2+eI2Z1fwhd5Fw0KtDHq8+
WOC13xKXlOxpZxJVNdJp3B6LzgjQN/F1GdFDj4kyRoup0XgA3dLuv025jPHuudTE
Hw9lMkdkqj39DLVCQcBAiIFr7Xq4bphX/OlejIdd63h8xLmhnmP+liObjh19IM1P
hQz+qoL72PBwRT2GreKbnKNNPceXiAzhABP+c7+GXrb3mTML5utO2FW/uVInF1jW
dTU8LCteoQIOSyBPDnRCsSHNWuIy6RgRO/mpcw6ikVQAJQ+u5VukzWwTrOyY1ITv
xNCXpVLvFwbQFjObGjv/6g3CxBoPfm0hEscjKKoTRzOqcgO8WF39m212O11ZxbR8
0LtWH4dsXGw5FOSVDq1CwlfDlrm4fMzpazEo9hoaq3i9ipzrtDMO23u2zicQn8ZE
Cfe0R8hBXarJ8hnC5puv4Sy6BsThw1qIpmakXXij2S6JmWI3DT52LJBTI9KpTTTh
VbrBdK6SbC7fOAEJeTVN/6ok9kW/9W8OwyrDYvuJeefX7X4oVpUvFo1A746n8zwx
dyeZkUDPcfa52jh1HxB3bpeNFi87qR+rYRoSQQrgLcg1gOCkTaGyRXvekzC7dTVb
NM96QNEabdSB2AHjPMo7Dk6ESuyzOalZ7wmxDmrv9K2eRg1qE17nCci9Zx3XXa28
67+chBi57iZsDmdpR72D9Eyz8O6dv+G8aFCfaqBAx75WlQe4oA3Xnw2nze1FAZvP
XsW1CCHXiCTwESYxwM3WiyZF8c+6AVHCBXh5vDqOQc9qfAGDWUnOhhj0dLRV5wbP
xmBOwEPDUxGLFxriEV2cnes9gPW1umoTUa4qJX3EOnIIs3IQ+Cedslbj1RLExkIV
C9WsUQGwXw88s1XKIePew43LWoIzH59HfLDWwHmgNIpZkqkVi28j9wOiVArhoayt
qI7ZP3d7PEehl1Kzph1ULbb4fC2GYh6YsgYfrCpQ8+Zo/w5Z/UDnJfAzbFYg0amJ
tWaTYHifShO9NQxCCSJWyLQavutorrtWgiz9LfxT94WjUMSWmw+cDd4KFe3H4Rux
kaXcMtdgMt6OMP+wyr2D18Jr7zXE+/M4rXJMJyRQ2i8csoEfyS/WxSlXS1MXiPSt
m1Vaik5uFD6mia0d2y+vsE5NVkTxPLQrsZnmYBYH30QNk3+Bmn+hadpuUBMU29O3
O/jsb543U/mGCrTdvqso4q+a59Bu5yXLGVbobRqHnwse7bUGi3bsdoCWJtXxlG+d
KaZFihU+yhTyP07ue4iNiObbMS0hkBPFebNdD7D4alfXzgGtFebObxFLS1fG/e+h
t4rTF9Mb5eR5IZK0rvPaPvHq3Y00Zv4uBAEONYUeD41ovgBlxuiOyjYdrWHrXuzl
We714LkngkkTHHIgCzMmLFLoTPdCf02oRf17fj+Fv5lWUItQ+VnqypXO1MAbSuDs
HMu+8u3Ssall1u/pIqnMHE7PlM88t95BcdqPSm8m7rNPxRf1tiEKOLb/hX8gzdUi
KDB9bwM1C5KKuCMMKSrQdbSmSl0YdoemvieN2bZV8b9EoNRVIILuY1caIAsJWNuG
gHMUmS0eSNN166Xg0wz9aXF3DOslqBhsAs19269rxby1fufClTGTQwU79iP1ia7T
m/ST5QV6DskN4TWJ3KHY1k3bv5v2pfYlMGjgwbtU2PlK9be5eRuzSDg95cc9OKzx
94nYlDSh+8dlV9HO/mIEXpFCquJWwVCvhubka6aetTIFz0pM8EqQqn7gOngzaFPu
KZjjVUlHh2e5r+LRTKVbJ5JBizos6x+jLCVSnuuO7hnxPx6S6laV33/ghfBFjoYQ
WJShUYw8t9AeaSrQQveqRZ8yRGZq0+d6HlAbTv9x+t8469fvWTusFShR60S6iuZX
Ldf7Oczz0O/+jwFUmqma2olrweBkQeNge2sNq4dsWKIhGkvrm0X3JbMErfIXJ1Jk
CAEdZjIDmqE0xcV+nLviWKlYahV63y/l4Y0GSvpzvnm4PQaQ5o+NjTKg6lGWtnqv
hxbUCOzk8O8rOLmphL9ks017/JK3s2lN8EAD/mjP3ES7rD6ZT0c7flNht9KDMz6y
M99nZtz3+Ry5Of0LXLusQD5t62H613uHHgCWgptfw2zrV+UFOJCOInF262B7ZGf0
PnNj5yY8H6Z58nb7LITWPAgSqz+NVW2bFk+9uNBbxNf8eSVW7Wm1GKQ1ZCByhOqD
AdiZsHcOKeGMeqS/P157ChXFwVWfM6uFX9PJP60SlB6R77WNvnuUUlr37u5jT2wx
JjVJlSDTIaHngVn+wQ4twYzNWAmgE9gUGJSmPd7K7GF3dZfYN/sCuZ3oarG48wxs
wF2m2Msy+ZQUvQ9rAgVwxWrnsIkXAbtwZtmXqupGidjQfBD9q/pXQQdB+tmKBrm7
tphNvPxsTm05E2tGPclQ5iJc8esO75BhDdcmTSL/i1Q884bWHFe1MDk5wDoR31jK
sFEWbDWLeHzq2ojaXTVbmUmZNEER1ceNstcD2qkKg6Mh/NSWOGeQG3nqTa/OXAYu
BUwe4r2OA1kLp3JuG66K4oo030UYcKxHdjTSMBHKBLXbgcaLn5tNdsC6Dna8YvtT
Rrrt8K1iIQG6NMM/Q3FbZiKo9Ve7UPhu2NW60GkM0VhdaWgD1luGO+ksSdtZpBLS
IRaWzxcH+APNp0HTD0a0vQoWK046K9JM0gyJjK+rJj9dKHwR8GF+zU+UgV7DCCdG
u9zf2o0jpHF8wzml23pbc6r70HOUX6qR7EXyph9x/66gpTdn7AJ7H8dI+5aAfqMz
LFeAAyRM5FaAgrMEkJTOPsAuD/cbocEU/jLqdd3gIHIJZPLot9li08+NCnWMteCl
DxT8KCZ35DRp25oyjFrbvLocPjeaSrRm68GycSJQDBJy3PY8i3J7B0Sxw4Iw+A0O
oLGpXnX2hxIpa9bkQBmoEucoMVB376ss7mHzDKg/tX5G/4Wg4A9Q8bLVXTgEJqjs
HMwkdkqhr8+jLbOlA/awQ1WLtpv9ixPemf91mhqk+ldFljnn6WiVbnntFW4nFtn0
VnBttBEM0odtZ9syp3L3ZZ0N84TGom/PMNaC5blckuAM+RiKdA3leDYuvLs9pup3
52kEOxNcAgfSFV2jDxuO+f54hqfhvL3L3yaTbuAqIq8u2GreQUFY+7aDZ+jTpiVV
dKZq3Q3CMfwEURE5rkFPWYdslX81/sXRAAgaK8fOEajXULniJ+LK7U0pVwm1Qu9t
bBgRIJ3QU/VGazf8Em6WdIb/tTTj8QEI45ZJuDZp9zhn9qk2OwwmUEaem/41yYMf
0q799WSR5gmNtANqWKcVq9qVZuZeZwEO/9fBNLUoAkBD0/j0sCvgv/Kn5dRT3RQ9
62kx9uPk6xYfMNFU6Otpv46RS4CREuu+OArTX1SeuDhS1FVZdZya/kJoWzBtKwX7
fOGKJEVh9QB/ojGGvZhzrpg/VjW8IkNhOeJ63socr38AHtIG5jWl566NwtmZWKm8
KzKmNPfJQxtc3r/f650aooxswYXb+rRsDjON1OP/4cCiOq3DdSedLXODvxM8MBzz
DLXMx6s361oNODVK3CFz3Amfd0VQBD0fcbz1M3ej5buAtzrEZOtm+6dh6Aa/wHNU
GvhWDJ1h8yvrnBwWVnR5WzLLnETQK8A7a23y5Q75CQhYXBj3lyrnP7hXI20zE62m
WTHxbZbJ9hA53SIRRWk8fa8bwkKg270FqNe3kMipVn6SiaUrN7xm2LCyIE0Wk9Uo
m1qQvIpDJsA7R1W4pd+Q0AVJR4d/igcM2WehHjmR2MDEnSda1/LR7Pz3IIjdZ7HN
AWmsWUCUVNuMED1E1sXtvKkozVGvXrySd2RVXSO82L+1gzoZ9S69xnWY3SjgZEyk
N1zN7Z+9E72Y49snELwiixeKN/yQtx1V0QuGb2DthVrruqgeFKVuxXZcxeO8XngX
dzxKV9BDZEAUITtX5Kv6Szb6nUt3DNBL9jxDi3NTZfuaHKPgsn+WpCAmLUksT/9o
R68OsNR+SgZSmSXOGNvNaG61zzDiO4wiJmOx7y29ZVPbH1TnOIeebdUMB1R1pm9R
ju5BVuBvdjA4poDpE5qkqmgVGfm+d1SUaftu+IukouJGYrQUB4Mqf4yvao+hsocf
C8JmQOECJd2CkLNZN8DzXNa/gNxfAUJbv0COmKAARmt/tDCJlgCA1wt/h78lT0zw
8ip/Fpa+BDg8XVYc+KYj369lLG1BqNGa4XlLDaJqQtQ6qRbdi/Nb7ccNRG6OSmok
uKGV1oIPNPA3BIDmISW1seaqPpgZ28BVAcSIvcXyG19BvWElJNTNNXM+NR1yw8Gd
7ztbiQEDF2nMfPwW2la1Oh/i7LXtzB+3RzS/ZWOW2IHPdTt+6WtyoKYpW3yJYeHz
xDJh5Oc0KqTg594y3jvwuI2yi0BzDFB5keMTHZdn7u9bz+CUqJmvnDeVvCRPPfQc
hpm+9py/1nq9ykHSGyRKNKktAdOTrl8CKt5tMUICTPYuy66PUCITQFx3v4dUWMz8
anEKz3zDECSYxWblF7mk0mgk8/wZ+6HcFDIz0fJzQnJPUmgNCnM8xhaE6RERNLGd
HMFb+PS+iVU+TPoNyRccUL0vNPOIvtqpi+mz/zen1KNXloqujDmicmEWAmD5Y5hc
A2tt4isqoJHIJIjNUC2xNhBSVI/MbVwqajoqjYFDSPnI+EfeRC04uM6cjmdmyL/Q
fEcNgbyVqFxc2We+NLoc4fefwqvmNPofswPOZMK8lrdS+f3Zzrwm7VjdT7RYK6Bc
XIPgs7I87GZofItFP5GHO/Ke+XGjGDeXASNMH4rUX9VmeblXrARe+oc6tzzQ6/Kl
rALjuHPuiCIZLKfIa9r/xiKq7rUQ01xkPwxKMRtjJElkPTmJAmz4v/iYQt9yLgic
968bSkR4QDVvRPzz4WQDXTip6KfYjT1NaOiEiCDzzq7qkv8Atdd2WgF6GHmWhNcW
+AwW9FstnEv1QGUNcY+FZzNmjISmRTqhm7liEk9D6EDSWESeXXU4rvlXhNa0lJnH
PeZveAHynLdeWuqwbWzr0r3P/MxeZoCjpILR8QA8i4GEVJnUk8zvD7a+w0abPZZ2
VZSixpbkJvnMGtIp1PEZxatLCa3G43QiRJrrPQpdQy9qROIf3i9400dr7VrLVdCE
vviXncFPa5MD2D0UAsFISe+OxCsIvkb81jTU64wB9/FH+Tkkpz58r9vpA5DOcFsq
hKUy4LE8uxJDhUcGglZOZOZmLFYHGYKlgL6radltdVFIgopSqq8EhexKA83k6kX8
MnxMMbgvSuODfUdXcznuHXY9oPeS2xrL3Dr71LKRPHIP5zFEmjXgB+sVltjzo/PW
lRj9py21FpDs+Qdk/SnpnMXCWf+JdOHRzb6ZCCax6tpgsnwa/UNsNOXcbqqaluI+
eHuF0WkP8qRXX9yti0h5Ru6TxAHfpWW1j09WPSicbVa+bSkw+u2OBlmkclBm4okn
RAQ0RZfpsHZTu43t9CvvWpirGJsJ3UMTjS2CPUwyHzDabXP2IezG3I1lawz1K3hG
1SbUubDHnOg9kxF3tNWHELfdTm6U/VE0M0qlBx0ocXFOa0WnfAmS7G4a/MNjbLjM
2hOc6DcDKb9hq7eBPidnN/XRTf4eKqsjk9aNDFRdr7Ko6cXOiQEtT2z8HZGi5HZx
jgJtT6IJIU6u0ABQiHIdKavU16qpkjCsLqTLI3CoWvONd3f/HASQuZmolH/U4tsq
porThfSeRHGqpZh7JS1KuFoGkqETB83f3/FPJFpewv3YMaq78pvpXq/GRJLx5FGv
c9AnMi8FPKhDIero4sjfSvMxtgXTWTkpNuT2V+O0ixyyDQ8aJmAapPZkCVNWsmKf
+4NNxnYNswu2wV9VIevvlyIhPkGk8gdtKQenEXsdWyTeiUZbfTQ6puBc03aAmcBu
GavIsWI8HRyXbkB6yivRmfazflzznKg/thJX2iiV38diUz+snp1pN7QBsC/bWU9A
KQiKR9WpUIWZVZ9w9P2F9JDAz4cjn8tJRQ++sndxBAumpi1gsqvLiRzqSRrl/kpR
xcw/xspA3zO1gBz7sAPGSWGcZx3ZFwlsk4p2zFKIkSxwAK4PkqwJqK0tWX1cCfBh
a3m4RdT+efIJjYjXZowfX3zyFtVJg5lKqPEjQJDj1TOjEnFy5d/0OvH+kNtZGbYY
47xvSsYJg6gOi1+PN4l8HE0F5m6xg/AVCXQZEaKGcjk83UcB7er0Gtd9luPjepBv
Ey8K6tCvatKBYshHi86xKhdJvLUZHlJg3GTq4PbbPT5bmasAK0rKh/gaa/ZcsKcm
OYsd3pIX3qKpOIllmc6ykee0xKFhEPfrCq4Jot9U73BcirhTPegktMXNjBk87Ydh
XXY4ti+CE18zlmh0a0eiVCNQrzu4xyUXIpvXj7jLmwEnO5438k8NKBghG6w5bb7g
GLVa37TDMphIt2flsVuEF7VO2i9a5Ww71I+ju+NnTDOhFpgNFviwi/4Cae35khg3
ktcDaxfyvyO0PycOvis76aZRVDe+orPB6IBd9PUbFo9AXe2X/+iM0QmmHd3agIFG
xTxWW+t5o9Njys11Q8/9187Xv/0K7oUqezyQTF5RqIsC1aKoed2hUlQmlsyNtTc0
/CxUFvRdQORm+zBK8ut8pfkKVIpIH4w5Q7aCby+DQdg51ye9ADb9RUHU9JPelD+5
IZr6fbNWeC1JIsBZ4Yw4RFaTjo4m0NEKaZ03cXIyZuUy3+Sa7pRDJCnXunrdgwmM
9KE9d89zSbsO3xlmr7FWaCLJk5gyBJr4ExM24h4SEOSvpRNRfbfv6lN/+xYyv69X
5O0af8IWFQBy3S/UDkvto6+aZOv/nHJtXbCe7Ft9xn7d8QrQExkvwXdeodDiaOok
p/RY6pA20kS2CyX+qudjr4GqN13TSPeO9+pkuIAwB8dlRtzDHo6FuVPA3hKiKX79
uVXJ64IEios0/knv1Lf3bUEp25ul9kl1RDrtKDe2Nu+DC2ISw6UwLc0ZE2PyEfhd
iWPJq/vHDDoSyr9x9J8QBA2kBGXhLLWmpbGiS2TF9Kn7puipuNuPUlXExBLRopB+
83p4P+jSmh+Vw6b5ELwgAOmdHACxAFEi2hCXnsbfJ5RvRmzBU+BNYJ2Vg4sO9905
troNmXkSLQzvQ98WUJPTPTCkNNunc3/Vdz4NQ40c96ndZqL26expOKziLFFRj7Fm
nVP4sXZHgWYPtpRtJMj9TBN/qnBkJPK3KcQj7Wsq0wTsKLE0ZYd6yWOoaFteyQ91
dy2qi7+yCpRrBAn8EHQYg35nYWwUfA0nKv9FE1QHD3UXS5TJqUAXuTaxM5jETu5D
q9/wqveqQI7nF9+TLMMJAc5cZAqHw5k/CQV/kS6JTR1JO5p6Brwa6yoRe1orGkRH
KeTIG4mCJx98NU0bulliZlJXJh8ErZ+CYF5oYAT90z50RbhlQDT/Elqc55quGBun
iezf02aVMKC1QwohsDdI6lnm5cc0XjcRBX63uXt3dhJZHxgm89LJCLnnMLR+FwGg
4tr4mEZy1k4KJh3EyW4LLnj4OpscCKzpwmV05CU+YxTNCLh1rtGNqFdzrSrstluu
0KpeMf3uZWEoxXFz76ZAMTPN7E4U7a0NyfDZboE5FndX80zsEE1FutgGX5EfyP1s
glpmu6UUZG+AhjTH8Y2tftQZtnV/VzpZpbGFstMDkdAHD4zOjjM7gtUiryMrUfn5
uT3/WudQFAZcsVOYrcIyK/ViHGMsRZn5H0gtSEHpjn+o2SwQbHB632civs9AtmZ0
8U1NwkJWu1sOA+MBHSGNIWNEy/i20pjuFAE53vIl/gtkpy7+jCXPGdWYFFhYIurD
SXevfpkRRk4bYQwKmSp7cWHIajYJsPt7gNI6nYqMooWCXH+DrIaTq6T012OHpKPP
5adCfL0QrFW5TBhr/P+nJeaxZpST4FBI4HOZ9NaqgNQBlMmlfBcCsD8DrAneaJTO
N+X8SSAWwD++xWjrDNaSxD8UqQ2x/ux/f3hb41KWXLbYE8SFlXjHJRotsPTxcYyV
ndhJj5qKFMwAjd/8NmRYkitXPze9ufmt4yNzwyEaJOIRdS5aY0Ey0+SeA369c/eW
RqYr+3v/GHr1tpr5OWGrz517gEPx1SQcLcIAJ/Wrv/yiheiPJuze6PVWsah8suqS
1+ZraAty+9v1Ry5GtZxJS4sOTOTepv4XTrVxIl5pcwb891jYOwyGW3gX3f4OB4Af
WglQu4QwjRsrLJkRaQyyTLyuD/Q446nrOjlQBcTZbC1Q9l4I7KzaZIoOqYjycVq8
eNJ3Fjo3KJQLX65Y4ngomlU4IX4nM1DQg6IGCI3u6f7oUkhKvb7tg9FNur2e4TEI
0CZrInyyAjDno9IaEAkJxNdc7iVGWnOQQDJ6YytCfU6td7MOW3OhXdCpCVupRnbo
Sc2eiCz1gfBcWFImXiM+KvdGgHmM9Rcsl3WjgCs25Oz9FhFxHHCZC0CW8FGBzie5
YutlNXsvTZhCZDRm0Lo7oyGaL9DCoFbNwPzai2vw7lxAqB8PiinK0OztcnPvKqlg
TE4vZS++USMKERztj8XkZimTDoHL8w3uZAlGAP+GpuuglOY6ti1vJ77SUHJ+m+dM
5D1Tip86JTV2qwRwqUMe3QmxdmiOzo6XXVc/UPE6bvrI4g8yD52ipoUKk17bO436
eSS00PH4k0ErWz8fxyIyXZ2zu156j4B5yUXVTKfQLgAlGnAQYL/JUsht1KFRdaOz
QvmXRO1EdJZacaDla1jXcuUzeZyDS1tRH2x7W4ovSlkvLuzZTpaLzgJnXJ6aW9x5
G035uqku0TRveSzQoBpTjTUVIr2lVYlwtVeP3fApnuQbd8eWh+JOHVDgv4Xlvm8r
zAzI9ise27D/KsuMEuU8h31p7gUhfiZdtddQmd2ptcRfbeThut2LLbihG+2tExIt
+o0f4l9e9cAdHdZ9INfB7GfapEWtivEaA0BkqRQOJc4GH5//ZxjnWu6efKFduG0R
nOo8g8ziVeH28mKor6dfPIluvHDStK13JRz9prc9WkKViGFvoJOwlVVTBoUTExyI
Qbs5YzB3g/mHLgsT2BlAeNeoJxOx9H051+dX+NbXe0L9xpn18a9YebtLlop+T2wu
FTjo8OooIUA57wcy/QBOQdybrLeOMMFo+8brVHkblgO+Njx6zMFHTWohvmEMuXcx
JEApqzOgPs65mrKlz4wwK99HSofymAJbvujAUjF4Qg/eMDSQSDwtwr0v1qwQeYji
LhmQ4pPEILKwvqXBAu/p+KxrZBWP6yRZXHgQPHzscVFxWQfyhkeT/Y0P6cnhgTdG
fInas+ngYlcbrz+P0XdHFQhbVr2ed4kMbpIAXpKiOKirip8ByM+1RdQxocfvoBbv
UJ8LUBpIs/NXdYlFf2jkQXcu66KOEKfvJTQkq4el4I+jkZAx3e5n/l2HxuH9M8UR
vUanK1iM/DsKfkjmLQdSf7pwWvhDd+AhSe5XF46rP61o2g8l/6SfFB5zdJ4ssqKJ
vXV+bOJcMcQldstX+XSyYyNJKNGVWkwlEb1zE0QUm3tJdnzEDUeYoUuQOsft+gxt
jAeqqlEhcHnYHOGWbED70Vu/R938NnhT8GL6JMSwAOK/KZcABaQVmRcUmLzwul0f
HUn1fjSpFXXDxyhnBYJ00pdPphLbKGtEQGgAiUj7croo7n0X4eDDd01Ag2vh61N9
PJgpjiN62lMKOXol2VFnPuTOtcR9lVGi6T54x0MYjdPtngw9P3GxGnciEKfatsPB
eI37PEkoKVnOEMqispKALsdcukErnTS6Tzo1P9QhSzCAFYGyytWSc47soeOAJ/YD
PS9PUNrM5BVL+UpVhiYcPpjpFakhfFCiCGkrf+j2RGOiJigdDqcAit1DC5vjE+Sr
qUUa+w2+2ChbhmZr0U2mEeqaGf8zS8HSfibJwMsfJ7kPqX9medcx8rttBzkwF34A
bNfoWTOUc7AwnDOxV3eVq9BVF0W+WTt4HqyZr9r4FDdx4ucVnNT7/hw+qGIAg7ab
1bkxXkmgGTwbPvlQLkSNmD6xw+jP+akJqcklOBM0G9/TnfRg1uLqzsFehcJ9Rpqy
rxJm/JIixNDWUFZ6lodlaGmEaADqVzXaH/nfQPh/RRzRRXXZi2IxOAgnGB/h4LLl
KuqCTlJ2RDmfcbj2jmn0B55IZ48zdgkcy5C91cVWo9aULs48hfW2Qw1X1ZHWgWfa
JAyJP/+Xo9GiWG17V5MIT2b6zhO8o0fQ+XStDZXmAaLtUPDewxkQ0rVpkKK7jcd7
kk5ZW3oRRcTOEYycYHKP93Mr15clCyKhkBhid9h8Xg6amJQCzOWXiBXz1JwBle7t
VOBA0rI9UQW975oROsvBAZ0p4DtDRh1kcWnRcfPVq5w8K2yzOb2kGdcA3r+7rjWX
bLSZi2k30dg0WrxrHsa6R11ypFZX3OMjNss2qvRe6TDY1N9C/mZsAzIW3Tal7qA0
ysUpUeNJmM7zg4q/+KKD/ziHf55UoOteq0Im3PJ3yl8TWtwSYV3G391puzM8kX/5
SLuatXwJkyrr6N9NdSm0HiCNtkDDJgwW8vS5gAHIhAw3ilmmiMvE5eTxqLjkHu/E
0k0BhPXCmsQI0BGXNJ/oUCNIvT6PWo+dm16RqTfcqejcaqPbHhe24Sle5iJUX/yN
vpM1njRk8pHuimPhbVDQMb6vMKfZTYJ6C1HLa5grPxInJNbNHLZhJqMZ8eCIqe0N
4pdHt6TE88ABzUJCj8VP9EfC4mQVGrMlI0AU62MilXggSTs2ZNdk8rJDouUFK1ay
8r8GpVSDbGQddagqkjIEb6GpVJ3LlrPmKu3ft+/x3czaM6XW065BpgeFf6ZohqUZ
50oSV57/3Ko/FOTNQ/gGReQnHLN57obT5jrt6nSauchP3QW+SjtF0n88EuIIRPPu
scTHxL0lnMNiWyDKc8Nf/iG4Tcz6ZN6L5AuDuPrunALaUJQSdUciKiGGjgANuE96
33W610jjXz1YlPfXXog5kym54/4xOL05UlZTTLZr3YXkR9Z3jXImLzVjKSZ3b+Pj
TdsecR5EqQoYpX+WRoqD1FJqYiDo4eeVEEbn1wX0klN+VMWBhMzvbau53uiEHUZd
7lg3BkkSzwIcVBZediheIWn+7vXMg+5/2H8TnHx/tRnbr5hj85mhUGkaVlM4fiX5
fIKoPk3lSodfVBFERn0VHqK0CCFiyoJJWrv2bvuItKPXVHrJzBzaKcBGsz/7a+sC
hdS8FjaPnoY8b8X+/TYTWGVez2vZtQxPXLOvDPLgPAKWgxwd7VC9/QY+MMJvg3wF
5tp0YZdwDj4Kn/AHMhVF09JLFo/wCCQVWNWZyDmgS8SbJq5yksmfjTQyOLfsdNhG
R4TvLqroPhvqY6vQhxuZ2yM7RtfDKt+bBFzvz83450hTuQqOiqEw7nULxAmjKv3H
gcgVRxS5aHj0U7F0KIwivWwQpepaGSGslyGWjdUkvdlPk9BlZ5vkaED39Oivc8QA
REqCqYJ81iCzabkKDCB5glhJ9lo27B9QRcMfSljuiKQmsKOoLXrlOEUyZU14iLZC
fizB9T6g47qSwstpfdz3nS0BRWPUuFYAJoW+DpFdo6HGNmLNZGYTBCqmEwo/aj9l
f4hAL2DW3ngOj67X9eZETe3+aRnnpHkpm695IWdY3o8lIz/UiGqkJXLCkixbT0uH
/Daz04zGcDPpg2e+cppqJwKEnL3/X9qbuc0OauaKTRgcOKdWxwsEVg2kSYTn7BC1
pGkeKTAZ+0Ken5Z1frF9oa9j3mm7RtMjGp/PEqZL67J5hEDJVa/lR4Gd188LLT6R
QDcLdANgPM2EerFQGMn1xkC6yCx9ehd5cuQ2xNsiJzNvkOttFAXAaPfcFwNh4M7m
P7gAz0d0QK4YhIYVVgqo7fNp0Fpq5gmax5JvSAp5Xy05pua8kPZmUcpIRazFDm28
a7rzX9wB3D4/DhX0wx2rfLtm1+ltc85V2uuLivc/284apZdwUhtn2dfljy/WLy3W
CyOqXI2vrzFHIEP2Qd1MeIS0goIa6g8McaDdbgUMzDUEK7ZH8ewqcx1AjrzOq8q/
yyNN+/0deHfHJdwvEkrT+2QMyi/COLBYS6SDTW/KbYHOsd6aqF9oR6PiiPJFC0zV
sfHPLPBPD/VpWbHh980PTVxY0rLHZBfrN/CmFy2jc6fSJ7pJTTa+AaokeHLDT2tT
BffEQwbLGtQ9MF6PuqnPmqV3Y2+un7pWkzqCloPO9q6x57k0dITkxITLXx1rR9vt
0YKjM/A6BXyn/hB1nlgtQhG1hah/nYhXtE+Avd0OjfFvBwy1lSYEyvno2sIZGyC6
+nXJMVTS2bITmcn+YN0LNa0NAJYQg5n5+J7YukUu6HRmHb5coGSJsYkQ3htSi+Xf
xhmBiA3BAfeyG1Im3Oy71cP7oxqgi2f7EWogXhZCIpUGToYOMh82+9ZYJtQqR9Z2
QP75wEgIIjr7uTrT5wq2n+8UCtRjxdYn+GwtIRVky8FFXiC7TXx+UZ37ucyxGz9Y
5UAK+r+L7Nzavmj3E2HDMjZIp5/XCyipeujbF20JMVii9mRaMCNAnPKO4GGMFjew
iH7JPJCs2A4w1n7nlGjTRV5emgFMbVUsX33Su0kZGd3sOEImtvvJU4X1u+qJwqES
ybYRxRDDjRmvWelT8jvMHsdjWJ1c96OSyfdZ3BuAL2DdqAuwh3Ph6320h9OWjDxi
4lcZjAuumOhimeO2ZD9FRAQhnkXJQ/Fh5W7sMFZ3/N+mZBHAzv9vSQbAaC0zhgCz
YPJp/n42GFbe1v2VOsqc1rPeBuxUTrPB2T6T6uJTXPf6eVj3Pq2MqxMZNcdThWRJ
PBOlOWKRt+bGnpOZ9ItjjEgSBRUtC5xWBVU9gVMOzFgJOvdbIonNJ84nr2jQjmbN
Br5ADN3VU0FWGMRMbTPyGIZvv0vx9vtJJFL7zd9KsEUv7w9AdZGP+j+gVsq3NLuh
mkP1/pxkAGE2+Heb5pDU8SVt+cBtp1yuNddOgrQuAsr2+md3IkyeRIWyk2WyK031
nj4ZjtdP8RkcUG8iKJ5/RWrB4D1+v11erO6qJm9cBdNnLl5UoaYEnITw9lWSa71d
hldTOUrkD8cJ5YqzBLxg2qCN2EvGvksjviRqS8dh8SkszvgcZwxj0x4uJyz+4Pzn
2Da5lbkjiwwlgvhxM0NmAr3snXe4Zpk0RDpL3o6OA8krWk6Yr9cYU3zxGUcdoEil
FP8iqiUm+oGNq2DcnBVTKKqIFbm7UGGxfON+A8+IjRjc8r++5Y/UnpLYI2rQhKlw
LFT/4AgHp1VJ02/lwZrlCbtZVnQClKv3Ed9ur7TlPDl5O0RwTZQ7hWJXVeTCttTU
KD/i27lpUwA0dV9aNf7xyb5hKlqE5eXJ/85HL3/TscCvUPsWCfwfrx0HhJBQRHYi
+c2UDFAh52flCzTRn95Ow5Z5e0nqyWNiVDmSNII6W2ne9qBrkygbzzWcYirDfXU/
KKxSuw/v0m8d37zGI+SJwqrAl5w7PQYHny18Zn6IbCW5IkwH4sN6DWbkCT0QYp4T
ygZApVA2w9jt1PqwW8Hy6yqvX23BvrUo7YOWxCGP9Wg4gCwOWk0ceEGal6+he4SP
EjLBhgLQvxgFEO1hQYmmJbrMhM5Lb3fu+gcyuVdrcdFZ1ELhCCMiQ1pz4OwShoTL
sk5G7jucbC91Pn9T+PETIzaUIVeZZuxvSlrdT/oVq1vO9ecEOmmF7a0R8Bme2xEq
ZWO4wOw8kjW7vgEdGJ1VNdfiEUe7h4IKcR2hmyHfj7SwTOANuID9/NDiwjaFEzjo
T3CDzbfC5tWkRAUv9MjAlvrInGOBxB9FqD8OuvssXAxKRLDP8cOJZ+5O/0L4U/hO
U/7vz5u441ctfva22kQ20BujKiDJFRC3HL7wo73WaReZY2wfK+aUHkAmakThdNyP
EiGmjx+9UIfw3WPHds/afbbYfD11sMoHcJCECsKtHqkDOR7CCmPl3Trt9akod0DC
PsE58fjfXzFllCoOiQnRHzazIq0mHa5YKlv5Kgzfvw2cSHeI/0ZD5Acb5ubfuOZ7
IeXsXpR/9uyTE3rvGlX0sVkS1AZ8Kv0+mf0csHxt+O3jK7yfk8VU4PtGjo+N4Uar
uDm7p9/85/bbcv9LudfTbgKPuqYk6rSlxzUlB2ht58DYrr6DrX6D1CUa1EyCIeyM
RVeUdx9wzjcngnhAvR5QWVC3Ve9cFIIOZ8VvgBh9ZR/LeuIy8a2EmYfjsi33G5L+
LsOGzr+qaJoiBFJMLtONGnWkFkD31rCR39dDc+pSCOUd1C/ojGGxjAjgoLjsGJ0y
IXeJ4rhS80K7J1S/iTnqtzIqBONAZJoudg6xjpwOpBQ1X/phCYFntyNAPxhGlRIo
zucMJsBfFxtfI0AnHkOakyvKiFtGqICPKv25F/QpoutV+1M6mfePcBiTxUHEK6rb
2l97QP8jqBTWfKSsuN1LK/SS8sXdRW5UgJydvq8PTXxtlKn7tFD4STn5+m6sO8sJ
qHh4ESHnuAVDa3JV5zd9rJJ16gH5JJ2MMiAVBD7ENuJcAux8lGLhfx9ENKmyEdKI
l/w6buqlHIKp4zHlpSFRlH3fIK0nWboFUqsHSIARyKofswmyZ9vfvjZ1hihl7x4/
GzVFgFxeRbazhzh7ucj+UmECBg7f/qoPuHyvvbr7cSCdWJRt1DU9sBb9GFhaxQIi
mcVnJueeI7YIQ6UXBaP/qgH0W+h9DIVRjgRmVbSoEI7PhldC8WxfNEQtWWSAtOR0
u1Y55OfyJCnzb77vJUp0J1pZvFh/J489cda/IpTMKRvdqbAJ1bcAHoC+sqLERw/A
S8XvX2Iko7G/cg1rdR7YGxd4PnQBFrGPEV3jL5RxB6390/bb6Vqryp2LivDDyR55
vNXJ7B0+y5WlrLul6eN0pFC7cPzHt7uWV20C5tajFiulY5no0EN/0S2jenf0Ams0
3YzNPh3qWobcWkIjEnOmMBll7nde4IRKZH8hcOpIUqjbQTzNlYni8FA1IxlL0rY9
+rGhJ86v++O61gGyyk7S8+7UR4XyDMl3uYdH51TIWYwyrlmPzBG9C0ASCy5sMzCP
jphzpD4Bb5SmCCMY6jmt3OB6BVPn7PByLQWElWi7h/ZhLGa4idgE0Ffen1k7s1zo
xSpz6haXTZz+YUo1iRbXn2SL5Gato9YHCD1Mj0rTTEcDlHj6/Ly2B5H2rcmerOSh
dMcnpIAWdMrO1VZDYUUZ884tEjsowJxHVzqWgZ8kVLTF1snb3qQYukKJfN3CFS0z
HdyltMZ/4IjtAYxE/q4VuuGNXQc3ZRQFQ0FePYCuuAb68vPz+CNWq5Jqhf5SBGJG
FizjIpmrI5jnJ09Xn0sarhIXfwzgV72VlxrQD0a56dUpILDvBQE//K100kJ2ixdQ
m0Zbhg3bimh+8VCmxgpXq7BrTd8edo+A3z7iDLGqIltatnE/6S34MBvg/CzeiyDX
C4IQWeyCWEB8lqk1HQbttHiM1/Izwwe7kCxY+TjL+DFw2KWkf89Zc/WAlN+Sy7tq
NFdBPwlLtuU3BD76Khd0UkOwTdnP8Ybb4tZRZL81Zh/7krNGZ88GEVoOvmKvPCVx
Npu1pz2sRYaLM/Zd5CQw4QaVtUajpXGbeDwm+Mgrs/4RmDNguXDc1X1qJg11mrux
VZj23wz7U/NZLzPgHg0U6Rfx+VTp+0HVh1LoSX5rNEajjMIZi7UY7BCw1BZRrNex
qSvq8t5XmJeIodppytW3JdqHQRRMvxbXE1NDoZ3MlPvuSqoDvzu8ahfxNpIBE+Yc
wn4SL7D4tf+t7tG1GZrCKGlVBGANPDwxWWaCeY4ey1CT+nZ7O3NiGyfkh9+IeHCB
WbTT5dApURcCsEN7ekF7uG64/hGdiv/e8gtu5tySPzeY81LjPuc+NzFgfxQSGThM
pHa7KY0nVZwF6NlIROQZa/Q8GM+XcMBD+27iweo92/FiI2RKrtllYAtpznbAY5Gx
Ni2qh7o4ggXiwxUGG3oPnmQ5veUirG+NvAFJpWVio6JugpRqg0aFck163+HIOt0K
rraJF1AC21F2uAfFocXMd6UOcmQ1F8w/WRY9P8JXLMmN8QY2wuFCPgIhem6kKgjJ
D8LOzqeeQWH+LEj0DQD50jCMUqd98Rdu07MJHtxDvE46ZncyrO1xWcLYVGKfo+Ce
6KiL1HrLoSgJbFc+W4R7prIDc1atAqXxLWd8Zbf6ZESwTYV4GJJuxihTd3OW1MkN
Y5bKrvv3YmTJTO+CRNV/ZOfcgutq5M5wXJcGORVxU8ofDV3PEyYsTgXT4DfWpflU
exIlod5ra80kvr1UJCyKXLW/OSSZPfap22lFT6qNGIzrBFuL4+METCnMrFfNiq8/
S83JtEJgRvVgLfUFWj9uxnl6K+BGzHG8oNLI/YiMyIIE5e15EI2A8DecEGnDY6EE
f6GTKF/2nK3U1yOt+Ma6mMmfkZNTpTig759iqMNRAkxs5K+useQxk54kjunwivne
xD8sHxyJIKAG2jFNnJ0hYJZGXbIzS+b9xWkAHcwm9zsSmt91Q4zEGIz1+Hj9Wnh6
dqhBNs21Zk7Dk59liTX39O7+5rCNoInopBp5waSbnkKm1NqC3rW4Rj4Lf+pB2TwX
cKzl8i9WMbNwHFjH++GJSD3R3raN6BGe6kQg/dHvA1cVkRBTlK4ZlxkwanGvnAna
8uhhm+6ADFpLeiBLbMSYgAaPIznwaft6Yq3JZSTqIg0jZKgBPWlrSPnPftgwhHUv
joQWCAZZwWe0+b0PBu57h09t0Tlh4UnNc0LmTwUX0lOhJGzWIqvStfiS/QNRklvi
hBss0OzSnoYZSWbxLsTp1V935UpqtjasQMSFuI3/JQ34TFJt865lK2ZQPdtB6M55
IZz/q6BlHQAewmwV6lP2emWTyHrRuIOjcXiQ9E7JMfLWVpq08Uhbp0L62GNSdRc1
YYk/c5ByPctl8s7yUDwYRCs1qrpgxtcigWd//XYdPpu3k0lshh0gJpuMs/fRoTau
NLH3b1EIBh72X1zVYM1tK5qFH/c7W6t9v9Kg2tTq2jq2U8h4Gio8ZiGWZSDlYvp0
EeHGWkOJSQf/M0/RqtQsj9573MuiEeDNnBr0W1bZS1kLPnUXcQFYmK6mo2/rv/dR
Eib6170vvFECo33FYGIsVI/nyHQEaU58hpIXhLQ/UeaKkLWuqJbGj0j/g9TvZuJg
609Q2i7Et4I1tigoqF3CGbGDI1Rnc4gMeWgM/SBnEtJMbcl7bzRNzyeS9eP8Knkn
iyLnCgvz5lTD+NxM42EI3Jn23Kze8CC5ucbE0gGtIdwBOStRVM+JESrYjEQk7grg
iy8ncYCFVgUDklYY6cr53SRPM+aCOxTTfReMRK6NC7zqrXmniuGw1iZyXFCI36GI
CO1stUkeLDJJhWFUfmugkTIheb+nougKp0qxTmxOUYEkEq2W5sTqnRMcMrlZKj3S
66TM4dmP0WQfsGKk3DVGlVhXeqYitWB+pt1zx3SgTOV+ZAaOhTI/ST+PpLI1imRT
1E/zoKsFhPvf31VUDxqrqNxqDEi/cVt6M1gMpv50m4HrYX2LNR6xN9nrLEVCw7H7
M+tb7OCTfU28usdP+j05BsgAIFZdExNIXAjcvj9F7QhhLfgPcTGJ+Qi0m3AnLNey
iaKNSyX4Dzflk2F13hlM8towaXdoL+7f0ZZkDZsgeSOtdlmLV8e7BLIyhNOSBQkS
XilZTzt73Yah+bwKabu8Q+m5qAj7iprrAlIP3P9+SKpJZAAs9ZLzqRwg4LiOVP9y
reAs5TfWN8UfMANxOj6G42o6oKM50MziOVzuiiWgm7GD4oo71X43YRoXJV5M1IVo
PBJKlNQcetMnaTiRDq3yb/Lb9jjfpxBAkNAgEjk8zggLRLK3NBBbkM9HSPwgsO8+
+7M8PvO9xINY4Yg4jc2TpqVwZUdVRCt6yOdDyg5TUkNqnZkQ4yCucSAniQj5LclH
UXrQs2iCEgkn0PFgH2UWkvNxbflI+7gzXJ55KD/B4VjXqSbWJ5Y8c/up1sC0075y
7R2XNatuLh7hgLn4IjyfCVyETScxTLlGg8d/cp7OF/xIElnBiHdWkQFK0cUsbFeo
r9H7pxoFA3xjUO3JC+Gw7H6++Z7AB6n+vbnRgIGLtg44ZHkBJgDAG1gkMtKBTcc8
PbT+h93yTQy/grOK0vmGG0ha1YzSDE44mv6nBGMasGmVOSanSdLT3rEwfGAoBTwH
OH/40b5iWo/EYxpmmDMRDKhb9C3SvtCoT8Rk/Fhbq5XdJdbFGXApXGkVhVQRZMQ6
gvgnYIY0IU8ICBsCjJn6TjERuva36gZs49UQzhDwLxiaFxTmDOr40v93gHov3j5w
4V67yP03pgHuzMVXPMdsQ0qH/EuXZLfexKl3EoXciG/BoLBrSVTBPfsfcCt+yeo8
iI4oTF+VIhJM4pX2if5+7PzqA6W4fWQVyOXtF9AvKisJZOzsW/FD8oj2BASINaCJ
VfLKj7WS5c0MWTSfLRT5ra+d1zWiwyGn6IE4qeljLACJti/qff8FjflVOOyJP33s
hjkvOSYUVt/puqIMMIQ9gSeqItuR5W1ZQKHgH5WMPue79V/fzuORkH8BTMYlAKJA
Hd92uNm3J0WgdVmlruz6H9GHfnwJTUW/0VRFl7NHGjlnvGqSDuLGYQUlaMcnTX4h
1KG1/c/0vvWStTCrGRhs3u+crBfU9Z2GsbWcYvcKdHJOHbCJGNnihh2Ae0k6stTg
plN/4uTOhnINy4/FgIm/ly2XXzn5n93heTmMwCYbcoegueIjopIm06QvgmGjCM5w
QjE1NDs9ZZ5YVmaaMcwID2F8+CoIHEBQv4gkilWYvbOTxsZuL02Lw/Nd9/IVKOg5
ayPmYzKxfGSI7wdmBybR5PsA5lvAfnOW/WNb7lsfekwXgH5I7XOGh93KIRCzNkRQ
XCC4rfoBP8qZ8rTJ5ryI3PyCJI0UMwflMUVgXgXOZduzMvfCcBUO7XaEEQvf2oiK
Ia1Hkf4orv1Ona+ByAMiWeEcapv7Rvp/2O7z4BFoCj3GpxVaa5/8Wu1aHoXKsgV5
5GdzvekYxvbxsOBqVyEO8blKWgiY/VEcxKSn/6FOAtNA7JU8M0IoOxCTIT23gfpa
SboBgeccykfbSR9jx3u6BLZ2PgoV1Xu2M+ZDLFNo6RrciOfw9yCv5rlEdJ4P+Bgd
qzTqpMEaRqwgKKY9/+3FCHsV6fKxqP3GLCejShZdbA15kB1ISWZrRkuecEoyvkTl
WgtzMxkX6C98Z649PksC9G9gAwWKbvovHaxRtzgYQY5gypaeFs4qKZdkPL36zLxA
Q2GYbGSYiPZdBEudg2gA/RmAuKY88rTKZt3kOS1EMIrHa1ZiQC2cWTM3LCbar7SZ
QaG7TNkPg9W+VoivwGl0HipaDmhcmsCSqu1C+ERlGU9jQqHNYXNbKlyrLPbfcsR9
7TWi+tUMamZLk/GZ4LugmY0/bSJMSZCSjXWJO6wzoOqoId2QQPnybUoBn0R3Le7h
nE9Udf2sI6qcATZj28i4yudzSr7rqa0/dmpARZs5NyDd60iUKQLZ3j52n6rBFeTn
RCfBGlYkDce2Zu2IoRguku/86bA7X4FEdZ3FERucc4yj/EixNKUHLSlqMCXYtona
jZ+CtEAjDKpRqPHTkXngb5rah52+smc+71JTxp2fwnxr1iT89I0AwjLiTEMUAgbI
wrgyWpb/qtnMqMVrWePEoOSooBiv9CqCxo+GoxikvXgnJ+hRbf3FxFdB6X7nuGLf
2FOgZZpGgaDw/tqvAm3cildoS4no0/u84iFaALqdd/pqrMazgXOQmns9Fiv3Hmzi
BR46qfmGSLO3GnwLnBn8mYElUt7nS/SH9AoBwJZBVfh4kltSVmRyq6flZYHgl0J6
6ZpTvayBADZhyiFGVkKEBP0pWDBZfuxw8wJbc/ZrawoORQpVIsjNlQmd+f/YLZh0
s+Vv2/aGR6LRLmeOJyEfvP7g6qfikqzGB4zeo1u20HYcCgiZc+sSJn+BYwpOhwig
FddG7sQ1GqsxCj2de7vtsgGmWeZvWGopGaW9CAWwoZjR/9kCXhJMDL+3AMO3tytB
f3bekSymecx4W8uTEcuW9NlqP74jLtwQawKuls48l+KBIs6FTbLI7/JW1liqC/cl
NfSa0qZIe8cYGul5qZBEHvSwA4bPqM+JL/Xuy9n3tSEal2PLuUYZHKpXWvXKpzXN
L//esHhsPfZ2TW+pLqIwOeiGTYo4/x0vvpw0q8pw83imRhEWTEPM88ufEh1pcP82
MKTQQN9c9jRRo9JGhHytbhg/GPtDeEFu4rkYXEY7fklAN5NdZkoRu3+EelxdoqP4
8akMiAjA84bdzqRq69FbhdQd3+prie4jl54vWKx+PGd4qDPfQwfOLqAGoNV5FY8s
TnEtaR+bYqUn5Jx88wrvI0sN3pHgS5fta/ANj6hYqdUIFFiUoE4VV1Ly/rdMfJIE
1bjCtL5gLRgRpGGVFPvPwdj88DiZ/5SCwkHTZX14D46Y/JID5MRPEVFfCc+bHXyT
WJQ/QYWubD1aIj5Pq2h1CrAPybRQqD8o8wvz2W6qvonc3ZF7nYOJv+lnZc5jyPZS
QNMMbp3hcuGVwu5DpL20e3gJDHHGjhlHjjmSkX18LKhEqWTdh5LUS8d6dpgZUUpU
UTmYrXXmUcgv0a44SYASlgAmVNo6kdcdFAcJQjRiEW0rBY0W9BZf+FIiu5HAI08v
GOVRoyxuqlx27Y0nFyatyj1nrrJ1kkGDn8K7X1+yopCPXbttDZffpfY0Ulsc9Dxr
gjRjTCo3eFBRSlKP+ZQh5RIsS5bHBE55sYguSsIQdaP70YvuzTkTr5i3DH19ICSy
GEfsDN0BrUZ6GQv4Yq48L2e7K4AlPzy4u8aXykBgiQ4ou8p2k5fh/jeDdAH5ORdE
lhhTsGFICMwWOdAY/D+9GIv1RYtj+fug7ejQReB4PWqQYKyqcQOI2aCLVlson6DN
wVIk0xBmp1pekOBp3E5uIvE+SsZOJIPaJOi5ikhv8LqA9OcAu2gn9HQElwENkBiJ
lPisjDsL6w5Um39hMSNf7kShBhz/Uj3U3cBqI7dc2fUhKqdTwk9wGwyL1v3GNsOP
rqIeswawRWnYVn3rKhEbllrj91SpUEPdBbsc/O4nINy2g9bqBl9/CslwXRhI+Vn4
hLuD2LbYDRZ9yFo5i+MPSbE3hYES29cG/R6up7JuOKTGjPV148xf3FInu+cAYSYJ
68PPihAWxGR8vSbVAKYgScTQDEjQO5j0Bb3uzHsdGd4XkL5XLZUeoYTYK+DSuSDa
6/AQgPQylefV37t7KKrmEv8DDRY0uavwlkgawhhou1pCKxNw1CGeLhPp4sxpr30G
Tse1RQbgR7NcztVwMLRlZBqsnJb214kFh9yNIjQr9QQTxVyULp8svABMgGnpjJ3C
Zi+7Qw1MpQiGDSUXfcOIFRBqjpHTO7XhXhdf/V+Jy1VAGpTpZdGepZxYqaABe4b5
xwMK67pugRwoK3rdf9vRZPbWh0ADrzBYk4M3gulL/cGVE0CVcLeASCvgZCnXEvOm
52jWNdJZS1S5rfD9A6CR8lWnVAUrljZCdwyjRxG8fMjJKiRZSjgpWmC6HIpvAhoI
Jts1iyvqU6Viuf4SkWBfMuqtypCTkBqk/wGUxigfbF31+51Wq+yXRyBsSmD4M/df
j/EDmnWJvQolL+K7tEbvGb7sRXijV9mM3Ep9k4yoP6oXJ2psoKWO2WfIaCnVnW2N
MdKUUC3rOfCcOYqHfj9yK3MAMC0d5j7j0y4cZk547u4PnD7SYv7xqDlxtgmsAkBg
Fj2Y3/gdvHAUDjupCZoK9Ia4Xux8djnXUJCVUNG178ytj2xmMfHzGsr5YJUkJHE6
CYgPYOQDPe4P0OX3UmzmlqseRWAMJIf+dRfDBry48EAH8LJhgu5hitZL+kJdX8QZ
rxuXSMqt6xeqnWa6Dbnn0xlbHD7kDEnSnDLTEuK3asAFy9R0FWmN7FvMoiptN79H
EgG/MLiPUdk0ienhW/K7w4S2nu6fJLcPqB9LAt7vRI7+Cp+ri/57vNkwMxAOuAw9
KTiz+i+WfMRKGi3qg7kFGf6hdssYGT49tmuJgegO5q7loA+VQ1k56bbaiwTf84Ya
Iuvfczd2OzMyAeKGPmajP1FRlCYZqtP3PQ1ORPYMNYcyy7TtMWepYmu429AzxgUt
GJ47hkMznI7cwStqLzAvVQW1iT2jouMFbF4d+ax1KP8JrcOxLN6q+4O7/sqOD5Ob
EpCv1/JiVViqd1jSpFNDcI68XZZNVzDJgl36YTwYwse8/shGgugpxjKpXP56AY+h
oCv9+7PTZ8pV8zULRvG3QOkZyGp6eJ+2w3OH59cF7Slz5BDbw/5RzG0YuRnRCizr
Ed5tOjG9v+n3QfL/bXA08vDIt9B68stVdiYnyy8hU/Bia+fldYw7JaMR237pM9TU
ujJlDfl8QnAkPc8TtLPyCEGfdjK/+fjLYqhdvXRsD8+qr4RB+AghhSPREYRTodL0
AaDLcgv/u/TwjZSgBPF3lktOTEU9wH+Uc7WhVaw3d0iHohnXunA9w4PCfgtOpWeW
6dmrBGX5yeosHKt6cwUaKCP2U5MRX6dz/oJKUWE7ERS9X5MptAdSinjtbSJ/p3rr
MPYxnFOiIso1JDgOkttTpC/XljtYePGK6I2XcYuYn5JSsxA0F/X2i+IBf56Dt0Z2
fsH6/INHKNaMOzlU67osHPm2tdh3Ez0sin6AJGGMu82uHzOTD4NVb9Q9YzzMTsTy
6gzp1yglg2T18+Baw1ySjBOpklFIrE+3n2SZ7P2SITN4YONZS8uYgNcX4ARowG2A
9jKlckBJM4v5c1Q8tkc9SLL9QSXF0c86X+AO/6d4tWQWhWPbTeameKYPWmIWjxTk
RMdC4N2b15fXJFhrPuTjODT4dj0bWDl6d4nUspfN7SVLy5lrwSdG2tLgXLhi81Ye
SZRrEPeB5bfrGQyhuhSvInFFt14j/Ljzc8MC3jZjoTuY1vMzfOY4T6j961azSY+A
mSAoUIB1G/wWaK+Ec3R6PkZ9JSbr9B55xo+PHz0W+mjKFJbZxGKZ+daEVexJzTyv
0nLRY+OjTb+1GL+lBCaRMnVexHt9KLSOXfldOs6rHWuZrJl8zSyM+eCrJgPpNav/
Ry5h+AtPdECpy3eumoP+4MB9+j+MTS46IHww+V5z1yz9JOPXxi0a8ToycybZyuuW
G0G02IppRNhL+qGsjfxkKM89KNC0Fe1zdze+xYgc9m62ESbQs1epR4Px3wpufZAR
c5WKTV5yy1w6Hl5avIbHFHUjgT9M5m4eApnaeFxzT20KvvqYIaXTr8UQDkd0EbIq
fNJgtuPe/CfVet1pD3BRPKbVuSrVGdoINq1MqKVdmcp89Kdahk/HefSh5ADyQ0jM
Tl/bUZyouHC3mEuBnzgA1hXur3pZZ8BafHfEnHnpNy3wrRAl6oVSiK7G1e+Kjbpg
JrkNgXX2iFZydwtvtQhGlgjgciHAi66pSNpszJ4TDRqZDwYYurQOXynNeZfwkuU3
5kx14w2FBTGVz058IB4L3Sr0SWVi9vikzbI6kqVnJu67iMk1YQFkDGe5Sj+WuqBP
E1fAqnpPn2JXlnH+VnMNagxkfp8+y+6u0M967wlVadqwav7SMYzrj5uRO0jggywR
lP+EoAbTIKbxP3yv29AKkE1CUJmiwcybov04z3zTuzY5xe+nZlEFMjshxtjycfOi
A9Agdk2QBGgC4OoH4hU0wNWdGRf0N10sSKQm1LxjeZeEDD8Vk7ManLgtEZgc8J/Y
F2b3jr15pn462j8gcisNn5SMr20tEjT3PgBGiCJukeLZPGv4lA4eaJNm6KGxehWV
+lNdIs4OsMaeOkg19g/b10IrrV0Phbd+M4LckoWoMqfmZ2D093KfBxWiXHTAOF/g
cC8WBv6GHjJ5pbav6/ND/AIArMafj6f4/CDaCL8JStlimXf5/7wY8YwNSwccgic7
myOfBoSLsJjErmsSpkdte2k5ghv8+eELMN/od8FA4IHv+Gz4R2OBljRqcnRHdlw7
0EWv6FL8LKmpb2jHoaNR+UofgnWWHcM5fN4kHwgv90m6ZZXGLtwbmkDuBZ0bdtuH
vVKbuB4N4k8V1TaJanB2Q43LiTO7ygK2mWD5gU1WybYc8EiDpHic7meJ3qkNl6Yf
OaNdE0I4laCEvCTyhpMZcGlsuwP4EPjEKO+47j/xRQyJtND85RvHXC7QXIMZ4ksb
E3gndMH4yflMl6X3P0F6+1PW1/nQ/LwRGxOzz+HL3jbZyBrTrFWwYExEP440+Gyn
RskEKeK6VaE2NiVgwFBAzfWAWpPY2PW0G5tUWv2r2GVH/mzkBeo3BzbfEoSOJX3V
Dtw/q5kFxdvGFXiiJsuERUqfU3KqXdjVuL0XDGBMbu/i0MZS79/5y0qb5P7Qhazv
hBOb33o5wHcgAusvvWZEexEjK5nyCND+VMK2fEs0PSyk6k+dUm8SMaDbz7r6QWyf
koiMmO7dFd7YTNgYu1bbNnuXrSjOoboeqBIDypr4uDpbD1ENzXa7JSp9iKQittLD
KeuFU+i8yb8SdhR/5MXX4bb6t0mzTccNdZOetBQccEd8ezoxAs58J7CJCR42Zm2w
F1R1KdLIi+an0g7mZo3UwdWZ4Nb920CahD4VjKVXtuMdnUSCP5CGVlcsiDzK7u2h
u7izGCXTHKgGLvBb73N60A4Sbwiag9MGHemjWTiPE61Ugq0/Ek+6BURHI/je52D/
EsykcwHpgGzfadHchPMbJ4ReeWvVMNIFI4D3HCUzCLqpWHPuO7Kz9Q0iTVZwsWWS
rVvr+WtMwuErSQ943Vk7/dgPAqdcNf6byl0WKRl/6YXFDuPzjxTt1xFIy8BZJa/q
fqPvepW/EscHIFxpDHMxAF1/jSEf7MMUuw1fj8AX/TBZJpKgbpQwDZy2AR2Qwssu
Bb1qEAa3dt1sZ3fashxK8Ljm3z9BOM3qAxK7Ix9ekjP223X6/AVnKt4iJowZbmUP
C4zl8nCt0YJbMEc1l5QejsUXLMBXrJofND2BO9SujNhWARMlz7dZNnAYNf22OfW8
W5ekrb3xqggCEg4dYR+q6X6ChK6csiWqdGBqXKoAwjTpNFIkF6vK3kD6gnsbBBMQ
FU2b0TQ8PoXJoNLR+EcHjcAZrsQY1PoewC0AWy+Y6OhbIkWXVqKrYTOPEbsk9VTF
eU//tWx57MNKTn2U5qidbXmwxdqHeynCIBb0VOvMjSZAWhfSoabF7C+NFtDechrw
eecjhbBV6bFsIFlsHvywK2nfoRkvzKE1dIlZUXmCZV8fh5MMXEEcKfLjgKZopZWM
D0CstTO7qI38iQ9ZS1tQ1r5/AIcaWxXrnft63vg5BiQ9F0OnCxL1i0DsKc8qQlQd
Vieg5SBMbtzMoBm4gawMW5d9OTgwfQJQ1rLPt2DFSktzT31SbBd9D6Qdediyk9RD
U6EkXUomvogdI2su87Y2pSubyeycJCYPgOfOSYc7OdaS6pkPjhe1RMkb+0hEjuaG
lFe9CACSeIcPR9/2uSq59MsWOu+Vp5xJdFdbKzRnsBajh3k93EiHu/dO37tZKhST
WmoT5bCiARTkmdzDVoRh1ZCPIEeLYeJMIlogUMx1IjaSfxefPIChOYvrqxyPLc1k
ZFYkiJt9Sq3lH+FXJMLHayK2/fmB2cx5XY9gB1m9Sw4+e3v3/SZQbzdTEUEX2OK5
0Tok1LlXJId4zqWcoyh5cm+m46r7gWIpHRsXBLppe9Le8KF9Uj3Sy0jMbF8HYWWE
zjJ8FbOZK/6A572L873djj/NMLKcFX5HPed/LZX44QalABfgnezbzXCNZhOw+q0E
jTrhYjW5GbiG5Og0owvUIUwrGi5jTb+CMewS/NYulHEL2hDDBO5isof3UJOv3GrG
zu/Xp8uppVWVQY0E6LFCHy42rYoPRO/D3oLMKzj0K6q8VGrgkcyYV+GIpjCoGoCb
KO8oTzzX/WVbeT0O+AdZBeOX46EGdOeMZMe1u/KisETpiHoMjlKunIscQh06gr/I
Zhy4/D6ck87EKRDj01BoQB9s430hMR3gY0NUxVjvWcYbWNm0qK4ALA1H4B01V64t
nw8b24Q33/rwGKF7BVHgKmkG55I3fH16Ep0Az9SKYaylra6oj8QzgXCZtUqmg4nX
nGwOVuYiE99Q5kj3BYXHbQGz+jbFuD9mB8zltlJ8HJoPqkgSZOtmOAIsnH6RZlBW
Mq5UsFRxmtx0YyP7vrjAP+A7zb+703Vgcpx++xWjmUHTbI9Kh+AL8FSlywRFpLxU
BJkMupvxKrnW1kApCXgqgiJzMfE/KPZlDa1gmtMO9emJkM3xx8JEARxa3/gDqifq
nnggUQsQ/YOPhOyquCq1ih4DdFMWIVW5xd7U/r/+DfCAFZvFvMJFqE6slU27JCQQ
r8cBCojoT8AD+knnbIP5hmcv5RwShlUwM3RcVLjuvmn4Mc9I2qcwCvZuiLSOTl9G
q0Mw1Z/vBQpRn5lpUOsoxJO2o8pU2N/k7vAtnFvAum+9xL/D2A/MiR2dbEcZECih
o/1Z1yz3waCtdGJJqwJ4vY+XzI5x+0ksZkeURbAJfqMYkMD+bg0J+jJ7wI8A3fzg
9Dy17HC/xDONpos4iydYoQ0yl/ccPK4THbLVOJykGkplsA/jC0ThIMN+yR+Q6NVe
ysZUCqF5/Ht84RRg6fMRlirkDENWolKcmZshlOFnzO+dXMxI6QjHxiJRmhUt0OvE
T38bDl4TYru66m+w54s7bpQfAa/tyZDU8/AbUDiMcyMa0i7njWlTsjmnNnSW2p6p
W8/Mojczh4QyDDIScAjpSkXR+bUdIEy/nRHYY71Yk2d/Uwq3qXIneRWZcIONrxR/
NzvOHJx3wi6U0hPaL9idS6xu24E/2S04UOqFGEvn1t1+q07V1A8xURvqtRFTR4pe
ZuUFa/VG6prfN9vnu61dFsBNpjF9/OPl+7cScS2HfoABL8SIQhIyqnOe2Ek9stvE
7NJdSJXuBNVjPHftT7verA7jjVCEVIryfoTbNM0j32Wdm8SCBSbhKEjUjW/rLrR9
uCcsNECGo4vKL6RNh0dRa3j0lAkiCibhuuZNwXG92BBbKhjIQypsxK/6/ow0t1ZI
rQ75yHgxEnE0JatuiUdsqdwdLD+BHSQhD7+mozdK9U8qokFbcsGs4ATHKf/PEB9e
SO/4Qx02uJ8hgEVFn243p303uFeB6oKkql1LnRlrE72/sqZkYdQeiouL5sjsNvnk
daQ4bTLkTsKaR+kGbtggOeMh9NRRG5bs32J5yAZHFD0kbQUgCLi9oOrtgTXmQdBG
T+X9LjOyfJvZR+GOPeXn48AwNCAogxEdE6qT04MiBYWDbZErrax5DumEgahMFLIm
GNhhI8IyfKk0N1zxa+KJ74Bsq9ivOpwWh68UKwvqoNfCuhRaqVECGiEs71/hIWQb
CqO2t1Jrsng3vsZpynOsbpyCqnL/YUVOouG1bkW5dyzRKXsPUEOZoyUpp6Bh5Ayw
XsbkKXZlXQruMEXFIxHQlpt32aWMSoG7YMBWRCq7r/EXnJPXXyJWy8/f/7Raq9TF
gS5kjCsW9hbekKVCfEtotdXPGGe1wM/qID9eD4aC0pYPYSsYKtXEkI6Jp9ppj4ll
Y1n16m/ni8WliAtVlLK6erTI9Of+I45y5QxyHGXRez9CU6bXhz8OVB0Gi+6j5BSt
tnl2lDjtnfQRnIKJ21rKVhTmX5kyZX5Df/JPyo+LufQZSta5q/RJrNXR/qAq1dT/
oA71VwoUMfcHCQlWm5SA/50iDqqro+IPRQ30Jrw2kuPvv8H/1lhNEL+MSts+72a1
f1kjVIcrCy6DlTcMCtecc7ydG7dd0B5t477AVDKHyHKm0w5wrveooMuQDOrki66f
pNWPPfbvi1BcNRNk38K02bHZUoqn5kCw/1hgYviBSKO7igubl0GFliPzIZuwWRMe
XF9gPrLlHJp6X//Ioe9fa/sEZDG2bHJQUrRGuPgUXrm72Lh7EotL7YrB3V36pxrm
PmG+lQRtUZ0kAVnOu0vp4DtkUu8oGkCNa1CAm2pYBuNaTI/2tz1PbzjZJ0SV2fXh
RWG2Rnc39bGQ8LrEKrYL5fIA6Bfox9kPRTXih9I9a/l/LHeOMtdYNm2OfQ1epS/B
8DN5gI5yRMh0WqNRd9PXIsWewMaNAYnpqh+acmAPRwtnr+8BEbxYxAMofJAT5SQ6
VZbD/hssvL/Bkevm5anGuoEl7Q5JgbNQpYSdkktJvF88M4g/BvGAunhrjD5cotAm
OOdQU3LB4RG19hXNN8UvtQqnC+QeO3ZCP8JuSxgUtpvJe/aA+oXdejLHR9PY3CqU
Ea4O76CjeJ2/TemNtuTw1b7FGRKzd60rXdgRZrS5hNG8A7jZCymIc5R7sdjyx2o2
qIh/KdKQN+xYUpVf80jjeiSgGIwzXTqTlcq9Yz75ZNlMuXfupSuw3kjVm+rTr9BL
j998uyqFfMTiy6fOo5IJUNAll8pU0/AH8Kyi/It/02ewMoR3mytx37DMaupFSysi
tMVnn/uXuWDDHZzC/75CthE8XL8IyYTlzPh91WybwRJ5QxnMjTpenhSu9ZBcsE2S
CbzSNnR99F/eZpnzLASIOcNFa/Fzc+SDA1c6wUbWEhgdDVhscgu+9BxVA8Xq9UXO
/qPpKSWxLlLSGjz6LOcD0cvimA/5NiaBliHU6ivHoAgCBuy3/jlvD466J/o+v9hx
0zGKpi6Wn3OZj4hfheB+OgL6vqBjnA1ahqNAKZ/E7enP9fgoff7XGaSTxla629vM
u49Jyc7hJN1ft5G859YfjWDd8eqEgD/gxT1nhJSm1Bnhqd4GHa1uY24W0MYGZDST
aFQRzmeWt3Vg3iINXBTqdKQz87baCe4/c2YHCFMkhcPVG41w7PzBSlV1LjqYrbn0
cirnjsBGRRpC5ymM+7tDbfeL4R2JjV0tiIutKVXfB3cfq0fJmyz5cHRD7VxGNlcc
/SsQnJxbFRGKApercwlF+bKWLhML74VCDlSBLmF5oOWVxgb+KXHyjLLgHDtz68aN
xeuiUvbEtxWzUiFu36HoyMJjOsSggvyKWwU9xFrCCmakKR5IXdhQ3znvB3uwt9nL
xix77jMaTmDuKcC6U8/GTF6Z//7zA9/6rcfWA0cgKtDPw41P3GmDqQnHN8Xh2BNL
ofx1oqkF+HIi6ez8oWQCcwKKG7lo7LvK2X3V9k960SzNfiOkJz/X7fxQbFLAEMrS
sN8tnavy70dFsGu51GlBaRaUt3IZvHWySVrBtV8ww+HtD5hFQBmQaGN+rvDNawlC
NU6z5BCxWoW4bKIm+sA4nC00dEzjkxuX3fkUe8hspXS4A9WUrr7Qth5C66VLLMkL
KiQceiX3jaobp7r1RJgUCgj9tlwxnqnuhz06sup456cVQIId395uCJ4jgc/bhg5J
XhEYD1ExspxZwj8fPc+GFUKy4TmiZU0fANxO2uBMHnHL18zx4WpIrdfEMm4SMzCF
o6SlnsNS4GCoy6nEU2NJcQ/ldH1NPuh8PohgFqfLu3KLJLu1VMferFxxyjtWM1rp
ree8acxIlzaurAd9oZAnUZzbwwULinVKI1ECXV3K79haC9FCfogV5iIgPE7pZxs8
T5uYd4XFYEjrvt74YS8/qK7X3xqi4xo2cFUULZeVQ6pMx9cCGLgCoGEKrod1u6LH
X25wVh856cE9T6tyjDvzIPhM7tBFisd7pH9lJExnhRSiiM1MjFFVVQilPI4khyuw
EZoZDKh+yUAT/0TtpJ5W3ItaBg5A2mCkzE3nde9zh/9OybT2K96AVozZcQeZCmpE
OSJYZe+6QoAZeyg1wQQmyoewpaStxT64gFNYpsepz7XVZ1ouVhN364lrts4j23p3
29WIo01FJ2hwUrGENzTiKD1JzsPEUtfSmCCl9+bP2RQ+alnXPBMALXk9VZ8B8LYK
jQaTCwWsTzuAanndP8jWsehIOB8HLZwZ56B+fzPcedXYgDE1rrV/FTSUTDoTX1ve
YJ2oDwR13quuqcNPSsbhjbtiwvihiZ9yhX0k161mDtFSqQ37q+4DywZQ+qUSLEHU
tSHYNLBtGMvTzvyYVSmFNzPL5/MLZ0P88aUMN1e4HUm4XlDWJYU2OyS9hmTIcC+h
EQsUIBK4vLrzioX8S5HicWxMmv7nd2JOsWSRfOxK2F6XHdxTU5C96cjtZqjsa0uV
N0BGABvowe/wJPhc/MnVCGqdJgbNKaA1aXpOOcdXu4PHj14d+mL7kiUqbNr+hjQK
LSTT0stVfqOgUnn3X4o2XmmLgvH0LEcressg9v6EXdknQaebS0o8XSd7i7w1nk+I
XP8A3rCoHZMioGBt4TA+44ogjLUtCPyJUmfXwKbc0LL9mi6OVD3v5q/vnhCCpB4s
7YYwgj7fEluCicXSVZCg9zrzZIdIWL3w9aQC20aByBbdL4P1VDceiodFZvzqFGoh
VCdrq43GKMr4QkTG0n11EmrzPAcJNobc2T1RuEIAbP81zTux1eN5LsTmFTue7VS3
2m+w+bvSPLwroGPIPM42E7o4M/VuBiRA0beQS1z7M7gYUee9awSSAPz0kufsPACd
4w+FBE62kLyz54CSYAjytU8bbjuiGgsVSJUmZHrzvOx/K+qXv7gvxOIwNDz0Lw7O
p/W/KS5eU+FI6sSF+pz3RdzkKZpXcNWXsoQ2RvmtQABwwmJczH4evH5GAhU25CDW
v6FKYLd2wGIj2l0frn/i/rnloiy9vB1XeUe6ppcRunS5lbXiiiFMqIveFVaC2l7r
B6rPM9l6QwiSXyCI0Hwlb+hfOJDum+BkoTxFC7Y6qSJtTVoZA2N0OybERSXuIa7z
1IkTCeoj6EDIxX12VEJY6fKV23GNA3mIJqvr3mhq+hw8oiv2oQ1SCfS/o5pRuEYa
xMb7ATRs2ea7wyy5LuzUqwUFRxaZZjP3rOx7j3R8GaocMo0hPYCijl49lmOaN2ua
DUzXzvhM1WSy2nmFHDVtj6RsZH8OtXaGAdhmjrfNPniHyGCM53gRmd4PsbWNjINq
WqXRLskwDLR8/jHb8kCw7QuESEMk0b2Y4cX5/ccWB6+FexHCUTCIbw5wImPtRRyh
xogbJRwhhe/gQtH/TxaKS7mR4rIGrxZKBhusD/5jefYZmlelHj56iI6mRcs5LAPt
gnV6fbyi6uXYeVhxiatz7N6dnAmHvcEsNEuB2ezS7qr+y6uLX8zfQA175TzPEYJd
/n6eKDOAdqSYuWRHcTn+LZAtNlFsxS+oCxHOEZajl5BMhANZ1f4axc7UvE1KSgp+
6rknqa9HkWu+pxTWhhHjFlIH2QO1Jj6Xp46cHoH2N4f1KZaFpKBZfyKbhcwsxsDq
QXUYsCV42H3gLMdAQLoQdkU1at+yuRYPpXIeMS7o9Ot4Ys8MUKN+2kkL2FxZ0feV
YhnbTR1OGC1GH/zw84EHqP7oo4J/tILT2URlaDY0z3Y5uVzsYz3ayMfl9dNREXow
VSfz1vUFopU9LzL12dLcQCOBhGOGrnjeQo5XpEFofb4I312w7uURt6QcLiGnXrMi
h9/LlsRqLsFb46OE++MsS9h/LViHJGLT7/hqMZ15lrwa14sBI0lob0VX4/v7fMpy
t+cVwpk1pCRYH7Oj6RaQscpRTZHG39M2AUFh8Ob1nk4KTDHJHA7aVIXX7WrYHKI0
XU+P5CFfMsDytYOtNkUrv0/5EXHnLJUKO04DWzJk9jS3ikh4TUUC+AUKPdnkSqm5
BNuRVJND6QOFtIduO8So+lp84baZ7y3EJnuL0BSxhFdAT72RDRjGYgjuC2mWwCsf
6xmOLXpJX4kX541R6d+SHV2/VMNG4NLAbheyYNSaWXiVXYdG2TyCy7G5PhLWcCoZ
gDxiTPjz1PNTPVXgIyp34vb5XBiINSsHvUnOKOtUCd/SSkdluczCijp/RWdAo7ug
KQJcxjoo1NcxS0CPflRN/D/hHOJwpOprZIfhIiJuBX1cNcWxu1rNEYrI/WGohLZI
PqyegZgSqU70dbiit9udMG1CGn0lu6R3wnKbhhyeegUphLkS1Wl7DlE0k25WJmkJ
y9gADiWdbMXEXm1DiQjx+yplShpHssBbNvsDI2lYR1m3U1eznxTc0VdUgM4EzYEE
ZpwAMGMBz8zRMzvbvpxP6qxha4YbxF2b/25Ysfp8jQaC0x7e06ueIF3Jy1IH+gVW
3dwLYxaX3jaMXAzyHhLAvgvb20jLFA5CNsJeXqllFyWEvSA4+q7B8/Pc3Bn92Ngg
5YOmzWfq0P7PnPulzEqcfYDUwUv2jehi8xtFzNoWGBwxNIG8/WXDrjVeAnE3OLd8
r28MqbaHQIeIYNslU6sgJsRtEfFFLX8NCMxT9zWBKujHkF1XVrhBzuvrEw13tV2r
zI++8o/dBL1RIOJAvTW9kgAQzEFCctBipKRCbhoWPGLgTRxZJTHE3xxvbqW/DVCN
e7lDsxA2AasYOSDJWxBVUeNeuvq52Uu0QBp7jdj5jfP54YtP0e2iGkJpAuF6AIyw
oO6UqgpMsU3uHqtsWYUOCfM0mbdA5KuqtPVCqK8zApPA5GvN7lQ4XRehpq3Ydqpf
PoIfsrRk9T+ov55tf104THPzg3YPx06subqUmTb4S6dM2kyBWk9xTl0+9Kce6+1Y
wiawG50Pjl56UkoNyOxO9KnWJLryuZOAD0zz7QQIHCiz4ZYd0ZbhkwhFSZUsmPaD
ifPoeozK2uuwek/uaVoqtUiCC+8Cjl79bY/LwMcR+pWPmRLBCi6LiMo8WTAolmWz
Z6PLEPjkEjK1ntxprGI22oZwgCqeBQe+9aLWpVG9QZM/2Jg/PtNDwdJ5bnxUoA9g
hpNUBgUG/VvqNwQXflmFZ5rlw03e9uIdP7Et1SkABnWigRYqyNcySOZor5vDk4HN
QAlHtqP3MbHKaiQ8/u3sfINd3i3hx7uiZIWhHFDPWdDU85/u740beGdRoI8o2rMW
aSU+zSpqk5SaF2j3xbv1F2DThIrem0ri/B/u9gFDM/oPO4UQNZz06y1OXXQW6v0s
kkSF49asZSCWrDKnjeUy0ThxT0l07gPsuzvj4VAqbNEDjvN9PYRHJc/sra4V9SMr
s3odqHYtS3wdFpAsNi/jfqtyW4Oo498dzCzAorw6ALsfRnYATLSWZLiEr4+PwG1H
X6nc8VaASs89lJ3JUiTrN++oZ/r02co2IcGlNcHQziru0IcD3KMae2gKGjgGkZyj
EJ+hiwj2t1s8C24Oz/dB+INZw4Z1LuJO3ZxlUN0LqXvuiKIRNlTf/a7JksdZS1bU
UCPGBNAIHNckYY6NsIqdgGdhcj1KaB06LRHkCB3Zea8rcYrXgd692sembdTqa6Do
PsZdGnhAhbHepD0SUwephEWEfuYqiDg5c0xPnjNbO94phkvg9RoSV64iJb1juCLc
vJflF4vhJBqaJzi+rWNCPOff9DivOTbHNDKN5M441UDjEWzknEAjBZzqyAsOyIee
UGbQSxwnWI5zyKOBlfuR+pCW1AQBUmPmn8lhN77RYg9QxsqAqSPC9eBDI1lkwNZr
Mtk727e0O/hQaeCOdu5JYqbf+NRp96KQ6eFUcYf/za7UAZE/WVM8HYarggzhiCuQ
ENQ7YFeJuCXbQIOTAphzDKt4adiS7fbNJITyMnWawEMT9reEmhwlIKbBI87cHG+V
sYXDH7W141lctZKowX5kat3HW5JZkAdblMQu5amMtDcF2B8BDou2iEj+erJFK58I
f4shCMBLXWqYamRjsVZwtKAsA0GQxlVLa3h2nl/0N6CLT4efNMibg4GPtakyIY5V
BTMB2vRmIlUKTds6EQ+UokxqYjOIz1ZSlYibKgoMLOhuOuoFzqKBD3NEZjLJC19o
QZFKmmK3E+UJfe/q+63lDcJSIjtAdquHzc94JgTu8dyNPnfr/5TgHYn76IP9S8cD
2UbnuahaneV4CbJkm0nKZ3jvvPFaFbQ6V3zYyumT/VAaZLL3VbUB3b+e3xygtsWv
ZAbIgScCNOvUd7xwxuSOeRmsKeGHxrO+cWS0bc/MLLVTzysiaZ0tTotYrcJfKbO9
Trc1gKmcU+pH/lhNTnRrEbXMnFdKekgu9vb3LLBnxaQFno3TFx6r80T/nCnqf5hT
2b+Hw6qMxjZ9Ugt4QABxfBn1i5qfWAhhzMTTinBKhanh1j4q4DM3e8beSrK169/k
thjEAV0Ha1MOaxrh7DOfVKUtL0fri6cgT3fSESqD4PYwSyEDBvoeLsbh6qyu/xR4
gyRylqAsk5wvWq/V9M14/YNVYHEpM70jxRU8YTkh+6SwOp4k8nAxJpGFVZOnzoxF
/ZZRS6sWZo/edbSTIDwrxsUHcKW/CUaDfH0pIcUlnAsfIX3Aat9ceWmWzszd5Z0k
nu47iP9iUp4GrVrL0oAJF31e2xEoY6Ogoz8Mdd9JP2xDEEAdJs94yZjSPdfKj4+n
G15B2aNYFwlP60uRGM4bbDzbHiEhW4PntbaDH1RGWi2zWQh5K6vUJxKMLoQ451LG
NMUOE6qkAPOBcQNRiiMhqGInJJ4ybu1mk1h65FftZivDKoTSgP4h7j9Qd/fUFb/d
CjUJy7xyHT/t5zwI7oqbuXDiQuX/qKkZoha7daNhp3RhYZkVSX3Mhei3+3LvSQbM
dvI8hkRHKJf6WvdA7LxEpeiJkQLJ/SyuAY63b3YKbWj91Isv2mcVKFhaNT3/1Z3Z
Rf3hjmpcHeSBFjzu88TVeXCuF2MbMsSiu/bVMeEzGxOK/Zyo0PcZ0dQgGy8tYW1k
x/EKeWQOcc3psGvDM1LnpwzX7nslJHf3TktTZnXRdzYAZbWdbcpTJvk0KTVhxp74
wQUghlQBgIV6Amwhn8r8ApxY1vK5gIPWv30BPcs9EcCAHuespEh6jYOWlwVosczX
eZ73riTkTrHIguuNPpJAkDz5ESf4HVl7BzaNPR1nNzA5+qLOEFPxczzId7IWyo3O
7mNE+XOiZSIQ+RjMrmGYVvfnDxD427Tei1LNEs6NbCfKPRWEUa8PgzrH8l2Pk8KW
DISQi0GPurdA0Tf4iU+HbGlNIYGfthcD7tUURQ4OpMork/VPu1jG4vt+CaMj+mAR
9s7+XffsblOIBd4Wmm64T9TA2j6PN862rhCnFPxtnN21TivLMwCuiAIq1Uuv4+gG
ygquXBJXm4htkWswBEIwuQtWRREgMahwoYgw4IiXfYKeKMrjWoxj2vETqGWYP3/f
qlMO4eH3p6Ic5d89Q6hLbkPHVoUaTrVqvGuPBDiRc8t2kYbfS2VKC4d5AQNmQwKQ
/Uwdd4dQ4k3YKeOAARaghbn6qHoPcax/Xp6PG4q73nHfcePaODwgfwhO0zb1GT9/
eq2QsNWnhu4g1AAQCXWx5rzmEt3j2aT+b/OTrZZyLsOwwUfh//EYMbtyyx0CeZZV
X1t5yRqr8cvoNURm5ZuZZtogkoWa+fBDP0EL5ZESXPglv391IOcclnTMvzOOZL0y
85NbC8CK1INGYkdb0VTuI7MU2LfO6DTdulHvqx7H3wwK1RL5tBWQqPyV7+FBoVbB
C+x/nFWgv0IKY00TQuWmRrgFlDmugxOPXF/or2vDyvDz0Up/32/yCnrdAWTQUkkx
XYmPsS1GB/bm+BdQWJN2zDFvmu+bC3hfwQ2VS5wPHfcd/SU0L5bbwSNWz3LCxOBH
JV5u2aIGpoKZVdHcLTtu4IFZgmmP7oz+K0ua67vMX/6CK8FjuNaAzQFgPTSwdKWq
9QUAXyzBIWdA8dgN0H4EAWlJu6+eOTXNMvN9Ld/pTMZcXmZTvuyfNeVL5Ut66gma
oWPcgxGQQV5FDOVEXML4e79Q31Gt60HOmCSOnJlCsY2aOcADlOaj+p8W8Jx7zDxW
KXllk2ToDJK5qQ3T7dZJYQdOpAagY8P/0Vwr/1x+i3jk6stHEJehJSekYBA/f5Kf
r5+kw+v+FLse5S0SPGbi5l1yrRbU621qUKRWd+L3kBurLEPy5yAvLPndtqtx47K0
udYs/Z+oiFzU3+gZcUJtCyI8aAKG7nb/ZXSPOl6FaFaVdgul3TL88QZdPElNzpmw
5Pz/4OONPRcbEh0l9bhkee90rq0nrlv6Rl7DJcM5nTMqKtdMM8aWwj4jxuCYvL1m
V3fj0z/UuD/+DeeNmMqJSo6NO98Ue1khyv4Z6E+vLOPzPXI+Vl/CPQxWihcZmYee
cVDh0UGnURhQZk+4Qx7r+5/bvRgrghzKwcUdUVvyUuZ7W4N0dy7dXXx6Ah6qMcH7
tANYoRLCkUmsJ/5g4rAmqLi1Eo40TS2+Zda/WlYh+jz6NtbSEqXewdSfxkalvxJP
eDQ3zKufv/AjvNwR6zBve25yI+e372mblKGOfZN4JOM7cMIDtWzZj/SKZYJtEGdw
iHTQJFcnr+4WIuhYysacUmqqEdNkWaxNYHr0e8j3AA0JiHS/2BN+f3aFBiZ9JnE1
OTn7sJk78x08PV64MU2URpXXDQR58nzAJ4rA9KCFnx0eyagze+mQXSMAvFxp4tMm
nknol9BT0mD/LSQ/FLs/iDHMQZEXf0n+ZfssuUKBNlCNl/XT8Is++KG4MuYnnW8e
iLnEdzoVF7+OrhbJi7F+NJRFcd7Xbufp0Rl24QXLflSNSNaKvRgQ57EeEHRToWBM
jcqjFmTOn0fmQYA/5KyxTLR4zxwmv4ySbqozIZpw4DturP9XYXx6yN4YUH1hOPmZ
w1V0NDl/q/Matjr/KpZ5M8FZ2rmbjHDKgwdOBe+ayPT4LPQNrm09nnWCxkNnxcy7
PqDFbm0GJPx8+NK00BV4TirUoSWmQxLsxD30+ThClCLYa9iLoRQdfwbZkGV2fCqF
pkS5Qn9kfVixHxanf8rbt0uDIRvXaF7cYB7RhUYwqnwxWyC9q93qxuhsC5pqnPDu
F61J84sDL/JsnH7XDanUZBa0H0JtGya8G40lMMAh9FXHxnPqKWnzq7xE9cFcIpqE
u4gsXd0KUDt4J+CCAPndAw5fZSBdRARFqcd8vgc2AQ030tGW3qoSTKOeNWDXB3Y1
u7IHJIkOsfaWx3V0rHVROHjLOAlNtZzGSHCY/ZCDMwPl+b9pLl/x8bxG/ShflBV8
bLdUUYGEeIBgvTIi3R08KIZntCp5tXgIBAwgUnlI9bOThnD4yvWqV5uSVYy8t9yu
MFXqDDsaV3sWGXR3YAJoC/3GT4ksC7icRPRsUMRaMtbBTD3qqUJREd93qp6OGPeF
z0bPJPdGqVlRtQOBmONtEdsaAjThXsSXPn2jgwZ0OFnRG1gm4KJhVwifPfoMyFGz
NSZ+VKrR2jL1V87cpV0yGcJco5k4RM6HCuKZpfT3Jj2+XqxZRe1FuOZguRn8pHW3
MLOsfsxetPSDA0Nwln5aHe+U+oZLVnQA4BUE51u2FIrqU16PY37ux4tN1oh3K1sG
xR6rZQDcADAY05b2I3eNe0eng3C3nq4NVTOvr1DNMsGopCx2gSln4QPb/0jqzZgu
v3YU590sGd94qDfjjcaZCcIb4EyMgl0J03LcEwdc0Fw5C3y4rRTdYEFSJrSmaw73
SV2sZ6rw0CEsH3YVPiznjPq0nOzgC56MGY5tXjupKCaESjEBCbCxlL55hpPXWrsZ
SZBhU8P03g4ZlF28DtE58lFGsUQfRGyzuN8KRgqZTol9qdwhTEChoNjN5SLFm9rj
CBQ8yGdjzokss9pYtgVjUVYXcVjGaaS/uIGyyHiH5dfo2VdcsP8gU/BJ8d+fKL7y
REX+j18nZsGI1C1lYe5nxxpVoawcdlUGDCwxPtdXFXA5C8Ke6+eJOMXNzywTrA2F
d9xEXUpmkMP+FPWE+fYKiWVUd2jEGCPvR4MJ6veiipuaQd8WoTcnIalzOSR9KDJv
zxIslr4tUE/EFjsk3oLfVpsae5G3mDD58KYgbv2BAYbuGimrqmiaYulZUj/HK3qX
k2m9f0CxKd85V+ycw4UHzaPGfQ3UAt9DUCsoHDhhRLtkpfzGt68mVBFRucM8cTwV
THJ03OoC/RqC9/hyzPqIgM+C/otiOV0GWL1y7zT+57iD0aTiz+xIDr21xgrIl4AW
jThbXvdTc5H/dtpBsTNJdfmTckvXhiz9v61czuzjmNnk/WQ4c/Tmktx4KwcqKV8x
ZFD5p1nh/og5moCGz/xMSvHPcb/dMWhUpqpFkImoLF5Fu2urRvR+ZKwkbD68ioTr
XFCWxpJJNFsxjoOqTHzAXAQImi80paZo+YDNgiPQVhLcT9wWOK63FuylMkwlecqE
B8PVctKqCfIGg5ruObMsHJYst4SmHVLKLuxnuCCwt7/WYOV9ykE22DtKrYrnSDFe
PdCERA67D8pgtndgPoMzpBAxdQhx97lu6ncAK4fFA2LJY09c7dsm0DKVVi5L9m0l
KFquXEAB6emjiJPJtqX38/LgGKEp/O+oWMHp4e1AQJFH4OX8nUtvF45p4qugOhDA
DlQrz7CywCifQllCr+nKI18lxJsrcikuFW7GC4VOxlOQARnBgP1axSXcmJah+EzP
NT2hIzkvdJjoKyohNQWC/k/1KYb9zvNVY1vE0/viGyg974bEkmTsfyxAt47X2fSl
1t4d8iA2JFvMqImocBae1a+yk78AfJ+qTiZjSE6vUKcdHVvGGY9uLU2rmm+rhQ+o
YjAyJhJ7/rwHRu9TOxtq0jfE+M31KytnHZCdyho9mQZIUjdHPA4eov+HSBTlupef
MqJegNnsERBzn7EQFCKqdlnklxkG4GZpNgg2eb0fXHkGM21oqLT28FIo8Qkkvn3z
3bEn6uHykxninOAV5PUpmqsOBeuWO1nQsNau3s8gOvWqbWV6WeMVTDUOAh7KikeY
dDqYiqrnebgHV/BaIPEQi+GU3NEuCQNyBc6avJ/7osyCDhEI0EEA7q6IrQ20LdZW
oG5lNSyklfUGRfiRXciUhBc+3JC4T7Pje+kZAXVb+plx2ayBSCXVWJzcN7DY7kc4
L5E7YbJLoBpfd6VR432qeIAyhPqxFISx5ybg36Oq4taxrfx9fz7DAB1X4rPqTj53
zmr2n0lv7u0QhT/PjoL1Hc1EqQeuQgcH+GMlsxqCeeYzDCh/2r4/97ilOjFsREec
1EM/4B3nGs8RpcGE47ZyI/EYcUSiG6V/abN/kEfoMU8iWJZP3PfFxvFE2OjieaYx
xFRRzphtYQhqYsd5/AQ7wNwPOojMlv3VQqqzoH2/ibp/abAzv1JuaIACmpf5It3G
COLp9Q0X13MEfvf9SWMyZKN0FjwEiH3WNI9/fSF17dRND5Q14VS36tA1y772mzsd
Jw47Se96tdKCyaPx515D3zd740svM+n7VrwMCNyWK1FCTS5f9rGpT8mBGq6duHLu
CGbtCSstYyySWog1POm6E1Ez1y6dDwUCI74eTxSijQ+LzXUHPntMWBWiObNfBTBy
9WQZqGq2EJJn1LkKHCTsF5Ox0mxPNVs56Ch6cfzyP0yF7kb7P4GWZ74Wia5HcIcW
HNmKfz0osJnX++ZvuaP9FB8fI6bXXsNjUNYwaHkLk2Jm2OCltCRU2JYwx9kNIt4j
y7rTgHNsJdKn9bVHjxG/pkoTqBAzc9jHvBFsWrF0IK/bFfBBPTtWEI4EkXyS/rKA
EagqXDlO4p07eoNQux6meG8ugHqlJmFGWgtkjtlBCW29+giqd5C/sWwJK09jQauW
nf5W6MOiVh5xNHq+BpyHKPm/oaA8XgIDIypHnlTB2l8MCquSHTkHrzZ3JjJFAtrd
bPow4OM/t0vqSk/N9yBoiowC75KPabmeN78N/v4LM2XlWioAvfbfh90W4adBPlyJ
tS7SohVU4EocdW/CzB76besShkITjWVenaORGQlRYKrDVeK1yhXOuyxEFhihRJ8D
vFUYSrA8NRHyg6Dz7Yn6Cp0g6W8IPkTIPqssSqB7NWfjhOacAiR3g0ZwB+0blZ+p
AjdJoffV7DBqqz7yHanIAMkCDO37Jy288ThNIxCvHY863CZOtpgvvc2lWjdFTrQh
D6nF36rxrOlXpex6m1ZKTYk+94Q2YCmHPNIc/ZAwVmRCfVmYCdRhq2gAOxAJIJMA
w9ChQk3dPLegWsWehKUATfwYxxur4wFBCA/7Fomn8dwgYM3MaOlP7TriDHts6O0e
qDm5U9p8+oqd5mLP51f6yBtxY6rBw0+191JlGB4UZjJzfN91fAHdsrl21MlDST8V
CLE/2PUc78W4o0BbmcL2suEc6hb5fD//QLaQ9Jr1s445b0FOwxw1mBhmPr1F4ays
GkGUn4MT9NkxRt0COzMC2iOQpf/bBxkB6J3w2ajclCr7N/y5o+Is5LYaieDigUzg
wjhHh9UGSm+ntQo+XeDjWav9VqLgEfg1shHFki9RthKcedtmLo5mWP+I2S3KKbRA
JRdcD8SLTensciXLHgUVe5iQCPpDGORM11fzNKYzW5VHuEid176iO+4S9MoX1xfY
hiIAERV6cgwoVHpJOja6B2YNoqBR3M95mwhDJkdGBmX+0rMKzR52Fd5vAIRT1dw/
MQKkrFSvXbKjP4n/iQJoaFv+kJeK2+v+jVSexX2TY0EuwJM3n8rpQKusUYEgaf4W
jAEYs77d9JVEXtqQb4+v392R1GXjGgULXLoR54L8t/+TaJxCDqgARD3dqrz3Rjqi
WccjUiXrvlogqriAznFOHmNT4Y7ljejbVCefKsMzGlbynrmkg8ABrk9KImwxnNB4
TV6JBPsW9bs7SUCQnqKOWdsZOZXlUr6jjOonMoSABA/DkI0ie6poj0N7za6OssmE
JlCE1cK+NlkI964unEk95WGbt0TzrMhbwd+r8jGX/4HIwnYfIBGbqkK7vPEApS3u
R9OuS245uXRhh+5rXeyRdDtXZkZKmVKOPHxG2HfzhUljAELCPhaQz06yze2KDwaY
BFX4i3Yo2nvezQQLtGHWy/yl//zx+US8/ZcqbyD636MO8ziOJDBfngxUSaUgfac2
Su2Bqj33BnZimzAxBbiDSSOb/NsJ5R7o8loPcilXnfIe1RBEmy6GWoU+XzTtcPhJ
ahnz2EfHm9flEEDfVVODP4LR5hH0OY93dstTrt6kt2X2FLj/QTYZHpof8jSXP09+
lC8AbAkClHAoSVG9fds7SGz9JclkrzYx6BYCjmOnmwFuxdPpD8W6jCqDJ6haeVjv
moNcxfYZVCjnK5VvWQrB8JB5Eui5nm1YyOnkFZ2LESghLb+6qj/PeYBbvFkQ6ATe
O+DGIOZrO6CYhwDbOheG7CQWEtjAMH0KxW0aqWFcbSpuAJf1F/RHyXQNa5ArC2EL
LM/JAKbtZf5S1bNklFt3NEmv2+kfXM6DRUSAJfSwj39li2nIHWvsMi+u/qNqVxXI
Q2pm6ILV/mOk+ZMlCKCyFVcfXJMFNoK8t99qL9THbJThrSoXO7xEJBz8fJXllv0H
9nNBs5v6MnfCpwXgNLEuGO6YsCPSc4kTkSQ55MhhLqZ+9dMxEYYaLg9I/bz1X79M
pSQMe2/vo47cZuItHv8zqUPcVji9ef5KSRmYuybkq8IykhuwqdmNwNcc85C2cKzw
ctK67LMkS7aZ6tVBZZjITMGhoLRRPH4wTgQlrZcLneQg7UCcU3XOQT7Kxpj1bm6R
je0b35Sol4yqhii6q2LXYXI4Z/HOQGoc/eJUbaYPZn0XFpeXoSMlFoqwfNnNeBqp
Iqf/AoALDLGv+FzYyNnwy+1V/VrDx9lnSWHWOG1jrQdSD9nePn/D9bamuEPhAjWy
QX2lEZKvM+O7ewXtSkhttJTly86VLZNuHYBq+2JizbjO1ALmr/eLwhbEj7/KJLVO
yBSTdQlHtDxlQ9emvRG8+Zaysa+5lfHgW27Q2s1rFSdwFooC/qu8yc9tevijNAZL
wRlmBexo+vAJpxOUpnHA4lqhjs7Xsf6L31pcpcyjk7koy/Y4S66r9rfMfFsrkNAT
Mn2yy+Oa61hi0o2XhUPw6oWD803XkKIHQAZ5Qp3gxlo3wKEkc8dH3/4dduAdv5dr
Tj9ddMkzQLB2TdkdZLOD0p+42L58aMCET7AHgUqCpX3qJc47wDZk7haLaUDZvDSU
YSsjHPm0Y3d1WgB5MbXVpKGlCjzvMqOsLcpc7zXwKIgjhWIReJKRk2NI+fZ8YHiY
gU8UKIifkh4g5JFK1CY5lYHAY/C2PiCn2uotl6Cl8yLNRibjFQtjyrxifoi4RlH0
7FXrUu8usTj8e5a3RmRnT3ltELmV07lRVOvmqvTPC4rX9mjy6vCPg2oN1DSe3IAu
s6LsRBnhZSIxTibihwYDp4IzyNT/v1Tc4PnhuWSH28oXGAviHyab91Iea7v66ksJ
ze0LwUgMVvNGaES05tUJ3R1T/KEMmZGlnqGpMRUQkOzr0+BppKfOt8zsuaMF54p1
3E9QMzns7jcvBWgyzGkrOZtsJwq7m4eBcYMST2ZeVXjONsNIWUDtilQzqNaDXy8/
jt5lK1eaiREaUMpJUBbw0k5eG3Jp3B31UrM3zthko4zrS27rg/prIZBABfqLFMxb
cOskNq0VFXZlG7K3Cuoz4rKxgc/1j/namBXXSX+zU7p5PX/8HqfF0kFPDM/nIm7H
NsA2yU4khZt9Rw6O4F+PQaybmr/2+O1rYa5hE7oTNH+zi3ShE79bFKUu8Fp0eRzG
J+mFmHm3eRPQmHNOZWzvIJ207bM1nATgClbraDy5053iA04Z+Z/Jrw4iNnIERufN
VDAqx7FydPY2HWWr7JV3xY5L7+7eMn0AaTBmleWyPq9MXDLaDi/N6ty4/bJ3FMhV
4aYft2/0K7LJo80hRgM7bE9Jst1zGAxK110vw2UTkDYjBM7yKxeN/HUHjTjkiTQq
hhBIdNhWYuGj6EsgtAqysCV1gDGYaIZGXGN46Lqk+UIn5nFoHA0L3hAu8WXMEGdT
NRghtrq5OFJuOAallG352+dUVaEPrKeuiIhWPQtgoOcGuiads/gDyVD187ysHk4x
E86wMF9oIlZJyVsMkzUE+SjF023JLroyxiPuwaSiYVVCXxku0yTCbY6HKPDeFV6S
vgje0b6vg1wgpEDDEtZ3oj5gDpHk7QZ36vgZKatAoXKuZp/0ubGSTU3xLx8bTfKh
1zgeJTFr0mGds4mcI7hudF9E1COu/ea0+zq2zCj4U+l8RIqrEvexyUk6mzdDOCkh
/sA4jtfBaZU6YMuL2DYe2Etrdh05cNs7TqvXAHt6aF6XnXaTOnhPp3LDnvx4D03r
XuZ/U0tyPJ0REMQpRqH+zvdZ2tJsr/1jJqnnzqckRIwbb3fGaTaBk25NDLn7kymJ
I2zJ21WoJw8qlPRnx0IhtFBSTmrRPVSBu3+X2JSn57Rz7ZwR+PPpOu9p33TkNn/w
tvHiu89o4SVOl7DvmK/YUvysZWKGXAk9PhNgradUF2aob0XF3p/DKJJaJtY+gH8u
9shV14qllTfJa2xmm/CcFDBg5A463ztixs9kGPss/HmlvacnkskfY8PfZSQrhK1m
H63Wbs6YerZQj/pmbDtcAnPXLv4pNooqXZPEyQW68FWak9GNggiMDahsPo4guOMh
djg4wII8/wdrVcFJ7dg+A7CyIQDOCfnd5Ta8JjlkIP7EkAtLP1UmbB4EFHyx99Sj
AxX5opezNtZKVgsDBq488Km3HK4DSEHkOHbEGs22fYl9lo+WwdXYcUKa5cE7EIAH
ojDENPFbepzTrTqh715iy83HuJcZ4tAxL4AMOMvM9/2ncLGCf4CnrXiq/CJEz4rM
EGK10KYgDXabT+lbSnwUUYNtnxZBp+OlvnPngj970NBPgOMY5U8PpYN6OXGNkF69
a3gEGsSWN/WtFP0qgXLfa6KHLVSsHL9EUVPF3X8gPnoWpDU2QeNC3OzThGdlbJBs
Rm1kcWhrm8yHWBbpNY1/qvS1gvkvS2VZhUCrIcr5u6K4X2/cGcLDUp+AIy5aXa+e
op198a1xQ3a3QocouImPg8KumDCFjR5apHiiO1N8WuBkfp5BlqnqTxXb2W1aQwTE
7YIB7iEHITSAQHZANczXlGdqQVwNUE9WHx3Hep9nT9Xk2yT+O3yiXumrjkIqmeuc
5BFJlqwQkeKVXpya+Fs++OO+euuKwJb/AootRN4lPnHLI9B2pxhcIy4zlya9eRPn
GJZ7asX56qnRBvP8rhXnBIBn/VDVr1oAzFZG/bpglEa8mqVVxuza2fvlIxxKWLji
vQKwz0PtUa3CYDy5BHXbpYRpH2pHWbJlczZg5lu3Vkpyc8Dcb5EKM3xhKTYJUQni
OYnvNi3gzBXPsQjRTvr+bvnVn8eLSh5jgdcbavqoyOdYsxugHum+kpoc7pyLgFmp
SW0fERkNMOPQdSzES82YgkxglcaeR8mbQDqGvi98pW01vsCr5Dml1yO6QKa8XhRa
qx2mMUbdcg5pJ+AZLedpPZsfHYTwtUekilHogDWQ+vQy3ufPktkAkLC2oN/+KBh0
II3pMnGs2adKOEegar+cK6BWBDrriTZd1FkcJ6RDlC2cjiJN7qoWCNpd18wTkYCv
SeHhwsdKaQPHwumtTF/zwAAfU5XRofIbQ2E3B6GHwKdVKsJ2z+rwj6YgJTx68wNX
/a9PENJgSAJSqGfxAIrEPPF6WHmwVNRwoUETBiZ8MZdJINv5DrbUSyNZOPXHEMod
pnTiHsNR/RAUE2Et9IEmtdB7fIvk9HugArXxuzqZdltIclJeoOiF9l0+ti3hL/wd
NtGaVNszHBpW7q5evi7FluUYd9vaeWCrYheGKCF4RAtCtQWVLb8xRGKBFaoPwfod
S3iHZzVWEPT4lN0zg7eOpRkAaucHH7+niyKH4hU6vpjWgzDUl3XQ+wCX1Yrg7j6Q
ixKL0gZCTPrdXv7o+nHFbBezFodtzXY57PE+VBH1r6vro7DmHQc0sIsb1ihmspFb
67WHo2Lmt9Ewry9T2RYVPeWkmOaKngPHOx9r/lyH5AmTougDAEIlGjAH3R7ptvBl
FminQRwnTNWGqYE8OfsBFKMIS/7gsi//maaReacjknOcKkk6JxBQta4VGm0yT4cy
hbCwk6U8lfTj1sPCKNeIF2kZdMNSmpdKBtCGJ3BoGe0N40k/wUcmMQYHIpLLROHL
6GY1Kmsze6Igsn2qdKaKwk5DK04dcLguZHldJQF59YU9iodaUk7CsOThUK0TgLIp
B8Eu1TY9T92OLRDPhpceTBRCoKk/KOYnP18RORZI79jnMN+pM7oaJq5JEWYnZ5qk
NIi0o6h/Duk8ut3L666IiQhC+VR1QjTX6N1zDXsRenDMhPDVZ6xuWV54GZVwEd58
Lozh91Qwss6m1Q5zO7t6wrwsgCKCF/Vt4iGyuRh9NVcI8ftcuu2XRbhDelb03wOm
uaGq+BhUQ+zA+tt6rIsPWBAFvJm2sXqM/LMS8igM+rq/mgRSyEr/CKhUZZSmzusX
Q0/QrUNQQYV/PgU8SNzy4PKTjQjk3qUe/UzHQU5vYek406192v8QG8ZJ9Xe039Ms
G055WGzPtU5uFaHIflmX+4g763qITH1nbe8aK9RMn6cErexDbFgVzWvwds/izYFS
sNAoIAwQpbiiagJDVnDsNVGFq3UmE4NCVlsJqJxNUvh8ZGtBGX3kVtOkqeOMJFVp
UXJEtpEKp+fZUnwNs+SfaS5z4f00U7GsW/0ceCn1i4Jc+GjfwTK1/Gw+CFmJnUC6
q/3+b1J8HCQP0oy3S5dV7zSJyrMNh3AZMSq72rhX2QHveJ0MXPC23huACB5l8RSe
QebplzFGRg58mnJ3oUN0AodzmEhUfxj2aJsJe3Yp1oQPYA6vqdTqSuD2DC8saXf3
d19txvHMZeJuaP4gzQBYuubHbt/SHqSpYDLitsOdCR+A4jNbNqQvKrHgsZGy4+th
w9WZYv0cMdTvV6lqg/BYGrDYP7v2OBP1VH+oB1KfpcWAZjlzBISr30JbDOzc4EJS
g92F88D0rvHidBZUnIzr9GJ+rwAh35Q1Ub6ydoC0pjn5IsOZCCSJCDQBWFmCOqdW
mQS5cGYUdNrIFEEm6c+x0U+ZBfljmk+gxVSSV0t+ORN6LDi1ZXk+6VvA2fZCoygD
baq18XYRhM8M+ceGFN7NiNtgkE7kxGM1chAVp6smK0kALIZb9XHyArqXhEQIiRFe
IARactT/Ss9/Rg+8b3CAfstto7ACytr3TI8fLFe1tB8ta4G2D6MWEmrKqErwDA0w
XJndKpZ1ayYr4KUCiutvls9oAKT3GiBP2DOxzNSx/0zt4dn1qJVajxJ6sTujlYII
jlzzB7MhyjUrF/s9Vbo2JNEXwSXO3vCMznmF6Q470aK2Mo1bnurx6RYSSENNMFje
d2kyvWlA8Q7xlyrLk3we61PTuWHii2/A/0Hk9952M2ryeSgbJ9c2CZJYlt3eN/O/
AmTJA0n/GXseSpq6CJc/8KdNtdsosYyhPUtr9JXW/1W5F/W1sC7FXwVaeIlBalZB
GlVsrkSp54pLQGlFD26nn6qkaLEBMpKITSO6Arbh/z+4I8JlKDDsjHUxLio7/6Dm
CadesKabYsSz2NEypVLCDrhPRfQT7HpQLn+usqO/2C+jxcVi1D0zWzGcoR4wksRg
5v4yASoiFBG5lQ4vGLnREi0Eyq8PCK+okbpXlKEksOnqqmJEONbe3/Zi+RMnWa7e
aJrCTNKPXDJ4bOOIM1JzPN+Z2624jjtT0KOEgABBqP+JobGI9lZZJXusqcLylGKv
BaESO1cd0LXgQoq3QOO4523FTeTsObefU2iV8ItQ6/ZIeOdzsC93kYNksN+sak+C
bMAeHRdtA+urQzuTit7p8p3NUXkEpEVXV9+pHUiABXorZbXUCDE75DjcQ6671msQ
1d4mBBu4/pLTMXJXwK2c6HtJI/uukuoK/myEsEoZayEYQP6XCiD3U8XwLES3u99B
vEGRaMEWnEx4eZnrmQnZ9p2iFTmGOJtjJRxrqHruDkqMNS0K5XM/XLDb7VBa1CC3
94BRx+qZ60s2k5OFUuJNYbgU5xZeXuarqU2DiZgBdLV3UResOBaDanZYhxIaYa63
QdyGDFqU/PZZkmXiakFc1ZNI3UXiTEXvOt4m0DjALPBNMhQmU1uPzCgacckaZzRr
s2WAs2FXQgni1WwVp7Y1AtEIfxs364mzDBzvSyEk+W1f4x+EPDrZ0r2w8oUTnTaL
LFZUTyFhzL5eo76/4ZFpdCGZ8+Wzo4a9oaJ5OVdXaupNQYshens898qwMilm5r97
1yP35vEbQ27Z6ESYrItWelLiDNiwUVL+SRxYpAAOoHZFJE9CyT0upsmhPjfvJqCm
Q/a8NiKWqhZM8+mR9A9/0YGoBDvvAtmQVDqCXxXdYQ9SOEaDZViaM7O11hP8oSID
8WCGcyqt5EV8dTiTQUXNwqhvoy0NAf5wpXTgDB69ygTYhphT75VWMK6nMirBRo+t
dekh/IzEM7Un+gAazpxAPeYrJYUKLoPtFckui7cdbooatFIR9L/XrIVMW33XNo9q
e0Wba6enZHVPpYIr1MEYSM+84fg82knme0Tkjv/CFGXjwQH6cdtUqFGsw/fkchKu
UPBiyN8gSBl+H6aklGPkIhBoUrZgQy7hs7lcWXH+7lS0Mm9zemyrUPQHMhqNbeF+
1Pj6cJhFo8mFqpozTChgq9LjtPebwuYSZqIkNocq0FAzUGGUWsPFS85gTjAvIJcj
l/5DCNVUa9Pgzwzw7x0vNkjANE8ICR1D5J9mpl+WSFPrDnGKSMVhY6mGjJFFM0fo
7+xxb6iqvh5Q+qBMW38Lv4C41LkOizEBUSwzSYuRdLb2n5toxdc0gvsVpmJwYfrZ
3tWRb4VywkCFJ7DyEOZI2VnxJnyfJ+kCdbpfp76HLDxy1R5Ekg9lwd/e0SNBwf61
gJr6Kr31k9LdOgsX9bQs+cERzjgF8QGQdY3lYUcyOtTOanNyvEQES06iXdFQEV7I
dyUexy+cs2VQi3FhZ4wUHCxkCTRw4a0oWQ019epIMoNCzZ3ZYexUtEIwFDNwYgf7
PR3RvER6ttF4r9ZzemQPHZqUVweI9RBsYOky+t1k+Hw6F5Bt4SjXjiBZijwzkxoa
1sE74bcxBLtC588KWXw5Q/Ix7iCSV34FTyI4OMaXcojQ5IRFyWqHVxj60QrZz20P
Ii7lvjZhg4jbLzmhwiX8PnZAEffCXEV8xjTSKndj0vyubs9zDJSYUZt61jpuFhyC
QnmPHT1OEWHfCUDTC62Q3p0UGIDSfYErYz0CdloZ4KWQJla4U5FAjBrY5SY67VpZ
GfHZy4AeSKQQ7FAYboGTak161pcyn7ED4VUUto7cD3TcZg5y/4mc4NtDMtJxoEfd
1VfsQ9WBwZJwFra5AuQ7HenRnLPZ1ctL99xzGKRmd7XntSOZdyMs00/ACIB+Iw8W
nsYQ8fNAeKenDWjiQFES4OUwidcgcK6m2bmsAKVOpz/FqI++i9SINXzMBrjIdToD
T6j0ayIiMCnMv21rpVsBvabyMWPos0ubnnYsPEdNATu73x3DbsC/sLjLr7r+oFPY
WxC9KV9Kigh9DZ00mONSyL+pQMd7r0TXKxyM9/ejsHJZsJYOUCyMWVa0oFgqjFcz
/Ugn0F+B0UZMQ2mGNCvfZ6fqrBboSbXT5cCAXVS7Xs08ExFdyuEiwj3+x6Hj4x7z
XHd4enLhAe9vwrPAN/zHjcQbZvOcYXt1xJEmaxIZTWwlShqBVli6tu+Q08lmfQlP
rmQ5bDtL+vTQPGvtFTnmtKW1XJD5ydCUG4vXxVJUSt6wEF8XZSUKa+bl1uvmSjDz
pO3xzubyUz/Q85OTnYXKzp90vZdSUPdyqpYkdIjv5IR9ro5p9pneZhqlr35UrDnR
lrv7SY9xYTA0B/8r2HMMY9RA0+LNa+dgi5vWgVWeINoqN8kmkm9ELhLTt5o8ofcN
eHrNn1JyuquGhBstcdRHqkjZHYOtzQTQVqI/OmqBhlIpTtGslhFYFZJLLRzf+2NH
rOCgYDRegH+xLOFi0kS9TfqfmoafR5EVi9uvWahO12afM+VlzzKByHqqU0VH+2CQ
TKy0RM5fHMbEMudvR+kEBscYs4rNRumXZqOeZfyL/oG9YtiCeS9G8Tsub2Vc1JF2
U4ubDSonlw7q1HLkPpVWOWz1UrkJ2DzyNmzrS4re0dbEOPjJrONyBP16x8YULUuI
jnN2qaFcg9Bs9VZ97p7n0SfG1HQ2j7G9dxTIV+6boZ2oDmiTqDcy4BXdVaFBVqhh
tb8V8Fo9u2SqPkq8Q3qwcrvNMvr3fhQx5yKbltd28U80RqchPTopug88dl/ZHB4D
xCy0mvunzARHfLE4ZyINrTvz1u3SuhDeMsvN8bCdaepEVpJOd99Wqb2iU9A4M293
3nYAqspF/BgDUMGhoUkYicy+eaXEOPCl6DY3hLoJR9HwhBKGV6XDPqoWaYBAfDYq
eD4mcd6z5UArWnv3v52IfFj1aPKlYi4HWj25NVTNGLAyl4eLluJ+2lQu4kDPkp9Q
Znsu8pHbttRbzPHUNRFfuWGS7gSZwe0CjbccBG+LwrZweWTOEnmGef9HplKE3vPt
gubiAhJeVFmTYBAnnXpMu1JdU5IywM4yOmUWwOmIj52OVMh8gVp56FeHrXGTJiy+
RiLA5B/TSIa2YSS3kThpbcpsev9Oekj9/hwnZm7j5FO4Q1+Senj18SGXwdByeLoR
D0h5aDeUKlqJleU3rQOG/FliqYXUdj8pOxO97z0hJ4Qcsd1y4y7E/NHzYW9qqbVr
Yb/tef72LuxWYpPBYcvkMKPX8p2innCmNxNTwmXBAQMzGSewlnSH906o2gEWaMt3
WK78Oi6BMnIW8Gmt8p05GhmC8F8iE4oCrEA6zOxjvYa/0ib9cIlj+ZlI9zD9XEJo
Ilmy00y6LoFd8H+tlvZFvriIAhyl28tmCHk+dVfGymxC3KTf6P2gcg8R1DmvE+3d
31C8kPa2zxSGIe3WiixwqlO6/0403dWwzpl3xxcfuVFwboKfgCUehlodq95Mr+q/
bbY663+wdYdYA1B4dkqkhSjyKNzyqzzZ/pvWs3tIU5uANj5nDwjeX0imaKJcXf7h
G+NiywGqFmlnaH5bZbxe4Q6mlTvwzOGkBOm/nlvvnvNFlo0VtdoeVpIx9sOjgMXS
FnGqflnxIeb/fsW1KrGgJto0/oJt4t20Ll8Xnfol3hi7HztSq2Nh458XW7VaurEI
xv13yQXwx1YMx1uIhmMLGzWk1Efei2296KEauSDSgJ1VvZY3ajRXy8+Lofl5RLRQ
GoNjZB0Pm14k8pvGoIcygBUXPD7CdTAWb5J55Sq7MipqenQwlPU49Xv2GZLbVfvH
fhuZZFHNdhiXI6Wtnqe18u+29uTNmuy2mfTgRMntz9dYsjLhtsHv3zkRGoMAIp9c
J/eMnhm85J5iTW3s9WyjbGQayFkEYRKupAZ6ipy/XptykVmPZg2KZ4FuuZrRVj4j
MY4umyImlFObttiK1HtZ1DXgVvLP1NFLBFQld1ppn/19lLDUOwpWN2rOuiomZxl7
dJhyOOLv4OPBdPgU4odACmXvMzd+4Qo3hakm9i7fkRmuCIesOVcsaRUYLeso4L0c
SQRh9LWatC1cEsgICCdi4vRVGo0XDW9EmomMyEEqXFfWXOe6tFwgh7ud74lzD6lx
Iee9sp+/e8Vco8RudHxTrgq7Q4NZqpOojOdnFeW8M2S/fkMeGjaZC75xXdQv7KoG
OyR5pnFqRYDJYoFQ/rQWiv87wfNqQex4rGHp4x0TkLbhL36yO9zmnS7iI314zKCb
oYS7v7EBXeRU6g9ol1MBHFgGa+DecIowtqYyN3Y9pko7BiNk0VQJFmF+oD7PoZ5B
D0dighS57CXJigm+OEgeOoLs9keY3s3OGPjEpi4h47uIGAD/HBsQTauYJ1JTxeWV
706WemexDbyczq267ss+geWubV2X27wsfsnmTTUX+9CeoKT2kg2FrWspfE1jw5WY
65UEgc1as5SpwMS294GnhnBVSpJR8uEj8Ukf4LyyE3sL8f9s1i9mfjPcTXb4Cikz
YlwAiYOjpEiQJ+Wm8xtfLiTxAi++O+BNgrvOn7dKdHp5BOpyiFI3kt5kjFqVeQHt
tAbgsFlvc9xvn74FU3DUbkpbbtctDylh8YF6rNFefWSDJvT9hxv/EQbn6PHWqwtu
ZxCk/MRRxKlVG7mwbtSpKfawVDgcwiNpdCvp0xRKskbHKxqwBIlaARMFkt9qW7iH
ww/+zlK1A5P5rlWYwwjR3RZNJvdC2XFz/DAwh079sXwBrzmkp5WTOrNWceuMQH18
CFshpg3px4ge3UBdl4jJwOYsyvxANFzMohwux46T0xqYqrmTD4sxJMsWE6xLbuTJ
1Dzg6u7GdoDmi869BbVmmhbn1LJO4i4ztQnFehb/zY8GoroHstbdkrt0eZJKJuqR
3dQVgVQI9fFR/08CA0SMEkTnKDVu0wUdRJkPAnvKGW0xGpQMhZvtAjAkxWq0VcHB
ZdXhvd1senkh0/ABZNKQLvtzaG57BXO55Jc28DTpw4xLZDaPxG4+DZY6yRzsHeAN
DiOTbgN7T4QZuxDV57ERPGBBZkk73Z/jsf/V0SbYyupOBXFmmF/SRw7bTuoxngBy
MOkGCyDb+IqlMr41iNjq5dWQWqT9b/gJM2OA6krLF078wbkyrDPAl+KvZKsYetVi
8RqxH0O6W32RWtoHoD4sYwp4g0f9mfjqvPpGIyhBYZfGk2bKQ9nZQjhPnhTWRS8f
TMhzAW9JjhGp86LZczDuY39124YKxdQhQnekM/x8W9U8f7CQt83sQ2D0pdkNUqcU
yfQLjGbGVmMzPfigh/qJ7NnosldU6eq8zxOcb6A5j31ewJieiRcs/vlL6zoaX+tJ
sjZDf4EwnZWNXWGVCtQtg/SwON1MSWO7hVlj4UiNFvDXaWxUdotNhGVw9tqDZjQg
arxjLk9fKiFMSKJWyHmYvAfpkE4sWJQxovnS68zujjsEq/2oDll4PWpnkK4tvbOg
s08gdMvS9YKQ6z8PzagTNsD/9y1POZa62xuSAfc1F9aISukMLcYMPHn+x3bLTuzN
UjLV8DfqV1JLZwFGgE+bcSZdUxaMIX1lNf8l/lmS2YnRELy92mdDIH9DgGL1l1mg
hAuPuDzrCTJenIgdvbikx5HiiJ9X/T33Grbp2Y6WPWBjxQ3/a8Hrqw4e4ApAHUCd
U6LNIIZP3/DW4snT87qyVP0+iAlTvk1HD2UNe8zHLhjpqLXElgdy/Qln6IzSl3G6
koQ4orAj17qHhtNHJHVhoYehHN3lELuCGThRpYxbovT52wnEWGiYZHlRkR535qEp
RpDpetEqjpvMGiWRnHh3lt7xPHNArqhmdLDarSGCAOsIn/M2pYELK+Xp/En1inDS
fJoK/3OkOOlCwYF+hLc4UGpfFqlb/Fp2gnl9ELXlvA8OMIU4tPaOFKdsb7fY3+Dr
UnyJvaDO4M0FHu86cx3D39Tnab2j4GdUl/lAsPSKdO5JWjypC2ZNieDLmAy8JJIB
tCp+xsiE9ZwGk3l5r4v4PaMmlBH9LkPeMre0ROVYBTdVk03a7mxbD220fO7tSUu0
AZLD1giPVOr61/RrLHUGbQ1YXdwgHHHOCKqhFBmfJEem31SmxOF5VNB8OHRlpYAx
AeQGf1gyRd3DZbMAZIcjeyomUg+RNiCzOt8YQqCTAhWqBh4W9iJNX2ju0BMhxpGt
0D1yF5hY7GKGmkD8QJdO6A+kf3LHdEfh1ObYyvEIkaRuRnfwF/WyobYFkd0Yx0u0
b7Sd88YcTO6uvMMRo7tUgN2U+jVfQZs0yv/HLa89pg5/JS97n1sqBnZG/jNA9DhM
IRBJMfSkcd8y9adqXtlo7AFGIjqSzLUk1Oevl6yWAfl+GbADQs9tMAOL+q5VPcvV
5ililzGzCzKzvYSJOWLaqUaMRCR5eiHDL+736OTtrzRFPUeNnsVosFXKf05lEvM1
0oFFq2uSuKnq1Echpvmj5k2CuGF3V0YPxF9Z7/oCbVcGEe9wgZsG1PL26VFJtVf3
O2se9b3QGOUmYNNtZqq/zdyNjGkCW8eDPDWWW9kvw3xF5xBygz9Z+ztVl70sqQHk
w35YwBhLC6qgWNuZMPwuoALFQX9RIamomiRpwVTCvnT/FekxgTYwARCf5kZpXVFe
z0j8SPkcZd/oxzQorOqTdhUzRAOI2CZ8mR3RXhmBdUEAnx6rY1MHwnMvAye1NtyB
q3+mjIg5tZ60QcKT/nRDnerPwj0VNk1Cs5sB7PrXIxO+5uWENV8ylJqVZ5wCsyxQ
eh0icQVaLAvh8uost/XEmFXDPM0nEXyW6NOEi4/gMuwJ1UY1l2bpxK443Auhci/6
IMUsal1I4W52sFTvfWBPLO0n7eMII7tSTfttN6odJ0vsmUOklMAybhjXUk3tTKhd
lFK7fdR9pchCHLzynLOR7Qt4BTidZ27Jg2sA0zhiOPiqXoZXhmAWRyX4SHfZg42u
JHsBDoFJf3JIg6bxp4VKvOVKhoCQZLX8Bdm+KKi3xc6l0a4Vp50BdpbbstCIXzr6
QuD7yG1GsoxwWVE8fygP8g5FsMttK94WjbjCD+zihnTjGiRz7H2z9nILTd0+5hLv
vlXUZ94plcjmrUNIh5b0+5buqKplqLAiW+oNo5t9sxrphin7NVRoywndWxpQcGLy
36K0P0dG1bw6RROWMBevEfrl/0Vfa8LAac1m48H+2cM1vDACNiAZUxxgmIKVb64G
3rLX9iW6AGQ2FwJP2DdpLPns6yiFww/MvwtT5LFa3hXKFKnJsQFwveTfEa9Gpqpf
IxoZCUmPVRkaPijuA1rsKwMsXiy+f71C1gP8ycmkKpEtR8mboJ9z7BDJePETk5Q/
CdI/CIZXtHG3jaIzSQKI6t8M/Z/kE3GJcj3AykGZZI4EcHEJMLNXUC/Q6tx7pRud
m58KN0v+8Hg1xHC2L7TAXSS3ipk/iL98g0QzVQQwRctrwGcjozFfjTuhGK57s9Bq
ptJ3+0E06v4aR3EdrfACNQl9nRzta7tsNEXusXJBP0ad3OciV+fktmmPj2ozWpiI
blcgbEty5hqdvt+Xk+/80FrUwl0dqtFBast4hilzDWC4aMEL/9fiXAA3kIevedga
tjVuzOYDhj3qheVlEdXQDzuBM5XvfCZ29MlDWsuzkj0kxYITbro2yMQh6liAsrQp
VKHrN1YIVFZnYldhRyBvQpkIaMOA4JGMMz0G/w+u3YXk3MnTra8FM3qKBwLdVWGs
q7zlBZSy1rEOtKz5+oqMC2hlGnjzOBJdhSeRhFgz7ndymrXv9+6MulH318h4CDeb
62gqJLhjXsxl6OoxuyD5n8QBvdwYzPwq/JrgaMAyIW8cH9YBo5sCOHS4ERmpuyIY
AlyiGwVGeXLFZ4NL8ETXHnHZJqYtEkBaIo7gkrVfAi3dPhemqcxgPABhBLbiqkXB
DrJ9NgfCh+tJarILRcPr9lGIzs1+3LD+GVj4Qos1Lw4lIsnDxoiQWcuyn3w4jcuc
eLzkA13mLIjUv4OFnJcDxPy1p6Ig+KidFmLN6FwEi7+jdLbDSIo7/Qgt0MpqK+pD
fnmJlDVRVwwHJfDwlF66nBG487ZzQHyYG0/M0QlFtjDdB+ZwxejkZgXNhQXFEj0g
rR2TKxUBcu/aU4hBB1reasZ78jO4SGhdCrTI8Gm/4f2i2k1UDI17HBzQomCXYVM6
qlzOZ3Cj2bOVCHQeuaqw9GYkl0OgYvOhhtnScK4ov/plTRzfsRx4SVEQhiSQ5z4L
WfP+j2SDy+2CWMc1wPVynE1VkxDqTfn3EuqttZq1J8rOU1b+qya2rCySct5k3RIk
TwQnHmDl5H4mgrzVDbyTIVlLfN90joq+0z0nVa3lgDQoKtHHFpXhKuQTtt9EdwwC
vvaRrJHPR4x5eIOvl6TgU7AD++eneMtYDhpK8aER2I6jsh8wGG1gzqnNRNFI5Ggt
Jpp3iNwWBQy/ZgSeNloFkxCgiUPtP4S4VNxOM1HhKEx3HQ3th+Bd57S4sfHWNhQV
qoE2Lgytjpu8n1E68GiEu3kyP5XT9TEevdaQ3N30Z1aZYedRUwhLMcWuFrYOqVRh
ZJXbTP/wHZclHmDr7y1zqwjL87vtJra2g+GTHzB3czFp4U9xSl6wkPEbIiK4zfOR
13SFD2bOBR3YHdacP9ZsyrJcu6Q7L2gGVcK7d23ACQbDLTxdXVJAIrpOcEYtpO4p
SKskiJjjB70DXf3N6zDI1VJ/nPH8oncbAksN9n7S9FlKRxKs6GDMLTnmArzh4qCi
N6kKPDlxSa05nkHY9x7UbdWv/tldLKf/eeFhAXh5uN1u9qH+YIMmxWjilpQ2tkxe
Q7ZkwZ+3kz9cQi9NcIrvBMHBACSKhKT/c8SvWNQOuzeion4Y5vyP3m2LNJWnJiRA
2FEqlZcivtqpXzrHY6uB+VMuk3ThoXLKGGbo+eo8aHI1b7n8KZecoCKwBqTLg/OT
2loEswsHf3H5i2HeX4U+3C+R8eDm8Ag2+vNgJMX06lnjdoeZrrDLbnRNfQ8yQqAS
bLMR7QnoNnUWtm2ZJEACKQ1hXo9rYoIROiprjQ78JlbnG2VEdPZYul26Z/0mv5Iv
occCmMm6OEw/1jmqdIRP8moA1KEXwm+LFXsy6GImR7s0OoRZQlC7rik0ztx+I7YH
uuNzKxPUA0wfw8zPVNdd220DRsA4C18Cqtg7/MaC8DCbaqMXpJB5XY4bKaV+vTig
4mDLbyv2Cf86jEsizqtQ0YZhZwbYZu1aMo6tM/XKiGz4iS1NsqIcb5CAoNadWo+3
eOwEoKe0DMVYDjzJqWShaciyJxlJ7g1+Wo5NDL2HWQbLCZpsqW7pN0yUSM93o+nb
kqEufu91KD64hJVXc6ZQyW6FKO1QW5+a5zTwiodiz2q8CfgCVHyd8uH150F506TC
IjzRX4Z0o0xnq5mfp0ZuXjpKGja84BWIEO5jRcwqSTMgbbKlGoTyH7S0ZviQUfnj
oWQP6bN0TgeYsvO/3BLeDHsnUXmCEIif46uxPDgMzomb++RUISq6euN2lBwhQOZu
dTH6q7u4A0ZglFHEHW6lVetmYeCbuiayDeyDpF/MccBgLEKJLvCcUrhpVlkjyjFI
aVn7vqcZjCQcZP3f4NoH3kZJ30ZNjk8BWXanwrfWjszI3zzjd8gXkVcpk7yB1mff
RJ0izvMMHCPLSmHqFqflwsQaFJ6ndn1KzFqE4bcKr5Mc8PxjrBCbWWV0tqhXaewz
5fRLr8qKzeieFjDAW/LZoG41S/G2b2OQj2CAHou6aDGy1jsWQfo0C7RYz/k/SlFh
1gcai8dlnXOFRCQc5G0gNOKZ6rT04scsHgxxYV4op6b1GdnqNCC0pZIFrO/tdT/n
4fT6PyQKA4rLjLhAEHvQIdiRcRxCSptpiqC8O9dF9KYZ62Ad6cCFFQIWGTENNKj2
CUsTOvy9v0ryS2qcW1a9ZRfe+4pqChMM/Xc1a7eMcLlpUc50gUJqY8OOHHUJC/2V
kwBE0OucguTwuzgDWBjS4mkW2H3ek/Gu+rJYm4ZCMetEc82fuXXTR9jCfY7IMa+k
9MXHRjI3oLqDX7cqf9dCtXnu86Ggk8Tc8JXbadWqaodk96nhijNlQEhUeEiysD8p
QSIXGTK056RCI05Rhqttgq0ou0XT7Bl2Rg/5ktXvPBerj4K+0ONNYFsKQm46/KCX
CrgEe2cOTLe/FdzfPpbFuA6V9+5tFUVKxiSy15aGyBbAQ1ZqTMcdoBMRwWPpODNK
iW5fTGdkrxnAvf3orv9TTsibZdDsU34s0WIhKuDgs/WJzJssMudvAP5FlcDo8PbZ
NAVZtuMsnx7ocgQgAmWSgwJa08hB/6gHoTlnY4QeaPL7uipfXZm/hdwEU3Ti9Snv
X39wm6OKvVNwsMc8+DLQhagcHLpn+KKA4ubMd3xMNaV244+jxvENRnneGAOJlk9s
qhhpMzXO7YaI3YpuTdU7MSzFS+RwADt9aN43CCHKKdibpmhTZnbI2bVYcW7Gh56p
klUzJBalJgyBtwHCCiPLCH5oCGEzqyUSy7Y5P8dckyyubCuWO0YwtrjujJNvPZq0
xxLM+LAsyRva42S87I4AGKnuzuxd+Zp5wOCbEuMWdr5TOYjOYslWnXTP2OCFjS3a
7KG6QxeUAHBHWeevs2Zza/oeVLeez4vuSJRXRc49kuct55pPhVRuhi88Wcz4/YOe
mzkj7ETIigBhsQX6tJAzzo8x4zugCn2QtFDHvUg2ttaU5Nto2cz6KAs27y37gTT0
TxPUQFK419hyvHuk5eGLcBM/1En4KS9pY4Wk1SWDd7I9NNAnsOesiENWiynfIagY
yVVAgfA2GGmdnxL8XB8Wi4Y2zlV8vy/AJit+G74WIlG12fpF/S2NS62AZ24SMpnZ
syl7BO9DYQHakN5WQUaTDGXmGbZZygoDDocwzNfe6mM9gREvUDMt75A+vAujBYCu
6xSHihZFPcbEWxQ8uroTznSTemMjaOMJo/HhL6fLcILTndSUdmQA083bnZI3YlFB
brQIipffXXrAQd200nfNAeQtuXRDyg4pzKMBtgjKnbA40W7WK+rnXh5O8ymLHg/Q
cMo3b0Ge0i787UyGSFKUtwmlNFrBjmL66Q/xHsBp0EThDm1D88VSKoGKToMM3SBy
pjEPNiBvuf0Y10Vr6y8UpgjcR/u97IdB3kLQVll8LWzSb0oYmWSsaTa6dSALMi6n
tcL0PQdvqD1u70pdJzzlw04QGArNz4+2f4pV94wlec3woStr2RhwuszzFuqBGKKh
W6ZkaJWlzFmR9TTjGxx8inU8WHfm6AKMfzRA8G3CmdO/F72GHCEqIPgCU/sxunJi
7OVwnUoggtu7XLXf1HfWuHdKg5TP0nvuzBKaku0iTWVz7gTR2SUoV6/OWP7kuCbw
/G2csuEgr///ya/CH4eI8lNEpQaU3+WjHd/vmmFAnq4CKO8WPaF76f2JcRV4VF5G
5ycupL5KfgYOowveQuqEsNnAuS8uNfvH+r1TzoIgetgU6Mlf4rRQ20fz6nepQ0F+
+FR4PiuXVNNb5jRxwplCTHeDnnU87rcH/Kaysx90SuRP9TcWT8RX8ziZfM9fp2n1
yP+Wz/0NvaF1yGuPsa6CHA/rf6Q7K4P1h/bG32vk9BtxPvbWBTCKGwujmXNe7r33
RXzj2HG9YziUbnhr2XirQ5OyWZ1YX6FLpThsruz3GEYQcANnp00XKoDMnVIHQeAP
VoFDm/oHCXiLrj9CxbGHArJy5UllSQU6U/UxGbB+FiQNQH6+buV3j+EDSXZZmbm1
BzgxdbUTPJ3raL2I8qFWMKm0MzllN4B4KGlyAXDoeBH1mS6or7nH5MoRGGGhcx8h
x10W8631+JqfxERp503kYDz2FYd5X8K91eD85zHxmTfaNjsTHMqJVbIyDEnyEUlu
e9ZXjf4CgNiNC5WauqDHEqRUqfZjzZFVyiG5qPxIQxgX7rICXWCqTKSTTP2XILF5
5pgNK745IOTPDBulfg8t6TcvHinLHx2KT2+htalqI5NldIjzej/bUkvorFh9dTJ/
fPbZ8csQDvJfZwH0NElGEUlOZ1dAC5PWXRE10MqjuDls9a1/SlpxABoXUL7ciNKX
02dzyKZPpyv5jRKrivldiEFhm6ofmY+VvEO7BQtsnIk9IbG8XQ1ADFTzm+IOS5St
zsKCWXVoTJN525bOp7iQERYZVrY/E30l4+RZqwcNABZzmlSyfZ2kaLou6/WmhAP9
SH57nxqsJvUunJKzmpV+gB7QZmcUj1hr7BylqNU1Yh6Wsh7XKO5/M+dayQfeMDmZ
UZ/yT8cBybAdX/ec4ALpqDhVONBvH1MxeVLAR5zMpW4Z8quG+4hMgSZbUd638Mbr
DuUjP1bqLNgd97ylTOws3IWQm1ujARX356ii4NJU9F2WgJIo2hJfh1zFo9qXpO7H
abp2skbbX2NSZF3YOuHRRSh0Wd2AeeLfan+GRH6Fz5/5fHo0v6pT84+DCQ/drBZI
H/kOrgx0xNLvspKBcU6jApYYjDpMfxjUDuytGT4Gwwgyuuz7q/pJVuJBb0uQcSst
hw67rdjcDHiio81iO01/OLXE2I51Oie2RL6UpvZv7z6cpMfxLB2IQWjisD6KgBL/
aU5VawtS3+baIRtYiWjKzs4yD9LMgvxKkVACpIitXkhgRjJhX5sivHvS2Gr2grgc
qT3HE/JNWTJMXZxC99hLNKQkWf8RUbtjGI8LXqHnVXbbg7ucA/CM8W7GvbVCL2eX
moQVjJHnoMgCNzuRwcqK4mac34mFAYGDTY7rmfS9RIm31D9HQBEXNnZfo50hwicw
IQZP9Aqiad7R+yzT2/hQvs5btJP/jhDlkYh6UyigI5pryB9LGc2qN+mQUeG3pcq3
Cz+xz3SdXDxn4pg205o1VGxGzba7DiWDZ5juDUeq81mKqgCoG8iHacjTpaYohEYa
YwbWwZo1WVWPSpumYTZRW7W3/D+ZoOvupFMeaF1AO5hNMJs4ljc+DZ7Kj6E7fU/O
ylBnF6jjKTsbSCjbI2YKUtJSN97kAs4sDzvQqU6PKzrKUhCLXE2D+Fi+bG52gyRF
76GUwWFBx3GGgCKVixpFnQmZtqH1/V+c3YXqtXvsKnemtwE2dwAcDEv3ngXkvLA2
M6JckIt6nVywKYNQ7AC+NzB/eQ+jIvD++j3cgyRuh7mQslCBF4Da1+eryjHV4g7e
Z2xyvqyL4UgoH5KW9RlK0PdUmQL9YX1UGdAgDw4StvGVoQtBSQnZnOyLUR/LnPOW
S9/Pp2Jm16bb4QdA+hxTVI5Vgg8PKfWU4Nm68mePfHLklcUCAc9hH0mJ70dyImTJ
3xHrThl1a8bPgKWBE1IE3NhoYfagoBhI2aQh0UjP1Cq2d2CGaKRb+Rk5jfc6pf2J
h3bWVA7EQqX4ijvtoagmvx2WXjdkuUw59hRxQKCOJfTSucQZ9L6/ejKO3SlIF40a
tq2akWqcxavibL9lIsHDdX+JkKB9PwKBd1mKQ9FkFaJ+qR+h+EkkdQHHbLF1D4I3
Sdx4sCLS9pCxgP5zCZtZx3Rqa0WKfZWq3uiypy6bXATAIxrSvMXPTh2QYvBtNKx8
MEYq79Ugy/0Tet58meMObpp3S9rp5G66JVEUyAU6PFjO6GZvBD1Xp86Yi0AlMEmG
Cndtkj9my76cYlzQ7FB97DGoL9Mpn6yOJY+5vOb1SV2pNjOOpapOtBgJkMjPtOs0
RyRbleVhrpFzee7ikaaN21doMSEiB6mEyVL3UeWk+jyQvlBRZUF31uncUe8u1aL2
d2vMzVTGQWmqmfcNdqqo85q/s9Wa3EpoPZucjso0hG/tK89ReQFrqzTvvII15O3P
6eI7rM+voO6P8NZ3WdnYXz/8njG7TVJGyESNnT5zaxEcbDaZoI62pSPTf6lTdrCQ
NK5qtP+6Fo/+cuAjxgFhrOGSPh6up1d82MT4aNzOxMzzTi7pHxxgVTQuVrYqWY/+
2pLMD2zppmtcQkPI3qD7JeZsrik0FT1bV9kkUc+Q1HJSpoMvCYwRDibIJNteigKz
sxkUdpaI8oeDn+ssT70UprCGoSXUlHRQblCfuHLRvYCTtmZq4E6RU4c3gmYELF9l
FLTrukMIdB0m94kuIINmT6aSBfwxOklvABbZ+pz7Qdx/Qu0f8j4Oyn3kIDNqMIMV
vC90/iFcJ3DcyevnPEPVmnEQsjMIymi0lB8qmpKu16X9kZEKl/Z3QdarrDxXu0d6
1ai++G9LGXV2v+c7IHqwDo+iEOH8YpqRzJPxFUHqX0Su231fDIquNTiHiYgnbRhC
I7XyyT5QFkHhVid1KWAmhYBtDj2h35jsBJLyDwLl00itIgclH0IALa2VT9Zdz/IE
mlyleNxz4G+cq3JhsK3LYexsMegvvRaepGWdSR4TIS5XDNlsNo3+tuXTUKk4LWHz
vdRDUoyQWG1ShSyVIoNaXrPdnaCjzCuYc+iGqF1vdHWQs9XZrOC3dRk7guQyB8sg
axSMta6/EmN/vHaXbfh0HhHFWz6AqMqVGTLit4qXObCJn4hAcfuDta8RHTRInSoV
71Ik3EhIRNt2t+KlDnRiFry4owdst1enGI9Va5GRqxCmKbHmwUmSzwsu3m4qcUa1
2ixFFtUoDkTG16d2hy/4e337RyiwF5q3ytT3m5LsxiP7GPqTS7SOfO8DXpRltNmY
3zudzgnZGSEJDUFEtnp+spAYM7eMU+DRGdFvhOws8rTlDloQuew41fy22togzdnP
CAAXaI0zWBwNJVLWHmusU4mn5+ILmPavSG5rlUD66wzClNQiFNvXBSMETYJowWOv
gAXfLU7KIietigroeNWSHDjSmzlKqpiyly42jSvuiWmnx0dtKrlOQxrknQCUNnXa
xnDuK9JZHUdJeKcCA7pIC46uFBMr8AdEcgm0rvUAJuaH5D9Zd+5UdV3K+o1DGKWV
MBZq9pd+PEkoXxWOR2GSw6OechkB8esdad0ssjtLhRAp1sIEIpQ3s/y6zdJdqJHz
vlft/ghICVTEVGXL9YsFZwhCl+CNJPa/nlyzer/gmGZGlZUj4kATuDvlCIQVr2kB
xhvGVIH6Nw0FDqnAUF+L/gQU5FoY4zzD5LidKnXGOnwQpA0eoC7R1ydk1xVnwpDj
gMvHf230ziMc9KtzVOHFJAbE+SQPsCvdhyTxUit07/o4AjrHQ0X3g0rnTmfY9Vmn
a+E0T4Jl/4pZwPq9TknmLDREPp0nAVLd7C+kJxgmoJiWDd73ZSoPeivn3B4sdr2U
vINzgtGbZdNUQLEEg/zYJ5krGYPDTMVswFKGGu+Z0G7OVXx9pH41THvrJyJEdKMI
uImmWe8dWeOpHHLhC7seOYwW/XojCH/kBw1cVizKer9p6701S5jqQ/GQl7aF0T6r
aM5LiRAkKXvJ4lRxBS7FzdgRSlW3hWS7o4f2I/iYXi+NOHHHIDzipFUxarOF8Pvw
18w7KFSy4HzBpBR/tT/UlzzX0cnOOtNN7JZ8Ij5a0QoeHo1lkH+LexziFJhWAapC
GeC5TOLrJHu+yJ4Q5zF2QcnfkQGPboPxxiJ0BZu28UMPc+lRTwdnzzgL+UWHzZlG
SNEKJbgmJpdjUkTldmn7g63RJzmojLKvBxcbYAi7ztBmofQrJ5hWVsS09K9hVN+x
vmfUW2+cFsc3xfqHi56KFKHQS6ob/c/powXMk4pjHlnBJilMowLAOidLOTlGU6kB
CO30b7C/HfKUyRFrADrgW7cUL/Wn1PzyfMZUcoNla1AT4ekoAhFe4wEyNVvL1jw0
h4oVL5jQphpVfOsZuo8e4OOFsAZhLtb9G/k3Px3GcJr0fK1iAVGPegDOwh3/L1Un
u7Bd6bOfhFlfeL84yuP2v3ikPzQrZlZy3FtCUlHBSH8dp02RO9PhqL5yId5t9GiF
tdbBoQrMX8bIgO7VhlB2dz0WYFwAjxMWwodT0hye/92gFTB0TwVQval6xcKHAJdc
fH68d3Y+aatGENVG3Yv7xiVDPQTChF/+yTnKfVKXB8G7lUjeU3NSezL/fpdJcD1L
cdzsRTxx8q0saAZhDpvB2AAuySanIvIFXVyidKU57n9Aup0G1VjtlhkGM0ukqcOc
oOmLshiBQjL65hIuXnQ9E7FwBmJ2zTMjc1xf4qirIS1dd4KiaQFfZ+uPMCXe4Xkh
q8L6js88qGbDQtnXy3QAH3WMnmLpV7wJjAq8YHXy95yHKqQqgLIFrM1XvLzlqVZm
4g/tKSuarditDyusfzsAjcyUyTQZxxpk3tRvKDRCHN07F3y9DdDd24F66M0OOt4t
RGlaZY5v0Yqu6RL5qIhiWyMNeBBR9QAPb4kVkI0rSLWNKrfNevJ/NKK/WNdiByuu
N0F86VE/BIozczFUM0BxnjJe75MBZz7W2hzEYbLvif7LgENmJBWeQglxYOCgytJV
LEXWNKPcT274Lswy9C7snMrJBcZ1OJdJwDnuunhmBIV76jWI188oGHYzrkt67sac
rXSdd8H3/uOxux2N17FF/CK49iFmMWaRnCwATj2qM0y0bxyHYBLwpfu9IfWUXVvM
CfsdSIX6h40+I9CMg9MfMy5LFauygxfCeUvxkIqxgdUcAMo9o7THKyIyT9715Ad6
LxfgwDWhaNAEvQeja3XdvuXCaG0e3d+e4S0dBCIIeqZOrSmyImGpZLNMO1LecMSY
Zj36IpzbhDTbhNFgqqfpoieTMC7rdvQCy3VAxiSjTZ4ugIqcf2/VTAhdM6CI7U58
6Zv9TVFF4agiYWxL4ZoHXU0R5sjJqB3IC/S66Vd4BDAfOZhElByyUw733NuWqbNZ
86p8anikn8+SfWhMFT2PNCXnhL4jqRpe8EPmElfMSA25+i3DTpkEf5Vl8yWgp3PQ
lj6qnncL6Dgr5z9UK6Gjoaf3lq8w8LZSU9pFu7nzsHaK+/gohTkQlnpuidql3ZUP
WH/094B91kLLqLypQMVQ+GkbzQHhMRM7Rw9gZTe784vCV2X0NnfpK81VGdtqf++v
Yi5RjWa5Rb3sgRZDQWboT3FX/xtxdlFxZqvc9YXrU5yTpvp6z0TxoXXSMZzq01o7
v73A+NgppM70bJQrjBVCa3mywbm2BsKl5on9PcMvtyG2djPI9re1MUrKUCtF+hwE
ln3tc9dvIqrJQbeHHX8OxJ4Fdp1AOi2wOulz4zWy5frPLVg7DZMoWb4cIhAWu9qj
KPNyC08i3hVXratw6hlM39jBkra81zCsVFNqJmCvEcNEtQYTyCy28rPdB4l6KU+p
nALgo1HDJGc41C60FyIhXmykUdv34kxp72X21x8sePyy3u7R3OJoK/vAUanNK6Ln
MVHUEtega6XnEkPt+PmvY5YCN2JuBwaj24/87HQ3KAFGluXWeZIMYT0pQzQCVs4w
QD4v81+5MuEt9HXy6jO/nOslYJ1tPNu4KwQ1g6i8qOe2VMcHfHTx9FAO8DHc9XAU
dMvpvB1Us/SaK2LsDhqDrKjwHQs7ZNUvPtLxur7KJeR9h6H4a3AlvupO2Q+gjB3C
wKvmfaIdn/iM9OT+9neFlyJSpNedrwbOr/Dn09DKOQzgmzDrxIqp2Ujv2vUj56i/
hGzq2N9RVP2ANV4jw6TlIffY6x6Eyt846cHvAIz+i2udpOxpL3MHN9gI0VHjkid5
hMOjtijngwsddNoJ1mtciQM89PJLvfsTFFWSl5cSuUfVCZRwpPGrXGkWUVkapaqL
OF3SSnL0afAyb2punJez84hLq+Ep5AX7auYCCPKUvHAn26T1eSsuaHksDrRQ/l5L
RoumQI/nRjgttLzCHK1YxTWlFclhzlGarmtV74GTozxXVF+6V6c7Ck9zmKHTsw2I
bkp9a5VK21zHAeF7Rigck7aBU8n2o+ZQM4Jr7uwGvH2W/ZaY86rA46WUoXJkH28a
X0xZ/XLmHdNV7nWID01b3dKpsv2rS3dzdoOYNYpLExtHZnQhSGyYU9+bdntcDRqB
x2AMAYg9/D4y3zHuZB1jCnq9bZgtsLUu1wrbX/RDfmC+1mxUYzYDzPdgLxlg5+/C
YQYudhHIundOBkrfscZQUH23Hs1GrfHFlCk/aieRhesSBpBUu5KSjEwsCaoPnEoH
nBkx3+qz/ZP2LNkuSL8ubUr39nXaiOQpQX8bPi5PzbEhIYu0WCwd3lw69MmArhEg
EJK59IWl6LOpPqKHc8X0+iODLt6+kEgX6C4lq1kBnqIAIptVspL3KysF3zxUS8iB
ySJafOLW3XIxOdoC5z61dzq+Nlfb17aUR9Zc/pJyYsF+C0WRyPP7Q+eEAH+BDPZB
IPnkIk37HoqAjjy6lpSfPHMJ5hGuokoEN7iqWHOv8e9w7J5x3+lqQc06bfVJezEr
/q1+5KMba3YTeElKLIBsoV0UUVTlcZ5eO1KVW2ojhzxwtr+9d65BOfSzePDqmYSk
WnII6wSvT/3v5uc91TWAnGYwkRM34IKLMQs2dY/RBjq8QQ++x+cEt1+XNm51oNd+
Ebo3fRbDCD5OMqOKVqI7e8wtJNxSUG+yAafdeZW5qWKI6696y5TR+0p0/2yeMsG7
AIiwKb1TeyGDGnGxxHVTCcvHvU+cVVIZfcvbY5/Y4/ghQQ84UdnPMTol0J6xKy43
Dn1GUvx41CZhZEr22Rx3olEiA7ZhI5x3LlX3PsZdo3daW2wh2s0CP6tAA04KeC/j
qGjFqglF3sJMRL+7ez6+2JrB3itVUpbT3jt21B23GV1Ga5q8nq5oECnvGKaQm7M3
G+SswSYnMzXLqXhZUPrF9OTBda4STITcDiDkMOXkV2vrBuHSAdLNNCGF7SIzpF8G
ldh8L8gh/RY9qo7Pr/n5+jJIqHhDsdJjmawj78mw3RfHx3Sx2jbkoQKCFAcuvnPf
hkS95kDhzDcxi1qneOa8kSNV8rtouKllLEwgblt56xYYJPYv293uP/U9+atck6h4
8J7WMAniUHin+74cc0xxoR/xBp1HUkiRwXSj4fvHLOrvlJGLVKRUk2efnRgjgcqB
0aQsdgdjHRnubauamZrBv0Cpe7P5q2UUKfxMU/VdK250SpWsYcMfBIMnz5mtogpF
vITe3/cujm948mgAAb2TzF+C4nsqMEMOPvmCI13OwETn9V6len/kVoBCaV8DpVvb
448DncqiXDGrgN36J/v8hyuvFnjDMctlCnZSHXxh4/9p94GzpLDoA7OWhSih/085
2tKmu3AycF4tUIh4GbmUYArTLPGhqwgMUUKjodgMLalTHIbou7T1a6x52QUb3fUZ
fxBK0kLFRzx4CgYPTjqhJ4ZgyBpb30WmK/tcggTahak15LXRDPVqEfq0V0MoTSBT
XjeKV407UQHUjq0h4NH/bRSJqGgkoyEwEg2deEjjYCkePD7UWafio6xRgHslRwTD
XnFB3wwcxsWM2PjDdh90PiLZP0Lq9vP2laLeNUP/VSPKOpy9y48ZTwzrL6aAqlnR
l/Gio/zVRlFU4gIbrFUzQZejPf72wvzZpW3WfD3MLXBl45Z3DGpZHHm8kTeocz4W
2bps2wBA8qig9bCX0hWaCQJXz2rNfE25fffHU1dobbeuRGcThyQ6saHKGk+2jIQF
jU7zVeIzZT6CsjR5DVPxT1L57KyebUVVzQbOPQ2lohRYpJsI3pVGXY/08LQmjZQi
cisyGcktyO6vnE3Mgt9fTK/g+2zhV4JZ2MKo6bvjxpvon7vf/qdvaMzllxKNQEIb
JM09+pzzpXNixGWGOb0Au23pQSC7GKygVVqZ6+orDVGXzZahcqhGUgsSiQsTRz73
/C7UJJQKy7f8Z8cWihANGnAzGICgnTg8ck+PEGX+QHxqi9lkV716jF2lUbEWWFYX
B7keHU5nuu/j9LwIjnIofKjqjUlwfeNMNta9SLfQ4fenRuv4jIQEFw3NhtyUSFYb
GbxJzxe1It+pGRKaZzJdhUD7aDfGpbE0ULzlKvttUHkHnAohg7bPcbQGgXfXQGdB
z+PDbb0lRSmo2RqKR4O94lV0bg4dEq5oNhgQ7qKa3P73rK92g3D3ygwEzjQhiWzF
R2IbTow5KEmWsUjyouv/FBR6sBuuwtletxgK0QB6uXbd6Qq7E+9yVhWu9Ht+IOgv
bUAnb0/38k+gTs6qbvk+kzUiqFZx3Dl/tTTtruDD573HbiE4JbCZehVHN6+KpDs0
TnzNaD4gGnV7RxtSPvteQDgT9SuUp5jF/Ummk0PwwjXocRSlOPCCsgM9S5E2qpCK
C3mMROMCRhFxjJXYk1aXPMaAK08g6A0CgPtedv28R8NNUo8+gAKv89qocwfht3PZ
2fh45lD+LOg9HWDnGXJMmCxcalY6HxxnT27xEm0eJ5qKEKAWAXZ4FSTFwMg036q/
TvXaNdC5IwQhACYpEKCX4HszPJ9cZUoxshtGGEisJ0C2aq6QOHAtIoXDL0aJN+VX
0v8eCMq86f9ciJEpesG+zdT68TowmJ53e1ZuqssfYdKcfswQ+bELjwHE3xGNW1nS
/URQd/qVdsYXEpMlo7f7/+2ie7mjQKkwR4bedUcC8u9JR8G9vlFw6aEaodViNEsd
F56DXJhvdJLGTxP8T7ikM7AIUYLWZ4PDNZPQfgfGlMXyqbjIE4niiFXCGmpKY9D2
fimIhtEegneNOj9vrOufbbMb3/mUdymtYxyv33zMqYrU87x4UAEOoNx9G8DatwaT
rMi2rKMRxnI4qVxsIDw7V+EjcboY2nOD+yhm0THUlJ3SKwqbXKcn4i8cYPuu0mqE
hLSN0lae1GqnAEPhxFEcT0dDkfFEIbt9UpQ81tZkff5dwzW7zjO8JBgBsKJa9qsN
o2MaKJ/SRzPN18QtNz4LlqqBLbarjFG8xUFElRrXSA4KZ9NZ5URGJn5WE0xiJdk4
EAY5ncxTE5+Kd2PsV+HJ6Qga/ytlM09tQPAMGIZmNJfsPLdckNr0MQC593iN1d/u
6ODn1la5gm9NtvhFp3P0qU90IwPijmfClGewCtzcPcrdZm+wLl8uEtGseJHHTCae
x2cHyRmR5RJWlHE2ll9h1efx0JD0L5y6ikzkQC9BBb9OOc/E8I50GKoEm3u3FvGj
u25qbCimggcDRjXoeiVoOejSCRA8fwNp00hXXILh2AYCqkBUQ5bHoitBEh9UgEoE
xI9lLmjnGKySZqx3xpkNEa+WKntKvhn38Bp1KXIFsJ3yd32+mmJnxoCkPyx/GpmF
iTljeTav/nlpBzljS2fMprzHP201uxswDYPHYd2RT6qYXA830uir2zmqDTdEuC8m
Q+hu63S9wClWywHWf3zbCTFQfffwboE1ICjOO33cCreBevfesiWi8TMIoC4VZU9D
muF98Fwnfwt2OR+NXK7p0cVjrDMPiGX5Ckmig1yBkz+FqRp8HPKzXQBrT6M/YTtz
xWVQYMWzT7aD8NbjKWzIJ8xJ5HKcHAIPi6pqi/lso1kOVb1oMna/JLUQENXih8iP
ZZtYjLn7aGSnQJ9Ymsp0TACBG2Oyko36CSWp5LvDwhRFg14AGGoi5PiJm3jWn+DW
baeyUcg5mxKY3CDogHL1jsPHc/S9uSmRsQpcqX1MxhbX0ZFsErFfOXr1ntVe7B6m
sL30zzCNH8+H+K7uJMr8kLGrMAAjeDhi8kpwB74M5pBgx4zwu3N3kFdsyUIR4FG3
XkZMVG/9OJ5biKoqOy0iLXj0F1QvIKVuwlY8/dLY214KKO83rbl887bF2mze0cLi
+0HOjKR43+n45k8floIgtTWQNccZyRpwi0g0EYikvF68XRtivFbGWYe3RMkB8alj
YPZQL5yuv+zvsPc+dcD1FRTqwd9dh/RD2BvWt5apiBVa6xk7pfyEjxHf8Sa4ZrHC
eK7q5KnCxtV5adiiqsaiFY0mBKz8hxQDktDPOcgD2ycVwX2H7m7/GKdufY0/tWTl
fMXDqSmQs6csdaa13Ni1LWq6iMl4mMvr65PVAaHNJ2P9rV/5TJtHG101ZHxWT0JN
WDYvO75hqvGpts/KOrBY+4ibe2j1kkdgtbOcjSJqRX0+ETjn+dka0ifmhzDE3YfO
vSOEXsyktY10rjyv7ka7WO8/WLr1hKvSOJMTeSrOPZIjHhJK8SOGDH51AchFA258
SZfWjPA92P9ybqCW5h/pnDLqUlGcREZoUUd7PEZAOw0RYlRubz54KLB1n+g6q9HM
KuMWOTUDtFwLqWXW1nvqbSBPebo20VAZfg3QEItoqY1zetYCVliUBldB1F7NEW3s
AVUQqSm0UZg8IP9DZ2rJ1rpvWopcXNIi0sRYfoMQKrlFL5Dy5Y6Eaiho4EkOogP2
hfihJpt9iHpm0qwfRwmcoeIklO0MyLir6FVEkMe/b4TMl+tKkC2ArbuPZjIWiiVO
u75kb2CicjQ9l9rdgxH841LXg9ZdLXDS0Mqk/XYztAMFF6moK+XN3uqWjMJAO+wy
bJHeh8bCT6GP9EUhre7pWLAdtSVWnfP/IOhCq1UxAukd6aTR+nVcoZ/PqiCj8w2F
1AU5y90YTqq5KKpzHO9S2+LAHxsal0Bi98HsfOORYVl0V6TefvY946ARGssUUy/W
KImdLu7O3Jk6djZObpO1m6AMDC5WFemeIX8iQAAn6vmxHVZWMNknCo1guSFQE5Yn
OFj5HrMwYeXVtimVdlIZmSRqcK7rNUCCCUhZXJi8c4hkAdzpqrJsDO8BCRztyZ/z
UI73Ev1ZnjJ9IppMB4Bngj5Cnf0Hd6bbk00Ogg3MlkO/RkQRXeREcvpC6VXFqlMQ
P86x+0RXFQWBbXroYqAsAs6y9w5l6dVsY57QxUW6zDxaaRVCE7lC9gnlah6unZMw
KNLUQ6In8bJx4nN2W4f3/BmvDc7DuatHQwTZaL7ToThgypVPqRmZdV6kcR260Xo3
FLcbceJWqso/4Gomw4HH0jqUIocReHaDGLTlg90+lWPOPbF0TaSyGYnyTFX7w9Mr
vm07aKEff3ImsN92o9Dj/Umw6quS6jQ2J/2O97cC/gHZlkql/ixslOqWO7F8cHY4
owz4LDzU3k/N5W843qwqSJwKNZw8mHW+V5fL6GV1PTYnV233lJ/e1PZ8kBi1oujn
PrevqQWq0gxYM8705wyoH1CPysh+trTNbYDO9ERNOapYvoACfqikBkqsrhvXv/u8
khmNk7/wcmWmrIPA4+e/wIGjTzJ/uOc7OlcMOsdbjJEWdkh3dMM4uAN7VVqnsqXq
Q60dWoVgHOREx43tmZj8cmVqzAegkp9xiqcTRzAdGGEd6OvPzkd1QQ2F02yZkjva
b69l4W1Ok5qK+A9J9KMxg9j1ANOb/ntSAJpMMw9RLaOnhRV6SUSq4WmuTyYgrazM
Gl+007kelyuXh8ZRtRj3VoycHSVjrXibNLwK6Fm3f+CHd9MsL++T+eRKUaU2MT8W
LsH3u3w/LON1DXFbEi2u9MB/hF5+8VrbnFNhA9khbAWNUe7SQ1CZXukIeStaitQE
NnyAXoCVUir9hPjFIAdYNlsH1QXhmId6K6rlnxbtRgsD8BLYHX0lUbaHIhKpmSUq
WXPezOGGN17e3ZOFV5PTSUHdtqP82SQgvLocHLMVdAx1oMx74f9D4BN9gtJY5sdz
+uTEEhFuttsqjx3MzEasfAePrcxLOmU+oAYGfkE6e2kVX022JqreFqdPvaZiQ+35
LytIghzOQarcAJBKUPUbkQDCId/QOE2ojRvBGJDRBocu9CdKfwFGctq1hF/E+kEf
5M7d5GL/kxsuZq8Psu1PdBTjfVcbti2dyxwqGwh2eEIDTAv/BNLxwfWJ7BM1Cm/y
OHhmetdveP12EyPMWsFbrUWHK/nW69+wODuqiTEGjyfq/LGKuWYTM9zU+Twu7f/Z
t+nK0hFAvDjJNyRaymCkoPfEiNroiu+Vn7gmA/V4DJJtttQGiEo5VWw8DP+yZBJa
Oa/J5GqTrPV7hlCdzOAJ2wYmYtNg/kblZbiRNtosFa0zik2R0DQ2+91Meh0K/lUL
SH7Sa9Rj5p62GEamTaou/qe/uoMYns+2ig+tx1Takt2IK1PtnWllOWfs9zwwOVhb
1JhkrCJQbUzfvuMcA0Iz4EdlFCuCJ6IYoFbFaumx/B93E3ayzCCKSVHJGI4l641r
SxPF6t5dosujg/qJsf7GnieovWxZ27nLjSIsQLY37/zt47h/rRM08+n0UBgzfQ1o
n5tYbPYP5dSO2trVuE2QII/Kp+FyjbDQ+2Hy0AQHYdAvGZjGUS7YV7uG5o4XMteS
JDGUs00Q4J38IAX1w6UBy9+d7c5aBxwBcqwxiHHFBCiNVnzcCMV6yvI4lUj3A6g8
2VeajJgkQQLv8ZyFE8fb/NRlaTDuoYE+7znsnDdZiYAJnFFjXv7ctmqw6mF5zqvQ
tC31jLmps27EqgH1C7BXoqo0gR4ivX66msxoI1wopbQlQW0LWemzS453nR8TS/z+
7i096RRY1b5GGuboGvgHop/hxjKER3Xu/TR2ob6Zfi/L5T76HuQTQNhOzZ+UapNB
B2anrTZDD4x/7uxW6+jLNsYMMopeqODXB3zNe43HInBWt1/JF4jD7kEOTAFvjF3M
PI3fp39XaCkD6CvmzQ/XshAtWH39XdWAeUz8f+H2i3TjMdGe5slqbUjnDvguSNLT
dGXReOVWB1bQbGQyfEa43UCbdqhpyF6gbfD/c5hehnWpiGWL9wkR516kKk7DJEi7
N3NmAbEXEZoa0jJgevfqfYDlUM0MrUJIoegw7kDIkD1h2SmzTKNNIXXczGfauu5W
ok4Zt16cMEcjM2fDQJY5ETWy0wbWL+Te0I74bsiyxP543qY8S9UTkvQsjcs1Rhy3
6Jz3aa+y3L22xelwpAmnMnX6xX+Dyo5DGc2tUhjTGk/cEyEqy/fbMuhXi13Knjqw
mb272uPKkOKNVPjGV67VZQnbvlb0cmTQ7pxISo8AbyTuuXiZgPunJPY6n4/HDcj6
nX9KFJtVapr07lP9agb/zKySr/cIFHG452XMp+4Rr7nlExH5e49geyVlx/i8P1Oy
frmLY5yhzb4c+QSa9mt5vUBcoyCpRG3Pj2xIDnKixoBbI8gkvuupE+ZIKm4ticYA
r0Q4Bh2VmXWVwTVTXYTVn5O4wxwUpDi4loyv+WgvvAGG7i7jZb4ecD98M08X280d
qBX+P2JyVJiN57srXn5Ridc2SNWDhphP5oIZ1C3gp/QnqCCBStPCbD5qX3reHdO4
pbqctqXOCZXVnWcezbm75BprPWM4tW79AF/cjAp7flXZ5JPl3Z/gh/E0AX5nXzmX
tnCJipORpe8stKc25V4+tygoFNIZQzbts4hHyiZbDhrI19IFVEohKPcUX4nY9unj
sPUe/gb3ysfOGaBB9Sa7lyiR4JTWWiZfXBcuPmDv9aWfAq7bwEAmtrdRenIpkpow
vVpDt2lVQlEk3KZhi0rZAPY0BCi3eyb9PoYY4sLh7ORMgWL7cnV6V67++FYNmWin
emffd6qmnexFTYwCtbS9y1c3MSp/ZCpU/ZnnoLxeWdkRZbyDBpZDCDrONXpMcLCB
22HeICjBzXzlN9tB8O9P916l6dn+mx4xHnCjc1szwcIR1zBUQQIwU7bj19YViuIY
T19A5JrtUHAbqWqQhczydR4SohMt71TAF4wAsJg0tly+++NJTKoUTxGqEXtKH+ii
GJQ/i0i+YAxXBZt+q/FYeF3ZG1cfG2WELnjMkzJGUYCl2v6BGM4m2dz0WBdP9qim
qU5wm3Wx25Rlv2h62eW8Z53TEClYrVQsF8WPEoGHIlaAPdlI0F6qH4hZgIalIC/w
ndEfAHm5gqcJP5ppG8l19SHt4OBY0VnHYTCuitpdVr2jYiEjHReHdrqz7u9fUlPN
vvtP6bXdVC09hdLHREVYlGsM0yaDO1QtJI2TQXCMxS7rrl8R4aX0qXpUNlGv3fO9
8R1xmwQbn4Gl44gCqQiqKQVVfN5Wkd5IxbOoPbEDVhL2Vb+6Vu3K1ms3rYYhCLoQ
Sq6iYoBuJ8qhG10Z/xNE7wZFmtXtPPjAx3qVvGQRSgSY1YnDE/E4l4WCa1xjTeJM
1+5+4Z7HwN8CQVVuAb2pTShXi9kKGwyUY+vMfDNzG42R+DtpSgAuTSiBXLbm0Ur4
uw0zByXd6aWJfs9mCNwM5envVn1TIJpHuko5o6fdDLg93bLl5RFLO8URTqwnVtfe
G2XKqCTfA+vVINGjtGxERMzT6TaJZgvNdZfjt3N+kqFtq5XLz+1dV3+Z57OvUDol
MbUrHAuCXS8D+xgCrLSFO6Ne84I/H0KUNUfD+VRzJZxj/ZdmzjYnJLijGrDs0WMM
MP6jLO9Ga0Q+Q359GaSnSwPMmgdLWajMYf0aUFEm1JTFbKhpNs9QCHVMu0kw/il7
Ph7J6fV87MAMnC+N6lTZcWF1WowdQ5Nekzqzi4qbf6K9xZiBJ1iDpAS9+gK4rK/h
K2/cPdQkh5J6TLzolt97DSF3PFtI34Jo/roZRp01wNBqCz2G/k4R24NyqEDXQdcG
LXHqLZxsf8a+XcZyOR5rcoTAX4CtqahfEO/LrCDdB6PlDPg4K5/LNRyAb0KEDymA
YUK72QCi4qgpiDilhS1vq6Pu3l8xmlwWrbVxDhv2dohJ/Dj4Yoghaj/aA/+MKLxu
YWoBZJgck8vwtcsSxux6VYYQjIyCKH5t/KohzeEwlzXtecDKMBTLhimLJfGxiqJ+
0D+yBgff4NtBrXlThQiVfXwOlrXgiTcpirDPv7F175p4Y8Daviug2QwU5Cy0Jo9H
Mn+7X9C+ghdgShH8fJfv94rtKri2XIIe5ZcGRfEOGXTEdoJegWeeNyKuvRzEigGv
yKm03zMD0kM9YqG9M5YvVoIGB0RXpHEcXyTASLL9efuwhXlyGlTFAOPPDFAbCP61
j/DCsOdXtC8S9OwDoQXP1PIF4F3VqqbSn0FaCXwFRbA7FkSWEDjFFeqGwzm7hCQF
Cz6Mr3XTtbNoGVsCknBGFr0H2wqxhxaltOo6mLd5VOVShbaxYbw1Ikry82KIEK62
FaPR3xEsCWQAE5w2SgBWuutzrU9wkst9s9t/3MloyqDKfGTUM0pfe+5rgFUR7Pdx
v+1gVzvOip0aiDdow/+fV9ms2iQflddIf/4P4YrS/tFcfQJ2wWIbtQ0O/PZ4i//h
p0t4Xvnep6Ryx44LpkXD0DWvPa4cNNevQWoTJ7/eB0PdB9WMN1uHaNCgaccQ9BtA
V/9Z8P74a+0TOEBFDIfTAurZPveihn9nQS3PnsykS9M1BCT3ZoAu/+w05hFPK16y
7DWgZzCf5RvtPwh5akf9mtRR++5WsYLePyCNEDtTUzZzkBd/+0dy1Xi/NEBtQFt6
g/5Du5onCV7HmmcgnGXlOrRdqdfY720bA0CZIjYwy+3QW1oEibVttPW9lMtNqiM1
mSE/A4NNKM77L7POUPbAdUllf4a9l6bltFadrTelzg67s4WuEpA1AVTh+Xwqc7+G
O1WEN6mYHF43eNfAE2fW8KhlE465VwFGpOXJNfrnxCnPR0wJ8GasIt+Xvt77jXDm
mFdIHUrebbDxi5jZ04PUnSnyZWUT3gBmRk4fhkyHnrqjV+f0E3FSK6fmcQL4NOSZ
uzMCCekogbhl9VqtbrVhjcg1zuMtIB3UuZl1L5iMShcg2x4ou0Kt68IlLfaeCf5H
fQ3BVTf1Orv1KiCgkfc2d9pCepEaFeA9gXouJzB+wRwOJ1fgEkVPRYRJcVRWKgfz
5lvTSysk6mb1vexpT93D3UlZ/uyuTkMSmZs9/0GJrwiuT6anoNvklDBTZrANocOz
UgO5Ze3OTA6WaVz1e84fVE74pk8c6fttI4RF1JwKpVXgGFGHk69YJCT8MR/SvTyP
Z/4tOvUFwLgG8NIlsj8P+7RHDXuffDa78Na0x/Dcp3f/hdWwA7C2RgzVim2ChhVB
ymvJUcGBywdhxib+CZtm54xS5Yrk0tmVKzH8AW5EPsVScTU1J2MX7AKknl7b3fVi
Tal+zK66R1qRITgg1SM51sJq4G/BJNGqGJDYJfVDEdg0bUq3By46pSvp/UNpaA4s
ibSWSxVhARIDP1s53uA6CXOHl9dqYUEBpXB3kIm2brstD8fWlCv3u0z00GxtxPNi
kLTc7ePDEo2yUT/uvwzMTUc2j0jVl1dehuYRs1jw+zItKI5V4PwX3nkftWr9Nely
BT7LcaU7qdkukNP78mSzRwYoezBY/2luRCv1agiwoPUvyM3PxOBf1TBSbnXYNMBI
bpouGcc7n6UDUJmldavYC5RbDnDpr4PYPyv/Yyeq3gRRhgXv6q52j3iWTObVuULS
Fb5Z/Hu4SYWS6k+Nmz93KINRUhluL1nSuRM5pNxJmMaTtXsJfjb3iMNwaC9Od8vc
YakBMGtO5y44QOkn64Uw4WBuA80+Qx4JSz/XWSBKnZr8+UoFnSHs5HMKkQ/lb/ZZ
ZcgXIf+vgKEKkSvaz2Q3aXpqkAgfD1gzV4FCnEv/eD6avtjzzogmddIjjW0OLUc7
aH6ynDQmOX17NOUpYYa4gMHyTl7adrUmDDVs3OhqQpQa2cHOGrQILXv/k704VCK4
jr4+mDTUZhOYpGeZvIqdf9Jt2WyPVn0GGkrLBb7ZkmjK9xw5ueqyjfbB6B9V4WFX
ickRI6y2iE+H+6M5siFvmZ3vs6chM7ukrRVjYyYrqIDgxx2iS75wksy0PGu1nShE
ZtqHLtpB5cJlghw0W62uwLuD6lcgkAiKoAET91s6hOyxSWYmRNEuK1obdB6+YaZr
kSE3T2GW3oaWi3U6nDzetg0FPRbCRfiWrpGjErGB4nH6yqybwsuYPeld87ARbLgn
Z8csUcfBfGPQ0SzWe4EoSApHBoM9VQJs047YWna01oBjFFZc4V6u9LsI8WmJzHan
p6OiMTiP6Rb9+be7fnSn7AGe9Z1LsRl9DmXC2TE3rhmHYjh5+ZQbgmJfxgUVATig
Yo659zcLLPjGBGg2J7vKvkqSW57/AoaHariCCdwS0N/FVHZzwkFK+U8f+oJshNp1
V0OQ8B/zBvtPNhIde4gBGrgsIkz79FQG2kkk6YJUQYxBv/jH/mIqbQKlt9lKf35Q
0S/t0r5Aqb7QK2VNSfyE2O0O5RCdcRDNDUY/h1Maopg/rwmCuAy9t0eVVi2hdyc5
GEjhFOYC5DJUU5WsROzmwRiEjMadGBdGmxAFOapwzYh/ydh9ii79evF2LHiibmt3
NNTQ4ALfklJU7tpkGZvOIcuqvx+JH2JWSCgdWt4byZU5nGPcORmjW+2SPLS6N4l2
pWeKhOlWVnQH1PywvsZEDj0vJ/ttghraKTzFG4HgDd/SBqW2Z6M5Igde4qR1hgVn
K7Wh9HM628nm6C4xPUSdi5MhmQ8l+i7U7MJr8WuGllMtY0morKvOAz4sM7/CeiOJ
lJdVWjX3E8xLpxOgUsGg2JgDjDsgPjXg8X6D36nu6iRtUtcg9OZ9ozXF5gUgTw3t
S0AP4H2aPqN9z/KBv2HDdOcb1aVaHddcHhG+2y9yB6iJV22d0A17C5dwNH401mz9
lqpf6+WwRBiYyMv3B9rU9ZlPnetqKm3nNtLpsR0By/3in7GeCZvzWtGHhNy1FJur
GLi7e2bq4fvYe+ZgcYTd1nVrWEi2OJXWB2v5aWEaP0zl2J0rYcwSxy1gU58qA2g1
h6PpucmiQUWFwrUFtWyQ+JfKMpMkWBAOlQaT9Aqhkmfx+Vb1sbyM0NK4lTkUeKe6
4fOUMyH2gdMeC2NcQU96leUODCL7D6z8BsVoIdhn3Pi3/3YMG0Yx8+wAOVyFdt9w
+ZjCHAF2fgv1n+UECIRdm1UbF0RentC7JMEuhYfHyiym8pvA186TmXjC7jWzEZnV
y/7KJMkxC34NMwBmZ+B61NIaF+ygFwWK/LOwlE/ZZjBkM8essBDUcIKoQXCvgMC7
zvsBxz4Obd/9XVDfv/TunqnDSHxOYa4/wNEoUfonqA3q/+qNGPGodW/0pmJjplWC
nsAps77oo8eUiHqk4+nL3H2xbvq5Ji8JtHMWPhdctyG1Mzy4jWwev5mZGvJe9w+6
q5wO+H7WXVlMoF8Aa9MLiXGyQk5n++3EDnvlcdVHDAraQq23Iq7FInVofyyfwCfK
3dVq7YOicpPl5AXiFsNtpv/5TyEo0AjykP3Kg2Z3fO+rQUddMwixBRZxqsJ79s5x
+xk2uWUYtkyr0RaM30B5jQPryAUJXIpTMKwkR868pvneYeTdJ9hirZbtQo2Lg6VE
ygf6A1Jpqkxj0QOJPlpRm/LxR6qY22rRw6WeqauSn8xe0MoMeXJ2hDqPEYYzyuLo
xa+be+oUyciGv78+Qed7YoE+LqPrstO2WtKQ8g8zzrWp7taV/o0WggLT97Zpe/ln
jhxO0JpRlhI1wNL9Z6bDQ/aaQ6y0HjCq5zKI7IvIsu++t2EvO8BS0MSOs426OUFd
r/By0FojCOgAbIWMzaKU+0ypvvC7X0bDuOj9rI64PuMyrBDvpjbFEXjja/0IVKnd
4cKpyrIUamFmXNEiwSlWebg4i9Vy9bqRyX6E5KAc0sB0ZzTzWgysyUSccU0aAOMb
lxqMnDHvAIFM8y7P/2Bn83Eg2TsOrr6Cl+7G8U/WjcC/iHjLz7IPA7cNCrEddvb/
XAADOQMeD7b9JeDlBmNdmHb6qjLUGF4TgYsEYdtVbPAhIf/TiO5aohgtgw1oHJES
wnavmSe9mA9Zlo/UD9dmlHKPD4z1YJ20fInhaf48i8OSRS/iEJ0Chle52fj1b8Jx
powSOtBO9tABF458nRsNaa06S+amslqa9ixuJ9hRCWQlCq8xsQ59gEDZh7h0lfUR
tQ4Q5jNnCwiEEILwTn1hl/qT4jhsx8wkTMsg2/MwrkH0DbsfjPIKOPiPvrVSNfB5
Xd1s/9kjzOSDSQ7MCYf+0V8Xt0E78e52AdpKPp6LIhO8Ip0iSiUMvFBEKQy+rPqR
n8xWjhya1g/v3rWjo+PQCtB3nUXH1oSFJQpd872flA6hF217y92DQc9q4DwpUY0K
rBL+h9UzvNJ10ktyVOcEs1FwxpRfa8xIfn/mAioEdJ+u0KnFv51FLIBcuySuuLev
zvuKLVW93vx4TB/px3wUe4yP14rRoR83feb/TzMqAPAccnEBvgafYruiG50Ogyga
bUlOEwUZ5mzyAo+7LFpdBiT1/81jhB8XP/VVmbd33U+Cfiy77cpMeNK5MxP+f2Qz
HkBz4dy28XSwMbKDgS3MuLg0ex79+/lBjfXJhMbgTetRm8r50C4z2ujDU0i9N55W
dq78MWm95mkQ8JEwDSpxf81zJeG+YcJ2ObepudHUjWcWdI/Yk0UfFThBXarbM5QG
0D5dT3Z/A4C2iLlftP3Uy1D86UkTlIfi7O3wuSlGTbfz342a/vBO5H+lg6UIgUvi
HBUJ7XwkXcQsturWbLDdXlfmz7tVWjq3ccLvFeqb/GnUtLKj2agrEjBQCEtFRAbK
Kw6Hr0/AWPQYfwS5kiYu4kSW4nJeb/ZU0uIGR5m+cskV7WEbnjp3k0KLUiqar457
Iht6fp7YUd4v+MvhpxA95koqcwBcZgJP67w23dcSS7ouPgdhq4Ljkv/Lm+X9Gejg
zHTAFprZqU6WYoX0a9tv5pGICjEkGh5ReKF6pTf/npv4SK1nHQmWEQxi/aZh1oLi
hJUW3Bms3NdmzfXXNkUj3xStZsS/J/49KrS9AwN6zmpNNhPiXC9hT2N09+2AXqMj
Nu6xJ+79/G39B1uWQuoOxKEl5qMifeYIuZfzrZWh09yHYf7ytjeA4PliS6L7WNPM
HfCcK3NMEwHGv6dTXjwaEPEW+BiC+3m6Du4wA8q5cVWz5RcgoMMsC7rTWgIDl5af
kDLCQjTJsWu7zEo3ujSv0pGuUUu1ByduHtIWu/OkTZXyUHf5mXLws9OMfseymSXD
zUVEYrfO7ezHAWtWJW0VtHvLZkLOLytxwMyXf2ZxzBZI9WdOQv/twXg5kTCJnz8M
HPFsB3zEfHjSiLvQiErb6UqiDsHdYh7E3IuxxEyMdfj6D94KWo1QRSlCUU8UN1eM
JZTC9zxz/nLjd0W6Vu+R4zyBwnbsZgm/KjStfL5lf5R6Qsed1CAIxlqsF6Izom4f
zv+UzcD1++UU30UEXj2oClVIxwDvD5caIoHgRKSo0zG4C6NyvP2+AkhlPaiAnUEN
5dU7KhBJeeKZ/9kM2LIWzdqTR1qScigIDS0K3lmVoivfhqhLj2MMVsRS3WqWJ49x
JMHJxsdu6dWdzXzqfiozudGOfoM7yj1TiIXvIJxjaUfvFptISf5uOUiiuMAIh/Jm
HdNd8kpasABGwzQqdfC/Izr1cFUMgwRxPhhBZpFUvQDpF+iJnBeQKlvs7SY/U4ub
Auj1i/7//Y5pV8MRBmFXqEskWH3vTGhKDbP0NlP+RRwT3YiXWvtDO0vTCItWjciC
C3WxPQbO5shT//MQ/hixhh4cfBZtEMc9/i4b9dm73p/LilnMl4u9QYGxZ5yWBIk7
OX5Ykgp+4p6NsWhhcAU9fYqfYGj2mXhsELr2YLt0ekxg48gMs+E4n2SuXMxQTald
JGPaFYC7vuiyUBh7qy4xPKLe9s+gYGiWUhJdbXDZWJr0Ro+xWY9DW2atDgstGK35
6JCoB+1wIBklSfWGEav0ogT/SDp2omf7l8/S5t+F1aBy0aw97iNACPQle2ScCEvI
cX3/baLObkREJB1oLKky9/GcNFhv7Q37ezB7cCz6SI/ko0u+WdvSk/mQv1Qd2mWh
CM+GOhMXb9SFgn29UWtm8DUOrKYDkjIqwa0gH9XlLGzw+iABGJqQmnl+QfODTnsl
dCdtsN6/XTsusTv3l4DlyANTqQmNfcjfAnhi2/Ha+MwDlfLhyedhyFym7F8TLVrp
+yRDfDhRqb5WrXqXD1GX8OzL5jfsA2Eqe5z3lzyPwGkr+bj+4jLYdyXk6uu2v7KM
f0VMs9D3euPdEPZL9YI0GhfKBFu7GfXDkRXOvxCwohKzrkYorxjV0v7Y9wj54R+p
p3jsXi7ljssWPJBARqVhcT+OKGncGMU1UTMd+CLcMAxq77NJdkIU84TdcdJLZc3g
RxWKMlroyesj5jpJ4mehHN0c8JKXNbsU4p18GllBE2Wnad7ZjRjgIH2wQANyn58S
u0OCj45fWa/Cq6IVS7k46ZfxKN3+623fyUCpK82mCK/sYBX19xXOKuIT+J6a9dIT
hAnIgZiLAncp3sot0JbtbmMgumHbzVRywa1TJePTVrObz2AoDKektI+In1IG7FhK
qyh9ES8DTGn9UcixdM0B0xqd9dy/9igOoK4BIo/pPd1mUmnBZOyBZoqyoYVRZvWb
1SzUrxagCWSqg/rlf0Kob2nHo7TzCjFHks+5kx6TvWIM6yvXYwt+NzQLD0jaYSCl
zJIg0t5KbQW1b/lbkbLDG7gjq64JdRgVdNxkFd0AejU5xJf4TsLSt4TXLwJMJiSS
Sw32nlzeesSWYFWNUomBvVzoZ6AHeiCOTqibT2wdh80ftSMA1OHsuLXU4qHN3F6M
Ng6cdfqs/JaMoerA6i2kkTznp/E5x3bCZu3+IRssvV+SPEDReLQQDL3Ib5nsFEUl
d8vmzCsdwqHyTnYNUtY+UWg3f8qreltzX0p2XQ0QJPCO8u+gtigO9Jnn7Jq2NH3u
6sBBEMlwSDA+FXcqp4pgokEKOjtT86oKoPmqVTcNjkQnSsZPANffjz2x4vrEvTOm
yMhc7i2tcNFdYa7WeTJPb2p0+63bxEz0jYSrT9CCOdfVAD0xGraRGh1tsQirq1RG
I2G6m8IkRj/Mn/429TuN814ZGlav/awJFh9z7zDqlkBLE0Dd2VasefKIj55vBsgG
IEpAU7utwMjmBuCFKVWKr1eYMjZGRshHN/3FgnxJhJNmrfHBIkjU+ptJcSHhjliu
0N27JdhKmsQ09VY+124At4W2yU9cNyZI9saGOoAUvcuhLCdIWWH83i8MHSNx3kAn
2ux3hPYNdw88ZUWww631XExNibZYkP8qKjHSJw7R2/eNKCM7FXNX/jI1TmuAgJ15
42DtoxhePELmftIL9f+6QRBZ+Lm6/P6w97JDk8D8ayVJAyEP+A3+K0J14U5O2lsi
Orane0O2Q8h/sRIini3SQDF10eITfKKj9Zh8k7ohC/IhZBX1urE4QD8xTUk/pnro
rxk6OQXRL0PI7SLGXKqC1WF6MzH8IswcNcuXY7IYFCJOECG1WHekbjq4xRUS5OKH
xowUlZKdedhhILarL7ezW+Pps8fs1m/AcAldhXbkFfzuV0n9t4qob+iDtmXlQT2z
5pgIDwdWqaflesspWPlNbTDsyW6MlXAqQx/+TXxhzVdYZXg0nxu5loz2ioYOeFQg
Ob3P41UOLLQ6lRinZHV/r13Dd2XkQ34qbm14NgIBs5HzSLQ2TNDOZG1wg6DD246u
ICAEwYEodM5JXKTYvZI6Nf8Mo2D1O5eT9J7POZ3yAMft9/zgNbSIpV3gJ2cvkyRf
Y2za9BNfXUxR7xrn3Z7r5foX9z5oa6P1UFkuVNnYOF8m6p8EVe+urt1GsXiPSO8J
GN0JxL4pMwACVQSvYkNZO/CPMhP1CZbFdi2uyys4XPmSHDew7SFlyM0oFWyQ88d5
508ffPKb+bsMNadJ8aq22EoBrAkt8DVUXP66r57jmERVlPmFxcnTHD5kygHOeuj9
9CHW6LD1799OCz8F6YbgDrv9ZMLveunjx8Ak+L416R9eN2/JXGa6CvH7GVW/NXOy
6jjr2U5hKiK8mjSDv3Ee6e3me45sSeOiHSg5iUI9uHNRRPGirUgfpFiSPl92EZ/I
WF2TOw1ZaNtf1hpwqRaf+vHF6yX2XvZDCffFchkpUV/mYe3o8dDiRZkKLUS3P8aE
0abE9a7nB8Z+ZUAPJEUvQTNHiMnVNgul4DTiFk5jYTnM7jrhe+TcTJNxqNwDAmZB
1PCOWRrE52bndddScNjJ0elSrn9puCsDR6iWiHMyuwrIWmxLK3ksTUgSRSKstmt2
ESyvHJIjHulEYrZjoiVW3RsZtJ1j3Grwin3uNUvujzHHaupXaYlbgPg7nkGDAFgt
GSQepjs+Vq59QIfn5yOWsmKcB3zORXmZFL6cngPCWwRK3Vz2Qd486v8D1RZ4FjIF
19G/Zq3ybwWT4kx86WWdTWC+TyXAdOMcAvKRXBxghbVZipJPbZ3q1EzhVp2wRh7p
RSp2AIZ04Rgwk0NwjKf29LP9x7dAmV/O25jnMAXy+FYA0PdX4avFUGOnhD+CMofN
rJpk+iGmE1EyuPJ3Zgy6i2joCyXQg0Nylnkf7dowMBfOy/vAQkc0eRPXZ2rjxvqp
gSt2JbCOcH/afr2UOjTC1Vz1F5vU/SdvDltvfqrlNNtGbYXijoaVrreE0CGc25Si
TjA6UBTcUq9QTm3NFkN9ftwkiiFhASPkvj2n0dgliZ5a/yut1+jGKmTz8ltE8fuT
cazxSfMvc7TVnpJCAcVFxj4+1kY4Um0boiehECHULcbx6mU2lB3mk4o1rsP1see+
ui84JKSKY6qsTRamcfrtOPgduV7e1z8R7DZaLFEG/F+99/4Z2MEtveHOWAjcxtm7
o8e5BuhoVagvuj04wvPSs8qHMDzzl23uu69DOAjX1TrRnSWbEIcTZEOnt3hl09YD
8rgpefayYMMRmY9SsZYldYCoq8GLdiODobi9v/1xcvbMm+ZRAivPiP+a8Yi6s3uF
RUk3dvXcTCQ/uUmn6N2cOZxd4EnhQyaxOv0t439aLrffMhOPA5Lt0JrtmsQ9W+OC
kFXJJee439gndCVfctTYR494fKtuUu/sKr3j2GdsLCuIKWu0puFRgLwk7C0MgxcY
XNPSCXoocaqwTHPoqS0oLf7GSunO4ySeyKAhA5wooMGGsoiyDsVP4gbYHLsr+ZIn
ceeCocoahfc181QtaHzFTbpgxHsRfFb5kkrzqgzRwasKdgPnXr9wt1SRTPfhOhKS
CB54j77gkh6UeogvyLYWGhfWFtAq8G2iAo4cdBhWKnZWe0/Og7reelR4qiFvDiZI
+FzTA595eX39ynOt1Symz7vBwb1oT4cf+UZsMrAkVEsnYtIqxE6+5vLFKKZi/EOH
RkZlWcwuAN8QFVDOqV+VWRgT/ylBEL7GBVFnrhVPWgkjwQjtboyD9TCVZgitMmJg
tZn2yP4V9FCPt70Z/AdM2Pagr1dri0dZfLmmISWGup7nuCSlbhnDqkzcST1jGxnW
3UHr0TDT9DQZ3L3Rcbu/jkGdGRHOfSB1MTClfrc4Y3qGAbKvPGXABLuR+rq8jYOv
f7NMoo+y3bLNUsQ4OOqA3oWGsJnXTmR76zCvorrS/zSVM/jjmbCCNVw/A663C5QB
f/DnxD84qrs93p+PisZzuDa7mChC9p5wG0B83dC6MSRCzi3RCEDJtsiz5jxkUHg5
ZxOvsug4PndpUBtjNxejZHPF/X6m1SMr1g9zBJvHL2DKu1nUkOdbKxLVy/YVAu/v
YK3sBPzI9wt33zi7ffSdVcaK6sPMPu15OZaj4An1U4JYhOD3pF+/KvutGVr5QzP1
eGGmoZhw8EhzHUBDya+RQ6f9H16F+7xPLhH5F/VMy7xKGAeZg7DdAg895hHh6wZp
XmjK49/JWdZIHbggNJ7poBb3LlUM0H9kKGYi4xcYkYNfRklofTHugfXPdPgvs0cV
dp4YaVFsd+ful81tyVMOQ9sH8Wxa6hd3oKLqtjEwlr4KzbdR4VMghD3N9xz391b5
YYO+IYmGK5qIfytqScSAnuQPyTtsfRGF8so8qNEvTWUqX3mnuZMEyw75fhUGmgjY
SRDqjHAS0aIiz7EG4j9csX3ormkAod88bTMYfZfikuUAXZ7T9HrIcXVFPUnWRmqv
Eg2ZCQwxaGTegC2TQn3K4pk+o0eUqs4Msv5oxQRBTRSijeMdyJ7RiB60GO3g4eF8
tf5v4nQ/ER+Yty5UtVjFN9YDfA9hz+ww8Eu2+MMYktUs9vbkLzNPZ8adi7Hiv0p9
0on6UpXhaUPeVjrcSlAcjiZkWO29nQEMeFBRl1LUZYhWSocfS2+8Sbgd9J+RhySX
HnxhWyb1LwUz4m9dlGStJtMBa/SBtmNQ4cs9t42I67KDnpbf/pz8uf1RAHw+Lh0w
aSaX8tIiwTfphPIhH/OyO0HM1zgGPgUbgw3gUd9HgRF00nuFSKyhbqlZUA0yT7LX
eo9MSHWUBAt0iT16URMW/2UAvV1NBXvI6SRRJPvjY4zbkBg+SqFwUzFe3tuBxev2
ib8m8/XMkhiRBBgxLiU0YDVS5VM5EM/gVWz4quDkF/+vsGrTvSuctDP35v4oyY3x
oQma94a8oNPn2m2VzNInCDLzEkcjSEDYL0rMK1tc4Ls8Bj0Z0pa3CKLaBflkKYdx
Kmd3Z648395R1W2Zp25ae1LsHBMHQwX5/E70g7eUA4asMpFhpE52/U/UltqNQiI/
w5YpV66MHlY03TxkVmM3iHlmh7QpSqOKQ78ovcEzWu6SViEAvhnke8d0c6lIOs0z
m+81dMze9630W7NhszZkoEwNDrNEqM7A8BRLiKCgRXy2SqfvFK3X4uoVtGdACVCR
+555s8beV/8NAp/5pMDei3waVLKdcTcGzSTnGfKDRBFrcPItwx3yM+Dhz5M+9PqD
3Sau8tWXmLLB0maq1XxaZ2b8g5tYAB7udjD43ZgniQRq0hjhdYDkwQU4tashVpdd
m9A9YvHTyhWahlRmH9OFfMzBJDscTbSEb8fnU9ffRdU8Z3supygZ9DGOJWq1bKlA
FbW+i38GL0JsauEj4r4s9law/zxRzge/R/eHKy3xjKhmRXe+czNbbLYoFnRCFYnl
vQQ2aejoA22ZVO24VVe5tcg7I2RDIkYYoAOePogdExwqidNFczsTmR7AYI7QGChK
hBfKFwuPtpbRo1m/GlhVY4r52NSYWJ8vCWhjAzmDGYxtW3QD2JWk9F9tjuN5Fxsp
FhW5CelStjbyBgGzk8gTenZdhzYNcHZZtkGDaGTNwdcUQabBVJNflvrE6ZQyBD9e
PJ2Nr99xmNJSv4CIOP3RxJSVdIEPQDCRULvLpk0bv0hJ9ym7YdNVxNiXlO7YYdrr
EbHmpoeIQ618rAyIafPB1ZchcYvrvAEW4Ftp6FT/AHU2KYKX+nFnpnBI9B7zL0P0
9LFxFTxSliZS2Jx/vsxmi0vqiy8C8pFoDADzHYN+8owY7iyQdjV3UPvUNZzVnzeM
i5O+diY4hAJrxnsJWlbY4/EWGxUrGQ1Xa3g27aDu8FHQJUAAkbcT+KTCkb6bN2BF
pqJNdGbT/gNUabw9j6Cv5rEtpmCp1HXk1d6K0Yb79q+BOoJmIdTA1R2XrG8KG3T6
LXczrJM30IZOPgTlCbF6BmD5hqvmMnwYbrBz7urju75bRuPnaAGbZAHsJwdzAF3C
X6ec+lt8/PVqlrYKBuqrjeEzm7a5mytx4SUiXQo7pP5qk12zXohNxHRddZmKTgQN
GCizTh5Y62w69WL42as/8StWkXZvPOD1jZDRsf0XSjUKrJsxZFPmAxp5LY9CoRY/
ehdDbPybwp5sFZHzD5R/7+PWhwB0C802mUoNk4lUV/qAaSQ6XJ+qWX5Xnc7eMlCl
k9UjiMxUW5j6U33eNx4dFofNB+wcCPrCRISvkZIJpKynkIcqO9yZ021IQxX41Ixy
WfCuUaUUb13xtm03q5GduhkFH8QUHjfOR5olvmVK9XxysXULi/32csHrnI2NMYSr
iw5gPtkpcBuR10xxLQZa7WTYTmTs3X86QzV11nzuPeDsaIDdrlJ6nO/iZG+GKThy
DSs5vjAUCMKcquIJnjG+PXOT5cr6TbHRsanr5Ni4XpSKivRzLsspeqykiFJhoMxu
7Ki98pVndgbfZex724woHfA2e+PAe3iR2bFgj59Bsg7PtcuzXrjzr9jLp+x28+nR
Tz3vjbfCWZwcF2UwsJONoGqUhKjhiDLRq9WqayPK9EBJmZPLYdlt/hpEseTk3mjx
dtDTo5OJ+eS9MYKP/ELrCkuZTPUbNEIg2mgka43nnVxLP1seD9u+aCSu6/Aa4D1C
bpClT2zlHD9KAMMeXbL0bVWVtgqnJV32T7sxxeDp0fMTD7pZSPPQa6uhhOCsHOkX
toqDuZz6YE+sZ7UkrEmceqVoOb8O+rzIU8R9KY5ctTP1+rN44VPs0YndLCsEdqOy
HXfiaRF+FvE/I4G9427PByanJYvoHnM3+1nXKexw8CHksv5lRqieEtyFhm4Hz8j+
TiuBTqrjUKtubS/355BE8CqeqxD9p1dFyTddh7YA12xmpxGTNsiN2eT7I4vHgfJu
dJgxvryPQKcSi+tst9oh/VAod9dnjXCndPsqm4ngrWFYxe/LXNIiDptlveoAUb2E
ht84YoX4kgqs0n8HAowWs3HtIdYM2y8ikFF33Djk2QNptIjNfvAdGcU2/KfQTuDr
h4dW7B6vaa3yiDork7Y3ZfCGntl9Z/PegZ7rtnCNgu72rNuHFMvjvGNIkzjecw3Q
FKZMsnNoFVG0uvlGGPSPc8HXTmp1oxwH7ncqrNNcVonKIWNR1nk75GfL71FjOnWT
HhM62MIO6I4Xwpke5XMOqymkmbQ/vCKnGlUN8e+w7gaJen2w5M4Byq4B8HSxi810
7+ZG5YYJLiU5ekS9CCHaEniuPVVEnzfNVdR8z6POqmrIvl/FSZ4Lmsar+CagLu+G
8J1kO+fN/gl4M4KPKfdLoIdbEkZKGIm6BFuAmjlb7DC4GUkWZ2se3/hcJtllmZoh
TLW61l+f/LYxNqLBXo1EjC9gEsqKoHdUFC4dQ7FxRFE9RbNO+C5WTwu0kgDWlTdn
pZ0AyInXY3knqeR32w22bn0AMe7XB6se8RODQUyLlRJcEXVcpAOer/j3sw+YwKyM
VvoQE6h1HHueTyVFZ1baa1Y4aaBSdqHDsttwwr226+9PM4UtJKcRngYpcr1VVMag
kpFCtMKF9GM0v8u5XIc/VNCfcqlnxG9ieqih31MDhUU/inVk7HxnMHH73sY3DyP5
HxZAnzkCvSzLquYyqIfqurwoccswnMh3Ybwfc9alZD8FvjjPqRUZxNv6wY4jZlE2
bErR4SdAbE038dnymKIrPtAfYvLDjor6uAXsMW8fgEcCc24bMsLFq2dy8ZhKrCt8
9L9B9U9aW24nAtHb67KZ4HHt8KgdMr12MtKVbSjLE/buLU/kS+TZoCKztqgfn8Z+
oLzLlBxc6NPdkrhEvjcG17u0rBad/V1EEsL3hctw7ToNsdWS6lJ1xuFoT7jHm4Hv
dUkxRMDKU6PKlbtTTHmsFfiUXqQ6xHDHZMK1MO0ft0+9R8Nqx0Ak3hwO96oIrISL
OetKGl6trj/qO8UrXlq9miqKwNYahF2kqKphVhRocqDj2mSvW10ZZcDg+5MaMZyq
OURTSpepOZ/DGmdMrtUl8aKlMQYcnBM01eUUih3nXS54wg06qSyuD0+NEz5DD1MD
QbMc5iIsgwLwcKBSz6Ry48UZrpXq62qKSreoiVJXJsKECc+1ZYpbeiIsC9zO8XgM
zcYnkM7UqI6AaBFD3zhlRX+hqRN7oJ1EDj/zTFwajrgN6q6XowjSCGLfC85VsJzi
1rW+d1ri1H3HPE90lqeQyInqlijr3JEJ/7G1eMtOCP8ww9COU1xPoKPWhq4jxLv3
ws05F1QdaaCiKVmAMmPPW9cw3UxREKfkEFWgx8QZ7a3Qbx+8A3JOnDcifNltu/Nk
NajJTeKVto4OGQbw/3i/tniOaWkGnu8VNeIVYu4/b+xvGioQec3+T7zUUiaygvDj
cfZj6keDs+XvwQc8v6s48YpPhPp4qUAph3Xybb35MQ2vbDfeOAC54wCP4S5kD2S3
wq89Nl6k8posD9nVxx4nb4gZfiXghHkBJQCcK+lAJz/0xOP8eslg2nv2m9a/hjeM
QI8QtgSpSa7DAn/O6q5gfEWGZxbQIdQOtu22z38y55Z/cGAex/bKjWjYCUbPvVf/
By/iZAyenOi3jj6Hdw7LihxJABPw5rU1iVoVDfNwR8fXrFtPOxFaBMFe6tncl5GH
Ooy5TvX/0BrLX9HxUWS/ZgbxenscoaJ1mzSqN74l5wotVe6Z9z0fsudcTTQCDnVI
+NF8c8nrhKn3ooO4NIoVgj+qri78MMgvMsOofWjGNTgirgExgS7dtcuzwLZfOFOe
Qh5tILF/CPTigm1Y4XT6MEhE2fVle55Z6rZ76dAmL2grRP9skFCPH443ZZ/eR75X
0HaTD18yskmN6dJKtoPJ8Z7pkc9aM+6QbM7HqxvGXkSyJXDJPEkkxjDQ5pjz1/4q
pAn+rQemxKCUUtn17LbyQ1LrWb1PbZ0NJ9A5b7RJ2EXIz/7t6wlpOf4taVKpQIJ7
xWEArD7GeQWm813iTh0T2kNTrgneYrlKti5PYxjKKgNdbWc3PGaFYPSRUrwp7LSW
HYSGGSnNEdvARG307yIijV3gnNcwZIqOrw/unD1apflYppZDz/xQvEnJ28G4S0Ml
zFSWZDcRsVrceevTovt11mY3K8hBGbRpH8Ai/YwUC4KWaG0OVobVysKkesErSpC2
yO8xBzbO8R4PlsqXadKtRJ+GC93dgnRAUEcz/P7ckFsJbc4ILOtHCFPScAUNZxMO
Dc4ggsYIHxzbbynEQw6Vo93GrWyDkzoPnCiIJDzfSQKm/DJn0fRXhk3Ofh3+8Cn4
BOJu03U8aE86WtJd1ky7gvZW34ubfN/CFbzwnDTj+Vc0g7pk3Vi/ZNp72s7D56Rn
7nOQJCLDPmsGIrCMWC2pFbvMpI+S3iwUDwoutThMC16roeMyNcItozsKa0tB3usy
05BwCFpaMG45PP7O8kLF5nCbYdew4hl6H98oswd7plYOeRHGppzVyJEksDnP24iC
8GbhO3kS7IhY9gO+uwBI+sJC9ORFN/24yhnoXvXUgzc2m1973vfDlixzThIiDOU+
EdcdjY1WRG/zQmzO9eLIxpRsxHedd9p2cPHIi9VMzJfYnNNckZxQ3xOHBTUrAKgP
uie43zJILwfR1fN3Z365VA2mdwIwN8mn35afUywHCcM1lhTZMv6XIKFMhmrIGpzD
ZHsMqCphihW2IV4G0J6ZHG/5wK+7DW5C9ZxsRyQyn8NPy4md+XjLnXadA1xj7qH0
VZkI53PF6CfHblXa1d85gCYgCrc+OYvl5Hq52zjr3BDJkixF7HTx6Vd3GBocHEQL
HqhVj9OaYGQ5RBDrSP1Qsd5N3/48XkQGcBlTsU2sC9kyd7MaMHvVQuXPfhVI1jcM
w8UXdN+CQ+enm6uIIcAG8gOb0JhfCzl82VA8RPFQJNNvN+6AjZsiQWfBLxuluNah
ZcEKbHr0nYeC+Q7BicumDLylvFGxoIc0jUZgPSF4dn/uETUkPK2YQfAXxAbBZR43
tadbf/omVctxA2OTCdn2X2ojZJtTmEeo9XPdnTcMZFCRctWkX+0vwhDbovCl4/kC
Sh7r1bkM/lRVH4aDfrEDatXlUvq3V77AQPAEXs/QJPsR1pNIcwb8gG0EVcnpel3g
w3QIVw4YOXaNSSdbVgEKkFFlS5VCQUuZkr7pLwdwPeFb62Pm3nWlBXDguxdvckDR
Qkn/8uHdsITiDY4oyVHjW0H0QRzWnDaxEzf9DbFappeCjbTOQIsEZPzMh5vw+Ghs
qtS8Ik0tabODpKlUbcIpnz8/7U/LTuBUlP+yM6t9qDlo7mjKpql8+qyODsqRqc5d
bnw+KVZngnYL/J9TU7orLT8KMoIutCG+Jy1sGCS1SsCN4ETic6+PE4tWsYRyPwUa
VFSLWOkvUpSgxX+uzLem2UdPLWVFHW+L+upGpHckZOTmaFllZv9ohtDwQm6qV54e
NVmLaRwV/j+SOiZBZPjq2oRSRljdAdKV76q0RpXL9NpyNOeRPTew3AqN0zB+Xve5
l+y3bqemN6MuXGKQlNkBR6zIngM65JQCl99LOR/JwEJAC5FrFPiSt4HwfuUun35a
SFgWEgPVq9AN9sVjsgLKkDMHpRNG7L8JgTJSr42wf1IOsLDX5p8JD2pxj+LQuDyn
FOZLTBOben8LbN6bENv69z6zUJe2z8z2wCXUz0EHvRtSCPlbUK/+7CCGhB5xwvNS
2kz6poSKM+RTa4Yr3OcHyAHLivk7T1OpFOE6ID0eO2b8VuxSBgr7KrRoGK9zDG6n
NfRv7DQP12dgl5Kmz0C5wNy9dtDXxojNvUHZwqn6S0YDgkqL4UsJgitqAcnfiPB8
p5Z9wfIyFluCpGFcKkWrMQgvnGXhXyVp3F+aTPQ+tVJ5vi0oJso8njIUNrV+u8F5
B4XSQkmWH1wFi+4dX0IJ82G5LVwWkO4lUvNQOrS6cQaD0yh2C6jC0WjJzaWOiPhi
7BK3B7ghE90+yLUWy9NmRIp5yEaAmQVTZ76ka6U4VAM9Lv4U6MNMk32l0vGdTGti
eNGCRLJmg2dJyL5teYntzhkETkw2wwMGNMu5oGjX7EN6C5V8Ia1GpFYZEHyNWx87
Tn/Cs4lqcKZL/BzjHVt4nNYEeAZ2C15/tZho0BZPEt64jX0iya8iX+0gdwZow9Gb
+IT3C4DVEIu4Nqy3bHCvWVLR2hwGDoRLhAjBIq6u16STncsAH/DGy3WIn3qvXohs
iuFu57wQkb5wcwU0n61r0sv8/8TxpXc0k5MC4uEN+OpPxFyo2vr18tUk29uSKKv1
P5C0FgJQoxsDN2qWDH8X2xgw9eJs6BFdXEvaMofk7vVWTbl36nHhrZ53CrYJR0G3
dMeJm00UGKygq4Sh9QM2g87/VamwdJduKNJgv9FP5StsWCDkktCTY6syFoADwZ9h
zvZfKOzbJyX7SBG0PYxmg4buV2ywsYPQg2cbf3JljI9cYlKMZYI0tWb9sLgkHUvW
LrBAQvTUTbWXd9rbTUG5IsWt/AQjbtcWHKC+5NUwFbt49NIFkfcaBkaCBPSzdwOx
lfM+1oBa56PNrpjyq0KgjEYxGvY2PHoHZuuFqb9uVavhFOysKoPgzTI1dqGWvBx1
0dhRnFukjjLInEsEJOaHDI396D1fx3dsq1oD2ULgt5/0GJ+XR3cOS/VAGOXDB8uY
xLzlSZ/9h9BE9fwhZLlljI7SH1HyKn0XMKkiLHdVYYiP+9gp3STe5kJKZeBjUKBS
tz5zuow16lgZDHBbdhArzflGGvwOO/blKBdoF4fRHu7fF4aMn47jWNGBw7qu5IHi
SgygXr9WPBy6PBSySF2Xxc5p5ZtLZGSRPpgnwisfB124ukGABcel3pCj/NNN0u+d
nMYhn//WZ+53ElB6P21btQA1fg+sKI/pS4+Q09a8GRlGbfpPuAPEESYG+Be+eLDh
j6lL0UhBBDRV8ag3+q9URAll7rRQ1TWsBU+ocAcCWGqj7ZIAJdNr7MsdL8SQnfMe
NEB1Mj4PFrswuz0+PF3nyVkRnb0PzLFdAwxGd1p25ESXjIxdnAWIk5TJGp33iSc7
9F4znpWJ+KKOvkprLKBKCGfWhpulutRNs7lftoYbaGXkjEDA9Mn4KTiJZcYfMTAT
npb4OcLXWQRrrUa4GhRIXYbF44IWVi2S0gp9mXRJZNpZ7nRWugwN3PGcnVu8makj
gLjH5LN9c6s4xk20KZUu+5z+cuvjblsHnZd+vvDUaltgOm3tYC1gD0n7uQEQyrk/
3q/6wWMbpfeRc3QUixc1O/EpdboCNmg8FDP2wH0cCdRUbdAKIAtkE6m3jm4aMgfD
RvKvgkOfM50y8DH/MP61hH6cREEm9Th2CnD8VBNQx6slp/z3h2oznQQs3gG2O+Zw
94ltaNaVSMF72r/zEvdf8lYYsyX8CWR6AsscoaVmT52ydPnF/5en8xWXUcirSDR6
rr0gxVOAXQpA2HL8Y4rR2zTKOI47hv0yZedQTIY2a5PpSxjKQDssvYRnM72s1V/d
NtdMkqfb0dzUaVP2iM1yS8IKauUToeIQkAif3saU9Mynh646gaCbm9rw/ztjKo5c
Rk5WRP5tBAYYd3YKcbhNO/9qy/ymjCnb/EhoQYlX276+PGseTGqkuyTp/vCBS6FI
yne+rVCqHmu3XUysPdyJv6AAa8H81NEJqZQn7xs7DhiQyOus14BR7zCLyAe2Jicn
uE9k5V9ydjAy41+2W/knjojYaoKPL/B3BWE/8Ghox7+cC+FYFWNtyu8MjRyDb3Va
F+jqJZgDJQQgUvZbF4sbXAgsSRd+1wwb+/Ly6/VOtf6P1TawA3jHbW4I0mBgkU6Q
Ulrnn8l51z6xJ/jWkSX3BGTxaZKGYlXj3rKYJDOXiT1nuHF/V2ePfr5e0PrEU0ED
oWv4LgVGsP2cCq/IhqiiBsK1B+e0ezlPugkA4L6uOstv/trocvZnwctSKRDsIfW4
d4KGOrnS8yE42vST7FliW8cZVsq4D66Hp4dSj8EXt9/nnr7pLZBvMLMB4U4Va0BB
2IFuvL6O28k7Yr+DBcV+aiPmpnXc/Ov/5Ohvi8nv2ZN1Pbo3saJaODVIsRCGvxkz
pbZE6o4NE74L2ENwfl5mGrMoGUCkg067Ze5z2yvEUbh1hPgyv2kVFvtChQhtTMAt
xcfH+aLlHU7zThkCQp26fPc5tmjWVFrkKCOrzmdeJhyWP8SIwYmLHp5ru49oLVhI
ZDlzZudWsULzflnVQQXXrKIkE1sI3BqnaisN/KDxMzk50ZRR8LZ2b7D78TzYpDNh
Is9Su+x7009/yD4tK+o4YaOThDPKxVqhaFPTpzdVy1ATxGwU/esJwGYu8nHKZuxf
pvh7nAjkDZfhIqfC04a6fYG2xp0N5gSLig0y91dH16ghrkYNgk0Qr6AsZEDq41gB
juSziDvdcG9HxdyeFK1KBo7LId4r24d0tydgUf8pEr9coH0oNiONuRkp4Yh1oOFn
PBTLgyJVIGoTVdtHuaEiqiy6qbjZ9Nv1LeNt+LqyuoUHQaDuTL0ntg3qQurrG7bh
zk/HMfEAoHdmyiPj7DzoXoq0++OiZoID/yhdGFLwPTGCVfN1jTwGH/l+br1uQGhp
AbkBQL4TBp0nH9lRucWGWiW9AmY7Rvf4470Oxj9mywItd4jxEHP+b8wNf8smoMI9
UgZGqgQYqiaSUDlxpimuFNeGzb9qICPvVOcGyFWKrdZ7Hzqu6Z3AXgmdUfsCbYWQ
w5du59zOkklrBFihtObFyKFhB2eiNxQI8NxIfj6bOHoe7DVJ8QyoB1XsyiLkmo/m
AlcctCuj+E8/13cS66+1fvIr7QDSibSYXOfEAFebxapKs6F0PvdHSxuAGXXX9dvL
2D7CZLkkvyWHp3bhQCsmIUQVknSDYQKYJ3YSUJZ2cfRNXnIZLRW6/DHtSkqs4fDZ
FCo/tteVmqNd8pRnKAuZnA0hDmsTNokLoXhzhbYaC6m173P4Mm2c2Cj8an839iqo
XRDoX6mt0V0Af/AKJncQVPROHtxiA9kVrGFjyE6YgL1zVR39TSJOrtXGuXQfvRiO
fWE0cndo1sY9BAYoRM6Q2KXbpG+ddSmw46GYqKFamAVzggFPub3O+Fjqc2Xn5U4k
NZ/cZc8Ne+TYrO0qX8gcpusS4xF8QNduoV1wyGcuKSL30ZMfgRaYD2A9h9LRWe8J
S/2jnnNLchxb9682jTi9ZUcqC74YQhFDVwz7BGc4HGIMAwWNJGvkZBLj+cM+JsHO
I6cTtETK0Zq1bTDlzvyzdBCOtq0jUFZ3m/k8IwtgxU7S6iXciZxZioynojG9xMX6
T6NKE/s0H+MknU3OJUs2KmOVHPiUYU8OKfPUPSFNyI618VzTy5YdANl8stDKRGxX
XeaTPAnV/yzyFb6d84xePcEbN3RSX0V4VzzAgqNk45wNdEBZBes+q41SxwTV7jBg
28dVOuxBmHqpvIcY9dGL+uP0yWvx1/crQxYIL19jlBhMIPwX4YtmqPm87Ooo+Mww
GmdKNmf6jWIJQcXIDHPk/zqG8++k9e8AH+VRC8TYUCQgWotA0BDvv5eN4WientK1
5KpiAwf3An6oXEvhjGW8floz6EqM2/FL0SLyS62C3PIL6Xb9eD3L3wW/qmVHIg1F
szxAoeQQdvuLWk/7embQrTupv+adDF0vXHWZfL0OZaSgxKhN/MZgUGriMuMt2cEw
D/zNQtfniKTI+XtcDms5KIlZWbt/AybZpXLWM6ghn+Abfx+mdWxre7rYPNsf4fcN
td319cMPCbCG1IT4UuX93KtJ0HWH2w+BwkUCczZd1dtr89xbx9iiq+Hf3/YeYitf
d2hUvmYlmKo9u0ggJyoK/BFHCqf+oYf7i4CGlwq7QQK1HqHtpCKMXJKBcJkyTloV
jn0FgomOi/0NGs60hyrbRjPjqXiAzvztYvzbvOjcwPVbcYzceNeOE0Tfl6ZhXnvE
VCbUYXVtzpx/V01RnCmd5BSmCjJU++6YuUbbC4v6wp3RRKNH2ajdhNcYdkPWa8xM
shv72/Z2ncYPNbtoLTj/XQYC1KyuF8xr1A5C18CgBER9Zr6en2iH9DSPw1lDoBQq
Zj92dAxYBwOJERiRrn6JD8p//aXQ2/NR7o2QnYXrFJH/WRmveBy0Jp4QEQ2F/MTO
+9OaaSlF8Cv/3LOmXgi3UbXZ4TH4WdONoMDcL5RhrkffqdjNZ67HP6FhUsiAt/6g
kl9wls8kuM29aupUKsTMSP9UiNR4duEQQ4pqb9v8/pNWDsa56o41o/I77OPQ0fDF
hakQjo3pJ1OM68rWSTcAD/5RL1jxdOHJg5vbXipAf4U0dNnFkY4eefa0JAv72CyZ
JO8UjtTURn2FAszzHBHioY7s0HvsFtdtR1Q5qOXNvGThFAlcIwXvaZcoSX8rrJxw
iQ9tnt5PSJ21vYHF7KgxPhQYY77xSN4a57gFf+OTKHO+UuAA5lDQN3ZOs3LfvoTl
4zT2ZezzQpSRhlhqTkOV/DkIOQ3frQn7hLHkDmTrEGtSx0XGVbtthWuY7LWiCIu+
mrtXThODukAuIjyTtfh6wYtceqb9gGW7eJCWKo3ON0XEhQMtgfSab8r/3S3MxBAH
s4tCZbAAlx43fpCFh43OSmWa5AKjxbqM6xmBgiPKB2peCmmWhYxK5MxqXL0XQNW4
qjpKq6c7QS7/dmUt/xSp5s5HTszVL5ND2vm8Zrp1n11u6DI8cKJQPLFIX4IHO5Bi
+IysdjH4yEJWmi9fGqum69tQBFxnbiW6zDJgB10B0iudEM6nVKbtEw1vw48LhAEP
1AtzhZfeQrgJscT14be14BOiENc8FXefjPutpVXGvsMnGDTkk08vXVc7C4ORhvVt
eJp29LOoqq78m8K5nLBOBslITP3uWJVcv1nPngCoZgm5O/uPejE86LMxTP1DjtfQ
ljSArH0rM7YpPiBlni8DbYOxm4Xyyi4P4+u1uf01mtHl6VDjbDP/BWa+BZ8vQsQQ
kD4xOoi9ho6VhGNv6q6RleYixG31QaNpwjBayrIw/KTJ3hRxJlqCIO0qJ1K6Eq8k
TE9oSoD5vUVnT40mRtyHOIut078NpLSOnUHdMIjLcw+ZyWrJNaAl3/RbV0xMBNUA
Vgikt9FYDQ1HVVdyxeofjJ99A/tAfE58TTrfKfniPH7wqKz4JFc4vEoxj01MHZmZ
GvaKn4/vmVka+aMMacGnvzsJa1Hcne4jModjG5WGMtEY/1nxKyJk1JJJ+1tgRnNe
j1PadOmBRsBeKE7iwBtWDORCDruhZvkYfL+X/bHz106lOBAf2E+RoRGB7Tj0Fr5o
lWvAuWOEBEbPKpGExsEdcT9OHCV+S7EjwB3n1FAcMnz4YfBZVYkZvBt0Zon/adi4
3MUwZ8JxO2QLPnUBONasfueAJFkb+coR6X1/C+3H1bWdG9IN2evziokW0P2mI1L+
JXXhly6thvlGeRGp+L0QTIZZV9RuwFmTBrcbWfWB0hqppqU1zeiWsnuxZtb4sFK4
oSOdeekDwcaNZ/XsMr6NbXmybMg7sOF5vwEOqzAi0ktC2xQLPw2xYgvdFV8KiMNu
C6/Vm+o8iXCBW1hC5NvoW22Z2s0JkRzyKtypsmMOp8tGbUqMVcZmAKzbo+kW/pfy
by9sCj8IDiMx697XOy/BfDQH8pi7lgHABHKDRxaJEUu/0HyiVrO1xy1fuke987MM
wkoLR8I7AV6hM28kE6X6uWGAdo5rAXtF5BVUXC9ZwXP7dTFNzzs6pxft1fifta5u
TrWg87ugo3YN2ZZGR2b1x3GUxYu6y8o5sd1r2Ji4KtGbPC/Ia5Ed/FP3wkLipaip
ws3nhwtsso4JEhN76B2b+PD26kFKtolIiDHblAjZH3i9ALFyIDxHkKL8IDAhJnnA
WN8XzDM/w5nQvmuRkPsOkbmtikfGZpeiL7meGQlIYztvG9umS9It5FzQWh7BcCXL
JKr9Tg9aQHIfwmuge/OVZsR8EqFJ11P6hnAvJhKCvPEpzo8xWHYYRWSK1MT8wHUm
PgQy6iqvTaNn3XBFCMv+oiPIlLNa7bW9SmJ2vgoZiOxNyqYAlI03bc4GRDsFcJJn
FZa7x/zggvOeZBZwwNj1TXP9EBtgd4VYEmnKv3+Dj7AjEmHCHG9xej9+z6yp8/mq
Zwx2g3RWi53qUmWUKQycPyBkEiIH955zqycnpFE94gugbC1vyhan4ThkiQ1YHmFv
S31IxBVrdlG39KJC6CJqqiGdflbSC1nGyQ7LwiKJ/DkXlF4o0KvW4UHXCsakLvtI
8dlwlsBXPDrA6eYqcq1Pqjl9FBqFOf581PI5fz4IovOrZbo878j126kLWA9PX0Ri
crUebuYjWP81s7zEUAfATcaQH5znjIbEd+EgeMNHfaxOaU5JDB0by+tiZFe5bTuT
DcJfEMGUA9CqMkaphy4LFcUN3Za502GAmsOdXW+ZjQoFwx6eeK/ZP6EFdLRR6g/9
EXFFFYKbS2akpM4enSb64fO+VGF4CbB1k7F6z0FZ1xP+zq+suNQYtSHmxpBC4NNJ
n64oJgvnt2cQ1yA16dHwzrY9Z9CP3e7aH0fozrLRk02zfTYHLWey7hcGFRYo91W1
Bhpg/LONPYPO2yiTrC7eZ9hHstKe5AKr6j4vXbZJ7z0hV89YIm3ZBS0RxyzxxYgZ
FUwdmS4KDbqu2g58gu5XRUopUZ8lhdsGHxHF2Of2xwNwtFyUAonxKxWjMcS4LE5w
pFm72nh7KRleclHczP29xfr0ICt8J4NOH5wRAd/so7iSIZ9O9qnirXi18+hLUCDB
aUaNamiiKblz2CCd3UPezGKkfRsvvWHmTGTwidbxXYWV36fy//hRVOdsHq/aF3xg
4KSRq+wiVZAug4xtF0WGQbLyUmjOrd1mqnZS5gQDCV2vpL+Ptq/RwilpCJSF05C6
bDZ/QveN75dbUHGF3jZy9y1VE3EL9yZi5NttP35rCmTiKKj44B9OPdK1WwnmqLqo
6vEfF54HsRWIGQ4gbzwP27Gbh6eF5n4aYHepFLnj+yBB0Go9TvKXA7UxPFPzNUob
GselUbbSs+Sft2+5QwrpcWPmQZgNcm65sy3+KkRgBYom7Jyy4hJhNP8RiFRuAzA/
mqbuTBVA0sZ+tJihzjNAt1Byh4m+vRpRh0rqxZjDz2WTcjwAC1K7mf2awYdtE675
yqQTLBc+rlWAtILrRKmP8ZaZowMPFpYIdGlaV7dzYE/1NQQ0LAPoLpRuwDYbjaCQ
++fBEvKoK24UVcG5ho24jSRWdGGbilCCmljhq4S6lsbVT7gcPgRtpVg4LlVsD6Pa
Hsf86K/UrHPNqzUsP0Nj2xE1d5kDfm9CwJADUOumCbxP972aNf+89A/tanCT/TlW
yvjA0M9RDzNW3leVdAjRZAEBrDf4ELSukXG5VH+Fbum0hVp49dtmzS4vruptbwHl
ug6YT9vNJDM+SONf7AuIuTw9xNdV53nTfyR400l1yTk10nhIyW+Nuap/U64Na4pa
++3mLugTjwSoVKSMDfY5iOQdn3pcfN88eZ4az+1f0g+gDV+3Lu170z4oI4B9EZzQ
mJxNzCMNlA66mxGcSE2DBhVNW9dGoKTzCc8+XqtqYsaNAJKjUoZA8tR66274YAlV
wwaYX81WLTkdUfEVJsmRp5ra0HdBHeQp9Dei2l3GF4M6pKOFluu+CIB1q7gb9ETd
ZzEHXeaPAR97kJPbGwkJkQQGAkhTk0dBg35/P4JNrTDrSWORh4mhx7azxaHlYr3c
JpE9MOIvkftlAdnW1ilhvuD/qrNIYj8uP/xJ5wVeiMvP7htZkY+LoleQLbCk41dz
gGtDqEdpxS9Dmxfc/9XAATPk7KvkeF3ErwqRMxD7dP5oM6h5u1a573mXjpb5EOv4
vi1NoWBcjBcvkWgI6yXOY0e3OOpusSi24T47YQkLweJL1N3sbDQMIEkSpTE4Q51f
PlBpSBcIjW9TqW8b8Wuci1e1iu7nyHNGk2xiKYwsELhiHBvZJyzjjnrSSBQeIP13
KW5UjaTt9+lP7s5Pd+R+6ZGA6192Sjr3CH0SMrU03TGh7e81SLfRd2ZIaaAOuYwP
d4Szlzw56DwlS9iecLd3Frk1lexUFSWZcQnrfeHDgjjE/yOYxJWr6ayVfrn4YWsB
mBcjVMAFjdGx4MXrD2p21X4BkR+Gl9eS4fxXREKjupX6tLw02yDzD7A+oa6+hA8o
r0Laia5YlfOysZ88HWThSTWtvioS5loJsx04HA+4juBHEqhmlVjk90co3EV8N1GS
CKK6BA2GQ+pHvjQAy3qkf7eHmWw3reBdi+EV9pDRfSvBjuctJUZx7Co8dQivIggp
jvCs7/9puM7aBgYX5yIFrMO8xxHCeo9/gfoQh7lCQYR6oBbSOuGW3ZK6QISq/eyf
9wOPgX13ZR5bAvl1GzUNT9lgyz+fSh2/DLNj0daZTmxynZ18Fu4PDMnQVHypfFMo
wBh9pQYQ1fqDjXn6zCoDKXYq4UAlE5y3vbwWmg+2pgSGhrlgZQTgQJscjtrM3+7d
9lzIn4sUJ2YF9kgo7xY0o4Af1ILPJy3JizM623ItlFDuCSck07b1Eo50aJ64w9Ba
YIfZk/2mF69kdPaxjep/JJP0N087r0r+p/TGi5LpeS8I5ZCL1XWj6OT5ITWizgRe
V+/hB744SBE4y5geKLKZ+3G+KvwONZffHvUfRL4a4tW5By7L3jq8bfx4wSNp0O8S
zOtfw4K5lDKLiR8XZY/YsIVgAfUQ6zN2uF5LaY8qBTiUBruqScHxW2ctarrXGy0+
Do3R12ZQBHB8muJ9E3wpJltjt88J/LeTcPJ+cbhHmx0elj/BklQNmi53VKQSCgvr
2/cZFT3Uj1IMVijKP4nYQk/pGzXDLlxVxb2M4lIwBYv0qmP4H2KJs+bk/jG3qNcr
u7vDIRQo55n3D6v1qK/Dmo3D4mIOkF7BbXV2EcCSf5p7CXXhaeKY2z/8V99rSmzS
efQx+jyAXBU4a3YxY3KgH/7dXYvITBIzBmCI+7PHqY0y60k38qJC5PZaaflD7xBy
r/6nLXS+TAOLE413dkvSqaUAGbm9M/pBxANtMdXGH52K2Lq4IYAK/uDGy8XyJPCn
1nFNi7Ren3ADyu16UOisjrBD5YacWUGU2G1JTqugky81S1dtZmq47cKIB/XrGhTr
GwXV0T5UJsibWg/wKCIeGWD/0f6XzOpbltI+YWZr7j7p3NH8fpPYxnk8YDPUVZ8T
c5/UfjI4hr3BvL5ydrx3R8PzjrG2O75ZgQOKBnPJvYxhaCuAntALH5kuCJ01K2zp
IoeMuuVJ5CugtYzyUF+YeTw+D3WxnDRimjcwsPsBgLSnEThVw0YWCZYyiHe7kHUP
mWyi4PPKP9TTWbL/ayh7n5M0bGkEdfu8C3UN7hSfjzRDIOXnx9gXMzyEG9HZXWSY
D0R/v3JoddEZr4TbRHI5HPUHfwyeIx2cdfzP2w3MivO4flxr04s/56KP60h49RjN
4mx/9z5vFrQOgtOvXvAZI0vJ3kHFHoIJjBK7gIr1TbzFKves2MSMIXBx6krur9zW
9rrfc/dKwv3180CX6Y3GnHPJGHrXfUyo4Ft8ycprJepugGyqEYBrgc1ba2jZUetO
sALpxN9D0P8HQeSFEHdh77WK7NEoj280dh96q5qJI9JZKP0w7JhVnn6Rb50UAs8t
6jp8lrJOVZGVH4/MJhmp9K1Jdjs+1Chi/XpsUi//HvIetLxa9O53u7nLVfaabbq9
i7l7aFvSk0a9kvMrlvI8/UJW68Zzas2YRTL2tVcW2H3yRXEMeLxh9y18PS81Cp8z
uZrj1s3dnheB+BT6B+ziCkFNA1ZZSYyOjSzhLs6qSNTiXoAfrCwxD6CJ0FZeolW0
xhevXbUeWE7Heh5GOu4G8OGm/bgjYaApNjLijuoiMv9dP+kHTCVt7xOaCFVygEzn
GK0lEC6IgYng7UNj0kLQ0aSj0kf/q2b+KYKY/p9EXKPIUB4c6el3dIy+Y+lZSunm
bI6lNtQQgx1SeUSlKkp93Yzi7Ib/wsD4kSzAlKUjxbREokbNIij/PnjPwlDVcJ+f
EHmNnpc0bxqtCNBq6O5tIAPfq1jnHafH+w9nYjPOgbwGgixwkG1yQYH1w58S2ttq
cLRC7lF36zSh6FD7ANKAJatu4ZbTi1R9cvehDesaXoolMlPqwm9xVUke5/qWsjfY
wHxnVU4pvsNCp9rlQ5LqONbL/Ev28FeiT6KAG55Ts8ddv3jI10lrTuxcgC+7RXhp
nlPybDfSJi6cO60JEoUzuFqpW3WwNadeqqtzcNqLcjdqdvWAv9uXNbYi9eX1Q7tj
6XnuTPl5MBuVZP5vNZ1xBgWM4UBcF4YFgnCdHKC56CKGl3e8C2b3wnmBlj1Md3fJ
4+SKhwu/hpDQ05PvLsVVYw/ne+eTnYEkv3SjU5aViH4327VoOLKoai2gD+oJsMWz
7OL5p8w9YT/8EbQO81pos7q+BZfk92TCkQd0W1YEEfE9T97lkxvB5Oqg/Vre6F+3
Fs79jMvlgChStk2X/y6qXV1hjAKdaLV4veMRgz3RNUCe9/q8wrgRxwSsEMyDBYoG
mFELxK4dq8wLKFUxm2G1B87s/7LY1Fioj8lBKRMKnZ/6vVw84UD4qzobXNePQ2+N
XV4u3fr0fXHCSAMQRuy3SX0leiU4KV0Vu/Fs8yuC9lywMGC3NTz7VX8akTYYw33c
Lkvr5VLgfrE5rXxkeOB7+PhFRZWKxqQtvB8WEVwzLbjAm6mZv2v9DxhTzB9Fq2dn
nxCYSDCm1lxuphETA9DQR77PoQRkdcpQNMtY5tb564N3ZmYvwi4SLCoj/v00tvfb
OStW+pGxCstyj+5vcyC6T0HOOKyhcBKdHIu3hwajLhwyBowZT9U3OtVfAWHjPwjK
ZmYJ50JMLlCOncwWWeLqFb1c8levbf0jurSh5YeFYyZ60ez2u92rCZSPN6rcxr6G
dwVQmzQz5c3rAsmV5JlN6OBm2QxBeW0IFCk2FmAAMXN4Qn6LyreGoDHi9Aw5e0g2
fGOOToafLW+Wsdsh3J2XZQD7DrZ/2gOv66pJ1rbwUn8AHJz3Z9BC/vyzTCPHS/kq
actc7DUpkl/z+BKg2zdZCknaZyUFshVZBYsZ8ax8sP6wk39r88mfb2J8HXlktal9
+MF0Auxd2BbiN5UUGNARHkOpDv5JhM/rMwUCP2V1lU6XXj6+iXkrYMStrsmZttPm
cYc4vek8irY6CTgVhkrgeqNE2RPgkMU19IrImBJn3eKiw9/7tdy9GhOunkPPRnEl
u1p/804wW8uy3I/ieDCur9Bz7VU9U7jwnECejk+hsZsYxIsb5+e3WkwWQlCRSbUy
Bog2VKuSadmRtY5uPzl5Yl4yJBng10OnNQfQcic0etZ4b0+GCkD0fbvKW6d6dWgp
8uAw5ylbL/TfuJelZKKnCdxglnKfHvLN6r/ZS5LQk6RWz8fa8J417DmT0giP/0N8
W63Gm/8ihg8rww0gfjgX1QzLaNX1W0xLQrK1Z1D5AE77axeLtpzy2vGbtXhYan2D
PqpBHfboBU5WoGIu6Gy+JhujYEs+CLt7RkJHPnVWehHVPwNeshyS6+A8dDSF0InS
VEhrFtsW5/2bD9nGphmRo0Td3cdb9dzwJ4pc685uyY+Y72Wqk3NCN0vr4DyAOkkv
FkF1TpjgsSuSBVr5skhDgYrvu7ULnlsJsfnDUFGw3wkMhgRokGU4grdjRDEReieC
w264alRz5UxFfnMsS/ZiBYXp1lAA0tbdLCQod7SO3Qs5mLvJSzoG/GRlEx0Se8fQ
637pcKs3IM+5jYs3snNsrvrrhcZaiOD5X6AGZrli1gjmy7UImvtoyPfwfschPCBe
XxaCGZIv/hW/g+ORxgDp4ipOgdORaX9x1hj/cGSDKhUZpMYmoPGgep/od4zY2db4
CusA4a/LtCX6ZT2NJhQzanyXzQ4H/3H531BMluerx51n5LlhXWPiPujeTdH3PysY
2pO1GAF9Gj02q1AuZYtq0EKbzvP30J9SMGjwylDOvUjxOE/RkCYiyTo6qa97cfgO
agMNNMa6Wu8N4tQGlRKN8qVMto37ZUj37PCj0MwmvdVZCgBPwGe7AVsa2dc3vBRw
TyqtGPs8NOD8dZ7ThVBvaqfX0SkTxCplZ1wNXNEH6qgpEeWraiaXd6afCepsesIf
+ZbM1zT65qeo+kzdsiD7gaVtdXJLPigVTRJx4gt7i1Zs2pK4SeZizZFzKQZURNik
E64kviCd5Z0RJczF7iftfYiXxeWutfGZH+OuTZFGxzUeIUiD1HWh1WtqY6Pswy8Y
GWc9V11vQSVGzUniIbNJcvjTsy7BB9UNFkq6zkRkLvJvPWluxJLX0q1wGT8TXSh7
77KWBQ1PB56NLXpbQh8bDj590SAHObmsGfkBQuFI9KnqyqI96eC2mDrN9/S8va2S
3dJJxVYOxwtN37eTv698uiAGsxIXSQCQbdwYerhFdnlRmD0pBi+2YyzYJOG9hUhk
/rUDwjAg1+fs6Wjs++CQ2nv/KlS8fON1+IYNZuDMm/QQMr2Ee08osVWhoduPdb9s
0UvB+t2xc1YmVCuzivnLXG3jc3IggNWYq+bV0R6C6LmHtE9IgfCW5ig0sxR8+qtg
hDcey9CK+a/sXf4ith6OzgnXEgdu3JYwOQxGYXERjnPYdBGtiOoZNMlbHE1vypyV
WlFSO8xhiuuQn1/Ag7SoBxKWfQ4nJ1KjfYzalUTesV2f78Q8g8X/LsBSM9AZmZrM
KaSK1iwMKcmHo+0XxtvOtWQIugiP0ZElQV4wTUr9x5tmBQH7BtvfaK4emrQWX3z1
Sv/bpC3RNIfs8+V8oqKjQQeN/zT0KMeKHu9AvBFLCwIrGDpql1m5Zla6Bdu8aaqh
/7kimhO/EG4sXK+i2bLH+ioayeHBoCqZRqrv/O0cEEgwc0ws4wF4CXl9qyfczxGx
nOf6u+wUf5gL3cQA4OxrRDDiC8LjWAZ3sorsjTlOZ7zWDQo8DZ4RKG6CWfWAVBWq
+SKXmx2AbNgcwRuaPSfPFJ+gsnkfUp9nNJO21A1OHpyF3OK7Q2qcSv1TSYOUgQgh
gl05urg2+2+e8utc2lCaIjyyIVYElkQnY5BoMJiQ7fsIHi/LFkrOAJyifNQyXNqe
vGO5HYo8JO+mxYSJyZ1esjwYxRrclGb9I6wjKohDLDIYZN2YOm+L2GWSPUu9yOmU
QRIpEXbnWgdpAmXK43UdLAjQR385Wso9V7F6caeIS3tL5Fy7BLCrXZ8cEDBbsG7O
72W0+FDk2JPRMFyp96rmu8Ap/oySsrn6lZ/qtu62tPlY1txCHRcGv6vNwhA2Lmux
iBLhiY24TYZqdCEsfltAOXVzCMcr3C7cwjuCKXdamLonhYETGbJQhy086nfHZfko
L/qrhvPkgQFk/cafZdZTIrjco8364pR27WaNfj5HLOeRJnZUts0ZRJ8xxKHkYKB0
5oWR8Ir3d+Es/vGFkjPBDXREbMsa8xLmTH+X5/d2v9C4iIaPLFq20VTQYF1DX/Pe
ZIuNA8ad80UsXSjZ3d/suvNbyFAO9/1rEkYdqbSENt4xnk2/4q36G4rlhZLe3knb
TmsRV6fRabQjgTIOQx9mbZowxO8xS6YHJYTM6LaGxF2VmaAwGj5hSvyJOXQIT+X2
JTc77MSmkj3OwxJ/9pXNQfNrlXwWAVXbCM5BSQulkrj0R+/+qgZ2Z7hM27xdlyBA
IfRLLrcsiox+6nFIPm3X6RWD/b+xXu1A8dGwHvdeCFMjZ/QQCTtrwS0e+P0JzPmQ
QXjqwv3hmIlnDdUNXmtC6YxtcJbIL9fCDZwh9bXmv4WyHHtKwRRQB1XfU+hinT3v
w5On/6vuyVsHqpAYttTKQZLWtq5EX79G/f/DZp4U0SX0g6D5QgItntZTYG5ByC1l
sKEZ/olN917fUVGS6nSxxbknUdBpGhAyLsqkb1GsYtwqp9RBQgRuh7g+xtleT6pA
daZTA4gk1Aqw9hMj5JPw01xF3l64QAeQj4j4w4zulfx8y9A6tGoPJZc+uQnUNubD
QKd86Ko92wPqdvmaBlTT2MnIrKmLXuFR3HCqUGjBAlhOAlUZUj9yspvstXr+DYWS
yk47OAHtQhUYfkqXGNd0Xiw4k6rBO1yeDsS6GkFhyh1iE1y7NZb2kdTfjwXOkgwK
R2ZnpNkB6IfanD/PgmWDYIvrmwX/PL3nNSicUKSeCGktfChhY0P5d5wK3wl5p2/N
H0pghTatF71jE+N8xaAtxadIoOEMU/5uQZ2MkuWaeD2snN8VUMI/jROAU4OeQXBE
Thcs3ydqPuF4yNDaL6GPbI9XR0NjDfmwb1miw6+rwoZSlxLObC19aRJjw0ATKCFr
pQxGLwZTwgd1vg6cBzj+9Gs1kYa8J8kym9A4lBEFAp0mSi6GRDxwV3XasmKsXH5S
1lfonl2Sb+9nODsTaiWr9yclGcY4y9tVo+93TkkCsnUsVQbgSxCoPAQ2NHvyIXGW
gvo6DTm2yAyNZZuUorrJz16ZgqoMOwCfPDhCRoJ53LI8hIEFDvjGlHIXo/PQmpHv
M4UxlH+gcMDK7aX4QZDVFE3Um5krqwegqw+bqCf2+MQd1rrAs6QJ8vLhJ3C0YKuE
bt1IN6M49frmx3vcbOSO+xC213GyfWS+vB0RSCR6QPUwWGdLaXyLVGFsWepTYV9q
2txnhJS0O8YCYdoIsFm/BdUgKNKh4Oj5GepiJ4PoCbH0D05HQem92tLloY1YZA+I
DV41l+Rrc+iCpHUI2g44MlxupVii36aFAL2RZsJOEVP/oz7tCfFGRh7vRoo1UdZW
lpI7BJiNaAZiZKg4tR2PIS4ddaTG1g4rh+uAYVqx30+U0ttXjqXRC4Pg9cbKf3xA
0opb7WOS4vqq0tm6EOvwCTf/70w9I6Gn8E1+HcmgoNlTDX4hBk4poYScdfLtTurJ
SEqmlbrVHKmVjIRC10QMqu89cr7iocqQXB1D/lRUvy2VGlvXqtQUQavmGblQ/bcf
UZVlQ2Rv2yGH8IZ0UGspJn3NgQWixIVMrGt7R63Pe9NAXm97sZnm0MbaItaMYm69
o8DbpWhYrj7Be0Fb2E3XD0kJZd68k/Hb0eNu39LIB+KQr5HfgMVJy7GuJBePwB8X
+i7DS62kU8YTHUQpJeIIyLAz2gEt7lGxwsQI09hkOkdaEVsEzObN8Ylq3deHmpTW
5KZxK5vNTgeQKZBW3VDxMsTa2Iq+ydxMhGf2L77i1i4BXZueXpi/IU1e2R6/j60I
e+iCOH4HX/chCNavzdY7u9TWxZNfAmOXioC5NpBIU1KMOxfT1F5REZBI3FMgVUyr
B0OlKqirNrWT1WeHdGrhIUj0cxepTywoihzPRwfdN7LacmrMqQ1vyXPsRdOdGpOp
AHXPhM7rLJFrehBtMyZ0apWZj8WMJ/dp3NszWD5CJaHF2acdzuPWjJtnUOeJVlSq
b4ZAisZ/rjFD4+yhYyr5Aziu/iwbcT8PMi1t1BVn4VFfi06fpLgryM+efYNZd7Ls
hOsrZ61hH6/1E4H9+tyRvRM4+XmKSK5e1M3Dj9Km/OiNJlkaH2mR4yodNbgKc91u
c/mxw0e5ysOjqqBSQ0TXNoOYoLavIZl4BlsolLB1U75CIOV6EzT7dqNoKYnYBJuW
ZTQd2OzcWWaSbPEvYhC6YtGm/nvkD/ZCsO8zIhi0NfJ++p+I9gc/wp8+3Qi3GfMA
IyuwfVE8HKQsrbZ+e4td00j9UOXIAUb1ItjGlNMgWU49hSQfuucOK2Idopp2Cgt8
hmeEI3rhU24VsKiuNFLphBFojO4UPP4UforJ7HUMcH0gjH2/I4KlJYUJpwVKh/O5
jHYUaFFRG0joDbZt/+j2NStf9jEugi24DViwLns0dIAEN2ypbK/Z1qaKZ8jKXeKw
U/QC7nCsC/PYxw7hugQNNuK3wdqAutmeMZPHrN8z8y9akpGNU324UKTKV82cJ1hF
sQPs60/GHknlgx9ZIgQi0f4SXux5TW30APgqRpSO9OfIJMhvaC9vZIhY/BjIPg1d
I9qE1r3b2jH0ssjj4K3mDhYXjiIwaP8Rckn624gi+5OfrPwGFhuwONoyu7Fzl1MT
7re1ILa6x1KHsVo9n3v66cEJQ9WNDMgJSQRROqgrgkzM645dPC8S1DuMO4M0TZUK
A+ipgyt0eOjjIN4BpDBsrpMJUcCZCvesQ/1n3gz5l/KeOZhCwc0DwewzUKlM2KKT
8LR6OGboNUz1AlB1Mr8GLgFHlq39JO0H+0rGp6EqFOTtDyETM+tNzEA3FGidX2+m
5eQZUHY+xDfspvANqrWwxr7vFuOPahYr7+NBqG1YY3gqSWM03Dq6SuMnnvpa6Ulq
69vN27g/xX5Di1GNUfxgteexRfkpLnKsmR/LqyRjdHhO+rnINfBH15teZp2hjVTI
IojVDDxkhxGAwEOte19eQfv6+AisuKkPlF6S7W77Fs5Ji5yoJeq+CrIHkvB0oNuK
9+D+sMZ1FhurqqlIp8G/XC6hNlYsfLA23qCPaS288+6Ug+TmibQsMieBt/nDsGnR
OJ++v6He/JJe5UxEiCjvlofKdr3/duQovxQMpmi3fitECnWveNWyuii0ZTSiik/H
olGNapDrAPpnr0q+fDkxC/hFaPoD8MR2VHuInx/AmjMmgaB6cdc2DbPTniQrlikJ
c6qBzfuIVSKX58XtjrCOUL1oeLMQHk+cl7y2LSma80bxNywKLuze9juK+MhpBYRm
HJafSt9EuB23whuZRkSkn7QS4tYPBbcb70EBNbz2w/BJ9WrgCxMctvZuko+LMwms
FXrh04eZlEkzS8XLr6OEuA17fXaYeg30G5hWb4EAWxXGRV4Z0qi+OH6lgiU1cNm/
JXm9GQp9yK9HXgFvutIsJZGpD6LV864tEUXqYlsPqq0jB1RfGhpP5xw5mCDt9E9L
tGrVawzDtTK/H5e2Kk+Q/cA9tFqHrLXSo0F7j6ml0GVJWuQDGJlExhg6Wnql28Ya
w9dVBvPxOQtoQ0uYm56F/DNKqBUL8y/mT/CZgADQ7FuSfpMh9Vc2K/EYCS0EhXmB
IWTTDUGX0f2WyR+FBnGIwGjpihmBggz40su8Y4OPZhdGVOWrUdicE2Bx4EPJWJ+P
s3iFQa8jBZDq27CZ5GKkQG4xhhzFDP05v0h9iS3Rv2clfDF3sOOlYzfbFNLyNHXk
LhYXNfcMooIqbedbT2KtkIIMRXAXlnwHT2cuh2bkEiPWXb45QkpDoN8mvArc4HLD
mtUMs56R+bmU+vTth3PoGb3pZsqcRHkhdagWxfbky43PG4b8hsQQjFSkJfNqVKVR
CAIaMQBF2pjc/1RV6ZEsTdDTocy1lXTgm3kVdYVk7anO+QLKPcCW0qq4ZRNIwWnv
e1TqGe0ma02FUuGHl9i0iTUC4Sji93cj1D253j23/VAjgmJvSbZ36Wf2Kg1HmUdU
QDUZn6o7xD5fyxXO+GWsTvxuXnBhgAIPFdxnHRvMP0AGt8Ov04oEcSqP2/vla6Ru
II4gaV4wM28YjODnwi9XaQeGhyOufijzc5eEJyXmBCuaTI5k8rEIIDm1fo/Ge9Pm
enGDzN/BPK1n/fqInOMuX4cwbRaWKcm5SJcnYCgbjJaxD2tKxxlK/kVW4ssrL6kX
r2YyKQ7P3/t+3kzfIE7y+9oxy/Bi65ddYqiaGsLi6/UfESgwmLlNDcylXMUfmu/m
ahAkj83Fu1Kv+5XH+z9a08mNX6HwaJEuBB6Bs+CKBuFBtXb5m+sEv2mpfz5c8BjC
EMqGtJQByBlYdV2NnJGOm349EAGxpvKes/DqKL1jtfQBCyWfQfv5VBDutXWjDeEF
Bo0HkpDbg+zHtGFhegx0v/T2l56kGluK0jj0LFbKrP/L14Ssn7kkVWhCM2zlqFZR
yRpL7itTQ3Czh6wT8hAX55emN2qV1X+THfs/xa/dlS8Y7BCap45bZm2cuCWt/6Ca
d7UjbOPivmbUOR4eZYyYjnk6QPGWHURus3zmI9RyaDaArB3olyTd5BJG+kFJiyua
jbFtM2KVShcDZzdKEYIznSzGN56HkIgSJfvetj7m5MtIbPoK6ybcbuApYdetyOFm
6BEUhsfE0PGfdFOkyZigizXyvEQSKg+JmbdotajDRk/xYRk5lAtLJ25ZOkDRBIVj
74mHZ+6LDV4u7IdynPFVfAo2GVJiSqmMZmRL+kmtjn+X2exohCvxi2f6nrhf2IRm
NDg3NX+gkeNm9D3E2+3Ga6XNhzDSAEIjnlKRUBWwXqYVoRyOJLQS0JvN+1FN7llZ
sFJzmU43wV0IRxejRDqtqmZPIcbYr82a+OW722H57R1BUjGKR0+11/vjwoPheppo
T4I2GvP0a4mizmR5Kb6xFvmuDYKzxg/iRhrVK9w35ptU/C4eoV77vz90ku3YHoZe
0ys/jXSMljYmZfyRGqIPo5Gwrk23/jaArRcqfvaDQ8PsQCl2qMBBfqVdDIKfvQ38
prIHQzqKojizUFKs+a3fyS7fZT2zGYDlM/bMfOFzj8eR4z1ervYyp4Ay4A5Vjqvm
clCNyJfjbVkfscBuicZCwg5WwE3bUzJN0kbm6Ma5Sap9QwV3NniBiWARC+r6OHp5
1iMFubiVka5fWGG4xCwx6BaxHsH5WU6/3d0IYsA7mX4fn36k7cjvav8ULmzBGhfj
in/FdRzDzq9vWN2zegkbjVdcoYueNWVJZGC1ADAqFh8UHRl+Tb0AsjkX+g2ZOaQM
tm+78xRoVUM9cHq714mEoFPAhCbvCHOJZQe23SsFWT/BtloVBdnE6o3DHawYWuYE
Rvu8KgVfxWWKeL251HIFbKdYDK7OyW3GqXjAgG/0SxdErSaC9CaptLug5xwN80rL
wFeGSmgW04DjtMLCecnz1Is34nk6UD/4XXFpOmDavgCoj+bwTZvH12d3Ci+purV7
QK6ZfHi/yxlpSXXWcF576lSvxZTjVs/ZPjkN/II2Y6QdLllROK9tzEa2ymrOl2Ql
Rj2onVnXH5gE/LGjyTCSiQ1ZJ4O2dLedIFrjFQ1YdadtUAWWh8k4bu2Z9iD5EFvg
D3pVQIm6VdCkwFiYP6UFCqQKhSaqh4Giq55H0oBcFUWZR6MwYB338yE9RVV/Qndk
KCxJ92EzRlLn3sGVOtNc6XjL6EeSYR6gl9+GJ952IOX4XDxTzal4QQ8zms1VgdQH
89FPOA837P/ij+xQO6Py8Bf9qiNDFBe3mhMVlHv2guHadmAmoTgD9YhCIcpEm6Bp
HVGBwgha2Q9EFTR5VT9Orhx8G7+B27b4tXs7dfK7SK+xWDp1Qf4G4iudjL8jz1f/
e816wFowHD93Lc3kC7In2hN6pOEKtHYZ+siTkFemdUbXEr1x73Xi4NTvq8MTDWOT
01ZbblxGFabyz4hmv9mCroM5dSQvjbt7uSKI4f8BECg4lM0VdIJBzDDOgtlm88he
iwyztSmFbLLM7EYxyZYz0469rXfeNgm15WZ6QSCNompptim5zGSjc1Y+S35tIddW
8PakD/FxLA7h9wrjH9LUt4ub7J25e45GoF/SghPJ/uFYKgKhCrCpR2Pm8MP4Ga5J
fHFy+XfcnN7/GPT4LAXAlbnnR0NS35tQeQjNLgI71Q5SnmVLLNrshXLv0q2aiHKo
5G0V3EH09ZL8dr3l7QzJEHcKFPm9tIr6WAQJdV9lVsRGYp3eUEs6YNhxFAYlNBzG
KvocYc3pI8+69mSCCrbpskpW09Mpo2035wK++V9pNzGkdYp3w1GGNOiRDlrobh+P
ChqkcWqkmnCNoitBHXU6JlWyIQI4PVGOUb6pahrVBF7iS94O7LD26lE9g57982Yd
V4ny0Mfkn6otYsBSef5NtZnhOKtHld+NjyfCqKeURZFZ+HKIeYu+tYvRbdHasXk6
DVJcLl7SdNnwiW/3ST1kgho+T8EQsoC9wnVH7v2qxJ/vDyf4aT8MJVpqaGbCFz8f
YLt4u5JlZvNH46k6qrtx87a6AetYQ7EsgJGWZjv9eXyTkTfHIuWUh3eGqrksDqCc
uHmFrHgS25Hy7zyAqofU8qBIZB8jD4V2OlB87FbwajFnBzl4orOk8wwcn16wcWUm
W9bZ5p2znimkVZ6tIo5/RpXn3r56RjLVE9oos5jDHy5WSI6ls90xKux81Ek05EV4
VEg3ItT4jGjFFZRLih+4xRPW9CcrIyVMX5swlwIcO4Tbj/5x+mWye15p3rMoJpkh
CrMPUc4/iNi2cDm4ACly4jpINxtVlhoyqHr+f8VVlsy4+UsgMWDBY9fxEqhl5CP+
EU4zsqCL8RaYmIDvm/c6RNViCCe/a/JO5Zt0704x/BdbllO86Z0dTlqGKzLiqnkc
3w7WiV4RpAxhegahoRhrx5xHLHxLXmzkaPb10s0p+sFmX3AMSSV/jYx7vwwTsZIM
5/lEcC0cEOyVFwRSIXsmdGeCTlCfeTCCRdotTpJgUbjsqY2imq+pGAhKVRq6KZkT
QNtwPmFHzuzkIqvR0P39X6/AQiXB7M0zj3wYADRNF0rLqUWP7c8e1XzW20Y9mCjs
op+1AGo7JbTlZ8YV02mTeKidtwRULNL6uMNC+FW/46G08VXRFDNBPqPpLlfKAn1l
IRmId4Bt5vwURV+ZXYkCsQD3jT9JAIMmT4snrZfySeQgIytAAxIWPOEyCnxt9Izz
JHg7k0eBTmkjeeegZl3SnkVMRwUdpNoGxuZSDdZn4/3bEWmvqvWBr212sNFjDHdx
NzvDbD6Wep3+d4tsHnmmK7XJCzPWb0GDaRej+7yIo9o7sh5LLqdsG8XCLYO5gBq5
euqs71mUi9bPXB0o226hfoc/B96RdINKWjZmAw3eE0pokItlhe1D1jnWthsEtz/M
m5KR80OdUK7xfxTK4x2RCaztZ3vQYGAcW6gD1+NgV9ynKGPPHjE4oILcm2oF2yzk
l7k5aesqerAXEBUgs9tA5K+YNJVsTT9THvTWK/itf6bZ0i4U7yKi+mb/FgW6n3qm
pNr95d/IP8YzYO5PPvuQ1uq62lTk//dWivmDMo7KxyosZE75sT2DtGIxtcGZWF0/
O8cRHXmUxRtHjrDIHqMrB8oXU0eYUkUKxN9ypzFOOoOU3M5rab14DaR/5Ix7BlOS
nkHuYooBHX2l7jVJTLj9ZfA12vBhq3/98gOp+zhsIzAgNPdgm30zKOIS/LlewCpp
+pIiduNiS+1ww31v+OpnZXZphiSTSBbF6e4LxZQZFHS/QIhNtxTyHmZEOieBuTRT
4h3pZkma/ojRHk/6KsdUfPjapQ+YF8/6wwSBImIqqRL+atOvPq4p8QKd1FideZHv
TgPLE/rShgHjLGmN0/RaxcwoJzWLrkbKUVeID23fwNjjSuKu0BArC9Ecc7PjpSMr
TQxsE9Fpvcw/obBZPd6BpbSlT/T1C/7h1fTZnWZ3fayAUP7Uf1vA8kQYufsDUpFK
Ze4xfjYK7C9+Eg8ijnXk5rR6dEVp6HsvbFPgPGmZiitg1C6yposP/q/mVzgbC+qS
q7M4Uv3P20BiOcv9J5QPHZ+XiP0zqAn3gbWYiS0kyaquRqMJCZwkKt0nCeeeMAh4
IRpyYfb+Scy+Xr5AUyacpyF5GX7gFXPF8UWOTE5wwZbO1Yq/vKtuPTXLuVZqORvz
a/+529hmFXee8PKYc6pjY9jftPHASctC6BSx/Zp/e6eOJKIctN1IQt5csw0eDeKc
+3Wto6JwUq/1R3xvSCf9fcuaKuiDStlCPpa4x5egfIeTDRzI5eAcHlJmFIiA9k5z
iexU1Q0Lni0DiEeq1SMdkjlHDaE5FtSHApYkaqq6K1YxjRhjW1tj45zczf7xboj1
sthAOUtYJ7Ox27xrz7DqAejBJKewOSgvym1agkhnuhKhx/5t5x1CCsZH8kieojBK
4dckUogk+3wr+ITlaKXKnBevrp97GA5hrIdl7lWXccwTMeNsLTA1XLx38v7PoL/p
9VKHiD21Ka4AWmUuZYvpYGHQyHJoGxxgoTGdqY7+OyzxzpW3B04MnL8lcG2AlaEn
vFFcArQ+3DQ3eUOd4JzEy8ny46twMtmIW0U/sfJbkIbCW/jdVDC+OzaWp6f+uGV9
zxIuDc+ir7yTw7Wy3I3WCBtiu9h/wuYZ/gHbvu2O8Ar5jhfeav6eQWj3bOBLK4VC
bVZMCp7vukQLPSOsmMMIRtdBTPO94KgvS4+QKYVAQyRbe1BWRhDUjB0ldlbXo4dA
L0HB+otzT6wqC1kJFY4HjmoDEVxj4JWg+7+EH8OZWmQmEznv4OI8n618zH8Z/ueJ
wm2tqiIf23e58l2ctNXmZYo5kczTEI86HCkpJtDylFT5ySimsmPJqd4vsonweMh7
SEXD7ojSaS5NmKjucxeo35C6XBmXne4dtwaUlfPlQlXaQsxJB0fJLOgn7ICAhHg7
uDgZMHne/Gp8fJs4o+uo7ddxl5bHAfCS7O6HwbVrCT/0BA9MSO5zm112R6tbLtBX
Hu827ZsJKtexfDZVCmpNsaChB+05kzs0D25IwxA3C07e+hC1TYlW1paLas4ODhPO
9HzScKlrLYjWsPEPoKS52iHl2zYcumW1GTmGTx77bkn/CL6h2gydlf5EC5TlXpgm
HqdGjNvVlkOEsrM5O4XKx7OF7hm83Bx5bdFPVvDS7RjZ79OUhfiJLfvt9ppesbU9
n9zH/EKEUU8cje+/G2pCyMSOsla8vxcodeeDarmYLXswTOS7PRD+mM6zXw+A48/d
BDlUBqxGXnYEOZQ4SSnAnCzySDyxJz/IF2goYAhXUmdp3wXWMJb1b03ZlJNPag62
eGtPmYzon4hbJWBVep8wbEkDC6o9jhdUgOr4lF2y+fDvxsj5XcJMXO3uheXLzhRv
TRoL2qJHkI2ViJH+YntaUYkdhYBSyQrzQFccLBk4WLpjzuex2Qy2TYR5qEryINkG
gKeGtpyWmWN4M8rwcdPkVIj8Z2Bhq+QEiX4OZYbpc6FAuSQJiQmt0l4gAtiG/2rM
d25XghpFs4niomnJx/GPvo2s/kK1s4pZ28jomeErV0WBS6EqDqYe77NBMSGHjL9R
cDzPFIYiW/YRBNfkoY+GUDjje0Y77o1vKzZ+51KznGWsauuCfa4XpXk5pgK6aDiC
H9j3P0ZzCgvZ5MttiyFs9YU8tucdNrsuAzTqaeFQwnITKWYMwXDSEYLbZpwxmShG
AZoehYjZ0e/7sHzNIfFtHCrge21zsvmxpIUEBhNtiGKZdm5pYq8GUnjXRL4YJuBb
NJJK6+4IORwQjUtdU8m0lgkQjmlycQwAj6hbu962pCfdrcDH7385xehmq/T22wSY
YPULGm0NNDeAVi/NPQwjYYGD3G539U3MbgQ0QaZ0vAle9Y+XsL2e2WyfzvtaW9pD
wY2bsh1NwAlP/REyKUCCzBUIcGTH/YigJPe7ylfCp5TBwZS43PAlgySFCe7zkLbo
p794FcouulsLCWdd9JiTzkuVBNoVJyK1TKWJo3qyDcYKY2Z9F9vdnNHcVDK18Qoq
luftOFNvn4OafJ4slC37PY90CNi4ByHM3PpBrokqrEY1BIzTwgvTpHN7rURREq3K
CjMkhpuiIogi/FpxZh/1F60MABHvViLNEiFF7+IcyTa8yu+RRqj5euEHqkukttHt
tzu1hLZVszMoPOaeLgYa90t6GZxGj8voXPO8lPYezNvfejrNLhLuIVKpoitqb09r
07HTu6uUNxrr6vIwjj+hbi0iiAczGU7ti/LH5QDajBBBFgjyoWqKdBkJmdAkfGA+
8SwwYzUIGvAsepXxoEB4tv1KJTj4wNTmtI7LlR2qr3hXeBuCeaXli79thnhOsL0/
uth65uDYgsKoK5vcCUrnrTO0eWCezHy+O6gKqWkCRSWnGJIHrR7CBvWxv4aNjfvN
OdOZFFeDJLYqIjI0f3iRsd43iuKGflSELJXa/b+wz6t4mbYl3ocjUiwC9DZi+AtA
xtJTtRCOnvli89DzVcOBWsjeFTYKMo8FpoSmV+ERdYmGcdILR8i8EAazL1K2Opkl
5jQl2oY2KwUmc28w+vMoH+HRKAAmIovO2pBetCLctzStTbDVXYsR4mLaii4229K/
1K5esuod9bT+ldxxbWp01xEka/fWf+XoueJRfH4gOjFUz+JRE7DGwcTT4uMh3S1w
R4ZrPjWT+IenzQbdEIT6iiOpfEN1zDnl59JK7uoPPmxJRvAhCGBgi6BCHMBT9Lnp
WPo6Fr8hA+LNvUGWKXV9f+DIJ3k910swCgmTeBz3WrHC5wlrOvrm0k6yAzyhh9G3
rfBOulOHSAgf6SL0skg834T0cyQ86q/KyX9D3eN7QtlmIo5GaNHo1KnX1rNBW4wb
F0YRcnh/UcPG0aIOtdv7XbraiUfWwd87RFItylBjVH8tlWPenyVa6qJzK6fr/06f
kK85wktUxdVKBBCAHxuzOl2tg3W80SNkfwVVEyN9DeWl5c7fp/+9vygv5GSnoT8O
mCZbIYwhvT5pRyQmA6fGV1YeGQ59/svKdExaAfDh5OAcZvnPQAiNKtdCNgREYm+1
tNWjRxIiEbkKxW2L2zSVWf3jhQrGrqraBnel2ZlCSbfdTmt22wq65/XVFqEvsoy5
56YeilhFnDFlbdl37DnNmi+0oraR8hf0djGEm2S5+rrV7LSepyUv40TKBKKQFTsk
z0XKtpH9nynp9QFN+raqVKMJ+7pBUSpSviMsxo87soSizytiLqsOt5JxhyzLPYsj
/MRUUR31FtWL8fCLjlvLQ+c5uiCGlbOMy+9liVkzKuMWu2+lNgLwiObcbAZIU6Jd
q/hpKUENKDw30h6NzjvlPccuLBt/BnhZJuVoWj85y3SYdSU6AWo8b7Pguaee5urp
Wol70qsFBvOAc+0I68E41q6Gcu7tijHMfSjtqrIPv+MxZScxxH7+aKGWogr2ZLmQ
0GPidaeg9CO4nW5lP+wit0jb02GGVZYUSGGpX/rSrAYSCsC1tqnSlofW/XNelkKm
FFuMAglbiMyFwDLD7KiTtMj+ovDJao6LfhxYJnRJHqT2aRjWdo/mFly1lK7N2N0+
U1UVRcYzod6NcqgMcsQ7BmvtYgXH86tM9OW3I5IRT4SuZWIx332uB5B/Y6ONRlpF
h9dP8R76ZtqDAFWFquw/rOGPbkSbPD2Ypl/nEAyj7hx1xfwzbMxG5hjTVJeZCQzG
+kKAGxcm+Mc5a2FaBqyXg1bvsv2x3B0j1MkvU64uuS4ghfAVAOKO4MYgEhGMf1RR
u6g3feZ4JtpDHdMnxZ1am6d8hn+iCHeTX3pXST6o15gCQ5cJkKK3AvQFuJn3BHO/
z1I47upfDyVsD74jcreE7drrn1y7F0Z51pJuCHML1gE8p+CO+D34eYYxzAGawPOp
RavVtN9IFwkvvnjqm7QuZyvbxxHa1f5XhbU+8Mkan5dWkJu2ozPcGhGAoTQSr/M/
6uG3N1Y4fmrEWkq8mFLIfkJakgvK8xmLwJBmW3yq1SaqQQoDXIkD0MN0J/NBpahy
S25H60HIu20oUA02sbfuK/QtPRSTze6IA4yaZ4T7JpF41Gr0I1ere7AQOG2LsQZS
HmqgBqZ8xOT8rT4+5eCFVVmYkQqTE+j17ak0X3OyNAdmUeguUZliDEYgrbaFHa+K
qwYjbA7vN1dMNCgsi3WatalgOgaidqnaxi4IPmlIeUDvzPd6NMmASsY1sHIalNpZ
yivAilXUwksyJzCgkArU6PLvL8hXlGAe99ixl1dsPW3KS+v+jZJNPxyXcDqq9amV
ocLXJUPEDbsCNz1khF3BWVrcBYEY4tjDJt1bqPHlkgVHRX6hv+9a+m6d8RiJPX+G
JkLZDPA9zv12X2pSV6lq8+dfUvTsTC6kmwXEYIb4n0c7mBye30GpgtD4xz5VBPTX
qWzIEgWw05MmZp9LkPVzLm23qHBxNreOFhrfHl1j1U0bDoI9Aerh+1v2x3HXvdMG
hd/aHGUaHl0zD4kmXePLaDvVVlAd3S0tcoqyGYVlP153fj75WYmuVutQMq2C+TSa
YHBehjGZbikmMgy2nPt4NKGEb7aDE6yxkyZcnpsCbb3LJngAPSIMlxSxDDjlz0fc
oV5e88fN47VXdR0lAKCejDnr38CcLQirQaka/BIqdkK90Yg04U9UgvwGrMOYPbGJ
7GqloiAhdz7KW77Z0qZL/JVPRiS3GjN3cRzldOu7NwdIzF7RzWwaYeXS9b32sr74
iMKDwCRxYImbIPUrhvAF/Qd2nhBY1+dlr7Yye20YvbXTlWJojksphTUtWG4TX9v3
MJuaQUbfBWgxEojwzmf0DjZRej7H7851Whx3XmcwHeXtyjNsydfcI8ubRVPEkcTG
BKwE3Kpl7guW73Ypg+uQxTd9wOAAZ52iM8we4oMc3CroLzTVMr83mAha/c1puHCX
mfod7Jz/bjQAx6HFWNru1FEDNjeg42GtsFZwL7gLdvgqIeist+DkqXFMIWb1rG4r
g4xtvZ4/9VigvDurOhHsA950SoMXf+JtfX1LV9QaybLr6fVbtsmySqaO8qOqu0d2
gRGpozSPOoC/UNCGl1n+r8g73QXPXGyVhopCOp2LWgg2q4Uz8QUH1mwgz/17f9su
MmYus1nv9lNzJQ57IUY3qULG/M6xDpdhWY9UtUo7VpQMG9Ryao6cPJIXHCod9Dss
qONubZqRyKPknau2IYdgKFk7XKJwlQNkvBlSo0a6m30kzo88axmhK4MxbPEakqS0
+qFMmQOyOYDsEf1H4mjpobkpymu9m4iPCOrFdJiTyB52sx6S5TfBorqGomVuc6LD
lZsWpGDmlx4qy/OPQCoijpTA8MwHatgSzEbm6bLehYx3UHOdxtvGMUDCUUq4qqQP
gij169Np34wio1JBQG+1zsEIzF7CVZSz3YQtMJh4fQN/8oUa0BC3+rF6KXznBXiu
JEDb98jGmDG1LY1+/INHOCJuJtKkcBaLPQoaF4jCe2XxwT8yNK8HE8e6aKO3e5Uk
LVkRB6Vfdeccw2BkC/2b3ZXGlRY2yUb53Mz/AXSxNJsQ8qwD537kzvb8sFWnndzT
qD5mawreL3Z0xdkTUUSTDfLhsYTO3FM5c/nNS0MT4capz2qo8/sd70ppXr17wExu
Gfssz2wdZdTMhxVFurv/N6QevmByuVxEBZxZYiKAoUCK2O9Acy4XvpgXKzX7q1x+
oyGM36XOi6+yupcn446R0C1slX/ywX2luYxv1LoEMnWRdhb4V/vaESKyfUVBGaqn
YqGoFjzoWwByTE8GtdVMpBlC9nZmY0YjgjwBlwX0aQ9mV0PpAUMUeEgjoVAxARNQ
zb66TzqEQ9Kmb0yxf/N68+pAeuTufJWlt4n932yOT8igWrkeBiU67YutwXGJdBjj
eoi9Houvh8TTeNW2JEvRoS8v9wjQG9jGozO8oveWmKbKZYoixEtXNWvayPJ5gpCP
a+QDmYwBCszw5la1shpRZte2SO3Fl7Byf8W+s5MhiB5WAcPZnHwweNi8ldd7IZV1
DvynNRVy6C2dQ+VhzFrloEWgc32zqPRwBL168dj6CNYWaXSAfWN1By5GGaWwPnbK
JjECJn9T7WhdkcmQMwCHA0tWNWA41/BbAopO2EZkFUZq3Pv1N3OGDxF8s2zqFwca
95r6hWVdNP+OgdpDjjF91FTIeC7vjlRmYGmx5yH9GEjakbB92jErCBraoRDkBgq1
d3nlV56xo3avdEBQINiOG0Tblz+SR5JkFxFqg0Wnk4ok7K0oXwaWusaFMmStBv16
XOaJVKBxMo8bprKMgzDQzgeWHtaFzDIuLoxkS7E4i8Q3228OfHTWcJMOdORDTg8c
3UHnpdrUDRxKVQE0jTc8/VSf3ojUmH+ow3mkRJ1MYEh4hVGwJHz5sVeXXccZAFiE
CBApVI8nh6rM/2T9GeevmK573o3OUhjBns45LJmIFqcNVCuX+8KGX5piNZuw2G3+
TRFgBPwuPDOhuRHlTnviI4l8wGnSZ36q6jMwToneeQaVqRdoFE++i0q6ZQC92R4s
JSFSLBAJcMQpP9NYG/njKVLHSRDk0Nf8macUM8ZGBi8ZBoTLCsJXtxLTUeM8sgiX
SWUT729nrRrp2ZdsEftRuzx0L6+71oVTL+qBuooQ3o89f7YbumXTsPt2ZjK1RBRY
QFVgv7FO0iFuNbwpV9MQYZlOvvqj3AaBG6FHcqQBhp3xSkxIHV/YIqK2TgafDH40
RdIZk6LYPlX5Jh7+OICbvJ1yWyhxJJ57a/ce8LmWlN5VN0NPkn9wI9W41Mfyb6D6
nRczs3HlRONj1aXAWBqyuswKF05huzdc83qxk5dt6PCqINmj7+ytm119Vch/64Nf
7H5z+Wqyv7LpvjbHQo7XLOyaSy6wW+h+bFaqdLLA1+ZBj9R+FpNO6JB1wo7o3vL5
Zm4ui8h3pycBIyMLmv/yH0v3WqHUmKYYSUPA9sWFtbL1AmzZ3z9DFgbVfNTzYRc+
RmQpKVMpSOiaGXnLH2oAVYUWzl9mZSalGku2L1vfXtKpTs0vshZ0LXv8fFm0Apnn
PPfTQsNo39XJ0vjHQ75qnPCMfnWy8oH3xiZ8hawQq/fbemz29OMMnd89BOuCyUC7
VYDwzLTmrLrtT0eQHWS2R1RrkReW83+bKCRkkOiNePobVK4JVNu1nr+GZpYWBZUo
f8f4jbUEqSsrjrlHPzLz8MGszrKpM+ITDjsdFmTRTzYbpVENQSbzWwztWgj8z07G
AQT4clhCeSVd/a0xmyHceC3A2l/pv30wC6k9nXkJvlu5LmGiQa07GLNumi4AqyhU
dvILPmX8bp1pQX8UgXt3wvlvnhecx5Pdmk5rGTf65ayda5vNhgGz9lajx4ieEgCy
+3Qsd9gQPiLzc+SwOiZpE6W5HMTBfqKxQQmAHH1Xw5GXQOy9d+KFRZ7dpVqHoXjI
WkvaVnFkn4/g030cLAZSUpc2xv28oA4k7A7Lh0h01UzkGf6JAvE9fo+VL+Dvqs9q
kVqOEmzhMH3N0NE/W3ZmM2nIJlIwcAYGCrrWJEy780nFw9AbEQAOiGdTAyul3RdA
KrvuSUTGI9lnptefOxeM3Sf0Udk63+cbv3lag5keZURtxLIwGRktF4sAva8ITMav
HW0s5rLeRwLxmrGSw9gbUnOSypUs5ZogCIIrunKxEwfUuI9DnoApzby/tWFHlmmm
0ejv/z7USvK4pG0X2ZEsZKFOlTiiWe7N2MOj/uglVDsYzT18wT/xiFVxtC5X7DKC
1TfmNrq0h5MRj7XbI6MpbP1hqKcxaIBf3frG0eQdo0/MnbdBeLI92bohUPspdAtF
vr7Ex/UvcFMJ6HcguQKwHF/pTqHyK1iBbu1kLChTmxKJhJ74kDeTvK1tznVeCfwI
FWs8sP714KVz7eHvakJ2FR4QDGvb3X6BABP/AVZ5qymn/od6w9Iligbq2BMpDxMl
r193dfBYc1fo0ln/aYmrh/12wxldpDmHnV31rKklBGmFXRJDk6l/O9IOIstZuSTy
vIbzagZ2BKEZMV6NfYht0CQIjgdrPTTv9dvFJkXoK3cVcJJ1q4WzYOBjmakJjHao
LCBQyCBPuEAG9fru1sz2n8b+p51a5UvJCYfYcZLxn7FUySOpfW8+718tTXtsbT8v
7RZ58+QS9/2S68EF8saoWXwP902pHEu/UuyRhixNA0ub4Gn8bb4sxbg8cHmnksmx
+qVRTWKjJzDAFecz6MVEXosiYKM0vJA7pHwLEdngauQ6TZYyYS1Lg4G411yzlKHV
x9HSSaT8TNEpAHwzdgWWlNzhG2R8LJb1EoJsSoLo8RkgbR+YPLxuAUhz+kidbndE
hsG/4AobeFBfak8UpckFoUCXpgm/b9rBWoYr4HKGbWskZs98bLDUx1RaehM6Iq6n
1r7m5mi2ib3sBnSTCZbJLTeQiGhKJ2YgkIkBpvPdgwyvI71RcLINYpP1Kwo/2/tA
mpa5WRDhk5qrYpqVlJLZJ2KWvcJVrzjnVep2TSvpRiaZO6WRnibXtZAY0Yw9gAk1
UTaDlSHQxsOBUZDh+MuOLLmDd9ieTEheoidg/1yeRp2gKzQ9okW6u+H8xMuXBqP6
KfBQkvCU+LNbmYpHfG0aCS5ymRMCnBkeoDWYw0mJeg3JuW/wf3PrOaDKY/euUyjg
fS95ZnSK/CUhKCXllWYbPOh/uTsCyPPxZ2tWG/omOKoFrJ51Us8DA7TAWb7l5NMq
gr5gJWjo4VTWck0abuce6uea1nSBHLuF+CwK8tR2eb32Fmx6PfYVdhR0Qs92Ustr
2UIWqBeMYzhTuVGR6nm/9Ck76oJsQi0oNid/9wu90GNuxmanMJ0e62w9JbH8NZuj
9ttrvir4dqLq5viY5esa/11F+I2ASOPM3TO+MzoEsNWZBFm3iZRLlwLPQUPnOvk8
jyewmNmY0Sju2bsd57PakJsmM4bqVxGbBz88BPTdAt2nLV/A2TMWCeCbKdwlSe+C
HxJcj0w6SmaW9Rgs42lMg8fHlGGDjdoAs5Cda/N3gBFd3aM4wiafrnRRDpWcBNwX
sc3QH/znHM3cOO57rC6uva9HzEO5ewH1U3MAnHVIlaaaeNY3qfKAMrOuV11iKA4E
pqVWusJTM5VZj7Q0cSBz+RqDzkWmnFc+Zonug1sI/87U5DQbM888x07ZSJs5bZdM
1BB/fLCz7G/LF0eBI1WWzdnkjoZcFFaTNnmnUJQgrUxej1xJNOGeFpJYMMS0U/X9
VIucoT5de/eyX4L6JSZv0LgrgSTbF9F6tNIvUn2pS70SjzJrd9zDbBmSaDw18UO5
jllFxkjz/d2eAwu2doycygGumennRVIFuv19ugQJshBv2/gB6FuZiKBkqhmtdUA6
HsmJKwNkqZZN++GIuDIA1aVeAXj6PTFdelVEFkiaM+iMcYHy3rOKh5UmW3rfk33s
8klj+aq8eyVjXyTGcuJguQWx3F5DNF/U2g/UoI4eFoE69Offxgjj0FpQMaBhnSj2
C6xM0npnHjrOnhGim0sd85Fw7lNkSM3zMycCQT3ObRMTz0Fllv4qIP/PByCf+HRj
Fnjn+UsKn0M2qsMDYlNKJIYdxBA4p7/qNgBg1cbuzOzb67g5w1a+1z9RqIhGb5+1
4iVM/FPOA+iKGhPK9IYMPuOk6TBHiv5S8VQhUgNb1IGfysAOGJFJn0hDdiGJnyyR
X8zI6pPlHhuYcNOkzyVieFSgSH7eAq8ANmD9teEa9M0ZDjUKWoDJ0bdsXv63YxY5
0SLj7oVh3G5q9M3GOtSCGMs9/DIPJY2Kj2VjC1bDHQEu5pYwAeYNVwKCQc4+R62g
WpZXsXVs3VliWY2sVbDrOuHBSn5SJyN4IsHqwRc0tXFHtzKnSJ1/EZzDSfeVv1vN
y/IA0vFL3v+LSVORkkJJFyu7691io1jljObv2X2NpI54u9vGpmOGbmghQhxmbdCN
oYHKGsacxOI20qvY5WMsPolaizfqN+sqtW2QJf4m0cyfDV2wctIJ4P9h28+DAvte
q6JRw12oqpB7Dkh4r6k2lcOWqKJVpmDBssaL8jamCQznZ4/8xau/8Mz2nQLfDl/E
dcM/1fLvIixVZUl4wDkdjDQD6w9Zxrq5sDujFNOoDHUymHPmVtXKoDKFtNGsQrMT
0/G5M6Kbpu+QGr+pG1YusOYo2mUeEw8lsic0eaATVyjp05b3s2WQLcmzcM8bhhd6
j1ZNIGOR+m9xNUQvN/oj/GPNK4qwhw1aixCh8h44pNPNX9xMgyYiu1uIpTS4KNPx
Y9zfT5lF8plSzJoz2x0ZALJWxct/RQCfH/avigXra87kHU5aMD6tGUsmkxaF3mLh
5KWFDFpNERzS3jWjryRKzF0xmqPfKH9B3NbritC0uFrAeMVfBUX5UE7p+zzXaaGu
b00dHPbYookbqZVscQDI3C1jGFJU9DP74X07ZpDXQgbs4mhliY0U61Hr4VFoQ0ye
UTEmc5qQIIO0S/oi0B1boKVd0GGiTztQa6okvFCGIeCOSXJ2J0U1+oFj19nzXmZV
2z6jrcPbljnNHbxkRfvVwvlNR9dYXnxYQgTIPEZeRpbgSuT0HlmOM3+ZQyBh4lbf
mQJRmF9JF3+8zdh9jCAGC6+KsA/5wmPFf6RPqNljjh34kOL7oa334osQOrTAd/Yq
EdtBL425eVyqfLnXPP+31ET5901sR9cfcwL7Jl8+NqJWnXlwqerNRzRVpk0h+PMm
6JNHhInaeZHZ7gtcLr9eXGlJUrhMBGAGZ3dc20YxWZozVEYf7OYYGOAeR8qRi6Os
lEIZ5qXS5Pp3oE13Sbg+KGiROSNrgOk9NKFXk8HQf1Z+1aho5H9JSljst2YuJHkD
/ElAb+cJqI3mHqVTkQMf6XFiuPxm4RGEDNOGGAR3+sMgognHG16U9XJxQNkUp3lR
WJbhI1oa0145rVS6+g1XotwaCF3e7Oc2wdT6mLDkJDUdhJJjd2N58O16zEuafoZd
mzHJDor0Jai2QxoRrlOHy2ZZ7+1iiGucXXvs8poJEOyT+RMthA6Hrt+mvVYWD3n1
+LW/IqcTQgUPotOTudWQ8YH/54rudYlZgFrh5D08XqaFOmLWUcY5c9mZoQUIko/U
cvEZGobyDuyLdZNRVahZv4ZIsVhuEjZQcpgLiq2rRNPFtbEvtV9a/AVAXC/CAnr6
1TrUfYTTSHngAyqur7HsOtDdeLW2xrj2o+52xmZuxo+Yq/tnOYImsXJvVwqlQjfM
JcyXTBICzn6eLdkwqM9OK/YCwKhmFoJMzv1iGKLLeuxXvz54IMgjyVdILCuokJq8
v+GkQVCGGlj0425J4T7/UEoicBbH/hzDzI4izSj1zho4CqVBcsCKZXs68AwqEdDa
1EvZqvESZfStEyFg10EWuCQKIk0KAUA6TwenxZ4fTFuzQ8i0HWnNZU8lH7pnPaIf
oDW1MaFEVyW5sDELP78ufAR8pNMbsTjo9bTR93hZP+zzN7hOjVz7RkBJU5ArIjQJ
IOHchAftMVbY2xtPVgNG3xw8ueltRw8Qbp8MTVGygcf0+T+GSWLRI63b4SeMHiig
fKehoIX7Ujoc80FzvnGg3GBGByYMdDIeqm5OwROWgks83w8C48CubATJhXHsLnJr
FAYuDMwByOkuoCp/s2fE/9qG4G1dDh6bMG2EIyb3wtrbqV3ijyl+sLVVM6SciD7f
cD1Zkrl3e0JQbN1cy7rlOsLBzu3zFSgxZghCKxWzFv7+1gYz7C/aOVz9Kd9xpyRV
b5bowSdgt50t3dPuUhVO9Mtr9krIa9H+O6IThxSL/xPLfJ7eVW5pHD6Hcl6fFhVG
iu7l2jEFHwkgEOXqvaGqGe+yuA70u85rK5LGthaQLUlakPVha2DdOAmc26NwQOXL
+AMADzoWs4UZb2DzADH70VeB0lT7j0ODaqgmL6tKsumHr4YQgk3UbyDK5iP66ugh
dmxjF2jrCL+ppUN+Wlu9pZsTfcCyR0Dwe5uU1YaEB4UvxjEP3FBKuY45IE8Zfn/a
uXKCvyIbt2zTr+gQ6VN4M+HBsAn3vgPWan4cSTRLL43aqFEwyZOr5HtUCuhH6cRP
xCOv7bRizkwRhVMbCkMq0EpdcKf3X60mJngNwQmLFjG2bGdOnVBJNW6TEBRWC8lG
LHwlwSY+Wwmf8/IGhJR9EwC2xqQJijX/ooRjzEMYVhlFVZGXeWpSHaO3ctnLZ6fc
zekgQeWhpiGEUwDGj/mC04aEbEZksco1hyxUX53yOhfAotkGT5EJfdDiMs2ffMug
iNI7rParWYQ44Dny2bUiGtmdu+MItTwM/FHHj8wJf2AaHkYwZkf5ai3pH2BfSjfU
CbdN2tbTRHKfKQRfXXdjFEdwQS6l6hQavJM4gvo2bLhNrchPS9nA1mRoIJtYOicB
B2Hhnh5u5bQn04hx3HS/dXeEUkcA+bC6zXAi/zjRUJRsHTrp43elIo3Dfu1fCRMI
L3rydCjx+1k9vtJl1fzivtJo1vrRdUY+Sunl44KCo1NQySg2B7AeCYY2lS4s4flr
1MTWlwMaThxTadwvjuf6cve3kwfoFJKJr5ikWrV7gk1qAiPD0kmUsXWPOY4W3NGG
mmBktVS9PZWRaLgSej8qapoKXPSvepSrF6B5x/pVIsp5zn1qcBPLTlecjqJzoWvI
GyvC3N8ELpQ2J6cOrZZP+1iZtOuuWk9uBTL1VnJtSpgMLMUJxyjRZnJK8IvZK69D
XIo7CWTT2voVxML8RmOjhYGxEzhq0pu66ANgO+O0hlwAjYgYUgSv6EMjQH1FroOD
tTZYGuOpOcwXoLttBSU6iLQFjod4JhDPHXhg59LypwAcYGznPbxVsuR294iRSPyg
tOVXYnjCPnvj1SVlLeTRY5opUfhW90UBBxkLuFnQRjFudwY4+Dx50WBWKRcMXj8v
0lrMjV7twUdW0B/r9OxQ8j3hsxOgpkc2k/eTPCm4N3t1k+IL8xWaUHAyk8vRoQwr
d0WumhV+82WLWxrHEx8wtaGDicTGxSl9uVwFa1rHQlyRv0LLn+PZEgxsa1LDL0b0
ed/x6+VRgQSrpziLckjbVe7glemgqKLCYUN1GuMCGFReGM86XWi5b2h7C9a8ZFux
pW9ZCfnr+n+nrTHWOP7z96L8LRJe6KChNVneFR4yYsUANvV/JNEwHwGXy/pT1YI0
QQU1lQPZ66RkLQFeQ6nII7CSmaT0l2xB8WWbsYSdHf8WBq+pi7OTln2+EDNscLBC
sip+BsJvHZybf59rCb1ofPgATtJ5vzWUNb8g0GWvEmVro8jaCe7NJGRBNRcqEsR3
vN2IHf3/x7hOkVSjAMUnTgBfcmTOeYOsx0ieQhW3ZkDZCG0wukEPwCtH4v8Tz117
Z/ohUgWzxcQryQxoFAKGJXX57ZwcCvk4+/UCo0o7tHO9HRH84ukd/IRpTujTbspD
BuPOvGrecX/MYLR7upMK1Y7FJowvw/4MqBIjMyBoB4wmKRYWzwyzj92BhZ1dLZLF
Si3Idm69czNvMQFIK1G7kS0KBbuNQqoFaCkvk+60Y30gAzsi2ZvBHWjyXQqTZKEU
GGXD5h/QgxRvwo2bYirqZf/xYnUyWbA8y5v3AikvN+yzkugaucIdC+s26CCnD0pM
Sy44nklZxv6hKn8EhT+daptH08ZFuINh/TvyxhF8T0q4yslFVp37ZJAHzdgff3//
TsP/jeVUvMuSH8apWJtX58gynpzQZY32/SUG+PxVzA/sDz+jICtxei6zB9kTSI9o
i8cPfJESmwa4ZfkRW3H9FpbvPvxuGhx73reGjFBXN3xhsFq74ewKSi4mMNpH5cqT
ioV2/dmQPcTSZwpeBbF28e3BBD7Wo2mKzDFsT1u2uAPEe5Cc8sEMdos9SkZLwUXB
waJHTSgVBx7QAd2DhVCabHZpbP1HNY808W5LhxgwP1Y6U5Phznf4RTBhVFHAJEfG
cXUlS2bWtb1RwcWKgN2EGVxo1afcN7c4lS72k9L+ZNZ+HdRCCFQv4TkjpRUoWNdn
D05tkg5Vyprbcm1okQP27blqzM+cZ25eH7QZ0E1uAVJ68julL/gCj045xxHJIO/9
lK8HEtXdiD12p5/gA+3/rhNTaaY7hxYb6ltNYxH53J19PSQ2W/o9oAHvvZxbPv8L
nTHpFJlB/dLJE3CHTPWDrKYOQfv8P3XApCsbIIAPP4IPpJDSWLzthPfrXRM8NhRN
ad1PyHyijvECkc8RyLkXGxPMu/Yj56c1NYeH4V+DHgP8kvPfyy3jmuCiavtHcN1T
Gl4ttQQAJzcb+cCed4iYhP5d2cm+qeocURKFy4phYAPJMkw8NJ9pB+K5lOX/Lm9M
EIxX6KrejWQdKZPtf6vgcSNkXDFHhJoU6l43ICq2z1v/NZZvEwuMijTfB9Pc/Pm2
nNqz4ZRud7RaqMiswOwCksEsYu96uuywqmClsOtzltz+EPLoCqlup2HyUEV6QgvF
dV1tmsxJo4LqcHK0oU6mjmzW1NdtcEz2Ai6FVwYwWMSqwEcRaqejf4+NeQhTd6ji
dI2UhDtoLouOXx1gA5ljmsYNgjx+7vgb7SoLMmFewrPdo49tbT3MGaZnuGUycNTR
az7OsTS9OFSEqvah/B4bDykAWhYd3GeUfiWuTIaLZ3z4PISUBZgmhlW6aqN6QHLk
mZPXUCgDTnR4t12NvEYkkdIxQjXsci9p5SkyWlR79ZmRGQ7p+7jRw2icthb6pZ2e
VBHULUskl2ONEqNHhqx5nqAOa9RBzB9lVPeNFG7uyyOlogVpMFwO3jPOkwfE5RGE
X+VBt4e5LdindOHrluWszrCVNlarrjOl7SznVszZ0tf9FStTtVnO/T1QeQX/J2xO
EffrgVq7V7t51XX/to6hA2fVTC/f3tX7IF2hWgTRRBJiMCReELibGCqyOJ0dSyiU
hxAhJ0fGYxY8Dolg8VlneslllDBc2fSNloHki5y39RMJd+bl4kQjCF4rvddWefBN
iGgO4IwlvTWIw7+HeVxUGj6iZcgGgfn6T8YjQaRNHfWwyJVUNUl7XT02BlmFZsFo
X8dWsy7ISLdH1NiDZzWPN78c9ZX3Vd7FNVFpuTMJUvDDAWwJil+zc6Pd2SK/QuTd
WnX92B8SoxkiVCSfYkKNSUg0NVx/kDkbwYrAwx+ybKrHZgPYm4uy8XiYRlGcE7FF
RapTFGdizVT517FTVyeCYvgHP4qnc6sxBDyioB69YuMIzphL3ucCD5KjEM8VnZzi
Qyq/58OTRmbDBRIbfHvhz7XwqCy8D1Tsvv+daxToRiWcJOg0WsUP/pIVNshbfEIg
e7ef6d5Szh2X97eMPoTij1VEcnvIMfh+v8MmW73WzVEH29hquOe0Zj/Y9zWQbyTm
jRmZ91yqlbwAQ1KIwmYoWfc1+8uy6acDBktLvc1p7NZS1RPDSNbFzJRjewSEjxw3
upZrzEG8/17vus4elomRWba7vBtL4vhxw/3cEEf4AGko0bNxr5i4iwi6RnbIyFJs
L9IfZEmBeI8J+rp+wOtwCshld7qog4VIoQl944Ozj/AdM2F4cSqvq4JtJz+/7IHu
2BBuDyWuoJP8hjwUzryWxkgXMUgnKGJd0cmAES4mkwOCH4d3NjGb1esjWQwZBgyD
C68nCWBrAj+Yx6RvRI3biM+/UPqi9WNvt51YMzTRRexlxVSlrGkA4UjoRdvfeyZc
YcMmbGI0xOg1kzqIZnXj8sDPOkpern6HNXTEz/U6Hxrqgt7dUrnFyENSlD+xIIqK
+gtHTOay4ikDJJfz7o8MHGqX6VsK0WGiVxieUaX6JSd3LB2adc5Bs6p8Ptk2OViY
TonzxBGdPsP4jtl5FmTJUWeZWNQj0XQ9VGAmqQpPm9NWrXSPeXFqWH6rT1dmUU/2
7+PuoHaRFSMdpWZwTUHp0pGG0VZoFSIrrMEzHDI7wxqAx8CH9LLmMrqHfYrgt0P+
FFwhGLGTZhvmGNZRckW2kBh93aOyWKGz+F/M8P1DFBCdsgaUbMGQUIqoSrelEmRZ
4i9sfne3WdvRZNF+ZU8pK0UwbQAGtWTrs6TefOSIf478G3CrW/G+BZheb08JT8WG
h6ZCl5f3kfuIhUXWFrJWHJuwosqjO3kEhf+2CZUFwGxYapqnUEt+Xh7az86Zxyiz
wPxrYOKpurZU32HKp1vNCSGdxC7bwjTtqU0Ec+6QM9WkpmugPknL/wyKBWQmxqnB
C2fB8O2CfcsyROb8ajybxqsMWBUbq0WWqI5TXyl+SuTq4PeZ0GwjO8/0LwekwPI1
OCFOM41/MosczWT9K8Ms/CgJUsP4RzJkJ1T9GstsuO0I1Sob4rzO2+ZZgmBfO0Tw
xcYNpecKKYV3d5AEgcTdFTUzO42io+8rfSKaExialC3dPX9LVBTYgQ7xdaaiLvyU
DWYWbOUuH79OeFXNkcw6r4Q2tcGpvIYrhaXoAY6/UayCba4N3pkbH9aHD1MiaSom
VpHONNiHa1/6N4uZeN2d092fmC5Y3M1ihWjscI5iko0zPUGrXpKMaG3Eei7kRPni
kb5N+o+wuYcQTWMfvOArQLmPvfeNxYYFyOnPbDzCz7ODFfPqZnvrRd5OU6ME+DgD
fvBYFcuIv1F/oIltu1EXp2ZRq2cjW7G36PefZlwa5k6oYkDB9wcefDzxSdGQ2Qza
K3VJ4uBnU63KHIv9gTN2XUDeYILSlSs+WitXXOay4Nx6D1XRDCgQ4YmhZUynoobr
dxMkfZYzkfF14W3Uithr96O4VMDaSt7rXWlZCI0hs7HOCIsnw2wbpjMt0GmnH8xO
JdoAq3kGgkJi8qJDksV44Xyblbv2L49DrVYtf6juhBTJT8GqqmeVUTKHuENYdrt/
7t7PS3eE874XfHbaZ/HhzT/RTLrzUXzxBPzABO/jksz9URnydLkad3ZD5z3Te6Ns
tWk1yebVgTPAW61Yv9ASa+OHfFYfJI8yorTbt7NT0vkuCgHzxt7mK3fQrxdx+oJr
Tgvv4OMlE8uLO3+/CbU9pxJQxLPVsSL5NmMDihTxOHIIdMfgS417D4S72v1U30iW
qy1f1aw/5jIQ4iSKjWMM9k8M+9HYWR20IypM3PAeefgNnfhrnByOO0hDJFqeoZvZ
Ov4zNhL5D3IdDA/muCLsI8Or9oQP2kEazqhZPnRyl1u5c+BwwdERXsHg7I4015+H
KYnocZObxRJ0+FOGlQQi/lFds8ixH6QMdkeET2+dn3/lwIsHR9dZRqUai8OpHiEZ
2DbjnrVN7mR/iodop/cib5DNRl8MSehBSJoBp4iORiyEhiMKLIexVfvAVHubNlG5
tqf63BiVoIPAg7QitmqBV82GKtkvpA2wcKmHeaYTAozCH76OozwMgOtRuLBtRG5/
Wi9jHpyKNJqbf+BW7heJPGjKE9l0e4bvrMuMDX9QUH0rx+eaNspwmhxFJ7HSZjz5
iVw0ZOwK6mVIpLtixsXBEsmABCuLlWcxVx2zK3m/YbvotBA5e5UCY7wxCVkYmq/f
CUUZ0t3nZ/e1JSYyUQKmUUULlrDgkkv2XSLlSK4NUsb9ePFBSYvGv1Vgo3Nx0qN+
y1QyOQEm9vVrSb5nfIW8U/fZ3b0gx0fOiyXQ9syCx6J1MOR8B0gZmNxtUSPhhPtq
QCfvzQIYEsXHnmRUt0o7SsEt8uc6i19RHlw7jql6JaR/t3xA3tc6nG7rSm1KdMug
Yvzj/VW2vN8XUYeqhElQ0igtipvcNiyN0IePrf6yoIiLT00IlSOjIrpKa1FDtV6w
VYtslNtLN/zp//t+nuFR9jzRc6zWeST+UHb4fwqDvi5NrdOoFMXtsTTmuVg0UdLq
ezyFn/apgE3WWP2ACTDaALFkNirmd8GGV3SfROffo1xMlj2Jlz6VwTuUTZ0GBzA9
Gzwr/LNXPxQLSeZ4HzUQl78UNKcPBgAgEsxAbDdEqwpNyxC/P7c020/SHzfsX7fZ
firx5A70nh3q/jAErNfea0YgCxUcENbIre1yqeVAN0g6AY/v/v8BaYg7IbC7vAzv
14W0T93YhmqRPjXYW9PNvlsCGLbzv7tbJxqwWJGwtmjHcDtnXCsmDKKlYjn6HU1v
ohXMdyHI/YXPz6G1B9170Waor1KgvJwPtiDIXxPOEI1aCNLLEYVDWQ0/dfNOhOCu
UTbhmbrBPBPOjRNHW9Ya98SQSfKTvc/ZWIwODdScuFLXRmQlYpnB1jp3YoJaM4cj
tEdZZ8Q0PATvKHzgE9/nhNCe8uY94X8Sc0uzOchparh7+CldErjceaT8ypA5tWnp
iemacGlQPutQbQrbEWC8kSfI5GdrDIS2w7EX0U/zmNISRrwVyYSzGxCerBmiWAEP
9AFgR5WWsCW29gzdL8+E4cBnghNx3/Cz2XBiBmq7p2md3v6bYDRwwzt4I3m6ez8t
fmTV8BNtcMEFyn/C3QT9mpTx+wzg7sCo8zEeEXdlYjVwi/OVA3SPPY/RUA27wndl
FoChK6mxJ+SjoYnWOPpGPXH3OI0SwG/d2jHiRwklBb/2KO52ikqgtxHRALF0p+sh
Tfl3uswA5Wgb2nPf0LZ3ka1Xvym6zWb1UZpm9fsgJChk6YOJOwCQaRmA9nlC6pvZ
7J8qEPfWmqjmEx6636oCa+s34dYIXz2KUvJPR7747vEGQsat5s/r8mQK9uCujnsD
om0oiPoVjvbANGk+xkoK45r8bGDSP3YgeaZm8tADEwtHPUFpJbn4g05ChNtHhatp
UMEIqXmvoLB5OBGYZLbJEj1oCcjMZZivKB/z+/7RjRFMs6KeVvXR38beyw9Gnprd
gQj4NIb+78qmrNiKJpNxROi3/Oq51t2TxjogzHFgcZxOWxjcvM0/qsDtVyXwkHLI
IFeHdUvhdiP+fiWhbCOblwzftF3phiTRH0WSZN5W6pfmZ3/dmdymfc15Gm4g/Uky
9+P7rkz+G66ahxKqaIhjNEi3H5aS4DZtPG5F+9q6hC2+7kDnDFAosJrUVM18JBhW
mbvbgM1+n6yxlZoO6L+7v+FJlq80/ZlEFzktnLOpV7bnQOj8gTXQXtIbxQ5tKPgs
CICsjS8p+vFohZmvzlWCeQeXcntalrUE7nHumvMo5+9Gzt80MbdFbLv/zCHxbn5F
/JzBPjAdjzgOSB2vTwYTACr2PmRKIKvApDEZWZskX9taQrQ5LadVPbMOtuG+rQZC
qPZYHuEbok69H+m/8GFDBswtVuJHwRusshQPDbyLA+cFcXO5zCUhBylKKYjGDSmr
aO63pIK7GppJeqMjgAzndsBiM7faAhFxng9+40BDyyKy4I0CBK93qvh7P1dlXSFR
B27RJiDfbv+d9Hl2LHbyh7R4/eCKTgpS2rtKnS+tDe/KYLBGpg/gO2sYnoCZ2Ezb
ZSPiSKlc4GUwr7HhQUYfvpFcmSvOPq8aHTapzWuwvUasQ0X16+l4laFr2qXjyVZO
+leiLd/bdgqZXrwQJGQ+v5gKK3Ya4Odt2Fd0rwKnCBdZ8nR/BP538J21J+6dxITV
58l3hcfKn9IvfRJ2ygf0XTFHt+Kdd1uwV4q3590RCC/NZRlHXdWMAJFWkKZJfM4F
PBz59kZgFdHzZb8f2G0F1wPxUbAMXpDecciV7PX3a7CYVmo7QOcDVVV+TmD+MiBw
qYWq03OtDUT0qWXxOKBx8+E1HuUnGYD5Fuvxgd6ARuvn+/SKqhf5sSxSk9Ls81mA
6HGozXh4QFldYkf2EQMTEGEkQ6YG/BRdRzI4BqwnWuj1Hd6QUPnT0CmzTqqnuk1f
aFDFEMuvYSwK6pQWDUlQ7WOQjfYAVWZB1gs28mYHUDXaSMOaaGejCyUC+YtTEks1
660djzhH1odaXduDkN4PHp4Y/hIDSatbtUInT/0DhHgzcDVQviM3fix3qtJyDEsa
PDeLF7TIC0Lw8/pTZyUtVJhrjHWuEAtYGncck2eH4K9xok1lzxCHOvEw6CjWlIzw
5wJsXFIzLObtnPpLJP5JL+8Tf+NFFiBECJwGi2i5sPNsbblwSac3i4BGAVcH+2N/
tYU8ROsOzQAnv98hx6HcTF1Mgkr+lsd7tiH6uTH5Vf6Wd0QLYXhIJH5yMJG5rRHt
egrs21xjzR86PBAYU+2c+OYBurCU9A5s+xFLQf84ecNETgGQPM6yy8W7qrixODgI
VHbGV+juwRnHcUbANy9rTmeCRN3r94hEcGCnXY2LaKChgxwHRP7jspnQ3OnEBSgo
P2v2NcNJAOCjwEIRzVUNUk8mf/xd6ELs0ms/H71UwefW73RSbZro8PMpPMSxUN7Q
+FZckHxrjMC17m+kkoFwL4/AOZeCZvWm836+gb3OKhxvcPftqcg1UahWV7gvGpJw
aHJ0XnKEbQBAEohro0GQPc0Qg1IyE8rOJaCPhwZyDgFNk5kecZP4zsNg3cRipu6Q
ZdvWnSPr3RHVmOjxRSmv/4E3/LAOaCk5VU9DbakcgKpsCDl43OgEBNQgjSeXlSB3
r3+FM+yNchikiOlekXina6sZqQey41BovR49HCxnfRmYa8D7kvbD+DasJ9K8nAgU
EOmr9wptZRiuKSaxwIcAZNxO6HyDaQcHFi7gBMx87gFD7ncG5pGP4RDgM42U+zpc
FEJO4X7v/tSd0oOx0Bnx08a2a9fud5MD/Xnyl2rudk4ZrflNrTH3WxLTjtM95Vbv
tFbUXl3Ca4KX3OjSm0lRIVtDv6dzEwbkd2x/+BcciRi1wEn712otBkeE678C8lpW
H7CcEeLuk3yH5fPlubw789prHz+CcOwe47JFZ5ekmMvfzdKcRUBmNAvm8z2ssX5F
u5Pyb4jUuCBnvwdQookUgSSE0H8J/ojL+q2L6VPXzHMQIS8Ig+/wjufU6FMgVG+0
MaOMj2aTRSN5DUPk2lRDFM5xmiXP0A8itEPzfw0yc+wASNPPzRTezStI+BXqbWZK
GNlibIzwNHzvrYox0Y5JKSd/DNL4VydfKBPIwV6hr7moyBqLU4/Ipv/WWMwQZC7d
QP3Tqea2r/AKn+La34N/ApkO0Pvji4o2tDPopbQEwhuQHBu69p7RUDhM2bQltqw9
Q5FIjBefegPcbg55aQBvqPi1lfAa7UkTZuHxtgWVBkxDTswE10TiglOHOwVDwPu4
F03Jd9BeWeXZ4QqiWclhqtLJsC4qlDbFcwGz5IY6wQvtyB8YWDdr39QLyuqmsEjl
xigskDxazOW31/uF6uwZ8c3PwcWdlneNHIICgIWp4pqSoU43mZX5Qx1qEvfTMdBO
lc3MOJjgCdFNMJwgLiblQf2YPtTdi4+5zhx/f65h3qBfxpsWPaeRsnE3vnJ6A4bB
soo8ETwmZdBjL385BiGrpfPRxjFF1dO/E90M6g4GCzyY59VIWceQYZWRV3E5DKjG
YYVeH0Wr0c6692zsdk0Z6vm9LXpoS4aRN3KPvB1TMVkX7/UGtikM+rNegnROSXKT
ePXNdRaed9pF5DX+WWAthAH/Minl5/OAfjT4xLL/mE5g8IhgnsAdj9MsPxYE/pZK
gTW+qQG0uNpdI/UNDmrM+AlUN36nVpgI96bpd8df1vuR0s4OGZa+OvdSuORRuXyY
yhMfm1dr+/Z0kglQGZy0NFqVF72zuhGV2Rw5TZUTOFlYgUKEd82u+X/EJN60BHfO
CoI73O9v7WfNx1yWlK0q+ElVHds5JmryRgBYTpljp7WLo2wE1GiiSRlW81u2bE7v
lbHg4MI1cFyFsG0CrJd7T0fKyRwkORRLUEoPZtKcDGJdvD4eC4GO9acKofXqoD18
iY1I/9OO3xLXHtaE/EgMw1Ykdohnt+/KynrtzUQGU4RncJUqj9+9pSsHXZPbmGCr
TnEucdX7c58CyyRr4CKwZz9NHk6gqT1yXJ91kLxlU8MGR3p6Q5W5tqeLKQ6x3a5H
zCkueMDU3j0/WsGbrsmII3dM+QZCH5myoxHbAikST+ZLq3UUF61ZKcLfbj1pMcCU
DiRGGhMOzvrikodV4MUwk2bKf0jsjbytQhAGV+CVliCkDUu2S8UQOwUkVsqhAFDh
aTsFLPkQE9HEuRAjYQ2UsXX3dy0FumzlZhMnp+711JO5eyBGbqPNJZhqcoSqAeDs
bcm5Lv6Nnz/RftfCrBt2VbEraSvv7+NQRKptYsSPDtJtw2hJhE4UCycTgxMzppMG
HzOYQruwLgdkTfefUdOAGOi5PDl8zgmskeh3wS3L0FRsH4YViOhUOg+JfsL2eBUw
+lW7pRhMA6ULzxrPz3iOlfz2CZc91oUMaecrRPA+hJWBy88MeFVyIBrznYR6vSSZ
URIMQu29S/X6yLXxqfroNhX+w68aNtseN957YdNoAkd8zXwOUkoWU3uo7M6L8gg6
OFNyQ2k90msD5ZivmnAzboNUuF+Lkf9Dz4VHV/RqJAzFFNcO/HH11i17tELOnieF
ZxjZYdTuHDkc32bxhXlDZ7OYuoBUdBJao7pCbN+nhVyaLryP8jjELB0uLvsTf024
3ei3X8LkBkj966zQdMRIyTdLYQUQ2TqBh1l0yCN4Ynl5ypqrVefz5L+UVKBci/wx
Jm0Of4GDW2ntBoe36/xUufwdbg7t9C05uA7TO1Sc2FEuebxs2QdlehvZVolYDThn
G07aR7UoaYFKbOs8pLWiNLipIDtSf9BTXCg233Tv+65E0Cz2BVpyhXFABFehXTxb
pF2a5q7S16SBVcPjEMAh3g+Ap2J6sX190KeFDbFOerBascPXOESxzqA0dCaDavge
hk8XPHqr2eGWz3j6SZcZllmO9vymq58ZlBiG64YqOiAapZSLwLUcmbPk2OnQCilP
HdXgbEjEZS7dNWUoGV9mUcByP30C8NYXs88XQcuxqtYShYkGrS+Snydof8mRKcz+
PgSCj0mDCb+zkJ21rbgiGteUtst7KXAQy31+t843nI1mqeJOP+Jzv371AA78t4Pn
HZfCWXDo+c4pGkaAX93/rkYzRO76p3BrUS+g9nG56wuvYVEe1UzJu2y8CKWluerV
gqv9M3EtADGNN9rgqwje5UJYAP/c2tkiQuSyR/cp781NhyLfJLlEiwlactYD3b/+
F0rMStqpxB3CdUTRNli53FtmYSXwNiJaoKKItDEHmKQgWgyRjs39HrmtsrMjwveS
qDzNJGXnbkECSfhTRfqt5hSS574y4W3M0agZll5ftZcvRXKXPS+j6BpHztMJWIPV
L0LvkW9xMSCRFhvA0pKFmzo3a4QbfWzi6Zi04VPVoRGBVH7pLETWeeNgCtIgN2VB
aYsiyTZxaJMMQNt6NueQvYQ7DaIa8nLddgR1rkfujDbDEuxOqM5HJHjNXelgrRiu
h3Igcd3NHFQY7LuAYj94SLn05usvYTYSJv731u8F2nYChh2c+MOov/HmEO86bO+u
gX6eMj0zVdTnLK7sXbGIC2RXTBImWx6XwejHlDCKXVzis2wR4YV7XXAhq93C33iJ
r1gMYfnwev1a1F2Zr1NpELtBedEy3Lk8/52irIWk6rMkrS3ZnvdGHTVPfUh0lnwa
OQ1HOgNTaH97z9nL0th/CaVAjH98dWIr+coJsSHNIJH7KvCh+s1cQmFiVTF87FTq
Dcr2PQd8RZzsG4BGnMi33nfkHmBneu79ovBHKkbak++3ftKB7kWHdHY+NxckGClW
0AvKaYDm2wb5kNcsHA0HUP7VyOQcv07lffAJ7p1L6phNoMgSacNBoKOtPR1oYS6W
J7yXq1vlBU4/xY7j3VH+XzQan+bSVIzAz0CNQEP9HSp/VWNmlWP+3OUhDQG00pGm
aAYW0IfUPyEIYr5WDWG/ysel2uTneTgajjSEvMnBjuG8Gdo2uXFQoumDsdiQx4C1
peDkDdAk6dKOiv+vFomekrzP46C8auPUJV8+9fq66Bu/q3gz+KyB6vBoVTy6dBeJ
H2NF8/Ln2RmmO2+Lqcl8mODb18XcAcPvrlfzuQLM7D3OHMQUXRD8HVoY+79ZT29m
YSM4JT3aW3Hj3lrhCEYpgNXxCD/69oKejY7o+DQKu/i4Z/bLd9ZEAplszFnuS78V
9kdTAbYAOE9aV0XrLopSEl/kVPW/rhazwuf3XV3KhsDoEN7pYSM5rZEareTfeTIR
hfwK9pR7vDx4RRAWf7FUMb2wpKzcXL7cy3AaVk8UqdZFzApQq0umhyWeQ/v1HzSM
vlRH5KB0CS47xjdrIUqTCjW4dZs1OxFDLs8Gx8Bg10BZ9gfoWqvuWfZnQ0/EaWwf
GrG/9Xu9pC6qFQxZCNECmxKjGz4Ou1gQSx3wF9GcZ7KOdcZvG0ycPhqmKjit/YLM
4C2iCJwOHzMPIk3/jpR1xmpyuIlqDf511a40wkbyKWR1TkLcoQFjmbO7eGetl1XE
faYBIKsnvzOT0dfJ3taWh+dmhwkwDnh94XSpQPdjuCX/hi6qSveDCxG7wuFv407h
edJgAo6lD00tWVp/53sXgUlHCra/LU+CrR+Lk5uvJ+6EnSuEpTNaczKKZlvNApf5
0lMVEATutw7zYoEa7Or4TFP/GlYrRvXVODyOUyl72WRW3Q5Zeh4Bvtq7VjcRS91m
YGhSf1yqoPiijsm9sWfX7DWxX+gsqPHw9+EFUCk5RvmzFSJqvubknjsVL9yEsju7
4Ijgvvq31qNi3wTLz7Y917VNfypkBKt3EXFWsTl5NKiyvvAs1s8V3pjjvjhVN5jJ
D4Ows6Rat7NX6P104Efbm7B7loxpXk1sp236YCyqUDWJPMiEs3zyt4xOpyH+/hNQ
c2M9eFmia6TDXr2+YId+Db0JZn1OaFKm8DD0OTL8iN5ouZVprg6GyDUJkrmK7c8E
3fexwgJ/6aAM89KojHUJC1JQ4v7XiHIjNTK4aTDwehaeVFqsCyCEmiGN93oakjwa
CietJm5x0tEUUaLzxQaGJj/0Gw6rq6LgLYjAZ5WRN/Pu9XRrWUHzzD2meiT/IZVO
aygVpYvHi5kLHL6nQ1MIrRob5SMJaz+ZVDa9PpzMCNKfpUL8yBkpff73uNVR2ooz
mhkWtG4stLXR+wlELBqXls8m1p39PPpKrcxrWW/ruFQ9GipSmVtkwktnKVSQcuPU
g6tNe5GEqUkABoAIo2U3RUFOTRH5XmzPGp5T4ZxSdtX7+iLcV1MLyiChYnT1PeXu
aVeohpTAckhfGzXEs82KHWf5Ys2q1SXnj1/LFWTBh0FFJrtoIKxRtwdJJYPyUxxV
+Lwdogw1jxCiLwQX7mLFc8+SSh8JjstTUYkrKCZuGqEvYGt/S19BXJh66M4jvAiZ
Se9Nd37mGHT2wXoeyw5ZzB4jnVGIuFv6encXWcqLSTN3SeXeYE5uAyIOcwLNP2SS
iH12l39MxE2MxjV8oa+6CKj71sw98Yw1/4o8k1H/A1KXXqydHtkjJU4kRKoOfqWY
KHQITd2F8FYjQYbIO5AICH/o3Y9rWut9Y5qlt2ShYF1TdnDKyJ2mImFjpRLdoTtz
t14oOaYKEaFcla5M5BuC9kjE51qzI7orWBnl3xH988nBr/sNGYsT1P2FbDpZrNa5
Q8fCCc51PCokJvxMYt9yb9s2t6UE4lywx3off3CJuPEihbUkvsE+CinpJLN3yIya
s6F+/QJkWu37F4rNFFQE+4Z1o3DP3otrT34YKNaszThoEz+3JhwxWZNYLdI02wOC
ZVCA2IgN7XaG+44uEX0GT1GzUUQEMFLSagM2hJa3+QTQuIRA/Ne//A8K/tNzyDK+
PO0UdTs3sRmrnFtjcnlyAOqc22hiIBG3xW8MP4KnlRqtqNI5NLM/AqdW28dFD3dl
K7Rd77e5WarrWANtBc3ejuUAkWLFkonab8Nv74rCsOgmBQlxhUO9/1ZG6A4Shddp
l/mme5LDFhgGVFdFvJ/YqgfEykjetRnAYmUVVNS/TocMX+r1/a7LjqQ7tzXQm8R3
t/qzMXSNcI2B3KNg8VcnY1aXFVXUMEuKUrT94rJl41KXYjQtVQXN97Mdgm2Zaz0h
2BQEwUZ9cWVS4Xc2M0DdAxTSNIBfgMOl8aSvKea5snjpYEnlMEQmfww30A0T+k6O
ZwCphfc8uxFKi0g9O3wW46BhBw88IjbdB1Lrai45vOCgzPdU39+n9wUZZOqPymKK
BsV+5edM0k/gdpzSsYwV2qOAI02LAPkHr42mi5yh9syqMMcxLPSS1ZzarqJS+FCE
gYO4nFXgaBp8O7oQRELABsSXyituzStVb0WG93glCNm96l+IaBM2x+WnTPi26YqI
nFibdpXW0S3smh2lKKFSo7qe/+HRYXE2GN5K5xUsib/O7Fzwsoksl3HX0vnW2kTb
WVyyfcrUl+xhGHZ7pU2oXBycCXNC68KyiYQk4Vee0qBqSXyr+8/9/fjGFwCnnqTU
IfSX3iCpe8U8rVSWjSx3jYI20fpozA2W99fltRCTjO+bsKEaclIjst8chO66DyQL
fl1ETyoEsG+2V7pOTIupuh1jRNxWmQxDrooWIUCLeIAcVf3ZkWMndLrpHqrnmKPO
VJDMW+5Xi5lYKhtPwOhQh4CNSKQlKvq1oCnm9NV1LQkroU6MFrOSMqupQYL3YWcr
laOSptN37gdYXEwChuJtdzkrGAHLs3yWxXuiJ/vBoykaVdGw9PYZxqYx8A3uJOFu
PrKZD8ABtP7a3KWl1lAMGrGAm/ef7XUJ76s8ABgyfcQ9UBWyZYRsfpoB+7qx4OnA
kzD3dGwRigcd5yoiCRZD+JiC2JyMvvm1L4ovEEfytxfc5hCGJB0vMBdi7fGxHyqa
t8MvphbAwq2ZCdnd+InwBgoSHTO91TZDIXGdHdhQySolvvptLUsIfy0wrDrUX0UR
sWkGqKYSsuXXM9AcWa30WmnNCLQ2AYRdSKs18xNptO41IxCDJBjzNSQtUQ+sad3o
7DQhPqoKWEP41RTTVCJzpGReoBkO+BC07oBP06B/w4dAQga5q13LgGqwz8lgDAK3
DnvvH4+wXsCFZRWR0McDgE7X2yZodCg+VF8baVmt4joZumwxbyuRL0YIDDdu/KAK
RAfsRt9KVruZ0S27vmR90xV4kxmtgtj/9waCo9yS3iOELcakoHMRfZDXf3k+YNNj
kNbC8P7ABauv1ICTfK5aKDh9EijQJUqSF/QrDrGzNS8BMQBajwluI3h5oLiw3t71
SAusBVAVsHH6sIbzC/qIWpc2DQ/dWnY7ZGtc6Z5uEjtsd9E3ZMV4LvXRnlGwGjYf
XohWwPRuxOeJ3pWI7SLaH6pRcBY87bJs8Bv8xQOpjp3M1lw3omUQwvJxasoYRGyw
3JIJV+QdTgxL8lkHcwOY9pvi6wuR0GpVd0qFqyzVYS/rlVX/nY0cLcDNNySw9Uj8
hVfTczQwQWMmRdbnaj0JXcbdKo1BI7imJzMLKfBbNl1GTNQCFI3/Z0sANYGfdNoQ
tHX2bMCnXApntYS2ew+Eg9DV7di7DdeRp2CB2C6Cm9TmD6bJSSknIdePgEgpY2hq
TrpFQVBY/rMZ7mMz+8LCDviUSkpb1ZUuTPJZry1OgDNU3sPFoBPHs3ylDJ4K+TVo
ubQBICvmZ0W9COJoUnT9fFU6hScC4AogiNogJJGx+QCQytPxCRBlTTs+oKWmypZc
3zRO0gJDKt4kisgqlmrwXv4lyt5I1lHheE9VbLcNKLGDRT+YYzjAnYI7A6fZLWPK
mgvGEbJfzsWmSfJlAXRfGX93Zl80oFVXcN5Dqb/0K8uJLxAgsvY9ukKQNxHCXCg8
3Oq3sMygJaxdcLU6XOPqOR8RaiQ1TZ5AFiVc5/AKTJ28zGWEjzOJ/3U3nLeFc+Tu
Ce6x3qLh5RVpl+unGYN1Kn8ZHRevv2fkN2lX62rjvNQ6t7PIF4LugK+J8n1WwyXc
atd3v3p4vsCs1hpHJ36wjZILj/5KXdzU33UQScJ8DGX9ForqHKBUhlyE1j40WXW3
VjH8KfNjlQsME5DlH+KrL9qnAgnoo4kQojpBDyXPc2uIfduLvclAAwHCVvcJrycx
le5O+v6e4N7UFyaqn9itfGh8W+oT/LjzyTnoqHOend+m/39VbC3GnTyGlhZaSrLH
4KwWiBwMhrMPYaYlMXhg7uPB4CVpiWr16/7HAf/C6q418uE0qJOo2vtznakRDysE
2LEoFf3dPcPHNw5wSa8Bolp5XoUhxetTMOh8HzVTQzTPH6zRlyHxuemyjlPMiiaz
z/l2wzPx2bKBhQkFosQUBrmqsBOEAyTZTDJioFL9px641/3oRcsCvebv8+grRpHj
9MJhB8OppxPhYWF/hjlzoqB8vJhCmGhx8/WnzUIPLzPuWx5B7FxPYDEn6gqant45
yIhBDNsEsPWbS/mgdN4ZZyDYlS0vrfzlGFVp0kVtkfDeLo++TkptpZJ3Hx0AUn/o
Fq4sBFmpHe0cHyClOWvUfNQ/2CR5pGqlIXqE5gf8sRHPMZsn1Hp4+QpT3KF8PuGm
OsQOaZ4VTNeEnlQbHIWLMamnGRtRARkCn65z07/+P8Jt3taIyag4y5az6kdKv2Pw
xf6v3GrIrvusvyhpQm7OdfxQdqdJqN54m6ZNpW09WlVpqYaaNqggB0ESMiKILwmT
1DeIx/l/XbFPqkZHewpF/7Ml85SwNs+TAnFodN+1p3VP5TNYWHOxzGtTCA6FXsZU
unvi8Ljq2KK9432hsRI8K1h2N0gDnamPf71Kpyi7eI3VNwUU4YK2t5T6krVCzOYl
6mndhfqedOYHSqu1bk0SAVM7F3cDK5CEeIgbV8fijWpvZDC0iy1Huz5NbBfWgrCl
mMTNeWcbqmUW2kB0f6kMz6bufPlsHGpfNpUB4+gKdFHRgfW/WuPLwNG3AQYrJKD+
zjvmoZg6X2w18PMciFLZtt9OYW0gSocHAMvtVcyhp+m3zxb8vr9tBVtGvr/bKz4H
E5AmhbGNJduDHzY2I5DDZdhAkW5IZGVpyTLfOg3eT90IAgStq4hflrDUtd9DXjiR
V58UIILAkegtl1kypCsXgoLoLaO7idDx/FHBPvtMnR6xtvOmPi2wpzLXDnnuCoCq
6Xgd8LQzGPLL323noaBzGqBoApBEUq+3ucwCUnpuTsrR+i37FcIB7SPhh1ocOSSB
1h+attHoQquP/WkAqSlw70vDRG23jF0vHPHWeyxDF2meRsjbmmHyMSKyq6YVNSXN
y5VP2jWF11bXydgvYgt8VEQgTHPgiaqLd+TkUIJ/1lBmVxQue8z4Nv3MAyoRMNRi
kVlW2JzNHCUKYKbOCEiSqLwxOAu/vSSj6SRAXZ3VXwABMvz3A7bMXqtd2YHJAJ9c
bmQ7RjY8CV/lkUvRdlUN/3RV99YkQvoQbGBnbotAdtmt1f4veAaxnmfI7wUAglyo
TGcgjTPGCQwqi5BlnGlZ8J+dDND9nwObpgh/B+Rcq7tDza6ph5ROQDOF18dntRPI
x/eq/5ghmWmH7ODyuSiAbzzBLlVzpkuhBvq1XYhY7CzFUvvdIKJjKVNNXLTjCzYw
vUQqBHOV9FAeIe4j1AdNMRDH150jHFxQ1924ODOu32Jr1XNEmrMFNM6kpco+s2cW
01WgdXToL+mNp/Pn3kUjCg4bxD70PTkBfSm+uKP53DuVToQzLrLKftI4bD/TMNXX
x18LRtazc6/AJ8Do88HXDz9LC3PrWz2lfj5ZENoc+X+zVMVXaqMsx79Q4shup5tu
JmWdkhd7JaJXQk88/V8dsFG/xt+g035zn8o4ui9ZuMlpk0B8ngXtQnItHcvbFhmN
LiPQNofwXE0NujdGWKs2MxRfL54zPjvSzOggsG4tN1dMv+1WvkrXNoWwXoRCr6sD
5sMTALZY1U+XxeuhbS9RdUvXEodegT6cIpPe6n44z6tPlMBNxfAylY4xIrP3jzYm
EAIYD76vrZfWCSu650q5JoLbBEDycPOMhNRL8xK2gX3I26XDOrB3fTJ8hqsWmsVX
b5tv4mvQdYS2ZAnBuoiL7RME3k6/qe1SHoVHwJrKCaCoL/vnVq5mic0qG3C+NN2i
lBdIvUX1pB7OF7GeT2CjR8pN6lgzSErEYhnNGtGQWhUCWZzMorocjEI+K4tGom2J
/sCJuoG79tOQM0shOccnYCheqvZ5x3SAM4m1LmG+4pP5sQ9P3GVVlSV4aM43qZxi
XqMf155JDWF/287Uj2N0DAW9lXf47YO3UfkFeF8SkKSkMiSW4iOsKNVODOEYkgPp
V2PgPn9LhEqErAKbQqEeTONKNn1XCYlAIWxXlEQmol3st5RCeqPpa3oIXpuPeDjn
qFl7jmZHLxF8m2+POtskwf6ZnZBMeSmU3LISFc0pVyMC44p9BQ4Zcmx9D/Q6QNSH
w9bSPa84LRXPJoH06OsrxlDVlhmpfbq2XYwLohSYzl4tz8x4XzsVYwnxQjKvwxfc
y5VIk+/1pYTWD8X00dXFP1IH114MaNPSLuQl+j7vLRa8rXxAaMeYr689CygEwPXj
7XtDQIffn7fh6fjpyrlQFEUc9dUOpDnigTksn40+UH8BUzFlj/6fNkbYSH0zookB
7DKfTnnh9EP5yF6kdqMFbzFhhSDba+5zH+EvmvJyEnm5EDr31uVA8vb1LsCijAII
ee0GicROaxP06cw0+EGaMT7OiLM12Ez128W3702oPq6m9QWDq2GiFTzCzTM/sWrE
XAg4ek/Xlpb6iq1XRYJxvuhj5q91Ll0ieQjCjxlL0QBZRSrAVemOQap0AdnHuThh
DiolIqJy/nJ5R4ecu1Eab6tHTUzaovMr5L4PYvuhnVCmeTzmL5waOfJAWnTojjtD
MQGLrzWlY8beb/qCnSq7e03/3WkhRT9yaQyz0V2CtdC1ZEgM7AJYKHjjEXsmtWCg
01eT0JzjL+ZtXMrPB3tkagA4m/p0DuGoIt7DbFtSiGrzmgH0rMEw0m6x8QYGt8qH
Wx0TZJb0oXQWXER1hNRGb6xrVT8zTpaRakDdo2607j/9LtgUrouJMV5FBSYmziUA
GYCzX2d1siYwLg8vPQEzXktxTVdMTUdRFU2QgbtJR+d7fI8wn1kpEWh0nFjWIGF0
MJXgVyTnXpZ+E1k5ndzWsjzMlJeZZ14UxQPX8GKlsztmgJt37g0nDmhztn5qzEpz
c6HwxJsHpJuCmlbd07CxOWj4BNx1DV6cmUJzlLjMRNFXVvFV6QQ6ADvg/oqofNrg
1po1yiuGbAgoJQd0fEWZgaouo59bz9RSXm9Iy9QPWnvx4/oeQx7i1awQW54i1LEQ
xzck/goNVG4Y3kRuhSJW0M2TuV8uk8+DabGEbflygItl59psQRnqWlEzTcg3M37V
/Cqc6sm+Nwd/30MgRXcwkK9iJlUfwY31522QHRKzBCUaZMsyxO3n/C/znVEyNaka
DNQ3sUVjf8SGdqPINEw+dnY7U4OS1Fyq/VtNIo/+izxy0diZ8z85sOUEpovFKUs3
qd6wcw41f88OzwvJQvnvWL4LWK6UlXS7L01eNE58GaFpxQy7jyBKe5tE0IEgvefO
mxhgi8u+AezQDsU5kYeFP5mp0gF5X2YIZJd/lc1BGGJjgiqi2jvqwsSs/A2Vkev/
ImfP1AkCLZbUu5afix1Ne7RZ+N3O7iR6rOb+hX1AkkfjsOrj0qWNHOKoiOqBmMfm
wql6NKFCv9hEhmgGUhUmqds3NfgQLV0tr2zgmMwfmrCgr0yAaZmsSo7w3nIPR/4a
kw1My1enGlHU2uvuTPw5V49uPD6+YMUjMf9/LsiEJpiEzDqphZyVeQcf/+MXyFkp
C6Pca8g+1v6dHwG4+PbKXSx1vVfbbRo5yCAtuOaeTqp2OA+MR1Q4WBI81tyqXUb4
0Y/8tTr5SbYxRlF76284/qo8Gbwhmu6KI10mPzwTBnYG0TvmZ31NZbMTTRteZvI/
lU7T5mvw6I02mup/KJQFp8rRlSj8clsQbXUFbKlhq8Wqoj9yBQkr8Kd1R/RByB9D
bVmQStqz3zyFtx6WS1JQzu1mX+OPw68IYpBPTt33GekoiCSa/dfyq8zqjFe7e1VR
NrD4ivIYDbALdOUcj/QKrGe3ZYDRW2vk9knfJ9oOB7E+oDaWKFiUE3A0vnfJPuh1
XXGP3jZRThbekkBUliv/ZDOxH57MfPYD2k8ujRZ3bEopx6bUOfidjv16fTm04q/5
WZkYVjwlbonBzC010FXanDA1XleMhrtxGG0S/nZv4NAWeY6XyxCKmKEwZqh7MHMg
YOx5nB29kObTToOZh6LtHJQ40PO8nRs7djjxybwDYts1wtLbV11ls6MrgfQ9iPsZ
N58qrOvcwqLwPYMKp/aRPoKhCmjaUGL9iw2Lr2dz6p10Fe1/fiBKzztCzjSLv5TB
iDXGBYYS2qAZJZG6JbOMMo4VgUAcwH8nMxzqwoA0MJCQfD8DKCIwwJUV1cpJywg9
rvszh/xWEK+xDcgZ/H8tH++Zfr+2lVTIRsOELNQZZ0gZoUZjzZWWRse9WLDf6ccL
NKCnGhu13kp5nzkYR5MlvQYqqUn18HR6V0Rlw3Uc81aSPHWGL74U5NBs1pSQbCC/
LK+ShGdkr3EoBlbC7tNTipqnafywkK32bJoNwdggcFTBTK7vNndxi9gFnVIPN1+J
z1NWTJVaHYYRQG5m3tuPSUiTtlketxNl44csiOEulpV+U/tq79xPYClx5wF+Iyyx
jZw2DY4oAdjjr7LzfvtBSo1gBVx/m+6bEuN0ER1ylDODKzQKzBvSuBwIpOZCbTf5
wsOp/q9lC0UkrPcJ+fSKNbvFpml7fBriUUJgoqDtwVZXg7p0n81Vzi1JUATC6zbA
EzpuUzJ121KLYO/AcHa16eQg6YlmzOOAkyQgnAR2wa2vTrkV76u7OJYquk1ORJcM
uuX8q8W5+CanruFvRbfOb+qiILpanRElX2onMhAwQwkIgHMHyxUgCFrMPJM2jR0s
Y7fcCrnO+lBKl2CgD3OXkHJjTVMKv9wGTtatmIRgoFvrrvj3l0usFenWwlUJ46sE
XmGbJy2o54sg78aCRhCPGAaQdI9Qa6CT9KT0RygCGyjX398hmayQCUZpV2aNCoB7
/d/tIhTDwKdv3QO82UH98k1ipBuaGyzCpugzBvSLNGG+I3sa7VLrX6fq7PU3/WCH
AVJLRWGpeGotSLnXbb/4j21UO2qRPht8GNYy6Bvnq6DZ5ugcObRs3lsqM9tW3h92
q83EkquYLjEdc7VnihsTlGl4VHhEtmM8iaCUHDCr11u+1Du3SupNNiUT30skE6LT
uz5KXuCkqZIo2/H+/+fe+f/HDankC/xXJNXrELikR5KNY1yrKWD+TY/wJGS9oKkG
OhL49i7lHYM77vvjDg5BCf72O3y9HmSjAr40J1/um1aFN0kaBcTupRxYEX3Iic4y
tXdOgK4XZDOtb3tnrzJmAtUuUYGSU/xgtESSll5SSJe+Qqs//wkbWfKNLenYUrJp
ZmfSEmOKWAe6btKhFRUZdpupQf7s3/l5qTsQlJRRNd/zJ2xyxXBbWVYgOdLVCdQt
DQqqf48hytGu7WAZTNrPkOoFF1EMJCEyc+BSilMQEgWpUmP3+pfdeaBb1XjfbodP
Moe1oFPTLIymljKpoz9gUM1KK7UDR59O28eCqv2siysGNW5cLoK+OtrZ5Y0nzHPN
o9CsqhPMKsVY2xOejSpJr4JL67VAiiR7gyC9ttGK25wHURQQKi++zp2OzQQNSsaR
35O/68a4mfuJFEAa98HswxX7jCy+U9co6Z3KEW41w8gADEm+YxiC0sY9dzTr7Mt2
c/m2JWzWXRowI8Gk8Tdnb2M4s9aC6YTgBQ6zVj6cSHt5q21297eP5A3gjVQvHfQN
MPI3mUSitYX/iOqoACrYQXarIlPEsjMTbM2b74BZH98InNkYMDzrtPxiOeFhjoKn
Y+QwBtmZc3nN4l64U3Lw5Ugx5JaiL2KMkg0S5Oiq0m062mqjReOqd4Q82OWmHhAj
WaGs2t7W27feTHiQc9Sior2I/9a2CApQ3j7qwkx8UAlw6soKa2nC+RcYFN+w6ecY
zmmc4V44zV7/Hr49DoqvnP4gSJcgeBVZwBQ0rGr35wYxGJ3JovdWzzucFOEA6Hfm
kNcfR0blsW4luxJun8U39OUOG3GRytK5PRaBnwn/QS92vwZiGqXfc67GXrAySiMT
11RXo6zTo7MewUs54cSCN0La2dxBLOdbkmQmGvsn5/Mehlgvh2Mdpsst7phGFzpe
RFnrRlBZfFEcKQdBRvSY5ZKAZqWSoCjxgqRfasgDp/jEtSW/LnJyIvig7q/eOp+T
CbSkj5898DKeL/mtqsfe68kRHs9rq6tU5FN1UjumVrtW7iGES4sE4OWxFqflkIno
LeFa7yRzgxsh0az5Q63rKhLylDI37DMeaYoASjzY8MtdyP6vws6psf1fleI6Bs1I
bkqSeqbkBBZzvn08uU8AVOBPWzqVO0kPwdWwN6Ed3lvRZba+1NjGtAkMq90qtsnz
CKw83zp91WTgrpHSSXSMXsa95Nb9DufgN+4Qyrc7kt7xHRb00aMK56HB5rsuPfgb
W7PWNo504v81RsMzFozxpnRqbjqB4M9qXjYAuE5pCEtkwUXIDIPp9B8PygTEMA7c
vyFPfWjKOqAV2Y+90Q+2H3RHWTad55hPk6oc+tk2w38IGlridY2rLaRKkuPro3sS
d7k6iUQ2bUkb2Qhx6Mb62oXcrvi2Z4MFPUm8CeCvEe3o45K6Uwjng/GaZ06omns8
Tg3pz/SdibysLrUVMBWk4Bh9e50qYiEuZm0ik5YLKOcIKvu6fo+EYIs8y+qioRXJ
POehX2leNbPgHHyNKIjAHZUoI82hnbu8Cmha0jefdk69Ql8koXDvhRmG/LMoTblD
mQHehNWVPK2gQHht9mDIZZ1lC/Rkayx9zYMhXMDZjEzu5q6M2I8FXhCKZX4/4pKQ
fkU6ZNyJRQsf6P+oErwoly0l3CpdHk9SADnUidXZ7+MWFz2cmRNVmmm4KgD5g7SE
aDmHK5tOOk48GeCoH+8QRv1rskKTZuyBOAO1xtg1Qx7otpxGj2XvKFcsR0onOcm4
nRDMMH4LpjPSg9xZ7YIlm7YzFgvkeXNXUX08/LlACZ3PWHpswpK+j+67u17gMHry
sZbAWbgggOHCLbkNP72JETo6+v+Omqb5ONJielEpuQDRLQs2mPHq75qkp8Km0fxk
oNLYC1Zg786eRFNKmap+GCQ9atyavx/ssoUmLje8r84rzPPkPQ21vgXCBbhaPXWR
Q6iC8b5WEism3RVI/7rOCFlPz8V2BdumTHj26soZhyhPBRtnY+3bx7NKWHGJz/KH
Sh6ttTBSq6HjHntP8ks9DksvjBFhNV+fTSO51VWKvpLnq5Uxx7bsF6GhHKvk39eO
XM91sjVyRQwZVCCutoPiM30zK/nVrQtWu34joc/Nhi+73c1EZktKFWI/54faIjvo
MJ3yS4k5vhwlgc4PgW+qHECN5p+oNAmkkwj0zMZD/FBY2SVZk1pTtj+dyYDesfXk
zPPoosDNtu7OaTh2R9zddZVpBkFDQYq1TBhKYp5PibWj5eZ+y4uAR7pGnsNT87LF
2yGx57RxyV29Hjhu/k/CeOG9+JDtprmypxJI000GG7BeQnX9cikeVLe8CYPaBfjf
q68FfVPwOgXxQoz+xflM8R09XWKGIOfjyuzSdduPhfR/m4Tpe5TvisSq3yrU1KpB
we1xw508sJlPY8EhhV0nQmXnkOn58dV0axyLEL3jX17eEoEdg8MfJsuKfU2VMKwY
tZMl2iW+0pONerkYEgE+KbOAxs7hyW81Qm7Dqizbr2IvYm30JSOXHEvyoQTCZ1KI
m44GOXztwztbTh3xk57cvtIPo4oHw5qJIiPQSxNzo1X0InaLJ7bc7tFYsfuRPeGH
vjGz6Lv7y4dOtOSO+AuniJM/WqbJz5J/fsUpha+OkQ0yA9ndhNK0Si8oCGaMQy0P
IfluQJK3OVUnfMgkSdO/xL/YAxkCqG2ZvNby5T8Ki6+XDi8g/gX3bj73n5jWILSI
12+tbn5mttJrynI8VtFY/ag3tukbKnFnD/aTKJ5UwfG/Z5vGstlokKrMyIUHnWt3
VsQASFtW5uqWAT/hStcCgRDnk9JAJituoAcrKmWvtLYn99O/b4tZKYxAOlb1MOp+
zejHYVbT+97zDnliSZN/KRCa7fATHc4nVGhuudMUxrJBrAAvie+CJIEq4tXUxZbD
H5cGDUbdjIrwbBrFNf/uhzQBVRPQqSFoXlHYqM5LE4iToEevzX4MYMZ7CCiu3KN+
4zqLv89VvTHPCHKwS2hwttgua8RR3Gr/ZEa7ZPzyS3lK9X82KGKPYXMbna4mmk+i
e6secVDF7vJCqO56AGRNLF2mhCOOmdHBfGvaMbzVvyisomCuX/j82QBP0fHqIKOn
BY68rNh2Wf6O6FBhrHrDVWAjsFsJWvBCCQXlA328OdZuibgU3zHDRec7NcPXdxLC
GjHXRIAhtSXr0VfMHjw9dy7HJUCxph+ukm+zhhP1SeLAAKEBLc5vLc62t426q0nL
N9SkbexJqBW0b8ATyqpvWfq2CgN944wDthWYqTUytJCBhMuvLDnmNZ0noGji/Fj9
YksDzmM89e/1atStSdGWJcR6/k8RjwDSN0UY12zLqAV2S6sEFF9nZEJbZ4JxWgAq
hSnZQ8R0u0iHH1WoIg8tA95nAfU5n/qeFPxLjeROq4KPAQjyx+s+5uw1m2gAtwsB
Y6GHyO5t17WnJM3ctLZE0kqhxKbRLTT65tRbyhZiwiEbEh/ZkvyW6WH/ty2mMlsl
yRFubF+8jWJN2QAxCTM3CqcBUgAelo59EIJxmEJ28iHWWIb5UAA5mRXr9IjqR7KG
rHdSQIBra4xO4pET5kYjsL8xXijJ1JDkMR0mmwH/4YXEBMWp+qi0P1bLWAtR03Xn
8bf/kCQ3w3JdAdnrOyt6s0CuIDtcGJNuBtTq64E2P9BRrlxb7n4GI0bWEI5ZIiTX
L4W0Zq0FT1p63qcrD2bcSd5+9maRPR9O0XltGPNRruWtTzv8DbpWc6LePX7G1JyV
Sz8t3B6lTwXnkClgEos/qkdomVCbqHxUIT8L9HobDEc0UImTieoUGZo4HxsjHGm7
V8yc3XwUDNOGnM3MgpqJx860UMllTmJYE5yzY9ELAF4Yyamkv5j30bGl+DN+mfNk
4jAuthYmvF83+ibKEG56cJKUoQGTZPe6vCXtt97v+jMSiBk2QhVARiNwBtr41NLx
C34PAqIr6K55fZpKG4se+yL0MV+Yn8Sw2dekY/ABnV3tx5IO8QD1f7aJNVYlcLD8
voe4qbiQAheFsoyvcq6Wm45EKlkOirVG/RS5c3MRZp5qAwfvhw+4vfDtd2rqM4bX
hW3TH77cU8qjuDTJ0fInT+bNFVtZ0NYc5uaeK8SxElwCfw3AoW7kF1q4oy+zF/2Z
CiYwk859cC1TOzmAdlC7NwUm5CUcLqmWSajiELE4bo4qxA5rmXSwB+QknfFfLeL5
8mvvSsmIil9GCTOv1i9KsSpZx9OLFN2+bEkcz69DkwTSfwfxYBW/B/B1UNEXz4E0
FIsK5tGox4tBVQFnvZZr9APEkaqPKQrK0OD5B+CssugIfT9BfY79reZqGhyDHJti
KsJEbGso4wBzTJZtcM7xEoF4NeZPh25HU2sqAuSWCyOJ6Hm2iMcVxOGv/CRvHI0c
mO7yDOfE5CLTWogiyTBT+lA8E4xjlVC39ueepe1Eyn7n27oroJUDsxct53OD9M8R
vY8hFPiuQW2369JsdCwBsRt9wJfn2spngqPpfMQ/6kGFwyRsjmw7hr1vShJC2UUV
N5NhiAq3ldbLarNeXnpPTdX7FJ5Y3Jd1DrNl46tSeWGEMHLGig3znW3DDLHlFL/X
CLUqulPSrJg/K9kdcipSt4+rk6SoSEZbn3bZ3egu61DNmvWlz03JSs5/nM844bTW
wAs37GFiGvcZ3A9ZKTOOdrEvRAoFmoJer5jQrxQir/aiZyBuczKb/1NnVOS2DvqN
4r5m7mq3avNIH5riXzaGWIVDN8ZLJP0iQc037dZZ67t5qbA7MYrYgcD+6w/hv6F2
orsARwTeEzsMIPBuJvxUrwDM5+JhOkbTrdsM7R1oPrFImjydK0ThEe2cy+UCrAqD
DZsnxIp/2401j8dGMcvLHrw29UfSympNeUzO2zzNjWqoyzm9nqby3jrR12nh/MPJ
pvM5L3sv3jpUFWMOBaKghA+PCydxAXwfnas+p979PttQl6q/VSmSOMRqYq2++15g
2CRwsExkOxwGI+EY94PNBGbs6c+K+rQElJotOwmXqNRPt6580irgjNY7fsXCLMut
ZuP6OgrkFtZEm9bpaJPAjnUNAbLt9EO3GEGXPKxEUKJvou4WKqRdII5oCJ9ttWE4
QsNcbroyLs9WJ6swYRTKMvMdq0WjloYQ4ugAJFkXkqCieIibMwAPBpJN4UKQ0m1O
Hfdok/PjoXiWH2KLj+ElvPUMJ4qYrDeGvFXMJpuz+XyMnMiupeKndYsWQDGYEiNl
kAPqkdvcHTjPah0JFoikTevNYHE+H/KmJnfvdjwfZQmxk/myRyv5cRF+MDqse7pj
TuLSBYPQ0cw/Jy80XBAREaamEHgqZYGYtnmafP8RcEICEZ+6cXnTD8NBKJBxCI0u
LJarrv4e0Gj4e2ATS6J2FY+xHc8P86b2tGcJCvEkLPaTAGBvaGMiGn+p+5BD2LQr
zc1J4sA8dCoURL07SsO3BKxHIuyNgaBgiOmyq2RNgxwpnHjknfu8sASoZIIIoKYm
uMG5qpjAwk2M9MPnR04fhKyQbRpItXvBnGsjxrvhVUIQLyZS75oUDlhcI71ko5Kh
6RxuvUaOuYEfH1zQtkYbw+t4Y39vZpoFZXrxwdUzNVcEduIcuWTDBeH8dZS8qnOv
3dTAv/s9l4Nes88liNTEbz+RLwByygCp4iQggCTG5tgdMI4agCqLmzINM1ZwhYxf
KsBfoddbN/oV/oce/o7mm/pUHmIwI3yNqV6v6yjFu5mnT97NLqyaiUKdKkirWOum
Frociy9PTDdv77IIVh+/l3+i9OncWo/ybflz3HVVo+KNgFpUlf9Q7962VQdxST3o
264y6AOaSDwLD0OOSnBMS+3a6QzBuHY1EGHxf0kOrZoiTvCjesZRAJVdloP+dZ0D
WdncRjCyT7Ny4yGDF9r4fbEi5U5YfzkzoMyZQluKU0HE8jU9rUelSWesMGBJgxdy
2e3yn4g4HhQCwmbkgBTxdKdtBPpaANs9cV2YQF73NelX6MUnwMYIY+K29l68mT15
j7HZjoR54wDwFpiy7x4582O0wOpuNsf5RBkEJ6zpAdyPYNeaOcxyyatkyNGSDYAV
JfBFNyKk6qGXQFcYJR/KyryVCIO/VCu1MS3IECTEwK3omeY0Z50L+hNWROlOgBtf
xFWKVZ1ss7FLvEenvTFFLZKpFc3/buR+xQJtBA/2l9mzhDkkMwQX4WSSx4amQQ9r
3AXm/8y1V04qmD4JPTQAVocHme5kk2x9ffdKhii4MKkVsdbPX16vjvVBf1VoQXKX
KmG7s0E/906ZoY6K99zVV7tp6JGxIU/ayxp+ngn6An3cWm/JlCvyyYi9Si66EPEX
x8pXyLjCAblms7r9UEmlpjNdjB7bU1jxlHj8glFXct6xb+42Zwtjnlz4iUwvOnUU
smQUUm3hpnX6yq1Dvlae2TfAyvig0f+MiBFTTp0qkX3cJ1jDnxQoCb3p1KVYhG4r
VCpT/v1ZClxswiQQldo8PfxwNmoDE/FbWJx6DIjeTEskqt/XnMGIfOzQMtsyGMhu
Dcq8mUFG3SpO0LDfI2NUr4WyBPRfxD6reHmdWXoteFDHLv2jIYdy1lTRIIkglkle
nK+mU5TtAgZhrPAHRDLgXvWKsjXfUj8w/zFYfp8U+qY+VDgzbq2S2UYzgIm9BMYt
NnjKgID5zFt03YltKVvrKNbeEVPoiOW95WeoFoaRFz6v61Uw3HSlekZZTT/jIhCP
Jma+reuzFpsW37dFiH7MYRfEMF3aBhetwqzeLLp1voQPstQ5Govn5DmZL+oNSJeC
DJ7Ho9Z6pE7pH2fL0xMY00goCuCLAL6apOb+vXI+TggRuWdCn46XI27D3k1H/Jcl
D8SQlPJNzhmW9AdTT3stN7B6AfJHyWu2S9QDtmKpwZxVOiuEegsJ+aRyC+kxw5f0
Q7UhKXctWwbICpPGHWbGxOezRM2u0olQUdChQLqzU/6hslEB3Eb1BuuvxVD81ZTC
AZmJRbX5tnCFqVYP8aeh5ltEsgMIxRqxFW93XHHlGNoDHjvVGNCsjRZRJCKZ2ZhX
I7mcpl4U0fNl6g8CI5/jtj6kdLQgF7+OdentRN1rSUMU8bSEY0AQOuyt+k6zcjqF
Uy7izX+2HmMRs88Cq+HGBzHG+1K1DM3mzD0Qd2xJoNdvgO9CQsIu0L4hVaUcfwy/
x9rk26J0JJUvGxgONX+vGPmNP/Sq1ok0jVoIbKmYao5tKfyHjLLS4RCuw6fCq3Up
GQaD3hjEKcE2yteTiRz5t2Hh6zx0KK6RX76RQ44O3MKixHc+wy+wsS3+K7iVrDDw
rPHq1dFzpAdrwSRjKN944OJ7SMrYcswA0aNhrGcPbmP3Cn1+Aps22CC/yr3n/tlA
gEDN36S45srLJrxawCKpVPzx4lXhbz7jVHoBMspR6ujmOVAWv9kt5sW/VYEHYxbD
2vEmv2c37WXZgIeaFIxFuLjPpAvuOnERNAjAF+DY6D298pnGfZ/Dxgmslh5XCxRH
W4RcP1P8Js9CTjRA9tlZYlduaouvg0+3ToxFl0hFKjwUahRUkVHBezjAzjfU1tSF
phIwxsLc/dUnzz2dDtrZ8E3Gm+t95q3ocbe7GOqiYO2+EyukYxTNwUAngO2+LXIV
SMKIk3+6Hnx8DxvrYxfpdXVAl9bsAvi+AmZp77skfYAV7vmMxKHaV7nReR5+zV+l
n0wZCE0OKhZ9gTOJjRlVO9es3C0RFYnI7PlL1wFhWS3n7+wLPd7/mYCyzKUjCz6w
rYm45yRjQ1xRD2jVkvw2+/R3XlXHJ9ve4h60CQn9wY/3INlUHtNlwotUbAOwerYk
OZ+7OCqw5vmcM3cBOO3R8ahI59r22MQ1Sw0jj2MAhXIJ0aNSJHnA/EWss9sFvKZh
pxd2+c9Hmb+mL6lT3OARs3Hm3fX8lP8gbXAHpSYu+1C+2U0eXjcSEzlgK/gqgu/X
jPvFb73K/q5Q0aIhhcgv4otnZzVdHpbPjULg5BbMpBSybezFLa8cguea2RBdclop
ZY8fqyGrXgJipWxRE169inby3rHVysr5WXf1Gz9nIDOp5J3f+Tp+F/hEfujASAi3
rC68fqtgOzXFjFLgRm9PxwCxohztirqsRq3ycTZ1j8h9JE4gRO7MoWQTCr1TLmmo
ePPdaYWtVABX+DQ4k0KYk1eYPnTEJmgKHFqWLeTVp6LCu+hW2cdky4XK49mmKyJp
JQpcihYHf0kQWato44nIHz3u6TIMeGXYIrrDHyyohyryv8LouXxE63SdDaKcsFaN
TPYd/m+8LN2Yd57xlrxTtq5Bx4YQ3SmVk6XfgTT3Zn9/PiY8t6JtruwnoeOzVHhS
/IO5vjep+LkKgg+iE7BkiC8JP5P/K1pEgG1suRUFNEAvi9fKjTdu12EzN9d83jJw
RwJftAnPAym1vGcPGfKLDQLpPou0whMf3ehnkLGxYPsIqLjxyquEgFxhw1vSGzMB
fAcTvHWp7minlC6nEkp+4LxGKTMBtHGeL0Z0Mt9et5gqHUgujJ7dPT0YrJgtZ9H8
0Bk+sr0yo/73nCOURdikXSudrr7sfLe3Ei0w9ROWo8ODAyzvSsYj06WB/DlFV8pn
LsHkzvaoWl8TkgRFcUgE7yvsB60+C38RFxGqT4vs+H1/giC21BaqJEn4hNHtO4WE
HPdtnUs7dzv6EOERchqMXNRLLx0xZKw/8sa0iHrP+ntvF81p3BmodEgT/cfb6E39
OpGWgE46BwZCdPKoC5lHTmgTdev4+8Vb72uOhw0xan2+4a6Cyto9NVM+RF/zKzjO
TWMgfWkBw/RSISXIAWJchVmOH1LcirWxYe95bUD7LHbsA/SmqR8ytWcbt1vd3Sl5
IlNU6xpxhvrGsdqvgfgWc8j7Ksg34noKPvS0851pd3/k+L6ILPdzLbZFGLPGYoXo
MpkjGDyavY5J/E8QTkhXlKJm9XW80g9e1dlZNil7L3EMvaPhAPv+rokypWcSlb6a
aR5c+SbXiFBKoG8uL2q6VguP5ywgwoZuk5mn5OPaAE+9ulbwWVpdwjoBOQW9iyS0
4365IqPwp78EaR/8MGXZPA/KJiYTZX9v9ADaLGCStaEWmzOLjNUAV0dWNF2qdBVB
mr+YNBF6HBZ7sCZUkS7ofz35aVxG0O9ujt/wouJh+/vFzJtUiipGEe1lfkCyvft8
S9/vp883CTDvgn08fMFTGeobiYO6qmEV3VFFX1lFp6a7iZgETeJOxooaDLo5kwpG
2+T1Iy/BI5WARwNvJvXRgwxWxTMOTLrOJI6PuYiC3r/uWftry0kgsYzhhu8aG4La
acazppHc7Kyaprwdi3Kg8DqMuViWejsKER3dh7OMCNACilncFd2OY0BMOav2PH5+
IpWiO/Cj6L//to9+KaqW55hYGuPG1GecK2ilByAemwT3MFZdSop/KTEriBa8zBah
F/zVKkLgGTt3rz2G4Z6uxL8Kc0nL7rzbHlM/z8eREr4E+pUWbXGnPmBgtNB/lOZF
3/A8PvD+LNt+pTxu5+OjsjRbRJJiECAS5ssojd6Joi5zPyE+ptRtcTI0qJWtAa0Q
M98fqYvkehdHfkL48/tHigHDmXliJr5dJN8VbzucwRNjWvQRTAXmqwFD3RNULU31
0E+ymJOo1to0HycEOtQlcAphQR/AkNuJ0W0djA4W6tYIkPIDZ5oaQtic1UCnEYCE
PenK5CLz4P4MwyX3MJ0Qp2tMbO4WFlaFkUwpDRJDzYM0VtS1KYmXIYxWDSCyjVbj
RCc98ZtPLFBLU5DRzZpyI5zAFYlGWwDwrgQYKFqtYVJxpN0NNe2xKj5xfc+95/DX
17cfoYVV2Od6oHTrap2+xZloqY6Ajmvnr/JWyYfy8SIEHXF3rQdvL4xZOrhnc/EI
wl/IHqMa+B8pt4QVd8R/tm0cNZ5VHwCIvlF5xSUtBUn+nlwXh28Iu6oFSXvXNmHe
1EFAigVOHMmo7A77hrhXik96Ptr5Or1GNV8hInHMlVZ2ATKePUrYDrumo56LGJdV
j8Nk1bKkuiA0jS2UbSFv8HepKemgNjJ/xeaZgfpzEoC9daMBpIpy2w74kqnpvPJz
G2pLUjvQur9jFvef52EPMKFA+xwcCCJ3mNUz6g9Pu209DvwJVjBDe8CEr8W+cpfo
gnQcwQWOltFro5G6vSAPpRT8E0cEC5+CKsOJMDIyNwR8Qev8lanb2I2HuLmzmwrw
c+/TSBwtpwjHCDIfY8THCc04Pw0c7WEDI99ZXeyE1g60J2mLSZmmLiPQdJmedFPA
frSAKVx1tj0vogYaPHSslHWEG+U4zG7s/ZG/qzfgSJv6p+pFomVPW6j82az2/XZK
P7jahQLC7pG8YspTXTC1SCvwqK3EDyL0U7kweCVo0e83tjejuA8Z17ZDFkAmh4sk
0RdnHJqShHzDdXMzDxAiMTA+YxquuJGbaKsCVCoIgrIzk1IIoEsnoQei5NrRqS1K
xVY2DEV3ru6gQOm9NHsfZfu/tR7Mjd2DXmUXS5fWqIOHa0aQx2fm/dFgybO++0Nj
lxrH+JMvlEHZchl7NGWn/diRAolWPeucIfE+II5jmF8fpi9Zj6rH8qBWYh+uhjPx
YhOYC58huI2XNxUEAxcCl6JTR7LUEfERKGKJN1N1GGuEMQjyGGXFIFa91mOCYZyC
oAF46e8PKYcM5yo1CWelxdMJaf4vTorltnahezmBs54wNHcq/JrOPBQBpFgtKRZU
Z9rZE9l8h5B6oVUtDkYVDNsidRmOPHRhW8kjgYeX7k914Ue9brXPUI1vh7du7tev
YnhbokLXXgSXwOBQG5dQLAgo4M+72v1sBYOAijUEc943QiuAzElB6iT7SJ1GrNJ1
0sSY9rcKg0h0rMwvzP4HU3GGIVGjxnCa9n4fn2dM4P01hQl92WkOnNOE7pPRe7SM
32/r6fWORBVEo6nS4m1ZEYPL2mRRIXHHu/MYAqn9YMpecCtvH6HSZwBvID1Y1L0B
yN7HTw7LxAmPSoSHMkP/BmOtjixzmX46H6ycPScQfu7IqPGPWir3N7nwSDrW7haU
bDp7+eFOrlpz+razX0ByOsCjZVWnCaQDaj2EhyG4qKPNJxJXE3PFfp0hoFqzLFm3
Edr94pFFFt6ZMElkbvkjdc+iCWmKcG8LJIsJqfU2IWBBQI203EKzsZhVD8rJ289x
wLd4cJ9hH6IOsuiKdTBahe8frWxYfs+xrDd6asgcAl7CV/5g0o1/Xgt5gZF9c/dZ
PCo/hKVyeHlxGQkSvPGh+t43iyH0lEaEcRnbM8SpZFUfL+w23v1fiWsvxhLXXDCO
uDo1gyF5Eq3LjR52wIrXu//TqfJNflIbAD3eeandar5GHEw5Mvr56SxjAQ2kbGE3
696Gk8NBv+kLu/8lhFel5T7lOMhphfZxv4i+XEXv1qN46Jwh1fmRpGGv79Xbd12/
k85ICDrWSWFqVQd/bGOUvjOKuonRaNhB4w1tFQpXbNwrTSwuiGxfDnDXLYKKH5wm
0b5xlzqZyaheNqY5LBqFKPnS7b/rdG1AG57PS0W8XwI6ttuDEJ/o3tIIowu1Fuim
uK7e/zNMS5BTLUVI4ZAMlNYQs7TwhxhLqRLWJ9XPzKE9eAQAy54hFegEcqsBOy/l
KPNipM4u4wGDPB2JbcG2/TGTM57VBrXluFnIswHmlZwS3mqbypVkwtOrS6AkQp7s
mgzoLhXxrVu+DkEKETbmDCKRksfiDhnMirREJD2kYc03RusIVLLRNyBFyUwyIFM/
aeRmAMIZU26NmhjEAHGacIlNmAmqQ+4j3UBqNknjQ+cXlopp3+IvyL5VoMm8aGIW
qcDEjQoGL1HrhXGE7wEMlMx/JJ/j69d5qdSu8wLs9WSuDFceNxfM8rftHziHVL+G
wnQtgNKVkrLk3IG0tT9Kbi1hAJXo7Pj4rTlEj0mtyjbckFSVOlbt9juRHhoKzfrV
qPZDr1LyK2ZExqEEdFCHddRX0c3yfhOSWwu8XWUl11+odDbnKwsbrQElL8J6eJwh
vhwQiq7leFKJvvDb/9/2jF8ls8S0fgTFMTrNIhv7SGvsJFjRoMRFmcvFCyvwJCxH
LjwDGrlvNFZXnvqghUxfJqTRcS5EvAqXmWKKXBKwft4Avks3r1svZhmSpzR8T82L
lQ/qYZ5wvqqUwv+JdoPZbbSlD1pHtx4lMYlHk0ssLPgV0IzdUd3IiEUCn2lbyebA
P6hF9oQWDHJMRcGqBJYWVsIlYahyFO6pp+lzmibmFejZlgvPVRnWCxcScFVVp0aB
lOMwDm6JKK33Q4B4p/Lu2iYQWiaOCejpgbr+QQ4HUnOQFA/OAr/MQnh8ArYB1Ml1
VxyTB2rS4ndSnnjGTLjtdU3SK4Zm0BQeWvkYOYqwHNU98L+MeXnoODNOkmLYyvbm
WY2M+N2IOu/EkWdX3A8b3qRWCDrsDJ/bf0iA3J9nuex4tq4sEL4Q7Y1WyDwRnuxq
m+lLAtP9HQREPNrTuGucOF+G3c4At3YTXlEKYyJmNPqL9/U2TXXbuVNAxraB4KtI
4c/I+/BI+eYMBmRPK8NDicMlcGJPTcdlxMDqpV6ZJrUgb/5OrtwXzTlr1Pr9KIYb
SQm1uUUigmzr5Ym/GjCEVq6Q39mW/XEVj1AuguYne0bLr+CwUmMp+4cz7MZJeURe
F/dlqiRy8O+oDepPM34k5tJVaj/KCkO70y3M2x1VM8AGBKjBaNBacIsTIOz4lsxW
NsmyPYl5o1X1eiZxZwvuv+710WBue47nbbTLDKv7KcneYrGPA9S1Y5i0XYlyVgXM
ZVNm/AfbVFIhsCO39JIFFsm9qRXPKB6nPfMiAnb4J2vQICpbItHqIyD5oFVNuqDA
+aAa1G14AmGu/60mCavWfOPw7uLtB4w8fOgDWCvBkc6MOjJA8YPmC+UK0752yqvw
ZqYkOST50OgGYth3ytYLjDyhjKrc5Ie1iMN4kXXZoSP+pxl01HMEspl4vPBtZO57
M2TiB4eX+8qbAjSIS5MwyEB1Ig7lOZa0hOa1yCAi0elOgx0+jvPxAmO8PLvZQ5mA
UPC7IigrhCDKk9tRj1xPOububYJaR04I/7BkGJvh/zFUjaNG03pZVgZ+ZwHfFwMa
MoC5CGByuILOixYiOE+9SJlsFHdoKDQXhCySqtwGT867ZgEySMxlMrD+vBnaB0ji
xTNq9jjbIFFoKeYeqnJrx5P52BqOg77MtyD3rRsAg5hqh36LeTNRyvMy5sykYg1l
MhJGGntc+T2dEkTN8rNfIlCTH4Qx+Id5/+xP/iwZp1t6GvfdIq52/YxnNeG2iDYY
hcLXm/yg+EXL5311zCGNoP9la1e762bIMvmP+ZqtpDl9IrrsMEL7Z9rCbjUe4P5+
Tpj2YLpHfkTEQS8c+u0Q3OmKGv8o82oibaImimVKYSqH/tAakQ0UCGe13yH/FsvG
BJnnV67NRovupkY/q4f75IaoENy4e3RyrBOxiSFBIMjOM+vAdnNFroTJKOVni+e1
/qjyLapUY1WTrKddU5PYVwk6oC6ECibdyCdRnbMVZITRWoaij16tD96Itd3e9MFi
fxQfrp9964VfrRS6o+qUZT/vyFbsxqUja5fBhi4/BdXTyYpUy3PQISN6RYbhfVkT
sdgctCGTpl/Wa9eWzRXiB1JgNGtjqgNC5PCBptI+8bcntwrqHbAm8N9iK/yYdYSk
Cn8cuSclml5+nUv/ajBxzxGvScCo7Gii4uDxhx4v63QMDZufRr5ZrC7pRtsUHeDq
FRaj4rQ/DDAl9cpUNQXZvOxmtWqpeIAu6QsxqrQdqG5XbkMVYnKyGK80IplaOdCm
PX8EPkxBf78zsQF0T+fKiJL+vMAWNWNumZrO1vwrrFP000KuzEdekxTVoNw1h5dK
NYESzbVVo3GtdY5POYjhzUOgO5dzCmfNjwNaA3Y/ajxcPydm2QgMICIXufcql0V7
aOyS0fQWiRuIYW8RLsKdFgHWRBAbrO82+rWfzdB+62urzQEemqG5wI4/ZbWin/r0
+BfNVb7Q2Uxnw7uon8uG/d6idxYmhXcFZ2Xa2ct8OP9WB6UTWxYgrOnyuHcjeEgN
bIYllenfEnUr8LfZI+TiReUPW55T8msoIiPOFdubtZJcj12aMqR7pM7wPYLRFCIX
paSRGrtCbclqj6gh8sAcz2WrE5xR7zxnhe6DndiLt5ICpJP0K3bSEjl+buuZPXLc
P7hQtchm5oOoioc54sgVvbN3hEBWdfgMLWUZcaF+12sxObaU7wIo+5RA1r3PLWJ6
KbnXM9+OzCxbIbNQU//0IzCzJVg/ktYpfI7u5ZXwgPp8VrrhP2Cotkz80pMXY9l2
z4zTkVknZEDOP4uBbsgOx4saGqSxeI3qnIuYcm4YugKyKw7k7M6O778MXbenurvf
D2jKpLxEroifohJuoMoBunQyIIAlFiAvjgn2dpBEbcE5V1fQvaxizBj4tpOpg8rI
dhGw3Vi2JbrpgDLcEdGoWJYXcc+6OLxH0QLap7OxmS1bB4RihD7aA9RV33joR0Bl
9Rd25wXF7b/SKevtc5OoBmYUBESnqUd6u2FBAKTZHsYT+pD9oPMSlEpABHB52k+C
jec/DarGs3AMBU/f1+qoB0R+jFnwyFhH3U7FuE9HPybx0l4Kc44UorzPMZbWY3xd
f407qUpktaqPXBs31p7c7eCnMH6FU/Ofls53pIOs+43CN/LCLObC8lbYr1LZp0nJ
XlRNYjg/aeHD0Fq27okQ5OF0JiTdN7CqvBq/sV5+b0yy2rPXjZbn9rTJERRIV7Ti
6EPXBi5jRm12LdKGov/pC2WNt+Ftd1TI2Epw920a7cbH15YN93TfYqfzkOpBSHh+
Ra4T8KGeItFcHqgCtd9lgXYCVnGGLkQ5E/sWPbpH2eVeTcbaPOVTqwYcEoWwqw7o
4E5rbZnEo0TrG5KVq1rQtS7w30SynieRtQ1pH3Lw92GDgNF5aWpNC5TDLL2rA5kg
BFoYLeKWirCSGShUuR5qn3S4Kf4B888ash7VebFM/OaTB41fn6KPH1GJUcFGFJcZ
/25VZgQ3InlFYdOVW+xfpsPlsHyLHtIcwiHQ1HiUpTGvP0AwPDjefq0L7epVtbPx
Wmbq547WYaJGtpmKRo8unga1z2pVpfn+itpJs36gUOx0+97ADj5jJhhBkiNs38GR
p5BZzpQ+BCUgTzgNN1F2XY45YGXSd3Uu5lg8Evf7S7xdAPVbfn429/kySg73ilqn
wZzAg3MM5P4bhWHPzi0kJjDiVnWoFX1Y2AeDDIxEiJdSYxoSna/XdILXZd2sd7ot
i6U5AVW5LqvqfM2KukmZBDe5RqesD19YT+jKVAW1zqF0DQC7XN67dUphASscMrlG
twahars5ggrqQ+ClMRbvNiR+9LdBdkKXOjyRet/YhhpZAmuyXE8Rp5ManLdd7A95
PvuUN/9y1PbpFDgd+DWtzSRrCGX8I3pBoUt0y1Yyt8NQoQsM0wclbpvNBUQFIlDQ
bjt4/xT0x/wLpwQkePysA1uaEoovpbZjn8jUteq3OlK2b+qGCUHaDY7Fh6w2FD0/
bQcukaEZN/1NELI8m3CRfSVBvoNvVFaPRCjD7UtuEgWa+z9YEqVcVDXb51oNKanW
9mbZAZZAzwVZuzNxwFGHxSl20wkyNVSJ1Ir4XElCHPiSdJveP+MoSKa9U9JYNvt3
LsiiKASt6nw7tnwsXkoTCnGTatbctUdtoGiPLIrfYRrRvd1Nzgu0ma4xCJGrrWAP
CpZOI8D4GcugcVPOExdT4C30kHirSI8aHHvkvn/0+s6FQsQ3eaxRbznlloiyYJTh
Qx2Ls8yJ5mNBrcSXgpNLXnWZ5LjM4nn2Kre4xsYWKgQunGaXQP+zkwGwjBmmvuZD
B68JyLJWKh6DHn349FpM1IjI/PuWh5xb8d7WD6kHmLcf//HNVYOOxPma/O2BLjI5
bSsY6jpa1r48JA7BXi3+38E1lOafgMGM+N5D9vafKd/lHDsXDu9vQot9wJAgwSBe
1jr20IzIz95r0oLjwUZwI4geHMWTZbQGiPM06PNDLwGzR/KYHiHlws1ANM6qzGS4
I/kFhy6F7Cxz/tinhUCITAABAZZ89S2PdobioRmib4Vyfz/SI4/hWMHwxrUkAtd6
btZpLyKSOWugWyfqTKsmmVAHlNraQ8CAePuO5ep9+T8RKsxtcZNPE0/NmACQZ83b
mJpVzsqOWHeeQRfsB+FmbvnwoiCaZJ0CUC0lQnvY/3Qlc5tNx0knEG0vggHaOTz/
Z1blgyZ9qcE99oTsUGUsqpkabkUVia6xINaLhF7T0UPMkFg5KcIwbldEYkPHb6PK
n4/VujfHXKUK1LGQPQf7MfSNLlqwedtM2bApkvzesNQgdO3pl0ojzABF+bNso610
NhFPzbBETNtJMrhhC0uqPpttW2Jmk8bG84Jo/nCVTguXEKEhxGvhviJiFx626w6U
NOFx9rZQ8PpIdpIlzigsFMJJrVaEDrDtD0cYNUkMotzmtdzmGpjFJLdHDv26Nvqw
wh6tURD9AGjqdPiNBjD6PCUiEtodtckf2AmXOwMWpc2DBdCh/5kO9sVcN7xqHMCx
1zQYnD+h9HE19ovl/eELR90HHFmDOdnICT1HlHHlc2y95D9yCLqQPr0dUn9IuLb7
VBJpHBaY4qoP492Rb/ug4I9ahSodscRRJjimD2ljBDwKVUx3nH/ZY4wneBR3bZDW
DvQqBOrxLfR28PeS74TON7EmLU8qqqzmCXVm9sjFmnBlEiCLNy5JfQxnq1aIw+wq
dCgfhEjP41fQt34JGzoOVkoOJF2iZGKjFCmiM7MWIfjs+1y4tvYZBIcLMwEhwJ2T
//Thnv2Y71QkqbzbMyRkFMWq4RtR2ikhYA/cLsE6oeLwh1TtZtUzoBh4rtd0N+lg
8E7iFSLYPoMMJoJvj9JLwdBkvYNBSrl3r63gDJNj5pBmktPecP8goBp6Qau2jKS4
Cjc2KBPdh4WBs8QNTEMEizOKXOJ09WBFL7frd5PEWXHJNeW7Mf5oCeMD0E/GWlTk
pKQpxJJPr2i9WjQQUBV3lbjpfgqSWih/8LJFirKL8YZsdKR23EUositeqpD9H+W3
iiOth9FgXBUfF+L2eFFNVw9etdlxEF7uXmHpcUW1feVvBvheL0rwXsz/MeDa++Pb
2sJH56zCbVE+3P+NaxemL7PbPwGSeYz0AFeOvENB1ZuMzlSf7nfk1KRHRw0u/RbN
ZHN64f7r7U2DQWhfRX36MdW1CfAb1Qk5CziCsRiLK3O0V1Td+OgtUmzMT4dTeBis
hIzASiwixJiM8c50cIAfd6T7VgjLMxfblMssS1vWJIW7Q5+raCiOLupV5rjJxL9a
JR6ln9NSJUTeIPKaiS+8ET/l1YNyOPL7+GAIJZnd9+zdQpNBJLJRkQPrNoVLepl/
mmryP4i+1hInGqf3ySOAjU5mnRWSCq05JBGzmX1Ge81sQA0gT8jQx//MGlm+5Q2v
lcDgcQD1ixeg6tYnSLDVUxOVeZcIx5jSLdszIyOae8VQ8oHGBrbILh5bhfsKBUf9
n4HKN8CyqmqVNqvMbEzCvLxE+HfWJ05xtt2xRSSgoZfToAo7F39QPmPNt99pik2H
ymd3JMI8BajgSqGYHjiTUS3DvmETZ7MZ4nNqZD983jHiToQVZ6uHW9zQbk3swmst
hH8Xee5iEH9ot5QntACm4q//YvaOVTwhK0E0X4O8HqWMOECSSYuxlEjI3T1cQXpV
vQCRNXE1Xc5rxJNK7e5E6YuxOu9qebV2QuB1GjsJ3SvrV2TItZKxphX5fkvkxiaF
2aPC/U1YI6hD+KcqliLXI67lnD+HPP36x1UqfS4H8M0EwHMBF6GDq58T2Ru3+irP
qCuvei6nouYY8UX1HtlZfH/GTvLMVGE1oZX8Q+jANgbYTBZ2QK9DvjAyKc4o/e5c
yUkDz6nft9Z/61yZI1zW3DQbLBpHeRtOJyLk4rRg6RxYFBbl4jkhww4yVSzNz21P
FfH3JmKbp6Vrf46UTgEaHZxiJu0att4zUcEYVYn/HNI/juQVEXAvF81l5NA0VM/W
MZ7Ku5cT073J/UeK3Y54e8L61Iwcdwkc69yC+n1vMwxUmUmVc37nR9HosWzogja4
UOTNpNpChEAT+NF+DXZtZ58K19AnAMrTcTS9jYyGsUGT2/i3EVHD6xhKMPo9tFlZ
hNj969j69VTSzvbK54be2jnNjoD9LBDTOiuE5ZS/cvb9CAXZBg66LMg/S8SFEyKa
n+mTE0CgAlo3TO2v26gNM6jPHPxvCky+Omw7qCbHEUFuK3ySPIzajZ1RszqMkJ8j
d1ZR55kH2ZmYrP4X8SZlKhlGVgvQVVPHe7MefyIGzOd92gx9K29epvZAg9m3DuEx
ImDSyClYvwv5rwfCqM6roawCdSWl8LzrfwekixjN7uD7tn+1H0C2F9GslPFTLgky
Hyj8WJdiGi+3ufyIP7bEJJQxL4PChly4GGfWiey3tVMuRVj+bainAp8WWu+Obnc4
FlDiCCE1UVvmlKmiU3iFXa/regC0GUf9xRx/0L1feGWv9dfGETdhbhk5/ucwxgAC
K89XlQKm47w2rljxsY/I51g+2wvZJg5p5YSQFsUCzfyCPCjLpIOrz874z6p1NKN2
b9qaLr6258SOtWzcODFm1Inihwg9PHMz98cCuCcD46osIi6N++F5eOYbeDA2a3VK
O79O/GFJ83+S/H2ORQ99Jv5k3eHXMPsn/7SaNmZmNo/FZ1uJZqiFHKAjWIZUFJNv
PGbTAfKIBWbwndsMFHsYZ39wWoNJJxzkgaXpC5SMUc6gEBsInv7MhDgPiJV5DMAz
uAxGvdUwX8vn9LRlrCHfAR5GIwzaWzPXKMge/Y3q6G0KJSfkp+w14Cp73NEpCO07
9ziH1ww+cuZJbsNsILmnOk+EgzSYFzPuokbwhdW7kCzBqEx8BzBepasbV2SKMOCr
UNOLkE87lWwRhrW+MEVIwcRJrkud85KIRC5Qq/JJdAmrlhVqq0bCn6U61RkKtgz6
y1PbCYeiMMKzz5B22EB1ffvg0/ulM4s41Ddsnch5HDLtcxdOltindDruCsQZKflc
NWcWc6Z2HVjOcCX6RwZszbbYJg1RU35J/S/RZ6s9aqQkVxNTuhDkuJbzIcULE4R5
pOlM9TRnK00N7omeYRrex/E6YsJhowcnVde8ZsMfakXV91EqRzUyDR4qKIkQ5K4J
/G+QqLWHxfGpMBycGLXgRQuMbEeUFrvkIpHIhxIXnL4XcVU/gSa6Gh3E2+oYecdI
CbY40ouAab00bftKI5jtFZ8o5lX0gIK767HHfyp0R12X4e4BaeLLgoDjNOkPzvoq
BqxJgZRmV8wAsrg3CLhYQ97zzDXxmF50z4hDw8Mvw6mC7PoFakWPs7WKWeb8Ap6S
gwDylAB5e1+63WWXt9Pc+MwAvojk5R2QNr/xarcksCRkJGFBUIh2soZrUG0nEVYo
NLlO47T4vDl0b3fSlvySzTl8iFpcgTX9lissXKgtn+kVqxikgpdsQ33oZwJN+EzK
tCHhhlheYB1Vlp30gifmNzcSqMy8dON0QJG2JgTu9HEo5Y372SL+OP+A6lHZ752H
1mUSaLXOd/uqYdbShNIinPTS4eVyJPDmPitXAt4+uMXXp3UoYTs4ewxkrol5b8ML
mfphSjWLcAcN49rE1JPZnylny7B7qrlor3puc0qEEe3OcOYRnBSAUk0ThXg5kGD2
ys8EtGB/XItOR7qllHj9tDT07mEboLmkfyhnPaP+6GAPAa6jPcO7k6v65QfLiy/f
stKduxY4jGsceg3oxEfiI80Woao9o+VnwqM3UUjNDN0P0dx9NKphEZbFGI2pTd3g
tMxFU2Z/NRdN9mNwpnfHrlRhkDjz1AaKoCZT9o2oDUsmT5Ty+SqM+SoS2KdNMpeF
HRHzsQV/QX1c5aun1zM/LKT9KzAlpzZNyzKcnc1rF2TcYyy7ziUHOkGbiRYcqljW
6sfuqTKXZYwDzHTsHHC14Cmulztb1yX623gHX+6aYiwSXSyL46F6mErr+qa02FyF
NoR7f/YZfBNfJwbZFZO9UGPbDa1tnHhKpoJAy/vp32327u5Sa0MBwMlZEP1iXPwX
pzSUIXwLqPt8EUHm9Vw5V5VMLiErdqy+F2DtVmy7nuszFQ7NpwhBVRYpNEzg4Mtj
QxF6AxZLRdY5dLWKs2GvrhrFRwmSBhgmaA6IV7jzfs8ArOOUCrlMEXkzrYLD64Cn
s8YvY2Ffz28EULxJqPtJiNwtXjtosI7d2XqLBIZBFCUrNEf7WUCBa3zyqN0vOLEx
DRhcP2l93eEDr8sHu/dz1mxUiidoeqwSK2VC2SPVHG+HKojJkhzYjMpgY9k1OBC0
itGbPSlgssW81Qx0KKNHW7l9yjQt64vlcNomhW7h3Z/lT/HZfUfrZiW9CvxlBCS+
fw3F9FgheykcO+9BxG6XE07hphgkDsmF9mNUOkLmNFpZIAkgTxJnpOPZKUglzmdM
xvQI++1Q/wd2UK/KA/NQNfA3/SqSx6u3ObRNt08wAlPULzDy+eluJwKWbzT5A3Qe
gq1ExDP5iITccai8oKBikU4DxyabJyqH9q9CDKREDiJf0+d1/xrIUQamsA5qKaiT
g94+z7+adLKUFfOMkLEKvfMuAxbKP/Zxou7khPakh7jkDgJ9ljTj+PAFtgKVDnEi
dUEVjLW13b8BAHOwv2lPlXKGV00JKpxNn4aUypx+D6/y7TpAwmOaXH5Gilq9wL5/
cYesUF07BxD0B5XT/9wG/a2w8zqw4k+vCaLzQLDGdn+PSJhzZog6YixXWoDXPtwH
M9c3swIunYAlLz63Iaf5jF7iCKBOG1DLYIh0k4jwceDQd0AhN7XDA04GT+cFTZ/x
23Qspbeo8R/yxfdbuCYpXpEJLA4rptp3g4I/nwgvrWHViLNShak+LvRD0/iBFyBX
1IGPEv+vyA9ODpv1kFWA2DgHY+Bml68KenyoJpgQoBCVGd3R39U5wpoZBn7v4/XR
h+McyJMe93Hq16sXc/dpK44sKQecpAFXyu1EuqoAUvczWgwsGaF2kwY2BjVsAxu1
IpCS3Ka+x4g1455OyjL/L+lF4nn3o0m8VCSAS1/Vo8u5tyWS5fhAaJHiPGvUnvt+
Px5fFzFR1eeLajAd0bwiko44QU5e37DNXDl/Wk21hc0vCsBoNd2qxOIwZDBXOAWY
r9d/v/9DNWPuKngVnhan2/rLv+nXq5Cpy3Rh8pLz9EevstrW5NJBROg9adU1g+Xr
GEy4AGvvgR2pqtpLxC8PeAkKpW9xP4HskcSk3FMqlcub/DyW6AsZQ3+HEtDg5tpU
DTRmsWUMXOnlhyQh/AJ42Odj5NmQ1JSSHrIyOXGin+CY6ErXggnx2N6yVcCIheki
shHdmxdzje/030ZEFqVPS4dlObWta1eI0hS4mqfY+NBs/zu5Z+8wteGejo1zr86I
1RbXpLIW2GWXULvqXSK5/P900RxJwSRRgJK9IbPN22BBv5PFjqHhSCBB+AZj1dI1
Oz+s7dSaK2mvzA1u7YLfhdvJVaWTov6ZRqkYZOVxp0+ZTdTTmm0UIfOQ2PKHdWQN
TsfbBd7bXykVnxKrzxbgaenC4OLDBgyE3Wup1l6brbGgIx+EPUDs781gP0raxZ6n
9x0zCMyxcZuKC3THoTkqsM/nPc9zyp/yjVq0s6uDBGhvAp3BuZFm3FxGfHRlPNUb
2Y6YZbmBk9yuWOiznzplrxNZGyDZ6h6buvjNsQuWcxAIr4OZhQfzl1UwY9rau79C
26Atw+3exBYuVKMnPOLOkKSCfUNqHVAXQqmoa5OYpeGuQ/1KBCc6U+DI+vUArCXQ
Kgpmh0WgNwmZCZeI5vqmdwkwnn6/aAiN7K2REHf0MRzt8Zn4A1H0rRnquu0cyBBm
l5jdIbEpyjV8Y5AyWazfDuuYP1djgMFk0zmuqDX5WbpIkxhXrHdNL0aVAQ0K7AMO
3eTWh+wJTFh5TisB7bNGFDKWzbGAwWwmetQGLC70UgZ+T7WB87jRtk/SJjE9ldOa
BWI/7fVO50sK7y/nBoTI39imR9c+TATYe+EfIe90IixY1/PjVc45k5KGVDJsOXvt
w7OgtxpH5O39BeuGsHRUdWQWv9WplZhk1/awGjSBYcNo+xncujKXBiQ+NNXQsBa7
SYxtGHGB0+PIRkSEl+URTUMm59Td0J4sEjz3jC8aYvQx8kecBqia/cT7JDJcDDNP
dP9WlVUuv/C9f4UNm0lmaeKO93pU6LsKPzAEbXwihlkxVmx9LM+KSQGG8Ju88rFj
XX09mcT/++QUzL/q1mMnz1O6674+a0F5ihnyNjQaBAichTQ5tRSL1PQXZDHabFEl
zEEXiDsBWOQXUje1rhDppQf7/xqAxQAzvu4SL4PT71JnOHLxJxKGryIbn6E0QU6v
Nlae1P28PUeQZ3LwfOOa5eM81Hv8O2JscChGomtFhJQEGTMy9mgZ+VD27blv/wF2
6+nNvLSPCmNXUTZTvKTmv5qofWdKCp0KPUmt/qRiiFQ8RMjVXJN/jFBBJ6ISSl1s
yr0TwYBzR3qDU5V9Tm+gyRtzBDBUe5SbHT27unFkF0n65n18OUO3CQU282vksSv+
D0SRZiNZF17yAQiOI3iDEB73dzslmqsIz7pc6C6FPROIQ1qY1ImsTK0tTxNfk0O7
C4WYXS3mzuHYY6wf0fCgsw7cdUr0qWf7pBAe+7AMlOPJfoHOKvbxiN7hcb/kS7X7
6Fcgc4BNBAmTknfDDzYPhKamOqdeNIiwI86FTTB9pPMNGUgq0vgiJ2Yj4yIFPqwj
UlD4kDLblDXIoooDglXk/qOv7veWGWaiULQ0IFUM4layZqu6EVO92J6OmjWzITRf
IzKZqzB6hETYYBFs04MQ7pVR96u9w+iF1GmfmyRQO0xd3nakR5LFlzDQUxaHiEWq
gdqXvvBVLAczHZdgEz9hS/5YSIUpJCHmPOhKHV1iPqz7bgDtgV4LuyF2jgKkIEKW
HXxMpk3Q7URpaNg88QjUm2NLbX8zbAKflVBUIhQUVCLx6pt/3eQ0D/veejwpJMBm
6GzziRY2La6Onx0SksV9DTsmEjVNb1sPj2izUSnb2jLtpb9TypqYBw58RFqSsQk0
pJiG9r9ksNTN/7ZQ1mQjJECYNMsYjzTcCcnY2zz3ePFoK9Sj741n8PMvxKdCqna9
IqA/WZFkq6c/bzdk9AdSS/lCpNiQpq6BdxA06JsXNUAqUE1o9WxKuzGHwzyHj98O
MEGbPN7roP2iDAQq0zqg7TpItnuaVb9O9OPPo3R7cJLOla6DbGxI9QSo62IBz4mF
uzdGFVGPliQj89/JhwHfLhx2UGJYiL3K4m/i1Fw3iYHBqAITKzo7m2cFG2/0VFOr
0x+8HxXoY8Qc8jmJPorIde96n3UmARhpHR8sw54QYsnWA7cVMYT0yCPhIBmp9UsI
4JrH/L4Uw2p8uRfvObTGyzfLegaV2f0/hL364T7/qRBI4XDzrIeOdg14GHXT+FLa
rDi5HFsiXc4Rt5wEoghVvVCWSvFm5+OaAZyv09W/rY47sMmFZGzsc7ouWZXWzKcF
xm1r42ajlcOottR+kVncEGo7ZbKkyYdu1uK7N1Zw4h1FRPz0zcLwdDSM+jxfrwfK
X9vNuCt4CBfJ63Fr82WYGi/6wB4ozB/XB8j8DeohEgAxnKqhSOE9kSFWWdgW/Qtl
LahXt6bfbdGDYJBdjuMWGg/9n2xihvr8Q3p4eoGmLo5VShVGGZCM+N+BHloMTjtn
Bmq19GjhPbBf1vFW3TW+3ib4vN9dRHJSYAVZbwReTdE4ZD1eB2h1bXc0LhZQSDYG
R5rk7GTt1++3bG6x4fAqGy+1SXIaDYPC5MqCt9NpYU3Qug21Gux0vSXIiIRyzG+g
iiHKSl1BtIXbBVfm5Z2oiLpB+9VILQkoHzeNLRZBX7ZnaWfv3+IIiBGDIPMhhod7
oT7r2avPrJYNrtVI6v7IZtKQTJvbtrRE7uPO6D9Xrt0oDQiPaU5xaG+LT2OY+xvu
wfQhfv6FJdJcaEA97rm+l9fIJj6DbAHQvBCkQNMA6NSMfMM7kIGpMwHER5hEPf2z
jraG3P2zbbpscSXz/7s2AT8OVHNgbrRIRsI9J/f8zJFgO8H0paXdF/+Nslf6wfHM
94l/bRtjkemUKlk2pr9i/60hkguqmVX1rVCIMA9/H1MmvWDSiD9TXFRqw70nl0l/
gzekG14wivSKUVaur8OrzZWDQ7IlCB6xxe5VQBzUi3OgAxcEam4TDhC25JFrTG3y
04k4PSM+6t6XI1keK470ox0fIU9TyH1AZNfxzQHlII2tSddAFD1tg4RJXwgIlmO+
OHAZSszKG8AG1C6S1RUGoCrzL6qWEULZ9drvV4mpIPKKw9o06YkCCUf+fYUAIkcD
IAJcoqeaXtnHD/jxEiMAiVVkSMJ4TQeJO2A4UV8Q4CJrPmQc6NPscN2XqhhYU2yq
AowHQgRoaynfRIPNdMob/tOYvLGcHWzFpoh7L7ga/AKQBgld6KUmzVOKkPlipM8J
6npz9eeFLx+rhatz/9DrKksibE9LHE+YIk9pEbjToL/uk3FDvWPF2MpJU78QR3AM
Wo5Ab9uQdgLixlqhkbCRG9zfVcNqDRY/phXq6KB7Lw7fI9K6l37YebA1l/djZrMI
tnSX+lp7qvqKpbZacBR4vDci20espxgRw5ybayG0krQenrznWHrAaeTgBqxrM08p
PCDLQzfT1IrBl4uHo/9RmT5HNNFL04I0QGMfjI0nEEWEXx/bzbgs7GG27x7mzKlZ
w7vFxD0Bbnv6DM5AV5hsMB0TPIot5MZBVOyz7O947BNdZO3dg3HBeE9RdRPV05Px
OSJ3dLKfan79gyuPIxL11BJpE39hdk4mX6N/OjrgqPNDOM5o9mvDDanBNY15377N
WmV6T+iVxtKqX5VKmtq3N6/lyzt355sJ+UD1Aj1GnRdL9bEBwPn4IFfguCCE0sec
Irbex40vH5A9WF0K8IwFkwKlAc7CiaBG6e+pKuS+U9AQCmShHdyGm2VVWBPOM9Ly
gCwSBE3iJhEEduyTl/BwNKmznTYy+tU2UuxKY4HWdbBeF6fA4KzvQG2CEn/DRfWG
WQ6DIFibKP32bNFCVwfgGhvw4KzsEWc90wY6K2QoQolwOMgJM+V6W9PMTndIQbq+
MWXLt0wKD3KRPdjypUzOHHOekyOi5SYeI9iebexB18Gi5c7W70TNmY6TUGLLXrTa
x+p9ZEs35ZPXTLHxSsBom94OQLCTksAX8YXSQiprQpjw9ynmkhXh9e6g6JBAYy3B
Jm4Mepi7YTmOnYsXVS8rqtCHMRDs3kf4WKaPj39zJwUq7SoFrLB/jIi48KVRtfyA
S/F0Ai5mvp510NQzxIkC6fuN5/A0le5s+z/GbAXcuZ9mD8GRtMLifRZ/WDvIBD8d
KqTGv7rNyP9XiptphHInNojxSHRXYVxtKMMdYhfasViS54LIgsGlx1gIj79PGUmH
0r/5DFXHiIrwnNG/0FZNSBwF0ads5wGrL34Zy7sSDq8IIWYt3TOxhr11WxV2V7fc
rrDDeIFiMEQgiJDk4nESpp75VSyDoqlJ2/dbJ7zywNi4eZNgTHGcoOSVlTiqFBOI
wzDjeOjrOe/CqrE0k/E0zvU67yqjUhwKmnjMD2GfFIjjpa3CMQHQpD+bz3ZqdQH2
RUsfUf4Xhon7enaBmNl6ce4HgGYX1tV3Mm0HNSSxUwYBuiHhItqr7ZzLgX0YSZ4X
0Prhcpmat9oXbrhFrK47WWbfAwWMCxZr1POBUfFjewvQ0gNMb7/BiP0sCcTe2gnT
ljI9iQ+1fGNZVtF/DjIkvYsoqp3VQBHvT0wx4ibfZhIZ9Y6/a7g3Jca2OAa2jaPz
hHG5InY2SruRRm3+nzsOI7O6kCkHzAcmgMWGUtF12KCytKw+oo9WL5TZ2rgWIycL
KYRS8ttHaJTpUmQXV5SuCUiZh7gBQ9hMpsZLrvlolROA7fbwhIQsvkTwJKvVXjTZ
f/4rM2SMcFjVoc13gnKUhqF8jymHFs0Hx1A/D5ytfDnAW0qwrpWC1+JpqCLbPdNy
DAMs7GbWzjOuo1p5WwlCINwFMOd6qMmvfpt778QIDpzFNQhKlGRUOFFU19Y9lzVP
X5BXWkZsuxU3pb1DUWWviJyv9UKB2lslCKwEe7TF0fKwJGJwXYo+WQ7c5JYnzmCc
iQPOCz06/Uy1Yb4b4hfni2XREgbBOdJhr5HnCDuJ8Y3SirlFdDlCPDOzYOxsZhbI
P9oGcBleMVDDyZOqiClIPMJ9+0Z2pnsuSeivCwM/toMYsS4FwRUDEHI+Y9L2vOow
/OR7rPd39Z5G+RxLkeihyMJlRVAMXJ4uY22VDjbnzygjvaMljeXP8b7P13v3aNh0
RZzq2fXZBdU4RC+lmqBXOII8nkN6gVN+wFDQMJ/09qOfTZbbFvDipdDzshXtJiXQ
EEVqs3Mkksh8hw5pOmIdCpHbamY5GXV7wsyrtpqrlUKOWpQX0gTqWoIziuKTL4Qu
SVUUlet5CsVl/0b9lmfWIVm5mJ3bgBg8OrjQwIFFOAExraMdm3v9fyPtTxwBzN3j
9Jl+YcQv4r8FSwh7H+NX4E3baWrBJM436JaVVe+yut7C6AdIcRDC17V8o82afnr5
hTj1jxZEtwXXY9EAEoITSAlTn6k7lwJ0iviOH7QWrsJO53JWFMYDvTwP3JI+LdCz
u+g8w5wUvEq7UM52E2MTPQMhvZWyaEza76aqQVAKQnO8WT9PGhOll+Dh56naRNOk
JnMmP0qOcbp9LgQLal/kozJlAZQcyFUekQNwyxD3PKH+EgvZBJfEtHhiIfdn58y/
OuIKgqQ+NMvdYaX3RQpuVz2rquoha1lDbSxqjQCc6ENUYLC51tvtZdwsaKvMoWaq
GMtPuYa0SocSy2JlYVJoTQ/5BE2Q2vaoRxYcrv164ixfR4UssPBt6g5D9ybgz9lI
R9v1QhFau5i3T74yv0H2J0vn5dQ+epvN2RH4W2rLbql1vBiOQSufdpo0zcVGDeyj
xmlyaT9rtAog2c+Dsujuyucarr8XlpuM0phPcC2Uc1lgf++vjTOfI8kQlXWMMhTP
FstYoqlMLqktDr1+5tS/HxK/3ujCW7TWB9zMHr7TcOK2nZjFiYrQBJAzDpmSNntr
BbVe/mhoBlfcMUTQicutCjp86IHGOl5S4Ea9NyFPI9kQVsTsRBX+1Q8Stuoln53o
iB0HVm1Xo3h4dPt9YAM3ORpmyemzYm0e2ppWzsgAfKn0oS0jTcY2WHIDmqRdsPtO
BhhUaMSZuuYHOi2q6qgarqlsNIttWZrsXTCitUzzinJZKR7DscHgzXQAndru4S4Y
1e9EBGYz/XBWJzVbIEEgSLTBDsYGG6h/8l5F7gf1HauPIQO3ieZktZ4gxyfe+5ln
Xivi+9nRpX/q0Gcbzt/Fg2ANYJaF0FfF0UuMpCvKK+JWjHpLUO826swbiSmAiPnW
enlarqZQU+K7tsONtxu0D/t9EmBML9Cj7PLxeooxQgsHFv6OnSh106JOik6alpas
3vFgercmaP+6sgxBegVAFaOT86H0WgvCtsjlrUTlVzk76tknaAXf1JPa+QW2+DQm
5BYGJMZZH/yHhQK+HeO0ic328+qwCMQ0QtlDJrnXgn/UK6R98F8GaLDO3CXApu7x
LOoKh8KNw21YhD1/Fl0Pfk1m2htBTb0Fu8W0MKCuwrWywk2sY4HoEwHzNfhutOZD
sra20n7di1hg2CPvxAWGqV4K4BHWFcmJa6VCZ0QRYF7vBpWD8RNoBmF+zajjWsWk
JwWtVMt0XjJ8fdh14AfCjIzNvcSNYQ8SuM0oVrhbYlFVI/f+7kH+LraLt7Epfqfd
27bGbvnDF+ptCQ54I48PQPQP4LKURnPnZIdLcys2zvu/maKySLESVCzlbOCx7Bhd
Y/sZr7JAXbTfk4uQwk28wInG1B0hCD42YDoQKdXy6jk1G8u2nTULbxfI64eguq3L
uzkVaSF79mg6MBGrTCHI2ZNE7jN7I379PBxxmc4WggEt3koVWcKt8r4uhYZy++t9
QnNMAoW/Kzm8NvX+cjTe1idUKZ99R0kvHr30vKTjG1jpEZfD0zE36Pgp7QxcZAhL
bg8P8QY3eWCSznAnujy9z17A4mOF6tawFHO0v9lUCgVK/1eylDTdLD9+SxzVf6/D
zFyIrX9uJ8vAmKh68uXEYvbcwurKubLJz37MFd0PNtGuUFbe66C9IOA4/gQXE7uU
xKyaTPsgqKqSoAuXB+gPoERS4QE4SZBoinJAMyy7ciCeFgsNf1tfo3cP4T+acGZ6
QSnD/4lbOua50R5OOQ3cwh9QpZBEyXb6LZmxsHhK5w8dHJMfzhO+GZxbrC8QXVog
NIgiQmwhQ2alXBeoBEN/ve26+mOQ89UdboNA/Dp1rdPTniHVbKlgIG5mTd7HwgSH
tRL7r0q6Nu0DUNjJiJaqwa6QNQg1G2yc/sCdVhvwzh4+jtFplaKr769E6orkOUEQ
7ywhuws/pPWamff4TUA+wO2gGesXKjnqRInRsr8wJo+te2HDDAPEygVMlPc8aZxt
LeGhYo9WtznRz7DWC2je9n1NrH94lSocunYFVFE8nu1gITkNQnBGuwY626Mty4Fe
IJg3shXujv0tUI2JVXikXO6vVB2M5m4N6hrsZbe8J+zmyEtYKJ63C0MRS7a16iii
SpY7QsBTtGoxqHm/avdzDTHoTvcTv+YRRpscLAuW7lWmlnxvP5IXiadxnEeR5/Dq
dUv2SkSHKmIQoqRjYnq9PwcgYsI6qF4m6LSye0BBLc+ynaTBBoS/2zR5rlqQ7OA4
Z/pQMgH+0bWtPzqdhwzlSe/mAT7MQS1acx6P487F3TCxpSeb/o08T9wnC2Q4DRBb
0EX+/+CAEAPU1awVnGDmtCEn9a52up49qsdXyqrIcN8V2BReajXRGHMAjw8LiYxe
9EeqNERO0/Y1BzhB4UPkt4T0sfSfjjm4vbJ6AS3X0W0IFb2P/QzZHwflOQyUXrmO
GZ+uZL7s+UW8Go6xF0zX2z49+azfwqhjWTho3kUoDlEvSEkvX1V2wqI5KDRMd68s
qkh9lGl4BxEPnm0++juCIwDaGlKRlkQ8VsHoEtGLPj/ju+VR1eAYrcfPC35DGNbj
FQ056t28cA3ypvYY/aTgRW7AUQ9PVP6ExptH1VOIH/uf80RHtsB+3ZsuqUNwGk06
ELO7MKeU+5n8Q6c0sKg8CjqahJx6ddv5Mt88QFSyyPd/5kBdddtgq1WnrNPmmAxw
w+gFL7tvIEt82ZlCCAPa9BTwBb1E/RFB57xwOsu0za5dhUItEZORTdWkQHfantIP
7K6xBNOTDFQSSZ5N7k6D791q7Fe6xxU4SD0NoZkzy8MAmTbYTqgL9V1cLcGxSYbg
HlNnOGlRLJAXcq8u+e9SCa8cjcZcE3kTzV73pJYQduvAdG5/Y5HYCioT7q/jj3Jq
u2V0St84pF99CWAHjVmzxfoRFtC3lLs4r24BdhHYsb50afG27i+eZGrznyV5fmp8
BMvZdczsUtxU6ekHlZykyefFGiRz9w2XpTFulKVDrNVrmOSgKTmx14pSOwlf6/50
oWg46uouyJS/iE8dGv/DwoRZqLtTnoU8QzsmyJOeuKLrsDbCaMwyZOc+BRKEDJnW
T8OH5oe4llPS6Y9Y2ZwaPFAPFTNJTSRWfciA1o6JRmgJA18Iu1bsEm2/dhfFtutq
Vo0y+Ef0ssuzpTaol7hQohCVsIwYODEqlLIffqFNyVam4C6QejbRshkLB+54hYsE
5XOqmr/UbNj3CN1YQQKDQuis9Gnsyzb82T7uD6MXWJ/I+fEvXlnf4zB+hWKoHUIC
1jwHjGN0UBcaStt5Q4H4xMnikc5QKXuoi7xs4fHBrtB+R6H6dyBmnZzRyoVboZq9
wtGGBOhYGl124VRfqbnMpeFKtZJ6hBWzbOFDP+jPNs3NMIX3tQb318UeIDMYCFJN
PzoZtbd980lQPRMTqlwMCP1WEU53LhCsna0sleHeg3DMBSnacV1onJ+UJOpdqXjq
31gyriMMfXaLy85RAIFkUzreAwLP0TnXeIpAcdynuwy490MmziecmJTl0MnnC+vx
GkPuXiazgmaot1bWmAE+rQ+a6QOEhbiAi7loQXppFmPFr4BxMqpkOPpj5k9uccc9
eaxu5PE3kjjIpjaWNPkt7nnN2CuwQ25CH8Ekcv4yceHbpi4S/pIx/rpjK1lHseZx
mOe+Hmu/wS8uzcOyC9PEnjDXfsaP9l/vme9sTWBcGr6JsYM/mOm/hoTZPr5Hz5Pj
TQXAmzpAlYS1fDzTfOfGim4622HXJmo+tOSaOx0A9GlqtUIW+Xa+xGjLUO2X2GQD
OdbIokveJc9q2C9tI8Elae3WEwK191zO4FsyHxh9KHO1YWRATsXK9Hs2yeXlggQq
O/GUL5TfqLK1PUECFA5hnrJPkJcZB0I59jp2QQJenegz9S8UP8nIumzXIQd1CB3a
eZgFgNfe6wWAMLYi5cJHISayXLASSyuKmdw68q80/QgX7HBE9rKL+2C50iseUb5A
/jzmiFa725tmqqijIfVw6gATyyO8Ieqlou2E5SSl27ufRAoFtTSc8XpJlPkey/OY
NLsE4wyA+uDvFjpwBsbQoAI5c5gENykGc711b2e0gQZ0SwuV6In9zeTpAH0u2kLI
PvwImMaF/4vKl48ASRX9IFBgktUSqLi0gIJPFGywAiEwnE8JJbAjP7MJG7+wNCjt
BjdsuBA4wtiweJ7IUhIFjfW1JRnP/0hXlgO/ho3RCDwpOCt799UUGbeq2U7kCh/4
gJDZNk539n5uA8swbOyzUy39DOewa59LpsgaFkUiptwZY0ew7K43iH3eK8Xy8hI8
n/sf3AqJxIUUzX1B6HuR/m1QiBdRTgkE9U1LbcTxpSaK3wZSRCUUsehX9eKWa7Ok
fX44+tMtT7puR3wZDz2xO+W4pCtYXSOc7Bl0C190aR7MsP7m8/Q4HFmQcajp00gU
mRHFGVQgATaJZyhZSP2WoTVkXvHb+SnS507fgjPyC0u7hOsP+5pmVkdJBpXg2mD7
wAMLZrWQp+rc2QkjHhHbeSWMsUyITrGHLizT/RKREgND0r5B7H0SnQcrV7wCuWj+
LVXiVT/HNw3TStVNrTPzEw3WSRgaa/Etzv2UsgppCDi8sIgXOCDDmawOjt/Ah5HG
ZkrTqmvQgPQJdF9/xRfXMwdIvYHgsDfMW3lFMQg+3DpJ4NmPYrToy6vxhRY7CaPy
4ZC+eP/z5ePzq4VAYxBi1hdKlqx7yE27uYIqs3sD2RvhC+nGYLMyTREtdfvdWATH
3tTURdw0iT/qiJzfXCuSZrOJrujjbuWFlqO+njwpaqmzMQtu5SarZTU48hQMsSJ4
OJdZc4Mmz6r+OLYM8+hcvr2ygeWVerkQcBDTKCefxwzNHNJyqxVL8h7Cy71q4R2q
Ja9Rs7SsYmYsBVjAUuIX05Kdqvu5EZZJLbTSXZAzkfQiIeEaMTt3dENoZ46Am6tb
LCJMlTB+PP83Yd/1MwYQMZbtWejL4EtTeDMDy5nKLhTsbc/zEkG16AZd2Wnn8ScB
TOfLd+1vWXBfGmIIMwu2EXg4oqWj8lxC/RgwOcXgUpaHr5U7MrDBrDAk93fR+Ue2
tD+L1cVwkMKEUQjFSGLD/kDwSzhdDa+eytRSTQQPYohNSbrEVukpipt8bX9wx8KB
/ptTPgWXlnaBplANd5U+mDhSLXgZkWMXO7T53Ui+MdSD8ZNxYNn9cGZ8LXStN2ll
t2VXMA5sMd22uPLZRdaDwEtavS9wKn3dYhzH+TmuxZR+kXhdkiqASUb6xHzUf11T
qQHXCkEezhiUqLUvXAr713l5Bh5EFPr7w1zbPSBHlFzSmgL3w1C/i8mGofnS1b8O
ExaJp7GQg7VYiBS39pWYxw4MegwfHdREGPW+8mtKy5Xyn++QMGBPOVkFH87RRoYW
dax/4anrxtWnR2lfPlKYOm7CCdHjo5FtPx0qJpf/vjLhauPHrqPD9QXNJ6E3njRu
+huTCFkSfYvA/txP3tQwv3do3kQw5HrK8F9g2/MQp0aw+XZMaTzBekNlgvA6q50o
1ubcfOQ9EuDK26qUgNDYFo5+I870zlalAUzLH4E4ncd90zqsqd8ONoCv7QoJNSW6
BvdTFEHURkcAEggitvVygwrjzRxZHllYybPleZTkt0XAlMoqJIU+wC4+x3qXj0b9
0NRt9e6uJrKqzYqx/NAYYG91OE0vp/+SvL7HnI//omRm26zNwYn0krxyxq5WLsX8
p0micPPRBTCJyHyuHm7DpffbwgAyaq78j55ZtTfHN11Nght56lETGKbX4Gj8uQ2e
rnVGhf6Ia8Zm/jvAH7Xg7Zmaqr9w5awGI3g7CKIz9vSP9mijFbXzk0YV7fG9iZgS
YDvX7gUD2gcAaRaRKfXv+/wqX/A/ZJij3VAvw2q8MATJpNg2XAHxMRsxmJZukOim
L5hZaC91ceX9vGgiD08VXsHvMRITcG+DXlw3DcOV0rh7I1uL+0RzYJ39YSuwsJoq
GJy+wPCzIgYezY9Po5W4+9y/pnlkuaBfMv+JiY2tsf3eM/zoKXlG0WrCdA+dF1bD
zGGd38GlwES3izC1ajp1vGAMqw0NJmEzAkugh8hUiFDZHPgch91SZzDyJg1sN8N+
j19ako4lYXYmACzb5ohOZAT02xC2UuRrBoe3pCZaeag77lihogI3l9xeFF09EvPy
yiYswkF3waff2NgcP0QJaSnMvqVa1lSsrL3rF/EoN+s/Nzn++0wTlH0uSSwBNCFt
Jt4/95iKdMRORcU7DAcMliRudfgo41vntX3C5P+9kWWLofrpwQoInHBT3LQG7I7G
1fNPRI+hSJ+JxifThisQrPOL3RJZWRwgWBcAxraT0C5I+uvInHyoKeE4Q1kzk18i
BdRvyGVIfZ0AEuPJTbx4czkZrLondbgVqSU1HtEYzRdx+gla5ZYGSaRuSQN8oc7C
IV9rmUsAGiee4s8XMGf8kBbdg4PZKxmV5LdDSlVoNQy2EBsn9zbK4AFpqO9b+xts
6XmcyxNEDcWZ6SoIz8tQxt3dpMaEYPyEzLyqfbaJBdFP8aHUL0DHPsinte43gCPE
N/ofYiJROFtPTdldJb1KIINZiwN6QmX83z9XK6Ljo0tuG95rhKRtshFNqTfnSGVj
q7PLQYl+Q6AhN+biUqeuCBwK3/f6Qeo3KT8hvmv2AGVIk+KAbBimOyb7mAlQFZvF
AsQXaWhEICZWBuSLosqX/Pzyqb5yo914Aya9PDQmp5HZKfUPml+dwAYXVi1PebGV
OqQNQxx07qRbSybrZCr5RIbPI1GJwTK/mbbWe6f5pFkzuVJ/J/LoWhjr6KqYXztY
ScRY+9Q7xWGHazJKeeePTiigAc1Lm7DDtCVYllGdsJPaDFlx6MUggA/Dzsfog0ct
DQJ+Qse6qYhOOt7yPNuK5ZGu3k+ZlFwBDMBfVqu6WdjbR6ZvTCqKhMKa+WY9dXbi
IN8G7LRe20N4AiynKO+JSsc2Q5wDojevFafmjKl+4Kwnkyz+72QR8ikMikUG0YWK
9+yxncz5IiJ1jlYlipTYzM3yAr9ocWcmgmLeKLfJ6vMxjx7Rub5Eo6ic64ZXdLAD
ZcN18+dp4x8DnmXxIniT/MS9BC3dBN/I6PggHXeTkTPCe4UNh6TvhIoYYBh4DhGU
nfok/596dUXITpfmfVPIuTwupcHzTRJBnUVUj6dZvLnvQDESCYdME6tl6+R0CN9h
sYKQUyYDpB9xeXmQDBSjndEgPWJdGFNWybWchMKNn9MHVWI+ZNxH/Yf3Ckf+QgS/
sdpJoBIj7dx9yQckRXJ0mnQVDOGcPJVBVM5q54ouzlMuHx8vTFaY7irgA/qGVOak
qq8N12XKwyc3v8PwjE/XlOeCyAfRuVRhz2mQmNIcseSeIvyNb8EVMLrVQ/6zzL+6
ddngE3kiclvMFmEpoBmh9Htc4y75VuYhl1vsb3mJ4sZY0TXCKHmdtdib7EnhtT9a
H6JRGpUMbDds9pF2Sqv1E/pzN5tHA+ojVW/XMqhiehb/PspQlFs6OUcl2kHlBfVA
cqykwMBlBDkNIJf0lm1anwhXafUFT5x4LCbFtGRjZNoXgA8TbxEPRV+mvPu5wSZJ
TLytl7Zc8E3//0NhhP5pJgm6CBpFWnpvtPpwbAWFAFTDRphrNdjZIZw/BjTCL093
yWLQCMOYIu5ZzQpBdeFd94KFR2zv2yg5HDoHp3udRvHlZMnO4xcwxqgdo1h2jheX
ODjUAm8O304WqpjOlQIg/oB7k5G4pQVklZnQZ0cybRrvNCjm4m0dPk0FR6qvk/2x
4dCY2tgpr6KiRGSGM/Id4jLUUj+Jbh0+wdAB96n5MXDgoP4jjG6Slc1jEuujKvkm
TmaypDw1w4DMvKJmCSlqBKZUulStyCNhGBkilTHcKXPwUcLXp2z+8cedL6U3nuLx
RgmE9fv4mTZG2P8OMscb6qnr6XLPqUJ8+I0jxcZLHHIGWFpXeT18cGfZnXL7rwdG
qnZ5vn8SpDn6tlRM2icy0Ea8M5TuWcnmKp5zQZ1t5yJVsGHYdyet+WxAd524KBjS
nZ0XO0jT0mNkkJta9zEfwMOVUlOJnrgVvo5KJAOrPbzn8+d3N9eb8JAlRv25Hq5A
5z2n/m+0zsq/8W1UbLUox6ZF6TPjDY5IcRkuNq6aV12pJ8oXqqsxEkrMOrEZ4rTI
tCxNbVq5o001G2apKXT7FHxR0y4IoGkIliHHdt881Vq55EhCbJOiOx+PDR2n6ZKH
j82ZSc0VEvuBWgwH7RLl4TdXdiYwQ/iqNA5L7Nx/m6zcDl4uzP0TcHfgxUR/brvz
dJO8xdiBMbUlOC5YsfUWGCtz8WnoQJXH2FCmc+qScg2DQPUgxNs+58GWubTGItYL
eGK/e7KFr8mswxot0Q7BYiEsrSKk8teIJBdSE03Ssush3xtKVTlFTxUC8heOT5Sf
Ng6yi0Fnppe4m2ZGb+2cUfH4acOcNu8GSeWULiachve4rt1nlaVPPMteO7N+5WGo
INZV4lQQr1djp68y5i8/vLhuxRNas6GCaaE6CW5F73QmtGSBpC22Pd6Fbtl+8N+c
gI3QToWWmN2FdQ8+jygLgCHbEAntK/8p7W1FBrX7WNDiMoSMfbWOXk/tjRcBX75s
hqbUyK+0XAmPWChWeLMxxws6wnCo4nijm0IBv26znAGzE1IsQXRjCVXV/o8UtnxW
8KojqWnAnxH+H4H4fmmvUUyJILoY39RWPmmiPiPaO+mnLb0VtqrZrQ/eE3jVkjOZ
71j/EXhDPT5Lk9dL72EC51rOe3HScv15WyTnIyhlJO6QN4+PJdXTX+zmzWjIit13
41ZEI/d+XqSZxyPOG9i4WP8WF/UQnc262uLE+CmJt5wFWGt48oJnpM9jjZi7fEJt
8ts758SW/ed0MyR34Gl5xoW8Q0+iaeZNkZ1Sqq1OvMgzQJs21r2eCemZFS/M+1QU
kI9XjFzoMrCzvQhQvzbYAVmxTnHZ3XJVZab6ngAkspQlcqlshJnPSl2FouOcBAn3
v8lhYaNi45WPzf4bb1Ll1jM5mUdFHZXgPdeLFKUXjdf86J6WBrm0yE5rtZg5HeL2
oT/M7V2KmluJ0q2VXf2Xjw8egqnFqQgCdwAdXFnazgXdmRTipFwNrLsM4//wIbyJ
lhb2AzgA6pBgPwtwBhn9mZ5TssBQN4ehLdgl/yKSnDgFFSVp1PsnSyiMXGmWbZm9
dc/dlwAya4P5yBmU7eHFmet46Al2xv4fyy9H+31vT7A0ZxMMsW8uEQ/N+CiIw29X
9U3MQD8wOx18qqTDYdhvPmaOAzlzfr6138RbiKYOAn1ryu8ONgck0xwdAM/lVbWZ
Il5xtmaFyJluQZZXvbkEXoojFMNEbWgGsfFkKEnkVvAnnCvGZ1BzTGf2e+MlhsXP
goIHGcFCafdCD7izJOgVDw/Nghh36y6hheYfVRtRRb6R3vnTxjFSodNsf7ccWs4W
kjiJWeY/Dt+P42YffXrnZJpozODymhrdAZvj3n22QzPF4ByqgWz8dRqT6XOf0K9B
JXDFv7yXfIUtEMfuvjlrbkASiiOTnN+KHMnp2LShCYPzgEtwcfX5Lv9p0khUwyi4
9CPaD3snlWfCkfUgTAIxpQo7eh4K1w8cbAHIbl4atCrBK3TK0MI+fdKG5lczn2R2
vYLGKcDElkXkrb6FmAgtv0YUEZ2+xVHlOiaTkhLpVLwU6kYfzdT7/LEMtUAiKe12
vwiJ2Ix3zEWUMjQJNEfqs9QxqouLyA15HpqLYBpX/8gwvxNNCbUzZui2Mcofvbl7
WJLxTY0stkqFrt9vBccluuUqGXeIo3kqSrSHA9XgZRDQa+Yzkh3XWH/cvbMf3Fyw
UWYhT5TTgN7eRqEAqe68uli70vn2XGSIvFTg2un5aeqrZ90WLQU0v/CuQi9o4cxc
j52zvUnWVz5c2MYLJOc4GlbLvk0f7cRXa08/7EZJs94zKIPl7rJbVmRt+GMMrrUk
Rg0/0GDo92DbAFvrOnTAe9zc2mzAC4CwewgKhQqH4pEUjYAPHguxPm8EfigYFM09
tge1k3BCU7dc9XX3Cf+zA1FK2BFgwBCRqN94ZxowZABmiS7iNlpF5/GuYVBP28fu
Q/7SHQF31IxjdpLiNRy8UNsIbuAscebED+wcMWbguYKqXjzm7n2wwzDdqWduri7K
8fcuORaOK9tHvROxch3/qN2HywVfw1lRncdbJezkhPBsDoVSWaCdycgnKVdjgxpW
ppFymFu++zUb3DPHhhbd3lVXY25LiJi6x0eU1aMuzW0HgTUSwbpD6bk1vd1UOrNo
oYezE98W9DHNCtmK00PdWQu3OA8CzbjVHMx5em68zBmIviuqQ2tXgahgXUKot5M/
lCz4mnPX6TQ3xiguszjXz+AIOw1BFTIEKrHs4OHTNJ3UKWlLg8uwCltTgAZbbj7G
8V06WBuXrwgbV0VLBiwuEJLj6W3Y38yjDmFdVY5r02KW/rUFu/wCGKsEqyb+JgMI
zUG392gNCnn4PtY5dVfzgDt3LG79KOFqiFlaUFaxa9batuHc9m/x18Rt/SM9vAsI
YP6yyhHztTiV6p/pvgyXf18LywdMDpTohG+peI2HS3K0qQX5Ml9YqZp/2akNieCA
6/eBGrSsbk+geovUO2PrWoRhvTVrEXpdwwumGvkBvfLFvepOxvF1m8k0d32wyKLl
Un/Oxt5EQnAnH6AKnUvI+2AGh8+RlFgc91TPQkCMCvGU20f37qrY/3JlFsmB89hD
STpB4kDo6b6fwA6WP4z/eUvxXy2I7AHXHX3jHZQ6AQLyebhPnXkdBHAlLkqG2/sB
F5fB8ajUmDIA5B2cNLw53fEkjKwMAtZaroZUxrr9Rk5+D0kQoE4bbqOClXpcNqkD
rqQW8fHGW0WbdM/gk1i4+w4ShMWhenKewZ9PVReI93w/wR8rLaU5vfsnAtl9zafX
N/2g6I+VXZS0L/7DD6zef5ytRreDQJ7JUZLAasKSKzbbmnPE2bjoZgQcetvT2fR0
zAPpTdIcVnRdA9pdBd3OzPsKdROOLL5ZC6DsgUpDmq8f0+GzXobgLbLEda66bAU+
Z4iLw9YsxKPTrRXCYHfgWn4TqHKEFRrfTbAVaz9sEFr5Oo/DOHvGVOXb9w6W+xKv
2YW1PZG6R66PWsa2P7my3it9KpUAeT0Xrd9gWp+9NUJCrsXFxz+VwFvfQuD3uDa5
DXg4HH8Kz2oxRNLX6V41emBuAy+GDdHFsAM8CXgcOQpvQSVSIBa+qcbookEeBy00
8mlnO2PcNsEHKE6RA26ewA6Fx0tQnryXOeaaZL7IyD+e7Uba+l38vHas8KyqWiY5
wbqTesVcouvif0Z9H0udxOATJs8D+tvSHRE+90geBewJ9dcyWh94TgAnFNCXDFi5
qp09e58DL6v5tCMFE7m//XpANjZiY9geGrHG6cKt74tCeMkdG31zot4QO7q5LEI3
B13U61PPSZdWg2Rho7OfkCZH5yErdvHFRNgvl/ADcsFhRFLB4k2eu2txHtm1a2Qh
7f4bCoRne9Othn2YHlNyXjG/VM49H2RUqNMzDNbdaQ7RJa16ttajC1da/HRPkH3z
A0nXXfsuVCUbiBrVAqjqL2ZnpRgIekMIOhxZGkivZwnCtSYHj22w6IopMDK71R7z
a7LtbNzdVDiByJFTapFPvCb4Qr15iVwIp63MNCVL+mECAjxKf3ec3IGc/ce3AEdJ
GZza2ui8zba3+BGriL93l68wa1rVS2DJop5Xrr7hoEnElZH5/cZRnU2yzao38ZDs
W2t8NbkXXP/7j7PO1Y1z57MQqIsuIHZ2MkLC0SZR1gYIoeYeYzRo5Qwo26DHBkzP
X80pIw39oZP9frypTmQ0jqVWxePvnACFXWYZvTq/RrXW2lLV0PyA86+afwt0Sldv
cpvEMPsal7UQmcWv2SY7zdiAsX3lQpP4d4pZBxR7aSScHBkNK5rEJuZA07PfOLyK
lBfx4i0d2d08eBpTDCkkr/+ItabB7OqjA7SHri5iovafO/5IelXIX9KCse9Zfjxv
2bh6lLWX8pkQDXcTrRVkHiPFgBH5Sa2AiFR5fzlnwhtzXy8tcdYNqCPsPOrXCYyd
J9asVLDKV3qCYOG5X9NShmt0rNfUCHJlEkM2ATzwP4kYpox4kgttyztU/1eZXq1E
JarMM6KG7KnO7/8RiiKsexbz4R431o6StZBB5p5fweH4L+41Yhc0AKY79e6+Tesc
BdRHTfNXVfVG6GLX1LT36LFiSTt3W7cp+D+lzqBQgg869a7lv8nJsW4OJqQgiK9N
TRXU1OzqztdwzZXJq2kHeo/ZP3QMVyOEd+CbhFtXZGdtrCGOy9fPct0J72Qk5VEM
Xacy2Z81UQqhB43vl6bPqG+M2KhSVKdejJC3LgmswepEv4MJEtAjGdQPdRNOdFxD
Bh+LjdSyCr6LA8oayg5tkadUBPYZosm//mgDtye5sFMvwrTfjFzPq3/EsAf6uNKZ
n7bcrIoL7IS+Q4aY+N3WL745/D24j+s3JUEhXTzh0ubvYLTKKzel63BWWdzqFu7i
AnUaQKx0OIehc8EDQsRjgAUCfXKaeyF+EN9taWG+hF3FfboVo/kO/HDC4th1szJD
bI0QnKbOcsaLmrZo/aaymcs9eBH2FbpGlPOnZUhH5+5/xSHgYzwFQH5E55/23E0Q
/7+dxmyCzNT9RvRFeTCL+j4KVkUr/N+zVAdMM4EqluoKR3/i6oa6gmBfNnwCOiqn
rKdmq8RLelzzuDV6T2YagBnYRk9hgvuUBC42PDtx/hrb3s41wD6+Jb9jCUEx+EDy
Qokvgi2P9R5hhJFrxYukmONtX/b91gl30QPQ6EOrcH10hcr8HjTwkXuac9u4Z3wX
nl/DiFI2UXz9tuPLyQU9J1ulXk3zwvX+MMTpEEQSjGUNYUsKUZxi7zPMzE+1nFtM
ROkCSeKaiTd7gVPB921/3itLIAjW5d2TJhr5kvcEdJmpIngp+hRLowik57VYlKaE
ahB6oXoKRt3vbCZe5KN5WE1kQymjZ3pfr+lIYsJye/4owPGV/xGTKw8ENGvSz4dt
CWmlqu33iWnyF+Q0sZjlrMhNjv0eRz2xtqvS9APUg58Bhf8DQ+m8ieVSrCudJPA3
+KyW8lgI/Waki7FTFfjhCuPPdMr5ztcvSegWTyyNXW7oUJkhlMdmdWfFVnHq/OyU
KXaG5EsSyRB2IHoD8sirL2ghXAz1oye7gXm/y5himVvXQaJSzVqblzrzCAOUbcag
kFQd0QhUyl8sf3m9DEqa/PfGDaDGgm7zCpAlTEbo00Ot++37L2nn1grAOb3DLc0d
kVfchwZ35gTdzBpqsPcmdymvH2rZUuvwepKmRiBiqghapP+CZRMfDTtmAJ2BgSl8
VvR/U16e4lifY9l2j7ebVduwdgu3nclyzo1k5uGHs9l87T7sHSxqE5uLKJBkKSlt
iU86jCE2MjhBRLKZT3Qb8LfQTj0WUCFL062p7iub4Kb+x0e6hdtqmIwwjVen2z67
95qidGT0oXqGoP/q9UfOWAEef8Lc6LNHgP/zS46rZd5kQb8+bsnuY4DiXtknR0Xf
s7VYu+KYjW2airjBZGuiBZfP9jdv5ujidKhl6eJx67EiU7frhSlUV8wxltufpqMO
AYppvBXs1RM+UqXBnvrk0gfTFGUlX8if5oeFMoRp98Ak/OVH6bTRBc6ej1SiB9OO
DtgzsxW3OZkU5dcU3tl07SPiAkjPUMK+sE1C8D+j9fk8CeZHPh6uWAxQp2X1jZuP
S1qbZXlbosAGcZjEw8DScfz6pGfFkUW+fG6Ckqm0YzJjhLLP+GVpS+Gbx1Fr2ocB
ECGAdU4sTQOJl9AzEVi/Atbj12NoKJagohAmOxo55Dk46WvvZtVBqL2wWoud1byT
1W8nwZE2jO83czCh02CcMuljh71qQAnqbDfcZ16MiyMzDtO2ssuLdAOkq5pBO9i6
el0JOGV56/zZ8quqUGdNxmWVfA3wD8gHJCuvpdWvkzPXqG5jhVlymg47WeH7fRrc
EhE0Rp6GP4uaEYLLQG36mEat6Du6MhwjayjdOjFwNNyBF3NZO6qM2qJw+MAbT0/g
JWJjp5dI1oBskYjEtP5xywW/nU7/kp/nWYQM1yhnWVh9KlQ2ysqu/kfrxxhtZylb
pstDBH9dIw56oG6X+q3Hb++zhJbMAo/Nc2Ihnf046kAQ3sXohiYTUYVeTorQyo52
14lsTFUOx4WThAGa5Bk9wpB2YnBnW1BIfRt0gGhWm8/6Cs1sJE/ZhoyOvhYxYacl
4ZDlN8lEQzM55BOwSVRb2Cp0dEynLlI7toNshsuq2w31VD3m7HamNKnCmWNQ0G29
FvOJOGUVHeDqihekxtfSL2YakcqVZJb1kvjQLxbfJLyYwcXQgs10/pb5q+cO2MFu
xb4xLczfqqJJM1wOmqavM4oHNTSDRQmGVFhZoeDpR06zw85FQgIvDjnLsY2XhvHR
rFuVe9jhtrOO7eiBSZ8nE2OYyBdoycl3fWyDEhiF16dj2XywD9Oh03ay3tRXRVuH
EB6EThGY+HMaBoFAYwIBmBzqYrtiY+1MrhAJcwHHb8pixF/UqH36I2KvXBEIt27o
ewasuCveptsmBEJNT4n8iatULDZQnUQWmwbohZpC4G4JwGgnQDhfJW1jOyrTxaN+
pdy8ERwkl+K16ERqC909kVUO9XInVAWz30UBlUq6YM5ed4nyeWhZTeFBMMS37Eo5
FkRRX5ho/gDsI+BdXN2ozuqaRB2j1zzpDH3w7BQeOfKx/uxb33mv7bsa19g8c1OR
Fiht2CQTBcbLXHYW/EQhkvydR0wP1WeS01tMAmMgphj1MoWCoj5ZAZhwchXFU0Vh
BLzHsVAjfNRnqQH3qvisLn5RTHafUYfNGnrpQ8FuJiEl7OUIygoNSdWRVN8r/Ne9
x9ppbmcxJqG1CZ3+J/JgfZJv88NL9+a4a5kS5ajegXyJo6yfYkrTtkI3q4HcS3Jh
z35Qhud9CeYzg6blM80UVWmY9624Lv0Z1HvpCJRZpv3Ea/dM0pShNRiwQjZLWgCq
yulZf1Eq5W8E8nfbbUUNLVip6rVLC8xDQhgr0iPNXJ0kQw/jkMY5yBMAK51bIpqT
fmHQuWJ4i8+914clygwecZT7XOfhQoslv03+nhn2Q4DVqaqhNyPgpWnv3OGs8UJf
zt2HqQVzWCzPPJpBKJJclv6Lhy6vr7csr8D2zrNS2bbTu8cDc+c2/FMzqkr5pc2o
Ju0ab2rMege1oxcibogV3OhWDD6zH2uQYzlLQA0c4+d4xpmqEYP99jTzIymecWbL
alKk1qvWYyn92v2YUaUtSUlVEbR4YzuICM0s0IHj/wRXORMQGJsaP3oY21HpeRF3
P+qRz3mGI3MwrsZZUshnmRKnUd0MpDL1F6+315jupiSlaeuGBpXaCSPGAPV9/zTP
144HRnUZwzNLnzw2LX3Q/vXtdfUVxEcP/Jpk+WIfUwbxZk21ziPNwH9iiiZiFP3m
XJbxFbaiuU1hy+T6Mcs0AknPOr3EqeRzH8dny43/zNbHjTu+hLLEQi954qCtuOsv
rrC/gbf07R6JU4QW4OJCzcRex3hddWvvNg1QxEh/3FIGWBGigU9DdgCdGyJlvddd
fQuJL/3xVIrbAluyHhKWe0ebQYBLByZepcn19//+UlaNdzxzvVn1wjazJQugPGTA
ola1a3AQELKDZGYXvSjNnP5qTCLFP7sRVTTEPkOI7lazMSNS5B4snY9ydohjoFmw
gSwXNlmKGdJQ0DF7gu7yRCR2zVSTkM1N3+y/SYvhbNNATSl41VdjJiBvT6v637tb
P5FMlcH45Th5IkMd9/XQdNJoWD1qrwZrw7m5kGdoeGF8GYRS85Li2j0b9lC05Iar
m3j/MdPuq6i/fkZgdcxoERV01TDQgqsz2EJlrCDFgRjqP754Uzsz+ASPvV35tZhZ
RNIJFRD09M24xYEAfwIGNnQVnTUHIDq7C3q1vyoQExqD5KEIuCiIiuIppCGn1AS1
zBP5sUi9Uj7gYpLdO3hHRWPBGMbn4aDPgI6G1sUS6bH3J7dmnwwmDmrK6pQuNJAC
WTPwcoDw86Empaax9OTd4grIYaTopTiwMHLVQXVlru0kuiacpaIPJvaKU4t0nCuC
AS/WWU/0Tqu5fv5iHsOhhRJpY4UOIaAkPBfMdOZyJItYLkzbLeRrvQqiG6xcBST2
PFDWgWAifkXmqDg2Qw1vM+z427OdZUXYAKa3VB5lYT32IKBbeboV/wghbgcVK4Kh
eRhz9Yd4ZK5z0/aY99Djg+eoIrf5+VcnxSpJv4x8FDW6sM1ISDL5QTbmIw+Fg9bv
uP+EKC1DommvAJO3RXDfsJVhQGiR9tRKQ7vR8vIVyrmR8kvLuMO4gCn9RhYQxcA8
DgpI3plGBMJtJCxYX/ZT2jJEMSN4f+ow59+be44ZjwQ8jx72AHB7cmFOD2KykQN/
PZGuc/b5DDO+LyZ2r1KWLM2CcbUeO/RDgu0bjW8ZlVYY1mgxW0bFzE9OacyEyK9w
Ez6GQRl11NL8YaDlCw5lwty1MG8zba6Y5ga61Jv3QkXxr9MoDETSmeP/hRMjgm/9
SjgrGptppgtofmFZjJow9CRYr9u+g+cWRMGw6jypn+Uf7AxEGCUQVU7s4ow/3kAi
ybElwjp3Fx8nC4G8FpdIhT2IicZV0pGC4EK1AuRj1D00xWUaN2m4orJtCBa5o2km
gUnZ8Rm0/GDNtPLKP8m+NUdOGhPDWnaC2LXHRdsH9Sj3zGh+jxnZPLNcFNLQosfy
pPAbKdKoddJrZneUZMhI9Vpr709aAZNuACOGfM6RrL7SIe7W/KvkAbAytqmwnSg+
iwyeJM+vwyAUpxWFX3YMYqSha8to9zAlCINdOTop9Y5Hp855ZZ++cUBH15KtLne7
Q109NiHcEbTjn2lJFm72WVlrhnQ5la1muc8MyyuDJcIBqyB71Jo6gTt/DFUkLjjE
cTnGt4gGxGARBEfvATsh1k2LiCBm0ewjATZj7A12rVxzd0YrPikvkYrTGiujO/wP
e8JR0ffMld/G5ECAHNO09LhlCzTV3TRjHrh0NJzKwnzv0EOwNUE6M2wV1u6/nDq5
OcoRxin2slEizlORbbzxLqzoHXsLA/l7AmiTlJePZ5XHrch78lzdtWT6oQdGVy2W
7Xxqlkdtd4Y3SJX+VD7PNJfYDtFAYZDPq5WCJf7Qgat2wfzM69ZTpHRmR6FbJ26b
Xs/PBX5SDqTSyDV+OLX58WB66Vk5N1j+R3zpNTSztulTNb1VsK7O+vZpulo9kOJa
vS/34sur8O3w9pP2X5SIGOwRg5x0MGo1rBQOjteW83eDxKgSFsKdtRU44i990WbA
mcnCvj0bb0nGzRVLd0dQe7Fs3nXJndNYSOHlHSOxOCN5PBmbAWMAXtkW8flGh8EK
EESja9UUhWm9Q6nNbRiTdY8KbgtRPZZPBTn+fEQ903fkgpcn+LjdeV+eO+PCYAcJ
cN09+UIDbuKKpR9lU/FzTA1akfBkKcrCD+20VpN+1LHLxPo/VHJTw0c9Fw1RXvxF
7FFzD5T4xQlNRevt4bHtk2YcFiMkA00Dxhe62hZnHgmRp8ftszzrbiayobTs34Ms
pfYnswnwRjKYF2ePKj7r1mEP8GVAo03FylZODF4j55z03OsP6Df7vRo7CQqeeMeb
0u+C/AzHtNmgCmay4+iJVdNUEvIJAl3NEg7AuJJPfIUwR22fdumyIiJYPKfPUHjS
Y4Rmj6t0p4G+kqy7yO04NQmO6dXxldzKOtd9dwu4DaENY0qMVu4csnSXajIrfb8H
2OnopcDwI+0XxYql3I4MyxKFd/kZpDS7Vb/OsOwOcppGBlx5ieK1u/hIjE/Mf1L+
QQvLHl6wbaIdKumx+6lvegb7VX9AClU6wbS/ObmtEG78/ZKfCBGXdLnG4OJ6ZcPk
R4OrnPT0pDsz571kA/xYyYl+yESEhMJTTXnjyrClYeCVelfnd6tugpeq1uup7Oub
vhTB7DBuEpLN6g2HZLZpi+xA6TlAEzCG5ewx2gPOB5OpnSsptR6hNlFoyVf43JXd
YHsFlJ7LGmKrOeK0zYVOtU800qDqgWsJ6Q8W3ebhdPwzVAuoCkFR8ziq7xBLfs90
f0tVjMcVoWdxvOCxOvlPlLYeO5+kTDGNlpD6sDgA8mV4wHp8JOLYIpmZIZVonXHs
l72QQBf2RC4kEo8566Y9CoyDDRBH/w40BCkTQLT3+3TCKtA2kAcVDc8scSnBJW5y
DbL8jhfoPMjTffMi5ouUlltOkm5nYIPQkzYCrFjhSje+rXiAJ46iW/ck9Q4BkrXk
dXF5FzbpVA+WGRf2CHxYvwjJWKBaBMESLplVW/R3UTV6QLk6LKX0SsZVf12elK4t
dicVLEsbpgC9VtM+mIQe5umOdRaFmOlE2H8AhHTYQJQokJNbsFwq+KqeUGBJI8FU
H/Rw4nlLmsQswt1y5kVT8JFcHXsinV7WNTdAddrmBxKlgm09Ecx5dQmnBFEpWpwu
EXKpe3p9+IktmJUZAt/n5YEOeUPusoanGdRt9dKcGwCgKQ0T5nI1Am0fGB2/wdUt
QaV9/HS/iTXEt7COGG2wHyrz0Q4r7DTUoxiSiyCYSnP21IpmUmHKwkzq4N3VN93A
/U07ATdHKWQpGvclabWKtmWOyNFuUZxRR8p6xd0bwPWYawqjuKIYcnSSzes4Y0GH
tot6QkQdK/3vqIRBvBkPVUTNc+TJXHryHVhvwZrZBaKY5AQv6APuu1IqjowOW9rj
V1Y/m5XoYPRADiOUK6VaU3J73+bCFbA6CK247GKhrUMadVqxtFWp/ALY5C9XNVHi
ewiwmeZZHw1x95IKRD4EDpL+Xxj6k9vO1KMZ9sy8b3386mSlmM66X3hhOGzoP3Ig
gluNgvta27tYj/i5Zf0HmKohY0RIIjk9RZlGTkDHFzgQUWisPI9185hJ91OEqbKZ
iBfD14koiUjd1vDbpwya5U/UazSPcPey+wqn9t+jyHLTUfY8LmRDN6k9i7X+upUw
4K+Zi6IOrz8IUwKYknwClCDDxXD1t0QsMzhUubIb3WLInQMq+LwZXiPpt9HOAbNC
IDrnqIS1pJkbI874edknlOXNC9qATFkISgWyGCr1aCjCGYvhtW94gPRz43zR96ZD
C0fyP6cm+l5pJdfudvbaUVyMF7R1o76cUOIuAHR/V+jUZOsqEIx3SEEEucyjRJoF
LLRPiko59D9uUfbiZYKXZc2PjCeILGjgcCFx1Vl6RrDO4cCTZ3X/DB1HQ14ToUb+
fMvyBdoOb8DYCbz1e0NfBIonZqbo/z0Rjx1wGhR7A/+iImJWQ3zCCIi6jv6TqLbr
fBig0TIqzzT4+ghwsDGLUYa5nTfIN4qvD6Po/WH5j2Zs5kVVb0CXUM1wCDMvLcMQ
xnd87IAQbiVSvexD56JsmX5DM8aY4ERhbtFNA+Pa4SbOFCHo5ODhL2gDAEiY5gLS
9jIgaPGWmNAl6SfcO8X8VWKe3GCMSKEmzTKvSMYEp/3kDMNpekZVDpPO6mw7XHFj
kX2J2LgykSUwFCW/Qjh2gqczqlKfdSwEa2wPKzG8YQ/AwIRfVDqnM7oKKAmJL4Bx
QHM5Qf186tJOrVdKgwD6LLNO1UFsWNTTpMH7pjFs542zV7w7LAgU2B+OLOaUdhy7
L4vxrqLDrZjLnd8q1FwN9SWwMDEdI4WlzXhU6isNfLRTxI3Y85+6FRe5EcwuQ2g+
FuUtCr+JLdfFR/T3bwGR7JzHmCyLuJQ4KcnEwZcWxla54dHGAFDi9UjVq65Oh4F0
0LlBdWZ//0rWAS6niHbGop67HoUCJT+G3fYiZD1ATlZIlt5tA+qtBB6E+M7AXAE0
znLCQpesdqqtrrnOPdGKsbYFpVrU2ca4r5adKz+MK3GiAID8/u2FSCDCo6nvZQ1d
Y9tyFWIdUoiLt3E40ZvVlWqVvFzwfa84j4U/KeB0RQ8PsJCk/QPHDmgjxP9PHJ2+
GUoiZ+PejDqgbfldZbSE2xE8zqr4l8cRdtDKUsoFolHB665iB1rET6pwa1Nof+QH
cYDlOUZbfvmiWE1mhXFH8DaChrG3TByWAGjqU2acpGg6RFjjqQOIm3CzyEXttKP8
bO5uAlXu9fabKdS8NRXbJH38+TQ73b6vXQgKOUXZSEOnT8emINLaWqsorRkjy4Ko
vPe8NdKdKP4VYBjw3bg1Rff3gjQuBa0bGQXdVIEZE6c4Wb1DXmA4RcDd6wxqnpci
z8eyUGxKd72CqvTV4IRn33cyi7+CDdHrvqQadNJCModl7OA6ay+y+ZuKK7XLnfzM
IsQw8Z8SrVmnu854XhwPvkVLXPLvhnFDu40rcYsVw5gVqY0oZ1R+WQTiGriDjDEt
6xKj76sAIhTz96wZyzD4TQrnRX9UrVJZ/s32TzQiEBll5hsalVyckTeDChAYJPS/
nake1Yq+ctACSI1Yl1ecbcTxMopTsG8vHwqG9waNrOi6pauME/arDaeZxkpg7iyB
W5Y04BJVcFz2rp9sEQNmYmbJq1SuohtSbUDWKbD3NuuoBtqrBWB9J4u8UfdeQ7WZ
X/t8xaGie6DgB4hkpSyMj2lhUX5bUad/baY2ZN++I9gyT/awT8aILUfxDrHiuXH7
k2lt5X5s3LW9/ZSzdfqGrN3q3xO3cI0RATMGkZZtI40J0SQYR0HfO6EpNDIQFnuT
7eisFv9T8wcqnh05sjwGI1pYzYPFsCHPkpdtlQLt5mjNfa5LcUubUdkTxCS+qnJ5
tQ+YZQK0hZuzfSDCLE3mY5oU8mekuKZ6vBb08WN57UDmXcgJYNSv0elmj3sEYxkS
lvN0tTE6sLUdo2tkLGMGDG8xgn0MsJlJSj6Qf8eWey0Thz5SCVgKi53f34oWnGMI
qFUJhEuBNDXJeoRXK3aZdhfr22+cJHN/KjSOPxntX2+5Db9Zh2Jik6OwalKC3kbv
7Ulon2Pc4of3CQ14hszaPbRwodb5n0BQ3R76NPzSnJ58I5g933rVIMKNRyZkdT1T
MOSiVEnxaL2KitOYqLJH4fzkIuQw9RXo6GErp+tO2WSmUHKWMLIP5WzyIKdldQ3c
Ze9ho9i2B4fsiIJqhtCLc/WK8+6KWW3CQ/5xn3Xn3bViJUfVeBxXyaiNxR+SCB+a
xkWK3IiN3chfUILAJgOBpMP5VjJX65eC21kadjZiMiuROcyBS2Qg4uApausOyJrj
ayffJzu40CGm1GRrheLyUoZhbGgJxBTeO6Ry/Iuf6TecewbBXLE7JVw6J0TnRaSd
oAozKkpIVVXo8Gw4D2XIdgXAyd49CL15vRjTgFadoMAeDkFcQYBKBiKIk+X10Vvd
rcY798ICmRZdJRxYQrYFixi7P/V1u4Wx5e+v4UlTaNwrmxqEOqCT5sWcamHE71Eg
t/8F/rYpNZK+ZERhUjKnjUvNSZLa3UNwmlJKATLzIXyY3D3hTf3yqV2Fem3C+Wkn
CAbHjWG/Pi37B2dJjvi2mmSflirNodqTHDIeQmZKvpPy9+UFUxSIPr3WqMwGKoy2
NBiBp0nkJIw393pICqntHeh0YDZSfoT/aH9nm16AG1GGApIKCjeozSww/tlSMh7d
6EEF0tBEXgVHkYbYdFFo+afvBV1UBeOnIpGTLemZ7K3oca7pvcuM2x0DqhliC45x
CA+x9/YZ7emXHFDov6LLbx1IhvolY7SJkXotbWeq+eW8s0gUcSv17AUX8qXbN9Mm
ynQHoxjrrNh0Um3S/Ig2Jc40E6CD27X/QOwfci3Pl6SOsIOO9I4e//Mahva5n4EO
CF4RQCqBL5As7VOym1Chlfa4IEMmLv6aD0TRLvnPmbxPTF7jIbUnoc+whhjKghtp
FcT7FY/Ck68yTZW6c0x8MD3B/Zv1i5w+tf4IUSg9Ex6GpeZQ/XFrF6k9JbGWzWFL
Ns0h95sgjKc+b5fsqwsQ1y+ga3P6ZBtAkrkjtwRsYSYqh3VKbHZpqfhQQ4QH7hkP
OQkikIWja6oBDJM7hwyfJjsWNWJc79WU3iCDEZN6wDss/UKdQr44aCSRUDJ1dC+x
ILOcR1dmSwrPUevIHdACOHXIYq57qce7kL/zEPPZH7cvndARQu6Gy4ROCksK0wbf
LNcOc+f2zwMGgZYO7nGMgzX+m/sErrat46UwNZ0qNcPRnKdu/m+V2H5jzWKxsseA
EkEZWUk70cEhzwf2z7t+0ZhCZIxz65WeBjlMsw4vHAQuiLALRPXOkUsB/hgGRm68
nlNsWj5w0tPP5nCcI+PO7FR4ZnDeVREo3qMD7vuemH+0Do3TpYLFwdFF7cWtmGaC
kKg60mUYu/NsPr9hNTmpNUGvTrC5i/1v+Y7ij7nHC+yI0F4QdOoXRgFAwkS5rjiL
gc9o719Sb9siSSBDan46uILNULivK08SyTHDEsNYFzdIw5Cax1dpZ+wikdI9X0Z0
LmJqRDqLRYgohaUuMBfPhU5MKhjzG/n47BpiVTol1wHqjjswPL1DGVmkBBgqNwRo
qoVfIug58qCYxz4z+T5twLwkG2WUodvlrjBBmrRcnIMIpNWoz+hUw2gMSeQVzlKA
/7TKniGZJTPjDOCLz3ki8lL40RQsSNNk3nJc8sHqHMhl9H7G/1uLi2XBFCzzjKhl
CBUFPq0fgO+qTrtSAAEt8hLHpeAcfVajHFp9vQsWbKGGujR9tWquqO9Sd+hqG5Ae
XjWFSmHFF5UIpk6i8cG+ZXMawktePIu6Htjb3QQuzCbTBlaxOzKZztNODIuOBNqA
4PW1oDCfpoXbKEx6ZkLWTB5sIiWOkgeIHL63rhnwSmKy8F6qoAB8Vy+LD4C7Cpvu
ng0X7GvL9c02jAJGa4sdQ72ZMQT9Jk5+FMyZxxraYxZEpC28I+HRuObk9yppCZBv
tYdtVgrT1OXBhKW9J3mkVEetyBnEexlxVWPoiS9GeL8vRg6IqZr6ZOwQ2JyEG1P8
KB5lMobBprXlgTnZsXzKoXIrFBBosrIozyKLG5Z6vKZmsR5usOuO8hMb8r5iuF9u
R7Z4KxusmaicfBWDJnN5xGBiUNyt5N3Tsuh/0VP6WnM4HczouE4HNlR/ZoarKpH8
8Fxo+WvP1O1wq7rnY0Op8PI5OYPEPhyZo1dVaFVKg8fdRuoWMWdY4sU22wNfXBb8
zBDJ6C1oSFFrRn68YNgbLNb4M82Waj2eFJYFQfYbnNaVsSa54qC9RtsbDONZdSzO
/zyiP+kdS1IR4Ce1b2wfnxB00Lp+zWVpmYPpsfFkQ/iiWW6HWEWNFTI/wE5VbF7H
OTsIqF0JJhh+/8S9bODdwczxHMNojfpRs6l7v5rpIWbrvbtX5QVIFsUN88VmN1JC
UM5ApdGStw9aB9FViaH73/Hdc9U/KZ1eUd1gbRDyOtiSHK28k4LmUop1PBtTACi1
4MNZVai8BllZT1w3e1evnGdrVbGXcWf4rzw4b9Q/rv85kjr5dUQO6ZARe3fWdG/D
XMHqweYwkSmar9i+p3cUgMvRVThN65ZshRlM38D0cSNKQmEejMT8KzK34mhvWrCQ
+nQCW1ORX0aZPuUJyUNQRWVNJykR78n/hah0NvTbDhlK7ohXipk7AiU5JsEPXQvn
mvSW7p3Bx9gKrJQIWEIXXba/hLwl6gmvFdr22drGr6N3r9hxWV0R7lriu6X1Y87m
MD7Q0v9+5fTrCB350FbhomQibDYyAj6esCbQ8Dh3CpIs65OKUn6wlZEeZYUC8ZJO
79O8OwhCY+nm7bZSR45u5nlPMOIw3uxMoTr3C42GcG4bWK39ZR1Ba308XRiN3WxD
VikuJRpbRzsUZKzgD+3jFR2ZVGuF4G3DDrKTNTIHbsORmfzAlq51VK2V3LxoDdW+
5RsGA/PBAQ21XLwjN8n0xVXxwPQFCDltm58+DlVuwYfdeIhIsZ1l4UWEmFmAzUu0
ZoeWzyVh6a5LbO3znIWCBN1MYpQ01pS/kVzEuWLuhi64x8cUnBMliyDuovoc8D8G
SMeQI/psz6zBgb8cNvzR2+iLV38kCX5VXfSStmeuRAo0S+Ob8biS6xbZ4HBw/01w
sWL+qCHWjlMNowEbJY/wS0GoMIB0iaAY5sLD3IXd5QD7tA6daH5TjPbLkHm0qSZZ
nrDGwYj8KOHk7qN/YtN7+hhiBXAn6RkYxDeRbvdpmJeKchiREBZt5N/sT3/1sVBk
nsrf70hvvhPkad3qDujiGGi1jSmUlN0Xetc822LdrmMOIscPZwgB4OxfKM8IdO1S
yH8vFGx5vw7LasEy8/5EM+N14fs3r3AqQgOc8pyeN6jo7ClqU1eRHhzbJK7HLMIt
j89/Rood355GHvUWQ5XD4zOUcszwn0XdqkQ9v7Lqoi7BpUjaw2qOhvbnyy1Fegii
vaVHorTBM+tNiY87hCT46rxfx+uq8dF6LqO+PpMdbuxoQLw1c2ZW3Svdx+1DlPDI
qBZWiB3t5F/lZHNjS9kiVV8vwG4+YX6uhIIPFKBgcyeweySLt27LZrfAykljF9sU
3U79Dl2M34Xq8tI8uc49ZvO7l9jD01IObqQp3WLGnpOiSbIwKoV+K/sPxPZRe2WA
wq8e3ABnpLqYsM6HYv/nnbK9FkvR8I2NLR5mlWCJ9y1yEllFfsrVHqdwrlQZfkJw
ZM2JvBzKSCFu+U2+/Z/eRQRmcMRuvEk5pPMXWNexPxEpemq8TAnOGqdgceknvyyY
fsbuV2ogZpsrJAEua+dhdCfqvd1Q7zhuIAm0P4xBhQuPPoaeB2owqcwbOjI3pFpE
neKS8bnTpAuEtGgQaF7W20kzThQ82tK2dk8iTsz0SOF1o5Ya2I36t1QF70b6OdU0
1p+Y2rhh/b7j+eCLz43Z8A+zj7L4ywgztPFimyhGGJaCoHTawNm83CtHGmGd7xst
QQ8vtgh8l6SGsz5eVD0ZZmEzgQaPK92f8nGh65zxZUpn+sMiBuMKapj+m8EnEvn+
/T3O7iNQtDuIl2TlfJv9bL5286845aOa8jx2TJlx0u8gMa2E6MXMnX9/x/rGLiCd
kCBqOgpYVF4mBdsfeOWAnn9Ma4/2THVHXayLnW/7ajtIyLZege1aPLzZjbRG8aIa
R49z1VLsEAwrYUzqSlBqkwpPYLZwXL8hJDrggXOL5xjNuhf0vQf6RaIBm71AuyzE
KdWG0jHPOBXyPCwg+50mhJU4nr7ARNJ+/3lmmi8eiJ60n/4UJehvDdXVeeTK77+t
zWRE1sAQsOWjlimHNcKKzdaB4Cc7390RroUc00EeQQd93TTwaSYiVsaxDOOo5Wck
+jivSqt9nQxU0SVQSApY6N1y6cj4fxt5yjuwmErcJqGp/blr8nqFZ8aPoLd/Otec
4et0fb5ChdPlzLlq4aKJktahur2aPb20mtKGnMtz0vLrKyNZkDuelObTiqcMOkgQ
BDCNY2JuKjiBFD4m7BlfWpySu88kn/OVL0H5WWYJnMht72zhefQNgLRhrz+C59/F
S5FMcH52epnAcr/vZIq/6P5W50X1PJsGawzwDC81Z8DGxc3PXczEZvkV6i4LNB6m
4hBUlVTtEsUQmUl2PiCEumypooS8h/COo22esKFU9Wlmr8hdYg/bgyBnt1VXYO9j
BO6xYUEH8ts8FbLFtBx0/djImAIVFPOpAsOM1zxozS0B06OPxBnMIZqdBZb5VfKC
Eyk3qfcgRermDl50/OdFBftIkgtgyxJPMdqTFBzxTP9kuREI6MTixzweb2yNmUcX
Ss77jAa2QicIqyPtd4HTde5f7hvrsGN8u97jdvrHkJeAuUjxfc8B3sYwHdTpP6f6
yVlMxqcZ1cqynC+qzDJrEHE5r7eThnlNFJ9LsCG3xwqgmDoy2/m0/MB8cScDbSAx
6COjy6tE1VJJO/dU4etCft0Sy2ZZBU3VwChP5plZgSdrO1o7OINbMTU157vxwH94
85PWXKUgJtAsWrdntF7/asbm6SIlQ4bHuwRhZYW+5ECvojmD2DAwwMgVUriuZFza
r0ZemznAHJJCfidqMw5TMG7M4gSyVRKXs3KK3DowLxFeQDGt883CW6XkSmY8DkPr
UX/sKO9CfQyjiFrO6fKIvVKTmvdzoJ45cu2y0NgqnhiOM0SqQ+Vsp6/Q4YMIMtVa
RbMEwmC+Q4324rPXDlfJTtqseUeB431GEA2Mz42rGFenX18jDDH3gJRormRmL87Z
d7bmvAWF5afEbcyKxLWXxw2L5nplHKU8fJuJEGlQaE1hjUDRqQE8DyEG4T/VhMp3
/pSCvWmeUr5iP0tgSZC/k+MybEJGdvI4hIdWr8k4b9WRclIqr/hbOf5tSGplgu0h
Ta6r+l0O7EXQLxoO7n59loIxu8SEiyuHjajdBs3AGBD3RqmlSnanrF+XFrfca7mC
jMA7eiScqod2SlD0tGHFoKwNVmfsXomtO6cisFEFe4MiqtjsXlqRE2RpPuK6BIEC
8RdWr6Cw2rPHQgV4jAE4+8iyVzYXKYabrPu53knTyZwFCKJooGZCeKHyDCFHlT4v
MYakpclZvjy9vivIueSn4vYF09kfET4dLfwVLuOrK5+awzSywxQcRCiykffe9UCF
ogffOR2ijgr9NYhr7fxpB7rY0id0xNepcYSoCq+0hVhbNUYgLDxYq5ownTR7ucPQ
dqhaTgcScezuINy5onjdrPrYO1fmpTIvniVhTFpFmBCBE8zzX+VksiM+fafeEVhM
VzpP3fYonRcQvnRArwqAo0XEahPJi4cJoH2HTvqL6H2ms9jK0Nrvd3MlbwAR8Nim
PpfzEzFWxWmeECYvwhwCZyd0IV0hOQzzmQzOYYfmKHMDEpTWyGRtqVHsbrKhGh6b
BfW6aBREvAU9UgSFnN6k//g4wqyTZGICwMydj87wCERjijEQoYasFX0pjbt5YqJE
GuoE73WjNNlg9Y4cUI9aWSd47b/kEsgn1VTcataNTZ2ZOzAzELRRIKJTww/eRtKZ
r0clLvjfvXhopWF9NnHhKgg1QhNwIQTG1ljpx7BMq8tBkeLVe1quUFMdiDALYDb/
gyD2qEX6BONkg42VA+ct2d7w7zOuCWGkIAHb5iRobbYmHiAFb8hhvMXnLjeMlE7r
LiIPAO33O8zsoWRyMO9Dto8Ic/Jb5vLIVc/nM6tyXmboRvveMBBE+0tuaXsb9R99
6B6mqRqfzuz6IiM1vsGkHQgLaq1qD2uxwxju2aNFiH63SKAxH541WILuZOLZgJSu
Sk+Plt7CInXJ1U3Co9MbzmeKB6/Y2TZVpmV9MzHNGdAGZsUiSVwmhUN9J6lGVIpw
5FZaQfWXThie6p2Kt5KW21Pb7anIxsFZTELgenYft7aeC4pwTe0vqEbTIPpRnTmL
/JkaSSSm1wsu7ZgyQho8mqxn8GY20IGqL1KdmLrpqxt1o7B3x7cMyn6SMCQOPzPB
uTHITRFhD9uJn3voywju2I1gheaBDS4J5+c04yMYkFrLppIRkyf0T5PmelOpgDDT
nPe+t9sS5Fp2CNIWdJy3devzA5WMYbx0NMM/VepLMH1EJLasdfUHzT+3QCIJDm08
M4WM0bSo4pfv+FPbpe8naSk2IH9oqTnqSjbNiCPI9kvJVoq/O+rfZ6SlNv2f5nSM
qkvXmhOUlNIyoyn/CSp5GzP+Ve90CxrFIOFm9QbWsm1j/80aSgOe44VcJDtRfuW5
vZOtewBCGe5iS0oCag1/7e5CeAOEEymXglNbIv/D5dimvbLtuEtFwkNWBTYJuPRd
UW9YYopz3F+bzXTw8kPWFlv8qKGvfBBJpqFz9MgmojeS9iEFJL+Dh7b3HtocTM2V
R2jFm5iA+krMSKO3XSHqiKzHK8DM3kHmadW2m4YDlJG2rd++DCvbuGHvV6R6M3zr
4n3yn+oyTC2ZKtMgGHrZvTnSQBQST8+5Omwd2aOfDTUsgcexxQp6zKQdmAxVSLro
m4zYuUnXM1zQXmfxUvkmgC3xRaS0ISOJbrsbs6JHPh7toRemy1/jGYN8BKagWXHb
P/hj3A3hY/LS5oMddGl59pMpfVEk9U4LfYX2HIZ576FhrEKVqJsA869jM3G9Vb1y
odpdA90+uLHkXHnpoRzoGTkAy8XReoCWqH1hGTdOnJr56CdyZb6FFguOZUbX0okF
Zbhmvwhbg2/IlPgDT0POj57bmd3W/ybUfz25YF8mn2pgazGU8gbaUZEI9tug1hW9
HnaRyaxkHRyJIZWpSl9Uc575HWytTnp4vGqCfDJuNGeACpWDQ0Jan6gLwEIxxrYn
t15aWDzrINJ5BHZhAnXWlIyEFSnj0N0gWc7VMmLOHI1NDN7URdvw88j9NFAZHp6P
VSITebw2nXPDiuoU4E9haARGMK3Se6hVDsnsGF5iCVJzq1SKV6AURNnLqtKv8DUD
x0bBS118aTqoSh1ViJ9IUnKSEk+6UfkgWxFP62+a/cLkyou+A3hxL91Lu5bVimcy
mjYVh2WGegaE3YQtndO2CLDLGUmUJ95aWiUyt3vgP28mzyeqwdOJrO2MZSo4bYiF
rJjzBEeNDDLdgRtBYx0sOVcn5ec9JK2RsaVGPPtWzn35ueGTOfRkpbw0dj6inFyl
nG94Rxwwjmcqz5oxLPAHSWsocCxOx8/Mg0PpPvYOU1eUi/GlM5JC+AzhnDs3CUUG
7J9JZKkbC58vQVYNq9yDQpEZWsfekagwkvBwuPE1dDtnhdTiGJenm8JJ3TmhafkW
yWS4AtCJgDM97xIVfK84jUImPaagp0j6eZh3l329NODLDzfu5pMq1ko+FoqVlKxm
hgtclGJwcnIynW0u0LbS5SG185ixl158bVzkJIIwx4DJhUXcVaJKjZylHaLRxUrQ
muyyjIV0f12+dNE8AkQUFLOkcM3kuwDpvfCZWScRhvYLNUjqVrEo2qwKRzFFD1FY
iCfzrxsPI5F23joa7vyW4ee/wnTUJnUww7AhG4WljRRqMsQ3K4KlXGXVmvUwCCZ4
WFdI3fQhQ73+rcty94w0bmuFrxC862mX+lwMvGhxDHoiOBbJj17p/NlXHnXjjW1o
a3YFLbJks869qyAjsTMvFkqhkoQuOST0WxY482LLM8MWAD2howVY+h05BAQGwhXX
4PzsCBclthj8Lbnzxtn7qcYkvqm3JXH78T1V1uY9a2rLPZ9yD3toYOUbDcCTqC13
pDm7EqI4sbPh7sTefdM3DORSMrXvMS7U1DTdEr/pun8uqVv5DfNlXKeuAM16r+ff
9s14c7ggjpHGc2heEdeW+E5hwi7WGL0Hc39gB7y3Yswk+YartOH1e2VSnt1d6yZY
OtHqbcQyBGNAddmvGrOise4qqKeX6WI0Y7vDmWivFvmWSp0cIaKLEUhmsofT2ntf
A8sNZuNfvikXw2FAbEEVtlXzZ6gC88fDxKAOwrUBMJjsZcLzgo0fyFHEdgTN6lwe
d7qpW5ClXOKu09UPDr2bD4yU/qHdkRUPPUiV073Q0/MmNXOiukTdpbnez7WuGbJk
4JO8jrhzuudQD6FU664kEsXtC/Xd19vV+7O+79f6+qvXdyklgby9pPHkNAMdXFrW
Sg7BWJygO6af+a5XUiEkeS05Y5vY2bMPWYsk4uR5gzAEUE7m9aj1px6UOLPlT3Hm
D7k6OmN9sW72UONsWdmDhjpXXh1n4M5ik6tZBKsJOACbCEq7VhOMPJzdxKjtl8bo
KjgtEj3nz/ltizyXvxb7KBdsULEPCPDjJ+gr3bw8doRxEXgewjQ2M06vdNY6Bgtm
87CPv8pVcmFU3GFAVu3RDxqeUbZyqNeRA1QDGO8YtePWRePmyrYH5EdB4Db3ktHA
/2HzNIAXcYxOWvSg17gIoOGbPElWdKL2mRsf+EXD6kpEDvOiApYjveMmxihg/qMe
SaH9vcFbEAavK43lR+jxMmAGFFWifiUutNSCk2S3srb1MDsu+JllkkBJLGOU15UV
Fv4usaQY20yU1t3tBqRvXr4+QX/5RLjPs9ZmICMJt02rcZaHsp2YEfvY70wm5gEV
A9InYJ1XX0kOMV+snKsyJrWkj4Nxwu5GzK6RsHIQTxAF9NXY91cXmEJ6TILtlnHC
Z9yR/VeUoV10tVPZ0CzM46xi3PHShlTZgUvk+l7IDwfFuVtNjPgzxUVeerCZhOTt
zvjdjDKoVTx0lqjcBqenwVNrj2lYkDjzE8PLEkryOhfPwD6lGX7R1SeCkweg6AXJ
0yyJx+oJeCz7+gmrSmK5IyD4v1/2Vm8WzDQEk1kxNdkLjksAmx+oconhrMUetXmf
tzUk6OYaN+TzAqeX7N9/rQB2i5qyiNGp+biX6z2MJt0nYqaC5QOEX2h9pxPICgpI
joOuQBMCau8izRnObVkqj5eTlZz/keO2nrgsNQXdvz+JFAJ2yT/8jYOJCOxGkl5t
aP2jP3Uw/0GKiEGYJp+98xm7zSbyyJ3gfAHY2ZPI/dCfmxii6DqbWUwaZ07b4ydR
dLamDLcuwtW4n4eh23mXzZIlqsGYgdP7SmueWVU0R59TbezPY3IlTu9mHR3gaeqq
OmpLfaeyCcjKiC6+KEzFZxboEr7Ztv107+RBC6DVmiQYO+RYysCWNPd00Er4E2D5
r1wCOiSwS5Tm7oJB3oHNtCNc/+Kr5JR8zOTh3Gag5X5BXi9szDRq9VrJaXyNhux9
NZYJhf7Sr/lnUsiksTMFt5pHyL3XTn/dbIzxcV1JeRi6ooaG4grvkXX5LAd8ZzDo
TbPEwFwu2MxU9QfExKfBX6UsnNW0OL4JZaMRAOQ0+5AkmfwAkOcDt+QUmzbb8e5H
MJ32iy1WXL3ZhzDokTGdx/gz6zPkxkl+Z/yndhIuPmq95LRGWzP55WWIeEIG5m9/
YFm8hXMfR2zjjQ+GWF11KZ2BFIz9fh5ucZ2IxWh3839Sjmh8w6lPA0luOVtvRcbf
XTEh0o3nOf0JxcwE20srR631IniZ3cQqmAiJEqs9XIKncy3qw4q1HLtWtO4nEvq8
+Jny8jAGJFIMtofNsiOtbHRQjjApxQKesDeR3j+OzZyJbrD1s7R93TL0uThovi4P
JlJE+DLofwnj+EzB6/JGobozzDpsTKiERDBUqFLIeLmNn8OIy/Bo3swAjTzlYu1V
4dVuKvk/7rEiQm0QHjgRvlADWhN8jQPP7DS+/y/i3zc1AZpNDQeWHE//AfzfpuUU
1g3mncufDWWvBiMjsGi/kD54YHE6nsAgN5bz2E98RqUkDT75oIzHhl3sUySYFzfd
D7c+FY01aSMMllL5WJB+QO6BN7rWxrFYxYdYWL8+2rwdYbboAsrCajsH5bzjLxtN
ViYF0gXfngST5jrCNa+ZcGZoGIO2z6akxFxSjy4Kq5bYpmDVcFV3gIkB/41dnnyG
YOfqt/CqUqJleBLpdzMENlh6cx9WFeW+mWEbnLG+HP7W0hGDTI9Gxo89jDQcUmvm
T8OlLk+oaGyPI2idrWmFT+7vHBJrp0LiEYJyDn/7Y+CODvChcLSC+0yVGe50I1ZH
0EZhxPOFEpqG7qbbLKzXGozEOpG+ireoNUY1VGnZauX0BUHsNcFTQITb3hmEteI/
ew4OOgcU1x76q0vbEvz+qdu468momclMKQPC36HIJt2fCGMSjs9WUAAppTOMse67
QsSMBY4ZukaMRp0FW6yr65hJtCTvwJxQXPxfRDUOnhyh57kIPn/a27lULmfQemrO
EIRs55aPy9Qt40ThSBdCyMrLfVgzo8xp0XkosRCPuRlcR/58xg5x51HQY14A33XB
of1CyexnIbBYanaotjvuDv2s5AneALhp8sWaH0IBmp/IkAtJ6DE0sLpmMSXuaAUH
Ml0LMD6/lBXsi2KvBar8UAu7zfU9W+oW3VKiyildQl8IMy4qOPH8Fcfh8Uo/I1md
S7RC4uly8ri/kzHmBoByxNAMKH+3BpTroB11h15x/vU8rZ8FOPFO5+8ZnUCYLci4
lYHLm1rSM/Kml1cu3VcymOl/HiZbQzsWD4tttRyy6f4cz7UAAOCeyFlpB/mS4m6A
rhPvbLMnKKYyrzcfnrTugtJN49S8ihlxHz9VW8GXMp2NHjVacSJ9OBA6lBgCPvtn
IBuLF4WBZOTnctEuOsCZ0l/uEzOA3hbUbSBmzF7pTZk4Dhx4sTjKrTRfOUCYs09q
UNLV+s4nQ+/BPzN/sSu/C2CYhbzcd4fEqG0b4yP4ZX14cYYWD8iQ8S6NVWxQtsf9
bqaC5HSUApfwTWAPm1A+ZtFtC0wjja3e7mVQjelfBtgTVJMIk67uYXqKwLaD8G8X
ZFAr/iS2pgKobgI5vKp/Jjvm9DmUlpqetccE+/HoEcDhEMUqj/Ik4NCeVIGwfT2O
vZSjpdFiKXVHjTc7HyaSXDvF+SQBr/1z3u4k258U9CHp4qvNVHXd+jeNLNf69lWs
W5hc8aYY8CIAzElPy06k6+eSjjJ1bgnT7UR5sKSHBQuq6X0S8sLod100A/y5CV9g
m2Z0uQMh3Go35TK0UMXZOTg6Nmjn7oWvEr/FSXq3O+pOYLIrL6t+F62Lz3e/osOv
K5NUun6hjx+pOhPEe6tKojcVeAVQMYRYqhforbtdqQDkgY/q1x6vGcFj94d91TDC
cTrmoxpdhDWCYI8tuSC6nD1Bp5kDm1ZpvO250SjriZ0VGJHZJGcq1LCmxXrQADcy
a6/oFnBrlvb0lP+j1OzNRLfl5znb+Oir0+dqwNkJjlZdmFn6hin2MkNQLdslv3ce
TLU/jrv14yVL8TlGocyKN0nsDYoV8zAO3wI94I+AoTDy+blv7M3d2POKq04180Hq
Cl+pY/Hwlo9Jx/4l5gNHe4fZvP7wWVjHPnfIK0zLaUnS4nZkMG/l63k/e9uQPmg7
Fsjg/p8wakipp6DQbGqqwj6nbV8M0qV8KJZTFasmMsV+5Sfd3TvFD09Ef/j5FI1i
QfsRV4Edyp6S7T+fn6/3DVui6JKblcFI5NJZL3b87lKL1J0FPD1Wm6m7zrfFbNEp
RH59fsKf4pcykI25xfAEP0aBDhoXG+LguLMfkbmuodBiry2oiw/Lhw49HSj0Ufz3
R0OuxV1HoIMm9p2vrAlSa19dlJVh/EJ/FgiZrdQPxmuikk/f0vAV1Cpx4K3mg8w6
AXL2y12Ucza4jPfJSrVb6JAlGNruGzWFqtqikJv8LGUkxNWPzUKwzN4zpfpfnP5h
35HNMbKxtUAkEYTwLVdJjkX4z8aB5cPiMrSviryxuSId2OZ0025TTLMAI9IWEit+
R38HTkcbKWbUe2qQddC8fN7knOTIyOQ5BUY3Q+wJ4MacZlq246qkYrn3Cb9kvGf/
9DSohRZV15IQOn8lnFnqvnIjEZoFgJoQNEHotlK1Fayz32+2GuWFI6M5WFCik9Uy
7fIt61crTxYMC/Odt2267hF6VTMMN2p1jVqLSBVEB2Sa0A+JnxeIPL3P8XlnxmVa
k1gz5cK19I99wt+W1+okz09aPU7mSWezQJgymV1gQAUAmRpnoZvIbTzODY5dEAUq
+9CnDpAfg4qFAzyIt2Y5x+vCrtckCHGus/5nPeH/TJJNgtRiu18TBHcbMJLphuBB
1vPx+OSqtUu8lwlmq5tB1zRAdV1yb8VdHJ/kaJZgLU2Hkhm7TEG7O9oqtdXBPOc9
RXakrd3DNV1zHwH/vuKH1PTKOqP5ju15/r+Bd30VDUmi591tHQRy+5EjlKwuU/QV
Wtky+mQ7erEGuxL7yvqUjYI181mIRETmID62IPvPHvWkaKBAHUUrnNszm47OO888
OYfXUyUFVS5Wrs+JpJYoKesRjpvOA6lc8EV8qiAxDIjecqROpbyF9/jMj6EDQ8rw
E4K23h76H6glor1s68yN8csKtj19JGf6Qn/w/sKxii67KkOzIRmZfA3Wu1mv6LjS
Bc1nLBQDpbpTZRj7Y2IdL/+6FL7qMZ10oWDdoXa1whiFRucRuoZtU43tWhuV6iom
rXHWyLZ+g+WsVXkhcghJI0dduU1yqz4XSIr90zJMVQCEriRENYQADdME0r6hxXSU
UjKDiJAa2kVxTV4Aq59Taww1nQIULahaoz0aEqj43H22ZVuNA+O1mszH7OkY9gWA
sXGOwul1+wM0JyIHMZR0gVQR9CLYXsBaHWaWnD5AWYC8OHtdePRiMeUZKLqNZcho
mhb7VvRgkJmp9QsxY/QzhR9nKIbmbhVZ+efDnS+f3OCq7rJSr0QbRnHNdjL9Evls
lSk4ShRZY9o2dVXjcyGigJWdackVd352AjVvNar0B4OmgquhB6j2bPL185skylhI
kGhPsf+x39S5DESoGnzwqM6ABGtMOXCYU1GKmTXLhmvaeilBg77odpXTcsNZ9Id0
ivKuj9fH3Ui/9CsS93DlIy1UdPkD2WHv4AAaDi0qJ26YFi24tpJP3WYtGFZ2CGm/
f6ugQUKyOdiVTu+qlZyycrq7T6CUivax+N1xJL3+cy92Q+SP9b8cmuBW1kGKUgVj
VQ/k364IhPI/Ry/swb6qYbL7618nGNyr45WxW3dIc+ywJU2jLWVXLJBKAzakB5Fh
qz0M6acD0J/Fid2GXha0/qJAfwUXSc/4UrAt2aYXd9BYnIhmD2+xhppmdPiC4dd3
1Gev90Bf3EGx5/FIyVa8r8uM3qgX1GQGexP+kRVV3iSH1bw381NXsZR4b/LuavHA
x+WoHGQDnCi23FT/B8Ghsb5MY/bY/hRsysDXiVD9yACpz8wjB/H52Q9wm+5N3bpw
qaMgwvYT5/W/OtmrAKzKA0LzBPkdYTmggl1hDRsKZsnM2iN2Q4/oT0ROM/suW0bq
xu+JP99wu0Xdv7GffalgffWJ1JP9A4PnZSgIXOaPE3RSNtmXwa0e+MbZAfU1nusZ
NFvGEx9aEjmf4rz/Ix0jj5b9dtLHs7ef2AuZRkkf1/URpcK7DP53c7lRU0sTNbdm
RIadaqN1feO0deCGb4o7IwcIwveIXFSx7Y1uBAY57sKn8mznrsDFDqRX/XC95p2E
Ajs7LOBIhSooLTBrBsmzcC1BY2AjSf0JX0fKoHWWE6pR5w/UXHzxghgtXkUVXdl2
+439sJWIHhJY5PrygkUzcc49dXbmekVJUMNDDOcpMgNvpt6dyGq2aM/3jk0Jj88A
S3Ysko0mnuHk6hBcJllX41HDvl2UtA5nRMglD3uKUD7pkoLKfYnnMEgMtpPqwECG
EOEqc5qDGtTSde08T5p739aOy2bGNFUBEzZmH/EFrlD0vlgWsztCEpXLa0FNFsAc
D7CL2kjwyPKwHH1c+E4fy4nJvsj+GT0tW7/CiC1MLvjHFAvgp4xsgk2fs4VNdhpi
FMGWVgwENi+O2Okmlecq4VmMkXeS0xPa/1/zhQLsLAd7fvMGt5qrmCXGufX6pZBU
+DcFXXQS49FppbngPwlQfHq3eQNZ4YqTI9tcPa78+o39F0FZpklgVdfi5aA9tdKU
BrcE3bAPZugZfIJhwgCjODMJJGp+6ndGxNtllhpvkF+U0lYNyxOKkGBYx0kKeVKo
U7mm/nK8n/mOwwvejpzueivxyrGXKd8BDW52BunoAIgcLqR4MHYuyNQ0L8q8Kqrr
5dFsHjYdPfqqxQN0rWn8NUfREPrAA6A1eznHSO9z5xgV3rKUxFTxj4T8gslU/GG3
TcZTbcbACLJyow6KkZsN2IRho+lj+b/janKpwSoUTf/uvg2UNHAxCEVyM8UglW4A
ILl4wJBScr6SE+WGCwr1RNlFboLxEw5BYx8G5xDfwa+ajda/hhxvTCGVXIdl0AB2
naywWWXoDQGPpHfGu9Itapq7wIy186KAkVKFIlhOYjo1emFshfc1br1Jue1gGash
IKjjMapS2yujEhFPnZQYtAsobRrRJphGZJkgtwba8jysICGx7oxuW0sX5W2Ho+lP
5nHF2vnPkm9W2pGLG/zKSCHni2vUHa0vl7V5Fv5OlNvNlkt9kl6IJaay+wTQUEV0
r29ZFN9S455qd4MuFfqVYhYjiyvsuk6dEi3ARYIoEoNMXSQqf0YHHtWyGzEOe+4s
IZoo0WFsZtgHKikpivWzKBVpfudVAF/SQWMA8GoCfPsObMCcEIWkGK5wvoi4JLnp
irnpWlf9tDa28h5ev97Z19Wnhavi1f5yguO+oK633rxydV4pLxXZWcggOI7s+331
LD7Gry4cUsKjFDeqgdPBDbADJTC8ioD787EjlKz73Qz2eARmm8pm2+ToxPS/urKe
Fc2LHbpLQCjSBSWTJrqynxVBv+c5MMIIYH/gSCtBN4JTJSNNP78sCnWueW08V026
K5WqXsqz3sn5Y8FOEOK5Y1joVoUQzb0mOLt0zm682UAI8Bgm4PZVP5AwDrGZmG6A
gZUkbYGJGT4MqDtzngBugaBf2SCNOe7UOV76cX3CKWo63llMr7Ie5JuhH9SMzw3b
FINFSCUA7MXDWg3x8KvLpqAqi1ELvzNbGttf3TorAuUvo1Sp281lCnsoEwgz+7Jv
/7X/bPvDejebKiJfcblc9nQn0n3KBbdZGbqwh37w0a8BHzl6eBgjBDno1618Pr+U
PKTqdsoX3TICi9pzfbx8Dho2srQO7zRym+/KODYr1N0fkbnmJl58AVqFfDx17DwL
jrKfLnqSfu+uqmhK25KiFpRrWxkgumAm1FPvUvDkhk3sDb6Yv1UvZ18njE2RGWeJ
bTbw6ULnLjx6sWJGv+VxAV30dPsQZ7+qHjgQuxOlmoqHQZbvNEzusyxl9tpJYxZd
DwibzXrnDxeC7Qf58MeCvv5kFS/JEroAhrkXbW57lDOeP09Zq8IgL0ki01zd5D5z
0k+xVUPvXCs78dsQvY/vUwtxYoC4NK0FvU6uMhSh//R+uzmELUuGNxq77Bi9lo8X
hfI2m6s+ZYY1pNfx/r9PXPSyABiDbgocwnLaU8Uy/Gdh8zQ9X8kH+/OjLZZV+1CS
cf18Z1xURdR7Ntfiwc4rN9Dzk2jvwQJnkmDoW6KbLBpqMvnEdWrqn4VwpbRuLKCe
v1qTHuHRKXm8Alfh1dL/YskKH+yfe1kWT8KuSffvQQ7OsXeGHzu1lURkovfthovu
FWYVfmPjOkS3pBCXSFzbeog+7VZn44ihcqubeCkYiwLFsLRUFDpQ/6NxaNFQtNb8
G6/EprShseUfVjywBJ4WiHuISLBIOQZ9c+HiNQ76u9p92cuKWIUBbbOKu6ZtF8tD
XGJVD0FzKgtTQPNiOP5nITEi5JNHJ5fH6Zxd9E/PoaJyUOA/I2NFeVAAbC/p0nmk
poBaxQYGxnWllVCeA+JtHwptbiLb9C5U2W3twa979jngrwgJqUV0HRZrkK48Jsi5
Ve0D2AD9htKcw34tB0Ef4AjI+JhSsV8XCEN9roV02AqChV8RxjGCyJxpmeAiBNme
Vx8wTJFo85BpxL9oAMCztEOFpVlFhlTXxLzP40BeTFmh+IZO7vDJOu4PNCb6gaVG
e+rOhzM4NuNUWPOq6zQiXuVq7Yvhec5UHGGi8htuOIO2XeXdAsqZcEBwZ5SuWLTQ
PA2LFfNm7Tz6CDZyyaKimh9erjEwSs2tvpX7WyoRI1GKTLiudghG4KLmzSorItT7
2O5jFh2MdKF0Uhr8HHcy5FiOFzUDKV9WHeIL7KiCOWo5205zhpOzHYOB3jqOs651
9Qu9DG5us1BFiQz38m1NvK/hA2jsLFRDzFx6N/e449PtM0tMRB9774kUi3IWrt79
nIHTMQbvWyN2wFYpYwV4X0BLTHs1bt5WCL/H/ohS7lKsV6C97m65BAgtwj0LjqVQ
ngAqYIj2zm2rS+vFTFn4d15m8Z9Y3HpoW/7j7DaGKUOgTSUKubrnySBv/Yfqg8jv
MFs9/aZgVbWO+Uv8nRcHoaXOWRNyKLjT9lzclukiHj9c7qqeVOK3j2+En0l38Aa8
DgvkvZFuPpuOCsJVZY2K84KZhGWIYe52wZUx9u6DKetd4BuIaCEwt0MWsvJlwO2v
Sglgtw10DQ+ep0B7ZeOVuhoMfKLynMfJg0hniVAvNmfKYSY0QLMbz8EULgQOehEP
QDyMe48NOnvusqlO/jt73cTlL+AACwS8NRWoiIhBnfVjmW/rgB9cGJZ3lLtnd11f
fmcDK3+lEC/0oL/vbQZVzo2tLebBwVzwiM8uiOAjd2m6Innbu+9mwbBNkj/kO/nb
bYuT/TEUB2sTUH8UXD6gBJuRMnw6rX1Rxy+a9tmYEAUc8mtgt/8ISZC/klBCMTaa
e40SY510dkIyagdBK4f4B/vhnlqtkyt6aN64XnLnIXs3sCedr44WSW2kmCg1qQNM
EfjFDSZ71ePdCngAIKrLTLGFPns32DwUCXJczUffCciQEri5DONsiKBkcr5cFM4r
jv2Osbjz7ppoM2AOtfTsMIAJfzdO/Wmh5GND5Bi5oIoNsCtP6dbcNY9EhxVV4I16
zW0ED3TK7V7aZ48i4ciA4GdXqCB04dme4GrAtRsJem/KHcNysutZGCALde1WGmqz
+yYpK80iVChvnsIc35PokQ8zexOefN6shOwzzGic+euKmPCvosc95FeQUTAwwaOi
vkbvOX6klPEF9d22kIJCRk7yd52OmDmFqKVSoVfUTw3Dr/5N6nCavSWzb+EpmVev
BsR7cD6NHPGr0PC7/MMW4IDgdSWMYE54TGxEfTKnC2EgXHbYAH00jdcrMgbsDbaG
UELgpcC08UtZtXfnCukHtLvBGmQzrPpzn6YAnQQldOOOIX4f8DSuYDXjKraNM3Ef
ESSKSTadKrXMipWSsackKylYbdVK8TCoEncHlyVbiOAs6opkf/JnipheEbsphFay
E6+3zgHXkJmamZCCKm0uTLyNVKiN8Gv6CSYm9Fuha8hq7YEcWlyyLcCGGQ1P/JId
v14Rv7goEWwa0WEALavsE/C8UpSOXamU5iT1ry+YPpwBtKQUiLIUccUjwaH8mZVB
OgROvPGjk2iaP6VcHs3Tx3vknU7vyqU5/uTYQr43sSb0b/FdCCsSuWVUZA7bZ/Ia
0DcwoWuMY8LgSmOxBmtVzxi82qMYSVLWSdLEeKXxlIBnp5Ve5/Ord4Iu1XV3i9GB
W435u+YOjBnUkyeD/ylDiRemY5LFeJbV138R4qyHRleehF6rF7YSdzjEUP22J9G2
v+ykTwIktTzRHv2GtiUtiQ1iz1ZXTrkREmTzBq0nA8qzucQkCYCZ/7fHPDBhLVs/
epHW6YgE+s808v5aUjvLoAS5uyZ5ixQ8mid8rL3UxqZIUCMWwCrMw1+YjjKDXvQc
Xpm12U745c+eUp94kpTmbI4EHXKyDAkbjyf922fOlA71apVWDqoKGmeIFywOxFvO
5OOg+kfjSvkSsX8iYgl/cMOcUnzERgvcBMPftBQDdFFzrW1Z1VA9pT3FLiceqIaP
k9x7CAyBQaG9FcqnYh6u9n+HScY2r7LDYwL61sLkn2UHQHIEgooUhK+AHLGyYzEc
pqMyZfmNZUbBxk0ShI5Ds0MgE7VVJSSK24ruzpUiQQLfmcv1/PShhZd49mpN2z92
ZgkWuG/MjQ56/Puk956BoH/5f9OV9qouK1NDoFwVwm+R9/3fHqWDsR0d3fg2Mrjl
iylHctLNwj3t618E/ODZ6TG5daCAWdSg35Lm9HOZf61PWduanS675Kn0jsxvDlUM
v+t5iZU9dnAoKz5g/I6rmaspaXhrOIqVbSprBvjuunLDM8UJPb/g+4WYEBQ90YbC
KcO1dgSDJDfkuKsTWv9pOIcnV5ejc2g96x5/RLXd5vGFvAJiyzpXcSEbUSCQ8g+R
3Wqih7ro6tHUZnTnUYLUY9NFGHBz+VnvWw/ET/RFwoFARzcSS3ytA5LdHLz58KKT
ickYnxVpAWp71Uh+rpf+ZhoXvDLrLWuk8TJC348kwJPv0KhW2nrq34KBJeiTdYjJ
tScVNV5HP9BU/XIJm455FD+2QBWL4B+AYa8bhAS4GQEz78FBGGSKgMMVtCsFcCop
ScmVHPvP/yuPIUCHj4lb2yisnWf6nRW7vEEM2XsOaU8Y4UVRJF7qDg99EIpArjEF
LWG8zpV6a07mSWRKBrZKEjKdRrJohiXzeE4JcED89ryM+Ebm2M6MZcQTbwmLjeYE
9mbM4Yrnj38lhho8CdkFHbaDddpBamgBUdqXw8oJA+UFi0zhsJqbkbJUhblL1P85
D8sGxidH47ugtNBBiJQpK0Fg/JT1jjgGLfNj2UHMudG7EoLQEMlF2ynYCZ0wWx6S
I2m4Y94Wi3XMcXoHK2yOsiI+c30PqhBo9IkDGOx5LM0dk5HLKxmZ12g4d6K2Xqcr
Iy4ecK3YnJCDwyON8Wu4p7S+3SOSWgNZ3t0gN7A8fJkLZmxzw7OEcNxFXDl9RXOC
tReLGG3E6jTESAmyBP1h0m8znAXtY9hVf4L9F1atzJxVHtsvLkaJfp12uNX4szyg
hg/9WI1mStidKh3ob5jyy8PmF5K2d0csej3zjFjA9EVbVbgxdscmgeDvwIHW4E/D
QWKTn/4WM5oMDNn4Uq6IWPZqJUYnUsxJ5sgKUcGC8pnnSSuyKp9tCYA2gXbrBwGG
ZArr3gcoy3G1RC5rx53umbbMFFkeovUh8iZwQSd0WT9VFdtXs70wfInNhxp8g4re
5djsOQVzk/QMsPCPrpi2FSiiHcyNxJgDqq6JxP6rqRqP/xvSbPpL56FLfMFgZ+Tv
SMKbRMqPlkE4ZrLJie1aa9L7nbkDoUO3/lAjCF5a3Cm/gc2NdC3goIess+B7kTfV
vpyDWfOh041nilDzLVqwoDBvZL4YEEOd3IBdK8aow1QpKnTKzbX8h+6VlrWaVfd2
MlYJCEdXC6YOWRJbYqcMIR5Yt6gdkFy9HsWqsyQ0kW1YEMn3htvyqnWpGuLJo/WH
XYX0V5AWar7n0f+ClcM3zG5FjNXFeR6dtL16B5UBHAog+LbMZ3f7vfbDpapiRBQA
JYj67XaEN62W89//ALyp6mdVlSasicck2kOUnUNw/WPmx8qq3tFdW8+dkfuPeClA
6uNQBSPltxsdc3ce4FcutEZq9+Q9kOrE/Hffn5XWkmde8ac74A7ksJa7TUWMW+fT
9dLHT9B/GoCrTAdb61WmeJwmsrTX5W3UDQSBSG4OtZQoLqqMPEVPJJ8r9QtmHftV
e5jM9njDXnDJ7f86ElKUPZkQBlHksp1/ZHwNUKkMwgoVOGLp3vjoEB77nvpzZLED
q64uTwCwsRZI+wH7cPY2GUMLQk8+xR4fYXBpO4dfukzw3rH8SQuUjmHzN5Z4jm7V
ATJ29pGBqL9irE8b6u75YLNR1+WRNoY2x2w6g9imJi7RPXQf8jjCVvIIAHSGHos4
YHKlN3mABI58V6hFK30sWVxfVnC9lvWNK9lktsU5Gu7C8QvAytT+x2EfPTmmxfB3
FfPD/caS4vMTovXkouDQUL2UKkh1MgtZdxM0wdlPCHlvyKOEoyy4m+ubmbENha1w
h95LKhrEqwu9R20SrenwT1q9skqvAMFITawaieSpKXkVSrTVYTH/EjnbQPveO/dQ
ssnmxP5UXiamzFictowUqwaeluoqCCdb2JNtHtmZCHWkAatbKX4TvF468z0U5ylc
fcgtZbSr8uQIyd62W5hQuckyD8x0TcI1/RubwMTVadWDScsnNHZ1FxSHJqoihk3K
M36GWEaaL0SCa5iBZu6Ii2gUATHhgXJfPDdFim8msZeGxKYqzi3x/ihNv3mjPK7V
gigBglEnLh+GBsf8FwBLx/61kiYm86ZBN057IblOg0ZmLQkVnVg0g+BXoqAF1SIB
2STs0C6Cl3HqpTXIlyIqBG31ngc+wZd5gRNJairlkoYDZGWfbZg1pLvh5RL34KLI
uk3lgnGFEloutCmL2ViCVoK66pDQ/aAWPTzM7hO9BnSIJoY487inHySGTbAxBjYc
z1pKQ97S+CcG1/KTUSkCYcN+lq/Z08z1+veZ6vk+COh3QskuRQuNUZ/Sf+dvVkDh
03+Uz4vbmQ37131S2VGPE0G1ChcAhCYPlrD32rutvrgO6nct9lquFChfyRRvZjKL
MRq8fdQZ+6giWEiXpIcKyRQhgehKhM27bkXIBBMwH1M6he/e4EI7zPP2GgQ58RCY
3sr6jzmk1+lrdw/jB0Xk3KKiqp22aLjFznBB7ypRz0rLd1yb3ClTKEf9Uaoov6AR
gS1CaJ/GWEagCXWdKkkonldmUEssH5ceSPlxc/iP3jvFGrpyIJGVb2TDx7E08rag
iwEK+A1EPQLQiFWda3D0z+y+9suuThAroxNbVH+urBLhUuOOHZMmPGjRs7IJLysE
k2BfX8SrPpPb3G6TQeLc1PTGcxe9fPRKaGSpLSIUzyExHaY0GU74LP9JtTs9nvuz
Po/6S6NKAwFhiigJuIuoVfZqBFejCYfjW6mzGJqvtGQT/uVzC/Phv57K9DAR9Et1
aTbqIBItICfgaUVGdDhEb7voaBJwbl8Kdac+dfzAL0HbW5IBhhnD9wC4ehxPJLAX
peaAth0zE3QdsGbz3HDO8fJHmoY29OdiE8ZzWWLJnGPG6WHFzxdoUFn5N52zLhgR
5z/YcaCFZUxKq1WDGFqQc+fRA71FFM7KmxcS2V511O3W6bC3JRhCET7gkg9UyATU
rUjfNo3B4wl0VvxvTSE2WlmM0ImO6ht+UJgh7bSFwslohQX2IieNCp8fcCXZNqDX
FIwenQPNHEZD70CZbjGl2oLgXF0t2kOvopfuoLZzwYzvJXZ1yCJpPfUE/E5chL0w
UYxiQDXy6VLwzVS8ODfRp0/kEG66rX61qojj1tmjXT6Ted3Gvh6/tFILTyZgKiMS
IzWk41gya3fToMlVYes16mfvC5bI06eXpBpx/yuXo1psrGDeX48hppYptCwsvz6I
HnRQKpRJriuu3f9MlqfUHH8q8bGqJaI59A+hEdyy6DmzU6oZ2NhrnIOXGgDxaGbm
ayQFNwTqjNgPBhCUVvHiNVz68bC9i6hwy+pWpDIqjTqxKYyVguND5gZOjCdUoFGQ
RfTHUWYTrZkIGnjVvo//tP7qo+xqYAVwGP4xzeyEVHR8URy+M3rbhKrGtoP2rvFu
eHBNVgMd4M2+a1hmyMUausmNbEpdyGuxXVVZ+wTxaB/4qemDlF67mmd6hfdPwlMG
UhYuAKBwCOPrDffLAWCgDTUUjVGTnJ5GRineCW3OGbBKmX8p2A+EqnVAwNmcCXa2
En+AaKa+Mia5ZAkNXALg+Rcy3bDiaiGLICKaj+we2Sv9H6+7H/04UFTSe6FdtJvw
09gwyJhlTUZG73iEUhnVbDbljzGHAl2w2C+Fe8CUmAQ9m12rIHqPkbvxemjON6Ri
c16pUPDpPGoGr0WSSUWcBRUWG3DoxCUtrAPNI9nvroNxyqdHwGnYJydkImT4qGM+
lewoqCLCRk0TAk18AycVRX+ZAjWV0Hbwt1luWTTaxkvUINUyf1G+X1f4swR1/KUG
aAOKJ1uPBBLl2o7iSVNRmqFeB/f3AOkNG0Hw1rQReuJpzoq59sFmDwh1AQbIy6W4
SWOYPZmFdHJHBiPEvHhLZ6+gjwUEn6FQIpRdYrWrMpwKpJGEiEZHmi7AL6pTjaxS
9RzDE2FBHLsEttYchvhkY8+BDSe+Gp1MlGNJwCNmicIiuNQnZj3WvzLtSexRT/aV
kavLuvqciqbsMvtD+JPkdaFgXMZKmlJUxbe7I1xs7JS5Z9zu1LG+GdVd6G1618RW
IFu/YkIJWIvayoJZG/pKSlkiZywvUtJlAKdQY+HkLGTiyaPUVUM230o/WwP32zZm
TFDQakbEpFISr/PS6KO8qMPUz/O1zwXa9a4ZndCS3JXBgsNIvZN4ecFBQmHkb+nn
OHaaA7taK+Y8E1PTRDwKMwXtP4oA3pWGk7odJ84trkHRQyXU2h/ZjiGKzf8Nx3FT
XqJON0ddRqy6clMJusjq1kp7rqGlC/Vvn8cjPiH/JDeSXuWhkNaXiTsnwCubHf4a
yg1d82i4xwGUVG8Q7OLEBbyUFGfXcO38xrhX85G3oG9rlrgu+aLbJv6fFSB0dp2/
+K/ZX7qnxhT7SKKXfHYoX1a6ZyrBSWxN2Ku6XFPpyUWudaKzpXp+aau/fzMpYlaL
vUGb/eGKZlmUEFRGywstfMTRLlsyZ76+7QtLd3iGja36hssH3Klb/T0tQC4WrIVO
4YCnD+HwOGenXk3kMknTa4+0RQ/COpNFlG65VUeA7bfHDMfDd1ym0mRYgIlc+V9c
ZhJ91bsjBVBIZq3v3guRsUFXVudJ0bNSe6tT7XzzI+6lg1x9BMgZaYFluajJw9Wi
nX46fQceLe6p0bTybVh1IEa/DRKTMXqGtV3YXZdLHJ2a6zyc0RyEsFTSWiORls+R
uA1XHwRf8tvx5S6xO5WXVM4pJLmbK09Pizfg0VUNMOs/nGn+0oq06kxTX/3zRv9u
GiGbmumHODFbIA0YtJUk9DkN2cYqif1SpWHSp4hIVGOBLJdWi4XOyl4OtTnLQXlk
zB2LPiMHFtqa3eMkuaHZAm8CJRnKrvHbD0+JdzvW5lXPtlzKyXqEq8CdJQIbUQ2J
wlIkjOkCWf+aV1flzlQDJgZWJpdRFWCRTZS52U7UpngmlsdorpAW9zv6NPpKnNd8
srKqTiOQbw6JtOTkbb3GodtXeO+InAxK6LU9gH9C+r5EH+3MOHOkGqFD3zNBfGpX
wfAkBZrRDdo3gXlhiHBtuXgvUNSg248C8EmoleDYV/X+hedJL4Hw0JLOJWIe1TU+
mpjiC4EszEmiGwO/6EE8uw6z1nwk3SNWfVM7d2N+MiIYQ58UZvRSN1pUZE04gwqv
9+ezqmEQKcH7Z/Qk2kTN6zdNiavrsdGPIT0YIJvy67QU+kQ6iit8audDPndyqKiU
Y8lHY8w0qJDk/7S3+IYWrRX+U8amIPq3LzvWQ86ZTxJmxukwLu2rFwTazBiHQcEr
smztnIMae9DlVI7H9sOdbpfgI1tHwruGabBbuAaCidCYY2x/ZG5fSTim6Q4+lvAS
YoMx2Q/4LKXMkfqO7eVZIJZjWWFITQn5ujh+vwmIto6ZNdnuRqYLIq0ZTnFxW2pJ
jhfboYtyVo80DGV3ChsQXBzkNwLRcqJLo9N6QvTR2XEnkhqHP9c5JpBhXH/G06xS
QK9uc/cfVa/fGkaB2MSZ0JoPTITiWtIXYvHP9MI0+wFqFGtGp2Ogvm0xPau0ri4r
UG3yQMxhzErp5HrLSetdvP/JXAwLd1xRX8nPTQj/z24w8Yw9gwBVBaSGZLwH3kWU
Unxa/b0UhWhiAhDx9dOlZ/jqtivVV4GylFF+gnR4vhDYkApxxT7VB2jwWHvepEh1
JRd4ufHCx5nebCGeIzq+mUHPieja1B3WtXWWBBOspLm70dOB9bDR2R7Tv+mSG48E
K6v1a9/oowOoc6YeTMPyythMl3bNa/XUVag6z0y/cEfO9zfHfecgNOVqk1o6tAPN
x/2e/WTI9QJcpiiq0inyLt4jlQGm4bI4V1gQNUOAxa4mqdfkbXS+mU2bNii2RBgf
hx0HorRFGEZ2vXhQrpTNE7924GK9hJvhf/Aaxwh9punyEkDN72tKBmLSmGQ8TJDZ
cT60pDcofHldQG6brhLtVyeiC3CT3Aq9IGuNnTIDWF/kSw+La69UHvFiiVhXoSHd
TCCT68D4zoP6EPV5k32jXlnO6Nrq34rDY2BKryzwtcMIKAmiPHUWpODOa2ahMOX9
r6s5sUy1cclan1pHHGEqDkd8K5YdETU4FuaLA9c/Vu4wPOAHusrjkeGPTIvaLLEq
mdZXVp4OBYv3ZIPj9m4QBAeesxCdkxtO1Mk4hOlBxSfoAhmT04YitBXMumLo2Zws
ElfofzdH3Xjovm56Uyy+6FnCxmLQmCzKAmMctYb60ULTKs2CRA+uJ/1+/O77UC88
EYuh8NXaI2JG9ORho6lZk9oUi74U3apY5gpiKn4hktnNu0HhWP82g2RSdsfvJCao
lSPFem1Mv8j9MovF5NdaG/zdyZ0vP3r38rT/LGGAwNLMTeB0i9EJUU9xsYDAth/n
RgVKAnef9XVY6cXEXx71Oe+8p+dPnXazcQTXceAesTjkNMiyGWVYEqyw2XY2C/9P
aaMqoDVVYnXUFboRUW4ULfWwHAxfV8ZGy17SCEpdGigDJeY6sbwa8xRjDh5LfoBO
C7lhSwDPMsWTyl4OX0ws0xrN8tEwHE5obU1N4LpsYxu1KY5yGJ+wfqB1cS5jNipz
Z5XUlAgF7YjWRbd6uweR/eCQ1CAONQhpgDJWXuxmTJyDW98TrqxRF4E2NY2QqRD1
SU3D7pWv61fGslKYhkcc1c4rI7KFLU7vZhXUJ69IjTQlMRembV3P1MuQvPJ/1ohf
keDwey8tAPVmhOcSb6EWErjzHjHBZInfYmwLySH8tjBc/UJ6HzoWXWpJaCKcBqTd
0yvmCh9BoAS6TbIpdSTQBDVTsskAo76KPvmD+obqqSTMhf/QWViKbOk5S+mSiODF
XSXzQYZeZH2t9ufb0u5ALDRP2AVx+AXXc9qeG3CwcuKyemOnIATUBMSTuDHq6xOc
ptzJFlQztS/PUfper2jjHIE/NXZXaxmpefqa6zPCL3Y/zb8Yp9nZKcf/xii5+uJ0
UY7RcZ3IAv4ZArRefi7/ZpLh8uWrve804OygYQiz1hgsqbcBiLUr+XKnp+E1XXs2
hGjRe7j1abLEufyaVDh4xuTmY3LCpV3EF9VUKC6a0xmPgTcYnC2DZCrvv27paUPR
qmUSzml8/FrVB3L0Yo6h/lLxcRCss/0pCSixBmDzBFm2yDCVorsmNauIp2vhKiYp
psk9lb/EsIADKW5aPggLzZCm6vDd7dTbPnIFVqITuv7ymJr02kCWBxZBkamAKbCI
dGkW8QAFfykQo6V3z7O1wBfUEEL7vA6u5wVto1VreqEuVxjDUBCZKQTslqck0DF3
p2/yf9NGFpI8DN0KJHac8fXz+JY8Qojm9eyvMES9wA5ymIQomJHX0J/j95UTEZs3
GdOs7FK63bkCF8gm3iYf4amRYyAM8vkPZYYQ0dninoVfciPEShJn6X+zFm4I+yQ3
FIt4pp23fEQxp2HzZWw3tiuWFRRlKRBRn+mgCPGKwjxPsf4Fs/QbYem8oeeE484v
xvYmQ44PZaPNjwmuO+RwNzZE6U4E1yN6kHXkYedzMI2Jl6RGs/HD/pwXEf38fU+p
Qemgho3Pt7ujcYP5Fci/2N30SnMgOovlQTQjWuCRa50ObM+vqLy1Llw8NgAIKJlY
fUg2U47a0EG0GJ+gFQdW5BO2nM+JjSaKmSTmYjNCWzKAIv5rmbhf1sddBz5HKQ+9
mw2sF6xMe24Ba0b1Z/ECFPsyYmciV3rl9lx6asaWkquCS0Y42DCqqzswCoBiy+mo
Erj6WKXHfqx8/IlxD3/2DUU8KlCxIWQpycNbNDMwK7tvDVsujUwqBrREBxm8iUsP
P5rcjpY1Mf6R8tWMEqVTOhPzPd+GBzIPTXlYUlbp7gz8We8MVAHeorm2SA4ntnrh
OHQLBfAa2fNpmMANRIiC3KdxhBFvIcP/KsuReVVjeSe8Y3gQjPxkEKWUmfI9DLZz
yQT/vN+bzZoXopwYQE+ZdOXJvVLCfQldvliy2+YsVad+behicQCcqNmDPP4j9aFD
Jo2XTRwMgEyPvinXZAnhLua8wAIgTQ1mspJI5wu5ufiBQrJbw+uFFIha34n9KZoO
3xotIOrFJmTNVAb+YmzTf3Sq10w0scll2zOVAXtLIy0QIXVTxwYcPWrKf8eep9rr
83Q8xG00Jub/ygbs0gXIZUPzWsAjKjqSald37F3xREI92YYhzsCOyAsiUXgcnFjW
mmod+thMOlAA94yjgI7r29Q02aQKrDMXISAJkhSgogIhV8CYnH/arId+M32dUvvN
xH/yyR9RT0pBfoKtVLlUG/6+nhg9hnwcASKkpexwt/qX1/ru31FAly7vjDlBxbri
nJJGU2flCLaonM9Wp08M+dVP2r1ycflxAJ0Q/Wz+vrV5Rj8c3t39XVYsrbu3XIka
pu8i1gxurx7pxzsUl5Xiy0hop27LJnxFkl+4B/fST2jgAdcb/0ZmUbYf3MKpk2TL
uT/0+aNW06TPyyuRd3WOvp9P2gERvFPhuf1Yt7JGeyNqOZPcs1mMjxCR08UCmDb5
Pia0d093ZT985nSqZUVA381KEI3JS8tm1isO023eJQIw1Fdj2KQOEYlN7/0FSJYl
sK6tCxixVtJ/x0URwqpqj0TGHYNSHyzFhyfHx9HUYd62//rlH3SnhhmZy95Kqa95
0WBJWNmJvAKylvHSRLS8OxKyhoPCkdP50dgqwUCvciLOng+rBIJDEj0lJVaoKTdX
TwmAPUDLI1DFY3xyPWsKeJCdwpb3R8BaIvIJqNoFJ1P53XTYZwleEpSOmnh1x4xp
SPLEkHJPVhZREWGmAqgRE+d35mYB7m28iIchaRakyryZxd1me9YQe1Oa9IKwSxBQ
S1a+O5P+wA4JALdk0wOXm5EN2+Xjk+fcrvY+g8PM4xa1z7M70E7YDkhi0Uno0t6+
4EB9qE0qV2mJ1SAJnkcWzwg2oxjNE5UUuSnjwyDkqBSwfDypAwJF4FoHF5d+jlKx
wuVMC39vl/wdC/flY21iQ5GnIfMP0EHPDLQIhQDbZATTfRtr8zZxbi+PUINt5DQX
ahOb7I31TEPUXA/VPFE0xEBLq5QXRuidHcSmDa2Fyg+rOHgLKEuDwIplw4/o7mHW
ho1Ni+DVv5z8iRc0SDTls/w4Ynk1dumglnHUMryhgHye2dO/HbdSfRZSXMe2AWtU
2DUrBWpZnhecTKmK0d8dK6OpaC8K+/kXTfecVupBr0eYtb4Umc8KTLRCy3o63ZAc
H7PjzMF203Gr+b+XZJjA+pQ1hEBC88d8at20aEpeZoo1wLLuIuparyxY632YRmbJ
GsUXu/r9aI8ABhT4PjrE8OdLDk9RULd6w83QmOBOHfuggSklQq8oF9Se4F9YZ34+
fn+AE+80v4OMTRxnF7htnzY1TDoyer10+n8oaaOsbEMQNn/hlaqIjBERLTXoTxuN
+pShtmu2ZK7rpyjsv0zKA1MZeGO3uFDBIpLAVRnTz3a6M7Xx62EHg1XEZIkZD/qO
wEByTy65y2U3e7ZQwuAZbol6wsQkSAYaScoJF5PIrs1H810n2RSBTNyL+PBgUcMA
hCmgFu/0zBI5SLDW3u6PaDRXDe1+ZvOVk4DAjV4bowMDawK9wcQViEnhZxz23FoJ
4wh3haQsU14a8KfrRnXCJ0NqS71/v5gUZukfDa9Mf3aGi/pb1IWWhZkSRO9cIFYA
n/nQUud0q/KNldU6r6BpIx+73HILha7ntRud7QNoDmiIDSzU9w5/EdGtcjEqXetJ
49RYUKiTbeUTm6RrknX84nI8eo/dgJ4h49pSnGlY1DxPsZpTmvkPi4FxBUOHgvEK
XxfiqD1MqO6/gnT+8ZxNYrvuso/avCDuu6MLhoBb/Ytf6FB00W2DM+ny45WCygqF
tAooKuH1GMhKyKKsVTsh9EX7h1QQU9CxrOi09JG+ZneSqzmxNOTN9RbfbSiyDoka
fREJyW/JJBKisQvpN2/rsdn42v35jNUZcs1V1fOfT9++TRurDRRZUPRrtQokR9uJ
QhveEHBWBLszUd4cFxz5g+4bO7C4eFZ4jkkIl0KGgQogYax3t3KRhEhAlNXsfQv+
jciOjGVF/vMeK0/QE0jrvSD82ZvEGkfTmWIdZefKvs/d9lSOr4oMHj7K230kCGNg
IK+iQPsdihyKtHmoVatHVhCbYv9BZNQ95+5USwr1dqWfYy/RIjTijoh1buLOIJ7m
LCbiZKDsjhAXQqtoc9aEeETUV4mzclzNFLG8hK1smbz19riqXjQIrR3+qkJDchJS
qSrdySGudNOs/tN0kJyBFsvQ5sOZdYmHF8UDm66C5xada1fT1oGfRxZfULFXLHYm
3Cdk9NwqIdyGcYri1Ko69aGoRe6O9df57Ok+K8RcEvqItRzKt1Kqe84sriUzdB2x
tWYT1Ws/KHJptjLBpVbldAsY1QPLgNCVYALN7xYBQceXLxuNKeGLWYJAOsPAIxW5
s09yQe+6vbrXMqXiRDSfTea+84THxlYzupkUQtD1CJ4zf80w16U87tWuApeoytlB
hvV13nPyGq89OBOMQg5wpBsrRKN3aArv9leAt4nEyQYeMgkiZw/cNR75gBdKQWtH
AwYkhVN8riR0FEgBo4/GEDNi8KDcRVcGQtQEFZc8foQFNm/mOFyQyi7JDTdiEYO9
OJdn8Nq2n4SqYk066eJVEgpKMepsJeFX60WKWYcHdBV+fEhwgwUX9Lil66WjOawl
e7Or4jFWbOVyjWe5ReBbM7wLB63lJtqCM8OQOYzWVtpNgIde/OjzzeFwZs7uxhRP
9/8qgasPrPEpk2w2bVG6jYyp4W3zkdYgKsxNL5vo4rYA+sPIiRIZ9Boarx0QaWPa
oNuIHzN98+L3uppoEg3j0/yH987W8rPWwukKzPq6PhfTH1sQIpJxZPeHB9L/YhhT
61HyyY/pxUpUd9lULlxh2MctCueMhgfnGfmdKA1TwEBJwicuOePFBpeuPD5LSrpJ
o1ZcfP0eq+RmOSgOKXRZ42Tk1v5FI3GPblJAXDn9t8fmTt9d9kuOm7aR4IO1MX4L
eEuSh3BzALA24zOzJIuek2pMPlJNZSv9cTkQ0XEtyZY5DSLqS5pFprYOhbuZ9kt5
ua5VstwLZMAvXsQCxbStoUGAus2AvrWabpfE5srKK9yMqNSgBS3VGQlbIrxvPyjf
vXk3PYwRg06+hUCjRDNOKMPCPVX4Qk0jow2nMQdQK42LoNchuH0vzWFzTURmt1kt
JL3t+TZHHHT2YZBxQ7wmucqeSIZcjK6a8fDvrZbjJdZ78y3fWpx2lnLgtIAidrQv
oZuLxJc7zkp1JKh6qn702oHoWc9amFLBdrE47YDofD/DVpcTGbfIgl9NHOGVmXIV
SVKWMlEupI1yZyDCdh3BO6wc11KzpMQUlB4nA0TUboA+k2GdFo0wJKzoFUr2HOLr
w8vOiEPdmvuFIaPJ0JtiYt7Q7D5E6xO0zl7s9EQJlNzAUI7aEUgjub+Cg8lTDZhm
u4wO1wIGR0Ez9ZkVKHeYAGhYKqEIEIX+35AAcQK3+P2stoarmjoHNTfVq0LnKatM
PHcZoz3cFVBVsuH6r7xWdPi7UleXqZ2sHmFv/L4tfSIKZAhM4KIodg6izMqlQgg5
ExMfICavdOkjnAf1n9CyIqZGqinngOivi/gNP/2t61NTisVWRtNn55BlVvZ0ivzW
9pZdjCfq5SUuZdykdgPWEzEPt4iE5vxIbL1pJZTNaRR/OFrlivjDb0GXqOrP/tT2
/cmxJl8gk7w/JKhxwpQYYEnfObiDmlPSfdehrE/BoHQo0NLxYqDrSTVDNt33qEGY
gayNKD0xU73UusHVAH/gzH9uz1MtdZFtLwDKJtYxszdh2IhxtOZe2PFpR6eVKhfP
lpb2hJFZwkG2jXhwwVT2Yn653RZwo/KJdRmTePcid7+aKsATRXYzPPHJxAqke2/u
2LIRFkTcPUmHYv5srACs384vJU30LlTMQHbHKJ31PY3ISexgx1lOMosXsgRC9UEK
3LCMwYyzp85R3oZlGL66QO4UePM5mKfBAgAZsHuNrcp09xwKwRdcXjssF+fadHm7
YvUd1em7EqD+9kU3lPY2WXeXqc/uo7pTeeagB77SMjgF0EkqnFyF+NqvtGkcjKeE
NOrGUkYcTuDQ1zAsIL32BJ3yKHtypxuPUNO+SlDaplR/kC2tLNLHnDaXoP/hv/ld
68AYR/YKf3q1mGiGFcDszKZoTD1Cfcp6dApXdSrvtt10IsjCYEueGaZM1bZhHoSl
c/1+/YxM8kmdEfQrhr+l5RYSgreA7lN39ojDPl+IeTUfBuJlI36/lGbaWurixF6C
XGc9+BSWgN0P9F/LFzwJi3a1x3wpuyP1t3BNcXDBL+VC5ZJ3uUiYHUWe3XUyS+k2
8rStDTveGIPl3chra9qNkatgqFzq2nyf54uISxRts4sH0oB3d0bUk+6JU2jo/2S7
wz0yq0F2dE5XzW3gXb8AV+jJnmZmXDNf++epFamw2+OUlU710jNyb/oqQemC73/U
+uqGhGnUL2zVDKuN6JI+SfK+o5QZDJPQwi2KM2RiD4dwGIBtWnAo6joP1vbu+ZpN
rkcHa2oE6R2eZGRxgrt5zRtLFZSYdLh8kWYMf31OIShDjtqg1h5oSguhlKGIop9x
3GqxHxj4zhtyCyD6SePknZeOM+MBSh8AD+IKjKy/tuXfQTpFCvx7H0+qJ8L0qSjj
HTllZ3jW7ArbZoUSGg5wyy286Mh1Ej9ITKWsuuXnTGt2PVsJv0+aGd2Xdh8oGI/x
dItdk+7UMbWHkXm7jweVT94HqyYh4F7bM5/H9yK5/owxpINwWVNZZ/H07R6BKW6s
jVl37LTFeGS01ejmbp8jMm58mX0B11AuoGwXGyVp7qRtmv9P4Ij71YNT3VPzw1JC
Q5UU2zn5oMRYe/QDDveDWfOyabR/yUKYujaIzu9Uz016eOx9APPPA7pRDTwaou1V
Fv3uPr2mTYnuIYbysChVrNxrPv+nG9l+hLluxI4nT1MxvsX9R0FhnnF9WQSwIRzU
WqavrMhvmerLyHO0WpExzHYroMF9qX2tQ9GBRuh64b0UMkTEiMgurMF9FzjJ7Q6V
3/RJLSHH8x4W9ibwguDVWVBIR4c++avOrD1/I6JWnGfr7eeQy6II60F8KAdq4y3d
usppNeIY6b0kltgYt7zyZbHCqDbuRLu9sVaAQN0pNut3Er7iOJq3VPnUQq3dQmEY
xfoRx0rihdUagqliJwxziJnDzbqrScflNh3TJYYk6VLa80c+TH8bgciPjM73Rl+x
ESPp9s81bVUOzu2aeRNkpWHgUV9Ahdk4TQKA/sErkH5UKKNPt+rjQ5DV5BFeWj9D
wF/UG67h45RDf1VES+WpZEurLz++Q2/dU2t1EYWB6U+z8nycFCQ/GAQ50vWMQYuy
/cjGF3iNWxfcgIT++RanxNQhCdxalaPuQv1RTSBFmY4BPnvKkGkl/N4hXzY8H/Jx
lA/N6f63TIsFW92EBPya2C8zkuDOIr01UGDNRo5Bgv6JJ+9of2NE2nmXF4F3Evoh
X0khSTIVh90aiqlYSoeg508PB5h3GrIlSh57ecW5S0vamTpPDYQkmPrJCoQVsAXo
zlgXbYZ0hKPeJs2TdP9LIuThgQyzI4bjR0owxexmtQbjO4BJDFujUytTbICqMQ6b
CDOLTa1zT4siYJnV5soEpYjb2GPcECIHN/Tb6fGp00xknBbmnALJv3JLjMN535az
Im/7Xq+nxkONJgJ6QTcTIENJQnp7Ls0Br9SDilk+jl5VD1b9sCwofQWro5Z1yLWQ
RFN5cLBUoOTfDWP90VKk6K59wz/pt3WF0CNXK4vSTx+zvUnzI2EDx7UW0HbIGInY
hCJpH3lbVo+Lg8ffcuZiHwCTwYcvSt0S6bNiaOzWfvA/y68VV+5ZZU50Ow6Meb7K
ZIaOARitESG1l66sdp3rpCy+kI0n4tLaD0zyuLHZVGU29OHx8g3vhgK+hSFk/Mja
pDbPkyDdQnDfc20lBg+hHDZlBhPWtI060bBebNTYqAywtsAOFPFGAKw1V7tcwPDU
W3EK5/BBt2dvg6x+Ddkl86GvU9pPMEU1L7XhaelbptUCDH4qMQdzRmQMvPaOlE2i
WgehodYj8lILLldlBdxi8ld2TxE1RBJnR1F9R9NsZKI7MHAjsjuGUDw/RHFJja3b
BIweMX7q00LAGyHNTmQBD2i40Rqx68TPhA2U4olvgmOgnhPGMlVwC/2WMidz6Mxq
uZ5Xy8dOSJDpJltFt+RzDlBe3BD/d1rZHf3NyIjrWuy17tZGh22Hs5GDQdpeVVyR
OMLjdUFktaJCFaiL6fHBeETlAtdojJoFMHXftQKa5FUnT+5ZrwIpqvstV4bIMnVi
yx8Zri4kFH8f/pY7UHjux3RpjqRdmdnPL2b5Px004KEa7w8/X4C2vE9ro34mip8j
3P2twRJB3two590471OVR6gDzxgOEAZXZ7RBmqkf76jlwkvfKmyTGr7u7BeC+66b
ueMsBkBUd51H/76T+3RHn1qTkHuCaIWX+7sVeg5mr7ypL05aNU3JmGbV3N9tAaMl
D3GwcD2LdceQ5Mzt2kpO/8vobGMG1SAQi9UOzniPa40wOh1cLNClsBesDa0qejUh
qXc30WwXbNzrPLJUuhEU1V6h42GYqQdSqkO48QebehPdDxCvgpN0gCsV5DhtzTJR
ZvknZsAWv2xNPg3hlR1ddHalYqS4Ach49rpIoXpu9G7bA3X4OEgoVkBt92Wd1qaB
S0uMAtyMXB1r910akQKzdcHUVPs/dE9Tfk9X2VkofRhWZ2N2PVrFGi0lCpnO7gV4
swaKL0vlSKFcn4O/RlBfqiISPfViHFaiI0UXW8eNRmUO0Nt0WYN6RTVYjcE5XRST
atMVtk2hzxkJxbislEqFQqosbEoceKfv1GvaH2fmyInb32LiSDwALkA4su7DmqgK
/a4f7iPHQuRL9PGDH5XxXXKebetlLHP9NpS76tc8/GEi43TpUWz5DzvbVUWyDAc6
hMIeFz8nIsqTzAndIxbmVhcgYQS7lp2nOqnuysEjFUETE5sxkp8Ly9VS8sgtg/DM
VlJ6hvmKTI3ThKIfb9T9T9FLD7Q2MvWFIGBqW+tzotjrJIp8/cvgG8sJRe1sGR/F
x+xibfOVYNJIewXh3zU56BSDe4qRE3q6R+cPX+6AxmzVnBsvgjY463VUU92adMD7
TKl/KlHtcIYT0oLbjHR2/mKBgf49iRnlPVrUV3c3e/0H361lOw1JsQ2bCdxBDCPK
lDAzS0X2yl9wJ1u9PhADwgx90N6JpDjhoQKXMq8tr9gFI9BXBOmV02DkxjnMg92X
nbLgNK4fj6Z5CA42jppmgHJfTMkSaC4j9EAjNJkSRzzTXIeKSQZWuL0/HaTrFfy0
aAIqfTIHwJKO8+b6K7oZCPehvCt/o9nm/O1pJDJa2hgXcBGbBF0LgoXw8nZVdeuk
KxFuzd7J4k46eV/UhX0HW10wIqWp4k4X1iDTlE1j+tn1CIAlOrvD1yc0ns4PuKU+
VdLAM1c0+ctosCrqtOsYdKz5FxNSc29E0WjAUwExeHJ258IZ5eU+Lz055p8fKYFV
BBSPqCEHpSXW0iP1qsLIvP+3R2utDkUKHFtJINdZ9GaNLNKe35YS+18vKcHDzwWY
yjs6t4zfqxIRtr0uXfFUUaBLB39oiOENH0fBGVvm4dPWVLdnxt2BKdNsMoSNiJt6
qEQJjf2G+xUtBoaEnH5Q9bLY/1M48yWf1KUvLL5AqPv7/VwVmXI/iIWN4kEkh+z/
ojmy+ObxgTgYoOq77H8iorLV08sCXFTqTGwUtTpNCcx6FitIec1zyqZKK/gjhpmI
DCY+5lmQ/i3t2oIoky0EyHaP39gAFbRDpEqNLPaAp7Gf5fSJIVsGq7UD3iRKGUiG
ySn6A48uydg2DRLvwXgviEMaoCtlouiODRYOQY38AP5hkjGSufAkXh+cbh3IiXcM
efxuqDRkO/b82//TO/m5NcxPy6lDJQZagetFxvV8Fy8roxEaQcCuE+Q2S/hxbVaS
OXs8Y8Jyzo6BUdUeyCRQv/3hmgEgDiKTqOgpNTq0rvYKempa+eaUk6T1UZmGKnXC
XMC/XR7ugmXfS7zwaXipoUoBlR2ifsidqKAIBYOME72ejFY66EtT/vIf52YNdQlZ
9zD5+uc0VssZqTGZ9+98jzjcA+LWsGIuCSIfaDijyhumsUjBmz24Hq+GWX3T9bB4
kXiUgAHKzpod1/k+Tp1cHpB5pU70R+mtFNHDDuQ9Zay/NDe1RoYImrz5XbWACMdd
9e/7tqhk1B2fhMAIbq/VKcJfWB9qYCsvdUu8wp4ABeXxGWzcFGiv7BuWcslTZmJJ
SX5AyTeWvJky4oI9afXPEez7HIFwWX9Ia7BehHX1jkefghYEjrxEKBpanlG0ehbz
TPub2YT/J5OUgo2/KGBH7/gtX36s+ZTHqjqczsFkET4v/tSyOPrHGGup3VrCYyI8
rxFQOxka2wd93P1bdEKktuwyiKx0CwEFZBqvOWv+aNbKqhyAzejFIQjRHTnEMnFN
IqMIHBFZ7c3bShe/q0Y3lIsbTrm3odyhYhqS+QtFf4b8FnCqG7Ps+KOXTESn/S2G
LAYXb8Nun0KH4YwPevAUqS4nUJFxQAEEmg+vrCWX5kHGItBD6lv7SnBwDrwoK1wg
NvLaUpfD4a55B1VcU9hvjfSkEc6Ew36jm4UghHHe2YKS+hP+UnkQlcJeMZdm80mh
sKDoHRViBiL2uI5I5sMYV4ez94B3GcYZMP62siIwMab4u23ItCiA9U5PYyQ+RP6j
F032ar0MnuodTXmXgCKNc9QAll34bZDjA0DSlGcSYK5fkaSiXdFmpEBXPifO7B5j
XCnErqNVW1qjPJcYdNJtNmkIel/xbajPBm/SZY9V6CeM/2JMnhnwYM7dyFAkwjsZ
t3eo2PDJVFntZR2zQjruvwHkL1Hfh1VzwiMgr54UsxmU740P2v4Zrt9siRvpOOYX
gElxpWmiYdrS9R0hCwqfONWp4QT5Tfips/rfnyIVqckebCsHp30o6TR/TDGdikx2
FvD1GsCEhAuSQTT3SlDWRB2a9Ku81qJs4C6Dy7Bip7CgA4b7d/Wx9GgSywtOTrpS
5AbaJjKfRDx5nWBOFdOgv2VPz0ESR6exMsxh8QLjdimnATkkB2omfgsNhaIvp/oQ
9F9aAoel0gvxXVRRI/A/cmctPgiasI1MNrGR8YZCUaAWcGj6+Kc3yVkl978wzRmy
KYDB9JUYgVQmaFot4wg0mzt+v//YEhAoANuPa7mH5CXqzyOLQxjVTmSbW3VRRWHp
s5lJWcJa6msOGo9Oxqz+Mm97IXRJl49RgnM8CjcBjFN5juznQd01S5lsBvBhHO8B
IRFQVzJqyfQcCWWQFYuCDKu+xDOCxgh++Suz+188auFrDGH46IUhhxVlrdAhQK+a
KNlQxSV9F5C1sLBIUgpaSXYYH7XWwSb9UF1m2yjlFj2/mbU3aI/k9B5BKEhtOTCE
4cNOmGpih5KXJc1qAI6KC6FdTpETQxtsslypus/Rm2s7wOAbs60U2uEmHPrG9xA5
SZGiLXvqvoSCb0w85XzFrbBD/LkUndxxqdvQ+S0lehnnVrldoTZO1tK/8EVwKd5a
H+TIC5409kb8Cw4Sd80mdU8GNQFoMVGcRs2q23phlF8W2mO8+dd9hzj4Cp5XGCVy
EXyZt6YSLbQLNDJST3LzIRmmHzblUn+QhRdX2SjsVUOtpJnLEQGyx0VB43Ao9+oc
Lx/cmq54C8HjaIrMeaIXDJZWPg/1qQn5NCmsndVkFlxhEdedjrrOfQuaRkez3amA
pdGuF04TCqsAkCBcLa8Shuv5CfiH6J/CU3avORU7X3qn9EaKSu3mzs8D8wLKsJYk
HBWEDFF9uU4ifBubSivYTudFjJXygka3TI1qJykEdGmdbISH+3Z5e049Zeugftda
n8JRCEWiXKUzllhKhm+q2nOH8D3U8803cj9D6UZp4KO0/MY8sTqKsBOmS/iPhdxY
md62vjS+uYpktbSA5Wvim/nA2hk3aSIuV5ao97T6urzpd6Fh2GLpZNk2sBdTkppl
bNz4hAf7sa4Tr2UMxhIDr7l0kzGMppZ/8q7fmPDvxFpUkzdmyclKkcS3/esiPXCO
yUsSmgzMb1i8ZjsX7MvHzbDvoC/QOUfR8TTPFNdvo/8Sk8dEADvjpR/vkHWZR641
ga315jstBSWvEUmAnebPHicjKyuG36UAmNtl5yuEEOXvHKHpk+g3wQfp2F++JiP0
LaCvFWexhTmjGfrZcJJ/tglxDkbomlZxSjtCCfgvKP2NzsaotjoFq4hgMB1Z7INX
bNKh6OsFqfV3bTtUVwQLaxeXtXXM5eFWuYqOo9u265w0wFn9nZXuGy80ksAZ83I+
JC8JCyfKrwWMCKIO4gUIBeoNGz6h3m1ZvMhwIE0QXL7UYB3xm1lvQTrDlC/BJIMW
ud7yxm3eDU1Rk3G447M2orh+Pr+gZ10Y/LRuFn62iTIZ0QuwEL3ZHaZJkx7c8ZaY
BIvJwmQofCM4JLf+ocYplFuXKbTpAf9TFUK/JEjU+l9aP2h3MWfyPBiSGjQi8xtO
KarWCF+L2+nVHx+ajkDq+DzOudVXHNAmVZ860IQ04F7rwiPhyE4z4HF7uy8pQSjz
pUis/qHU58HnaTehvHuY5wpZbVL4xjBfVkNYEnpUC3WIcxeUSfnMoTzB7lfl4rBp
9INB10YMXisJGLcqbA4y9lFQU6D9CWn/enh9Q0tcC6m84iqeHqU7CtuZyjWEiGHC
7sPMyAJkVhHIGS5db/vv/GicwN+14afsfSo5/grWKBjs9d0vUz1loCTQrHwvjkxw
9NY2UIqDHQW4w8J6O42wwBj/gGlAw/X/gjuh7cIDYhxTU+RQWFwtRI2II5RMzw4/
xamMv1pb0SJUUUd8ceOj8FyTtvCKr8RpfwezwyJOawLSB5BT1+0cIynBmAu7e+cP
C2hInLq8WQPkL9AKO8Wxr939aLaiXvi8pFzJmPdj4QVJUev8C76hdramg1wClYfi
bOXMXZE3vpDxoDELRNN5T3S+03D2U5HkXm26M/zC6UqPjWszk6BEnxh82Nvnuw1R
ExOMzwVp4ziFrvcPDhJxBoVL52klQ6YTi4c596Zubiizii1Ws+0pkg9qVfEAhrIY
fbrRc9Chk8lN9TyBCUa6ZhfWa7W2Fm8q6jK6IGpFj01b63BS2cRzXxeJmqwCdn89
guFJ5wKrNKRbavUixJjjvwY7Jy7LiCf0odrh+iizbcN8VfzS9GxwLVMmNzxxxfrP
qcjpmKQHUS9rRqj4SIk3ZgpmIZ9dhbisshP4TjXHFFQpSijjkBKvZsa3Ej+kDaTB
2kxXCB6Pbs8N1F87v3W5HZc8sNM2Or78fDg056ji5es/jb0GswwH//qBXsKTNf/h
43U3HYoQVsN2niG74dVUr4I+R3hA7GmbC8lX4kuTFCMcoVMKp2uhDDbTdLrEdIby
t2EPFDL87oi6OKiNH5JSDOXpMabrx5bBhVaL8P1zV2rZhQ9dNngC2yGIzywkYj5R
IuT9QopOAc/E9z3J0zORjGgjgxz4S72xvZYAARu+wcMalWRVPUD3fw0xlLZPPNUN
NOYXmGrEWJ468Jk4dd4GuIIqlYhTjsIP9lvIrz4jKgdTvVtTP54DfEQqqaqOi+nh
CTlPOVhita6l0EIkGYMbWzuWPZ7byfnKpBVYRjWLzY6Aq5vz1GqUOlLavD4kwUpA
Nu0Nlzso5ilzZQdMSCXIpHzmY5P5azZgSX2dLE8JrkVVkW4HHHkEbvVoWXCxxm7S
D2F9GDvH2p+q1/SiT/CR59pafKbL8jyu6q4k73eD2jceqolRzPzTYiMag76VM8j1
EqFp9fKOvAAvxTeRtaMIepqbxbU0F+86sLIyMOmsk4rpeGfGLjXfXedUCGZkGJRy
XRtOb37TmzfLBtUThuVBAi0uJ6dRFOKYm/2MDVQSGm4/A9zS0bMUMT/Ynww8DAXD
cjrJGNfpBaHisIb+Bg110VCeRt5Zooznb9cR4G8XxXzIAf6jSjCuI4m47ed4Kp4i
hLsVvVNF5gSybX/1UwLqZU/v4UuGgpEjB2ssZmfFtkvC5SCNvfpSJgIGnGkoeC4i
9ZLJZ6DQnnIV/8cz3PHpeMDeCfb+3/TUKWdz9X8NEwanVFXAwxU4akoS2k+NF8G7
qxJ2suFCwPhXf2zIdchz0stACI3vbgn69fMDjy6d3sNlfgDhWe6SvZbb0X5X93uv
5nT7DXt3Dp/L/0voyMuoLGxe9LdY4eKLqZQ+0jQ1YCcff7vYB8f+h4NThl0AxAQr
uqIZZgtIA1LGEUFYxiGZ4oe5uVI5/hMpGjeb9qEKe1KWi2DeH4QbsKZuCBrEk+Eh
8z6WZvCTUQb5GnaQYp/fJLlU412u/iFZ24nGmB9/vgQnBYCIx3USta3xXBKr71Zn
VS5NnacxJhKcPVg9aWAU2zFeq8079S2hdaIefjKVFy3HF0kfBDCXL1KNGyliFpbm
IhJ+w0dEStQGzThpSvG7EYrGI/AuDIM30LR9QJW83kBwRNDsA2xfiGRFG5oWWffu
QPjjBKavSecFezWkwfuVWLxRONI9tzyp99saDQKsg66G4+TnkdpH9MGE68eMyhZ7
bRAQU/E7CmevOMKKoqV/8dk7z8n/KcM4LOkxW7Y5PdKUH2q4JPOeZ4NA72U2r39e
Okw5Bia9svi8RbuyIVOphNf2+tHCxfQF6avg/vFIy6Zra3nOV3YjdrHROxkrIh7E
dAbi0WHU/g7pW+Zcrqa9xv9QC8g2Jse8hA/XhS/JlHS+nhBROLLzy1InQj1kkoDj
VHPsPG4OBLy6S8ga8AOONZzdSZE2pVl0a35cDxURJZqxZVr9v9TqID54ebXESEwg
SCvtZOiRIix0xVXf+o2HzXtmSyQuFg9BYoiTlqJKKCTbbKnUY5IvVMHChXzxhYF9
jClRjfpP1SaepbP1foPc3M+9JjsiXofrR/lSD7hPTb8Dw+xE468kJFaXiQ1U0YgY
iGgq9973nPupdSqKHmpSjM2DsQ8wLKGgw2M5fjrZy/9bdN2xt5cyhGZFkvIXFU7a
NPFS3J+pQpKOLZEa6S+Cf2mec0ezKpvxDv8AVZcj+3kRTeENKbZyPb2/Gldkv55m
dBoCo677vkvu73lBPzVi9xrEDRauADOIxSEsSCVMgkAvy8GIIMjlOPjC6bopT7B1
u3TSP5FNwSM5gJzY6VaCw8/ZeN+xGk37PamNtl1S5po7mq/R4Z7BtKD8bimQQkNM
sb+w6RGcuUuECab0Ly62osjUPV4m/9Jquhrw9n5Ok2cLQheiI0Iwl7+BGuj6jPDq
NspZ0APWN3XqMnA6knPjolfYPtFqmVIYGEDJUm+HDQFSG5nsFXl1b//+XwcDOInI
rIKstVnXqC6KPLmEgvtZcWsv7ZZo3etsZqxNOx4jBTwZaCGZs8fiGZqm0W2m7EQs
xqaV0BytHdlrYyqGeARWpR0gNl2BmDWmNz/UPK4xlV5JbC4yDmRu9hfwoBm4DQAh
Q7U6F4uz00tHz76a0pquDUup4VlCTtGliZjMiOLiP6GvUibcHUVpLSIbq/v7OQWX
SFvoMMhjsscpd4cNFmvqjRrOvI2Diit9gfHSQ5ICZedQWiJNGosoRC84++/GIKvB
vbhuSRqW9QrP9+/jAjL31pg5jSH0/D+iXr1/6aMA+IsoLtgifmrmTg3frl+8tV1l
0mW9u12T7hU1ICAP9Z4MlWTLiJk4GKcZCjza5MDWqtWodnyGSQkNzF70Rh5YPKQ7
HNiSYExdSjoxyyogMSptcToH1FqLRPaAUfSpIUAjGb2EVYGYSJkH/Uyf59U/busr
9vIK5kK0ise5qmauHEDJroD4Iu095q5bXv1XBG3plR02W6A4P8cDnOsGAjV3xhRq
gGe3lJoqjc4djYsfiw7LnBAr1lbVa1spVotYsGQXwjISmlDY73BCajkjz3Wa+vQE
E6y3HN0ohbYl9jf/RrLJcN/tyXRrCYTTEIEmOib4tIkY3Cs9N0YE7qd4JMolylAj
bxSOEz+NpFu8us2pTeDdMYsTGnYXZ4mwxaFyCvq0YsfAhPCiBxODTa2ZRr0LJ6g/
TVc1qrERCxsDpuQnwKuotl5aoIHY1Staa3LZ7ZGmuB4tzRjmA9liP3YOmiraJdA6
Vkp+4IF7HwqKFOUTvDxCRROLx8PIbFRVew0IOnRkyrN40abMfqWQloZzNa1VLTBU
DZQ1a7CRdPde991bX3Kwt+vNxoB7dQ1WCMj9xG3pfiGKGb5A2dqiJd4uDulMTZ7P
FNtaDZ/f8EKudD9dI/J3PYCEFj/M+Az47uO7wVkfvJuWh3rcTyCD8K8CR6DG5PrC
jGEYA3kbZ/r0qtTm/vvr4Kvr0IJkG84uZRnFMSwwVBo3tNvoqoK9NXmI0DW0r1pQ
AHhMXWUM9sgULZXPfrqAXHp9EuxgN/Ie7BjlQQUKkt2iiMxj4TML8ockuWEBkdl/
z8+g/hl5KYj1HbATxFyciMjWPaZKFGv/hMopL/fsevXRjvUwo5MltItQETpc1EI+
NYZazbvont1B8/qf3rR/Tq2e6ttrem0q+JeVJZq1efRwjEJbO0TMkt36j0oEICP+
aKwH7Kc446vJbHrf8kO7uAqvEj+Qzl31Jb1Bh+PxIYx0D0TiY6NJkCr3ZLd8D5CR
ZZCqkV736qgj54CvfEfopoFw+fP1vLQ7h9LAVFLKcALnBYE4n2OQh6BHZc+C75Ou
ipyiYG/lQpfRVh7VWt9AyMRJueuNeIpFkv1ubhDszK0d4vNhgo9dLJR9sC8ryjMZ
X/UiMay7GRG12UpLFrWdxQziwHCNq7tc/vbB0HQHsoIBILEbihRiQMTSLEpAsyjU
zFFFC3YzWLO35JxycnTwv2HlOk+Mx7QgfoX5r6k2JrP/uq7lwC3mKmdybe+XwEJw
BeKlWLt3bT4enjIfEpj35CI7utWipJNdGoRPXoxPDL6N8PJRQib1d+UssB8w8Y/W
Wjb84cu7R/fAAMec9V68Q6bjbcBGLSH5hPBkgkK1BDD8GqxB2EnBRKvrJ1a70C6T
GBmif9hNRvnNXOyJpA/INVALK91rTRnbAodiujvAYN5MuAiEhM5kasXjQXCs1HY1
xl9M/EsR/XO+qhiCzVZgxETwfvzRTVlU3bHuwplFhUE9dMt/T8eCN4bJLstvuV2y
QUxESdCFilbHXu1ZomKpSFl9ulPz7UoQPRFX7zozTq1X5cvlfHnOA9n2rnXV4APG
rqtN9CyjucNk4nqmRB6iwaL+y/+Sqk3ZSK/5NUTagdSKGoMDWpZyfVdiuFLPId3C
b5cKnwB9iErDH8N0amLoQA8t6BQcaCiZxEAqG4GarTMd5zJr72k6i+mwULHESkff
ILZR2Sv2/HZ/e5RD7Va1oLIbUZzQNpdHlysSrgD2QZJpJY5YKSVZMzhQvw2FYYE3
PPno6HdjWekAqpMzG4vtdwZsl6sTUvVUE8atT7FwK/iCqZWrU9XP94WiF5B6WIus
LL+EtwETxYdibSG+DN4eHg6rNSSjKkRguH00u4EtDuv6McMSnPvYAwvp63ct1lrG
n7fLi1hntUfczYMF37SPd/ewS4F45B6caqPGz42FkzPlsWSR1qn+D+hFHf95wylN
hJja+JIlLoqjv94tABD/uQG/taTtgNxdDOMMs7Reas1VSwI1062U/NFRRCvC4GOp
zccKqI8jR8WvlkkxdCj5mtbTkcs/2nnnjqg8KtG6z9vdAmUT9KrQN1DTBoBYLml+
Bw5wOJGbKrjSgKGCUn0CIxOTKk1aVqVESg7QE/TtNiWcEub42u6ez5fjfenfO93p
rbhMJlGN651xvUaYb/l1ML9LThUIUgKzO5sAQUU62g4LukUIS/4B95EnlJCz5IO9
vCjNmPU1NzvE8WGLMR3Tke7TC4JixVX7omjbHpj6diX6Sd5OPQac4kUwLoCK6bvT
QXnflY2oc3xWAdWw0CE5cpFf6jWaY5VYDF391oERd7+LS2AUnjLpC9FMvMpXaqRl
DND7i9vPavJb/I/QswV1d+bajpS92IAKIHcu8RcXPogvKuAQWwfZrEhsVp3iPMOB
xJH5AB0xZ8sugZDfbQQ9g9uycIwlcgsKxDBlhsyjtxZn+rVtuMkx8yZh5bLq/nOu
gKZnjntkO5NxdE7sCmcOAaORmyPMAyw30kMjySWei6zCpiaKJzioVRHnQGgs4JRL
AOltTT5uY172IWT73Wl3ECdnwwQJZACp39VBs3kmtbDr2WJNy4T0T+jEirWCu6gP
k1A12D0p+TREB9uywKvceKVzTv3P+z+A4QTv4RyM6kzfM0b+ayQfWwMMcLMSmSBm
Hi6eBPZ3mRgXFkD2fXtTrIlCR2otwN9KT0QAYNiORNhla0ZkxNkMFE911e2XJ1JR
rKNxff5nc50IykbUUMfK4GklJmYVTooJpxPG8JMlXKdCZg5CvBFIoB8dU7ZY5oz3
2QgaTHxB2T/E1hMnQmVCAU8tcxxPNTRHTQ2qbhTegpTqQGwzqU61a1bO52bBWTcF
Aula5A+2k2GD6+7AfuIS1hOG1iM+NGvrW7NjmVhEELeqTiLMsgkDIknOuVzmhZfh
oBImqig3ANrslte3IXJbMtNDK5vIeGTXDnsM1HafozovSC4UU6gM2H6r4Q+gS3Ci
Klrp6xTtLaFLoSIzkaKqadsb9f+ixTvFNOx9n29jvU+Sl+I80LmoeeDMOL1W9LAH
dSo37V7QEDVVep7B9CQLTeTQY7N/lTKdNOQAQX7tddzmY4J4J5+SZ3wbm1PNmcJU
jrI4AuQgDlLh3DOPsCDZTFoGA3T3Pl0Q8scOWZQCCPT4m/nsLu6h1N4hQxebhQuy
mN+BgyN213QNcbNAMpzyR8i/7lqSu9Al8VxQolSrOGEDzZv3qZQsxLLd1qsRLPYe
kZyBLB4OWI56KuyJ4tUr5OSMHcL3zVQxDjqNdH+58DvzAyrUwlJsZwANsvmEiFKA
/nOdgcpLOAkpeoYhjmjTdHWEduRfRqFdlt2UQxRqdo/r2i9pgVVTAxgRqQFnFENp
26a6RkfzqNjyA/XUJA6806tmn3ZPZt8d/PM6TuOndfNkHsX5VYjwVYLTUZUQcEBk
ifus8xHhnnFZLbUodyUnyCntLfOCgO0ARWYLlsfmn9Ymu6G8mUiSHiaCiahLYzAG
xyoWbdQ5+gGjqknAsKVmkhAI1xvfcNjAxP4pBVne7geDhI1edfAdZJ4Ty5E7vq10
UtyU6aL/hn5UhIj+ASVJfYs6bGZVwCo1GZCf+bUXVwCWCUkI7ZXdCzBMqauxxoKA
pmNOvmprD4lLO6/QjFUjOH1Xp5ARI83hreXAD8GjFPe0ycek85iCB8FGr0uYgFfP
jUe3W3exdtjPAGu4SGMH5/cG9jMFWttI3bIULrWkBtAus8MWKmsjYU6MdPNKMVX/
Ea22Nu/zAnq05FFZhO8+qzv0s4ojqGMM2l+Iologn9vdxO2fbY5kDjdG0pHDu3ap
sR/5S465qM8GJjzlZLgP7cNt7Su74O7mpdLiziajQK3Ft4SUGB9gHL8xLBuGaN1N
lmCjlmjJ69nqVWdXNVgKpjHofvLbBQ5ySbvejkedxetIJV6fRT2wascVdqFTBrZ3
KDJWRBidJ7uvJ82GB78HIDCC1VOQfY81l868y4OQYUkpgpRH3PdbagYmVgbdFucI
1A/2jaULJRbE1u6vQx49fbDB5wk8iFUSVCtZZoZ+LocOKGNQ72ot384ULLOLHsLX
b8kP6Z4Ntqa6IqG9zaZF/SRDC5qbXfaAGTzUUHIcSyFzfr05FT2APCO98SciN4XZ
rYjkdPy/7l6IfpAYrOGvLdxfiVC2zqlJCMzbSY/z9O+amh40QHpsWo2h1Oh0qAXe
6xMgNmLTgWkjbDIoLY1B2QKZa8TIknkwNGAVbS9pf4XkuNK/b5IXEaIzXe4Izm/x
9HGnpS0BWaKB0JNnh1D7WO6nky2MY0vCf08vJgaj77yAFqP4Q5NGWCNHzwwzBisl
pQPNvsdQs4waQ92eQvXFa1ibM0Zk2/qlG13RFvBH/bTMQ0qVqQHyBfNkW/8+Dj1k
b0iAZvIITnPEiYxQZl9nSE5ZyUpx/Vcl+WJPXUpMh2Zw65Kt7HGlFb+C7T4gfuJh
by+uqoxjr7r0QfMBRzhkHUek/lQXnI2w4TmAt2NCR5AJsoaEiDnwQzlKCMbqrvXe
LB/hk6/Va5w7zfor/vGH60f9PDbIJ/Eit3m0Q1DCqqpgY1kfqDETjtFf0OqJvS0k
gt4CWFFTANJtk9u2m1xdNRpsT1I0jdNeXXVswoD+ihKpdLDzL0rfKIVOPVDUT+Zw
rGupveMWt6W888mf67J3MwN3ywKa8C32desK68AWRhq1uwF8Zrs9w+rDLfeLYb6g
PVuSwGtlNkHdR31bMvsvwDPWh7VU1JW/5HOP4M8btk7zfho6qBuKBFfxz20fs+2L
XMd8SL3N3k4K97BeDSGi6OWjCoRBL3CBJYtwSCJrKX9FCU1XZyaGi9EdfZGNtbnB
Z031g93SkVK6HAnUgOOB34SXdOf/BCAIbO4MACLK8qW2ixNdd2pcGkAWXkz74bqV
poIutCB+rsNekK8TJjdhdLSqi0woltiwM04VPlvjFpIGC/1mCsrGZn4zBW1QQF36
J6HNA4HSA+keHWtE3vYnV9y42uX9/VFT8CH8AJiubFYsVZ5ga7VIKDFaeybNFl1Y
FMTY1KE+z3c7HNGcrPBFl8eh1ABJQEkLRDknIzrkth8GL4xBs7nGad7ULSdBrwSh
FA+YNvuKESASA9KTHNxZr8Xagi2FDW1qWq+tz56fGLB5r3rVhge7Lgn8DvZ7bJgI
oNZRmvZydyml7cjkZamfo9CiQZ2UBTx4JaALt3yjzYzJOqq3vukNwMdGh0gVMGbh
jM7xvUtafA9a+PgkXboKUfcMh1A2+vMR0MYkUEiT6Ihgq/9XiAefohRu6aV3Q3O9
VnTuMlOkZJ/A2FCzrDHAfNhJlGX8/9pxAhDznZv5HXInzL66QybVoeVAbJDMSS4u
AlFP+sEYLl8bZsUK1Gn1juqg0hP2erph4Zivc8Faf4IfebGAI2BA3u8G6GgR/enl
fE+/ik6K0bID8rJHflF/UYKPBfi2r1N+2/sOD+bFyq1gw3s42ji5UI17prfeZYcc
Se2zhOiH+dy1R5aOJdR9UrZjCqQhMDt5NWT34I5R1YBUe7je08CdHOuSZt8iAeDz
yreVFlAikm3xVYtm/eaEFeo+lqsJjc88LDqD6Sef6AiSR0vs6wze+zzXBXvCDqmN
TZ83spfqbB150l1kPHTlbQjziFl9oARhP+2NQ+6QmSxGcW7+Rb4zNzDOLuxsrygT
Ky2EgtS7uUuJSDeTrt3RcHuvUHkb7kJVy91cvkIN5tHczCFv7TbePSr4tmZ7TbKR
lVjIHUVeLhcVAB0c631gC/GRLJI+5jv8YKoi2vuSUdWhFRSAonMqf+weT9Z38ab7
pLjUNQx+OIoFiR8HP2c+rN3c4Kzkr1jTILbWfeXZI8S7Ym44ms1YdyTo5MPT+4x/
vSoLXpImmWpacvlNdpGo4sEuuUTDpT0G7FZDn8BIBoojvQIRnZM/ArfG3ZxKu3hZ
UaWTtMMzrrerhBJoxFnoVbC1dyhB3RFNWBWi7A/cloKkiQDvptdEb4u+DfHSRQbi
gFdHAz9SI73j4uOPntpvOV/pxg+fUtaXM0dx4afv7klzZIRgKIOVKVmO6wMgxDS3
DuM0SgggjwXf/OvqlFBIWhlAxmZUjWRnQ0r7PlzIoS4K7uSEopeHFipooTK4vvTI
PqCWLZqTog+vt6PyCP3B5VTj3TQBK9QZarOVPd+I5zzlyPJ06PHlCmGJx1IklI8O
ONAFA7hfPisQOG0o0PhUSybz6RTJCgCbK3h8BEAldsOTynARfmPjpTiGC4g4fvVS
oW8Hp170zihDvQOBDm3pjoll8lYqMdOBdAGRQbGD7jXKHrL9O61MsbgL6BPyb5fv
Xbec4oao+vPBZhiOZR4ZJvv3W7ArDs66KAp/ey9wAeFKRVKhNsigaHhI50xsMi6U
Ooqbfm7Uof9GpdSyXoNigVcH09+XJfgfJGcFWnmo61BpdwqszNx7T3PYJBRxaAZE
sYplNK+DvCL1ORqcr5Rp3HH3I7jtNfyaPtws9lcyx9Vt0gpzdKN+fzjiiuIS5ekP
Pnd3q20MVzLvkXYaoJglS0I+1ZbiQIUA9ebyLfvPGZoilx42ygZu4KTQaAtB+2Oa
gW4OOw3IQVfTj8alTV8+2UuXHjRvW3fg02Ar6d/E/GFiC9qw0D6v/WoXIttnzBY0
z2x5GnvuDdWr7Zxrdk8xnaZD/yRnTpxfTK7gu5s1b5QrH50B+fIU1XM8mlbd4Djs
Nj4ysQgAfSqwZbm3/XKy6S3jPnoRR6YagZBVy7PJnpqguodkkfOdYmanKtxuFoVL
+Vdp9XnDeFh2NWoJ6odecu9m9cyzQ7rcrPomBBHZ0MhWCRrMj0qqr6asIqtrD4sR
AFO1lsWfRrecMxjCLtWlVyp+EDbppv0zTZpCs7hLSmg1LKa3sgEQ4zDUHl/ateKq
EBK2iMnPbz0Crn+cmKKKnASBCXMERLmhKLi12/1gS2qHjRq8z4UVpGsrPXLaubMZ
bl3fSpn3wdklrvtgVhFJxDDQChsApwoApzCtZ/QEn4Ql5+odyuZuun1QumZ4sLgh
PkmIsDRdg3v0n0tWdH5JrKQOPfsI5PFlrNHwTt9MYOjK+a6OzFSpcJxk3SOV0IjM
rL9ygGe4QUftKTE0FQaqh+IWbwXvet6ljB06byUgv88dPllxbHPesE60JtM2dRLY
v9AUrJJ/MUrswM54lY0RKRiZwVrTTRUFX5WSAbQxWhbOlHDEXw4um9HRJI5u4+zV
OdXc3KQ2ZHMEP6Jpdg5uKVoeB2IpyZPPnzgE/W971TsGB/zwmSgPNLs1FPCSq0m0
2CXxDCUMHFyp3ih3+EbS5hPChZrZSaMDNpZPqM1A71oS1/M4AY1jT7HfYwK4IE9a
qpv8sQoSaXMlAI0XbwtT0rVU61ec1azgY8/DxpwRKkbk9eLnaSyvwfOXOFqQAKc4
bSs6WgtlrKVGNl2EiyGcGUomlmU01uytvvie+38Q/n8nAcW5xj5UXixiK3Nj7qTX
ppWeB2NjO4a6K20v3drDT80gd9vmBkO0w94XWNZXNcV40dMGzuaeJmdAguPtrYCy
dUina7BMy4m0TqBxi2HFmR8fMzu/ynSP0i9F7AriVRM1rh4B3RWV5Ty+LdPWKsQ/
5EVr4Uv3eRGjnoIahgkvkkvmKm3jTVXLHoLktoMp8P8qeZhB/dJ1iC63nBESRlwQ
YM+vVBL+ZdQsAGSyJv92medmoSuX4AhNF3NND+3en6CBqi0SpEla+2S7WY0EIvaz
QbKuWf1csAfaEvF7sCczUpljOvtVilBCkvX7wo5GB3xUDB4N+VOecJ/yad1wj0Ai
VLssOQz7YqKLVbBjdwE+WAm+ggOaTeYZX0uTaLqDN01q47narbnpvNJCxC8Mnvco
G3mwdYtrXsPwB9jKDq1HggoktXrt2/62mYnSNGA5aw79qaRjg5z/3Xd6d8sVQxK0
7z3KfeK8CjWfbxLItEG8Vs0XgVbHw4sbeIcsQZHE+8VnXg0ACSklK9xZZlhmg6Pc
+ls1Lp2rlF2YxydVteGjEfGlUAVYLkbdYfjfYbC/r5GBYg0QXkVgJbs0V/zP5KlU
vYyG7ZiPHQsU/+8IyZ9xvww0SqKcxz8HYGbGTrsG4B0nsL971Xys2aDs6bZLWZV1
R+YnsJoKWyW7Hk6JPz2xHXrnWwbgmKhyWml5qd69Rvo03EywIeay37Icuz2vW+et
xBln3VzEwsG2WYJttcZLRu9OovLRRP1CohsWcB2fUOZvyEaCQzREOaReZCxMVIMm
GdkfW7LJmgriW8p00Jdg7S9Z2+WVOSdZ4B2qVP4C2YEQtHuwmevZ0SuF820H6yfX
CrWIKbQnn13lw5ZqQKRSjw/UmdReQlSZxSGRt1O6hRy/GugLmB9iIppSTVDLMMvp
7pEe/YnIECiEkFaZf+SLbBk4rUd1ZwAfm0dH2GhfZB52/deniCjI6Rca7hMGxwkf
tJpZRgVUy12y134gNOaB8lmP2MGEloW1FXt+BZGb5OvT67bUlMu+wbWaRdwibCjt
BZr5rOWQDyWtjVd1HVEYRnypRyOfmIBE5BcCa5xi2XSuAJiglbqUXCNV3p9Du2Oy
/Sf5wGcSn6p6+UIu8Azzshu619ZLFr2+LZyPsL/Nm5F6fE+WItutYo7jrlPd67Wl
ZKwow2aa6zoUnzSfDele8uBE1ZapH+ud0y8OB79uZYl5ifHlmMdJ3KX3JU+iCOFM
amxoE9WRjEI/XBtcgR+NsFt7pG6Z8EaJub0rjYnQlLD5n6Yx+3au1YgpfE2G19Dr
rk5qsV30/jN4X5b9fFt3arO1/JDqZbNQgIMGxUJy4l8iRroVLbg+at0l57QxZmrv
O9/mDo/XiH3BZQf7jza/Ale4lMJ200p/DOe6GS43NJgaP60+1YZAycuL/RCpi2GG
+x+cX7DsKdwJdMR4QfxHPW+iCxUYQd6rSSkFuiaKk50mfP2+WmIRjl9svNoJjn6u
qYqaPXBAM9EXghZmmB+M9RaXkvcviWHJLTNnZYVZ4lICW54msPh1cIKDdx7tzHM+
Mz1lSQhIBv9b+UA715keVTBVbqdak5CeCWHRW1jyEM/Bm+XLDdDRUOm0gEDeIPsT
eJfT/+wMSRs1DT170+C7SgCKRHtkbmFjnMTFmDxy1dJJByiGrwkgnlU+0WGxRFxu
lBk4wB53JzuBMZPAddRLysVgQwVcverYi7oBzQb4HZmp8sXd3X9QkbP5bVqzExZp
q4felUD6ZiYhkzG8QaW53DE6oXSF8fosNW2xQ6Rh3WktDaaQZ7hfPM5FTGCdJJny
WSSkrpEKm8UYi3/EESX9E4nTmfG9PzrXVpzm2MN2+j13G9hzKX0AuQLoHkRVDI8Y
fAr8dVdGzGPM3pZDE5ypOPhBsZzrqOBofhSKXbWdpYA/QAWs1RwYCCCDW4w4pO+w
vpCVwcnTPzo9q66wlblZjtIoi3XfTe0dcHwXJt27uvJZ/53XgPLh9YP702+D8oXO
9GEKdtVZXZNwaK47/+Q82+tyP8ScXb1zEDjJGe+UqRqlf5xmK4QBq2cikKEye172
GlPVBwbHACt2OGiOgQVRnScp7MsqJDQMiNmjfJ8mah6WQ+QXgbW+EAauMOsYSVzV
cZ0T3GGgESK3kR+LVkitG1kSiJdI/4uGWB6EUPwcCCu9g7q6qV3PrgaZ/ZYax1nW
A1TjS4+Bv01tVi17dJ+NgdCHUBb+pQBRaX2gq/AyQwNqOoBd/bhxe9Ftumyda9JZ
zhWaQE245wvrvEOqbEWtr/SO1tJ1CL3DN07OW9aN6peZ9v8Y288PHIuBUmkgLlW/
zsHPd4XmAwY17Q4VDpfJRUeboEWbaezwtdNuVw55qBrVTPFRRmkn6VOsKMLkG+Rw
0Qa2EwfEs8JHL4KBmjUDCg1qwrEDWGtCK+Gbge7OJ77wFyLWB5uxXKZY+yFuLyMS
inrjGkXL3ug2f11nBArwsqYtnUhREWlY0ebM4a8aRsejwg9hu/lMz9ThsYWtTez8
AemWjyGT42IbamWL324x1whXdkYQwk2ka9mKjoBwzs79zHfWtG4UPvbUPgR2cLEq
p/cqEkde2VdVV1pjdpdyyI+Yrwq8YeQDRvCoUy4RigSy5zQtDNNs3sea8WdRCub/
THc3OiSvynup4CT+EtBgIFgKW2XizdP/eJN3Jp3zIarmS4ixQ/6MaQHBJbd2Q46F
rhB43HhI1UN3oSZyDJRQ3VCpSavTXZZRvarBueK4E2oadSNttdu6LqIaPjGPur7F
GdI7IpI/xw2aBVZetvltQ3mGa6Uv38Dksie8NlE5dSZvUfikPHrdedjBI1ekMwKx
ic3PmCvH56p9bm5jN65/8UoBv6h+E6SvTptfPZ6E0X2iPuyJxfCPHCHib1eEXcQ7
tUV+xoifJKVZ3/wAEq5OQuYRCs2VQ08CYfbwBLldkKSIx5ThFAcW6UvWQ10K2azB
mpkRRhtdeqYIKco6Jm5E4ThopdfWYqjD/JWcFFxGm3BGfA5wfxwf/KzNJlW4ZKki
A/DLIrQn3gc56yVoPGIVfql2wRM0pfImskYXtluV3YvLj52DbjZq0SlmyjUmxnUt
3IhpbeqtBEpUcd1h0H3N5hIoJJxzrxzDUFckU0jSsSkHwvxPlUWZqAhYhqtQnMBk
yUbx16tJi/b3mKW7kpfw35D35n8JipTd0cKTNpVzD0/MjL1WPL+8A1J2d4Xj8L46
YVuWQFLBICCcqxxqjdd8QeE/w+AUka0zXQb/F60AVOlrJNALG+B8pmTH07qPYGQG
vG9v19GzstIGVuznxwhPS1WmVAh9ALkUNeLishjS9sOwoLNxliD8Sk1Gpyaj7oPs
8GvG3jNahTGs7Iacp4UgFNbrKNvlKUQPZkb3l5pd0BJ6UAuabED9H5OacY/H1HvU
mEdtgr2dXq6vEuH2DZ7+T+iRBLJwXxaoJmdOM/+qVtyzZDMrgYD7+3glcQTU30pI
TuN8LvNXbbQ0OcfCVTnLJCLp9/+a27dP8AT+VUUVvn18FCrpixsCdee44qNFFxzD
aDfqkMKIn0Oq+YkfppSWD2VrT1txV1aqyswOyub8yQVKqIfjHB57OQH2hZPNK3py
hHMhFvSIw6f4lBZO3tRDOs/Dao+itA+6vfzKtsaQl3B9U/UZwrJXygy0XcLKzPc8
NSN5c9iurZTMLaSb8ejXpaX9QsahSGLpSCI5ZD7xeJUFN+jSKZyaH6aEJhKjc4LJ
A1LzTqcRO3gS8lKuw3mwYMc+0dDhoH7YeWBe+bxzpS2YaApvUbdysqzXodzIBpRd
4Nhhy0QyYsAV6KWF3yRnJUka3KShIZIeNlRn6dlD/l98odKYSnSDMiiFgRc1ZjuB
13WizjLQ2qiahpYkVcvWJCzKNpE+GO+Ji8rQoWBItaC2euzoxDnOg1NtpW9buSCx
DWKDe9hmjRNgvwYqI2OnS9S85UmWmH4jeryEwvIbdO/MJCyIRn0m/baeEfB36idJ
q17sWmC2ony7MEAx1Oa+e/aIKTFuXKVTNykgBhM3bVMR/PQa7QIAAivj/I/sq9WI
XMKTNb6mdB2WOhdPNC9IwdKvePi1A09iycnWpbguI7SS22qC/9kDbf8RjHb3E1T1
CiwG/2c5xTkjd8QRu0x63xcfBTYiIFBROoHDhAbFzBFDINyXsIRlNA/f0vsiD/rq
ezSzRAnWmTG7bKBa34lSbmn0e+u5Qs26SRc8ZtnwQ/Xigi2FNk2AOZNcvkjnr0ig
R3T7wedM5zLEaAR9qKufxvGZQTwsIBLA+5svFVawQlQ28/NPIQHBzMzwg1QY2Bac
yl++Cm4wM2SAevGc106Js4NVNhzR7BKafm9yFitEpJWSs0A65vdvFER39R5iSpDT
xcB/DslOmjkqBM+PQUkgw0xu493kKYIYg07z0RKXL+cwEVRrOmlQDM0/ReQlxovk
Uj+JNufXIN99WnY22jx197wcJekvP0kPfjBsCX3QEG2ygZWSSoY2yE90D91VXFQH
u6r9y4zVr/eIJ6Yx22trUKmM96mI8IHNWqRFSQ7Z/OZsaEYUSQkIPr9sH5IwlnA7
gVUk21pKPYzPWNOMb1y19SvtcV1g79pR6nFFv1xK79swPVq0gTcrq4WcX1+QoK+s
V6YSfFruKAXgH3VRWUg4ah9EhtFfa62FRH3fC2U5JydIvNa+YKJEiFXeC7BejG/f
ou9pcKgzbwtKWKUc8Krxs3zCvl27qGf3Gg3Y0fRC6+Vk4R/H5eQLHfFI9uPAf9w2
qON5gVZIkevYJ2zKXqzWVUU247dYW4L4iO/YMiF7JI69NWExduzH1r3IsU27y3GB
cUd5uR7w3Dzagd9GgIiTFxiLnhp+DZbAK1xSYKliYSctTiUdwvFkLiIKFEq57MwS
bpUB/aLK9+Z1pfU83IHmVE44n7IwOexdoNkGqsBEZvePtCHSMtRq9yC9LUHn9gRs
mHtf97AwsyOU9UVfblfZR3LVQhxc/bJeb3ZlRnRk6X2DfzpuwEQpZEIYgcLwGfu7
NOEeZiFWOjasx3uKXNS1pMJZOlvJqx9WZwWZVqxLUBupqQ9cfkf9CUQzs/LLHdmA
r/qylma6pryzo3g/tAp6GmFWdFtKP78tZE+zhFCCIN5EJyybIbYBP39VUP3FbyQk
NPBP5Xqi+9yyC2kJRqfa5qZH7Gq7GQpjO1zNl1tcWpLUUChXoHqlosrAuUoPO8ZK
pcreY9PlIJ+LIhEKr9q/xyzYVsmQY4/qeGs1wXV382R4tgtAHaH/e68Hs5lYSUbG
cfChC5yWoFB1Ii5QDaPh6WKeb9deaLFYX8DZfzg7S7o3koJZeIqTpZciVFAUW0cO
8cz5YY/SiTFGf50tbHZcl0NshOczDX2i+BgD14qiMaKcYgx/2RPwP0XVuIaoTR1k
BqbvO4+LW4mXj1gmJA/OxZLcJv4p3fVRVm1uIH4k6Sn2QvpSgqwqhMfFJKEfxzoN
KF9OzMhTDpTfBD+R1A1fF5mxpznLmiFt3ob+/QboTqt9/sQtQry5vKc0Y0zSvx9P
7ervvAxPZuNfWoV7bQzZhu/G4yX+x10PM4h/sLs0xoNjpEfvxGxdeehtsIWKugVl
4T6PyVgOJ4FTuz0cr6Zfa3cwUbCokWMSW0iYWRCH42kxAM2gr4E0bUgevQg6iMio
E4a9WV5qxSbgvIkQQyzRHLd9xn427QYJucQz9FxSkCUflu5jQoVvVEqiiKEYcldO
Ccan0sCo2fJLWk89g0DIsJODRy/E93fAmgN3Coo6scrbHqoWcYsh6upsYiv18BR1
sMiw7ROHBp0ynpi3h3ZcJ6hDWO5yyyRawybtzGuAPew4emTyH4om0CAdvV+3o4jG
uNMtACwkhF2TDUqySEZbU+aQiqYylaI2J7XMr9zikNVa0CJCLlPMG3mC5CaRcSF4
ewMjsV2yljGjp5hKCb4hMtxsHyoE/0T4m1e9Ydyz4bs4UwEip0ALjcLweqj7LfK+
+S28XxWeKwketevl6LFK1rTalKxovsFt8ISsM6fQTFoqzrw+s4Df74SFNDwZzExw
PKx0lj4UCh+FqsFonUQ4uYdwbbbC8nwicvKFgCqx4dE+lJFLiaa44GeuyrDKTQJt
ywKWE0YGIQBklYs+yCIvSnJzq9Xg1mh8zM7yTdmmCSjXHO+TSLdcqMlPUpdW15C0
KGMUBDfv6aG/hVHOfkftgzY3w+g10vx2pqErplb+7NvJ8iZBWWMLZN8vKvhyHHOm
A3Wn+QHFktylElm9WQRF01EkMPsPoJiF7R5atg7Y69XavuPypxK4z3P5xt3qLsOc
ZrD/62wkMfkbNIhSvOpQ8uRT/fwEJxjg5GeePFlsnJ3QWX+weYWVhZjGLjguoG8v
QSiI34QM8wvyR+XL90ESQesRwBC2g8KVKAPA989AI8Uq4G7Oxsy6gHaDNqI9ENEg
T+aZUrkAoK7kCrvDEcaDu8/BDyFbaTB7qWD3rUrxMXjjM5gjNrrA2M1qDcJpemo2
f+/5mvIe6T5tPjmCEm4XNVYQDHq8Zbp2w3ZIxuMOWl42M/QgYbktEK8/1qj/Wu43
bcgmxsPvXu8mmaGoWp5PbPGTx3h3p/yihkWsG0aBKY9hEcA9cfckm5qqzTgrM4eJ
G+p90JLZyNjWTtnr6Kk8wyNslSH79jRaXNtuxv4eTF3ncqdq5stvbTN6D/dUI6L7
A3f6e4WKnfOO60rSNWUIYrA8nMFz4Kei89zGfi9b8+VqUQxKKec0m6fBJcBXc32j
kc0ll3q4BddxAwFCjsFu9kKyWRi7NlG3N0sDwfjVz4AJuFkC5ruH77fWkukGtNc5
VhHUCw924/jSZSYGV3EoNRgpzsQKf/IfSNbD2aTwkfL7jGH7bq5u34in9OZ7ErVF
WO3mMe0Z/udTwXF64r6Z3K4wGwu2wW4B7C4SY7xEDRLXIc/EZCi5ogU64JQLJuCi
wpnDdR3E+bSFlrZZqRFRonXZC+Hp1e6YZnikHHj52AuyqQSiIjNOSSZQqYvaEjJj
500+HkeKmNM2Hfmy0e2Pahwp3QkFcJA4ZhV/1nWUFpxb0XGmhva2DdOVfMNmrzor
/8hU7D9R7ahNFr0waj879Vm8M8fpLz3rGrEQkue24vI/BSLqdYxJNH7QmQ/YsZ8v
ij4oBKPY2l8D/njj9gESNxdIdQXwP4MXtzwhtS/xpd1LKFZ2suu/GflkwGZF0yEw
sEbAyPucPUb2TYngg1MZ1jArZzYLqaNLhrzPUisLHaz1Q++dzDM+zsQt8XlCvy5v
bmu6Sgq4WzU0b62Wi9EuiuhescFKgVMZZPGlk9/F/I4mTQq4SW6um+CgTBrJJ6Ar
MSqUK5EaLokKhZQTCdcP4BskJYRlItUn8zh7wX2tWrhJYD2PWhdQlCYZPCObh12/
jTPBCvdrUApsLvBHHAqot8U/RmnnBeJOP18HxiszuTlL51Q4Sfv7/GVt3OcI7kpj
O6CDrB96ppFQpPE+6KXxcJJff1QXj4BghYOt0TfLw8AF2oRQocrOL1XBZ9c1cNNY
otlRqQ3EGsU3krU/Z4TfCI74I/aIMS0HQxJnWhXupCu1j9MX87wlmGR0cX45bd+R
C2TmgnVoaLw3qGX93sF8ntgaSKY/d1d6wExkRIm4fz2gf1mHLEI61Xj4CCCloVZ3
HFxLLlAJFUGUbtmLftRi1VvjRusWPyqlI3vlmQDRucoC9mr2O4GGURnGLFs3b9CF
u0a4K2Q2u3zE4pZtDum85gTzDX8GMe4vThTN3HCD9ne45pFAAdZJjkd3gTMy/oYR
SvXN3KiWqaNzKUX3lvSc/Bp6hNHGwAcpQKsU8xvzNqN5/7xj0ldNuFEi0Cydi0cq
dRjZe5vF1lAjCwpkl+JRYID+KP//72mGbuaTZhMvtsc6m3Ya5vyDvypTOHoUgA62
r8hLFMhwJ0IsnpAOvw7jlrxwxlrkwgy6QS6Kdj6cE53i7TV5wGBIhfL4NTaGa6F2
xQRWRxu4oKGCqrvQ3tILp/li0an3vycFY4rpTZPyUHJJW/DoYr8pVEuxY4knpoHC
NAE/fMjxd06TjCkkXr1nyj+gUNqupC4VvhCum2S/xj+2XcAf6Xm+Jyv/NF/4gxMm
/XMScTAfxSnia9FAPH0vw2dGa3FtAmwXguvXSfnb9VgQZESA9kLw17t7it8Q0pSG
78qRlpexoW2Z6aaGqqz1G/MvDth7dfmA/cZnWCcVMWuu0bXlyl8VpGDIcUGQSrz8
jPyBk1PkKzw3a2r4y9/pAHDzLxatG1tenHPhncY96uPfzu8nfQYPKM5q6CU/rcNv
PrxpiIiIHhacV0gpymgPb8GNkEqFsqDYP9oMqzd3BVJf5VM8szRpWQh69iexCx5Y
gMG4t4VOk74vFL1F7JJVpRUnc8Koqy84mo/2GHjTZvPSYMsUtcdsnd7/bAdqYmp1
ka9CzW/RNL5UYhJ9SLJ2OabL70ROJKAG/DOXXsWQJ0Z0daVOF1qjSXWoU2wciJJ+
xEjfZ8LZmyLXR4+nbR67KW7ZLy3aAOAtm04lzIT5VQpYRAThz5o3S/v0ubMjztPF
G6LgbzXijT+w2YR7CDFZC54vs5lDyci0m+ysqUSmGDZGuSg91Caet9BT4H5wXYbu
VYYvM9k06uyyYnBfDYtcBBwdE+JeyvsGbts56901x+zSnmBe12e/fKv/SvDdb9Ff
yae7mcOKq5rq4q+gtL4sg8hCN2ZWFdo+D0iZOO8Bzudx90pYLWlaog9LfeD53QCZ
SzSjReZFWqNo1rPfjGyU//+uX0TKQBDqydnRwLjWRDYZ4mHwc9Bs81IJlGH6HpAD
s52Z+aF0rFyOWTtXn7+bj1JmaNQ8kKSS52pNVLtaw/xIxKtqnGg+5OIE6+S5ZncM
6wiQLzC1FfCBk1CY+PUqeN4sb5Acp5hLukF3Aa1GjlL5IoLwnTarNY3SVQXUAQHU
q8MhAjwABdC0g/9n9cydUuE2dEQcoSBqAMuCacw5jQJ0koYO3hWyBAdeX3YRlY8z
lCqakHSi80oo7VktTQedaBd/0nd9uyjj6Py0Jt1GXyuH2u6nwPzT3oPwSaox4cCJ
T57MwyCZ6EenbA4ahSf3+wWjIEQTmVmuSb5OaSnlg75+sgLS5ZBW1JpHRweJLGfH
CSA0jBzPb28VROq63UYvS2iZG3z0yhqBHb0Wmf82/f9XpJmE7ETt7Rezd0w0Uw3v
yWbH5saPCyu2Ptgf8p7smdFDH9V1OZHmup4Z8ec+EJfyze5fmQ5gGryoXUci8Bht
mzG6x6+aw8BNbcpe2/NVHMCnxIAvRvD1nFyxkEGMJ62nWhQnUYkCzYQj5OT04hOt
52n+tPyxohH+wvIVd5bD0vJDy3age6s6LDTEThj02ub+z7IH6KydWl6px+UD1BzB
+8SOoy0I39Ym3lYIJPo5YJ22YiaiEL3tdOQJB6hIWzKGKbo4NGPliC57aaJkcSGn
XTpipXD0xL6IpjKIaNekCXxaDjnIoi6u82inLSzYu7LvoEO0gT12alCBft5HGFl3
cV/YW1jIyyI07YCqi9s47P935lMumU/tYfGhwjsYryw6ZxCQ/7TIPAKs2iZAXYH0
Y9s/1aAgfwEwvZSrQpgMDp5UoUmH2qK7Y6o6P+6zE4+zyUOVreVnDtxbjTNtqWkl
ld7r3OGpmItO66caTwXu73qlzjBDflvRB7NxCKcMl6hm4XyQ9qZ39S4RV+oabuxX
B/uvqFtA3R+j3Op4H2yXUCYpxmZ/Z4oj9QCJEo0vpGB6njDRSf8iUKj695S7BmD8
EgIUkegXKOVawy4vsJphARi7PslOATIN7IXm5/Ge92v2WS56qQMN8A2PypduXlsI
bQj2fgiHPf8ENX255VLMM455r9769clg3B/uZ2NBPQJdnkOApRXVXj744isT61Jx
64BCb4/kLJ6w0cA/V8CSW7ZfFGl/PGf5fpMjXj91kH0FQdan+AbEP6MnrDbYwLQr
zcobTLulCKZ/wWhI02KX/1ZmOgtZQe90h/K8YlLsTXrQbHYoGhs/V414YypszJO7
LBVORfrgVAlToQrknbhg4LEHcT2u2zBXsiLtVANKVZIxhGivqcaizsVgAN2jdjoe
pe4Up8XTPOi6QT03ELfLvKMd50QUuGeJTE6OqsndoHNprDGFFWk6e4RFIpfpoaYX
gBMkW0452rC20tScnsSxCLWrFEwRKUk10V+H8CDD7kKS10cNpjwUTaIuxZaCJgjT
d9m6oOL3kJjAtZeiwImOvCqmXikMaWfloL+XxeyYMTKpgqoErxcK0JDM2k7bN+Mn
4+Kc87tcL1H2KvSjHuZEynLHu0smcqrQ7dD0kZ1c2A6ip3wgAX/jAWuUBb+/tcQ2
otTUwcMIHScolMul2RQMArVqQhug8aoQlQ9XSQxKDYJDBCGxVBoG2raXQ2zi3mWN
/NLMyjc54KqCEe9piRjgFveUq8ZaR3BYB4CH9d/uFjOjmIJhzzBOlXMnIa0ntEWk
nDJrZbnQIOyHMHYZO6vkfJRTux/CGnJiXOAHeKwYoiaxeS4PPzWv/q+wmGpbAvUQ
GIkiU34quxjf4CcZCrec4K/xTNNrW/+gqkfNMVB4SRk1PRho5axsqSEIwYW/+Zac
V38rcpsZl88dSB63218u3sKtN7zBJZhzEl434lpGm6NOy4E89GwZ03HW1x4ZIEhT
gq93HGYPjNj/y/lhj6DTbtol940YJYB4g2F8w8XO4xm88YtO/MwR3ZpyjPsGTrAI
HvTj+oojAXP21VWn/jkR2BP8Q0UwMh92pA2jcRs2/7u3wtXcZCFDuqJ6dWdd2ibD
9PuIoLqVMAeR2YOtIHgVbVRUF/AS+r8m4Q5cpmQS8qibzsjNNV3d6wOTbLf4q1ay
N3Mb13zWHtC36XPQ3YJnJignKbh0SdjoeGL8jvwEGa1Cn/IRtvDJWhOKu4jsmi4H
QViNW3tTThacQ4oUYwW9bzR2CrtGGbQKRR6KL4KhbG/cpQYIQyeI76nIJVBbFQgF
zlZgvxSnzz5sOA3waMqZxMFswBVnGFBEExAkQ3vg+Q4F8AWXuGrlPo95yDqPgl5c
CjVfY5+qfyCEeGG5OwHGKzElNoRMLh6C3bSUVZhjSHkIDMn7+Spbm3u2pTynSWlO
qCBfvL8AOLHAbkFLaUE9m8F3KqTns4OakCLixmVnEcNdn43oCiDo+wSmWcekUgvD
DG/83rjUQTTxgnW4ShfxMydUIp6Cej/4vP9mgiKhopi30DKP9JkCcRd3BKtyn4P+
yQzPCcgZZ5LUoRnUUh+6BDXYdZYkleiyaEERSbnV+s4VDENvYO1s2H0xdG8ntHO7
jmVJFtrj2Up3cApMgnVeudtrJHTcZ9QbhSllxIHr/bP5pPSuoj2Kx9Rt7Us2kwO0
yt3ItO2wJtJYzAbt9x4Wat6+cVOCs0sAvcM6h3lqombOozFrlio9EGhZPtHgE0Nc
aMYrVe+jd5mlVMIs77lbgUliOt03Gug6ifkWWb4I6AwKeltb/RCanQIoAH1q+HKo
N40b5d2UZ6UiX7X0R8ueT+znRyTvKNmdmwLTMgDhX+RAglTDP6D8xl9UVGKAYxkx
49HiXmrC9w1nh1RpKrHHkoleWvMRsC5FO8B9YhUIjFXFd/L665t6Wh6XsWAbcf/o
3IOYxh2klX9jPcohyGTA3CWcdn8xGIAaHD21V3bghUE/0TRmCs3yQyGpdsDY6GfX
XzphgojnSBkgD+CvGTl9We9gp/AQ1wTUF9wbUzzukzXBtPPMVGOt0hx17ypa3t0O
fJXhj6SS3VJoURYz9pV9F/mHC1RwzwvZR5LiwOQLAud/vSxnS4b4z6Ik0e01b8SB
rRzsySkvvg4nYEzJYlJXwerWxr8I+RxZw19K07FWW/P4+eLbRGjIe3Qd53bk/qgD
ey/KrYz8+JlZHMRot9P9jzBDm+OiGACD+qGBy+SeQjHnSa10EAcRV+kSNH5SZGOi
HX2oVuCBDl+P2SSluU993TFyprbynR41+ic8lTdH2oy59kvTyKCAhx1NWxglSiCP
rm1A+JkVTWfQQzMRUl7a9Ftzusiua62Z2eZMrJ+uIgR2UkU6LS0XKjxdMRr6Rzvt
8dqsJYxvfiBjIqvT3xgnSeWXWJYRTibxWGDOihhJDMeN7/yzXK3tmYa8C2MmGgjj
RhCWovOTXUCX72AYMHg442mlbaPPmwFGRKn800rO3fUfoOm9nnyFOMeFE11xG7UR
2qCLv2TFHQHLy4ASVkKFdctGZu70t5LPaGYdoLWqTG4cDfLD6ZScHT4FuQBFC+Pm
3o0XySHhBODmaaTxBTA7yeBaFX4kcfuVdOA7Gmy+VPpqgayfqoYuhoLwU50+KJD3
MtWWbSoMjX8bfvoL5kIiCr3hiP2LlnAl26/vnnaUvUZigV2jZTGu4KACkuiFy/+Q
RXXGFPvLcE8IFeOQrzmH1LgvlRDXyeCIILTb8vLdNpKD1drFcrLJB0C5hWx40M9I
AWbuETxZnBsVtuSXqfz/dBYGurXWZlS1YC1RdIs0KKrcLXjJGK5yyGYv8y3QsfV2
mTPLCFQ32OQd2/8R+8D4ozHRaQQcy97oOezw51SUYTX9tNZ/austAXJ36ejsKYqG
HWpkmiGrpf4irqKBApqF4aTKs8vF5vTOFFapk0tCBVyRpi1iJGwpI2Br9wlR64p9
kSB3e5gs5L00MLlcCHWRHUJ/GH+fqsEqZV0Qw/oVeWlsmO5U+rOtfqBnNDeC+sfQ
CB6cmvZzHy9DnAcLU4YkIcDWWszOCEsi5UO26JmIFTqck4Q7Y2StMcv6RHO18Rz+
20tUdcplDXV6NPcyFke+b4utNmgOt1TkF4bZcG6FHhjP77KFY9V+Srcr6s0Lo9iH
/eytXRlhxjAEVqJf+XtMMA1eN/OPORu6rsGIQ2bu02brddxAY+j6vTg2AZrPVEre
4Gwoni5dLhFBPcUpW2k7QI68TdjTilsNkIii9sO2eRDsW30N0++x5ZjGXVIuHE6q
WPo8mE32Up63KSEHwAWZgKWmAUBQ6ZPQZf+dvJSmDZZOTgBb5GTwEyXnjEa86sFS
ee8GGq3Rbg4QHcZJKRVjIiY1m85DeYlXSEa+tpn0y7IdCQiPBHqPN9zUQCYyDb7h
ekCfaRvcAfl25yR7iikxjQxJhdjRzz+7UrbfV0cs1b+rmHOEgN9wkxGjY2ECYu3v
6hZi2jhznmQcsbfeNh6XYzXsdrhKxWIYkSnywtha8r8i4WGG8fleUbyUcnvLsGrZ
YvFWojcakVDMrjm3bPgaryQFE+JgzktgJDtHNhZ3AoIgPx1n8BdA6tu4QCMfB8GE
NytKSO8XNY57qxKQbdP95gCo8dqiR53bJWWVNqwu/ycc+XMayDt92kJPJvZEuqe6
W8Onxu8TfKmdJGq1k1Z7oiouIIEuYqWiXtiJ0IPgqZ3apKG4DzG2EWBDzfUbM8rY
aCOINPR/V17uwxPjjPLGEanXOVauaqj6nBogC6AXhBHtJ0jp03vBxuDXz3MdAFCA
8Z5yqK76zL3eI/72wAyAZ8AYanrTJ4UQ7bMoD7O95ZS2xMKvMIZBtaAylVOhI6qN
q2wBlvkFGVWGCgtUp8LmzNFjDaDEJJuZWybRnX+Ecn/NaWGBlZWKdUpFgpJVTfy1
4yA+D90jJ0J035Xm3BAkAaHoeZ9TqMbLGoDzuaCfUfONmKCvpkH87fUdYFVRssTR
H+noOk0cJcHES5Z0heAz5xZiH5rlmiGakFyJMg6UVgDG3axRSg2bRDF9DpRh866f
7kKq+wzYpkoXB4dNoVC0OLI/wYBS0fjePncyssZii/36F05A473ydz4gPhODsEjW
j6J6iTV2SF2RzRXvpX2HncklJ2kZX0FWyjfAsWJcsyIsv2ZC12Zw44ZVmKMTwmb7
ti90lz+XaR/pWA+ZxLWxStQgisMXYf1dru0TPYdNH6lR/UNKnOnJu6bJ0YvKNBW6
rTm8AIjA5e2lDhHm6Nyg5V9acdS5vKbMRa+AV6ST5BNXbMtCX6Hln81a8n0Xh5KV
YATQXeYZWoOmPkz0k2/ir1sLMk4S7o9kz1VBTV2Mz5T1NEnn2dsi4kikep5SQeRS
tli6CGWbeZjFKFYR0gMICRgRUxUAex0SX383NeDz9fvNJ3Sl3behLmHD1kf7SxXO
wR1lpLP6CFPKyy8ZGh34yGAZXxhR3JB2KYWfkyEsNfqH65qE0TjZNQFvR2VTF1mK
jaJWm6/yH31/shwAZbblWK1pbH+79WkfizuWpFd06QfRJ9D8lCqBLhoyyh3rnaRb
ifvnIUVJdmoqIhT3JWddrleq48DNcXKCufaqY5qcgk8vrljx+PwyfqBjOnELD7Vp
QO44zlYyW+FWWmS0z/GAOlrp1FJY5Yu4npCm4gsMqHQYI7Zgudfebtc8fXegNX6+
epL5rU4PydgPDoSz9Cfhp4YMl7RPtLBWJeEGVPHUM14seqn+XXGXcaHyw/aCDDkL
KGit/R2BOyyjF7BtEs6K3QLQxkb+RI835EKySxzEyVG0VTYfSDPxUL0wD8AimS/b
Js5KOBTN5rX73QP2w7Bizp4cZJQkB9Fs6APme3AXkegZ6HGjx5axeoxAfABHeNc3
8R0IIKomYB7G5cfYH0/5D64/ccqvP2K+IEbt6CFVbnZf+QBE/chqVMUbk9nI9czZ
W+2IZe5/fmfyP1j4UtgFX3FbWkCjBvkrAlRgDtfHqZTL/r//zdAmEhEmeXs2VPJ6
Xxce/wkHQrKi2M52anKYeXtuvMMTOybuHwvGrlTQEnvfZ+M/wmFehNlcqMFhOdCr
cJHtHeqXWc4YlK3o69MUqoFxAZebDwjJQUINhC/gQINgqirZojfV7ngHidt8w6xY
FaX62+wEDham9OWzV2cHyG9Plgb2+08eyVwjQSPzFZDUUTxlCqdRXRBX2kazaGEg
3M4em0G3NudO8Ot7srnaFoyLCLsTz1TmUxuaa8Oo4qyccESraqnaLD86W690D4BX
eQxS2nihvD2VoWPzVomG3PV8OuxbgcnrrsI9aEbB/kLIgpKOFXR7oj1h1OEqTkVV
ycNsiRkJ4Dh2BIT0Y200xSzjB3ImaTUqIYvZondbLoZwd92IRyEwK2/vnouXXTQF
rHHpWoMdXnE87YquhuSVrRmM7K7Qfuv2zbUocbu6Wsu4wMw/sUYyPNrisiDPCg6H
q/7lktEdbpYKoQ7PooORp2Y7rLOSLBbFB3YX+sytEgfpwXuny2oeJdP2PufClbtD
byw9S7zULg07tUTHEkayJTTS5lTk5jlPRFywv2kDyGg2/UX/d3xQawuATXlRnJ+5
InNDsT5p6KZrB6lfoUj9Qt1q0CHY85tfKc/zA4MQ27Z3ElUfgvAUv8s1hOij/LNw
9wTM8vD3j6x+fNmUz7j3EOYHFhT7a6pOhOdbbT+s4w08S6Z95CnQXIJb5UqX/38P
N8iE2C/CFQaSGTvGLfYrMDJyKOYSCsYXCkG0uKEh94bHohznN+njB2pqfohPzOVM
wkc56RYVcWaHAEjiL3BWp6JxgubnwhYoNGFz3RcZFZvipI16SsmnOw3cRliN1UWb
wU6vDYmCoWTw9lXZO2UKANaxlmhCa1B5QNEwiE/w+lAvzlh6TBeg55f1r2jzuYV3
Mnbxu2lBXWQL39YBxQfJ+jf8JSh5rQmNBtX8WHA6iux0fNHdOcsfR2RQguO8D25P
2l0gTEytglK82vVlbd1OOnFaibC+Ins2FcMvZ265uq/awDP5ctDuIqSveImvP+lt
x9zh7XrpU0F9kfqH1gtXMRfb2QpjVEhW+SvAzI3Pw3OHl2A28n7T4JPgJmM7K65Q
rgJWkAkUAuYG7XbHOmRIz9yow3GOpj82MCVhtHrTU52QnhA2PnMcV5B1oVwePS//
DLlWsYBfpAI0XegsAWWRvYxGsqQyVu5eN1l5dQsqb+CMb1N192cJA1ITzvPpFMO0
xE/6GFZ6bBNpkTGcHmlal7xxOpTqxN+vneKJyMkyRRHW4Eev0MsyJ21MTOBf/qsK
AtEUDdIyoWrYemuUZUue+SbpV3AhtQd3cq0s/+DoHUad+aJWXgxjaMes1mjXaQ14
dWc12Xx8dRkYdBXndr64nCYi42YTYQCQ253t9dkahjjHQ53ACchM3YNqUelOEYKv
8FxS70an5Qu02XWeYx/AZEvqMvSRzOHPkUSgeaRer3vXywUYQZEC0D1Yi2HxxanP
j3IxspN+CthvvESgL0cd+lwtxsGMx6wiXzuHgleUb8fdxsAs6S3pJTvG0CRBdVCM
2Sof41K1gjSoimuezxy7aZm1UERlrI600W7hFE2j65jAfyc6LBO0sopSWdFWQy5r
BYtjIODx6CXmh4r1FqacxbmF5eLdugbWfd8SUJ5F3ENfcPX26sWi6yBDNVMxV3IK
JiMoSgGstIIgqTTrkBBxg9Oyo0wsOZJFiF59kfNHbCdL/dI/KvH6SbsOdy99o3ly
UDmJyUVlUxWwbvgwq328x7ByttBZp9y9DjHtD7Kiwe0v9Izz5FvchuNmXCyiPlmk
3jfjZ4txc8auvb/3Ru1GwrmVfvnJBX+9dFcDW/Ip+jYwgfwo/JStA21/gfqe+Jd2
D6ra5ms0Z57TDdE+ue/pnVilAl3f9EBaRaamSFJoLzbiLDpuraOv8oB+WazHOWNh
V3j2iViKEdY80ml1pLs1RNsQINTkN2/FBFjxHAg7jC5lHmBuhI+VeGk5k9VgwFIK
aJKAjKLUoJbLIKEXdK/46aKaXues21YMQh5YDAPS6llZ1NxBp9X+6JwXzg2R32R8
F4Pab7k+EVeCACBR80L4e7bbOOdP1cx1YZHFmN+qyUJJljx6avcHkRw2GBgsuK4I
BGOWK0wskaMYz8NLmnFnQb/waN0Xu3LQmYMsKAJE2XNww4Fl4K+EfAS+Dc4ItXRP
oqgJqzDuD1+v6YqIThgnW53vbm0m9LYHM9BDnkIZ9ph6KFXyqo72ldN42obZ20kr
3Q/OBc5Vi4hnMAhjxIb+oCE7z6aHgKHObepgDe31a3Mt2btTJ9YHUQZPXnZy51cu
XUx5+QjpSumYMRF2ifBNU+gnYnzvUL5dhA7KVRIqKvf5j8beV5jPZONt/hoAI6cz
Qu8cffJOx3C1xo3HVCvOtvFlhR/GK24qHnbTp0gYHAZEzBCYIvOpfPKQPU6ejl2B
TKdKIQDD1Kswu+jdaOB/a/DolPu1IdBwYuuuBBMN0d/AEY4vZMym86gQJUqa/gOc
pJiAc8e9Lzw4dGMJRXp8hIK9sncpwdZautvO7Xo1MuoczQkFtQzqktV6Hmgr/ici
/EOG/x1z/lZi7FUYJlo/yfdCj/AL5j/5KHvoriZGdF5p4PMBGgy5DuEsYzAidQMN
RFu51yX7AtFv2zstsez6By/rhrhB1+B15W/NKcmPe4jyx/haV5AevM4gMcsRr9Pj
rsvtXzjQOS7EAOGZiE+y0TxOUk1y8WaU18h/hl2B4LdtIADD86/vv/UVLqqj/lV1
/OrfK8FY0dAdoSAt9yr5SkX0XpMTxjs7N74mZdWboVDy1CPF+GB+jxB/7tMn467l
YxYeppvPu8FOvRhoVIgsKbYY1jGrwzCmjP/vnTPPk7dwhjaIW22KBTjZqszHQ8T2
U/ae8YtBK9ojZesH/kPrj+dFm5jwpfh5xdZMUTXA6b6eB8krAgLHc21RvWCOqPvB
g21uOEb0mlmw0QenBWnLvZFjn88bqZ4wM+lV3qQpYisv6DJPaeMf+Ug2M4TxN+dW
Q4qTEtkE296UQg0MOPwuNE8TY6tx9j52rJ4ojr/D2swV5de0px3ICA7hzK+xIzt1
4abyDWaEaV1K/vqibP8EOzNDqgbnE0eEPzJDa4K4DzEszvwZM5GbZ+MQI87ZJmhj
0MS+rbcjQdJ60z2w374GfSROpQJZ9i+ZleEAWqXmaiQA3ZASqSKf+3yxEbtcyItc
ekK5X61Di8+uSTTw5sbx3aNvjw5ZdhPs1WN+1Sd0MObJbzSn7XG70s2XCLqPPR0h
1XI2BOgy0oZmLKBBsNVtU3lGUioIZPzTN1NOHxbkAOU5JZs+PcrmBZFQ/WZn9w1e
W2XNqdpgs0JxiPgNzRREf7k7N21Bnx9gOo3/cvVWztcA1HLtsWr6En5tMOUvbWsW
A7CygZkqcbDh/UsGI49oRS57Na10Jr/+GlXZN77JiVS8Bw7OKDCFMha5lix4bp2i
UYrMcNaKbaemXUj7BE5Lstltfd/orHeSXX8llp3FJ9GpuWX6Oj9jp+EcBaaNCOuD
t0QnpFmIHdlBVjZeLuAYMHIcd+5nQ5L+HsHIsyD4J7zvryCy+pAsAVOSOISBGT9U
O0S0bEThYFU0Y2EpXZgvC0dZ/fgpWNGeOIOM0bUmpjWL0E2gN0wT8gnoDVzmSzNB
MJ83SxndYS1C+ehl/PlQ4cQP8XMLfWr8fHSqlM31dEzVnh50swEgfihDARnkQsU4
AeL+6WxVQVUzEfhZaaEFrJ6RDMUK8thcFmxdcsauuxT8Fi9Go27UcnX/sdUp3b4N
vNfhliokgWItJ+w7/g8ClFC/A/Qb3ls1mthC4TUcVcfKuZLt5NuBYzfDp7w30l+h
3YV+UZHsU/CsNZXT+dQPXvZPKdTp29l0tu/3HyppLIi2JrmYq4PM/QDo8cKklYFR
dp3k4ZRBxcApx6wIqQy+lIq4bJ/6/yQaZmBkNZIB0J5N26uniiGSJMWlkehnqxh7
ZPHDNjhllIXwW/odfFH8BK2xyBCYCDKSfimqEYNDSFvsDL619g+Hkzyi1VLsEN1l
rC9rOSKQntLXJ0ZT1nYspS+pdyJ3qMcgxlpfLfHLpCngEY5MOy2vAqEgUlahMNwJ
EI0D5DtsMNwqCx+v3PdPFnd6pxMVEuX37naEC7i3ysVZCH6GhZagqKBDB5NVodOH
N5CXgnBfoeQ9QVwLYqtg19FNZLmiOk0bfVOMnNFV3NkQSObIGRTDC/vy7xh9RVeO
UnEsMhmXnNrCjujgzNHmKkND3pR//oCt0qOa0zm+RbCqEKSOmnjLS/PFbC6AzD9y
Gfgma1ce/RD9cfb1eV0R0dkM2zKotzjuhM//ze0piZQ2FyTBlzfoCANiHxHbMG8C
jjaA2uArQ7CbeNzy985CoRttnubmjooo1K0LIMYz5LD7phEVnauWghZ/NotM8UUZ
SAOEdnPJ+S/Aqa6Mz6NtzuZ3iqlcHnxdreg6wsRiG7oodwt6zSToZiOlTPUUQApn
/d3ISJtwcBEDgNyYLJOKsDiTIcXrDGBcfJDB23q1paogN3h6KcHqPz5fFug9wr36
SbmUKjEuONNA0l/DXBfhb84RJUOmmAlWUeA8xq4G1tnx4l/sTK+hc8m2ChoWxNOr
IhZV5QaJKb69Fv3EM73JVgx1rPWJQH31MLLtZtP0qBb1NZ99AS4VmPUC0/0oCuL5
nQF7JE0HwjoGUpi9AEQ+ZBtwJYpgwP8m683TFgQWxRCoush2rXcT0xx9l/MBj2bn
Cbbia8HKMkwioG2PHxB7DQCjrxHmPzp9uRy0GuS/pBpoTDrEBkeZ+Y1SWYHU67pf
px5GB1GOGZyJ63gIRX6mzJl+oyc2tXN/aIXuXjIVuN1OPsGKeuaCkw8TMTuR6OEp
gSXj1NnI3i8oF28p7GgXjsby/9aZ6hjj93woVY6GpLeLU/mAD6+C6klMvthbLRK2
2lBmi7alIYdRVFN8KkOmcmT7Po7qG+IjWpCKRatsr/bOFNQqeEhhR7ldveJPL/A+
HM2Xa47GCvUTr1NNjw5/5uf84s1+I09Tv7ZPiEK85EiDGnSQ7sHjSJybIT5kOr2A
bh+aylOgrHK3t38pKaDO4HMpffWQiA662Rhqx9I/fHdi8GBbnq1/ObWcwCx1shTa
PsBYd8EWUuPs3P3ooNObnLzs3B0BRL+lZflcvg0wcfTrbf0Lxrh01tLu0GGGa/Xu
eKB0G9NKmLSRvCfJCZySUEdTnihsm1D+3xdybdGMQ+nSiSk0tI7sp/xCIRW7X0No
lu40wNQ+7ncpdOFOPnfKGdpovoYOKJWAfRL+Jxt9xDDKULxi0FGowboXFaVZBRZx
KFw6qMvVlbhiA7x7b267P6DWmM2nlVsxMtd2lY0EWNbjBCCZ3kLKqfVK2W6r5I78
RAj5Z6aLZG1o0QXzJpXdhqpFUMZgYU7OEucTDF4q8OTze65oXvVgQFFpv47mcm+h
6y+z0HnKtaZU/BIxmkSLoUNXE72pAcK0lEj1nCaSTZH6ooRPeGWBAWFqbXhp6zC2
idO5KqkEvSyUhlni3J870raJJAZrgkrOitoT9qsYT0isdI889zKYAD3KKm10GjUL
K0DRY2SnCTIMEWPo1rUZydDfLXUaUEqtkSEaPwYw6H13OZRLC88FLXR4aPpV5OuU
Mp9gpEqp4EzJqzcCE5dbXupkPvQhjSn+Y2tc7GvZpMQbiV72ajQP8UPiArIJczLU
N1VonSgTC6NHLtM2XLFnG6q1My6+UBo2UQhqvmHxerNed2K7j30qWZvl+2IjR1Sd
dh+Mg6+nurVWHekcMit+/lJ1LXf9k1/n62DOepd5oXP6ckxBy4Zhm1N6WEqABAjU
s/Fy8hrnna6/NMFg41fnMd61U8IgHlYiypJduXbROLgm/hp78opX7qNS7G4ijZ+p
1qjVW4hDNbf+DppdYv9QbekZaEwd5le0EOyTqTUZ8Un8rFjs03Y3vtCbsgUj1SNy
SmwSmtHyh6lWekV8d8JuwzPMMeWO+OEq81Yio5N32decAbz4vwrsm5HqGCkIiegX
rfevZPvGAibnPpun2Y7/XMkF/qqSTjJ3Kqgeu5U6f64jctEOUW+3XCQc6QptSYR5
cdIvdEt/xv3/roCLoCpNwvHL+I9vzBt0xZplr6GLEb9anYTUIzI3n+WBnLzpKVVF
0lwt3oIC0gRSoPZFCuPi43jtWRQCh7j2GtmacH7XOUa5VE0qWODOyvDwK0xDG384
JEbGditiwG1drYLZ1wtggsUO8UlGXyvte7rhcvF9BiE/Ynlv13JqXFkIbpaMFix2
3cjG+j9qMHNTqpUlFON+DtL0HW+4d3384c5wW3zPSDfmzuz649rYYFqBMWxCzXew
2lgy96LUYBuoOjwvNhUxMb1igaQ4Sb5k0hcSi6EIQpcwhUtzbfSr4iuxuFA96URD
mpNEcuVpfivn03MCe8HGyW6/fTj3WqtxFkWxf8a7eidBWr0uSbrieYUsTWbVxuPQ
6RxJ4+LTkEo3eThrcZoXC9v0Ij2Rl4IkUtXf9wgFLQEhHGmeSEttznZiERvxSHzc
vJTE+A3XOJV33FtGevD5ixjdI/0UEnMTAVr2wHhrqXsyqNrH8wpk5baYH3/QoLLV
Zd6JO+eUmJOtyzcoAYvjM0pqPqjE0hs9FMpVIDIW6oL9YT3ynsZyqC7Ih7nPWTir
U2FklvD5zzmA4SbLye76DwTKOVf1OfOqd9TUVZ9ozHVR3tKCeAPdcvL8x1h0O6L1
/jfIhUyCfTSY/KZhtKPfe0favPPX0bw2fL6ZGBoOIWQDpXCevyZhD7lCI8U5rhB4
DSb8uV9C4XzTcSIBbWyXGbq9XS23WnvONao+MynULElGFalkMZ0uuqDTHNbT6pQV
e8aD9t9Jwy33QkNWEsSE4W9ISTGHZ+685wffZ3I1VWOA7rA4+bJ2ly6xdAbu+OPR
b1Kzjbq9i0W2uHFfKyNGIjrWVc3EtwGu9yYHrkOUUkBi0JGNO/ss0pauzF/t0xVS
d5BVXKxVPSUc3NG9X7Gk/Z4uVPiido2neo2aAo4tumUIAZbZzzAJcHWzY1T6U+fk
32lwnNrdWC+jKOhEenfqgZK4lMcLwLZahuuhLX7Fw77NAgGHhKLzTzZ8bf8wedBz
k32JnzcLlZtt+r93EjiopU2a5Y6bqEVMmFWs3JdO8hOsV0QTdKYbu15sT8eHXNsj
iJwBcmE7G+hlLJWrsY2IwVEBn0GMOZNUqe1tJETx78w6J55Bdjn8HgcvmjC0aBoc
8qmQTM9Xa0gQCRxWQJL/TZJvQIaZn37jhJyE9a8ZlazTPn+AHXMT2ncag1lTENDc
sT0G5e88N3UUJ+02F/boHBFgNKlTFnnc2XHb9D2t4WYwVb7Lus1mveOb6PD53GZI
VX5UVyHn1Kmk3yBe9kg5GWYjcF9mWm7u3e9kU+okPjogtGJ0ACpDMYq2XnhDUEUP
4T7lDsR77Ca9Jrs9NXhFxgf1Kk2MNBqXlWL6m/j9jOpwBtnypkxZ2o/DshBMki49
ADCFEplcH16nam8bJOeP3OHbMGpW9AnVMzqKMpsH+uprz64LNb0Bv+tN3ww4d5ny
MlWIRy37kZ9K5OkWmoHTq13rrENykMp4mvSHmxD1qKQ94lNkfuMaISj8G/gOLKyV
b7h/VB2OQQA8+D7UEjzd5aRvUhrEfI4PKkZtFULfsbL0zEkWyOTAFeQjviB7avvs
V5fa5tquTKY4/tQ7K0D8vuWMMvzWtL0UQ3X9wb5r31g0Oyr9fdbixehlYSr2TjzB
tIR+AvS4OCbQIfRzLAh3p8JsqVawba5OukaBAM1DQ2l7Fskvx0QzpGu4pfKgmKPk
QBK92+Pkf9Bue+1sR0/bcAzP1+JYD2kTWYJ2YSP/q3/fyXqWb3JK3/eccRKIeiF3
Rx5MsRwz/lyuxjuMjHJuOM95JkBShuZ3/wj71ocD6sbaDOHF1LvO1ivLwWuoyARt
VxCT18jqVpFr46nIyKoNrYDFxE7P+OPlE7rT7cQ2CIbQW5bfa0WTTAjDAKvW5Ibu
Tjp+g1ZEb5/h/JcqEXacmLob+KhuXF7Si0VtO4Oa/eS0nmr2zBUoJavI6jJx+i/F
QSaBd+5VgFCV/6+Ewe/orj9T09t+gKx5fqztLKzSPo09HAUuvLtq1J+2Zf2Ist9C
6uKBYX/tV+i9rpo1mN3RjV9r0fNUP6+xvxe2Kuoi7MFuMHrOYmlbo3NhgctGFAYa
cOsF9hIoeuQSWgVQeY0YUgx7g5HXN65VhNybAEeCMSrY9JpGv3GIQpH9sOP3DC63
shHedpesnOOLtFRDTgG7Ylaq54pS9GCBVDc3GJnRlbxWuXPpRCm3JXd8TzdHC3na
xlhLAlMuSGwqgkvfgp43B8SkpSHM8z++HvZh3snpfyuFMxmysxtij4Pd/LW4v9AF
EoSYnsHqFibeZ9mie7LDJHlct64apodGqQmc5IIqus8xBUpDCoRxssb2bh+H39IW
XFBk2i7SikiJGf+f2FW7LjOZx5BTpTIWiMLTPxXRBMYNCJ5G8nepedl4YrvEgmvq
uIpbv1BW3pgElsGkAHub96Qnrfe1BwST4ZtvNXoPW5FjOi2Pj+D4obOTn4XhXKn/
/uorWeT2u+FfM3aqpdl9XMvN1Ub91d84WO4sXqWKTmnzJP7OzUlhwSr1dbx22PAb
7sfLkS6DlAlBXr1mr84nUqoIIcOywvsUVdqOM2uHOjDBvSOiz4R6ofl+xW9N3rxv
a2xitdlg1fgX6fgrWalaQ5r7meCi4JLgj50t5t8koy8ybp7+RB4BmNrmIQ2xUt0D
tcPCxEFoNymhusA2kKikXsS2d2M7hEEbKrZZuy2/+yG3KETHtrVakklUMuX1sHjL
zcLFIw30qmyfiD6WJXr3l055500XDupsfkeyaDPGbdplWbvrZVOnDkJMcfVVmBnh
Bi8gs6P5OpUQ/RZ9+gRwU2sVlDOeBoIBYIU6kUaX/RYumTTi2P4a4j7Xpx04AUQV
1UcFA7cqIc45KZMfP54aN+dQ3KdqxgDKeCzYjTygRIJUv7uLxK3UijjBz0Oqimj3
ae0o7HmyUK9s1OFzPvYN9uxbdnw4FmZx0gLBxY7zQ/8aFYfyS1ulv1Rs6mt7btqx
1pcyLq53yFc0J5+zOnN2bvz/4DyM/nixNT6/oENY5FPMetmp7L4eJhsetmO1eBUb
X9aPL+E5916QYLzuiFR/4wpVeg4gaMABeEHePq04JghHYeY/NXStp4HlU98V3PVA
ROd/I0WVyN+TVZyUNzlSP+JGRgqG1jFfIx2ReHhhNsoNQ2scrtNVuRziid/wrT5i
/u2gB8j4OdTQjL8QHqxFWVT8Z8huu4gq7iz5ctyXzXoEMOcDbO8/r9KsoUZlko3N
5tLCWqUDzqq2bO1R+fjS+u+m/nks6LrlMeX/yCfzwB2q0YuVvREwJWZ9i+tWox0B
3UyMxjSxEgOcB4PLBtkltg2lHbagZjgDPf4bW70YOORpQnV034QzoQAzi1eNC2Dk
XBBIBgfuuOWlfiqrHkaoSF0V8YEB22XvlB9CUg/fky4KJ7C5/CBS4rtZFd50kxVe
RqDphnTZ/OWpfQAgJDzbrNkVbNWuApYn6LrNR4qeQ6c98LfM5LWYoqJyec9t2uh9
w49vJp01sIiATT6/PfZEQLD+4bUW3FS+er2xYfbE3roSUY3/LqwmtQA++6gGIbYu
KSLZGmrjZwWmrOvKo32eddVJycJXlSyHgbig7jpCJOW40Uc25mg77RIJkZWj7QJe
ZX9TLdmUuByqOUV0G+ZLOQzqBOcYpT/uLXUbHVjpBm91j4a1nPL5wv0ZqdvxjsDz
bMP8/I+GgUwsVvQbpKZgpNt8J9EK122P/Pa5qjHUq3V1HEvUZoAQBnSLpMSe20MW
nWkcL9463x0IH3LZjsvUCnmHLQuEhpTidNKi2qCdhsy8I7z1IHFdvFbaFIr3o7l9
pfukiK5Ky3rV3d43oij3Rr/HYCyidQOqPc9bdblZNCin6M75WQ6F02oCqDD6aJUq
y4BzJ79Iz3Pm0QxvClbIEP/uJkRijmC3QeTmT/0v8zP5pEOv0HqVl2KXMlKJ/j5j
EmjFzaWTgKMg5H9fJtxixTxpMdHfCSHGgINsbULhxAsfawUlvq0XPFqv0B8M5OxA
U67yto+cF0snxbWLX53z9x2233YbVZeSZRXmmxWWlzewCY/8F/8nX0BEypF9+OIq
lkKKLou/rZ1DI7/r17v1dLEHP2cDTRlLEHEZQyoCVyXtVqtgN8jkxbT+jJPDTwWW
7DE5uuLjYMQQtTn7VYFgVQ2FIzHRsHOtnIlnkeQsXrEMz9/BpwD0UuAxG5N20zhA
9EdJIFgNgoFUs4dkfnzx3SY9J87JR4BPmEFxIH0pDZIK+M190/SoSV1yF2QkgNRo
wCycYpNhKyF9XP44NK4PjuV2Zaaokwo84x2DU4eLtaEwTCs6pAHiJMrz6DV8myWn
AT08g1EHzfQgb7z/Q1KVvtMY8V7UHxN4mPFzgub4J3YhA0zQcGXM484NT4M7ETOR
RmeUK5dzTgVGHBOkRhhzDo2q2UMxpWzT0Qsi70q6mtb8lSWOE86df+m0efphFpLY
CyTs+rSiScNoGJ4asDzwEVyK2YpJyPjXG14Yh5ui9Gw3iQOVPJMyAS+P2+cgX8AN
xwDWHkftv8WPg+IJd6At8zdyg72Q7OxeL/vMchTEr2xD0hlfZuvgQrPw5AhDMLkH
HKTqjCIOBgaq/DZuzXfM1z7GGPjNynC3SzW3MJXlMUxpegTEEHuib1yxu8z2u2pm
rIUQ3FFc1cXhlfMQ4j3u8bjIAPtels0XCcjCgnBjXsh91uU5Qn2rHnd4YxMHio3R
yqO6y3EpxcK6DOWm0Z2p2AbubtWssvPuuaJPvnSMgG8j0wg15lDGjI7ivjHFk0gt
e/apjyj2R7xLqrE8YViShOocKmcm21N34gxL8BPu6JGeQnO+g9dZJQtJ4xfE3etc
cnZg3YK7R2PWHlothI58YBbHEzIcf0mWOJQLmaIWSnfmNslhoRroePXRMqo/+RQI
xQ3YmEClWihnBUkKaN7JoyUa8R1HjkrBtZEGeE2zoSxt4t9833NtHUr3FZn1+Z75
iG7ivdFGIDjHkgGlKX+iQIIQN0wiGXwioRMcCmw7xB09U2dvcnWO4q5JWUmDSvar
GG4IIaJL4AGkYCN+2PA8TqzkOkt45kp1SeNSlkj4D0WUnNinRsHdF80y1WFTd/7I
X+gYHA2Jp2CjWGFGO3pybR/z4wA0ffBnoldnHI15LL1TEu/X46kK1tuCxoEuYSFC
ZDOXM2blXxevGonXua4RRD41mXz6IW/t75eBsQzk5L3Df1Y6ga+oEA/PnQpYr7dC
+DpwUzdd7ek3t+PUYMSt/sUydQJ5eU8nTTDC/yl2yiQHhD/Nk1oW6JrIPQa6Xi9H
TcCBRQvl3OckDbYuFnQo+LKjlrFYumyswRhOEPHOvKB5CNgvx8vr7KtwDWK/62Uw
1cOTHNzW1OAZvs6G/0uin9P4CHWrq/QqC/rKiXZWFqahgAG/oBhu+SHriwzm3h4C
+sk0JcVnPWXGnS+XvUEP39sQekWEYyEM8nLWP+rxtlr53aZTRv4vwg5qfYiqs59/
djsJRsZ4YHfm3t16A+LJi1NAZD1uJmlgLFG5KkWru6zImw3hOePqms0Md4BMxsAJ
G+QkbQIZ+pI/QnGQ1YfBj34V60RWKh4zNivuHI7SJYhz8/+ck06jpyEVuzEjzqgM
SOmuQStfUHvfHobG64c/zv+lBVvEAQ5GhyzFKeM9f/ySgSR0gLjTFy/TpQquxX6j
qLXFwwuIKVDoHAmv0Gm+fcJ1eFPWzKdDKcBlzBYyHnNwsqbQXWWLcLXHBxskf+S/
doA2zrygn8sTIAG9+HoULVFzHepm3NjhoWUtjlW3ZeeIcnv6bPHWJrORjmzipMvl
QJmvZtySPsGwZU1Nlag2bh2/Z+5Q1nvKl8e5PkP6KlK7vSDucOJ0RGh9kKXGHCIH
/H72pDBTG8++9h2NPOaDbQd77AVQn1a276PSFzhmjn/WsnjKSmIGZCANhjPgzWJQ
Y37IW5iNqrE7tm7x5c2Rst93z5qvv/p08kULCR6HN9D1zgYp8EhnkH62wP4TUrof
LNA5rSqh31S0u65jte9+rWhBhfheW9BSh8PL0sYOBVeVnqK8TR+RaorLHuHUkr7K
LepflYF1veO0dfHp6RRBRy1WLaETlRS7+j3TVkWV62lYOyXJQkTBj0r+RVhU8IIT
f8kploOC3YAget7gMvVhZENWN1W4nMiwqDyK8cO/8ZztcpKA6CLGo+6rUHE6fcHZ
ICF4vd2aF632IwmcMO9kRaLn1vDO1Zs6yNwy2HYNXHHoWRxFh27rtXskI/hTp9xs
3K+3VyBZnPV1lqQiOMNDhqci2OqfbuGtaHGipwSihLtE3RoA1SmEM9VH32I4VhZe
neSxWRpFD9HEhz9GHapjiBWYzs8eIKHkiipMk41PtbORIrwCyHDpDLElb7oRoVoQ
8R/wX2E9IHPUJ+H+5+dqv3oIJ4/ECJQsr1gz4LZKbkP3V6FnOYU6DEDnYQi/QwjP
tS9WSGnw3YsXTbsVYub4MaZXdfCEXgtxdPfTfK8cKECOp9SREbMcrHNeTlSsC0Yr
4okaan5Vrg7KkKbRt1sWXIOVm8iLBFN8HWPcDgtU8HIroBhaGP52THWh80BF5do6
0k+x3CKpdNPMmJ6ln+iFYOmyTvx2gxiwfCq/vnUGIJ7ZDcFcQfw3aR8l3YOYy+87
omGafBM4SkuvfsB7PwvDX7przoPyUGHZCHpMnYX3hKzK3gAhuywDHbX8LTDg3EwN
/QbPCiLCNGBHY6sTERRuXUd2sE4OaQvq03Axw/jpVFGZ4yVQsJn9b45cJSnlnGBh
ws/R7dUSsb7yCukhfNqGgu8a3Djpjv4geWAAq8yB20Tv2rRX3B2G1/WmCE3NXvNK
B5D0b1ebCnwEkPrblJ+Dzhwnx1dcAxowX60BX+NuCkQEmIAIYUGbk0KCT4DJ8Xur
vrCjUdIdCvL0I9b6ram+D4PFXeMaQNH+JtQAaylenWW2B6zD6FODC+oyh2TG43fG
ulOulkEwaXcQDSAqBr9ucU5NlZLjC4+on5abXw+P/f8JhodLbrAGvdux9dNwbL3Y
xqmFwv1t7TGkvYGNOd1XqRTwcg1JNhqTUv2UKAU26eGP0LjCy9ynWeer6tyHNDJQ
s8gkxlzhJ22SZYL3ymZ6PtMI8fcdlCw1+J8MaEuzcJJIPGqWcJq2IS731ZKjcD3g
U6Hpm1acNjvxy6Tyo9CuPy9HbEl4SWOjkKkk5I+TNfE1bHkajx+H9wXzFF5upoEF
SVFPjQv5uqboq4MJBwAXLw5FZYhcC5GfFniCEtEzcEawVzThmbvWyX7suY7gw8fe
TRbdgZ1MaUBsaXSQUOz2NmsGkKdAnGsNrLgUDaLraMRllI68lRaf5aXh4ZDBXTmx
1ZVNdj2WCLt3dzrtkXGvq6upgq5A8ccZMqN5OGEl8we/soTcC5zp+7OYBdzjf4V4
3GuXnI0mTO7i89ojx2kOwd8tScR6BQfHIa3biYqu1E/AsOHjO+fKY3BDFIwMYDdv
yKeCGK6Fscht9WklTGo1hHIAprTwnCZOfd/5qXVR6yPK+NGP69IzLpS+U1Dexqbf
8453IAxBV3M+qtpqoTz+WCsBzFWDJgBEvaA/mwMFO0o7s01QfSzjlekxfuyfdGvb
jJOn661xTYiPmjBWLhjvdkCPX4TpZzNGVu329ci2UKl1avJ/evEL/c69vPqPes73
+CimvHm8l5kRDWQ0tyJ+6rui9nXCfIrFKQWTXH5Xr/WkVsRgXiG68IrCstnBvPOy
LDbdtrj7U8oKQcWipyUXx3WPjLLcop8GlWWO/WwW7xhj0Sb3jmrRmoO9BfBfb4nG
ziW+tGD6oEem2/sSXi/OWgb4uM+8Cod6PnaSEC+5DNH8UM/EbVUVtmkAXul40zej
O3o1GI+a2vTgmc05xwfF6AR5I7vmdJdjwO5o3Z2Mv9IJ4q4FWNf2ENlVwcUohBsa
wjGKXn8CjREDYtBEM5LMPUaZhn9BwiSKN1wXCO0uFTRIU49/l5VOqODhrEmsx4vf
wbvAsFuMFFi0J+Gl+wlsG3DvGNB80j9nFvNTcedxOCgxrX/Mt8pJdckCwV1eOWYV
C78LclDc1VkBNUsDjIqgFVWUhKrxVLTqARlw+Ag58ND5kyxADl68l9o6ADoJGyKU
tb8TT5H+YLMdAt0xtxUzqTblOkA09i/vKsfIvyVnB4vUOK86Q4lMcIJ4CyP9C5WR
ZQm6JkJpO3dwhtvnDqRzYuDh7EwxOpbl9wEhPhk7tZp6SZ/ChvsSiFMkY66UfeEM
rAs+sgx61X4z2B23fYmEcPnsOTT0LqdpnBmgJ9jBTmwZlK2m5hwX175k5A+P9jpJ
MC5pSVd9tWC1XmrOCI5u7p2mB7U6RHr8Q2DgouxINSDMwDmdZPnFOb/8/Iwl1nqe
L8AWdCdztmdEPvD/M/FNc42Nnt1q/sHWqJd+D6qPFr2RQ+KZeOre8pEYQ7eYcu38
xGNLO60pDdZORhPEaQi86ZVNVqakvs6Lxg99mXTja33XcZcFXem5bycA6O7ATwDL
X5e1kwXtdHxRfVdbTPxPeKBXFWjCYXDBGJlX/yGHgkyDqsq8sw0SuJAR/yHUUJll
amfYWSZjO8EVW0Qua6oKb03A6zphBM9tn03RU1soKL6PUQvuicSMO+iNvPIROjFD
UQSUkMPQPKY8TVVZgpec0MCDDiOYtLz1Mnp2PsMLOP1faHqpfeVOqrZ2QtHgtWf/
AN6glr8jkwGIP5XozY4PcOwgEnxIZhX5aX/8Vx8duj6VnrVgegglAVYGvo1UWCj5
GHoZ2eiUgjgHlD+IAPLhfWO4C9cXrBM3uQG9fqFMD1LV1wd4pC0aluH0DlubMRo7
ptzDsJXLg8iHu17053EI3jHpCkXLNV4n/Fanfmvi67zNPU/UF/+91Jxw9gX/BqJ4
INU5RBeLGAACqBVzHwpSWpFT1En6j/dhylUzSpNk2HODhfPmqDG6U7fWnCSr/hM6
iMsTfa3JBuNAxNS/Hu4282Z/i/jh/oHzDZsAK7gLyAUcjlVKzPHfN3mMR5522GgP
piXnHYRd7m+7SOfdp8pgk0G2iDIKhta8MVORrQVoHl/D7K+LfxDBN9q7Dn9rFfNO
SxHwCSmclgex6nsLB6DIVRokmoixNRXAI88K5MBTm92mpuszWl1dR8+qtblOYmsV
zZETMG6F/kYOCWysJnfy/fpWrrjiR/9FPTdlEdEiiuNlEx/nUbV7lQEEUHK6r6IC
PgP/Pq8hR/XYMM9vtNrM5W+mraJcGB9DW/zskJTyRNQrZLbyAUJsOD/galWLTu4G
h7W06VapTsW58O8HqQWFRhRPW47nxaA2xHMVBI9jehdJxBr9fyED0nq6nIlLSs6G
XsFcriZ2SdKid/bqpBer9GbvjY+0ozOOdf5NVZ286C+2ef4TyVTvpPGDomq87N49
JnZO89aJMILFHP8vxg5c0K3i1J8LjoMLkQ3dl/Xhkd1kplPz8g8apLDs53TkCG2T
0JVM7Bo/NsnZpF0RsK7LmTy2h9tY9XsAhMD3KulYUQAMSQav5TqWGzrt5SScpOBC
iwh1Hm6cLBxfX4YMmt1gHezqEexIKURlOKkTtMr6xPiH1fDpOHYGWxzrN2b46k54
XofOsdyY+GxS99psR4YTkZh/3gF1Gf/3pK/rCA7WNWVz1N+iQ7KYJNKXTxxXkZB2
66GrSGkA1eSA0XV99k0HUJQ8BIXiT7kac7LUI919GsFvfmnsajQypz9vxaOJLmXl
vdsR9PGdXyARuNga4+pEdLFznTYspIDf6K7IkTEUInSf6J+KkgxyucdyVavWvKOc
LXxY9dajPUO5wKkYKTaZDoNkrRXePVzI4/Fmy6+/9eDIu7TIBrmuW3hj2VgKrK/9
wd/fRizApsQhiHqcdG5LlX2kZIg5tIVP5jEhTQxbxMUFGyIlpjRMz7BLVd4Yw7Bq
0csMPrTHPAx9y+QADKXRzn4+hubfiPOeDl7xYmuq3q2JiT0iFRtZKWvHc7HdyECg
2EVJkeI6FKwZ2QVW4UFBleZJhSyXTpWoBe+lWj8qaGeqEtqle0uT+3BA3J8SC93+
a7H3JrMQz9VsGr2CFgwoSCa7b+q4kRLJDYP36TE42HmOlSWiKdKqAhrTkQtwLs6t
A2f0xB8/HSwPpCbuzf4Ug1JtG/+rc/Lc1cks2izuHfCeBeeYsGQzBuhiIJHOmLYL
YPSSCTs++rJ48XT5T3CCxylbwZvM1ac8keS/Fdgjbzk3NGgRdsazq7ypa/9lqPlX
hWm138G3rbCAsOWme6iFgqB0h7vL/AAWVo9+UOvtOMFrXBJYrW+FI48k5Py9i0NJ
4lr6EXAxGeCXRWalyhxCEKXQHpqxemb5zpevHaybHCigIw0jyzWRkEU6/IncakKV
OLFzcXomy1dJ84zwH5czExl3j8CRwk8gRVx8kNyUD9nmr2YNk+0NpSDeIjMXI/X6
NdMKne6YAv3/fnrqdrIOUy9yUGXzVTauZHhZMk05T3Hkaa2J3yU7nTyUy8EfVttP
DN0R0LMvpdWU9l/dR2N7CHjS1uHHPwzJm8Uy4LwdQJgRVGy5UUsOEsAFKZ4CJkrL
/PvnDmcHWB5wk06r8jRE5a1FbcD9LbcChTfBtQlhOl3SLAgB8sG3L202QP0n3IrL
H6aCkpQRXZxN4ESBsC74vVzTskjL+Kzc6Ng1hTIB17Bw7LQ3M9JgI3n41X2/kfjr
zWWTuWLLrqAMAeAS/CvtAKeOfmVeE8jFuuA/Fr0VzOaJXZzE+be32sCtmiVV/Ggc
aL3zZ3MEy07Jco/k7NGCoIox1wV7obfkEapBt68wp5t6jlpVylbA1S0Osn6S2AV9
Ea6wfHbVU9d0JiRBw0GNVX3HjM/86E8McuL/2cl5CPcQrQRBCHKm0WluYOXlugDa
MjAjWmVi0e5tdZQc1yaNzOyIb0I+d5pGAaErd1QisXjO6kUqY5DkgkRbuTixXEXK
vGV4iVgOdI5Z0Af8jA3taZrVQ42daVjak/LZmTUK0gdcjcs99aUSCmzElKT1v5t5
9+THvUHS0Qvf8VSh4O+50P904mIjDhZIClbHEt4HugUp0bKRynDqaVapqnWMqFGV
wS9bkxP8G9cey2b/qUzxRtNj10zxQnMByO/7sUU9F6Qw063Kbq1XGiSPic9PRqDk
k6gm5t/N79iLRNi2qriIW+9vSIRvHKGg757LTNjRq7k8CljMOQguSkgWwskzamFJ
B4lGb75/0HXZTN4YJALVv99zpL6IGGE5o6CHK5v/rgtINLbXnxaTGRPnVOUqWMwV
F94WA5638i+HJylPvq/MJUZBiM/OavW5nJC6HkdD8UpIfDqt/B1kTcTFZxXD1pbd
jDsl2tMXAnfON35y2r5/831aphn5rfYXehgn20zmOpoekVs3Fr7j8R49syNz3lbX
uXL0cmNSi0VGsM65nkH/EAW5MpHkGuW159Ti/BlACCD3DBf7aIlLlI5YSf9T7UhV
al+bx6/NgVQ0YQQ/x8o4DcXr1oyBc6YgBuyphJWELSUi2A1+pG13d/Q/Rmxcz+Nb
OcRnLEF1wPp0VZdVI2YhLL3lsonOk2rsf5SF2IoNPQhMFjTTzvtpMLpRnEHXB4I6
7OG0IeNh0W0qRhOyKu36RlFFjxdijAsN4ueHmRQXwE5gIo5w25jF9u+VH+a5AoSt
6WvMtFsDu+IreH2phNx6C0XH983NIwMMxlAIYTDCyhIJGadgIMvFweD3YK2HJOfK
xIKKTQI1hfWwh5nzaY0agcK0+CwzqwDmPCEC9GLxZLCi9u+yPU1A21f41dTZu71G
NyNi+kN8l3zaJyLVX0TJWAWRnugF67HgEYtE02N7m7ZNi4In1zHYK+eJeZaCETCY
N93E4FW9t99BLHhUOgOorwFzANJzSQjQTXg2MsLrSuST3OrfpvQazihJsS2BP9KL
ZSQfRmk65BVhCh0FYXHJypYeC5JllGyHUX94WEbMqmfCbxGtbH12ZNszz1kD5bkJ
0gQCSEwGBwCl3SAv4LvKQyi8AB3UMjeO8XroN/17k4SUsLhZjUZ5CIs+4+zWkaxQ
gbhOBLQB8NnDGeFoHwDxkoRiZAv24Zyqc6tzriDTQ53ZVR3MFgt5+suDPIrW9RZe
YHZAS/J7o1pN1FHGq7KE62M2y/W1unGN5v9GKf00pvhCURmM8Lq9U88LPyC6184L
VQw7ikKp4/5B1YGeGxIU3j9Hlbv9lvuOH5fRZQeD6Mfs2cVynnLjVR0C6/pwkiRV
BLvxRtdBSep8fujehtvyfEqW41nC7/CDFZIGdzp0ph/fnJFqhXCYInqigJxu/Avo
B4rKAzTRITjTv/w93s8PE0AQ1Hhh53osGelYiAK47AjPDyh3pnhpAwv4fkgUmJLh
FdQAIn4eKd8bkFYT3fN0OtcfdudJiU5LoGIeZrCxEDWGu89NHitktbKUjyzU7CvD
YpXxCpUQaVa+IK0zi6Y01ovrMvp5/Ysy9FW3bCEeoYZwdo3/I/hQH9bhDaMicSu6
yWwuo7TFUQQM9279IBEDExo3ZhcsN4N1ce0QPmhrEXC3+PDG1lhpaCAoLMUGOYS7
BXna99R99oznMUNtLsyyoGDkzDcnDaNLgC41bkqCcj/G0gOyNiRdmfDL0kj462TG
X3Pzqz6K0nW2KWHfyGDfsUa7MYk+LU9e7l/oB4WFUHBJMyNLrlnQEv4kgr6UOD/x
ut3yI7Jt28qD+tJpqX/eyzupt9kvmuRDssxNmqoEJars5fa5iICrk3kx+e0pgNak
RhyvTrMKAPBuYsRVE9+IlaCEG+toYRMQzg1oI2Ots+fP0IAMNjx+F/rKLdD9YimO
nbfl1rOOC0wdZdj+sNpGK/lmOY//qmtFqdONCCTEFQEFUOf+o95FcogDK3PTJHhz
XwAV28LoZ7KDC3msmzwLVsPzhSxY0XIzizDULNXwbe8Iq1+lXiu3SDWjIkAZQ4Sq
AFc0R5xG1njK/9iXbn2lF/45aJ2FleXJ4mQAe9dqAMKfEMQq1oTFh4zp2OqJMAMA
83xI3IVjVYUyy6RIv5nFw0RFIauS0SB8xKZSZTXHz2jtFFztCNP60P8kLoupYehO
NvTT9jm8TQ3+bxZ7Q6mrMckiCg3ouZ51a4NZsx9w8A3zdsTWJYH5VVudmNjhHPkL
EYRLcbZHFxsqJYVZ7VcHpeJTPcPLxWBgEuVN9abCO5GpCDN9lDx5OldVsf0PJhRb
8+5DgvIRGKKvEXQ9TRjLNCmmsa77BS2yfR+UvI5NeG7zp6bzI275Fp9h4C+Qlhlg
lHUN/FNCcx6sDM7lny5Agvrk8ZD6pO9NKyKIMaxIj5n/8B9+QCAvH3VKKa3MhH9z
zUZ5VewuMLXtWnWMFS7gEYZNHl51b+c7WZMSzVEgNewsXYnMP1Pb4nHYDFojhScj
rVI2us94Fw3t3Oc4LtLwlRcSHiSls4zkwlfp4FpMKsy0qOj8catEhf4k3APbNWoO
O9RjUx9mCzkTs9WzaY25BUH/e63GW17w1pBJDe52qukRFIPli5Pxp7uWs3YZQt5O
rLwerPpLTHqcb9twC+FtmNV1apMVVMvS8OdgiOoaWJXOfxQ+elgKJUdf7N3AtHwR
FTk5G0MPXqGA0KxZT7xrJ4zMRxWgi4Cw7O69t/+m0DGZ7jzPSO937fqp7gGxsgPz
XFMySf90kByUDGx6BkkfCawYkE1rRZTBO8bwYWzwNt9ODPFT5aqGsoFCoHm+j6zo
NSaAjp96o57gnR1dYGV7h942lyMw6X94FHW171e0NfjgjekOBW2pbqBEA55m4KUP
ie5M7DLZiLyS4BKvxTKFZtt8teXsnJC9z86IfwRGNGUz+OlCo90UZJ8qR9lwDTxu
5S5WAXclgtI+Y6hvHFtYqdrGShIr/PZ3K6khDKG3awzBHwNgl66Zgewep7Wzok+4
1J/ZIC/vE+1doYwIupD6d5WGnXUWrpjotoCYSpLq4BcP9JxFED+3IH6Cj38tDb8h
Y0UjZ990XjK/FdXsAJeiGYbUz3ko1+UQJMru/+Fw+86OZ8Zk8FLodsMi7ezsLXJn
T2Zac0OoR4HWAhfi6XS/nVe51V7L8leKD+ujiesXUpZh2G2BCyGbcs3PvV3+T9iV
eKzRDxSbxuI+q2Zj28lRhGBund+tdQjXQHrkiLcHyJ6BfCy7G2p0dd3aaxOFUYNh
CqlJMgyv/zT5excgujSdcbd2vAY1RNwW7DJ5bpw44nNEyJKwDQNj9/MGyIdoO+L4
akSUeDdxU56832nHJ0T7TfybEQXOPCsOfp9+9Kxh5X32YK12cPy0CHxcp+XuOclI
K7tMlajWxHJZTgozhdrFgKR7YWC7qqYycQbhB/7kfYIpBfLNmMw0W+eeIcGB6W2h
oozi4S0ZzB0fEMfpOjWv5MjP1t+gZ6o/zU/EPHXuMTxq3wCVW77hXk/qVsGeBc+Y
YyalN0ywHhCWtPiYVP8geUpv/jVhRHNZnw61hBZziIHI0FY4hWSoB7Lo/q9Iwv1/
4uHXdNplhJ3DUBqtbzRiO3aQQQwzOH/maRx0LkJB2AqKkiJRY5QjBcM3RoTfB8ep
lRmMa6iWI/JbvFKq7hTCXXC+pROA9CxkbBBVxWnjytDAWR3onfnWtYLsyP4sl2ze
QAQsH//2/PgGUxWPfh5qA2Cc8dGCuwTt2MG117OOqfiyFvJEFE346E8ONShkdFnx
72pJyZ7o2iAZ/8QdPPJsBDSqff9ARelLGVzEEQ9ZT1OFZ6S9UI4GQy/G+aPg1swq
1gR0sqGGbs3/HORT+3U+4bIKcd6gtyfVOyN9TRfk6Tcwa47XpLBEXlnZiQgAxJHV
kV9dftf8e9CxCKHf8RCn2Ty3PB/nAGg/Ha+ASY6X4Y8g8XmGLJL310wUxqvLeF/V
B3hOhPvy8CeMhwIbuq/+vFc6PQ9qIqoxZtIryenW8U/R39AG+ox3Ywtyq8KRp9nK
gBOjxxCAC0CTWMj+lelQ8upoENC+cR2lqDyVCaLC7Qz3tGM0Q75zx/vHXyxXqAdO
tua60ss/fDO9h6v1pp6ZB+/COLbK195kiBzvXSDCvNZNfePUfT2LFOvLB+WZn7rl
eqTO7nu1mT9aF3HbHcDnYD8vwQSQgw9SqqKic7kI8tsrENtvO0cjB8FKMsYFo3iO
1RVcWO0hEY+GkX7L6xkVXVm6lowFenE6y4a+HZaoOJ8dzQyFcuoDFvk4uT/ePo9J
7caevQZur1aKXvfDQVLtuV+NJu6Mhaoer3hOWxvw4s0SvuADoXPwintaqtqMgRVN
uAo+2q6s5UISMQSOlIe5nz04cTH2+XPIBv+FocYSepI02j96f70nMgTqudeE53IQ
YZCWris4GiizJ2MkzP3fS7xnXqsXpf76uSQ5VGYkRChmtytrG7jbGktDbjI1ObkY
oLoxR55vRwzEF4k9jFKDiq15ZleEelTYjNPe2DCSuU7GmihdPczmqtBcNrDAuah+
AL0n63WREJNgfXJCQnPgBM45rG1Lu6XnRL77XIugBTDKV0tNEKZf6hAKdkWysT7C
XWE08oE/ehay/VxFY6OoRfw7weDRvQvBlmgxyFnG3pmkuU5hhgQsL2gH9VeBU4bv
MYZnFrtSVX1QPcwAWf1G1hvQgOBdbJ2ulU3iYS2EilzoDRwmGmR2S/lpYPGW3C27
DNbDhrO5lAKsnyvKOJNeQ6UfYrSxC1HCEghuinZV3OXJmDfLawqeQ2yKU/SwvPNZ
VzNrwFLtCjx3nTV6f22opFMMrRVUBGbyHtL1NN9h4SNYPYfbzsORsXqJ895V55nz
N7wqrq8lQQMqF+EFGeOiE+qIEfECpfUUln6TH9FPQRylofUGJkz9PEYbmFdpb49Y
lVPoi+Y9TLBB/K22PYoon0nFCvqnOgHzmDjLxocZ1g0c5rI9XOTsIb7dsuoTniln
hYXwyzOPYO1eUh7BECxu2bFqTjADOGVcIHAjDe8uanU2Kr+ZnhNYoM75uuJ7Fp9A
MC6lxF7p0LZuFcFrRgn70NkP0Ie3CmT86FngYF10L9UcrhYZEl8JK3zt87aaCnvu
EBaqSgxcYa9SOdA9wE3jANESsdd6BuoSsGhrwFeDVDEYPkY0Olxi1O5mR9LJKn3T
Tu48RpZmiX6H7tDPADXjvV+WAR7jcmQC0MfXffw1M1F37oy9KYncIyl66We8B7/l
w3m4l0yFGdwGj8TNzcvODU5Mo+jqz4LNdPaG68JGp+nccZdGNhsnr+ewWV8sQf8f
/R5/RNDG/GUbymedK8fVZzmWOcFojAngG3WK+doOIcWi0GzNM5PeBIGB6KkvrzPz
LIoOFN9WIS5KwYKpLD/B2M5QWDNGB5F3oZYsLxezPFukEGMRZdhRCzu3r6O/4U8l
jakuwRc3qnw3OV9pbhq76StzGIWGp0ZyjlC872qPhquu0TA1xIN4cJ6sjMR29rMs
PRZxV3/s2wD13y/io51doXVr+N9sSI/minD32h4iRfw3JPWyx9PkeHfMYSoJEhgq
mqpVsbBMUdjZS7SBFxK7v3rw/STDXYgz0W6e4sz7hxemDVgFvYPefetRFJUiU7tr
Awe9L2do7LOEBtdzR2T+4zI14b3ohf+4/H4s1kDeveIo0sDvllQfesHWI8KtygQY
CmkJT53V2UwW9gvqB8KJqoJz04SEk2CkqgBOvGHqiJHkVqYEkDysI6VsjPA89sMo
1/VOVY6zLd8DQklsgZBcP9EV+e+XI5d61AKpsnR8+RksgS7uQVcQhKdqCJUnlFOv
F86VwAS5zdocib3FeQNhqtahLJ0NPVuosvfUxcxBkjjD2/YX4ie51muN+4pOHwU1
URtFv4e7702n2N/QJ0C7Rg95z1jgw/Jlj1vYxSSUVYLqOEO1UtJOkDlkQzcapBGs
sKJNf5Q72OeQmflETJNwcuIzEdo8u7Z9zeom/R9ddW5ndM8XpTbXVToiyXbekra9
6EPkf4tyiaEwJH5bXnHSMuZNhIqTTxCWS3LEVRmzix1dzxhvUlR5oZq9ldkEyKMp
mXJEz8mAixjfk8ZfUpgmtAriCtmV+JSvcOWofh80gcbD8Dkzajt0q+NIryEOXdy6
SMw9kuoEXudM0sm6KjONFZPXak0G/Spn/VGdGs64i74qP5IIORAc2Rt5UDZ+JgCL
eMCR7+BsSA6sgjucfJLsNEY8TIzO/mGmUZnWY6s1sS29SOJ264iLqSKzorDkMeZM
DMikorGjd0ztoBvQk+/we5eOyi9eJJClTU+VfkOjgTWHzSPr7WJ9ikJzt8RcXvWC
LjEsL4/BapgI440JYy9U67Vx6r456fW7qE34M9pEaOR57G+NuX+tQ6W7Lrl9Ygn8
Bbl05YmXPQBsEEAEYttqX3EVanpGv9QFvNCS9wXafZNkB5bvWcQ8KUNyYGV3ZWKj
O9vELAJop46wkirukul6X/H9YPoTZYEQBeRqwvZigPfeItCZt83Tptug7XD3Jpf4
kSvPJi82VR1RyjvTGGZoOEEmtetxWhuuZIzIreLUnRzCoUiR3RR1V60fPkM77kqK
/vYpadM22FsfLSWbqAnwE682pxDYSFpiKpW+Qnz0QiOddKMaC3yHG+IJUDlteMnS
HW8VmXVp8aCSlnjLr5yf6W7as9e01+IGxLXwT7MSzW1z0ZrRAftl1Qe/kqY8Kkwz
PLDRh0oV2PILHiLwfW8ZIb7ooVCED2kaeC50/AO8+XGQEqyMu1p7kacir1zryK19
wJj1rz9l95HSWwx3XwFRh721/C0YUCL5kATd1RA+n5c6J8zIfLwp1jgrOZlgjZta
UdA/j6dxF+nSlkGE7WOs6q3QFnmvNt183qxGA6Xx3S1w3GQj8tgyB1wTnfvlkURn
ADkZNdNdmSjS3llThXzsmNoz7zY7AUVBMbs1yQLoaN/enCNlBJVu7YPcfKm/Tynx
j8c6+tNXZT21R30JuxmEhgoRWrYqenzEFCKl1kRso059L0wVMX4SdmcZXmA4c5J2
T7d1kq6VjJ24pwaK+ZAt/+YPolaLi+dq+8tQcmWtuQDm0aoBtBbs9z74J20idQAs
LaPcxMDoj4IfXkedfqJexXAHx64RJKnc70UltjL4PCEGk1ADRcfuGpd3Qx5Rg00W
z4SsU1mvRnuJh0M9jjTz2d4l+A1/4vGBoy3LioBPbttMGnVaN7rzO3EboqUr0NfR
77xzjH+Dvak75+qSiBLtF8y5R3pjX06lb6TipKEY/lVBySP0qbfjjsJ7Cshsph3q
NB5ANSs6miSuFHrHZ7nRqJTqZNz5Txa+604PHM4Tv5nx44yB037kN47mHFhZXQ0V
YBmUOkLZqqS65zVUwF8JEvEwbISXiArckF0+/nF5J84G0dA4KY+EOIaDOlHt69fR
dZo9MNDx9AIg72OgN27+qdYWaeK650u33XdGB79IyHnM2XP26VKdealjwWP2jRKo
3YCPiJGXejJ6yomtgN8iSvbnH6o2/DWQzncKbuKb8+ZIJqZ91ro6YXcBwrjecn74
GwtHynuwyId3tLYLx6yIqI1QPC/FOUWfma5qOU6R8dNXsmcx7I1LT5J1r7UAF57W
sa9ZZ11wiGwzpS5lk2/C4bLwcUxH4xl81irxI1ejOU8qqMFGOZ5ywewWRiyoOYvU
+RfW6DKr2bsz/87dSIwsML53iutAbM0FCCJYIq1o/59yqKYoAXbp9d8mk75SH1xA
pxvOwSiAhHOp+6LohKuo9PeSOLbIDbDmi6PP32pxy8BLpPcMAXyRPBfNDwCqRoEV
W0a7ka6l/c1lZT88vnhPbppPcm/lIz8bLIt1dh/eQnPpb+liT3U5xZnSCz26aE/8
7XVVoSuhjT+JVdGeUt5uypBKMYEtCClT29St6ATCAgVT6vgkM/tjmqM44iblC8z4
qogDoL7S+QkUp1obxOUgNpHtC0dXxQjKEpxC4D6ULDb+PM9Ym+HiwC7JPNGGKpDZ
zj+QeExgdMhdf2nE5MBRFuq8GT+/fcgAKnuASnnpvtBtEaX8xMJ6AqkQbjSRUJUE
N6QmlTrlt0HGTfSlJgjgIXMGNN0mdIhkRhuV8OiTyv83bEAcKOxK8jJp1SW4EH7f
R70sAQkTi6+JAohKySZ65UizTxQrkX7VwEo7VBomCNwlha57mpuj5c00tXfLCMnQ
X7stj48wf4PvB8L4HE+d5DHbQiYL7c3hundTneLl+F1D9LYVRwPLWhCP4j2lWMFP
zYE6IuahIcZzzhCokrEaSIs2gUJJTK7olXw/hQVTyzcR17GTdt10OpM7SkOY9hCS
yb+TP2Di6875SF7iVyzRqSNqpCbt8bbDZ8fM1XU2C1zemUPH37VhFnYUHbGKv+Gt
VmskYzTbLxrHWwZHeXXeYQQc/x77ETuOd+u40FuOeJOMLD5Z6skdgpHl3TnqOj46
RnwmYYpovyFU06Kbq9BN7ArefmzDb4rQ97akyURlfk9emzMQSAXS7DxoAKpK8CRz
i50kIB8lQt0As0LkVCBzGHZG+x8jR4weX7kfHMnbhW3EJlQL9sxD+y8RB3ra1qYY
shS1pA+qZEp/zBKxAOPFk1uhsJqmMqdaajNfJh0dqYjDBu5IymJp5RWOwmPrKnL8
NalisCwbhI1Pq45ZtshSY5fv41y0K8e6dwfdpESAb3rmIJ38FljECztEhA4g+rv+
urYpJvnOGZ3RKnaMEpFC/YUEsahfdJpYeBGSX7NQn2AjZ6NWoss4mbtWgTGUIcb6
ZSSJiVcTRrE/w2aqkYqmEvICnoKhJm8ZtkemLfhFWaFRHdOd0/u4GbhGJZD4MxNs
v06VH6PTpzqYq7SAxWmCvZC7gsPHv11bFjJdcc1xYEF53Go0x4a6lAMn86o0LJML
fQhSatPUCliQKCBAhuXp/vg8H1e4QvJ3z/UIY7pPQb7hqHuQnVyyH+z0Pp7wgIw8
uDfIi3egDpTRrpNa3KKGSo7wnwSloMOH8N+Qj21lcH+1aZk4AJ1iakSc2Jo0ogCg
8JUBd4IuaozZVkV1vlV2/iaocGNib5Uz98lP7WUJDE5WCHFMsJkqUNyLacrKGLJk
xhnsBWA6cNtWXdnPA8t3Z0J7qgPc/fZZN0k9Si94CxHi8vCqoBYXtC7gQNC8ogA1
337nN1xujekqEn2LksXVXc+IL5KCuEQcdcKoe0TeMDbJBO4c8dAft89H4eAj7SPR
08qqVTcx3riXQresMmLWIQoo0x3Lc8LKCW3rFvwHxVK4HkpbpDtIP638UfD0sYzv
+DCHZ020xWZdBEbRxcel1C8MKkzVL2r3NA7vO/xMWkX8oCipxceNFPNk3t+DP17q
kShosf9x1lI+NwC4RXOmHZnawMBMVc4dVfz+yXLH0Aorad/oluEe9BcBomktv0a+
l/rq8+yIypfLPGaTjsDdnDDTW3vqbxr2iFA1hxvzAmSfr1ix1LlPYr0TMxtCQ5AW
Zl9wRZHJEFRMX/7MKuNuaTPUxusS2bxMUBbzKqV598Zgrcp9Au+anbJ5VZnL0t0B
goGBVAmJjebtxi5T7J0PwtneDMWWED71qI2gV9pdnBnRD9bt0nJx/1kzLUeZ3diW
kdVlmMmUuMdwztls+idw+RM9MUDgQ2+8EMO/HhDfIEfoybWBkBl7E2eNj8tJru4N
6xlLl3JPJtn+fA1VogqfNDlNblzlTd4NsoI2Alcr3M7rmQ4nUTUpW1jSl/eEy2lj
BSrZbW6ML5l97/tR7vYcAxIZ6hJn73TQdI5eM56HKjqWpJVxW0GBu55fLo05otoa
+RSJa5SLHiSLyzgoqurtP1ZlhldHDsT8Z3ADHJIj69zGZ4SehNv7Vpqu8ai+XQWP
NQSTrcN7MYcRFpym16g8PggAj3cd0UBWsEoxAVD76sPZTGY2sUZLzE+xWNJuOnhM
3P+fjVNsE5UbmcjvDl4j+CNmdd363SZupon3nEo7mcW4lyAVVKihDv9SKhntH6bz
P2r89TOly9J/ei95uAxoPUK+bpX8RG/KQyGMMZC1o9t4uxaXX6RZDdsi9+iwvZcd
7+J78mkopFrqMtQvpOVsdYWFlu9RYiUrma70TwmfuHpl6QLlfqJqEiO3alzXwrKH
w2f91OsbTNNwnVwVFY+XQpObKD9cUepLqeFhDOUKWAwUUGBP/ZPrSWQaMQntfGD7
vg/8+e58dIb8LXssg7GUGhevBdMDMqsLihWrJVPSOOCn8uCfGlVx8h49eGfb50na
nYjDovRl81wKZ6lVekIigX6U6OySrpkQnL3dE07L4J3JnT30bwvXMP83EZfua3cN
RizHTw3Ie77tTWdWUc6NIk3BiLe81/MuQMUgYeIbo1JpXbV16Z5IeeW2mghzYhB0
9+3/JjUFD8UmzDDZ9IjjPzZlP3Y3UYe1LcZu6inKkTXm/JkpR0Nbh2sxm7NTt2ds
Sxr3gKUkW9dh2X1K+01r/wCFU6DwPmdVp4DDiWA2fsaDJOkwOH01CsS8ODNk8KO/
hMtQWZNOPjmorH7hE/6pzb/nGmTuadoHlkjxS+KLrGoIg1MJFLCS1ibpu6nh+pQ1
2ArSWPmdzbj6ml7EAehKnnQYloLEl6Fmpnkh+peChNFcpb065Cp1ROz1cqns0yv/
9mkGdSlXUGJ9YPcx6YsexHUNwcAg7iAU82gLXRfTJqg0INV+W0kaFTXJEAyAqKDf
B2TCBciZrO2h5wKCPibBb5oFlZJcva0PLNdcTVTWl5alRFzROAgSvsbAdAGAwB+/
62BHX3G19hYAgR5xrWjxWEbs2iwkYZiuIg/L/ucGccovd4/1jwIPkBisKJkGYb9o
zPIovVFuKJAYcd6wjYKLcdWjuyvGedBp56kBJSl5lZC5EhuwoZ2qlSwgPO0SoJpT
7Wl8HfmgVNxrJdKHhp6JLkeRB38vWMTu3ua5aWRRTe6XoQ0/ezZ7DtxaFNq21a8+
3ge2czlubMkbg5+AZ1xCUoDvor66OJ9uU1biIYBQ/BOw9Kr6WPYFiT2MOkL3+l3E
YeegCgUMtJ7ck/e67tA4uZGWLn5l03yi1+LG9Zw6ScMKvfrvSah6b7jDgwW/y4Cy
0J/vXn+W8vkjq3/g1QEJ8F4Ys3NjAbee7Q5XjhJEl2CU+wFliTH9ojS/fowWaGBn
8jvJoRTxVlCIaSedjYTLICGCcvw/OfWa429jE6KolENZqpz8OYolXSbBaBC7x2gH
UNaNePZw+xEUxKJaQVxE8IMKZ1nGSi/5Po1v/0KQXUQ1MCnA24Z+R/Hf8qNS0uBX
ZqjYx6Od6CJUXCLfBjOTzNrUSBoKZcwzlXrd7kPIHpj44lcCZPluJ8w9q1FzTm3Y
jzyrpkADqsJc6RgMbXfeXwMz3jLw0+lUVOfDeGmB9iG7/H9by3goMngbPGzJv6ZA
lVYTVZx9uB4JfDRrAcb3S3RZrQt1TLIL3PIu6/mdFizkF/UWPK52ZtGG+UYrYthb
verEb49w9DvFDkgSx/S2gx9+cOibefiHDahHiYe+HjJ90X89cmWDLcIBzR8GIo9c
slVP/yZneZYihPzj3G9Qt5wUBvOeg0+2dulVWZiQea5/eongFZiYMcharKSxs0j5
+rBGTC9ts+MyE/ybCwiO+RjO8ujLP4u92iTdD8Uq/stmR0BQNPlmkr1q0HE5eWvJ
A52C9kJA1u44uznZ9xi6abGBFt0uxDEWvhoE8xMBQwCmMqI2zz6zgnW6RJ9Wd7+i
hlfbrtmPDaVNRG29+8HWPVawFBdSkdZ/tRjRw0hW9cevVtdVEmuquO63j/JdRDar
dS6nLv5oeWk6AxalF4MNuG7mmKahWcAfSHMrexeterDCbWevuVylaF3k4ixzkcGZ
Guv0Q2HmVhkOYP6y3/WMqJL5PUo8tDg2IQ+P3lBCbGUVSULlJ/wY7AxTwx7ZPxRE
22y+74Y6pvgqLXv+WXCYiWkJRqqbButA0gXP+jiN8j/8aXbIl/sSvnHJNlg28WXB
ZFK5lu1RYY30VYZtNcGGtvDZOEHXt4TRxmwsSPPmWMY6e6G5/cAzy17YG17BzY6s
93ShZiRwXSen8mU0wp8f4j3gruY1Pc2cMOtGEeuL7EXZUAlqFhLIX5ifOLhyhXPX
8LnBd8R8X+61HVmva3whucLJ9PdUgSNmjLdiFoyjCub9psNBWPMlIGZG6uu0NTmO
4Fn2PhOkrM+agQJSnFFdRuXRSRKGpakJs92i5sDDrm9qCM826P7H2PFHUMTWm44o
kuzpmG3VkJVI4p8ZMPZ8lUwalE1oIlr/43Hb7gnNiPoHTiVfE7QRu3mLm/0dyEwN
HaJ1MytR8qGoItznMskPVQ6ppEiF5d58fJUnP+rpfSqcYYmkvAKdYSTlgbqR3CNh
DG6JtgGcHIfO5q9piwCNRkPGx7/oFMqQC3Yqm1J6dS1WCpC/oE0uwCPA1S3/RCCD
rdLrBIhzTbkB4+legI05XzanO4bliOIQmrjlv1xmm9CIIiTBp+CfpgT2PI7Wnqxp
9G8AXNNqTPtpaquttZ30nv36w+b6aUBJRgAME67h8R/my/1V4evgckOZbYa9yH8a
vTTcJo1V+FmsL2OEGv2lA1PC7WIA7W5YPhVsuCOCR6evaGcgmkhTB31A7rp6yyFn
xbiVL7c1+Ntv6JM+sV4pXqexSo4aJgzcHdhnH8oYvxK6dz82Erw2Bw4OzY9oyM/J
9mqcGirPjVqp1SfSca5pc2ROf3Clg1pDle1GfiHNIPaHBHrTF3SQLoXvs4ApwZkJ
e9H82id4iOOI3vo2XzT1mZ80EG6LZWVgdHgIQsVOTg2sB7ozG8dD/Ph7MOrSOdlI
Wpe3E+YfCii3Q9ijXQpX8oisvS3g4UQG/UGNDNw7KNBeOXlw3LGU/H8HQxshSSt3
LyWjitjso7EMYJ5gzT2b9EGzzL4ba9aK3BsK5fBxhP9uT+SY6WigyWLDF6dUvWDs
S85Zhi5rlkC58p6wSUQSkmzgZ06TrT0q5uXNlCrbLzrfkMd4cMH0zZFYncCGH/yH
32M6WvePQzKY4xXhrTpttUpgTwVqcz8s3+sliEC3JLm1iy/3SCgB+foYk88zOI+Y
M2P4BErgBFrAKj6kCsufZXlZjeY280F/OrUZLw24O0qtTk/s5EG1QnP/TyEN+uT0
/B8IzdL/I7LrvHRv8odR8t6+SwKajTiOAEf0fQCwDdaNyuhaN5pE8FWQasD6X6ZZ
9Pi89sv5Xrv8vdZy9L1nsBd+ZuMlNFb4BvzJXCRwv4FRjQt6V7bKWy/4hdYonAZG
JLBuvwKhW1hW9K8sEygOcTP0nlUqNO8MW/knAnPrJoFu2wg/ef6QF2mKg8+p5gkU
GK4ezPXxLqYIyw4+/Igr4/8p+5BEFVt3QTYfupMZzQr6Ij5L3Wg0OirmkW1frpuQ
1Ugc3x83XGt4RwFb4mL54gZ2EzKUrOV04x/cbd3w2LIDQbOsA6dzvLYJMErb8GP5
OwSJAqHU1rT+JgoPUz92rLZu8CWygKHEps3RRdiHcg6n0sFb0qlj55hlvk37pj0b
3QNJQirNdstN3QwUWdiaRJwGCQIC7wQUcMk5CSsybH79yLj6jLCnZZoM9H3FvmhO
v33iCMsCxb+loqoZGysCA8Fd1un9xV5C9YKpPne0GdFlkWmx8SG3r8aPETGW19V9
G+byvPvjbb4uw4oAEbTaC3s+rm50Czd6OK0eapQFSkALufq7eUJxmOMujhSO+PQr
CQAJGycw3qWNt7boXCXbs5IOs/FC5BGyE1c7VpaalCgrCnDC1QQe9laGgd+A49c+
ngSv0oDutXZkdwUa1+fopWUs4btXJzbwHMBY3pDKexk5kXc99Y1NkGbVypWczFnL
mvJdanWd2qEtpfKrRhGmM28PSb+qO2T6tfpc8ivPu7Gc9kKRhbblvxY6CmvfiAzK
dh48n4SMyGKCWcUVDmnxEdYOIeDQNiSeMoT9Sa6O8q2Xm6WQ0Vpu9wszgZxzsTSJ
Q/10nzpxfFrdczWvz7EXSVpCXMPzefokL6PZOwQPHTeeXI211UKSft910SK+XvOO
Rgm+Gol7qpD4aMJBCf8fGwcArIMpPy/K7Xz9dq0IfC3ObGIT/f8LadWojl4mwxCq
B9z5jIJos52Z7xhi4yRbF6qg0U6KxrzOvCxwTbpQ7WALj8qy4P+E2aKEkOTbPhOB
/3VVhqfXwESgRfM+W6DXgj2NC8RntJqATSEkgKfqZ7aEvsYQPbvPkO+b+bXC5dDx
aPRlwJWYDOxWy3DQkoSP1UYUyyL5MPuss9vF0NV4OgnntjbyNj8y6zuavPp8nYPB
66e8jBy6RIvE4lkwZ9mWW+g55IU3o+OEmPSDP3bNhmLuT5EynRM0HRUjldnmdOpl
AhbBTvLVlssSQS4XHW+zYUTHBkQhwBoG3iSmMTmShzo9GCTAZdlHnAo9ZeqeHaOQ
HqiS4DElzHbFZbV4kUmKp4vhEC1iygUig0FXBJGWcZBhnUe9y4Hha/lsITGPJaAW
8Cnud1l1g8JJ05j6GhzjusJ+7li3mWwi1xzmFm4qX6MjVsitcd79qjfCVVjzZrJ9
pdlH41Fvqpz0UQRCL2VL/Qm4cUFHaTbhz8REDeEesYX0FqKfrCOCIZkNEzJqxcW7
oK//bk6cukf/DINMDIpJ10rJySgb9Et0EQJ/taYQX8637bVKO2gpMXZgqBP3yNbW
W6bCnroXgqJFy4Xj3qwYZHPLmOkDGA+4LMDtpwBGcDNXVYIqdeAXGoScfMI2DPR5
Ub5yY3xT6rK/C5uY/zWN1IymSHD/VcS52OJfwXi6wSd3mCA2jIigeA+AzKS4pgUb
0JdzVuNjBzkVhFIMRROdENeiZcVOAI4IZAO1CVpUsRZPcWsi21Vt6qgOvvEiMvar
FfchE0kJQDq3ytdXTVF+ZfyEPrHeKuJ2to4duKjBckd0TI4YiNP2V6mI5GkZA+0C
soAhrSS3mfODSJ72xwkRR0cPTGP4xLcqr/S0wdFcbS95rGDS56bP9ilZR9MbGPE+
z+D6YKEeWNdePQBY8yMyqLx8mcNzIISPF9W1tViuoYH0tLxSweBcbHKnKkwhwk+0
u4P2pqZkDQ7SPFcIcahM9evE/QgjCTrqPFvFbXLoxqnwkXegSACy3WoA1OWsjq1D
6BREOnZCK1KvvxGEllrvUlEGuZXqVCiTWyzb2fF29s751OpqlVNndXnL9SnIUAF3
1EO7wqQfNIgHl9xDKP6fMjHQqSBVx2ez0mVArb8pqMTL/lb/Dwgh+elygqXdmsod
4uTWBWrpLnHafThjwdyWPQLCH+rDFWhJ588/sE6rdPpzvVHxS/8/Vpo93RogTHXx
hXrUNU2grfWUpR0Qe4d2ncudNt2dTdE0D0A0kxrLR0c0DGuCQcr+/hkqVHnKlal7
ocErzVt+HDzq396/S56VWEYbAvsvorHvNxvGXIm8AfvwxMaYT45eApc8Qoi7o/XM
uzvNwXaY6vJPxcTghrW+dnTdYq/QOdnpByyUR7nQShJiypdhzkFu1CKQeXtzb5Uu
X7lWX2KMIXxk83bT9aCP9zBoSGoJUaLB4reC1dOYdgUtsedazfcJX2NNxr9/PBYX
WjteYXXPlr/esdVoWExf5xoFseIWmJsxDS15eWc8Gx2RFvezILN92VnoDhdkCPls
pYu9S3MOUKC3pKluV3qiVQi9KgofF0xXtVvwWw0oMXR1UEWv1rdc5Kl2bW4X6+of
07GgWkc3MwQTpQoZ8krphj8DPzIEUcW08ShE5puDoKDajBwtllR8YLXuiR+E8pzj
Q9MkCSusO8CZDMO9T7GKuiX81fEk90lXWZDz+8TL863MsjU14neq8wx1Ec+an42U
q0SGOMetGFnEnhPEKVAtfVU2NOMKP+UblBahK37nAPB+zSvVMyMLjVP4HzLJ/tXL
kSz7AwJUlXniK31ZYJ413q5Se9/7dl0Vk6tKjiuJYk51eDHz/wgDqr9EPrQiAn4Z
afuGcSiRV8aFl9dw5/E4OUNFf+rrh2KLO3rOOnoL6JbpcX49JVYtmrZDcUUEzOFe
iYY03LcvXCy7lRnE2d18jZo2siglFUtjIkRPK1Ul5PnCxUbK2mT+XuAYgbE19XDy
Vza//uDffihs2e7jIdJq426a11XgtvwOFD9XFsVOIQT1pIxuStbWS4U5v8yY0azl
jGNT/uBdQBKFqICYZVJt4ugnBdnjwrBmgJEKALBMqkXX2gNsygCeRjOt2SOdvZ9t
joaQimOvOfK2trTuv4eTAZcQwqujKIKAhilcrPW72kuvZYogu2Ubf0G5Q7MRlrgZ
a9PuaTliZUpaz01CDG3h5XMF8WidL2Rg9uikH46Rj13QasvRaGfoFdPgHjalR+f7
QWgfSsDXZ6dwenooeWCSq6gL9DgI27E01rN5IIUUT6h/lBrv1HFtk85V7LH7wYu4
9oGVv3aYhboFtxUFum7DwECMnWkLasf0iqLVdmG3XkQZVaaY90WisWhOCpMytAtQ
FxKG1ju2JojvlBFuBBZj3l1rLND4K+Y65LLTprGgHhdJH7MwO7ddz9uCRutiT4rf
mQ9BbX/YLGrUmryYFilvd1pEXgI3WXKDzVj5nxccKl/eb+C20PnAU05RoMdSmzAg
lBlDJaJqgMJ1UOZC/Z9JiJNI9geoipygZUOzdFOx08kcPJBvwdUdeJUNl0HPW4xv
hC2su4oIsmEMtVVmDc8EnKvtV/gGwXHFGNVaCgLXgLoZ6NobZECAnRr6hwTXXxfd
Ve4/LFqjQh5jyX2HJxHqzwI52JVeIYWrra2e6M/hEM71q9+A0VRzdUgn/gk6E8NL
PIF/HCgxZDLdohkf1Cvsgt/DH30lLKjComgEbJlWEjwCuWgnWrnFizaCTBchE1kS
ZHutgGeCpD9etDp4PEf0Idj6Nqqdcnkffts2R0PDz/hBxinaAO2MPukgdcv/y4Xy
bW+iIhJKszL4x9/m22J8USCF0BurK3yKwBHINUioSIGkJ6a4MqXr93R/vbndD9E+
W/82WNp2caaH9ScCozkUcMOJDUePAh80MdnRtxwJb0aKX7s2jcfrLDV4mOqlY90P
aZYypUcNNyIGMJVvPaiDa2Apkc4Hdyvhg54bRTwrarfF+7YA5hFr4w3/V25XRkhr
mLj/byPPOEg36F/uN1bC7X0S2tFlUDvTLKbAUrJp6bEgXfIkpTGGLMN8ecQOJUzL
eu5tsb2EHnioZYoCAIvhuf696L1cLWW+5MZ84vMKO6Wl7i/+x6ZYdXk6VNGasX33
q7u2B8a/KtGP9uXs19XFHJos3aBuMHskLYZkfoDLjzMpwOeCE7ujqz3WD5GaT3pJ
GDFTGoAX6aAx8BIPGP6+olaWtqMyGVEERZad4wWSOpsLpNCmOTl6x+D1JoCQxLdn
E8e16nSfU2nTETqVaYOezF3WLwaNUhSd0mpbw4HBCTWfQNemZcKSxN1+TTGr4Abq
hZHd+8VDfzk3n1AMsakm5AWHA2ra9AnrJOcAEIYdVnsEQWHKIL8MCD74VAC7A+dk
f1BXckRQv8RRLS/gBk/bZU3oO79Vz+rfcPVYQjRIsQPl7gCocXPynO0duIrRULlC
9WR6Jyr8NjCGBi/9ft1SsuLcWwSHRffv52bCgTeOM0dy1xLfP5pRTiGuwuOjxxFB
x0bavRu7yHmHwsHY00wdQv9vr0+Xpyai4xOh+RmobAy+BTqXJT4db1d3j70lS3L0
l+xikcRexZHQmWQcS9/nFkvZLDx29C/vYzA+Kjcacadv99pIOZlwo0Ua/QaVIIV8
I1lywNlFhHJKn6VVzkj9/Rt3azHPwoOTQWK3ph4iHuillPAvkH+xQok19ev0vue9
Om1TiQTEHfYrhiBLW5iyIEquFZ8mmFPYeWPye8J/+BW9A/3lwlmhzHeU7mvp4EPS
8w8dH7rpPsozVlo3k1zoWZKoEkpFSlbJq8n0lic2/hGW8q6BMTNBtfHxwbUC5SKh
E4WMxe1u4eLsD2gTwik/yHozKH/PibVTbc2kkU9zvfvJfFjKSGuwfcROSsYOAdiU
wn08iLuTkYrDjYKwAs615Qsl7QfxFSWEPn2+aCeVpkKH2Hbbv2xBVYJRnGTnQ8RU
ngGO5D2IQGJjaAeuYzb5WUClVncIxI9rQCkX/QqRfD9bE5f1aiWR4KcRnwDTkira
oV5RbIetNKp9uagLZyzV/UQwjIxDjT+6BhRHrkdCq8965S6TpJKkLC3nfEdJPtcP
P8OdmvQlgwLbh3qTy/TrdEOypAM+ZXk9lSi0YE172I+0hZQnLBVIOCThOu6C0WYd
6rbUn1tONXx+PSOZ3w4ezwMnr1ShgNBsm0S41URgKg6YEC9aoqz0JrX3mDMaiz+o
RuqcF+JzTzQe1mTF1dakEiv/jgKO6eB2Ta/l2FRBu8PRA9ek2qi3oG9WyZmZCsZ0
5J8UX2DX2dzQoMIw1HQqR/4HPkRGreSYAe7txX6WSyNFkIOUMOTjFeHqWP0bpeDp
A8b48t+iwdG2Y7pituSz/XwUgz7XQPYA6kAJg+txbo5pCJ2fVsTGJtYNeeXBh5lT
ZuLmmp44Zw2WgqfTKwtx2Wd9yRXDhB05hisHHewImLP7XnguFI/CiatAg8vZuxnF
FvN3GyAezmxeuGkMhcvdumGBHvyXy5q2qYwolBGi+WSltoa/eUwYnEZ3IX6RCB9S
yXI6MRciNpai4Umm0fLBgbpL74LG0pgLvhIOFFUzI9nQOrw0lKEn8SnLlHBjesHz
4NdTwXlydpJQPKAieP1BhR0nayLrIyUjOUNe3LuvJAv1bw8jMXTFU6QI/mILXZp2
ktgIcTKfXPNFLevhbINrWFC3e7Zc4IR2CaZYic1UqiCYOYmQRsYSTkVbuvxii/av
RePTOQdn8gOCOnHoV5RwJnq+ngmDXTIRU54hCW+xbRGs31PeKl7yT/mOJhw60h74
HaY9iOP3u7sQtkWVTmGagjsGdJOLvsLM6WWDNEK42Hd4tHE/coHhQSkv50CLr91+
81hRzxszPJytB4zlEln0SlHwJenQO/RA8xnm0CHGDshyAxEmSov0j/UEhk2GCUDT
YxioZ6FGHfYpwGLJTpKd3P8IIwQHewHkNCTCtY+A5UpfMY55Dt8mhm+mQoxvqJyO
VI9X0o1FZapBmuLwSOjDYbg0wfvtBVng6acMTQ3vSko1QF5Vyll41RJsPASDhpJ6
rzdUlucXfRaHzb8B0FnYOG9ceXqNTeu0pNaTgy46LcYv9ryVXq+kiGzu9hBoeyeA
X5VrzID5JEXR2Nk8Q+aqI5UVGZu13RdpvZLyaNBzDURgBibvhgvBlsTxtn6hvvJ1
+VwdnlmMwCAHL8yQ8zHc9HbEVedR6b3p1WpWj5lh4XGyn+qvHPzWHTatZHh43gvX
tJaN+tiwuRSJKgxUrs3+DlL8Kp64MXhrxeTkRrVBRJKmYIrHUMgJVMF/UKCPa3Ot
4mN/gaWZcVLlDuOIfhLDDhOKMTqzneJzJ0UAoURoxsCgAF0iApodmC1JCHDfltSi
uiU6Iph6Y2yRptLv/nTu9chVhZ2jHM+e4nNru1Vk2swir6VoMaSwEXFOwm4Oauwf
9kC4U3hJkP3YeiQJvInoW6VRhWd9vWf4mp0ivQqy+RLWWt5CoMkNdvHpXNw67NKB
8COPb5mCo3oGC2822u6j1wcmLwmZx+BZIpOff+IYU5YWEQceDCySbNL2ZHTiAp9J
dXJV3oIu6Ada4N9kvjyr66nfJLj/ABdA+6HgwrQuftqDxghRwfe+6Qav6gRNuxXD
hodSOzXLY7ShReIiGNRwBcqxpAYqX2Pj2gGNQomK/xzJAHUtPKHO8wy2pnOJ9YCO
KPJ5PNBlCf1kdGnSdBSp+Fq5IW/vZRWMvntDPdlhmYbJNRlY1GBDYG6h45LfIRij
uJXO8UWxohfGMw45d1pUNCypvrOfRRRKDAVX1budC2WKhj/3ObMLY63rLynU74Xz
rQ+kpMzMNq4cLW4rpAB00O9ww/kxrRbMRKyetS+A5jW9zwAlIhGPn2kF3JjIHm+q
OnPp4Jzixy7D2SPHMEEIoH3tV9B0cHnjMiVebTMp1sgCPgwu5odfQKsaN60C2JtF
MtecfTBnjQCaw0suRC5N+G2X+ochvl+UIqMCvJK52kl9Q80Rms8b8KFaVGjZ708n
MiWELF8csN7CZmpaJKgS4WWBGJtbhZ8mTKYYA4x1t+FkKp4Nnh5CfieEubrgFJ/i
RiUCAekzXfAK7neR8NhjNggf9W1oL667puKgmglGXvW2iGZw6y8qXE+jBUQPHugC
Zqul0G7xVwEx8A35o/jQUIcy5OzIwOhQ6bVYhNdRXk9xlDY92pCekTIATv0JEEQi
5kNshNkzLH23maYT9z1JBz/aXAdnMKPW7GSj/1uPlkowBU0aSzzw9AZy8suPCAnj
s9JLpSc7dprMyaO3pr6lSbY8sYGiNC0zafqn4/q0n1WYsrOD6Qa44XDpm+Zvd9an
KmhIazKx+WBUMBS/wBNgbGSIwLMPin9oJbLJdR0IPodSKDTERq75EB+yTvC/MXb8
edVsV9snRUmV/Nwq9fQveVpIR0JQF5LqN54t8dff85uvGwZcQcVnz8x0SED69Guz
DGNA3gSoEmLFu7qMqWrsFMjQ6T7dsKTHGx70Ukdqmam8fQT/S0gIkVtWTVGGmOf6
+g4f1LfsKdRttdV0C+Zwx5O36tXo4kKOiHNPhorxWrs4KUmPf1HG6LNf1wL7IHc7
PqV9ZW8jKOrmmQJ/lOlEJD4JNAUTDhN+KWbTAyydd+lFyS3VKOrV791MuMVZRe2L
FksE19EFUkAh/BQqpj/D301e5nRml3tqfAjf//WUs9NUC9A/k3VQ+Kq2n4iR5t6+
uhd8Wsdc6Nmn5dqk4IEQBZqH/m+tY9vuwnHwwJ2M9hV6Udplbn7PRt5RMskXzMyF
hd0YaBBBBv0TqKi/nTOP4xzL9SfyVFvP6wmAYNjiIelkZVnqS0nIKQmQylCn42/b
thip4LcOdYlm77xYAAZkMzqBako8U3oIr6NUfi489kF1tweA4Is2Nmwh0g9V8ceT
ChWjU4ubpZu5YuKk0+fb8wmKEqy/XeT6kTedQt+JP7GOZ4KsQ4pdeVds02NKYuug
vXL1GWUz6G6NtKNiHjClbPJNY+M0OlG5TpPPcc3Y8D6/Rpu/KpU2tc7SqVADm117
U/TGERh/s+sPoHvdgl8OWcaX+Bu7de2uTLJgi9Rdgvb9O1N/IkFx2Oo+Zbsd/WPK
a0MZFxV8KRUjDm5Z8y0eBWdqLohk7TVc5iwhB0s1T0eO26rxZJA5hP18qcH0VhLu
J1o7/TD3LCmacicZQ/RiVSXexi/OMikqZEft1XYLDgL+3W9rU56FW/8Zj1i1rqha
yxeqcUr9H63T+FwberamDfUgB/kYltFMwPBF6pCFCax9bakmS7lhTIukto1wrMzX
hH/WgvuCTY82Y4zXrcOzWM8qVPC80nJTTLyH6IS2zhAUsnfIEpRe3mgUpkvtI3SG
rnVIGN0r4d3jBPR9w4CE3fx7ciDNxcG46jwF7McU/PqpKxpjvAkAtlFdt5Dl3eGi
7sh8hQd0XGl734tTaI6bHFO5H0rLEM8gEZHykUhTWZ99ItaNeKYOW8kIDFRKTtac
gmXzI7gQOwDhxeiKjwVRdCA7Ojx1EXClUIf3lKssqg4pQK8F4/RSP1pFbahl3mB9
Ay5QNfAQCaOQ0zRfWI4QROCRbhld37cI0B1jxqCC6zb8VIcq9xTy22gTQrfR5e6T
lVCS4hJkA9g+/rMBCNHZq3VbK73yokrx4xugG7lcLkY9ekh4FfCP+k8Z/e5sIBVh
gKs1Cmc/MCNbd+0nSfFKiJDbAoGD6kFiHR3Ay9kOceuA3PwH7xZOm6wN801aPvtl
fhkHSfpB7vKiL6Vq8qf6V/KCLkGnSgGlvSmdaPi1hSVhqQ1Qu9j1BJv/+EK3WwDA
/k3+Jy7eKNUme6ok2vDvM4IEks2NxTyKgOAHs/GRoW+eOsUQiYZodVagHq+hOgfL
iEoVGGYkdfnGguqLmhdZU1QsKMlYeMKvoxYPKocQuu8BWpxdDcsNy8lMUHelei/f
MMEsNPMJ60qewD/9Ef78TC+2gdd2JsK3BkEL74pQVaoGW/Z6nJYGTnoOoMTUhIt9
d5NjgMtwDCaDBR4/SwBFiVXD+DpI7kVvTbp0BqM4hfOiqHeKmJx5B0B93Y1a7akH
rkwOG3ubuxBhixvE8PnzH3rt7yD7QuHYC1Xm0yFojriwK+tQCJDnUZHKX1gKoKqn
QkSUHggyuKfNsCga9yPP1Nvc3n5RHuoujOJXE0Os72RrYBe9kS7RHn/ccsQ2UquS
DEgssNJpm4u9TosNoqK9aO81YFl1/frj0uxU1NzIVlFaTah6eG/g2zn7LzJoa+8u
5mIobKpdRKKhJvna8Qr8+ZLD9kavSseEEKxQmk2NYwm0+8kwEpbk/ZTMXGxxgaJe
uK84VVOWfUS+0rPuXbxseUJHt5WIr1zdgbb9e3TDF897rmMdobz3tpfP6MYR9KaO
kUdhZT/X30l/ETILnZZmmQwrKv2+JOp3fbZxA8SjxjWw5Fr7mssIQrdVeJwwDTKB
poWr9g+4H9hhfWyK1o/BYoce7mASVUjaw7eaMcIOJqoiPaco6/64cdmi/Y1sXGGk
r6oenqhN2GMopWLPtyUciWj24DhwNJkLs3P5HhjgM5mTVjRlFhrka7hHo0nZrd+W
GeGOa+OBRQ/IJy+773sSyXtEkeRxc+hlM0S7Dns5S9ezmNG0CiysPT+VunH4uhxE
Dy7lWNK6n/3EaQ5o6rVRetwKQd+vzeZ6ckXtQK71IUJ+yldNRGN822c46SUGFyqk
8BafGNVwEsQNHyL9M/ukFauWGvTrjlxFuiGlYF9Zg/m+Kr14MA0qLhDtrLztci8s
3UXEw8BLfbPkntRNB5SqZBGv3KO1XxfYYz2Gvr9KyXFbpjIbap/QKm1HfJiJJR4+
58C1nRJa3aNRxudox526A7Fzgv6SiNiV/0K4rogvMvhCwaW74ctYeb6Jzn2S6elI
9jg3lxTZnl++EkrCNkSqo39mX2RIxwPXxlA49WSk8n2YSxKWaWgPoSeNMELGf5cw
IZmfFFHuz08UWrO6DnNkFK1uLkXgJJb3I9c2MPugCFJk5FgSXEwTHFP5OEEqu2mQ
h1lTbYuFqP43KRJNAhfJtwXZ2qlYpXJ6NXHmDoHCHRMjhRgEs5WhAJyNA7JV6s3l
63udnYJ9d2J4cW1A5vx4hTArmPxnK1kJvHCBAsZBd/oRbFRklEV80HS3fDGRQmtX
w8wmW3xrFS97M2al0Z5LTy7BSCzQ1EOEDtTbxO0f3XmgoKqyuXPyWGr3zFo4kk4d
w3yUFhuwKbW18UCs8gebfikDw3XO9cYqt1Nh0IcWj7FA4BDdofLIitTjHo6ToCz+
MAZP++7w8HMv+wYvhJPEIg33E7Jt2hfx4rbldrUQUg0vVBz1hrUu8LVkVmCn2AlN
+ySw6X69vRypRq5Hox559XKU9vMhWYAUOPJCEtjmdW4+07Y/5oHyM8n0p8fwjFzj
mvrllwIVpnEQdN3PiM8PltZc5wk+6lojDnlp5n9nb3aOm2Qf0SLVdijUbDAgOmLF
FmMUAJ4TsRlB+qVEcqD9hRzdw4LcEw7DaffiWMQcKWoIPeicCEOhaw6Gq5wi3z4o
B4CuMnhjO28+ulENnqgGUwKJEoAaacJLjt6s5WF0BteaPwJVY3vIIz+D969OqjnE
zJFnSedupDDCo8TpuRGyX0vytEX+7wizQn1roTFxJUB/tqagJDclt+P0WIjzcvmn
ujIEWOvaqNa4qQdQwIdpjPOYNKdtjn0qqe4gjUjkV6I8CqsDM9bRTW4Kzq2uP5gu
MCtWMkKT5OyxjKv7DIIwmUavfIPuJR9cPLY/qnxAP2OxTCXRLfsKBjqkrApJbRvH
eXR29XcegXAii0iKJRDzO4XUvX7P0CPoJAPJv+EgbX0+DK6Z/+1AP0ea2hyO0NAQ
guWAnpLiqLSLWEoUv3sAXv1pat3EX1hcKAOuPlBynmG/s/wTMfyAtcX+pkoVUede
Ty7mzbR6YKhtNiaw5H1cXNWxBOckTID4t99b1j5oKU7hbaDOEQyKBMze1b1Q975j
7VBst1cZqhwIDUcIYCzpGwSTmD/scfs8/w9ja/AesYRISqfct+cY0wrSHapkfO1H
eMofybquz12LtgD8bVfE0/ioDVErvljjw+DVMV8Ozwhp8DUIAZtM8PghECxqRYZY
4mKP0c5V2SNsCxdrZO2myZKXg2xVisgTLlI7F8gVrsgSSz/8pKwdDevp+9zCf/JZ
kUphy+KLroX2ENqpflDV0Np4EmwBqMCGOSy+E3pWhrjAYjshPGcB1d0tJsApumJ4
vI0kQXlUuvKwynLwAyqBoPf667tLLmdNKulQuyjr2Oz0h8TEY6be4dXPenin+VuG
ey4pZsmze/PNfpY9aza4VDUsx9SRjmmfFRzYJYkJ4uhXwLg4LFrZUywESyIICVKo
46uitXW0QgiaR4ybH2eROREhEYmku/ljg4+F5xJqGcyFdm4FysCPKkumUdG8e6qq
myir+uT+eY3kNMJnbinWflzZrJwkG5KTlVNcNVTIE9ClzcUjFiZS+de5qTwEgf9W
u7veykeB52BTusMiIfnU+aGFX1y2l2FeR9/1dDPrqlKMkU6pLaFG0I8M54Kl7Goa
BUMQCYW/L9AhpLs00GbioWiJq+eH3+QAcZAIk+zLfFOnnWQ4wD3OBZQqpynNcOrE
Tvm56IhbF/qGsH+ywU4f5eL7OBWZC1TKXns4BUGCpGw8+Snc/TlkrAlpxNseHICP
MNl7RU3KFFwnB71XGJ/jyc78R2fKt1X56LjSz7DlvJi2WiopUiXCaatxnBWw4WYI
Cymur1FlgYJkw62p9U5tiFrEKIzvwE1CDp0GVGmaoBgZ7XdZx5DZvpeFtLuUQQxs
iiIg1iqohl96+KnBYxO/GKRzmhjyIa8nkStw9UpMaioWllcA9ERZssc+zCtOTG3i
AlynzPpZAKFKolNnO0fXKSSkd5+VaW5JGeTk6n9ldrL0BenLNh+iJn7mZzDwHCNM
NyN29mcyQlMxk/bdQvDW1RwhYOQyDjapmoqvKuL/F8B1GvhX46eBxs3dJxW0Vr7V
LEO3PaaK9tZCJqtG+blWWO1PSAZWTXDxpg5aLZIsAPOfVL4tFA5w6MQKA2DtQpfI
rpOaIwwXkWuSxYHnV6uTNmgTQuvCPPuUcgVNAqTB3YxQr0nyXgeirBraDCmF0uMM
VWHg/+ZD1XoGzZGlvBUu5qOBe/UnQ6GH4JjXGWujTtYwV9/HZQn0rPQl9r9+OPv0
p5sYL+w/gKoqy3Sg9NOu/N0FtUn4Mgiu+IqwBGxFYwBs3I8J9sLZL6e7bPNZYN53
V6ObnmAAqyWaPXQeWIa3sa08QkPlrP3ALXPxPa2Xf2EbAzo1GABoVKclqbTcMD4U
KFY6V7ZBtu1PiWSwZ9Loe/S/0huEE8sPcZFaDtuagnsTxYRvvzJ0f06LebUNY53G
Jaj12verq2Sk7hk4U/J1Wzi6x3XGjPqz0Uy2mexuC9yXzACLCh6XU3eF0fZcfJPM
MIsyL+Wyty7JIb7ia2asjN39fE0NhAgL7oxikUvlqEo/gJMBp76HVTZc3bWaEKFw
c/tKVnRSz4PhQ5kVHJObsDr3snKFT3B5hR1fxgSMSVvT0LV2492EFjZYdgIkdakR
MWjEGIKFkuxlTGEjGa5GVt5tlb70tb0hllM6kHiJCbWTuWaP+sgVs8UNuF7b/HA6
UYDA2QfuIItuXsQMCWbd2Pyq8g1CXWjmTDXSnCY3HIzAVdhE7W7PydmD7rtdidIf
ttlNRULGmAxb96ExJYbT/aLug0sKk+bN0NHDkRO26J93XyZL4+H9lh2WDX0M7i5t
E1yvAQpUHQJOJVlkGL88SYoHFM1kPeLfY2+6Gy+xs2J2xHn5LwuOGRuUk8PDxeYI
Vo+hkS3ruigdbezl3mZIeTu2iYIibfflD4rBv3j8RXGITB8hueDGHh2KZfhFdw9A
WZ6ZieY6oxjBhi/Josg2b1T04sOCl7NAJmZ+JLbKlKxwOwig1O1PTfI09UeIt88w
5i9p3X8OJiwzf23KnSky0Mz7vOvQulVqOP4j84iXoDoSN6Ji8MVGtii2u9RcITHv
o8SqCDQJh4WKxerSuMHU+5y8al9KkB6FcpoXotafpdNrxtH5DVw595Gh5aB8+STt
Bavq4y2ycm0n05IdBUZ2+mGY5jYZa5ya6xnOhivaMSlzwSQk4OJuLNNCxRFYmtsJ
yE1in7/Rs5yumQTjF1YTpk9IEFS+VlPWCTu+uqB3x2t6OoeBPIoeThFu0NlhSZph
eq62WBVKwiOw2/y6Y/hwz0MBc302SAOGPfp+cLBtDThurb80TH6oW9GEZGmZ384R
ApY1tkGAV6ejyta++mhBTSJ85Wxhz/XmoaNvv3P3Mki1aVV8tkZHQeLu7U8sLCP3
+wCDJJ80odMnCuacxwkDQotu6bON92/ntKIUcyLdaYkIzyMRmxBVTtHIEqAZZFRD
lFqAFx8DVe6Ud0qtdtu9/ZSQSF3UA/BoccSCq/3k2CO2Repj6nt0w98C4gAnVWUi
pRImJKAN0QDivYclkTF2KZUevO0WGJ7Bakd3kihVgIFDHcLSa6YNysK8RYV7KSmp
zP+fmp3diMy30xeYjvn0GSlzsD5+ZtEN9b8wd3NK96Ed4ZXm0z7C/6sAMvr9/Enp
vINbOFCpWfDfy+o9EpVvCCyIUhKFGO4Gnih4uXurXjhuft+FR8Z6WteOJyhEvUXk
fdnVnAKhyu5VHhQr2YBtbM+0H140n6RavW2dDBrSg/W6TipClxXXEdzwHo+AMvIt
8iedQhwPxCdRUK2z8lrm8se7J3Vt4uMLbvg6iPnEag6/5P7pGo5Gz748PkeBGT08
IWyhfI5xmjAeVKDfgKwBhUviOwGOdAPL0YVWEJ635L26k9SRPtLBF53i3/w9Pa+u
82xD+JLUhPAw5afkgSRgp9zifktxNXBqqmG981/mSEubm1cYzGYaahOatBqj2+4p
c8gkX8kDV1vvIoA1BZfZF+8dJm7DjhBUWEvs4O3tSPwABg5jDggc5CEI1JNY5CGX
FTI9235LjSUcj4ocn1OWaYyTdSrndlgB61bfGwrP7WrGrIe7hrX+z/PFp90AJ14o
GRObbUlm4zr8HMzqJmZH/JvKGn+hl2Cb3jZQ0zODf0ZqZ/mR3KUm9+cGT0z+0jqf
k8Q6nBSTqCHERS3DVeq+NHWYuR2ProQzpltukF5S6N0/M+3NcdtRx68wm3SEoXQ9
blt+mZ6I+D+WM7demb98izDebPsIypazJYrkxo0YhofXNrxm/DXXBvVOyEfEhLJ/
aghRxTnnOhlb2c4wTJeaSyXnjr7i/i/3HK8uS15L78RptTKbw6UtlLyuQ7ko8WQa
GCdmuIE9NmZ/R13ZWR3iy019uaXP9LQeBsJbp5OOCYcMSrVUR196hjDFvj0lb0no
KR8YXJobhAIRouf+AGxl6RKiyaSxHniOODcVxdWpVGdtQqrPY6xiOWGhsd0Oxe7+
SETQRC2m2YPyK6mnhSpQlARuP7jKLANbqsixLUBaG82hWSMiA0jYr2Bzqy6NkIHG
OX/vcdRiYRIBwadMztnPyfmibUZ3IyNzIqxRb1wOo6bfSH2bOzyQuibzL2ECqjx5
AHLlPc5C3JTssxNrisZTmIrderUOQYeP9v7axxJF9uQqZuXYsEsVRZg1fGfNCSvU
QGySK6FYclVQzyFjHrgq3gna+4GVj1nsNzI4TbFG9zdvT+hGUs/cQAcO4jVOLj3N
HNEJAnxiOIJGAtoO0g1lCRzKscTJdl99ZPlWQ0nT2x/749pJMxtK4RJX+GxMuhKq
jxzJlYLejdSd0O4VXVXBAgrT83KGwhNMjup01ljToRWYJIyoa/VJ06yPfebHSEIy
n8HDU7icrG53JzRtFSASR5OPsIzikVf91UQ3kZiIBoL2XgOO9kqgQ/aDGesxyozc
QO4KdfjcMtquSQTPDTSPnLDeP8sg0Ied5BIkDt+kSmBgj3FCU3Km2U6dunrz7P7B
hTE6hQFd9+D6I/HiYiN+XKBDEgLCDTN3VI9pAPG8Ffx494iZeJDrPokRBix59HA1
wmHjXvGu5g7KZm9gpi6eJZrzIN4juIPLo2O1mOG+3hzHJAJ6hodUsdY36HFxNL0y
sUzqvRdXu2P3Y0BFoxG9zam4BwLMUNv/QXti7lY7uCXmdioCNt4BiJouXz/oNMqr
2JVOR5dUm9Vhj7wgiqgsc4CsLdq8fS2391SyM/iLeuGNm54OP9UV1Vqj+sOJneRf
e2iiRa2+AcImMlyS74EybP6iHAjBuBI/TPXy/lVJJayxRh9HjtZruvbcup7NN2Dm
yirMS63EG+K6E20vr60BoLHJ3I+NpqkVaTZbFTKqUtbqtlwFgaVIRw5sbQpYOavu
51wI1cTOBOzwLoXsVzRScBDjcioR3G8tJIUkSfiFJz640JCxgt+Rlk6y8rVunXmF
r9DN8vBoQDpBuYNuT+LS0W9Jk5U7JngyKAS1IfoTepBiRmlbvnFlBtAhpuKJDvVn
d1IlAp2Quzpk+XsKFJeUnEx7u6bNFUnR6hwoz//2LhpuZt9uEb5aQwcs6ppoXbcN
ZzyR+cBDp16Ze+yFidV8O+qMr/W9KLDiwh/z8HN1D35X+6hvcY8vHrsxIZLGpUT+
8smKnt0vKkdyRpDzQDihOZ762AUHtXCWHjNZsczinXQxXFICreGDAWBs3eFO8fBI
+gYqrxDwyDkT0l7+rJqj8Q12sG72srQCrZq1qfMsigluXAa3zmEnq12Es1x6PomR
s1Cx8OegW44urGSG6Z849XJmd+36VaCCHTz8+hWIq5m+hPSoztPGQPxZI16yVURS
m6WBWxDs52DrET35tJX54SofkFqnSahzwl1af8Ydc06rcI40cmpxEq9onBGu0d5c
JxQxZYGdmie3b8l4uQ5yVVuO2JPk1Nl7iIycTKCtnb3btvDik/tgS9fskqn7yevo
qZ8O1zJl7MEeHGoBf5H3lgu/xnyhEkzQC8YyxMjch1QldBAeq/Df9XvbBnWglrya
cy1EUbHifs6L1fAClGVCkjeO7LGI7O1CfWIAeVZaUVXV+xHcFuh9hGqsoyQtUNEa
swaQkNbuwUCOVa+dGLh4REjYdx5YOexKPd4ZsR3DvR0AhHkDJJ3ZlKjHu7IDvtia
rw3PZLNN/Lm4O1cQPTIWj10RFPpe2rSX0d0c99h4/OZ8CxjfRir/t6byYfRtXw3L
RK9tnXrQ8t+W6MS7eLYJuy3u/SZPtsEFM8MH19jrrKeF6o0rUhz7tN47vtnWdIMD
6mFi2ngSwB8/kEhs6hSzRy3v2qmrVotdX51q4jowMRqevD5wvbzcBZAtkZABB79h
ruIkGf0DaONg1H60oNR43qD3dFBj5ry9tvm6N34/u5P/u7D0HtkTwvXn09aVlxMX
wJdYi5n0MZrR0Ho1f7quLTETy5t09+skY2jLFeWjQPRMDh+g/epSxjgxs9rRQAFG
PzcQLSPlJpAqImzmRQxzb1k2dbhrfwOZOEyY1O7jF9dqgZHY6lxc7SQqZMn2eoEU
syF21YBwBRE+QG9VoValWqRGBWPVkY5zl+3uRI1VsXXwovVTsA4YB+BGNMOFz3Fw
3JK/JD5R9JD4b4BhzGycOOkp6pOqwQ+goM6kV2yr2W6r3KXLuWPID7h/Yuo0QwkC
TcHdVrwKLRUmiSTblg/UngtenScZ13PthB4vxQC41LLkPFMxfYmaMqEmt/Tegjym
Tu1fdIp8KFM1KpggqXy3GqGebmssfsRE171+U/iHBKwz7Pg8N83Fswo9mLxwR/Q5
0QpE1Lkx4iRsToPYXWrOrqfFz1JPLK4Gt1Ht7k+AV3zk0qTANL8DkoAPqM3TfDqb
Dc0/LuKcPVC9M6MLyJtTfm8rq3qi77H3owaNFLRmORpA345LfN3UazueAP0fDJkE
yDh19RwTp+OKyORelQPjjFzCJyzh9syiS0nPdoMwubG4zsBsJeufV+ErBCB74MwX
CJLAeZ2yhzxkPD+qzpI1Qgx3NXuvUEemeDWWQ2+Kjf/bWsdYzu9O5nfUCAnHLL9d
J49EjXbr710oDZXRhPRv2VntTCCLBXPhhLokpX/K4cw9lOeg8Qp9dl56OBlZY9tk
SRWG+U3zkbwZLWJVK+IdtQr4TW7Zl68mug3AAGtV0oRTVl6ENkNwL9rqwhrKrVYA
YD8yOanqCldy8TEgihPkKbVtJs1Z9O9hHd+Opp9kzwdWbE00potgKGYD1Xu2dwvS
TTpKAiEpXbRvqXqKlSqLw6pVvTL92POaIArnT+VTCcLubcb71TMlEXA2BGmVa66A
YleO4EXym7xmLzHpLcajNWYuleciE4CV35gYa8+1qWizXrgsMkPr66NnHE0ZKhiB
tyE+iIYraU801GgTwhanGJpge6D5fQ8DDug4f4CtVxoVg0PRxVpydTmbxP/mc6pM
dDqbg3a7dnIdYPWgcC3F07hlPyGJxH7D07xT+Cvy+dNnuGoz4aH00MWJh9jbTgYQ
NQZ/szh0eOpCWzglToI7uBXG12oGjQ7mqQzkdQrCk9xIcdegBrcCIIPHOe0UF/3A
iFBpzYu5IZgKza03F5ArYbv22TWFS+0IT0CdZUzrsGh/vUejQuMfi/iLOmrNBgdj
pgvuShy8IrsVMEgzFBHXDAh8kzMBfgC6kl+yWqC7oV+BDOS/uVqj1T8d+RHK3SMm
3eLLNXyzXYafhLA4xeCNSH9zptBs6Q+1F3W4so/R6ILj+lrrnSnuPo9g5etVA2Hu
uA4a6DyTmkE2tZ4mQ69IknbdrzM5WS6lrffdSi4OF5GLSBmbFa4L2HBDBdOdTHFo
xzu+58GiZwR2w714GDS+hZDnqQPciX+ztGDkmZ0JI480760ZQfctKUIF660nyjqr
eXh38IZsJlhHZ1/5r3EFDQ6uXnsmIEW0wKfUOl7EYcJdcZxK1g5Pdi9I8TJf8JSo
Fvx/6iBF37KSitPbdoC6lJhzkCQkntQdeGQy8OOUgZuyYbreEA5K3TTPzR2TpPxx
TVl/nPTufpvmD6impwMUjQeOcAD91/520Cbtx61grwf/bjbSfFEJZtxvbd5dgfvh
u3XNNG89cuWiyUv6ZYF3ptCBjD8RrEufzjc17eRl1RuVgy5+SA584ri9chcuXo02
5sjTfM8TX8ynlptzLVDRHz1FR6plR5ixw5Oa5oB9LXhdYW0G6Zf3XQgZ+Xnx3P2e
oLo8AEkMlR0+BmAhFcSvrn2H5ojJAd1fA95eiQ8krdCqlBpjR2ha4OtSKmRz7N5D
OKratK7rRzZuhPABbbcwUN2qHhubx1ySyXhf1x/mnzV43umAGzcppzV+NmxJ1QcO
Vs7fQGHf6NOoNfy36iirzdiIw8Epwd2/uCqIDDA2pP8glR2jak/74qLnpVxZBAuo
gZEhbmKmAa2JgJLnfoGzXud+NHkQ3thmAX0UH/KTxrFkBoBnLRiG5oJe4KzGkn2E
RBHIkxfyze1kqQUau5IHMr9dD1FZ9H9TpmK/vrNX2Y/LWSqfAhjovHBqmgUOs0dB
Q8825/WPwtO4FXxH9i3JBeY2uqU/W86UcfrtMaxFkoc/EczNSy070pB+luhNdeeH
JToMlzwmStyNwQe0XoT16aWz9AyPzeDSlFWd02Z06xfrPHDb/nzQn60suA+RCwz9
fyI5FqAPbmVEEp7Rts6gG6coX75PuMkiUhXIxIXfilECT132Bt7/HykjGRX01NRG
ATHdcc5WnDWPvYbkHjeMIYrlUwbuYycnSweQp4czZM/AFLED0tqVE1XlhNcgznL4
t0T/3QPoNWe60MbsKzcdXagfRGASLiJT6pLuh267MNFHjd6p3PYnAwT/2WTMCZTK
4w4YT0adYRx+Tz0aYvJXs3tZ4RtGb4whNgRKNWbSYtYGaUAunr47piAPxKqmnOPv
HmsB7Ki+o36CvgVpbKeBdCSDLt1UwPXh9EOz5c3898/3BVbVtqLR/L92euUONR0v
8T/jAvI1/pPu7a22Hh0rbHcIZRcq//B1hpeR7oU984mINTPAmlf/klxyysikIEv1
O+PaU07mdOyX9LCkrRoF8Fp2tob5YY9cELu/EAVGt0LuKrzrw8kaJeg5/kLaWCnN
MIFphvg8OprhO9f4jFozPmdMTz3Hz+KYsZFWJm8Gakpy1p39sUuII+E+ZmHH9h9F
y420iUiXswOjVVCttG0GlFvFRnluazHQ9k0zpZqvuFQhZf5muV1U2vOviEMqpm+O
JC9cbzio4Q7KKjVqQ4bzhO+mnSMPOalYjaWZOMUyrE4tDXpc5shf4Ht0Jdrway35
29a8Obmi8WV1wC98Bzim/loFu+Bd6TUgjURU5I9+jhBmOh6A+wEwBcsL5U543Bbd
CE1kldsgvebKcAhL4eAnTggwTp0PZFPKC/1G1vMGameciK1Eua3KGQONFep9QIGp
2uXaq7cHwBdAAFUf1a0wMKFWlrpT8S5ZTm7rWSA0Q2OQq+l/wUqJBZamXf7ymFAF
wD4KfB1lqMU5k9YOEebl8vE6ErbvLUK8TgUyp6uM36KpDufqaOYqwkKQ0iQ5kd6y
YLTSpAcN1PktFjJSQOwDJXfgN/8vScwvHO6KnWVMBqK3R6cMHn0JhK5sGckVwykx
Ag9O3dWKsRlU31ZNdJX1j/CsmORj97Dsr/vVMYrOLyoZ+OQm2JDbap4q29h9XQDZ
wu8dPCBYMdVJ+EBjGKbAtA3g/SJQeTU/XcUxBSHi3KDLeB/ENVHnfhBO+9qNBUlx
WFHEZOli4NXa3b08vTCOaCAchqGJdn1le4G18oeqptGOTYZQA/NjCnHZVo3bcoSs
a/E5JceJKwrPRbgITIuAW/zHGGiATS17zX6BFOgzv3mXE9EJnCh8JNlHszJP2PJa
cRCpM77pkUgLc652a0e5+6eqUergZjtcDs5RbuNpWFo/K5VUrUyfRUT0SPCze9N8
HFIJiMJogRvACVrQUU2BU1N1zkup4rVn8sNGUILLuwdZpxAo4D9kcq9/kdcjQlKq
ICBv++EU3vObMxwX4kjZHLBx7p2dvY1WseaaL8Ojk5+rAPKk9jVgcP16+24B5rKF
ku2KRDnDPUl0tlCwjFiUeIPBMPkW5fmfWZfF8+zrrxa/K/KwWXXqTXBYAscpFUp9
fdvUEqrwgstASwOGuW5VLMxMF/D9sWQowNaKHbkLakiDbqBV/BNFEp5Wn1I+dj3A
QBOJCZKMs5h2CkJZPDGmt+O3iROs3Jz+/YcJ/7Xlqfz3g41mOQ2kI4fDdKYryCwD
z0wjDaaxck1FIRpsDNn3TrUQvCN1cv+GveLifDXegVI8vaSv4huHfxCOI+JneKxq
sqRzTNouqYhlc8rM7/akLDRrH7inXWHNX+wn67HnQgxE19wDYTV1k8BbQcr+Xk86
uvxxmEqv0yfEb3KvrdmyuO5rJxUt00pENB7L5j+7yfPZ9S+5SuH1PG24OstQf2yy
wOSFRYJQZy02N6B1SdE0V3Ly4eZvZD35I3R5pFyteblSw1rCNVjDqfNKD5IT0bLp
5eaURfxGHc9ZqhFrK21N8ThKdbVzWiWXnV4yvWb1/Hdb5ijz7JAfohwiWKh9ICav
sHi+fvu6WbvXeyvcp0znXVnXlHI7ektPJEWvcoZJHK2aXBgiYdIWrhKkflHwwsLo
JeD3gwTNusPhAbNY55ikPDrFijyinrZTGkYe7vA6hXvteRxHrJmiR3Pj6l4p5Qte
awyK6mOgy9kwFXb+qlZQE4hVBod2xZBIidPua6AGpwvLqtRyYoQQbEVqjntNAg4y
79ucBVaMm9j2KjKtL8To8vEGaJrUnX9K7RLbufnA2vGbhmDSa89VafAPdzZGMOxk
WZxQO8tGhjDiKje4AbZlgzn8lq6VV8f6ahBgwkpv2RmQ0lZUGjtzAYI1/f0+3ljg
jWzNc/VK0gwoYEwtvAn9SRkRKz7qSu4QVobOg1cAEU7hZ+T4b0VyXolu6nioLds0
1xEX/Pnhw+DFhBaxUzNr7DozNvdvvkYDOdi60EK5huoNbK8+G/VWh3CKg7uJ45lb
wXOw2XYGd3Y9olnTQX4VPh9xklbj6phg9u7Ai2OBXt7nwqxCRFgLCurkosMFBuXq
IkE6GSdy1ovcvWgKGF9XoeQMJNtxaSPxE2CDaY68UoMnOEjm2/9+V+NY235snP6b
RpvoruvrvR+9BD4gPZ63GPLWy6y6umlQ2/xLgFRHolJ1k+pG7TJF97RW9elY6bCn
E8Ryj4WvwbVTAeTTufYC5Q0XqUj+vWqj4EEiNZt6icTgc1Y/7nHWgiv4cFiQhnt8
9m95mXjqzxDwPmy16JTWrhbmqLgHgGuYycFBbAm6+X4Z3nL1dnQLwFLbmmmLbPcP
Ap9nwofb62pUR9krvd4BGFnjl1pEWeMuFRx24MGOtQaqBKrJU/u9AS0pZJ//MIU+
BdLVmLvCJLS5ggohMS9wWWNgB9Au15pBzOF/+/XWk3Lw5FGdfWgIz7iva5ZyaYlb
3FboOH5tWe9Dn4oFzG4qeAHNDfuzh7ckUqpzA3ahnxQqQMV22shZo19zQLWlfJFa
QgVhn4h5hK3fqP0c2LLVsHktZN5atIiBtsGrJLwxy9DCMbMMAqMl+vgx3UYgtrVJ
epjoXdTpmsw2MQFG0upFuBTjxmksKExo38d9OOBa0V4X8gMjQTJh6yPRXrV+I/wz
Q6nf7vlAeLXmOlyQIJa6n6X2l7KJ2n+85Tqhtsu3u9UaESwv6btrPaFVcwm8URXy
Y9W5QefD78Ck5Wlr0OwZDI93m81LRJjK4tteyhcgqdQCkNZP+Cy/GGet8x5tVBqB
RA33x/F6Z/7UoGlDdDpaQvZazQU2OSjLfEY6J5GxOxveSS7QhNsY3sKaGNAZwQXT
V5N/lXuhYiW2LSoPueqM5Dq3sql9eexw+m3+tCMh93x31JICZ1ssNwf0BX7FQ8FL
PfQKloPC6VeWYckYEOnizrtG+Q36J8c63IPjRXtFDfIfCcvk19iERDyzqSweqqQc
olZc9Vhx5akLBkSgarElMtbZZK1P28wCtoWIzmm+9WJh+rRNSTOK+vuxT2f20lBw
JmxDApVa75utWsdPiudGq7rE7IfI0MZ2bUfH3dJFchrTBbXyziOdA8WpldRdcheZ
CpCc3NZFMvf5Xto7uOrIIgeft0BUPaVJZ5JDbDMcpc54i73QgpevDI+FzdL8xpxn
UAL5qmwfWWTzN8ZoaC9/Rm2WQ/FC7ruBN8+JKorCxSOwCGMiRCmZP3Wux7nI19vK
bWIQoJC+CTlKMkw9tyij993kKE2Gp+oQW9vFc0oDEtuqiPfTkZlfNTLgdM1ORgA/
az0Kk4aNxJ+a1ZPfFFWkg0bHh5tH7vAnI4OBnBKhSw2EUQmoy6hYnJ36Yo/PgfcR
kFrRaBI6U12b6gZlauBu6vClN9kPgRfE3VjQY19g4xtZAen2cGJzGMFchQ3545iq
78Smg/FfQ4xjr+ZiRRPY4wcGMKkSqupk3ha4ZKn8HBy6cKfyOp7NcosbvF4VKekU
N5ofBPYoJ0cha9IiNpP7MBlkjqb7BcHDO430gF0Iqt2aNHMNde6TJXPHEEJ81XyR
rhfTzD4c5Leh3zdWdqM0tHeV/sMigB3GrFd08P2KEXIDce6EXKleTwzyQNT7Qmrc
adHAwvIapzNZkH67jKvFqMDBgVgOuK1YZ6sDadBb9yEXjkWPohfJ3NrTPJuob0/f
cLv8c5YiV9Qe1+p12u9xfoOcMmwrgzIo1TkFfjm1Z/fHCcVutlvrVtu7yQbhgVJk
ITqveP9szfnnbuibluIi/BJWHBn9IS1DA9sVuISPXp36JuQysETBbGIBldybqJCS
JRdlvidCRU96QHPpKkRIw7jYS+cLiNZUhQfVqGehq+NUKIXUJVhSi9KYTOECVCe3
vS73ZtirhnUZuqHNI94ZYFDm9dNIdmkf5RMPGTLer34kR/j1ghqK/rdbbzC/wNZ8
gzOnmOgnR3KmDNHp7TN7HZjLIVzDK6lckxHBrzo5GNsaU0ZX5HQA4WV4VeM+Mt1O
MAWZ/lDqiK609H0gIjiPG54lCeHzL09i7E9WuFSupqz6uItC1ZvBCGzS8abOKL3a
ffPJlvV+PfzgI5T2+gXXcaZp6YW6HtgPUrA0hZa1RbIpb+feaugTalJTFDGZv0pP
LBlW4v9WXBnFljkWvd7b2fG/cO9oYK7JPLW3ojsGoMjQy2TsbmQR1zxAjAt1HE+t
9YSJAmbKPp0ttamW+0QmEXBExBRvG23SrQqWQNdV3LLMXl/FCBki86p4wHurd4OP
rUAsKSHGBMHlYZstmzYnCdzB7DUN5yCpGugxRCFlj7XPh9cO/kzspZkbhBlcUR4E
S2fkvFnT/hB6CAr7K9LLwf53HzpcUbOgaQ1EJInWfETzoM/6Ou/Y1T1G3OVoxN9z
ujLwPplYR4yWNowLpTvthR0koE9gI67A6/SqAq2oTvu7P414W9hZ/+OjE6Xl8DHF
j2XZOkJR2+KDTGyjM3KNrqRDNkLHY/48UH54izvfWVotI4fhSbUI8m49RP9QBxnp
bCEoCEqe/H0DVOr0zw/7kiIty7uI5AsSNnnkFrFFsF0wXTcMnJPtkziZZNkD59tK
tOjxlEo44DYqKB8rwoc5HuXYTWGAFPi3jjjRiT9JWmpq9iXurEmWEkgcF8tAnGhj
YH5g7ht7EG2wV6cW6S9qosM7XYbmF3jFBpJ0MkmTj3DdJsgw/z7vPEbxhmB0bS9s
7MxrOCxbIygjE80kxaoOLHvPXDHGa/rUzwz/czQAU2BzJrXoQz3fvnn4zrPdNSfR
mkROIECBD2t/xa+ZW1ghoE5Hi8keywYVf+HaN9iuSYZcLGaci8sFRCm1TRu36sLj
8io/yWrwYyCdhvqVwGq+A6CLvJK1kTT/sS/PKsyhaQcJTmfly20Z9eZQOpzc930L
EAez6aiLkdudoGTvvPNQgjSO1UlyWGk92oXYZM6IXKo+otD/1cAC4OEscAAZuG23
jFbw5qYHEldIMPBnVSDhAhTgQwKh4QOA1FF5/7m1ixaybjP1X7m/g9D76DR9/tRE
iReODV1/xDx9pEq2xFFmZc+whJJc1CUMMTEfFnPyT9csXxDmMUexub/dWtXvQOKg
o2vwCneCy8Cpunm70hZJl4HiGzPH3qDIWruWAzTUY8cCjhHj3VDVF2bbIXZNiV0H
/1orhSEsSIwhsU5SDQxm9BcaHL9z4rwYUPHbLO5sqHXh/I2YDSJbYs/PFDzsj6Bu
VPIgQLRwrrizE2zbTaiIvVhSljfCosLm5izP05Y7S0y5JX7hSSHJO0sUEamnd22C
w3X9ZBc3fdwhHdxzz7rSF6UVmRRggPhiDam4pZ2y+zshoypaDk/eULxcgvJ56y8y
avC5blCxgG/kMhD+LEy4xULgYaXaC0Jd2UsP+PL4vxYCoYCC9FU3sYTEf3WKABfy
TyI30dw/nhGxdJkyLuySIcjya6oX2vZP40bdxiRJkQqodfvLSpdnXfYEKPuIDmL5
REGbtmWRbOZcR3pn6B8TeLFlKcCqinY8zQgxwXfVHSHz+wEav3PqN3w/vuZreXRF
oDm5UrzQQyQ3LcbEZVqWx4tqyuvBRxn+BmmuzwyNH+0BpU5/cOi4bcDRoO7bOEBQ
3cIbWeifMrnp4wEecNAI1Ns9T4lyS7kKZzX48KbsrZXL998uic0OE5+AkxQmTmBW
UkxazWqQBVDEwdr25X5rtZCW6wHI28tmTx70FiNF30MUdjdj9fOjw4jtIVTB1m0j
psfD9KTvvmwjTBznvbegRmFy2TM/oQ3fgX5HL2NA4OEjPd053vKG7RTg6fjnGOMc
A9cOLPT1fmKnjp9KnjanV3OjR4XG08QqEn/hqUud8ZpLoE7bhz8XjvHWue+IcZlw
Kmfvq8v6TA8g0DEItcvGHz331gl1TGA1QAsCpM1y6Pz0En2hhBZ94FdFSgD6NFiu
uKGe4V6NdQeO/VYemVn81KsPhSEx/Vu4dtMx592NKwuMCNV4pIeftIemFbNDRfAH
AnQAlra0HlXgvLRgjrHusnQbt5w4r73Yb2gmj0fqY6uhvvBFY7VV3QSRWCQIYbzV
dN2qAP1D2jjllQeP7+uSVKsBZobrMfUrygTs21IXJKeu4e0B9Qggad2i7YYYUwRa
LaMRR9sO+/qTHdmpXnUtJArd5crtVxdOGcAtVMINX/OpMVEL6Wb7PrZCOT0FUiWG
685WGDwLi4l5j+wYuBvRjm3VKDD3vrVta60Cd9vWeRRR//6rMc2f/DnG1IBptgUF
KDvm5xTWlSmEPTtxG4yEkofH5j0Q2rKiLeZ2OQd2JD8D2kLpQKXnaXA0Udbv3rDm
eAcFybagwGQ0LyLmHq329UclwBIY4IgY3iBnrNk2kU/eOoC3fAWYk0DfQm4njN7R
KDXe8/T6xauYswIeXA+cDyouJjvdK0McHmtmZ9gu9iWnuM7DyD5/3/xBnV6QFRQy
T2TnJzifGwOEz5xINx4rQoKB1WBwz8bCDqrCl0krdjAsAOw3VFtGIjv+7KzwBz+L
7m5lGCycNgCpwVBLKB1fAI1jw1dfShWCXwuB/Hy940dUZX5OSJ9mljuObQI13/qD
aA4m7gtewjlh52JRhAtbSEFZBKZi+eZu0BfjZYxQ1bhzLFK70Oc2tDkZqOQzaj86
HrBJqV+hEcqcaJf0K0zXHAh9hZR6C3MqdswqFMDV7EyLvrlM0lTJqWUwnZrJFRHJ
mHSyU82886r1kJS/+V9hrYdw/y1hxYxJfhwBKLEdbyiF0M1C1Nsd9f9UmVNz3lyr
pWg17F6tguBYqBqjThIAP8rp7gWooEg6bDL9b7cS6437p9ORNHqPotkSV6WW8wP+
d3Ch0rSvH8IdGu+VFSlX0zwg1lCSRwV//qU7R55NU2yt2jMZuiny6sUnOtDYBR3K
GIIBXcWIX2zJMbmNjdqNcC2sq2XuVir618hEh6sZXCGBSmE5MKDIfF+sxBgIllKs
RvA7jPvWQTZbZfpIhC84gJzpmIrJHPaCzgxeKhQQM/Z1cLBP7IlUrWGT9AKpVosu
8qPUSh9j1RinfRRfl9fX7CWIOOy5P3QJLJUQYXcu6NoCQW8LhMby8brmAhUOvN43
MF0KXEF4CbFkdyFKmeIGyYqI0gFExftsCyy5uvmxtFG38ApVB2e69u0BF9YfMFPc
IV2Yd3f8J254WqYtWkiYehXRpmto4ep+8muLm6MCON9qsZGlOIseq40qSo2iAY6T
qeEZGAFAcdlt6avGbwezlSDtuayHHjcatRtIFhjocwI+navq9NCEy+2DmGQJi3+w
nZDcDbQ8IaiI9BI6OGrUQQjAZ1hrre7INk7hGU/2FYR3Dlpk0sq7BgyJXCsiHQre
kdCN6gT8bg2/2zFgqIl+KiCiYn3UlziRY7LyYJO5tU4kJJjuWyUOPwbw1D7lkrM2
OhjuAgM79/poc/yYCMxCWXhsHayRN3sstmXwSWuDErJADYFp/kWaniVwsGZv/5Cs
0wK4/A/gpHjT/TN0rXdseaui7HuJNuR80yrSC2yfBwo70fljWAg1O/FEwPU2PYon
L+9p44sDzfi0N9vR7g78lRwh/iU9yVgUP2xn4DnH9YNJad5Ks9efKG92O3T452QZ
oShVyUP3MhEJayNynOTE3Aance7D+t7trxRZF1et+FKijoAQKr6/lSJ2z9PudLiv
ntv965n/yigaUBZKQIfvIyt8D614b4qJTCy1BiNTkox9WG4nM5NTS0AmLng05p5C
l1P3mFot9zoVvDGbndKAnYOGjiaCrLg3QuEqi53b7pZnb+8lBD31LCL/mDEfS+N6
Js3e7ILAqdayMQqA6p0nSn0fSOUnHWHw+vibONfMYtzyVNAIJeSyY9H3OqdwfGk3
4BC7JwDaFk+rARHwMGgAiCaFS9y/l1kBw8ipfWq4Yx68sPVu8hbXdl0RHG6wsYRk
ukz7yf9M+wMqLHEbPj3tXcNU+l9tlTU56Xy8Yu60x7Sbz9SPx1dDVhzbcRJWfCI5
mqlK/r4og5Emv9dN1QEyyIC3IycKetvO2tRhB7nAnpZH5iafaSb/XtwkQ8Q/D5tX
VP7lmYfFDCrDQkhP7etXRSkSIbMmyoJcRzx3hK1hhALi5SI4xk46j8p8iV5iO/NZ
1FbsYSPK8Jq8n6cdw20/d1pnb7htASHXdZwj28yszGswzUQa2sYuE1VMCkExBTq1
B3WrCCaK9MfIQhVBtys1FIzYAN+6GYBFhONHeTbNbh4pVBbbU8rXF+4dmgSVcR5X
n2bWVSiOqhHJ8S0Y7IsNzloIBFlwzNgq60n9acdwF1YVWiqa1AMy0tXXULHZP6LA
24KHudbotV/96QkZ4dvmzt5OU2X30zsVkX1UT9GUGHaj8wlj1bFya6klu1F6jS0E
FjdM6r3y8hRt3sd+AZA4j4ID7jnnQUBch/h2Afk7M0xQLeUx1Ii6s5Q2ZLe0aj2W
ha9AoPybuTD4S6LbV6FTLSSGxQFasf8OqlA4UiZFe+ezwr6GVrY6PqcOgsWbZn32
HrtMYgnHq9EGtheGCjTsYWn1wkoGfafZJ2HvJ546xfymS37QxjT2aSJXU1/6lrk0
OiImGmf+g+0tI6jNLDb3ViQT7vAZcu1nYj9xxgqvl5x7tG0rZoDqwhQ1rRthy7Jc
zgDxWSt8n4lbydftuKowPC6uqk1zCkeVzfy1luhxPtaG2ANTVtjSdXRlm998kqvz
VRZDDanc4Gy6n+g+Rlm0QP3wCoSIDjmX7jxfqLf/Tx/D219e8AUcLVm9pG/qxnkh
nLnA0CzPiqx8m6Dze2zxsUbk+Ek201Nrd9NQTX2DH8JHrBGk/Jqp+Yu/zbBGwxvW
w+zPQ+l0/oV/2oSvaWx3e5Aqe/mUKZoBGEtI5/qj3bXLvJJifvTieA5bvtN4Ipjx
3rzCYyFcYO9nOqPTtmnyMb8sNeNg4xGrxAKlFQdz8q7PIjjCcFTES7PwzF8m9P7m
2TitZDj3klJSaMOn9Ums1T5fBDaWg/s25xnHY0WHH4GbiiC07+8Y/s6bi/Aq1/S0
WpJhjekghoeNEXzU0wx0sCZOx81XdpQAM09azriumJdIMVyNFxdrDI1mWxfg6jOC
NfJjp8Lcn4smcwaDnktlvlBxnYEvraZy4n4y8Toh7NrxzWlQ08tX8jj/xdptUttk
EqPRxGnSp03Odm90lDSqJpgGTMTD9faOLy/g5eXQOaKSIaPMXJ5029+EIQzAyFTn
UmodC5B8u4/r/94JjTKp1unFA/peiybhNhFbN7u4Fq8BZ4K+e7jZolUwk2UIh4SN
zBmagz1g3zNGYI2bvnQjw/s7jSUk/oJZoXAb6yTNKZN4nPmyy+4qqi+3khOu0GDR
DmyHjHCBvg01yMSw/jSa3e+DrFu3q/FFouoj95a/KqRsuPpCG0Uo9bbpNqFNQYAM
TvQhFbNRRQvannAyX2b4Y6eSlnrXCKibXl0/ueA58bGTMF8r0n2KyoJzqbBSODHk
+7aTU84aq3tBQQ8h0xbj2Mp4ls60tZqe/4J4r24K4gS8xII/QJF0IrBYieE0oJ0f
r5naxVQD4f6/FtA69Mj6w9cODu2yW8mWLCJXo8TfKgPehmRED8JRUA4CYmEtFMmi
enwo/QYArQTCdDOSP9xz8fo1zMoAWKZv1UJGqrNIrm8l7iS6XqtghPYMC1eQOZ3C
XcnJ02jfKluV1tBXuXYiUNZV0IdAZ5zshoD1/DR3tRonjShq3MXWfcWCZQHfYdtS
YCSwINHAu1kEid6YVhYd+ryLp67i1//vRs4BO7UpDXjOrfxElFE39gZZs79iiRa/
OsKHgnuRL3U36GmlkEBMXBouVvzLHqH9++wERHJXJ6FS1F0Vx/c+fPoMt+ARGQKl
GFsOD/Bp/vvxigJwaETteARSsIIKTbf2xxPmIH06+nvwiz6SKHzUxwRxFWUTbLkZ
8wbsro9gevAqJS/es/yvP/abFgBAuC43RoGWyKrxdLKS7atKLXQfdyvG6Uv3W4N3
WbF5Bx6Bjcl/606i6S9IM+0YpzCqQ+B5rSFciAEkPzAX2u4qKjTY4XjQRZiE+44G
vCumasD8JBfN0G89S2OgbVPm2S04eo+lG9qPiizuiWnpgABASm4mQzu+tfJ3F5rD
QSrvEZqIY4NpqvfxEbfg5jwVsqnkWBUJn7lEFRqxx+tO5RbdsUYFI1biYbwhfZPJ
GSevS14VY+spCKb9lhSfqj+bRhaZ6fvTUAFALgStuyJ6Hx/3aSSTEa6S0xQ5QxJh
AUC3fmkzqP2unt3RkcGGIb+50lXaV74p9B0Z9/26NStq9UcTMvlnpudzmYj7cMgq
ejpu3W/z+z7IOOBQAicEpWf1PslQlPETyHmxrMWZgdxd6YBlbrYdvzAS+kalPpAR
gGS0QzezVYoT+XZEHI0fzz7J0eRmVuhfltkkcMc8itL/jqfyx+8cxmAFq0LpafHA
dliyHbgfVUoP/V80Bsp+8viEfEnRH21L0t68yXZwg+HsEkcuioRpFmtUneUxNdpq
eJj/gVYiEksOPYjH2CcA+1wbGLp2+yWU5g1V6Jx5pXvfUPyk4PiJqhHxoZosY5zM
v41sfV7I/tHW0cwavwZP+/FxmBNEpZ9Mi+Wu+zb6JW/FFK4mK/n2lN9tdTF4ziC7
X9X5ppZDYeSR2pUONbNkg23YTFMtfu9cL8pFDkdAjO66uxNIKMPXDzE8lKV1Q5B9
BZch/YGdl0Ms4b9ANSJQEzz8Sy34Yv22bDXUPLpZFLqSm3EPlw0mrAnBBHIkeeCN
YDJL2E7o4TkIzLJYKsF3s0LyxL+QEPf+9WTqiyszgJV7/v9GO9OTkQ1ppvtoR+cm
OF/6X3TjvRt4/TWzDWyV4VqOmIzynNS2KzOexezRkwM1UOYVA1Dr3n9Y/u4GhFVd
JB1+D88NQFKlSIWLUp6d96CN2SEDn/WExAr9jqUSFyZ8id3BNauwgbbryiFYTZEV
+CO9XH/gX/gcqQgOuE0pXz0QI1vc3oB6Sx7PM2evrbGhsRy7oCa7OE0Lb4H0uf92
lBVcoNzotclW0pmKh2xTEU05aoeg+iOH4q2mNZcJv8Xi6KRkEHzgC/EV8OSnw9rg
P0Vt6Dv8WjT6rmEz5xp68ovobjeXQ4Hg6F8UNwD4aiYK9+bRjH2GKkYMWLdCOWsT
b5+Wo619nPisperKWkpyXXdfxlsLaImTbCWcHRaOBSf0v8ImScPZ/x/+zzCytaJh
nvyUxrF6cVNvGqvrUCZWkhgmqIpdJkszeYVBxvCovoKiE0bzXbJqCrl7tI6JeK7O
HMWZEDJND7V9FXArVG8W/CuL3bKvGBldp/zuKkHBPsuIz/sw7wadMyVzCHmDhxHL
lrhxHN5q5+OHeXyyZU48FEZ/ISfKSUIj7p67fc43c5Vf49NpswMYVH7byYazuNTd
KJ3KaBfvgARSUumJ7+bO+2EdDsqF/ynCVf4ag9drhdcMgn7dWisZVsLU0uV6VAI1
Qioow/o4RujYfHfJx503RqzpxI5PbQHiLtIH7u1CW+tWBsmsf3h8ONKPBVV8imwR
EVrm2iTRax1pz7ZqJiYvWhgPK+6iP6lYJFj8tt0/bOYOe5tJBm0U7UL9nwqting+
tthpaiD4BhoTyKiK5XQ/TCvkCiwQgN7twXpgiDDV6f/WD6A4SMluaG+SHsD00X+r
/zuMbIxaYcd1xC7arZclvJUPhOqV7EW+KZf51Fup2aWmUbbVKj0MbA2FyxN1Q79s
O0Mk3rUfKDeXko7O5JyBnc6ayDQBS7EYGVo45OwT2FLjQBwaXls4PrAJNJ9WyrXA
9m1yCmNHUioinpJmndLfbrhPNDwwh/bWqwRTgkfZKLCen5Q7CNOmh+vj1qr7daGq
OCGyRJaHt3jfkf3mzVVDOqgh1skGstaOTTO7p9HWcVDAYUID0yfYkOrb19ZZm9Va
pv1baOeY0/ayypaOunHXl4XeQ7tIjUmoHpAp53VXNRAB++gfJm1Dl2z1avCHZ1/v
REcTZVnkrPNWuaixR2IxSHpaxoaCF6cjNgC5kIQ9qr4uwWFa7eaRxWwuXM04jcQA
GD8BsJZAcUZ2P2BACbG2xFRaPtwyNShXd3DnhR2TU1W4DefBwroegg/4C5C+eGrT
FUUsGTdO7UWclT56mrhXubTe/pzcMMQgRyMJMG14q2qQFt2Ltq2MjiFpIm/WDaO+
xn2uhXTzIcSqfNoPhi8akNd6bXJs2TSDOxflOqO50Mh2+TKeMHyasBASRBCkGu4I
NkHWRDjJOCWfcJ4HREoegdyGfwI0DqRNiJkCa8o6Il8mn3o8yjSNBaCvYt4DSSgH
Tc0XQQJ/6iJg442MWvWoS91SsH6EYPHWwow/bEvhfO52BMS/t27Ce3LWvjKT43dD
IfZqk/QbbLhzTvp+7paQyLEvFPzenrf4M6xmaihHJOZOq0KrJA/yEFhi4yuAAKWD
HQKMg/o8MCaZMlzXHHfKsOi4pUkJIQaSTCmiMSl4Mh60QiifGrmYCk+PJcm55CBw
G8qZB34RsLgieqZkZbYfrTxgI0QixXObAutNDmt+j6Z1620TQTtBmWZUwDW6l72J
izGuVrAlOcz/zC9vf6Xtfz9gGbDGmTb89xb8ArOdIixqdrEtxl5OX+paHmaeBv11
6TWH+hRID47jV7kRV/xUsdOU2/HV4B+4HlEHLJpbn2/Ik05kxr3QcfZVOsK6xZfW
NayiR8QwSsYnX7tuPEnmWOlBgGAtJ2QWV4BoDThVSbscOkMeDMPMIMxusknoMRCC
jx44bDBP653ovO7fy1oge0tKyPRXI0PQr5ftWJfslsEBFj1ReVrD+/9+LQ3O9Bly
XqjF7gICBOtGgJwtbxG0rxMvBZNIk5rwM53/u1I3Hn6IKBECY29j76NFsl3Au+Qf
JqtLq9NARDXTBsIxFNuCkC8nwKAGAWl1fWl162IrhQnqmuiEcRf2Z/h8Jp4OdYHe
8S1AZkgXVwtEhA5mMxY881EJe6q/XweHYl0u7j/9hOP8pS57OXxc1cLMxNoWAflo
uo1AICqaO6SXZgti88bp13oMLrcVdtNDbtOaVCK0SHnfHkju8hO65gRm7kQS8QdU
o4lLyIpfYGq8dNvArRzYbQHdNCr4muvPZV6uHNRjEfRomKA2aXPk8CfQH6JMx0ob
suPEP1pTOmQkqEplXdSpkFO2/QPvJdmXZBLetYwyfgX278ZP4LGMZvNzi1PvfrKn
mDgdzCT1voNxdukIBB+sVIHkdtMjz+f+w285jWLQz1vhcIwmDn9M4l/ldBw+sAe6
Eb6QXI7vLSJixvFPbSEWmUNegmDk8vhCkR2u8FCQqxg5ISlIccLAfHc2aj264dlk
d5RL6YuT1bbo86a6AW36C2h+uvpExHdaU9py6V6R1LSFvTN/9eo8LRsvObJHs1gi
GB56IuApnIa4koKgI6tIJuNkRf62A8lhleOfF9YPkLKALGp0k6pY/Cj0Qi0DrrID
x9Mo7jSUq6GO51FZ3eBfyecS9ANHVIoYSulynk4ciicfh5bAlkOiag5wZHuYK6Z/
8u9DaNuIZzeXfizvWFFPqTNldbnqXLnP7bTnLLiVbag2B260jWkLq+ecFFjYv6p6
vGGyho9atVTaWV0Jg8/ZpTjv72V6V9/u4HyDbsAlXA0jxEcb3g+NJHjhVQllQvUt
ESNPBh/kb4jfDQWbylPU4PyRcSECkvWqrsLAXYj3z5v37xUaMA5/a8dlm7SSnRNE
CzKVgxNXKOAeWXsZmUNmMZXCB80MMX0D6W0JF1U+WitpUeKHqGxCukNCQMoj7WSY
8Y25RdURstOYKExcSvSSoUZSZmv5hz4FyGA7+EFblnSQEuAQ+9z4CKu6+1ZnUW0p
TyYlTgHbna3iJPBCLsZd4lsBWXmL+z8VG+6Hh/RlwVOPEYrlgs+Qi/48LCkirTCl
ASxbdBHi6Y3nq7umPQvXcaPQMBeg06CqyqNsjvci3vugBW0K3GjjuJnftO7LlZDr
DH1W/2HhJr/BOQ/i096Yc7UAMjEguaGv6vfHAPWdsT32OLX254VYzX3sblThWGQa
ySTog9jSsdh59XKkH4vyBRuLofWR2E33X8HqsT9UPUQ/macsh9M2OkA0UwaXgLdC
0dxhjLo+crugNgPKph43bU5OL6NupJ1MEvtM0gED5EveA62CIm/JI6Zvu4wqGwSU
jZsDtfr4YWd3Vl/EH3sPNbQAP3owUvmm8MqVGU0YQsDCEW5iupmykf5/roaTmzfy
eVjqS2oVg9YCV/62czexOxxb7xzMNorbZLUPwaknjPm8Q6lGBet8A4s3lrLNKBZV
dWuUT0JZ4rxMebnGT8j9rVj+TVqTJxqVmSS3secKa9gR27YHxbMjzI+ybEaGyUXV
KIRXmF7T9Wv+gAX9Hdgf63FT8trGIWBYHlXhRslbGXTbymi9egajiGO1EAYxJYqO
9leRzcDjcw3Nl9uy+uUXF9AhnlghrVavLIPHkuGcpaxpfusB+nnevha2lyaC7Cu5
d41Y7YZG/sKs4cKUpnYBaW5pJWa9pvsUaDN7t11TMVqvceJL5TfRLvYcEwbl0q93
2vHpDXl87MYpF5zGb/pRMtkfkIUT9lnCQXGTJWz2K/nWX8JENf6Hggnw9nhCNpOq
ZCIMF9S0uDc5Mc/UoqemraM623O1FobyLNBI8mi7qFBKH5L0qWII2z7JoQ4lsUwV
Pc9h6jtExOXH17ZSRpy+HSElHMeVqmi2xfjlJ5PWHPa5k2tBmPWE/8rLgSoBjdSK
SgQr29oiam5qm1FVerYQn7T1FEo4E6Izd4EVfHrLUuLXcvN22qA7ozGD+AJP5A1Y
1qvEo4YiKCgOCGTjg8iAXCUwTIdkoPT3x6XXWjCm7cwHu3UIIYV7GwiV/8AYPVWe
r6JNCITUswf5nGeosCuNJwQjE/mlqAOrUJB1sWY7cc++il3mQwAt8sMmJ9VCfZhY
5QQhqWdtAuxwV8hz9XszR4eJCl9ub7U1Vu+MEHPEwFqu4/SAFOOuN84sQahomyCQ
2Y/FhQ9kgUHeJepBtMDtdFIaaM9D1Ex0ttURgXfXUsSQsWToX7QpdOP2roF954MK
EMokr/L5WNuHdBo3B3qfwLpEXF2TRoDQs0LYT3KavpOFKriYe5L1wGlMsgAZtXDD
NRvzjzRnoOF3I84SF/4q3UHSkOba3WSO+cZPhk7RrDRGdxQX0y/o5gOaztHB7NL6
fL/Wf6F+qldN/+OetmRao76uYLLZE5bQzenL35llLzJtkJvpJ4xGsk0y6uWm2Vy5
6dnQN78sXqkwWnEjXAPR3nzTrfxaF+qQCirKogxnE6jk0BpGbvMrDFQvQrZ6l1DO
z6/iasnSW1Tq8xOcg/WTDk/IwXJP/wQ8DpZ9NFubF5AfIggVJ0eyFMZESQgTB0hd
a1+k3s3YFG7J6mFrmAHshleRiOrMOM9naIONQrTUfsurXhRPkw34Lf7C3S5iA1Mq
+EiAwRJsbpqlAhZV2v9VR0CftHfmGxUYoYXo91bK09HID5eHRZBfuzxqmSnOhvQm
3mdeGjM4H/4qz9t4BxmDZeeG4f4bugpHLfssaIm46YgKwVT8bZua+6lJo7e8s5zd
rSKxzEGWbDYm2DGTVcHskBJxul3xV73nel4j5t4DKs4xkIRm6slmm325Mc/Qkmpu
R8jJaG+rLVwiie+gt6Lr6Nt8yrXYt4P83dFYdHL1SJcGEjYjr97ubnh4ofPUAZb/
AHyiG6B+NdkZnzwg9yjsKeeU4tYr4KW3QHiKIgeYHgSVQbjToCgqCTEBdCJ8ZIiE
fElVH0Mn0a0H9ZLULqcEI1uJAwNITFETrNS3yvesFXcCNdKwK4/3Vts/BL9aKGSg
OAzskY7VwAH47j29irKwKa64NOG7SKLR7NdwKGUeJ/LIEZyEMHnChuOHDkqjS3Pq
D/g9aNj9UDOqeclz56v1qWpuQyqe9qg/jcTgKAZgxLe2eVXZp0u6BojOdCpvKHJP
FegNarxyD2lZacCf7F5liy9YFZ4BkBtYx0nb6xxaYqokvaxfqzaH7y+a34XxPp5i
JKCPxHBKz4rrBvsGLGWNZqoWpw984K6Off79feeXN9K1CUK1DP4syEwEV46I3Ic3
V7kFxDZ72s9BQH256YvVTb5RUkyeV75Z14GIlOxiQwnlAYgkPp3+RXi06tPgoJz6
wd2iQokHFyPP4upaFkNnA9LATqVxE4lWopzXPdBeuXXYaCih2USfu1/I3UjKA1Ec
6VZGIlPCU+1gpjzGdtBcfvuqQU+oiCaiguwrz7FxSV7y0kPfsQmjhFaRH5+bCfB2
AsU+J0yXWZ95CuFrpSdyiVIYJWTh+EBPAbC96UJ16ph4mvHwUebXuNnnvZbcTLax
y4f5QYc0ojKI65Lw11lWX4OO0Br1Qnz344EIR/aDwUmjDxpusK2Pf3DTQN4zn+6m
FO5MSEBQXVoi0n8A/f6BhcSn4VSdGh7PuF1sl8eW469BWZGQx5a0prK0WbJEtIwx
recSdr1afQepZGTjYiOkHQ+qgWPjy3HESB4j35onhqDmEYbdUh4vJmgBqFzg6wGG
5VMtGdcWDrn6qI9mCSdluxKnPnnwxOEFKnEicXTqEvZyHd1I4CAe5Uy39mxqCUJI
gbc1Bw69CMhhe48HLqrY1n9nL1xLmrqeuHSTLcUvc8OwSX3ZAiulGClziyYhSv8J
3xfspmUYdDi0BHlbD6RISrnIXi9uULKz1wG3w1Tao7XFeyEicoN0b/GrJUiPUc8g
JBIR0usO//B2hmunfesEG7W1TpMBfMT+wJDrh4MRIkk8XkGp6VgNTbmBe5jFBk5m
F42wDHgijaocm4J+DLkHdawEV4/JBVqjPsTOTzGdHwLDYAitHXDBBEIiiVHqqGUK
1cnHZ2RDgsRkAhWRpNxpSDQNF+vKBCXiig34gNG/uWOjuoaZYwuXA1PEjQ4OgrKn
Jys0yfEIMtl2ca8xiy2vp77h8XEEkN4KQRsUGUYgPwux5XeOp1zhv/W26DOFsWnl
G9bw5ccxEm0nDtjIiWc2miH8T0nQTmtWvPe4yfWHzFn2hV2Jv93kuJVrrnLQByaI
pAzU5owbrmxkUf/MA614qWjwALI922DdNlB2PASoNYtjGac2tA/Kvngab9vZ8WqU
EKA5prtT+LaIZMjfpcZS02flrEFdxSdFgWyizxVVdhsJts2pYpdI9QrN8xnv4fzX
unbKiUcmM7MYjTya9wUEyZYp05nRyJ3jVyryzXHZuBh3OFeR5S7zLlY2OmjpH2zE
2+Tfxl6S7Np/1alpoc6HFePQWX8TPnFN1ckhpYPOeL2YyuLKbqnK5UCXe5J8/rIo
UzIX4vmzLWZcg8j1E30DNmgIYHC+nPaLecvE43Si2iUiF/vSYEADMXl3/ssef6Un
aIUA+n//2R7Qwb6Jg9O4U7rExHwmjqkpSs0OHPfr3OoZq1fpqNt+g7PW/xsD4tla
cqH5WNgnWlmuT2RgN6y2k8kDyJFAmObFS1a4Ed0F+lOlxUSKM1R3qNY9DbhME+Jm
i5CdKXVgIoqS5GaLoraH3tw7nPe+2J+soMhYJHB+qyPcFrlpDnkGEx42SpN4gPAN
R3he9CYJzIINQGIqB4ijUcxjcLpNCy7Bx8EP9Kow40RQJI/GFdOtuyBsBag3Q7XA
dCkcL4BOyAEN8+EAaXKTOskQga63A+GYaP31/dYGjfnFt4UokV/xZFRiqrSHpiPU
5v8R4JM03LIxMiNzHUHHkrggu95nvVxAkqUfcdgMM7uyp+CobAZdlLhlGVA12A0e
6OQBJopIO8clTUjrk6ym/6Pz+P5+dLHssDkM2tzHVfB3b6WK+tCMhTYew12/pbWm
GJsXThs5UZNrLv9//r2o93MM7wHZZiWva453zjQLDwZdS5Ua8d61Eqa4M65h4BV2
itWonrqJNWiK7Jt1Dm0au2SEio8wJAFdrlHUYTCO849VJBNsrzNSCwwCg/xdqV8U
NJp69tvDla497Ci0O7XcXqg2Re29RM/U4Dp4cxukDtXurNFZrkg/EO9VqpGjzEk0
dudgOwKtj4n/IlLWomnmWbGM0z0Rd8ioi0bjFIqELCUL5vaGrjyL4bSdTeOKDrb/
lOLVwR/wp58wueutaFGmKvXVoBmI4vRkH64osyXT640lUEZA0wWnCJ9FSOH4vZ1p
QOWI6IlewtelbuF8zTtOPjc01Zn+QaZKb2V3k3xlBs/lm41/xV2p1q6jr9LAjCfs
hUX5eizP+24B9aJ1I5eREAsI6FerMNkBELw/ceKiXAGpQJ4g8k1hv0l0f7KwEGuR
fP7EmOhEYFQxtqlwViC4SfXCxIhCMo9YxfE+CaZfri/hNty+E+u1mXveAXSQ4mZQ
FzgPT1zPEYC+fsJYFnmNCu6vFvTT53TTFdH8jsJvHhbbTw7XQyWvd/kd1Pazksp9
2+kf9X8Mzv8N7ETFUIiGz1oscLMfjaiWFzf926cSj69NDCmi2n4aoZ0yN17I6kMv
LXkWWF6v9UkYcHiG1jbWsuDYV+puJ3Bdvwuk1j44RflwAOdwbm1r0X/Evi4rAQwZ
Xb5aExuVsVycHgr0gFWekJHRH2SEsygl6/vOOgM7NMMeht0ayWGHDhSlXPu0NjSS
bSCRGFfLgd8X9DwjH92Ua0Nkx7UeCEwSNm3zlZ9VDUKRMJ5QQfbMVwCekBwqCdeL
59tr6VNl52FgKg8pY/GrH+MKp0NU9uA/aLlNOBAKw5lRXyICIakgnU4wUN05h+Cw
GW8N6rOpOD8/S4zjLfV0d5Rw9Y3hucqbvP58YrIc9XoCNah1R0LBC6ryuc6T6/fB
9H3kIoXTRzuPq4QsuilIyu+aT8NJsoxzbpaH7KLY55JTdNeWF0MYif9ae8Gklsq4
8oWmB98kzLGcIEKsicl8EnLmobISY9JA8uH+F1WX/BJmB08eLnhA1q/xApyG5fgE
lSmTSD6e1QBLAdoG6ZrDAbrh8KPnVH9TBMg2/7hoq9MjeMdSAqrXRpaRB/+f2VPO
cL9PO3Fpw+HsyIXJcJnoV1ltXEXSv85rt0b9FUzAyTtPP+IL/uQxEYw693H8qAK+
tK8TOC54mW0vbh4Wp/da9sYU7wjlCJiq5Yh0+I4hiiG6Qw1KqqK6LscI5efaiwo/
49udI8pBr+kkMCOeNi+P7/s0FWZ+5qf2KRF4xXvnHuEkBhro0Agkrhy4JbogysL0
rbdDT8YJFkTllFmOgMSIOFr5mQSAGvpH4X5WQzwsaSa/TzXdpWDqGleXhmBpuXqn
Upl1phxDeq80V+UkVgA1EnfnqCUZo13Ct/BmCpzzAZDVgAxWBtnQ9KwGhUXQK4ug
xQGqQeoD+fhcFwg81Y7EGkkbe6kIpEkXKH7Ov/HNpFhFnKihQfoZqTs1vyo/1S36
x3zjijBCSFaZwyMIx/zclFdoSd2edQ3NylHen+2nUT7uCrHC9v0vtktVi5JOSMbI
J6uLWWm4wrmPTQBZGbsmBLQHgn++NyducU26zz1ByxZFNpQ/MpwkNi1ysf9i0MaZ
wvv3dmAyr4/+7kYZSIUxjZ06OnGzxRLobGhlMXmfvSO8o566NFb8osbF9CxUUEFj
QFamQn3NVg2kSuGH4nkaD5KmaKWeSTDkVcNbtYJ6dBS7JgHRtTIBmF3pAiLqypCS
hUMQyqRZJBnN84+aXC3Yb0O+CJO44xP2CBRHeMr/mIksCqVP+LnETuSv/bkZVQ8O
JE8DlhgfnPRc3dIme9UoRe70GqW8A+aYd5BbGRPaw0cB7xr9cfmvJKjJ9Cb2BuSj
8gHs1XCoV4uaobOABG3eBNHUBzrMFrlbsA+Qna1X1DsHRPyhGA/tB9TGWogdOuzI
wvtnGSa/CW78G+Lo8//lD7t4maDSqSPWtDErQyErABRNsJ09sBMk4B3zYCS4wwtE
tmCaI5v+F5KE8auS36m/AJvfrJho9O8I2duCVEAN20hujADGJwPsPdziTAntV/BK
q3dQVv6P+tTdNFTWoRmEqisfxN2oAUTVt9PO/dj/iZwCGCBaJTie9AWqjxo8HJLt
LD37Czg4QbWRiN7n7zJNrfu/T8gKj629mAYKx4IExrwDxVQL1USiQuBl0SN4Vkxm
gkeU8BKUHqWXedqfj7ITZqUNPW92t7pxc1+Q187u6O5FMhI4lT3xm+vSMyyFdkFC
F0DA0Zoo0Cv4BUM7BxT/GQBoEerSZaoyClIqFn0LNVVAoo1YMt3dqL5JUMwhmL6t
NqKKaDUp+B9kSUHqLZH9mD8Vt9aN3Dt3B9a6kpzJuvnn8i+49sbCl8rDovBluTT4
+BQqtG8vuLTAAl0HEquGm2FJe86LpYwxqNXg4lqDMQGNiHI0y6q2SeQcgB9ijnBc
jwWGdKEyONVorSPVIAuPXiAGoV4jNRQMj/1p19xT1SnjYBOON+V3K3np+jBDnFru
4q3oiibHVmUlPHLswTbLnLleXCHKPN6tl9MHBJqFfHVa44ShWi9fL+dMrSyrum7h
00AA8EyPoowB+W0Msh02QzjdduT8ScbAxC1YFsI+ho2tdvnlgQx+uZj41ZUF2OiQ
RG+U2rOM/mX6kbtKMQqpj3KbpSSBeT885wQC1656juMTWNJFTB1Zy1RfWet5v/Aq
MrGCAfsU/M/PCrmT93A2KiBtJKWwzfYDpgMxe+ujgfx7Gb8q8bN+Wb9kByZiYv4t
MWZeCFO3wp3YbnqVL0UgO3V1NDGrkHl9BvlqA+/W2QAlUcwA6KiXK0zlwtsuoyls
D05+xxxDt8cJgFWOcAnzVbSqNEh2Xr5VHbCmwO34/oAHu0yw2G/qzC5BeBywo+Y2
YIxmaSE9HZfUss8pdYx4e97zUHoEWtsE9IQI4HTPzplWBohPxAqGiaLPRfDw5adk
nwTV3HQuZ3Enbq7u2HJUoAzxAezVHzORhhqNOlyHb320laBMjkmLdSQSj/EQGv3n
x+QfoTAf2TCMOaor0GhkD+14xJWsjn4Xr16QNtxOKoWyM94NtM50wb9oIyTkOI5h
CKCET/u+wi53rlLxm4friOjNiwQGHUitRZoZzJRXS0i3a5C/tdO/bZUbCuqF4UBY
8THinkXnHmciOB9r4aM5j2+wgi/322luUhjiukb0vtNL7L0BMKYltB8oVgUM5H4A
ail7hoKwwlw8SojBrGfbusd/PXPIw+Ywut0/P2Idd47ywxQwudfJkj/ERRDCi6bh
1WuVwRdhplfuLG8k0aEsYJ9Ot/mf/Vkll1w4UwVh8XU6UFf83dsfMF641+/PnOl+
zblBpz8GD9JH+uMKQMdQK3FbBvsDPWzprJrwEhz56A/B6vkYNUsoObLpyxvdiuN0
DcAP862qTiCszkxYfaI2NjwoA4o6vex5BeFYj7F7XzGFv+95TdUHzXd5JOK8+veM
X57jRF5fObe1E73y6Y0nzMawsRtKnH1xpy/AQDF13QNzDIvV/ibFyPcpl/OFlZN3
7CwojebF/MgZRs5NEOUb5oc0TYFxhyIufV5Ta0N4aDBQ1I0egZy7v2OPGtvakBmT
D71CRuwSg0K9rdcFocFuWbjI8Osx2tQNi+tOHF58SnkWiYQF1ZM1rWWX4tKvy87i
FhhZ9f5IRH9DB2JhVsNK/3F8z5GgnrrAksL/m4+V63GEre1rKhxfmzcpuddwOedm
im4MPxyefE05i1eHHMhMOsXJeatoW+HYn7KnVqxqY09HdcUVUnXObTRVTpjD/yAa
0HR+oCwSGxEIqX7SFFBaCDzqs+TPSuBacC6lL3qf1oKVNGUhn3YC8RC1iaDSQIzQ
3KJa1r/P56TUQzMWRlzj62m6dDHANONBVtmF/3xYAr/IKdv71T5MLT/pBJ1xMGGX
/zYZXnuaOvdHdpMC+In+UhikDi51sXaDG/YtAK+2z+nVwote5fkar9e9fROiiwVm
tU1spP98oFVewjSXuZL0+XaQsWZltrJHbGpey0rriEOk7Zfk1Ylfiq/6DJoiofQD
p+YHXsj3H1yFRXzpH8YP06Uzxif75jeNIQ+ZjvrcqeltfOlXTYSaf+O7ctwOy1BX
Y9cHVGIaEr8t/8oFDTebQ8BZK09h3+OfYKkuRnqpyIFvQl+NQTDZE6gkEkeHmz+F
fG16TZ8SHHCTDlhRz1d2fjltbX8FRBtRfWxQ7aRDEqj/zfAlfj8ZjpGDeWeSF3+o
N4/LRn7EESd0YysZcSpKSnhvrMKwfA9Nu2OYKCHGc/r+ZMYlckQqstQQK2vnOzPS
P4a8XzoB01CtObA7ENlirrl+fxUFllWHdW0bEwUTGebUWzcKgGE1xaGG6PoeqdB+
YZYTRn0o6RNmGIUuDgw/+orWt6tu9R99UI5A2Sk56waXiJwFotcvP18eRaxlKIgR
p8mKjD38qrWsEI5/SclaNafRV8CUPdQ52RKvExXEaas44N/4JJ4qrC8ILDdzjKLO
0QJhKkzgwYmmdxvDioPvqwxak/xyNUcKz3PPZJzC26cYgS67rOQJggdYUWrNtqbl
2V6xEjXKMeO9tJ8VeEc8y+2WjwgDYccjKdrT9RM2i8+Ca42kQbN8G2MMGJ3ptF6x
7nnonrW7uyRDsr2UDTZsg6AMB+NsnTrdBj2MdtOEDpzui0YTD/dAdAOYVtQy3Icq
vTtREUhdQhsH8HDSsQrNqbOTyAmn15yTwOLt6jClxTD5DjzzMk1yQ413W1QKR1is
q8xoG6eHhqsCDcPAR+///VezDsZro7w7PZe4uwMKHKj1s1bUUvPI1APSbbpeDiks
HDzUIQvcyqTZP0+DmYGLFfnQl77p0PkILWfVn2TeMlGfp3iZF9K1ORbxyNWb8L8l
FD/Buq9zjFczxEm304mj0ZYkJSqmlAgQLZ0yXei3f0kzXT8YdjGPwvBzcYHyy0F2
RF1TboFvgA1srjCGfmfrpYY5OekgwWvPUYC1CE/5YUm4Am1G5PstLu7MEWSndbrA
SMX6klAhwDNp5K7hB81PFq4f08fzOJUdnD9jQgOKxP0V1wxG2kcPT9LmLJqwhIuC
XCWvU3y/Qy/REmcrdoMehnC5AstAjsRedNzCPou/A4XJUcDFDZZJ/X4YM7m7OOZb
NF0PRfHxkspFG9H3TcX+d8I6H3UP4xa6By4rPzbsPgX0pqFtOfDZmuaMUqYRda6G
uotxBYgrcO6qi7GRm7kezRAXXweKOrNBdmoW0MLUAXuz8WuZyitvNig4i0ePMUE/
z06vsRTQ2kq4fd17TGUBfomDGHXOMEOvqPenKMX/vQZWqE+fphd3S7zlU79ROEEv
QSV1VDDeKd6irFonCc9N59RvkTWrzlkvkI3hVXiWFOzpXfwBe1DjMfyhKuEwnqA8
0qpvyGQhkg/X9LsjTW6w4Nz/R/NkVsmOF5WMCDwAo1SOqL25nuYHtfhDLZgrrkcC
d5mPXtD5g0qkQqjn2wkw1igO6mGS3cqZgupEC35W32E7CKqJ4XNx1Kmxk/ePIWdR
whL9ks1E74nM+WpLZRpZxLwGxNcs197CwgTso3yFYDaEuuVGz4/vrJbDwnlOZTiO
CMdsiDiJmuVXVUiYqnggBnlaQI7N62KFzljoujWEhpKHF0lwg1x/sanPIO5dkNAZ
TDMG3uRbyxz7qx45V/i7OPXipegCHzlryVWdP2u7tSUbZ1u6I4u6/DLO/j2NgAlH
NsHZDtsWbVzIR61FBLS0kAmvLeX6NfPP0q1UDpXssQMB3VlatVSo0X1XmhGoJznS
Aj2eu2UKgVNaeXiDS1khdG/il/JB0gNGk+ckZoW+7zuCO3TUAFtjNaJRD8y2czVC
yLL9C9kOFhnjIKhgN4djdmk0ueKMb4p7k5kKXOQNQ4nJwL9Kw5OoeX4r2AaZGcEC
Jx6NY42wnbX00WsClC/4ZPkzxqIXI8Pqq8wjK/hi9Os05dpxGw8yOCrK7S71DJMo
VEsLz4S6VfNuGkwUnab5i9EL5Jl+HvZrgsueuwhwgD5+ZLXCdgrOtryxpxrHIm1X
WgyOLruza+RKAofLZKzuxai/5Kzd67JK2kd5VKNVwX7VCEe4e8JcPCLDU1JIXqX9
xS/05mvWZRZwPG8qJ1nIz3RcOJCokmpgfXv/wyXATubkRzqgDyiCOgNVHWyOQN5w
w1YTzpaVUbAEMiKlQUX1y+YthazUjM960dV9/DsYkL+rR58oMxGkNqz2OMRcMCxn
04lDwzBeZ4Xd/aVDuLYRRCdr91lxpoP6v0TyrafE2PfvSwxsOTM7ulPBusfcASlO
t+6AvMP/kMdyJnjOQTLM6RHIsu/2KGjMGkIfKXn0HQJBVil/sGi2Jpqu1jKwXUAj
sne0SOcp4KrSZGJfbOEgvuucSJpW3ja8hTEdvOu1FhH0JOZci5tMe/Dm/PIlGT+Q
YpX1oYVdhvnWyJ7nzcibQoeQ48CnEg1VsyCiuQy8kEmsjVWpbdZpais1tGBua9Dm
w1FxE65quuUgsp1xPtdFOva5ZkI0kadreUJuFuP0nktLzEr1TbjvY6yBlNV8lHdh
auVnQPAwTaEout8vvg3AU3VMo1wNf16YZyorRn9Jt20IVPAEw53nUu7sbdx1ILsU
ycdnvoer8Jca31kpwpmNZUWDVdLXn/rPnMMTWCuYLarnCGXn7OD/v93Y3FoEJcG+
DsLXoJzJOJaAUwS3t1M6Bizt5g9BOM0cz7UBf7rFGEbrxWCZQS8iUIptf10//V2A
42ex2MhjhC4wQIhQYy6VmH8ZAPIqvJHaLBohynIWxMs6u0DYz4Wjd1HpTQ8AVcNk
nWjgxJIVAjcHd98sqeyBuZiWvOeFWmYWN7ouXzBuPtbnhZ2gJy/NU5geopE6bC42
XKx4tu4w6H1hha+Ne+OgXpz35ZerNxJXeJIHr7OdPe7AgrK1Ky2KN3Y+FhtoNZDb
VQbER3yR0g++3vlzabTwm53L9ithaJHrfDXrYJpePzLiep/OhE3LFQkNJzBsPaUC
zLSzcz7mGYBMqlTnkxX57uSOuDKo/yGif4RvxsOBlK2YmybBee2mVoOBtn/CKTBK
OIcHkgdq/cmpMBwsg8q6EFpW5cyQoAYCZHA/kGTdU3rf7BeUINKgWor7vcnFnxyJ
Q0/lXKt6m8eysUDpITdtRvSk3IFSsbvyq6f9W7RdMFMKNYXOWUYWA/Z9P6QY/4GQ
Autw5bhljOLtOo8PfZINYDIUsJm7K03B/ZoYjaHV5KBCWK1RuA8Jkb9tsgJePm2T
i46ejkBdUFncCvFrpgEU3+bz5evDIaBjY6cDtDhOnVHvUSFXAKh9ZgsPZTXFJ9+G
34oNStn6EDSrhDWqQhtl4KZXclJc1FiaOO5yRbRoPl99kaKAe0LkLc2JczeNaaFI
dHRW9SvFmGXCNtO7OHpI3PFOzcTiRJByooxs1b0d2z52GI1ZNI0PCmtgYbRM0MZY
df1nBIXWw5jfwLVEIl947tSe8s0uD7yFNYSfQQ0ZmXk+Vx42yty535Li8HTn7nYR
YLItKLo9S140eNFTx2qgs653zUmXlDfWgOjRFeQ1YxzuHe1WYombUMioT60cAoYa
te70gl5J0a0z/tqpybVVY0k/aySFFQEhnJMLifgMRP37vxQ1z36wcMHFRu1yVwLq
otZJ4DuqrlG8ByFqucxL3/7A7eifqZTK/ErgQR25W3ZviJnHmscJmS1jgJeI0Ujv
oKm99EapBRCIsZPS9w7OJNx5ULaA7JxpIkFieP+safUWmhpolZTwoof0sAYPc/lY
4Cj8k0BX0dMLXQDj+OxWIzT1bYMFki3ZhdYe8hACZRU6f/wj39pcAMBscS2FTBue
RYqnyJhhI0qPBcsQPwh28dYrc5ztxUa2tlgbacz9wi/3J64iDWdp5gfUj8OJ1AT7
9VNMHYrp8A3XhRg1nej4LL7WHOlLuxUvdkutHrY5rlBms1EJZnU+AmKCg0nfOA7P
sG8/JZ+mqFpkD0V0+xOfRvdQylAuCjOvTGb1d0GQHtvr1diAePpEQtqS9tj3UkL4
EzZCN5tUMeIv2eijry2WMtiyxiAjyv964AEyhPsTVPJk+POEVnNIi3owoWc+oc31
ZVPc915xkuDSanLRe7wl2a05flwKGiqFDp34EjSM6PwtILcaPgJKO0yAAoMld6re
ZA033RZ29S5rscKHjQzlHH6Y9Dq4Xwk2Pvj6Ak9y37XMKdTg73MymHPJL6/9c9yA
X2JbkgCN1qKbeRuCps4mRaF1G4muR0v4ngQTm55PIPya3DYZC5nXca8y7pz2pQ/N
jfVCEPeyySaQhcsVehhT5ai8zxQW1KeUOkf44IKyBESV8BeHqoK8mPj+bMN80D4t
CXOh7DHp0itPXF1FP3KisKQN9Y5OvISiZPcNpQ+oQmie7VRDevmJvO1v0uwHjBFN
TMSrxE43gWf7qQf81B8m72wAaoqyoaPN10Cztkj18e5MXPAA8ZiTf1VYiOd6Jcho
ItFjRD8ieefNm8/2c0FytkeQzA451PzynFgnVeFZ37PD7ejaLRFgsdfh9Sv011IC
gM8z8MsiTN1PJDltlBX7o+xed2h7G10Tyt3bB3KCv6VIJ+ebpiDnxYiTltM14wbw
OdiIWPgkhYoiqtPzSSpyNR2I0jZLSBfjRVOAJ3ODjSIScF86gSD2tPZaM8VVPcgL
43U5KUZy/5l9zE4yokDOyT3FMiLYhKQoo97MzYw045r4HxqcODYWA5q0x5U/FSr7
pP36oKK49um0G9IGtP1IeUdBtZ9u3A2vcmlWtMWBEcTbV43zyuriPPJ8bPdLVowb
lKkkTfPHMUhqAPajgxpjLwN//g0ViWYarDO3VJWaWN+D6qmQhdKRoIyfcIpln5+0
3W3HQnomj1UQGdrgP1JTu6EMLGgTutkCNJAIahBq+KNWSknFZvVG5iYUzssh6shw
eDkaFe6KrRtzr4BG6yBOlqLhTTYhd8b4LFMGrJFoiXJp1lei8PYDrzxYLwPdC+Jn
5goCg7vDjSSsiTlkcTdpLjzbkeeJ1851eFxcCLFv45XNCHU/CXha1BUqVQSsRlfa
JEIthly7EKDq9NGdfJDTyW62jLGdiidrhCMCORDiOk9LgGv6qb3aNwnJTXvc3qbN
R7D9gXZTHlw65Tam/aXX5D6LRR5/bTdCgDmr1bdUVVriruRCVmiDhE7S1aaBgNg3
BRImjqGkk1vFX9UeUf3Pb/0un5eAB+VrLWHzNQE0hOAxgVOC/k8t1jEPmm18yimU
0/VSjQoZAB9q9XA1+zs0dVzxyCN157V3F9EkRW5I1toEBrTRbP1Q+HCVS3KCNfxn
QXvcD6Y+GSQzxUuDC6jh4ayUEaDbDF8GcHZ2V6XQUSVgbYc6dxTy0Yk6qaWbo5gn
n/O+RxtC0VVkNvjlN7jcV+/ctagBPVQ4NiAoRhKmRkgIET+qtzb/LurjP2VZX4ex
6Sjqa8OOEh3rDzonzphg/6DKUml5hcJIZQ1DjpmZCrY/7cNlGoj0Xh6isBWwY8nQ
7sPlPqaYRJSEZtJ+3ldptnkAtjXiCyWoYsKL2uafBsVsFhcJWQ7Qq/GaFU93P/VQ
UPd6jxBaGSzKjMzswq+/FuPwfzQA9oPoKKfXl+qZ4Ft8B/1DRd1pIs6m09QW8y9D
u9hrxOY8b6S5ag8H8QZkQkhqNam1NqHRPsudaZvZfrThi6DUbNouBNnJWktaETOM
MZBpTwDEDCjE+NuMo9uYmVhTiE03/0YyLXaeZQx9gbTa/WRKbMS72HeGme+rABLR
NSsRjEa3NFAjtbzmvNjZb5sgJUtYsoRgVDLf2r8uCTODcXDaYGmc0SBsvgp0gv/X
f1ac392nl0wYKxwXlLMYY0gIt6L4yrCwMvN+UNWwVB3LoEMMUqiJPkdaxZDNENI8
0aUSWB+9goQiU+/jqukj7MzPSWhoaJAvyI7+G/lxHgGbu34JYcFb6FAq/Bj0lzCb
VzY+bB74mtwwTPOSUYGesSEsXiXc6JFxSZrXvSwSO7zHvrT0Pjc0m1N+9cn1jVpq
WfLPwRPywoG8I6IkaAGlKtB0JtvGj7K78FwLdxmbAK+Zpa7s9y+NFuqYTSvByI4E
EL3hqdFKJnT6pxsRq6Z+uQlYsLcsn0ul/Hss+9sCWAiNB1vbn2UZVD1X64D8NkES
ibaeyVnX6VX/eTS9Ac05+cGcKuxcKZE0e7VHb/HHU5N+J38cLr3b55V9MU72IDn8
ufbsNO15l8eCIGm1LSrKOOEbXrCxPHeyZPpDI4LQjnUF5Y67PHpzMNO1hcngazvQ
6tGL/wPS4KP5U83LOTEmZcDynEzmk0jtXy0FVtr/G8kbTJEB/XTVIbvScoXvnSBn
8wI/28F8c2nWR+bmaL3ztmOHmmm2wmwicJtZK9ih/dKg+ja3GgUbHSXyGq/h5pRS
x9Q5JQDihXNdZN/YmkVoCP9P1WdRHk8PYx3w9zD0QREwbA4x5fv7F4nv3dfEnjMR
6z9GNXfaY0LUOuTwYP6blnM7c/ZTqgyD+dMkjHtnfeqOOpgERDRX+58qI44651Cj
vG/kOKxAlUN3QNMQg7INFD094QMgqJVNRtE8d01KY0X7lg3CMCnrpsfMSFtuirg0
wgrH/vkYOf9n+OfO94dOiaidPPkQeEbNIsSoVosq491v3v4Q5aaQ4OUoM1N3Cdxz
YrSfUPqbtyHLRVmnyNMf92LOUBk9FMV+Dnk/XYhZyNfzw5ucj/4qvocHBZG9eh1R
Tcg46RXO7EQo/V9RpHmhZ3zYzg2txZvw6SgRYVXY++6QqM/qqd23KDcyo/d4iIXY
4KO+pc1bHMkvi3T/XHuDlmePj0crUxUvEZaHuYvAiMDM87ql2MklnHrt2F1ZC4Vh
gyOMVq/bnuj+SRRUQwK/ykyhft+hDMa2Td2Du0MjMsCp3jLy+o6ktd4P9sqEM7gC
IApgd3wRezr79pGU2woULmq+AGkyX7q6snlKLYMmyIKmW73lOn83GvSe209nMdva
k+vmV8rKaf2qhZobD16sFXxQICmx9GPD1ddGw50Jxa8AHaWF830M5Bv31XhfZeft
PkhwOOmubaAV1k9jkCkw9qaFiUH9bEv5Q+ta1/TolJ2xHpxbFbUAtE/utZlC6VVx
jHwlOALyV3RlVi7vkT+THoe605lUUyS8n2h5+IXMGBWf3dguyTFs5zoWLKdhcNNH
QM25tTe4Ik9uT2gLabtCUq/2zf447+PzlRNmr8gqGJo7CpQDdB+YEy6XQNXjS7P8
Ofb/dSTSAmgx/kxfUd8Wn5A0s+QX9l/ZJlpaZzu0FMp41cmb2iEqznJ5Bb5e/ufk
GahY7jtkfJoVuxroL6sbHb/DC9+TMeJl23deSHg4aFOZWL7i71Y3qqP7ejFArkoj
ZDhS6tYfOjXwZNj7hlQHwgkPifwoBnayt9Ql9unMvJkJa1gznqiJ9V6AYAIpEeXo
CGpN6cU1Ed0gxB0+vwIZ4Cj8i0+rfEU1DGGcHB8XhVZbBIJtXgTtOnDNaycZsKsD
BuS/mlmfH8QT6BjOBNLxskjvHT6uP8NbjxdMJgmduPXYFhUGQtBIR4T0fP4YuCcA
nHo8t/eY1qcXk0sQ4ImCJPlV0u0rgofhO43NJEO0BKeVRf5Ti1jNG+BwX1pk+Hd1
vxpAyNP3K27T6muAWJpBdmXh8Kmb2J7owQvaNehcJIUKafK5B72GxQ2OOlqo0e6S
5wybhayt2enjFC9a+X58MvViymWDaMAd8H42PL3CmZhXNSVb87Cp67jVMStWec1K
GyQlFCJ/jCukX93zRrc8TVdpzNmRJGb3jOg+yWAaNTc04Ks6Ot4/pVVily1JnBsl
41RrCwa6syCIcp1UpO0eFDnvgkMJVIZipra/QRDTIUBuyErZJikRiI26WEjBlYmH
K19fEdPcxMWmM9lfcDnUGuoyiAPFKUDFwBtf/bSnxiIBka/zqL8DmiRdEpaPVS1h
Q0+LWv7ZPjZHybfog+Pj4jqvmitQ89KTPojVT/yROAeU6Th1R31ToroBWG910g6h
rEaPIsCU8VM5JIXjejtKCa6g2m+Sh8QThBzDQV8PqZpriTw9Fg+I/jBzniGi6dpv
yxl/ohHbmOp+fQSsHbomFQCwQyJ98fRkqgQLFLQ2qNMoXua6BvRwrCdyw7egJGCl
cUYd7DxrIMIz1bmZRNOM9BsDRcPtFW1ab4UFNRj8G1yiEiknKvcfNUvxvctPdDeG
sc3a4EeFiLLo353JDYtFwYjfX26NphrRP/w8WCuZcW1RlQm6ldOWf2UBgem7PID/
grvy7humVdwDLKlR4H4Fs6Q67xrERwL3yT6rvxkIg5SWBfy79ZPefaA3SpujgIf7
IuYl9Avsk/MJ6uffD9XwywdGiLjiWY/PX8LOk746lqx1QUyJ58Z7yLWY+3VlaqbC
mg6fuaLHh9ioZ7PKKKeCQMw24mJmdDJruOWYQXh9KSVPdW+J6SlBDETWYfWGWnbs
iG6eBRJbw1DY1e+Tna86PpF4ipOJWBYx5MMrf//EHay9/IiwOjVX7EV39GhjoS1Z
qNR+CwDHbGlEihQiTuMLwHE0XxaunG+HyDD/0FArLyrzbq1ZLLtdxk68Zo1MMsLT
10Kl/rDYNc09dikHod2eYZWn0MombPLgwPQk11mlWBcZbCY+G8JNThSe1UPjzVh5
zFDO4sqMFFjdesJ5iA6IME+zZ8p2vK/RCmbwuDTPqJNrabIEgJiPYqmFQe/AyWYX
oUpr/hhtH9acqqEMZ4T3WzSMX51yhJ0WZ3qraBE/9ry/LWlzruMcfRA2ARWlvWzH
WRElQYni9PCSuP0oTiBVVABgR8yOg2zNukXOTcBhX0TCEWjzkBPQQOu3LG4XdeNZ
IJ+yNgGlJ/+WFYSk26lU/MiXEwx1nyJmxDcDDk9JvRwRbQClINYVRxDM6sNLbumP
Gc0F6XqcBTDx8Mk44AaKeuP18o/WIK403d/E9dQquGYrcrDxe8XADdL1wR6IyhLu
O5hanc/Ogpq/sRnIb/bMmAJNQJervDGNgMGI5PsmAaW5YWCbWc/89da5E/dfpjZ9
555Nz2od9v816PxE2v4EY2nRoYx0fcxTqBR3Jdzc8d2/vQVqXDXrcAdidXlm+YAv
mwpZAq8LrY+nL4ffnY/cRxneX4XsCCRBJhnFcf3lpWryUB6h0B0AntTIPQJ/A4Wd
87cMWevVbox3ucBnq/NVo/SQ+QFwUe9IKfWV+SqC85Xv/EH7zISa853kZo+I0ZDh
oJtUSXJAabzEsCIAs8HgLYQuUFs7HBkwIuRD7N2RDiYa50GT7LxT8RDhoZLrM7mm
8Q82XNsW1DppZwE6JpGVIHe/ueCeYs8EWK2lVEq0qmc2fZuyTAeon9NBjOXs10iE
SXEDGcSrbYjcu6ltP8N+eg6/34q1idPpWEIkW94/rjfKWjLC1eH9kflAymwcso+8
NSLOE4/KKNZlpZ7Zd0tWoro+XEpz8CE4k0P6QCv/txlmgwdWiUYLDVcF00vAh3CB
wZoyqCAEsX6TQhNqXuq2RPqi6gabYyLpuTh6u0gCxJbC4dVRB6jNmGi66J1XMYUJ
N5VFQmEU45B82c2daoGUhdecqlaLAtQ9rAlEOkictjG/5vE69f4mGiWOA95U+aT9
iomhz0Gu1VygzFWEsR2zfVrjzZCBTXStKcBEm2NVq/CqiZjZx+vbJB6VlpSFANOO
65aLS9SFqoJeRpqPZC0ZLFs2mhEEkoEnWR7E0IOHvFxybTH6Ci7vpcDyEDrO6H1b
Usf01JSQ54IoKFQpD+cajk+l95IDBErzR9X0Wrt2fphda4NQl9nfT3S//LEVuamM
oH0gu13Geusxask4p98F0fDub/u+1atuZ8LNb0zPxOWxdXEnzE05EsNs6Ba80d/J
g8LbvIKyBVE6tJA1NdozMZRCFDhVMqRmKbPy2/9mfXj9fLACqXsmV+yQ9/gZr5Uf
G3rDrahf0OxFclAn2zPSENbbNHU3NkDnJ9zH23BtjAPyNhwDHFUa0ZV6vy5jMuTO
sYRRDGKMkJzXfRgrAB19U+gTb50XCLCZWoilUdlROVMB5leZoZq8mYnF2edu6usw
rwH4IJnCc/vWaqRU8iApTZ9j9ce7Q22qq4LftPrmS61vDaDoIVJ64vKIprNNCGar
pJw3YQWC8LCJN07i/bbmON2xZ+GF7qM0K0VqD9Jm8Rz2pmAcwl9aE4GUE/C4IMAT
/HUmo3sP+ZzU/f4nzu+6vMFRSWH9DpHj5Pssy2BOFHIYtIbo6Zbmzbsso/1jy+Pb
x2LKK4U1aGH1V8OJdlu4Ux1hY8ESG9KLnajGRntJ6vjJUpleh9S7EqmmYzsLTQYK
JjZJlljQGrlntQV8TcC2/dJWuqyhI1BLzXpSkaudpUjzVI4n/mnQStowZZ5czHmf
JD81N4MQv+7iaeYFZtfzz9Umi6By0hJ41J9fXpdDQMHhHuWpjuLUxQCrmCsPpVf+
qtWVLM76cF1dbyW+WjpqTpSi000zbR25hp118u+6Fhz9qQ+6aoaf3EA3flhklxKb
wZ58Hq7O5XE59iQrwmlS8dl+qyFDyuh/fnJ7MG/+MWMkfAo4/jcDsn9pF1C1kt/6
VsaTS8RNpGjMZYJuuMcdnC+HLl7XFWOZxbxn54aINud1OVncPUA3RfX6fv5/nLzM
ZH7qRX43il0sT7FYwMTnyjEmksySzS42FEtD+xECzTN6QwClJfz5PavT2ElA5Wwk
radjCQsbvlU+lN+ckP5uvewqzrK0lhOl2v7UgrdpDlrFRBVQi44SqP7aWuZvuoq8
HL/nFbj15B/hqeIIIw9SfJnNVzvIRBQcf2EMSdXH+vDTyK6LiR8H1ZmqF+aKQMwA
lme6VBmljk1rjiZX/AAOYU5xQpIyEOQwmoz6vSy2M3dW8OBEs+Swq3dG1yPeMGSx
e7GTvZuQzjPIBpP5/mQOE1GthGgE0DAuZeP9z+7FcJclS57kb2Du/SQD3USfdYNb
touqLpW3bQPjQKMlieXh0GNK32d7TvQBuMqSBQEdiIM3Zkxq8gxNXyHfmc0VmGi9
FzLkHJZyPS1V53+QQ0guummXQ5zcSBYyXTFi+UW+rN808Ozw3+zV5NOs2LzvHulL
+Sf1fYrQ7G0MfqWuZsGcBwDv7kpu9AfGIBZO4T9KbEn0GWq0bpGrurDnEJosLWx9
/TFjlFijS8omgCDl7RqGuJfBynR9ME9GPJ42K6tAvDsBfj8bInBrhSxo9w9k8+bM
9d/esjJkUrFbKXVGHgFl/Mj9OErGn2rdj9kH0V09gg4hwoR1+CB82CItu3pabJZl
P4d9FqwLQ8nuK9M6gGmWy7xdcVM8H6qe0HJ4WnfHnTMDP6i6En/orPl0J61fymgL
rxZw46d1r9n7IDkY7mH1HhvYcPgLQFaZSt7k6JQO1vNq5kBSzdGMgrIJtmuSdi8q
LLIKDFg2iqkiUJBdENxJy+NAX+msbxzUHZxSz74ANRcl9BQEOI4h74h500SxH89Y
boraa/ot3PMdSTK5T5OPx1SCtuOkjFLtmIzch0nIVZDHkzffogQOyQrX2ua1daDB
rp+CvCmfSt02prSBLcq6CY1i2E4RS1Rk8wl8BddAnofybjeSNttlLNmt/v/cqy8d
QETk2WKAB6Ti5LcZR4YY/ksYp6hHGW3MZ+X+JxMw3uixzq9RkV2Taa9bCY1hWwXq
EaTFQQniJZ9cGbQ3OdiTMwU7fZ3weuJPg/tIWO1jBaIGRyOImpziNnjtsuegMNs1
474au4SqepfCCZb6K7PZbeVpS5LzKUP0WEJibiYPV3+tUWWrU/GZ13TX/bmuIoNP
1JUuISYsIduyD7e7tNezZHzuaoFWkY16xei46dAP4yh27LDOYkOifp9fHPla8gbt
R2+b3y2++ooC9LZLRjHX1H16Z4puwwWYX6s9C1OOn8TNf/RyPTvnSUUEx20rzw8n
I0Ewvvx4i+LRQ08FitTaTG5sRtoEREw4oYo8Rf9GGBucnxxijHSxqonqB563Pr4v
vLy7+jwQrL9BS4hJIzUd0bACn3vLpoi9BzF/+7+/kBi+xSGzoQBuO5ON5b2E8Hxm
ULAufFFLdtDYyexM1D0eqpNiG7xtSzHBWD0x5aWEKftPSQFCr4+wv3rH5d+0fzMq
JuDxFBGFTWbjcfnsv0vqNpQHM7rQKwYNK0wbcRpj6BqwBlmAAmAcZ85x9A9h7L1T
1fwqr5lumaGX4MvnnhnVKELQ1JtWvBRG2Ovs96ifW3yKsIuHSm1pki20glAyGVMQ
KbO3zr24y1ywpL5gwCvH6jH0nR3AzEDSEND0Ecm5O0tUvQESy9BPzB2YMXCpuDWw
OoeQmofe5u2q23UROC/DF/x5ZdC5c4ExkycOAqeftZojpyguk1jExdtjUI/clWCR
HL8D72XQHIsObhK+MMufSlUUnJXor6Ggu7MMiDZDYlKohorIbEWjNgdpntw5gAJg
JULAFxkeeF9bSA54L9lvxKuFkT3b0DdW5pVYxMjG6Cgyf5sjgg/vBu7jg/+6hfy1
5f5nlkuEyq/zYI64BgK82JXL1AqrycT3Ms0g72eLFB2box5oyPCHvbwWSfPJEekr
JTS7LeeHR5lFQ5FF4vEIR7dpMq3XBVwz/RUhOTLwxlN4pan0rPuN+jGH3m2tuDpj
t2DBFGsP1Dv8/IITw9Y+Bw/YNHx9cUrYlgVsqmE8DFNiPy3VaS2hv19Tg9vEllKn
rsYKV9d5ky8UHDmRfBFK0ZnMQ8c913CAwnuzxaHvRC1Q4UPbDNcSScC3y0TotspG
GLrgVO1U50F7S8aRbm4QnFgD8qw4cqJm6KnxYgNU3RbyDZzxL5B7yfQtqRU7CzEG
vMKnOS8vxvveotKurD+RZthejEqot0TNa1ztXlnhtXFj6P8+U1f70RGLyhIA2eAi
NsqpFtmmQaR0IwNRJDS72KYR2rJiSA2F/IU2blagbL0y42A7fOrHpQU76BVFx3Q6
+Uq6pJ6Py+Tu9nCta5jqxcBl+CzekkdhKFiyxEMD4u8zTpfLbTT1U22m3onqVr7E
XNbV/e9H2Ns3KDRtg8yqk2+2hdPdPxVJt5bJZK/3IaqysbwMDYMktgd5CUdjX3YR
alsMjPMsZIaZQUjWfz10nNMxEiTKQIej0Q9txelCPXA2TKpS9D9GFdZcbD6VDrh7
4n99rsNFWcKTJ11ipUKaCSlfcL9pT7+7dO89KeOO4besD8xSyalbZI7EeWN5uPgl
CU03mVAL8QjB6mFe5gwiLbC8gU8qbhdJNEfxePPU633YPCUZOgb4UYw5cVjVq+G2
FRtsuHHfq5kuN1zLTGHOzKrJVCAAq1uzlGC+K28zfPdJ2bD+zUC6c1VxLqzPNgXh
6atk9uf18D6aIKkhVO7EDBVDQG5EbvN5rXuhE8Pg+4OUKX0SmXJaSxdLE6DENmnb
Yu03NqTv0LJPjSwtZNS6/uhDOcaDsbhpqzw1oK8XQWB2nr/IRNQFSQeMKFJ1JHwN
AJiMrg6avwxISP/ElpBStBMtgFNgFDpYYdFlEZB3bOarPYdKwAkRXhJ1OuiT977L
8gy4hCRX07P3Dv33t2R1FFhQHrrjq5cV/GYzEAiK+qSAS9tsi+WqQ7/ko1/DBcAv
sQzoWWDj0R/I8aFBRCVuzkfWchSJ/pSon8oAtETp3OoHiTBdxO/NOqOkoghfA2c1
Er0vf4wUhygpeXm3Xo76pF9k76YpiAQ4cLAmkYwCicEABcK5GdmOVB7Vl5D+gBoW
PxbNxxJ22p6trzgsJpM3krr0P7FApdwQu4T86FazQ3R+dREA4sVSed9Wb3/5fKFV
YvwQ09Jf3BSdS8J0mhdi/W4r0dGKaQC+Pmb5wRlqENtlf6v+5pBRkSFw3ts9Rk31
Bx6UHB2avoyy5+oaAQdyR+nRqq4/TSFkqv/VKgzcNQ9cktwyesyz+8UGGsF9ZWjW
4wDPI2k0R69hYa7fa0TXS+AUpQsdzWiCZ+MI/2tueZGMf4k/OYlKvRsmau+gJvOX
ZGHv5uRaMw23qx1T4RgS0oISnJs0ZTGRrejY9UOMwpiI6iTpk/K9nLW4MYxtXK1t
Y4+z54Xlb9pAsXpMUTSZEQyzk31NaDFwo1OMj1V+kXKJ+BLs85AFiWRRVuhlL5wZ
d9+mpsQx2aTH33ijih/01iWoiRQyPNSx4JoactjY24uJOMjrLuZHSyAB492y3Z37
Amqsq6yOn/J3f7geNO0+abbYpZdyWwSaZszsQpeD3g9olGDFnB7YEkVBDNLH/Yho
DYqmZsPu4IVumFr2MpkWR8oe/0Ahwp6CfbNrHCAKJDkq4acL0zMfiP5YXTX9jZVF
Izohm7v6gsJmDOmdk7V3+UCwXlxANGhieDddU+/BDNe7mOrXY9jJ/p4pHs8ZkFKS
AeSC4X1DyQAwSoJFlNv4cNbeLyG8fvZDx5TEXYiA7YHTxL4I/7OE17lHhJOmC7ow
ehsJ5aFey8sVrtbdxV594Kfo+xCMokKEcNymo7EYTd4Y/uk9gwvPUl3oXbCaSLtK
vEkicuWe0dqQGtMlfASC6azOuy0AgGNIRIplnS703ZoCJ3XQhwCqZblb+wmm7bPe
ypGtdoMYKcrBhHSiPhpcybqjiYydsvpbtIDvW2g2t7bJn8URZCFABqhLBx9gtxWq
8mk3mb3HE96EHypapJK3If4Sh+Yb4H8bzpOelK71fZi7M4aaPBpZRKNZyOf8GkNF
A/YFeBZRHaF47szbeUywISX1lITE/dnS54Qzk2UMPvGs9Mc5wBYJ0ZC9RWEPOjbg
xMG561dTKTXrQbwGQqHBOQbRlB0M/FkHo1dJlvQeKOyoi7tFe31jQeH2L7wWWEUd
Ubo6v4F/7U5XMIE/rdkHJsXdfhiHpPT1NHZvb5YBUHDbHwEH5vfM5D7Idu4THXSi
snM4ToodEuu2ii2vyXKm8r9bVjpfiNcaoZu1DMn1jtvQsAFAbyh7KIa92l9LhGg5
hO7h9M1PYUJr7OR2indsqGClMm2VjWosGdDKZZ3geBqHRGUZRCXpR0N2hqQLDsiY
frsQH10WXP6WKjkcnYKeblmYDenV9gy36LzrziApvD2gv02fTZuDUUmzSjKiFoUl
g6bwdaZ2UOoXYhM5NfUTRPbrqYk6sBJ1cIqhgddMDF5S6fDXOj72vt8JI4BVvC4l
kQ4l/msVNsg7wYT6wm6fIRg/oBWDziFygkKTQf8yvFKm8kkOVWxewIq6q2Ki0pZa
eSQl1f5EfD4GsvfjTwh87ThFQcNkyYaN+EfiLYjQAfoJj7DRbsfncaEhc0TrjGFd
EjftMTJz7NCoj6d31GFVg+JNiSkqFcUk96zfmGzvHyOGYiIgk8FPKI8IaJQrEei9
X+zDtX8Ea0aml3rzbxI+4C6qgOuU5Bw17UbAyxNvp3aBhhuuvLXQo27jJkNfwatV
MzKbQAvgmiJYdCKh7EtT39opjbuyIYbvKb6rr/K1Zm4wi5sDR5kxAH9HR2DSAAGC
JUkcPEC4EWnbyme6h0/JyY1PumkbDXsd8XcbrtCqtaaswyT98W9xVklh3kWyu3pG
Z6PttZIZB10w24sxgGe+CkStO+7P6RF3MUP14s9B0WUmOpcxEU7KKUwJXwOyLgb6
AOk+VEPAYqqb7eUzFdx24WOfkiXT41ylZiEWcTNlKRCKfbOjfEGOFK+FoGZeB6oq
piUTWD7uZgtJw+8qCMer22Cb+MlxCPEMi74OnllJDwUVy+U/ebMI0BANCvuU7gJx
I0fAwYyhUIXBnj5Z7phYVCccDL/o1YfFpzNx1Q751UHbVxiWm1ZAQOjOI3uvocvr
a4LEJx0ww9VKvfoUHdRuEjNft93JSdF3zM5x4vBzh10OFpmhEwYQpqlXT5BcrGvq
IjJPpYwO4AcIV+thRb1UsJxeiQv27CCTB/KrSvZHi82uMPx/J9z+V5GUjzX4p9j2
ddc3wW2wOmZg5nH+rs+9RuP9MXjRFSXB8GIQT5C18173W7ZV3/GOa/kI8AA1mb7f
TyFL3ubbHN6XGC6wddlOXYDw8fWtyajTSlKBlVTCYIij2liX6X9YtKitFdp++7F4
oT5OocHANZqzoQJDKR6Bcp/pO18X49INeSpcyliTpnt2VFY+0Prth1jiiTBtWm5l
0idS3In32HnyS14HWV4uOjL4o4f5XjzxUI2gea1UG+a4/h1zkxKYE51cqqkMj5AE
hEi6bu5MfztvbxgugvJF2/+w6czHouR18AiSaZL3JanWWgCfSN71ucU9zrzlnHcR
oShzTQLbP8+RzAeQYEZz1Z+9ldqdGvEecca4pPrcmemGQr5wWmFol4E5SlYRAgxZ
lGhQK8BLdzR6ohTPvAnKWhOWArxx5l8jReC065HVR6PjBSf67rILDyKHkMnbfa/n
imvB+WTsrUO3pXLP0ygBv/uDLmvAKnOtiEygQyFJxVOqyWdONdWx6czwWf6dLqmO
eZbvkLS5AkEgoIcCxHBPPjvSvWipUjhhGPhUBejCU7Z1t6y8iqi/Ok9an7UQggfQ
0MsVvj/Li64BaEriyETas9b86wei3CkOlCKZQyWEV4e5pqFn3k98LALNuAaUTQgH
OJFE2qVbbMwvYptC8QcHoLmUdkyMvwqpCEhOY56LlZWFyTMvslmoP7hsKh3ckUU8
fwpZlFOZtTsqzWqrsQq6SQDrI/NSwOQtN6eNoYtPGfIMubcrfa3F3c7J1U3nZ/TM
2NUfALigdbV+KYqLwhO4muCk5OURunpiBlN/tgeP6QHgxqzsOrhDlSgYnNRY2knx
Rq+RU8XBSPrRe47JXJKK+Bht70NQ54olGkGDtI7VXagYd2UzJepfRAJsntB5+fNC
5m3u+rlsWphYjJEswJgTAP9NQ0V8Xtov7lqKjkLusY6+sHEVgN6Yg/pHoZrTXJJr
Olkfn8WNDDb4JydSPhnFGOjVCsR6bV2KUIoc8THRBU3mseB2ITaVvon/fNLqwdP/
lOa/lo+C1SXOjN+g9b8M2vtNJx7uXoKgx5R7oUiehuJKT0piwi+mB3/DvMkGoggQ
Hi8tOekRCeaTJRYZdA5l/2ZTYlSi+ahqn3VZtYdumxFZkrV/LaTMK41MZ4wbdlE4
8iT3l3oJ3LBVeMh6MSUoUIK7oo2dEwJ5pPKflq/ahioyvv6uMn4MpEZLEDK/4rIp
Le9LL52zWn3f+OFyBTbF+xav4W20rrUA3RVK83TaE4+fCvsquc60FCiQcwMHRIH+
W7W54osba+JwfPdcZBRLfQocA5lTq9EpyuMEIfEqn3YbQd/DpCyQWbpb6MKo7MHw
UNDWxmrn94jBLVZyJVAMk1icD7fFqKGjGwYqkj2N5td4CttFJea6J8huSlana/ph
+YSedjx1iQHiblMTELGQlDa364tNh/DVQfAyWMFekzJw7xaOPn0otbgmCC65hTEf
Gv95ZKudztgQsACe36HN7f5NgpuFNt9T5D++nCovj1kPNbklnSwSKOQHYxFSHQOb
CAINJtLb57VVQuypn4F0rB7aQUEq4JpW+BGArtFZ7/kqHSTXQ2MBZRePpPLofxHI
yVxEO67GhR4J/OAJmKbTI0AfPS5jDioxLA9SAs8B+2XGn9J/xzBwpGguc6GNAvzT
WIOCpz1Px/gNRJV9EKgplh8sO6uIKjEwcsA2IqyC6aM/Owo7z6Lopq2gj979mmXp
8/DYsbsyjHZyObXwaVGFwnMcRBRvrPVCWPMbYeZyRV8Wl+DaRZbkljOAoyOmbgyz
W4TBtFZLTMU4XxaaZgonokRQxcW4yDwyixRa+cPzkMeU7Rs7Q4cM2XJqi/p5eVZT
8qHKyJAI7jKK9FYk/agwD5C2O4XOpwJtGztx7OuSUQsytXSHMv+J7bpWWu95627f
RftO0wNux24Tz7kuY91Bqpw+8PXqG1dzfepczyjysSIZkdy2VbfelhhZGTnG+e2J
2b5oA5WJWJvTsSc7L7Lraj8QAJcrKlv5NeHKZlsA/YnRMRSGqfjKoLdjAd2wlNXa
S4pJN4RhIcgvYKaOIjdY5OvitYnHotwugm3uq/8E0b8Mx6/pP3ZNd5WKJdaQmys1
9G4oVP41adOjLZzTvd01B2M6B3MOCwqZwL9kyRuvaD9NmcutEnkCaua63JxxCCef
RBz9lBI9nbIWYW9qvX3IPf5TIMrdt34qx7t1YgZl5ixaXnDavqoaOOh47q3AULVo
zFI3z1AOpIO6opcP2E7/9EPAeyoFMGtPzEIJu/7ixH279lrmL7jKtgl4lHLT+ZjU
BCnx/g6JnrDWQ+4YTFLcQYIgJ2dGufWULZ4dwtLpqxAli9IPGMLdAiE8vBOIylKj
EOxHix7d3af/SyRvGyOJh+QfqUrgs7SQLIAxjyzKb+qxgYTuEufNPjlrq+OloUxK
6sCy9xpYnteYiGYItaNBWucvieJzaZGiqtjBndgQPzFQ0yIY9MAz85xxKlSm2Nfi
ai/Lks/PbC7A2MGNEmjBwheJrNU0CTk8ELRCd0e8Ipj2rRKBvrpFjdD5foC8vFWI
Vf/aXBJ8bd+z54jwHJwfcdyFjhjyW102Q7oTEKaibmA1Zm/A4aUfvnto6zyuCIXt
MwJmUWK3xJI9OzYPlti44ucGYLfN+FOxUTHPdCAIws4AkwOao7a/iDCmp8tG1GK+
nJzfdchczU71en+wQBClLOxCNOO4niK3XW870NriAOPyeyrDNNacFqyYMWeiA5Zc
ERP9h/0tgd6FFu4CHgknP6DTuSuDc8yY0RShuBz0Ld+s+Sk9794R1bYdEDieRPN9
hz4KlVA+fhJYNeX9JgjiPO5242agefFBu65IMc+P4lEC7jzW1AxNBC0SWYXMHAvb
ni8dxiqsrMXZRnvWklbm9Y8ZbLGoWhtIWLAZCxVVo6u55KKhCb7vp6bXzOGwAiyF
FbRZO63v3dIjSdkLi62vbyhIqEyv/lxdmCcOkAV2V019ThLg40Ai5XSkegSnrIWe
tC20Zh1NPpwCM2IWWCRR3M4NBNF3ufQ4GzC2bLC9LqJTa66lCz/xG5k0aQf3Br+9
/rZigbrPY6rGlmeULUVoREwTsMVYreUA2TrWaRSWZj9B8MeHF6amS8CtHgxw+4rn
LHNkfNSvY8SZUtBiZ3MT3PTQ72vLl/8dEakIohmmmet74VjdbZhiumBJBoPr5Ft/
85ZPrXwWqYyKFkcBde8j48zekl5cWxVYWJb42XCpsvoC56opbhTZ0hQP88MApkKc
5VK/x4ixHj4WLrVL7s2nSCq2QvJ7iVhE1VbbHFOxO9RAc2c72SgKPoubeRy+uwmk
g6/ax/xoYxz5mxXI9rMNDT5bJAQXLyExNEjGc1IDRvKnfWBvfMFV0HyxIahbmlpO
T2HxsK13NdUdhRiNhe/6/pFoMEjcxWhV3GQ2hpCaCI1tLB28hgCJx5S171O8m1vX
OQU3MTsCjjWGmRbhBc43vpubHvzHHb9CdcHCpKyg4YZifGyJuyC66pFwcINyp3QD
roIDuA4heA+T1I+jBJh05i936X7cJrz7DDXwwItpiaRzEjDm92nb3GFTG9M+JhPD
Rg4nGaI5ahzH/gMfqv+2SiZ4s7/wPQB0ag12To9+uPCDY9Pxq0qyVv4Ors6qnoPc
XkGekQgky4awiIK98OKMfsNCI85QVx1zzrP2xsH/z6YZ372Pn+/vlJwxmK+Mmqdm
laZaiVaK/JrYjr8+6Uv+Df7cEQhudsOmYEb8GSC6NO5NLKDmp9W1rUU2BhlBusEE
pZbBOSk9pmiBL5s/xk++Tvl2oBKrJY4hK1gjU51n50ZrsWf0kJ39/pxMwOAIhOLG
5s0tuK/BGD443hg6WQcQJKlakXJ/HWYIzjAY5q6ouxU/Vcv61j2BBOpdswNecLy1
qk0JqDxrwDXE9/RSrIoHIcDXQNYJI4nX5QcsMLV87dypAVl/NVQ7vMeqVL1cEzQF
DWvAcye5kNDDrLI7kZEI4SeC9qJImXRpMBY1sLR7ereIl4I57j4uydof5fvt+Zrb
elzwsgLoYTYwxGGs5xV0Pkz9kHdDa87Q3B9340JTYgryX/pqMZzZoZF7Eix5BClq
RLxpMAbCAIWx79gx+CIp4PY/W+p7VViIt8pOAp8yqqd+B1iW238n42E8JBvwVZXk
q1yDIrcvfHf35QhNSyrL3hsN7yT5xXnP6t0lj7kiXwQ/sRN+vnQquGu9zunW2QBI
zy0TACkNFMVb3mbJVo5DUA6w+AZU0L3eYk4MVA9f+azyT9ujG5hX32fwym0G+kjJ
l+5NvXoiGL1JbfXIZ9Krkp+yujkQwf3RY1k3QK43VZMHc6UxjpUry1B96Tzqwwwc
9sl6zwuZ9VCKvaQBfGqzWCWOP5pkQoOufpmeWcjDj2UQhbk5+8jW7D3l+7Yfcf4r
fy+IjQmMMyezYSId2sqtNamcNHMdlEO6V/MNVJqx5H+jYFaY+XxbQ9S+AAUTPdfk
iOvEV1+SwIxxonoshrvGLaPkr/wnwEjEpggINkkC/Q81tfCF0sgMj3x0uW5yiqre
nu4Q8IvctteXLTorTAk8jJMvn9r5ljjanJ2rrbuDUe1j4Fpz4yEHALLDV0Q5JQrK
34emWokEwAzggBQbOfKWYu0/LTF4wvIGOSmWV7rV0gqaFlFfJ2QyUWf5xHpaZknT
xlJXy1nEWZ9bp9OV/iYKt++gjKTYPzFHWBvCZXOJrvzaCJ1QJuTlVGhOAzrti5tZ
fd0XXTO3wTovC8NqpuRLgSn4gYEuRgh3jaEb/h9wMP5aH3Cv9Mi/XxR/DzGPQY9R
/GoGOVxDWy1N9yI+qT/knJeeMHbgpPP4ojwBiu05B6NNlQId/qmY1h7EpzIts2w5
IghbIrNGovBdp0Z8oLZ17mzN1ZdLqYqFWevEwuz3esJhJlbB6BIBFm1eCLNiVdE9
kjSOkGubcEcqI2fJo2C1z+wZQTaqjrl9e1ZkAXWAGweoVcB7ID5ZN71bwJ+QxerA
B4UyIfhSp/1kgZR8q64lOvUqe0FF/PA+TOidihw+CJQ46K3+9Y5hB4sQS0R0a0Yu
+DaoySg4FWUBpYm49NeIPtCtQub3Dt0xx6emHxEbzHkZmClwqNkiJQFCA/2f3Bhb
wWGQshIlKCLunRvf7ljr6I468ftN0KzyLJpXMhIifX07APXS+BoDj4QbTfOh59KY
jFHoT0wdmrQdH+E6LqCg63al2EIhgr58UlUPSvXDoMcl3hOR2WyLLsEirB85nxlj
wt+cH0ZMoPr1+JO/5ufGGSZNq7usFmdG2Lj6n3KweBfn+2y4TkNgYHM/5N+coGZ5
Dizu4vnRIbOaRXc7dnjA/X9QsW5lMPY+CtyNR71YDnhB//Ktz9U4cvNdZJpDCtnh
MEP8qItKjqpuwckM0qJPNs3emY2Fza/XQchmmEjw1HH6kmNcdOLa02obXLWv2sGD
dP2JDmI0/sLSL8VggZ7RLGDnZrSLmwwquqKvZgjkjxPvEG+s5mATpXQkCBTxGCjT
H8buBCVeblQN99yjPgR18Zu5VAZKCfO0vEDGD1WM54J6jT+ctR3LVBh9ED6GAMsB
fkX8/o9JXRMjM3PuK8icmOlqFWJAnYjOXVVQSBa9fBzZGCgb9lY+CfkQjN7A5FeX
tsbcgxJSPkV/QIVqBsTQ125TcyaX3w2yA5fZZnFs1RcNOVuCmTEaVbUKnrdrtK80
Z4aoxeC3xIcvXxfLU9H6KMQMUe293CYAzr6ZYMvaxMPYkxRThp3UjYraFOkPYMgi
e1vn1420dJchz0QJxBjRAS8Z3oYDeGKTRw0ctPP33ThkhwxDpewj6poTcjFEH9ab
4/8KXO5zNi1OqyUH+rrpToz/DWD7KmY0SMoG+JIWVs0HBpDKDUXwetHZ+uNhca4M
34DR4MPkuEkUk3z4g7qCzlyeeotHeNN/A9kXizvn1BbNevOkqIm3uxVBaQT/Yb3N
pS6EsI8piF5eeAaOomD8hmZFajCBR8Wje7Hb70dEqHWWpv/poCoYZqZYRH+HLVKv
xP6GI8durOmkUSOhyjCK7VEYAeRV6WLnOuAvtI0Cthq3kPXe4dzPEA6Bbb2qLDAK
dTb8uP7/r8A0jBgtA5IKi5JbjaUd4XJ+l8WDoMIZr1lAJhNUiT4gHTNOLWz3wX8t
JfCWVae9s+CsIn1RiJ8PlOB6ydZGQIQfrk2wDdKMG6JEQUV9GhFBmvafOVfEwXEq
NYwgz4wY5zjRYQjUPLqSZBd7haCMLQVsLSyGJCKWBCxk8tFVc/fIWH2cGeGPgo+P
sVpZ2WLWywFrNJwGcj410KQl3eUknmAz904P6EIP0OeW0p1zGoJbRpwQPzLmVpsB
YAaZjgLl0eWhKSN/eZBFvUq8LEYUW8foMUEhDEpDZDAf8zDzKcG/XYvasEku+Z5v
et6KJ8znXMSSNQ7C1/sHPY/qJut1WYYyBW2q6MmyACfDUNx+3v01mOuqPSV0Dz+Q
61baiqUOBHubqCKK5CzzLKRmIKn9746ME0YfZJ4cNmDlxU3RvJMQSzhbSc7WWgXU
SXTZtjquedlY19EQUrMTDkMU/UClIFvZzpnLdUBfi9HCSyBJiRjhBW1mZe+AxzKk
CNgsBSoYtZVnbwwRij4Sz3p4yOnta1jsXbQ682lEAZgF7tYX8xe33HOsO44auImv
y3YOGs6yu5B7d7G7fvWrx5COGZNPD71DVnfYlvcluR4nh+lNNN7b46wZglYZ0t4o
c3+wxCEtMFq939Dk49pdPr+Hy/ACyjc0ZXErQcyzcWNZc9Uj1BqTtoPCKXMacWmh
Zn1gU+3u4T5paG8tPPsQ/czt0qzsFIFIKfUasN6Ow8qtJ3b5b+zmPyDvt/YoPCMj
hIuwIpav9YV8PMJufqzAW6vVfzs5GhbjCZRNNeBcSmpZ6vDvC9LbB2JfRJVmqier
zFh9jiToB41faTmdBSUTvcGdnOsQjvqNd8B2lTN7IfGAMBcu9b1FYDfQWcF2qnz/
9du4l+f7hxMxQrXpJB7ET43KTz6nTn7js8hwYpN4YGm/wLByIp3pGt8kxZsFXyY0
nS4IDOcuGJKCvERG+UyoR/TTCzIemHaLOLIiM8mBFgw+dxHwMp8YN1gVXGpeq7SE
R6dXuwIYpGUI7kQOW8OPmtdNVKzhawNjxra63FmpmfRjCoPJe7O13U8lBe1Eutd4
W4LEfTRHwa4/9oucH8tK/k05TbQ4oroFt9vjUq2woXtTxfGufsLv+vNNq3bX+QoK
/Hjg0uf1hMiXKTugVQOD1M7TwhK6hOAOOuE389ZgWMQzpsGH/Vxwr9+F4j8T5ioP
LOn4LKHjjYH/PWhmt9caLjGkGN7VSGklHzOyHRZfv5KlvzbgD+VRw/kR6cqwDmw3
ezzivnawwdLblidk6Bi4QCl5pkfxLFJSBbSaVr9a1LPamgZHhzFKsfdloacTbY5x
o/wPV3tcWAznsco7uO5IEIq2S/s5jbZkw+92x5Dp1IkQZc0rYoIDLezaKeWdV0lh
zpqbSrzQgflGMb4C+vO6h5bg2W+2Jovm5WGw7etZpmalWeQdASSSjli9SgbaMRvH
bW9emnEu4Sca3ivXdqh9LNaqqGKR//m8bBXlTEaOiZsUOtSGTH8O0eM37vLnU1Nx
tIsjt/ZcZND3yxAfpU41JI+bk9nUTP68yT2hf6YLDCzDPrSPnqH0wZcOS5haKa+M
nqb0S/OF6xJw2P0UaaQVzzNbJEuVSxFKAe0Ey0ONWbY+VKX0G7Z6OzlhuFrq0Gmz
mB4MiaqrwMan2wnSj0IxvzxdSlGqBIQNyJWOyV+tElFPcGmzEtS5jvRKmUHDUhCb
5zx+LAyTrGKFFK1hJJ0gtCdwXdRbEK92cN2Io0AOow4UyoOkgVXvOdHtA6kfnnwQ
ijmv8qVCx1vMWhUSb6rWOQds/bGO2mDGjPvKfXnFYAZQtJYXmL1FVd0Eb7eEX1n8
bcI4Jbc+NW7QvUJccxMih5kypzuUqOUNysajZeALFcdoPnrztnknOjj3h5OigZFQ
5ZGhNFONW3Tr15sq8ZAlpOce+sQqFs/DSWwK1tQ07PQ8rZ6bXzI5t+bwrSNCjYKE
bYvm9vYnXLB0QucffrCyMzEsKYTj9m9unmj1K8Zk7qiv09qIcuJh1S3hWT28HFmg
1BtlRB0Wvnyj4hIjMxL2SiaHoFF+MrgLmBJdWxFxm2MdFlLyzDVPpIispoUUTD9W
cw3jFRGmFfmzlYYpAgdlTTNGyJH6e390jPBeuczNCdj+iLfiTfD6VE7UWaxwSrvG
FtudW8mLE8ntcqwz+WSoyu0eyV2PacSpmSycl+ARhgS7TewETR0KIPZAQJGsELiz
u/+2iZitmYYfyMOdQLesQI1Th6wZWVEndEXDtmD8g4C+eLknH5hQKa9khvjEE+oC
5Qc2njo4E44Mpk1mwTQsQTYkaCr48OmEDJ3iKypJwX+KyVhGSMof2dsT6GkT5HIK
YNS4mwLdwAINLOc9pIyDbePDTG/Gs/B5xC2i2KQpvMeUgDhDfFfqeGoxzO6+fMce
90Eh/1d3EeBppUPtMUabEHdE3H5Y5tmXYHezaoFfCW8gcOko1miTcSxEvHJusCTc
mr8XStPAXd8BY7PFeu2GrDV8ACXLA86rVxR4Lh/EXWLcNm1zykHUWdohE4qdGVLA
UUkshbQ39xLwr8u0y1a4yrVggLnzipOXPOU8hpoa3Q7sbq73FHPg4muCOo9EXQ5H
SG//WX3BYriOF0exY8PlZvS7LcobS1oq2cHIkPUkRNLzwxWwYn668E2SA5cUjE12
0YjbMQ9mCL2PEB4a0FRFVFOKzryxeuV+XupYUsTNCvo7DwKWAF7GblRboW/X5jpF
8rFp3yXfjd041QbWTAfB27C+KCV4Cs9KBjB9eKag7Yh68TM/xutkqv2+LtVnj7qa
YkEKyIm52i+FC+Ix6Tlii4yzS4mjz2S4f/N7UeJ4rVleA/UQigaBCsUmbQhxxcRF
x1EHhH1TVu7Y5EUJ3YJgXlg9RqJ2fMYGJqls9mMEgo8HvCCuFakTeRqT1oUcATet
qsJKcrTeKZQT3qmXYjgQfO8t/I+JorY7zMuVHhAP6arMtQjxd7RUZisMlSQqprmQ
WjplyeT3huLE5kKmhe1+m/aaddNMKGQAHXUS9bj7Y9qvrZBBVCrOM84a/R/2wRUj
yrYfWks/wM+NVvTV5bIAcieFrtBiQtpeGZTD6nizIj1c8pQgqXlnJ8pUTdrnMTlM
Gr4CulElCo6nFnSCSHGEsqSVqttGdlTBpCgJgzAZxMRQNE/DIK0IgsATZkP7FmAM
iF7Pl8f0aKjykbdW87Qjsnq0cAX+/N1XZgVMqbM42gNHWLe86JRkdFVTd8fsbl/A
M8bxMt+LuSg2ltIEtea6zJWu+LEcG1N6tXtSx4hVJFPPYbYh0/lZ2vEgjC7bPjI4
Zoo7/zlF2EUE3N7Hfe3yZ03BzoNT2dCk9QwxC8xWJiPbtD6FLoyrDGh8YSU60B5F
APqVtsb0+2MKB7Wglro5O8L9KWY6BzOd/Qkq4y+VPqlC+IXj7Zfuxtqg/rwekfs3
dp22iFOYzjeJZ2k/+DyIjBx1zzVft+sg8xydwP0pFlxnss3iV6Etp/CcZ3XMBAp9
a/4j9IJsjr4HOm+BI5aOFYOVUrfkjsK30kA4cT+0/Ko2B9XzxCYSbhdSZyO7RHoo
3K5w3yk+ngbt8Y+Z4cAhJKa+BS81tiamD36z7qGD2njhB+A7Qf92Ri7eTD9T3+IP
OaYz4/jIfFwrO71NPJg3SwFvXG5LAu5kGdKNOal4BJ60Huc8U5eJ2sxFQPswqZp7
yeZxIPA5ZLV0N1oRoS+buEGf4AUA+v8arCSh1Ep/i7TMZn5xojQf/4GhYk0poIQr
6FYKBTt2rgkk01GgEicxdCR+V379adkDS3xwpu+Z+tnRsJ2750FmKfifLlafM38R
RwrMIKTnj43ZnmwBVOxmnItAlgrHycjwaCkx3y8EtSMcVrXc8BPHqDEmVCA3WR25
NQgAfqEQetMcocXwq8R5Al0IT2LCzmZ3ndZgwrlWbhHLqAhtb2I8Y1DR+pcnZ050
DhLJCQIwFd/USkmmnz7DGYqyPBWTYNT1GYTVoeOUrTqpXfnTesoVYNG8x9Wxa4fb
2FZMn4n1LhBs8bqprhXnKo9hpV9tYnmnrW3bI3i5O/VUCdv6R/K39MkZzamQfVUl
EF46wiiu2AcH92cIAnshjNw2ZDHpU8+X4wyZ2TWSuT0BquFLUEtXlf7kWOWG2Rbz
F2fTFbVny26pWgAQhRpvzgx1dgQnx0BJ8MpPzz2SPaLFi4nZzE979fvu9ku1bFYz
JHMholgERsATkXWRtZexoTP2+FQXbPApq36oR2NhZj3JF29eEKzw0hccIppP1JmL
OMksP3NU1vk02/Jxho/9L4ob/CO+ax2+t986A864YM/crAiHb7u/MOtJM1rkHpaJ
swOKuMa0VpRil1XPWG4l5iBeAOKmPdhL7c9tUZkh3G2gbuxxWpEuiKmFUa3BC8p+
R3G1vbYoVPnsXd5hfoc7/sQMT0SQcbjzGfQ+Ei6wScngAczv1T6bFTkpLXVMAppT
guDy8iQNcQsEHfxjmEwHUVpjl4mq7WeRKQBVfBF/cyXFFARM7j4LMTZdCtTIwrou
8dak+k4K+ACdD4PWZW/P37DuVP0rIQzd/o8VcR9LLX5mojuFu8I1dtOfpJc54mMk
nnTrarYdNCrlaQZl9WLadeqBLMfbYL1oDvb/Fql3dtq8eImLBd4i1Phf0OyvUMo3
+Aa9znqK0QEQbK/0UihvnAsqb9jZ27b5hSkN9DFSEaZ5qzkN8tjPZUYYQcX579Q7
Q4cqqq5v1qRhuV2z3u4FxW+I8xYcUP/IvTVFWMM9Y6n4md4FnyfjHYyjLquGYqov
ec1wvbKDgLsvEFP6XFSybvPwlhBSWJ7JAWqAETjW+htZUG3r+mI91+AjBUzPphGZ
I7uQbSIhJrQSSyo2y2Uo5fepMwSwkpm3uVHuWXaUl6wLkl0jbixyAkcTFHIwTdGs
u7KnJk/mj8RnlwXgcfj3khZ3KTOILlpUuba1rXD+tqKeN9roORedamSBwy3Pnmb7
Bk5gvWa6zkH7QYFD50DDyDq5JrKA2PoxJIlmryADLFxxbyH5SNgldceQc6MZb9Gn
TeuAwt+wx5pQMa9Xo9ajTMJ+rBpjBpfEfr4Jv+gZJDNtpTqsvQsR61mfSCGg3hOm
Co8GrIT+uVzgRwh3TECXhBkWAaeUQQWf3DYFyAhbEzPM/1qmDlo+UnKnA/PYlgQX
ski+ggJTYi/Hngm2OORRcFvKCwnp7aO1y0X4Wk1yg2EnILFmBG5vSYz//m/ycQ3K
SEop9g+e/IEG7UxHGvDcKf2fpRT7SZH/qaBpNtYJ7kJD2RcyQ8bdg87J8QMxwuqO
5DpQThCrOVsG7c4v3Omw4A8H37vBuSZQaV/N/Lz7EUMMrJH6yJb70o6sK4WmYf59
ZLhmQLXc/D3o5JFB9pahggd5KIbFqGD5X8rpojDNjpu/VdApiujQx+p0RTAcwo8f
oXTTKn/cwEgM8aU8rKcTuKC/hQr5kYcjqPozfeb6yb7f8sTXrpH+PjtbRFLGCyWh
UaI4KBVTJ6fT2XmxQcSwUIjXJqnCe6zvSz1ob60Jfj5yzS56m7pZspoSaQ0i6301
px2+H/UwldjrHeKWQa97ZV7weLnNYMcy6UoTvyS1lNkHYmngSQ7/ioR8HBdCZvid
riVEAO1uT04VyJS59c25cM3ElrOsPv3s2F8qYAnBX5y3uBgYNM230Pbz+xuVkFxG
SRcvVcRofTSvsJfxTbqvYUEbtaKU591Qb5bsll3p5gI3a1MlhAH5ttV4kWVyujeZ
MNWP+KeX6EGpraakKhet5VWIM7Cdt7AP3lpVRBxUBcFZRVhsCNk7SOvCSyrLfNtt
I04lDGrZZD6NAjJm6zjFzFRDY+PX/aP0Rwwxp4ZpODqbJ1N90avPLAGdEAcrS6aB
zXMNxq5McmpOT6hDdmDdJSCKMtJ1K9dpuXKrSBvohrBR045kud576VMt93s6blZC
76KfQ4PcvWfBxcww2537tWUjuKYaqviKA4IOo0qolBa2cvWwtwU1crGJwB6IF2dA
e7W7W+fK0ASwkr2fIsd+P71e/hDqfxfGVo9PjwvARgQUMvlZCVJRAujxQl0av8aV
CoM2ZMuqV5l4yFQ97S/CoKqvKlrEV/haFmcyh3y8mckPvZfWxgGwmmAw1SB2kWm/
41qSNos/lam8TYw7PIoExVFe+gJDEnyzyXiXKuxYBJYoQEokKGcBc7nfW82RQHxF
0rOMwvlrqr10xNIdMJpwi6n+peWq7EZ6qGm0iGsZCtpnpPhjJKxdbyQg95r7JR+e
/XFHbwYbSgC6+q8n0dAOqNXpo0BcVN2eR7N+tlzJAFgFWU5c/OmoO0JvXCzsVXxJ
veeRm9ibQ7hkYb6S5BXo0b8fqTFWAT3MSEbhcBXmXXbHO+AJjPDFDdzWikeu6QmC
/mipMxbI0uHYPR4aZxTBBSAJVrn6TjwlpW09ypqlCXgG1LYkuV2B2+qZbP7lJLTO
6VYfVvsLPqvCpTcclexyrjF1smOIPnYA+EH2UFUa+egG3b5G3oM62daSF0rz/52N
baWjWik9bW3646a8w6+5AY0s6ixp1vQThSTObrsOOcE95qLaaEm6O9T7YEbotzBE
7iwUxkxQnEZRbbYQX9G2sj1fgpB72/7tQ0LXtdsDC766ZVXRJengQDRwIxKjTNY9
CATLhD5qB8Ht7LQzqvl5BsnopNvAe4PQvuiDVbN49ossKOFc6DGia60gV7EvaUpF
TDpY6hHzpx7kILOoQgF8RNUDmqPMA/i9kFHJzNT5E/vCxLQE3eDz9NrjeYJWrVhM
rgqGjzecOb+m5F7x9hT9G8hsdKbqL8cCiVJ6Wi8K2jyHDR/JxLybYbKas36EFJ3S
w6c/HbFusX/0hv1Cme+6Vy55HFhe1rWFmtqVmAYEaZ6LACcAjfOtLBYl7UEyhP72
Yg3pchVDCd+JFiZWEu+WZpcdBclF+njCsfCgXJKCCttkwEfcHDk2bT1eP/xtocZP
CBS+4hQh4UnefttxodN1KTA4w9IsaykyKw0JKU163GvT0ewg067oNsnpIBoRuuJH
AeB6YhX0smLrfn9RZoD7iIagAJVc6TSzIS87LeGtYpOUR0Bnr89BHGrj2qy6djHy
lZfIiAJd14S13mDAPjL0iVgxz0PPd9u9f741A9fBJjWKYdbappWSEV4kaG8PJHeB
Ux7ZSHedHNRmLmQBJEGZIc4Oglb9B0zPq/csdEFKEKMRGF6VTKPeYxc9pyzf8InO
P2WIVyJcWaEJCB5LGDITJCYUOencGSrpPzyvm8bZGd9mqqPx0Koh9VrrBp+UWbzJ
/dG9+mjOCqx+xX02AWZp/X8mh3bX7fIqcf6qoy+hWW8Yco1QckFUykLfAI48yL+p
qtdlDvfl8utvoVWiixOzg8siPavCozAE1fvVd+puN6ldiz6e89Rhv4QU98i/XQmC
lNC8dsBgqooBP/cUnzx+5YSXRTqtvFJGJfnZlaZeR1m8N0tPGUiyyANiLDdxBYdR
RB7qN1YR6+uV0/OqE0wvgRATMfjQxwqdTnyrRAiufv/++z3kt6HYeF52waB774fi
n+uIae93GLdAd7EnMpHQZwE3fxGV+HPbDqwUS5gB24ZbF87a0gOOsc2S/WI05UBb
ek7jfQS2TK6AxNiuu/XuOVWV2PbTbPr1P8YciG9pdhIqBbBmD9icxzxph/VUD+fS
amQ/2WEoqgTmiFgv8yIRL86Oq8eTJKFCh3NcF7Wp9BDQPd0Bbwt/+8r3HWEOJrGt
I2Hs75gPP/+P+df4Jqfa3nDsbjOA1chOf4V7CIWVkGiLkJ8V+0lHWskhEXp9e2A7
L+Desl98sqh524hMBeStAWUAyIy0LpzH0HUfI+SNASAYi9I/zZ3PwDekuNakzlBk
PWgxeyOQjL6gj0KQ9PaBA2DLVfp3Hh+Kb2lp1nGHJLqkLgKgtaxColE5JMCS0la/
Twz29IAwB6Q6TUjA3KkTxHDJH2cRnBUjNhdPg1GJDQLyOlAZ+CzdXKlO5Rlz4/Va
U2oYtGI3shWfGUL3Y9H8tq9QZr8uacb67KZGNnYuGm/DBmPr3F4qAhs4BdRFulNd
W7UgyR2TGJSS+UKCDywkVw2V1UP8fzfZpVzOhXjcFTuhlhdC7HyJvTybE4P4SNsZ
CsC5R0+qZh449YV8pORtDD42o7GwCTuixg2k9NulohwG3HAKUkK+yz8a1rMdfuLx
6NpMdxnmI2KRSad9vdNfLurWfa96yCzPX4Jsur1Qg52ryqIL4ns5H/CPw6b2MTNI
AOmkRZ4a+hYpo6h7/AQXXkQsXXAYLAWP4bBM6qJLh4pJ/2UaPPsEAAFVpRmZ8yA6
nNbbZ6ERvWIM5E7zUVMp0EBRQmFpZCBjzEPuSk1g8FkIyPz28Yk6jTbX4j3/EjYE
98wcy1UmK9Gmir5Oai8o+RcAJT2L6wrvUqG0LXdkiQCJwZZxILHN+Fryi/esMzKE
Jl7UtfqTY2+H6hsYKaDOUcrILR1C3ioepkEWbUhyvZF/0Cl+M2KWQvrBwosl+MVw
bJ7J1I4+57VNAjhKo+3QprnKa5aiYfGo8SvLxuwvbTvNVA5PAwWhRyAs9UbcBpcf
92YijjbX/Vjo28h4JaSA6Pdgxyduo2uezwIVqkzBig/f926hzSXWyni8bAcwwhcH
t5suu6+JPncIGSgsU0GzhxCWDzqpHGwBHuBrlKan5i40nVKbcc3aiFgk7kSnKorZ
GyMWSgaVk14b06WXQFn8tc7HLAhUyAV00lwXICRbyoUSVVbgWqZt1xxMsV3QV8A3
0EkYgntdn7hdq4/81QXZmka4JX7SjfcJKmfvO/b8IzLFsG03bS0d8owRo06Xr46l
zflekRThhi2n9N+vyWS75LswN4vMvzlX6/1FQ0PG6njZORDiMiwz4spCsXXJe7jr
28KNP5o+QyIaR7Zl9+Gwvpo0jDcCuK9PHf/UrNxwgObEfAgYhjdukOXgfSaZfzTI
TTrcEDv8SRaoVWmmuUTcokt0sqpJ6jZMWLIBfXuJn5CE5JcN0UeDx0SW7MXLmmkI
N++THlGY2adIlbbpNHpiCgW4Yy4k01vcRyYiwH01sBNQ6mU6pztwVD3qwbBdd0Mu
H48E88mjT//78p0gFDYSboV0fqIWf8v80Aar88bv6UntXcOYaxADM/ahSjp25sf4
ctWX4np7UNOKgWirM9V0CR3r5DGoRUM7n7dpo7pVjqFbsvxYTk7yVmB5Kh8YQ2q0
NkUA4TfAfn0wxyQC9jsX0D3MfcRBv9dtDub9n2qLxIE4qXXirqSD33qLJgMVHkfu
02Wr24WMie7u38g6dnujkxogyM4X77TSv5DGmxNnBidcyMCDCilSu18TH428FMAs
/QvfyJ2/JmqwZDptHMHL0zMZnrDv9Oi7NV2Rr2X6hV/KsSFobsZ1DCG3tdMURosB
+ayiZfrt38sJttJ+/H/sni/nMHy8rUzhtaOzzpQImIOJo/W4irhMmUmMTqxjQo5z
xFop4OulWOcScI1qoyACwPkB7Z9mRv2LP8yv26B48P3E+2/JSWenXvW5B7E0YfG6
VFl6gpyDoaNXj5hNt5VLbCSkZLBR4nS+bLqpqS6qxAgGGsPIz93b0WB3eTxzcnJq
ssEKsRbdNvaGUH86o3zafcr49knj17iVBc0P6rVszFyn8Dj7Kh+pL9FMHeCqj52b
Yy+jMVCjRXsNxlcqRgxRT8zYs0cnMENr3lDRrEG/t2mFszAqSfLnoGq4mca4IXmx
W/frPhJaxjAchyo9Jy1/WlktJl+BLczB4qcFHy8HxhU8Xyc7IUT6zMoyo9QnRo7Q
9JCyHI8SRKEcU/cyE7hrAcETLvpqVBRHCqJmK1sO9a3pNXxCjRc2Xe/f/nX8yX2m
4nEZIriEyISQUgd6qxWgJjznbNIFTFXqjMBt/Z22jWSkURSWB2blUfBTz/zwu91E
V+BMpqHXVWfECnXQhcyIzV2Si16d9LGMcx2IzQ/hAaush1MZqPpxbL/6mjtyRFqF
U8DsqQ/JKvC2P00hxhaWLbzIHH3TpMbMZavPlYxaTzJ53VUDvm4EHWNSnQPajvKp
unw4vOgzDjh9t6APBJC6j6Al9tW8qUfQMgj+FXIf8ZcYcerXzRzkuCFgP+awBlTX
BfnYck67p3stKS7EkE6NZn/Z04s0dSbsv1jJ0IkTNMi6DQzBRYhSIAhZS2xkVS1+
yJDjZbPxGyn1OOXCEC/OV3TP3Le7H5+Qb2t0+46piqDTWC3yHNotxOZ29iHn8XlU
r5WNVv/6QyC91GahmTCqUteN16WnDiIcmXKIVSJ2HqBGKQkuVOXExg7a2uBJ5kaX
uLBhz8FiJQEcsANFCJMDHdgrmICgSQYTkHs9KItOi2j+WeYjk5y+RwqSoaxLWqqy
BIkACIc9IIk6ogbtz0KhOsUxv2jX5zMvA95haDbz8yQB3l3Pi+N4AmX+1JkQdDg+
QtfuDMhHh72MlLTxzRSIuRnxOn9HnMQZjzBGS/yVP7xrebH/FH4J+7RaeFztbx58
w4ASY0H2TW36rQ/B28Jc7eouiiOiw930Klk/kKGr/2KCKqLhklY6QJKeRkveXXyS
qCzy7jkpi3YWCt5BoQ8HP8zk7Vf48Pa+Od9fB50FGZ7yiuc+IG+QZkjFBZHlDdJd
q1kYGDxdFnLQC95cuTknFi7QLe9gJ7jr0Pkp5T3Viiv2GZknTnEeRLqbalNPK+cj
lzbZKrmhu8oGK5gB8L8gJ+3Mpa0hgCp65jqBbojkMePgpBUtq1O4UaHVV3gWhZKe
IIhTCwCgYc7rdHs5355T3DdJp7ZwMKtHcZ7rUHRhRZ3batUDC/faiwpv8npdz8ov
SPpk2LDuGh1bK+V2mTGQakeiBSjm5HTxjjn7dfjQ/aWUCNdkWxrz0shpK5zlw2ws
QYQyWSS30xeT8bFugMTLDRxR55UaQ82pQgFkQaxyyypt29/pFhyWhBmMLyVTDCK+
2iAp7cP4rLy/jxf1ac6pkQ0HaiFy/kNv4cBThbLCKxvZIRftv9DXX8V595KGZJmc
j+FjZqD2Oyv6Mmv06/s9Z9fFPv57ayr2/bi93rzrxyymuCl4HjHlz/OumF7B/dsZ
zY1vkNrfvefjcpB/Jx5bWPYoFez9UXZjaLKxrAxfo12VsSTxr5omTMrytGv8iW8f
UQQsU+no8imNml7LdOna6UwtBoiFK6f4yottbm0/1nDjT3bte+1yZoDpVwyiHvaI
/O8+RarZKvLTei2UhETYjRVwZiv8QXY0qdoBXwsMtyLL2V9ZYaiYgtbIxqYhXqju
l0M3JKeueB7DYhOVOpaEJbugl6MphtojimJkgPE2euzEuTQ6ejoLwmM1OokEtKw6
75tkIIU7wa2ZOfL9/n25Cy532JkALTz5yRkoHvq8bfZh6lPHw/s1H8H9rKvJtU35
V0Qg1/X7rwRBR/jgnKcCsfdbaLIEbAqTcX2/O8f5ASfcXXstjSYKOPB2qAs1FnAV
8OtuYgcXBM6JLtE7S9ySzPKibbT6JHFsTFTEMPjkrsvEDWilr6IRu3QzQ0Npgp1F
4878bJ4OylYV9wGF0eWRsj4p6wNu+WKyIJbgHQnD602fwbDrz9GWnyL7BYEnLsJJ
m9jwkkaLV14ocYarbtFuWl0V/5berqLaOb23AEy4N0FGSqlhLgLoiUrbG99Oknnx
jnLFMsZSdDYrvjWBUjA0guessnZDMZP4qjbnadmbVsgUyEnfVsR9XTIi5pxPuazh
U9jf05WnIABGivN2MsW2Qf9lWqxxjURyHKspg5eBrbce50Otn7dd28/IQAg8j8uu
yZ9hnBDWcHdxyjF9Lt/VYmfbkjRHVDz4FbuUHCR694+2tlihRJSWkaV/1VBXws1g
QS7oC5RzABvPED59lsZUVGfB2qHiiN/0Aaj2yEjG076Dgf8nIPjHZtCKsCzFV7/v
7nPycDbxzd1nHxcxKe9sdAa5aorE4B9JINvtiirWWd5MblxFWi6TyWWCj84GWTVo
/eYH/CqOCSoAuPzkt9gCxWYnglIjO1NG0WxD0KtFKUnJ4mu1BASvJvWrFG/qVczc
ghrPW8NKS0FSzsHKiAz/5FDIRbxFyx4FhxAYzL6G46ta1K5bZap9N8qRi3G4AE0L
49LntuxCuob4AFnlKxITlFDOQ1iBkqH86/WPEuvIfft25B9Pi9kY/3of052cnmoU
ZZFoQXJFRRnJ+8/ZaL5ckAcWNdCzzLoO484c2UdLSXfpoPCMMIc/2KejQdCacQqZ
VYz6h958b08E2Z9q6vfgrqpB6weBMUADdcV17u5EMf6qhpIKZrDqdyGh5T+XGt4r
oPdB30up0cQKYN2nIWedje08ZubeVQONbPKnnNXszCGBiUEcZaLovUQUO3SiqBn5
6tbeuA/pePayrd7C/JxOTUP9+Z3VjAx7F2s2u0mC8hzB0OFH7WWNwRGJkoI5IntD
pRtn14TMcQYzfBnJM3ZMsU6bD9HWPNkZXVNVrrUhwGNOv99ULkyjiVfOHxlruQrx
ZljynRYHqKREFYEuJb0I3l88Gwf2Po5cwZ6DSEJyutPhxIQW5J6H0Czi8dRAplO+
xXmiTfG2gl8yVNnxjX+UA2a3Eftjautne/+kB+ZmiNQ/iCNycASVJgL+ThOGY/F/
WanWps//LEIfsiIRzBJYyfYFDGgDvPGf0O6sRvIukg+8hTQx9T0qwMVrPaGI4Ezs
NQYt8kBhZYMsTXjh6ekPUwWpuUHtuDrxho/SkDJYih8BWN3l+duAbHNaLKVOBmZU
X6X9jInWkZj3iD1EZDB1iyIV+eoRwrHheJCfOJGvLBdQi+hSJdO3feP9m/Bjv5Io
9qEcuDSTrl40o84bKg3SO++htW1LSYWPR5gT7QH2CLhomRPJOpuWV7BIPqKtf46b
RwxR6ovZ6PQ1GqnuxwXUDKD/EzMMxFm63cosE//raKkZQJHqvh3UenB9OV402+cc
OMy8TxvwNut3OtDXDgdmEApEbj9vKCbr6T1ADIebUbs0LAw1zTecylPB+rW4FQld
Gzms6LcE4WRgL4QFgQImHKgix1kYz+Gsi4T2Zvy+EgiZ1hvA8MSYnSQpbFuguSo6
QKp/bWS1rrZmAho2GxS47QrYy53sxTevWWNVAMCo0Gzh1unUENCNNGHjTNS6CQjQ
3gLvkLMOJySC1G5EfyvFtoDFV0dk6wdnG/VdckcPZoq6gsV5z3wxmya6yt08AFIZ
9Oy7fWSor0TSJRRse+xZDqRif5kf2xZcqyflTbjP2HjgSvGtFA5HpWYsCC80+bBl
8IZg5VgmUDdTz/nEwiP7YIqVFbofeTWxRIKLsEbLIoaUaTLZQYPM8Ypvt2Plj5Ug
8fj5YnUsyTXcIb/tgc/ZPV7ktiUwVhIJfLYlWzx8z/HpEgo3zvDGXdt45PvIVplY
l915BKjtOCRkcwOobVu8rR2vqYU7Iq0xe3Dv6JdUfLIW/pGahZwnSjOmdnyOfGZD
2FKL3l862kEkYljeKBM8IQ+VFqOWaJ6iuTvqsByaFhwyjXLxvLtO3B7BY5iMAyfM
UmTGQVoZ2EGLj/VYAgBa5rPMhBAUp+JLZfU+Mg2LqGR989N7tKe/HIRblBsRbZ+d
5T3BmFrjMe+B5YDolEOQixL1eQy04PROEWZg6wqzhIPtfzu1vxAdeKLPlHhH3PLt
TkbNRFjfmBb66xd8WP6Gf1mVsOTds2/xFPDRlgYkjYOyY+3jRpz82J10OlOMyj5Z
XJDI0oojdkaZu36/gLfWjzSgZZfxmxTSbO7UyJ79Ez72/8Hyd1oF3e8w5LNsCuow
vGL9sZrGTlAloWpWQ6b7XeOLgVs5gox2EAcN9osyjaXBTxBVTuj9Fewv5BSy1xpn
2lz/Jruinp4P6fRDgyd04gq2ADkTQ5eW0hc8zphsOpEbgRgtnHO4uFWAfCSlIH8M
23DOWH5wYDKqxSTJ7wg/e2WK3yrDyIdoOpFIvd5zKyBDjDdfDojRHt7suQA+NfKE
U8vBcdcULwju6wVgk9iDDn/WyOAxDNbn71XtFbe7htraHEJLmlKVNQ8Jg0HeuAPs
zBjVdPPL39PRWTKAxPJ3TfnqlGu1ZU7mLH8dE6WtAhl9vd2ipVePBopQ1eETyIdR
TFJkxs2KO7BwRueOZ9tuOHkIBcGe8C1kETsf2XkzTZ5+q+zkKqBPmIbjiFKYyD3P
Oqe+/uKVgQlUNLVIldFslu1PE6UeVywjNyO1MUyFv0jWqRMqPj1b+4L2dJvb8eFr
N8fjv3Mc4e5AAxc1ySZ0ggUxTiTJAwciTTUj5bQB/no3CM2vuFW3wY/3P4afPa6C
dG840rFCQAZA94cDB2oOr3HipyJYyqnaXpO/6X4Rxha6FMXDmv8jMh4UMRnQlU6j
pQW2hB2jYQJvLEzJNmpMo9wyCnv5xac6HcLmB3bPOw800UPv3LvsBxUmL5PFyDMC
u2TN/o74yEKTGAVouEpaoum7m9fbJiSa8o4/uvhyFJCGJFXlSjry/dMgqoyabq7F
0bQtILyH5o0lYVeIDlXLnbwc/iUk1WeuPL5PaNQE1jRsrI6ObhxId2/T/NkQSvQY
JNfsaDAf1dd5ypDKOMUw3DlWsDsIAhtWVX0cYVZF0P6mrdSovZrh/lnLnoWX7s27
QZK6LAwqKQIU0lcx2VnKFtIFADewmh8Kzq/Eea09UTgDeQCB+GceB15n32XyzdYV
6SWVZLjKj2DZGmwZVpbVLgsKuQkMUf1bY0xMp4HmbE2O72XJ2z/qGsAHNNXzJXYc
ZzirYtr/Ju/iGRhMgpv2vh4uZZIFhBUBifuC4VcLmwrh0k5bPWpZ9NCbEEGDAwSy
rXJvsdPOK8QCrf5CDqoOhg49usYvazcMKLzf/uKU08xczyw8U8QXoxaLDscRWENw
YAT1RwGBAt7vQmux8SuwJRDm8S4E2qLnh/jz9EI0WKHLVA5sCFV/9ZBBPHzix1x2
ta4aoBFEqFjkBg7FH/p06jVX6hen0GAho3Obz6UHxs08WVg3iJ2gPebWzZg+eqtH
5/zP/ILKE8fqx/2KRtHz66CdJUrOTr6MEvKCw8ISFfo5tODmOwnkXzmc/lkvCh/J
UEnMdt/X5ZtKUNxlFngmPfFTotlJ4zRxuk2eXXJe+qkelIOimMqZisCAavGEMTVN
ddyjx6EmQGBdlgfOALZ6OuqhCq9KkB/kRYD4Xgwt4mV7KMAQ4P0XFEh9rs4ei+Qi
kQbp+3xN8Lq3unqowDwYKIwYjRga79gDYPCfsVx+8kPA2SV9nHUNYUJ8CV6bum66
7YOCbLZ2GVsrvWi2kPeHAVA2+xyJzkCC9xzTlKdjKFGG5u4JDgHJgX64GIUwdf1E
D4WI139+SXmPlEeJhPsGDhl0Uu40mivL+wmleiCV//fkr0mz01bY56zVCojcE2LI
a2R9NW+TriNOSGkmq3W+N9pkkwmN9D4RBGaNRVVSV21afFR0hkAkddKxEMo7ZVkI
yefEBKi7bAxNFxBjzvNWJixm89QtsLCiikwcutoZg6GZ63esRS6myZwMufROlALR
GhrnEnpSz12naxWlCcPG3tlxfIe7AYP+uipW3OGPIoRmtba44paM3MbC/e4sBgJ6
MGRvKFY2ZHo4jZ7z8abpxNDIZZe+PC1wdH5nhRQ7x8X1s8RgAcZaEV0oPsl985rY
hhkkXyaVyTlEmhMtd5Y475ZPNwt3GJNTby22Svk1DfcfFi1XLSX8h2AoRc4cZCQ/
G37hvfi0/s88bCvcH07gGqIiuUHW+e9UzM4EZTcaw8HQkJSR6lvSfUbmgplcyVUw
408NbxHzI4OQ/3PZ/P9nz2LeWP+XJgUN8w0kZF4n5YmJ1b1BEjuzAQCmfL1Zw1tm
0fkJKRUOb2+aAGQwM9Q/XNcU/2YHPm4LGsUbX9x3E8ZzhiOPZ892f8JlyLr0gS8p
wXePOM3If7dUz5KQ5gV53kmwMY1XbQRT9Z/GJ0i01PQxfXKEHVT4hzttNVV/QlH7
sPN5Tbc2dOgV/S/jSwcFmtpW9G2b7O9vMvjVlsbPorpRBFGMaaKfMsgwKGB6+6kh
2mLn5xCJVmzv8WmDt14nQ3Sfk8uSYre82+r46f6GaioIWJwOzdeGqJgreGT98gS5
ygJoHTUjXZ5dCSGFEgkfHSBJjGLGaSJFmKpDXni0EmpdF4FgYXe9Fydd2C+/xunz
TC6Lw+V1bBYqXyiN0Dg/jIqRO2s0BuQWQJFuMgo4z89FR1iBp7mMWi49X6D04iiR
Nl0bwCg4duguh/2J13a60E5w4FVb5epNk9dXv82ZLk1ZXrqPgs4qaTL3b0aJ1LdJ
qBPqT7Wiz6xS5e4I/KzuRtEE4IG0L0pi79KnzoMk/yvpMs2HF7LgI5wXIVm9RBr3
8pXglec5P62QbhE6hkQAOWGDE93B/XadU5RZaOFLgk2f6eCVcFa5JDaJaedr2t4E
8xl0w+PZ3p5TuA1of5f58GmW48RdX9/Kg8H3TeC/sKfaI3BFqTXXJZHwmboFzez8
MqOv3JnoZNJPzIbgWRvDA+7kp9KGas3zVfL4/3sL4ExlV3H0BMic0aTE1a/ZvFjR
QvRemm9FWG4DgBrU2dmR16qaixkMusjvJ0cGpjcUMwAFbKKf18NdZLhtFv1lajnA
0hgYtkbt/Dw7pPO4nAQaRCLrYMaMWogT6uuyoyJKc9Htjv44bZLIbHgBDSHUPKH9
mU15meU1XlqQ/KcuL56g2uvNKhhhb7QMgfSa4+kh88IdMS+VSjvPTAVbJ66IP2L5
JXNYA66+QcTy7lHI+nLf5tms0fKE+Thn+b6Wq1/n3dN4dQHsIGUgBLl6OPgCLKsW
fj2YvZF5yQ9gu3yB/RgnP9fj0Q6Fvn70cS4lCVAVWzSh1LixQ6Ehy38wr0BCrvc1
WNzy0kSLh89T5gKzY1bGO/gDtD/HPdav/DEkBgHsfX2sGkOxpaq6wfvolwtb++M2
tg49gHCWdgf6/ezr4CCIy3/9hwh2mjbPZm+VgNxpBoEw8fagm2MNqaXIiSILymiY
CNqiTPYBMs4Rn/rLFg1QhqzwtTB43E32aBVWFhMnMkijQSVpixR+k+6G2VvM6cPo
lEKifp3zeXBs00qlNo/++viOb4J6HHaspnhyyeIB+m7K9CfohJKgfTVxsP9jtv1k
rO4Atd5XafRKlu8D7eOsr19QyA9mrMdsueBtt97Kq6iAM+jByc9MT1erG82ZOaAy
gIneYeAjgqkHjCkTBWIZR2FW0p76+oimcTNvmRToLB40+U79Sbp7d/GXGDtFYRMc
vBJhctzeA5viPVNYwBSDPfzB/SJSRYcawvhK3UA+eC/651ePWWp6KcweUSYuT+c6
yz8/MuVHgYhW59/KSFx+aiiz9kDFW1B/yo8oWm3uvPR2VHPZPPRMC/sLM65KKmE1
FHmchFjHFcFOR05GOA/u0BsyextwnHzAu81JpStmkyMe9dN0Gk9jxj8+HUpawufu
D3+o+wAlDW9k6H4iUoE9jUGE3N0o/KsgoVkhchuX9WA6jiXvR0WSSTkfUGS9EmK0
ofSABfO6erJ2aJtWv6CwQJq0Ic+kbiJhC+k3NaEa+u7dD346OWWtgj+1bVVBWp/Q
NEJmExT3N5xk57c9VE5VklbMTQAYFYiyeA0xoQQq/2aN9btqR4OLeobVL/epBV4V
T6zJ929eOv/Xy2Ta7i91mJ1T68CGM58PNc9PgA23dXaqBxsy0PaQOLr4QlNTPqk/
PQ9xoRS6sBf8Q01wLQP1zzWRPXoR5SSYLLkI4jxTvppfenzVRX1PlwSzjoqrmrfX
rM5UR0No6EHKfFjuwQp08z0IwkBQ9qHWnHUwEOr6knMMve4aPuWSgT4j4BetLU17
TRizxN6KUCmyMKZ5ksygt/hUkuBt5/wkFsflljcquIgiu8NCYk2gLs6a/Y6WE1lr
eiT/VavEkIAHdKONeq2dMQ0nAD2BFjaAiE5/dOvZQSIK6rpzY2Fjwzz++lds6jFd
M5g0Aa0XefvyLz5q6SapUkh9iI1H6nZrGfvb72KaP1oBlcwD59xjTT27g/O+b6oU
Lx8gpe2c+IUMk16BlkZZoIjNVf2ixH9mgrAA4iPGq19G6npNzCmss/6ukW3WQLLd
kJdrL3M/qTpfG25c2dNgKZ2ANWLDRSIIpUj1f9emKUaWBZcbKb5Pyh1uGvorl5/T
ooEXv6t7Djg0f3/m4ukWO5wE7sR1cck8mv2PednJXbCPUPdr49x4a7A1F8jLnxRo
C6/HZgasFj7JzeW19716BTp9Q7YTKaF7jtIHyDiirA4Ty7N9W2pmcKDtLGtCgqdM
erW898gHQsIzyTlboAjPSOKudkeweW+5buUs+qi63K9iwvMOt1xan8Ab6Hc1PUBp
pE66oplb/g6bd7nLSszI0oTHtZKZj0EjInnIRylex7gZpeYIiU0lKR8w48iaU0Qb
WjIlq2EzP+zTzkZoaEanhLkplsFKWxGSMTud9TGQ+eLOnjL/udzy8P64KZiRlBSq
WCOg5p5tDkpIl2qDFnclEey8AAFbhE2dWdkVycF5Pw1DeptW9t2VpxlJZ8mAoXsd
bLd7TNZzTizRK2M3iGhA45wLgrQHFZVZJHoizUMXJYrWixEhuZ0iXPyU4GlTYD83
GTzlY3/UfZ+jMJTgjEIqKbzu8WyCp4vAKQx5VonXFNL7p8kO/tXQKsgZvu+y36mc
OlvJrAWJyJuFvoWMiQUTUO1b+kWSQl0NUfiohgEeQaVUh19/Vco9Ff67zAzOoRf8
ksvjJBC6j4IINijwZhcCLvfh/ZkXCjDXcPXZEnkzRyPz4kgartb8FMwxytu5hueV
xhdF4NuJj1X3QLOyKXwnUIXrdCK2PmYj2y5IReTXqeU6BaIQaCIUF8xV6//iQ7DP
S4tdKBYaluMNEZqpsY8sqhnTVMJ0xdG0RpZwXjEITyAJmp6mOii/niYVUTIAgVlc
IZqiP28TBK9CVUyoBAEnYZEzAEyFLv/iFVdTs5Kk5/Yc1jRyNugZPXzUX9cCRhwN
JxkpNCNlKz4Wi1pbAx8LFvK39jgzDijW6lW41hna3L/uaLuLHzl/U2icKjrtW3i9
jAqz0jyPGJmVjU55M4uqg2IaPD3JH6yB1vi/KNEmu6PIghdDc+0TUXo4RtZHmgho
J05j1MT5GDZobZ7GpfpXfsRFTk4P8isvSGj579QtPGCq8ewQe+2K93FpHofVgQ30
ABjIdFaiBI83FFUpnjYZ1RzrkBzEqRDFZy5XMMt8G5X9+a5g+2mcE7VDcOKa78Pj
d7x1WGul+uVlNTJm3M/rfzFbj0bQIOitizroemxaIfbfFIdEJMlnwJ5/r3xnZfyp
aHHlZhMTF/cjlh6c8C8+GmE8c4PIXiY7qUZvpfJxAOyVZu/EWAVktLlctJwE0bTW
2xkH2iC3sJYr0HCXpM0g/vhAc+3H7F1PhRk1GsBYsgchf3VtUj+85NefAOwOh9nS
i1UevyTmX4RjPVuItcnaOEjPae7sQUljulBVSXnk7y/O8u2fazStOE0WGUAixwOq
8HN9W70bGs6rnkswFbDJEUXpluqfkM+lb9MKGzJBVccuLDnx7JEnq4KL0Kx8TWhb
IYQwGqOyCkyk54h7dlJ/vN5jqqzNfdijl5hYw65FdDC+2SSW9afQYNcVhXmoWGQ4
PdTnEpnoij5I6Wt3N1nvyOM4ioYbbBt/8InD2PechHm8I3axzIxB7MLdVScMkOj/
+qbPYvceCw1Q3ZLBKd4HxGlZWBgaalvgQjm/uFNm7VF/TuiqIavcbYstNKtszDyo
6lNzrYNXU09WZF7VPVB5SwexMZmtlDnY6LWY6NTw5ycd3q0RLw53floozIpG+PGi
50oL3CcqIuzNIDV73fu6/e/G7zurf52jO+lK7qrbHIRmvoFs9QJklCZQllT/Ou8F
9c0cfR7qb5kVN7vRIRx31A+plGTvuNoHEOtg3o5qm7gBqrbCj9lA2G+JulKGhzhO
jjv5UpILEc68F3+b47NS3c/lCQ4/I66CjrCGDuJB6b2RhZIlHkwoCorPwEGOsy7H
FWUYTy493QZThQ131hMj2rATRX7LAwPVcZYDjWBseuKozc/qSs4JOajbh2Xm/kBO
7zj1BMrF416KDal92P2bQ+XOParahlXdM4uAfqxtvQGmpUPkx+LZBIfb9t5I+3dQ
bihyjnI17BXCy5PxSDGtILcwxYZdcOBV4fbN0eK278Dp0VQpsVsjDGUqMGgI8ahm
o2GDATzNLmqSiAnFV/8H80UhSRXRU8AKHBUvirbh9H1o8AS3+RsyK/rCQRT6dNKC
jOeTed5GPWvndiAHmv4uTLXU/hLKuDfUjJVSozXAJZssKi3WJUA8N4YFcTubXnnL
yZZEKkGTGBH9TF6pYaRikal+lcTN7GCh3OKPkcuFGE8udAAQjXLmOAqD9uDBD+gi
8R0EnFTZgnDhrk1ZSRU8xavdkiMySjobM6IJn6K6/kgnqrtJ/xhl0+lwg8WNhCOa
jowSj0ai6cAqJ+DTZupPk5pxL5w3Cxqd5uyNxkjgp+gy47sXMpAEXPNxhS12c+vz
bfQYijNnE28Q7ScBzU+k2ZLiBgbJdteV8pTru95jzdXYOSwzjmcqJEHkHa37LAM2
xJD9rOe2jWEm4t83I7YUSDHkJP2cc6p6azzaKHUk4Aa+Ql99yBIbGqN+8jL5qxPD
CF0G4sx8xfKMjABahP5kYFtNE5f0lvdKjaCdciK9lilWHTB1ClN+bAkwBU1/C9Y7
cS2HAyiKn0Z8xg54Zgvo8YJ1M+ON6TMCSWuBbEHfYn/7CfmNG1YGnMGOLO6yIESR
YQ+r9Jl9s3j9JpcFodCCzEbNwrUwzIEXex3Bh4sssbpuFC4AlCK9MihOUKy5o6q6
Kx4sSlBSeY/IdNvmXrq7ztl8cib60H+uhYJtX/sMRZoVMsVZ6+mKMQ6UdaYw1wLX
TYpLtzslOUTH1EI7PM+pAc+YlnqYei1wsakMOtG7yd52IHYu0zlowi1prKBPqE7E
w3KFM1V30lNY+5Z30qfNHcG+gQQhgL86bmVLE+IQs2hr+lqhPyFLLG04lyWMinF2
MAFqOmQjZ5MmcePitLDTnd/8ap21cUewUtKtBcpdK7kklG2o5RarNRp0+YIsbwkW
9+LxdPureR7q+b94AxmxAJkEH2OklYqdySf7hH71QHmkQS9LFf8g0yHCDd1Of3mV
URpFJ0zYQfNitaiER/d/XDX9rWGqO+TkhQyPoCI2tanGPU3Qzg0EshpQdTFKfgjg
dW3q8I1LOZ6LhcC6+grQoFKTFX971A0q9p5n6aFO277geegCVhXuwCcoXliN+35B
USV4Kgh+fFVjTuMu4QBWqQA/zrHBFIFfxMybUhyRekN/ZRTMkL1T1y5q6Mr8+0X9
oQRyBuGeexdQPAQVvYU4ATApw20yNKA0el9htC+3/XYgGrYQyV69Em8rJyDa4l9j
yyADu0ZVnOtl/UzXlQQwU4s5FemEyxg/W/GsyDz8PdYdHpn7TGh2XWHwVLL1aNYO
J+vA0bxtZEoI0Nh8+dd2CEMGh661DvaGj8IGqHmDunvT4sUYq7z+xNafvk29unf0
hwT+uwcpkMy5MSbROHaJF0uzIMvrCAyBzM5x1GjEBNXje4hoMB3qE8sPS0bU0qjU
6ico4Tbl7wgKiPCXVEcw+bi7C89kgr6DarAHhDUu2c3PsusJkgNyVAEYNt5kdNST
HLTSINIWtYJUfeJ//kg++/NCueF4Udick9LQPal/TmyPPg2ztcLOiN0iozCqFb19
sMUi+bHP6wqx/bLWRNBkKmr2qhQ8YnL+MhLSxrSYYxm7IUA4QctlCtUXHiaNAYbZ
FWfg7NKiXiT5AQe5C4wFS3yU+Ma5EGFZUHqMkS3UXKq7eDWE5ZdQdcEixwOLY8nC
fXZBht+wYHnkQfL3wyXC1SgV4Frx7zUo2g3vfFoBYFRtYzWI7tIIK4y/fcgGlMRR
qwo9w+T38xRgBpmQrCscx37LVVQL7lk7PPWrHappLyIexrhQX5BDGY8coxZFgyES
rR/v9x9OF9uqnBx3GbWkbDzMIs46BToKRxaI+xOaYwj6tfGACFZWn3BqWHNsM89c
ZlF5XodQST+5uCJjg0CdwhTZk2McU+EMMu2dOXOCxfRKBTma4AFnuFnivZvSKsN3
Oy0Ty3rYHSkYUmFgMzpBb/TacovrXBSv4XW5UELxck5b+aW9M+o/I11O/9esgL2r
SEo+CMWF3IYAERlsVgFBj3wK1bAotG9+MSSew6Q59zqMBfarZNFgXksB6XBHvOxy
6Hga4bv2pFLNOUX6+uH048oWl9vffidC274gW8oqVYcdnemKpPPioIEGWUylBYBv
+DU4giwCPBihdHsyiBBUcrTL5KFyGl9BrefRqzsnSiPsbBxmZMcoFn5EXZM+0P2G
S/zhL1DMqrj7jDW0OP06YmoGax3xelvoOynAR+xFWCzhiSoUhmfFhHoWf6nzTcbR
iP7kmBU9v1yejFgMASFeYNLDqAl1PwVjanYflOh8sAbv3UeFEqZzZ+B+OyQopZwQ
nXa7nK8aFVQijvO+P1CJGiF2di0lLJ0X5IxQq3cXxSSzohx7vrsNI0KcRY72rkA4
WPzZ77yC9os9EuKHNEqEHq+hbg3gGku21KUCZLLcJjnBZ1iBIYZnd/VtKc4Vx0S6
eB0wqpZa7dpDCB/JZ64xd7m8lhPMxklFicpeRiMgL4eSlxeXeH7rjL8ENRDzQloP
ccPiKPmCjCDzq6Effp2fIrsPsbauQxpgIfMguFdAqaFCisPvBtYeaMwnGSQTAbji
mTbp9V2CMS9M8ZSPwtIe03OhGs6g+mvibrpl9UIaWjxA/ZjwHjJV7EDTee2G4KM8
h6NsfR/IR83Zb0lc+o/Q4wWCH1V/pdjDCd51KyG1yBCxbQzlTmy3hf1iITBL6hTH
wEzVlxK3R5RBfV+Rsh8AdBZz/BztsV42KqMLrfirFbWIdEye18YPhm8C/97D9e4j
k92zjWrAhaLTQIdtWOIB+7ii13dBSv7qt3Hd2Ka219QBtufXXKGqvDe2srTng6fC
f2S34bzDnL7l7ipv7gv3dAwc8KMJvpvTmUl8eXqMZR1b7TmGpIUrmKgLo/pwp8zj
LfDELwnpioVZFKatSb8DaDvgVvP82D5RzF5roG4zSzn3cnUrbdPJ0w/i/M5ryt2j
tTT/qN5GhdMRINQLd6a942mZwSWB19xVIUjLq3xoCrXS6EN1WryQW6jXmkNFu1Db
9aVPLHugShfqJOz4Ev5r4+Ga5h8Y2Czmy4URylEv0UkiKvzYSt3R84ceWU2Z2aSm
Wl/VAW1mXtDJ7FUY1l5vlnVFuoHlE3D3kn1UE5aoUWZhBU1aD7Y2ylMq+CnTvS85
GDQ/pvxOkMo7ukigPq1nL1YbKcUS/3yLsDTTPumZQzv6FOP8WIvaFzPqHRctZHvj
ihMeKckMUWJc7TCqAC04A266796oFLfR8B0N3AeahavWcZ9fLxYtC3gYSU2xdj1Z
DLqJUtdUaGs7Vz9wa3TuJ1VbYWKXND3lV2jSwUhUzMXEGJ0zHfui6FlqP650tzlj
WdqwrsIcE7JYatwW6v9vj1TwTKLnCt3wqCFvO4PO7eC66Mt33DoNRwihH5hTYxSR
MjRC5Oxg2vGvrpF+YcDpD0isLYF4bjawo4eBnUxKy70nhurNigwhWUt33kTZ+l1p
HWBshGHnTHMAuyvG3p2WrIKRYuoDIfduMNmIt8/eGIG2ZfyOIACpvATeUKJMDEZ1
7TFK55EH8rOP2AksYWOfeyk/+ksaK9h6uLTAHZEeSRKxJN1IH2+F4i95lqUvLZdu
QdXARIBzZS2uJg4l8vSTwQMTK7Yy+hcHtm+nVjHJy6C6ooMN/tqvPsQ8Ny4L7L6H
A3wnebo+Z7uy+NhNx1RF2X/fkqtEfaMcuJmPgyQcrad1CFDiHmTJ3TTqWpkMc90n
p9T8vzjqXhzvKKPfpRz/fdlUIpcstPl63SsjCeCqHjjnOoeNJiUJ6nDLALXnuz27
8WGG5ZKhQbioo6W2fvCfDjDtkXanPpw2+7U8hJvAgUI+lX/Xl6v1YLTNU+Z/Mj9P
TsOjmavgwblejh5i9619rmQ37l9x+DZNF8wTBmtNhaO68/htcjPkhspZLtvscIg7
cjQER8GYPwJdJbJFZoxXByo//DjeB9O8DNFEH7IJSR4rAaBf/0rnFmjTBmjIEnq+
awUS+wvjqYbMvdcx0ppkIue2/w8hMIKT/FlVkI+M87qyScyZyDZt8J8hj8xpVMR0
f4BiO+GPJa37FzjtJbOPWildix8gJhCakl9vQ6UfPc/jC9lOPHLCmnvvOrhVKMvl
SCQOAawIJuF9yazjogxSZQgQA/wX22hbM7iHR7m/f1J5WDo+2zi8Os9N0Jv70ejO
Yj93d6zG6jfQAU/VTp4cE4lRIaHEoOYSiY/jqAoMa6s0bHj9yQZY5JXQ93dfaFxv
D9zHvPPl/7TPJjuUSf0OK/bK48SK+ICukzjdrUDOHmueagjvTBHkGYfuV1oXPF8g
3jp/4iB4zV8hVIfZxE3Faq+9iyZcXkIexu/IQyCBLnIuFYXBlmR0nAauFmO2ptK7
P3H2612WoBhQGDDMlZoG+CBZuH8853IZx51wClccQkdrKgKFA7YXuRerFaTOOu02
DtG7+qsz7xEydsEp6TPiKrNZE/ccW7Z6xsZy/WTrHANuCnnfDGt0iB8vH9Acw64t
aRXlqLJhiWgcy7lFfhwch1X8D8N+siykrPZPUkwHgV+tdVdHbDxp1MTojgQYTbtU
d/Sphzk99KDY1erePEQzsiL77+i1EojWgTtUDCaVMJA6xjh5ZdiBsH4l/sIS1z4G
Q2mSI9bj2hIvxjTSts9MPhSF4+tqZDEf9QzfcjuVDyVpGmbVSGNRliC0EjBQG8op
cni+YaKkn+kg/XjPl/YS91CApMEKP73/V/u6ehHoRsBuo445NSa9ez8lCY9b3IKu
SGJ0Ny5mWD4lIAMduOCnomtxduRbWybhRC6GMeJ/obyq+7sInnxie1unGzZbLjwK
mliap3VgmEt1tuOypAYmpzRZcEaMEHkpo8JxTGrXSD/MtkiefHHB1f0I88b9JFH3
ACSwhsvZoUmfGJ3u07l3kvymzM6/ZBKszhi3olLekg1TTLZQ1jt9uKn2bjEfxzfI
l6lLLoYZHfL41XQUhrYfsgORDH2vUSj1YuJopYvOFd1YgmrPQAausP4CNN9dMDxI
yJvEi/R5njfqywUoT5x0f4W3rwkt/vab5ZKytXv0QPbJRt0JF4O06MHDJAgZaeht
4OX0iyHjXQUx23lKPVVcXrEsJDtKUvYfVY2UjcwcEJ1njFkNbQsRlqjDSHmdmdG6
A9rI+gaEWBLIXnPD18FjPUGCqegXnxILc4s41VTEZSZUgJSsmhGamePgV7wS0eyr
VIlCHhTJVXuOpJUn5nYbaSzZZVowmNuxx6hHFshK180Uk0jfYXeYiR//U7o7ViPd
d7mInUAzV5dKdff9J+6MuoN/B8iolak+eKjZaDaXcsQR2Qf1qKDt/fj16sKWNfVU
1uWhoCxe93S1gZbdmqQDOq32FP8Nxy2j5PONvuLzQByNvb5UbyKVZq5fCIUl/UAh
VPZKyjKb48jkaLZc2R5r3VcoQkD7vO0JUvZQFgBpzyEcKzp8A+gnnwNOaA6ob4nU
A4lE8wK3+FREtuIWXSBArIA02SkmjFZeKlIQmyi3UkxIh8luWWLthkWaZWOGCYCp
3LnqUVoU/EW2sZgu7WbNT1+R1RXo6yJzkF2bWrw03yNRd3h1LcmZfMh3ISGXxo8F
19z2jNdQzIE/+5XOf5Ce4QEk7fgXdLVavr2E/GLF/0b5hkTXCbTfY5Fk6MojT5VG
tiHHmn2O106Q/zdbCioEDKFIZ6NkeRvsYUDV3TVua8SwvYdYzPha2UiX8WL8T65c
6J7RU+WfJrpat/KQZ2PYTsbqZb9hjrGK+6OvHkltbeLY3iPRokqZbaQJP5ayu0Np
FFMjpr2N4hhkPmBVFDxgmmhXOYgOBvYuS6TNjski7lNR6pBKnao932RRIDTXJY+Y
PLxx+Y4ihUOpK7LPygj9yoFWvl9MrkN5hG/aulPML8PSpZG2VVAvAnF7kJrhPfk/
x88CuHpTotJEXazY5kAkIWZJnSmH08fLc9lyME3yt+sIR+Tzd2Vu+6kydu72jN8x
10L4FKnhvD06xXG5zSrVqtdwjuGSxJPg20GNzdbmw9GlwxenKh3VzmlLPIKEPWsj
o1eB3AE/I1KiobNW8+hgeJPpZB3LTUEfRn9QBrCWN2lreGTOtCcJpidvrpPdDoa9
rj30YWhRHiK7JNBnslglcpdXD+nVGj+K/hdPnItHYD+u2AhZhHPOVWwru1hhr8z8
UWsdIU9Fg4YfPdOdKz6Vc0/BYJ6QVFPU4v8L/R/v9h0sm4rJK65DknhcUTwranIx
YZNJpQLEk27QvaQIxCmheG6aomPQpG2EFe+w/wutr6ebgPAvF5TCVrhPctJL6kGM
N14ghL8BrBXvcWgbY6qOir0P8dXQ5bzVSd8SXIiTcP/ZyQiYVTbs9HxjYi/oT3/a
30T3oF4yl9ljZSt7+cNb0+6cgBHWJEs0V6aONe0AJkWHo1vycjBGpy7A3g8LPpX7
FD6qpViS0VnwP2EZyjcyPmGVeWdbatt3NT5wWCdBLaw5bpozHpMTOtpcGi6IFOQp
IBnmGZqu+nxVYTIdxNN/UbdB6vjnPvocTJq9PsoGSEFRGARYMFUSWbt2HZ+NUeLK
LPt48WndtZM5BTEpttvyhIW2Gt8ecohi99HJWj/22VXQNkjmtUUQiK9IMhF3UlKg
/TMyDNXbaqqwxjjX7XfaVRPRScsHOZ7ieELqT0v1H0GLwn+3bTJyLdQW7W6Sso/V
SxNlO6DCdT7bbcuYaUmCOwy1RcdaORRw6vSGqQD8ysQUXao2qcucV+hJsbzbFBpf
m3t1sK3pE2gRFhS5UWDanciO4liJQovDBUnsEzhL59ZfqzssFGypAYVOsWGKm1vF
7GXv3hQLKAdNiHMxhsSZ+c9yf75wzr74SB/KLcO1jiTrHY0PqrgtTft2yA2JtuWx
9wibbPFOXiRbgF6sDnypX2mdwiqgmq9isnCNzzCnKzzxtFGyNecFkh41cvXTxjSb
wpu+ht2BA4OWIi3irmW6+PYfo6sj9pzSgNgz74sg7pYk9sz1eJFXG1jWlhzXNkyQ
5GprU5xH7+SqmXlksYaAirqif6QeBcSjw5iVFHCy6wywP0MP/ebCT5rT5oby4Mmz
Vr0L/doDWn0Y82goQAVRXxxLvnNL53R9xfHwsZehUskLiNJchLZG7T3DyuYayTJX
NxEw+JEChMCJwBb9mDuGBPD75Ay06sxbHzz3ozOLQvCRCNtIqH+vpkmLcxCFvRxw
P7BQ75yfckTvzSGg8ZBWT6cJbIfINu2EwV7dwRt1zJDPc1/Z4C/xrRMGNPymoe/n
KRBU4Rct+4P6sEj+1AbqL74qd8c+qZzV7TUvs+ycG8XYZpKIuVECXz8ajUEbsGjY
HpkRQ6Nd1qvAdjEvVd5ShG6E4Cmo2UfQq4DpjkOkOzaZz33AIk361J8vjN85aOB5
g0lZveqagirNw+fnqd5q+WFzj0L1kcsYmdYnm3OfUOehQ3hk4MS0tdY5JjmgTwDf
QKsjL/tysBfYBF9xYRSSb11vsI9GII8SIOhQfmgxVD9EWZjJU2nMUJbkNprkH0cM
+KgrWUMllsQ4BxhUd5OW/QB+E4M4i/ddpKlQaXNTi1mXF4kKaQkTY5YmbO4V/scr
BXdc8afNC5SrC94c6VMVX5rGQuC/Fs602rNEdKOVb+bdiFdYvfp5UtD8vDXxIa5N
bezC9bWbp0I7sAuJAP1PE+YTqts97jwLmTYRiEVg3iWUKZ12I5jgllQ85uo4QHu4
H4q3ZwKSmKX/FYupTkYUEEUqmYKcuypxeYqeZMKWo3ETs6ZVvk1TlLJ09id8ind+
P6bdcWYLUgmlQZ+sQI00PA6XMNzyjrUduaThSGweFmu81KnQakagwPio7sNA6KeQ
ekJk/mjfPwJzpqL6Ruz6cwW7N/tSmQ8K+Kmt2cbJ/Kidg1NpqYvT6evfMvVxOP6J
o8odwV27ZteundhZ1xkbGUKptE6UzrnW5/wxzaG6Y45tVUNFDLGkvdq4V4cOH3cR
uocZagy/+H9NnJlKcdDEvp4z4UbvbYEMpO3vlKAjmuGlaNXo7QWcCLiPeIpneYJc
GJgSpqSsnHYeXRlsjp7ViGgYTIxN6P7FzOew9OIMX1bF1LugfYCEiTH7KLSGAB/A
l6kp5mGAeAqaJ7jo1e0vqoEGYy7Ls3wztCa0Wqkkgo6qVWEBBjdVTbiHfXvSMN1U
YxdAgCO9lzbnVNMD/pOThOX6AJDSImanc+JFJlfyAfufSrLQDGEoTy6XMCOjL71l
rJcsFL1880nD5oGkp0IYqRLBs5pE8eCoeP/mVt0NaVBS69q5vM4oZm9yfgq3b+/E
GA27NUtqesK+bAVUh6L4ufS7pgX27Mib9leXJBpBkWXG7c+uIvGWCofvunln2vHp
d5F2AcUe70KQKpx9C95wPHsUUlPnLw4iK7WezzpTE9CdUJKRucNYl9uHgaw0nnNx
jKQRAB4pbe2UKjfuNccD3yVCWYpjwc85xEeYCDOw4FtzETl2Y0/RfLlaRIXYVwFy
OwuWEEdvfWHgxvGesD5BKCcBKtsHdmZ7N/7iwFawkB1j1xoFXKjDDbmyPxMLsb0B
6N7OAItMZazzXNxLsdpFUPi21MCVn6lplzrJiiD+ZIt/EhEninoZbLiH+suMoqLP
rMu874TbStQ5RAMufbL4SSYHiqwnzeK6jfJSPJt3Gquh4maE+whhYmPc1R3QDpzY
AMd1yVtdKQSgQbkGca2gu6t7y51ZS473QtP4iHVMlWc/p1BPWzeTnJaDDhstuRj2
fX76309DLNEWsf2GB8gKxDyWaYgfXyiOhBQ23tM6GuGZJpsdGVJih723avLFpm9g
eZkodneM1gxDxufoWWvZfWwXqDNm/lWQ/yK9PmZPHpyZc52m2dp14u+NsAPwCTIk
SmOg8Nwh0Os5+XCXpeSTGn64am2rnTiD8naDo8lvkNx3j5TYWIEbNso5olD6UMQP
HTQL1CzPAKsTvDysAABDE/Tc0WbZfvc8/t0lNCSeON1cPATosQkNshGNtpar063A
XZ9D9/n/ePjWSFJzR2DYQn3bzEjujJa2wb3Eh54mqX1yUqvLd97wq7Ju/yCc+i58
yFKNWC1XfVU9MXrtpgqOqsH5PCG+D7pAmjVMCzBaXgGtby4ifGqD8loGogy80VkS
gG8uuGudeJzJGGNb8uMDrpSF/fJV1p7aKtHhvNuCq2FuzUYU/kG1RGlqRPDLeMXZ
cjn+lznigkZtIAn8VP0r66seRhURa15KCdpTGZiuicJQGxxLWJY/iabWVaeI/unG
dRhwRR4jGi54YPKLqRj2gGWh+iyOhiNDgMFDNHQQLTkvTriq14XBUo5H57aNxDSN
x0PxRSXNUcsrhmsRm9LNJQC0Chhiq1Xb8TgtS/zncKGiX+TTzrhxljLFKZ+yI64t
LqBbIGEcKQogj6VuwGylDG3hDjEUkzoU4l+NNtRfcekWCXx8EVTtzMf2STQxwQaD
PenDanVH6iI6ysojo/sp6/01/X2/JjkP7JWb2igPn5v2Zb5UX+URNPFRpwWUs9iK
nIn60pYj7JZfkrwsQQwOJuPyg9FF1RhQnhHvmc6WRPYRGTDv5rjH2lMhDMMYcPwL
nQzDqENiLxMaEGZiho+h1lNd0QjKd497oJGQgKGTEnQwmzadpQwK1y4DRQIMmGjN
t4+v6Hp2stb+re6hUeZIOBfUBKtHNF3w5StkJIVrWmtYzawJ+fTotsxMPyJY7a0N
rHj89HD0ieFIFQPE8lR9TJRB9reklaDBahM2w31XFSDESLafO/KLdncSas19oAd6
v7Oh2j7LzAyTRo5iDVEAReUdLpOzXOW93DfzqdBwX3ngJSy9PMn3NMR3xVdFln7b
YO/cLwg9XXaWL4zVnmuT+ySeoCjPkuGqFalp0MBNj+LNCj942ussieTuALYskLMQ
jHad8UyfRMywenQraG6cTedvmABPi5crupCMMnf7jZn2Gf7tsG/r6iwZmQNAx2eg
wvgpYOF3p8ZoRFIQahiqdNIChJSC0nQt6J70J2KLU8Ij4+g+Klh/xvwPeJThhCqN
A8HbxpY+0OhoIMDVkq/FPbb8PB9MrL/zQQ5hZ1ePAgje7MNn2iwEuRD9VHjVOHhb
zxX4AQm4j3HBhgVtd3UZWiEYPkGsKZnZ8G14UezDJXmHNrRYussUNqY2M83cxTDx
wv1vdWVFRMctfmayN6LJ5JtAQRnvN+KKKhgpvuXl/6xpNEnr005oqxmNMLzwa8/K
nPvQnKzFjSdZ9KkreAoAON3sX7uWfDFUuf8olxqPffJHwoIe5Cv7Vjkfmg95m1KT
Wv0A6Zp0WwhA2dljDRbDLU/NJMtHXTjnpwt+fA5z2MKsockBAHPUlZJ7jnzybMN3
wYC0s7XAK9FAy0Nmp4DjuVL+tsnVhDMDCeJm6M9BQ6beYQ0M0HUO/kfVVDgPfRRN
Q8YBCTIQyprYr4GICwOScP0a+jGSLYjlt5+M9GmnoO00+ANhPKOFeFuQOLMTSrGB
yBNx67CBIIO4Ig1FPAG9y6KWHY3jk0ot9qN6pJdJcgtGnpu5yuPk8Ln5mx4/78qd
GSu/cJ2NtCKNy2A08TtBwXCO9KskEg7UkcMC6YYJmkV/UF0/h0xA2PCNrOm/YrVZ
bjs9LTk9m6kU3UB84PtMcH1X/be4r2+RdBx//ZgmYWymakRfB7lM3IKaAlEKunNQ
7mSY1/LuulWbDLqawD9O1LdPmn9Wt6BrivmcMvlWN0fFZYjubuM6rShiqXt3JBhp
6xggn5iU/lwPXjIo/CmLHQ16aRSq1VyquaeOATI0fRae9C1JSLG75hpbRN+T2XIu
wGpBq3mjATvwFpgRJ8ZE5yFQX3zaSr+B1RJ9GV195pUIgyOxpfc9bVUEW423Tcum
R5GEjUL+TFu0fcQUOIg7Uq5GyaZ8Qn9EBeiLb9Mp15EBdj+HU2B3LC1sfaJ1i1fh
GrW/Lpu6cp74Bb8ntCBHfYBv07Y/zgXq8Knxiwwun8EdC6OGoppLm5BS1nVWl29S
wwUNpqrHOX/uxivw6Om+koX60tqH5HFY8ZHDvSmVWj8UVpiDCwtwDVpADNaC/G6N
iJCpqQbZKSWUsuyV3hTDHFaH89FGQ/asdHt9Ap8whcj1171nXSBhurE7Re7Az2zE
X19nAJpVkso3N/7Pu3sK1D1+33V6G8T9HDugb+UvOolSPLOfRfPTSbHfy8g73UQi
+t+3TuoEh+dMjxDXiG5aUStsEQkW7lI9+s1C4OMYn6lj3o/XqfpdnRl5fpgCgMAK
/4emX4cMpeiy9nKcfI5MawkdtqPrnWgpT/FJOD6UD7+qQJF81G0CFC2As+M7IXK6
plzsv4uh6013hl6JIh8G4wHs7S8TvcZCoKeOc6JrsdPwYX14o0+EsxzP644nziuF
19hphDHIaf7ptZGVJHa+V8hGSX+T34QAyGtylAmB9KAOsG3KS7jVdrx+k0sdgUIu
u22yvdgECItBn+6OuPlsVGskG6Z7XibJErR6QXG/uSTHUmrcpsq//Y0SZdmw0X22
n55rStLuusQO12lVq7MxlmKdGdEqUlmy9LVWbnUktJHZgVvs1mMaeIgNqEFK2/pj
cL1C5WyGtzck2sZPGm9Q64sKOtqzZuOWM7z6iUdtURdajK+JeIQ8o1T8nwdWBu3W
/BSs1og7rAgd3GxTw1KwKn1Xi87k3fOtAkds0N3uVPTTn8+Ll+kplts4X4bsJQwi
z850X7NF080MwsMqVnix4yyofNfXEkGV/XOwOLIxAVhR7tfGEXwnQoqfk9rZet9F
XU52UitA6bjqzCuN4LFt82fJBSnhyfXmV0j+nxIIZwfX9iQCvWeccimp9csGDSue
KOS0tdcAb7SC3cSzid8hI8pzXkGnP1IZAreMx3ieXeqI/Em8j51PL8vyPq5GBMbs
cWDo/G1/bajloGCuSgDo6RdKQyxXjxddZljVfp7NTuG8dG0IYapa7320WjT5TCcl
2cycK8V1qoEvLb9yOLWDg0Wp1MS0yVjQgrM5jSg1L8b4JjqTnqv8YPECnMn4ln+W
/YShhwlNjNXdXUaATzpQvX0srzfvY2aXFzQP1h9pmNrzu38542vRssEj++3WpZPh
qOlWcFZlIjk5ngoDY/PU1lBYQvfmgYy/m0XfVHtRkz0qcMrXRHjvZYbrRsJ9MkbI
ACvgrSfq+ZulLJ3D98XBdHrCSMRHXO2beXyioJDDdNh9JYuJeP9KLRPRGFl+8b52
yhLin3gME8D4j0XZIwBeXEvMOyu82kx1o8rF036IJMbSu3BshR/mZ2/PYRTflN/X
WvQxrNgoNkW0ic9/fkWiTmnhJftvOly1ws81ZyGFUZZyaSI8Clupf8rYREO63XPi
Omj/rkLb15mDcfJllzWhWVHb5zpwwB4qiDf32ipp4W/RiCP1d92CXWpEjajVAEgy
MNLeEXKcAnK4Oy6ERcONz3RcXgmS5BEENFm7+eaUvT9yhoX78KmxIUwGaffzTihY
CX5i4/o4qkx+wzuOtfu1AGqquMcYH4xaM1g6ui6zmKZMYRkLfDzm61k8Kkja9u5g
tHoyz2ia6ddOGOtakQ1Owa/saNykp92iSvib/6/dsow7B+tsDbdPvG/okqZ8mnW4
qcujKKJrHBj2ZIUrZJh119cUyZd/g6A+hYPbkzJHXR9+8EkbGzNzmYnMAgdcBLzl
Vt2B2fvcgrJ+ZOafqs/nSGqRvQHjo5W5YsgO2bkzNU/vBxTNBN7fVr6wjql8jY+1
lRWGuwBB2oqwPaLdiYfttLU7laPpVt+Y2a2rGK0CCG52z0OPM4i7XSGBMZ6VZ6ee
7EvByBI/0iXoXAZ7883J2g+SeZKW/4WdZZPcsPbDkhveHop8usP4kS1pq4C/rulO
8UctMorZCGImh1H83g9y1waSaDJAINQuHnY7uTf4uHWYvgqfNrAFkJRbIL8EDTzM
BcnirMS2GIMCZnJOT4CILcGuELY1nL2+j+OSPx7P3FY45Hhdfji/PkNErl7pSc90
oHNG+mBvrYlBUMa1tnfyvm6om0aT4vwxxbuYi/12W7dg4plA4DxVk3uUlPL7B1hR
KJE2LfcktNxRhIuFjxf7PDD7xPUZjIW6nKYw3SXYF+uMWADTqh0b+MpWH4JcWVac
ABeqj8KrQJKsOpDO8AIVpB+Hd5cc+8Pmn7802fwm5hZhYwsu7mel2FdS/GGEDhlu
Jm3+m9bXe1Y2X0FYbZWFc5BCFwD5yD6eHOYLxUdn840+jPi9Wnu9CAxQpbyGL9N7
+iUWb6TTfAmrTshtw60t3XcsPINghyvr7dK12Pwofb1EQf4OIDHjNWwDPiF3EaET
WgS3HOL8j1q99dcoaIZKPhHQDcmBxlIkn6ioMbdijcm6G3PJc3A0mNUjRpmb/F6R
T7oKec5lwrmCRhL4Z6weNjbqYJA3ZnnsVT49pvtHspokN0ulD6pNo5Uo2FUDY73l
e4PkVju50GPatzbM0R1/XzAUXUrpqqQPhH2/sazx+TSOQneK6C2FBLNjD+fuuu7t
UISuFYab0rcYq2B6F8xUEgV51J4KUe8CiwNOBydkQES1/zjduz9oPztEvLZ61Gur
Q/8cbUEUhQwrLtFm4IWIiqpt+J5z0epbADU0xUsCLpNeS8YDxsgrwuoPnANjYybW
Kly1irNO6WklhcYHzXcYD4MP21tkg1/DimvO7L0HjV5wxY+fxeDLvqepbSkknk9a
F7aUELORj6u2EphEp8tMQX8JJUSyeOfpQkBY8z3Ue/66ToawSqvAPcX5nEY7969w
jJ2i2GVsJQxuKlppTToI77hdAxPzMzp3Xxd8+6lsTg/W02u5t/5iany9ZgdROxwG
Boz2eEmtUeiFpErgy+DoQBrXVMph3hlqpGIrnfowTaPZb7KxJwq0YlqAUvYaPtjJ
49KYGpp+igQHK/WvavWpYdM3vKC1cUpYKRO+X7cGlPytWmA6m1xwl35bmHlHisUW
uO4LKrqZ6cjEmIR5N4qfLT+eABBj7tjgg552QcE5OpOFSTGoaEycx3hqepSXhwEP
h/5c2DFzfF01LsYve3UV+MStDygjutLHg9bXIery9p5WGNT/chcsCrDhLmRSdJtS
Zl9+KSAXyi7sodSiZBl4bfDiqIwnSIWJPXExHRYP8UaJSyirun4tyuVeoOpYXiFy
XzR2zVOFamU0jhWJaj6Vf1J+rvdEDJfBQ5061zBMsNtDzX9Sfu1Ko+8S21np4PCd
6kxjJGYW/tiyG2pdPBzqEMw2JH84M6+KOi5zbwGJ2iwy0EurP/ewL1OZcqQ1GrcV
w7GHfH3NjOlFUfjgEL3kfjZ/EsO+5ESOFgaetyV+GMFvpgWQ/n+YyI7rIa0kAwdG
NAT8we461/+VT2T/HjI8pS5SxxnCSJe6OoiaGJn0TWTeWbt00Bba6Ci3HV8sG0SN
g2C8FfYeey9nzJetlpnIvCgc1A1Z0UAkty0ve+4ZycjOajzNwhpNrBithaj0LPqe
2d0ipmv088RKl6T87nfjkQFtZ34s9JBLnDQd6bGrvH6QuTzioRRwOB99bMgRnOoQ
/oQdj76d9DWPC39w7gyrQkflIlR73769FjHGsbbDMc/KuWlcp0s9VAuvEDGxAXo6
6IwLOjKRe+a317jalRCm+2yMHJUylDbXCAxtv7GEgktMVQUSskBaPY88G7UrS3S4
akRcsl8P8pYyUY3TDPN8sRHGnSJ/bCx7yCwCsyaj0dM7QiR4UtAZquN3E+16sj2u
ZiiilQQa3nxPIxh9Neh9PteJV7dqKLn395jCJUIMFnTAEGwWSAzEXiZJyIEfmgAX
0Emwq4kCJ7MS5rXORty0MheHvY4omvE6UC6ERtDXGxaHUcN0lGqBP1wxM9km6QN5
DU/vTA/j01z4knFnuiLARyctfEvDYGSgs45bn/MKGdHa8T6KCBRpxnyC4PmIsxGj
08jvmxJi6l66AAZozxdoangtE/THvTceuGxzB9kEVU1emMOitU87jvQli93pRRL4
Sdb+r3anR5S6oVnMm1kd5UqprWZYqSerS1/DDKzejvoQnfsYXOaZVrOwPFFvsm62
eQEb2VGRCiEhBzJITZgUYTYYCMD63IbC4/BDUHa8qAQxVQ0QNnXlufE6ntVZz4fP
JRCtHZhUUroRC1Qc/1Ml/WKsIVLqV7MDAYhgELGanD8A+VZXvg88VXKkQpfDF7MZ
EeE5LkDmHibuCYEyLVaI+w9Z89WEbDh/vegLc1FJIBv9HUtt4KUhCR8RfmHWTcVE
aSGbQivGSGb2E+sPh+lA1G2OVB2JM5LsLSKZyYLzPOZm4S4n4LL3eEfRWbND6rAW
m3L35dwtju5D8eBCRgC57SUeH75p/Ue5t0AUSeJx1uJU0uOrNBGCoLCXTTaTMejr
wal2KaLuq4f+JuRP4XD2W5Rzb3d1NOV39BQmU7p3QB7R/zdK3vhereuQs+3y1C9b
io59BmFr4uBfLVYqYhPhCjOHFTxkBk3ES7a66/RRcdjwp5gkQ6ZboivZ+TYu6/fA
bFBblZ4HfxMZZwLdhjM3yhkV42t8urMwaJzioRbRMTEr0XGBY8eY7LyNZPnxwSP8
pWjZd3FG4vtHvKXmRvmOviHpi2w6yJHCUvrZrlRlHwRfshnx2jAiyZWTrZebrGjB
ZpKd+AgsFvEQettgyKvVdOzbV2mdVItUO0yZ9uolqKzUqp6GEu90W+4FFBR5Sadj
QDZfK+Sq9Fb6ExS9h9o0pD3GouFcgeLbqELxQsjnojsNdtIFP1iT+9qg1ZG7y7hP
LiA8+8hJfvbgXsJpvqOAaqsd4Dw0GuL3CbgRGRq1hcR55xKjNH7JfOtQ3BPSs2bw
DSzv2yvqHrwCIkMlTdJDgFy/VffoJ+bhW8XoUR/J+AiTnSnGESCO6toyD52eLKC/
+HQhLQeqb29l/RInZLYGr4poTq+MaJm3S6vkL0gFdogVuJHHJrEA4XL5H1dah38o
LzBKwYGfw1tKTN3rwaBCkPGF1gI8eQExBBZdw+IJuAYTBZzZp4AvvYhpYJDc9hYG
+1TCbh8yHQgEidkpaq5nG0LZBvfRhd50sHQm8QLhwxmawzRT0is81tMbrLxZtFAo
Ah7egOmb70DvfMdUR/DGOhR+B9npxg3NfREDQ/GfhlqMDK9njugB8x9NGTXPmp1a
V3GJuC6qvpbjErOChdnDDKYDyTlsOXrJbjIhLgKFag51/1UW5DUM40bYnB97Yccu
fy0i4fHJafQvVw6DslQzrLQH4J8F8Jy5i/LC3ks+ClovXOSdh/h8etO0i3onRJDG
NFn3SQNbOO50WQ3KXfQNgV+D6d5q2Nwd7dlq/J5gVQrh8ckXNv4AL5Etms2nVaD/
RrB6Qc7BCDUpLx0Bekj5oNYBvmXwpBCZe4PgET4v+bgPR5UKEbcMgiL/GXwKFeBK
RPM5gLWubkqdn9UJUJuDFyc2cDLXeGleCEggDcjcbsVJI0PAACh3U24fgs/NnC+S
HD4+rG8pZBTc50hjtnlQlXAbjq0fBt3nAV778cUCzoQOLLRyXhVB1hx3b/45drq+
u+FvVrfeJ3hQTtlDtSF5ajHFFI+Yd5ql9j+4NboBqNvz9KY05fW+N8Ls0hosIszp
Pg4OGJ5f0rv0iZ4qg8JnF6eMHvHTdDBH+FR/bnkQoPHBb/B1oYw3GvgyJcqIRAYL
iRUM2ygfrlyIpQPxQ/IafVLpajeDfLZ37tV0Lmp9fxtfOEqzqs3mN3Yp1LmyXi8n
xEUQoQ9lX6LPztq7zF7FddrnA3Jf2wYC/AagXBoCEX3F92TfT4h0hu+M4VzVPH04
MeF5mnEgYJw+F3V0J6U9ZJ95Nt2T6dkXY8HPCkflu5kgAB7ymGIl4V2DQFC6OsMd
1DigG5ifgqrdoaD2qfAf6zwJr3jGmlG+yV2ZOaL9ixG6XaWVkO68ux3n/5I7lmfA
iKCEoQGVBrJrECbiXnCdIliXDEYfxkEfdTGuQeRnF/x80KF8hNxJ3FYw4jQLCydE
1gAgwM3KZ1Ka5c1k/tjpsbN+13w1ImqbNNyhweWKPg5kVYl171jYbTITp+Ne0zXN
LhCkpIQAAzJYwHx8XunqNJDKvcAqXk4fR9iEzfLS5ZdPJyftsqgzyfwrJqpbkW4c
Ze43CD5S/2bfve6FwjAb41jdbyiNi7i4vlaix5NXszLnaFtjhjhE9lcqwNd2sii7
jkWVjRpXEtU2plHfxeOOT6X8ircalE7tLKCnsC/HgEpEYeky8rpwHb76QthenDNo
jNaFwbfsdigBXjRA6Et0CSb+5c34IYmjSF4bqlb6GQ5y/4KBwa3TGKjG4EMmXGUW
RRhD3ULYTQoZlShnMC6uEXR8RlkvKbkdREJwHcjV6Jj0rF7oTEOx5tN0fJxa75zO
hNdXyqzgSDXJ1CrXNx02SscocyETa/qgTcSqfokO9QuaYPRCjnYwhq90lxhWOSnz
B30apS9VOn//HSmg2iaWG/45xxhD20DQpefjd40K59qSyWQUixC65aYKmiVPUnkL
GT0lKP/X8A9OPyMlXXKCWygNJzMKOcpv2D25Zcg/AX8i3/104kV99PthDrwUhXNB
oWytdWiiuZy31xaaHIzDn3rr5QFy/mXRLVX+PYe1sZ20eZPpRLYDQfyzp80K4hoQ
K98s19egriSmtcnyQFFJ8PV3G48R9jAnipxCi7VgW3SbckH6ReZbPU93EWNIazvu
AblYlhMOCVuc/tJYM4W7DNjxleRR/a/nOM+9AgOlM60DdXsgEH1mwudDVbN8mtks
vvC8JAFxS/RifbcC86P+UC50+E4Q7DiOv9bjx9MzY0CkF5IaRC+/ash1nI74/iqZ
Pasgxyl6LBinMuP+oz23gykNg/RfW51JO4HEq/n775bR+NvM0b3K2K9KkaQeOLNS
u12pCznE2TjBeAhgB48BEjrXo4m02fYC8kbQIm5m0puIks7xDZMuKEdQ6NREcRKX
6kkyLRldOYVbrSMdc/FmnHespd37iNUicW6J0bBCWxaqzwGwU1cnm5XiSG1/n5qH
qLc/sjMS1L6+AFV37CLk8IB8ljD0hhVc+OB9TVzSivkH33SDw/p/SFvGHsYqq+QS
KAuXQc6T6fIaiFFziLP6ulp6sSmbY5TZXVZFqQfLKvepL2J8M4aVwkwczALTB/cN
f4TpU9bEz/YTuPL8RSB06M76DCgeOuBVbK+bZNJBYUZX5mBoPtmqgjB6cIAhCVZv
/JslQkYGVb9+f+Xu0DfLUtXku7/vbyUBVzy0ZPvt2e5pDtbBHk3lCl8FS4GIjWCc
dwxg32pY0G5iRfFqhP7Qz6SsTlMp7woHG54beQulLwP+TtpVwW2w/ngfFxEahfKm
VzTXf8wyDvWNKgDHWDqJ9Ab02ndVSzhvzf8S/2dCUjutMisRAlsROa5epZX3PyeY
y+cFTRxypF+5Ho8Yu+r+zNeAQtJln3BbApzW92jMQpcTzBhFqYnw2DrH+7+LOW+D
66F3DC5Km/B/sdU7KAnxBDjNCfi3bMeJ78W3zBx3tRz8ae1AUm0xj5ZsxfD96m6U
eJE6MV5NhSexQ22Mjk1K9ysDx5L9Fh67srInsqd4AgdS8fB4edZ64AxliplutAVf
p/bXXwZno3EoP649YOznfFJ81huJDCKxht6rBev9nzx7HOPD5zms8Xllu/90Eb26
0N1iML3tSmjL3xXlxGJCHhDmmX3TrDj7A/k+aIJtDCgLiExiJH1hTnyzK4OCW7v/
yRGgOnnA6TWOIu2McDYiH8ew5DeW0CQ6mE/Diy0vL6FSHAVpF4tXM9XnlTL2lFfY
gRYtri5fFmKd0EE2MorfjlhV8eMpJsV1lVowq+85bUDWp+ZMwyeaGSVbtLRmSjUr
c6Ybfxp8gfTrKDUDUOqGcmzxdJXZjVvwKsMMc46zHMU9wuSHwuQWAdYa5xPMwkx4
CSbBvAiFa7+FXoRrjBRpuEp7M6qnF4kGNEnsxCOrHLRitqKphaFdQ05q4dR7NkeV
v2L0HXmZWA/dKrrQRlvBM6ASsWoJmin+nFZv3nr7g+LWXCJ1jKI4DnGzqQDx2xWE
mKOAQNJYKt7HjXJukyvy+cX3SnxOehLr9aHJzPjvftq4QlP5N0eoPRItDgX73bOl
tF/2lbM7KUQzf6ocpOqnkajEOy/e2vQ4dVe/joNKlF8mcFHK4H5RcLM9VLMmJc69
ghAz9wd796HWHHLatyrQW3f4vIc2JfpPNecFDQpLPhk7v4h5c/M4YgStU2Mgy0SV
YQDkuU6FpVNoGfaa3BWka15oWOvYh8DVWO279NM8k5xu/F/brxIr3nkPnlB6tYVS
lE/2cDjPThB8POEQoTXB7bkUgPQeO0vE8dkn7JcsSnutS7HZ8FhANgiVi4OfURpE
S6oHLPJe05H4xtjsA/+SnmbOI7kRW07H+1gcBpb48kGargCYLruIfzJ9hla1yrgi
Q+oWy4vsS+q+1w9vzCx5nU5D4Sx5vAoN4qjn+xNS5Yq3MF21pSoeTPouA8kYZvpU
YdacqC3DPA9msTvFYB10mA/ZPyMx+YkxNtiD6UiG9sO2J21u6be1vSM8pKvstUCC
nCDoeWC8z581AQZNNTXoAbJ+nI678Y8ttpWA3z+xWw+vOw9N6pxfIqbSIChFLRN7
meAN4uY5Io2B70+cpSA86v64Dpkh0URxRWgg2C0GLMp95Y4fc85rruDYRSNJqarQ
2W1PP/f0m5ueXVPRfBpzitpzuJX5Wzv4sx36wo5tSCcR8hI66XN+7Ix/t/i23rNj
w5gnHA6dFc2mEgK+7IxZhffKit51shDfvU/LE3omHjMH71UHN2qB05VUr8anYeZ0
hQwwkTLkiYQzSrLrGJfbvpESFEMBXKUqbxc2tqY1wiY93uU1tFwnjC94r8ksBAOK
H5ewRYU50M4VufpPRbZNu9y3GP8CDoE1ke2xcrVW13wa1JIdbj4RceaD0G0FsOKc
Rlk9BJUa4VYSLemZlf7A5KDIBL0QqxEq61b+prlkDjlM6DncxqvjPEV0PpE3P+oL
MTLrMCuFpJkrHDC5WrLoJwAYsS3zYHieWj4kcfFTifalemlGddYUB1fasQB/X7uV
Ic3rPh+1FMWWqKQmkXBPA5mEmgcpkOvTt6rbouI2kaWokCaAmvlOolw6LLcohdx5
yrg0tWJ1acwR7YYrUxbFOUCzXdMMxyJHrp4aJJZrAtG4ZCMytz8BoW/BLhDXxAeZ
K9UrJy9w9ETIMgfLusCGbvitijnE+ttoxAaSspn3bxyz23YkKk23+QDeo0ze8pBF
7mHYokWa1SNaZvdN15Cid3LL1qqZi9wLL64efEE4guJCnIipLSWC2X2rsVYOhygg
9l6WCbWOcHRh3lQN1ZdBSWmMgb0J3MHpokd++jbLp5SwMkDRCx6WPhGkAr86/qZ/
ps0RAbAuUsLqClK+0S2ptJY4yuv5g8DfU26kwrz1G6HIi8OGckLNlkuKSXp9HfGy
5DTbX9oZNt7jn1qFmP/pLLEqajhnLEDKgBmAg9psTBvkv/pIw75jkzXQcxiaylOn
n9LAky6ZJJ6i9mv9EjMVO10iNBLOmoK9yUlP3xTzKQwmbP44+D0lv5V8lY2rXT4c
gmTz3sSfB9rmnKzy7BtLceYSP77X+mVUZiz61vZjj8Cj0GrITpH7qWqAgPsErDHT
gCd0zZALS5k3kpngb53COHHaGz0AB8dUv5UkX61UorWyB5BhDDzLtb7uI15MA3Ac
vYWRmT5EtE+LPqTAVK4zX4KiWJ2mEyGG60qyRG9Am21F5OFtP0wIqVnnzbEmOuVl
YtbXwrwV6J5+5F+hpm4VYDOf7dPPmHPy5Pdgu7N17f6jxwmPNdMpM3I8n6HJeAJJ
bGlKGVwWT1j7IWjhIo9nxQ73XYVafM7+TuphbnNyY6hRM3T7r9yVFSShwvmGqBSp
kLxcA8quyigUJtoCQBf7esAcBoC/ffbflzb8bxeJ0Co6RUar0p/37IwV1smeUeRt
S0xnNVIle2whdg4xnZG15N5dLrbvNjRXBaSiuuQuURWLXFD0wlndJ375g4EJh0kg
H/u4cWYeUmrhcVM2wHIemCj1ZCB1YEeBIAJo83AfGuK0bAEMe9g4TLu8K0QP8QN1
qeBkZTs3G+NluRf1z5sQo0eG/oc6pmtIM8+3qqRtJFaSIXqTVNmcJSlyCuSvUKWt
T6j+mvm+f74JMaLgKJynmeEv8O0uMojjwMby8SQBSv//dc3f6A06CH6nKyVWmMc4
kXfNaUbWhT3c2h7/89aOjWSNRVks8Z4yaVHgJRIgyhD/lZmBdPwq0nwgG1zg7MlA
iU2v6zGFwlgLctX+zLQZ7yIV0aeZO6V2O+N+uNXI5Of70dvpUuAAX9hq3WRF2YZ2
U9yBa0l+N7mU9L2ZsUUNJAfxrq/11ZUq+X8JQ3XKTpoY0K73dtHtBxmX2TQTzhTI
9GZRp9yDBHBv/BZxtUMhq8kJakxocQ6sOGr2lkD0BTfKNSh/Y6UwRLBa5PNZUaRT
nwbxPUdazNuifukRktiMu7upIkNkQt8uwOzWGDLp1r+Xhhm0gOEYl7f8ukBjNGc2
fnlOUcFOfVtvrbw+WHB9zFfkB8lmQETwEW8R4KGmCb7xW2PGq+4tOzBfJ8GWPyqr
1Sl3K+JNU5tzPZGGpE6nsDes2S4zaus+q/9tZaitD3w0g0iV0ZRPA+PW2/ZZcqEf
5XmsbZ51cx+rJN0bn3qWdaue+Yj80Bcr5ZW8rnP/1Dvm8axuTA4haycYKfOxfrDr
s5cHLSe/FDGvbWRYo5ElkMcNRdBiJlRqS0Mr93PWxT0hbRAEbnk5KzdLnvYUazzv
IIT8V8o3EC85LaV1Ni9zI+w7U5rKYTwlhUV/GMgDdR6KeqVBX26IVnSs2nuhHtT1
6UvuHZQqYzWhrxbKSMr2kWe87IbT35T5vYSGRy5/bVBX1jGwl98BKEwJIPRrMWqh
XfIwMHd4dLvliFieN5m9t5VR7F3SQTsoUYmkAV3oWHX/f3GOOt3nZ8RgWmwU/Cx+
nMHjs+NNvMRFbXyGXvK3op8RHY53KTldyU9NEntzWKWwkdLcAqurvx1rdlyos5xL
q3ONsRUt/23n4J34ANwr/043LbUpr7IJYHrr2BF7AqQcuY4BNOhz+RVrH9NTMw0W
+Fy+uwnAgLA2J6HWFB+XUz+Ua18mhVgcrpti5wqHCTxFyxCb4HjNTLYJCLX6mAY3
UwKgudLTN7G/+HBw8dnHh+wcuWtjjwJJ2vNKosbbNg0lJSDk6C8Yca4uDC9H1+Kr
3qDpN11jfk6LcSYNf6Zg9LphAqEoA0zvz18J5Gcw6ikGgf1KU8+zJ0/uVEZeGL/R
a/dCOuqpzKDakPpCkVC6HM/5RaXJPbLXbSxOx56UGLNeAv5exXeYkv764Hg4ogZ6
Tpst5Oy0203k3ca6P/Q7SMOOCVOdUx6w0u6drfdcB8DVoD1Pchx4ot1brVXw3rvT
PmtJit3syycTFcYAjdTM096ZgWcvpcVOIcaNNoIjvATNcT6G5APGGqHZ3e0A9B77
4eZYOuh5XYd30YLKt8nid911smJOrRp2zKpaq+ZQnj3nAjx+UTsmMZsyLIlAWFZU
hHP+b36KNlG6Es7xKQw1QEmomyTCeObnWywmI9M1YI7gB5hMqiG95+h7ucDd+MNc
Vky0CPGGJNrMlgm7PLZhl4rbUZe5sCSXbacJ2pnxnvcRsAP5lSupCl62aNtSK9B2
KPaxxRaH9nPBFXhIA1BCVskW6x31swJ2EO3pduHJvyV1i9Cx6+rapcY5S05Fk6Vq
EghZrgKjoqKYEdlpuTG67BxdZ6/QdCqzLXbZFT5YBjzKoayD5Lsbt+WeeJAE90Px
+jE1+236fFDfeQw+Q2qObJ6iKQTpfUZDx2ipDrMSKYzS14SfkDC3QPWC/QQoQ8le
Dgk+I4BfaZdiXDLm5HhQqul9JdRuqxv29+MKwmvvgKm30n4iYBgl2SNGl5GGC5vG
1JU13Wf0lkLDoQpJzBEcklcXTNmMpkepOi9Xu9/RIWd3D2VJWt/T8N4oYFNuYdhe
GoliH1bJlHRXikpR/6fD5SMDowUqIqaiPqBIN0IGnG/iNCkxSW9ikazCySHwTfO4
l9XfKiZ+ekR/kxzhbkeZFGo4pwgEpMn7uWmorsNF8FNr8tD7TtZIfMMgJwldSv5s
fZJcpWrf5KihAq1d7DirrrOq/jipmAbr7tbIvprQuwas9TDxhLB/kNldfGGea9Qt
kEjCisRSR6NmVAp+IenVEdD3EwjodE/PIKow2dX+NCap7yda+zvTTcIsapeT2Ru9
nZGwFmE0D2OLeSZ3T97mOY8g6AKF7vG25ZQlpanbNPmLlpyppwIQRivGbLtPVkqt
kaLnq4I0d2Dk8wf8e1AhtCp03JIOqbB8kWXq0/ZTfBoBjG9/jsMuSBC4TxIbxeP1
6D6yAVvYtVPacUWSwOCFOw4OF2mMwQooqODusIFXDHgA4pfaVZAIDWLG2ZyPt/4/
04ILq7X4ZhQx8pjiWdGyLrYB0AYHNnaIKPpWd6Hfu6687Oyyp0pl7cPwii390UKe
026Dlup6oFAM/KDpAL7tntu2dysT+nuv/NzoogAaKiUg1CFy8OSrSI/dLUTKBg9T
1pPRbTDNadgpHkuLttVO8FEDGwOmfoknngLbPnoNhBOjIJxFKMuEla/gj8i++Ptm
VtWBpJwnOM1SGVVeGO/U4S4zBj+fyIpCdp8OtTcC7v5/ildK7sdESRtMv3s/H+Z0
f/RC2wHHkmea9e58yC6ztAPGR21Ke+yT3K6veFrfA6KXHQzWsyRvIak6o9dWZcra
zPgq5+CmxGiQ/bx7xFGRih8MlnrepngNScmYZI39+InpNLP+9bjrt0to+qxgqQGV
+vPZu7sYfvJy8+muAEf55n2E+kJPm3/Yxp7xsAPloKIRjsvDqTFlU5Q2s3EoVncW
p6TwYRZdE90w+uucxodj9TqzyAFg5TMXKXUSy5HKup6QZ2ROz0XLv/CxR60eYfpl
IjkU+3VSS6Y+K+HR0K3O9+hJTNJ4vqClWEHI0xIaQ3st0++tgd14zmpKmc1ggs2c
j6yffsQWG32cH8VP1kMsqRXDonJtk5NF4Zt3sfS8HbW2XfzqevcHmACAMCu3GdT9
Zjjor3bWrKrzrmrG7ZLVzBJgBu6j/gB+K62Kod5o1mEx7hja61hSzfiRg7KQEUgC
5ZLYazlnkBNuCk6Cxg6f7XsdPNemOkBE7Nu4oQU9QyoY9ggb9GzBoXyxygPpPIW7
GOtO2bWO8C9a78+xICGvd7tSwLR57KMh+LZtaEw7NVjqKsYtrgsCoHrPJi/LTSTh
aGT330qlInRKQz+Wdws5awiXWLNV3ZMrCMRBySwOPiA9KPLSEmG5cyb45dIjhh+A
DHT41pd+na06PuHd72R0dqJafwSErOI9mxG9/Rmf/P3RaHigHLjWWFHKk2Ik2tdu
rEniS8ZJzROvHtgYkRmzYPc2UIG0e/BY0owW5DbO9ilDx12/2Nph5yK+qTHPZhPK
BT5zI487bwnR/qNoM6BttlT/GKmxFXDbFk76gwl4eAOQfHYbEk3m0khXdlBt1aEN
fWuujfpZMYh5VQd0t9pdd4ibHFarhGPxWVhGLT9d1tCMffwf0fEuHrdKrqnkpB5V
ChURuUZfzNTfo27j7p21PY3uR/WSYpcH5cMk0HPciC2eznMuLnUsHT/ssvGyO/uV
nzL6/oO9pxyDfPLhWNSI3sqoypRriokT6MnztlD2pDXrA3cnTs7EjDkZNBAyH+Ds
4zia/+d6UIF/IsCjROZvMPM7PfEJcbsKapZDuJMAltCvFylPDQPGjDn2NE0MckK+
K+k9DAedQUZc35XkOFIk1kSa9DGw6A9zmYu2tROXhZ85yDManyMqF+5A0NpMe6sP
xgBlHwQgdszZ2hBvoEOAsrbpMppQnJN+xRGXpvqWfO+xU82u9NPqBmgJsELPl0rW
SkivMeS9acVb6RSYZy6438QhxNZSa+fRqDGWA9CvHzFnQt83umiT975O0l5kWtPL
gUKGBDGBHcCFqJCbdxqmirpX/+5uE07Gf7wjdE1pwyZEisq2Q5YJTyfQ4+AuP0DX
ouyi0xDoDZuee+/loV/QvCiOm0ChK8HjFXnhy4/f0+PPk49PfRIXxk5d5JfUmMXH
I7RUhG+ryqO/6AIPe4lDj4xt3QLpPHQUGoWZfnPbnTgwep38MwUE6k0h7XVa7WW7
ozumY+X61QveYsJ7EJOfCNyFcOT3I/0f5CLFPhsI84M6ziFVhwCnXPiUNhlFJ7hE
IaIizzmI3OBrftle4U8oqQ+QGd/OxK6/G2KO+9lbSfTz31loC4wL6MP3QBDlxysu
9sBO0kkp1phT4R6rJ8c5PX43a35F7n26CGXXaRo0u3UPxuhqE0jSrJA095zQTFqC
qIL843TSCzrpChy9E2gX+VX66km65G3wRL+fu2Q1sXxCEJ7YB3ZE/wEWGQfs/oFq
nNL99dhZFN9zmyNtL9wh2RYTuuPPeQXRrEjbGQfqQjsjSokWFUdOsVBIQbhv52Lk
UZn9kzTqWWHT+fwY2iMyxbIZXg151JgY/x5IV7yZydJfoXhHIKHGdu3BSKR7katW
Py3SGJ270TSSUYSrFsxAKCyDpsXGRGpOfLM/2VpiLJRc7dUs5/4jTYjS14JuPuuM
evrsr2/IqnkBhZfg3O2aCOzHv0RXCXzniQU4q3+ZEV91p0gvMX8ALosvD7chlcbF
WLjg8zN8GJLjfvny1jE3nBq9AI6d7r4JUkrjSL5fL24BkxZ0ygJsHSw4eYEfxD9y
6KfAL79p5P6MIHYY4ZZHPplKA79bMcBv8d2lAC5ENwSH1mxgP3OIc7zGmdEkGSzJ
W1UXvKqI4I+I9hDSwmnU+i/B3F6z+OZpP8LuecmX2NaoX/TYnlOA8CUBEkRCerJ4
K2aeImC69ICEoceV996J7k24Dy1PmljdTFiPUdHO2mD5YLdVVNuH4uVg6na24sHA
jYiPfR7OOksfAwGe0N5ZZbBTXO2STswhPivRoIyfcoCtResCPUpmbrTivyqYmEiM
V5oeVdaJrzC0NcARp0Mfj1uReJKBv5yl91NmraQI6PgmQuaXnzeZ2UPszkzyMwpE
Xr/us6SjxAVnsacPoHQOswnzhoB9TGNK0789fXECFwDkzPeaCscWoWgpRbgYV2/D
PmOZaKoTKCpmpcRZIzZt0NwIi2Qqzf6KVd4wE8F9/7kCl6N5KUqmqMbxvBy8I/Zq
9aqRCgl5MJIoc4ya/8+OWgMZii3BKx5n9HR3H3TPJrCS0358QbkzBfVYYkQvwJuK
h6cqsuKVLbp6wmwRgNbc99WwkMuTltQSBNVni5eMRfrnKgXoZutEKNqQ7no0q+sY
ACa/w3qQPbhnM7hFP1FXoXXHI5MRx2Wv//cdsbVn6+xSaRRldjk1bnuB97D5A3aP
duvN8ia7sp/+EfeXZM3ypj6zzdubH5vVD98Mwn2/YeQKHfntUP+rMs+wjrB7/7gt
cZQq+jhj7I4x2/kiip5eqcOs8hqk7hlUlCwJ8W2aaSxeBK/LKTDnMb34oJWn4WXC
I3um8Ulpu3iVfvWdsdYIp0dHrlxRcXZapJNyA87nZdQWnJodWbgUhHDMtoRRh5tQ
NqnB4cQdVnzgZ1TPlYbOaiRKn2D3dalxWURkAlU4UDUMrkh7CVMdsS42hs2MYkis
rX3KTdpwT8LTIeD7NeoYNPcJcnvg/Bb+9cnv4UsLLdfeRWpWVzP9fTGlBGcnMVrF
/E5j9A4dL1CmUUuVJYVIXL4gq415YAOmYD8bDlsjK15/mOqvNpEyOWd0SQb1AjBt
M8DNRrqOY8MLtM/k1iITpwNOzfU/a8HfT6qf6kUOFnHZNGm0mlwWY9BS8nelOi06
jldbRbnxR9DHOmACYt7TS4a+rzv57Pj9XamTF0ZTQRfmBEQO2Ax/XamPrvBXf2AX
+NlHKvtV9XsrO8R+mqpskyp/TM7lwWI3C8p4oy8ejYK60K1nnyNCYqX46R60W6Nj
E/4zLS5GTxbuC/PZUrvhOKxNVfJGYWhG2FJjSZDdcB9XFOoMAT7ZFOyTrTdLBcgq
5eGZ3T97dfDEgmUbtqfGEdtY37Fk3PlHyBN4AnjetkGGMr0bEkLIzY5BPko8bkgw
sw52loqJ2mvKyjZx2XYeQTP7lAWJQ1Ib7agsacuMbEQrNGcwFUDmrAsZqTqkSZUJ
umpVBAqExNHzaIUviZ5YXqjIdtlty7t1rasxYfJgTN7XrvWDZI5RHHGDAjAP87iK
NpuOPbpg/Lqgqf62Ec/aFSyQ/gpeGBnWrB8DhxOtWKVRUwXI19nxH5mkQ76SQG3U
0yUwcdDXce9o6vAVAOXPZwUSurDCp1YKb34auAjJUWkB3WAQTJx/G3U687EGAWs7
L5uxleCRsKTDt1Vu3p1QQUrfTqOrkHeDVHaeD80ed03tj57a7VYQQai7nSW73o4o
2kh/hrMwbs5N4TCw+/0uU+GAQ0EY0ZtdU9ik63CozZ4ut6HC5VSnhSrfyArP5DWy
sB9BcEFfofcYUbgDakOqRb+FSTTSu75h4v2LtbxHnFSECB0HxAS6Zg2ZLEJ4AIp/
SfJ2coiMg6IeFm3EvN4ToM3Lb73eLhl8eNSdaQGLIEDB56tKRl7D9QFoiy1JV12Q
qJ72nOpIkAve1ODJF7TbOXy1DM91faVksoB4zOeDOW/rJwNBUD9jGc98N4XKEstl
BrSj9zO60bIIgoI/Fhjl75WPnZNOYsQm9Sy6Nj/verSO5UJXSB2NxVRAP81j6KuT
q4V6Nu+CK1L9z+UY1PFCU4PbLl+Q5TJRTYCNwEDX/+v7L4vXAqDzmMBGCbEisAc0
sHdtti9vBmdGBXYua9ZtARUyyvnWbeZsePYaTS9iclQlbsT0hVU+04rFmfuyHIJJ
9kvPZx2KLZYHi2SB451dZWZYNHciv9e/5MEdjdYybZKnoMx+ZxYlisg/h1+aC+bF
V7KiKlt5GqkIJs5liV9zGAFIzik+nIP6eyYc60kCTEWKPFUiLf/bHsU2OLtVKppa
ZweneLOuTaUc//e5C7R7OYbnQxfD9vFWoV3voLHIpw213f4Umul6PHcLMLgcbVgx
my/To5Lz3/5Wcx04oxpV2Qrii4tBUfrgxudv4E5NAksRY3uZ7xS3+QMv7bHLb/VD
BrAwJvbT6icZY8M8YbDI1vejD9pEIWLK9P/Qk9DHgMnZk2ou780Ih1ZnqRbu0/j/
NASJ7Q4wt/ri4j2pnJAYcI3Acyv2yE941RGQ3x/7+bTlBDUnP22gQAD7xZOOTtWt
OCrZE9nfcEs+fptRdE/DH/8I/cwuMln4dXr7hTxrIIygLvOWNCe3AdCB6oPFXaiN
0+aLSEdqM8W0idHB/znB+TcSh7TzRZ0rZpMbgCquv40FmGr0QkJir8PAfBEW9jfI
B/0qwskm/E30tSZtM/pVQkb+CHlwBJQqZQVN6gWuPeQYH6mEW0sqByk6dBGWVYlv
nMjd4qf4vedGrr3lsBEQYNXUK4w4hrNZDkuX/0U6EHYbo/pFzfMaZ2DxDi43xb9T
m73budpCxaAFrbjegI59hdZnqtvqs+SwxMzZiLNXNGuovejUKBAWHH/fOCP1M3Gq
sxtIvLIAn9wR60wRWedAY1dmbA72OrWHRjQ+prJE3ouie7esO376d3dsAowNRuwl
maSNR4tsXF7w9KJgTfboHGSNuZm2gMyVHdsxv9z1UKy6Sy8S+tUSIxmdjGP94CiO
+NSTxTXfkEHTVXI7QCChKOLc0O7bAvnFIfvd2c7DxwKPZdBCWd4AeHoudTDibX0a
VfjyCcr8jdCKDhmsHK7LfkrZuBpW5eumjpsOq5G3YMyo24xGiZ7V3VoOD75KL8GQ
/cvsFpZ95np/UAyesc14h9mxpOPaSMIunOtFetSLAdgX4EhELDkmss5FMo3ZkGAu
sH6f/PK8AMThTA333J9GVvhNGCoeTXI2qWpGH73Sqs3Sk8Th6gKqNzaWC+DF6LbQ
HmRmwK+v0CjWkUJRRVQC7h91YG6v1I87cfHYFXx5O/6ncLmzIm5siaml+HYq+7v3
CmR42ZJnXRmFZQHcczZYvuD5wlOuvgEqvQ2kn1qJ4RDkD5EblmbG2N4QIE6deQJX
tF1Jr50sRxeKNSaViY3FuqknBDPlS70O/J21L0ou9x/ORoq/iZuk7evmN94TF+Jr
TwiyFq1GtNOORLpIXOIJ6ILyNljRKmHZWmTio9SkRnzW3ntfwrkoGpdhjR5UaqRw
8uu1ewLPPqYWmpQK+mDApsD1tLFV+VbwDBoTN0qiMPZqy04hTnqWTXHBHFNp/jo4
a4NMYQmLfN57PK18AgWnV7FWCo5rwF0oGE5ChCMEqjNidc8rFcaxvqgano0w3QjV
ZjmpojxP6t3/m2o6Z+31nJPBMOfzYcRquTjORMrhZPbH+dFtH1Ffkve5clm2O0TG
VM4XTFxVeR3fr3ePTYwOazivmiqKR1cbldniInmfH7FelR/NG1zpjkutkpTcN0g6
0xp9YFaLiwXLpbc77sfq4VKLN8N5KErEfqBUO/awbRb8BuZIzTdMs3HYH5FFIAVZ
7f9vGP1zoMAIn6EHcyx2f53aNjIMxt2KsvY3FYVgFhmsBIGaQxCi6jvFXt7ye7dm
QELEytnuaOFKJGvMfKB4DFVsOg2OJ2uccaZR4YdkNMRjxW7OgVAdZFHil+siD8/A
+xvauu3Ho5PVf39uu6UnwIHn7F8VRm9ytV02mxLspWIU6Bw6Xz8xmULPRXfXauHx
/64o3UfkQWVNlzCW65yVhlATZSughWtnlw6NAjOaTDBATLOtbnnHDMldtrbptkzr
110mCt7A3pOaVt4/BGWH6LlfbxVmWPsoamMR3iRoN9g+vSvc53knzpeXuJOPZeH7
j6P9qSqTf5d4SCI6QFicDJoa3GX5wvDvIE/4QzMniUGP8d/VGW+ob09+1VgKcX9X
JHF1PPpEFONX9ISnxc2DusMLeRB1Rjw7cR5kpbjMTW/Vw0T5IhOpnKXYAvmLE2+E
pJ/QLwpYlwll1o1zpNM2pAWJ7KSvemP8O22UMWBqLPZYeugUrkC+RbYusQHKNwfj
bkiwPQNZYr0eMKbaaUAQgPc0qocdSN2pmpS5i4mxjETryz1RNSRtBqfRX5IHxnZ3
Z6N74KErZUY52HKYBVe9WQsw7rRF1e9HNZFoBYcq/qWajr15g4ptgulGQQBH7ypJ
UlWJP349cmgnTvS++NxSeZEYaZbqytwCnNgYqco/hEef3oCtHOkTGvvPAD92B4iX
zPkSnTKKGn/rpzDjsDzYWDOvoteEwH8V+7DYPcuvqKJM7ECwev99f+9kmUv/QhkF
52LJ0uOY+t8Fe8V/OA19OXopv7sTVkj5v4eo64uhYt/0KrWCAAlrqCeCgAIdMGbN
ScsIepc0P88iIZnmb19xUIzg6kQQp0N/rraqjfYWpTkP7OoMOjDjPyU3xLFj0hfG
/P9IJNcigtYYefcgNy1ttZ40MXAQIUn72m6w+xVvhTgQx6pP46N6jMR3+HjUHDuo
DNbKfWIXeq+bh5RGOJe9BVzYGPJCp3gY1taTEgLzqFrtFEJZr7iJtUFpf3fEXiBI
HjCBy78hy8+dmj5a3gKxs44VRilNrD7q5C0z+fdxEMOxZxKq8VPkluVy/ysmPHNQ
0e2sPzusTYF1Ew1fu0tOQktTdrVuEv/QRyhSvAJsRlUJpPVM6/WO7wrmjstZ2KGh
lnAWt1GmjyHKfguOslf/pbvNFXvJaPPU6WxK1rh1NXCv+wjv4hFUwgNvud9lHLgN
6WLEpQAQqUSS39W8dHVR/KLBVMpLwBDUovRXJrgWBE2Ht2yd9iaLuEDQ8hvkp2wx
NoBk3CRQXiJ5n2swgyv1O7ghOPv9di5LMlhW4g0r1B/zdUCnK7sBqebNZnY8TCnk
wNPxFH18zwXTOTshLtE1ks++iXWcAREzNTDL9pnMwqT2FiR6I0gPgH1L9t2HNnjP
7E8bBGSj8ES/SNXS6YUT95Mj9LsmY6pXT3YCKH5HoYkeY/bnkS+Ubf2yWUABSzRY
M02xvSUqxnNoitnogyo2af2Fd/JhW+4lrRiDZdXdGq8TSoSh8KZ5TTxFQ7mPtm1m
lh99C47fx8TV8GPYVvZBSMeasAHWkZR2QHDtt4JM9Z67coFj+iayNM+3us7znaOe
OYeo+1AM0yMswhsSMBJzinCNSNWjb1owxiW2YOHLQ/X0ewRQTINfBybdza7MHsxs
UJMgnTZANA9gye3RiD9q/vE75xGLZ3hvYpoUlJPBPp6ql2emCouDkz0JtUl6Psuk
7PqBT0TJag+xtr5VQtWQEJExShdraArS8jfXb3NDFkPEPOav2ON8ZEqPNclzTV9i
NhYq5ERRPsvNlV05zOOu+GQub8GEM3Wb2t30g4Ec+PdI/JBpVuW+7MXukV3/spAI
yTTdCjVD/y/45hPvikbzzvFQ8AQ3bfea16sWOEeDTyFDt70Qcmbta1kR2RQ5PuP6
TgKhHMLWl8JCt83nxE721jOui4K6fv7aj4tHS/YJMT02t1WHXlxHMXgo3mtfdfs3
vy8TATKJ12yHI8VMJCTYMArlbPyM3Fn8B2vc/zO/eVU4GHaoOhQA1hXypPEZ5yKQ
3V6e17NOr5P62gJzA6a2fZPIgR4QK6t9HjBrbe7UmgIwlNq7zBuvxRGufxX6W+ql
J6N9Mvyi1fFFH06om4GjWmDUx3x/VFYmjipWCd8bGrLq0rMhDsGfZf63qIWmmWZQ
QPM5MprAxIfGiJMQZ4O+FMCTkA1NCAFuC1IfQN1u+awBHkq0swkDf6b9AZtwx4Ny
Q8XcSgxq1SgjWFsz5C77jQb96/joIleAKdQoPgThj2L6hdbfjb67RpyuedL7jJZZ
KYG5wkgCtNR73ir/0gVswG0RCnYglNlk1z2ehLlpibppjN3mTbug/VMYw2sFHWvR
um+WKCE1+u1zwz4EdnJAy61vm0xDhoy7sfGh9IQriEE8yEF6K9ApIS2egE6mB3mS
BVZPySZp0FNBam9JPlkC/ebfPVpwiIeXIqF/wt/kLZM2z/Ymb60D48hZOZqOpnLY
o3JrQN7vUS2B+CBakSPuUtTBwulOP/2KaE+tONX3BSFbU8b4ViI2GeoYg8w6oxJs
4LpbQMG0lG9rp3+UMqYyY7HYgnJd3QF18Y5Ew5pTiZ/dWlm0QdepZ1h64a7/mA69
0mCDS7HlAoKf2pGQba7q4fu5eXmDChcbbgCs7ToPdvUlxQM1NunLJLR6Mx819qdC
X0MnircTb1PfXSmWPoiEDIHOGr/oZ4ngjL8FLxKSjozOYe0B/9Aom73bRtHa6VwP
1EfV1s4M9/QWxib9IduMc37bSXQFzm92PsIrcuQSydOtO6t8zM2JNRoGSDHZaa9z
RI6NScgExSKjHlzsJidKBTLAyjR54Hnn1xQpxGYOm+V9CpSpc9P4UT29OVZgSCtG
hSnVo/FP/PQD08Ub5N3r7sP8fUgG77MKllI4RWo/2DtgC8NHabEBbBpU+84HpwBV
aImfg6r6HyYOfOyjwWr0KYy55mEGaLxRz9m9ei+MTGlfo/JS9G5pcWxbUuENbZWH
cczLgn911qqvxU6id85jYi7GZlFnwdxA7SonrUYDgmJXtMF9YKGDZ1ee6y9h0jqL
B9TU+uil4F4bazRxZZumy/6i2WFmAerwvm9ylzPjOyhe3HP9Bbzs54SHlKl21E9v
m9xiNoT1AeeNnWSTf1WiF+sxirVjKKsMGJatrAK6UcGtOh0rJoi3bqkeEwHh8+k8
HkHUoXlW7VxVhKlSI6TXh35FtxxOt3wwRojttRXxkO1iLNo9pkuv4WQDS6L1YAng
6io4xDh4yle00ht7wik7Yo9NRz6LkJyFLADfwkS3pFjLznFupp/1Xg2xDpz/3PyO
nafoQJl8/Xcnc6msu8VGNH9mrbFj1vFW9jAFPFMuhBU67SYL1kcY2ZE7no7jW7IC
qp9Gh8SG77WHksGbsQVtOPw6fccz7UozHOSmwSaO0yrtOjIZKQJZLEdFMkMJvAkO
xa0I9ByLqhbuG71T6lFHws3KsPfMBIHY4Qoac70mcshBUCKnHwNbJidwC+qSE1xV
X64QswkBplGrXo+MZ7kNV80jR4yXFU73yjy1A+DhQgr59olEuM/1XzQwvsRiJcJC
PukoB3Rwz3+NO4K6pr29pPxAhujq7p8voBzOvZ75LO+JGPaDiriFdE4UzzWSLdE+
zKvnIoyJRDrOv6c6gBsnodX5TyojLOgX2ReOxWZ5FPP+eV8E9NoU57i7U7NWyrbu
ihH7pRBOKSi6O7osx0t2W/Sglq4ddX94+XC36yh3lyK/ULpsoFVA3MJ35U9/yoGc
ucuQ6tXldNhBDKpvuWAvNlIiZjcj50+RTGOnMsYEtEohijmDbxkmyJrUfwOj6XAp
6qh1EEeTcwkWtJQLghg7Ml+UenAUMfsGlQjVJN3OZIKQaIURrvA9LW0/0Iv+WaLC
kHGpr0SabgaQkm0CYyeqZ3w5Wpu3a64SpunppujqYMzJhsVmS5IRLHUB5G5Y+3U9
w7Eehpzq96Ib+FRIY3c8pv9S+mRcDnX7R1aU3suctX0K6oRpEGJPEeDHPU4N9eKj
MEapGNcEKRZr8Nrjutzcgjfqu33eZo8pNbs6Cfwf06mgQO1tOqOo6+Ca9yceXodF
Q50PsPuk4Z4EfMXqfqZeo36Aii4SydU1yuiADENTNS4YHiK9V2CpBz7OqI0tkEZy
CCnWJLkRyqP9+qZM3TyDtaHeX6odyEI4HukLbe0apMiIFZ3Y3RF7fHL1VpAhEKZD
/quPKsGNpskSSDkIslyhGQqYhZZ+nJjOrU9TgbMFoxBrnCO5eufnIvR0xX3N2AWQ
NA8h1hPYkvGB8lv8s7NTJURFPcaOXB0RaWU53cP9FczCuyeESj+L9R1w+FiyeMRJ
94RExBjgQ1AwSM3jUnSJx1vyE3a+HvqyFcrfQDMvPb1h4gP2HsSoz3m8eRre7Wdp
iI6+BfT0e31HZ6JwxptYMdBmkGUQKtb4sP+3jvX9l/IpQhUYu+v7o3zTV8MpcA94
zsxJyphbXPmW0eu+J2v+8CRcv/fAC/mtQva4vyYs2BjQ2nZgn6z1KojuTiTx9BTq
9s3NGvISQbZ623o4T09gaBFuCdYpnfWrXd8A+Ug/FoCCVDY66nk7yE/T/BFDLvtD
DtHL96fdQMo1sa7Y9lDsdLFrnPKB2zvdCMTfAyK4W72pHflFzuwXaKO0B0G1nVXE
aF38TYN+LGc6ir8LvB5EkPMVu/VjWjzPrhdNndGyt5WJMnQFXSma0Zwh5sB2j9B/
0bIgmGprMQt5jQ4DbA2uZfr2eEDI8wi4ogfRXPIqSMknuGuk6oddDlbetAR/vDGu
9PHQyra9FSV1RXzt9e/A7crE3azT9p4CDSSxSY0PHtqX9A7kd1nXQx8tU+I2/MlK
fY0oCxbmfoUoOJ1VkzcurznVwK4pReWfouw8wC0nYW7skWMii0FF21R3GGlPZJ9H
n0Pu9gy3H4D3W/eKb4CTo6ltC6NfbKccSDZg+dA/tpFcDCJ50/Lny5rObueiz1O/
67q1JDYvaGME2T/EyNwFD/n7C6uYgO55YC6Ty6s8vMdjzRYdcv3u0+KbmILpSiKO
PiQfm3OAPFfXu3NR9SdSigH6sONwSVHbMm+ada82ayx9+6urPt+AkkDWAWsRwape
1QF4nXWKucBTWJy530DZSQRXwOGi+OiyhOz2Chse18CdF8tPZuwpodeXcfHssLqZ
sQcSstEPWLeeU6h0qB910+JUFG/90Y5XSZuadavuzTqT1l1+aO0w21zB/kGjfrE6
i+P2p5MraBK7mQ5MHt63L1o1nDkzYLfvxkZ6bksZhtH3ULMoV1Ltcib87QaMwQHQ
aF8DS3mVVZXA40bppdUnDjw/jMAqjMhDXl0E5xBoTugc0ig4BHst/XdxoHhMys+C
NEMugQqGh8nTk//aOYQl612e3RF7eW9yCeNEf+ghj02OPgy3mxxB1XRPRkK7egN8
Sa0O57wBlY6nBMnh8+Z81NZV2DRnkbxrywmbVd4I4A/DwYsMI4pPFkYOSeGZZ5+H
BKoWJPzdIDblD8MNGFTyDJPUhzA1V4YSdtx8FeQicoMyq0osAG3aZLxwbsVVTWKr
upt6dWY75HtU1YnVWaUQuhWH3WBiLenbWO6FQGtaN5yKjDfL6IsA8BWdvgWK7Agx
9uU8KanPzMDKR8Wj6Orc+jsZ6L9k8nDppiygKeNLO5ZOn/zwtHdJGyb4t9PrMmSD
eIDcpSu+x5uDlkRlPpQlTfr9RnhDMV4luxPL+JN7hF8JfrOgQ1nadIhqapA2kfcS
jr0qIAA0uvEMRH4C60kXWYAVxKgXmfuJ3XwB1V6zU0ABWqJPQfc7KdOPuG3RmdqM
PqiMfsEVlGnRc9g8gwtVOM9OAKucUQ68YcT/FwEur1PGticqBhFxfxf+mPAJ6Jq3
H6yV/8/vPGkrqsT+B+ffDDtAOHl3mh+w/eQ5twXHkSPf54IXhbKAhVhZ5TzFYqRp
Nr7qQTz2m5h2ypspIHh/bt6dQzCRO8GBTDtBWA7eJM/3JvP5YASm0+aiZa+gGWnv
eYRi8AXe3gUIGiKcK9gtb7TE4tE7kzgemZxa4h5Oydl53Q0zX3jnv1EjEINiML6F
OgWHRswVwOvUgbpaUbK+T8ibQ6lOq26B2j+Jyf357AdEqSC0JI9c2IL3B670Lo/y
nsotOmRSJse8GLvolD4adypG5Ot7XrQc8FSez3QAIFK1G5XNiSXQQzrPivPCC8iY
iM37xUWmIEb+rsK6/2vZUW541ZrCUlmE/nLvVRSX9Pi9fiaAt8Wlq0PPrZ5e7I1M
x80oecabXq9CEGQ2VjPJa2FLo32Cl6JkRbOWC1O3/K7d0yPVibz4CKCFCIsCufIU
JYqErJtCQbOca5m+NCtSjCt2by0sal/BomLVbsPwJhThAFcLiQ8CD1duFXR+JVVT
sAYloo9FJDSmZ+7jMC4McFiceFTOyAiWfptLnAOkscnbR1L6WqKDi54zYG1o9QoP
EMEf3eIM+fCiP2q2DZnGQognEZPeNoAu+6lpChUkuURcKRjJVMWdHdaaxBplXA6s
oDDTogdIlnX1hs9exe1bddVc6p2LWoAeyrlWQd45QEKX3ZKoJi1TNT0SNCyo1a2t
yGDGZykgwQxvnnRP0Vb0hMYjW6g+a+7AyJyqtIEUDLhHqO2Cp5pkwg1FhHEIuTAM
FkIquqRc7RVbXyBPBlqYEdCrKbw22K/TN7wnQqUtTVy/aDDtBGBukxpMvnxWZO64
ZttIfyAZrwONFfe87drtljGnfCbjGjWtu2cLTJByXtchLHtVUxTbok8LgYnxPcLz
LepUNZimbpmJWJO8ZfpuCh5YH+q8agEp1dHsHPcZoglbV6+Wv+uQwwSCaFMNAr7u
a8BKnip/xBB6IP62pWTtnidQ2cl087STv043qDvkI7GRx7fMs9FjsR5yScKR5P2S
35t8Qis/QjCU77Tyj6MlRo0UxC07Zj+Lfr8z+L9yBrHBtA0G61mYYdO7cQdN0+PO
Ch9b6KfF6WlfA30yodUz/2vdVcxTqUDQBc4Mgm8RXajpIDV1xAw5vxQI3Z340dqy
/pBz/zMIp6T01fHZvaUQ+D+tCiAdX39K5Z7rmvF+SaOOMUmkPe2mpaz49V11mBFd
fmRR5shkret8rHMOY9gXI3m0nW1Frl0s6xEfmBbTK96DIeMNRxo90Ra19HlrMIyP
eoW1DW+547AI8ZUOMBfAz6ENp7jUm+hmg89kFhF/rB3nKxqcmFkVIOAj8lehRL4x
qsXBPwHiGhyQsgz5+JuvbZZrSYSJAGdjBE5/RYExpjwsKDz2Rz2Qlh8xwGlVHupX
cBGFA5E5BX6APVqEronNFY2OOwSeicgi11E5WfF+yD2gJIvzmDHybJzK+XzhG41F
v5lluCKUO3f70ECL2U9uAI7McPRP2t0rE18xur7133FVJo5yh9ZJeKhfc+NblYrr
KY+Xz7QfUZrAgyc/GdXMOHe+TyATT6d3HfaxnXgiJsTBcCoNfcEAr3ULbaQFI03l
Y3i2U3653orsGh/+FC/GXl83uQuHBkow0kZmNgzQ5eBkcE+QEuQsLMplehhtzhCn
5py/W/TYt8JjeV2ahYwkwgF43ZgnjgzH236EkBasAGER0M2XwV0IocU3ikzfiB5F
VEHHUX0UyZFvekMV09VGubcmaT1rWvfYTU9HMscIddPgOjL/0OpAIB5fBlx6k1F9
pght0mdUrUCJ7ihwvq7PUhNMTZ6fBjItEZxKwCLtXiXtNAjYB61yMKspfjeNAPPV
GqidBpNt4/dGiuAghx2DWQxhg1Zwtvl6TfKbPXixd99p/w0ipTWqrvqhwxaHiHHj
OFp9tzn7grFGMR3uRaI3YtvbQCLCMK9mTicd4O29oUW8RY4aCRh71uGiZBwZ5wH3
DGuOIUtmlj3d2m/CmT+4UBuz06yS7Etx3ucFL2h4UH8SGBAswG6l2hoafi5dzecg
x3/Mc3R+M7+hkKkws8fMO0BSxwhQ2vtd+qkDBlo2TXqpC+F9MSu7oFwZCzeSlwBb
svlOm8Q2v+gyfDawUILACER86PrPNwBsaPZghCv70yNq+Lc9JdQFCC9ylWSqc+X5
GvW9G/AzR1UdWFIY1h70RHqnOXxpzWIZU0gAzV9+MFSNa177MozVmDHaWlgTqxGY
tAHMWq6rCkEQGki9MYpz8M+C0b0XO6eDvRJ09MaBHK6NSI9FazJwyYjo2OW6Sf9a
t5QUDxFFpw7pYqJA1jARuK81Qr8cK9P5RpFW5WyDEG+Li/UFIqtC+zlA3ooA019N
UOJv+lWom/hJb+XtNpYZjVhbfIGX6RBggHDQ6VfZkd5luCXND8fveE8B/76Yao9i
+aeGkvfe4dqf2tPQDNr+sqEfcUl5yUU8a1GBZo7nY63gth7r9H5LKRMNBUC84Ib3
9eQfcPTBJZ5mVDUBm04A6nbyjQalZbEiE2BNve97o3yk+nOuOR9EY0bAt9NSeYUj
xSq9fj+O+h252Y6BIVag9LEahzCUZa3LsapLhDdUhANdxpezZLsQn/obq+EFVEBH
Bnca1jodB0iv2X5rRpc9Q7MTe3AR2KWnhh5NnlzhI9pCOumh2a/1tlw31iBTHGWD
0CLeup9sH78AJpCsynggkJNf9kys1YvP0P7f4VPSDAvkAvZ4W8XE5YiPT40Tl3fy
K5d9lkijqh2Dm6okMjWkr0ydtpAIkXg6kNmJbE5JCoES/ks1MJaDKZS9bshXtaLY
MF0y0UPwV/6zXTUMGUM31RgkB7gHkPtH/g52/7VJy0vmTSBaDfFsWX+Ux2ssyZds
cXnfW/nxg0GF9n5YcqYVyRjte6ufWlwRddWgA3QbPlzdOVooQ+FuOG6N0EKCwgxU
UR3uSnDc+wvy3OjBE0Zr1u0ZzThrhGfJiu6k2RKrke5nzuSoc2K5WXZC7bhyeWqD
1BWc9QOSOiBK/ZN44uBkT0543AzQuoECcph5TLpr0JD9+n0QtCvQrOUWNhZrCl9p
xr2vhh096L1z25MQ8mVhuTuHUh/+h4gsWaGXamrEWli5yLC/PgqWJUNL6YB7C/+z
6w62kQvhvyqPlMJfA3R9gxKKj7pBAPUDR6mTq5p2L1p/8ZDZ9W+G7boYvn01jZZs
JDei3dcvP+AZYkE+b48vsekkKx+soNjQVzoUp+/CxHN3Q2JY2Ks3fBI5D2a1zwvf
bqAKYJBulYoOerNagC6Y5Z/Dghrf1TXGH5J8UU0Pkk89tXvqlXl4h6NDJYs+Uz57
v439NFYfHLCcouwfrSAzhJPZXdjrQF8YHXt6JCzZLFHGR+WihtRbdcIhjz+pZuZu
vQA0G7Rx7qvyf/Tx9Tzj/pY/KNxrNubJkn/zS4j/RbX8eu8sLJiF3uxIGUmTkFd/
VP6GEYf1kbVmOSgTY0h6YcZci7KRrYozJtpCkj2Ka/dPAZCiDYtfPqDoyQqq4x0B
fdkfWHdpcRsTYBNI3B5TKlDBqcvlC+noQb8kVKB735I+lfNY6ziUxVE6NBpJ9HZN
TzXoLO741cwen0ep9xsV3X5Kx37VJ8bz1fpwujnrCh9rhtMQiIDYQHodgYac44Bj
OsHIC+SjizXzHjFkdasw/u82D+zlY4AFBfcHb54W2mMYlhXUmJdL409h4/9FqX/i
aQ/vEDESaS/V1nuLUcG5zzMz9YqAQx/lNArSyeoPdB0YXWfLQjFcUW3K3nDiCkUR
pj+ZSU3pHejReRHgNxQRtK2JC/eNqc0zhxZa4UYpsezUh1CA5q54TEfYzh1o/3fE
e3dvF1JqIFuLLXkk8F41tMVYKWH2GslBnOS185pxZu5YjmqRYdhuMLwx8dwMJ2WC
kWbPArZPECHvSdIPX/Ol62Sixy7Vd3bUNnRfHKEvjJC9PovXAYJAUzG6CQZAjpRp
AQBX1adYixo517YCP4RWckCq+cyqCpQqkPe2uIA+P3/mpMu3HWs9gEMTvamtseD7
BOWmlqdrQ9Io+nQ4Mgh69d0aEXyNeFP/GdZ28OvH+f7hPaJDu7rvp6nGRM31n5Za
H6cBL1BzSPgDwPeAGKXMqNDYMgTxV0KGxEKUpdOEt/DuMcm0HggRnBvAJ8PBQiiT
zvw8/GqIESHq8QGYMrinrayGcY646DKy85R8QSP2TDBZBtEkmOclo919DVZ1xzXc
SxdtJg94XdLhSr/KHAO/ZjuaPx73nIw7iqaj17LVHXbIOYMX7nEAno5dXjQ29SY3
uZDOj3OD+EmpCOZMbLD/LaQpooSlmmeTK+hfmLcxXB8whmS6YPwhdvnd15Dg7WMi
62RdR1pyJu8/By2SAdAvyguJ6Xkq7L9Do5R6PXCPvu/FPcZu1f/bAuRwuDxb5fvJ
RqIYbnwTkEIy3893hJCOQkXcLvu3WcU8gUf2YsHIapYOKiCpOTRozgIz7UZfPbuZ
9r5t05a0mtZRD8lGLLt9reizaGGR8ZN7RZFmcl60ttC0FLBriJnpFDbTFM8Bg+m4
tH49txd1QikSkcWz+MQIQtBhwUMVf49pGHRhFKBWV6m51khSJwy4tGLFjNmBkL0k
xiiVRB3abxXb5wtq8tA0PlB5m76Y+ZKuOI4RoeSdAtM9Z3zXpX2Swqx4AQ2w6j7h
h1HC2Iy9mNRXblhaFYY35J05s6/0wA792d+asqQvhyjGTel2EbKxAMSkf+mEL4ik
7ITFtFc9bciTJoOT75JsKof2ztsrsmDrO1TzUKtn+9GomKpjuJdaa8QhAMbyiEtj
JO3aei/vvX0LjiqXpC/tdSVYoVwdbr3jEf34QoZY3BGvEHO31ATOBv9DeN0K51oB
fLruFGVkAcND9Mc+edq7MW6ZfjkFL4ftHr1FQrwoED196TZOyp/73u+fe6VUf3lw
dXNXf7pdTTP+zxdO1D9BlRFECtyESYLmQe+ySuqdNU2YMpSvaOGVDR3yH02yB2KT
sxPGABIjXt9F47pHhYsxP6VBjRDVC6oAl3BH/AnQgBLIh78LJdZ8lhXdiQJFs01h
KFSfD1Nsup6dRVmw6LoKy8vEytwJnVwjYZP1P2z4Q96kBY605d7yoJoQLpP615rQ
7V+y4XltiOLCq0GYp34kdzZ/gDuPYVWItZmdGzmr1OBGBrQDmkO2sPyLPjgCydIL
I1G7LPOetTgyeLs8/RyYwOjJne2467c9MqEyzZgPevb7F5THiO3dicUVjl3UUs2m
aXbYRT3cZG8Evi5XlBMh7+9BCKm3Dk3hBd9biSIP/C9TrBgHUxK8lv1rJGKxyzBu
kIzPyTrCQbBBW2CtZUQTDY/xUZHnDlz79Exe+8AO8FsAYM6DPxzBRw/95wQwwhiQ
UI4cf8UMTX1svazPN1BzbnBmEOuUjUq9Cmwd7GuNeZs1odJKF13pI74swsGbqt+w
enxvgR7SysBJhogn6XHqNkRUyEHptw4ivVMzvAvEDgqKHFJg77KhuedFM9Ps9Wl3
A0Q/Ch7tjNPByPQ3fTfHRE3ll4/urckG5JTXjtOBHZ/GeI+23Pp4hKpzdy/64xrY
4szSWOuVMnkINh8he6Gy2L2VAsY1xJoCsdUlqW1Hy3YkPUI5GyW07NNWMv6P8Iqc
Eaws+bAwiCyNO4V1+aLSad9GsP04kHY4xEoM+j6OXmVGhVwaV6sUbcyl7iQeOi/e
RBDK0Ookaf6tnEQISG9Vq9tcB4eypZj90/F9DOsXJxvEU4W4/x/z0YKhLzKYsQaN
tyi6ute2ZpsXLgQd82diUnKM4EvCxaFsuDbAdh6RXPlvAXcWAgI1YYYPPTNHdJj1
MUTlgDz9+ePgoDYLYqMN0l8w0JcNPuua2EFQp5Xrp36Id2w4xuQ2dxytxjO1Y/EA
zZK+R72Ma0Kx2pYDF4M2lCBLD6IpOaCtJS8OzbRnxUKznleDu8bmrSGmuLIT5dqV
UE4bLMNhWU6jpd15oeL5A9uNcPUsr/WT6fhD7GHtfAoNJY80bARQZRn/QyzvbJ34
0OP/y+27t2gGe5y4R2N2kLlgAuFPCA/abOOO7dRznzNlyHbPWZMGApcenAWJCxwf
tTIwAHaDpJd1Y9/7agtginDBErizCt6OmyPHb3ZcBofqpONBRne+bNBH38c8V6EF
EoeQfQRBKWk453BgGupxMCpJMUoCgO0F2FRT9QuWrU0DN3Aj8h6cn4vPabXUon+a
E/0+6yKboMy7t4wl8TyZDDj8yhok3FJcyoUbabbbKJZibV/7HCq1J6FmNZhWNI2z
vsTDjEBVRwWmjHiv7m8aSzHDmU7PPbCWuBOmftocCfXOcj/5qVDFa8J8UvA9932W
W0tgfatF2zFp2QBneXPzQ7Y3zNpjF9ZP1v3oE1Iirbo14Caq7lVzfut2+qOMKheN
1EB5eGsGJWWht7oyab8Z13PBDB2qp3+hwSv2ICNclGudIbxP9S2UYzWh+MJCGVF4
CGj1lT7PuhOAR0opYl+P5PwlnNDiLVgouZHoaJNCtZCT5OP4dSFtx6MdobP1apVh
25rkAB9PzzjlwELce7SuXSqen0LhS4ZnUqjmt0Lo1UmYKT3RbXWtQmNDv0ZZ1u4f
X5EXTqqe0pa8h+0pxtln0cEmaWHxaDRg5CpPQb50+9sfydhoY3KeCkhli0klOiho
Yqcy+lrUy/CxHNUIeAIjaNUO7Wrz2TwF9LsxBBsxsFgb2L55g1KrExIZi0FL478Y
Hmrm1G5N7ZshsFVcsNcb1BfCOk/sjuESCiXPPs427ZAG2a+f1sOlWIg9jDkdR2BZ
2Ol01OBtnv5YSstVpQ+fgMXGXmMeyufILoBtxyLKTRtJeH6TgI4rH/us7sM5UA2X
pv4lB19NxR1hD5rCcRyn1Pm4CcHnZevzaiANS3tuSSEfDUnRI7EaSPEFOYrYypfq
bH0uqjzMYiHB9xq3D8suzW6pL3iG4nvE6ASE9oJLhTvJsfgrVNmBUF3TCVvJ7pxI
f4RUS+5fQCgZGDWlUl13fJgvyIqlVCUDUta4MeuIe/lHqXpGNrr9oIE7JQZ4JTHO
KNDXyHDqM3tUAdaEYGhjLi7VqYLQN77V6MZ9hUXiud3e2rZ8Jc0qjlHyM+sCmbvh
qaclsAxIQT8j0u68ufHp8KEvJTngSTTgmFrYa3bIwWwg8aNdbiKKsCsUOJk+i4p2
joJsiLnVk+cQfNsUYWUPrXcGpTelnJK269j7Hph5860KniCmqoh/39OoD3T/XSCj
seAa6WYz76GGeS13za4iy7aDwUZOBxiZO9kY3g8ae8CJ1ibn4qcCaxMVDeT77R4j
DH7knxErgJxoVipOuU2hUE/GQbQK3t6scBdgaChiEmYs2A7hb8OaUV0PTyf21VMN
WFI0YS4zx5njfN9HmqPPWLT0wiK+yU1wQYj4G1prlFKmsvbkKcL7H/pvkkKSRvP+
L1gWDq9/OcLy+FYM6ZTi3dTPKlSBdbEcnTftd7YN+BUOTxKP9A2AROOUKnE4V1xW
qj9zWBUGjrHp+cHEs1fBi/jcMeUPZIerxGwpfIzfOQfAiEwlFiuZTPcsE6sdP1V5
gSlkyFcz5cPf/mVJoW8GES/BHJIUcWKc9RVdHogf3iPIRDXG9wQVUE+z1lokwZJr
TfGJWJ/OKlGiXvyLinaSuXjtwwDRwPLV9XHjdcKTD8iIiPoW/RZF297a5htlySUs
S/ksTypshYcNh3pt+6yf3/8Ogkrkcs6gWCR45ElyNp67mxs6jWbLPuZy33iaDnj8
cBshllfA0ZM0atS/YJKR+DHKQuvMQRBsHCXS2HJeWwb0fovMaWsOkc3MMjRcanq6
biWdy8/9Vpb+fvRO9WSu4RQ1LyYtt1fgcf1YNxPcaazku4iO9l7VJwEiNind4bmn
6aqsI/A6dY85SRsv5ibuUW/gD2Ty/PjkrFd32ADK3SlhvpzRZlkpqs4NBNfKM29h
8/EDmK5XxTz8iOt93ObE9oBIZrl5foM1+YiQfBVPlEV2VZvlHGHJuYyZWHoAfc29
39UOxmat1CN8E7acFbKvgWF+o2ar9HghTmvpBCbHbYelCFIn/02mOMAj3dmDxw8o
/7FyJwpiv1pXhYyx6iH3ChcFOuxLrflYkzKXfy/mtH4Yz9tHzUcsbyOP9fdee7kJ
4/AzCRvNa4t3v2zIoY1/Yzpmd7cqRPc9w7VQyn9yACd4O+1GS4FPwMncHPgNF8Ec
6qYIczdNdF9omZ79RCbcgfAS0FCN+oEeBuuvMFjmMsRVfdzGnRdQpyHN7m5xszpb
Nn3hi71AWE1SDJiGH5bOQtQEhw0IcNWw/77H+lY3HDIAn0fh3l8Iynmr4SPg/77E
KKn/06lkkQJSnXl0UiHYRbencBEDD6/KcLwrKyQTZovBKtxkH1qDKdztJ0LoTETq
SeRNJGjP5ZFHwdWil0VSOyL9akL9frbYQkbUKSXc+wzrYuzBZxNSJa5R+BdBC8QP
ZIqrhzrNkAyS1n5qsJXg0D02i8dEcIwchRTlFqzrIv1ae0Xf9R5NLmm320mxehFV
6jSxxZYmyRv/Oi4lIscr4JP4kcbTtwJokDBwJt9BVC4vhAALXRXz74xLYuBj7wv1
X98sp2I45txMvQk9DaV6g7l1rSxEi3QrMW6Axmg0oU+F0/A0FLeZTfv3mkanpLPW
+brejk5zeFRMTwNavm0fLzimZgmnTAvLt7YcIjwRoKasg8XievPJQHU9IJGA7pUt
QUZwMguYJGetvSEM78J4P3QOscRfThi7mSNVTWTmKje+/Fh/Af86WQiHuLZYsZ5U
myYlt7ATw6m5c+YZWshveOTWACJYkajVQSYBLaYrBQdAExgSmFae3a0EYY/OP2gH
SVaEUAbHlEWu5ywy58wiXd86mt2NTjMsqWujcNh6H+rcSGEER2clBAeguWUaC4sI
9NCNno3WmiC+0zAUfbeJsW49jgl0+jbl4K2MKWv0DzjsohW0B53EVunost7yLXSc
WsQLtwHNttuSbSG78STQFh09NlT3qi+p5xP0o+JZ8RgG/hk0rFvGDoWoC85QG3nR
pE+WhFPKS0Kk8uFxEIfzrCdxTt5/zJWWqV9Gtk34izxcYI04mCZAFkODy+5pBqVR
7mV/X3X0kctFEYEFbSS4TzqEeftyhFfLtsyGx/hzHWQQE+QwlKGNW+zxI6ibDwxt
HZ4Gt+jQ7rkv1pPn6D0MSHppYe37Dc1nxkfSYgYRSWowLb/Ew+mDIQBXCWEnLFXA
pIaa5NF+MrJdXFnniFaMYjd5UmFwB+jpY0vd9kBfS2U6EWkrO1tPKqm/mvIJiPCk
ZxV6SFWyQbRGtzbkNWQBswVZxKHA0c7H4zFAlk1QFGCG6+3yLNRRMRd9QoklsxlP
h8lSHOKTqhWguuYeLvu5bjkJXBVCjNew2QEdKvRr2zFatDWKQw/VvwbiIyJdVEsP
r4m0aeOQsfwoJxlzJLKui0K54L7ytkRsj2mAadVoUy8UXpGXVdWEy6XvD+qW63fg
bdnqIxJB9yVWEV+liAMz8i1SsayeDZV10hM9K9hpS321Awtk8SXLWsO2NuydN+Cf
oK2iE90Hr2tMBFsWAR1s4BFIPYAbdEQYK8fwCB7sTp4TlEopZ9jUPZW46AdLjWM5
ltbhkKovowpXjqgCad5oraU3S7v9IWzGpfbh4hrC7hyzpJcXL76ng8Kl41O5q3yI
+L8qKYeXrP0Z/LukLlmPl42SKhli2WsDeiUxzs7JoKCbOcoOClWP1oJfrDSvj3yM
Z5kLcFT03f3UDJG8vR1U//9pqhZAiFbtjYNFPElhxnSoNGpjsTYu5Fd4OQKzfIhr
AB5Cfych6/ZDuZdQ5IT8K9iuv33BxU02ajf1PXlW00wTphN8DPhuATrZ+oSbiOAD
urEjOkRMp1ZjvqFOnaNeInVeUJ4OnQogbt8L3ptYX3tpgT1BcE7nzcBs9IVXZPtS
30O/BRvnJ5/7jvUl9gDu5WvtcDK8Avk9OMxQEYGTNLygOILO/EzWQjFI7oLXyq8x
wDORm0BJFmXQZB3YllVXICT11oaALES3IP9rJQCuVNNxHAfDvNMODjrN8hLx4jqv
L5BkZKRWoqL5VNumHZq+hm9jH5L6w4CMhj1VhHTTjPmxBixQFpOvnH7pK9vtGIM4
7Tew1Z1tdUujBPaWU3e51Q0OjyQr7SIXlFhLyKEBE6XMvZyeJpUFs5zDusRad96Y
o/8FvsRWevMov1umM5MyefaHVXm4+T8pK/42GpOhsdI1HfqbCp63n195hd6pJDlt
jPZwwlwGeHgQBC4J04nKGyNBPyJU6hUxhW+RB7luOMetN9cpOSgFRYFkMs6IeE3Z
qp9C/AN1IrIrK98mNGHYPxTU+nyslk+h3BAmR+rx10gTSKFW2LqbS6cxxF9GYjkv
h1FRLOJywFrIVh/7mCR8SxYue8JliyTOkfxh8zmvTUXMBQxCzmZvvdf8srzVKlny
yjM3+/2Cswg6JkHeaUPUh37Xg8Q9S5wzR+poqCzra3nwu/TrnMLiksU0B7oF64Nc
D2fblP8bno+wPSgXUJngc3qeLqLp6Uia5pQ0YSMmOFlolvaJJtXx1F4wntSzzxzu
FFR/eQxdCT+O0oyNvsgTfLIiks3nxJRtti2aRSfjbWle4wElGwTy/srIKIsc8qPK
HlxWvSN8e72lpvic2rXk6KdS1ZpTBcV1OP0NCHe+w/eRIUV683jVT8DmX/AOMH67
8Z0U77sQoMnAAN+s/rzEs6jWP7MPOtSJm3tVS2Bx2+1FJ5zsJhVXkw8F2nE4YzAS
G9hRkFXFNkk+YrPld89ZotyuSAKezBdv64LoAPgxi8B4JnTvz8wTzJlnfvKfxGN9
AX2lP73j8uyyOC9GijXld0kA4TubRwEeNvKQTD9Sf4aBXz3x3PTdgmtdrkfu+/Gi
N50rwVH/pv5UzymltG2DIIGEWNI6DRHmzrjzNP2Y6m8mE9DlAOJ+TNm7sjXWTpzD
LjZBB+78ef/NSSv0ksOrlWqABAjuiX+WYsT3qDFEB0OQN8UFOmZiYckBZhu9t4Xx
aR3Djb2DKOcWL+VUyilmxKrHufGiwR4lpZfB9NEPhukD680anFYOlPr/SbmPektc
C/T8DeJw/+n1AP+HRBONch6DITkDr+QhxIS654/81mGFBcH9rXuUgOOmIjgpNzjV
n0Tww/5caM150nu5HRZHrVLNEk+hiJ2OHzuE/ZwBgT9XQs538tdKF4rtzJQ+Cd7S
IwEefERvYLxbNSHG6P+TZco6cRmQ1OOcGAzGtoYrRb0O4GLD+d0+yU5pIBmPsmRe
gDYe/uRTTwf1eW6ZgDM93nNYEMPp8g+ApEb92j5AGCnwlK//dPKFQ+VJKOZBVEIi
B/QHSRwGnChYepJ7OrcNtjf239/y0wPRVU6VNhlIgSsQ84He5kxX/spiMReAngyx
yfvlfemhqcSflyESUiC68HhlyieoK40v9k6/8SKKDcEHa/FRoJ0yuf2qiODqDQac
X1rnFakqc0bpbzx66ePqv4ruHIFzEBBzKtE89/B+HwiFSVZ4QCnOVAG5rJkXv3OJ
x+RtBuayNVWeBbFSYnbzRq59bGFzsDvOYTAgi+emYD+V8xKvZSN67etgbzgwiMo0
3kq3+CcEKeR0oTY8LyBARmZmOp+V3pZRxP6uWzQQqMUslBbgkdfOmFdA+Oi0H01t
MAXZmqQtD/JhO9datx0UjA2on+VffFMFcVQI0OYxf8MPmZ0Ia6ZrFo4jvlvowfgI
kVJ1KHk4YNIZDKmzJbcwayMt4smtuGC+BVELROQlUzs6iwolnH67xW5cToRuIV7R
jibVK0VkXk07F11GPGf6dRKaR6T3NuFZFGLjVSC5jQi/EoR5UdwSdC/4Y4Ca6haj
efUleNdjzmIB2NmJJcvhZpS7hpb1+GkZXg395wMlJKk739GqOTZL5fF9SbbhwyQ7
hhDxy5wSSsuZvZa3b4Oq2gOLxwYInsWHLzdxErRxlrd7GEqo4HFLi9/pTJovFn7h
3B31rb6qPCoybhhDmguj2di/JICZYxQD8DZYJM6hiQi07iOA5lxzbRHfcT0yEd1u
0+Y4yaIrvBzh4F17YFtYGpjtuOaq3Gk6QIV+uiX+Fi5JrvPchKZkrzicQDnlz5Fe
UwVAYNvhfrR8MagV3Z1F5WpTqiI+DVaJjQ5pFDnP5PhCEfZun7edqZ8dBUfwjFz9
Lcol0LINchjoJvOLWWJdOsNBM5NmkYzDV82w32l/XAMKSDB41DmoOeBS6ODJTm/Y
wCOe3+PHgbDP/DkZYoPZbaqows4iKfrYK5GeDPsEKSM+6rQKUCdrJBH3PPikyzYC
EADq33te3QsTENpJsU1kU1xnOB4618Ihc5a48PqEYp+EQSXUEtiV/TGcWE6wZfVL
f5X50dB2RoQXqKxedx9LzE0kIQ25MyVGUtO2urux+z+Xb3cfhqC3YyjFRqCqTFlA
tmpFLTlog1eB48/SDOu1g+cnanHlTbavk4xBKbE6owvGkJvAAJKXObNEWxPj1fVN
VPrktqx5KqSm5B6thiaQMLEHSVB/2W3a8LbHxQUqIr/P+6kdpSmqPgdFgxha9L2Z
BVMJ3bjGb9uj9urRwwGRkz6cTv1nB3kd18rRRUJDttc4Pej3PMhlbaaxg+D9IrJl
9o+b9rSiwzWVT3L3t8nkJxynSpRTpwl1UPvr41FZ1/ukulxiyMqIl8DHRwYvs0ck
cyK9PRaWUtCaYBwoPgwa4hMXU/tFHyr/mvIUrFgRC5O3bbxjvxo0VTFnh0sH14J0
7XTolF0WEM/Xbck5jLUo7ugvodzCG8ZQU/eSat9QA50x3GdfDSTNcUH4x48CK7R2
R5LINpRQYwvI6c6tqWdXgtvhoZg48AcuM6JXzwf49DOk6K2Je7+62+FtbONdPDkK
qh8LjSTdiDs853b7QLQccRd2UBr3N+mn/Ht17DC8KyADY5LLER8MO+Be4Eq5sc4v
9t9njHcc1+jWM/Te5rxOK3DnS1M/jlTY+rOlRnTBURIQiMwuhiY8vKHzW15YA3Y0
QkcAQZbLV0NXTWZ6c+iPNhe6hY9QigLQHw/KdoQnegKoKj30LBqEOVJ+CjI7ajxO
S4KKt0VATCpINBGbmrQkkJI/D3C54ZyFJg6YH1lgRnH0O6JzDfCNkFWcjU1f2z3j
C2WDxsFVdPfuGLq1vK9AoYejvevLeri+9Y8E6KdTbQpuU4QWSTJu9ISe9sdSJ7tT
h7YwXXRCoxikzSBLO6bVl7v74SzZ9zk9uI99w1DpztGpg01Y7lJBS2JyJzRkEwjB
iueIDnjqu/akYmKfYgx51WFFustRaBqvV+YRIFwgO+szHWahDbPnXOI6jVgtfwCQ
yinStXDJiwDsRLGnUdaKcIn3CjsnzVLMb8veVi6VIXgO2zi+L33sAgdpqByE2dzE
L7wS7Yh7pw/S5gRRz2qILRVLKvRY10x7OczpUmVujcI93AzRY4og6BNGSt7zdbNK
/3yRENu6yr0vMCpESiLxlFTFoC/mQ36uglpL5daM+KzE42r1XPpehAHdhnQ+cZj7
yY1LKNmxcVw+imJ1eMcNp4BBk1OszOmTRC1LP82mFE14nCZGTMeBkc0y3/c/Z2yy
lUTLYg+j+bzatFgfqx0xKJSdxhuPH1oySVNZTx7N9D9svm8bPdx37wM793fkZzuz
aAOrwmosWzI5n8NQte3GXLwd8q3GS2NooQWfTGX1+lXaT8v+8wFWzEGmQY9LsgR+
qj/cKKgqOczF2YLmWaJZ/CC3fkVaeZhzgwhUxEmMYuR/UlIsjQtO5t5yLomDmx5S
dNTVXazgY1T4g8gkYLMcP4MX+lR3eoCdMo4xbY2/TwcPJVuPh2OKxOXzIl1rwJ1u
SWkxUQQCrQCs7pjAtJUipfdmt2KIV0DcRpTwiFWfOLpkFJ63dh8XZPEGR7mlVoFH
1i1wITD69N1N2/ySGRg29Xah0MeQMdp8vfLHICw7E8u2GHYdZnnEYwIL2P05ZGgX
C0F8VdNJBhE4tRhsbK9sYJA+ITdSn5yyGAt28krxSpZY8i4Eh8nftSKdav3qRM6Y
y46SNwlvGRXyGhWFvIKHi0YPHcNmwKgKm/fG6MCAU1zd/MEVgidyKvKvdmQyRLPx
tLC8xNDb0IJ471b4SMk5f5/TfzbexYGmCUbMt76FFOxlZVWHtHCPcyWF8m3ahdN4
O7CwrCoN2wiVcAu+XWjiaAuyOs0boayZScn+tQE/W2S6P4hNBWr4DWcYNskiqY6e
hEw43bhVaLlNZck/KsWE7WrPh7TM9JmFE9qAMcfRpqQ5WNMrUUFesaxbsbHi+J9p
C30A3SMfihOKYzIuJiF6p5a3yC/izhuJ0VBccXo7mgeznzgrHebIFNv4TIl2+A4H
bSo/i4vy6gxA9XEb/oYVxU76OEDGNbKseAfwW8UK3E1VrN4P8Ou/ayVFKFC1jlNv
z1S6c+Xg14z4nGJWA/WfiZFKJWElom7QXZ5PWGS61NVKiDJbY+pRKeBFb/xkWM39
vKu3JSfHsJhsJf0w3/KucTJ8CXgH78bbYhyR4IQn3YSb9/E0UD8aVcoWseTIqxb6
B5G6qZaPXmKNs946J+NZ9LJeTVKjBi033YFcwnvJ4yc6bo4mMBTFkZVsqeliTIcU
zGxdFhLqkR5Mv3peLHxMurG2grKtMdBB/vmmsjLSx5wEgMvdaoyrlWkjgijeVFEy
GVn6ckYMSB21aQtKWHa+RNAx7YYkQQFyf9ySVZBMBkP8t1u0419W7V5B/rmDMcQ/
SBpsg9wdhLrNE8y53vYrOf1KT3vRwhki4rFn0d0kzilEkHY/gptWJxsWgmmC7v6c
b3/xT+P9gRap2y/khmqjuEy1/JPVoYq3i16IdpEPlpY4R1l6pJeggVFwfTqAJxGV
RsbQx+UeZnoUH3qfwm8Wz+LVRBiiRfg/DwpWQnV4q8bfg0e/7SzToKb0V9qhYhBJ
5wXMLN4OyDLE4QKFIMgYFHv+JcNypzw10Y0RAdEuIBrK1JLMOWY++sHqGf/jgyxk
V8o0fzAf08Au8ajnC45QXI0jbFKLPode04Ma7jqA46aBCyTckZT7Rl+U1pQPefa/
E+qayshVX8XgwDor5yuOsIlAhmDFSDnq6j0qLQRJO7Q6ZegPhexgapkfFDinB5NV
HCSPSvMOt3gEdqE5XsGRT9zBlv2mf98SBneSCwjbgWthvN2VnzvNKvQFYhTss/P4
SFE8lW/aMb0HTJrSAzOGBlCIx50owbm98/HDiqs4KEXmLJKrCIbgOnCfQo2P/BmQ
+A5GO1ouXPWfHo4xRPxktKdl+pQe6muJc2bm3RXejGmBopyO9LcIo6JKQlxRrYMR
o6pVbeQYEOMg2+bD7zWcN2H3Ub3We++/cX45ik8Ju7zLscbq7tuZkSu6VZh2t0UK
rORKm/Uf0++DM9m7Gw/YhSdGGsM6xV66aqnSM4oGOzKDOPBoNEPFyhQYJMccf7rQ
dW/OhyXiqPaqeO5NbNXJC5zSKSRWus+vMPnBOWOf+P4EFao0lDNp29xT1UCnPzgG
eRL6JgsWHBizamSRFLc5AQ7Wz2DU+3zr9EjudRAs52KZnQCiYpcxQ/8yBPTAR4RH
Pdvu0BLuxMMJ436ObOaeL8DybuB43jkmQxOWDBsTrOeuB2ZfJGE8y7/A/sAWbRX0
2ahzuQqNbt1JsRQRhibTzhl6Ajmok2xjQSAyhV32IDnR45Kg/oRkkoMqm8PN3fG9
AV63KxEZnscA8k+9A1y4cTQLMLv7vZouPugD6C0d2godCQRbXjOpt5E+EC72DgwP
O9OnjYKrMTwEiGTwwSaQKYOxrvTl/tvCRU6t1E1xjNW4ozTycF0aOp0K88q+aCsy
A2reh8xg4OJxp8/6b5GBydpNee6JRSmI3o6qu3ggMya/LiMrKxv9CimpWMFOfDT6
VwlvZseCD30svYPPWEDSpH/qDRHy/6M70Qt1DnivJADzXfg68PeIuKDeXa0/2KOx
PwJpASTEYRxRqSG3KLp1QteH4DxYQKqaqzzUGM5s+5ufpt+gxDMyKBQgo3kRs14A
0u69J9mDtcQcZ5zec1eOSKrZ0zbThDeRXVmYRzOBTcxM3vW96pWkn8R7K+KlNR/q
4dPQbcc8VzZOTdMOyN39mtBWLp77gGPDJ7OIk0D9WaDUZ0X8fS9O+U39pA7pEvvv
wiJY5yAmSz4Gq7whJhStRMbT523mmjv3/J87wkP9slFimUAkzKHjF5NK7fWBhlLf
TsSwYU/mwTNivUwFkBOipYMPwRD6Jh62+JnfAMRDEO6mJ8JH2ab2qtgaAK3islzZ
Q6xUiKcdQf5tcqM1eiUfMwzQMwIEq/Rw91cuJwyHODFVlsG0S4/XIVIfrBASpsu/
ucmRmimMCcTydizoanmNriHunIOO4JIevsep3+DfbbRl8AE3A0k7uQVTPZyR2oPz
SFmyERNlw8nDw4xdZaku4oPMbCDUyBvbAq+NEqMbWjYEEKbB+BTPZ9QqcMT87KFp
Bm2lmJPJEsbxdExQ2h+4axDnI5B/XA9rRpn1ehIcZsWTe+osse/3GXriKO6xUWMQ
I3P/nmb9pFJeb3MjlWc6wiNrVmFs8YxrLMBI/C0a3+GmsErsAOjMOwjjQdjqQvJB
Sdx0KTbWJoY8mSy/BjDi7EpGV38jCwVwQk1cNWRksI2CBzWAkBa2ePoUHwB+vtA0
YpbHCouUUbEZ4933lNo2ZQn5Oqpf8c5UXviRIbGGYTRpO10zwLNqOaJl39Ycbsb3
Ai5JjNPq+loPm8+6U0FlTbY8sUoocVPLZh31wyGiZCdRPZtQGpZfr2HFQN759dZ3
Howdlgotu7MyTpSx6E5I0hj9kPHx47ma+2cJX6uNH9lySdzlatxamZPu0C8AP1KG
IjaTyrvy+piW0QU1z9fjN5aJDM6IsieC9iOc72cPHQ0L42fTRMWLnDH47Oyl/76P
CbbOxg05LwS0pKchNR3innWgj9LzWyH5Q8HckGBj50PXqlmLUr3ZuHmeUzGAqpc1
CRSQAEDaZV5fCuaRuF9e2/K9tW/s8A7+j+8H5w7I+TKY16jo5EVbKS/tNmQyZx9Q
tucTTkB2V+1uvP9cCRRu8HivKPc4VDI7C2vIvgL/kZUyNLpwqC78vlehZzck+ucJ
3daQcYaIVwsqAONj6iDctvoRuqXQYRNqF5ZeM9RHWkbJpvmnEDn9qfv/9LPf5g4G
vJ590toroq6oHUsMJb24VtSc5K9MRFHg2xB/+aW5CPrp3AwfOXsMjyUfbVJZkseq
fkL6rlc+R6Mr3FJearT3TnbiTwrB0C/CLl49E7o4DgRfX+3pRaNY9zKOvg+6oD5+
moLF1LwWWqDLP8ttJ9Qi+YCmFgS7XNI3Ao4ZkJpPW4YEgzNvjdILyphVAiMh00e5
/QcF08G+cwBO0YHoCgHpal6Di9f5BjzocMp8mWk4T784iQ8R8Fx6FtcHpKswfOvs
dkvTYbxDXVwbBQDDPPKeaismWxITkC5LDaY9zaD5nIruvZ4tDMtwuhqwqQ72MHsF
xA/Kj8UkcJ7Uvdpsm+DKpPJl9nbgUfGR7gi+2ggEn1AsbtS+TzrjXususJqkP5/B
GOIXl1maD5btOChs62UnXTjNtNvLx0hkxAVF4ntCfitm/4cJ6CspU6HkX9YwGuDD
pKisnbzJyaPNVKfFFhBNEtdwrPH4TNF23GGYqUpZ6h2zAePGL8USCgfA+Bm1J6Jr
1+yyIijR8JDjE6wUUfGvS2iI3PwXkCtmaeM+mkefP6YeCgZ/j/7UvqrCbFs2SVHQ
x0MlX7qLZpjr2n7YTQQrv1epwdi5UMEnvGGwnznw5ZdlSQwaXOtJms0YTawwe/SE
4eH7zVSRXz8yFMFsy3XBF9JgrTNYWzLoP+L4HCARd3TB++LykLUko4HNZX4uce4a
1CGuIa74t5R8UvEs6W+5k7mRS5lUiBV3+OtxW5uyR0f9hFSb5M162ftusQWqRofH
kanGfy9qwM6O+Vl0L2gHGrbHypvwzO6FSDP2JM36GuQ66tVfhoZqJY9XLhAIBQww
Y36jUwKT3ILZUD2zbaAI2N8FrvLmZOs+5SUtrvSLPnktrnbUR/RM4tVbMExLt1q9
iEztvtuI5sTVT1T+2qdQXC1WqvMNQp/b0zV/r1gg7/ynPOzjEvE64NLJ3KhzzsiQ
IkwkFtvh7eqM6+Au69OQe1z7yRF+UFkZqWInBxbvfSnrQTeGmc0c3bdZITPopwwd
AHdhhphUQ22wvVfyqx3MxSqeMeJ/28K23ecq7hS1VLXKHq/CjI3L/9YH2ILUPqk4
LfGn419oXfmr7rDw1N8iIzgyFS9J0y3BWEKG1CvoJ5vQhj0QsuSa3Q2+1xkomUAH
m4u6J4kEBZa9gIflLrAU9uplzmFhXRDjipShd/htoulmAmWk+i6K/ESuAFy3TznC
spU7YVaibUrX+HTRByuDKTegOaXdoFAp6YyfNm+VjlKwrtsudKFz7bLA94ChRDKt
QSFT5RNFJ4Itb3cF89G2ylZmCwyzci3yry3TFpdF5H0E3m0LtN25pZ83IPI9KfN5
zLfefPSb/QyK03W7oNGHRwahqP6iTeHa/0mnNR6WEsjTjw1cI9LeTvG8kcLCB+gz
ONerWZGDlHV5lnqSU7qaXU1/x/tLPnHuTCmeWy/vLM+5esUsOn341N4zb9JBkj+X
f9+8rogO6hqxwELFl4l6hZ7AIwuUP7kV3vEJaBuKE9X7S5ciC5G4S4nHHQhaNmFQ
R9CCRMKdZmRMCvJsyv9OYOjKc1DtmAV3eD1x/81+7bsQ/eUqIN4+QKHTWFeKKsao
T4L1XnNw05buWkjLDeNIoHf/uxuSJhdiP/hRALz/zngIVZYjroDU7vffSVDSiTdf
oR4WQF73Bcsrl/QAglBu0d7pKTKQn5UDkYq7YhYUJFlhvqfsedoEyDr55IofqaEk
mpJuAwiXnLqENLJ4iRlkAVqyMHoQOhyMxzLIJoUU+jlX938eFgIZp7bzAm+zXSe1
+NRCRmxtIr33IqQ2typ23W439j0NpFISYBty3UFZIJwT4elB17x7lc6bCezqdRDB
McCRvEiiADAOd0yGosQk5kSmgZTzzJb1dYCXHkO14ilNID+LJWhnMIA624+u8K6w
SCGbeOgpRSwryYOFwHlBBDT9vfJ094mGM3lAy6UMBof/OKuzTq4rxCFLOB7sJfLc
ZawMQy65/aQWvbJLSSLNFM7aiNQdI4rjNrt9pyn4wrqxlE/D4OC81CT06hvi3lOP
jSksTfnWXMk9Q68n6biAUaHY7T+zaSlp8C0gNaEZ52on7JL57FopgMCtj2leqOwi
55aSblOvD1g0bmg8u/GtUkJOd6cSVkmCbN2mwKaVKoXU/X/kdL4vKk+pIaA0kbSn
A47SnybHvJspoh3aXwVHqzOHLKhhNu6ygBBXNCWs6p6zCVEQNKERzqA3H3W2UbfC
36fq1SwbOiET9wdFhMc1SBLwgDbGSbhyxGZ74az8WvBCuWE/Z37XWk/PaUeQEDlA
vFE+fqiO6tqRj5NwQwfVpq6UeyGFUrEDXJee9w434un+c9w4aEyqgQSw0rMygxKr
hhYNW3GbZw/SoWv5/nI6dTyRDdQamQEYFCh1trWIMDkIn3Grxna86fXS6w4rcftm
O+s98jPeFzB3EK5t/ioUtJ8Scl6z9BxLmMlq104qRmUkyrQzojMj5qShwkds2FSF
KZofx15CLxoFBMr4a39luctL8hMOIq7P34SRyt4YnAD1dPBqonPUBBCuloKHdnJz
xBHRZW7bfTNqQvgpGVMIyoL0Ntau5NvK/dCvI1bjwVn6aXUtLpaW5VYsTP4djQdZ
p2vXq7sDhE9b/Y/wNzI3v4eXpIlga5pqgE8pWg9y5TiQGSn00058NeEBZRezYAa1
w+2M/AaLkdUTL4m3U3QXH9oijNs8P7k0x+4jrpSJTKUVnvV+XuCdEA3/OetZuql+
CbP6j5eqMY6dgatkwN2x7g1BnjbsZko/Wz4NA1rK/yYeJBlnI3kxrfva3e0NPDR1
pOngYnxqlmVYhvoUVcGuZqCozP879clCBQ2G5t0deobliCVVlAPTFHvpbXBei/mw
YaOr9oKSWwc/B0NEctSgbIpRX4nxCJ2o+S8953sBE4dK6SOCXlwVsEUZ10nab6V7
Bg+mKSzfyNsagQz3e6g6C+Q9J0ozDMk2yOdMoDhfDlAsQxjsvn89MMIYnEcO3Q8m
wzazfrOfdMXA1xawZW4hXIWQ2QRHmZaP6NkhDFjlkI394zAGfGKhduD9CgLdFhFp
coPXovZZsL3nJ7E7PevvAR540iHo7TsQGvhQdokvzSAGMIqHVszq0NOJtAcEWNmB
RA5DO+xR6YaaUcZ0Q9ydRT34LLnvFANPJrWjDIAGpPbeXJagoVLlXM7UvQKk3eG+
Y4B16C+NAIKiQ2Wk8y6+Efjof+KgzWXzPL5EqxTfIgZd55P/S9jg2n/4wpSvHpWh
AzvCkinb+hDoZciGG5MCust1QvKUo/S2OD3q11/jKZLl8/9DBvWDYAZBXOaiM13x
1KDX1WSo5N4YZNFWhu6oMFM1f68KJJFIsjTCppuDhgFeFDOM4eUcHIYZbhdR70hH
d3uq+nND1gZSTOrh0LUCcvwrqhsZ3QQsMAStB5gZGf9GXkyR8Qu5YotcJ8OEDlsD
jEfBTXg5x2gb8jRPvG+qEfcd7Pvcof85iLc/K5oe13NeO0L96Bg6NgDD8fZMvjlB
b8BPvIWlRFcbT9jej37rPLZI6d/CeFSDQw3M+hYZEqSSGn6OF28sRJFOmD6K4Sco
KoECyQZeCu0sk0RhJN40VnTAd0Qn5NobfEPXgvaONz55DuabXI3Ej5WjAJ8MC0IX
JV8+doNS9Irq8FR9BcNe0EH/LJDmN+rcCeMbvvhHyskCHodwHsW72rLAtD7OfnwK
sgnbhGAioBMz71YniaRpSgtfUlP0CkXNLwg5t4Zz2M+Wczhrjy6X1UglTz84j0Lt
rGrivu0lOBn6Yb0AqgdVsOZYUSzvYrx7JNUPy1GnTZwiw1jn1X4OzrDzbSWJRMvC
1tNMldLgjtcNX2nLLV26w+u+VEw+I0asAiJpvp8rADhDIsozRayDnlHpgjLNVgnR
HJ2oIwCPV49wl6oGshDbTdO4EMHLHFcT1Qq5jStyFG1kLFx2mHW1JfKcUA3fppSQ
onh9H/oflmYzw90GqlC+0gQdnbE72ZpR+Q8QFRxdwxTI11UpKiDjvKVs49shdxT2
h8KW7F45TJLwcEsPXeeg0gy42jqvQx4Poz+SN4/gDWqoQngvPGdiMHK9XFJUiFQ7
KeAKs9bvxVoXm851zXZUb1ZSRusBDEOJ/SawfNmmG1la+6Z2Fb4eq+3vnyn4EZHU
jvCmpGSRYYAGMJX+EWyW3SWCna3SZF4vceks5MVO+bKLxlWMUOHlJEj/g1V1Pyvg
Ze1PGja8QYpFRpLjb8Bi/kvvnTow+wU0g4yf0rcBE7ffXQjG4V1IixUTkpgpvCkE
Pt7jWX/9PS/ad/74gM5g0JeckY5RmmUsPSo/xoVSg9FCmdWD1mz7NJJaPuNacc3H
5oK8BPtcovJZFtYRc1/qIQ3Q/5RNJjEPqKRrzTVKwfJz1u0r71SfygmbzxHeSg24
1O1wgN1Mj6ovku7pwGZoDxNf3EG9HUIcP0BInVWBkHDmgbW+8kd5oi6/KWzJdY3/
et/6eD5TyPXNG3rx1HDwgezuRigjcvgJTJP/EH1km4/Uw1iqNPM6Hrb/vkC5y7lF
jWDUzM8DzaykDQvBe6oOCGJhqDq+8MbSACJSWx+r3Ska8Ge5SBfo6To5gDNldyEu
sLM4QH4ZtpMnnhWVg2mLsEDjpd98vfrUJS1s3oGOd164mgT5HSCRgv8GuPLq+G18
H7+0w9jJ2L43DyUjQyGVe/JfD4muytOOxpCxYTN7dGN5FYjgDWUo7LmiguJP5Z1e
/yvx2Q+5+6WG54a1sS0OohH6NtgQSRglklJFZ4I65KLSRc1G5QT8DRCA+TRXJyX/
u2kwl9cbP41yy0R0QsqaObW61svmgykGTHbuy2Fjq0OZJ0WhBeFu43dJRHOkC6C9
oK2Lj+gkbJoRfacmi4maKiE9gps+yueUG7pp2r25j/v/qn4GlpHa8nKqejUfV6m1
L7151nXGwk8qH81kPWx1NMl/WBYkzeEqUrzLjUMlp0HPsshZtkTEff/ZPP/xG1Ff
hRn3jjzm3+pFqudkRdI8+hI9uTVbq2m3o3AihoO2wJCjb7iiF/CAiDg+ZGp0u+7m
hn+KeuNsVmsEEJY3xr/26VgCuTyBQhFphhtRqGynZ4+VpVYWdN1VmjI3qrIw+EUk
4HqfTZwoaxeCayvUzFOILDnDoCBgvojfTCm+xTWotEkFncBRlKvpjOvETQGi2bx1
Y/0QQs+sCZuPz8k9W7K2iby5E9d2/X9+30u//gHORYO5rRifPwClTYCko88fVet8
P22g+nXllki8MbQxaZPcCFbrysASequ2zwiUUaDNMWKL3O0UsMYlw0qxY4SgI83d
vdlt6dY1EHPm+kZtw21JxdxQddKSiZEM9gvY1jthObkoMzIWEe2NXo0qWAEuIp5a
wSqxZGJGdBKoepPmbp8z7pYNqXc3JVgpWyiS676OpNBMkWVSxhFZYhhq0DQUDdWj
WyacVaKRquIx1AcexY7pQOWKZ6kFiCX+8MDbWmghWBK6/LnRpsuYJuacWeD672Pu
UYLLonVuN/h4plupNSbFYa5XypS2R0NBw8GlYTWziqxzL+osRc2kkBtqkT/AuViC
h8yZqcL0sUGLMi39Uul91rtIcZ7njqWI2GhAnnCW8VYa2tzaJJzGGuc04gFX1RHb
xpwYt/zrK4qbNb1PtvVmaJtYBgUDScwW3afXfePwNnGJMYirneFLgcr1rZVZ1kl4
KFIHXtC8zwmJdokcOgULHakpDhJJ3nM74Xndmd15KDvA+yTyqtWQW/0iESwrI9iG
fRpY5Bhuc+l1gnxCiQvDtzJTRXOpEWS8HiDXAkPNvgcXoG1tJSmzkfgC3/rG81FA
ghRCt/YqgQSPS/BRbDFOsx8AePlzzp/hyGOdzyBfLD8CCjJ3xMocHY9Sj9WJGWOB
9iVIGZU9pukfBrkeU8JS8Tuqj4qzYmib453xelTREdgnfcniib2+Z9iJthD9wDzq
Jan4TNhTbogRzFJwO/adP1ZAXWY2tDkJU/LFHZSDVOgweAPoA7RMkkNIdUxF7OEg
VCRcOoReUgnTATw7/qpuUPMx8sxL7vXQC8nectwxgp1eFAvZaQVV9lVNzWNJf8cz
p9vjyKVomdNo9L3qdzzXQa+H3p+hXJnLDTelDYQeLQDsZNyw9PItfqNZDELNGuLd
q7H9jNGxK11hRtfVXChtwQi2ujeeUsv4swj1wQxQT300JKLBKnsqD/Ikldve89Qf
QrJHgqJkP9UzWIqf7dZn9ynby7J/TJimeZTPEKgE3/oUHRstWtcmD2dpGxdY+JNS
Cfd2DoOMzGGeyJwQ7ZsWQPbOojlRaQycr5y66Pm0mcGUPBkXuT4r5U1/AfpSW4ew
27jNNBCb48Pr1cSbF8S7tep1tPkRa8DSA1RVHpzyKXz46o05xJ3uw0m1XBT3I9G0
szqIQI5F1RvVSUs3LCcd2AoJ/YYY51a6wix58dyTYJm7LbgdnKUcJQpRDOTVY7Xc
G7d7c3tvTSGZT2iwgITU4VEeRFYyiL0gQX1e5VIIiAwk6T+cj38BiRl33KSAnbsH
dgI9LupXlho4XmYWk1hCH3pCT5Z2uboSRLX9So3hM1bYKsavA93qjdc4izUOZN0/
WAmfUwE8fv36bzIeHnWtDiKumEsB8rnKzOAo9Dit+qTIznRK+g4yQG4UL4se7teF
7ZMqn4dSiqEJ+koXNT6b969zPlucNGbA0NaauGdhb9v/auiwFhyOXu19xWUHnlIm
3Y6zRZ2gtSush0/2l32H5IcDblMW9M/jHixCk+F25sWvXFWMO4P5imm8LeKRdkRT
Bvs5H/jUlhd6S5gLmuvcNWgsRJqxaFen2EwX1s6lIxYTQH7vHiKQnNh2CQie5/4y
+ujRX6QBpYHfWqY5K+iQrkxdb22wydXXJeRkjWjjbTsGrIl/UgTEsfm30WjRRKt3
uKXNfefWEze9BPdcrfRJ4+GHfH0HEqkQ/tCjpqLmz3l5nLbMY5P20PZ4YcN2ZJ5o
SBFG4/NwI5sXYZc58YDaoNnyw+FixhbPGxOcyz6FJdPUXmpsAOdBuWTDLh8HXdR8
dVM3Uwtt5rC79pmGMN5+pGG16VBgCOAbF1vy8iFgfdZ7Gfuzil7wuzpPlygxrZy5
JDmB5qtoaP2qqtDUvcfc+gYTtXiy8JkQgH+NS//MuPjX4lhKKeX5tdttBh/MsyXL
TXYKk4VY7VnVuDj1iwaWk2n+RAXM025AI/V+mJfKx583bbvH0ivU2h6sk1/1MEI0
aDoeWbOY+gNr09KfZXsGaZEIDNy9UmTpAW3WPd+GYlmvgqr7QBPfoolcgAReVGqp
2zP2FNIHlKJWqhW4rcG6UtHSeuPrVd5ovKTjLKRZgHMvO3I13Wb3kYtifNi3jHYw
aqeneXvKl9zBScezBW6L9twPiWROYrYUFmmKYiXs9AZR2SifVlxRnbAKqi9qJaZX
xMS+EK7d75knYc5rc2LsgZDOBcCiM6toNn4zCPSqxp5rFnRiL+O3WbC1IenawscI
+1mDRVk+ldaj+Qpz/4sahmZYOdyqxDMB1QA4CFNw+/4B+1tFsR2LJkx5aE2+JJTK
Zz/h/d7PwrWMaQOlk7YL1F4oQD/cE5W6YwizqHAYOVQf2BHrfxut2bI5+A13cGy1
FeTmlgAIk5Tpy4VoIPUNablmazd4oR2A9TTxmZNB9E8ncwr2pFJNq+VK99JlDPdY
oY6GlcmohG4ghOqHaCdHEssmHRGcrItB4z2JkF+ECJ2csxRjk2ZOoyksCH0OUcj0
4+H67pNRldnziRasXUmXqKhsNQet9AQWXA4rTPc0SRaVmmC1QcApZtztgeoquRzO
Y1OmnMRWz4dqh90hDy5in27JaDQ8aVqvPzj7W9snbfaT5Btc4r+fucQ9/y+MVGD0
Lvwz9MWHugYcdH1hPyQSsmzwYr6OmgU3HCFrVipJJVxKd8NqjdX2CFGelcwTlzXT
7hx4ah9nXjkxefzGv9Qm2539WG5FXA+V94ZmeaaN0SJxD3iPfp1VSN8cb20eE4Io
sBJbXihOiHenynuXsJeA9O7fyVcxV4U5aWgq3FD6f+Ddd5CY1iH9k+D0OTW/PvdR
b+ILK/9i+zP5GpyGwvr144ZMvj76WD55cbcD6Q+bdqn3PnN3Njbqpfg3DyKHNEyk
WMyo0gIpK5i0wJZObOhUi+FYPW5jZtD+j1CXVd1YG317mNVicoU4wckiBULoY5FB
tT7SR2iQysW+6xZC21kFkV12xsLVt/9hgXIu6w1JoBVxlq/KcM8+9nYJQwJ97yEG
eVVxpZBRv4nsrce33SSpHowK/FYOM/s6T1Yy/Ev9pvOUdsoxykg6l8WP1SUhzMao
6s2JNW/NN9gA2JgtpPfdnEdQ61BCVEuf/n3+U8yh3cnD7PqxMks6hSWwr5r0kVB2
g6y1bKCmaHbOKL6kj64fUcAB6Eymcqj1onAyYtFW24/oFML6zIg8sq4jjAhwWQbl
uidY8ZlQk7YuUbAlXZz47QLe1YspGNZFZZ2TmCBku1gmJbMyvghg0pdXThuSzdW7
OVmzzvZxE1QFGR/YYrYnCTo/fvhaGacz5TTO9rtstsY7mL6X+UvSxT+mr8sXxFdo
BOa1SYYojEi3ejA8Njn80l1MrfoODL3K/W1C/MZSo1IB0q/qCnbviyquZ1OP82nO
Zz1H6w9pNqmLg58DoQsCZ5TblQdaMJdkCNXQgf7wEVNl8XeJjiXbmZNKvA8XSV4C
UCK6fun57xjLV4PV5yoTAmmsrM4zw6BglcOCApenVzQH8qN3gEFkj5Z8e7xAlQXj
Ck0/TJwaohMOE+uUrbzcEdObSgCj7SWO/phll/YeA1LoNsOmn1ZN7hiMtq6V3vTs
ZNnEP/CTuODL/wXsFp4RasDvd5xsnQtzfi/pWEnvwIeJ0WJyEuBSgYiZHzKhq39t
dAZjjn7oIBE7B0Q9Mp3uoNeRmPuQ++nAUYzPNDKSXCYDS8ZEfljgIZSfONdu/asV
/3sJVlrKT4qG23RFUHUdocywJFi9wQixYW6G8w1+kV1mGnWcHA0QKEpOb+9Kd6AV
JgHnXoiMV6W8wpi8N+/OI5kt9h38PtMm8rytR22e1Y1J/jRPDyx3xDMZmpzJqoPK
EIeY0QIt5F5GO1hTLD11ef40EPvpi8T+CHdkUjwKfgWs8JP1ID/v/cCpUcun2bvU
ZmfWpxIG99vt1vg+drg/5Q6tSZuabdsjnjNGO1uiW11Rs/8RIIUZFgfY+oKRwk8e
5aZFSyWhBt4V8KRib9XI8PevHL8NfRktyERrNUjRDkCopib5Rwi7kkL11g9a2f0e
+Gh5BTsRZ8knImJ9KYvE1doB93bEmopcMPiR19kYLSTWMiJeImh/oBaeo0D252xs
Wmq3mnB8RJIL2FCcUpvsJ33AQNQXbYaEtqB6mgB98vAqbtPMGPY27v7KP4QIYpjC
PhPWlw9ctQ7QSCZLHfnJEPNB4rWHY0dkbwBwLW8dJcl+SpefLioaE93kJck6w1iw
eBy4JTH9AkvUVUX4Zfu/7GLDQBOiDyvm50jv8XJmHm5Jd6Phjhb1Z1YWL7p6ZWbW
5+URsVbEej7Y7XUcRIrxRXNriYlHook9mHb+ROaRozRj1T/qf+NXWGLHm9+zA8U1
zp1b6zzwIEtBU3p5hX6rxZQdrOGC2MhJslD/jdEm2O0rSl2tJ/ZW1aCAwarqLhkA
05TqLtzDHNC02KKQrIa/zGusNMTfNtMrgsilgcC4/jIcwWyQmBIXxr6XPyqX5/Bf
6G0yJqiUaeOYs33/RNPx8689vvqnSBWGnhvtFEyR2ZomamJXkka758A7FV9v7URe
BbVgG0eu16fRiv0uL2n6duvJdaYZFMQjXff+pOp2EAyGHi7akMnkHZ8Hz3m34zAZ
4OjSmpt5/jd2DSrLuDJB4okyyQuciiQiRZvLH+JvctweddXE19kslO/xD1UPfkoz
Mk6JyNW3OdJ663JumPH0enaypq7biuo3JeWDO8ocksKqWzRtTYusZZnTSAugHp5C
KP7hVSurO/nMP/4CJVN396d9Dm4ZaOL+D3T0lG50RJGUIMCvnG3qUWzyBYcwwQ33
GONKkVwYxNgvrDgX9w7lo8gx687Cl7uuxuOGZo06wFr3BRHHzFmwb0KNkRzdn1Xo
iOsL8kfWqZEZ/ouraVHKxT8diOmLrrYI4FAqFvYxgHwLWXhd7T29sXmOO7mbZbo2
bAtkJxC//Tc7vl5ULu3AEL6gtfBX0ZeInv0LaE+LuVFr5gp87z93T9U4srb+v7jE
hMTPQeF+1cJyQtBvMKh5ywnJvRTG0dpPrY6zQU7s0JCCutWpbbnBfRm7ZUszYiol
hVh7GiB7qSHzfH7idndjav7jo/+DjLKAax98cHXwqZk21N7JFRgkpp0YFvfkFa0W
v0J/wDVg6XbMDc0Bzqrz0rb3q06svhaI51X7gh28CcrQmb2it98SPoowb68S31oJ
RJ8jlXbKQuJwFFz0nwxi65VmnxP3nO11JYEwC1LBIRER4qBTG654LEa9Nm3AVHj9
KZv33wXlojwUrM48QArja6vVx/HXi3FNdDLrQDprL9kIrULhV2UgYMkQR+VDd33I
4kp9fM7kCcOQ8UoO8bmGNe4vvm7sdAnPo2ClV/FZ+HaEUE9MC/BBYOd7oOCkwAJ3
bYxKc/DqPMrypumuj6S8KXYRCUBldebijHrUDYvNB05BJF4ydgsG9+ZgrnFcOK4V
ZojoSUOv0HW3Tylgz2Ti8iomHFQLoALF/AjYq1JF+9ZLMYm/raBs9FzNb5Pi+gfs
YwHbNojZIfrVy7u6wKBEh4owptHDh9p6+I1HQLz0zW6fEzolZuAApFmrmZ3F9eAQ
AHC3JiZoz9jvlweereHcYb2rt9KprtI7yvHTZ6QqEdsJ75AdNZh6EiMzNsXckpd8
QW/kA/4h51ZOdEYjUUHnnCP7UvblIgtLxoT5U1DAz+LtUvRq6t9eN86bm3YBmYgP
sXgQiZN97LyOLUDtpL2JZ+d8W9Hh6tQBMy3iP0gmCz4Ua9+sP8/N4BBUms+N/RVS
7OyiCWoh007Bg2oeZYcKf0a8jXe+l/7snXTai/t/ychyhaRkqW3z6l7J3XMN8u2c
EPXQCDhxA3bfnWtpz1l8aLqzVjut05VBK8Ln5qPnl0Vn0dX8WNpzkSzc+Ajg//ws
Q6cEAjT3XbSLjbD4XwWyTpwqOEAfWApzc/VhPVYErD/H/LhgYm4iklsuQwaLZJKw
ppq4IDpiz7WWEIi5UjNBfkQ9s4nDeOLj6PtEKGmdJjxSMcllKCTnnnFwfgGjL7v3
U3B2PU6h3NoCFi7UVHVJ2GPckOCWtO4lPlbS8GdjQKllVAsnrjitgamGexAvK545
dZYhT/JXflUfiJyWHG0+iC1kngIvTYGYmF5I9LzI0wWmptNQMkIcesFl4E2NWczi
JiN5ssVULgxhSgwybSaJSxVbTu+osJ282XS9Pf1X0MCA9TUBdTiO6qzWY/ek+CdP
R4RTlyobiWEL2Fb+Ph5sx7dpZXw7wdURdQ9UcOvIYBNnUGbGLKhbZP5A3vi/+qqM
tPxPQahS8UHMFpIPrDQvxZa3ZEyjsDxuQiWUBxgWcvdxZXTNW5bFjgkGGGsOZlpH
e7zAf419k4jAo2nC/SJWMwtDCyg5aqjjWZnmZ9rLLBc3Xn0wymRjy4tTOKmBd2Xd
ZWHXxEvLgpcaXHsH/0tvb3+jVTVDwYM92YaY9zJvYi4fVcjsVOWdM422KiP/5Cef
qi7gYCoJcTJGFulUJonfd3t0bK1kNn5d8txp9eSQwjQZfJ4h53napiMd67s7TLFh
qEM75On/ZFLfrShSH/d02jOwI77iEvNE+Y5wAHA2FB34gLOu8nIdCp7xtHgcuDp7
LJwyPbK9HR11mzWP2Om6U3PjAmkpqoNrAnE2/lHPX4bChRyVnI66XKLMcpVEfhDw
fj2ylcoOQ2YUj1DtU7lBrW0BileCULs6E7BUI2d0zVNFK7reb3176Us8ITKryyzt
hhNTtIuR2cnzfVAc/SCf1q3JiB+F7ZSli8QBhN4UtHCwZIws1X4kEADlfObGjFWG
wHmJjmk7y53SRu0MZpVfrDOxlQj20vkGLZUGajKp2WnJ7+eV25TDfEIKj4jVItRh
8dFbyoIRPe8d12aiyQ+UqiuGZzB3xBFdijJsr6Fs7Y5b1eFIrib/4Qx1f1qgOHrY
CSVJCg9A42HEmU3SBkGGjftz4goxNdeMY/eMp9ydf36uxNnDXDWuC7wXQh75WUqY
WX8KgqXpZR/6/SR9MVp/L8/JPB3ysoKcPI4V7uwiq7Hjzg7PlN0Fo2ov6LXGTMqq
Dv9SAIai3n0CX7aJuMHoVD8cYMgewu6QW3dcD3QjWZo22/uYk3RMgDK4tljrbYr1
ATIuTTAQnj0cV6Pmzec+kmMyEaReznaxA6ITji+kerERZLrP4YICvaWzhlnNGFxu
xfcV1zH+eJ1KA7zQF3h58tkbNvEahqa+ndo49etlgP6ZiAOzqs2hUWFKSIFVrM+F
wkp2HviYy3/6AMlxHNtAaFmF3oW8FN8688PgdetPlY1Q5ZGFORpqVR3y4VD0SEBD
bSrmPqUzBX/uP6+rWwEdgke74728gEdBDqdDeHg8lFV7iBBeTy0VcihnPqGm+0c4
2+EOoZv/PCM7EHD+xUOdVREgnIU4yPMtRuGu9o/6h8iSBC3pT141aV8ynv56cE+d
0Vi4VOaETgiHqVj9hKN/lwGmZ9w6/fUhf9/QXPPMbiNJgAy/VR+NTVkauKzxyK3m
8XMXN23f6xCJXL6o8ukdPYaJQolW0OG0qgD758sAUcQFIWwGLl/jMshuSljjB58Y
zr9wEEEldMTbuxfN65H0bAx5fMSNiHt26RQofQCq7oegm0+ngSk+/0zAL/DncERc
GBY6kpLnUVJseqD22HAlJq8oMEqay9TVr8zKnTX+lJ9Oi2+QjX/IomTxLqQ94uEE
rHp5FoS00QIkxx+6mjAUijENd7PFHPMTmqvmddskz++l1+Skq22VC2C8mauyHDed
eNHUk46kpsV+LqC3v/vqsDw+i+KLhI0Brf6DdgPlREEsAStWy8ornsSJTgpOWALA
lc73a4VgNKQWvril2p6wXtNXcE7qOVXVumzITGhC1/TeNrON9M10edfpZLoW5llE
sc06PgG8m9FixJ9zUDr5VNOTI1xfMkOWXZAZaB5dD2H4y5tr7nf9s+CC7L5U7xce
s7yh5yY0yOSiIUU2x3XPX1mhAmD4ex+jqlPXVerVZfpK8Quw9XoE5pPPhKBoZyA1
+OWBZ9dlgGvRwU+r+z6ZBC4AtJ1CNj2cVZq9lI30V29ZFlK3icJGCj4ryqb13m+w
57qulkie+1aKyVKOczJN2Y8iTmNAuqygUJB8n8FbJ5lA1ZQJolbuH/Thj5vzkuy9
Z2t4cQlIaNPp3E2LRj9YSIV24BH2kryqUlm4C60kyZGz5eWIWLah/IY/OebEnYA2
8nX0eAey9MW7Lkpqq3SSALmcxVrzOTMRyirxjPhlmKBQCqrlox5bZlqGGBfMqLuC
SeqAjGYSZ+sygI7qSB6K+dP6MstbapvXuzTFQ2pTpgQOlKeCiZT7PCTngWDMc5/M
gyMKpzwoAQmF9gmHDztyDp2JWy7OemJg6om+VmA+gpx+08kCvuKVrOUhufArIRHX
LkN8NbIVtBfBkF0mT45g06wgoB4zCO0VPg+2gdnv9Confp79FpeznrOFuBQ/SlGb
aei/T3F2Q9FD+vEbactFuVwiyTFv2yKEwUNTGLjtawkdoc9F3xwG8CpT+GAsBmgv
Ku+mMSp3EEIfvVPoiB9Cwm05RkG4ndLh3VSSr/cyaLBq07VPDzFrU1lnVZ3BE6hd
jvnDiTSzXlDdjfxSZ9onlJCgHqSx+vfoLZvnIMpeY/xH8adDXV969EmPmDff53we
ZNdmGIJZF33HOpqdRLSks0UNgDTwDIZc3+U8VaAiWVHhgn1kEqvmkC6hMQg88ZUw
b/pk3BojYZIVv2Rf41l6NFXcsf8WHi4Ba2rWO9NBnYNQcUEBJNtnjWP4EO/FwvgM
8CwXGwKECwLeOboei71NHi9xLJ8DA0S40aN5/aENEVUooCOxjk2HY2KsQQdWd3SY
i9npBgpwxz+R6hOJYpx71j7EgkVEFQ3ByqZoj3QOuIfI+uzS5vSdI0QAbKtZWsb+
WyqSb/iY7vuY2z2f1Sg3cujlIxpiI5U32+f+Cb9reXBZoLhj1mnvOznztNEYYrOF
WktLrCm6lHObtDek2tElwa1Xlx/4ElVU/nydlDvbv1P/aG405KcxUEHl+8XGXZIE
+sQuopb10wUJCU8cQIqS/OcojItFUUSyW1Wjnf7h8skCRLCY9sC7nIUDEu4QeBkZ
5yAev+anKxZR60oU8gu7KAnLKhAzXeqHKuE7k88qqLjnbivL278PwE+CyLcgyHiN
TLL4Ua4nR/BzC2hMbeffqGx12H/BBjKu+D/eI9q/GGLCOcj0oxCPuz9MHhv49VOY
zPovizXh4aHtEEUDeRZYcYKjV8eyeFuWYzC2/qdnNkJmTK4mUT0E12M/5Ba2mVhj
tnelvCDx3Cy7CduojguHpsbpU62dIbMlqaAUfBdMDOrwhdL6amPtGZx91Ln965op
QV1AAjdTjgovMICLjmORa2OaKakSJCI6jNP4gp8I1xzwur1VO4WDh3u6DX6sJzGz
7Bd9p1ZtJcgKF6N43Dd9+h0lj6XHpCq2kxcrh2hJMrEo3XZU2Sf+naRvDvyrvux/
ropFjjBe8rXOM5u9IUm+n9VkeY/qqsg2ox3L5YRvq2L9CcI1jquFWy0gWOHf4u+m
b/BHWE3wWU+6XE5BcLLPwHp+OK+Xt3DmBmo8kNCXw/7IH6d5RJSCkfw49su6gWkD
8Ic6IY27Ie6Vz6+C2eZDultdI9dezE/xrbHlgOY/LKD347BCkBXdkTASW5sreRDZ
NsNGA+/Mfb6E7FWbRQOoLOgpshzIF5LAKfoM14YpjDWzbZdTybjZ8fMdT91z6kko
D4FnUSNylIEh5hpoEGATF6Ox0Fy3ddcULAiCdcpJasNaCuyTezbFc2MqbG/dRTlr
cJYruS3m90QtvU4LaI4rSBWYko7tJKPCYozKN6u0wzwk8OLJaqEyq/Nsj9w1B8kR
B4kjx0rDOUxN1GdhkZ4XAk20KWOUmng+cqkfav2g7liN85ChZLUDjePN2+p0Ad90
MYdd4UEQCGrJRlSXfiImj+z5QjjzfFh5wsPkekyi/OOKGSnDdmI3WUXWg/UiE1Vv
qPZn8nH8zKT9sdF1tNJPEW71F3Bon6RovscllXo++Y6BjcPon/SaAxXXBGlnsEr0
aaIMPl7GiARs6XphqfYtRZs1AuJsrhxogucOyrENiHwhjb8HHdphuk4y5thJkX7l
zEEV4qeEvGSzlPVJB4f1IyeuRsEoSWXa6GfDZaUkpno3nKwJoHaLmsixtArrQ1V4
BM3m43MC0eh+S2PF8+E6mjVpI1pHMCid9JfVSQhHUvEMz5lS3hYRYWl0MeXinHmp
fglMlrd4NJJlLB6/nGpMXyOd6kCTN0fCVxGh0p8BvXw52OyLNVvRAZtO+YgH97Br
qhZa+qeGjvFY2iPpcPT6eObh3VBkNHnj6Sqsf++rPZnVaQ6GqsDYzGSyEHP2FWN0
Q3pjOeqcuLFPfdhuTuKyrqAuqUpoB+uqWgptUkyaEkBRHdfp9LZJQITijDxCqweK
QvE69isPvmKFcHOZtyL9WAKmM5SDK2Cm9ptrCHzdOKMgISJgBoLqay85XW9NrGJ0
hZN7QQXpckECbIplBvL3XHqSDN29JpkodzVK7tkcXlqMwrNhxyZQWaY5e2ug/vbu
WzttktGPDdUuf/bmz3CZeZDrDGwQ+DBUKaCGXIUzMXSo4Jlpf+iU+N8H0kRxE7Pp
z8Iv13ZnGG7Cj5iVHdFZ92Yq1YpXgJRgT0P5VAI3070Iy0q5kHHeKnPl89QLYsdk
c145VENFeBelMKSfF3UKCEbyraQzaUBMXAlBGk8zRaabqweJ4qfSyAUReTgMDSk1
XqRgZ4ChVYa6IwNUFGNtW3iID9RLxOywkRvNF5UgGA33AaKojGd7nAoXzcwLXJhg
1yOtZLhlDxtiFBlnCakt+jFnJMFVJ/TF9hNxCRIMlLxfePV7zHhVFtqF6r1Ao8Ba
VmLDyf8OaC7mW4e6l0RSmOSWkF2X3VvQWFSN7oC5Fq1XZZHR2QgobQcXaxAPMWN3
nQZzbzGXGPFid1MhkaTIFCIHib28+H66PzAQDbtgs2taKPLyPQfUvUB/KhP/RoXc
Ncd6Ib2Rmu+UKZ+wUhNWOq2u60Jfj28sY0gAj+mir6rbiux6K4XP95QGsM9Svmvq
FTJxblKbnKbdn1Kw2YxMWVMVWTtnMy9AZUMzNTWvXNHDOY3WjNvX5MCsYGDBuz6a
KzZBp0JKjdOAkMeH3oC5MTVGtpMgLoQ8/3bLBUQNu+WksPCPErdPXW8n5cOkq7bn
JNuGSLcE33MMXRUJR8COZiFkBaq/ZKaxzvmnrLmKIsa4pz3RAYiF4qaAhOtyKcew
RSspAmwKH/o62kWv/64hm+E9Gdo/x/hP4oXi7eU4DaVj0GW6MYyHPrCXli1cv8Vh
xyOUP9kxyw7ygfr+A1x5E3SiNfbxnSrngogRYVhGgwsokDLjWaHTMxEHoLOjJxzo
meYNFCDwpsxTBD/RRapowyDDH2d4TCawy56BM2RBIz3+5Xcfay8KXifGlXY4ARft
dB9jplaEVqCZunQEt1qJNpiGs6bQJh9d72jXr/FH1DsrNmmZLWlYBYIPN1Ee/LRU
0x4t5v5y/Pdgt11XyKD/7qY9C3kRKsWc1SoH1mvC+LOFvM/oXOJ+7XqManGuI8rX
IZshSHN7J95rzRwapW5wy5Mr/ImJnSlKJUTSq7FnX5gh5JPMRI5jUE8kBTNv1nD0
R4aODxReUUNJs5h8BiPINN59BiSgJKIdsif1EnnMP2nYJLfM3UDpw8rMXb6uAPwV
D+FdwdfdpWEU8mTqEKFcyhekGA8QpykicXaOyl6nheJNm4EhkDhoJXEpYVcCYlzp
1sgTuadhqlAPwFCRv/mdtv5hRxibrAhl6GG5Qr2AMiwGM46inGs7jXCjLtVpdEnf
2MFt3agLDaNOVhk8AXtRsK80BQc6iTByFmhMuSP3iVnOGLZ+TsGrAlnNO1BKdHZp
o51Avlp91RYgzplNu/rUondEXH8ydD9Sl705RnNjITvfi/CPea9NM6dMUy1KEoD0
8O9hTZqM+bjIug3h6pPvPVXmdLj2pQJvt0VQDPMvHN0fbmh8pDfAJ4SFbKwdFI35
c/7FU28Jb/HgL1TxA/KVB1iIZekGMlow/OdX4sZWIxABDT0hKC1nN5sCrCRiI0Hp
yyJYncaqD1Nhau5x9uBJyyukXCmKNXLTQC2jeehbsT15zT1/HIbRAR9pk//6xeTI
r6Lgkl1F/uGWXN24pD4rMFQ4Z9lAKdvRjkJkBZgtDJZxNpfV+6ghZniYplfWR107
E8wkVnyLruO+vr83TSZbdT+WpK0dUAt6/cZ/f5LPGjsu7xDTbhNoFAT4Flrt1JqG
YS8H+k1CHLhf5mFSl9pVC7FcKKlAKNAYUpv/aClrCEK75pUbkhjLYCbtgm2X4qWn
cWcuX1q7Qf/KwtPhkkJZ7vZgZ/e0x/6QzGGD1BEuBK7GeaAHIMm1IVmCe9RsIxyi
/cgN3Skxv8MgIl3cJwaeJFIqXwy+k1GpYIYrH6sWBLAClmPKUr7icBc5E9bGFL4Q
hw4IVpJXAfSkixvMcgOdUafAA1ft/tuHDlB5AKF2TW9q6TP38y61olD3Jl8ddbJS
dB/kEKk2JqAaXvcTJI9lTD0cdpMERtIICS5Ijptt0hzlqsFDJ3GqazOtsIxCaaIH
mRu2AkFcSqirrAbIXZ+AX667hY2VPf1NVj11qZl2jWLGTJpv8yxMZ9kYTpVX3Ke4
iZCXj6+epKnl5jbaZWR0mx2UVExENq8wa/7xHnHbxId85Qpa/m0agq++JVMdq2mD
4+8GLqTMZzvVvaYcKwgnxgmCOfWwfzCegOCIBZH9u/W2teHe9i3qjKNEo5nPRpwu
qNoDIbXZfrqRMF26c4pXn+DH/UK+D0GDsQWC0Ee9PnG9lujfPIlz542f5/qdd6Ly
HTJ8l1UgqMxx/Car13nW9lCFCy1zycQwGkemiMbWUeTq4aFqC+Nq7qMj9vkd8Q/p
nHZ5+BGftQiIj4xVY5/XgPCRvowShlA8y3wPpduIDYKG7VTeMOikNhFmlbBk5DoG
DSh18+BXL+Ie3C2bROpdPQRnH1T1Yer/mSKRY1cSfWWVu1GujGWeVvkJJpj0pcIx
m3mPINYho7ESHgFdBbA9W0hXvqYM+yI1D5A16MLJF+Fi33T2Mn/2wYBCVT8u82P4
EqQYsknyilo1377prM6S8sqoqfVH8vm2L8rl9/rVCuEmMSY0/7K6o57TDsbu6OFe
6IVgTa7ZqVbsE3T23VWhZDqGblkC0lsTuQMGhh+sAY5WY8apwCIno4M/4rh98unM
qYYaQI5JU0QYoKHGuu5Tofi186dZEwW/dky/LBpmOByzuip76Ozmy0IR7pkiLmcR
teqhMUeIFHVZvVjUelPM9ugJDv4tJ+2DwIbvS9L5bNj4Tt/FdLiJLFErxLpjfHqf
7laN5fjef8VqFtMocuRBxTM3iAflFIuKUgD9npmE3UQlVL11qIzH0Xn2tvWrEu5c
wq6zUPMdddcsdQmHdNGMrrzq8Xceh1L6zDVHTJHCOjUV7txTj1fuAOqhVnhwoA+r
IlAuU6N5auxCgtqtTaqfBb7qcJrDlX7L0CAAnxU9R26ldTZDVI72WUHhH9GuomqX
MXu8DkJJNMjfntQnV/kS1hORGQjP4xXhEA226uqsMCfsYK9cUcLpW2f1zv96+//e
KFo6T+bPcL88vRUngZwLuhhiZnrdqWZfYENPBjk2adpCtaxgNpV4Lf1kGuIJsdeD
TEZg+f/33rj63pc+nWulVNbTWwzUvwNZ+lmNS++NYxb+Zkx7rVxrSCLz/pspFZSb
N+Do4y130TF1L5oKsxlAtZRSntac0dZkNuvlzah7RHijpd9RIut8PIe02YYTNwPn
bYMZhhZwatrQPE6juVbKMI6O+Dix5xoDGoL4dTqs6rXQpr/UYGGY7C1aT9xnaHO5
3ZRhsv+wrBwF6HGipj5fV+pSJ5N2nDYQsei+VMoBPbvjD0LlA1jgTAsV6eLaAPiO
MbdEhM+6vZ4R+0VkicfRNeZ8LshiNlY4kHbifsbUi6rJL/ZadX1K/a+vV2ouVrvR
N2SrUIlzwp6pOue8EarOhmzhA14E7UDVKxD/c9j2AN/pNmpFdXkxKLveWceLf/rc
1sYBuwGzU+Mk21raxJh3eTh9+D9/M32hM34r08n1a0uhYcdoVzNkDYKJqkFP3Twj
2v75lpGDFmY78NtL3itXXjcfkpXxDV7A05mTniTubgN+j0ZUAaIEjTrwXfzwb2hX
8HUc31OA5DWtftyy2UGDl5L+Ogzr6Wla5xUA0VhFgDUqkfejfiezILasgktbNBUD
wMrLbI24RM2AR5xwESwErHNQXeWwSBGWcWrF6WMQLqVX/nPdh39N1iw48s6Ff/uW
6UG+u02BMI8V5R3CyFt0W/3GnT2hc+jvGyZpD/9mDwKXwHsNEMEfZ0JdlOb5CesN
hpf5iFkRSL8fkLsnWLqvcY7miCzRSSl1n3DbaOUPCgYhQx+eNPRckD6uwle0Zpf/
sb/gezfEVYTTSB+ScNfntmwiNkworA8jbDmU0hYPFI98JMHZY7K6GWWuL8ps8jyI
cjJDIAWQbkH9bizszCQa0xTzyTLUOijXbsNXyoxgLcJbfsr2yUonWywlivPVt17C
OiRX2ChkFaVM4hD6X47l6zRTn5dLt0WXzbVbZNlzR1eydU843gKhpFZtpowwtz7d
h/DWuxpcfUOeiEYudjA1u6oza4iBkN8RPARbpb9yqbA8prr0Zeeif/poenX8itVj
GrUETaxGer2iM9DHGWsytW9JT2bveYhhNd7NryDxwzeKRnoB9UNvOqWiqyH8usZ9
YlMHzUhUXqaUEH8qjD3tjLM+akpjzt6pOUxf9Ww6VPuW0BbD00tJvfMlw3O87gQk
QBsc4aSw0OD04L+B9nBRjJxy2aAtbcK6TnB9JAdS15V+u96fK9JTepbn3fQyx8kj
4oWnCsR/wiTl0FgY5TibY3itBJWSpNbEUelWplV+/1O8ssdYAX+VSBa10U4h3aoc
/CfMwIDtFGm6tTdGuJtfu8rAEJ6bKVYVgPXaALVMWzUW1XFym0E8yGWGxNZfYeCX
ynRG6YxymR8qiaiwpd550NkRdfqmr8eERMHXAQMHvhH46seqf3esUfPPxpcccabb
Oa1aE4J9GEBZ8NS/uZK6ERSRD5LVUnxLSUY+ZuygjXtfVlbzZJwkAR7ZGqFXE+YZ
EK2waZDmdhcYg1VZ+jhVgXQudosXENvC3i3n8VtS9sQnWaDSYYQrY+fGTSdA3qwC
j3znAeWgFhNHQXrgRTFi8gi5GRGsuapplH1+5Qu5jULSlbn7n4g5At3ujS26Mle6
9MbhYSTqtW+loOttmTRGcch3OO2DxRag268C3M/FoVZNi3Ko/sFEtF1mwqkXl9fY
oxOuaiLK4f+MeuN7y/BOMMhaMxpOY+AwJRVkCEp8ueuGIiU99btNd8O0JS3dnWYx
lkkD1n9E/IlGbKIkog35AcVYX8xAe2SAAWgVcZkaunfBJonTl5HppJzQ70dQldGR
8RGI1kfnsLuGPcdM4bm7vjQiD588F4pnqpFLgL6SD4RwyRGBRjhkH6J0hal+9ENl
EvunZH82kfZxSvseRBjYg+vC3YkywJsGfACx6kVksoXFQ2zNNaiqVR4WH4MmFiou
cYpgHIcLhTxz7y0QEBhsGPDiRPJzV7jh/NY7fgz4sbsFWqyPO8wPpHQtUKVlsY1H
5gb3oIk8ANKxsGCLXX503o+U8TOHKB5vC+GVRTyijC0VLkCFyQxWaToNi2PicOJ1
NvoIbZpd/oqYiBb4ZpYc5Yw745jd842KrfoSe9vkR+1UeoiDDEAM6zwS99K59Kbr
gaLFpDxgCZT8u/CFUK7GLMuM/08RZ9NZR4mkAb4GDU632tK013A9QSpb72xP2DnQ
QvwcumAbictKGh7BoLZmOBs5aOSyVVITPLhgMuZA6mupTUqEOVMTfGPzzbRYbnWS
iTL3Ee1jBeFXD5uQGQpWaLtoUPIAt/U9ORcZ89S+xifjtvepxmOC+QZuixTxmnzs
S8hTeghMzztfVqNPzoFUDuUd4jOLw9reWeV5+xevMXpWwYISylAZCHJ3/SB4UmDX
7WhPXJcr+rd3GIX+qLO1XV+jUmw9Ca8q3ZS+5Ssdxvm+142Kxvg/B6kTZDKqvYc8
MJTSDNWB3UW/muwRxPRkBp2CG8Y9Deb+DCsIjwqH+h/yubA3kNCU+lP7x5KlIMIC
jIdaHjmCobtN7e9ybMEG1Th8MB9f4AgQ4OdJhAveSlCd1dcgYHS4Z+MthUCEHX0U
rpJDfutskr09hVvpPLZRp4FrQF0n5fFh0Y4yOeKN0QiJwyWKyWuoU38nz9HrJm9m
MwxzL/sJepxtXkWBC51S/WPFAy0oUewBRDYgikyUFe1+HzRy+AaNu4YkuoaPeruX
zGf87Qtr7UKSKbr0958Pw5WxwbkLpRLaV6K08eREZFH9zV3RRm7e4xfs32omgcsd
F80HWISIdocu9D4FkDNX14amtOj25F1O6iIAzdYEo4Oqg+l0sN3x8QehB2tSOYQa
pidOsBoxtOMsHQP2s0fgWRnZ/ZKzVJdvqP+Jac9e6zn1YY56+wmodbTpIZyiiDcf
gPNrv6WNnTvuHyl+vZTNNSdGWyWRxvg/mQE3FafRNV7PNSebF916tLLpHged2yD7
4rUv4iokSf26T+sXcnIt8mozuyycMB2y0tfHU5c1+7c83qkgggD3IuN3uFCptmXd
NoYFL+O+ZAC2+qh8i1IPsonNqTxTmMTM68/ZZPnn+xmrjEw8S6oLTv9quph8cLeh
gGXsh2YLKac5Mln2QvQ0+XXwWlWl737PFlA++hFx7lNzgfXKwuE3QyFDYPOaWPqO
EtPGW2+4J8KgxADpk8er7u2WjtZQ0GqCPQNeW3nKMunbnPEWzTOPzGj4PxPQDEsJ
W5Qj8CCDQnpD8N1c5DT8a1g76kzhnly7wYKT5MZV/bTw4K+4ZgclrVdrA6Yc3kmS
jZlExJzqqdR7Dg/2DHAsiTaT0CT9Zqc2LXKGqZEFdDF2u3iNAKlcG/X7xAOEfm//
4p3MsI6iBNlyk/UUCYlPoXRTBwBk5OCWQe4f8jrKg4BP9RcDYHRVFy6+UhovxXFk
8zlsQn+IKx+eKW5zZl4kpBYOCeAafGVl9wOg03iZaAx3MUol8fiPeVbugljPv6zx
qrNk5kZkNEL7Yk4mmhU0h3unvVkBPFldvtltv1GG1u/R75fd6OB4fDBk22tJfg0s
f5Hb+0gKijyKNT2k0+TfaZkf9knOLmT5+IEC2zZmTaknSrr0JzibLO1y4Zcu92+e
DYzo4UfhHGxd2ypA7IwFErm1dPcO0knJ0fM2pieo2ksQgwR4ZqbcvzV50t7TblgU
RP8fTbQWaDzNfDVf9I+QdwKJRnCbb5QuuueYpny1RUW0ufr8aYaHS486s4dQGji4
rHr8+xAK6sZHjtAnmSUwVOMpLggYCu9uPGVQ0xaWK/rkLoyTeI/FuALqj4iznLzp
f4Ua/4ODj9TIJ2zG42YAKnmRtt3VFFI7glUQXOrF4hYBbrtth/SZf7PZK13ECR40
6lBBeo6g15iyVP6V3Dm+qPK6Bwg1gBGgYeCF0yZYDWlmtidFQzJyFkf10rVmLh9n
a/ZMWx/+wr+fFnmhU7mKbBjEJ7MiFXVfhQCDi99ZtdDJQLmo9mWtIOiP5goPBR7m
4B26b+BUipuv7x1NkdtYZlr3Z/VlY2q7SOo7zZmWAvD6kcjMxZVUyAyysgnXAbc7
1Qh3msavA1xr4xYqi/ymB6G9iIPQYetHg9SXuZoNpijSv/AVih8s+2GDL+/3ffQ7
KA0kTPyuSI1sPNa7MY1kgqgPaJDeE1DK/NRH/RkleGUums40rLFzcPakmBEnXEye
/mMoRMI89a2ElPWKWqifbZ3GB8wixnvWI2Y1rEJ1ObqYVT0a2gL5vlAXsrW73XkT
4nAOUimJ4bt4Kn+7FaELndNQ5keDcfO1iux18ujju1nv4cVqnE4tLEMFn2JTZ8aR
+PQ4HFBb/t+/9qLKUJZCJN1/Y+PeDPouqOqQbPFqsiJTluLm93ORxhdnryCXkTga
qq3QCS99zrnUCCYaa1qIdhpmMbz18Z7fL54gYfRK4c3tqWEAPmUbLZcOuw+zXYp8
i71uOZK82hqV5ASju9/truyWHpY0U24ZFn3mFjTECFTdOSgKKWlPEX/o/mDhOPUk
eTdsbQDTpMDg7Ab2Xxp+WmNbXyGgdIY6GK5pnxXwaWvEY56mHxzBe2/7E4FO4crn
gJd792hbKgkw9FKq+eBlN4t93WSqCjZ1TCdcUc04HSzHUJYMlcLsW6GkL+DnP+Fc
M3dWYjftkyQsVfEYldPH1r2RUDdIgCBveNDNvJaylFODN0KiRo3ZdSbLw1y0pepE
rHA/Wyt8SAAhLxWxLCQOtx5hWzzHpKMtXRpNtmWiTUWilEyxqRqt3S5zpotZKxuv
RbuD+szmjzfgq9xFokUtkC2zHqlDX3pFMJeRA5fYqzWW4j0EjLWeg9pw8wZLqWWn
l1oKf/VagvCYeRXiWJAZEi9GuWDWLvKeLgqDaZObX3gROhrmCmQoWs7vfWizIJEY
KOuzU/gD/DbekWOaggBKDWvocwvCgiDCAH6L68/fqBMawqG1GownZD7k6oVt0aUE
3Ymq9ADuE8rou4zQYkSx2Mgn7YJbWeLQUwdzcd5lBC2SghKmIfTGKmwyTefYIbdo
oTkfgSwmoA/Mu4o0lmxsRq/GVMqdgc+APa3ilAtb4iXeuq5unZyJeMhnFVBatYIp
lTLwqboNHS45Ajh6tj62LAJwXLikaquaqxC4rWN0WJIKCuly8brJqIg/75S5ljBw
o9jtIbCkCqzZbAWmwmhJ7j6WNq18RhWg8Ig4aO0CkaJNEHlxyqmCwqSQ8pgEKT5c
hLuEFTZfeIsPZQTKtJTkcCUvKTpoo/IApDQWN2hN3j0CBof097xpbQXR+Bvpw+Ot
/z6JO5T0n15sCP+iVtdkW60HqvLidknobJgjULUoFJ+8GUPvexu7grdPn5P9a+aj
XNcs+7YBmwfADodZVZ+Qha3pa0/pueBs/9u78glPI9/xIqSJwhmu35rRMOL+S4RU
P5srCSL4SMYURULmPcwokiBYfO9V6jkAxvPkNPd9W7KR2rC8Y6SzGEVEhzrLgjA3
9KnwIYyjF60P0NFFg2APE0nbgih7+iScgnIkPkHe9R2CAjejYzEe2NEjeDjjtTNz
+zCXytMJbssF/MU8E1L4T0e0x4Os/ke49rq/ggDUPPFkTeTB6AMjmfiapR1xdMIX
2DsC6r8jRtcHrKih/c1ucPY77b519ZUTHNmf2pRWLsvw3L08bamRnheXm3ldaFfN
KGFpIzyXCKvGAgKBGlrXEb7mkRsnKLcBdXp9fUfz5inNHeHjq0OKD+8Gq4t3Ly4m
4ZftK82xlsRn+gIuQ0LYxesPlVxrXaQlPe88BHyB/HNpffnRjXG6pgx1azK6LBwJ
RxCJ9vUff0sNTHwqOMMfBwCXWIq2dCe1BaX3zQyv6HmmpbhkZs7SMH7n9MbGhgQ6
lhBt1HetSmyYij4NYed23v8gHfM5TVEsOfuc+e8Z2QWTFNtLKisKTDNZaB3RfYKT
0U5IXyEve9C9SpR7h3WptskYb9/VdfcFmXoduML0kCvitmcxqcAB2cmC/ON1lzcE
yji3axiENBCJ5yt/XQdvuxyG1RPMXBbLEN5chh+n4MUksfP21C0UnZalICvCkeAd
EOv2BM66l/MHeK9DBFy6U/YeQQF/jZWS//gSYRrabXL40hEu3s1Bo8DTIOxjuCiv
mAdN410jQBiSSqedgF7/yIf9tmz2lwy6qZr7P4NukSj6KYyLXl7im4a18ftqVPuy
w+vlo/nXJ7gy6a16WVgkUhB2NgoMtDRlINZXS8my5Qmg8IXU3gP9pBpZdHq9XSU/
vyAF3rFl67ZmD9bJJc35w16Kae+S/PggzZLCFvDgP0QU+l0Qe47yCO8OGf6KsqKX
MPd/HOK0e8yl+PKWjYjxkM5TkT/Eo9YyzZNYBuSIRb5C3tvbeQWWHAG4M4ivcCY9
r+/0/d+6kfqEnP3H7QPofhEFtxQL9VsWJlrJDccPTjg0XMH5a/bfEfwd3VQBGMJZ
ygFI8myWubVZCRAHxwzZtSshRL4Vm8RUmXvoHt9Kwuk7puyiYqjDcSDCHIuz7XN5
Bkx5MAxKAgKieQt2H9enyXLeSP3MW9KedqzgjvXAcnShf25SzDvvOwd+J+Q5f9fq
Cq9EnaPHwFYmnSkkBT9nsEgOlo2vjpxFMSrKtr2ilvpSCoibBFI+dlPcRcDBlO8a
SmjBDzYKCfW9uren9S0SeEKCXnCUO4/E+Wjck0TaqbLgfHUyDpq2N4aOnRDAS7Cs
8Aee48J7orcjCYKP7Q5anLH23x7iEnkpY31La00bmhgLOFIkxU8gCKSm4qTAr3GD
+WgNBSek6j4FjT2YYEZ1IplPhsGaEguoyBXQYfa7a38TZpcS6AIhVDk58LNF0f6z
OK1KBkLmd6ImanbKhulexr6t7xjrospLeox/nVYH/wot+DCoTzfHWdsdsntHSHmk
ZnRmAG3DGSMjZAuyJwXL0qYW/M/6PBeQQ5meFjMMN8BS8bmWvnqFvZ/vO0iEHpMo
j4NcqtuCwCB+yPdI4umdL0rb4Tl1JLqYPwTpPrdFVrBDu5Y29psMRBv9CMtVh5QQ
ngF2tY5/mn0gHyic4WJRxz4oba/fu9jzycZmzFGPSQ1l6X1GfuN7TWOICBwkNooI
If1/vdAviHfSNILE4/VXPbnN1mQYiZmzddPL7xScAUDxPWykzYKbJo6p5S1gpArd
VhBWQg0eNEbvaCSBueGIf3V9+E0EfMOg34nU9LLvCYvBDwf9NhMnfUEY43MC6Vl2
swXV1VO/xx0kok9uqei3Y7vm/0CkGgnAH73eRkV0XjgG5lEA3EczOYsK0txiGvjK
OpOUF93+8MWbwucgRksGWOqiI6SgmVhXtQDvej8WEGiUJ+CZTJ5UEQsbMQKXDDO0
ObxaSKlc/nNymMTsfCEhTuicnrQD2enQC+GbPRh2X/HH4i5V4eGzaGBc0mn+r4SC
LeC1F3SED+N7oD0S87etXFUuR+970z0VXYDL/B5AcOwPHe+YvqX5xlZA/U3Kf0gx
oGqcdQ9V+tXGFAd5EH74Q+FdNXa6V3VhDivjApe9Rs8suYNjgVUE37l7BqEOmC6d
KU5FGMt+N0W1hVXPm0kecWNaNLeArLAAjM4D1GSfJLRJyXCwgrqph7o+BBTWv2V1
xBCTVYSVKfARBKTQo/4EiPgibifnXN2qmniXy07tiomFEIMLannqBxbDLp1Zx5Gs
f08s4HmgOPBce9Ou4zNhw5FStE19I3vsjietyhgjq00RdeT7Ie4xi1eeTDV6zzVW
BC7mC07ffhObHgGBIw86EincfBRWkVp3/dwQF+S5NF8CEKJBfzI41XEGSHHvWB8P
U+0BUk8S7f1xeH7r99K+L16KjwTFMHZP4oHKY11pptPKVldjB6LKKwzmQqEHbt2d
dhXwvFzZ7Fgs38A1a+QjrCUtMuEX+In5OTed7ZuGdCM5n4ZTIfOSqQxyVYjdyiMp
aS3Kpbi+5V+KAEm/fMcKiVifg8mOcBs2wta5VK/Vk1xSnKPO29RlbPEAgWMUymuh
HaY2X2Bqgj4RGe7/JRfS5RSV1hjFzG2oE8llQ3qYQp/R1Rke1SeQICaT6r65yYsu
UvCQBMwJKnpM797z/BkgSvcDnURi6HM3+MO43zCW6wLdxzptE9KtQnFtEHnUJxHf
ZUffmxTEdKXQlFGTcwvTQxm12zFuEhN3G0KK2Ocsx2Xv5aEoENuKtWbhn779FEul
MjGGnJcUwAS2uuJ2wo7PzwaLAC6Xe6VZ0EkiBBfnaslWKrlrnAUGRgxrJlr0ELRm
K1CgQ1bdtEWUGPjvDqDcwtDFEqoEKiSDOQ6vQ2NYxFEcSXhOkgqp583a2mojZUIS
gO3z8atOLgi6SqCfGTNl97VnnQw+bzuZ2/xkLzPgKsxqfvfMty7Zq2TBaqUfOVDM
3B483eE6N4H/TT7D9jWdzdE8wCmepi+jBUeUplCJKt4t4SEXsiDVp/7Lk9k55zmC
cgRaW7kMuX8XHuGSG2KXuIT7yOTHX+VlXY/rBMHvqjmNWE/FTdWLkuXCcYqgfExI
Wrb61ZLDqIjXEg6xvh6AeFaXtnn7mdYkTDmoRjYNTfll709nXEBcmzVxwcaP36KO
K/g7LTyQkOFABcDQMOnf+40bzLxPiPc896RFgKkXAu60LxC3BEajlmheIkaKYSYE
VYN59ougQDKQe4LwDth2B5hLlUC8YTCuxeZVpeNjoKjUeB5cDTi+s1rV/q8vJrk9
562AHYCjupzDE2UGHjf3Jq/Sra+q/EWGnZysKjqloFHUmQ50SoqFQyUo39P4YpXf
LSt+7txq7QC+cWT8NW3NxVwzkjXUehgPPap4eh2tJoe+1oWEGAZbgQjwp3BPlvcW
lIaBxLfaGANCDDahqVsCnpX9yqfPNQmyA2O93QX9ChH78opU1EElZPK57snVIh1o
LzV6UEw2j0LfhzyCVgYfVLhxUlhOvyugktDhNESsYqDFwNrxDT3tciWaI3swMkC6
Vmn2j4XQKmHL0/JjarN9RSJU22yvAr9GH84RPdYtAP7j72ZTttWqstkwO0NJBx6N
NKYw3rOVMdO/Lg+JTXWh7Po4mM6yTMehBqKiqhF9cI9bQLRR1haCAx9VdTfwzG8b
20bYJdmx3rnFHwKm1ZJeNbJf806nqIA0HlaS8EL1qGdP3UIvtwAqS1oAR+mGtHeP
AuFOT62xlsaf4vU916nh4Idc0yVVc9nO1sEJeP61HGEHyVgzty+Jdg8EASXWG+zd
fMb88qofpyeXzfn6L2F+3RpVHRzIk+hGUxvx1Pd935d94UoJIAHumnUrq3et3Uk5
6KPpTYIho0Oe/JmDI1RZgWs/b39uTLi3HC94ydd7bhFVXDyKgE7lCl0R3du/18S+
CuKC7/ZFHuGJjqAWwXHja4kzUq1JYuBgU8ylj+OiY9rsOAjX4vjz38vP3hSPMqWb
kXYDfTDSAlZQtWK3snvD0wrIJrj47VaSupM34Wq9RmRvBjjFaaG8GFl+k5b7Pqxl
sZcLoUSMoY3MxpxWuCvHCtpTkBpDIICvbIOCXRykI1poqss6Zl5fZi/bqYU25kgj
bp0dvT+ftin1LCFs+s59gvhQzMUPVArTKo+5JU/OtLTFEjVsarx6WkU+JpPC+xMX
CjDyHz0YAS5d5H+nk41X5eNUwCjuqn9+olXOVvPTZllfDZZxyChaLiXf15kZWy1z
pYxmqahUPU+ZJTq9bu1Yrg5jcrf/TIPdaRFc4EG+q80P2W9l9LTJH+55JcEpmHFw
JR4S10CxAl6p5vE1J3q2O9O96eknUN4QkQaHcvHKIkTT7R4EELm450k20Y18sgnb
dXydvo0zgYdqjonLrQ+p8i28Opp9yKUeFG6XKXCioxmqORtc/O3v9sxQFszK6b/W
6OAJhYrxT/LuFRBA9dXC9SJLT18p4zyGlAZ4D2WXvmFawVY2GlJciiVs4XLnOs2p
CcONdDdVsCRDL3wvVLLYQ3241yCGJrxeIVVSgFwP3GF1GI+rLC6jLThIqjzuhnMF
zPXmKW6b9MML0YWAEiTN3W1WUJcSty9OzReK2ibILlRK+KRW0tAyDko+kv6ZYwRw
NV8x59D4iIBDUqwOWOemRYEW2IsEX0NJCEJZn5XaWc2QKleOFbJk8wyYhLdrSLJq
5ayx83RW4H8ZarefkPzAbjFVF/CVzQS+cQ5XWpkvWOSq5k6E5v+4euFfHHyTjlJB
DIze3qVu1MWjbdAwuNh2mAZvCNcAWvLCI5asZo3RRlMgZ4ke43FKMXnbFNW6e7ZF
rhkcU+qFpL4UDtNi6w8wpF7R2ocVB5T7Yo/mXykCQEjFdWejUSviVKyLEviHdMRd
HQpkptUzAnbwv91kD0Hxoo4R1Sce9iz6vnwmQ5txW7cDBaO6M5gUk/w0KAZYYjeJ
/eNonwa+/Rl855ufRvHGH7ylZmczCIpa5k83WJYnd1/SEiMgV89sSMecpFv+aPaG
HEra2biorDs7wG478K3aXcTLn7BsYMCzA1zYGUVVrNYZai2qjE3+9/6OWdhqVV+M
SmaEKTJChL7e8AISuXJEz7g7Qh8kOxK07Y/TduFXvSGon5otaCcNf4tAYv4NAUTc
BFpe+cDYwPYQj3rWzcBcbYAhj5hwkyWV/RREowansCFxNNHCr2Tjl/wd5/3W7dhG
DU9q8RNk8V+zEt0MOq6pCgY6pbt3XPKUgEWN9/D12FLZlJXcwa5pbFOnBIKtgt55
zy7RzCx4XL0xofhgtspcbHkc1x9DVbk0s1uHHI43LaK5eotSSrAIk7Of1JvJw2z4
kbrlN0xeSYpYuLpWlTbkHqarGvFLhb8TrtYp7NUNWyzhPsCQLNeSB0CvE/3ttfgS
sjwHgCWGhTfzVa/oH+BAAooa7QdMZmgl9P18wBHg5bQpxcWTd3uIUyF2KOipNOyy
DmBnxyw5ZG1ht68bBUk78PYfptocj6uLHcG0A77EGHB9xGW2ZKbl7Ir3IPcwxjtk
/2bSCSf0QDXcKgIYMFeF7brcec5pTBPr1tRzkwaW73WLv+dTnxp93s0yH+2pwnFE
Xs9hJJuylO3l8/C6/BMxxxfXq4a50U11Gg/ALUkv2tv60XUaV3UXK3HnKowLqrM6
1NaDeYZsfRJnlZpSdzA++ukpBCXNMkVJMUeCb653efmYCTYViE7dUDgPO+O4+drN
QkZSQYrI0EN2xR+S+MXVkhaX1zkxECuJOkSM4JIAG1CY3LanP02F2wv6wh7sbyZR
w02jvInHKFyXdd6MyoLlwte16ukS71B7HfQKR+b0mhb3cQKpdd2683WwkMWKBbfC
aNJTynJUbd3VKcmP+k6fXpR0hsnKNDPtZS1b36Jy5XHZbwyx45GHFBwePR3/p7JG
LXtwOQ0ky40KZ1b1/b1VKqhj8FcaR3bKJMQyIzB80GTDAI0UqlMo0YVp8uClX/4A
aCDbGzw3roa/39pa5mNxE6dY3nCjrakiF25euWQ0AjqY1JgmIwi/3VpzNl/7v9AC
9Dlc9j0U1oaL0Mz+3fMpPDYCFXBtF+0T81y6IijxtDp2TToUhZFCmlt2hRjByu9u
K0Fhwif+x/w9AIv6R1RVCCqtuVGtrepxgyYVtIkeEMFn9ishbRYNHHTYuM9tmgFt
3LzR5AU4iqwskTgHd8slC37DvUtnXVklujdpMVfcvNsuEQ/E1F1b4r964mp+PJge
Zp+pC3GeHVs1bswbr+ieIkIky4AWI2ZcGmdDbSgTcES+CfNZiuP6bjpDu82C7HhZ
hESiImzpOaYJT8N/wQXnUb+ccTl+sum1o2I64r9opSeSIjZs7AosqK3gceqrOhAd
J0FA8BQVLLVPZWEEnOZvtR33TIr1yOUcXlru9WsKLkw51iMF08f9U5S2WzcX1mf9
K2Hp/ClUXO8I7fUExeH/DQydD2ZLL3Se56q8XxiigFKXU/XfW1uXmgF0P43SrfzQ
silGTcXcmEPkK1/Z5NV8KyEZp9GPk9e702urdX9cxQ/75pjlBiDYskNs16qmDdcx
bOpXwfUF81bTbmkyFN29jOM2tYCrVpw+6+FBL0SAdyQKsfxm7COY4T5bC0umnEgm
gtiP7WPmv+qXWUjpOA4jTCc6/NpIbat4cac0meb6kLjJTr637z7/EvRLNXpbIdA0
UvXFnz9/4wz4lOBIfDPE1nTS3KH0xSNBUH7jxQCAc2LoIy4mHiMSfa5NCkeYmVxs
yAkgVOkVZe4ZTE+vJgxIGi4k8HwLyxapZVsNwD1ag5ncwzIQAf3Hc94sBzQi4G9a
jENIVrSIEqndDzTkfQ4X+MRo9/uc/rGUihJFt4ov/x4sj9xwHfKbp0UBbYzXSjzi
hMlC/bzJrYOT8FVrSOmKrxpSEhbXB12a52j4CVOz944EAa4yLNInhdjbZIfUWJlO
Yne4QOMV3Inji+5Q+sxLOAWcb5fzE+i//fJjThGNN7m9FradvoUHh6UnoUucdRuC
E5FZWBCPXXl4X27eJmpeJOfZRllGG86zjB4kbhedsrGrqCo/S39DJz/mhtXiadoO
1vI2104s0rGgfLRy0GU7q5PxiT0Vx2H93AV517Wi7zddiQmG9tpclx3Ngj8EJFoR
8hZm3bSNOZAtc7ksViMawMetRh1vadWmR6Z76+RJVT3YEMbYr9f2y0ROrpuNvRkR
3EtOwcz9oKEuaPEm0TCQMDVYY0RM4Z7e5Uckm++fOyoDF3Jk8Ncm2mIfxePffR7n
i3e10yjbDNb/GCbIoWD+xUcynF3JJL1y5RraVTsZ68HAadgm3cSypPlUZgBk0hFO
Qm3JHPXBkPqFixy08s9Exd/71dqtihjFtqIjllSrl0mLIKUjZtvUygxYzpcWbmjq
/vGmiO3PCRj2qcujmmjOdoqAEczVoOtREgWfLQPRqeeBdy/0er3BPUwyibBUUuSN
hkjHndMIUhwa0V/8FMiEm3/zm/figzO1yGGFJHpZB0XJMZIyn7bFeMNm4VH6OZR7
qtnX2cTq958ptaBqHDb2qDkZXRc8wlZ9Cd1EznWTsdrmVs53soO2IzRTnR8sjCFC
Fm62vu2iNIaLQcXMrjgnbbsAGY0qcGFMaFmLTmNr8Drfg/FeIy8bZo02kgxB+IiF
Wn64HU1UfUpCZRsB7khXCO52fdw7PRpquglyr9orvWF/CjLFONiLEzyEruTTznd0
DUz7B3EgCZFekY1llPHqO1zBF85aBNGG8suLPxp/zXkrX/5Cv3pt+rjcVo17C6v+
CugU9NCWBzmcmhLFkNqIpULZExEj6HoUiyscl3IpXIf3D9E7reNj+wj5H+rA6n+S
1JdzaS/8LkQ/wxui7/MNw7btba/whrHyy7hz2EwD1i/LrtwDakLWebiph8jZVJCC
OgzQeMQwQlumCIHH698ydp8ReRwEI02DcFdHFjRjI7iVTinIn71bRCnKoMIskdtI
7fYZhItmMGfOdcHMkHi3+pufAVPodrtrpXUAqscHE2BdQgKBgoy3/qxsFflE+ODi
wLKyeMqwEcpZFT7K/U/C+oMuk0kcuaHqKgKg+aDkKlTdzfO7JOuF5aVFbsd8HyVs
pNYFi5g7i+FBAtt5PBoyMh79V1jTGMBlzu1qkNlzBHGm8mLjVeSoSxanvkKVHDjr
cjwLmcWYCB9ez7dee8XnUtuUa+JXpgzM364z/IF/fl8wsUR7+VJyARN+qjfr6zeE
FUhCjfizlt266Pog0fICkIzO3zLuBRnkvjEatrFGgW876axFWjY7zpELgr7ZEKRd
IHNZMO/pxaIsEmEGlLe4l2U3UWER3YlbHnTmJhWCyDvsatWPpuML/bJVBWSND7YB
N2EorLYwhURPJ1K2wG4tNSzXs6ZAalGW5I0JG3f01xCa1Bf4VTynsOFisWE9ULnx
aYdoWq2jd+44E8/XU5gkXonG4x9Hdz0vPrPPbjEqvZPfQCH9nPE5uoo3rFzlrdq8
vzoNgRyAX7OeuHiTgP8cKs4J0vpzgijElxgc6menCqp1g+qqlNVX2iK72J8TVCNJ
2q7XyiRluWIWV4fAswa4mnTVoulUSFOMPXZsEaTITqQ2QVSp0gUW8Bm3IizPPvgi
IZJrOO56AfRc5byL+U6dK+Xvp/fAeS+mwT4S+udyL5/axqf1a8mbeD2+LthJxMBh
hbwM1LjkOXgRAWVzzqSgsl00F8BSNj5oFz+ge/qFjUAMbAhwFfYA04u8Z0NunhSp
x9YhqSVtM3s7Cjz4JO8KD+ihPACdH+zhwkjntEO8ImB0tHxkWPwB1m/fNGW/lESJ
a51YiMyst63EVHLSUKID+J0KiEADiMcbvv9n2frlG8B9TFcPLDuZsCz7tQ0siS3m
swx+XYHHbhTFCDHsNbWgiQXLmnwgpCy+ymWQUO4VUU/N2JaJqHWkI6PkjWBRRLiv
u+P7dfKvAuKc30fe6CBsiAFVE0I20xLsgdmra93Ld/hnpZR5SkiuGgkskxT1HSrU
FclNe3I4znacPmCpuy1o0y7tcb45FK+7LxW2aqaFVGjcR3ICyXmuRf3kFXMQpH+4
BxQzWh44foFrMPWL4ShsYEUrx0NrweOWCf7p5xQ+CT8OYUBvJpkgSEoeZvYqz0ZV
oBVL8auVl6rUd65sIwdEqr8w4OniTtq21N84aD3n/2vbjVeha3NSClTKr9xj70Se
VegszA0kSBXVP2bwQZAD7GmujtxjNOFydhaNjFH7vtVXXK4gvNlE7STHraxkvJxr
EdenFRIBYGYdmOhgD7AMii6jb2/LecAgvn5wZSDYy7iPv71H2sK+MpVcoyn3Z0pZ
u52wMsyhdpilsfGn6XSD+JfR9Kp+MTah+2CK8gd6vDfan97cKsyrmPXByeFPLftF
ieRm0f/jCsitGo+i4VM5SltO2mlSfCeMwbC6QfT4z6CpiBmlc58NSdRU0853/a9J
j6Y3uT9tUJB2hnX69zPbX7y3mW48QDaeml1EzlOwsaYND41SpxVrqSauEjnl8m5y
QoLHUPOWc/0TkERbKrlDbmPvitVbJOXMwZsMymYQWF0ELK3kugeBnX4Ar38JcfbN
9gYo5tyUQPrN4nzgMLINOmnnbxjcIQfkOIrfJz8s1EaV+gjwNxhNpG6qx1Wl6I4Z
tdfXoijgzhPdQTsRqxNB3BJLAzYwvZiclyvHw2+woIDVX6C1hIVghyecM+K4PDwZ
VyZXOaS3M6ZVbdkZpa/lM051etvKcY+KgXsn0A2uEmbLwJB21ruNoNSBYq7sO7Sk
UAPpuu+i2LtdF/lJHD89/YRsWVXMje10nNAJh6lxSENg1n8F+x2tICjncVlaD9Vn
nsd6iBUiTJ+Te5nG0ACKgqRR9zf32gPjaVbpRSvBrXAinNYkIxHApBJFDVX2pCKU
BO3lx9LW8W8dc5UOBkgq/7Q1OYnY/opriWr6mg6D06T6unGifTVh9S605JyLUqU0
s6VB+eNsAJSqM5saMJFAyWA4TvM130JVbxCWFCtuzteYdvXZUH5ec4HPSoep+F23
ZHMBfFvFrcOafJjYcr2f93AbaK9OFWlJ2TmIcCZMoFGyW2+n1vynOtO9aXakOrUu
UH5AIWR1X388KUVHI9VJ2CfjWrGfDn6OqHW4VJjbB2X10EIoZpwAVMcEWL4+5IOo
shsXNAa+4ZJV9JNPNK0xTomBlIw7XcpojAkwNdLfVtJVHwC5l8pwAAgyI2kqSDiR
qI+2S6+DVWpUV9MrN0ZXTq3UmMs4txKYGh49I3JoRyNg+i1O8vyRnepzuy6+1qbg
Cf6ZlxmhyUhBk2iJaICt65jhQRNSkSAiiR4ibTIXq6DsJIBYxlS6yCqLums84Qd9
IubprmaI/AFClyB+PpENejHbtWol/8Q6ZCvJsqWXpJT7p+VTbY6NtWsomXOUB/IF
swzNyoD5WUOAR1Iw+7gaGOIFqe05+RlkSEG9m75ioL/tt+qydg+URGGWZy9kMgvf
Zq/hO4E+YWBKRJJ99e6aEGNXwxQ3yX6DHe0tvVvAQCIqQGdVDqZRMSeV8QHf0pc9
bK86HTH9r7QaDySIML3VT4GZQDWhQPQB+xCVt6u6jpff2QCuiGhto6Na+MHU5emh
aGFzieUT+JFW9ZDVFmrzd3xoYAlCzovqRrBFQgg5HdcUBvFbFxVOQIXIoMcL1963
ODF12x8shg4SpVoeVXuRwxtcqZm+J7YIdkIcj1VbbymFgYjZONW+W/7mU0bDkf1s
ff3EITCwtcpEmjPuKi75Q6+QdBIumbLkIZG5G6eQWilWEHQc9+mOtjE5YN2J+vzM
NaShXUJSQK/8YciyqDYLX0oqNGXiwTQdU2GERS0FRmqeXeIHb1wCrZ5kfQDXXCX4
TMUoC3DFflVnOXzGDIfCF9KXsC1o6redphde4nKxsq8eSe9nnofHcu0gXFbNQv+l
I/A1eKcmvOcrNrnS7KQzL0tUSHAc4m/nxwCYmxrDWw3XcGU8Pio1kmBuqTJrezQc
ct9M+gJLbrzMreyAAkv/F9XbU+IUi23pYwRm3v2fi64JNARzN3khV9grufjL8qJx
oWcN02vF+JIGkKaCLq6ao2c/rVLEM56/zy0LYqLei5cCQRsZMeETrJ53g60vHnHf
WaP81cwjJmEhoOI87Kr8xROwgO3zCu4aAvS6Z4D0jtBajTn876pKT1kUI/rrTrn9
i/QVqu2srCoSEc88JUTeTKEkOi1dTrv/Xg/dS+WYwcx+1sZsfCSaTGQIvo9WKONX
soHwkPG6cHmZPB5fEgS1X1boZR+zcwXPtc+q/cFwfM3Q/LtrEkEel19uVpa9nawT
Z8ODn6sqShpXsJux88OGEP7rRwc2iRDUmlj+DdftCjwxEAX+VVjoaojuyw0VNMNe
NE3L6MmDiGrS7qMg7tz5Fw+wrLwzqD1x3khl8GmchuLhmJkqbCcDsmvu+86GDMSR
Vb3Nr3W3KpuMfJZv/KaeBkIY/8uerhqRs9bu6BOwBA5SQLd0ACEcH4tXy5b1msJh
WXToWOi/gUdr3PEPdnp+rTKyokIxrhMB46CXjsFoCaCyqvVsFjH4g9FWxIj1rpRN
q0FkmsldtUQsI+gpoIggV8YO9ZtR6jqIzdooo2H+fKs7Zp2voRWusFXrbuq77FrM
EVD6unm8NJILWZxYYRzSP8SYfa/8FupffaPwNNZyXTJKhLESNNNIkrxRN1rKowLq
JoXqAQzcCyzNpQVoG6pVHHsputza0HgU4tVO1ZAC54gKruZc/M3IRl3b0mX0FepL
J9u/Z9+zdi/QzPm9/H3kG+4+cAlOIn2JIarvZKpLVd5obDlImAxo74fZ1uq9lJ7M
goz8B1aAbleHN6Ak94zDApBuwVx3AveTCTEZi23ovWN0acOTMjeli6PDfeK2ulaT
yyRKein0SWnCTd5U+F/V/LbqK3rGJm63mmAO8TE4LAEICLcfQkQr8vwH5rK7edPQ
CVNjo+OMCuuex2pQQEUsIzHJNu63R7AKdpHtfbaJrRAUzPnnM/Octx9Lb65/I4k4
mPlUj4Kn51ArxpMMIxIBLblJqmZ9NpN5+8Ydyjj952zgl+BeHOLOK3L4AQwBz2v+
uI+T+eU4kxvMvvXl6CYxE2KAB0LOSK3LwC9DeAuGSpNFSlx9TzYRancEhxeSADdw
gCdj5kyfxIUzYceGwYZrtWE7oALxmZEEhM6Sr+XU4x0bdqbX+vu0STtcvvnfTEKt
pEk5vGy7y5JymN88X/nJa9mROXj+Eipdj6Lxa9gYBANGx7Tkgivrp1OVEYIDV+uf
jsUbk2FNyVvLEhgrAE+L2Dhbwrhv6KxLwbGJYuo3bYBQWO3pbl5FJ5sFDs5DBeY8
m5ldoNluAaFNAgVeH+Zs8EnCyL3yUokvRtMzCqfzR4leHr9gtd8RplEyToCtyXZf
z90udWZYYyRphGEEauMY96pJd7cOq9otrMC3u8t5Iksj/rQz6jE519jnprh4qli0
rLs2+bJl6/kSlmz2/mVh2NRWbqZ2HWpG1HC4y4FigpizscAbHKPi27HtVaNcPvZ2
PGtijTbKPzQVOSZSvtzFlAW+1ksYfUYLxAJciY+/RM9twKokWo+/8Vj7Jsnb+NC3
8bVpPLvcxpVnwRrVfiMixmcbB2grHE6wUdzpfmqUfBb38DZ7QqARkbnc85LyCCmZ
rVflZ7U5N59Xmmi+65YI3WydCEDVEJUyFI4nH6839UNf3a1yOYYT4oNzSSJpMhWd
eo3ULeb579Bqhpk/1/+fX66zVVOROzDdiNh2fQ6/GiGp/7eGnW8wYCDig/az17YM
8yz53nk6Kkm9MRgIsQyED9ZdmVf40uZxFH+yKv5i+kNNMIjLh4H8Zk5yW4ErwiDF
MswcdRayfGRblIxQfjkomiawdUx3XUiNajlKQmOmxZimXxud8VP5BvOTNg+D3VxA
/oJ8XSBbuL6KaE1KkFDMW+Db6GBgBiCfCBBO9kry9U0HI/x3yXlWGthf1Sdl8hyt
+oUI8sntXS8Jayea+N4gl2oxJfcHHlFHBfelowSzCpeoIl4my3yEwTCGUK8eLbii
xfdSqJaRw/tt++uJFAwxo92m1rAt5Y2Qctcrr88x0hE8TQ4a2lRhVDEQD01SFhtM
a5zJW9ugkg4vr7H7LM4KVt81suxf4g70CxDo5xAvAVSKdhLCzHUdsMk5qOmt8gcB
V80cNIvT0Vuwtq4qwQVGfzjIAOyI8TRD9GmNtDejMlBAgM1cVoKNc3wIHudIRc91
HGsDzecg3kQjqQ4rDj9dqac+0NCgUxfYSDP7NwB9NgnhCW2BbyYYkYR9e32mf/ah
0AURSQ4stbAb8guOJYSVTsJncqo88zXV98XLxAl7WndcOZaPzQb/AS8W3ernLmfb
VIKMhNdF7a74nT3/H/cRopSKb7dnf6IYGEmKxQjIX2uPb7T7fFItGAMxAz7sXtvJ
THpJZknwGCPx9qtp7VqvHpozDSBvmcl+uuPwUWpFov/LhaCIu3zv3rS/FhKhopgz
OUlUD42TPe2r6/oOzKIi5eFtDdGiP0wJua2yGCrqcBolhIxzdsjiOVHkUXCR4JJZ
A0LB/zz/+fCRbwIoUzPbzGQIG8XrwUoZZzYhcUi+Mcttj6JWhsVOG/Cid9pyuhdE
jlozCW3sGD6q6iLnexXuSECVHZx9zHSnEJS5MnTZEfSZDQ3Mu49WB8rFsTMDplvk
1tBZE2Tn9ijEIJt0ukodAOhpdiBH+JkmdNQZ0EuwmWmlfZPI4uBsJVR+Ah5TCIaJ
4tqCzYXnudPMD4bYRbMz/6sWUxqKFad5gPVgV/Xu0kz8Fd/uKWp6wnoSyKOz3bQU
KtPSCKNZk/gswhR/qSjqoydgIdapa6fjK2WsW9ZEyCE2Ubsi54kxQfo5QEt4QyJb
cG0M08yYrw96Xxvogd8giJlLMTBzUpGxq/d4drUkJkmx6vqBW+K7ZcXiwREkBYWr
DJ3W+rADwcH9LCfB6mBx5oBPvGWuN6bIFnv4GH0NJWTd/CMx7RQXSyCcOmborIyG
V58GH2MmRvBf1Zfbrq/HXGi17Y7c7WUIQpmOO4l0sVHlZIHQa+TBsMQmirBjwvMt
B31n5C009nQhjeQbtsCfHDG8t9Sh2FgK3biny0wwIwRr8/zNv3TqT/9DHxd6K+0r
nON1QdpIfT1fZqq5ui3I+qgd788wJFzx1NNWAF0QcoA+hPtuEeL08znAcNb4fNfB
MtbK1Xa+btbKRGo/TqinylHjjPDNohM7VW2sHXOExBm0RyTm3Fp0hKSa+RCz3v/C
Y2QqailwpULViNAjjoXCb2xtVgvSBmevT5zuEoyzhcuyVrj0xFQann9HKFt2em4z
ohaj4ea3Z5V0IZih1/8u5MoKTPEbHwbiwL+sGS/TQNmkaVVicF6pQuyA0ywlm1Cn
6GM0NltDH5avQ+BVGS3mts5z3DpDAiTWFw92HRyOpBXFkOe//F+vDDiwLnFj/fxW
BoSXEtPaS2eqh7NN98hBstpEMEo0xwJdSejgyUBQaQSpwZpzX2l9F9e8HuQPbRAU
XUeCug5EIenlWTMD5ITxBCKGQ+kId7XurRu0wthh3xH5cXhN6JzUH/M/PEEJXEXt
Jcf0IRXbMlrfJoeMlkFmw8ttEGYcniTygAapn8G02SJHLyMVF3cr/PILKj6UHL1A
TNW1b2ZYt7udJfpD8xZMWy2wDkM9PovsH2KHiMriwRGuJpbm7U0c1UW0tYoa+Kas
EtWZ+oANT3vJ3IPQ/C4DRdjMT/R6dZKlotkCldTtYl+DN90wcjackp9kxLuZOrVD
jVS6yGCNNU8t1sLg3uhinHYD7kYvyT5BIWjRMSHAGlvIH9tkcW/gKJYBZxufGSqx
ZDW4iIKPwvwtd8uUSRTw68elU5zoX2fqlrIpBJimH8mCVqMTP4yRq/DK+grv3tnl
oKLA4Yh0alxbd4OsaXpRtLwdWMM5MA1TxVX2BkiYiRqJ0RLokVeP2Rygy1z4eCsd
wYep72GKwi6GNvg7SqPB0qEwhzfuGEdTe9GAMoypw+zlNyGs9WGxkTsd/B+N9CvM
uOwuEKm5h2xGHqllsgVWmbIBLB3zuKpCZN+7m0jMPj5ZU2IHlw8cFLE9tyAhDp8I
NwF8V9LYFgMSLdwF7VjR4bf4YBMgdG0DiJ1I5i/sxhItl2YNRN27TFB2RTEMOQMY
6y7vsL5mjWce1J1tNQeKMkUYH3DuWRG6F1VV4dbAXkxIHTQLkj8cIC3qcOrMqLnq
/u/EPzXp6gKJT0hlV7wb/6uGihrjy/CUf5z7DGvxih3xM0RrwmYhxRbXM3yNAKNU
p5gHuRn4S2gFKura1iXx7Ci89mhv8CIS2UCUdIFWsZw0Y7OC265m5YmbsVchhD4S
iEIwS44eozbuwqBXsfQuFS6K1urbtOH9u9iHB8oEMOSBmpvGwOpQLA4hh1sguw3M
72EYmopehWUD57hT1vz4PZ8j9Xzqw29TR7HgJ9ovHhO5Y1yJOrT0gcgapCL1tz6u
eX3IlNrdWyORENq4Hta6b2gWhT3hd90BGEhTAPRw+kfImSmeFXyK7c8KdOEe22kj
5k8Wf0nWvy90gN9qaZcOYlMQpsAgNAFS+ZvrURfkREV28vlXSsb8iXkvwPbf3kUO
9J3kW2TBpKT3WmAPRU2HtiDxySCkC/WAMTKAXj+Am+3yKbgMXad3g1/a3gw//aZs
ykb3r9Nlx0Zj3fAOTZaKmMin612BTiaz7z2P6L+aEQIdL999TZBrLthHbXMUEcLZ
uXfD66aXF0ijpvHs9Ws3dNNnuI0gEWqdCm0ShuZxnvlYU08MZ50oI57zX5TekRXR
F+XHImr3k837cZpqdiWQqwTRhFE1BzEB4CdARprUWFn1q5Du0E/V9kqfel4MmQHW
Nmow7j55sJmTFKUdMfYmT1SVhjnfm0N6fu+5SUujB3aHnia6bG2M+LlZtleENQbj
Xc+OC6b0+2p1FY6u2SNxfiK61cDcgkpIUjlcefpBWl/+mqBr2W5xpPeB+Ac4Twyg
S4CSDmoaYs78CYJwslxMFhMie11/fa1hrWhXVGZ751hCgAN5s3Bl5yZ8vrxKimOG
z3ZRVaPMNIZBI5D7P4IygrF7G0R7bTmhWTx5/R3IXJoZ/mhDmzTF76Z7NhlvCcTd
dRJ+JQm5Gvif2pmyHBNiiyRcoOADj4ab9s8HBQNlHxjWM8WLQny+3GM9AjOHRNu3
zIn+iFTtS8eczXoD35lmQ11ISnR/WDxs2p4w0mEpPh0qNK75JwHU6UB0aEroOBiL
ilXwnai9G8MyD7q33XG1CGYz8ys1EcHF2MaXFJcY1tfGYjOUByAa5VDeufQ4Moms
NH2tUVVCqtA1aOpwTd5r8l/WDXABmQEuZzs91S6t1Nnzo5LX2ypEAvFYFWJJdyDx
1dYT9cGBeXpwxWmmJUwgmRj5g9phJmLvjNRJ6XWmI7pPiIy5KpGYRe5dQ+OiLHpq
2sehFkw7axQE0dyhHuBZMcFKHJ3LglX98XyLSNPzzieeOzR7wgN5zsKnNRKFz6Or
RzpBEUPLPSyscrhRTqKB61NykVsCVN52Y6HBhU6O3D4tUKMUzwwt5hvkz54J7wbU
8G64I2aszi7rjxjVdzcYrDxkDCrihfcT6U9U7qCAgrVuFyDYAWJy5gqcX3tVV1mz
4vsXhN0xonhIOrlrLrLmi8TU6OpAHCuNwBrOlc9izTXBd0hECtEIuewP8dw3A/u/
psJmEMqorvnysDEsQnf7zgExmATa0y+FdwNGLkyMl3mvfKLwZCgjBZ7bd+BEdR7Y
yECn1GbWrjVooyg2P37NhoUXUBKby3Of0brq1YbtGBH6f08TK2JdlMbZVC80SfpP
lz8qFJb6URlVI9OYp3GLTnRjSPRmlcJd62qmnJpg7d8F0CVXVqFNDe+Ccp6vpKxZ
uZ0F+zIRIuX9T2T7QpbHt0sORTlHcWEnTusGXhC9yKXVwhoI7J/D7Se2UTa3vw0C
5VG9PnbHD/0yW1seZ+yNCOCFkm7g69i020vQdNqMLkUnaGka5DTQMOwOrEUOVoa3
Oy/T3yeZcPOaZrxjcG2YDno1Uw+GXNc1OyxRRpa7w06ow7Ssdasg2BZNtlRod+fe
cnlYmn9XyVRQ6zhzNot5iEVv4D/1ULJt02bQSNnD6NxEE0ijcumgWi+AgJnLHqwr
99yw3zm187b5/S9Z9hDlXIUU4Fre677kvM5VoYzOzaKleew2blE8EBnPezjwufsq
yxqMI+4Sv680i6RrK/vFcuhBnPdUYYxGtDlIF4UBX7v+4W2DVMR4PEF4YqK3uqNV
9JiuT2JxkxL0zT7JUMcX2jVl2ELie97CJ1p/tmrtKZnLzcXhbDximYZmWuJuA5SM
UnVqwB9aHOQtXu3fROCaEwsDzj6BRKbhl7y7fmBQwA70barOxw0bTO+76ziGmio6
vLOIXnW39boiMrN1ne268LaemxhT+Sscb/7JqYYXCZwTUhMHjFaQAce48U/WuTKl
YQwYYjgiV5vHCfhiE3Hmjm5x1XZccP5M1UUtXnFgYd5ep7E9P33FqvVYZDCphBQx
gDw8oXq1QxdMszE/A044UqSa+4jthVwzYjWz+2yG4v+tVRP/AGW7eTTO0dnUX0/H
B/aB74bweX+x+TewscA8TLALdGveSS9ZVC0q6h1jPRh2eVhBacrPJSz+o93+EUA2
zi0k6o/er2k2c1R/2izT5xcxZIIpYO/hdvENPy6gSwMm9Tbbhe+oBPNBwAT+fk2R
NsWJwzaqhMgx3tXZBjBGWMakFet2mB/kLeEmhv7Wvtn7PCQqXK9i/Ez3qrnRVKWd
3o+fdlly2BWxjIUGNgRotslmuLXIhRT3+YcyKeSupIFZW+jMDjv+s70F/jypcB61
4i/pw8RnaBd+G/tBTlcFrr6jha6l84EivEICK3oE2E8jwMbKu/SRvSKaajJ/kEuk
k8aT5cNtVBs6Z/Us7ileOdnqbkjKplQpHXRBDCN/3eBRS/cAI7LaoGeyGBfoSsHj
GgLILKo70QmVwZjEeyX6T6ZR8/BWCoYMcpLzbn7e8e6eosBVeuvsO86Cd6aPT0PS
XxID9TwJYcODugZhiKjY1A9Ifx10AhSOfmD57CHaOt9PUwgADJ4/6iYJpt/nnt3Q
6RAQCG5pq7ZFj8CkuFrLa2sii7auaMHkVtjZa3gh6CjMMTvmARlNad9HHSB4QVwD
ZHA7SHYexAwYAqV+QAsk6IL+L4uz+DX6OxGN5WdZ23M89nivrERhSqF6rh/Ui+wi
VxsdfufAaAfDfW5lDN1SOepBZ69tEvae99Few7S0kIM4xeyX4VtLGwS+QfAVs3Y+
KMHqp4yKGOSZZg61w8L+NKWg6Yx2CLxvbDVPSPMU+0Wx69qgBIZHgajV90k/BoM2
PXJI8M4pf6OHoGeuKM+JqjSXhwDTXF9UWA4YHfBbo2hqczlRd3qyHcL2gOfCtabK
x4Nnj0ssZzEvy4KCHS9Uvc9mobQB7f6pvosnjAxa17ThV45pIHbOW0iADy3y0Se3
7HhvAzue3EUWmzoNUwFM0rFSbFMHJnLQWNtusX73XwaNb2Ka/o0shBUX6SS/N3CO
Zut0h4Hffvr9aPFTd+4UYVBfortkvfLAzMEna0EPFBbSp6IB/nZUgtjMnLhoeAZ4
ESbVHU2Cl+IXW3UAV/reJpWXNy6uVZvAXjiOAz/LzIJjHfEFUD8JJ3ejBoEtCOtE
WO1Qsyrmbm6o9KgjxmVsTgIc2bjcvS3iiZRKS6qXq+DqElvcPjSzQvgWUxYWaTDJ
kkCjt9aU0STxU6dYGhUYTMyK/616scCHhThjlElBX2lV18XZS2lS3Zi0gK4HcVeZ
i4EUgN8JPKMQOVXEQWQjnJt3aq3LP02R4H5sfeiqdB/PtGMAfWhLPfcFp7E9LqxQ
xOuwXetNsvGUTsMi8UDFmVB2Ek5aSaTmJP4JcE5IfVEY1QeBmy6TEvFr4UUX1npX
H0MdwQ4+q6xEDhyQe86T5rzTqQKLst/okr/2HVSXGDxaTELq1+8qDfYwkbhjR9KF
JlcABkRrBWhONEdGqcE/F2gqvjzNwcvyZwXOtv56PYfY8GE6+EwFomzDHIs28yQS
vY6b+tU9y/Aev+Il22AfxHAcoAweiD+8haxu64mPblcT39XcGIZDbD30I6p4Q3/F
YkVmGq+rtIDxJK6VEpxaXcLsDSRZpvVXvhriz5UO+hgC8EvUjEPkDJmL4t/k7lEg
lhpXZDZUJNghFBZcVG+lUuAyv7q+ILAUyVqTo5sUJrq86GH5aJfNItVWfJEeiTBc
Umz2xr9Q4QNmWhxqOp0tbk9hR5ov5PcbJSP0GuTKuUzYKUzWHnekCbIYx6+NuNWy
fjeY836zt9WjsWo6qqk2UbZmSscRYTpjaYkCewv+T4ilP1oUcHagES1uJfAzV+mv
IuQejwUPKiRsiEG6cejelKsyWBLVb3QliQw1Nhn639F9hG2bSs0iaWDRbXrfI8h+
d6fWXKJPcuPB6s0rxB6u48WCNWiYOMABJEajQUWkdKm5ynCdZNNNJheMl7ehBeHP
Ixl+e8c7/IWTuw7V+HLIleT2TbjLi+Ve0eWUH5aVLdOBkw8FfVMQc0kMMEcFOVNd
rj2Phi1w2kAXG7ukyEg8rfI1L8zs13eKsLEUnUbNcN7Ii0iAWw3FnUREfWuxDuz4
FP01ABsFJ2Oe5cBBdwgItp7csjT1pBQdB0vdjqhdyHFDi8yUnxOmQUU5CtNvSOQZ
L+TnUPFBAZZPqsRxBTcprxsVa3i+XILP+D4NRpiKHJaO8wuyP4MvK6sglqAdZOW/
NLr1bC4S6l9o5/or5hE/L25/Ac5WR3nyV3sDHWvrNYhSiSWKSSm4ycNGquF/eniU
kLcWxCDnpPEhz4eJOqJjmqSiXnKpBdXWhQPTDRBw4sd1NE+UpBppf1xXBoGMDcJs
Ig4YBezwwJv9J+pqfTfsSY44LYsLBR2M2TDkbA2AXnls5f9JvZebpx0SQlFeK6H7
Wr+AuAF+jYg75yzm+UJDqorAVAcoWKjTglYhr6O9LRxwtuvugfg0TG+mWwBV66vT
4EIEcq+M0Zvo8A/Hbr0xnaAbqqOADoOMdCJi5mKStKdZDremUDA9hYu/cJ/IRGIK
tk2gnG50s3C1eW74UX954Tyu8eEjW7cBri11D8+mchNd3MF/Keob7pN2BImAtcSV
E4b+WlSeZ1G7T93ETDduzFItMey7JeEfk1GMhiHBlB65komnqBu0XKIVfuDjDJiC
nRfN4yk068RlMo+l+gE3SMDdZ22l7qzO+DwpDtuf3i9PNoDKw0iGRBl1Q/O0oBwf
5p4luSJhRCHXaTWWc0HDDMYoi0Izrof1Txtmwi/V+qLiEYBiIQnZEKDUqwTfXGcx
YdBLAJdrzHLiXIP77nYGF1K58AT89SKdMg1Iy11E+y1lRbnt4vztHjfe0G7KttWk
njuEJyK6sCm5Ka1QGS+48i41sBpfHRVua4bHrBNFwOYXZ+NsAI4m7Bb1ZOb3t7vs
AeAZ80lATZ1/blqP2Se1HwlVahMFt/x1RuvPJEREsqI97pRYc7w4v0vGMe1ojyWW
4avl+BHFP+KZ2ieJb+HDYMRORlFYqGBaYNV2lEIYF8tVeitnD7jGTdc8OYApv666
brBVdyge0PeAY2eWgfiku62Ji3lBQ4aFg4KqYXFnz+EvLRw2EBRJ78SWB/vF4GN6
2K7vGqlRZwa7lJ/6pr69I3YEoayEeR4reP+POKe2pYfMJpJvoKujgAxoL41XJDAv
l6IWluw9ODOvEEMhL3HI3Lwk8nW2XunJ0Fd+mSXf8V+U87CTdhmN84jqT60obwEb
Bw6Zj79XCHHActYAhgf2DD+khs3pT3tOs5F0VMKEo2PXbqzzxty9Qtyn5ahYMwSG
+1+ofPlf1xNx7bLCpOXwA58ZkjRg6P3N8pV5Ao+BTPX/FfZpqv7IbR4EC7dGFhVm
zjXzl06TVFEb1l1rfcrHrSsLNAbmOcLmBdurac/NDO3KmlYzbUAlII36v+ufGFR2
adKfLbkDV6arfIsdLmwfKwSqNO55J7IbSDsBD7mZmuPZNMvh0s3Wb8U85PwHpktr
uUMzGA7YQZtZWpohpa2lrQziB0WrqcXoe/AUapjEtsYO+UW6uRGdR2H0noxKKdCk
nQMytPpRkeRaTyKb8dCAhRir4FfavhLMLz1rA/yAVcww8yQTvmixounh8S777mer
T7soXtAdQiPRgQbHbB6RFhO960QpSGDcolVBVG1bgIJ87GLV/FwKkE5eEsCX1HIn
VJ9mKd2HRmhqaPinR/herUmBI6wwVgHU5NqQ3jrK1F+ASjyyL3btMLh1579+/dhN
wuRrmZzlhZtNTPeZAM02EkrX6VjvqoovPH/lEVSNPd7hgw0hPuIy3zQWNfdI8qFs
82XDZe7kkSD3UYfTBArNWKNTRyldZ1fc+nPPZmeJTxc0UxrC7xlAbgpvjTFB81hr
N0u4gF0nV9pFBwQxIRjUGjlURVqHmhZYmGijOIrts5BUYMArt9VP7RkuU+czliCz
rEfN3ygWvvqJwtP7PmTANTud9K2+NHOXN1y3I8UyVybWJy60xl2fjD/0KfHKYquK
PdJTIak5qSSVEQzjI3ssQOFIB+kNpqH+siZNMOY/c8oHpt/s3WIzQRQ3hGtOWvcE
CPlMYXQodIl0ySXV5fl9civlgSmJ6L10HxUiX4VAcYzX78oe1b1F54COVvs/tw+9
kRY0PbmdeHydEVZQst+AzcA6gxQtahdm6DTsniLFnSEX04k2Vyb6xgWoKh2CSzIX
1OTBx4SmtkgE1vbojjnzzZwP4smUSgB3ihUqervgfm7I6y8ngsIgUutgeoohRYza
RTzpNx7Rg7woVR2qMI/fKW+53pTB4+Lbz8lyIvGF5aKaBuXoObf4RZrlmTrZLOmF
upP98h6Gm+lqp7vmvHSCEqZIZarbTyABOK9KSZPnCOKqp6pkefsXiZj7pqwQiFWJ
ko3+uBRXapZKo2AGtjJdWQn494ggGj5qhCTCKDySfn3i3O5a5r2ah1lmQMFFT4gc
oaDWuNzZcHtJqRRxtAcjyD/NdM8UYZhRxUJq9MZWHc5ZDIW+lG/Y0SBsT/DvZKCl
w0Hq5QuWaiGcsV77AZ2BM1I7ZAKiRrmKLaRtwiYPRhoJcRaz53r2teUt3SlzTjjw
5J9dqmUfpVcGFuttSmWrpLpIHXFCY41BITUQs5ycblTttEaIX8nh6QMTJ0QwPgxe
tLCwsoRoGPkIeqXrdyjpk0mbtC56W7mDRj1Xk2CMAyMI5720UmCddJAy4ft3hRpc
TICR1ZsrN/z5MAflcY4kEli7s8eupl/+sUWphYORb92Lm16G6tpgyO8FsMNtPWe4
ThoGEIUGgpaQfEbrhHJlBQxf4VyBw8pGX9JkPyUx/rXvCxnsaKLDH5aKDS0+AGeJ
Fmt/rqFmVmuqDaHjH8ltXoAQ5IGj3ZWML71NSII6ySMDD3WZuEfxhN5xI/zKNosB
R8zU89l0twWht/w1f04mSGYoXrmQJOIQyKBrbbUKmGeYM3Ihe0qiNuKTA2yLVcvl
Xt8dNjjShAyr2TBH0qsW7Vl3o1riaqhQSTKFPHZ5GfARmbUd9up6oAkv3vo2VRPd
i5QfJdl3Hj/Zlabhu6Zi9MBjh7XWQYCb8Wxf2ggtlJAAb0c3zC+aDLNKok44Idm3
1Wa2Qi5d8B+8qLbUTA7s5Lxy2eAlqsXmib3eXyBz/bG1ZO97FHA4htpepq2RCk9H
3aKVFeG6KW4IIJ3S8wwJ9zPTx59/m0ZqjTfTzIM0paOuk+lCyLWWsRB2GBiCe842
3d0v8IBzlAxWCSHNXdMXr+n396ohz8A/RZaM95Z9JcLLsFT8I7+l35C1WufwTbON
OL+GhZbWfAesCd22BscNUdAt/CfVyCIVi+yWcHHtM5DB79GdJcuxUHowG83TGoYC
xyk+nNYZfOtoJttV4l16MTM/FDciIIKefTD/lGFOjwggk1DyncUQmiG9YITnqjAE
OHXUD4adJsqnBS3yz7joldna47BUhy3KT0kaxtiyehjZU/KLdvlMDRygxLpDpKAx
RO2sjuIyrV6+hEypcKB9RAKJtQ2WSGcSy79iMzRvtAlxIJSXuEUCpG7pHe2pxN6K
Me/mV5x4pCmWkRCEqAEhKmOxlpDVEFk+sb8oLbrjhf/rudDpJ1av7rwvSdIW/Xk1
Js6kK/WOLWh2W7oTA6mybtBP7pNDvrZl8RdW/fvREVZdT4mqjtheWcbGunb+zsX1
BP8cKIngtvrZ37QPj72KnC4VJ7plJ52M+H4fwMDGIjayXjq3agJ+OjZC1ZZdND3+
7XOlQaxZs0AoavLEgc2Va5N8YlwDcL42R/cQAkprUY8XBIDy2hvvl4AusHW6iXf/
AMbhcpjSbdA5MeXcLYsoCcvEuJnSWJLm2auDMDILdDIWzE0X6Su5dKyCCpXXhtNZ
2nVRlpe0PnLcdcirBSqfafjN9YQEWBRE+kq42VQWV3bAEB/En0J5ynB1ZaqDbe/l
U4tPtgXcfr0nBh3EWlwP8W4FDwof2kS7aOd8dUfwXTxjsL3pVOFiXg1hpx9Nq+8s
B6vguFW4SG6j16WuYz9xsrBriG3KNm9948aAfxd5ReEafuJbNp574lsuyxZ3BVXM
LCWjaa+TBYQifStl0PZLiMFTluahcOfmWRwd2pp97daK8iZoIuR12Ks3UjDMJNoo
owqSOxJpyQlY6HIFINm1Gz4BDuYfXN6Nw7kKsYgzRzRR+3DQFfUIbEQAIR/f5u9r
o1CAjRpHaOZ07ChxktyRVyRgLeAnhVICbvkeZCtwiqHdNhW0mC1kMtT2bj6XZgjc
u7DDqUWj6Dyr/IaRPRw6AcVIktYEM/hSTxv5AlOB5POtUoVNE7pE1qVTydgzVAzl
Q8WDBDD/IOoIVRpuIojqxNdM4WnZLnrPYfUqozH/fbBIqoOmWHkV4AEo7EeQLYSQ
yUu5/khJLkNa5rZyaIQPz+9ukRVBlz9YeqtMegXeNa0MvUAt2VzePIkj+qHCEIm1
gLZfdP9JOnqnMSYDN+NdNNCI3/c8eKkDC8LlXvLZqwo0jPLEWWUo1h6iAmTyHfih
Q3xl3jvXwyFbJ6tJtE+vGeEX9Yx3TuaNafA2nxb43f6bnwQ7pSoWhMYjUVqUbfVA
E19GIGh5lzfFrtL2JlSKlH5BzyMrtBUO07l30oQ78HgzzV7niC4MAEh74soip5vd
osCXnT1L18t6mzP7fiiBBYrK7fGtHYBkEXohw913/aac0spaA2FUTu0ZcKSnQyJ0
fWRRrzqO5qa9rxN+TV+yGp7hPXvR5A7cUtj9FDkRf4VGBQV6genRMwbsJXzRjmQj
q3BZ64BFdtVBR5PQFf06g3GdYjb+tVyEQrXP5vhxqdT7Do06vql8sNHhOJXUwI/c
QxH8UJg+aJijrNF4u+BsqVGB8yInE861o60e3TiJ9fFOzXLh8lvJgCuAbdNfpftL
8m3dqv82Pj8mFvJ8SDheBQWLAfgB/AIyGNHuCHCbBMs4fFCC6iN1w3TvKptRETfA
pXmoh0l3C9uYK8MVtSEXcfApl7yThB/N0QoBN/eNWjRTFqfQmwlt0umr/olfkZ/0
T5DfrytMx5eOjfxfI2ZLMTMNxx/OWByQSHt1t2zul/4kVzJ1gR7WJF0Rro3sS9DA
rjq4mbTqsVtw5FYpeBxluD7BdIy/d/B9tUV+sHrhD4689Rmf666o1VlRON0/kQ5z
8a7kWsDnfYatjvTTPO1eJAJWgdfc29OR5KkWaPOaD3mrPk3xBSIeDya/Pdp0a+q8
thkUDkicF4GGH0nYzNWx6+kkQQZ5lFv60pBtHIFFB6moU4lTwEaf07cA4WguCAqD
vhDHJH+QFWPzv54Pw7/V7UyLQ0WLIJZh3eJTX4pN5bAKbuqTwrYWpZlCStxeAmpg
ByVdFs9cUwqrU1AQtQIpFdjTLpTsB3CoMacZRsq4QpDuIlSoD/oFOfckjc6mF2pE
tohUazCF43vu+Ji2HM/FULR8Z5t69r+8+EDKWH5vYox5xU93WPd/GLyCRVwxQycq
SczZ0hypwkq0cOWV2xlIdF7xIrzfzK10A6VOF5gu55uA0NYi/LodiGqduSyXcx6R
9YebHaJdYkMeI/WR4TVOvBF/N6vdwyZ3UFNL+OfNmniG+bwQF4jLC2WTiFuhaGT2
QD6HzwjaU22es0UMFxahBOUarWzuPEFLEbScbbvTnTr6zUSGKcskfArn3znxxZ4k
7xH+kTT8tl0Zgk342/S30yujHlxWhallHv4d/5Ly/EdvGb3vAlfCFnWi5vIhBCBh
pOUjh63kWbdRsN9qWX5hkkjwSm0lZhG1rhyvvNXZB8dr0aJ6HSTBOYMhvM8AO1E8
6K8X0Y6xE3E9EBi5ddwaTcV8VsG5ZWJjTUIpwCELBR9uQErWGuZotCKN/qxyghrf
oBc+lg99T4/f0XEps/ZB+A10WEfxON5qehYJoPrNqJuzSVbOhfVI9xLwQZGvlTjD
8FxH5HfhPiMcD8BPAK/tGNLjQp5GCF9+HMU4tJZsk8KGnGW44qEuvgtJO8d0CDib
JlR0Vmn07sEvASeggFCTe41oqWeB5hGF0dYxeqmJLPMiDRGzB6QmqNgI9sqzkrj8
EUcRywHNDdTLrOMqfSPKrjhx2hjLfy2vxgq9FgqNQZxroYgtQGjtj9bBGwAzLTac
WEAIYhsZ2jPN/jHnzKExzpEVHdQ8DWfRnmpEaNz7ZOUTFS1K4ldP36yFL2ClRWXW
Tgckm6iyb/xDnGq5cFSgkbp1C4ytWEHgJ8c2tzJTsXOL+QOqaMxit0MHqhAN2SOa
8HTcPC2sq6Wg8jqu0aXjVb4aR9iQ1+mz7mmB6RV+tRFEYlzlkGl82h1yftN60WqF
j5rk3I21sTScsPYa6ephYg1wjNyZOtxDyzKclndr1I+5jeZWsAkAv1R+x9OXDk9E
v0IH3xLSdcvjQuaamOsHpggThHbmcEWZAckRk/kqQtrWI4lJ9xvolwCP/qtr+N2T
nhd701h78bienPJgPgZw+5jM9qqrovcyviYcah8pDzLggcvpsbXIDgyMuXUPsAAA
gsy+pSHBzcmR7JTVh9ruXK7BBah5UWrr3XaYNrn5TFq3BbM8oMHa+deYRgIrzR4C
8xKg3nVEsjcXDVqTnV/UxzvEncAHUf+T3CRfo/ZLV1ymF7ZO0MMwiC08nM6f6Q26
aVagFIYrZMuloh9Pwh0ozsRnNHRkm7dowoYueDxZsYJrCtRtEwzFajfPo91GdekA
XWvrsIye5ttjSdA6IQbIDzLhzGarr5bRN55jmjw2lIu9jJlG5VDyfzTp9jwb/GxS
Y2XjB2M2qRqtjK3DHFiJJ1ldcqG3LzSPhntuDnXmbW5qhwI37RzrJa5RUo04bEZO
00Uqm7sNCOLPJa6b4GTu7uDmjz1QXpjBn46BZpy7tEmWH9ij6l4z9kSQyAHS62En
/6kSeXHokqJyHBbvygUrcepcLYoHrWcm7yrtgocfaUI6e4S2Lv80KeinZnJOZbOG
Z2dPNqRVpVNxVVw45oAN3eczP4W6D61RBXezHYGUbK009JmdMU29IcmFXr1XGKwt
KDkhtv9kKpjCbZvnwr6e93EPFd/z4w+M8O1/D+u2v6vqkkEX9MnL3Oj04+a2X141
bH6nEVKXpT1N/qHT0J0wTZn8jKfTc6OT4BdyAuGcdtNk/WQkcCCfjrts4C9qhhRO
wqzitaB/EQxC0vfZ3JvkFNgukbaJfw/t7Z2qt5jNyNnlqQMwp5d2Hne7f0/RwJnj
k1Yu4MxwxlDHRUVOgJZvj9ykrRMvFpTqsflftmUp/Jpvhr6ICOsb7DdMRJuCZaqh
RvQP6U9wV5NN1o94/NkhVJctHFgcd+ZW8nDOJk58jJd+gVfBpJX5nVW6Ut9pDmih
CLZ3LmS9lssB/wPwemQMGeEOHxU7WnNJE2H8bZ8/tOkbO4pgdNlmYbhyqr3SuyKL
uyTDtUTOWByLoQCsJbE3XoL4JHJx8u+8jyA6hOJXtTxWkZX8B0i1zhHvY+q3w2X8
JVdGZGZ4pOviERmiQpQ28npSG9q7u8epsYt17NxUKC9ZX5xk7FeBjz8AgFK7W+wp
P6D4WRsOVNwp/JErxUNfa7XAttOboepRx1GZrwNqbWruPeWXYs/3obvUYCRsiyWa
WYSNTd3s7Jcd0jdhHD5+JnXoxdfreTZnWTAy3woXRB5Uw29IOq0/R8oQnMQJySQC
UJI+d7EgLLBYHJR9XYfj+QVOHVBrD25PC1TaQCsj3PyULDTp0AVSuSI8wChcp/Pz
y5SStGUkYws5gLS8NuPb5vnD3eCs50PQ6fUBlBU2K9M/z+bp37D6Gs5Y0HMXdx96
QxbeE8bauPYd1MTaP51TCZPGtF2TUcHWTz/yUZ+WtMVLkPVGYkzWXh1gg8InC7cK
EQRo0hIMrfA/gQscWRV71Y2db27OKGuzXWYSdZTzhm/wWu4h0c7vo3DZXfhk24vi
hgF+y7zHmqBESBXDvzJWIpjT9kT2nIjSHhfC5c+1cjMO5WqRRUVsiZkvY+ovKAc8
3M88dKa4qwiSV5eAcbW3LuXGioZyjnLZn5X1RuHleSQzpLb7wp7bG0xenkdcDpT2
DH//4y/AowgB3kYRFXykuNL8GFAn38EIkZ3ikLzIVU5kLHswARdKPxheQpy79STM
g8ahS9pSMw8kQBpQalmLGWekuYAIyLCjh5MvQZJHApdKYe5eN29059bYPgkXKxYF
M1UPIUS0y2ALkoWXhtLyGcCJzYrBSA/ybqoKlWgSupjQPUlOFKq2+PWzo+dmhkr5
ibuPu2u3AFe1GiiAsHNLKPflvcE1Us/nq6BKBtY6AwrJtB0jSkRtOZ34vn252Hqc
0AVuq/HVIvbpmqXCbh0zD8Ic9oJ5I0mC1bFsPvXiYAldUdeu8pEFwLjQEh1CP0jI
oKKvCixHRRN8Owl+S6nJKUvpohQRCJMgG+vzWzM0Vy+z5DQa1XBCqy3iog8o41QS
yVF3Dk/Bv/Gp2lhAG/gTOd18P2r3+m/ZKgTHWsTLKldwEqVU8N+SK3blVpdtrUf7
nQZkYZQiF+PpGh4MIk4Jr2lIpyZN0GlhQn6QPQXAzL8e0OYQgNZ4PJ42gBHkRlRW
VXlum1OHrYyrp3L/a89KBE/lDdwtqbHctc8Z/mWHBV35UQN62Xt/rOkTeHtUDMsU
9DqaMwJZ+EBWh4DLrsO2mheDXVVx10gmhNNdJkYVrs+vMVxuxaTAEztw99lhKFxS
yHJqcQ5ZG0sRC2IUr2q5E5c/4nceT942JdOLIVAH6CKtkP8jy9jn8jD05ELaBEw1
Y/KgdDkf9f3RAzTjXjcUrs6V4WjnxfN9e5IVJ4ermyIO0vMdhLRLWpgPN9lZ7xGU
Xus7ysjSX+mgb2Wj+72hAp0bc9fZm1+VCBmGEqaZDAvecwog9dfer4lhAlyXdlV8
u975jT/P5q6oDieOvxWSkpAAOLpkJ4WIMH+S0CSaQ26IPSII29jHcjkqUrY0wTPa
y/qMlxBaBUWhnpLpjgaf+/y683ONtQuwIVdhlDb7wB3ZOt0YUpxz9Wja3PDlCCSl
voahLWbdg13hF54X5AvaC9HnFm6a5HRgCysDToadIsLvWMgI07RSeD/mmb8ordFo
GalZq/BZRLz2e/jktoApOu6mSqZWNpJ33T+LsIAWgLX+NHdNPJ/9afV3KhV4l53j
2UiOc/zv12ZeBLgT/hBKT2wvgVZuSXy4DqHkAnDrSsKFzD73EO+At8Sxns946nEx
a3TmcElQaAq5VxyasmnTBBdZfiEL0x4s74VWzUTYvKeOVLm61VzcaC6wKx9pee11
PRL2gRGOPpOHqmbkoLM91I8/nOzCeTlrJLtad9pNwevBLN8oY7HLYc2a6jzh6Jhk
90ciCwVGadS8pefC52711DJtGGKd7PqlGKJzMrfQL+BRAU/ItLNGSpiIFQh7O+pr
xIWqwEVSm/NUt0wgFpVANyUDRrGitLUKJ1lEs9dNVoCXH/TtbjA22VWlUeqcGsAx
iHBeyyTjlyuGuECVytfZVpA4MiO2DRuuUTjgqwdl1dbOqcr9c/mTqzIxEndmbeNi
OG+4hYS1KpYWQ2mM9mtGQ+6v5LaHuZn/cyL0e9BwThYPhuUV4BXqYY3yP4UUvW8i
9TEc+34Dzrygk5WtXsbfj4Ax+bHwfwgDEXzkbvQJy+BdMkZ4fgiiVRuIwbWstGJS
mtpeQ65ts061nag+pFvMDQiIPbnZaoRe3GtKCAmPhUK10tU6AKDLgjXAA5j/slY4
Mg4TFXV6ZarexHSg8QqPSQQoLE3t3Vr3p4A0WI/7XM1ds2CK5EiUs+FA/kqfAAL1
Q4tV2OUsqfKv/r3ZNSqiwbJh4RErr/bu9kN7qfwhLSd+n1pgtMuq10ZC775UGvkS
o/iyOrMFL3795UyjYXmw/prK1MyUBvEK5897D3b4Q5p9ei3WTYlQ/qnkcJSWHt5e
OM7nAoKj1wUnC7SHt/oEXXFX3/he0IX/v5Dc4BjYVQmwxksBh1GzMyFsK2dqdVFE
CBX3E+a/0uKV0BnknlsbQgMgqcqwo4BGtzPKxlCyJOJwqFiiDw4wUJCtqmMhzzLv
R4fME2xqz0MG6+SkNKB/VfC+LrctXgnMho064KLGzGbawHjm7/KnoDNOlAgDDEnq
dcJ4YUQ9kO2TG35Yy36qxAs0e+ptyVZwLU1sKHr7iSyrrPrq31gj+rQaE0A+Cthb
SbW8P+4X033dBie2Km4qyA3qUDFq++Q6RRi9m3zH2AqPEYnm76GaoS9SSd9ODSNL
NrInF6SXhaIZvwAYkqwO2GSYq3dfiSasZX3WXFUqfB/ywq7Dabi4X8MPoDNg0CE/
HmyXx9fQc+PQGIfEvoAhUAEwGX9zKeUDijFgs/1u9Njabm6MtrcbbMFjGrUluVxR
9r/FLf4kDEw2urzAi/eF0KfHUiWAB2NoWAmGnRRFSNEnEhzOvRFYEJdomDtE3OEh
WtlU19Dj+NcVVSJIQ+DlMWZWi2hU4cdj6dsICOHqlyzYUPBMc2NKc6laPhfCEDXt
SwrATQfWOPjSHkWuRJM76SqYh3wSb3hZ7NpGpVG0dEgbStRDMY8FLCg65K4GPfqQ
JdoLCWkvK8gWlMRcOi7clPeLudeyc/Wpj8g8NcTQmY7/fREnazyAWM8uLHMX/fxh
/ewCm880DS2GN6jDcfago1PvP8oYf7mZ6bX0h0t4idjUnWfs59CrLXbGlGI2axwH
BsedErHY5mHmAANj2hcr8XHsvvnGzYAnO3NlxAnBy8nB+NskpgVqTJMfkG3MaSLs
L6c21AfstEkvtX8ueCxvYinL7gs5cKBt8R4Wl75CDbCUlnKzyAPmjHm3qbhXxF/r
dH0EpPxqQLgtsGSZ61em7+6i8o847FqKU83OYaKAn9P5E0H8QfHvTYyQO41pyqMy
CDmGAzB4Noz82utoMfJw31O1jPirFEzfzA6SNdMYIsLGQu1lqfro6AP/Uo1ufKIC
B9RYJrTLM1QkkpeN4xa3MREE9zenNsmGnJK/Of2EcEldrHzQBUR1EC9GCyzZGVLj
7OV0gxmB/BImtoKEzSKAKWAs+3J5PUBcBaaxwXVghARJMc8AiQva4diYJPV27zru
rVz/+84GEEPYnIzmSIS2n9g5OuoITxAIZxFL9UZ59zN7Kk1Y2s7IXrOIFjmTDnzg
zVWgJJttIRp4SW0zzTvf40kNMDvqx6Ub+u9vjQoB1zxJpsUdSo2NhFgHxw4EX5XJ
9neJG+vJSUHNLYuPz4msC55dVCbSyAEx/GaN2L14ewjsWHxDBN/H9ldKDxVa78hF
IMZ1o+U0ryy5meoWP89kjXteZlygizrJOBrwKUpr3tntiy1LHPI8QjE7ZvfEEUx9
sc/hCAWY6Ijxyru12yk9o2VzXfGK8Dggz1+qWJJ3Z5LqFZTveT+OWBVTFkNKnFWW
gG8stQpYua8ssrBAkbVD5uYgOEtBgngEOhx0o5luM5PedVJ5axz8wLkCVnAb1KFA
gIbhbX1RqBQw6LldG0jmQ0mD4mTY/xb1dI2teAGQAad2xX6ryGgSrA1sJg2soGKd
Zu5jg/IO2OzXvPgDo6akoNh7Xs3DtACoTSAf7JkeHMoro4Vy3z3PwaeB+QZly0iF
NgAHC1+0lFDQlWRIPcCQMETs4TzWZC3GHOazSIIUK9m6BH5Wc9+XtdN6fhovAt5+
eoI44/9zpOtkMWHAa2rI2L38g6z0awE2Tj7Pfxks7k0UGemt/iYq8EJAhPvGx3bH
QrGkvTynf48xS2XHnKz/J7TN58bvxwqJPGTJZPtH0VcW9LkWdKyEmzK+m+5NEug0
/oSeIt8qJ4xMRPSdsREOKT5VQaA9dUdxbyA4o5Vojq48KO50uFnPqhwSAyZfZiTg
s1oWnVLdT1f4kdXEi1+AZ692cMY0zgGsqKEXhw/QJyhPpQRYWhARl06haVbPN6HP
wvIcrhMl/Q3jEYfNPUyI2BOieDizIw2pQqa5U32Wlh0uYNbw5QWfpU7R/Nw0qXmG
gjuCTU4Ma8UtxB94zLp9Z+1gk0r6ylTVEpAa3cP2IXE5wenKa/Xvf0y87kMKMBkv
UAA7aV0mPz8LYHWA1fMpwL0Z/xvnHT2/2VLtsoJVg+/Xc/EC1S0XXmGbHlYWY6pe
mHCxoz1p70KNtRvH9isZqBCA8iM8s/Fg5EG9VwhlfYKQwiGVgWl6f+5XDC1uwdFV
/0nayN8KGBQGKwzP9spw6fzE6NDXzF9l05AYlXHwMFwlX0TwiAPObnhsJ0OnTskf
ZDWDVu6E5qIFApqob2fkoljt2l0Bhz2/2xCwf9bW+bYv3WDnl7zJFTM/pbRTW1sg
qwhj2ro9ntZ7OBHPn2B76MXxELzCQTDTo8qA0x66UiV15vLKLh7oNWx5wSc8X65h
EHJBsYdSl4PE+cGv9mdYlOCy01TakW+F9g62HrYen20lgcM97qYD7HFs7J42y2/W
PoGQAdzI4gPLm852tH1MTN1vnxZnzLl1UTZ7/xQJNeuDGBBLqqcmozrI1TVmmcyY
GaR1/zFTGa1p8/xXA6UKrJ/S0rYod2Pbzu16bsM1FiW7sNmtQUqeiAHB2fXlW7q1
rUFhoqoPbeikSIQVyI+Js/SR8mleh+cG/UqLwzOKAP+9He7IkgN1lS3Ih4MFfOUw
aSfKroANlOOM94+VkH9aDIN+TWTfUep2Yt8oJgnZynxNoQDNzVWBGXrTQ2rwdK9K
6BHEUjtKcc+k8bHsvrcKM23Iz12jrUnfqcpggyi5SN6cHctqYl9WDA6buD8ZHlRM
UiYUdtwJOJhQO34EjFpGDDwtcLeD64EXV92vVg9sXCyujDA4keJ4GXaYVJ0plZ7O
qB9TX7hxvx4dNO7/rfVdCqE/r92LlewSgwOtXyzT9DAinpbwzXK9Q0Pq+tuLcu1i
2ECNmQAZz5QDWpNiDvVxA68ihlxIOY3wHyDhFjfpcoV5QJoN3bY6rxbSxObqvfP2
2GJImxmsyoWogoGHqzELWqIA6Nx9VPake4yOmGetGYccYH9W3ENauZdCHlXKiFcD
KaY68BNQ84yAb2AdrU7e60VG8OhfiIg729Ku6OmBErFhm+Qk+MY9douLZd/kV3v2
nnZqsVbaQIFXBldloiPwA4gPiyTsRdx/0mDAy4ioFhart7SaUKIjMkbSR/m8Z5Jd
07ycnD/K57p9EPNDNco/WGt/dz5nNtpqBP5oEe5mnQObFLktNAlaefbqA93fVyoF
IozP8EZd09H0brjTIl0ROWl1GA4ygPuJpbICVSYA22Qjo1fSad9FIZhwzxTYoWWA
CKAM9nB6RYdPsxmoTsfxuDYi9f3s+cfwzTm6eBWhfheulYTnjoRg4G6D7kVeeijX
cVnYzS3PJmdQSGixh4CsCyIGEyNXY8kqx0FskcVYJyF7hD/vGCkKx3+UgItPLpet
CXL3E8LmjpVj/te0tNGAslpTCOSlIfwhX+RRbMVs4wnLCUPVKwbG6V8KOF5obVJq
rGiDL80pWFCe+fPhHHxBcVVVbr/ahETXpvGh4R15giYYZOv+tGmmJXNVAhw5kQBi
rMgGVStVG9elrokONPGh9osTQmX7YmgpUGCzxS2NbhV6yz9PgkPiF72wpI2KqCf1
7cOWkqVLyzVGmlcDL15WNuVz+Jpc8cL4orqCmCO9gar6KBdADshaP205Qkf2+VNg
NRdOYgSAYBKzs2NY5LxPDosxUax0bFnec7SkbHYmb4ZbtRPalH8q8WTQtZzSdjMt
moJE5YiAvxRtRSUPw+nOM0FzK+3QSw9WouuKkBTWp9t0PJOlKxp+5L8JVnEIuneO
A+BKnPsvHQBRbxa01L0jUBPq+ZD3ZtC/yDfgQcGnqWRzdCYaFKeg6gv14cQ3H0uc
5rgVLWRWPIP4Jk05ZYpvS5+WeykO4oUuE9++Aroz3SRxkM9Bil8EeacsZSXhhPD+
YI5GYsvDDLlSAfvdqppA2PA7i98xQuB8G120rdYjyJYRu5ThXcu08aFihEo3l4UV
lVD4SRbpxjvXvMCnCxD//vdTFfpDS++Fvf7DY2+Syfxr8eokUymLbYxRyYdZoh62
7u6n6sAX5GP2/dAlsjFCLssntlAXA2J8FRWh7OC+BVq2a9qR8V1fj1Svsro41no0
OMz3Hd8YUkNnH4Bmkx40SNo/gNgUZ4wjSzucpIKwxsTmO+3sVKj9Di8bOhn5BKbr
POy061eZu1eSuyGdnanLnLt/Qf0XRfgCBkWKc9/XqqtiVfm4hF0FgvI/2NjtA+cf
Ihk1hpOmnEXIHyprxH5m8/X0zmo4LM0G9FmN1R7/0VQryVX7/TIIhRDZvvEKNpTK
Dk3v1ovLwoEAkVAK5iPzrwhD+Phy2OzgVBpeyL8Anyfh3MblTkxnBFdrVXYeDHmx
XfGgdmZ1Gz0XmBr12D4L1hP7BOr8X05CWWJVf0pFZCOLcM0nCRX6eWSZrKjjgbze
W20U9gmS6Uw66nTWlWqwK+nDHqDSirtHIxtdZoQLK5U90k5PoZRM/SX6lF4TQNrY
ZvtYfBNNhSXtX4Z+enXzwSUBntTv9Ga+vbKZQ+vwB+usy6RNdDSydJD6C0NW/yN4
R/hk5J1DcX+xpNnICHsnnGECYg/pSRbCLanXmVZrSo2hlTOfMNnfmPocda+b6/rx
woh8XriTqaEi2n7w99Ff76a6iiZ60kcCLbWYFOIycF7zS9uaSepf6GCyuFRU8y1F
MGI3TgMZ/xKws62f9mDZOc9UTz9Yh5ZTUAKbyykPmmDMCqnnTuuOt2RO2ZJ6OmaZ
2U0fVLSp7JNDo/04ejVrChpEAPWSucmH0Dn8ajbsaNEbMLAWCCDNnc94eiAC070q
wkRxPzYGsBp1cJ5qY879Q3PLZ7o9d9s3m1ti/VKoS9lunEIxO318A84T0h0oIM64
dFbOnNk5nyt/ZTC8jtzlXgE0UYv7FyCOAf7r/KOUedGQDyFu0veOTRAwpSWryN67
sbqcOW9y7bbeZ/t2/srfy41MZLbBBNc2L/q2pbSGqF71Ft0wP/sxuTk6R7vDvaE3
YBi45K6OYrhn0ZgJ8mHgqFX8WoadUESQSV15B5HHBoyesT4OSprv43uQf/xLLmQG
vr9jc8tEUBlhQhE8t7j1sV6LdXgjBYUxVxt9GMWXFJAPMnE0ZfHFE9kSjfNsWDH7
xMfUvdY883bFUTqsqIsxZkCMmVfm1NlW63NcPF4i+wKEEZm+qcjgOzi/i0o1z4of
7XXJDQlT8DDRgVs2Qix7D4MRO8xGGZN6UfxIiEdc+y3S7z2mJhoclVJUc8pkMQG1
CDWbcVRe69vACow7fPn+XID7dglS4AKWe54jF8JVul2deM57oWQ/4rPLlMxRvrj2
SeEpNl/lxdkwirKxFFmJKFapLQ6Egyx+Qj1/19rzPnzz0BM5Qcjlsij2lsBkUPWo
DVfFaE2/DqAPR+4cYIJ3yb7gujC1acuWOVWzTGlOywQ8rVx90VUgfnBauyr4GA77
MZg0VcSZr9UKIArNPr3lmuInUASC9f6THfm72nYnBsWnLlfbqmoDnPs0DjyxSP9i
u1ilTIX2hq4LR+wZnrgDKPhH0fCUjBrdjmN4cgrCR6cHaDSU0+5gT2jjYPtEto1c
Za+LM/8Y+N+167MckzfxJRYtpny61/bgpSRX+UQcQeukimcctUn8O+NlBkkdVDPb
H5SX4k+Hmq1AhgMHSsU8Lwz40phSDEnJsAocKA3aBUYe5usktEe0ufvtdfyviD+T
c06mXpkEtdZHm2A3W2sBTNQLNAZKkHbPh3cFooCw6hcY+fa9bSKdAXQHQccUKG84
rHMM4LFFsfczl+aMfoSnBcsY0jzpXn9DDir3B+LFfE9V3qdoG2KTRs06oWiVq98F
nSs0mMc+JxvLwgoIZFnDwpHfgT0VdzFO8X4OUoXvNLOmsPXflnLcV0mmhaxJxB7p
4/vcCK8z+/Shlg24awYywMB/ZE6lkHBzxRWgbJH7FL7GwKTK2CU8uTrkXf04EPfO
SUCRrTLUH2x95pFpnz98JXy/xU7IL7ofclo1wmmQ0j0uZVDy8H28fKWh2EO2ZSlG
KMwfBeQqRQL/x0gHrKMWKXWW1eYLbFq1xb5PtLTs8VZ9QPnOclAtalZdJoe9Bxsl
hP9iCxCvar+erb3II0vLMng8i8kmtRhZR6PVaX8W08auiptQvIw2btDV8a7lJv/b
uzZwriOU+k/jWIdDag3XR3OoF9xUlDopLxXAZ5omvb6Ol4BobDWJBO+KuwPPV+Vt
3d/USrIWsiccDGwu+hbiPwT4Ae2ngF7orL7JcWR7WK1CLBnVgJbA6d8jJlj+rwPv
xcKApW3Vs83CHnEJZIrRyZS2Y5CU+1dWPgtBn9ZyNrrjw6RHzhap/S0B/vEvXMRg
B6YPfcXz57MK8sNOQE/p77v7JojdyI6leO5x4TwGdM0OgJj7YNKojQc92/paasNI
VYgrRSzDdIAW5OqYj4Z//b+0XFhYX7u2Dd+b5m+bsE3YQCS8CBtyn6/Kwa/DJ6iH
rFS6NzAAwdUS4I42ahWXOA/A0d34iU/NGDfLQ3AHj0o2P4TWJrTP1/VEjT8jF+LL
w+J3l5uBNYuTIhKW405ZBN32Kx6qt8RaFk5F7SxclCm6y1lmKY22L7PUMJDPjPMO
Ume482OY9Mebf4ENJhN7S3V3YX3n0qAB6k8LYYiz+G2a71JIZVaDMJQdsjDptvue
2t6wqx30nVZQ35p0kZyprWqC12rufbz54gTqEzNrhHcDEKQbRlBiG1hspkw0KtHq
XnQVh3lrGHwSf1vU+J1N0qBsgIyNiEiDqh6UyzFvlp0oqlL9CKmYyW6J1DlVPo8E
Zu4Y86Y8fLyjMGyGxWX5VU5p1jdTAtAOVnG/d+3Lta0JEe/NP13aRySBxyI8SfJ5
R6vuIf62OlyYrxPSuUqCawPae3uzJcZ9lUO+yFU6ZyaiClKJwB8vfqA/rZBcAgU+
zFe57iyOFF1/urtAZ1e9yIEk+dNByhsFn1LwMU/TZHQC6fvCx+S03jHvjK7zBq9i
jEdfK2sX2JNvkfxU0vYgflRUQcCB9IsZgRTSgIDDA0skOGPppfNsrTPWv1hXJJGL
KWzzkHGUwLE+/1npr0/erOl++vRZWbMI+j5/qWraw4GgxE3DVK0781V/TD7vmlva
9oBZWwpyQ0b+dgy7Kgn9m5hq74AJ7WoqBcBvdwpI/+U9qoVVswUdfusiXwPB5pEZ
RD2fP7+CO1pyEiLh4BE9YTPf3+cRYTrBIxlGakdjrqVdUHd3D5NeZVOjkA9b9ejb
FMmVwbzpE1XN7cm/Cezqx6ckb+ucOZUL7xLp84VaICYSjtYeLTYybPiTqa1SBC8i
siqD4kP/jTezV4+fmr/kmkT+toEJ5TGXe0kkPa1FUfjlqlBIEuB38q3nCUvmWybR
owes0oZlaByh71C7SdKoM0da59UyMvsLlvzGEYZxU/81EokhElINBtXklyh0AYL3
xL4ApppzYmk3h718FNw62G4rk/tbWYeCSt2AsEavGqtGaQYSeUUa9nkuIEBdO/3C
T3NHFob2N9GbJmKY2tKzxC20GavEVLnS4rvTeV17eo8KWUGIWbhNapjn39vbfjFA
kPWn3PfY0EKN+vMI4BBwcUSZlbn+2a35oBgbwt2M7FUYJqdf1GIs1PuFNqy/rEpX
KJedHEAdoBhmALTdaCV3ZVGFxEo5EBzdYPZ6dl0BTF4kACyl03DoSrrsx4mXO9ua
qMozeMoEx0l9otDIeknMu3HpzY7oaaU/H24haTwfCEvJDQ6Cdxwmbvdh4SlxaUNn
qvCUlz60Z85Tf4UzCeI2TeoWbt4312xYDHtZdRtcRx8DKdfOwc6D07IxOtER/0Wj
E6ApG+O+7wO3ymZcuX2LqbpeALtUSq6ZDmaSYWmR3tVUfRm8tp++x1kq7t4d07qI
/1TLd+JPwhAOGzRaZBO4MtOJdDYTQJ50TA9AD/oDRXO2FLSjHcy++PtC9ALqmC9p
n/WCxtzh2IKyZKX4Z++DVtHk1rSN/Akc1VTCbcRyUiHLiVi63ZEUZjV+9K5YSBZk
7+PcmTqfJyxWJKnWo05dTYmQ7pr6+3fKrciWOc+prcShiGpXhliT5EXpW0JbkQyA
ny6uj9TO6mfsnuOj7LPl1T1mFLp85VgE2wfM6Cyvok28esmCYzbgEz3t4HRGNXMI
zCTamev4j2l64oTau3W7ZaoQ4dF88FvzzJS+JFkk1cKdbybwyRtSLi/oTtl/xkYx
5GVFDZGl+AQlZdnt9ThIS4y6X/KxDgCHKNwgRIbLNU2OAehRoCqc8TnWZn6f4h9C
FU5WyGCyNoYPrAorSdha0Jbaz26h/EyY57meSnen8y4n6azgMZHtC5hBqLDQCP4d
T1ob/B61r4DL7V7anNV3IjoP+GIWGZaDE5ZbCMr+7sHHrUcqAEj00Jarr1CRGqm4
X+fE8HtI8TwIRWkK8VozDeaX7s7aGG+zK8HNmQdvFHkBO+CnWocoe7fK+XFJTl2+
wjoWF/tFn4qXlsQ1PwCSkOgqSa91tOOTtNNGxoepxZztLLaP/Y8iIUkGdOkFpq2n
wqV9VuBbb/vKERfOPIfO091NCIOAUKrbdGNbCafayRaxV2xU3A4u9iQA5VB5ldnn
dIHkowG/jVvJ2C7FRGeQpmj+vRAEFQLGJrIfEBilCu7p1dwauvTV3EWKcG5cwNpO
RUwLbNt3xGJdlKNLVAH6r+18Pdakowoet5Biwn3tjVRuoLP97b5HKAPMVRL9+fLf
E1C0E59vK7gfbo5unjr8kRxf5pvtw4dOrEYS82bBpRuUUXYbEKMbmNqLyDsQWxVT
sr1VzWuGy6rniqOBGERBwhD9YBzrJFSau8gwhS7CW43rcAwCjP6cf9NFtj4HMumR
OxqSneqf8R34z3Nh39J/hdADJThldpJUzNMyAE7HQfy9UGbApyfsCJH7GhYsA2/4
I3pmIVJv9AYuHdPj8CG6eEbFE6+VNZ/YvOPZPRwR9tBeWkTPSBqpHDyMdM/+Z6cT
dY/dP45kDHA9MDAwwTj9Oqqe0REHaMqA76GZJzDJ711Q3MU1VyMPJWrR/ffO22zx
xAuK0W9KwWq1tIIRX1J+36dkw784iTz+dddi9OEKEAmxbT4b4VJxHWnnVo14lLZ/
Qrm/Dsis6pm6n0ZMEexcw6Mi2TQsfdk2gHGg117SEUsk2GVDjEmQXy/cQEjKSHvu
eajneHHlS5uxpdviz1Jpg15/ZLOxfC8aV/mYvsBQxkSBFSnrX2aAqyLAhUq+379y
F/PF/FLvyiOW8hRS3urgUxOmHTD8bL7eYNaCigeaR/zP7wg0RI32X0VlSKZ8JGOg
E5TKIG+aH78SnQ0EYH13IpvCJirXijGnrGfLwzsQ6a1RUMfTz+5ZrV8hiavPCjo2
4kA3OSmw0mSTxiXKXV88O9pFDNUZ6ekFaY+ngmwiW1u+rSpCuEWdaKJ4incjs0fl
eswa+lnt5EHRoPuudR/QfShNQzTA+xVsFVQYe8vnbX2/UgffA52MZJBc4AdRvabL
TlyayYr4ie1f6Jfdux6NQ3tDgt9ADtRuyJyDFSqBcCMRrgwS4MJ8hQ7l71Mf3FzZ
2XyyhHomDjSKD16N5Xoy+hpBm9auzbq0kcArddF8gNsXCxIVVj52gONYtFtkzKNm
xILOgwj3tyzP6pubnm5CHJLQN/SB16reo6JzrAstdaK6adfu5xDgkSY/gvTi1TqL
UTi1q5iCampbYSaoTRtSMMEVFTq137+RNMm3v9h/Iqpz4qg4UB9qqdEJwmyu2EqX
mWSTxSWbWef2BvxNsLp/jW0VWMayLXPHI2i+8uHrEdZyjYJjipN3Dr8qcflT/bh2
+ZZls98FQ3INRh/+VmdiXOWs4sKGHU8l54dPLKikZG8T9GIQZi4lXZwVoWBawLKL
CusFMY5u98xHPRcnE9qK5iHQjFfj80EvzaK7RAk+ifvr090lwxZiyvXkYvuLMAXZ
l19DU4OtKy5z3e9nyP2Xz5SXBx/XjnrMALyNO6jgYMBhk03EPQL0amv+t8x7Eivu
NYPg1U89ip9BY1J0vALn1lLRRJQRsPIGcvR7dMWRD+1gEZzsf6rnpZIkbrlskNDO
tVptG3UvSNvdMSpKMkqHMUBpt+bA295d1ygE1cDkZOWOJFt2xlDVl8qNVmF9dGpb
0N80M6IpfGF9I9kSwW0z2YflqBMRumQnQAGoggFb4AwMJhaZsre2RXyedqEbXRaE
kYH+ol4q1PupsgstvfkBfjJuIqJbc/WsoMR9cjfwHUW3zjsn2R9nQKQBBMY8VmIk
x/KB2/XP6+MYJRiJX8kccfKcL/BlF8QaOfKGxucGT3luTDkJadX8p1kPb+wwlxhV
JlZNMK9wug8M8rsvKvJe+T4r47VFs9KVUWjSATWsSE55vS8tze6TufaE1Vx4KJ/a
RMYRjHeUzrtbnHrkhmaynJpCeqVz8Md1cGz5+IfGaVyfVg2ZNMi25kDNylv21Zl7
ca5L8O37zpDlHwIgjNoXd6trJFcAnxt9G9fnZAvicAS4cFQGogARPBYFlVWW7Ltp
QAm4104fcaTqdfQ3w0qvF4RkJ79fnuIZioMtzuHjmbUiDIniZTyf7MALEPAozUqH
KGqrj2MxWJNOGPbZ6A2a72DI/QPSRN3ejodSf5SxvhgdcJGQpRnn9n/Oru/jNH42
dFjf5litEg1raPqFLFU7HkBoasFocpo+OOS+k+3z9SjpalD7eQFDXwnll9SuH11m
yr/F5XIwyiCl+d3zkbwA1D3OeQvCumxj6luXulZN9CTvnGFsQnfMpU84glZ6P+Ee
cnK8JvCEYQGtuAr9TGFxQxUr8GwPdXUxTXMaEYXOCEuwQKrv5DS97r3s6uKxv0Gn
mqg6dauheOHS0wQnF6p3nuESw9HYIGWugH+MAzSAeH2OHRqLSGBjBtWrwyLN/lTr
5KExFsEoGJNyUUdKK+MfFOsH8/wU0RkCDqeOhubB35khlUAwhQxjzxN8ORmfg6vC
Lgdqpkud5TyvPnV8DwBv4/lUrNU7lVVCiHOnVeZjkTJ5lsTi52ZyeyStjAWvH3UB
zoitlsivrka7DtiNGdCwHsz8vfspRgZz1LuOz1rYyMVxZ1wQ87IFYns2ItiqzTkq
RTEwkVSEXE0I8xqmKLZw0Sw0zWAlQSuNnsGsV7CCGdU4lgvqNjgJ70wD1XZgu1lJ
d4xNGRLFWROY8i6ZrbG2Cd3cpaQ7Kny8oxGXpABmDRyR4YPQtkw6IBGEdpd3KxDe
V/Rw+l4vnkUiQtFDi9EKVwdl/anlmK6OJiQZcMII2umP4RXg68OWZPvAjeeXHSOF
VwpyucskTz1LJySzQaj9cHHl7qe8CegZ3q6/uvTH6dU9InaKVZCDDHR68axUrHmM
nHTZkevjE2VxVNxXjd7GDf+oNmiB3cvwy+r+6KiaAuKX4lCoyXYVFuvhlFDGS//n
a2J2i75DiKOb3nj4zUAhZFAByaJNlcWySCrjyOLGIGUnprV7uoJzfYwTp+uWLNaf
zXso0PRapn31qXoE7GoMUu5Lfcctp6GzzWlAI7/YUljPNWoy96+6fpwk6zgTb42m
3huVhAZy1zcr4puIxkIS3NWdqFKIzaf0/3We7JjcOF2H5TBVckM/ldjme0t71E47
rAQTgi0sxzXr62A3LNu77Ms/c4Q33GrJcn1E1nWT74IGz9hJwKTnTQP8nBg/WICP
CvwowCXxQBrE5NxDHjYdXCuFrP2r8FpNjEl281XDgUTlCv86HJTbXT/1XxxV6MLc
i8UZGKiJzdox5dFBO4GZaQl8kM9BWF3E4Ei8+ooE3Ztd9PDAIwU62SDR7zESCRrQ
M0FimkfySxDaGSG2rsdOFoCiFTrHqcOCkmzEinX3n8wB/JPod9wsq0KKny6cDlI3
1E0thm5C7eHwwGM5sjB7DfTQhYvXzXGu+lLE59rC/8q4n0EFhX0ar6sjC/mWAhU1
OvzIjZ84eeMmQNlsB+ZCP2MowE128GFYk35Jko0siRmK3OoGnRDO7gXiVvMrSYld
URf7tmPHa6f3o9tbEqcBAlszn317Tw6Bq/9J/c7/lyK+o5WjDf4T7gwXgidY4IZE
wJTkD9vF/U0SOr4OkUPYQgO0No9WWGIQJlOwgO2QjMRwMIzp4W9xOhWSFmmvr3CJ
R0UvyPdqSpH0XNj6iXH1FRAmb4Fijr0uTv5YifYzxGZwLUp9f6j1EOCORA6FyQwG
amyb9TZbYg9RbBiBfUKDz0YA7XyqxHhPTXCExwy8EBQcKdJ4Hrx1f/bGUSlEVmHL
rWn6cZbnoPq0g7VP0c3qIziZoo0GiAMcHvfl4LAQ3o4KeDZ+hVKDZu7ZycnqKtcr
2h8Wxge+nRWJ2JW/KJt0KFZjQ81wuBWCR32iypbx5+t7t4/fFk2Rr2nQmtMBgWT3
6ImO+sZX2BKUQkyJ+CwQkmgv4KstcW2IcMNtFuh92tP2yhzLbR5yz2GEwl3mtHkC
cbrMwXu5jXdjo/zyFLhjWmSOQDYJWZYA9jaz3kBuVQmltA73oA20QP0uNgkLdqky
H+l8FS+TSK93iJjC0W3BQD1zBB+Pm55+9058tem0GZHpeQSHRy+vdw8IyxovDANB
2tDtj1riU686xwEUybo5dD+Fr+VSfPt25mMd1whHO2Yw64iIdXqWTR+wbC/g52fU
aJU9H2cplIPU7r//TDsM8ZgeV6y9qTm1CnEFgdwfuGavyCd1u8+C5vryRMZ5s7nJ
pgmjo8X91Rb4GOq9vDl4Opcb0EhdShMh+zev4qyWD/7XBh+S1UiLipslVbhhEF8q
XXaYhAPxM3QNhKP/MM8ajcn750tvIWXNZ5MhPyB3ccK3fFgqzuvp6lhtNUJaVsor
7vvKxj4IFtVM3QQu9TIKWG8P1Bb7MJyXVgvOedf9Y03j2wGaV4Lf+mRJsedA+l+F
yBk4xc9UKYPtjVqnagcVuEizFzSXsD3dGVUad68HA1rKe+pyv4+JjPctTlf/Tm3z
XMXTRjvcC/b++2XsTxL/R3f4LEW4l4yG//u/+HThvNBT6rZlhFquIPaEZ0/kgT0D
ZVzDWt4ZXlAm+3LQ6AeWEeM9jby85FwBgKXmIuWvDgHOT8tqyGarRwfRUeo+M/r3
VnP5pemNQyc3YQY7V4Uthcdb/nFGcOBIt83BSIMPB8/8pv2+wctJEZRm3Ph4bVqW
RBIKMvnR2ag7e3eCSJX5/7DhdMA4iRtDNWIMz/nmzChkmprhFxPMfYupoEsfYgbB
srVENr92WEFo6FWawFzmxV/eY1A3TMf5oa5irP1yyjcocNIewr6Zubpn732qz1WJ
itCcucI4FEe/YP0GmBPjAxq3JfRxT42KI98vIEMasSh6zW/XOoIgCg5pxuz1suFa
LvujDYAUbZpnedfKqSolvXO/867H/lMmF67Cn41k9pCO1mU9bXyXkNgPM+AFH0Ah
TeV559IH0WjeHW//izc+pBuI7OBAgwolCTyrFq9KxxJkZL6926K1OE/v3b8aPEC0
TMsfgr0/ydgbOCa6AyzRMW8AqETJmISLg5j0h8peyTmYKrtIhwf2WcAeDnLWqYDS
6/zfcgcQfe1ufCn8OFgM1C0qsQRNdyX8RYtwtejs+PydOEQ4oYOwn6sTQSWQuwt2
qQ94+JpN/gUD4LFYXAAMC3J2C9cMsH2n64HQaAWvWdk7ccNtg7gu7v9JmCSHwjne
8zNXHRvvu5dvGbqliftRso3cQN2O9uGgfBh16fFoowNoaFEeh1N7b/6ve4LKC4kZ
e915d7TKpyhYLH/Ylkrf7P1LtPMnBfuN4U3VgCaGJijPAEjhztxYv2osTywq9vDE
oOswrkAr/v7eJFr2BYbFSedeoD/OPu8mq6BA7K5zih8mZoYk0qZ3u3ql/PPXe+vQ
IoDeEJP5s/1x4gncVJ5kYBmDvtkQdgNaafH4z6fQIcSk5mTSCRQ+ytklNxJsHfrU
2q/1ipv7LJ1SR0k9F/6hJsYVn7i6PLmzelX7F+bPNcqqgOWsDVK2aacSOhLJ+Pk2
Ycm4yFWLe+WEpGPt4WoPkPGj2g1bRBMaS1kusQuWGTB6QRpSscEd7L6m8//13yjk
dXXBY5DPf7U44q8XVA9FYguMWJ6b/xY9AOeDJ6JNJz0NV5sN8E7BNXqw/SsUWf+Z
zXvjLvlgl1Z3dTM5P+ud+HqZkO9ogz/6P9bPU/eNAjU3/08hvyx1K9T9KKC6hSLL
9wzSrK9a0ujfES6J1wMP6+IVPS7Qbgs/UbCibYpcl7SU4vuyQb0gVOSfV976t9ya
Y0O9vwgK6al+So5LXI0DVsgvQ0ZoeaJM7OpmFu4LTo+8eXky6gHVCh3Egmg99XTa
Pan8pMus1FWWTju+dG6FHmiTCTPoMSK9g4kJulfpgZ0J25nsc2Nokmp64WBxM//e
ZXz3i33MRNelK4bEbtuFmgxvwooA70xAJBVlcLriKtmikVXIhLey4sVwGjUGlaJ3
BwcSCDJLQQ/WUI07XbHfTN1a1LIWnxcv9F9Xysr6rEDrb0mCspiZvVl2yPv1nNBx
8jRE3Hmy3h1/RYgHGqBoRrUL46upv9GOyOdxXNEg7Fr7niL25Pj2+IVsb9NceK+R
F92GbfnZLIpzfr99mvQGbeQFktdjTxG/MqqNYGdu9vx+cJfbzuT19nZ5oObjq7/Y
DtuVwd8zZYatH8HCfMB9KUDcQegPzZYOdY6FOo02KsRt7ou9urjrLXQ7vcYJ5iFF
qolVL1LXJ6OW1sPd3Yb7V+x+fJHKkqoB1q7DdjlHW9Eqrx8zdcivJPcR/8m7MiOQ
GlWzmFP8vo5kJyhzVR7P3uEBrSljFIlBkQW4B5YDRcgu27qysA7SraPp4PQqMiR5
TLWwH81adGN60e5E78inVyVvbydjdqXBjtXe+/XGMFX8qPaMe99j2wnJ4Ziflmwe
dTVhtVOsT95fPFeBiCKUj1wPk/aKh2wlsl51evZ7Q/STpDYzChNIiRIjc1397bo+
3lEUoqMtDzcUe96i/sCSxQB70/1Eya5GW6sKJhbDd3iKMuf5d/rZ+bgukuaqmknT
JOdZGTOUpNXDPz7dFvY2zR4rZVHrwFUm6FcU1cFqx/ydpkc00RwYzFSqZNmAepJW
MhABjfb2jpaoLkAK1onTK+SwFazKIfa27ybp945SFyTEFSnsuV8V44joNbaIoeBP
KEXRWU3nmQCLqrbFIJ0ZHp45K/JStv7k880ERRaoRBDkGtgJVTGAjUpIRg4pIE0x
6IQcZbl/79MfFiTfZlJytqWJJLNn/GDtRkDsthpdatPP1Oh8QGymgWH7FF1iK+TN
hf6e2mJl7RfLE8tyKmgIfnP3hokB+/UyfHT+4JOAHh6MFLfR+diAyIYuqnLdgHhe
7LB1qDTN4IUIf+HalkPaZT95FZ4Fh2qklbtOlv74lvaIH7p6W8owIfxDtzCgtUDV
Z8CfAA+VxcsL3Gn+V088edIeCvmo7tpzmLalckfxdp1vAEPjdEZ+Z0bdWxIqxJgY
JRswVswXieqvHEu5/QWnlL/bRpkYYFhtXAgMUkIhbN/QnTlPCbZLP3ZoaF2aD0VW
qc5GXKcZXmK3iYy7h1pgNvRcuuXCGc4vRaFAu5FGMjbrwE/SNmpH4NzgriFjZx/R
7MI7GI+GG4Kh2yWOfO+wwtzQTelkhKFBgoHpWoLUC/93GSzqn2BQQjoGb+pyihvt
6+Dv9V/fLWNXee0gV4qh3z/jamUZL9HIjNJfyl2qsKcK7ByjevVAD2dZpmE7tbnH
JvSYFi9BMeETVS9424tZmbcgaJ430w8Pe7ZAh9pOHkkpReETl38daTGkFFgRQfSH
sOZXg4GIKpCHeaawLLEDZCytCbpKNj6irkFrgmVqhgpka32BbJvaW0CFzIKSLRjZ
N3RMVQBRYPagQ3drDlZvkHn0PsHn99OXDBkBMBMBSEkH+Xc3nUxEF5G6u1Asnxs3
Krj2wOZLei23jMviE7NG0Dtpp2WI+G7Hbv9OZwOPJI0y++nxXeicfYthJBJwrVgB
2P63hwqnL9I6YVoYsJlV2hVXIYGpU5jl8u8TyC25DBDNQQXR013KFkQsch74BPrL
+1KqWEBVFWA2hhuiGsVqYsTmz8jy+WUDRKKT0iLCvPd0G+mQyIbjVQmWOg7TJzFE
issCRAxKQnyjcfHTncwziU/7xjNfo9z1xvqj61c6JnblDd2JqKhQGtknIdpZzEnQ
SKI0qhH1TqPUSgPYQSIsdlfDNflb8GkxdUaz56IzX1JaLSEtBtt41ckBWWxvthlM
GlDw7JfKamcw9v4QvdC+dbO8IGiIV/8UGYh5D6jYEAQHFGA0RflN3/wVbCDtHXh9
1TqLA3Scl3cxkeE9c/kaZaFqxkr1IJ8XctnZr676jgu68Yq+SZnKFomDhABkazI9
LLQzccl/rwe2KCHZpso1klqZc6c3R+JrKcVmrLiZx29ILtDFmH1B2HD3ZgAdz5y/
wLN1A4AOvkMAI43PrGiox8qTJD4SPYS4kvXnQuGSsDy19ma6HYltKpZA3mE6uRZ0
XhLEwnQe5Wt0gE3sAs3SbVPXOldT34FkqFMdMaI4LBX0Xp2D+B1/5MZ4GylHA0Vc
ntjWHusuRUE/CGtrNzO1b6F4BtfDW3QUB5oHc8afnDhzhZoCHUgLXFYD1JpXMoCP
T5sqlOfz7jcgJK53P3i/C3b+h3wPTLnY3LszfdN1oOU/95nj4Cmoy6HdmgoE2Ukn
dD5qGN8NGmKWMESNCO50xrVeRSSaOLhC4fiMz08maAHUPi0NL4BWtr3WU5OfFi45
0jqaIERgjCrMllaVpx4uIB0M4i5dC14CpSeomEhKeTFoXaw2/iVb8pvBXwy/8OgT
elqfSQ0KIW7gZt+GiXcyOFzrU99BTGtQ+aCjZZwhRa5VomfNigz/oeaucY5xZpr7
1Cmtdj/SI4rt02pkosgZXSlXRhWr40pILhP8kCnGWFdnbQMxDTedhVHMS1cyrB4S
eY4rFSn0c4PcKsTAzivFx9NVYJLXykab5KSCqqI2HX9sPfaJ9azni4NUDWsEoJza
y7QRg6HAv3ogGgBS0ipAM0Qe6Fd0fzOpm5TodnsD/GSAq4YPpMN3rHWXIymEPELy
9YFNU6/iu9wvB0yqjVvcX324HfRY21MA0v5+EKkf+yN5Mq/IOktZ68g+Qw9jpy90
jXzFeO+ys1uNwW2s0tAJkg9Q0Vajksreun77prKjgxxmtTJ09RF7Mu8rdDFrGOQf
+dVQXWwCiV5xZj5+3DrbnvCQmByTrbbydK40bQDd8tTorL/NIRbMoL0GHfOM6VQk
jEuhsnYDSqSToJNs77Kt2tfYLHVP7wLE0WraprPdFfS7HQ7dWHCZt9MsvCeB/U7i
FVU0MBW7ejL37jAdXn87sfUVYAUiJ6ta2CkCGMh27CKhTwVwH6ua/dOsUb24gHpF
x6aMuwOs5bd0rJ/K78B0tEAIM27sJSVqR3BP7Msr9WW5zjbmSMUi/F11XlV1b8Xe
WjF7K1mZ2sIck4ma1W5uCT4WsVSiEbTJAnAw7lV+DOLTpsYBQ7ZTRl6+Oar5wnyR
Mnd+z7hg5cwZcVNXq2lLg0S1/ClxWTmWtN89zAF7y2P9ef5W90+ytYt2FnmO2xaF
VA6kZzKBvFFeef/JA84bmmfNiHuMLZ83DvUoPo+mVy8/C0UV7NKz/XLDlz7ssXFi
QkPvoIQ8HbhTcpUbG+ZzrDAwZpGuC+haQKKcfFiN7YN/jpupwe51CCHiDHuVBceW
DkUkRjPRO6kcj3klvzGFhWm8nWoPTpOEvcQkbemWV4kpc8/zUtDRBeZqKUkYV+Y/
ZEY5blMiviM4BWerYSlxFfhPSbbUU973S9G/LAKJyUL/7WQcxgoCPtyAbLxv/TCH
tNT7Oz4x1uJDRelSXPrVnjW/8dneI/DIz7//0lMStalXWeb9O3zOWx+Q5Xz2JeFW
0EQF+l/KGSnNOPZRLrTqIGQgT6F3fE/yUlJBpfD5vj7xbuQIi4Qz9UTqRxSzsDXV
kjaifCmVtFI26p4etzBEufkfCeCUK8fnK78OFakBK9/qCOo67LtzHoVqk4F9SQF2
HDtQ4XJ8O8ArgrLSOYitFrXrXCL8s/RjFhoH5nCMntmB6BI2qSz9ZyC7gSAcHTK4
3UR1JIv/WWDONu2QghNAk050TeXoh+ZmFtCUq5jwuS3hLXoE+14ogv/Vm7+sAF1t
T00r/I92UJM62bF+b4uHsf6eb6UXC21sHa0m0in2xix4rAZ8xI7HOkEynN56U+oT
H71RQ8V5I7bnQRf6in1Hp5eLe8D4qisKdMPo4dTiKp2XSQuUXX6C5abhywqowrVo
7+PsTfuRiu2ROaIAPkdbA7/3kk5Jta4KSJ2NinGK2xxnKAFDCnNhroVpJuULgvtb
NiAQz87qCzTCpWWoLrSb9D2OtKO6kWDwU6Kau4heROZ3VzugWyuCcSZ58oMzib9s
OBAlrSUwq/8oqbjTXEMW7hlsxIM3ECfwe6u7WJz4zZC7mgEBY7CjHXBk4hZwHUPJ
RMJE6lWV/9GieuA4DHddJN7gMCqHs2Q4iHWKWBd3OY7cnvU0fcfNakfQGFEs3BPe
J9DyUU9wzjXr4EX6/+W+StyVyHnKHJuiFp2cp/S1n5/fnPasmyYgauDwNK6t9ls9
K9aAFfPIaFMewfduIav0XCE+HxuX1D4woMLnbhQ3mvySsdYQKBpmJyrNM4bi6Mow
DPuCjiP6dCB0jfLS/XRLULMvabyQ2gPMKaOj0Mzp5rgCVYoNIu1QFVoQPYuqdxFX
8e4L4jJxpPHHqJAb5jCQWm5JFzg69RZrQ3XlewIKbtblSOZ9EGhlWuFDFkOz3Sv7
xg0RyRk3OtvlThf20a5fOvev9TKwUpdi7UhZpoUYtQjTgiFi733YPV9a5Y1fh8g8
L7Jewjm0diFe7PkSCLFoSTDs3F0JfvEIIaF6lYhdtuwEQea7OnPMMOqLIqO2RMH2
383/WDLENAEvwELTZ5pgN1FBFbUv3pcEGHflhXNnIcUwn/MFkyVO1eil304DMyPw
IVI3otiHM2hkDiRi0svwOvv2u41ue2q2jCuUx2pssNormhLWTS7MxZk5YtoiiBUN
D6ZQ5Xzd/RxnK7YjMpS5VuMXQkOTZZO66pveVfgqwYp4KKSVjf8obFtdXXRDkA9j
r1D5/3a7IJwKcjl8JwN42+NuIddH+cu0e4JOERLFHkcDbHV1wJaO1gc9NucuSSbS
vR9R1jMpJXP/WMl6xEkLt5vCi7kpGbEk43MmZpGPb7zJXvSkwPhuJKujcghaDgE/
WJmCr6f2tH/PorhI0rFbN8J1fxjjs+pHnjMWJuGCCei3KH9jdgdwUdr+SO0HK1eL
z6S/gpBfRuFqFgaWSLBzo/PZgEDksYcSq98I+UmtRw7B70awpin9tsSA1J7hP//W
QK5RlH90MAv5ui4gLghc/sHgWplL1nv9pjhoNk20r09vifMidBVKr17EYR1mw1iY
OPEzcT0DTb999BCatZ7Gf7/Ad4fuBHSUzpvlsbBBW1F6b1pQBBP36cPccYfyHai6
2qfTIoAqyTZmrnDCeOuCy2EWQgVe8rNoiEZIlry6BpCKLpWgWRFSOVb4Akx4Ss14
lNnN9WgIBoojNSLk5cJ3vXMIL3JVjHFxB4FaSy1eEtbwdbUFOuSJJoE6Svw1yfvO
YIw/H/6MEfSsfCHstDqS1ay8MHfSRLyDP3fHeI/uNCwO70jfDzIwfLPJAGmqBPGu
5dRXdJxH6GapLElmUzp3cgXf0fami6ce4n8nEUCCH75ZX/1OmdJv6kx4cgp5bUHY
QC10yII0xIHmXw+giobGbjTj7/bfJDOWRjxFDmF3DSRbPE2T6gXItnAeV6YzuWT/
8oGdX/OkKn75eQoH44hMR1TKGy+BRRYGjn7lChtEehN4GNFyf+BIUdWcYmWz1Dv9
ElxMsR8ypibWBp6eAklwsHjRxBqa5yF7XX0LD5k+rHhC8vG1umbpHuva8kvLin0j
wquNSjQSHg+5YF3wK/Ll2y0yEfIHdFNT65IVwDsni/NhVV36xWBHKHMBYsVKvpv8
X1gEtx2S73EfyIsqQdywOd5VzYiaq4GwOOkXg8dKF8/wezMPL7oZpFYEMyZE6iC/
blFXQCMNsoN/pVK/5OTDBhUYALvfCd/Ozch9nNuebHJaS7iVLflF9u6pv/6a2pPR
qfvKA6sZZxbg8Q8j9Er4pJbERro7X6EWTUp2FSxN5FUPso4EBt+QtCo4qGccJIqS
MmvYlXGXQuDoVBoFVStbUMpki32DsLryA2ce/ejKPJyVrI4NMu4hlO8kRfOqFgWe
YLrUIc1eMYZSrzHndJQwRiH7ZuTmBCVXwgPv7B12nbcuivGorb+m3L8uGbNQx4No
vamAdlDy8eebdo15NWRyDlAqGEqg9WbGwzgYzc4YbPq8bGw+H7sy/uuOf8mYXHof
0pfpIK1WjB4Bmjmg4vNFIu5cMBe+7Kb6aVDum5chbj/4SKgdnjH1XAM+W/BUSB+2
VgHLu8B60Ak//ZkXwBtrtP+AHwiZneBQz25hR0O1DEIEgqGRgISL0HsZB1cJMaBZ
G5fJlZY5/dfxUvT6dGUosnD76PF/yS4RyzP0TZKGYa+cbyQaadBRtDT3lqo+vK+/
J7BHOO8fXiINkDeUn37dLdOnCdv1kSp939nKSrJ9Ng9papKlsx8sW3+mUXMa2cyW
1yJR1N+vn/IKdGksgtzXRNXCxvMoHbc3tMgFefNfSrAtdTuWtE+A3RxWo+2HPTHl
u85AeWX4T1Bf6rRG11uMIOLWWPlO8s2/5pM8Jx9d/0h7nkO64yl5eQoIjAwaTWGy
t+EnThn58jrOT1tTRzcm25UCzAUYlWKd5n9P8vVxBwGLffPDL+sIvf6SpLnm4MpB
hxZ9MJniZbvDtw4GNLdxx6fcnNeWQW7wujo/+61YqJy79IYvxgW43TraN0bXoYUu
eI5213dhPdCv8FDQQMFot6z2d2dg4qmBQUz/mRSTs2OYoVHK8hpiSnN9J8aycj6H
ffaTP/2XHvdI6lx8d0htohd9Luhz2B80FCgvepTm20I8SYvGzs2TbxFy8lPUTsxw
0w9MnRCIbOoY87OvDbwmFs44bMD31dxrijS8ot2XCGFDnYfq9/SM1mi/HVTWh6cl
NqPfw43zvoO5ZQRZPzfsgLfsoJ13TRwSCejrKDYtljkaZDDwGvThAI2KtVBZ4daQ
zWRL48SBDaYmpTfOLE+ExztEJ6lK+Lj016eHD6uN8UL2MmAfiyzlZwz+VCE+OyeR
ZvtdnrHE4zh/8BwjaODovbmWPXg7R266DWOG8LzScs8heUdOGwce5bAS6lvRk1+e
MT959qaduvlpL8dY7JKEADmz6CQK0VNHywm8lyECuBydBtsC5VEqIyrjLlGGbgwg
PfS0vK8ZBhZxEmD/txa8F6jpjgFwFEXd2FOJgyUpPEdlHBY32tsu/cjooqDGuzs1
+7w9NWr8rIF+ee6s4Tzt2BPD3mFnD6Rsp0i7ANN04+8z7jiAPu1jQcTYU9qThvuH
rBRNCJeSvjPUv2iBjGIB24NKBpnKlzXmSNFW/l/4Z3RrYwo770VGmlNKTLO1M5zY
NehrdWqEw6bveblckAdkg/jZJjmOi2/fGcwuEnwAdCFjjqB4c/jRwAM2vYXnIaso
RCC0UCR9QorVaVm4fnJgxcoi6Suwps6wEACy86DHS5e1f5I3SCVIfGofAn+Duh+k
8NBOrnSAUavDbKiJFPKKbSDgqW4TifwaLfqTXNcEuI/grkYtVkGox8CvjdF2zarM
4VoHDCc9lhgNKMoAPVfclpYV5PsmQIbrkt0NaOFv1YWGdQ01KCwUyshaOhZUxYom
M45MfeGBZCZkjX3pug1ZFePBcPFtutM3p3Ur8Ld4+4U+ad/S7mdyde+p9ktUt7So
HMrBtSvffcuglTLScKoHTOvRQeOIXx+qadNJYbfKh/zGgDmfXirs4fDvClzujxJd
YcwQixgUy3p638/KJRbnp8ZTqyQfNpsUji4RJcZw8B+tC15SZjeiUqrHNt1m0sMd
wMdiLYwZ8vgNXoV9/hJlHjmOBEcO3yIHlbP0l7tuLbXaPKn5n2y7T+Q+A5oeLmOB
lHt1Ou0RRp5FRqTlmTsf3c7rGOfKtR5ftioYR44lwu0RkPzlrTosmaYVPC7TRJM3
zpmXiyaDn2nizm4cJk5HM8I+di0vpb2NSY15j/kTcfgj0m8poZox4hblEeWVKQOC
kiFOLzx0Ho0l8fc+z5H/FigjfI8VIf69MfhZwTqGBIOYtKT6iEud1nVipMHYRdMO
Q9hHiH3w86U8EGunxl0y71UPxtEUZsEyDDW/OUz7VRt/k8iYKsuDG4CwH62RyGOE
9dqNAjaAHt/pUzip+8Eyc1hFs7OstiR1ZePUu9BrB6adtuZj+dqZb0hAs4JK+JPK
dOyD6rM1qN2rV/VyqBIPA0cLyPm/6v/rwm2QdapqyW+tJXJVmP/CCFBmwsHakCPq
cmotcyRIcJDJtYi8hF2QOtNQXB1WJrKEwlUdFdJEoxQC/uXosaod0l/EbCiT1adY
1kftA8yDGaFpyLsQLWsR9eciU4w4RehtJN97yADi9Y+PlyJ5rTRR7iAIduNWy8Z8
ZAIt25/cOCevivX8/UbtWAmAmL835KO/bbAPSTVRGQeIaOZNUyOnIfoAIDxtJc03
95JWgYATN6G5s26aIaoD93PpHSHKqoau4V36qLI1N4AdS+6sEVifXABq0T8Jfors
b+QsfPWTBK2DlsIm0VZDFxJSu2qjZZwOQ2du4H2tSRVskUfcvAGIgkkdJOeGlD2G
nmxcUuTDWDUnBwHBMvh9XWyF4QH1RRlzBEpkUz0GzAHsMhzvdTHT3t5d3qkCQQ2L
eitn9L4qFyFQP4ipnuF7R10PlmGn29gFNLbAPdWCRSUWHcjMok1oDrGZvayW5ET8
7au5HbSs+57PNC4BAnTJS9F1NEhcegyUDVSQcrY3WW/DvDV0BIErJiGOC4E70MkK
Q1F8jkuAhi/srcOY0Pty/jG3Z2Zgv4kFZHW35ANeIM9hQS1CpLlG27PmeliSpMa9
+3hqQfJsJSRnXNIOzcKhC1mXFuaimVoNiadSFPvtywrzXTQDcyGRpGLR+N/MALe/
WYQMf8preu4ItHqFgovJRWTWWsCUxDg/8PWz6YjxQF1rd8TNuDDEXmrmZf/DBaI+
U2MPJ5e4NlMWylyZcjf38/eJ3Ac/2AfjpLDZ4s62aFkhS28ZoqdRs72AZ4S5wLmh
ZQVMiEPFqHbB70c4ZM7IQTUmH+1lQdVcZ0em864yxJswRpjFwAoueSZIlJtTFEM+
z2wR3sGZCozWt5sBUubYTXD7SDDmtNbVU5l/qUsS4WlkF/x69U4pojBiI2RM3wcs
QXM0o6xG/vEM5O2BYOGrzUdrVcJWhybpw5XX8HNPzvKJc8JKY8yK58QozruXEITP
JQAPYZVZGkWSJQ3ZzxvZsl049YPQ9oSNlgIU21MRGtpMls4MdiFnarp1ZMr1r+s5
TdcLFxp+pFXEMIdKXQt1Tvlor/GFHdvsIRDddn+hzRDEAWqz0u2Kwo45jMtuyNMb
4uxWiiPQcyYlmGrmKvt96D8j1FT52cYnGBZKlWFKeHzGC0fZRoPJUsAvKvH9UMZg
3/ZqbP3ixoaDswAGqArQ1c0J0zGKVE6lP6Jhf5ALeyffnl0Szn41aoFKyH90iyNR
zYWjNOBKnGDvKa4OQJo9VCK++xJDdlVcK9jeFTv7KJIxV9u/XUW3QefSSUQfuanB
Vpyp1g8yoJGF1t68IyxkKOpno4jYpgHWyyAvHreb9SwfyJaIAcFq6raCXm1zAHNd
dzPKCsOOoi/NF8bz+N8oe0bBWGrJSft35WFjwY/3whLkWOz9npS2707ZkdBtVBcV
m0yhpTO2iUmOSs2b3sHAgu34FXdAh4A5HNsVY9Ju4LHk9aqEDWNzeHLQgZUpO58Z
wBi74FP6WMQmrFiVr6GXhjozxAUyq4fd6JnLVjwBwsFexNd2JpvGvlmcOoaxy5Gz
kAeFCpT+HeqVepVs+aG3EmoFMK+PR7Hcw+DPN7CTMkEXMpPdx4Gtwm5F/8tCzJcF
HLmIXQ2P8eSpg34dtV3tibFrfxuMo6VQX2vTX9H/0ypuRqwn044ud4ZTsXx83wwA
fuoj4josXBXV6KZxqIgvGPGsqhRG6urP6YQ7yPmCPQgLdPsdXbKIc1P420/1R6de
8N7cei5iJZ2X/gDyREQ/pXKXeg5GrxO6z/52TBxk4Q55QPLLj839xlp0aS3tlBNh
ow5/R9S6ShP5vndQ8SE48jjpKiPFMzPHd3p9EbAOEEiI/uyAjmUu6EEiTGyEw7MO
1ZaII+B0dlFWnlaBYRFOTpMVCFQXuJamtwVhwuNLFknWtRnq/MtzqwMGxzjEJqkf
XYvSSZfFJEZ3HmzD8DSuRwkOEVgoB3UHkYKeguUlevkN9qlAg4s7D1YBdw28YTRB
ampMWxcajQc7rry6IP6hGrIRHkFr8NGTw9rRQ/b3PhfJvW/DqOjLkx4qpH9YTeNa
SoPuYFIc5B0UxsEFORl/TskdYFz1VB0pl49PO6cx+OMLHKKWwA0l17jLso2mXKtF
sVA+0QYvObEWQrKgFX86A0Zon7LvimcIaYC/4o0Jcr3xdf0lM5E6hPPBtHw+ZzRH
PzPdKDI/E3E8SG1mQys/5VnFExL0rTDtuGBmJlWIrMe1u2O4nOGcENG6FV6WhDGC
oSrlet3+sZ7q8dhSCZQTKlNO5jAM44gYeWwVEH6XY7noAnmGZtrVWwsO9Um3R7T9
Z2Pj1Xi4/jbQsMyr9/p7NJqj4CKEityMTjzsxm7mllrsfWCs4EwES3cTIaD1STP/
GxcTTw8WTrsFPaI24v+ZLo928RtYmRc5OqC6Fuk3AFjGGeuZ+LcNsS9l1k9Sk+J7
mST8Q006Slj6mjb+7kOvVEx43cZqiKXVtbvT3k+S73Nv3ACEiOFTiB0ZtcROnRHW
TCU2x/ZTTRJz2sQka/lnFDeU6YE4oQtz1HY1BvNzclkUaFdjkq0KhTfk5ac23MHR
DIfCd3TnmaUDsoh6X6/XVw+mjnZ/RP+rP2vAegtL+Z3ndhPojIL/VMoM5h/QtKUX
oO9y/D6FBhGE6kjqsxKJN/rV2707ygMwOITHSBE3sW1HlQe6OCpLRZTPebbSLwLS
FdXrHMKuJ+6GdO1K5oF7KbOwfYrzx+4cvgip8dhTLryVnPeuSLgLunuUBdHfExk/
7oP915qTV1kNkZA7jvTUR5ZXaT0CoQg3F91BmIaj51XI6ntHWcYorGFfN/ogsifS
lTNK+TdO36rQi/j5HBjrR5s0atjI1EE4pGw1+FAra7mSeeMmQ1FVspEqPacyLSos
GdRnFhL/CD0aFhyTtRhfnfGnvQIXfEMBwIM2aDJN2fK+LFawmF+qgMfOJyiJaC4o
1TYeEIe+o5j/6aZKxLvu/o/2Rwv1QUq8d9x32GtAQbUTtDTxbX3CqM9CbeRFhLqI
bwnLRwAB2GuPZnA6eoSOdwQRObTMkr2dJ3NsEtW0vwBTfH7vGQsWHqf+htu2pgZJ
0vE0CxK+3KBNirGF5vkcDRRVU1/0nF4iSLJSqj74qcf2E+LWNBatcKwWJqHihe9Y
Jgd4bsndIpA/MRbpLHpXz3jN2f25CmxVAyJa5Nk9j6d2v7o3dQOLA8ByVcFD2yi0
IBEHIrpBSh7QjUgaG0Y3ATl+dKFPAwFNPFF0Hhsf1uUWaEVmxC8W1/jvMzNnZRQa
saFCs8VBI4AirYFofgQvD3rSzGq93liB+K075NgRoEsFFwjVD1mhCAQwwgaCtQnh
aEFuyfsx9seU8/4YjnVfJWtYkvYtte89L+Mtl9k7XDLRssUSpGMY9Crh8cYvFxK4
dSXrz0owuRM8dxn6Or7NfHs1Bn7vuvKiIiwOuLo4+KLcc78czmwOShZGhUIbbcbG
6Q6B6c1KdbMykBbr94oo7zhZtyNd2qUK1UIGI9BHn0Xg9fq6yBMn1X0JWizrDUpb
/ZvqF3WOFz49gioJrVSGsxw7uMSkBE3POGQXC+znyzRW7XMae/TjoyFRwoQwhaR3
JOjOkS5G5pk/QBK+vw6wN1GPOiVEGljigcAQUApgBglsudVU4G8S4Jouis7jcj5I
QVF5EdZC74yRX4EiAYZg9zro750iv1ohiiQaY2wRptmwj6GI6eRUin/sM5rnJAVJ
fdNIOoc2vqIfeFoAtSksQCVd7xjqeRw4SgG7m1GtmDd/NvIWn0Gj+r0UALwFjRUB
RUS6n5nqs8X8g09xo88cEIpLSEJyhNTyIn6oc/wXIJ3g/6t8XcX6/h8P8bml7c4d
gAFdPkjbwGJxZIByrpdM6vNDeeajFePlVoibop6M/TDfJrYsYaotcEcFNgzAcF7n
f2TycSwg9EecqlPtTSuVVej4D+Q6Z2fpjOalkcCBeds4Zok15BrcrcQnYZYQaYPA
kQJrSHGRpyJ8nwY0sY+ESxXH6PBq9o1Zmjj/GM6wLr802suTW62FMFYHvEIkmD0A
VqmM0s+RJdUBrUyMC1HqjrK2OXpAH2k9eM2eMUfqHfpkumB0yQUB8PqAKx+ROdPV
VguIsx8sAyahscvWlcqoG/YUePNMCTbFMbt+z+4oJ8jUASLJglFU71ENsBn1Ete1
VqvGPae8tzz2KTq6iC2FJRyfhJ0/TPBXKudSYlFyy//Wb0636MsvnsdPfHeREsgl
szMywgwW66rREyPn3mQNzygH1DC+HMUXtcmVtf0mTDiop7vyAlrlcHIj7nBe80+8
/Hvmlvh7Rjbj7kd5Zbh9i3OzTkpM5OGQL/wCrbn+CnF84BlOmwef9EGTq0IJoBO7
PAcE7r3JCrLLUUDgF+i7WA6EyD99uAE+wk3+tJadHZkJ17qfRgfAZ22vLAHhlcin
VVueyPKfA+RA4gaxxcasPYv2OPA4AHZcFeM2vJI1o+/8jNGmGG1Hh9iiBz4p1HiZ
YnnEaqhdfn71PPaVLKEak4qCCL1AIrVGPm3RzZuTHXhye7IyqlgWko+HIXVohVQF
cMPkGpUhSCwf3f+PDkXxCwheDfukNdZY+fI1xyuKgf0wIWmCE7Co4BzY/EJFjneP
wciEf9X5u8aDFAYUTEqrDkpszf8aoEidcpbHd40joOckoEwnOyKn86eMcB8C/kRA
6IEhQgPogSCgVKtg9GKhAlNy5I7HHTja01Wc++vL2P9NN5+GXtyz76pOPC9IrkP8
kwA7j627CSZJH+t2Y+iFwfTBnILnRBXzWAH48qTHelbUzzhIWt1a2I1Lcj5ctjR+
sVdvexY4Ja3tcUWLyXhaRAn+NbQ+buEoS3OzmUUB3blsn9I3cm7HvL9kinq7PrqA
Og8Wk8zesJKCo5oRpDOnVUZH2/qjXrG7BTmGzvdB/ANnijhysfLGIxnqpAX2QbU9
SFAeILwbZVrB/tMkK+F8gfMePPOoX+2kIMOt3hz42ShmPsfC8L9TZUrwzLhKDnhf
T/c83mfVngNZz8PUm2KpHT1TIfKfqnN3uR/wMjOeP74eqi+Q73FDZNLdLc7xwqDt
2nwSRTJKUd9mgpxd2pzWxNONMt8Kn4ouCHR+bPUCD71UG+xhlMDzZiAhPQqbKP06
cK/mwMYKY0PRw+yKYXSKZXd6Hy4jeTTdCuEIIlaLIMBc+QrzxvQCYe32ZfM7vzGT
VrLi7divp20OeWKwwfadM4FhGw4dCzI4LjBFkL6VFNx1gCS7EUvxPCChKPQNXMye
x768BAnngdo1G6Ilwvbu02K+1JT7NSPyj45XJKLvU9eMBO+1UxZuyCPphqoMuajR
v3V1OHF2w5e0BzBeXRxdNa4xuWX6+U2xvRE+8EIU1Pc9UlW0bxrZsPK0QbhwW+j4
6uujXIirTq4SNerF5dG1smdxz+v5GAm8Rbj4Mm0hre6d1sJ0OvrliKlAOdY2AhAV
TyWDy1NuPIRlb6OE9bYbR8UOw+XwWIWA1chvyTcjfsfpwdwqTv9v2qF80lT9xO2L
t6VekIJrnpnSrxTt5RwVzZRsyjTq9SbqaVcIbnKt1tR78lWttKvugnBKaSJVrm4V
qvbmyJNMYmfZ78lS8i5AYm6Syf2mC7q52ozOX8vrt4vWmGxjrLj3byfAjbwwiqKB
d090izqZung1XuuyVTSyIOQxUXUEuPbhnyKB74fKQS1oGA9bTrUMDcKAYvNO1VBY
PBBQI5e2fmS4Z84cTsqzrrvU7g2ISS4f3lrnepEX7PaNrG877VcC8MUG5jdQpi8y
qxyfIJU/q9pCBtMZU91uJqlnmht7uV4FGbuR+FHHQvMYtYKr2G+jIB+djHuUtWSg
3woVGp13g17uZI+iliRplNuAbxuhw6HbIgpVM1Qj7MPTYYVlo0/ZhaPgpAIpF+Bs
+Am4zYWoi1ILJZwjePVGVI00YwzAXzFahAo3D5tyU9sOWbRdWEgF3r2zw3ukPOKn
6tyQCoLtbsNtxK89s2eARm2++WlrVo4coY94u52dEFmHTevhDIgz+frY011E0RK8
YWZBLkIagGs8v7wcIEHNBHGHdpvfVQb6N6LoQ6WUuQoZWT2rJz6QGBR40f/gN1BZ
QwXKfY3CO5AF9IwgvYf6WtkhL88p02LdUmh/0ZWJs2t51wYElwgOLT3pcDWd8HAl
HNNHVM2UDPbTE8/FgF3FKIPPmZl/nQ8/9pWQX+jlpZuhQlGcrvVkOGwXl3PiWYQd
Sijb5ChNcLsD5SgyZMQfUsUogDJelCE6P543sXMzolVk7QQEr5yyHwxDmVbmUG7Y
hyfhtPn8CQFycni/so8lchbHCOz8erDIS8KjMVt5otEzZDlwOvRu4qHrqo63i627
VLH7u3SgGY8mJ44WzhnvGgxGRnjSzSqZXHHe3HWEPvyzpcnB3ANg/k/v4lmzkOPP
WmAw53XfPORsFLVtRt6x2MUALG72BqukYnYvm8DU+rtRUyYf6LCaUvzzxrssNr4E
dre3LavFdGddhhsYLzzOgxDcntxeigFTbzw1vDyvO9jFtAX41vAZXUNaRFHE6OmP
5l4clsRQEa3pmKnmr65fYIZhMUHNKlgEPKNQ95UmotXVZHRI7tFDqFqZG+vMjPDu
+x8oyrZjbhl4OegCDGjJsknlwrstcoBKvWYyaNkkEBEMj5Xt/RL75V9BtVH6VFt/
qeooBGndsf/szw5OQWkZWc9RHBEtwkbpRIeCEJO6BwusmaDUJnghiex+DZRKwM7Y
XrBh6/rKY6mojJAWExS7OQCTfYp/oDfhA7KoY9ulLbEHTSFo/yPqOJDGT2NSv3xF
SE7g/MHU8VpNnCu+gXiiu+deZ6LdC5sOkBGIyrqXgfV/NheU2Btwtokd/ZYCNccZ
LdqGImqTUIdGQ+/3P98oHTib6LjCFEKisahl/Xcag9xNrqgf9Th48zJszmW1n1Ej
9nGviOdYzkFpPlO/150DZB2Q/Bk3BCBd847O8uYGpsyVzMMM1w3/A3x8ehwqKPUR
Sa8tBTPP+7BP12XDVbimYgbdEouHIdb+8U/WpMioz/hrSgnOGOIaUOAvevFapg7l
FM9ziNPrrDmcUSzKHRVg05wWq5cLC9T5ihA7/skU4zgkkHHRipSgMeYh31PBP1gY
d5I7OVsWAJvy5MxSXxa9FMNZOV1+fThZVP/xX/oTsuyEoiT1Imd2CRjC84PeqZOu
oCZqI+hXV0/zmfVOZAOpSkf1Iloc5oRHCRjeqVLhcQC9rIn4yhdVKwizMIyDOJE8
aOUPQrRL0/XqKX65brwG5HGcQWoK3XCAXwhkdBQDMT4ehNG2JEtiCOdIs0dWgoBB
7aQUNbyjz6RokRQ0ytQGxXRqB+bxI6PnvpSvVo72bu4gSJSzB97HzzXS/sXVhmgv
3215DEFW8Vr8GL7B60vhCsLm/yyyEypgFr5SOAi2YHhrejkgz1GVwADYbMsUSrLj
Wto+BUZs/No7Lz45O8MXKQVgBIwd3235IcKxOYxPBDiByhz2CxOaFm6xUhSmFJ0X
UKLc9Z6XjL+9s9SnBmRUy4FBDvl/hZrJehYkIfWX9dMSpN/fIuFnPUlAnfdZ5k6X
r5mno5r486H4Cw1J/DgaKs+5TyOnww+WTWWH/eTkwRT4bmN/OIOvSG3lSX+q3lpk
Gif5pBqQ16SKUhpnNaACt/YhzM8xbxj5BPBgG+cK6sySPb8GuQSydtfG11y4PmKF
WEENmTW6wg218rX2jHbwJRp1Kd3kelSJgQCzhYJs0DmezvAiVuzqbAwIiws0nJGM
4uCYjsu8SXjLlW0XS83VQS16c1omojWR9MVTf+qWrVB6eyNIoVdlG4MA6MSBpCd7
DWCTRg8QIcnkX1ZchzXzh6yyoIg3qHFxFDPJ9s2rnSg9a8IuNjRfj8siNN3CdQFM
Vo7dEfxqUHLL6RXjx6LKh8ZyysOLPd0Cq0+0rIczoaRWuYTuuv0KzqZw/1aOFNQB
4WZCRqpfA1fpAuL9hcaBtAA52NlcSiZKteSCrVdu7S9C1UoGQR7lv5bYsgq5VKDM
6Pa4JC5uBE5H3iwe4vTLMUn7LgD02ygTdj6VthhwZg444WsasynxL6Z4A/I8W6+W
zqmepGzl9zoaNd20e1/6afsP7X4dKiv0aRQEXpeSCDyUAI9q2sEnX6iyMfmf+mgb
XQiB/+zBX87yBhwZRmeFktgInLo1/eZ/GlGqDRXA9GXWJkSJyhpW7OCJYXcjUUoN
yMnrUCEMIvFoC07q8v6N2qgNtVG+ObqpORSS4AL/yEbQYyNLBG9wpbKUKwN+tjsX
8h4stLJ+vj3LprOyFcRteHdCICWdEFxLiuvxmneL24KGHAng4mTl7+LTnMBAgLlI
SRLTe78Te0MA7yywF6TeOk0A/LVZ1S5R7rCp2ekI6OrqO6dYvMv7zKK0L0Mcg+Xa
dzzI6dQkP26ttjdnA16rbzvWf201KcZbW+/Wyu6YF0JAE3s3EUg+qnY2bcPZU8mJ
M/pKQVkGQP7fNY6z2ADwvi66FpgNvAAe46olUJ7wNz23wT5bIilsR23YBxbq/jKv
RIbTYSdzQWHmwIwWTiyEKwUmXZxtu5RQU+9UbWhmiJsUWPuHpjnwniXWZM4vR/WX
a0wQfOZb+5YaQQ86JFZ1OBZVOc3vF3PlMn06nfSoT5/cs2FmPZLK4J8usEOQRX5w
Zx3zuJI44afHm6yidi4+fVDuk19z7pQ4krC3/fxYTTvYxm/PmLReZIpxPOJJZf27
Nkdu6fSeL0eL3Vscw8a1YTH6PwPAZUOLyrcavKIVG3IUrt1IMmNmki+3XFZ90XAc
T4azasKc/0VKV8QCSEvJ+7lwtpPOqIbz0TUARAVzPGPFzalWZotUwgdNyifyGJoV
6XCgjp4fLqG1xfsOooCEoOO1Qvp5hXaZQyGlueuP3co7xbWUP3pKaxim+vWhzX/g
pEUWOhRYcVU/20VUJFs/jT4RA1ijg8VtphUWYFzA3dQD56jLM0YFK52N4Pch06z6
m9Tuy0dMxU7ApU1jG/pvvZGJn8moAa60+NZ7uHGTAbDozdpDbGNsUXvdGzVTZF6E
Rm4MYCWtqthoYCqAdJA2FlmCsiM5MTGzgJ38dte8OEqvr337E2ZHxUjVv3026CAu
X9pRCq9Kq3VKRJhMoHO5vfhCoANBDXj+Y/gZvETv9bdD6yb1BYQo2wmqeVZXxCds
LuKigd9lIadCeJUeCnzbjuG67RZheFl7c0y0PqLnue9YscjRPdnxyrkSp6hDVicJ
fMMxZHvgA4Fsy5bLvf7ENup7vEr6hVLNaCvpxWthEonTj68bEszDudeYXi87H/kf
s7T80LgoTGT4vwp7oNX50+6AQsWsRJbhn9yAqe12NSsXchxPe+iXXQdq8JCM7lWU
unIEkkNtVax7m92ja/uxmKaMw83jT1S4y+viDxRKN540k5OiZBuOrtKmgMsa/Naa
rSn3qZNqCbrjYjeGi+6RhEmUzargPcHxQJ4wUexqr1VLjCWm6iGLQ24z6WMFjCjX
Q8Ht7Q3jCdEkg7IOjs+G41fi9xj6quU1UjcfSuVBUKBjBUhxMiAn3i7n68AYeShL
IMOkAgtl/VeOu5WT1KjCVd55q22t9yHR5uXTlaE9aOrKGES3gwiYYUiR9BVvmlgj
DoK69hlXSE+7USIaa03fCefU2FdlUwdzUYhKR0Uu86rODhAiCPKIGLeEAQL8C+/U
Qkyx+z2/IemiGUkhLLIXUIRimPo4wbW1KOsTqVRZ6fWVNfiINgXN92YKSeWFg+Aa
QcC6Hl+fZ3Y6mE6l5M2cX9W+Z+0IU30X1Fzhs1yFC4C1y8rwJJ0MlNx7znKd6MK8
xfV0Hl1ksYoCC6WwRhpzmJBVeW5v3+Ax44QOZf/02F+LBRWQWBb3hk3CO/YdQcxz
dFKe/6ChFXwBDJmXGREsAOF4liV+nCo58kqPHipN36144N00mB6HQ2puVMRJ+Hgv
4GUUB3Vdz7qkcadNtOOFaK5d9WkXYRzxVoJ4hk94Ae1hYifArtlRozP9yERUFi+K
YOdBTiX2UaJXrIUQaXDfO5O2DoJtzo4Yf5spk2v3yL2ywUwIZdSqUh3uN5mAIfp1
rbjFRQanbn7DH8lSotQY2RrI8V28eV5V723Ks0vutPA6PAUc2lw/ksSsGhd9qMxr
LxqT/Iv/RmRhgorH6c1tMrPM2ov7vKn3/p2row7ItUZgFo8G4fdo7tut2YpbTQN0
vxpDjLvEbUXixgGLmAJlzbJScDJAwE/NJIkmSASXFbGN+UTObhBTPwic8wh9rYZM
zVFgcBaoJB8xwS/+gv7zIksccPq+UA3eqxyueELp5x0xFBpoWdTyjEQV3sXFh72N
rxapElL1XMRwvr5sGsSPAi6IGsW3j61ha4sDkz3iKRAUPonQ9oxS1vawX3YiWfJU
wKuCQ92KXzrWXPhkuEYVwbOG7bJmOBgtXLL+qxhv94B/98+PdekjXi4/BReBaelv
2vWDhnA6BqCjup4IZu9kXwZDBEWzDIi/cww6Ll1GqDfzVb0Q6UCacElmP/sHQxNP
FJR/JCb4KnSBzZ8UMeWTKamCxrUgYYN+RV4k0cYKMIv9K2UYwzEXytHWfyMo5ejZ
MNpaStgaIDXCGImK7xvs/Cx6eCsZ+XMd5jWtJWEr5W2Y9pf3kRhy7ABUcPFgWbzX
AR72fFZmTV+Xpgb5UCMSmgVv0EsQrFn/dlm4spLAifw/Qh/P/U1TwVutC1SktN30
eD0AHAFpPGKxgXTRtUy/W6rIldvxsxu7k+MZWYCxvV489kgS02p20oKxj0CuOM0G
7CgXJ+wOn3FomZa9y34bPAu8C9dSKtyqParz1+Zdz+sWsYJO//SN0epYh4IOnLcs
R+oMVykSLIm0N88NsCW2j3qZpgEdVNa5q94hycm/LecgdN5f1itR4T9bvz49lXS2
HxCYN8uv6MlMh+2u1dWmNOb7+YxAq9RAZhctJx8wq/dBXgOj4rfFo7DUBC7aWOPX
o0BFijJGqxw4vDMjF81kFrZF1kjH23qWszKQnsL40WvwST15XHzLONS9tntY/MfP
T4D8RRmhA1AdSFH/q2+IOet8yQ0PELm8HvOWQwwCfXScgCrYeZYHCCFggpkmMQdt
sGRpOWrIG56hW4HkyOnnmSGUAllHlNnAZQ7xpm+teJ186BdgcXxNNpjN3AL51bCE
fA01Li+wd3oAtBSecpDkbD4YSgszcdKXG1qknI686ry7lrYopgKmXHOVjr7ZFdgE
b11c+f2m3ko/o5Eftro4NgyekhAK9DOIsUFphpfDhAsJJO79ROBgugLcM4dLFOmF
lhO6CJPQkA1mt9qPHEvSYZ4ycQUEuGVEvR1RXX3ib72YjlsCb3JBV68F4ES9oCT1
Nrz6tsCrSi35HfwPmPv11pd2Bz1h04zlJgIy7iY2Gsd+FfwQwEG8u0jxSG9okbCd
snqsqmPwNfwIm6kjNxVwhzGuJkmcBuQ6TA4nRmcHGd3ZPTGJPRaXZSN3gHTTKQIK
1x5uSj6PLuWq3e0Ky5T6TH0iRS/UOzz3wN/mnixu/2szJ0kPr6vdVTTg//o/crB3
xGy7GTuOXc4gSREwtboDjnuy/glDmTVA26NJrcdctwhCaNXmd12gd39+vfEK+E7+
q/Kv71zZakzsyqM4girSecsRa65zRtcL0ZfflJWG702AY/smgLFciw3WThq+0BkP
Fyf4tyZTWqA0iIAP0V9wiRFj4/6e8bJwqf6h1BaT4HVNGbYsus22I77LAtezBr3r
SeX/Y8gyQpaDaAJWHWY4KwlptylsIVi5Fab+TQ5yP2E8DgDRVigospUZRugMR80M
WmocAcxDqxBs71zAPmy5e4+etNubomA1Yq7w4Z90mI6JBRzsWVmSHs4/uJ4OlMqb
TqsfDgRHm4flaPSwHZ5CjeuELR+8wkFzg69T0z8kvSAySV7Iivw5W7TkauA9HXkS
l6fd96Vtku1sI0n960w7BGpsglhnDbUE0QhI/kQPQJQK9JwbozGoDKhTAYGmIquZ
204swfPDIr9gcdXdAMYTwNqIuQAAHxd7JBWeE6e6nz2lFz9zQNUoRXPdC9QRQZ1m
ml5wjTrZTFrRDDI+Nv+fldE3RzPAMGjjqr7i3ShtnBIO3vx/bz5CI229TVgR1rhp
Da9zIkAtIpR4F7i75J3mRBL4s/Le4mCxiF3ewPHbLhZBWhYf3ykOruGapkmJrELq
rcTqvOPIL9Fb4LgpUu1jAo7FbFJ2BRPCchcWhbUcvB37GPR8K5f9rN3kMEYsby8q
2/Qh5jIOAFMcDbkRgk8m6lWKeY8SRpkAAtkjyAS82+bKuspy0EY5edVgxdh1cDc7
3SGZKYT22hosYOiyoq/Ih+900pltMfnA5w3PwS39wWFe9qMhTVIzWN+9YTfiA3Gi
m+D7XV91kTHVEkjhXmDjI46Vpljhf4UOWWD2tTuVj2dqXldgOBPWDzTvJhxyfpMZ
P8BnEbNbiNz+nlqyTy8UASCy5ix6dxbIC0lblxe330V0RafxVpT9C96rez+Qy3z5
ZEfJoevKHxgXHqyDyqkt7ESUTHMmQL2N2OvscPfnCaso5gW9i7kBYrcp0fxzMgZU
pYUhRhANTsiCK7EdtiDqQVVQeNYcmm/igi+zI1T2bd0AZCVBZLd+s4jPccm+yHL5
Noq4FUqYjC/Y/aP8SCwSaq+6KAoQhv6Dla/1x9s+9OfI2we2Kk1k8DqmLh2spbpw
SnQUxQzknuQ2NJ7WPGERkehLDzyk602q2uDZIC+GZE+U5YUZJScW6JOsnFPQ/iPL
mQsLmLKk5XUnzneZm2owW/HP5K4ld6ETzWC4D6fD4ou6swUNu3HIYDZbEIdrrdPW
eHJTSIEjsVfhDf5B4+ZsxnKEB8q41et62LAiTQsOZhJH959GB6OPzCpvA2VjGDNt
ibbnYl4KI9W191+mYnftnviEJdrFjlPx/t+uiDZP+Mg5Epbn7viduVJR5WVai6iP
+iSAAbhE6SLF10/Nn911Q1sc4kL1B1kXBbwZ53Od4h8woUlEeDV76HvgKR/h9gpj
+3XqUt0cZ1jlgTXQP3ctufYw4OuwMh05DEuytsWHMGHbeJqWQKh31xBN99kKHUR1
JKGcr8Fe3OwXji0g6bwR6oCwhbago//fDz5tcLqXDalnmMr3NvdFSYrw0sc7BoB9
My7eE74S7cs/PN9Vkws2Y8UiJaire/om6CzsSXTRDLt82yHh4i2NQC3wRy/PTj6F
0R3geFrjIJCb4GMONFHNBqIUu5XpvnwofylB39BMeBZ7T46Xa9rgWD+4fvUejZph
PDFbpMWeh/bUjsa61Mjia8rnrjxlITTCAirxT9+4+JjtvcjydZ7s3DSvBoRIyTSa
UcyL+4U10YVoheCkWyzs/9JZZK1CMgo2M1XduwFLiknJHwT5NMwt6uTvV7ARY7hc
D3f56eGkXx2Xw8DQkaeUDhwODgMppv2hEC8teBnXMo5Zkjldz6UtFodhDHmqukiL
KnqA6+24Os/yEir6w8lXfI/S7a7At92tvxIbtKHVDehugKmKNNGjH3eZMHej9Tbx
0WB6qmry3TJallnPsfWK3rRb9BmIkKwxKW8pUkg9utzt0iu+MDqXlg8DXiNTQut5
/mvLHuQY2peiiY6x1kG5tFAH3FvFa20FbCpXohVOM8+VAuubQ1QXHChgrXjHXftp
XxpU3q8hZeKIQvjEnn8zGu1OJbGApf7m82SOqSyqvsXjuUoph3rtFLEepvZKKr3M
nAOAW6Noz+Xg9Dxo6Ci6S1E2wb+tQKXAO7NxKN72vKfYsLIRG7jwnXYRMYNraBdB
deIrGmzS+onDM+4WGfDCQGfh+SA0yKoSbHHquxL669gLaKlOD5Ry8earD5LzvVrr
GvrTy1TtU4JsPfS/b6/Aag8VxbubVpJSKOZTY1kk3bgOANRFSX1JIgA1WWcMWtNG
EGoYHWHeXMA7O82TQ9OwK6g9m93oI9gsJENkWnXkrYgDWYjd7h/TfqS5BBtGxAHB
/W/NBFtgWezZkwkVDKonRAmXXtLi4t3NldDRKnJFNCdHu3ND4e8TtwPQP0t+u/yd
jwBPCrDoCSZr0cSPZPye1TbOz2n3SIEHG6pDUhOZY4IVGwNDhMD9WmIg/MB+mp6A
kKE5QR3Jm1tWWc/5EKyOS6NoxBPPp7kVHEC9WAsjXC5/yUGMX/1zmudMyn3OLdAR
6GlDmg0VinGlC7/JKbbk6ogWei5rCKba3wLccoxXC/5Nw7/QQCRAAUgSP/E3olr2
+GQ4l2/ovaTPToWCDPBrib101NxeW/7lMyrP3/t/Ev0PbcacZdPxSEOLa5E8r6B9
wb4it/DPgOl6Q6qyqcW67hKjjCEOEDLiFhRWVITzlSzeZZ0+fDnCLFqOSqz7Yd70
1n7LV4Ub0ROhMXdbyj4yqNwnUylIDglK1CEXlWoy2V0M6H5/T4dXRo7MYjhG4lo4
iVoLD1+7DRjrH0+pGf+wH+rc+8CiErcj943vQ3derfjzUvgpq/b8gcj6BmQmXvhs
5XbAx6T1XOvUUTNQVahsLnAwraCdXL/DRoqjp3A3gfkHqMBY9X7J1snIdhO8nZQk
PRy7obbAWR9AduB6XBhCgCZiZWbIu+pQT/GTvhKzwMT1bj0tzvgnDn/oFPJ+Uks1
qdJ3rcmawRY3nLODuqi47Xla6uVMHZX3AsD9eGObLAaODrb1zfQ1X0AaJ7ZBHVdq
MsrtDoboEytKu1HBC0K1OY+g/XZFYUrwWNcmH4Dk4dgLXYy9GDzuRAu0ozFAqFkL
5ooSf/4vyTmJXpfINpollSfEt9z4buU23zCQSTc4NQ92jmwluNECXMPCiWjadSWb
o33oT9yGqiGUSEvXcVer3vwZ/ZrTiWMEvwzg2VZbgqjeL43YtXTIfzXcweG9nZZt
kQZ/8jwI6v+DtaShVGSIj5LmoNpvz/+/mE1qUJOG0BMB9hO35SzLMn7/G3u/Cz3p
uSp9fiDbKQnC3bEl1lLskTth63foA0nebfqJSZYS9ty6J24LCukCPM+z0lAyP5hW
itsE2EgU1iCZgPoqYEM16pkEjVlXycPyZf8vAxGF0kZZQCacZL18XsZsnnn1oTzX
Zl2LxxOl9FoLJDe0lypvUv5bUGviItzyNSlTN6/uniU/+y8Gs8uVM/VSCGXUwEYn
sl5u+o2HXYcnWwDtiuuLa3ZnpLbAZbXD3dpYGEpOy2EtDVvbQCecLm5fWkrZmKY3
EWEcDwHoikI4gX56j9CoLEhUn/SZUZHbAOPZ2R8Qct1qkvDBuFoQfC0rt6in7dny
0zgBP8eJ6UXFEAXakfrj4quDWEz3OrpdVD3VhDug4un7NwlBNc3P0eHMj3B4jV8n
SjAKgYGUvk91zmU5N/KbfYI4VbHwvT3e4bQaB4SkIJ6b3fjdvIlNxHJVgY0sZ4Oi
x/rq3qj1yTavPVnsMA7ByOIwZuW+u0Xmqy0INGKWzPCAWGQBTtt3GhvAddwxnQ10
04IGl/FlLEkQGyqzl2YX1I6JrJHmeIPc8MFsrj4QBpZgvm0mR/ArHk8OsbblOUJl
qCMhyJjyMS+BeHqFOqVC3VB20XbtMZSmyMLHR22eZx8nlRpRYKe/LTb4dE6bc2KE
xACZYqXzF2yffvVPI6fGuvBASlaH28AJR3BKCXvls4gDTRz240R9sgL9AW3jMtPB
zQHyiao/GXJkKtnyhUTd3Fa9Wd6pv6PxCnw1/07knA5220QPRuw6zov6w9mjUqQe
9VvtgwZ7c6eFpaNf2szc0UUZ1ah63SZGkXQ5fP3QybDSd6vuUjzmmDgh50gCxrzV
38tAdG1BiA8vdgpWTuaYM4wgBFTulXd2ZukMTxH5IFCCSPyebuwzyvW2fel6gB8j
6m3+tnbNXUlOH+TfsFOT5ICJc40I6K396RdnbTl+kMuXgzF8pd99qd+yBjLW3FK7
6XutSi+KifTmnW5SlpY6uzrdYftYdAgQz6Ww0Asbp8GcEOrUwi7k7fLpcEASajlT
9dGiZqScXYE7kqCmmvQ/h6afgqTX8awn5lR0kvANCPYDkDRdW2bmk9K1a2kOylAv
lwipL5Qrj9E5LqtsCmWF51N2rMM+UchlmJwarXombSVjtQXvC1j/UV4a0rec0xef
52cn9rDZ0LZsNmFv+e3k1YVjrsePCvpOQTdDwtiUl0b2nI1up5dN7Pt0Yx0rJWG1
HRI9CBpYm2cvf7jwq/Bm1KA0GmxihKtfnjiQqO2yDNijY91VoHcpn//uzfPBSzeh
IxJWEth3sniETrKIhDhXy3ILKn6xSkF6FMQVHjyI+6Lrv0Ey3PNsdVaWiF4m3PFI
Ct3BTZHh5tIMvQQgDSPXhmDRhxfielehhhWDhfQyY1RchS54l5SqpPOtIYIue6x6
ewjqQZKrmnajwxfJZYH1YnGVoVkUIeWPmXeKmH5LTWzYavgfLQcSZMkpgVTeUYj0
A+/14PA/UZIYioHe7wbvh6pUDIy/b3e4FlBmjxBMorJ0oj+T1IQG9o7CMbxLE3xm
nVpBizVwNB3FIXJD8UhIPDOVSNU5tUMp4WBwTBe/56DqnAxxIYq0IZPywaeDIpRA
p1pPrRPu+mQN5fZnU2jN+Ge3SJWeU508dYVgNJYYd8gSxVuc6gytcmfygpyu4esz
oCiavA/44fLiftEpYjOov/8wcIDzTpt8JIjw32jmCYol4TyG5mF0bSKsBIXVKq+P
zhU6gR1FD/ozv4VnUIb30K7B6D2akdHNPbxBP0Pp9RCNOPyA1nuhE0t83bZbXgng
RYyndg9slgbF8dDxGvZQbNdR0LGnfz3fAomk+g9tRejIblczdbO68d4nkMIMWnK/
kJzlnRvWSTvgSY495LuVgNZlhbQnDKzPMg1NemdraSD99QB2Smh5F/t2f9CITgYD
TrEUptyQMEoHNDNNvaHDVQFLbysRZx82qhK6VO26HP7Me4W207TORmUMoLNmPVVz
knjA+lLWrhMRTdnZ69ljFUKs4mq6lCMzZMa6QWXutBtWaK4d/jsGzC4HLMP8Vg9S
kGhXGagMf55J8vxrq0ZMkBXe4CXxQHNaMPk805OfwddpnIK8WpD+iangSNyy/KkR
VPD0PjDbqOd22ZThHWQm2mJUNPxnEYarrSAMP4G6HXerJXs7b5dUdxDSOj2IyPrd
IV0T4LghfeKEeK54y+QlwSrt4DJXykJI2AoHwYTDIeahpC5lyf1iRDrv8Fvk0jx3
ezX5DFEX8QRrjq9OtjwT/yG0eALCBq84HBzrGzWTDCaxJQXjGrXBrqS7du/8OS+C
N1DPenwsHjSq4593pJGcXoZYwpQv2ibB2apBKhq4qqWKta3kVbRiJmZT2TGe80T2
+21Ds3PPbliMtzoLPPxyruVH/bK1D4DeOjM9tctRO9dparOkMr+s9X/wfbA9lBdm
8thdSOsX3C2FSkdZrV8d/Q01Vbw3JAx26sVSpqi7gIDsjjoACTSiXSD8xYgBb9cd
p8iiRJ11Ov6LaNwu6T7SgXti6R7AmthrUwqPqnvFtulNmrkTuGKcAY/CqRbTnlLN
GccUNFuUkrB/xrBFwl+qCZkjYjzQlr0Y/ndhWViEfsVwL3tQ0dwMo/pMtaKFtoaR
7gDt9ydEeYdlZbo+ER+QCHWUXBY5uX9gljsEe9k5Kwk4DXhGr/Dii/cX0z469jpf
9ka7EcztbTruJ70yVW1AEPQDlq+t1YBSNPF3B5RIpVXwvL/82iQKz3fc/UD9FXid
/vNeS6HpF2YghdErH36CCH4HxJyPLYTMcr0n5k2tOVfVoPbe+4Z3/5SQpl4eUbR6
gXTZAl3c8+P3rD2z/Q7Gfk0ssmQP+OTK6YPVw3iVVAwirvlsTYH7GvRJvQtUFGJ/
aB35Qa2aKxDpT6qZReMpQLaXpArfLZuhXmLa1aASBmnDQYaTZCCy7VC2EkEOr9Vu
WAq6oj4ZBT+CFQwpiftvwahdI5PFCkGEB8Boy7f9obKDx2tVXTaMsFcH+jvIIYbl
nGDmhESO4Kj3mhDS6H7m6oxiGlYpxmgo0kn0D8rjOwJLIcdAgv3y+nVeYYUxmN2+
t2X5d4AxLy/Lz50i5O6udIlYuV1d4IEXLsJ+rtuuA/DYsxeSFN0VhX4QA13usb6r
jORRilxrXgyU1gHzmANniBN99sYwIXQihhTVP3prQgBL5jip5KruP4HqXLRM9/fJ
rWFqlVc3O2kJZAZi7Oc6NiFJpMqP6cYW5kQFyoxHppzznDIkFJWEX2mSn9kUFdjv
4m07Bvkr/aJYFcu8PEcNxzBbyt6dJ/8NGPqh898cXqxFfC5VzhvgezzO+FesWUAx
lWSekqVdEOnkR52pDBKOuIJiN6nX9P85T0WQNJLctCFvTTjembCbbUildvMK9PB0
RdYtOu2JS3NhG2AuDnd20otAP/HoEk2VvV2KimRfbQKCoMtaE6EI4GHKb0KUXi5G
KnidbeRNc4b6kfT73lO3WAOOig/1y52tzA9O7HQvqTz1k8P918mAiuadW3lCK6D1
1Pl8ztA+r3oTx3amJLOma3F9ZBx33N7do1KwKxSD/0JUN1AYLDPKaSl7uppalZAc
hsYVb5mghyqo8IRPjMuq91WJMbLhCanZ1dlopLtcoUy/yBasYJFDZPRecogwZdMh
osEC9bZeTntCOgNHXwtA1+HBThmaakDPpwVMdjt3A9B9TiskhuWKiu7D0/+V6i8A
jBDM30ZD5KMUoq5gZIQGgtU6dz0uWBKSHC3pdrVM3Blvt06u2ZfrEsolfFf1u4nM
cFIf+TxbMXLAXrHnyw4wH6oW8R+k1ABJFnReOD5nHZARdezT5qrPt6U9pu0uCsss
qwameaCE3JiFDqi0iDAlg6co25iR/wHUrcsLbh3z0SrAY1cvUTKwOd1hAzJLCBZQ
Sde/pheZZhxCOaNkZNb8BuHd5tsPwMnGSNkQv3GL1j0VyxekjbBNP2j+F/K/pbK2
Xpia+dS3tEwDjPBy0LvlH1XcdvwJY3amX+tsXP1IHP1jKgmlpe77wPR2ciPNTsXf
WRNVc462DJ2FwoLv7rPczO6UJjz45XEhoy6sCRNrPLtTRPce1AxcoNurE5hVaLgd
bx27b3Rt+oXGU5GlmU0lYXZDSKUCWc/pAQIgbH/CH4cvDids0/VffTYQ2Xj6wO3R
nrXiaGmdbmpuGiPQBjHHNw7znByUGfv0Ypv0CItFzs+FhRwby78K8D54NDMq/CXp
j6zGeukMNC2oYuQIRB1WTfXKQrnaOxjroPZccxOC32FgbjbN9SPeA/zk9jTP77AD
V/c0LyTRp8bagHkFPHKBRGD3Bqx9aG9hj9u4UR64lQzaaPaCHV/0uj9u2oxgNUZ4
E3vZ1jT0ahKuiH4zZb/lUetgyUGeoWtdxHHotT/BTtZasImzm1bJPr/NSVHKER4g
4l7TpV8iWinLra9fFB1umkcfkiy60aS42oTRBfUHp5Al7jIcLNodfxIxfkzlWo04
xEISA8sz/yQ1rIdV8O8TzodsMSr7bRzwDrxQOPU8Xt02XIxKRFQolmaLnBV8fcvh
QSJTZCmpceUvqY9iJOTeIdSEUrInv9eC8X5/VEqORUqYwkR1iHrLrhWnUS3GwDUl
5RTZpe8Tj4o/iDSvDRPW71Wu/B3dW218E9mEnXVn7skitWs0ESoGhQ4DazHrQ4gT
8Oq+qSmIKkdDra4Z2WfjZb0wPlxVOj+7M4AboGrw0fcZZH/g9lRn1DaGW1PGNZC+
ic6n/oXWpATRjbtFKeyq35FQPmaXTw4ta+LkT+d34NCKL54FRNBfMQch7ZpV0n9n
ObdklLb6nvsTcuDuxrxPsWJhUbanUWVq4Nshb8/PMKX4snLm6g0fn0ZC/RAqU5x7
mQZySYdPszs9dgtmMXLMSIX70y4VCtwDDR3yFoeBOoEK9fLILwpnmnQSl/duc14t
OYTL0/mQlfkIzf59YJy+GdEUg5KFN6q+8dbTsS1gAMH2Vg9YBFYPsKSCUQopf0jm
z8k4Eh9gK2Mp+pjy6UNuP7UOPKuJq5f9wX6UYVKeAMBWtR6zIH36LuP0ntK5yCIJ
+E1impQ0mKteiRq+jNgtcZGZhirftamT3pM5X9WsAmqV3dBPH0spWFQsjwArgOJj
8ZZMx5AU5lBwv2hb+LG/IHlBICQth3NvVd+HHU+XUQ58yUx9Lwfb/BfLMBwOhIq7
ABRrrJMO06I7UiMl/XJd3CEXRbarnUISnIHS5ebebxD4/cMSFAXJv9XJtRHF9NU3
FdCQYzBWju2hw8RL67EFyis1hUYxb4i7JGpcezyQYnf2Zn8RhpbypAOLMKZPXxf7
4Oc2d+HcBsn+clPkA1bZOQEHnN/IPfYua2jjr0Dr7yLiq3Q1pod/0mVKo2TbdNWs
s+bqtX3xfP+y+RkTGxE0NyXxhA3kWohy8frw9x931ieC8bFEsUtpYdu5eLTdJlMd
AjyvnAMiEHqYwfMOIZ8bMdeX7Srt0obtHbmrS5esZk8JSDcIFExXZq0W1kSZmJor
ssKh60N2sMZZwh9c+eRhVcaHwyu2mqbGxlbI03Q+9MJR86cvJJgeMoL09FVbCvz9
6SPEEDJoaL6kmTKzDjw46+RouMfw07gEFpFWkOS4eJB7q+EVtXVXD9QgQZRct5e9
QLZBP+rfXyB5OVVRe+lz/+9vtoJPX6oE20Im8f2b/QoqRm/Uyft4bbsmaZsdEbLE
AJHYIAdLrcIO7gd2K4DHdvK8Kx80YUIQDSx4wx32/46rwso1mcVwM2mh+23Xun6D
0V35BnQcTQiSILLwUAPqX6A4OSYOiwVUKHQbqHccy1VLvAo8WRdllGwRsmYmp1p3
pvldSc34nkQv8hm+O0w67X3qrC8h2w429s2cs+vUu8vrf1mXpavjEzJKrMAQoxkL
YsMOXTsJ1nVWp7Io2P3UjSAFO/a2OgjC1NEM9MI2SwPYg/EiYdJCNAj1YTeW+Tqq
1fRCVpzftPEQIyDtn7aoHFfFXKBNK84mByTGWA/ADGtXUaPAC6bVc4ML20Gj2YLZ
0/+2HyqTSgudwEVXdStTD/dPtfhOWna4gs7EXr6mh8joqPKLCKGzDqmqRRoKWauM
cx2UwWau22YZ+TrhyK7IU1el5sN6Kea90CyrBHtJ7cm8E2S7TsiV0saxSMgo2p+B
Gl0vV0A4Wa0t/Fyhv3pluiRpv2Ns9Aics9aDn/QJWezSLFaKf6+r4cZ8uoFDEvpW
emhXfe/+TFXTqAaKPpLWq9qCt63VD448ABlNkP/MOln+/vPUREtG5fjLTNvBRgc1
bc7JPvM4/iIbukpgWxd9SWqMcibGcSogiIINcJyr5bh99SvC2yF0flPqykplShxw
wpm0oWKeqtHWGEMe+2CBt3SxAojNoJCjO/N6jNn1VzOzLqvt19C0LaGZeYzu2ZZp
4tLC8qBmcWgPqR+P6DzdpL96sD/T5zgS190HCNBfLsWzVu9oErCPqWj+NxgJpAIQ
g9IKy07jqlbi1MMBoeJL2iiZbbdOjzQWYJzxLSlz8eoCc/+phY5JIEis5jvOjSvT
w5mPUUslbTKX0BCQLiSdVevWItRUTsiPyS//bFg+l+vrrT2qf+OzDQplLg4oUPCp
k2wPQKqTBGLame1v3ZkSUfG0ZjEljxhS3n0JEqKdj9YKe9Lq/CFAkEfGtp3qM06l
K0H+QwY+jqmjyB4XJKlVG+UuUBgqzWIOq0jiJWTZ5cmiTwbVtP9pQfMpejzztsH8
OEzVTSR8abJYGpq5qSxkxPl7ssPFCk/WnOWm4bolXPv5yWJvtVbpmC67ex8hCWfz
DTsp1zvJ7/HMpeQ7KkSxfx2VrcX3XxPpdmALjdY9wnSCSkZMNH4lGEQrIS0RE0u6
iA9lm7RB7EGrDsatTTK+H/L0Qc+EkI03SfbtyC3lSbvSejebFfdz+Kop26/vTi7M
GO7hwV7co4LgZ2/XW/ZK4dXfAehSNnUw+bZp5j/KAuStS201zFEsoIVViFlwu74d
xs5dyDM5tIdhkco7SvxVJtI3EdYh0+asd8VPH3ZC5/8C4QmRJKttYHbKRZj8+e5b
gW59x2swwt04jBomtonR2YphFFt8hZtUmn3y3DcTED6qqig4XuF04qwHRZt91m4x
hfCEe+3lzTW0KdnI7mXD8PfdKDP+KEMpVdaJdgAsW5y/6KphlHPZBlFgYmDoVFfV
IDulbO8Dv+w1+hvXRJ9XyXh9PT37HuQ2XD48ZbyCgUP63cdSR/xRgoKKhMndPqxL
Rpzs+xIjRZUzVnV3VK/pXwdSH4BvjJsAbkeqsvfZixTNlJZF3EVteN38mJtl4dKO
NlXuS4WlZWS9XaerQQks1rmOp3HZmxhyH3x9+f9T2RqoudUKxxQ9fB5Qhdlj/Fh3
iZj+I8KpVBFZuey9Qh+P7tNVRrOtXsnoV3K1iGEed0dVfydvJ/aK05D8VjzZu3p+
Q+J+yz6vbkQywxnnytQxby5ViKdnNJUNxjhzpEbR9n46M3cqu3YocldOzcLXpCpj
B3k3GZItWnqUdZkUkq7ev8dyQOSHXqKDNGRx0I5dN4yI9DBoxP9KVixLjtzQ0yMG
MGR1gL6ZET6a5jhevZSi+QGRq58jQbwlEfc39C32Lxf5OXwz0cIMrx4sbct6P2aA
BIiAoYglL87FvGlWn5rTga83JOj5/l6bVLRfeDI+x1+4pX6wEh+rHeGrmWwBoVar
JdK0CDLrZTpSgmQBlVkQPJl8+UniDOKFksrB/XtvYI1abI4cF3pQjtp6FsVfScXh
Ip+tvhmX9GkCaHmZz9TuKrd0XoiuIu306XfT+hoX1TmhKU4mKmGtXstsSw7kRr/u
Hma4fevXAFnBt27TT+PGYqF+sIh4tq5gYZPBRdcnyO+Fvn1Wd0FVDoB9vtjOevfs
mKGjcKZodSudbNkgkCFURfcc0iTgiZ0//ta5FhqikgSyXu7njM9nh4Va31nwPnOV
fVF0hTXyQsfGD1ppa1Vvvd7VjpIav/sOEvusEQ0/bbVSi8hVpnCNASC6wznj+JPs
mfpWu2Pj816xjtFv94Lr6qyhhE1F9HDTX4aJooyJEi943dvfz/dPIdWAzdIWczoR
lAq6MM1rEt5e5rLn5CQlZK+yxP7WDZaD1DOBp8JntS1LwwMCmwEqwKN/ZG34rtP7
K9xp4QVAf/4JOQ2DnX+d2EvS+ZSJYrHNxyIx5mlGQE511lufPdLEr9ezEZi07GG4
7tm73cl0vcxiSsu6hgH+c1A+dYsVEhq5DltzSTlTx5NjUQyjWPwtLsOLQDQIX01y
oGb6Pdwpy9VQwd+B7lK5l4wdlZbTaz7sZJNgdovjN6Q3Bjblf+CYOSb5ueJa/ADz
XuvZMc0/ZUwx/8lCx6m+7+J/3gFJvLOLrRYhuT9hvKwZZiX7V0LsHBffoxYZYIK8
tqv9To30SedFHFHPvUOJWHrkNfiAM/lOud5S26jGA+NiPpD3znaGJCbASurp0Bu1
76RC4SwxMT6GPn+qf8SOCoMCOEXs+GPrl4+4ePTx5ZlgwNXjLAsX1HrjovJ+3vSY
7UIq2nZKJWrW9h+ZtUIowI6Zg3EBa4qixSmyd1lc90UT3/xJ2ZcTnPHdcbdGsVJM
+uhiWwQEHcbJOCnUCgwbiUR4jewCrSGHsDuI74PUZD/Rd7PuZDdTuamw9ASWgG3N
DGTt25961USUXj/ur3Oy7A49RNoapVq7Xp7IhH4fITW6R4J/lr5pm/9nvgB59XmS
0WciwiWpjVTD1YH537SN6ABK7yz4D5GUwKHZqDz1LnJ4JMWLUQ6Tpf2VPt2ltJxO
xs7Mg9YO2ZyfvSqwLV9zCBVeh1dusBW4axSkmVhrKKDcNadUzEq+gK/795i9wj83
Y5ioJuSJnbQNHP5j4L4WPdrjJrMWLcM63fq7T8Y34W/lSqSQVSIQazNTp2b5I1Ef
Fc221lJIlfgiWx4/jnljIsir5kgu07W2yvtzpVz5FZPZlUwgrSSrPtNjvPVbhH7l
jtWlS4JCmHJxvyv54hlLuJxHxq8fOAAYTyCAmhy1imF0xIu78Xz0SUFRmdGnRy94
inG22GKG7Is1iLYMeB28bvJ75d5AyvTroYkNXZRn1re7ESQ7d9Cie0+3oovxD41R
IUsJcvwYDe+nOjjTwJpuyKziK/w9loCm9GPZqaZ7+uZmpQSiFx2Vpdc9co67FIgi
RAkTEXnPepPZ+y+xOw84F9GSBlYC9q3J7KnL4HMbnfNea2PZdwWmrGZHOsW0TMIe
duwMFZRIYuJwjOHh8tc2RB4HPlqDSyIe9WOsQGSuuodVvUyBFjaf9h21eVRmq/Zb
jyMXAjuWw7ZAGm5ukCz23mIledWMlX1EPuuCTm9qm4cA7e0ZPW6DArP27TetOqA7
OH1UwXY3O9KeOHRfktKPPrL4XMi0RqJL6RWu8p/801diYc2J5EncSMHSXpKKCF77
+qopJMwJAeKvWGR38eddQVzQDTCPvVFUoc6LlIVds0Mt87cUJRduH0XVUqaQAqcg
szjCWLdzbgz5M6fadR007q7pu8Wf4O1wul4vwsB6TJx/VOwzRtLzyk7NP9zQozBB
mI+OwJ67bRz78auJm3zSaXnHRJ9K6ivyVr4EPSnIENNxwqFJ2099ypRZ/hoj4SZ5
60OlGZw0YvEtuQRM6Xd/+Vkk7pJ0oZZUBrrG2/8k9CfSw1rmjX1NVHlCyhUaHtN/
9InKTTpkPFMNydM9aZuuCaki/R4JSF+aj7Zv2wc+qYSIiifXSyAd2t//kxEd9yEg
i3/Ngk3fo/Pi05B5ZVYofIhB+lTp9a3ATHAkynkYAu36vV5cmY+5xfXJceVd1W0Z
rnDfE2PJbiehYJGZ9hSPh68wdO4Y5E1mAOhbdsdP2v3eLeKSYWo25ZHk3sFvfgOo
AHSPf9aInAPpJdjZVsVmAcz2VQ89oY/yp9vOXo9zFTN1cf14ZdYmpiReTLivJgxW
4YAz4gGwwLPMXkgRswBe4hE7infgbcDfb0x4y1EQEvBAcfVKMX0YaZDcWN9SE2M4
Kah9dM26YDLFW9c+szJ5Uph8PGIta8DmoQOxIWvuZv5kB4bGmQ7yMF+myxRcbKOA
24Js3zseZpf2AMOr90nkAy+jD2LE6H8RkDVP24U1FQkcs2Hg66HsmulgjmbalzbR
/3RcSZqM3mkrALuJEVcgbmz9050JGRenCt57WaHKH4nRkN+MuU3xI55raPcyRDUD
+3BFrgFeI9zs/MKyhl8GNNElr+K+nUgeAB8WE3LBSVI/wxvuI3EwCgQFgTJ0PQWs
KjJH8WiknRnnbZz+CwG2n3rQ3WLRekmqi4qY5zkfloYfNaUBix0mlmSA2fqMT3uu
vWhwPDeC1rmsuT0Rut2OAxyB48G1CJCRKqnJbszufs+fqyfECsvRbubgpxTBTy/J
qyhSs1T4NN5tMTmUAoqMO62YG9o5XYuQKvRWnYmL2ENNLLYRcvF+5UDJ6lcHfc4z
eAaiQq+M9Lqrn2Np40y65RIFbT5oCMe+4ONVbIYhBYn4KrJkSh+MhTOopJrNfUmo
G4pOW/MBm9fYl+4rwW6ooE/8R9+9Rowcllbpo0hKVxhPh5TG8iOUoezWnVO4SI/Y
r5u6AcPx1YeQEpG9JRaXSGatYGmRndSE3pZCNPjQsMG0ffW5cC/TEQyDdfAlYk5l
iUK54iOmtJhB129LH0H02bkPRWmz4kEUYZsCaiKKDOW+Cuk9u5SsfsEKCfvs7OEP
Zm90EqF2vkNqETk+UNN0sVTqbX8KUZgprScriu34NlwjCtOcw3fe1aNJ3Rc1ZSPe
+EtcpSUdjL/B4YVTUTJxUUwwvlzl5SENd/t/o86u4PKulm9+mgNPdoF7x301il8m
+FLnz6greAIbQPJh5bxXekQi2iyhvnaWFnjjan62lZBlyUcBEUenMaGhmbqkWfmC
XQO8bGlsSVbMyxzXgikrr55vsWc/m9SuIApt6PQS44j96qW5UdSnYp7ZnKz0F65x
+x5fCwjArncswif2f03TSjImYV+y/tK/+PCxWwQftitMVhCMuKI83/OP6Xk9qSg/
/Rx+HqK9AMcYzDAdQhto1rHAZsjXtKbsk18mmROanZT0Pbu7QgcPZ7uTwOzWFhmF
zcO6cUgREqfh7YFvu9/fm0J8EjBaTEwoPJpONnCc5pM4juqw4vCB5sys0CwraY0U
AZ4ePhqKvvYGiwcO0XWck7kUKGrfotD4PK3nzi5NjjSBziIVXT/1ZtAv4wzWzrGf
zd6sNSP6QoLQVmYcNVEUXx8pGFSBlN0nQKXI3XYN+/BA/ZtWenBM+Y2GZ2J5gb+/
iO6RaD3yHRUBLXtgMbidlLRnQCkhsaOdhF4xIkYrcujsGiENWgyqg9n/AzfxC/x2
pjrALMaHPn7bWePQz2YtW0MkhrDg1WGIjzhCCL5hfwp/a4wJWdRekVW+ZBV/THs2
B7s/OW4pnEg7RzQjBABl6/C3zX8/3TwavPRLInSNDmYpe7FlG4OfVoWb/Jieh/fi
3c/8s4zfBWAYblLt5o4ATOX80JU/j0dNmf/KSfdSN507GGhrsK44hbClMVpvoMY0
aDuUnQPyh2Na2KtegU61X/Bb3aQheoTuXnwsayx3+zkzQqOi35CgOVEOeiCzm+Ca
gqc763I8F5ozR5p7LS8/4zp+QY4A39k4F8HOYbMRLzgXfkK4nMdbokppm2wlLaX0
D0jIQr4PyS4BUD3FbZYT8e2NynDbjX8KckVgmEXAazh8BfEnvoiOpUPMQAxu0GDw
Nl3vizyyX/VqgGP/Rv4NzD4f4DrNafSOmdusTYPhnHBmLcSmPqnfaVhZFDfj6c2F
yvmCaEok6LjxIaasNcA1WVFVpRlVxqvy8PSbdV55Cfo0DmJBLWnTMfIp/X1C/e7n
D+5vadbFiKL6+fujd3f+wFoQHUyjfkcIEAhcsjT0mziVZfNHgEOML+OBAzPA7fpx
vsJ8cJLrqqra5MyuRGOaXc6AiPKo2GOZlHR7NbXQFAkFgagtTfNkDeCTC9mJqCtL
o8eMoDVtj5RzrPzTVD+mYFxDul7tQLauOX9YndLqoNpNMuwFTRWQcAJq5qUbYOsJ
y5sWL24IsVk5hQIJeIaVMzsUKcqe3litSJAS8SmcA2udbpKwRdxmiyEPlZr4PNEe
33BpvRNfzxtIn3rG/f8Gc0P0qHtzE2YQ+A4SnserOXz2UuuRHZC3XTjLu+9uou7f
LtJu84xzhhKO+A8rlYUX2aTN2B+OBBUIJfigJ3vZl13tIyaryuLC4+J2cKsMUi2M
YsvHBDxqvGDjEfC9hYcMRZ3AMEP8EeLR+ZoYoBb2bGFZeIWbo1XpAwCtY9TbZzXp
3mI6cZiNKw8oooXt73MvwKSkMN+Xkd1gPLRsjtkuw5WuzTRqIRbXtoX207D7zsv4
4Q9sqb9c1LW95lcYCf8nO64AbomeGuReoON9pXaUpGu3SBp4k46zBLnNeYByiWVh
LJKPbWvLtqOp2wlADfpQFQ6gg8KL3Oyc38J8zf/xWUmW5/X/u9Fcp9bU6GLH4x3Y
RdAtZTvpnvoeAK8EVVMiGt/PxB4aVBCOnYuKAHRNU1UWpgSc99Q6lq89g8uktP7Q
LU6E0i70XZ7GGCLMJ59KQLXue6eCUlWE9KXwPRwQ1BrQBecSyxHi14AndH1EKSAn
pnktx93T7bJ9p01EbrNB3EORHujXSM4mvF6BGIIRpyY78caQIGYOjXINCJtx0wOP
Ubtf9iUyh+FlsGCA61f6aciEFesm9jGJMnK57MvZPTEflE7WWduB+ueNa+RgIwtQ
3T2ZS6FHdAJk2tj7uuKO0mXHwYmBtqPzBrRIjrRLxuoCE6HfAWBG0Dmj4bpXauUl
R8Ks0YH4gNLw5RR0PUwmWBOWz+X6fC4H18RR4OTUOqSVYo+LOhd5acHpasq/CQjf
UAbNRyIzjeBYW2N4hlgUbDaD4IKKXv3mPLIGXT1lRgy9v4gy1bxGY4VCBF+F2qKT
9WMk0YLBRUyFudlz/6Flt2WaRwdetfgqKkI4L3uB0uYkeylPGcUxBgk3xiBGZtbo
9ChA3FBNE7mTo/RTtOjnCMqVsM8LBRVEyLoFK5mKXms/38yJbOvqVlLs/aXILU6K
stTCXXxVKZrU6NJ4bUEtlAQRRXLU1p6DR1kgT+MBbB3WS/rWp5x0I16DikOG9rrl
v40Jy8HdreXaV585u7tUeRpZJWoam3LrdBAgqIF4Kpgm1Ykklo5gyg9+XTlOUVL+
FDZvNwzZSyTIkYdwPQCSrIusC0+YGDg+E3iAD/ioRzesorMKx44iauOv1xXGclqC
oQPmg6ESf1QvRi0LLBrygyaqEyCooP2y+DBDwHcpf+XoF2xr3rmi1ewtd+DUQe2R
ddsPGFTI8eWzW5/v38YtXG76Tr9JRSYXSk7maSAjsUin8lcj2fAlItbUFR9KLSHb
oyIwVsoatPLVu0VMDsdHxNLJS1P5kdIolwoQBRyaVjxV2J76PeV+XBxa6U1eIKax
rvq711eiuXEDA8wCI6PYJ6RvRbchyRLDQrRrgTDuAUklJl9YQq8dnbPBQQGbs40m
MXo0qTSI5cDWmqn4PJSRUd+HlfqjEGD05D2S0MAtSymEqsu2Kre2UqAKOqIDTyCh
1AgSk4WkpFiDirFSpYGFyB4qG52ndpiF4SbaOKph/4zRKK3xDDMpxU59aVZXMRB4
f/IBzrNLUPtXzxBnoDJux2CMG+ex+45Oz21j45hl49OQMAqECjH3m64w7wjyhJ7l
AMp+FdH76FXihgFpbTaZmr3opBAQrDd1vwKIZkQgY6Du6Ht/VD91xOZ0H+P3iHX7
0skOhm8fatRY24w+f7KWdOc5K6ekGVI7t2uI6J3DwbJIBxP3iggybB5HyuDhkd5H
Sy0QPK+XfGWnVWEQx6CGc+pKzYGKMjidhin6tqK1lgV+NizTQYqYv17HX5OsiDvC
ZB4DIRd0CIyVRKZ+rDfthCa8f2qNjUbjw4HC1Bk9xDNWwZGX71H90Y3AsxYWXlkF
P97q8EGJloew8YpJmU0cDI9yieH9+wG8qB2xqfI9S+6rIFlh1tM+T6Nhppr9hIew
i/6vJsLjrACa+aiAU97qegRBSW9GyQTs9AphVM/5m2sO0LrZECTPuG9ruQ2l/rCg
OiUWnoklNsk8aiOlO+ZM9saGaxb0P7X5cyopB2B+8luiK7iHSCIwzmR1EMyiiQNN
NS6M5wgX66xY4bkEJQ9l/Ja80haxkWfnFs3T7AlMCHPpycWitACGgThmbCTm9GVA
w3Z8zvywATQkfm97ttfm7Zy9Jsw2onUOLTu/cUsM59vjvNj3Sai4tXFgtY5VkyKE
dHz0RmYJ2HiuMCuh0n0MhYsHcw7hVcr5g181cBQPSxLXG8KbKZgzXEe26BHz3Ymv
P60ExR8hm3p2VPpQViVSZ17dfet8wB1P4zmbhLfdnTUWOahmUOqp0GBt4HOpImMW
R303IFQ06D/8lNUEwGqauoLWaGQh5/vTU6CoRSqrsiARGPZEtZw+totek8TW1thJ
49kGgLZMkpYOYkLqX01M9romnlvPqeI6ypuW+2Yw0gkHGxs9nvy6spTkg3aNEzLs
qAz/PfqksWk4fF7JHhEXNT5ZhTl4AhBIj3/goxYJbbwRsgr0qd5ecGRhNwvgsCws
vir+V6wJkbOkSDcLM7yTeMKgyaaCxr1wt2D7GduqjJaMTmyVGa3rgP9J2L8XMcZ1
p2wUilnDAjBqt3ckGFsDJ2Tlh2Sv99zIbWzToBwv0Yq5xifpL31gZikhDNFQOjHB
5JQ6ThsqAeSAbHUN4TOeAlSiebnbdIOuBHxWEyQ3wgNNMEcU5ZFwCTS4msuXyhx+
dLhCIEZkZuCgyGqq/fue0Om4hsKACSI6pf7rqWR1D0C1xZ/PuekX/NXv9/GKQllF
vM5BiUE7AYOiNiuyYFh9QpfHCO2A1DfWVP2V8/wW/gazODHabQjF2sPY2qmKBcMj
eDABudiiEWzijpHbVk3/J1LkcbP3TkLHZFt5nDwLaqsfBNltzevJhFtnYPPZB1v/
pY7lZdLAiF/pvoQNY9SYVX0wCgG0Kmqgi84NdA9rg5T2Utj2cNhPybcLRw3nY7X5
G5BM2rMrfyh5wXpcj6M0vMNw4wN8VRaXXb0EMjzXsW3rNG7M+Wyn5vr4MYsbPr9F
84sgHPbS83y4Q3JHMlR/GFRr3tIgu+QRgCjJLxkCBlNxKh1kIpzLs1B/nCeGaUkI
fEF0NVdrOX9He+LSDbQmCesucEaaKxeeKETeaC/qM2AxCZLNdtkXeE7sFTdpb1/C
3QWObiW8miEf/koYihe4a5Sw2OASvm0ORu6uoYdZaqMYEcwKPnoGOJbrKri7omdt
O8Tarh+JhSg7aziefW3QX2creKDqsdKGdN7HeZS7pypgTixMX/P/AU0mx00GUCmi
SdYVWmA02gafLK1B5wpgLBOAyA8UgORLCUViwDrZo61OIeI841xMFwDOZsn9/5On
U4eKBCCtC02azYw6SABE6zFBSbQwEjOfblRLc5XYcj3i+VZu/laOU/tZMw7Dst0H
XNSqmBN+920N5ekAITPkKjO5RaC4uTeraSZY6sIDNLWVQBmbko9XTBqWKxON8k0j
DW5sWMnSaAt7kKRP7DShfRFqiFYJC3x+ZWFxuYZRy3dc/nWteQwqUufYGM+AtwOL
ijCiH4CuGgehhaKggzEXbnru5smWvBY4S27zPXz23SVHAnKpqgKmpHxBGD7myv1d
n2j0X85L2bWhX+xoEhUBqYgos25ziHoy48/Op1YtRedDI80FYRfflpOeJpNuRx88
4SfYS3AiL9ArlskGkCX6wQSQALa6zYGIf4d00hkONNvXwZNxfLC4sZRxzIud3TS+
YhyxvOELIv3KdU/UGWSBaoFnLw/QGad8hh5yEFHadZzcSwb37WGIp+57j+X1wLO5
xjwFjb4fiQRtYUjv3VUDYTcQZboANrHmqJkBA7Aimm6i1Up9XPBU3oh7LluJoYRP
Rpi3NoGEtgEKzY6jhAV9LQT6joGC7oEHpuoFngTNqGdYOtoZEJDGL2j5ytSQM4ym
9weo8KPr1asjo0tF6M2xv4kbLl76zuyQlXwr69w4g5sMwgdC+d96fuAVjbo6ewcu
uDzkAS1CN24w3DrEtB63bE4W0bO9TknU4z1/dIATtNY8T1br+Zkfl7GIrMKKfg1d
6qchTGzQqYyvpkX2H4ZgsNRyivJtl8k1JovxTpJGOl4Si36SuRcwELeFvQnHeyMN
xuM0l8Jh3KsGOAabTMMXemnNbSa45QrQRmB9xyP5r6jzOPKOGeVAk/uGvDRrZUpB
DwIMAvc54u83TS2AhlsDBb6mzIJjImYb8Qq7pAwBi2PpiI/pZH7kR2PNJPn161s2
AJDp70mDO1737vmmW+62os7qknP9h8b0iKJfwHo0r7pGykw8rBNHRXrFOqbilMJK
VLbT785MM6MG6Uk9kypJIly5ZarAyy3E2O9RPo6AA4kNgsz0ZVLQxRo+Pm4r1PHE
nT3mTWdO16ZVw3Va1Ok/qResYd2XPI14LKbiQelo8LneQZyvPsTAfDBcH1qlwOrl
Blo7fy7TiNudQ1QI+QNlUd1YfFFx29Yrnta+6dfPeALKAi4bALClOQJocNJ4iLQD
bNVsORxzcvbfj6ndDM9JaRmucn5AAHbfUHQ9JWyCzILNlhLx8XW8vn3ykL2fFQHS
DQPlAbWFp9uHRwgbBXQZIFW589g82I9xIwFpXhDoSvZgQKmHL+JVtn5UIgxNDTuT
ou90LBQkUuUctlSso8T+et8Jm/tcoe+gzd3JSKbQHr9a07z51MjUDq5JWiNzp2zk
9aMVK8gB4KpnVUP1bgc0p7KTon0xC4jEpM/MCHp/cUBn11W/rinbzD/rc65t6iLY
ao7Bu/7Asll1aFbeYiOvL9w9V8IgPVGFmKDQqH6fpvbf72J9J9PXTjYRmiMgzk6N
yWkJgTXTgW+K26JlpvbveVwd5mIOp6NrT/JmM/fcj5pe/guZBLmaQDV79P7TVzVw
QcOFJpYpe02fAAFPt9ZpY0KGRS6XVn+LWuraYtiOjm7bieq6oNOJc2l4PmJT3aui
s/VaV/okZDvt+4E/QimRvoAtPF3RqZFDsz9VYRD5NbAG0kTVj+rhyWBKBYiJxTbc
f6bH6LJthrVIjUeMEqNVLsGLu6UZGV9PZWgt2NXaGwSh80PtVBjAMBHi7T0bZiqy
/sDC9S+UVQC8k0AL3ERnGxDoimswbwpxjxU+zf/Ty/h2N3oyf+DDPKpwey0lrv0V
ToKEQRYAYjuI+C5QCzlm58h2XLUXGD4KEPYjVIHSKS8p8wzRKIte67HtA/0nuln0
NAsXnEr0iugxH+vIzgbhYoz2w8SL7BXp18H1Its7yIdvRAfJjEK/+bnfnrkspHZS
m6WfO74NW2DAinQMUakXl9F2bL6uJsifgDQg/KgvMMvkMqTOsJpw0DRDvrj6hITQ
cGLcv5rN1UgdxL5kY1plKcVGqJaoypkXU1smnBIJYhP/sHN1kDxNmKxKZvlP2V+o
WQWfL8nwxvWS4/GBMEk43qnib7S4ueTKV+k9ZoqnBIXR+U+hlFJy17nVPwqBtkRV
JzARMlex1/m0yw0VKS3BcF2EwikwUdC2B3Ar2X5p3oBzgsbAb3dmKNu6Hm7RmoRL
3LyK1VO8CH0dsS7pWNp3oI31m4f0W94M6WkjuercUw8q8xscBgccUtFHxM4FbQ7Q
A0G87mw5cXB+55jKmwjKZapQfjV7vqHVJLhNwJeJJ6vs9UZV0pxPa2oQEDBp/gvl
jz4s6vVgIN3mgTAbPr+uJwEuwGbuZ09JAvHv+P+MEzlae/6L1XFzk4YyJWPPzXXV
2tmUZFuJDjaczLmKB+vZ21t6y9tUVpeO1SK7QWQTFu5zudtZpU4Fnu4EJ5bO77Kf
8yXqHGk0sDP2xC/8fSd+AWgY7/XXARnexskjGmfGOMTDMQe9b7o6XWv621dQt1dO
KUBHYLxa4lPDNebgQrarZdRr271F8gs+SZK2pEXbCZngZ7FQjCtVPenX5I+TRTMa
XeLdg7cXzBmAs9UCK/VY+x2JqG/sPIAliF1SqwQsKkzRcosdulnEUo0k0ymODyk2
aeyhX41VAGUGSh4XZ2i41kR8poszPIQK5XatmqI0NAlcPlhr7VXLS2Mp9Ms3rnVX
OlhEwRB19xKNJid1qxQcxIzKOeKT1Vs9OB4bI63RccanO9mXw8Lo0gRB8FJJqoPh
DCHzKa9os41VljrQYs418Pbc/eyJPh61i8+IkjMg68FGzkWqH8YjM6KFscaIT/K/
Jrn+rly8tCXvQ1HZggqItZ1i5Ktsk8g/hPEKoRfmX1yQ7ALrt/N+0yKmp042odAh
0bFGPbB48A6A2lkKeic9nikVAAfpitCGDsJfJU+YEBtT7gxAHLGLDKHC9QAMXvGY
geuoEpAEgxowJxu/ajRCFGpXAHCJNdfTuy7OBkLXTS41tyNVFXMYJEL25+v0OshS
yWirLqhPfAxFQAqKhcXAU2pFLGrNfd7cFaMGx6GrIlcV4BIpdRlxp8nogSy8tHhZ
JMcCRDK2zG8wTQOvM5MeF9WQDhvM5r59sW+kG480f8oBK3iaiYZ1rYe19IRRwS+N
nuqWOvlO25x1ylNdUVSfJPS+VnElVCtAQGbeQg2xW/QjJGabiL+y/0yMlRzst0h4
VgZlJxXKzsFchkUGpfH4MV5uTVpxkqTjiPK/lNUps4PxcqAMeWIruxsku9Cyoc5E
z3rsNvrEqBmjdt9QNSl02YDUHU3G54Hft8biMqZEoPAL4k07Jjw92phgMXg+sRZP
PRvce7LBh8njbGNiIvZsoxNV9U2U40pDQxDr7MMpdRSF0SY2PRDAWz0PG5S9GOm7
7LSPSMEhpF/3bEpeCTqeXW1BcoyK/uNPsaq+LqcUe7HPEggJykC8zs85ewLBo1Wq
iuG112as6PAtoB+SbvGSj2a0snGgMoHeDg5s0LFHwACyGt9VHRFyG1VPJivT3YzD
K6QWCM41c1npHWOxkDYdbU+7G9XQr+Op/4/ELnTLFs414MZfkX6wN0+Su6yLpbQ+
ETDDfr98LXWGVG8OBQRkjmGY8ALOmJi2qqGqsbS+RaBvLQ0KSWIYMyHIfXWL8nfZ
4CBfcYVmERsSRJAYanXKQzcy64dYFLAoVgzJsgZpTYga68QLf7iDIFMXDKLbTst2
r4MhRAtwbrxFAE6PmJ1npjSanbQEIjCHfz4jGywQVgdubHfplqlgoMqoLsZZaYOd
o/M24w2sGvJPEoSYsWl0Awi4aVqSJKE9uP+OWxw9OBBrPcYbu2dTkQTEV1bP46ga
geaLfcfsUL7LrphDS9Y4Gd8pB2epxJzCNeTcDu7Sx7W3LckDsgN4CWHarwFJV5Tq
dAJ4romdMJ28N0X3axrslfu8VYTsjc8gYB+a31c661pZ+/1iadUhLTJkRtU+e6VC
l/5Fb8FvGF9eI4F7kuzGT6BCbNz+HIifw1+uwhT7ZvnlH7E3S+7xJGKnlG46KRlA
TN3Pr8Ss6KR7RNsiRksigSixycRw/z+gHrpFweT/EOWoEBuqdGa8fL9to6fJzH9v
OMSa/k/zd2Gabyn0xxd37zieDqv7nN1u15XTlnQ63I6SjzORNuGEEJtPL71CS3mY
d271aw3xnFziwi97YFq9p/v2NqbhzhE52fsAoPVoJcMW56BSudLyWFLisN/GtSKZ
6g9DphABLvA8FEJDvgJXdwj+I64e58tbWU/cQr0iuF8VMdFxIcH/D8yk7JukwQ+M
lxJTe2/HH/DEiVCk3um1pre+XfcfDuO6brU0q108TDvTGWF8kCnSGyyALlFQZkLs
fcJ+rFlYegH2cFUiOtwF5YkIcJVmkdWOMOfgLNbMy/VjkjPTri/qEwB5DNvXrCMb
ZrbAzmYnXTLVj5Rwqj2c3lx8kkztx0ig3NJM6V4ftjAuxjdAPiX1216UOqhua17y
RITNNnbq4Su3DINLf/TFHpZfvvlP5CiQEQdnxl1WGkPcHx4HxJwrBLFDVAK3GcA7
/8DHxK08drFwtfqvYLGQelqs2yh1L9OCH+hmeiaU5ePH2+SnWtHfrY5Odhmmxlec
ghjVQHM86nnhUOv4qigxDJ50l52ERlDDNmaohPGmRZSJKFEAnf4HIzGs6r9vrg2B
qM8MwKi/jk9FZDRwu1uDYfwCEBufwFE8F3+9Q65+g/gbauUGJ8AZ1QIf26Cnx3rM
AGUOKj8LRAQwrGI/lB5dK1eVd2FIIAxB65D9n+VTTmrnCP2XOuFBefAiTsf2hEyP
ruqaUkFNIcHI2Am2Q/5Gffcqhyv8AG23KGNMAxcXNyCGFzUfAXnhLwp3lMpxnJ/J
pPiQnfI/59sAx9aK4M18OxmOTTSIm+RvwHxBUCEX65K1+wEZObRrE6Kb+4ENa5Ie
Q9g62HD+0Y9SGSTF1QoKpknYPg2QYDTU2nhVvcvrCGTKFOYBflJnGrepmu61rdHP
khUego/yMCnDKqZElTYIl/It0h/wPr0D0ufMYBvfzKRGKmPt/B8VxvWsxUvwzSup
kCxyhWX1LxKdw0+7KwT3KLI6gvK7JLJ13NLXYfOKLK6U4Gpl9TGJevURRYaf55yf
F7hEpe8CtQ4LDQl2rg3o75Ov7/vCZ6sTkYIlrB3E69KwegRvxdwMTA0DOfljsT2n
NX6DvajWm5ckUHxnd83h9zhZLThmk2w8NDwXKRAUw9OcSDNB96JZKz5jU5X698b8
MPkpXYBv/u6XRwS0RLoVMrUUaYR/3Ok0XUlq5yMfqJNT2qL6a2QyVr4hAb7zFD1F
LTr//svS4yu4WzrLuQ5PITLenS/yA4TdBwFkLvbZvEt7M2bjqWftOeFPBSEoicO9
6zoQHIXpCSSWJV11QbQUaLLe8eLeAnxSBZF1q8cyuPnnVvqsXtG5ShOMgY/hdjt1
v7LrEBRfRS7X24EAGMw8Jmy7+AujP6tSWddDvdcClL7DT3MPeJXZxsYTBCeiIH0J
NxW8n2g+D9Eo0wJ+/9x1K5648ERt20t9iaJ8AZwelhCxTN7HAVOzDRgl7AoacqPa
EqkZ5crtvef3uru8iArSpUyDTs+wZSaITb46r2044oxNjTnLwW1oNeCDtMaB3t80
RrHysbfQsFNnnYQwxoGPVdEVpBkhj/Vm6BfneiwF3q1jwEKB+vUpucs1EXiVaQ2M
jTrIEkg9qL7WzB7IbqucGvnxQCiwn5QAJteAhG98GD20LAT0bnYL92nuTz15Eiht
E5FLzCB6qf58x9tPowGU5OuMpupL0Dgsei+AWyzLrE/XXSVOGSkOEvRPAYQdkmKj
AO+zJr88lH8PLOKh0JOuC4cAEq/lSvHowkwhbKSnqE/WIn67q7CO7QNDUTN6tTxQ
bIPaPP6YzLVypyaYYCZUuFs8nYEL5uF5UpSum17pX16COqeJzQFTp7tzolwSZGsq
EdW9Tyd0IrCRB82rDkFu6EcyGQligxKXg05fFk2I65K/7VrUPqjZl/fojC4pGMUc
tqrPILDeBZmEBYwwKpnXu9tMVHw4H0zL82uSoq01vj09KQj9dN9A8niy1D/KyKoB
2htTeOW4ICUzj6uMAa4M01UPMpkCdrD2zhNQjvgh24ubtwNJrFNy/6hJ2Fog/yHX
nkkbh0eWY//HO5VnzXRv/6dr1n5AulM+9hPgAt0YeEsxwsyVUpCzAWDTzfm1JO12
z07cu9TST9bIRGdzFPq53/X8nskJv3IZwomGilruEK9PtsE9jy8FZshta9nAv/KA
EvNkA/UWCWtv05lvO99arJHQ0+6RBzwDO5ZMeMdF26KT6ZwG68cOQ5jy5Y2ivQt/
Pf7m+p7bYmOKNQ4mg/ar9ea2BKE7gl7UHZ3bh7QEAG38Tn6dTwat1/Sh0Ne0HQfm
LilE7wuTmZa8WrjIf586bbMBxXVwJpRYulqPcbHc3/Uk3dz0k0odKQUFaw31ioJN
eNCdcg83UD4m9qYUem6C1bmaZyyO4cquh0ewLlLi1pJt3ugRpRFGRoCwryfeSsfs
TkiJEgV3C5UhZZ6kl/cuNeFaH+lQbvxJoaOw/pecEbdX65VeboKIN+RGgr2BFjAz
6X9cLfSTll5WPURnO/0zpBEvMHqFFmu49naH5ALhdU8UptTqbvXzxOYxZIi2wq1u
HpuYo1MY5KeZcc8mRnJjpGZ0mCNQWqMKHyUfIOaUBObOKi6Yww0erHFH9exei/0+
wDCkt+XepXsi0vF32N7w9BQcpYexA+MysTkE9KHKZ2JTEQHXAFbLM/JtUIRlZRzc
4rjCpn2k3UzCC8Abuw/8GKBAUmCCIMluMBAh2eG63FZ1lHsp4NoYmOKO+yGtVlFa
DAaOMKoSFEH7vB5wurTg2WxpfD8LjBtiZAwbYtZFMrxwimHDqeAi+B5vUWXHb1TU
XhVMa/VY0JFC0ycOxynj9A9w6v0zk4sU/d9V/rXL1DCLWtf3uAKFq3vFJvRxF4Nz
yLSPZ4fiMlY5VDi69olMpNXrLxwrocreVCy0BEUF6dwpSB4irSg9SNtXOk/m5f6l
yknKd4iZVpS48bjKLUaJHhUv3Me7LTRh1+ulwggQJjLuQgXSB52Y5XdPo6aOQhYr
fEpgFZLPyPzT9v7o8hwd/Gy7qCa7KXakW3TIn8i98myJc/tGM7RFn+UExpaTMTGG
jS9JhHOt83PUYRMqZrVIJjIbcL0Lm8i/n16XA9Y0ataH/oV68w/GWpW/cQUOJjW2
nKJ3z8jPJL0KiSuf3av8VxyFg7qymvPxOJZzoiPdO7sbgGh33vcjydYLRjhEA68z
ELMUk3IzDel/quQ1w4V2wTPPsKEc4k4cMJmoaxbmKFgXpLbYFu747yEgXLPsHix4
+wdJNjsbzZRyemBSt2phW07PzS1Cz1KNNq8FyJkMoTccz6WUkQGdFJ5YfX+3CDfp
tlkGNj7UNIja3eDy2c+PMSW3vx4fX4btHOCPyjmLsVLP+Ab5GRd+JJlVZbFXXVVX
au58fEom6YNAf+eTssvS1bO9DpC8fHEAuPfIPjwcmmsVj99G1z/QeGTc17qQGkib
tp3YPCJup1Y/3TZXa9lKlAnBH75G3o4r3x+iO3taaaaUrIZ8wlSRmY0cEnqrECHl
32BWkygBejBINi8t8EJEuv0Ssf/VUpH4kn/AI8GGgS5HFiPn89R04h24MOFzy/pZ
c67wvYeh4+3neDgvlIMnCwet5uLw/t6Ik2GleFddShrC2rcbIuArbqeegbFcPlFY
AauW7KQnRt71LR6Mzia1HselbaW+JhBpwwFZanRU9G1n52n+2xJHQnJO+gkHjLSr
w3R9/XXM/RP0BMczGwWCCbV/eDVA9HlmFMKn3y53zWX/fT2mGLgyN40ID7jykNPe
pre6BLWyPcMXvba4BOusYZiwhSmAyfwG6AMBL2rsj4noi6ImG2u2fp1Tn+WpXR68
RIMHvVRQ2u6HZG6omcmqX54JHxXSz5f8zw9gcJ6LwUUqWIN2lW3EK5it0C/8qYKB
TaT5pwrClcsc27ktVls4JEQ2rtDIdEAlBKu2ILCU8gGrq4L5HweltWP/xp1HtMDO
W59epc7J7LnF/KhZfvuaqUEuENmpYH5g6CmNPGe05oQ6WLZ/qvrmmUyh5hMcoboK
+68MzDATAogL3iDwQdv4PRmyxIQJ1G3YHiAwNtSsK0ekzs3pe7KanFBAxEaeXRQY
18h6F1ipl7C6DfI+9RCa8G7UJtXqcgLt0er/EUQ5evLoPTCT5CD91O5XRRr63riF
qGqqUiTSyob13xFNRiF+pQD6ZQjLLAlt/FnIdpXYOYsLzi5zl1QxYiREeAQR6dVg
HiEImCeJqPiRyeVVLxM1MiAwOG2XuJU/iLavr2KGti8IK8kSrlUAayvwMUPHaLJ9
4TEtfGiGTxHQ8hVpHBEV4A6t6YsrU/GNbXVBiY6CyjANFeze6UOV/4vvEcdESKat
UN9eZC93Uo9soh0M9d2FF4UaXrbWsIcXA+PGoGGALtU5yvEdcwG1YOqPQxDzwiRX
LXolFkh8fO5GDe1Flo3g6xUtOj1heNIT7xD0WTxXYuQxYCyFBTk+y9fl/JbmOkqI
2uVWn21kGa+pNjSxyDyGG6CNn7+RkfIABrhStqokK4GQ+08Lhwp7OVZrRDTn9rR1
CDwvQ9aw8kTgqZzNf+flKy3WEWDlEaFXeAPiYduu7tZOBqye5h1VjqkKFHuyZYtp
a7oC38h+EZz+8ld5bvKgQ3fdZCNd78McjE1bBeeBB/DyP2FXKAPV8adnmXEPCdqQ
RB2wPKsLhwRm7YMhd6qYH8MeniU7PTea5Pin0O0Xc8JsLvjmOhVzwhY/Hpd5AeVQ
65QJvDdyCTHPfGguO5rILsNWo+UZ4FuP5SXklPaMWTbrMiW51yMff5jqLnlT4T6m
12YgwRnxl+2OdPHraWVf6onVcCiYWXqCbC/0FwwtHkK03+N/W3ITciL+tigh0b61
VYdklVO4XTDbTuR13fvdw559YIu7MReBGINqVe5GLuSNzDUNVsnZIZnUpDAm52GT
uDb8ymKxql3Z4KktJfwAsDcLbkRtXFAbv2M6OOeIE+7Gz0Q4xXABipqEwdJEzqNY
LQuy1cB/5nkD47wzggvInUi6eh/qvwPr2rmDk8oapsJYvauy3fMmLkaW5P3n6VDq
qHXC43hgWaSnMggimPSCLkoITFub+1nG4WqkSV/7MAMvRJamEkVbIzXYAoAccKpm
ADGSi4Tpb4am9D1oogXm49xit1XZFt/pFJF/tkIrflSi13tOZFT740N3xKpTte0O
aKBDtU5NIKxLSe8yWCjRT+Q17LSbAy8OrYghDXC6Fk/FzOrMiTb6FcIyKBblopbh
OCf44RJEOACzIu0V0Pv0VdyJd5o+rSRWVhf476u3nDbMeZoG5kpDW1GJcS/GBNDD
TwlmE0Dlc7OJiQSdpGV7okMwAyloogOwg0mrcsykSQtf8ki+qSRB6b/UMaiPMWx9
fHktOMMOAiFxRSQHWB5DKyulzdphIX69JcXYW+4a9X4X0onI13nw+8f2Qkl50GlB
LOBnLwyak0eQ8aKHURvqzzejmfSZvv3DM+EBGAuRKhQ5vFD3CMSY7gir5owkvTK9
iPSXcS5kc7tjUlK9Ospu9aR5kbcOkJ0WDRC52CVwF01yWuOQFOiHp8urposoSpG7
aT72i0aTS/MkwhxKJDbDdsebUBE3Dok5kVCNaATd42yVqp4YJnf5z8R7+z7rb4I8
epZXZb66ktmIbrKouV50rr++suOpIRDMT+k0zdU+dxXz8PsDMQzjl8QOyynqEFFy
hxIIrzO4hag9pZJitN3GyN74svsHjwUq/IyvJKdH3TBlJ/G/TOambrwyL76VB6V9
oieRbrbo0KANrIbx6Stx63KnHAyoXhLHgAH/gq7XOmyOTXzqxK0GwYAurmZ3CywU
4dFpqPZzDa7aj9aB9GDQQQCHpzTAy5GaK40cZEP42/0BeBjDZtKRCCZqVAOH0y9I
GpObugDXAuMsvjeNsGVvuAv8e69bc1O5AoZ3ICAfWFNMe0GeT52H4YBgtPlfrZrR
KL1pbrdUPhV/TPGnuFrD2QlxJEJzMW4WBj42E/3bqleBlQr/OvaeEKMzFay1/uYw
4dFPptyz32Q+YnbjxD7S8nofEm6DqtxfYvXfFp7E9YaJp9kqtEZf/ZaiaMiVDuZt
kCi90RNyk7LnHnsGDXVoQDBIo5rht9MI/rg2aWapzb4KrB1T1TRtpxT4eUdKM+Sb
2qRc19O+/NdJkkWgEkuzKjZ2MMRFkobRUhm+Eoq/rmmXLulOwm8mTqu3KrAkAa/7
ADVmxjJudedIOH4t/3qZWPO5HUXGFgsSdoYPr6oz7+X7PmHEg/B5Oud8J6Dp57Kr
GzZY3ds4hwVKK83+lj7j/6xSG/5Lzvtst/OTvznAfbYG6O3BMtdoVv/C82lWAeY6
xmeBgS4guxp/yS8tJ1Dj8d7IxvDOilQ3fQdH7KtsZLTKG5JDTeCJkO6rGl42c7nN
QGrof+7P8vMV0T474bqSYRN3H8jPZdlVvRw1Dq7i3pSOGt0UE7hGoXLsKf1QUBcQ
+YqIiYnMsyAPLs4TqQ6SHuPGgVPa+w1TBEhsp+ZPP2eINKAVkx3OlAcfQR/D2Y+s
lRtZDCK8oQ624WWgwq8ii71pTQoECvyR0xMxPzeSReZgsuQoWTktqa9cZaU3XFP6
uJxvsXOGBiKxpnwxgCWnsOoAV/5eltY0ijGs/9CQnITzD3mFlf9BHZ7GpoPYYLRf
StDeLNPOvbtW20EGvQJ8az2ygEuZGIAeppDRCpMrRM4iBNAFpQlV+b3buVN6WW97
rMO8tz2LQKikHbvtmQ3CmZ14MZ1+KrNWwmhp+f/YO60az441bcY6/8oTSzUjhdZJ
J1N8L6mhouyVSW2gy/aXq/1Psxw7hJlJadGNts4KWBq427S5+eaCTP1Zp2FEJbfd
4AKTG6xE38KbyCbeUBa1lxN9+6a5Yd7GpviWbaI9v2uFknNs4jB8Msp+EqrBWUnM
3pP6bzlRt72JwA2YqOrn1ta5DEU8dSyGaYkyu7eiTRMlqjWS1kUiz/TbArTrRt8L
9oxN+ddDYkNl44CukxCRNF+g0ne+irbq+mwycoW0UwtD7F0LfwS9QOLdSB4zJnY6
O1LCm2xHY/RZw357ORD3ITnFCTA8DCv1DUQgrv6TYuRh4c7kFkzx5m/C+KHSmfeS
4s2e1Yg+K7+Eo6lf0h4/8Eiy9jMEr3HQhxfoyEI39QFSxMEIax36Txgztc7xqtgB
Gr8rFCLPCvDFjmhDrc4MS6kjIeQRZ6MFe7ftXeVh6ZSkh0I1Y8/xfFdojN1xqy8q
Bm+0KnPXCH6Yrti0n7/N4t2RGnJ0RPqbpZovo0ao3FF1Mu7ov0qMxT/T5lUD1HT2
Af9sCU4O1sEHqImdalDnJiDl6rtLYWRZW4a7U+LqUh/jBnqzJ0YFbIKg+1iLqmD0
I+J2NgWVys7uzRQwtv9B3CGEwukT2XGxQQSA6/lcu1WU3b9ZiviOoxIUwSJz93eH
QJxKbrfLmCQ8oSEEoIXVdGyNooT6cgm7GQypC/J1/PS3EN0xb1PFUzT5ms4TuURX
r9VT7zHGSxAJBCSpnFwF9RPdCauWwqthhSlF5M6ccrY/anU/RFqtltq6wa1mtybq
QNJlrydiyJehOh7jtxD3CiHoPPxYLQg+g+zTg1YENYkNsj2OVEzy/bgD2H5C0Dwz
gcC/WJ7iSppKFn6bW5WZjV2wN8IDpqFsRQ7oPz7zwKaDEKt4+zX+204jdAq4carx
hfAA4wZaDOWZjAzwUkIu/NfwqPGS75T+vx+kFn/+Y12V+caGkFs3ZlifWnsG4Oyo
p1pQC5+r0EMoUjK/QJU4nVHYUBQ3bnmAkH5cw/5/opm97AdrOu+H49IvIlMGibhi
dU7g8qfhEacaOiM/u/jmJKKiQhBf9dlxeFshpVbVh2u8kjn21CC5tY1+VKnqj+kX
KTNRZ9fWemacdnp72oSeTZS0QN/fb1VTip+gfeT0P0T6cVKv810zhzgv5islTae8
t7DdkCloSWlKPa9xCJJJ9K11/C0M1j+QtczTlDwVzQ6aDS8qSMii3QMdqcFJQH0Q
TGOH1hP8oCFY3UxwOYcnaNINqVobL7/rmVPoV2OVlbOVpDXiBZ72hjDgDHPHVVfN
HcLWHH5SCjX5uy1esdccbCwPqsI6LIqPqFYMRQV+8JJ0Gy1+XFy6idaFtr0Iu8/l
wSpltSXGmVDgA8Z3HpaZxGx0PdDGBVkR0HqEh8fhJ1Enjl+3EunsY2IzgFHDb1WU
WaRcQPjwUnIQLcX9pziwm96uE+sUsQlYGzWTrRAOEq+LIQZTT2ofZRtc5aR3+n4S
3ur6rvCw0QOh5tcknpCvTMLF9DO7dDyyCJX0NOWeJhvBrIQjvKMzcEUrHxSe7gCo
XqxlUVOwAf/LHMPC7E8KlRGglaHwN8f9HuTr29XTzzXNW9lJudKv8/aECU2J1K5D
U1wIAAW9NccN7eYneK/skDhglJtkTGMs9Dvjlkqcqk8sswAMeWmOP21s1GZDd3IL
lvYp5yv+/oTGxia6LNlOb5M9A0BLT0VXYh2xno6suk/pixujn7RQ45ZtUJsYUhS9
sQDNodaebC2Q0EPSCrWNXpL9IxxNv4paPssRPytOBylsx6slk32f0azO6pVABF9l
7djK0sp++vB0L6bPxBHBnu9HjKfRNzCa1vmMTdD7VtmhDDVOdgT+KhurAEtCD79c
Mgs4x7dgnXu7jF/Narx0dlXx2J0v9B0Stt48KBNXELZCQ4ywuJhRPJtGMWW0nYqn
0vxhNyDxm61tvDQ+SwDTW1QpehuViKr4/sT0KwrruZbs1XKvM7QZPOkGV/iC7dAq
BwqTmCT0ItDn+ppRHuddkcsJSmpcJn2HpVaFyTsnyaluANIgNfoso6p51aXdOSP7
URA51bWnL8BietS7OMCFPK7iPxI9ysGZmlB+hZjqAECEMjGV3CjnL9zXYLoLTZ8o
wb0Zi/pTz2nwRteTJvbKJKJgD+DAUmTHjk81h6dM/NuKuBENiPZnfr3XyrVY7DOx
WWsw36hKdgTNr9G1TwoTuuVfasOu7O7PVNFRKlq2N1pUvvhui/HpohMBG+PFBzxF
ecBeYiWMCLUtVw9drHfo4wsw6DzxNENaNP9qN5ax+mNG+KCYDdoUpgtA9/EIlAUt
mQJRi6/TZUzsYk2oFO9iVxJhT8LSv3HxOIJ51LMOUOiMHUY1Kpf0nzveBtZxP7Xx
TRx4KGthl0mpeOtXU8f8/pNRrf7ZwTlaBe1c2PqpwzmuMjd47UhGxt/3mHkU2MxO
0RlxZZj55mBQpuqodM/tWh9blJWlJuS/JcorsgEE+jE93BtJWueqqD3N+tQvuUur
7Fc6XCEFXIR/RyR5/8ERDXfMFlchwRECRJRqoJ4sfVbwgTBAMKjBDcKYt2RmQay9
QKV7Zm0IKaxZiOdsEfPi03XYWzYuTp0wgI1finjDxEkidTNTTg1HBjvPdrR7aMEX
QVJBO+E27ilkYFRZGx3ZhEt7PzSP68wTXBNf7Ojht3i+ZB+kQoRDDC0ox9dN4ZoW
KZ3K3XtCWbYuQaAB6s2hMeOu6dQwOdy2RjT7HkqMbMU8frSGPbUQ3hSMxCxaEqT5
aZzgCB1hP2cec7wvpgWckYJ5reogeh20TtFuplRTQvdfdaJiMlyM1xycN/dsxRSN
fyRJ7Oe0p02KMtf2RI8VM3nWHuqiRgeRa4T5X23llZIwneRRpUD/4lStLbs31bYX
/icySE6nln8oMRkHQylP9pVu1T2rg6C8Sa2Jimhvmb9st19E6Zm1J3ASyQ0YUQmJ
PUJQMJ5d6ShY2FhKji12iUa0V9lZtTUPOTawGl2URYgj3D9lDU/j4aZjpOzn63/+
mEkTEsd6xS4VLvmL8L3/TkxFLe4dqBwyDAU+MqAZ6qmxMm6GDLLP7hXm49v/aMIB
LnOx4s+MtoG8kPQU0Fk6YMhF72hsc7OsGP4K2eJRpWiAZKs50cAWbBZL3erooV71
YUFwt1ys715AU0CEh8kfReq8lUUc01EmOoURRoMn7dHE7ILU2XgnhexQQEchYgVt
z7UMFUseU1KXgNfiDI0RyhS9J2F5vcowNhJ4ZY/ZzmIjFzwuGq6R5CuT521+ipAd
+ig7bTEIHaNg+fFQfGGRrFWDJcdvroaz0xCqmdzXl4XwDo8Nd5GUw1ARLXvgH/oP
kNPwrx0IjAfHIiOqeO1Vl4qtY3pwQD2VfAlB+kYgMXMJkr6hBO7bv8Bpaq+9xTsf
j/mP8US39cf/J8BqhsYbxPIeRYroc8d7ysey2n1RSz8s22IGiy/MC3PfWTKRBUiN
AnuwiQoFoUYKsvnZvngnSwx6FrfUtSOB029vNAoZTAJ5OqR3x0euOf6hMGeKnr1h
ltOd3mHcGUkWEQkS9fzLbzsGQzZG3PPIZ+jkJdhFaG1X2aaUJdsEQ7HLmnfx1Xul
CMyIVutoHjtZHREbNzX1GNVGoKDDQ9ayXmEOt1YB2JwgzpZwDqXVBfOR3aVWGVuD
Kz4fzdWpaf4/EvBZNff1zvzsc5FRRfPyiByytBdc/FZ4mPNTi0j82RyiQ3WXkXA2
bmiGcFmqzXohk3ibzG7g/EnmyzLsMgMVkpB6Cs2HbbNK8gfi875OThGH5npFKG1v
++zqwNkaKXQLVrrYLxw+ymkcUd6N1v9CBqGv35cxpIjB/UpUql41H25ITUllaH/m
Olp6wWgc1obe13FmmXvnvPq6ingNjBxear2lo1XXFjo72+RdaP+P5BIidtW90pqe
lMr7yuxGmh1og3KcXmnzExohAvoEuT/nIW7HYo+p54IS96VrAVuFLTiTmX/zgFlR
qYeK2oSFm2XsFz5A56i35QerC0b69QbtGdjbnQgF9m4d4hAyKQ3U/tHTj1GGZAz8
TqSEDmR26PfyoUqhFBNc/1U9lzPoGxLd9JbTeVZ+yREUC10MZaAEmbnGGpvJYWPQ
hoY5620KPc8lTjjdunipHL+EtpJbi/O+sGGe1QT0dGlfGcNQT+tsbkBY9mpDaXgi
ht98I+x9b4pwZ79oX6rwUOhjCmA6N8NQMCvaQ3MPmgfoc+dZWVm6U4wokTEdqLe7
t2VHoQMUZgFtSqM2PM4IhFzNCifEIiiUVnKe+LmuCmFR1/xSu964vSf9iMcNjMvn
MDBBopWDgYuYdzOXIh4so1Oet9x4hydZffOZUQ3ORw5GrX7jtPUyFimB3BW7ykFn
d4CUQdBe6PShUSJqclvnhVWBUFq2/qswprucpfMSySmVoB2qub9kwU59BN6ek83k
XpR00O2YoxkWuv+mw87tluMYfXfcRhuEFmJKTx/7LiIesD16UQyclNjQ3b++ZbSZ
4OhL1dus7EAsdmx3Uyx20Bgeieu0zmFL/Rvx45nNp1mGsLQFYGSNWDn635A9G9CO
auFqBYc9zuqnQ/Q4cnwNoY5jt6MqeFBxyz3zQYOdagaI4JLpO4Q6PAwSMIP1ecNr
2SKrfPOGDOtucXiaxmeAE03gq9VJd8TGqn3mCelguRC97XP+MDaryGyQTuMpzeJZ
zXYuhdQRX3Y3CBuI871nB12g8+uI8AJ5OsKX7sMrD5zVA7IptXexAQdN8vO7am1C
42szQY7scb0A0slM51OgIe2IfhLfABf50NaWvybaHX1JWqe4l2ZJrDjlOLt9V/7C
zqFekbvpUB/2gcWZcudEzucVCQScG1aZGIDQqhDf4VgMOcJNdSgOKH+tZ/ogOpTO
ZkmVvdk3x1dSTyoSmf5q3naeRwgWRlGcDRgtu4ZA7TFsD9eD4CzO7qGH/MHFwLNR
ODi3Kb5KQ6XlE9iLYoTX00MF/4Krmawib2Lodwy+t04PB5FF8me+66r3pP4fg0NE
e+8Jb605aokKOp6MR5LVDgAf8mHUe+X4y94n1rNNg9Q1vfYUivbDC3qQZQSlUsM2
bFOo/ree0KdbBpJT3aYBTvR8sq2DtJ8Lgh2mVxIeqt+XYeUPWR9JJD7t2liYQSjo
mKi928CD6ghHdPXtfeeJLS/3lTb2309k+vxXY/dCCVhzXGQEwVthMR/w35jtYf8A
47UBp0phg4vgwleGT0Z3os3m75yRKg4nGVLqF43VxMq4XympwV594r7hJQdTgZJ9
1kXFzMnMvFdXnFf70MwrLBPcZahR2ukRHYNsfwGVGkqAVW7GgXH6RqWBLhXt4hK1
+YhhvnbZVtC92GEy64fTd2IHPiXlekXHTjyIivx4xMzLzhXiqe+6u2Ac3XYzX0Qd
t2FeulYfoaiKWr8UR1kkYb5MH1qsPnALvOSDpB5QWdiBPhDnjgjUI1YxSIZaPpz3
IAx/WH/aWwvTvWXGp05lOBsBTebR4l3DgGQUWLj0LJgFWtnDwjLfVOm/s4CRVCt+
YJyFrXL4A+3Ot1aMGBOdSddjCW7WOWPK6FQ8PbwBtOLmgbzIH8RyXCxNZ0GKF+/t
/VB8S2CKQlTpe4HIHeyviF8FhSpEtlQOby6YBHU53qKA/TkgWWcZFZVknCGcTFRZ
HooKKYnrCVWDjNZmcM5Frno0W3D5srfbh7NR23FHdm+VBtED2Q8HvAAmiwYgC2nK
ZVwZwZGeXyUUAMqr797pfRhR41mYk0wzEGaWoQq1sLmhh8HZYBYiRW65YVFISTv1
6sS2L1s12qbrYZoGLMEFjV+fgZWdIJxVC3YlW2MVpo7VRuMKgVZ0Zbkc6hcjlSvh
2Uy2/X8ej8XpgHtDAlVfHOEhXa6Vtq0n2pibXF9jmlgK2j0Nld75WPxOaTO15P5r
FMkLRY1cjIZbM6cEXhEYzLIxscdjebMNSc9wsriscpA9J3fZBjaLGs6dCekOhiBm
PSF1b+xqrdbIxqbO2qwwOfiRLVXNe+Se99kg9jdGiNmiGOtdHWb6MNDCLPJRmAv/
s8y/+9IIxhlQOR0p3Wp1ypZfz7TEM+x+iHmzpl6KVvZYrfAbviDPXu375eDSETU3
Go4TZRbuyOze+Q/RTHZh1HYN1UQqz6tuuB+uL5swNDCyLsRftEYmqe0hPMQIsZ1x
yX1xf+/MJitGa3m0dKfcnyMkGMIsCCX8R4zBXkvu7BpOl1ojb/LRmTSDSJVMgVdJ
l5ZqZ0Zl2GTDLSWRQP8vdu6ht90oYuJvHb9hIKGUNKuG7pobBCY4kSxTJYtDWkI4
RHCsNbhHWnkkgMV0KfjldwogZSNuy6RW2VXRJD81vy9m5cUw9WpcSCopszY0aFux
WApF6tLE7LISS4A/T1mzB8qRwr9/wPX+m473um0mmVOIUbLAR/toMb+/u8ZoRlP+
3G+qLU1LBCrAq2BG1WDPAnoo9X5V8YppeJMEDhjsoQkli0DBd4+zJB5ZvNZ+qfex
qago5UZAwwZqj3AKixC70FFVItAbgpQ0HOhefgCzm68TlCRQJyPzaI60szV9b12d
2z8rugNYrFcqm4Hy4FClJuPYkJZVt4gL30iaSWUIa6kJ5B50JLCLpnembVVhSVEa
VvrNKO8YPJdbBeRrhuN79yigkTq15UjFiUlsYTAWleKzsLuPhkBpRNsEJ9R9ogzS
bXADRDKqe4PN8sPwmQ4EktXPvyV6LtNF6wMJ3I1TkMvUHqrQez7xjIMn2kr2Ugju
dfHlC+3QL4qLT7YepZdrGqRN38eWTPAxSPtgWIqMKJIq2LB6Hd9qN+GeGCw8HgVf
4hgO9CrunsSd27Ymm7oYkyzljrAup1AwMzKgQVm4ltfEpedwvQ0/YGbRk/TV39N0
zYgCa5MkYu/ZKY1vieImKCZijaAkLJ3DogWgmEmsQ19HpIjB3+wahrl1j48G2g77
jJy/V+VNbxx1osOzbEb4fXsQM8BiXEIPqmTyu3u63ir69KWscpm+IEniAJ63MQaw
eJoUw4rCh+LDKaRWjNQnXf7kX5cqhr/He2yFJZxLvlX/XydYCDvoxn0db8Jq01xC
E0/QekJH2GIzhwdsXOT3qkcFWroZkA7GMv/7jizy6knE3R0qG8UfBjsNKw9vqS/9
rgFCWq43pUrMUslirvtqsURptwtc8UV918U1JKRLrBIGan1KCP6UV2YEmsVuNH3P
fYbF77iIqSXU6VFk5AFhv/APZMdrrWPVCJViMyiFdTdx6v1ye1Abu/95iGR68Vp4
rKqPBc4M22t5zHtjpD3OC1PgeAwVBgSx5wwSiCJmP7DVhwcqueQ3e/Tc2QXQ67UK
igpuuzfsS9clCqp1Y/OHRDoL4HLCma1aALbJqyN3tBTFIdBwXn+Hnung7yTa3F02
gsFlP3n/IvE8y9C39WX8jWDX/4q3T0NuU/YUbgNpYuLIO6CbTYMYv/GKfLvLGToO
ZfXmsn4p8XDQk9Br8DBbdOP477f51J80wAdXKI8NpBbWwOZuVriVpIrTWWfkBnMz
065qjyGFvlYoREe1mA0DQ8Ijw5PC7Chcwotk4Ma9DhsFD95xK1l4zOJ6tqEARJfi
0B67p0DA6y+AGG6smvZDT5L0ixWE1knXlyS9Lm4olUnT4MKTYrXcYIewRYgjPAZu
/KpVUJd127WD6JUu8/u4aJbI/WF7QFiYUQjGAVMfg1Cdd9Xu6pbn9JRYtyQOkJTM
WmG+PyqDAYiFIiEtEbPQk8yPTPcdPf0S9Ht0zJ04c1ziQCGLfiLPPoFjJzzPrcBg
y/+3d5/D5oAkNT2ffZPOxpD/qjMZybTxveayCjJItoLtAelVOuBi6jm5Bp7bXieI
ifMLna2kqSw3atjX390cu4er6Rhp94xofF/8+3nlC9LAZfl7c6d6WE3cJczXAtdi
G4auJ9Y7G1TPHNTJgZsOGuReERVVusOXzn83HA6Y+FwLjOIHTwxYNFe0MT9cf37H
ySLcyM16reeqP8WEPzvzHNKjbfhzUaETozKFlwS6ySTzAUSAsmLUXrapReoXLChR
TzCFzP50kDkf2lmlie+kDwSIvsj1iPChoPGHWgIdIIlJWiHN3XwIc07ZkVYLV64W
AIEP+dtocNVqtNR6JPdBvht5gDNdrrUUE8QuXREO4/EosWD45p4S07y90mek9to8
junwwzpUwcGx3njsFlmvjRwWBv0GmDEMnsJV9zKo0uT7ICSQM5WwxohjtpdQUCYO
SNTW4P1SQPT2ZmFmN875CHhRRsZH29tYPk4cVlsqxyrnhj5QHYQzyeHOtsOb5EaC
VAc+OfimWQtL2qSSEgP1OSE1KnHb1owsxAFoKBOVFtMVu3Rph/H15l+x1Ktdgxw0
oTOtklvZS26ki4BmrOTGR2cL9OchLQPVC1TglFjVEPDDWyEfUaEFtkT2GsQxGddK
0bLQj3r47RgYAvXRAYESgVRCtpI77CoMzHX6aQofyzDe43upvZew2DCplEfUYEmV
D4d9S0+qh6/5wVx3OPXifmJBe2QHfUE6mRCdYWao/Owe54aD8coCX4hnlxxRqXSP
UPuwYnmKpUjaDjcc81Xnn5gAKXLOosWQPeNejoXFMixG4TP7VLCi7jV8WHytUgCY
ES1tk0ETgaSXtrxVHyABaJWrXYM0pq70tFrs+D9/9DOUmFjgB8442TQAIOjMMdl3
L8PMQ8U7jelB/XOzElzJ1QUvkm60gv3FxhPanyudraY48t/HJFvg5Yjuh9Qc/b/h
d4iob4cpp3TDfbb/0WPCzlVvpcYvWh9LMjomT1BdRuaF0xaXiy6CHggz82uXg6eV
w5TL8tytoMDXiBvTWWk5EUG7Mee0CMPrGWqmqty1J/4bUfB+5w5DuwjSF5vo7m04
+QNfOf/6Ackzn9T8Hzc8NsrmTusd9Rw3BfDJLnZNFTl/Zp+C0DylMPuJdWAlVeFX
aR46B8lFUpVc8kRkgeQPK/prKi033O0J0E0AMJeK7Ykf1CaftxxWEaFyUNP+geXP
jzLpEDyi4Uw4kgk6QhrDiJTZnRVKJhRHt0Y4d6DcxPjgUVYfPwpQMaJOK/kC78DI
WuuHbvbr2MB5FvIfgbWOlz7QiCeLOrOAOc1azWV/N3SSJOch6oddiaa8WXrp7f7Y
s1bK/HSu8vruk1tyXpfsP9EOJUDM3SyCFHHXW7XTEoGfMhVDZtJib9wEFnfb2q/b
leT5i0gn3lHMKQ+bNym0ME5K5+TEk8m+RSZLMZ9Tb69tfrL86lLMM0gs+lD3kYgc
pO6UlUtSpJR3IHWylRM3CInS6rWTTfYEVHQ5J8kG0PlR7srP6Wog+SboEBRVzlPT
Vba8nhEnMfee0K+3CWSAqKerFj04ZpqlXSpdZbPvkGdHcv6TbL1X9EXuCqD/Lng1
nCCYxcI2wkzdKpbAqhPy/vRODhufCpFAcnQISXHpgslbTi5yAKLovjDWJI4eAb4/
eF745UpVFrjcVTTgC0ZEcMjsbPKB34Bt82Ydlq4BKYgOs0BZRJuHVURfvzMNDBqv
rBdagsVn9b+RIyyUUMLowZbWO7kV+YWW9DxilhimQDE984dNVRBXHKdXvjKY32JT
mwBGAwz8kzfXnZolC+enxOOxLLGqt9tE6AfLSEXaPLWFWlwVyu/aI1BYY3KDDUnh
iBklV+ByMCCNucfX4h61Brcnh17lz20yKwfZvtmzol9xKRrNijT3N2K16L5JhV4l
lxQ/I2bR0PwqLrRcjt3StoheIJI4cUh78T+7JekYRC45O4+zMBk/WNRpdjUx6c1I
ncdyTDxN0/nGI6vY98U0XjscLSp68vHQPopBLla3clneEQaJcbXsUMYrNQ0SCWkq
vja0ICEAzbSwtPQequ5LCylVXGtsPxUmidBLnH9vJsNkgGm0CsD9UibL7C0CvLBs
AWFH4lG96HO/Rm4KLQKRq2hzBJTI2nsZDD3NAMvhigI2m1GeQnqvJVOibEf2JhXq
4YY8KBzl8Ml4R3N8tVcQBLhbqUPFtkslT7G3x5L1t7rlNaAHJfFQRRucnvtrYNmd
FlgmZNvvr6Id/ksm1FWQwrNhOe2nweTRs4i+4W986c7TARksZyXJoZsNBTnx+Gcd
Yk99yYTsSLsM9MMY1gbktPzuwe0bUeF/XW/U/uZwjJ25z8OefsXHVqxgr2FbhHDb
0z11W6pO0Ib47A27UIekxfKZHzGd2hjtJxe9GlsD16rE8N/zsD8BPOzd0jEV9hz8
4z5jFbCbTsZMPYYr7X49R/CWMoH3mpy8YWMwncXdSdaE995UpcU3K6xYawAAvui+
V/50L2DXcmUQi1ym7CMFFmUvXOzp7GVLIHQHAOiCjg1Gry/RTVX4/K8YTz3XnCiv
EwPt8UMABfsP6FzgkhBYc1wkmHF7R+eJZ1kuATqw6F/5fpmoMi+wY/gIxcbChHda
nOOoGQz7rv/2jXl1yc7wr4RE5O7CZT2/TXau3XZKhOdD8xdpQ4HvDprIbIn51we5
EnkBxaz6hqgv9neEN4wirdbl0iY94Iul3L5e6J/7SF4fxKy7CCuoyisFvqCxqhNB
9KXBHzOKrrg/HG2arT+h+zZwC6Mn5trhRVFYjswZpw2OsJJ196gBj/aJT6TeWMSF
I5Sd0R2dxPfjw3IEz03bU5Pp6b9ohffRz8ZwuXx/ZC5ExvnAjSu1Hnc4IYiM3r/u
rDec/bDwsz4xmDZmOLRsiyiMwLlmja8bpZm7lR8pDB57TZrAs0jvc1/Wv5QKWnGH
KjD18WN4CU8u7gdMyE3RelHVtFscSFN2fubRoEFiB6FuFH0ZioUi1uG3DGL55Wlj
CRqH+zoCYfMhg4e23Gg7mlhk+weNjWMvuUGsLyMrLIyqV06KaQE6ZsAqQ5L/Oriq
xValdxRr11Fm5KH+WSARcYoGXm3Fna5xZGzwTYDMCdy+c81+JZnyTtP124H8z2EG
hyJaa7HvxPoI3rne67U+64QfVO0u/dYCQVHAIjEyG1G3Xt0SM0J3L+kshmLbTx9w
ehbSju4EN7lgMYHigskPJjP/ugr6X23fygY6vGFPrrF+vjYn/Gj2XhiKsUEqn4Sl
OUmsEZ9vXSgIBmLkgdQv0bMdIAGET7xKDNID6MTGoi6/ScxXB/q93l/ynPeflKWz
Sz+m9DsDCYHx7HNHPub88oMuoOIfb46y940K7aB64ZVmtlVk6vWuJ1zyajFV9H9V
4c6fw7iRag0gD0mKihyA/RGgpHwRFiRhJgWDEOTBp522mMiKnuCv6jjRVAJSLtEO
WjA51rqcJVxpYADdCDQVp2yrzXWaC5g0KrIp6NtHHQgdL261bcH7CI0zK1nNlPEj
Rbk0c7ffEsKgXlk+K0pRppx7NiYwQMkr91kSsDhEl19QXhJ5iDgCUaY7Vysu7qww
xT4Jt830ckG2e+19YhDhKz0+Lb5UmBE+3A47WAx/8LUQMQk/8L55if/ZoPFG93g9
yxgua75cP7b5pJiK+n9kwsYkAU3H5xPOeA3G1DlwRMwl9EEuF5ddg1MO37zN6dd9
Cj9llJStjqeFaxZyx6NRm7HcjWR5QgsELIFlKwTGrnAfmm/uoqRWcSHNfdAC1q7g
SDyMuR+TUq4L/fhwB8UkMJm6nE7Z8zI856v6nW4DMckFQ+dGa4UcHEZ/DHgxSN4O
4pFNY5zOUaWcerXk+dMqWKIDRh9eD8t7Dlsrlqsfw5a6qa/SI+/fUBZnCfp61aL4
4sk/XXMRFhi8I/keMm11bB7TDvsdzORBN4MrOV56pqZbzdcb2T8duMOS3Qe6FjyR
E2E2BhPPLuJBQ88pgjSVUqHRtjJhf4FnILJEUwddUf+G9RPTWunjMQD+C9AUuL8u
hy/zNU5PnS3xY3zFYux9dscy56sDrJ0T8AHUQaV9qh9QRDJXOBfHbTvDrMs3I26k
47nBrv4m49mRiMAnzdYasiQuHbTFBZZWuicDbqaaFMJTfNF+8fa0bpX84UOAvIOm
Tpv7Qn24Orf7jkZ7SjnLx/GxD0/UHCMcgJF+SzE1F9p986vWU46jRUxjz/rrzNCb
0D+RihyQFPSrBmxwM7m+qyGQbRLbtR2ae93gy38oDGDpDoQTu4+6GVMnw7kCJ0FS
647wZvoqR7DnTSagmMs7R1JWalvil125YG6OPiufOT1L8nJVa+//6XA3HwyNFgJz
fUHy7KvLk43WFcpPnBb9L6Dr0jdcdrG4wD7xcz4/v56NhVCxg5boiDXeMN3Hvy1a
OmCWIpNp+VsaDALeR0AMVq5P0On6Dp20M/6C209HbCq+6q9RjH/NzBFXRSTsCNvQ
UZkwRek1bPQbPuLhP2O0EuksQ+PywrQjXYzevMr27/wjTRZhCwbZxQzzsNG7yCSR
fFv3FzEvjXY/0mqkU0ThTi7QR/TogyM17Y/TsclmotM95z0pavVKWZt1tllghsS7
6JhI/T1zVETSAhKe+AQupIiIlj09aGpLksAf/b3DiIV4If/8lEtku6TzWSjm9Cn1
TuiQmMejNiR88sSQLS0CM4avSO4IBPtJW6glQ3BRsiShtjItb/6NSZMHZczCeWWk
W5MFQ1sOsexEblE1Y9BLfrWMZHBlCY8tdsFtvITUFPOyvRYfl2D8GAGQ1LWcDmDJ
qxfeLl04gVLxUF+kNCsg0CNE6MPOHEgwTNp3c1cJ6R30Fu/0pc07GUk4cfxB+GNY
izK/cmf9mdpBdcnOuQrGKFgRXeuu8DuwMxRar28MpJ2hI7RUMJ6an9fqVVyKA4/d
g0fqkK/F/a44Cr4NdQ6My2H262CZ9hjazJSn0Fje1XhPkMzfTL5MrWIXC5c5e3Pp
RbVgGMATD+GoBbK3U7+UV4UFwb7Yc3QqT9xL95CrzKJiz+3JiEPicIUHNioTLkVj
vWlRXO65PQLH6bxLN7RvfD2GA0HfPA0Hms8zKR+AnBPBldXI6qhdXm+Jklr+wp6+
kwfcChnS+2CMHvFtlX4WMLMiNKsF0wej+HHAiiP+dxyTBRSUDUYbWFuH1vpEUPZ3
QQtj4MCCIAG9S5mQmEN1NLXwks/5MvOGuAx1/FZvFFkSCWavIGKhqQcS78TmZ1fV
dFQxb3YHRmBfLjl5TSWWKjqfZJm0MfW+KV9G515+Gjvv/AvjioQi4xeiboRw9+BK
Ms6RlGQKkN8FKewyvbYFMc/huwy8KFTgoXsfK+r0DIh5ZzG87fJDFo0XPuYWQfaJ
bjC3jZ0PymnZjEKPbEY0tmEC/6LRXebV+VoZnQ8+LXprLjIwldi4lWrLNMByVhiH
sMx8xBwshxoA9wwjHhQSqUMknk3Pne2wDPMnrddHFn2+Xn81puPjyQn5HK+ZOohs
Y/xT2qAABUe1tGAdSftewf/INbbbaBEECHtFfiL2VSCv56lBxYzFXogX08J8HceQ
oIbwurtk+Vp5RkJ5TomOv9U2Iwv7wGHO8SMA8wI0dxfQEZvou1TwfSeuq4EMmazJ
QMAfpEuwTxhLKMApXndSvfK3pP3/hPflgh+5xQ0aTnGI0m/gt0v25MVLj68mRS6+
RBggu5goYFGRNcPa+G/XWJNv9By+U/NuUz1Or1Y4/e+S+c4iK+9tMKHW2eDDCC0D
Ta8An84E03ZpL+NSczqoQw98Vg2qG9usWu5nWL4hjG9BylKfAr9wx3kZ7c8XAoSd
K5MD0XBZkkuB/ZcCQ2whAZeK4+9uAKAXSRxbzLh9YVEB7o3YQTN2VZdtuwvlPrXl
ML8Kg5VqGivARp5T1JeO63amUduiO9IE4tN7ob3Twr5MLTnhUDwwMbmrYuyLT3h1
5u6naehmXGOHz1XMR+/FBhENOZ0uHuG4usfsaZW/ENprXBNqV4IInUjtL2Lp4sdk
kKhkn1Tf8r5GQwUyW2mvsLyI+GqE9AIxa1lK62mDaorEIJ/90sE6BLnLBP9Tqtkr
3cXw+TGS6zIYfg9wcw8E/i1MsPtNh+nbZxM1crFgw2tQMiHBZXg4Zf+QMm5AlqUp
Kf5ag6IcKqrN2whw/HIc9cuo/zwcr93+aO+iVPzxWmKszYWR1wzsI35cQZ83zfdO
cIsA5iMACoj3XAT4P2ojOxftWBTIdbb2i+zcH+Cl+3KZOXTtkX058qeQNVRSBnkj
+RrPRKj4kh2aeDwP8uGe1EhqGwe+iRAYFa0s+BCpuLloFsnod89PnHK3AfIZUASp
jZw1Xm2PH6DUDN6EUgtBWYGOscplW40pbt4wngbvmYZn5cpk/pzXS3h0dY8vSIlc
dznlCOgjE1hDZM12CbY5TgXHIUuM/MhtUCGkUx/Ny5oalnx8xxB7grbTTbnTZRFh
CdYCXAcKZ5TnUVmrEkXD4dUzIdbOv3RN/MPndAJVZAFVg1kYRwCAguJha8knTBE9
XmfQiZlSCAcXWb0fzt4QLn3By0HbGXH4ikYLsMsVHOuzKlXwxhIENXvgbyA//xv6
lm5j/HOuc1zHKfI6L+LN+Q0uA2sc17WSDKS+ZM+paO/NCetQ3Klr6mu3mdW+YRTA
8kLgRxRSvP6/RaVXApmBBKsuQYXnPP3bEQUrViLGGchC851K8lx5sk5vlka+poPP
tyYHtpHAdGOfFy42KCSiQyhe4Skihj+tqt6+9AiS66O3tnasK/3NpaM4KByTkkz9
KOlDVWT2J9nZckNDOefzkUSmPLr9QfHNegSS+nz7ZwtP6oOTC+XO7TkSsGdoeNVw
Ko7SUcGBHesVtP0372zf9Ag/nmqeL9qu2JxlKZ8sN+v7XMdI6wqn12egxy5Xgaac
RDwNWCYJ2p6mwDJ5jkMWXOIr8aX972b2DfmbVfBRVM7gDrJJ6XuvrHKP31rFiiXB
CxmF7YJPEZMxDOV0yMAg9MoGvZvP2kZQof8/ogamAWJOG34nt2bCd08ezwM7b5c9
i7fBG9B5cEFA9hrhYxro6+RE8DA0HZ688k0A3I4gqJG4ESfDZ7xocZuN446BRBUm
3TXQVkGin3gPHBVTawebtcyDvfXtGEj1i5w+vfjcsMtIUFsxl0CEgsenL+jxY66T
eK4TeQyFBwilEZ4LvT1Lu2YZuHxVAUa1iUJLkOkkN/AbZ9K09A7UCEpmy5ESgGwh
GL8UJawfePCkasFPP1E61NZBmSjv+GZ9waHIXFo9+AS4f3PbUhBX0sj13HIBv8pl
fCkDu37J+aRZZ41nxW2llM478nNbdTQkEGjkZ7FCirJPzTIOhaZO11DlxRhSOieG
VV9EZL06x/S2phTAzqfQPqo8Exi/uZTYQTs1QoVm/gVB1VZ2gx14tTFDGA6jIhop
N7C/IC2r0fEuLSnADiA1HfvCDoTfcIJV3EhOkbP6Jquni6bwp3hogxBogODyJGdv
izejNokx5RUk5vIr0cIxMcycrWx8fye9ugC0d3I/soPrv20Wu4I1JI1qG7oiczHF
dgACCLTe4kXVOKpY8q0itgSfsAFQRj7Kvh9iOMhkfR/O40gtkW+krDM5BGiy7ljU
MPDdM7DBemD9MtBfO/j0rf3GbzQLNmhV+91M+CZslEtU9mp6QKuRI/j3g4aykUO6
YPdLLVokYrLHvW2u6Du0csi1koyvEorQVpwc5ouBK0qu7BpX/B78O3w+4bbSoqfd
DbR4ngt6vMROkPrYCg7Nrso1LrZx56vNKCbOfo4tEU5Msq57mhrHvBcZ9ONM2Unl
wHENUMEptco7Q+b68vbCPQOQm33UBymHif6O3iAJbS25fSuzrVPOHAX7Ra9/xMUm
xOwdhanmPDilF7NqkmB3/3HmIEsxFqR2bKc0y7jRwsTu9GNQGZNS8wZecIY4oWl2
wUTaHRpkzrv+fuSZYXTLDhtsv3+Nwuk5eG9A90ENNVVm8eGhJe4hbgtusrDrhEyI
QEgHMcg3/2xUvXiLZ2lW7uEh3eJl1NlZ6k69amKa1cSHV1g0AsJOcqKBJu63oV3r
ujcE8ueZEOzUYxOh+lXz3LVQKzki4I5zyG6jvXu1xXO1WZ0bijztcap5isgfho4x
XnLzC5fIkYMyResZzhOfueSwIpgye2hRyiIVkt/+QiT8c4JjMBqaDa9uggMO+00N
BP8pKVSQUSc4WZhCnZPa1ir06dxkYbsnCrM+53D7hPWFJe4ZgLy97yqLt6QYV3SD
zQ690y7OHB7U/Jv0qqUEdMpZnkgOZkhcrLalpIXHZH5exPtFqU//7wk/6OLXdiZp
RwUf91hJFzHILr8+ZuBM77DebiEWq0F1LZsGd+JEz5HOsiZVqDQE0+KB17QGgMee
p6Qjsz6nqpT1gU7E6H7IjmvwVttQ9B21p6rWtlbYZoiQwvFzBLXQfA99cmN3AQe+
RTXKsoS99apg+4T+y7nu/jXMLM17bfZ200quvdw9lWKRGgSpZ9JbrcXE79ObaExZ
0BRtmKIXL9bDijwcWTMBzxD97GNoKNOODV67QDdRnLyuMfOF4PQXzCoBQNohn33N
ulmREjpHplEmMeOGy3G2gmssWDSjpxh96Q7mNxzOwqFldkBSUJPWAKqK1dDGAehG
qu0VzwUldMxs04EHoDKu4LoILfiGuE7KI0rpIA0VVDtz1WDNqrauh/pdRromyZZ2
RkdxgyfVATyNOdLnsTNdfv/e6lySOjSN0K7vwx+qOtmULzjFjYyvLzrP1zl6jH8R
W+/gkv93eP65zgAJ2QcPYWOWTxRSxmZNZOHug4ofBN9cqBtW9hmAQjj1qAsr7LkV
fo7hT0NZnTRosVoQGYEw9Pt8ZGwd62TbJOMva4g+KuhehsVlimHmFTMNJemPhvyx
lkhU5zdVHZAxkTLpHxvBEMCZUzHuvV1gxfDVQRHVpPGKYTh/BEAOE/Sye9Rg/yAH
Ua9FdHLwKJ3li4PXjLryQ8zfE5zVawK6ITwjbL7o4YLDkiisp12l1cCu/BX7sQ0y
xoojWt82ABhsPHnAOoiY+GA473TbRhwggD7b0rwFAfui0J3DuFK78tY5pSPKr2im
IZRc8HSshgplXT7nRauZea8pLq9uJdmSbSVkPXoaroEq/wiaeu48Zbshrx8zCBn9
JCvymsSzQ2Xfh/edRbyYj8HFl2JEJL9c6tYJbiNKBAs6s94ve27OOecfr/8XWCnk
R2RlavO/pNraqxTCOqDBPTKvfPj6Xq2uUf8S5bxwDBKF5vgL3a9uzwa3IK4Rg7ZQ
SzOoNtW1q0KIbA0nQpd88Jtplnlw20J9NqkCIeHsCN49IyF3nVKPiICodLTWiNJC
ezxq2xib9rSXEXYVuQFG8vFRLJOoTbqLHh1vo5qdWA1S2XLSHjZwq5I99YniCcO1
0BVCXMWBc9dUQ9D83BSXlpsCWbpm2NoSz3BycL/IwAk7sU24rGk/lLp6e2L33bgi
K/pAqnA9lC1fmX3u3yOQ6ENXmVdb/9X/Vw3jXfxzA97qR9Y5FbRdFxz7Z1e1VLcw
qS19M3kzFLYS/SNbW4xj0+U+w9z6Bv4CIl9XV0GglrDQgOrknEqxGwEjP9XWxo/T
m8T69dfINE5K8/MReatPTgMawb+zXZMuWQ9QFPr+ppB/j+lsav6c3RY9ljHu5fxJ
TaZEJANakO82YpIohExgO8FnFpYB9cQKEdF6N8am35SbSafV0WT8glkJqJOCc9IK
XY8r7MC2cUq1xJtHqi+Mbz40dFpCqYASL5wpW2KHEw3WsBexkwCxT4r6oTdlTpzz
M0R1beVmeIQQ7jQOOe1vZYb3kv33qyybKYlTUCxp95QuWTCr1JcUGOGJZvE3N6D0
NShmGaXsxuYJ6yxVzHGLdT2iGrSFHbD+a4eAs/WLoTAR2YOJZpc+a3CLXlrag3SL
QHEcG7Zas8Wh/2YF5mzGiRUW18qPT1uGAHsOnvHVUQZsjpj8B6yaHIi/orPqSm/G
kbDAgJRnlMm9tCJIxrHsPPKAyCrQWVyCQo6UwCCIoojjSe0BJUnmACkn1APZZuNO
RCaYSgJ1viCGZmP0C5/8MlrXV8pRmJei/kX89fG9CqSQkyAy7RgekJ7Nsf8NBj25
W3AjVaGJY14LB49GedeEVmyiMN0RaFnIiOw2xFxSZ13h0kvaLKQ3kk4x5Msg9Y3v
oRvjUKgUZjM/DhNPOYe5wJ2BrUeo3U/z9IL3XqT1yHlur8D5vYcfZ2qQpJRHE549
rC4VyZ0O8h3G3CoP/s6q7lv4N9RnWMg0jWvfXCcc1dQgDJjDpF6y8uUeATzXmwEG
47vifybu9l2t8YjJ5/nMETcaGRbQxhpNjfks5qt9fdkMjeV+gi9ijg82GF5Ma7EW
GEpi5Gh0PZtXLSApC92/lI8nzGd+ufQaifAChZ8u6TRO0ZCIh65H0yvRjQOY50Zv
jXvyLojHzTnyytgnhW9nJ+qfTCT9tEKcYq/Lo2KQRupm0noO0UfsPod5I1tumraK
ixWKbMPRtd8QJA/wgGijXiHot0L2qnsqbUUpfs/C0B8X88z3Tr9mfXYV4ArqlJs/
dDgkbxfOU8aup31he2ps/Ges1Q1qUYTOaUaXjC+0Fqok2hzmBNOKv0vcztkn7xjY
yE3QyF7G+JTqMWsvutHMjs+Vm2UNOEvmrg05SVaIX959Hi2LnBfmSlqR8WfORubw
EDV2ORXnCq6nHUvfWktieZGeLM+k163k4t0A9atHJKAQwfXe8bHRSsabvZgwRnDm
av6u3n66Dv+o9nLzxvkZZLJshQTSSo7q6JBMbkD6Yo5mMqvra6CIQmw4OS9al+su
uauvKzf89Zr13BCcTLsH6p/mWbF2ufDQOrsIvOflYmso9xiS0tzVIhchq5jKlBml
nqd+zRjYZO3qN8kXeqbGlyJgNuu40Ncoq+8/xwE/uDKAkkEdt4HudxfTT5vcru+J
v3NG03zUeuSfHz1xzQ6isDVGvtTIk/4xXDjG3XIY2yHYxRsT1lNFUvB6wopPujMW
aMDTpWakQ22LsucwZ+cCtvDlJzvKfYBYX82oTIIwtX3pKzlFUrRftbXkgeGnaF7a
6nrkK0sPTdPcxRuWAew76qYhbdFJAyg5snrJ0qgW1M+J3OM2YSi6Qrd/oHOhe2ie
j+nf9luE/bsogKsQ3JlRTNVTxtZWAi/ryfhVqsqV12Hcde71RLJQClWBQ6jc0PRO
i4RM2Js2W64CzeqvvgiuICopNyOOXf19IKoodhwodSZpumYUMw7AX6PRqmE7VMlu
xM5Mn+i+3GImM4iM0X3akLhyuuaYq31HQQCx6jOVriRpWxCf3KZCsAQ5QtBLUmfZ
L4LZCZVMHbnHPri7lHe8qnAZVor7qUxk0jJjdpTSoWKcBlWO1NBWmjYugNYpNXpO
Jbe+gVGU+z476fcFK4FgdcGjdGk6e0xdpahnZ6YKdbFl6q0nMi/qOdm9xL9h3cQo
rX8oRZKP5R+icrT54NanLt6ih0LiWgHjHw2B68AXiP97iKtyE8XJ0Gf/RsGT1jCY
lhHts3EIZPx23jVyQLl0PAc+1YHTGcvM0GukG1OTaqXQ9/MII66W8UUU8NZbdWH9
poRYKVXP/YqYBRm7L2tCkvujbxAdNKAj1v14b+bShmlMtXwv+OoyvmCVhM0JFBGC
5a7K0ZcDICnpz/FtebEf10x7ca275G8vMW694Gn+peZDI5jz5zZEp8xzR6Gn4JGC
A9Kld68iPzzQJ63ZPSOmggc2rA+SUEnncdQlD90uG5MpyvVEOsPOIKuyWq9NF6kn
eEMDSu5zeyzzj4FiJqX4D2d/Lvx3z/2O/xU75b4oVzugv/lDsNSqqof9gS8kZSN4
mvW+Obo0ARoOK7z0C03NLGXBZRXIzNc9JB/WJ5vpcjbkFiZ3Bk3mCvWqMka9eoiR
7hZn+HUKxzYOYSJr5OukJLEAydNeCda/DBBDWuM6CHaXbSn5u9TZ9HPBmA4N/Jxl
Z6AtpwWgEgk1pRLNgYrYxg5CJepTZCecFUshhVi59ZEAOUw8oXxdDlCWEnCbrC7Y
gNmXWdh/SqH8V5RLqPFgFtiMelWB70utGZZDjL6wYDNZY0ILicz2FrATAqr+NYf4
95GdBnG73axJCbcyCqOBqVjvEGU9nBoxa2OWq5c/i6mR6ltd33eeTa5U4tG4XE5R
TyerzYJJvFJaI84xUdq761tRKXAISTaoX/gWc129+Ey5xyGxBtSEwC3LVPsJxyde
14uhXobo+X0u+Gb0QHXNxeacu2HzHYGRaZlgrHETr/t4CYvUaFgdLKljCNNLc26e
Eavp+ObexYFy9mdH4ZWhi8YmP0zIVRXXCNk9PwyM+JOmW4N9+n2s5GJ8NDRTMm99
GjwF/cZdiYz5vCdTZCKtva5Jpft35AyDfAZwggRXtjrLD/IEQkiLsax1uhulYmon
LcnT7kPLzix+2EmeyrWBuoXPM8VURI5GXvcFDapva1wsRy/b6kAQffYaaOKrAeFO
FbkA20bO0KEfl/eta1UM8v/3EXNTlWYfF1gtcXMvhKfJNJ2aMXF53kTcpveUmoV/
vCn4Hpv3bFQ3d7a5BakQ7jDtlcnBuK+7j45Doa/n6zW6EmBvT5UPgodyKJExnRrx
H/rFmdRV57kBwDDmty70AZs5tK4nTtNNOv2kWR2aM+1jihK8pzcCgsTdtktWcRcL
XyIMWYPCqxZEzg+DuNyV/kDvZj7ZZ2M3cBFbaBW+2QnC4ZMRe3+Bar7/uyyfqLSt
V1XCt3EPrqNvYkh4jj4boUDEbQ7AuRLabX1uBEvVqE3AEss2hSYVHSyFA0S64B0R
xhlme7Az9danfO+b9yD5Fh5tMv8rdkHA2q5RENultI2vtdfVQWdEcLh03wXfVPZW
LtJ7UTwL6T5l8Uc5O054b1beCf0y3Kj0umNUAobZsDkLxHr6e25lIDRvCjLWcvr2
+ZDR51keQglU0KTRTdfenOfuHO2b6yesWBmSG5e1a7mDmOfdNk7Ys2O+toKzNgRc
PWbh2kf+DWisTbj11EoFoUS65LUOIUGnomlhHqG0KGfBLMgfYw0Ud0kxnOlDdv8y
2Mu3qiNfyuWI0VWo6oaklrJkUN+w9TvumS5LEK//7DuXs+qoD4J4qfY74zwkzkMD
9TSan9n9Wx9GGgrnqy2iZjRnd3561mHJ+Piu2sTB1BOe3y75YzNp3LGPyap7Hi/6
DEZgfWdprxulZIErSOqxar+INhHY8HTuDR3l93R2psm9tOBXVoRjjsvWlVXLK97K
fYWC5QyCTyV95dml5SO7wTgluzmqv4Vr0hJ68HkQ027jjcaSAHpDIn/E41a5lR6j
4FlvQox8ItHcSlsNp1yNMzSDfMqN9WrO7/+FFC7Fjosmw1zQn8blevUGtIEua3vL
xXovXYrH4/JLPhJ+AIoRjqI3pggJ1aC+QhrikD0RChwd+4kgRw/al2FHQThj4ZHt
VAEjYHNQyI3MHFxm+lC5LAJj7OcOaQjIgyPEh7oHv+9H/zvHCzPLU+DkG35TPsyM
JsxUfh400PMosuWkKSm7NBWWRFz2wtbWh4cScM18jrQ8QXe53/+V4+eNyvgqPQQ2
9OsNGKP5TFBLjGEHdCGXOQLJYX4mFGF8+TS4Xq51OW3bgzSNx88atTceb0gaJ0Dr
ih2rBxZ6U/dDQoo+2+K1vpfadVaxI7JhQ4ipDx3/kc6S2Kq06Si3RKg/hvwIPWLU
kPZjA6YGpy/s+aAE0eI5hSs7H4gbNw3KUWlnF5AFrQztz7rl0I2CLsstsLSG07VL
qy3JQpuO1AY82qLMNCnYDpD6aAWsBgliQGm+3WQDPutht7q2X4Z7H0oaI0u0N0UD
5zX16dqo5DAuZQCpquMRpU/YC77UCzbW22A/IoxEE5lhZQiugnN0XBiCbSIXJou0
QEvs2dHcJR9w1Oz7LJHTLnZLr6K3Vhgb5h8c0lPJ5QM6E45IYWWH9MZf0uYRbO0g
apOSo+Ja640H1j2Cmm8JlgYCKwrsxSA4dT7BFmvl4MsdXw93He2pqf2JVwwc05Cg
mGRYrYSI0nO2rW9FW/2c8TECss55uY71kmBMjbykOvcwu1Zmz0PavWYlWD9RDPYo
I/nay1viSZrZ0LzCaGC0hsySAzI/4n5KzRj7WQA0yIefVhfamzHf8ow31mjzCWH4
QtAJ1FL+41Oq/8rhMuL3RKAayPc6R5IbIj52bNK23vgET5rlKh0JaKhE8KazNe/E
n+00Td5A8SP0FZO5iy2e3gdlddQYkyi0BtXoKk1AA4qHMvVzbjiKoLxPGbZU0AZh
hrfVuplMEHEmkyO0KpP6uyNRJni6U14Uzk1y/mCJ8LpK+lfddHyuc//O25c5MNFO
0HN1ZSs6t9SbG06xYFUi8wsMslwRA00TjFfC+OlmdPy7ym2do/KI/Uc9bbUtFrEP
azVFjf+fOPDZCOBUKREW8/WXOPO49a2s0IrFGpxSbaJPFPu1/NUH1buQ1bWoQOX2
fMpVYM8uqc0YDg3CQdCsbogBbxHuYrCur4T/whDjNKqka/RzVWW9w1O3Qkk2ooad
bkRWD53YkVutbv12oPKrjHFyjCQaeNf0qkIVabNZWPthogdISJeSxGHpTciGsvwE
D8wLGb/MOyVcLCFCLVIosntBGExEKkYrJLV1s/NHINiDfQC9brw8qKfqQJvRq8zY
RByVvOUEYxAP7NRcu3fKbhfriF5K1U+IFjKrUg58dUrstDYpQAh8E8K1+OPHBR++
sLOaoXAd8XCCnk1oSDAVpry5XyQ4vv0vyZre122ONziBjmFkqT0diM7oDdSiau/K
/5QfZkHMM6+LVqzZaSCS7Rd5UGcKkzU0OILhkLJgcIeGlIpPWaUyGhH6eVrqOzqt
WcCCDu/qY//gBMfkT8VKdqPtqjL7axUamP4Z+Hf3ro2T4i9//b0m+JF88N/uCyYY
QLei8AIQLCBa4nIACPdwWOZdkI2EkuuAn+LoW51baJIKbNARJWcRNqg5Zv5qeT/Z
/U4QcjA2mgGiHNTs8DiGeABY3Q/17CQUhJfOa4dwWu48KNpEvGv1M7A7rHAolttG
Eaw+H/bVF4sC+mjAW9soh/MNvDzerYNNmf6cmpmg2EeFoHU63XhAqjYjuDSjBxfw
kVBwoRQ2x88clNf1JO+sFJgY31j6e5/JDmM9oqvbuEsAFzZqxpG46+bgyo0bFBVA
adktMzR7UvTTo65D8sNm8KkyDzl4LpKUf8J3TZ5I22lXgoaBBj0L/d9HwIxpDi5r
8oBQ5gE0MIc/+EOn5EdRSUpp6JTUmqf3/LJ4Uq4pm97C0MBDydkTol8POiq1oBqO
tDSXpyYp5osIUEelq7DwX4kCsqu0YY56TIMBJrjtBFKZQw5ZHIQucRznfhey4Ib7
052LiJJLVSkOlEJF5lhuUDpzmfSe0YtE7dATrL4lqsBqUevNm8zILOmIv36AQxL3
anWANpp7ahw2JAHWQCPVqIZtoJhz79crrVpztirfn0gZg8Y6UOJDfG5KXm91L1Uq
lhOjX2bFnhHvWqUxZvMTh4JQ2Cq7ICya2e7S4aa1SSfOKgFeEnNPRQcziPzhxnbQ
I5VevhMkzBVavhQDSZgxuFXblQ+DlUBCmjX3Dbv7bx8G36L4/m+tatVXbOS9n0qq
tdoG9kGQEWdETuEkAhvKqa3y6XFYcwpnUGqBf644Kxwl0kx9OJzBS2Eur6T40Si2
0zONXFbvygNFCzOIuGosGWTCO0HhdMCytUTtaAeXRIBvfL0N5ABO6fKRP4IaqCrp
n27J5Yry9yANW+JB+R3WERqmQxF34XvUPCKQoMfZx8yem0lJsonTj+J9DQQssUk6
QKJ3+3NF0fZ5lUETd8LDrsYBiYxz28EoHMWrBTuCmVZP53ccRNWtKgjOWjE2utQV
PIY68COAMXHVsS6wtXK+WsZbcPfDs7dKZAxY40gEJ8cpQEXE9IQbauIv8XEPnagQ
Ni60tUdD9lD+wx9sifF/UjwOxcg/4r4JNgvFAYHZR5c7zQpmobbO5a5tQt010B16
eslW6LsqjvaHrf3NRylaUxnCtJDKebEbaUymmK7XEUuJYpe6xYJQiuuHhBVyKJvK
HZ1zyxNdERayWCLYNNYVZBed52NuDoezi4RqwEahLiYCyiIhh+gQLzWr/FX9tpf4
8+9CKd+AfgBr1VDeAIP2VrA6t3UVEBpZrBpz00ZCbANUnfwhJbY64kFpBFpXBTmE
LW7wbKdXJbQHmaGS7o4wRIf0YL20Hp/ByVFo5vWU4alDuiN7r5MU0Oxx6AFGwGgI
sJwDCz1UMbnm3udWwRhc86D8Hjzk4Zbh6S7Gxlpsh3zUkOU/c+KvgTg9kV8par9E
1dA2ASvKfwJNQ5+hT/gxzrMN17nWPpYq324ylfDQ00sOfIYUs6k5FP1JtHDGFupl
s40nLiRevWVwA6selEdd7VU2Q9ur+Ik2lMLl/gm0lX5JKxm18nbIUOVSXuceJlDt
uQ106dW1XUyZ8FhasHKRAOyAw/a5D5ihBJH/K/yGl6qAVpGlp4OcWfsdZ2URokAO
jlcdDrW6Nlk9tWQK6vI7CmluZTYIPmCSV1zJclV53UGHOzg04FYki9tnBFaJg77C
45+nf/71aZqx9jFamyYdYHiikIiIHqE8dkz/snymXeMooVa9NOJqyCSgfo21de5L
X66xgmb3ZEeBtgLlcjHZytFiJLR+Wp4i4zzMUDGsRd6XwbzAnNnMecq5RGKbJj82
cJqx/T29M649A/CvN82PMWoHvaIeyJyxHIHzuRTxTvUKCu/+yGpt0lYDPVBGTx0x
8awyjjnXGMzIiE6vwTJ+2DAfO9kJB1rniuJHuII+yON983t86KFHPdLq+itLCgdN
JIeJQzTmFTeh16jA7gSN3Ri+MAjSUGD2h0Irq1MSRns6C8oQmRYN1VjO32Q+OaL7
lQ0DElJdlyjdfJZJUnTkA8PTk1gLFxojWPegRNEPVul106frvKliedA/fY5GqcC4
tzhgpJHzZ9TtXLG5YWGS3Y6lmTYDJ6eGqe2yLaj2hq0XetNS2WwjMPKB4Xstl9IK
iqWAUEbMTfZnboNpC8uQIMw1EPplRsy2JA78C9g0SpqC9kl1472/rjihaI6na23r
bEA20Kr7jvXekeDetTdypiFAW02+xoZPrxEgunWuSzkiPMuCPwwIzeNPPAk4myUS
hHzcwLQ6dWkFaqXMMPX8LcBcokPzf3sbftK044lL8pLQSaSz88V5WdFAOgoHC6QQ
0K/DfKXaLLz2GBJNuTBMMMHCSRU/Dj6RM7/XdGyhpqqPFnDI+XbWxFg8DDomepW5
AATnjOp8JRATzRXLOBGz1iLoHjwdNU0d3hMBaWgvtA8bbk79XMzdJnHqOmSHM8G9
0De+H1u6fb2teElclhCjlcJMMUiQlcR57adsGfAnz82E0y9kM0ulqtUm5zWcnbkT
/m3ZcAia37z879d4DP8w96mO6e5FL4+GoCM3HuXQ2QlJ9wPjEirRrCGgAHpWJJjC
6TUsIDPRepj7ldxY5nVSAvmJI+zhbDDGhndyM2tLyoLE2z1AzR4G43TcUI1yQZPG
EDj9330dS2ArNCtSqiWXnwlORgc3lMgWS7HmM4MNbJGY0ZORiw+qTciIiig5G99W
+iXIv30NmkTwtdT+CFdTY3H5j05bi3G57sT/Ds4wlclvlIuf4/ToeeAWszFEGcLo
MjgJf3CX5UA55wKUx4cuGplUY/Ffqq/8ot2YRGlTmjN4GRuw2kF4fgCtgD0U0Z2a
ayys+jEQSAKEJUm2XSpY6TrsPcqq2YpZCOUtm8bafCH2P1ayypPWxEPF4ae7ZZaD
DdULxkxSedbFtI4gM12/BfKUkpIfBjqAf31GrcFIDdvEynJLRMGw4YlP3Hn4WMEa
khB4Hp02C/2ibiCQ95NV8GDDw0iODbiEXy+HVrMgXI2Wi6S+bSHhl0ZyvKl75lsW
AxiZsvOjdFX7Fsvt7sStaLI87X7gv3kXCCzbIpfbCVCGwLCeGG8urAFfMrXSxUXA
D5v3UdFWx9fJe1Wl0aLVL3xukdh9XefDrlXzd3Ak0mwk9dVo2KXT3ciZNZmI6IrV
UwTABu0ujQwWTjCMSGK/c4fLQULgLLqsSfuQ0J2YZ/93ZlLDLFgvmIU0uaN7m4SD
M6aBuT1euWWTlHdi6oN1baF4K3RNljdU7ZOE+TCbi58Gjp+luz3e4PVp6Q7OUp17
g3QuoUsu4u1/BLGWPi4yMpi+UUrBMTkMrv9Y+HOunBNhcV1qd1Qo+wFGqhAJl5Y7
D3PFzOxUB6NPyqjXFq4iu70H5Y3jmiz5/mdMFpQtoAs7LNOPzg4UzRcLJPYv3bQS
w6O7qY7Kks0R+72xJl0FF5sUHkf7Pyarsi359iT2SRRao6QtMBYeZVxr24hGmmx5
eaF1zCMtWHBstcSW+tX+y6ExtZe+w7WibQtPS3aY/e7Isrz3hJ2z1oVc7Kq3M4ym
KxxHM9HytZHPuhcn9EXF3R3dH37T27nIACAZTMDRKGnMSCKaWMvBqDdeHT8z/188
JRJxTFOLA733j9bUTmCSW1xf7T/FgPcPu4UqdwxrORSWNIpDMqXEajDBo/EjCUWs
IxLOGAQlAlN5rEoCAaoK+2qAEAt/w/zLSL3ufURug+PjEm7KqTE8bArFtYbRe/rp
MrwW57Bwoo73AC8LLrNJtAuUEd/sGOdTJiVeGtLQ5Nb0yO7TDEay7AgN9cYrhxqa
cRaTZuh0DvlIIUqka92CskMEeBrWsM7PTdqqdniIAiJv4iqbxBzUuL4Yhkr9lMBy
p67TCxiZEnE8wBms+uAC3cK8W2Q+qsqLAoJA5TEYfzQAznxm1vr/gKRr6QzZMDlo
WL9XXfPawITmKHj6kzZvJJju8cfZH3zbKfrq7WL6xgUovnKupyNJU1wdT0Zw7PPK
YJSSwEsl3Oo8euv/rCFKueWUbMUbwCF1YPiqt/t+WXvaGo8xNlqPYtGtb5Lpjmjn
qAqgr+i2VrbVziDKDHK3fWnHKSbExrcbpf3qWq93EU5XXTU5SghPt0M1bCpAIj9e
kyv1EfY/5T/sPQr/1LffGOuNe+EkuF1LYwz3Xfzws+vEZAyPz64M1jnSs06bAEiF
HkyqU/N60hRKQW8wFkk3VoZK5Is2v/zGHz3wFn0DoQoMlfoz1Yk37Uk47ZC1OlfQ
Rvy2vm2ThH6qOXBgTzOLCMJUvjkHYzZJqpdkjbNDRSDUqox6w/PPILel6gFGjlgu
hPXNnJU0OFrg81ux/j0ferKRX71TfYt6fFqU5cYFNTiGzuvSzOmGGQI30ZhvoZAG
Et0Ok0gCn7fJ7O+aJlJBfhC1quSrW9VHvVKRoKil25RFUif9Qn0ZnInmUKGGfwdk
Kmi7frqkS0sYoEX2VaTjye+2L/GoczRGhhuE/xLooltj7htbO8Ae70ehcGS1AeNB
LPmLj5RpAEVFCveG2y6MrJBsXaMYI2nqrNGW3B5tliEUd2S/KNgkLpbM7A6JATch
E603iYiUjA2XZUAawMqpTVUFFjbkcxVDnZ8mL4rCJhZuq4t9d8w0Zdt2KxeJB0Du
l2fXy2fUvUITmu03ZyKCdNEouxPtlPLjn4diHpDgZl+rrwJ/hPURKOCAZ7O4gFt2
np8Sx6++RFUoGQ06QsNp7zMZOGH1kRybaxUg6segvBJnkO6QtdsZf3AHVTlenRmx
ifFEqiNFACFBJix/3rkzac5XLYZoE0YA1Q5CstC59DL6bgEwkS3Zz7TVyjIFGDzO
pbTeagmTzXzpJDEBSzMHNu+slgUb9DLlGhWiFQicpI7hxfL85s6cFQyhm6Xyyr2P
H1XiWg7pPNknyH9BNJ1rArdVFIJgzOGMTSw6s33ll8GnN8mQdH10M5tD6H0RK3m8
a6OoL077HL3tzucD0tHXK97lmJJ05p++UOy6XTMb+G/+2ZveWnvWdwVjnLt/z9Vp
Q42K/CeOYYf3FfXxz1eoDu7twwtVjGdDvWpj6M65EAJ7unufsgG/mYsrC+PwlTsh
dORZ/gU+RcWevMXJhSElGwNpvo0b6LOgvWF8rUIqKf/pfHZF9A46fsCyblQWsJcV
JHl03twRqakLlR9vwNzY3abjfxearnqvYTsnknkwJPePzbzAcD6yLaqQVZbaJ4v1
Qb9rermRzQ52tITGMAARjHOD2iX89Hzs7xnzENbFavbky3/AbLHa/iFJ8RJJw8O/
jEM1+34i+Wclr1f+z1N29CeNnELxniamQ4TOrs2POcCPrR+hW7dVcMY536fG7pzb
cQu2jgNC+GMGtOS1pC07r6WYyli4td5x71PhI6uohFaaod7eL6hULz81jB5M1LOQ
LGDHq6u1Xwy/J2mVF3AwPWZM/71+Xfjq0y3ZaNaXC8HPSbdRTqmPfFGbHwsKQ+MN
BSQmWKUfAkie2uh4K9GtsPXOD3zy8BhecKxsQ4kzZuTJlHflO/n6yQyL90t2wM54
5nzgZG7I3n+0DV+Jgbff4h+WNmgS1x6Jx6ze9lRAbYbKswN55mqRobD6lJsI1Hr9
IOv4pSwJfhqkNWR+juQNPqWjFb7itb+4wOlxBb3wqa8RBMMF2Nt123k6+VWdeA8D
ic+4hfzw9DXo7NT/VQ3Dk1Sdc+KVGtHWvLW4vj+AUj9jcDsQhdOSSewpH2eb6Ufo
hMmCmjVnd9jmU/pDAOWZtxDSyCX4fwq5rfNj2q7HQHmIm/6B6/6+tvA6UqEe/dfH
qDZ0UnhzFVT/tXXD2BODEQuXIU1qNmHUIEchv+S13aA1/xNDKyEt5W6UUa+xOIl2
ZsIhyaTZPM9IOhlzqhkzDkG6oo8t3YOa5NajTVuFyflS3Hj/QCsRRE7qW4Pn3iuD
gshK0TVWvT0FG+Ut1dJ4Tcg/U1h7fbb8Xhm+lRFrbIh89hCl4mWEU2s7enXM80+Y
i3bbG2ce+FZecF23HKxk+o81xfhmzS1LPDdo+R5U7Bhvsf3PHgSagnEjbx/ulM7P
5fqRSfhf1z4Hd6aTOy0L1RxJDnxQCQt5V5VLoExYHFAkP3FHs4IrxboYHE4gpi8N
er32Nkwa8fIPif8Vp2mX5Vk5LfQWx+fHa+zJxSoJo0emzh89HhunhrI0+CV8E32S
64171g8gXgu17kNXnYoF1GqPEF1rAMcTQ6+hN9ZkWtV/YIXziCSz6MzOwE8BOw7V
ZR84VH8PKQiD+bpLTPaS1gh23v6haErkvq54W6yG3iYXcnt4JvjcsuI/ZQ9whzS6
0T8t5SLwdnfIqf/tJDCJpxcFncQhxaQ5suYQg9VtqCFmCo4DftCbwS1T5lkdY+GY
LfJHch9LXLUV2i1389j77pjuVcBoJh3FYK1UaTCDi+seo4Y/ONF358iVd1vfiqaj
hwJ7oRsZWcnBUZL1CZ7zgDwTGzuoxYp/QSPk+B8Wct1WOxF0AvW5gH3hypZJlsay
o/1hyR9AOJj8xXuPUbwA1nf/6w0zcLlHw5LktCIn/vBRIPcBVrIE6x4v9qPsTRU4
H74uCcGeOGoXxzbUxD9CWpbcMGPxYURAqBxJYDRZJE7kCOt3G9RT0hf5yC5fv8OU
IbFMEFBu1LsBdaaomf8Xii32emNg3fWNn/NRDS/6mDc5XOZEdA7rQQKM8Zl1z97k
BJyxLCzhRP4i9Ot/ZP3ZYu65wTORYGIjPR3tHTeXrf5lxec/Vvxy/2SZwFvIv0i7
LIluNnzMmlyrprW7FbLROMUAw07tARvAd+n4J8AKnh7Du3PbvEhMMLBTuvVkP1qz
DLVzKcxxg0+TYYKsj2pbD872GzQr7E9jvMI5doi/DtWQ8fa9C41es8pyNeIueyVw
bCselUd1gKQkgVTVjd/nVFABMwre8ftyPdA/8coP2PhB48p7zvbxelH5JSGGOsPL
0hRzPZ4ZhiLC/8wyHhB/yhzuJ2mH6ScnQhjmD007rPpN7h8+zGcQzqRsJlJMLC9V
CEFDV7gY2NfIgx7HbauK0MLxOQmOTMF5tG4TpwH38iIwursHBeV2gL9TjgjlP2E7
g1mf5nL39V/x0MaqQOHy8kuuP1M8kflGfej0Iz9j5TEkFMZdHz9wf8VbJgq09Ox7
6YINDX/c3naaqmF5JrWTfN6jbRUX8X1fOCXQyDBMTJlXVlFf4b//LstfncPukVB1
hcAiOLM9fwHK8pbKax9JRTBYMWYByNgrefRGSQ6H77uTQKz86wz2PkDoeaFItUNB
SZKjAzImuA63k1Ha77rzY7S0DKh8M6YZaKwV35qCQCDvSFLEm2Jc12Hgl/W5FB6G
g8bxciHIsjNr6ZRy9BwyuI0jYNztGZncB9DSdTXkYZMs+FjdLNJ1xLNbsyEW+sh1
9YQ8loo3K+Qu209JOHvRK2NVCIfjq59enmgtsYByrY4iFphHvNYT2yrv4SESEJZb
lGIE0UQ8dwhX39DeGC4lYWOoIx6eD6j5Hh/IPQVvzmjsOtWL7g8rqN6IfvhwpSJw
+7GwDvn41WIu+i2/Gf/ECj5122MeYVXuT08WRIXdHbcgOQS1IIaHhjATJLFKxZcQ
LPgelgp+5LpeuKVtEjWG/jMLiXpoTkua5/bk/fQDOotOFtYe1cG0VQYyv2MEk2mF
mDXQx+FuKkUhgWCSHNcYm77QKTNHms7jinAtZkCPYTgnaD9CiQYNaoir8F7WQKo0
1PrAtzAt+2+ixhwgR03PCTyZBEHbbE0JeBA8K+EZVWxcvAZYTNi0lDTKgIFrbbiN
98FR0K46mOUfviv6v1nWYLzQYO77vYfpkNeAO9f6Hi7GL1NISR5HI/V8G6dNlr5/
r9qzPNtK0vYuaz1es5yww9WPr0w/9xV0uKKkCzJENRod1ZUqKalrnsFApV26oyoq
fONxcIRtQfYTbZurlV0HyGIUd9AMnR1DE7OXuSQEzSP7MxPYZGRs18UFyElbWPwW
WTApxWk30JYfOpuMdM6qzAoxkcDB3ujIKfoHgn/S4/dcUBkzgjOvKzaONzOVeL2U
Xr2HtjGtmweGwHMJSsexSgyUHKnRJctECl0g+WaIMppMoDtSUeLboQsBpvIsevdJ
G7w3tymG9Da4uDIRGAX4TdOWs0Wac1pSxvD4sL1Pc5czmEr8lZmR2hvieulpxafc
bhnYc9WMUNANhR27stl4R7arTdZAWDzy4St7Kv+w5azhgyT44EXM6IoGz+5Jy1mt
4TffrfWimxwZM/KKqULqasDjmroNLoLzCqbuxBPjR54C8iVUJLULlgU3BML5ej7H
JofQHAfHOsUPvHE991k4RQQMYCfVzGWD0O0jmiNsRhvh8lL2eCtUT0tW/JC7VJH6
6EeFTqmBIuCUkYkkG3d5Si/4Zp3xUqDITvEGqKr+Wq6QEACC6qQTuHpwJOHk6uIZ
T2gLomUGKBf0T+iKIvCZ3LbhurCNOcsD9RqQ94bSiV/fwR1dS2Ewoqy3my0R48Ir
kXGeoRXlvZEEiKqIG24EDMVJWXLl5E68bqkZ47AqZxBATMkYZHJ1edVVauxgLLVc
57Zz27S33Tls12szOqlLZhADmmWISxF3a9Yfc/bKABWi3eNBA/ZJWG1NCPlmMC9W
dd081V+kwKijso5PUqOLUnVzRbb6KWLcIO6WBne20A4q7aQMr826j9LZZ82z6EtI
+9gF0U4x1LK7c6VYN+vqsJmeAKNprxaPMrMt792JiB7wa9gnC4W/VPVVFr40DSRb
pl9My6LXcAMuWrSFqKeGRYNZxDbwF0cwg8JZb51hsulyx2wpqWf0LXbX24zw5nSU
2h71g7/WiSDOHAabxKPjVsAit307pENvldCoZOPZsbUQNjiuEKOSXnE1wdvF9gCT
cCU7mY+2zXQAnyTnYG4nzDOJRK1nel1+ytfEyIbEYnMEpu+xl1qZ5MufwXSEZqve
JkL+ptGzeBeTx9OyPQIh6ZBxhYkC4ljPICTvEpS8yzf9ZR+zyiDa1NvZ1b/Bxs36
chIsMpwSjydde8q6seYWJR2GMKshFJHrQiagVhS21QQuXxpoMGWNEaooOxiKkBWw
LaQvVUirHVBTAzofuZK1ck0At1hTnSuiBNT2PJl7J7LNLd7IBpLIPiJBOXNIciaM
KB7ksXd1QX3IwhoCvUnOc9Add5W3Qbya5NFJJwwQSfV0TsUjlYVT04xYsAe4Zo1E
mRIb7LOX9lL3b+QA05AJw1nqD49B+yi4xNAYseywGpvzfycUZ2YsM65XYZknkUZj
gbBm7NcKPJBZvqyZ7npihogK1uHtMF7lxY997Mx+hiTi/46XMJ6piIMXr0AUwBbj
+DB4NcQSzu3jRhWTbUOLxRyVJIOw2nw9gIj3zcJXkwnTGo7midexlBA8Qj6EnmF6
j1MLYHI7AdlISuqxLTYzikkYBhsRv92ELjSOuYkzx6U3UaC+N1tw7xJ+C6xI0aLe
JyGOZY8U5UjzPWGN0wmz1kmWQluLpCL2fOA1M6R7jvYedBdLEz+s8Se3J5PtonVM
St3bNUxCG4XJ6FVATytIxgCfDKZiF+/8IhZ1le0YDaYiHvU8muqJYSoVZki8U65e
yvtmhMrJQdfWQuiX0XLlHUo6mzDyzZmRqapWo4mXKCPKHjvvs6sz3ukBivlwIw9q
EQv2rKMggs3/n1iSxxgIyiY1B2FNJsKUmsQbOu8cAg8k0Fe0oY2Zqtcg4SSHXra9
s0L8hDzy8nnah+bDjXqT5SisBjsWTUim92eq7PCtk8P3OLLBh25bp+rODyXu5Lw8
F/IPKdLqWvaHZVE94EwNkNSZJ9qNi/C6qogqAgdoC4NTGR4T1crXlp4kWVmdvNCX
197g5usUUgQ6ulyaBU9fne1FXIPNXWY8BcOGI86biHqI/PWRRfl4QVUUVOrobreH
Qr7YhJYXp3is2enzLJH1v5aE+HBHzi/Ec+vLHgDGhf3Buuuthf2M9U5r7SnfEoO0
rBIMungdoUUxV44dkJAby2eCsRvkhgKV9RPEb/GGe4bu8RXzi8ALUz9UBarAHfmW
I4OOJhEASfTHvBrlCqbaop2dcvcZrYoufe3HYorj7hxqqCJL/VNDhSfTmGu+2jVu
qIgrQ5qSr1zih0u2WgiSGXpP3GJC6xpLQYUX4SQ3xQ8k4jiuDydz2vfOUNZ1g4ws
YENvZdzzJCBGde6yyk7/lnKvYszAFCcwmI/7mt6ppEXbNwMfFq9lImXEot5p1a7p
CNR5gryCGoseX+MeT8KEriblVPNkFyTIVKtEGJgVBNBPxraHKfDnC3qY09GF3I1Z
XAsXE6FFEld6x0Zn4KCHEi7JvmrHf5aVPgyHGp9bIgmZnV1TpoQN3U6pdk5KSjUL
7XaW+xoS32ewXiIHBnmW4Ei1/0JsIIL74Fx8lQBlNhuNu2gFZLyqLknh+Ti9KOyl
e1lCZA4bFXyUzk9uDfvfOoxiM2ZP4DWHIY72ruzFzOqo9o1FKcItAr9zIqnBOqLl
L82EuXEZ2z8Gp+XVzNGG4B22RjBE7PjY52z/r0z58ismNAvPqHIpGtK4NZ0PqI8G
seBLqh8LGdhbz7kyNANSVuZdRiFqjmr/aiMD0Kdk6JK6gIFxJRSAPT+gnv5EElET
m0p2vA2a+aS49LMUFd7JIB7p5iwChTNuboPvo1zEQtMcQF4ye0oEgjuWxy3BS6BA
aNzp1kSo+8NKV5RAwYxu5TyqwwkI2Lzshf7JW5qv5W13XVYoaDC7Q/Qmh9QoVDay
yOdzFTykkS9KYwXwfhZUN1YmeA8140oRaUhfR2CjIFPTwN0eHtsFymLAHiHYxHnB
heg88mXbKxE57HdJPqH3dusuW34Zodbv223aCn20+bFYsJKJPmegWV+CnhX0MM4Q
/U3P5vyYkIyGI1oe0QlAnwgsj+E89mMQRg1SPaMVGuy2oLZpXRrXQcbdxvRGYiWZ
W0oBI7myvIWtl8xtjGpXrrjkoE89hSOU67I0DHiizHyweqs4ff+yCyesEpCRdCM2
GZocIhCnzcAgIa/YnUwk7ijcCtTHovThFCr9wFd70KsnVCxR8SwsLXPtPm3YZK0O
wy7Flg5EsXeZqJZC4fPeDN/Kr6+4Y+4HMGS0k7udxqZg0fks+tMtG4/QqIOdS2B2
crCiHwJ+O6K+KsZRh4SKYdGtuxDZfULOTBGOO5431Jf33LwcXyGO2aEjUKaprZOI
7zgfeKOdbLMZPGzEhFv1XlpPRVd9uHbDVjIzj6shlxv+bTNHLwbY/KQ/jlS5U+bp
4YCw/qlvTjXF5uMdVlVVG9wcKr3PfXLUGLjrfdqr27KxtSitGMDbgmI/7l/hLbCw
ju+9s4vrJ4kTkL5hsiagbwmWrKuCWu7G/uSjujUtkubjhIPaTIzPkHc5z5pKeqXW
4soMTWGci5bobqZEP/dp14z8yHsjFcJd8F5pUJ2UT60jljAs4sUuj+C2Xx6Jy5Gs
xEviZc/qPHOXbS0HIZTvgswvSm9Cv2tNbu4S89ZxtxP7BdM0j1RgO82FiwMGHvPY
leEbn734iDeaj0p1AU/7PA7fvmvYUFx1cvItdfdaPiRSeWvnvGmYl623jusZsOcv
CT2J9bLs1ukeUgRG3nVB+sqwsfnmlwPpNgIqwrpR9U0YLi8pky1/0Wu9rgKG9aFm
XGhcAWnm9EFiCj0/BGUIJacTyu6DMK2XEXkTzwNR8Te8o177ONAi01bDndOaWUN5
IxL4TkwVh9X+6kENbquM5sz2kNbQ4r8N7Cm6Iq4SheN013a9oiV56dRDT+Bf0ubt
TNAKZP/0kd2J+4WWctcqV4Tme6SMXThLpiRK0j/Eoeg73iwJVV/kE2u+IzeugW/T
bz1a1kQYWoEeoJSS2Tmp/WtUbJAj31ZM2SmZyAgb7z115M1Gegj+OvsqdlWeXkbY
5glXtyzTMlGIQC+3oCuqA0dtn7yaHPOv3NzzWKBeTmSyr2z01/VhlWL8DQjYa7QT
Yy7o92nZgfrGJ1P/k5ROP8mHcvS2y/ABzAezjloGBVmW160CKBarmGnu2iDEf5qY
VQLt5Q2ZGjNOV5YcFpArntCyLAVDPTuV0dhng3Lbu2xIKjlPm/uBweWAMWzuPAE1
Qj2DjO1+FGckboilZrpsJf1fTaVExczhJdNICIZWJfh8GxV+ww2FQz6nXSgb7B1+
RcOrNVBX0EIRq/Ij5yVM3nBhRmHv6i2eVX0NYA4qyaSlXCFUM0BSb4FIndCcNY8v
x62hBHnhLYhPk5xT5gZi6WYxxDgcBwxXn2Jvta51axV6A9l93Mt9G1VJalW5MI8x
8MyCJz4VBhev/UTqTv5lLa380+JBST+SpV5ajMwrDSMZGJrXoZus7J6FSNhSS5EX
RFKVco81uh3+KnFjPXLrCKsyAsrJX87KNiNopdvLFarQUKnEsIZafxhe3i9Nj3i+
sntV0T6U/UtpHBTrNtqKzU2+syz9mnEj+NA872UW4JKWrLF/9eThPDhYP00nDcYG
EM9GdEyqhGfLBOC7WIFnMGxAwzvpYigRT2n+2U4VOF9PMoNuc+F6c0tLsh6H2Sj2
VWLsE2FzNLOdgQQqFLZA/tYcm6CiKbkZPGekk+teli2VxSFMbecJlyT+nnVjDYvA
ktc6asTQDjuW9nry8C0hk9Bh4XuUO0FH6pzfot+/Fb6UtkrSTfIpDUAUuLMzJc3A
uNPx6C2iO8oZU3DVW/SWAcV17lm78CJpP/kEfujcaWcBWD/K3MJ71RF7+WcJb3tH
EmqPWNF2+/LK/xluMGzetQlgXAmp6fzRiVan5Rg3gDdDCKakv3tbU+V2vG3DCcmi
rsCRzFoyY+r/vHBp1Qa6HfBfBVbQ5E2UADAj+zZny/a5cVSVYHOzVh9Js+TKhxg2
LD/lzQAtQz7W7VVnO0BOyZeaPnikx47agUNoLIlYQ3XXkex2Troi2OyVqe3160kj
0k1Uf2OlhlzoJxNP3z7Sq2tB3HvzRZCtLwtNMWaYUi8H7xNlrMHUpWm4j1+QutFR
kEi/Y00cITj4kgPtfDrgDeJhtHUlp546wtM9QI3DAi/2CZSFhX7PNpnZzOBh5fNK
liBHhy0OeR5Qbv6gld51VVMColN8hzNX0D3XoxZTIjsePFxp/Yuq97qzx9NiPQbD
GiyqNcpvmska6zH0S8SMtOt1U5OzR5S+x1+zjf55o7SJX2YX1ow2C5zOOfpF7sHZ
yhvIpECBtnU9GCPBjtYsZAO9I5w1a6PIqSBXRIC96v+MP6hb/gLRCZFXbDowftKL
jOOZdQ/KSXWfVJxCE5XIe7Swb1Kj1gbtSGHk7qWvHKITUPxbd4N4GKMHtgdPBfLb
ZZMiiLLH8UJfMwCXvIH0k8SqohNOIugugiC2b3csn1Atazr68q4g/56plmq+f9VM
MQam/FoY6lBDJtlPwiBwz1ZJ8AdWqtyCxewVMHk8sS0MKaDqtxrTqORHrWjyZ/b2
4eadkGO855VvZZE2ernO8Ybu6vhIvk54DOpx/IrmxQZskulpEYcF17Kk02Qlb0GW
yn7U+cMCPqtkAfU1gTPM/yyKIDcxpl1a38V1Tq7+No3YmPlcbhCivEn6w0f39RjO
whCOtynNRwpbkgqICxu1GgFq5xlmylEW86UhdDY8AthZMZLSeTXNLlrVcG9n+ugy
f3Ps1qS6be0z17In83X2Gzps0wTJdiqwxrwWolrzE5f0lNYv8AppnBc4+nYoDvgJ
e/PoGvKMUdgMkxUMwsjhBZg2KKCQu8j4HK6P3lmsgbsJkTRfZ1gi/Dw6GT3P37pg
r4RQvqccCsqCN5yXxHkfht38O8m00mlA700K7El8Lc3uiR5jW+CDpD9kWTMCwJmt
2yjPTGwtPNPOyzaHLsDUxZhf3FIroFjgZ0t9HA5uX+m093GvucZcrPNZHZRCIkrR
WHnfsYz8I+n3OkjJ9LNte827nAFDSkHyemO3MPepBCibOmuPxdpJUTatD+V4Unm9
GvS5tV96kwLi3rT1zfI6PSy6/F6XX+M0QHFhfa8q/bBIPEW+LP9XfsHqbWqG/9Pp
xbeZU51250AaWHOK0GGxDdZF2QIEIt8p7bydl/Ax2+wzY4wojpjzC/G9janeCUPl
mF8tFSNek89KJzM1ezxSuUM2HajKQ04NjJ2yegdTY1Rz5U9RL2pNe1gFU1pTUGN5
QQgUosMC+SNY7TY4aMwhy7F5h0bDYIV7j6/rsmqJ7GD2QYJjOpKLvTXpqsUtEQBH
ZYSBaS9/itlHvTK3ybckFGQIYb0VloD2uih/02nbPux56j0Ae+BO6QfHG3ftLGKp
r9JB37a+erMPgbPXG94B2Mfrv3I1+8pJUA1UuoUt3pasDI+XgaT9rw6tr1K2U+O2
1bzwqVi367hX/hhJPORVe2pewuD9aRsIzMAwBd28O+hKD9B19EF9vY2kuyPtRFIu
98ZS6BJAcwDcBV+tL6/ruDxIEozR+rtIdHizInO5/0919JB07FVRmJcjcF0BexS6
4/eH0ojLsNMEeM0o0foomogdMLNt/iYJZOjQ9+UHC5Gj30nBzFtk1A9MT1CUKVUx
8DClFHk4P+s+EcmfRMR9bUGqdhgwGlTVA5+r5GTIkMAPQ92HqBkw8/QbAP1fuNJh
mkZZ3kJCpP8W/YK/LHrZWcIMrPThz0evhlNM1mx3Fgcrpe+oGvQPGtDVRV7sBykX
ctJE1Rp3ney3phr9JFcd8RUDCkLraUrlVJHy0uyuE0YmMBDZeQVgxNm2KYgsAGZT
SpSB/NEGpvIv+gs2eJ9NGeQyDKB71wcOnVVdnF0Al1iloCZnTPs4Oh7xUB/k4R4V
II3kgTEc/KXvVDkFYIgcv7HetweRTJNpSIABlNDFMq3pkem0Fw9tVXzEqLLnjBco
kuWTCWhWO5Z/VmPocomUhP6fKja2Oq9vsr8ruwOXu7f+40inegGyfuD+f5/XCCUq
KNcJEsvX3kolB3LAiOjr7dy51deQ1UnxROoNt6mzx07N1+e52LyvtS8iYBXUWNWt
7zvN6luU6ac2+FIUEQ45kKvEXj6U3rIa0HpExrJKaVM/jBB0GKz0D1wgdHnNyTHL
Me7geo/0l93Z4R0esm4PiZCvEaB1XTgKGGdFyNlTZE2QoGmZhq74ufHBKOen72CV
8F6kpjrjlLQlpLK8DvMMYN7airN0EWBI8yXMPwg9qPYo04Ohdjq0KGm6IGJlIsYr
MIsdHnCgPp0n3wKTmaO6prR7zt1+L/oUvQmQG8bTYClnGChIL3qHVKcNO5xjqm2D
3ggkSRA+dGKWZtKLebfxSKHaFpMS56PM6GG1pcylJAkcr77fxbNo0a98xF2lkpp3
cse6d0hpUCv8MAtirsChsTvya61cBrbZaFsNnseuwEVA6gRc8xgi8QURgLcCByKG
/idaJTIWayUi2fF36zuAsSzzJZT9Ru883CMriQt5NWR7MUD6R7XeUUOGkMxKYHys
R55eYKI7B8yMWrqh8ahwWhXAddxkuXJI2aN30k+q/kLzpdPYAHeipw3MgrCWM/ka
uZpqJVOAeFp+XkdbNTvm9YTSKLI6dBaPuFhRYmxsCLv+scOPhHUChewSijKWXCYw
BbLdCgdvWjdHILjtYCK2suXgac247ooJXFE1BfZzmStqZ+SSO510TdbVqFDxH+1R
i9IrKJRA8AFAu+zBMwJLCG34CkOUaBumr6mdkybFozuentUKc/rtRi7fc9OF6lUI
ry6j893kTg+wWTJNvaCbw+sR2+L9xmp1bnDHRGTzPEgtzsWJmWxamYyrqnWVP47n
9G3AE+u8w52kkGf6B/QDxfsPyLyF1jVH+qKkCMQQgCiBFwUvR4GK5llxGp8dRcIm
9B9m4AKmJIWG+edSdit5bUtkrq7MDh6PZyZ90KW7lcxP64v7fGF6Q7muAWuFBePp
Qifh6HqEG53M1N1Mq7C00truKhjIaMGsg4ysdTQJIr0LwppkH5ZT5ptJIj+oJDGH
DvZpeaYQRmJLc9uIFppZsQhqBZVsD0IYvYI0DzqhABNj+ciMhtFkM1Ga+VkWd6TE
vfqCRNHhkVwCJzhu1LEr+aMKrHkvtHF/tfj02ue4XKvkOinLbzWkC6ROsIR4tTHt
BbFCVFhDSvQNEeUipg81me9rPjuA/J5030+csl3k52B5oGmP4i+XrP4HIPXee2Pg
WOqH4xkt7qi/I5X9r2aNPGcALd2dkhOo69D6a5NxCgVJWE/hKe075ITI8qQeueX6
viI7FbxBzld71eMYEpRBZscohu67077xTd+n9E6VwjtVrbOPhZWVKuKDus8MTBIV
4FzyZgi1mMv9glYWGs7IkqjLE79+fawYIgXLhJ2VpMp1n9eAH3V5T05RXUbGURZZ
HuEInhOiwPG5oNjktrxrMNFyuU8LUKQLgmzUynDSMG1qY+qLLTJxbXuiILsuuzMe
0IMiDooqjOqkoGAcbV4VyBEN7vDFAa0bQXI3Jy1MealnCXiX+nIRPUFEaZBr/RzU
tvEhNpyO3aQAsNulDTRLPTWePBBiaLEo5cH2TV0/kYh/ecv5Md+zHIihOphbnv6p
NVCXXUelu0IZmMOnsQRUmKAmTkhlYQMJYsGT9NiJ3ML0D3F0GkE/LrZX0F7VIzKi
WyBaoEUWAYgL9g5sj5BGHshAP6pHzYFZoZQawrVvv8S4UVTaVmHXXTmk2tfzGJwZ
PUQVg7DUFfMCrbZ1WvbsvWKXBrQr2iLqAfwMWX4hl6mkaz0OAxMkmT8T2tlFPTJ/
EM+AXbc7anOOE20Ti6x023A/DZg9bctv4Wr8nhElurCJtAwJp6zoUHoutThzoFZl
eg2XHs9ZDlxWq7FtgJ7qP+GXRKtYN3dwQplLSF5h5qgB79uvSH91oxoJJf7zmWNv
9A7869SjIdt5ZtwWs5JbLpzHchOF4C+FaRCj6AWigSR/QH+jug0HLXG+MsOXjhP0
5D0q/Ig1WTzI3wC4wOdZn9IQw6r3nDCvqhhn9kx361sHxAcXaMEHMhX8ORLpuA/z
fj+AC/pVdOREg3Wpbojs5REWkENu2G5w/eHHuR3D/njD8T6sN5e513z0q1e8OGeZ
IzbOTQjHnUx/70Tte6WMv+W4vB1CR0vHyEJ0x1qy02WJA3RdVnnQIP3UDKGKUwu6
UI2qA05H7fzpm+Yz5IvjOcn1dcw8I1S2ALoqfXU3YRUq6IMJ1nCTcrZ+QGUYBYc6
dmoVitd5YWlLfqjf4KCNVWYO7bzhpYPwgsaHIaZKXzw/dwjPfg50wJ8ZZuUWyVVM
GSToiJkm4iDzwx/sRQsX0zp2mooWKPz2VLZocUmY2PpupB/M0YEdpkod6UOE6WUE
4lg4RCvDmsWYuIpV2AqeiUcv0SUVSuFHoQX0nXoELfSN5OO+fv8VQsAUed8VrEI1
gcnvPLXhT1KH5kwSVIeHV1t2KQxWQwom90d7VdC9ZZScUpwzJioc5cJ/ISKev2k1
joKP/DRuB9O8H/V6ccmhEonoGNUQZLJWfvfnICZ9Sa95nbc6/QmfzqalDcDDPpPa
NrMmEwVUpOnZ72qf5IutCAOkjBCH810kPzUn5KeOlqtYLyWgsy+1G/7XujzZLee3
Wlh8BfejauyvYg8FmlaI4HQ5RrV6vn/puA1/MNUct1imiADt0OdmkwN3JczVEQ6Z
/AmbsZt080mYmyeEfIDeFtPZPhfN1981d62z7XCwC8894lwbkmG27uwYBo01NWM+
F/FA1wxXRKy2QRqqlY6762JbUiFhNONlBswtjpOCJnCYVn7S9dTnBfDlSIklyK8b
aTolJfj0B9yafTH7yG9vfJ/CDQcVDFtLbn+sD3SS0R0JCpt3ztWGXP/XgPECFMMm
lq0a0oKD19MOKRkJvrjch32XqWEAYO2H+Q7qTOMx46ZE9bDEYwQEan7Nd6wb4kU/
DjeZj2uRGzemxEhD/zT8msT9+UidMOx7oZ+6MEH2b9Toviutb3Bp261q+NyBbASV
kBwDrgssXt2NXFmq8XFnPe+aywkhEPkob0PC1FYJlr9hpyozUrHtWbIWjdgjxYdY
t9JgZe/pv756HAyCszT+oAjQKigDRBg1zvEmYNC/4mi07d8P+xACErhCGg0RKOzB
I2g88aLZm8DUaSDJ0rz2ToD+X4wtlnOYs/3nYjZAxRbtMm1NKKMkqrsB6NoriuoB
5Lj5HwhdDmtEK42lflJwPG1+0T6KSJPEIO1sGNPo8g5PDIcXa3lD0SRNNeOZ5gRN
iTr2iaVjrnnohH5HysxDSFRPGFUJCBB11uA4e0PQsYaeS4H5LbGdIvyy14p9vdIa
QkfhZtaoZbmwK3Q8yIxtnVRxz5eMjtgTtt7dRTpIXvhBJ/vWTQVn5XNuwYG2QEeY
dquQwrdsFlMTrBNb5fE6ppDFDCWwz0If5uPS68bay4p2lOjrYV4HmvhcIO6ZnzQs
EXpN0mUcBU7L/+ZOXOAVwicQTcVcPm8ZSog1Z/Pm+PIhTQxPosT9JBFYX+yqv6tf
4xi0cDA/+c1tF6J/+k9OCH+eA5d/vxBlG168KxMA4fzeM4hBXxOBZ1j9IQLZLDqh
MwwnlUPpkBujPjX1L6yrZQ7QxqCFTrwinetlREPeZF4PthiRVmMSMV4X+5Xl7pcr
N7f5FUbiK0BaJUWhpwTs2rNCn0ULlWa0L4nQgFpGOKGO5lJDXkYtdxITNsonmceW
b7vGYTVycfXfWWVlt09g30DenHT8DheQo2Rk61gJtxLpHc94O+HVuV6py5e6l/yT
gNhcgK5SVpxOr/ZXluNibl4aOR3YD2Qza1kJwgnirzvK9sASqgUxSCpZ3ufWSwzC
uXEiKsIjt3PK7QuTv8QDHGsGUktEf4on9Qe3BzmNiyUOtg5h/ba+ZwngBC2JIRpK
UZbzsHNzQNJVhBRWdgg6GswnbW3Hy5WuJPbxxSC+3bkxUEERQhTU2w/S5a6SLSSN
FxVl7UkDJeYCdk6M0HeUxvYAS5rvSC1TUHT+XfMDaZdooS754AJHbvAxeqqUGSCw
GbB8WaLI04tuSaolDeU1/EQ9pw05P/qfTD4GzGmI6gT/G7MW65uEYiml15acYqZB
0zejcko0hVxies3ap8IUZcZn/rWFSeM9+gRdAfPwgIAhXFYtEpjXlTFVcQifwI7+
h6wk7GrxIQPwAp01ZLmXyjvF6dyVIU0xwKA6hE6EJVVuABIEOz9TQorSDUqbasaq
lwckwb8GyPAAGcF5Pq7MwcVbCdRYw2SjVtxvvd2MfdoH6Vo0APl8QrKRQkPW4e1f
uZ19PB7bCOsFXjd93OuMH+z8X8buLLhrNb2O+K6QAirn+DE+zyYZcPmC+sMd5RVF
RZuRP7/WIc/zH5VZGYxT+FTOkfnqJjObg8ffrlOj6mVc0edPw54ZRwzZBtslEWyY
bK8FbowVyLieEuw18cRJSSugO+Q4UvAMKtOfIuEwCvkIGSS/ubhb+QZTrk96CbWh
yv5w0fakE1p7M7CvqTGUdUF7qz9rKyENQXxa8I9kZlat/qXRM1QKnk3JjJ83n3Mr
FxmLASWEZRFn8b1PPZqyRx0pX32rS95BpQ3gnwlvQX6lErjM5GIuaBB7OkHiTnm7
6Xa8dV+gJCHe0gMC8SK32z69mVS4jD6uWvo/2VbauIqSWCimBOU7Ti1RBsg3UpJe
P/sll2pG+5A2tKHZZdDnkdjUffdXY+eSdoabA8jILJaBhXw+AZ990gTZWbobZMPX
gCzIcHUejCg+0+HJR1yDS+ifgnFzR17KMvNXH4cSyleI9lTp+27AsXaug50nMqv+
HtO026Kz50+O72X+tPIgcXsfRagThW1tWU/ocMkQIxWurLaoniw4c91H2aOgDYM0
e1mgO0iT4sE3LdoMxeyUbI7I9y5wxWCrXIdOITcHW49oH7rziBDBo9MAwfCLbsvi
jYSIYieaz9e+j5prTWkIOx9nAU4of0saVjp7lr61NBTQDJyh2HM7f2aAvMQbGANo
4WBkm/32R6ZN0RUY7fRKwOYPpRwhKeeagtPGGmI2tLt3EhcyLYFPJFAAUFx/hHij
yIB2XhtJss3F8ErTpHYp2n17gBA0XucYmazvvybRUa5mbOnYKXvjGGCcjQ4wyj83
gW/uZDHuhzEbOaBbZGRJfDMKteA/NBLb0DeUlmvP+Wa0cv6yMA8N3MKnL12lS5NB
/1yW0GS86o7q9kbO8Z319a+ux7Q5gQn2zN2r3fx+99uid6GbvZEJuv2lbEI/EsiX
/ye/tPSyeIfdPELoz+V3knPk33LrP+ZhEpfWE9e0mH8POENzWaZTLlUbrPQcf531
udE7CcRwc7nE/wzRl7d4U86yJnJfkEU8jTsh6ktdPlI+sPpVVE/qcyxLp/rPlUgX
KAjS3PgapowZMkwhuhM1gxMKMHLMrqdqztnCzSRXGIzbPtDMu7w4E9w183TwJbxc
iU1ORhVWcheJVJvonqFxx5jd0uusws+htiPmTB+rVgXfy53CkJj0qqHQg0PMk9xV
jWtjdKvIBIv/r2m2cxNzy0WLWtzLsu/5826OP0a3EO7T+Sj12jJ5wejAoJarwybR
jqBrpnR/sL/0R1x6juoZznwH0p3X1cpjtMWZBuntEP7ZGbcIAFiy3T30UpAdgaVB
C3Wm99nLB6W1A0OxgYAkSSMM6B3CoB6YP0uhTJ6jHtZR4DQsJ3ZCv5a8E9tTo5H6
/ZUSwezj5u3yKeh853wZsn0UHk/MeuB+4IdygAuhXOSTIfjiP8SfgSnIFuog6HmQ
+x29cLawGDkTxPXqpcqhUH3Nxm0yiOr2TFHKdS59jYOGb3R2PTeKzx0NLI9w/plG
lefD8DA/Cbhy4iS28dlDjsy3hy7wHUtoDfTrxZcrGpDLsSDEOAzsvBNRZDNcaasG
23Hj8yxhZ9dQ+htgmid8TcCi2RCxlvILRq9yZ695dqRERYSPPtLYU3V6aHf02n9x
nCYcAmlcX3He0OzMVqSkAoLG6BOsHTFWweI5pc94nkjVi3UsGIMqhU1CxzoToOTk
HoATIqS3KOQiRqbZQeklCUK8cCEXmqnkuV42mB4Q7ZiZuLiafrq15j2IY0qZP8Mr
3EV89TSXwek2SznWCMDCRdYE5qSkWuri7UNieTNIQsqyF4SaoeLwcel8diEAcvYG
ag3p1cL6I0rcBDS60VjaiO6RWntzCJyuC2+fUKKblDFxH01g8w5Mf8IsNz/GBwoJ
ooLsRDcSTLC4dGOZnbGdMso8XX26ToBtm2K9NeK8gvj393gi/tN0ihr7X9eFP3A2
iHtM8nzCEn7PZ3gXkM/G2Z95YbQyBRIEVuaPpRSYrRRA/yGuyNk+vodMSAzGe8Yh
A6bGhWzXn8vNB6LlvMb7GcKFcSqikU0a0Q3pGckhBEc60jiPZINfbZBr9PsgXrW+
+dqCw3MMKZXIAve8h/pVSw0Qfn7TuTrBO3lpSnTfdW2klACsFX1EL5bFeptu6h+B
V1gZyVoqxyEj3CN+bTdHyM+3TRVmZn8yoNrt1f9tsJSTqxPFXNelw0jyEF/gYpI3
V7TENMbKdwTmzbtV7a7yWd/L2Pj3N0r64GEbKm29e+mBs6AHpdLQG3SCRoQRmLpF
XdlCTkOk0eEOoPstK/6OlLcPXTuROJuD5YX3v8g3o+P+Rk0UJCsnfCh9T6eQk/Fo
k+11ycu1mIFK7ykCnu+/imc8XEIejWteFRqs2GkfTHfZvo4pXV4APlmNMkY5imih
Y4jMElr4Msmzg+UsWsg6lYTob8pUyyhXlIpX7+nDiq6oQfd5TRVT+JhCwaqQ9PgJ
Wb44qhlejkWlPiDJmIElvy359yMC4z3yYq142m73lX1uRsvR9eLN58HwlxUfhUkF
+LOmekudM/4asZ0IUAhOsoAMzYkl+MONcSwQsn3M33B4fMSOQgp5vi3qbDLCsCgk
IwcIrnx97gmnVra3WiwCowLkj3Rex/33iI6NQ03AVphe/IeX/njHphzAtHTBCr5Q
mgy6eqhIgqAtqxfuEtJna9upnni1MiJQ3TLNiBCcZfhVD5cb6MGxJtMiTy52zQqw
8uXjB2k4mGcSrqrIrFu0sN7tjamOypH1Uom/1IwsvbZvc0Xw6ji/B6QQKyTP/7fB
ZQlwhbpQaUjI1GW0DgGJNcJbrRyHxbqO4M9ddHco0u5epCz7iQnIV6ldVcpKBSg5
VZDAqKLukJxlRR1ttRpelY76ZtCDPztIOY5t6TUpwnn+uNV3J3uO0MucOws+rBDT
1tnwTq+LtguLKtGDEIxUhemOuV62POSh78+9pFROivq13m5k2/buI+23iRucq5dl
pPuGppnTd9v1ddzNWTSP2UsQ+WA8udXZroUVg8/9mXOJZF86wWbmwfqcy8l0IN+2
/JkgudeYEt1GI+LZzfSbEE65d2PczXJJMltH6epXtPA6+nsHW7iGfv6vK0LuOq8Z
y6w+R+SfV9ksLqHcKyvud/ANe8ESpUnDMG0snTTSSsxWEfQDkqg7Vf1erFLb7Mt1
vaKayyNNujcEzfl09kdIKbqxDouarpFd3b8nAjj2a9/vkOSGCE8hteFmXbxSE9zw
cenflzMvQn+fCOcA+dg+RgO2pudd4ys3ADom+keySlF+z2TXfH0PeYBA6AvXAx50
p6pRg8UN2RGFBy2tNhT6tRzZNl2neP4ugbqqWy8yRTcMMTGGl0y9WtuiJ5k+bKcI
+3X+7pAMeE0ytuTEZfMctBieH/M8K8B9CS60Gy4gPyuOLuErkd4JRDXzHdziiv5Z
nBwoiLJ0JdGRZLvJCfgRi6yZMR8fo9ec8JTMvVcERZim9HpYRInoq9rixpHpmKCW
vIxVGQA1gOdYxedkl7HaTXt+IOIDFMtymlp4LY2WlWERqdA3OwmNOLDV1tokQPk3
KLW4Qho+eppBJrwJENoYofDc57Xg5Hl3o/b0rYfBQRGCqXAhHkAAbow+fNZKOuKM
CL8Pviczz5OFXPWfvIxVebVPkCOMerv+U1Aabebei718EjJ0Jm1Dfu5uXbWjEwSA
vXoDmx7PfdFr37nIoigZ7/Edq/ZbspcktyI/Bl4w2q2+fJzUklNiuUSoCqadIYqj
wplePKjpPdBaPZ/OBxdKgFq6L+FpRRAU7JfxsQ7za957WU1Qrl/3VTBWxCue3Oc/
oGgbg8zcqv2/dAsNiXDoiyZvOBpEIcZQk9x5Btz7IZz8MWQfgk4Sbp6+Gh0++Hpt
r6qBlkf/ruluuQtqHmT8PUpjh2tb0pAMXL4Ut0PfFegO8JAl/ZUNNP7LYdzVniCg
c+aMZ69MvOPUHnMWRbSeGzBS1UJolp26H9iYqdUFsjQAAa3czPK1ee9Eip2y+/Kl
rzs+ZMXTkvStFfiIJZCk0YnHFRMBUWedcX/lGxrNvNRfQxYR1DBRKLLfHwGinCsF
nhr9157kZmC3uueB3e14q8ttd9vRVtJUBnl22cII0sTiw7quXvD4pyeoY4m48VCC
Ig34tmRR2DIpUMX3khkAmWmg4az7z7BJ+LP1rg8s032aRwBFRbRZzHfXQa+eht8Y
vttHv1qdY/JcuhngjuL5kq7+KF7X+14NPaSaTuai6KHG+6g0xhbXqwVtOa0XPRCA
BmGzyDqYAG1sJ5fmwCopnoeCMwL3e82kd6SIf7LDRacKX1/Wk3J2Byb7W5oIaIP2
C1bZcaSrYva4ZvtO8KdHVsjPZr0bIIeHlK08HFc3bbFyRFula027WTZTmRH1v/cs
xxLqBJNhrQk+HY+cPKrUnbyoTYXt3EMMJR0SmBgQZFnKVDQ8W0fsB/a44nh75113
xNo9h0tGG8UhAVl3PbPJop0sMuUg/+37FyNhAWVUXisYwMncbzuwXktut0kphOUn
wLjmC/ic84Tf30621fSl+T9Ng3HKAaIR5A0EcUNxu17oaCIpafHob9XXxWVOTWyN
7sCsmAe74yZLVy9SSkc6C4LN8/Zfo+joyyuxhJQ/t1kDSXA+DGYEUnzWLC9Tf3xt
I3cDPsMr4KKJCBqD8wTsII6gt3t7dvTDtaBnVM/jVePc5x7hnHRTerNozc7Laodg
yfevFy3EtPVwFt+bNT7Mrqk7Ns1ZK6qM738jSlkX8ow/+9Heaud5sRcPTCmX7JU6
b/3ZCKBItu0UxtKGyfbU1QotUZ8G1rZLsqhnWKLh1MwUR0pPkH3t6S+Z4VrLwrVM
q3olb18pKnJIYsoD7ahlXRIkuAwEZbVDGu/pRYTLDxy0o5O1AsPv/szXPI4zuQcT
Q1f4ge08BOV3RrNLhH9buJcSCFYDYshYqSEsM+Ajqe+GBhh9Pf/75WPqyA5rdj8F
0oV1xE64E58ffMgg0EJlNzc8dB+honJbZer54qo9IRMqj91BtMG70XFpL0BoYgWw
6htKVsHsDAsnbchzUYAh8llNHF2fTQfbWHPFfWIyxMx151TsTa5NxkENTFw62y1N
4lSt4S420+pkG0cYUhJ8E9VZuYppnrquET1xorOdeXOQ+K6so07n/rL4Il1hUB5p
vixdaiOi1aqukVZf+rqndsL2OA0LcmVxkzi5ApVUCusvmXByHm2u9vsPgsoRtn89
fYj9j4yRIX7+LtuT7ZxndvjDpDMFqn5zUnmwLiLZEGbIFmdtDgfZ6CG83s6A5ZuN
/CXlB5DUmgRv4f6SSJ+s70FxLrOt7lFTsBhwREtofnbtq2dwcsJFzKOsr82USMwX
ASCMKvww8ILGjnYlWP+dFEIAon7pOfeWFCAjR1wVG82KCcpI4FuuugslMFNfMr3p
XPCNxzlnzu/HAsNOSdF0NCZaWZWZ8Xyod5lnk+LG3PUaAMm/eHE1iRRpKwGuMEMc
B7Wy3PPvQ+S06W2sk9kSkdV6GDzZuSFPaz581Q2uifjGEbP1PfgnpZ6le933YaTq
ioEB3UF8pS2SPz5EojZLviuATT/WCMFpY2EvfXrPXqbtgHJQiX0rHLGpi35rHktt
LoD8ivtKlyc0Wa6zu7G692RCSxNPn44aqQH4qTKJkZ9+Em4iqbR50AfIkx9T/MUq
RIOFeSudB8BTaise5nCz9d4xXDPkF3Z8DawEEGurDaArvo2Cu4d2do30VN7a8/gI
gyYKRvGasKTYwhEBzdHjqJQZII++UdRKahfq4MrOnPfEg2l5OjNZfuwEVQNkmePN
51vKMYe4/jwr1/7Z2YmklTRKmg7qOYGfIjcs4Ywc4s9vwbd0qKsr6WyaPuLYs0Lv
FZeZJANgqPkq+Usx8UMdqhSii3QnjjKOJloHpZ5LgmsL7XpLhhW4rXV1/Aa5e/by
WaNms+HQjo7xcDMx3d2SkhAJ03cKs+tzQ1O9tHvLn6fbOI3SnRFTMzl6lPredzxI
QUxbA6NTj1Mu5/5lJuNwIjHG1l3krymBZNnCIbbYj/g4VxtwvzPR3w7urIldShy/
n+VrUtekgWGoleFUWKfJtcYvyFnFxlqxHL+jvYIvXv+B8vpsbO4SfXfzs4sodVrN
p0CzYk008YGhZ8dWugFib3zfjEZ5occ7fi5KbxcGm9BaynNN2gUXaPNo/vgzQOmJ
egcvW3FTa0Bmjgi1Q/ALpfXiAaIdlaSnor3zi19xVApe9mXbTuhET5DsYUCv8adL
rOrsLYRnjQ5bZf730zrkkxtXJSKwGJ51gD8/7KuTLwGfpGBP4Ni1Dc/1U1+2WrOB
GccRLJWnVQJfn5lqjb+bLv694HZ8Jkm6MCKlgojMc58pVNVtOHQSYwVLr4KGxXzc
uWVvbLOpJ7zVHMS56h8CX/fA66VoV+Pri2wFxeh3hxN6dMg3pTpoH5yZgrMFz8UI
+FJ374DsAbprAjvippzOxAvFZylmknvSn6WtM/1XNxoRDXMR20wylO20ThYf4S3D
MSyKktgBoZVyVbAf8zwrIG8ESINI5iusDtx/bs1rSc+2dBYfc+3F5NfYavCTSTqA
qrxW9Cra9PTVSaRfOrDuo09r7gWmQuDr0u/HKsazKD///fHacUmM2Tvn39eg89YL
89RteyfsWzirR8eQa9XCYIx6OlbecZL3wLcAI6KtQL3exUXnz+iV6JvDlVFEupKg
caDrlk8jnmEkHpo2GMwaGYWfIkM+tU++SnbBvNNNQE417hCLXAcoUncxgouLUQ7C
x1G9UiFQVrUUrrhYHsgHM2/JS5kNyUwRzdvnG7uEyy7Z7vGAaLzdmKipS3GO6/fJ
bNYfW94hELVKhY7iDCnK4rLVCBzBQCnF1gDWYQgu6jvwDfnRTCBK3V9k01Rmysit
9/anM5mNn9I5ehf0m1VoRzZVqGbOTbvNBEI7vpLf4gki0A3eeTMnXPx2xqwA5zff
fYLxoKaXWkz8u9LfjpL0Ei2qC3OoyORt74cFPOhKWbUCf/IUOr8ghWURfaNQ1KhP
P2A2eGHbD/p2KT4fsMRWZx5cU0aszG418jWn30YSe1+YuPAfDVIkioYgRAXGWbc8
fFT86GHXcKz0SWzOU3e6Lk0Ox4EPn9JZhNiehCToUBA6oQlEmz5GycWTezcTTq0q
iz7tpQddx5+DDxRgBmJT6/l5Er47oCC3NTwHNeQsWQWUY46Scec1JNDinhuF3dZJ
ucVxPKB2h4x0WKTLMapNqSsTobTaCb+mx2EDKvOAXhTWXXTed9nvOs0qh2BYFPK1
HXPG1CxD27c/TdXOULZ+pRdWDMNkrT215oJRaxYfeUZ6b7NOwrxpAXKIGnIRmcrf
RCBoMk68SPe+QmLCGx6YjnEfADvwaH60QyDpcq22a7I+JLDJlnNK1Aq8i2bVftSq
NCTsBfik1rfjdGtoQuwyQbJtvVQspHtxAfzkDkOnX5WfnUa9BWStRiNh/VinUqS7
H0XmXEhdk2DrVU1BbIMhMcnYtb66776P966qaaM8C1A3MP/PN/jvVPpZjS0CLJ7s
AVqgsAHCMmQRx0lya8ssFihIqQBYX3Oxn5AMMn0p/fbwyBRPRiuyMGJy3O9BfejP
+oiWWcH3uBPC0yywlVO4HYI+wYbzK4LoZ0rCZGAExMTshPuTGCQv9/bjY8MgGG3R
Nr2E60SNXPBaGzXiBXpK20MaPsf7Q2vzmVLozCjpH/1rWH55jgVip/8FPkcM7Gns
nZ29GRWsNhtfKOR9j0AaHf+er0aQCW72RmDIrcOBsKyq1mS0KpxosMnFarTrsoe1
es4GGd4LFNReGr0aa8TM+z60Ekau2NrB0w2ihnigQxxTdNYKakSQ0tKxA9efBD5I
hs4MhGhpqblJndptKMSXhn+f3Ej0Bm+mqbfAvFoBy/rBEqCO+yneDSlZNxslq3NS
extKKccaZV3wEUC433rToERa9oPgwEYuf1AhvoAECZK1N549zpgpJVOI2z11l3AZ
nGct/xw+CzcSZ5PNqlOUz4ZcaLvrnOEMvmbTfiqs/ucCJhwP6Hp62GIKLLFz5SYi
KOY0V7N7ui7LCYiOVDa2CbSkmNSyZXAcTRtLcMPcI/dbw9AnzGqolsb/0pwSasuL
OFsm9c8GZohozQK4YZFcqeMjDMfu6kuIvTK+mcQsfuyjBb3lhFcVngld1d5i2myL
hyjOlMTXN1B9leoFmjWHh/BIiTQ/ZEmT1JkpIrfB9giX3k4tCEpO2J1IkP5aXO59
kw4/6lLjVvGdNrBKNwez8L5E0urrGQIwHnSq1IGDdN5GHQ7M2auvKf8E79qBTDhF
+L8+tH1rkzpu/7vVIAZpeHRl/zpRzQdAHdi7E6a2iXVys+KtQijaKerC942zKCk8
8n7p41L4Uhz6HLnW1qH8uR0sX6fuzZ1hkYGEDO5NhdZpMgK2HWkEf6MLXmXG2j9e
ibW1kYmmBkd3CHB8idzrOWSQU9BfmTnJMsGrCXbPoP/mQGQWk1G5vBUSIYazDI8J
yO5NdLLeRbiVa3u4IKrlyIXzu9NTAifq8Bng7smLbO7vPFSrqoA/q14Dka7hQR3Z
J32eEmtifAR5SjWI47TT5jqd2mit0LIE7GOsR8AOGIg1xK6vo/K46y+o89hzAY+A
t52t6qkvW4gWOBvljDd8LXlfkD/EwRAfOr3kDNlESI1jhrin4bvpTKXP1dSo1uzO
Dywj2dEpOMSs02n6rmENe1HVbY6N6SFn3IEiC5b6wtoZUD6T3Mpl0vmHqDG/x2Xf
kxIjswDPTShVWAoBeH0rAmzgA1jcuQoacWQs6AfGmjkVK7fj5NZXh58v8QToUJdh
I3p46NtoToJivB5zlpPDNSK9ZyFsoWOAyBZo5noc68lI0+VLH8kmGop030s7ZLdP
R/LK66cUdyKViuRDMGHRPlIurkU05EsYnbUMeZ0Cv97KBVlxC+tCbrZLLG5i3vlN
1aeWwbfQQ1TbiNPfZp8JmXcx8G108+RbRQ9qLYVhpLXgZpVpZroXKE5diDg+fLQ9
7TYo1t1fHmkzQhYI0W6uX2nCCDk68J0r2MsguyHSmybRla7rCmrrYCsiTjD6YIYY
DWXyweBFXCZUsQNyWdkwAFdiJVMpL/3kkjosR1v2jNz1+FY1NO+u/105JRAhwiVx
hG0lYktS+so2Uyv5o5gH3yCV6LoZ924jwT2EW3yz/Wr4ID20FP5lckDc+JHCA7iy
VuOqbgDcV67cYBBAw5QqoMeHQupAzwRo50hHftReZytgjTQEsyQ6QMuaxPJ/oNxp
nu34xF9drSJMUCQayZOBDJuDQSfsa1ceBpDFtHxMIBfau/Qx0m0w0ic6praSRMcQ
KfrPeYe2iHG+qY44BT7WPN7P5rXdiV/hR8kr0nn2BOPq1t7cXxlj1OhDmeHhPCpC
SBhclC3St/9Sq/fx0V45Ae139+jMUoXM/l1cJxq/dkWxV8wyv9gArTIGAx2mcogp
yoGnGyl5tnju40+RTjgXO2f0nxWRnv384acYBn5sd5BQJ6l6MrsqGsUwaJebLJd0
sh9aHFnXvSid19b4svg6PSLKR6cX+7L+bBHyZbC1EsnQIwL+gd3xVGWkFvCV+5lG
xHUg/swfH+y3C246TC2rgyDGlCgqT8Tg/MqSDFZJZ3DibQBt1w5z5BhdacGqjRL+
h2oi4pdITMCkMtW9ZIOxMsxdf7kJ3YZlg9yEszV3AGz9GJkSNYBMi25kuUnvmUav
qgiG5llUMri4V6CRjl7GOWVMLYRoLuljSlQZxtYQAUm5rfWn5feCedjhHPfbUa4+
x7iT8F6xKs4WnVdXmFxWsOGGETJKGL6lKQFjW0SCX966xu7KybdLuoxKS8UstT3N
7bHci1JzZnnAR4LrRjztTD9yKTsqlhFlyZNeLoKj0vk/7Z89LD7olSbe5w2bFLrL
kN9124btJ9qtJDKL4LGSleXUdIq91DpvZT+cpQx+K2Ak8/Lmu4Ix7u3DX3oRYONb
7WjlfHitu4yXOXBlLoMMR0o9IJjwuVIHiDwVvEQDWRne6U/xyBQWfCLqH7KQEBqg
ge+UmLT3Yo4+yUeQLS3xd1MsVSyTeI4UZ+TkalHpP16QULL+KKnaLmRHAl1XlwYY
hEgnAQtYd5EM7w+CBhRxQ2X2YY0PiWXkRN9gVFjXPpK8tirCo9wM5158kUp5TDEj
E8QTETHUFFfTSqGPtPjcZuOpuQe/1yWWHT/dn6+fp7Sgd+2xlRxSlOXTjs1TM/ZQ
RHz0tisR6H/5VCEIFs9EGCaCeJjJYrEsyK2fPUvJLjo0iDPhxhC+ixNFUhUINdIZ
RySxdcFzmRKRPBo6Ao8BqB7VlcDGGrqLafEPoOCU4kwDX4puNYW6XIsMgOOuDcSv
06YNMVt/GhykN+ptStGlTTSoLPI4nXIa0VTqK9d7y2t15CXPefx/cZkd2sBLaVcZ
4EmJrPRw+sVLHxCD88nfSaC+MJJQZL17UvWWAhr2DigfMjPB5YQW+FAdU6e+yVg5
7JV4fxYihzc4O4vumQumPPa1WDUkk4jvLkRyOg56W5O/MV1Oj2ogmOvNiGF348x4
ihlDdvPPgsyChsGxhm0tiXqVeQTPNVI/VTyWASHoMg2rrdvOerhTWR0jds+k0kxy
QJfiqtvSpNcJ+wyJeDAkQPqR21EQKg6l4v2hyf7P3qKl6QZJSnn/ON97sBF/71Bf
dxRVbz71ytPDaY6u437eC+5D4JXNvokxoM/ayEDn8Y2NrRrKxS43YNKQPiJBTlIr
qQueBxiw5UFsW+YfLgrMmiRhahDPdTfYGZJ6kZoOAG0mrB5dJ/5DvjHFcUJyxhrL
C5gzGblxtyVvxePYsfbceydc5HQ5pd+eH9DUCa2F8RVwmb7YoOC1KCLCc8k9BKui
DpUg57FwpyvjIdZGAcdWa3MqjtA7B0858bGZcFnvIpBwKySW7/aY+GkLwUkTzCkX
FHIiJWxya712SVkwI5XhHx1GSC5J4jm5k05isbloLEvulyHa10rXla7L0GTPTeJ3
GTWPIpZ4l9tMp8lHv6sOStxbsHA4xuvNlg355Y8t5hx65WZBGNZTTswszG7TpAzN
/VupATsX98MHgHsbJ3k2aQpzvtCO+KCPQ1Ih85+B3eT9Mmrs7dfoNnUfl+/nSNQq
aZG0IKKImzP+Zj3yaMZL5ycOuIk+EqVXL30a96t6HTV979SYViSmdLZmh2mUF0JW
MCBzaBwBaHfc5V/5edUkkmRUwPJhzc0GHh4dtOYSt0H0wAOqojfGIJYFto4G0jwA
NLXsGlpJkoepvIf9Wh4ehyer5w+d8ezoD5B2Zw7hoTP24m77RjfQwYptmu3E3Miq
SxWUxB4U8CTKP6ZGFAtQH9T5tJdX4JoXoZLnEdpmgaLLi9HRgxHCLCD8DX/330PB
Wc/YYNmWfHBGhU8CcTWEszTiTl4cBixWc/7mXBzYGD2dO58/neo3o2zcCIsa1GL2
Hx6w29KBNyJ9RdsEVUfBQb9HQKmGIa7BJ7yNbmrGP/hfWhbSgh17ntrMmRSy/q6P
HVdE307214GUYgTEeDxb1e/X5h6Jtj0iZH+ljuaZ5QGDCWVSBW+ZrFfkCvMw8a0j
YVptyi7j/9yZaeKCMlmwE8n/HQ9vnxor4Kk76LkV2qOzLeSapK8+O2rVLmtg/4H1
DYY6kAwp1w8VG1W0O/XE6cqTxtEB4SrMXaUWjQZQWWLXOrv3URS1ZjfTXmH/TpCy
GPiI65VIHE0LIpS3UhhbOE22q+TBVnXeW+pL7nxVv+WVCC7KXaOrXL8lxN8GV8CT
kmgULAnBXYvTIqEb30j5ahOjB7lqoyjpNZRvu6mtt6VgKjwuuvyzcp3J3X/+ubx8
rsvWYFNf82XIlQdB1muInV3sjAKTNO3fO9hDrNRjLKB5LTK3k4giZRYOpQnF5wax
8SIyXo0LgcTXbPceXYB1JGemlKRouAgM5UUIFXXO3kGs9d3YYWJ5mVX/cddp3f/w
/36lJMsEKL2H0F5Z2Mfii3ZlQedNiSD2+ebDRU1WsKdwp7qb5f1PiEdqdg7sHxvY
JNW5ym0M3H8vttZOufMRigOat+oKD6Ud218vRc/gTHol/raZYYKzRoCIvmNTh/WS
1RzXtrYXudk6uVn6fC2eyAOAjnSsZnwYpJ5xIUA2lQ89r4NRt8znX0dt7NLIPpcH
RA5i2mwvSrXqoEaNtxpEjf/235Lj61L04Eb2Ny90ydHixFJxesh43EKV7wdTV4HV
WCeYMxgyk1q4qQRqyPoEyk6+g5kUEHmcF1Ihp5ubgMICB1U28GTT9WoXimuRwkbh
PTHaUtDW4hVrvZVCydyC2X6AXGMWaVOyUdfZtxSH8IL616uLuD/sLZppuD6ajVuJ
eHVBurYOVop9924MvsEQDGj25LBtw4FMvqYvflSZ3HLixcLPouVWvowbMR+YprBk
TdmTFFsP5lB1nVkIKZB2czk+uDgt7eYl/8ly2FCpj9lu+eI6pn/MEPDbYovVUPLO
xz21RFksmvtRq2IH9s8UUjMgrt1OXwftAl3kAwvyDj9yqB6+pHRvjS40Z1MxrHkT
g8lqsBCWEJvkkTbAm0zEK3nyiZuKBd7li7Q/gMeP/bL3uIEgCdJ6F51BSvGPHyxq
mVAnoQL8TAxSXD6itgxB/jLt+/nWh/vfiRJ6MkHFeWK7vlQzKItlpR4KD/G427Zu
hyVC6vERjx+1rdjpu7C5C7uip25E54RxdAKDnLgAN+uGS/x/+8IDFFlYnuEhqY6s
PfFell3HQ5g0NKzqz9dA7r4rcN4quq40Y9vFr1nSrpC5V7/Rkk9CDUUr/yKFmaK1
kST1h0C3joZAg3v0IFoqZFTM/tuIiUVVaLELjVWOH5fc252uphrU+3ZT4xo3pjIb
GCuSiup/yNRGvhCAM0yYAqAjv3k583Niut8MyvDw9n6CJJISe3Ov59iU/nd6/l1c
3jxBHUGXbKVZuOFuLW1sVb2VpAiAZo2rxZ4ADQTabbF37CGppe4ZQC8nGs4Pvv2x
e3ds62mvP5jK4Fg1UDvbqYDwV0LjP6nA8cDYxW7J1NmQIUxLIfMJ8JxZfI+H1zlB
ZP3gGZNGUH6za5wubf1Rzu3HGB67qAPlFVUfYMyzJCC2auQvMFduJujX4nM7ABq/
m8ax6+a/LM6ejSvn2HEkFYZiG5uGsWC8Y0f85iKH6r4nwwXisJ77kXpM7aeLaoky
zNUPxiTW5BEPuG3hQ0/kkqZKOd74tAjUTLVyh4VjvjQaDbou68J2PxypISzJ5hGd
UCh7NzcuMDVyoOaBDjakGpusQhoYLyF1bZjkLwLw0EuGVz3/1FYMw1F1xYWOQJRD
eFjknmFdC02moE/w8FR2db/HLY7ViDuzj8jjbRlYQZg1JkT6TayzRUCFGnXOYDql
KQS4UI86ppejgnOQCt7jWKprPCepxTJJlcUpewVKLnqm0ovWMw9okHvijPQxm8dF
bR+4yAB8dmThbM3gHJGGT3dqyF/QfM3Vi5iJ1C1uI7VjYHnI93ZzskVv6NDV+ZWI
I9J49Xl2tZttoJopJOlc7JiEZQhvyiDDUuRtMrYhk5hqLOkeJx4J1LogcyEKqTfw
xs8QtwsEwlm9TITE31/XtYgl5jDljSx+44dZKGPKKP4xso3cYk5fYk3qx+FlW6yr
mI1S5VfbZ/mpP0hASEvpNoxyoLkEqFPEOEiIX43VD7kAhutuT9TaW5xv3TdBJp6H
7UTMFkLzjVCBw5w0oqlkAxWXCD4uuJiBo+NftASbEpkgKX7kAfn2D69Gv2ailLn3
MMmwCJdZhyt+o0FdIyqtZTlIIxuagDGkf9bs8UBo25fGivSDibRiUwytiXinTLde
VrZGA90Ez1EQUmiz6Xosd/sKldCflMoaaRkZ5EXVeRABNEzDZwATPFOh3ixCEWv/
wSGYB65nT/+M+pM9mo9N8rukzcSIXt7btyWxgwIDb98oPYniLvNhlT8NCnnAFJGp
KeFx8hidXe81TTBwms0VK8pfRSAv5EmKvBS69f0fFg5rNZKYIYqwWkN+jpqS6Vg9
CUsOQ7fFrloslHgkqZo41nr36+qua1lhHlv8jxo/FMs156DxNZtb0Ub6k7rZ1ryj
FuBGDeJpDIB+xiw+Hx8JJgbqnVrr3vJY4YpdKXVVvx/+zT1eviGV2IIQ85zuHsVs
V2y7zKRoB8i9BPEiSjy48CmwsK8MFBuVAScFsmtVJN9k5qI34uxhs0VoS6vDJyqP
Z6CBqJlMGR4W31aPTBZpJuUiuuEZGYUeDVfhPCbJdcpyjWJEdgbs4o+6RBK1Dyaf
Zf9dtEAAfdgAhmm0HJAy+FL2loh+eAvGjAY3ppcaUJ95C3wUk9Jq/gpe4LxNSSZY
35pjcCJSgjaZtxY0SSFZhnUa2NPrrH5/b4NXIbyPWVVG6QdJFT0jUO+Mv8ncjM8O
kBQeyC1wloXVAXrAnJv35K0Bk4kJRTWnQviuJM5kaQowIftlTVAEQ5ZSjqotvget
kelh2b0c0SSKLC79ISIlOSGsteswpJVhi1QOl+loIJ2qnYcvihpkjOG0gGk2FftP
w9OUVbQSy39oWCx6YOsiVEQlk0w7PC7iRyzSe1GUwfWtPon5U/KOXTNxGPPDwTEF
UsEbrcX2ZBIXB/r1hC2YT/g5dvInZtKuNkaUsnd81NdE1s7wi7oTKnoeW/BYB5Kb
4i9+X+QQLuJZEERrPf8GXNo8KkWGRHES9VRHlEHZZZthkDOsr7JhLvs7lsvgO4Zf
C5HTA5GGX+wGc8leARh9CG4rHgeMqqbSkNTICtxV06GvGs8SiMOyZ01xVRnt4wqO
Y0cGE8EMQLDvbJA1PwquDi+Db89QKeygleGEldJkhy7pbZuJpAeREjVoSXa7bE4z
AU3JQte8mzRbQZanmfHQR+kaAqXOx5hoxaOVcV1sUA9mra2kRsyg0T2oyk0nITWV
CR7MDvnA9A/WGflp37DsCvhEZLDZFSDe0RTBN2bKDstEaunh/DZd6Hcaso0dHD/Y
qjHEs2VQbELr7/Ixa3gVQZqTx26DRh2vTTXPxtcoFiRfj+ogpb6fRPD2eHBOSGO0
HJju6wJ+33R1JteOeKR8HCHbMpR76YsxnZtbHizbqW0kGKoYpWdGTjx+85nQWEJV
qHqjvjRLyhw09IzmxvmS/hSm1zYWOY97Ewmjqtd07mnJ75exZTMHm0O8yFRlxBGf
5z48zESeBLz8XeyMZ4KE+EKU+FuBdta2O2CZnSAJIbpJdSoFEu0Dvw3I3Y8eAN+y
IYVDe2KP0y9LXK/793Racj6Su7nCenAwuZ1kf6PdKj/Db11Of1u26ElCQEqREHaa
xFXSEWa1+9Cw4Vu2TWUUQdBkz8r2KlYSjobF1JhnYZ1PcQx3k1MNUX77gb+kxPWw
nU4uN4R5Yw5BEnQTybB4yZczz/BsmmJj/ySpJ37F06OLXDKoW6f5LhWLFzZmBbu2
hyUtAEWWRD5/ONWJq1e6/xLAouXX3+7PTkGume1DigJO5ixqCj77scKKCRy1Q09z
rpzkq4Wqv/VvoqbfJzOpV1RQKNDvnnlOscWgDDm3ruODgeJgg7xFwX/EOdfOMlio
/b0Akh/Zr2Vk8nqt+RqUf/FexOkFVl/nS7G52Ff2qX1F7KYe4dzuW2tZsv1bZlhm
EGx2LqyG4g/wHjWFebxLtN8JF3QC3h3unRQTy900eb+/PBh0x640ATm8+ehXVB10
8TdkOgctbS++ZtWyPDPVzPQt0FZv/8qW0QwB2H+gP3nXOBlxvKF7lJKiahMOrHlu
TdUNs9CsvIxSoeJIgbSKwLFcv2kliLuuts346IYeKPM3BctcgvDZ9+M1VMSfzIoB
ZOhdmZBOimG/xmCTWwQ19lHxmHXKpiVuQg3vvLAkGhJKR2c/afXacCklrBhLcGuy
3losuPfds5xxp0g8/cIBeYs96WHOZrj+59gClgDaycAqVdNcQywydsFMFHmKOpLO
w0NJiaf/O6e3GPJAZzFMvypsTnodx0B6sHVoPXjDeTvDEGYgKUpqlgJ+GZF7wTH/
B2gquWiWP+QRKPBkGBaLjz9tnPP+zWmTBxQAsJFjZrHYA//rz82KLFgXsU1IQ1uw
9Kf/X0M9LorVPgB/dlkc+y6BIQrODfbgwnkcpUtj+mkBPj5YtGnh5Bu39ImP1Q02
PQuLWTbqVCe1i29EfC0Cga9R5eTLOThR74TldoRm7OX2XC8CJH6pajGAsA5RgdvN
YMBS5VaApeJONt9igJx+5K23/taLXU3Z7AxpKGcTIF5mXT/3wYN9ULuRn3TsQGo3
MqcOTk/BEdKO8sv+hzEnq4TyD6E79yeyiHNsPsCgva5Ffwwo2p0emz7Q9d1WgxAr
b/a61PCJ9pKoDqAK3kXz6HZN/Fxj64JA2ud0VtrkPx3TRYV4APRZK/IHu2RNkp29
bWAjwEoRfO7QtLjSmKcD+YXKFMbp9TMXuIU618l1U52xfKaoQV9YCVBoPfYo06lm
beDflIiok6GOaELr46AvjAQ68qTYj1AygAUDbyOk+BXwn+wbV4G1DEYo5N7gIXnf
tdQ1ISFfvrB+oyckpxZxEmSnbV7jQwYF+cvmp/WYyo5xgpaTjy1bd1qZkLpVgGXU
xF0mFXvlCGsaLUVj4jIg+5NYwAKqnQ/RU1ROvNiecEMxJ+jLdiWZU8lEyKmwpQ7q
b03vD/b8848+Qn10Dgacfh4XpMSlTRuMkdT6U9LLVHhdZU7HxxQhFULa+V1rsN9i
vo83+ToLIthaMpAwcvIxYXsVxgdfkoWNkjhf7uTABfuNUagMwiG1VR81KseZQPXk
/BWhLa3ilAAgLJ+Nb83Qxz2ESoDk1kNjhL2UQHu4zHHr+ddSHpXaHn7C9E70kML6
+xeqFJOh6TxVVI5a7BtJ6uQupNPad1e02uZPh/7v7qfiJ6zws+GWo8gp8Cgu9prm
hUKzq1v1SAErlCCt5rEXkh6okAFCJ7HKj8HnxUGWHEBui+xI1hzSBCYcimqClevi
vMRQvYPS3UYGM6IWscqHbnFS6JCBJeEUta8CSS20K0DU+ZeBs9zqW4hNJuyn/i8S
nz7ivLh9pYWbUdkIrYn/ZiR2+w6WArv31BrJiNPhZY53jB8dumNiUU5kXRu31JBx
eGCn0eaY8IXD5xlUmAMYDk6dhraK+0U9cjy8WILNdX4LJilCKp47/QbZCHImgGzU
ZJUyKg734PJ4OUF09/l3iIpxNlV70YhCjh+DIQzZqZa0FVrFjnive4oNovxdtICH
0BnvgrhPsoLRK3ac/LwdcbxQvrYcuCB8zNOYnCLsvrKqBOHw117txYza1mpaLkxn
yTN/PTzao0zy7OMvbWr8L9hkA6tpQl3or144UVH59LO6W72wkcFhgY/OyAyGBuoN
CXMjwbiBcKApki6RcmfEkoVl3goU6iRCNgReig/IPmskxzQ/kJkkkAMgaRuGLA8N
AYNwCnltb/l+j/mqncOyJg63TZrq7qAAK6NT+M2PtE/tbt+v9s4UZrsjPIx3lQAc
dpmE6ad3phmulu9y7Sg36KzZHy+jpIHnnXWRYJO5rimAlQgZRj8rlaCMzIhZyG0e
bdRy/ObqO6w57gsPRwBWRJqMxzmUSQ2RDTsG+MIZlNsltLUI2gugkYd2MF9EgOGZ
oL0f/RBVIEikADrK3ayg+lsVFKEcfJ9UguRzpQhzTDqjsFbiYaV81ReOnICYLCI8
9VFM0VWtSKYk48ssU4cPFWdbHrZ9tx+3dxxI/va+uSlzP16B9NrgBkJ0GeLyPcVL
yVJZMS+b5bIFW2A+Uuqi1WGfotBdzWpKs4NHXNbty328PHOV7dWDqGf1XW3HJAgA
tLtt3zIt875yPL2r/1Ux3sx5iBjP0IiANoKsm7R2rPrDJiq14eahJHqgc6ZKWk6q
MlwUPtrw7zGZvwJO4GiF13GIGdBjbXFnkl6hp2/WxrAdW+SO2TXD3GxB14eR1gPr
8U8Ly7cIIgdhzUpV2VY4owVGs2mHNo0kJXfuVLxbW2z6ql1CQGE1RsBCJEELsmxi
QEPWLYcjoezECv/GP9LSZZ39tMcXVz40orPuMUpCNLwXME4L+2DTgvNoy0OXogtH
1D24qKpGfwdgxmJCDDye65hDdKs5UaX8pItsJ7M6RH5NnFtZbVlUzCJ09ECg7Xr2
0BAeJQrEehXqtgg+xRfxLpQ86CkBx/0tM4SZeTH6eOOzZx01/Sxv3tu6T/J8lDMw
rqJ2DYuxa67mCn8S28FoKqjkE8FznkVycq6wNR2QS1bd606FkvETzWHUjnqCxIb1
WYZtHsbMvppt7csolmVisG13BX6Eu3s1Lwa8wzykc1OjbDgtXsR52LTcLJG0VmjU
cUh0+RqbzZPsHnXSHc9Wm5a55t22iOdr2VQI9irLGvqEXPsA22eUIxtiIGh09wLT
bq9XDDRx8ffNA62t/ubWTtnj5B1Qw3rPf5fwNZ/X5TVDJ8W+u8jPJSn6sWbDi/Oq
F1GC0HV0J4IxRqvRtsK4EaXNmU40gZGUtb5jrZLaGPRVJskZEQNRa/U3IJ/hhSxu
4yS4XuTUJrElg09pMwosSYQE0rAehC3mQ2eallNB7U7CESWayEXluAoD74PnJkVd
hPWZPgOXhLsZkqJPXf2WTuz1cJ4CyG2NWcjC08wL0yglN8RzTWfsstuw1SQ3pSDr
yclaaWdJMj5pNpfaMa8T1yopLtaIJu5DuFoKYKECpbC41TMinX0DEQF/P1tsAnVT
9Jso84hc3Q8/H8kDQJjEOr3cUO9UqCpORIzVmdOIQ1tQaq7zaKKbK8FQsXGYxfbw
fx6OJIYwvoxuuKPlj29bXYlFLHJL/VHXzLbWSgVEtTmPTgvXuN6V87MV1a2RUePQ
2Z5iZAIizAoNKshrnLjq9ZvgAUbxLAcxFMbOkiNQFG9qPz98jdFAi1UpYLf1C+wt
Q+t0h46y/2FUdM+OqkSOrBiJxLF0402j6SmWB8ShqBEJcMKup15VNJ97kl6y5PS8
FYobweN3UXcINDvG3Qlq3slAwhFPID3Pfd8RwmF4Bf04tfDobPfcI4gWspFngjt7
cyMM+1G8avmhYLTJQAPaH19hLsAFfopmNhxjpBqDP8bntNSw1FTiUlSUEofweuKN
xiM+CIqBVzdNz0YIK2YqN3aAKiflZ9WCdSP8ejStJ7QP1rp+y3/044/jQURzo7pw
1gdr6OXYpIOAQStjGwEy7du/LhqOidKstOCvLZYb5ggrEuGJHkluBCjgRQmabhqe
g3hWTKVkG9nAEUb6ndRLDbdmfUXTOU0fIjVlqdWSEMbM2Vu6wL1X6+Gszq3l+Lh2
RL3R6NSxkq3RvFmHz7j+tb7pVNG+0o+WVmuOTpBXKYuUpik3+scrUAHPVft6AzGB
+y5dakU/lZtu4zQEi/YMBsvt4tMy5IvM8HdDqh/+0MjOce+jvoyxPnQAdfUVUWgM
3sFl2Yk0CiQQlsLv4ltPhBc339sEhr26Yd0rJ+zMRIjB/YtMgzGDN1nLmkcnR6lB
BIsoOcvbd4b144WHWNBR6IApO49aePDYzMddH8xj9aBvKihJ/n1at/kIDj33IjnB
cigPPrBVqldKGjQX+ccZa06tB7o5VlKcWnKLNE4SqVNctao6RF+8N2xZHcdFKMWj
RUwmmwPS7rrUit8mMSobWoxffC84lKL095jZcmlzXHp8zAFdeNBqdF4wQbcILqRa
2WSi+FIwXTQ79AFgDwHrxoarXkJss8g9RFozxcXJE8Z7ihA/zgf/gDg3KQ+J46aF
xCY7hGe+RjZJUivN0n5Wk7V06cMSwZeLgbOFlhbWp2VQ2CRayYEqVrWmfefEA73K
okmcOdxHfijAmzrrbJFjQapq3mJ9eeXb1JUfBet2e2UnSR0solr4fyyyadEnTr3L
VIwCkjh3X1/t1GjF8UFJrN777bdaXdRXA6tZ6Bb2uO9aPpd23gxgmpmqL8Fn6XcD
1i2EB/rixgfN41394CwYgagBRUAZG4oOqy7n7EXK9ErDLJgdbp2MImM+VBoKVCgC
W/7T38Ss77VXD+JAdaIOgCVJVsDHa/EXltrQCNvI4MakkxQSsylN+WnB9onMiDA1
jmeK34wdDkxWY8lsiIFqSkkXM+jreJsNL0KkmY7deOU6VR1JGuQyRM952hh+f3wl
7qGPpYZzwawbAF8DNzynf7SE3l5jgEnj/+nITbtZ1BKrTzM4xFfIuAeF2uhp5m0i
m+SWylcPoPldUcr0529rDbTmTq7T3Osin9YSNrzuNQTuqheYz9yL0Nykxh+pZ5Qf
p3lL4F2nc+ypAgXSdM2b4H/91EKQMH3m8JQ8AFnqNa/9yCRpc3zQVZIScj9cRD0n
O6r13oVLjX/zDyuSoMl0Il6V8JbMFQGYLKu6qvSAA54MLrBPexlEckUfg5r0z11c
OpLk+kKf8wc7hN1IbYANmPieeHeCgEksThJb8Thu8G0WN/MxamPjC+2L0aW1lbcK
OgjenXw65dmR22Qb0glVbyq8KqZYQsQcXp4ku+mEf6tD4rfKStYT8NtQNfJh4DKa
jNtrPOXbwOiRUTz8lSL/YAha7Ml5O4iFM3RlKbdMvw+gRLRRABx3mnvnFvPPwuLP
pAjetFfoPOgxSWy8Q6HHsOa9rFB63mQ+lVWimgoJp/FqafPLkvL2BumNLoztRrYr
QuxNlDVhRvcAC+PCUQPrd0HX0n1vxfJP/X2a8G9OAP4J6G7TNDO1F1nWUv9gVNEF
BslGz2S/M8KP5hg6+BVZFnRHoGWau9GHV90ibvV7JEdV3hqGNDGcN4kSYKcfilQx
dPTKcv6P7Io2WYuspHqo9Vi5VXNk1X7a4O7A17I94EOjeF1C4qam9EQDEuNNki0n
MyVNZpsaYWtZDDPOqmzyLR2hA2ZqT7/aFWPZKRib2LRoX9PrxkxhIsNTCfeuYsx9
pGhznlfsDATn6rA5hJjG0PYFViWD5tHmnV8oWaTtCEZFWdDZ36Fh0NnjmhhK2bou
sqLk6QGlUtquGRcRO5BNaG8kwAPOxZPwCtcgkvdtqge13PqWQxzOBMUjchV0R+3N
nNm3Q/yHtNUO4g5XXP45aCY7IlPIZ8ByxqXTV5tH2WmJ3ip1ZYvu0hTGVntmwFKn
T1aXk78cOGxgtRd8AA2cXjk2B96adZxPCTTQkx3rLMZ9KijbB7PwuyYIaRV9OSN8
q6IFNiw3qvZtGy8CTcFczXmYopB83on9yLHdWmpn544O3UxqgrHXhEpHqfEL/aLd
BcZ+JIkHrwbWZ3mLfq572QADbO0evtHzlGlWvaqSPETqqeFs+PRFutyxHV7Abxaa
1ketMZjJl76hx3VUJjY7+V3tEEmW9j49oYg3q/dBGIvNc2hokghdLDsP/NacI2dC
Brm5wBzEhZ7AXzrh/qobIaIQLKFv9h/r7NyklWLJWRznj7voagvbzsOWvVZlKIa7
YP5gAvWrUrbJu8cs7GvTr5w50q9GBGRgjfs8Lz9X6gJcoY8PT9EEOShRfiL1RmdZ
DiQrFyQyuJgxtY6Jd9MGtZKHRYsGMY1J3lDZ5Az0rpaOHNBGDVt6FlUOm/+1BSxp
EnD+q/7q4b1b9rzYHNz+6sOVF/NbxvCkgO18q/VKBilBldLHkuMhLJX8Y0+f6cev
M42VAra/zANyWtDdbazGj8BKhBy2nkYnNn432d5OYVR57TUhWSsf3XN1/qyUCw+W
1DOvn1oatFX3nvQxt1rYSHpa3+CKCY3OEOhmcNhnOXWMCuXRv7VrE0zxN32CmFpv
jzgH1OfUEQFLgK4hH7K2sd4zeer6yMxNqeUho8E1zm/+2f/LoRQz9HJRgE8lnww/
NcuqTHgLfWbGJamaOtmgcogzF9lxec6trcd8NMo1eyg6qYivyLNXOOyd7KZ2siRg
YoZ/yIpF5TmVe1IXEruKZavGoAVxMV2gFM2/aOsm1rNiNeoLeF+RNXrwxia+sgFY
IZtUFLGuZvGdZ+7z0ZUhfSIFrh6RdD0is7CECgkw3sYPJXtpFq90P2FSZhgE7OsS
Mp8A2ahSniTqsB2NiwqhHPJjcHZ9uiITcC5uRN7uKfLWpB/cGKoW+HV4OkML/caB
oVlCVxFzZEfxvaTKrwCFy6UYM8D9avQl7bpgRoEb+LdLNEDYjCqQ+580FRPVn/0D
JzWOM1rambi2CdEy7Th66zEZsjfn67noFj6NyESjT9NCJWpD/tOnXxGoNC/aDI/f
iCykKpJu3oHrVlhwoO4s4XngPeyNlY8DdwkvQhw7bAKhgWkND4ySbd01JFYcTboQ
JrddO/DA6NT/M6PRbkYns92wLiJXsSi/G2KYWfZcPA84uVCQ+FTfQ6fuZwq5nuP3
y/O1DPC97uMOo85uptVLbHI91AjD1bx6VJYBNoZJg4TVZcbKFThGG9TCuX1Z1XAy
Z+FRLqa3as2R4JUBpt/nd+f92gkV4oUVjN+n1e4V17J888pweKl0YFNYRYl8OH1z
Bk3JMm80zM22z2SrbZCqSMfqcnrYQ4OZ4qHbADszEIi2ytYLDCy0IP4AKr7YeZDE
eMnVIrWlkXZt99FbGucZbPVQbAN1Duzj3MBNPsIlGuiUqbT7foSq/RsaOn6XrXL0
UeREwK9dU6sismvHO1+UujOB5/vVhhBRHNzBgqgPWO14xyAYTPWxcwKdBpqRWeFX
txTTwYCfJYoWipXo0CPhij1xym4Qt+PH52DDuVtuPl766/a37+xfAy3pFvsDF4mE
K3NAmZIWMStiTwch4c+L9I1ViVRpB9u+tMRwD7ok4ZLvzqArQ7ZL9h83r/UASBYF
26ufcaQdEgN8Hui5NE+nzYUaAYc5jHZ+sJjO8rQBu8Zr1fcBO6WXboxfLEo3UMaN
yWCCD4G0E6zEUQRyOtK/noZuQrndjnQLzUOKH/P6s5dENnmeR/35+g8GU1LquRvl
Vs41vw1I9of1Mvs7wAb39iHLZ3pMuBoyfmaXN34SxmZWMuHOBsRGxGobitAB9dNX
0Ybf0VkuExIjZo/JDa3I99nVExAMYHtMiPU3jlmLMMukMbI21Eobx2gV2ls2dkqN
LTSBtII4GkayDUCd4RLxiSKN6uxWWFp5MNE+//bLfSL3g7WTxV6l0Wf1CksgxrBg
FKJF05LOya0M0GoUSFqaCVrwCrHe/72e6Ivn/isr1PyAh+UC5YbIhtoCsdY4VDLc
3XKgUjtsjASiIOd0DiGwf9Nj6qLcQHlfMo9fEQgdESWLOz9hB0ALRp9tubiqq0Rw
zeijI51vjyxrNy+srwX7A6gVqlAn9ghpA5aibTmGp6Ibl2kI3iRs5030RLXeRExF
RC8jV1Q2gj3iEyoXuOqVBkHJ+XBdLqcnOqC6Lf0QVLXGajLHYmL+9xL16PAHCoql
6engDFhTCvUg8fe4yMKkJhDlwS1uIvBtP+9WMDWSP4kCaVe6LZPnM5Sj7c9s1PvD
XFK+iZ9mEs4QHk+3pPBrhDCMMk+JsRespOolqvpRm4jzBr+bJeZ+M25Ei5JoJnUn
XiLFYWAslnJastxuAG0B/avlZpNKNVuyyJ8no1QJEr+cFXf5AO+r2+KFZ+Tv+j7+
IDoW384zZdqVp4Y0vd2c9jpiUdcAo0LwU8+g0qP3mm+vOpb3PCY5/wBhXnPmbM2h
S1WK5cr1pfTXH+dDF5WdNQejpwL977lAWRWeLikviDcITAq9ARlI8p/wx1970iL3
kf5qm9dwQJeUQihv/LlbAEIcxJHKyQDXTOY1LJlWneWd/p/Jj73TTz0Eq9LOB/1H
aBnMNEE2LJDGOGrzmjDhKxsBALx/vV8Vo7GkynWAGgzit0GXqIOqq2FWKJrqXZwT
/DJg2R3mQpyBp5zIJDBQDps6SPUi38Sk1MP9mHQdaerEQpmSyp2jTMCe/zbbZzXS
bZExmU2ZOvn8Nk8O/uYeW3mZxwq57+KmcxaqT1PBH6DBDjNiXuvm9iCR0StO0M8T
0+e4DoMrH80FnmbSQVQPIKE2h3LUX52HUztcKQqCViwQS0mqFyTChdMnP0PUFKGP
rnYjrcytSEJ9KJbjCFhB52XWGRXYICV6DU+a8+UADjoCYgFQcId5vJ2kL6/zFbMP
fLUW16GuFdSpDNFG3PDNQwskrDDJlQCj3lOEmw5WOg6lm0v0+jrVKR/vK8R7cQTV
qB0jJcG8vmfET1KTpjcS7gGAZMczRMnN6xEBM8EaznlD0qUT2rZOWs5lR5tVcMo3
nDJfrbkCORODipGtozLTqTVMlNxiaMDjnRZGUBaAEF+D+ygj7u0gSe/8KEewRRK5
yi0gPUrPSIeVjyo4ERgCdqQEBGduBRGJDsTlNFt5eDyqXuQlmTFMHaA9XoSgxD2a
fkhgA95ZNtR1ow5+JKOgCMHAjDMOEXxsDOvLVKbr5obmmYDtepDDaRIXEMSlI59W
ZRKcyhLnEYi30ZIlfwRMmFw+i70IisUMM8SUEKqbTjgR6kj1EZkG6gHjp0FcgAfh
5yoadxJx7zrUfxbc9guA/ZA+kOJp0Gc0zhvsgm5VAlGJjpJbF7RM5yaGuzWxEAh8
nAmsxei+R5PzQbblqq1vlnRyaTn9iCj9TwNyZ2QWa4WvyKBLg1RYtNNEPYERnl79
OH99ey3NkxVvFfqIisHbjKDLtLPsmaEdVleQxzr486QuJ1mGvDZhCn42Yp1a7JTV
D3D6YszdwfKT+A6sle7AjA7qxot11zGvSeUPqV12rFS+gyhJCtF0uhS2/CP3yrln
MmDhNzfIAkesXO+o7ZyzJMkNTUVrp8GNJaSkWzFlX9wINDldLTbXwTfCdN2bmxer
aUmqqou940bmQsyh6okdFxj7OSf1N7AhbE2WY7wNH3glsZVm2RbGV8b1/tieLuzz
EVS+RrcATFjEii+SNGX4Za2A2sFxYHydOvg8Id/YYDmAglZ7xlxN4i/zSf2LgGYD
Ks5Ck5Fq3d3+wdXHYrqdFNqA7Uz0zYhGuRncehoSRHVF48KZHQLNhJV9U2aQf9Bk
BSrpfbmnzxnG2dAagdhVA8kpkgNee19QStOCapgwUfKCZre9/NzBdHZ218ZUqQMZ
+pK2+Toe4atgwF1Jz6INqeBjsRRvJAsdkc442boo6zam9ZXLf/E/kdKSeGLxfeSD
orKPu4Yz7UCdwwTBZopdEeAJm1MFGCy0omLPXbRU6NUSM8x5cONktfp/gI7Kb/wS
43iK7NOM/yBLb5APOXc5WQTbwR3GKoV6CIfZbCzEXlTxUjwRmFEZeqH/6fBHAhLa
Ch/ZBaB4nmD5scvHtA3Su0wp/2gLhthf1iVhvEgIhqy7JwjPf0xgA0lcXcv8f5Af
lMDSCt8V+e0PylBfSCX/EpvkY7NCjQKxyT1+otW5tJzphoA0FtDneD6pXmk5Pc1O
1YT0S6CSXmZHjrie22dnuyfW4oGsrgYITOGUopQ20U2UTL3im7BjI+N/5bXtuCPW
ht5oprztyo7GIRUSYzsykw7LWSMUfOgeFsiC9F0fyuFZz65+jlZ5OvFU0NQn4q+a
MSklaHT9hLkJkXo/AwtUXU52xytpkvVLqbcXDihpb+hkyRx76geB4pn9+Z4079Df
B5R7yxTnWF8P/e5RA5UYUIIHxzinSYT4wxZJrr+J9Rvd9WsFp+qgcCRAF0/8I3i3
QLgwgA7DMB+u3EPXjR8x1MrkptXtwNQ9E8L256gTbYNqhy2jf2xuC7/0ucKLBGkJ
CTZ1sWz84l4vtZ5I3gotwXLHnyMbyVWrOHG5JIR79DXB5+JSKBtJEifZe/e5gx9U
qymnOw9c9jIH1wc0kLunzfRYmxMfKFVpIsm0scpesvyQtY5JDp15dqgY7V0oqVyU
mB0YzUInXSz6IkmJh0RofXI8C2tQysjokawFQ0MhBo3scrIpsV6Zyr1AkAws1adZ
sxYRmB+OjUkX03Nt5xr4fNC611lK9LeTAdTjp5lAavIy9YOyNUQvcELLZ78SBAZZ
5j5eUjDyUy93jrADHwLXrc7yrgh9hsZ5OYAMozrnf9NVEPWxlIpSE7VeChblLc6V
n9RrF/3GbJLjh/hSdhEIL8yLr+pavTlVXhbQYSFkb+of31XXjZnZRnFPONZJQrBc
U4vH8wfhaAYur+sCccYpdKS3sMYiSJOPAsPCBP+9EUPstRdr9t6t/mO1bh7oacRC
OkuujjDtcAfm9+9nsP98i5q4attMfNyusUNzafV8RVnw8tV9V16+Id0pi8djAPxs
SxhOCH9EsUVp3lJw8+Z2Kj6xFFz4HIP3IAFJ/41cug2xDbKtXr5pvbwX/KjYGj05
kwkuOZgDbkzxeW4qL3J5IqpaU/tXPR+AdpqDpcMb/T0NY97rUIgsNB+qx2+MsjRL
LYCQgWYQqruqfwy8/X/Q+XkvaUolrfvp2Rs/7IdUu+NRClSFAyC374yik0LKGQjv
Tup7SXC/VvZDxCyAVX6d/a9A4NGIsj3AyaE+U7q/RaZypJRjkP4SPrZCLPwxSK5m
+mvAdm0geS1Rc5zB/aafj3wv6oEOV8UrRZum2vBZeCgt6cO4chI6fDYAl9iY8hVe
dw+hQQhpnRuZjCsKNJ7UbcMRQSazR+jKc3gYBK4t7psc4gpktujXbHw03F0JjGdR
/DvUqCfNRPH+QBM8i0wHlCznGPESlLAeMfksPt41DwTNCtxq5kfFGWLtIpXA1+KJ
WeScXRWDnzTdGWNFj4jOZTGPnoPNJRGHOACALmc4WQ6pYzhdgGrU8Tb9+JVEQKaj
ESidP6pNscQwaoedkrnG6QnJfkWwQ2aBm3AdPOyYcoSGkez6YfdWlt06mBVDOGut
MJHAUnbMSVAz0QGsJ3XP83TodKv3C7BuM2awcRH55lCkl0ebhs5AwEgAOfZRQxfZ
xzO4gg8rVrS1q528kV3ytwtzopKQulXRg3GHlCn2nQLxXx7eUJGAJYAzry15uwk6
RdvXcw4yZIIJ5iGIpJ3k66ewjhYrLZUdEvtWnUUZLgxlH6YmmoI/1TADOA4NhZlc
IHckMjcf1Nj9fiFnhNPvIaarzjwIgPGvIUa0zPa99A8fqa7AZcRUBBkKPfmf01ax
sb06GX+JPCM4l2oHds8phmJFAVSDkpQCJoTlwClFFy3jDWR3LXlWQuE8yshM5RJw
sPV/eiHazQTwI8OBGUvjTbV0ezfYO+fCiE/acq0K6KjlIJfHCQlgpvRcAxbPEX/I
eIwZFUUbHzyCMqiLnhXOOwXAaIHelLw92Ef2HO3J4TjWPGpS5sDU0H8lyEzV1ozQ
pltqapDIwdptM7OnA+ctQzjiF0ORTjSRpdRndZ3ja7gpI0dGyMScjF5eTr9dhtrt
J9t4yMZ8+BZx1gS+Gesg8fpJtnC+RW//5ZbbQCYaJEm8isM2fA4ZsaTj4R2XJZi+
PABhYJbHMS6WzbRlj5JsHq7L8wJUvsEDmW2LzrG0DUPXzvsv7B/UHdmfTptvlACV
qXIRquI7C1PWSE85g/fSGr+qyLymnxW0EwKSWbe16MzbLklvug2Tt5ecGTxgfv2N
mKXy6wGhXeTQ2j/5tv4JPICMDNGsGrVPrFGoLhHj9GMrFPM59XkpNcCSH3IwMOdg
geFfK/tZVKK+J6naKTV9UYlMED1JOpo6LA+mtq88CvtjDrdrS0I2jZ0GBu8BDLPG
x+ko/AUk+fNgZk6bl8FFA44BvdGamWL+/U7baWvA0mv2YpJEhXF3imp/og9pEEh/
i+BiVcxf0G7RtTT6iHLmN+H/A8usAD5SssJ6mQFM1+Tme0QBmTU3o0fT5bJmEWna
vB8Rr8OMPV8+KMsg6pJ4fOEavCzEjn6oD6XcetYB1Y/1dPJQu80N+oXMtAQu3kt0
iGVeuUQSDkgKoOEtmK9nthy1+CxUrwdx8Cw+4+fTB4aTZIzq872NNLtqXoD4dj+z
Qb2qclHls25GN3Wj8/hIfm4A9wQW+2XwvmOqNEeuVEQJX05+Y5+79GsMDV+TzCvg
moARMJljv+etcavJoDjEmKC8thGr8vqhRJ5vfbIqxLpaeFiYZReN37yW0CWjMTvK
N8xLRzVpm/ipJIVa6MDHqZgk0BQL3tRH9YgSdT+FuD02RuzkjF44JwygrMzZXRTy
wb94SFlp6JyLGQTNT+nlU33h80QzEp8E7njBWj6l7bg26GOgcGnrF+wp8WXoFmc8
8EL2AfZfVyOPcPPGJO7lzuxT4X1VfE2oGIhmNo9x9bfzgvoK1d9RneJpdsa/ODtR
rhG91kjrnkee0/i1VCc70lmwAFlLYtIvrFCbl7+eJlft6c9O6Ubv8CiUDB76/3Ra
M2vto76oKsPmKRsybucKmGhMoVGsDG8tl0imuyXgImCvMHWdI5UPLpMjqVDhYY8j
a6C6teOl6iv+9+A2PGuuMBNPpuqNAZ/216qsK6/Y5WLGYz6cYrkeu9LHmZXu4PV8
A4pbtzOozgT4nkg4LRbkX7v32rcqmNQhnlJzSW0cbGRHEx7irHblo8+0kCL//r3h
cUPJ7gxKZJDSQqIiF9JaMGEPEkvSUzNQ33X8EqBotQ0yPgcDW0GtOSSTBdiLTJY7
6XUOTbGQM4zhkmBysXzIxcxxBdho+aRG5za/dl5kbOKwXmFFdemAf6ouXaNrlbGB
hKALV6NPG3zYUgRrpRfHuuDOFSM35q2pLEXJjwbmh6qg0PzDJ2DLqIQGYfFwSyOn
0eenYP4jMRh7opCOPJ6H1Ry+k3yREskAielIUUAPB0KEwI6TsdcsNiY6XyudDJ3j
JAP5nDvJZUVf4yxIBb8xa/wk4sJ7ccdQIv/aDuyq1dlvU2iPeE5skzQBvBtLCUR0
7uoKhoDR0+3OIYGBjh2/EamQjaBYIct43nPX+kUBTMg3JjqijWZCtrTh0HdejvOR
9Ida/kOjB6ybiUW4hvxXOew3PGlzT3qg7MtCOhnMWf8bQtWX5ddQ+0Q8mb7XifZn
0K0Svxt9NE2QS9K2o4pqkJzbL39cFmSJOcaXnBRDwbqqH60F7ZzWVHUmUZJk65h8
SR0zD6gtd/g7mvavfVdcj/6Sjhia2F/T40nePsma/QyRy5Ia+0dj8ga6HLMvpN9x
DP0NdYh34DrQVICpuYAtwAswWEuo7pEdXbQHWhQbF2ieS/Th49UJxTZ80IlUPdc+
bQsvNcarBC66CnYgMC5sDIqET402QKFVLzEzipo2ZU5WZ8j5fXLOPxRtFyJnVOrr
XS9lFJXBfwCqEGJacfQcRYI8LHUDeFfHMsQJPyKsOwe8a49/nh7zL1pgCZGP8y80
dZKZPyIbkxHajXXv+xDaRq73GvUm9imeH0GqIkRwBSaibhbCalMRhkgZnBBQwKDc
z/UB1/r55qGKEJ8fnBDaKKWzuaYJ8TDa6DBP04fviS2Gmo9GZcq7P11glwcfvs1q
7nFTPI1gvWk5fdRxVX8y6sy8Zo0qUHQRg/R7xXeBr60JCM4Ihcc52HL3zKkpO8N4
/n6+vV/incsLkdj0Cgcbhp1GHG+pKpbNMT5rn295VP0TaqQ1T6/XvfYrRbWmUf0f
qxyx+JhZBA0vbNwEn8npILbb6CPzFVRicM2nD1xC1xmXCA0S1AbFuyc1unNnxVt7
QolE+lhwrC7EQXyQ7KFkbNsO4UwNW6DHttd4aDVD+HIuJ3/Uf2V7pUTK3HOYXAX8
5eqaKELSXkyXv1KFKrWqPajBUhg6jnbPNichm6+wk2VOE2ssOUq070QbJT/nm9+n
vzi+bLLIn6BXPVUEjvdkHpoPKkTj5xOLEE/kvsG/LSbrQT+Dqy8JXTuAG7UdmUKU
OJzVQtFrXj+SOBpzVfed6Wi/7GpvrvVa8kvLm14iGMxdTzj0oD3yBeS3CeFPAKf4
RoB2960KaWFqhK7eUsBxB7YMeMyLTR8H5YvfIeQVMtbrgfkfVFjtugUdP7MgF2Dk
+HAi7//zhHRG+umpFG9PznM1ga12PLCci/Ki6gWVKuvr6MJpdzsCzDnfhYeSyY3s
jV+6ARoWq/eLQN/2H5nIL+Zj40KcIaV0TvNY+oVMLxrdu0xQKXvp55eQM+XVRbvg
ZEHLRZm8Uong4UiHWjY0Vmq6/oSnYyUXDFpx/kMAQl3EeV/EwE2oBB/nxDUEm5B0
tPgxFyaZaR2m2y0gHZeF7XBYetMhE8XQut9478bgTveRfsiDjLgMsvCXp2yyfaph
w/IgGXJEC9E4sijSbFdug2UGWSFPva9hVRifR9sB31GOMM5+3PScOZ9Sgw9WBbLl
5wmRQUdXotxKQcwoGnUhwxjjivBfP9pZNkxA2fScsOZwl48lk/GULM707OU2wHDk
dOW+5efV1MTzZVfw7YKDPwVk1O68HvzhmTrHsNwF4dUdovkQWQ1BbmWHSQMYq6qD
NQt2JyPPri/8neEbCPoqpILfRUJnR4Hj2DaX4w2GvvQKNHsA1eK0iYszCMHwwPwU
ENzQfKymqEDVk8V4RmViqb0tGOZGGMIMPHRX+BNIFe6MKM8RrgKFCH3d6LRSSprm
BHH8EAc/V1pW5Duk8DTwdz9nBfEvtbwvGeLvVzhDNWEMwW9MNY1rbMRkh1Ezgel1
V9S8mMW6ykm/J/BeCFUJQoYozWVstDeQ+Zooa5vf5/lAidRHebZtiUc5o+JfxLyf
Ug8MBEiO8IlKkyptfQfXEc+ctfIS0NXjBxnKMYhQuxwoAMNfVG8Wk/68D/dYcnIy
GlsOu1jyTCHE0N39+i9/lhoS1zp7j/UhqpuSE9ab9GKOMCLGs6p0SpAL0ZdrR9lC
QJEMNjvSaR26vNFjqEdGjfOlKXMwHnBMNpUxM3QAeSr1uMmwwQzty58YVDf9lQ8Y
mnuY4iorDLNeP1xMm7eqZkiWjMTWTZZCemm7/ngWEi94PEkRHn3Lbc5tjv9DvOuY
XFotWcQezXHqQCcPpKD4FWVIE4FwsHrOv9UWDhvBvx2f0uUCBwM9ZP6T/opcu+uc
IEGKtOqJmUtZ0DF1zp/Zx88jOwpRV2DV2i8cSs7Pa1UvMVPm6PkOpWGKpPMhblO+
LDo3m1JOpMjLzETuhO+1OxsFhex/xr/X/E8rOZ5loKH7ee09x6MuayeSh1SAnjgj
JDnh+bQKJ7K5j/q9PrBIxzrf3uaunlzz7uLh1NYRpeoKL7zm9QclPNARpG3lKmeH
Wq6IRBKZis3wFrQVbHBXatuY+zLomdDswnXiY7HRHKgVRClRNsYfTSe9GEO4f1+7
hARMY/x9AsYP+UoBuIkzYs3CXZ/Fbkh0+N6+1Nc4ocq7pKZ3bokw3D5SdrNJ3SjV
uBTAbnBvKdSKZYpVj06E+o0wCJZtwF7vFtInJZDxUd4Y9WDO/IOXV4GjplwMENN7
+VJ/rbwZC9Nh+hOxhMd5MdXqqqI5vWznzpZzAqLoOaWF3U88z6xaLdL6D/KA6d1Z
DVkJUQzPgeyeo2Ko9QmAjCstHTkzoC3PRl8icvc11wANX7c/Hul7XB7gwFw9ArLi
D9noz7EHqj0w7IoN3ijv7c8xooukRxr+wtVdyMXRSB2kyv9M3p6imyuvoo5tIQLl
xzKUBfXzkVtfBFE1B2c85LwZkoDWfOvcYQ8zbLRWUg8IcbxnSE6cxgRze2nP5Cxx
syUAJ0+PGY0ozSPujbsQfOyRlERmM22Levzx0tt5LCNXFasovQvNX3ORuDswk5S7
OYQUJRgYx/HxAg5sGnf/JzzI/uDk9qiLHbs1+DRLm1ukM5BFfNK5huI70bUqRj/5
srtIrfOkehnLh9VVYJc/lLGoFKNBtgNoMHmf3XUozoHpA9946AWvrN2tfTz/F0n4
OwNn425r6PGqjdMnTqw3UAlIbfNa8fljK3Wv4uxqVR5+jSpctPQ9pMe5kLUpO8Au
gU86uxeXwA14goKcDAeufNi8w+DPDK7RRRyA5as3ziHcVIAVm52QddvTIsjYetds
CJbeJ/Kk48m/QCoKMZqHkYKWls5+eXVX2O61uH9/dao2RaloBhjpKrWtduJQE8xx
sEYjOhqjuvPZQ2jcy3SbGZUsvJ5nkL46J6jI6USS3ZhJcg4c6nZQ+JGn6Z4GQrUg
pqJWGnqyfCpNJfbhdnV2dv1kRgML7YTFw/pKjCyj+FpFTfyxUOXF9YJE7gbnGdSW
NtYjQPmtK5mGMUpk+XaXEGTB+3jugSds4/V5I/V9EeI4dcTiL2Rb5aN6CyNMBH+b
7c++wNka6K/++cH2b/20itjsvxfZNINho1GC/ANU8g6vstvbi57Gy7Zq+kyxP2BU
Jy6Smb/KdsFSyl8OgfChtbFMKTetquN3AI7+GnRQfcnOPFyn8Fd/aEUxZPy7FVbb
mexQV3lDO/uqU+ZlwepcgjASgfzmoZwaXDNA9OkR17keSRp1UEMJXmy1I/nHBu14
lOOLxX2Kz0HS082eagpjUyIqfPbJVqI+HnZPWfx9/hOPVArEwt0V+dMXCTmG0w4G
ktH/JGrkiGjT5Pi2NLUi0giqFAOHA81nBN3on1S8V/tv/0CE7D92YEKtzEpWHrVI
QXZR2tG0TlS+ByHSj9geAUx76St3mviS6NVabTGJGgKBuqcQhlH21LomthEicv0z
hRbQ1LiOOohaJGAEZjOxo/3QNrM/K5fG7Pnh0ACr7eZpKBo1fDAfA8jmjHTcgGxE
RNtd8VV9lhMmqnrG4/gMPwEez5NWUEwL6jYObPDIOlZHirr5z6Xtjbm0k9Rc96l5
yWa6zDZaIRZrEZLthoMeKn5n2OyB8m3EsHVI5KBzYpk33FdWdIN0kHzDAXuntZGd
406hNSMFcJbwIHrZG5dDFvOXT7k5KCs/j0COL/cDtq/6tckv1xKSpYRLaqndiYLR
+8kTZFqPr3sBHx/0/8ajCTrswsIMUcJz0N+v4d/O5l+tSpDEW789XGk+IBHQ0lgF
BJiHccejj6mLFF7Jmw2ZkZ+VkGbZjlWirJn0/DB9VWuLibvo4cUwKUwWqB2SBd+d
ENg0MzGhwL/796THYsfIN6g3e6nCpUTN/3yxx1DQWHU93KfnByE/J9d2HyEBjlGx
Q7F4VeEog5iLk1/qdPJFNj11jH23WFDpho3gCSG2OcyQ40xXe19KmXDddZtkXDc2
X6eMZAGA9j76bVD/lXETVyY7MowBJlGkKps90ztwGdykkE4nFesKFsInKwUC+NwX
uegM4/KjOWeZlRZA8mV3iKrEcykJA+hw6uYf7xRK92fX4g+vH7DjdpQ3ZnzqtXlk
KZhpyPNgbB8fO3cR4mg4n8JQDhyF3rTR8pQRVZKezhOEbwEepTkUQTnqxyP0gCKw
ddNhVfWHYMX5pqjLlMkVHgHOg1VhGv/cJ1h3W7hRg01/08FF9mr0lfYbjEV+msR8
hfAKUke6BZlfPsMDkuY+UwHsyNMZYYGyvClhxlWxZU2aywQ9oib3lKmUNAJ2UAH0
Da3w1VlMi2+EW06AK8jvJbc8da+0gl5p3E0Ec0JskiN8ZPgoL287sTJNc+mLscLB
H2k8VSsuKTDBoJF46deWKC+M1d4Wiga3P63PSZNj8DtlaSJf+I/VhL5SdGrm+PMq
K5GLcr1fGwEK6y2z7aMw5zRmwqPsl9dCMsbnebRwwwlUGMgzjf0nDDniv2kYomUq
Y72uuLPOWGxPJhCAXSHhzVGFnZqmw2YmaGB7wObeWPiFmWk57b497jjYq1FEqPyL
Kuus4Zduscjc8SRgGEfAbinlu+UsR6EE4BGPiyz/VDHs36biVxGsi/kBZPJjxnvu
TA2gGw63gaJ91qJAfMs5m9KZMCbvfjHcWyav4bSIj5Z32hvDwmKkOJBmBMb6L7HD
Q8uLJiVvSHVIlFc2C9B3vs47l5CAnIIpEh8CKWlTdAFHSL/VfWsGC8GsTU9FBPkk
KeywHpUdtl74rZUGBnmICPp11fZb/QdhTV6Yg0W5attaJjVyobMjYZfES0/wz68n
HWd74GizLIv/lHZq+wLWuurj6ygxz2BV1dB4GRDb3++Sd0Md2n27zn2kBxE98VeN
qlkg52WL0wiisRmxsNsA9DJiSPsaIWqzrRVQUbQLFlTwh24ncHEVnIVQVOfQ+RKe
PSreI2VYoeGdOooTc2rrzEt1Uz3ImdJpcGHvB14fti9AlW0Fp68Y/o5U5kuekFzD
aroo9ls4/6DdVC04noUAuoiil3RiPQHuuM5UFt2PPEEKnnSKGndEOH1iCoQSIIRB
jJg2bVLPqH0J3SIFb9I254Vkot16Jk5FLLRQJAc5oPDlrabFeFGR00i8rSZIBwGt
Vm8J9Y8PGFzy/LZ/MCQXVCc7h+5x5mh4lmgSvUiITRE7h1gFZK6/LEG5LVMrAPtr
Grl1+LFCX6xaz3UORt8eOmkZlZlyEe7Xhmvd5tGFeZ2KKgnlZlBh99/GRWv6NVeZ
10O01jqGA0QIg9Cwja3Ys1Nr7avY6FHBKyBI5cLp+GHOJv+3aKltikNYnwCkK2Le
If+CX6EXMKIoEyz+Go7Cm87+dvgkELlRcUbxj2VN1vOpJwDt8GqYosQW7X6VYIWs
U4YZq4aXs2vlVyePkyVrUiV56fsEWwFkjebHyuHikZMpcimbSMa/pRNFnbPJvVtf
5tH5pjnpIsB2DrDt/aPvb8k5JOusapFvIj4qLh6i7vxOG9U8CtahvWH5ddYygwpV
N56OMeTlqLzTAhE4Z+Fp8w3VuzPuFwfrEeYfamptTTNbaxw4kzyRuCcTusZAZAF2
/idC7hBt51V9VsPyeFabai8lfs+UrSrrFs6I+XlhmCnnTAb0tEDTEltwF0W6q8AO
9l1OlVP99Ermg/9sgnc8OIybbcaU4RhY5k6xNF6oxg+Vo7gFjyFh5P7+to0W7klC
CDmBuyn0ofMlcwzvozafNCfptlQkYXvF/CSZ/7QoT4Wd6If5upwKZRVXoQBQhCEP
cFKFcgGdZ41lHT1nzqfn+TcD53yM4HTNFAboDnwbLxQwxhFnM5i0STSI9Hp6bXAo
cHDsnOs5ImQlcyuYE06gQ+iar4eh3nGVaaaAi53BzxouisoCrRS1VwpaxiNgY2dg
j2Mlp+G7Ierj389xVcQuKGaM9b4m1ODL0CARf6e70TovJrMxz91rGkuSAYi4VsqP
5j1KIyZrV68K3oukvAfEQuDVRX2j2Ge16i8IPLyk0c81SVOozcM1XLh/dRfXsbTO
V16XLRMwMrRTWZfF9EOhz4hcj6ZoatJd4adoYRkDFH9VXFFI9uuxPUWJPw92qFd8
AYTLu5cXSoEdUqK93nNzJwy3HGs1gWAawslVEqN21eo43Gi62JhyYqeWR4Hxrmhp
PCEXXpScH8nxyuheHUK7oaZhWnz85r4jz0mDFoADRkoUI7PKuqgiEFra4J6iCqE/
3cMLs3ZJgMdR/c2wWeF08XbM6VM1aOQxVnWsj1myOUJzR0K81CHFtd5rkdyvJvqc
NlCHQ+F/ylzhjFlChI08Kv2y6Y5avxwjGHh7LcoKrFbVlAEtZiw34KlTPgAV/UCn
nHx8yh5EIcJ2Aw7bKmLqaQouvBN58GIrjc3I+YNOc7D7uztjZpLT1Y5BQzA2C3tz
JpEaTQiIkU7qXfKTZMi1UnNR13Xp9HQ3sDSgvowE4MFrhBZHFoOgSpm9293WlPmV
ro9JopYwbHiyHDyEfTPH063mtrLfCj5fAUZg4Lihkt4mBgP4zgmGy6QJlVVs0SKe
tFLBDo77to+PUDCsKh9nAaky9jYFMRkkzw0URwfu6AvounVoqy018y6sL2/trRFM
II+OAcaMmjbpxbhyHvtG8e4/MQ+bWowD2E81Tok9LAvKvkZE8m1pfUbXeZjBPYVh
UmAiff2Oxow4bxIceLRzezb8nTtcRM+Yd+KYBYPQbejWDXBwPQYfh2PXmDdTl1lc
marKNXQQEZP1SWP7B/rHLBSL0sopIc7gSEo5I2MfTlMMlDSPbwtDEdlmr1mpknH9
gPWb5uaiWEx5y6No6DmWp7SjC5hoEa4H72hdrtgOYjEkvlBLx9kH4OB8EEyTOowd
+jBFqO/5JR/hMrmvCxEIjXo8XTDWEzjSVCkJuad6KBa4DGL1NX7cIwrsW+R3F6cL
2S+H8gyaa0q0QYQDePccfth4aefQIf76nM3Njr/Ap7lYuCwf2M7d6daw4qw8aJna
O76wHW3bHh3ZcMK9Um2se5jJfPNvmEe/wSl58nIZb0+cutLI55KWMnoqsQmKbUWS
M+aauizN3Oc+bRsW7TfpUONmNzIHycKTViVgGfbi2YXAfmDDOf/Ff6BWHqfmV69x
AXd5krUM/gG4VLqdOXi2fsHFIT6s4eYyADWuKc0yrpwlgxUcwWVeQJcI41HIf0r2
RcxDKtacc/RONW2tj1aex/kVKL+hqJqhRj4monVhg5aM9i/dOryYrWcueXJ/e2Uf
P5RQsox1YnY/ltv9b+fiZvpNZXgzJF9aDz7C3EZPn1R+8b3p60TesV4lBsugc4U9
MQGdcuJBZLsA7/wi8iHmMtr06BbGq2Xxji3n5s1Eu4faFtY4J8mIFvm5GRRCD3Qa
HUOb7ulRWzcdHfKiyHRymkdltYIfTw+I4Cjy/av2Azpgl8c8u2JKviaAtgTSfnVB
4Xs7URglUuWXUEwtEK9iiTS9fTum3z15FhqmP3aUqy0bcDCyc5nKom/QHU773IC3
rntkHHAI+aLQ6BmV6k2LbR5Kj0ZkT3uA9e8+iROak4qAIxoXXrdUBVKKjfmwECdq
p3wZ29KvwJhoI3vVxGSK4Q7mBy5doNfZ++KCY1GuyAf9xPcF+U9IpBkOW6wWAUq9
0pQRZMOdEJ6ZNF1TCfEJXvnBTHrBABvh9ObM4Ti8itxzAnkYqIUax4qNkhpavgS/
Zfsd7Cih8htuw05zc+Z2jOIoGxiDimIiKLA0hSjPsEZ/f0/6L5ppGb6YGO+B7ayi
xUINKHHIaPBGI547/wgfyOg9c+Foj47WvdJIc6MyJwvYJMK4YwW7k1XRT32w7Wgi
vCilW3c+UX5EOY9+OQteuI+alqtQ0tH7xobcuKcBdt529sFmeVk7ujTIF2QaB8wJ
MB2+v/nUXMjuXUCy8i+OQJnMhaINGB/gCqM1h6zUU/jQjqPIBAC+RihSt27nrBxW
Spcrr8zIASqoRZSshbnKNiaiTcVoTLSm/MDPE6Ma8GvmotC9l2nSslaGxCYNMhH7
ZUNRfkWLnvWLfJASPFubEwg+QiOEOQxxCIdw+tO4uLobgnI9ZrUy517tZVj7uNel
+FaGaq83hxCK3/hbCqoNCGSCu1cGSQYlzdxXQ1ypBpepEfGiYqZr0UtptKc61Rqf
VS+LjQEuG8HTxG9Kq9jSg782aN6c1qCig5IAZYlPALXpy870eKYrP5DAnouNAV6M
faNRnd9PQOUvDRv4Sig75fG0bdgMkoU1aTPn8lRlg/ND6cxEBRwah0M7BKTfrv6x
b3a/O4He3FYMsiYw9XY27Pb72jTHlhtqGaQKqY7bE8WmdA/oWlCIc25JVXkjMfWB
g4bSwH3rwGJIivPV3IASEfBLcPIq0akjgt52rv5KfqaCqPBdtebf3kjhyxoITCvo
5by6E//k+Gq8xc0Oz0SEaY2kq6XRkVQOPTAO6BKGdqLqvIjlO5ce3LHJ0T6foSPa
gfJPgVr+Akqt0eDd69VEeItt/uSuECf2oFBVzjCddR+mjgVhMhWG1vY7tIsIV1/f
UQzBlt5NhIgdpDQcLO9m6IiDqiN8Sq0P8Mscoh7OXz6GxJspmKpcYWuy7p2W0oH3
kw3BIPdUreEiK2/Xu5ZJiAypJ6OUtq0LknozFdAGStbp448WZGAlK9HgOVP1fHex
EJO1MVaFxDrKGhTVy6DcUFsgYbLUIBXmKBPA6Ym9PJmQRE8p0t8kJ1KIi7HxNt3D
BBDc4+Wds712DVYYf0F8ISJZBuniYmpgKdq0ReI+JPGpxRNqtZ05h6eumpRhaRCG
Y8W8Ve3jDwsFcmqfBRAOzJY9oa9+kZ+nAYwaYowucuLL/JqEB/abewH6P5HNxO0q
pcjXOpFZWi6q+quXpXMxQQ/I2V0xLjm+cfvR9KPi9ihMysDfH27cQTIuGyjazuIw
JKr9vDhfZCbP/p/+n9iI/cZALgG4V59lM5PbAEoWn8PSgmrGH3FW3fuxtzNDT+BP
kDIAwJ3SUJrpd/7eFdO/zjtR1Vp1vPPpmZU0glU/ETCQHVaZYeSscJnVMjzeyMGC
COMiKklGdqUmMWZGvaOTkZ9q9X/pGwz/EWLMavoLS6EwS0u1KMlwEyfFSa1y595l
ManDkXwRpbORUiq23ZDNN4xb0+rz26EVdp1d4/nXamhd3a/O85c8PCzTPd1UH4C2
FkkgR2xWuhK3X5uGUDTCsssD4Edk2Sl7kgFdhuBsPnwJyqr46haEFiomK26bk0KR
tZIRjTvBrIdewjjy5+iA46wp8iqBRcevc9cLxD+BRI0ByWccrMELnM0svwguMsZI
1+iJxQ12v4pxnAMyvKV4pvkaZIBRdFp58+XIS3pu2/MA4fjs1vTcOV5QN/ERfMNY
le9SrS/kr/5G+NJlqYoL4v043BoEQzj6Sb0WdhZ+veuYFrTKPLcxaatLVmmR+8s4
lreHm1mPXQNcmeDBIOrZX69iVQeHwS9y8hYUf7dNd9Bnv9s820N1TuzFucIoAu1A
LXBEeuUqGPko6FBbq4dyvCp88vzwZ2e2uznapFn1FHEBa1m4UIX4GoueRXTV3B+K
h132SF4ZLRSuUkPTePnsiB044ORk2sM8lLmTE06k75gK8i70aGhKnJcI4PdxnwgF
dfxcddFD1y/O9S+2HTcbHNhxKbytt63ICgvxFeSM3OFIgkUl0wBKokM0EIgfoyeF
utz+EkVctW/xGHvMNl7uZhxEIVMvalCtwp810TjefP0KKy/ArPErN7BkK+faehL3
INg7bb71mV30Cchr2f28d+pqgG/wtCCJsFohER5TSoGj5rZMOplpjnIXIVpT04DK
hfUe47AJQZKMpGrEJESpZlxmvI/dumVMQaCJ4VEGebfPHZrzIFI79zXPuU/s66Ia
ac9+/A5c1PrbncL3hFR8rM2hrBg/p4qhCLLhn2OTU9h6VcAAcYzo4ErpIoLzDrzC
61V6z0wg/ROPldMLA6rtf4XmsAVEPKGXQu6B9P8yaaOID0fFCp8t0jDRO0hGH8MS
1RtoO+PuDFSsI+r1nt6NPchFh35RpWwXFD9wqnnIgVoxMVJXKJaTW7kCxZoTDXqt
1Hw8h5Wj3DkQmUxyYQrkta3kpnZFQSkkbdU+dE42Up7svlvpLwmoy0pks/FaaYId
XYXKzx4y76wvKKzvqyCLgpP/ip+V+Vy4vHeakZoDbs7stFOmhNn/xUf8sOYMDSLK
YtoeZj/Jzn3YTUflFdqvLS4nzuW0IDp3GcrXd2Pc/UJN2rRYJe5xEixnlnJhK9W5
bBe7f4WEZ3fpM0hjaDo5X6c7WQZgfysee+2Vrna96lmoCLj2w3Sw1MY8y6Wx0Lrq
qNadfx8cv45h5+W1a8OjlNgfCmaF+gdkoh51fkI5uF/BKF+JofCY/DjA582do1KP
eqXEP5A8v+UYm8wbrcTqjXEy8muUQzn2/k+WYe7ua58UFapZZEdFdzuPoHH66Lpp
tytFenkWxWgx2z/amojN2vLlk6oTBAeSQhfia3XELVOGtbl0rC1L7Z6aHin9yxyY
LEjk9UgEz3NtKLyL03NW0VS9JWhwhcOJoOiGcSTsgjYHCMwtUAKWiyptzR0bUwgp
c0dvS57EP4w5hbybnjCfJNgONrrARsyU5l9GYbaC1DHIiW6JTFgZvTBfhRWCo6DM
JNvnpdSofO3qzcWwX6Lfn147esjHvCt3oSWtzULVkq9AIPhrzFHwWxKJJnDh4YS5
fq+hGrDZUAyVWLsDfu3SQpOWlmlVQiECKO26L9zBxw9QRb1xRlanqC5yjuSl67gq
ep8TeSL6y6IFYx6TsD6bk2yewoKOk+miW/Fc81zO8TznUPlR2MrtQ5uOhtC9lr1Z
adeFPQEml4jsdpc9vDugF0J6pqYzQ3aKzZsaM7s52SJGj6njDR1FWfEZGgsGMQkF
VqUwWIOcl8adPQ6Zfw6ufqtM96YnHIPF2PpSnPtIQz4CpTkOVC5XUHmg922HOIYB
0w1DgbEkI9autZEB/QjjOhot9Yy7LYLk56EAsFnFUh5jV2U3jw+yss5b3Obcim/v
UjfvHzrPD6qahrJT3QUTmwqjwgpi6lOx8XfS/LlYc++x0MYv+Rm1+5XwkhAFyaUC
HN6VmWKtqvP3EJLDvE4asfgytxOPN/5AAXwjw43Beb8cjKiCdrIqcGD/i6250MwD
fzh1OV1wNFETCHhCMpUkbiZ32hTa+2tdvjY+lRaKmHMqWuBwM2/F+enwqqQ8D7Pd
aBgWjoPVi+WeHFGq4cEGRrTGhFDh+WEGH23U1tXWxI8Rbumcwp60Ur74NK3YOBgs
Cfl0lAOc31Vvshc/aPszKxXbqsdvzBAtU5EFNljGsDBDom54SyHZH8a0QnREu48r
LzaMgvRYptqxhcPKPWrHNmxLR2deLrkGZ8/+noywMF1Y9SvZl08DwAZGSxb9K3L8
ILyvXrD3+/Urga6FQYVjcLvzAolRdtW7TO6/3FeSwl/sOyBRoXSapgkRHcoWhAPC
fbEP6z8aRIGao/W4JlkrKmta+UuGYrjb2DIouMsg/b5/3RxifU/EsBCbsd1EAFYW
y+gz4CY3ewHSUFl2CX+3cC4ZcPpkYC/awbJuMRecVPqldoYVbN8PKcwYVWZ9k2TG
2jncZXQ/Ul07zL6fCX8cHcxpS+l5tRhXGauzmTDKujJZTYcRH9UkMXD9XRjl0yYK
Tdy2SJEFn8NKRoT09HucF+FSEzOg9b8HSSfWfJ9er5nRvtEhtz6oRiWz60i0KOxS
6CbQDYAN+8PX9pIG/YNysXy9snDL52srAnlIKT2zPNz2udXmTJy9pi+67ssrZXYP
pSauPWK2gNxQVQA8WAjgmbiP5CtnEBFZPrjbqEbjMNN0AiDEUEr8BdqeugV5rJm9
Dhn8XEEzcYYQUNddx1B/dA7nhK41A9E4JUXpedTpghg/kdOefSgspbid20qXndjx
Mdp06FGhhUsdiJUzhq3POBP6ogYQAc1SvmxxQIDaOgkLnkqI7rsgfOjgLxfGGTba
zG9LWZOpemBKybTd6Y8faItX4K/vfLGZOfTsmiDQZTI+G0vwj+OuiRsBMMxkXS9f
UrHHQwp/UPAiFAIiMwex8LYtbN24dkV0V0qkosc3jc2rGZ+hh10sEmnNOrvAeOTN
Btpi/7VQ0Z2gKlsohQN3CIwoGolmkFVjcgaT1gEAl3UFnEhcJzwljpJIgM9lWB9w
L73LwH9AoxaoNLcruQD42+E7hAqfnco2i3HMagtkKOvqV0++yy+OUeliWjUPVkB7
IXCBcGUdHW4A9/SoK1svltZCfVRUVbcoyR4zfCd+2vUdo0QR3mRYV5mX62KcuWpM
ehUAu7CdW7GW0qdr9woaXosUh2b6F9s4plX8bTQO4vvko7RIaP4unwoDAzl99y6V
CRE+s9EHUthkCLuGpdD2+Wrn4mgFmyNeC+ZX5O4boeThdq+PxAoGTKEBy06DQmQx
uLCUt4878aoLZMMLD8EtvcaGnkL+XqNkhMvxeLTko3rY1Vhh5To8pWQVly6UcrdC
v1ZEInZCiwtsPyE/w7MxJac4V3f3bFUhLdPWzkoLvCIwWxnH9KxxdTR+e5bDcH+I
qzICiyAbJFcNJwXFgHzM+nF75ThpNxd/ZYj8Y6kG4cyW96s3YEBrYpr1jJoRaXUT
rNJCaX/meJUikgwLtMWBulQX3hq9UBWfcSFOTGjo3gYmHcz4nQJUwiuvYcga5pCs
l6Yjmy6MzgHMwCV/b5DXlMcoMC4yZQeRPxZJbFhqLWiwe0hEKQJTBjoa/EgclhYi
4es04FQVGjrh+HsM/Fk8ncgdIe5lw6dZNGnCFT36j59K2c7E75tEydM+JosD3gnZ
/wAL4KDv/Px9ztfpvw2jExPI8M5mEtQM9qyAH9f2w5x7YZWXt8RmHF/H5MgLv2Cz
pooqQ6Nk6HcX+XxPV/g8ZdQiiZyQx9S2YpaU2nxxFnTMJyA/wXV3V5qs55Y1KX1/
LxMhYclyweiQocBb/PKRsWm7ZxvxXuRyPj01ZNeuetnj6Zzg8TBqChjza2+vFd+y
QMwzaTFl54ykJup7CSv7P3x1aHlEw/DxWkDKFyNwnc8a94OTMwxzvyZlNTWrsmG9
kZthfTrbMGAfsW7cOstGnSit1hi/hna7si1Qo2rZnFgSkhvz+5WSZR1tRce4DcSC
791CehOWSplU5wFJVjV1BnKbe57C0wy37Z1q/Jm/XWSlv0i17C7b4ELpxk0gjtM+
aGoq+hvpXQxfMlKHghiaFFoVJiumrDv8QcsxNyQd7JiWNgalWCVL1++hGGYjYqUp
VMQ+uv/F9y5qL0S1OPb4+Anz+0jnYMocMFfQgQ3mCZiw8oxId/5LR+Xlq+Io99Pz
iD0wf+72Q8yHL8S8P4Gd/8YRiDHzNWHWg8qz2kjgbdEZTedBu5TGgjDfaQ+vQZZl
sKPlJrNwjmav9GnUnuSlVrrF5pi5l1QW+/UeZFeaAKlbqPZcRp30dVCtDUgMxs3J
stI9ekBJLIy+MKdKZ3qdVgMzOADvs7PW1s7+IQAunq1nI1R4FU20aq7nnJHlYf3f
1NNCjv4lSxERJeZChj92TfHEiL8xD7M26DQGDDxr4wO8c/b0kBEyI/sYWQcjgNDQ
mK4gJk8gD9AfiqMaMkSPljXMfe6hWoIrZBo+HrwWTtsXpORYNtILaewOT46eqp7Y
45hP+o3JGIdi3MxWE1bW3ycNsV4Y1365XOEXipLcJRSLvZbOplTfbHHX+eh9E+l6
kXQPJxvwpXHsQ5+T8gYsb1odsKQzOH/p2XOv1UQ97CS6prGAxWI1+5VVaeJAGE6j
9MjU1v6RX7TiNXeQRusqbpl+XdcO8uGhAK3e0JyB0xaLy8cvDCk85F5Q02O6NK0z
sY/fbXj0Hwaz+jqzSi1+eX0sIWQkpqvYue0LEoq8oeUfAMFpoLRZwpbU0+1lWLAt
7C9U7z9ta8d7ViBQAvMuQubZzofgnHMRGDgjQMg0Qh7Ghl+YJu1vpF72et1UokJ/
Z6fuhes4TNrNlwFVVZcDsqPEr3JvN7HYrWvE6Wtmem30Fqd7bBZx8mVdZJ/e2uO0
/dtA5Jv4fqzXc8bkRAmiU/cryd5DuqjOHpG2ysPUzX6jT5v5ah3MxUFWD6rXYhNF
OUqCCU5sHa4S8vIXk3s0qEKcDlUU8CgP3Ud4H2CPTAHCbk4JEMnosccQ9q0zkNKe
VDjFrrOdbcLO45atRetGQHiNO/791Rwh1lqUw4mLN8YBLAVMFs1L04XkgOStb5tn
xm0otjnMIGYc/c7CfOw3m1vV61qITsodEYvDSoItDU1k7okm6N2aOt8BRiShNVgF
MfVgMbvfFKYqZBXm91J8O6uoOIYB/Y++H53vs4ORHjnv25LywlZvI/AHjorP3ds6
IYfJad2u9jCJYdThGwNkQeR5Be3eMfvKODviOD8ly1FuhnLTjrmmLzkzvqWc+sCH
hzpehQqW/4hqQFw1tHzY0e4M6H4dAwykIGepz9uCDPCL+AymL+R3iBvssYgQsFx8
ofCCSFlCBnY+Y1siTvmZNeryoJwr/xOxWcXyBmqOs46mwpX9ga3Kz9epeDnaLYv/
zRMNgY/xgu99omGU3SBUXUhQU7mhtIx48dJWUbtS/OKSXelt3F+nlB3A8UDoDWPo
huv2uDeZsTblhK7yt26i/RK03dvdUhkDPSoN3UJdO/TIJUGilO/j+c9rA6IlFYE4
jFgcjRokGnQTGDHvttYj2GlvEih6Z5eKX88uKZyryBzdZejZJ0n6T/O4ThwSx/oL
FajiffOV0ayE+JQia8Nts/nzAunyXZOPsAKrc+icN2l//ZApn/oIJh7yXyymx3h2
ccINZtt1v96hUKSt17pAtsQOvhuEkP382yi6CCJPzOP2b6xBkAxTVVyN8mXShqX9
PFWBBfHxzp4xBmmVh4Cu8+cmQsHLtSWcmEJ6k5SjeAyzyluWJzwVhZj3WCAWrKZx
hegGaVAxWIaL1Q/rSSZeBtZl11tPZ+9BbVlQLNCwEDRnpNg1fuyLK87cqYtOnbUI
Ohy1gh6sZHBCcuarbyiREghz+l6uSK2E4SP7AIbOWdC7tfJOem03nDO/vpVNlsgQ
07UpjKnNyuAUkIGx5G4YGUjgWYDWsVoSyKYQzsxoa0NfY0WI+6hJ8NSken2nEoWv
/bJsHGOE4JJ2JsUoM08TrvIFWJK2Ms+dRv0o50NWc/V9qbj34taetQ0xneyy1lue
nC2HN1CjNM6EoqgTzUZ149I2kVx3gBFt6Coz8mOd2XSO6gy5LTPTpyq6HuyaZEV5
/iVaOe3Xps5iYV2OGnH1D2WGu7rnjTpGH959D4Q3ND3J5+t3a/JVhGS8YpidJ2c7
22Y8XMsCcOGXQIUanx0uCkeFdsv4erfUeYsjrrAmqr4LI8NN3tzOjRb82tAMDSb/
/WFyiAUIscMGmNf+8fwlzgM27Z9JwWb4oC0hAxlL6zcp25B7Xz9PMwaWI/feAt2N
vF76NgaiGCJKXtBX6AwqypQEpgBVL98hhDmVwLBtPJYbmpgixrLUkBQexAYgpN06
UBn6B1ND2T2JIZ7iWPV3558juL+HzSj1NHdwQPre+ofGtFJlvp0Nm/e4QvUCukkS
ylqt57ZX4emk9G1kkaB6At5MnUrcVU6ghjSI72ilgwMGtFMvJ+hdEZzJAZEvHk2G
sDKFyXVpGw4o5jaqEYxP1xrp2t7u2h1KwRjye8y8Hl5jKS2h2dRxLO9svmqKGZU7
UQNaf3BosHCQB88SNXgrwK5pnMHEKj6y37BU2mO/8EXIYkcYiJGAOyXhtMgsUpd7
GVxRsMlC2AERdmrsyZNb7jBgQyHIDZVh7VdWCWieIylquc6MEm4YjmFSspfZnV6h
K2Pj+ruDW0fHnjL0R124l1fWXldvTPra0IuMcVgDDbZni5VW1p2wmTzE7oYK7/4T
S6JJ78DTi8PTl2idMcgFlc6Mh82zytnuRN848B82iStqkWl6XoMDJYz4q+iL34N8
RdthniAINqXnmVGdin9gU/W+WoKla34v0tUEpJGxnDhISrMhDWmFIbtDlxb50Qw+
N2LT7SHOdCbITYkLgoTiRanNEV7/2bxdpSJbhxHeX6wFCZY6ymyJev3CVUl3KCJH
+qqjY75QFuKGaBXgy6nYeQRu8tGEeNHUbJZ+iTyNE6cTOuoEs4WtqhSe+D796IBe
aeu1ZNHSlFx5DrAi8zYud3DWKajn5sRN/UIsXeLJSSeHWXIby/CYoW/TC4qDCLeh
zrywNqxc+dmYLP/IxKzo5gXTvGHetPnTTrZ7VYIHtnheVx1BKnX0tep1B60GKXVK
x6/jpeESlnDo8Kj12QyriA8N4rgfuch8zPqE204CG8s1WXOT8c8RUtjLvemwMZ4L
Kfe4AW597+JjLFW3hwAljOucZ4T5LYr5BUbXw90P8rNZxeRL3s6SfUYkShvv1Tly
/Kk4Op5T489eWvnIuBhDYcCdwnCXSXgsD9VBAUmuBh5jkXElfU6KhPG+DchQCatR
zhEQiJUWjfCSpsZGB/CI8hPcvfy8D/MjEEVOnOlsqOD9ZdV8vpyD7+oGlHoe2dcK
qSjtdLqUhT7TQf/ZTzJ0/zIwgw8tUQGdF3DHfofXnixfEA1Sc820QIUeU5C6rg52
8bLtPqfhVQHkA9lsqhGxSaVtX/GYwSdZIGx80YhSBINeZnbJwCDXFH59yzAdz/EV
oixwPWB74IqqWPkAxynMn916Xorn86GG5ezY5omQma4HWRwnz7BlTmFmwutIx3w0
sXdKiHXS5Ak+2+ob5y6SD5jNuOUzAQElMv/NSWXh52xrHL8RyVrCQjM1NyQudyOF
KFnNGPHSB1Szl+OT0k51mTyValT12o+jNaZ7vfV1hMK9YoDeq+peLPhyzAYP/dyf
SYD4zGj/W5C9eNlylyOoftOHEuPQ9nQ48Xm8Yip74kIndQy5WiLxMrvsBCItWZ2a
Z7uQ5I4VkS3yy9GaZh7uCKhkZddlJrM3DjC3o7oOy2Lc1jNQlxpzqV7wyIxD8oqc
JZv/pm+VgZdKmISSU0Ln6Sn/SoTg6m7t5FCb/Qj03q9XpI1BKjOaFAumeh0gtdOZ
9b3kAY+GZb5/1dEOOs3FrU5lrzg3ymRw2MwXArnhMSP2Zi5gyez/QTpDuO/S2ddL
JD6L/bQ4vQzE35sOdAnQ4GbvLxSBQhKdZR4xL3PWBUN2DY+ym12bni282KrKFEw5
XGKeAim6B/jIZTG/+A+iA65HMPYQ3HCwVvJtyHTImJJrJVDVJhE76Ntn16G+krCt
GadrDkqo5Y9xMiOXw9X+zKHL1rm3fdh12xdkUW8dzTOR8QKwgksdXy8gjIXdtN8M
Tmz3+DOM4hpQhBMs/7om8Re2glnOQ2rqMScnSPoCNNwdW4taUOVASjLm+Qg/YMoF
jVY490mAdjr8dswLMCKgF0K5XZw2IsLva5qL0/jKM1GovtcHSDMP1SnMr8jzmf14
oJ+bj8UKYH27zT0lxFw0ylWsai9ETjfugNtR5QOakTGbKvaY9tJdMLPYRU7iJxxD
zNcf1ckcA2/9fAgFECanhhOtPvzEKOxqcy3Xnv856PWnR4oL7JIGO/h3WQ5jfGZF
UtwEJGHpFoOj68M5mcWxn1jo2R8BOzPPfTLJv8On2s/UKTdZ2p/amxMqOCwmtfbv
rN/IifgT+XTaDEHn4+KXtq7sGN9kNiNKvvp2msNAYQEVwsZiMXW4B60xV7AUPT+M
uH1A5x9K7LWTQmcRwB54+JTb71aBh2VNGkRvUNC/M+WEc69IYlU5BgydWewbjxAJ
w3Z9AUAyKp2qRhoZ6ORJAMnmse8VinwJT23MoIzVFFBicC4faIU7ri7LIPhc1dus
HolXN2myckfB+lQybVWtaD1S399SHW6nxa4Jx0XsQUCW0+GZPIj5U4s5dvQMV3Vr
T4F3tzZDY45FNmrSBw7SRJKpnTikatv8p8ykMu8TQ8DMPv2f5xF5T75FB/pQX5OV
7Lipk0F1I+l/idHFW3ciSBVbTRoSUa0BqAcm0Sy1O2+RATpnHkjxySJqoL1f5L03
CzuS5Tsxa51wlQ7Agmym5i6h22F5jaJauAugD/MYx7G0/MVyojgpFHj59RryZi2v
mCXR5IRPAVDbomOzPJhznHwfz49zbi82jHnP3YCPhwtARhFpKI+sRGJ8/wQ7M01u
fSI0u8fuSvP14ReziD0fyNOb9Ta63Nlj5xqxFJkHkjdHpnDwpMW9VocA7gBPkKQG
hb1TiRPIHmH7v5aZZKX+Ssf4hN44K1yG1miYpQJPsflfB/RlG5f2BOvAXIu7sOUa
BPWDs+oIw1QMoYA3KX8g0eawXMpwOnfiEVvWq42N9ajvgpCPRPvDASI43GoYUCwk
ATeascNNE2sZv5OpaflknR5vOGpb3Q2VLpuQKzZItqs/Xm+0A/UNdoWvTxvy07aB
+/KielFAeEF0IxrnVo1zPwdCXFNcDobZt3ue+gOvX7+hrifl7vhl7Z8uCPomhtKH
fn9G4EtJcV6W9WgRZZAoBE32JO4sTqFbiffR12B4oWSDaJVNeOp4OWVziF/mb7F2
xy89UrEN4hN95E81UHE93l/FgzbJS63Xm7uplIcsXPw/I2ar2XSgtKiqMgHXa4ER
9Fq7rhw38EFjfaAf/fnHLR/9GbWsYvJav+PyS620S2Rt1DxuIYPSMO3Kp5jremb/
TBqoLRGe7OucyrDfdtpQu2d682f0TVad5Mp/qIIvMbAh/3Ur3OX6klqrLeCfIKiU
ovfqRtOMnX/+OYlDR9kXwIRDH/etwqSNkcEtOs42pw6xTzlhWMeVRwDWSg1NM/Ch
JWBMhrhK2h9i9FsPDk/STZdgMyoe4XQOEXRrtWl8qhTkaB0EyMf1dxZBeRiTciwm
VRzqRDnKj158rHWzoHtx6yzxP/YhMV27Uf30bIqiAzVgN3ep7J8P8dM8u2B/zaXi
bCZugh+mMRFnRBWjr7+YnezunL6aDvCc53iGkcfrCwXM3T9xW442OY/cjM/Qt2Nc
b1NfabGMVyqEvgckjRJIUcOgXIRFDvIBeNAIL/syKj2egqtsPYOf2ihK1GeOPTt5
3SFzMso5YRYm/9LxYunPhbKCkqQLL6oJe5TY42wTC940Ujvm94N0W9p4t2Zx8UQZ
qbraHRE+PFHJJJ/cR7D/Cjh1b4UulGnTCIPQDYoI3ibWwFcVz+K62Njw0ag7lD0J
FwmRCLak6K4WOhbgtKp1pcEHPuaLjF1lboTrUs3N2hPJUFtPiDFZ3cmR+gOFlbhX
M071A7mUu9rQqvDt2ZewxmKNyciwRYpHk98fPdAnNAfeMtu+o7QWXbGqtneDPfhE
JY5YR9SkCvRruOk4LEafggRF8b2LVG1DSvjX8Pdw9wd7v1ORFZUmsmqxGM5A2o3l
+z+43GzF74c1tBTmEpHj2il0q+L00965F/GgTNdjspvU+SPS2pNqKMG/Mzju+j9m
8Y4f8zSNW0ykJBFtX5ZLaHCZl5UQvWpHaaLfmOTJ+PDgT4kb1XpaIzcQsYIfL3Ct
P1pxEUCqpclin+s1Z93YQrHv7Lkqbv17CX49sqxF6pmrJLk6kP0relrwW8cMwIzQ
WF6O/SwwQ4deckdO/6wsboTcgb2nPNwN3War5JuZktHYje7rToyn1J8yYKOH7vkc
9i/A9vDuM0vAhpFBUr4gk+nwAPmk8UQzq+ZNoQqojHlnuvmjFfhRCefwwNcGW+iz
pIeku4kdymBPjdd/yU8lt2xivB/qPbalrG2RgtQjEATMejzVfrpDVs8zX1z66uY8
porgaeJcsRaFyZST1SvR8muf9mR38vrBKk408RtrpZcUt9aZeZnSn8qmZfPF1hUP
N0K040S9XUh9y/vc2TwYcGTQ/0cb9DhNuwxGzVk6+JVEP4rW2DOm75hboScByWwe
s01Z0oIkp3ndWOf1YDN/IAKEQyzFWvU0qDxwVo4aTDyx1X0QEVO0WKMICZbmKAKs
GPRvpSwydLb6iQbVd3Gq2CKk94nVWCUKN5M3mNPzAUCjmpEuXyN/IvlT90jvnIBy
+9JZCnhqTs2UwiYCskZtFK255+Lzwtggi647dm4fo+xfJ/Y19A8YI6yqRaYATI27
fanZXgHaU0gG3QDkJcdCmCNBzqfvqS5tzzRPOZZCe91zFgYzSs+ENxSsjCPOjoNq
21Q2VyWa/NoV/In0X72wiJQAxQhv58q6LkIrBV7b9uKbHlvWv6K2vBqaQylegBQt
YVvko9zNN4m+syKN919GoCx4FlLXcz1jnpHcMlgxTnij3aQZVezORU1Rp1gjQuDv
sIe84Mcv0OzOxv+nSXIMFj39kpYSXMBzewKmVgcLf29JlrbEL/6NhENUTO/M7e6O
QZmY6XXnmgXw/yifNrhc4OWicG6rMPMde0Y7OC4ZpQr4rDFGvVEHobHEEcnKnFFo
wtr5D5ltmjubeL2nhpcpRavFqkXiJFedSzuu0FYlUMiCSqxZb9X9gBJ3zoQ7uiTU
T+zkIu6MQhhqTyI5JMTbWbbP6MDPwkPgEy2sHsnJE9iakcO99pGGPWs3lnqw8SqW
l/uy/XL4umgsro5veYT4L+41tam3sD4XIM9hHno8I3CAERCaDwxzbxBcrvYYlCsi
K4+kgfGMsqmdWwBQkRWVB/PN+eGFtVv2ypbNe1vq31Gh2OHLvjuowFVZW3vbNz5v
L+YOvykoF2rHrm4sMqOYDP4tWJuzg7lsC1N1b5OEmxyls6fds6xyOa5kj3Cqdg9Q
LKvC2KhTX9+M5gr+ptu7CpyUQrjazQzEo9dhNiC5sUpH6KSnq4U9142JIMhEv1pL
QeVJmvaA2IGNZi6UfiO0DceQVuvzGbkFHSogiwq3jjVNMQ6aBmHlw55N3e77dEIP
YnNSPv0kKpMkWTZtVF3EjV5vn/9cXYn2REh4qdlaZM/izTXqPMEVps5oXrldsUHk
23A7veAC34ZjnmHVQAyBumghcZEtOkmmkwdgPicVluYgxlQmGvP0HcVaR3478lhA
rM7BIl/rpjd1aDdzS24O3oUeN2cQ56y+byP3fQhzojGN9JwTgsAxKEi8BWUmf6mf
vedLO+axq2VHbDVC94k2TMgYWeDQYHhZ1orONaVcIoTMqQ5wOwdSq/lG5VqBVl/f
Cb2DEtjbQ1B8/o8jBJgleHBLHgIMlCH5PITz6si+KIxqychoA4xRHEQ9V+33bF9D
MVSnOrhuLWFQTlzCBg3gUSEsgPVVSil2Q4xburPIBW1Ww3R95YJybBwU5mwbHI11
z8tGwtWY9jlsD0IwWcRjerxo3bVfUOsFIyikbJPzdaaiTigXCk2x1R5XKZ6fihwA
BRED0v09mpMNjw+1xYbd274tQcwieP8HQ59OW+Z9c+nE2KdOkOCCbkuhXNdkqtlc
tnn6oTg5QD/e2ExLiKBLmHNh8PMhAX8JfxYSrLAShMBfFf1s19s51bgIZhGJw0+N
BcjdhmyH8USDbBoo3AO0Np95bQIAWgzNTZmmY2FWjx3qFiNxYLZ+vynGFMhfgbkj
HTNn0VxvNc5e1SvG6DhmTFmVdJa3f1dEms7e4FEi1LmBs8xBEIvrbUDbQRVsJ1aT
ilke9dwKMVZ+IWOKWgWnYP8MwO7DYslkxP+UlBJIUwYFp/+9C3BvxpajESf14/ym
eIlTyG+9ZGDpDy4llu+ds5ALSJ2oNGsE4rvURyxuB4qPD2cfvGAysbjlcJOaghTV
taOjnU5G9veRrnZkAJ6+BqVUcQG0JSPHt9QO+GjMfayH9Lhq2RbLK6RyqJ1n4bwH
QXP7oA4L5LkYakWeHxG8h8rnOHUnuNNvQ1p+I0Xz+8kSeNCYb7qWPTBShAth2LDQ
JoPJ3+sxbuP7B14nJYFaWmMVetbGvrq1Rogt8epZszToz+xZR3gwkSWnS5mcS5FJ
zV9LXI8K26U6l/JAD7sRaxJJa28YmRjzkXmAYWBCu91MlLmuCI9WJsBd675wPI6K
LI/QJL4ryXLd2PDX6hCLCW2T6QuNUIVVZIU27nEwC6xdmNKFzgO3a8Ew8GM3KwAk
huMtNT4KwjbK4G0hj1Qd0TdhPKrvYDpOdp2VqYL9XM4JY1wycLm2cQrs70gUT4FA
DwC8y/Uq5m+8cYk+xB6DS/y7kvlHsBpPyDFcO5pIOWDLdhi6UdwuLkHLYz+mKx61
sAOPNYBkWErGDIZ8VEv+WhPfWGFzc31r7c21pWKPlV41kowxHdXrp6M5Wdu6xfxw
bbscta6ikzimkuuaQcaJM0VkctwXhja04w1CrCYoZdErN1aoBwBCzIkFF3CPm87x
lQ91q4K5DCzo9cO8YcxFJuj8e6QhPaUzl5rT9ygJUTC/oOi45IXxfHxA49AFov0q
xKptCABPMIyrydQYn0h5drwjIH8BMItrwJa4cjouQ5sM1NxlmlLqsgO0APKAcgl4
IV4Jox04uEPau/SG7Kdu7rW3jyGJArdwdBphNfV3Fg/inhJ/QfDiqCikwAnJEG3U
golFpwxwzfnM58KcKxcAgfz12OgzcZjXH09hWx0MtV7fptjpyto8gfdDGmCQLHUx
THARfTEDc1raRz4WRETOQCRVm8vo8Rw/mfTjcVz0jzCkmXTR3xP9XkyeUiWZKX71
AjaIAGwg/kuC/MY2f1eouVU/7PTJ5Zrf3xx/3jPqEcLswrZtAJm1IxCsuYrDKM49
YFXeHnqA9ve04iQoY92JTMPd7vlQT42FMDTQf52K/oLDOAs5DzG6DzMC595ZxQ/A
oiDGxZwfJfMRaK1Ps549J3L12rr+ISu5U2LX59Yr9jUUa5XLQLTjJ3eQA8DqO+uT
aNCuhHQ5JlyQO9Og8ExWNJvegUBZKu7MXa3+657pUTkpwjib+OI5yu9CURBQlLAM
rsAjgwcanQZCvieCodpUYDqZrSk68N/7uNLdc406hOoI52wkdtLvc5jK3eduwsbl
LH4VHmlUOmrwKuUL7QdujMXwg15R7Y9afZ3Z1dREHL+f19J03YiZ/rKBtm5NaI1m
KwMfTlHPuIXiyvnhyKDwa1Q31xgU94SrGnwP34C/na6JYfw2I9y9ABIxiXc9qfpP
WvdP7IcKDpoaS8sAsMNAZ5X6Gy24R9SBQcQ11w3FiQxAdPXYFylKaP0cKTX6z3MF
yUmi3Girh6c0uVDICUWI3TLK3FsHOuIBDarG51WuZn1UTfcOto4F5DShCZ19HcPc
L2CUd0SHOFx2MizXdegzmrM7vFEjtUfBtlk0/qDxka+e5LJG7gTcZ2iGVW5Y0T2w
LuKVV4KR+2RGM3WvQFrKI202gW2T+OELVvgUbT73LyFYFNSv+35rlDCNDp2G0bXE
c9gswypM2HjFwWRvPqwqJM5DuYAdx7XKpiMJYlVvgHgd7mJdsSDMFijqZRpkgFrG
Pwl9CJ1P0cn8Lfj28TCGZR/3jL0F6ey7QQD78hvRNLeKtqUZP5SURVhJRK9rlDNY
boDlDTsaWVxtLEq/oZ6qgeWZhLiDC+Llqc6tJ/X5ctCHIDaCmcNsibY2F38AgA20
Pi3iRnq0KkZwg7VyU5PrOzNtLAXSIz3KMlzJWxcYgrZ2QWpb4XvRCI2XKLYBqz+8
gcNxnRlJKDfw/8ZxOTD5OR0ut58qywXTT3vAB6iRBI+IUa2uZKHExUCsXDO9JHuh
xKz1cgOuK5JUGiuX2P5ZjRABidPwO2l4t/xZYNLRyUx0yxGtyS6GwkmTZhn7MM3r
gVxXLqvANFd9hzbH3+grocGIvkv73ycVbtk8hrc0YAtL0H5m03K6Fjlj40Gf+jzS
sOK5UReGaiIcgcRq91jztpQkBv57i9uDNhcr2txAJrbkUSyi0mY19AaPtZsCEGSy
Gq/dBZRc2egGfczKQbiDJq26/atiMTAiaf6ay/52t1n8UXOWsnemSy00P+yo0Ag9
ao/aMP1kZLowk8uWx6b64CVID4cG81KkQ1cS3iPWZBTM3B69pqZ6ZBkl08TROsnZ
FKrz+BvdbexLSOzWolp2qqozEJX4wBZtNWnH6QSO7Y2Ao50en4SuSTcQoER3cNfC
zl7vADVFXvmzdSSjzl0lqqvU08szulxNKybR3FQIow3LIOSnDR8SQ3fxrmZvpit3
esSdEpHWDFzVxW3lv6tDjHphJDKNWPwiOWIX3Eyh4j2kkD4iLezkIUSPpGc+SRFK
4hQQNda5oH/bnsyBczafg73Few68Fw4s6MWstWoryUL34pO7UH/Anp3H56wLOkax
v7c/qohw59j/5EysCBhZy0bJsrpeJCK737Av2/NkG2zfENAfA+/mPrRQZN+zvQWP
Uyqn0AlxZp4O3Lwe2PkZQ/EJm5syQ9cFvBUWLAPjDQVXW7IjLELpMu5ngGM5C7E3
8FB2MUvrW86VjqzHnknRXd6sOGRrrL1AymjtByxHhKAfdptE/6wMHFFf1Ljr3N3S
wV8AunG4+jCErVuqVI1rHw3AS76xPtcCEbGGduyrym+2IQnESsUwrbXBG5udDzjA
zEwAvSdeh9tK2aihiH+ZhnltTh9U+RgcrMLw6S0U5WGizKGJH/Od86RCY4cmss7P
JQ7ZxJj+cd731nywd21HwAgJUILXkAdzwmyfN30kpROhK35y8IAjmUEcRbqtaNfT
478hglIg6AeOZGSvAa42zjzxOvPa+Ds8VYGsVh0XVSKxLIzaJYuki7x8H+jSjc3P
HZFvhisJ8s+mMKj8+0xcc9wmjQqyJV65AzBpDj0j6Txygx5tRbp0/iQQQvEKPKlm
JFNOAgE+j/Ci7paiGu2WgpFse1OTY2HNUgmJyuJNHCsPnGQ/2aPsO6MlQRvjIGOT
YciiGmU/aOWKybr8MAYhFR72cjwS8bF2m9jCZHagZuZBEU0eZi+0jcLGbvRn6wsD
/J4oXjRdEazp1wNivSRR+e6zhmWH6ThYsrrQRG0CSKcW09hzlpv249j9+Y2e0TyH
8/ZExtSmbtkJoCHFiCcqwfijzad4Qv9lCLHP8O11NIFxzw6vVzq1+Y2o1doSAHoB
DmYGD4MCwTtikQdFy4imSWjmyPhcNRDeCDe8pfxKQScRSWwpN3SIQGnVu87kXuED
RJRNltlZdUhHhJzfrn2omSHwPe89hVOrd4e+bDjcLDYuFqss8eIT0rKZz8hoNVIF
2GH1ifTS3ot9HCevzT1Eu5nmAzQKkBBREartWhiIkCuzDdniEBw40C2QvhGyM7Jv
iNLwvB5esZk8q3m5V3fsDUFJ81e24asNMdE0QvSNku/z6sH4vXSSZk8BmnZcufjq
5/oN8Zqqd9GgYVP15KMNklDIV02/7PNDCtGMP6obXW/wiVzPS8O8MeCa5YR27xN7
QJJZtHhML2KIQGoc4/ChJhdnDMiplgBrOz/GSx5zdogoM07yoAZoeGyjdghY7Z/U
e9lZjJcI5wNhH5MnbLWNJT/epw7+sWCC03rSYYHUkHsQOlINMPtoGLZc5HAsl3Yd
N31j0pMODjvM4gusDZYf1SjC3mvmkWoyEHqT6n3augssol1bHzXWFGLmwETZIicU
j4XrvkNb06RLmWflwhazUayJN/83eOg6jMSOBzXbAOmAvBJJBwwZpR7CHaBY4hnR
5Kyq1eE6+5yStHHy4e2MTCkdvIwtA27q9X00o66/sh+PllhG69tspmcJCAcc5dII
ViEWooPPDgZQn82N0oEriJJD7iqyDnZPQ2f42NaNdzknCORH39cyVieZjrXPXgxK
avsFxc/QcdIxOFtH4VlaVxqK01mRB+GB3XDeEXdrNzdGa32N3ELUfOfkn9XnAGIq
EazZaLa6st2pwy+e5wilMm2kxniuK1hacmV9grPK4C49rEtwzDl3Ntuhi0Ox/zmH
/QwwLqqqav4Kzwevpa8iIiuHNQMU4Nyd731hiiwmV8ncxzUkHWbF2w/sOxJsjPdM
6uqYBYYlSLADWVkvANtoqrRNd1f1Wl5pgvVTQPpx2I/RIMJUOV91jqZzLa7jlQj5
igL9Hm/ted77Z1jD+GpgmCiQq5Tnq5T38I7S9rSm0ZrEOQ5Q0iqc1pOLoOP2yvFP
F7E/7cfO1oFu8URRFWlo/LVHl+tXP8ftTvLPQo/MBMWJyVrgmpt10mxIFJJQ1r0j
/eQiNksykpMNSjtf96GJB3RIsElZ7+IFAeKYuAbTQLqVBI5HGKT0qOTzg4GAQkrX
RoKcet+tJR1wpG22bEqaCCtPbWRcVhajB2wu8KajjwhI/nW1jboMA3E80vEu3oBv
8jQzWCXSTtWMg3617FGiz9OJI7N4tC+5Ta4bq2gyxT3lqXVsLEOkLNuinOY3t5G5
7xmLQtN0odydEYmXgxZIFk6DLzrj3ZGQw4ySqS3AQwUC0v4oszLeQvQchJ4KegNK
HuKcNCGKTFQ6b+XIkB74BPsC13y7nJ8Yiu/bxOoLBCueGWCHGBpyuderC1qh8+/o
4TGg9cmkq1vBM/L4/py3TlpqSFKpYMFXqztGxaqVYU/ThBCptHS/AyBSHMtjf4iy
YekKAGfFY/uVdM+nXg4VeGMEfPPw3B98HED71vIxRohMyLuu3FjJtBFb3HVGfJH/
ryZ/tXrUKBwhvB0hJnZT1xtWZPJoo1dq2RhKvzSw6X/O3DS8iXwi0B/DJ6Cge/2L
1EE4mtif+n4lzFCKxtchpROrvE7y3ulqFKHeIaYJKZwuyWDd/ROTyatML085kQSO
Hc2F/HnpL1QR9zIe4LnsO0lcf1QEpKxhDQE2EcySzOTuONrZgzui55y4rC9IMKCf
w7r7t0F1v2tZi/fKQMXEjk4KhPBIYUMuYRGBhpby4bYC/NDzKzypD2G1s2YBbTbr
+lwllXl99bZFDVOAL9BC9OGi/DbI7oVJZknClLqdmbWjiAFQLwzWj/f3iqFMJCOR
ZiXqJnv2k8wLHnj0nX3WXE7Y93zMx47vKDxWWR2V8WnodZ+eVmEtGOrU19SST2Dk
FFviimsrT/1BQl9BHytSjLBiPjRa0NKaYCrvt2QN2d1VQiaauUthJ6hf+aip5A3+
Aeg00E1pzvNBOxA/HuwT9bxZ2WfCcwZN8WkhdwdzQYSgKDpaHNAzoo8Xq+3NYVxB
YoVo59skkb7w6aTi74DJ7BcEw0OZN0ndygYxHd8mj1BUB8EP5u9ZLenHFVSSwRbl
aBtFx6h7rFNxtZQiCoqph6h4Qg8FvOZY3aO0XJf+CcRNVSst2xRo4oUqFL98DnKU
juo7X7DerghOY27isTJ58SIR9cnLU81r7GEjNmqzyulH+WnLk1xXfkA4KvnS8dRG
8ZTt7IEs+0WDnjA4B2FzienELGT0jy1BMWXFJRytcp2Au2r0BkRshgKiLRqdTLde
YQ3io93C2VVr1FA0uG61RvUpzEEpx/Llx14xVWBuWmyVJyEtqtWsnZR9taZzMw56
9R2CA3VxSNneiTich+Z5cKe6IjIXrImJNYMM+MjGvd6pZ/4HE/ZU7os57mRSgucy
+xAqEnrt440iDCB1pN/fuRQJouaAxCN5wUCY+en+TPkvEytcI0CAZRtxGdnOZB+9
DWOdlKLPUCm42TXr/FuEQ3cIANPOe+zdyye5/FzK+xQZJzgAlBwiPJs87zEcGUxO
e+6EFNcBpLRCXTxcgx32fi4ZrLsbPkzunBlEzGSiBGzjCq7ZzmPfEjnj5p5FmQsV
U0a+mdEep0VGfKJ1IfwqitVIXCbvTKPpR9sS5mj4MECDNvIoN5EL4gqquoHon7yf
E6+8iHDWhhgzGXKWAc+mdpNZ7zB0/z22eLt5Zrfdu7X78k+D2w1dRPvjt7hgyIVL
n4pUN5Km1CuRoWlHdgPitbiSBGiGToJz1Q7IpN7SokXIv9qrdyBW9WXyMl680o1X
6HekOHLknsuRTlW2xHDKKzTQyDmNYWWQYn9Ew3AzkcoEglClDxOWJNDmdPbhKm3t
cmaHY96lZ3qLrTLcYHVueDzV1clJVInm7EYy+GJs3qhMm5K4Bo8FJlLWC8xlreTh
mmoMJvOR5BgScmO1/kj7Yqmj0DWybZwgrF3jcwsoRJLEUMneRFKHhOitvjjJoGWZ
o3tNkAGqETigk3ayPKV3CShgqH8EsncHBgSIbIjuuB6cUbOALDNF3DXo73M88Ye/
+evkjhji/BN5grFsnYccKncEkd4/WV/4CvolnfJQ9TTp7jdB/kA58y5QAQePO2Wq
alL0iTBjoo2UQfxUXW3WK1r+IzAj4indwTNjRTuXAAT7a5QYCrMo7lkkW/vzCb5G
St5m4i5PtwN468g72K68Bkz+4JbJSYRKr0WLkF9Wu+a5H5nkQtkM29p6hq8ki7MB
TtJEHkZxQZySNLcPzn8V8Fp30aAsJPUeVEhcvlltfdVROnZQ8V4JTXry0JQYDRik
2Knd9PjqJSAVP5AjbVajNX5qek63d7aKQ6n/7yEIeh6nnZRMFZTxrdi6Mi3voTMf
1U9nOTWs1pS0ZOoDNIMDVOJGMerBLJG71ldw7b3OmYAcWTLwXkAWwziYwj8yurBj
wY8lJRlEe4zWTczumVQIbuJ79GYTZGbcNRJLdMRSnv5kn0j5GCFiMIvimwbTj0dK
QIMODHxDoz3Lyy10xUi94UoK+MyRDytL0JAb4gQaB4roIAnkQ9PzNZN2tyXts6qs
z76MnO91DJPcst5H2wMANZlYK93Mhx8FOI/yLjGU6l32RFhPJN+PFZ0qqWBCWObg
5Eoe0Xh6hmI9Him4F/Gm0yYhKkBsWU4DYpVFi/IsLa0RpT+fvpob6CKs0Nmgdl+i
i7Fc4NrYigS3oyBye6o3l8Hnv1bBmDEy6mFnvhFadFiwvQ62x0uNwHf31YR7FPLJ
ftEC8HDtSSiN6yAz4BTe8um6G8Qtuxkm1nzYJTLDOikvmDpYDW/Bit2W2cj/7d2Z
FmMypLcZmDMeuCs0FlNv4qVdbKq+FeUI3dSb7EeyJpY5dz6/zkr4ZQrAvnlqCYFK
2Srru35wHnGrMLIx9G4rBWK/Ep422Zjau4TaN4lmIsI+KsgQb+2jJv17cfnMsWBC
7DBQgcmBFBQ2pJjGaaWBLhx8yoajLZe+kDi6vG964K8jowoW12mPmkA1uGa+5XAa
KRwInzyZD7sGe/o5L6OgfRfNpntX6yQnG/99ZQ4sbeEfrHUB+uvoW6kkkLGUySUu
ch1Q7mwBw/hulJKOnG4sWf8KeZWFDGyvigCtGdX9Hl22dnj34IL9ddNvlaNB6CCt
ES6MT74+Og/e3XU62cwHJrhLCzmBOTWbZYHCOS2IzijjUfZSZsCiKqtkYklkd4ec
3MN4JzpHSDbc3/K0u9f6zjlc1l40Y+Onob7FiRGrkZa8UNjdyhy0Ca5prhXJ5C44
ACz5CXSCD6dIDEK+SPBoqJPhq4fyX6Cd4InSzgnjltPjGqVYGIwRMU7inz3AH1J9
OzoklqXOu/Ct2c5Hnv6eDZ0sd6yU9oJgFANt8JTeEwTLZxZaZx5iwaU17NtqGXaK
svoJfCEuFq3KrFcaiKrAuqSqVSbGd+3Q/P2XbtKx0KGUWwI+KRrfUqvscQfbv+wm
PeewbYSq3o84sjb+HN7ZYHNypMUvIC4p9gIlJ/JdwoXAI4t3Fq8akRFqGwCL4leV
AFuz1Wp+qrJ4hYot6WocR2J3OiS5PVm9/oGWYcQUbY928i9AJTGfnvZ73rf8VY66
IKsovUrAW5yOLf35lSdH/1eAxmB0sKKfx2c62j+OH3kQ3HmFIH87EuOEgWQE5jEq
03DxXsomLOsQqFHAYThAlcinCP/cZfbFuYD4qrrodCN2CYsu4j5uGT9ycwMew0AD
ifBcd95Thg7aM5/rGmSKGT4azmn6G4KZAXeuW+E+t9HPCbD1ik8dtrsNN4vxYeCH
cGceafPdkzusmlH1Cq0HEEABjHeQBeAFZxwaKl2lYtGHGt0oERebO92Djt/Z4la0
7o/VrcX5nCF0y725lh3779C8xWIVmMBpT1RGS5r+eJ6uOfCBjW2j1rncfvnXHzbf
Y99XUFlgTgrQRRpIUTiLDz2GeuRJhHXNG/rEyEJwZrjzpAEOxgfnCvClAd5B4ihS
/pVE2lmGafLFXdqZAiqmovORcGizmXP4vkwoxOHfLlQYIohB1cLNCQltoNHkSt5G
vKkf34g/xOR9FyYOFdgPwZz17P8NReVBp+88XsAI92l5IUAjrSLF3DAGfJ769Q7W
M3ratuMtDAYgSGEnEG0SB5fATvKS3GJoMFCPKNokTmACCpcZhaX7YmQBRGdT5A0w
ORpmGN4+RFJln4VJZzS4MmvCNF+43wOItZpgvQU1M7JozxLUydNhW/nPC35yN6uR
48wi2xg++jE0d85L+Fv7CEiRbNhVblvLJpd45Mb7IEBe5HIST0ApbQiFeeJY0CXG
HGAD5KWDBrReYsgqRkbYkX1jUVnRTCrYlSQrfvykvRsUKbpP26P6AAcwaGxr/tII
rN/qj+K81YaNRqc5O68GWyRxXZM8LK5TQgl2G/O5oejRKbcbc9tUe2PN0jY/Ch5A
PEbK+pS5q6Uh8gvD0Ga7hrHOQS84tI8aFLjiZt3w/2BG5fO6MRW98syIa+lbFrx8
ZYV2GUEnu/QD9XCDEIHEnCla/K1umLn1Cs73gMv9F0xSPqw7pYI3qQj440PKblAJ
5y0txXDtFVsgqb0Dx9JuvePsdDaPp76TNxpu3jSGldgvM2LAUkrl/EE/niCesixN
HdmwuwLrfT6MaOOPdLvguU2mnna8VxJs2WQImzqPCKA9+L+ouxHlwhRAsA7HNz+9
qEajl+plaeCwLVha52Lppowob7i8zl8xZZ1+dJkNZxBWJm7qydLhqrVle1GoS9p6
SXEp49DfijIT5WRhfuERANygEC76VcR4Hu6yRGMIIYcsxrZBmcxkfqVlxliCOK6Y
aDB3W4inUMwWkiQ0p/fBkFinKGl3EZaRfEkc2tjNB8oU2ceXzXBFsyI37sH+Gbh8
OK8WwsRdQYZuuAJ6ZB2ouleGCSXasoVRweIHnQA8CPk6awMrWr0kMvO/vtrKZ2Mp
blNo3WxYhEliviulZ0KGKNModzQlMvBOXo5qTqoX87V3QUkdVxxHXFItKmNNRbPA
cBtPxOHYwoJSARFR9DQWirusbb/1Y5MROu/ICnJ8Cj/ZdhbOw21wqphYU20xfuWA
BSU9LYQgp8BmDfCgVt6a7YHdtjYRILyz/MYzkJw3zZiKGI3pKpdBu16fk2eHCa1V
rv2lBZj6MuxFDos23UAg9avXXz5GOoqtDWh4Z+MEJ6WFUDMwq1KNGPGeGWSyyMi6
I8DZrYDUcxCEvdnQ079rwKKdhqyiaDtkfT/EXtW/I8jT+V417nwP7nk2StMPxvBr
zVcG9TfUDrylHHgYLxEwruSq7dAu0w4GPRj+erkHKRsirlYKJjeXkYxnBUj209oK
C2eIJ5ELBuURGbdeoce0+ohjUwQ3ySRzvXaJFM/qc3wFJ1n9tSUX/GRk6p8AJJ0k
6iKUPn94K43VTmnxG9+YwpADV4Zsg+9XoL/poO1WbPXVpqwKPDLlS4SxsOHfv0mn
I5/tMFMJENv/KmPmZlp1yfiILHOAynDFDUUZ8Hvgy5Kg5W3IJSiU79jcngUwIOtK
Eynqvs1gJHSfSEmqvI/qNGSzqE7ChBfnf6NUw6xWGs9cNvB+VTp05YsOHP7ygQCl
yORZLDKkq5C9YIPX96CwX/AVzy/qL6F7X7gwIcF3DWS6o12jchPyycx99r+6+QwY
RL5jpmX3pClr+72Ya0x/k/hOE3WTDix3GKjuBA1XKGUDPCvAs21THKWFcJctbtfH
7QNgaGvrr/jAcAThw65vuemYus8Yo3yutKTWgrm+lQW55HcJgz1eQ6gLwM8KKlw6
bZSX/pydaao1M8xmYikXynmPpCuAe82iRUj24M1zV57mHC8gAa2EGP/hUPVyplkJ
zG3UrRARHKLJLPJn40YnJEHnyH9Sgr7XWE0Lg/5BU2vWwZC6BFAcYkiUmUTmbd5G
msIyjYvuLmGPRXu54FZltyWBTtWN+MiOsRhcFCxeFWB6lWMnOMAXP3ItJKCIUI27
LNb8170LjLKyd6QY7rvx3krtfbpIo1lKHCbMFMh4Vo1iUBULwIRNKtco7C3YZcFT
2Ym4XljuwQqFCFAv7jKT0ZjLW0Wzj1k9hHi+1R0mPmUWMvR7OoGZWMpo9Dt5mjU9
3y+2us31bkzAj/8s8Bxnf9nngJ7GsVrglvAOYRWBvhHbgUyao1wdHOZMyjssiTha
ggDvsYWVGI38mQe3Zf1JM+GP3bHyRmshAG5mmo6Z+ERTngC8adNBnv0xA9E4IqMY
QcFyyDJctcloOA1iNhFlsmq1ws2LdLs0jDJ2uVQj6JVydl70JVnMews8Bfzcc+V5
Nxp2AcZLrc6oVI9lmSCTYPsmoaFbsgrzzRWFBD6JDlIQqKmABljIdQw7iGgFNd8t
6yyIn7/gbc9f5QZOA8WheiXiDO+gNhaIcBokrc9CPiAXZDexwurzUc7HAiPho/FO
AlcrO8m74HhohtcbwonDVcOJDTCeachgkCEOJ2u6FdejtuWQQJT2uA5hANJfScRp
bwO5hF0pEjKbPzSy3LXh75/1FbnZj+ppVfsZ/ZMzLtuF/sZfu9Spj63EmhtTJsrb
epH2Wo0XeNNrC3pbC+30MX6Ommf4XqgXYw4C4uamgxz2VrIR0qF9DzqPuSQ8QnYJ
im5HTVwj5mz5gt/px02yOeTvRncMmH0Pcl1uiU7sN9e4LxTLBII48zJt4I/MV4QX
SDC0TBIfVq3XnG/by5wmaQbrJSXIWfTTRBy1TgJr+hUnTqTln6O7lvJl9IdNDdQW
o1yb1VYdUHCkB9GVaRIZ+ldieZ3M0jRI8PYGnrNYSpNK4/QvKIwCSSU1FgHpPT2g
za0fbuLtGR33BbwRmvPtWd9pzDlFjZ7m2g6ZnbwFbi0gb6TmWgrgpGGaBZJTzslu
O7F1rcL+bRW7K5RE7P9TMmqB6mx0zBY7ON94YigXNVQcwo4CJIrihxrZ/+MKHL0z
TY/IsUDtDkwXDR8Vf3bGN9Ig0jVuegUUP5wwTcs8tzu1PJTkFzrEgoI9xdL8DG50
e0AnBiUnxl/U/HqoFd0/b1tIDqUsWy6i3f9fB6dowruhDGF2FFTv1xLusfAcficb
VGXMz0+rDiNcYYH/erKJIYQA3pJZzqXbyvfoLf8I9a+J/zWebZeGOsqynqLFs9I+
yGkb3LEU+76nWFJP8/2jZCCCX2/wPO88ZniLp8E+yuABxPrzw21UHsOhqCQSKbfS
PW1fllOQPGaLmz38u1dPx/mF0KBzRf5WNIGqO6HO/B8VsW8Vgw5PGl7Z7kxfA7Hm
3KME0rNZOFX5Haj18qQa/1HxWiuLy/vwSeOt9PCagHW4VnVku6pJ8mlgOlmY5l2I
4bteNHl0BJYmI6i3ovnbzQ1/OJCbwVnj/y/hm/yfdqZe2B5IVZv4DSAP0jRf+QMd
SGs5ZYo9uKIHuQTN6tuucJQ9eRjd+HtqhrUgO4hfY/p1tHG2zz+6OXBaXcfyNzha
CsiS8yAjQx84pYi1iMf+5U5SiyLHh1KYVp6vLWB+EY/C4GIBI/SgEPllG9DaihV6
OA3AcLhi7x3aPao+/QYfSpPZd5XvC60pbXOE2Ok41rnVQTC9URyS9y/6JiOW66ej
Lak+PjAqVuxNECGNTGpLeLGCc0g0psap2spwrfFzvwAs6ZLSO4FZoZaHcAlNFyZ7
muWgH9b3qyNsoIZGRNMdjzweAEM6stQyw23cYIxvL+RMPgAORg6mN8OyTn4HKvpz
9W+KXmaPDCwBQbJ1DSPikn2RDJ1cIA1lugWpoejRuC72daX9VM9JGcTLFTfye2pe
yjdpv5DuRuZlRAoECrDgrT/CQjtAz+Z+0FVytIUBzhFIfqEIDZqDf1mzdKmdrIAy
oONwxCz8NF0BtowHYW+Ti4NOiYtrUu9S0X8uLo3nxibDbQaIT+LkL+5afIFvHVxi
M9613Wy5wtq8XxqLWZR1y6u3XA6zi3bDT5A18+gguH5k4+ajzBAIU05iLSCIOh+k
pGPd3YGCLAmpVp5PNnoSCxWYuLyIdBQy68vKcN+Xbe3aq0TWlcHlJaoRJcaqEhUP
jNoumAEp3rdVTxDdUOa6kTJEvjExFrZyCNI2rGksKYuNAoPVR93GVgj8tLWRWnP3
0LasvKLwBNIfEgsRwSeXAaB5IyTWV2ErWYDgkwRyJ8TlcFObjdlOoQxlChwcFEIT
XT8q4jJbx+oW9mJOrEjqZxGgQeC4UB7ftUUsB2GkJVhd2jk0zAZx4wtgV3p8FYW8
I0zyZC0akWW8tb+Y1WUAX44MKGEGT/ntK5f9u+3SolXyLXmo0Pj1j5oiMyagKRk2
ueBFAjNuGKLfUptlBZi0E/SJ/X8KOKigYQf0jP/+4wr91pudK0EtkqE6rtJ8l8Qi
jKs4HM0InXvfmg6IJnL/LOGe+B/w3HUMEmkhSW8ZLMejB/Z/56Z7IlFhhalt03/E
3Dfao9Q3Vq51Abj9q6LpSxu9ooo2pbEoHFPP0QBJKDh+TdOglBAH4V+U+0z3lLFw
AgIHR8wV22HfUS46I/f+qiIbRc+YM5pHbZt/tPOtu6UpBHIitTpq1IcLlnEB+lQi
McSjuPcTLqYM5GS5BeTfhy3Aqmp8aEt/imElJ3nOXudaBzXPSI+wIxfR47+vncxt
VeskSpXtQ1zzN7/vRrloEepuWpFDgAxbkC1HaHSDvfHfFChIy5nVQkxxUYVcvVj0
x7fgUnGON4by4pBrpIa9JMgz7440WnsqnhlsdepWVtHXplRWQ8DJQmD9Olqc1iP/
0UKVKXkHTNfLWP6JqWRM1u8J+hi3hCP1mWWJTxEf/HIORBYdiXaFV75M9kMsWUta
IIa1pvzFflCuTxC7sJLzsXDvtbqaL8Qw2OLUa/0kNcS/KC7Y/ELBcyPqJRZBBwnt
Qh1DBG8nwd1s92u4vLtDk5G2Ops2oCHbV3T7CA1C0mej2L7tpeUyEbFmQELAno1Y
7ARJYnrsoc6uqZvgDkPBM5Z3YJNw6n3ZA3lBZ0PxRhPrViIt1xgxnLTsfk1J5gRE
F0nqT23BrFih9eMbeUJLuBQpSGZSKelxyvdpFG2cZRfc+KoAeuZDBpX5Z+xT5e10
SZJXa+euJlroZbnyz3UFaKiG5EfY6DxvkFN5QdfkBfz/78UHbrW7TD3hKuOQQpih
sRn7jqPER+3zb+I4YE7dECiCRdIb00gYoObVjjzW95Xe7NxNDuzDdou8yB61t99e
lsMIGzgEXxh33TFqv3LNW5X9ChIKdP8vcXgmqK6Je97U8q8HLnlVomgCXfeGBWZq
pLJRpW5nrNVXERNLm3+pg8XaJ0w8he1PRqs4+Eo0riJeiXLZrqWUs/1ru6+pAhkF
U1SGMy1mfVw7p5xmHOWXwEA1f123datKg3lJvgMvxI39MB+68SicvBsX1VLoD+BQ
/ArcvIv/gcOOeJlToaBvGAZ+l33CttULSDxn+IS1H2gneG+1v1P+2DseEt19STEz
6LQRiQypzOV4sjoJzi0S1ZCszwG2RW7hiT1VSRoCeFkTABsgEZj4uzrOzgMXtJ1e
iEQDEeCe8xdqxgbEBh/+W1aLj0rI28sfGa0tQujkTtpjcecOm9g2YusLuqmUFG6d
SY2fK5EzFUHy1JnZBaUXSBgXBRXF+kUkQSsYXx0IlHwofR9UUWTZje8B0KrFQOXj
v6Z8QJ6sg1EBAfcjdVA76xoTg7LVaTVzwOwXJj5hZoH0VwluxM/EZCYY8D62bjQk
gfpjnsUw20HP2LV2zAV2C0tfCW3T7aXfOCPHXvte1sMzGTwlxn/ZE5ssOvT6wAa0
IOxHqiWFkkbQR+9Kz03WcCIo/t2hUbSylLFJHUWpIxpkCtL+z6mfkFW7m5cD1NGx
EJujbVKua66Nqm7BS6f0hf3WBAguazL3O3dTEaCyuBRI2sWGjyMg4fcLdLkrm+oL
RfkrScNLh3GF4xLA6I0NwlDe5m7qQyXTrA44V6tD41Skb8LwYUln+/sCzFXBGiWY
I5Elp5vefk8oAq4iTlmn6//SZPZC+MKYA1Mec17hTd5XBBj7JA7CG1wx2A746zkw
u+oiWkuvZ9WvWSkihWX2o61zx85+2S/uOA3pPj6HyWsw0BpbOsd+PBDWCXVpmow3
lWStBzq3iI9smtqNW6z2Ge/sL5Pl57ym0MFSTN36Cq7FT3Vb7aTvgj184CCypGx2
GHPdQcQZvlBh+kFJahIBQ4EhP9da8kH9Ri8vwz1SlZdTk8gfLhE/lhDO3rTpK36V
dnBRT2HJ8STXhkQypTOfcQ91NoUpslNp//CwuxKkfkuqeuWxGMggj5573tWRYxzo
FBFz/WrYPt34OhPoYmT/+Pki2mFQ4hB0RCI3lKsSeC03IZxolhj0k4DtxTNxWc+l
fw/KLydQ0C5t6dnulLH5WZ6/ht92Pco/9RKZUl1DgQGBn0AxB78N66S9Vgi1QUha
daO+b2XR/8B1ZOPu11HKWOox5GLyFkNHXG/QGrMygdQFHl2IP0QiP2XY/4moOo7e
i8Fs1QiUJ760cQJfRb/YinbHImnH7t8qabfHkaWEpjpCw5uDmXUtPCcTrTvFu+Ka
LN8vdVyRsdEoscKyEbowwZSvHEuUK8k58XxaWbCCQqMB1BZvXcF50uvGFM8Ts4vR
5ZkPetXR9PpI+ZnJ2qS/HBEP9kMVDgJC+UD5LGk6cCajb6wN283PA43iO3nJ6kXe
AWzV8DswAkbu/mO59h9kg4YtmfcEHqyGazC7peE13P5yg3eiOe9b5Gng/l1yyFjq
f61b6/eJx1Ass0ssxKlTg7Vsl71srnm3YecPw3Z9BuvMqoPQQkmGPBV6LAEe9sf+
3DcdbDVKotORljaCSWFJJbOvklI6on99k5GBkfTiNzzjHotcv6EMm5rGbaKtbnTD
ja+zgcCIkE9nYDfFO17wtF3rNx04ZZRfVv2nDNq26gSY4zRsMpFyFYRR49OtsaJv
JQ3p5kdNv3iwl/7TjCU+xswEbZXoEXTL8DBWa779B4lGlXPnsStrT7DeNrPSuoVV
QtOS4FqCaBkVzDAtANEeCsD9LpNEzGGbl59mzwOzX9huiK7jK/578yCC7wza/LrH
a31mCwJj98423xyvvHwQmXM2ebF4nRbHhhnYUa088Kue76Y6hf2PMk5UkosFtaTI
avOtrFMCrm0R+lB/gzcNbebC54CuyaY8t4Y77M4aqI9Sn45pYgyYmQOs1dp/ZQwy
0f8NvPzT3Fiks8jlDjs36nLO7JX6xD3hQrZNCctLsn24dPlMElivJ6vjR7+F2iTV
vD0k4MWi0DWXsFHdJG98xZtDgdDgP/1Z4kCK2VsSNrmI4Rib0ZZd/kEAfGj/gdKl
1LwAJk0N2v5sr5Sn5BUTW6ST0Rp2xwpJj1ljs1iAlpOtMuYfpTNnobg+7ZM4XJrF
lLifNTVsp6RjzZG7YKpPqtAuKtRGWw8aLz4dE563/2k12WP8Fh+mHcyyhdE5ySj6
Q5qjiA0uVML042pWBPb3EaqYlkU3Qekit6yPs7YbdEd/LEpIjJF2QJ/r12daLfAI
M8Rh/Zw5V2qE8Y3ZPI2TOCE+lMdE8z+hNOmatF0pispoosEwv1HDe3njNMzUEy1+
F2rAGSy+f2mWKuB8GO5XcuQJdCM27CZkcW7ncsdrdoN4UzGzmU4w0fuH8EFz4c2Y
G1xEKvmt7/7Uu5tAtV7MayjYgAb2yrroNmf3wry1sZ5M74VumK+ABKzo9KIOYP+N
s99JWQ1TABmIc406DJLmXPHCdEXyKe4QpFOBtvQfadM89RVfGyt8J+qVemPDVJpx
eTL+9u1M0Z6qg1/JscSh0Z5Gd/KlGrKCjcXZIdtA0x72xaaBc6Y78es/vcz8V0iO
pCkY8GYRK6a6htXVnVpQG+fgiSgjPTREEjfRPpKD7lNoRvTqzVcHCdOitV9ligqz
oKtu68RLzDt8cewtmNrFRRtVrS006/OwBwn5NXNwjgvQOiVM3rjEgyoVYG+e1tz+
ij/pSOUtt9GtS43qhMOIXTzpJ7ZOaF66sV67L5D5YmfhSWQRxp+CkQzuX5nwLL6S
cLNCJLcQhyer6C8E0aPdh1jQ5oAl48X0QKvUPi3l/bxpbiHFJ1/12fAdnfBLPpLf
dIZBhOw6UnfdiAP1Tc9gh1Ko1/j/e99U5hf56QDhpEUmxbSRyuBEBC40zZiNrJ6M
cI30fO1qlkwckDtWXDpeoDRxjUlpHwCr1YS7YqN1XLJMWZSSSNdfUAFPUZHPHM/N
115tN43fz621EVzqxfmyPX1R8Tn/n864GqtfLYnmiAQXXW/PXdHoI41+GJtjkxkc
IbfAVwcIarb3BEhuLoBb2yhvJjFETb/+dj+Gjdpf4N94mO5ABE62Kr5dFUqCakpK
8Kd8zMcik5lTnP/ooZZbMs2H50VOgPnIRMkgNZ2nkWThJjT0gaLNXajC/6dF+4Mp
sv23d7o16FnzYWnDg798g31mZ18HKCTQmaP0THtX89Ehu/7CGHhy2bFw1g7cU+Hn
+pCmCnBag3PTdPIiy9dIUz9Qg8paEjyIbbRRHBi/l7K3lbnRrPQ8h6RmXEQacHgw
gpBqgyxfLjmRnJ2ZZnmGVWpApI8jTf1DTcN3qw3FBz9ZOfjGK7sbkhMm02NyrNm+
chF0khn8hUkqtrWV8C2hZf9+/RDKKUhQWuASOWQw7k62fwuXxMss8p++j/WWEm73
XyNKvSnNhsEy/S55/2q1axElguIfT8PODTyCfVQ56fmQftq5db+o5xrBwJjtU8Fn
nDYbt3EfoThQqKE/DJ/4acisfxECSh0on55mkYkCS/zCsEJsCCYBdLDvvqtnx1nD
OmB/Gb8L//R4V4wbyI/IFCX5gRFun8/gT/47pyO0KmCFoPrQxHL9I/UIAcRh3dy8
To7IkIO6PhLiZtDklGyNMHECxBCq3X1HvyIzNP8z9z8vs64dMFBPTGG9VeC5IKhe
m2JL4p2IN380dMXILP57yXEbVfeRH4LvtGoTqFrKi5V5yTX0V8v8Nh5dPVuBH542
9o+mn48xyLmsxvyX4Y3f4v/2jeK+K8vzDvu+S8eqw49hf91LAYW8IpaQ6PbGasoQ
VCXRv76r674LqVjO23AdzVOe7evMOoSA+Y/2Or6UdSE6ko1hiS3GFdsYjyMZd3uF
A128Lrb3dsiC3F8f4PEIFanMVjAxSrzgRkdT2u2laW2HdjCOi7ICVtBkUg5akxbW
862gGsVwim2dxVCmdGkDDgEC7sCX8NiosqSaOlNYHqpSzq1zB/s12Kke6/Jk6QKz
0iIbHC/M0X+HlZRzbMKawtWbtTiHH+8ppRWaxZ/5NlTxnapb90IogSVAbmooNQFl
45Ak81RwzyU7wv/lQspzKlOC9Kr4xiAL2IQzDO2zl7PqBgbKLAa62IiasuEx67ZF
91JQSzb9efqPmlbVDA0Xtpz3Pqn9gLqS7+ru5G8/quP2OY3dI6dD15rxymEObRFe
6ctnD9TvG+mzOeHKm4qT8xaNjiCsRyiHgWCXHTzTnPaYiajgdUPB0YPch8ZWq+Sy
xIwg2OxWES+0yfNKJkbU3kX/7o8X/tp00iBAT5urE42ZL+oxapuEUgZe041XGpYe
2lD7RAJ70B4wwuvgae9/S832b+7v8RZhyPS2nc5yXVE9Ud5kjqK4qysnja7K1HhL
V9P5W/TZUK+XrKyCPB4wouicJlUsAcyRloYNs1Aw3G+NBPndQSU7p7iAf9CaVO5e
/Q/xvDMxyIa+EO0bVRppsxenNEaLmWeolwjvkL88oxpamFzm0XWNsYfgBbFyOeT0
2xhjJj8MscMGb6YLEC60VOFDkWml5LWaCvku4oFTGqPotEtpvmM5KDVHDvi7RiYz
YNCUIzv2dwLURf00D9doZaMfDFG+RpaBN+TnaHFNTVCVXRWZqVdEy7jW1kBQlpl0
YR4RxJ1X0LSLdOMGus5lFF0wLG5ihtm7hxxXq0fPcyTwxMwAjuOVPKRCTQdFJ6q4
eeBoGzyX+sR6DbrLvEanoLOk962IiPsU+bxPj/IzZyPEZv4gRkTlp6xhazBzAuH5
+n1QLUYoCf5gfqR2vvCCBZ2/fUQA1/FQbv4ZY+ShPmMtCGA1gUOFkFxx72/xKXnc
LL8hKGfejb6+izhAQZGslj6JA+Maf6kuVSpde+3JM9x7ADKwZNNOBV1tMAI+ivsd
PFqLmDiOuvRCYEBfZKEoQsVD/jTY0MaN2NVnO22DAHWRj+rIoXkzLMcYrz5PVVjO
pgCgmypI4H+MsFQBx1Jw6iE2XngMGJP8Gez7c2pM8TNwSyQKnkh0qKud478ZGHy7
4hP4Oeijsx9/kqmVNEpXOWibHoiOww/4wBaLzl7DdwDGcY6Br3kjIyxDDz0gzmvT
rahTDr4+sJOqyF1cSJr5dOlyTEiA8HONMco24eiUmoctSSEz2hBvmwldrWFsC8eS
pzS1A/HAZL6oqawjH4SL2Q+z5cvAyAUm2jn3wyYxbBtDUz39n4k4TJ1HTdsLF3E6
mwesOmE/FmvsqahBGMrsAA0cI7epSZwyjLh6x1BzgiA4BkXP1rc4/X/+oCM9MD/A
ChuRCWOLFx9KGcRaaprAKtLtDvLG2qdP6vbXdm8pUD5Gn/A3wXuV+UIZoDGopPb1
ayiWjUyJcxbp/GD4JcroSW+MTGRDAjiSi5AfbRhCWY6W88BOKFqmMHauR9mvxTXy
mRRnWbYbelHYRTd2MRgdcpteRXjQftdcaPZpDcMWrCpvGNqJrXPeDuLbhM8832MY
VgG1hhi8JiHSGpX/s/ajTrmE2YQvpFG2PuSP0wlqHGH3h8JlfoT3CvQ5+MUPMb3O
OeAv1m5SGkyStbDOmcYR2heBJWEeS/rg32PfoT9nKGY+Fug2e7rcUKtAdEvOn3At
O0JTM275CaEEki1/mQIqwQXGK/lkGg6BvFSm+p24kyIsiT347aQTAgdCxCgDY+s3
lUeVBxcPxDUXL/2AlS2HERE0DdoTJBW3Qv4w++Umw9VO39vN82xFVJA+EvqlHzRF
7CbtB3hKeLNnP1172RVerGEkUHiYs/5uQCGVKEOsJUXnzXSNQM5k47EceWjQvFlR
BksDzJqe8ag9f9h7oT4ZAAFhDG4NJoe4nZfUzF72V8zlDQKHi1Y4vO7oRkJmuuAC
WA4GYSZ7u1KdCc4XUzSdqgiUN2ntgsuIw10SuD3jCbrki0yotvdbvz4jWomwBH7h
D0PSOH9ImkWGeMpvzaJBBtL80AQ/1G0yqkMzycX+Meg+thtVCZMvzIv+7Q6a5ald
GZtfaQyEG1LhdFVpH9RNsNYyFDvwC2ZfrHJnuNyRsK5XW3X50u+xY10cbDdI9j1x
i5JzjMg8DSzVKO8HhyU8TJ+6dW+lJSDgDVJ4dslkz+fhFDT/puSTiik7xpwkUoNQ
sFy5IuA94tShmxXpOnamr0z7yim6k6LyOWYqmwkO90g6Swa/8HSImv0QVGzrxHbJ
hCwXAq1JWhQpER3/9EGRh1Nm1Xz0XmeVbqkG8cl+5BGCaKcI1qnHA6VwdECDPCVz
3KAr4O9eWxDJa/zqtmQhwE2yCyVS2FGZP0CzIyvRY5N4lkKZ7Bv5oTIFFKPaCoK+
bKVzbXF0JEPCgwLBKztwf6+M8YK1mmokxnAQsLDMPHqt2A4as/9vYZ2qu4rY1TUn
Np1uSHzt6nOzgdxOwXPbrAX/2g+Wn2/pC7LYMoJAId3kFx4VJ2cAdA60uGOFcf76
8B73Yr7skmoZmDWp0hekAengxJl6T4rYYz4Ni7n/FEIFP8iRuDHd2uVo4VsIo845
tOwWfdCNtvBE4dMAk/xtTBZSvdcguBigHJ0hlk57nCX9kmJH0tM+OePozIGmV6uE
cKamVh43NbR0Zr9IC2o4z9prroFP9o7BAnWnuNN8LT1rETvj90IvdqxvLj2PFemR
Nb5M0COaIaIlDqD71Dx4YwtvajkEwPeCXJFc6WCedbCj+EnIN5BORdDr6J5pHYh/
6NsH2zwMsKV2xK3BnRjcoDsgnfndPanrcg0PETMcX5ZO4uRtW5erJ8yNptYzBfr3
bwviI+qNz89e6AZeXucxftrv2WZubywOAFz6qm6xDQZRJYl9fOl0HJDvlu0ORbpc
Iu46BUc36+c/hZtrkcaBHzidsl1NRtmZgl5dyslNuzpdb3QGQSnZNxq6pOzch98F
zBwinYOOXoTzgh9uwCwp3qj/OZtZdQR+NXOcsfnBRO6nWME9JzP74uCvjA80bgiI
bLkY4AgRatHGr9dyQkwYKINXbG0K20Po9pGB2uByUeDeFBT11fiv/JtJMSk0qVsT
x7tCbFR6f+m6YFw5bXWBTRwB7o4ZYEhHfcZRzXDrpXGthz+Z2LMtrLIMvJ9xoBGP
X3kMKui/Lb8PtO7GQbC8YfXDNB92Q44Ea9KAk/VVr+5tZUDG+khLhlbBreqrRkFK
M4zZuKZ/Zu2PpTplkRlrv7EbYh35y4voL3CkRhXdnQG5Hp+HIASC1KSur2VjDj0x
3pR0HoriAQkJjoYuvhl+yvouhE+AStlMVwVnOXCpe15LV+B2FSESK8Y9517Ci5Mt
okW+kPoZwMYrhj/sP5dUqT0XPDS6x6rIyv/Q8ZHFTNTd7kj8p5CDHdWNZyy5TWGB
K7mSrmMcHuJJ0WZ4PJWFJ6kOneWCtD+D8sewmbQOcg0f0UgoYqC/b1mNjQS9qMDO
dZjXEV3tT7loqdEveS5oUt6aFGDOivdlkYHkj2UQun1GBoxTv6ghC+vrdAVQ24vU
roiGKJgNBmmTbGOSIIAxWM0s+T7OHyaZ93VliZoGz/2ea97zulLcQGSAbZDmw8pw
n0oQUt1wfHvQtdju8zIJ1AhEE5zIMLmmfQqJfrqGwqsNNwsyTw5IdQZ8IJE+5U1d
pwWNWHqqxrIQ9EFBV8X7ypkzT3RXu5uPBrcuIKAq2QjuZCwUHqdtu1PTIt+muKFl
oMQn+ZF3VZRDb1p64/T+2cK/8jSR651AAHvlc4sZMNmzsv28JXP8rHv1Z69MOlwK
Io4Oy/1nIn3uMijjc/K4BPD66tNtVXrl5pSvYmno2bUsk4L3c9ivahE0JJWXYWPF
dH+ndJkrIJy1eEsfZJFqYQE5SNYjeSSf0EfxJR/d6DN4c5mdHrsZWT6Je6UpugHT
BJHPw9dgPBXJEcyRd6b6cYpEFEg9Q0RXsohqG0OW+JOXJn3Du31stkoHccV/LG2c
3SAmrzVtCT005glOIg7ENWdR0PB4jm7UyT4zexTPUD+p9bcFFvPldK8VXZKSRbAi
jj4wnRAj+MhTe1XrYgJmhz6/pcrl9JoE1+V1qETCTVKMxKs84GHLOJ4RjFSKeDoP
ygWMCCvuuGYxpEWFGMocHbBRuUAci3zF8EdEAQ6x2EKcQqiYtMzBfC8Ad6TfObnt
SO9KXb5yrVjyrAvYDkpg64nVa709JhUlrXMb3siPhNRYSEdQC0xJ6QZ9MzO9ZO27
Nh5IAszWWrLn332bR8CbPZrjigJwVQmW2Dw4ihA6wiR5MhKyubvhhs4RL+R/W1Ph
B4Lfj7tKQphuiVuLrl4s9fe5QAT3XNZROi3kRPCSDkUdN1ByVG2P4baK/CuQ9o4/
TCKXvbpyADnFiCqr1B0+8Dui01jQNjFkDtsPcfsgeoqlBFxEFOW08bYj54kMkCX+
5VDI7ou8rpHNwf1K9y99HsvuA9TKRZAravoWDiCG0sG5RODoOZVRR+9rxXPilx0P
nSrb4kFFczVBUmPIfzBMF+CzQL5719z6FWSrOhftJo2Fx8LvtkIpF9Bpr5NoHvzy
EepMgMmTo0l8nBEaGdoqbPfkvZBgZhIT5ennyYL4XTWizL5glAJpufzWp5whizLR
PwVGapGFGfxs6NqHm3DF+3udIVF9TfrCI0e9xBHmuQRuP/eJK1LO9cJ1AaUImz0Z
DDg5vh7w0J6Get/DfH3vtAOqzsvdsAA+d2NG3vsYuWETi+cym2Fc9T9l17uKNXW1
ocB9kI7wNbUVK7P7vU7pqzTXhN+a65EaMoF4rQPHGRX04VDKTw/zkq5tDNglpt0k
LaUouYRWvxC1RrY03oyje5oR5SCxe13knSWxUpo4n6UOqrRxygShIWYNY2+ytxtA
H8n9C+UgPq1ChROqgSaDxlWJntVJUMI/JI60fGlzAozuzzNPAY25vtgc0zS541QS
deuo385VJwHlQZIWygjBedlZjngyGYTmwbGwJQL/zfAllcYHEGPi4SvqfQ1GltFd
nhttYduY72etTuBmUXqDEmqZh4yxg3cJLttUy/43DoJzGSC73CDU69e3mhau6EkB
3Ya7FenInTu1v2wJTZaNYReW735gx5TdZdo147F3UP6HsOKEwU2jN01nIs9hmaOQ
77fB0khAQ7f1Z2jubYCpF3pRGDGjnduYdLl0ixzOQicVHgZZbYALKU4LBiDyNViO
z/oh3uNEbZE3adILOz+xzI2ia4YQeatgynOKWcQZxLzIKeGbiMG7kEYJ4PDyIMxn
5L0KkNlg7QtOy+L03eIbcd7tfbCjn8WWFyGo8z+pIqcmJMJsGf4JxwazCJkA/xB2
E41B6YUTJQ4GpiiYUPnqPepe2sO9ApyLQr+XTjEKPqaWLwUCB3Aa3XY+oj9GMPFa
/aVguR6qnkN4kj6+fr7tIOR3i+3rlPZCo9FLWzN7LFeSMhMdDxMbFYJVcSzxFQT1
s3iZlkoioTidgF+R+++SaX95rZeLkvC1HpGIy7c07k1BHSH98qgVX2I0PsitYUzR
5XLYffz36mny4VDJSSeuIkV9KxpR/4sad0noE7smcS7rQ4EAlulYoZXZUF2wKpNF
O2zCE2eX5KQkMIKEk3KRu0xHjS9yvV+1QJGm7IHIK2VpqxvDkmCTJe+2IN3XJR8u
VQT+kzbjE4nznEuKOAv2iIpRFfdxrOE9ZJC1S3FJ1ZInjGXpmyVQMokXYO2ev0Xk
qp+0h37gbaanFf10nPZnS9dvcf1E0sVcU79FpQr6Za6v4a/kSjhQcnVcwEGTL5et
ugbIX8c2ty24yiXo7ba8LzDypZpCXMXXChAPuYWixVGLtkgShC0wPyCy2XHU3kdr
mxebIQ0e3AcbZesaLVQpjxvohdWlJ+QopgsyIy7uv4z9yKDkO276cYRf9TxqqWz7
QYYoduoEd7UBofpQlkr11A6PSNhO33lI1W49DH1IO5we4V/kdypfl36HLhXNFJXb
GotU+vPjpG3URiyLt5kI6W5eAcUeO9bF2KQIndy9IOYRq5NhNGiI65Ej28C89fFH
ReFIInb2mhJCQldkCxyu9BWrC//EHkqjuaIK/T6f4duAMi6eW5/GYNPpKPgyEBwM
p0rmigLweW5LB8wM4QHSCE+xweWkCup5qPilhXjtvrhZX1+ugws+aeeu3gQhebv2
Kxl/nO1vo6ckHWJ3ThHvzkZZ7NriYjfIoyxx+09Wsp6ZW4629mlE6cPISMvmsret
xxIFmKZcCwa0OfIbn02eAYhix5Hu9bLWAyN2C6QSlJhUrnbe13vr1ldUvcnXTk/s
/vhinYk7zC5TagaxDMq/7oUHqoDa/wWqx8m2BOe8tk74NIZQPJvYJhJPfLAkxG13
61MpwCfJ/iRwAHI01QbyfZ04S2MvGpJPzRy4odCKeBHUJZdKbPrlLB1Y5AWK1gd6
Clm/9CgNOdLafE/DLw3dmlUCPTwra/C5sbraS6tRNDXBgAh/m2iqGMStgr39odQM
C1x18C4yaob7iSg14KLglg3N/ducq9j/fAYVNX/q24xKvmc9N8jOVA2+EeQ4dZg4
KppFDNf8UAN1NsEy4HdCor5YHtpSIcwaCcJG6B/4m6/UsDQS9tKR+pmymOqwqHfd
DNxijOUpeciN4gM8xOV0M6epzk/b1VSEcshPoHpxHOgXXj5SBYsAunMLdSD3zDAA
CbHWF58tge0+tk81TyIe1syVx08AGkn4QKW5BmnWgJEC+LEnRYZ1X2JIUIGEbakI
hRZEOWqJcoxeUHFQVXVOZHcpJ2dNgt8brAVBC8b4mR7JUR7SQqI98dZeV/iqInkV
xS0IY/EUkK0OBtJgppkCfiRedSvmN2swpd8YyHKc5gQlB/0pN8Ww3bctKFYxXHe1
4DZJc5D+raWjxpNmsJiRi0AADzNMv5EkbookVjNUR1z8wo2zRM9RJcxshccop5Sb
W4Alg14lVKKUg6cIMcC6m98sL6XUMPHvQPeWwQ2uzW/skqk/Vt1+uLxqVksGccVM
3y4sFmEA/mCXi5tkfKUifmSl6F4DAbYS8sBJcbEo8H8DM6A6y/gXl7k+i1BU+FbW
lm6uasju+O41RpXIk8489JFAPXKn8Z0ISS+KmkZTil3pJ0JZWfajp5yHVErmmcHK
oNeyNxYG39zN3EvN4F/t8B8BTedlb/+5msyTKDbEoteZTbKykUpobJZozK6UfMxO
RKnoxols2dcPz5eutkTpT88bchqxoumj9+x8U35+J/KOAlD4YWFy7XFvJTn11HUk
MjIP5TEwcanimtGiRtysVTiI2dQiZUOdp9XtgXV7LTugSNspM0zI8TUJlfYaBhDb
eRg6FtZ8Ju8Mb67g9rm2Yo3evMMpK6aqZHOCGtxI9oGWrQ32GUIPUVNMp7eOhxa1
OHa6JtxsOdLHfLxGp4yCj5ZViL4FAxebBOO61i8g+ENM27YyLNmx59aui72KeV57
VQJV2E5rIFWReF7zNKvILB3dOeHpTNOUWL2Ulv5Vv7sZOUKhCCrnDDSfwxyugINy
Ta9wN7SFvMF4xKKuZBzQMuFwizkWPdle1QZVZb4KdliAJbwy8ayb5FBcft5KAUwe
Q4AZfVF4YbOJUTXnIjhbtDK9MeSnXgC896SEhbdkPXapIHzX49UxDn1lG/1qTH7j
IPySKK2IKBzvc+5/2CHsZEM/Bsrh+nM+D9ncxIMhPU4sEM4PggKjUGyCeYhp36AL
0Qp+hCdl1X8JvL1/Ws9xynsDFLvmOMlU54clpGCPb5Qmq6MqPumlCbHA44T5fpy2
QJW0BnQsEONHnfvy7c7/lymekUO6Tri0TeqH4zIv1mTqP9aN2mRbNUAI3yRzYG8p
2/ubjSN6t7iuwlMUwoISmOQg8K13vseZOKPO9Dk2FxQIwRsJfV5dg+TGk8KYuW5k
VsB9VUuQxfRxNyl30f1925wq52jP1NpfoQgIxU2OeCMzwZgWC114EV7MGJqhP2IX
4c3CKjCRPe5nYhPo8mNEemMwXoZb5iUi6b9cLubKp8rNNqW9M5J6hFNKqn/nQOJi
pytAT46LV1Fw6yrtEXpBxeV7ecf3qwiq2+03dAeUlI70R5OxlfWgLu7Q400ZErb3
8AEDBR58sQzINpsuxLkeuMloTJXxV/USzA0mrXNDOsgSpDLy1mHLEGYQa1Aae2Qk
4MpNdtN86Ybz4vlcQiKtWGGkPTDazkm27j5dj12eO7/MzPT+MdCfSd7OQEpqJ7J2
dXktY30G0PpjczowoYw6Yjdy67XkGcZOHaS0ORHJmuuBbW7XDfY+oRVMWBwD/P0r
h8Pr9Jz6vPa34lqFrIBXrS1EwqCo0dmONLHuInpGH/Jwrg/HOy72DHC+9jjHRXAd
6HEGMaYIuAlpduHj7znzPjNeJbRjSL738xUyLP1IvjGCXQGEwafMZrJCHog8NlIS
gLSRqD+JWH+0y/bPDtfFSoP2D/QKHi/TdrXWzjOdE/6AYUucGx4ckN8MYOPhSNhD
2q8TQQp7fBQxP0+SM+sVW1LxL8fzrq/se1mFMzAt79qmabZpesrGWLdEAbO5nfPX
2Zb60aYXYQVS2Treln+fM7OzQc2BbjRXVPYP2eeRfsO4k5asT0FNqSzO7ZzwU9Kp
4Yqn3QwfgblvHLX1SmGK3/4Gg9H+7ZQ4paEldLgo3ETWP9YILAvIp3+ELjv8EAWh
LXHGqpwMRKgvMN5Ro5KfAJdY2zekBIUovRY5xhr3fZqUbzcKXXUzAITD9a6tqU7S
ZqRO1F0sJvvE5W3hpIT7A1iAOTSvF5rey1fMsmY6vh3d6xOl1LiKjZf+NplwqFyl
yqBuq8iRZpya8ekKOg2oySMXCU400NArqz1eCUvVHGNAeLpU2zwRJXeuao8zIEYc
g/G4bKIPpiWvH4uIdyFA0YtOnmEoCYxSAw/TeTohYxQlzi/qk0LKxnoppdFv1ji5
W3a3/rQVsc40ouqabiEQmMq8NIOyrvqmVVOMwZxYrYUdY1u7X/4y3XH1GgqS6qwX
hRXe+06gR2YxWHiVgEoSjKP0XWi5ZQ/7ku9UZnH1cDZ2TlWiFWQunoUkeBQTxc+a
Q67ZdImccphcy6E6lG58oDpOVL5KBZeQkIhwciQ48m/TCzkhmX9WQ0x92ZTHXqZq
vTLcQ7nSQ4gzBNT7vuGGjR8TSyWnASigoCsH2xRpXIGNc7meWy8REskCd5BW5O3e
sIi2qi3S0UZ6yWJdUr1Ujwc1Tsf0ZZhlV3WkV1HInJQiOT5IyPrRFyC8jd6w1Jck
8AdcquS3i1mfVi6ThSl/6iTMwv0GyA+N0PDMuB4JudS989gnzZEZ8SnTukWevBB9
xD/WDUHXT+lo3rI8E9DWY0JYO93qWO+4f9xF4tll41qPhDmQOq4aOiKoFL/yfsWb
xdNc+twqVTmXOtTR38COTPPXWhV0V88ZwpWE9XZsmeksLdplGYs00W4w5N2ECKlI
i216dBl/EeeiI3U66RicilBIJbgD0aNf7jKGnyB+Bl3B2GF7eW6QI8Jsewb6+4Ef
gn7Uw4P6xiq6UdathKBJi5u/USYYyF4+4ut6w3ekECWwOqw73yk/ZovvXFMLnLlV
VIA5gOclSkOxkYn8pePFy22gMXqimHnN3yrWKRdUXQJDHeM3MWcQHy9xXK5n4uQI
MkPbZSQ7atrvITuUC5p37i4itpSDyC3B5p2elArCTjs3Qo5FFzdexfux9MukAuIk
FCGQhHtjJ7xMG9vUw2c0LhJ36J1E6L85NE7gYw+VgHZvqK/L3soH7RGJCB42Z4ou
DAB0YedkZCXkpQrVzz4T/dKWX36xB7IoCy9XTEOLpTglKHYSJoeD5qClEhTP/w/z
iwFMXRzbqlR7h11qUZUc71A9H1aYu2YAD8G+w64Aub542mQ18jJUoG4kbG7pnOk9
IqaVYvFSFVjfLZu0sva1r6c3PauJ1iJcUORqlb826FlXGqmGogvknmZ+zs30adGY
bf20bFWmZdSFWXekg3ZAj2tgCsfRfL9J1D9wTEOKtY0jMLr4Du/oaY6fChGHMuZE
42owo7M6AJWn8S/JFh7uHNbmymYimYrg3QTECeXcyd2131Ro3zN8hhaJImm6QWVN
BPBCOCc68ooMKuJPMV/o2+tRIvw9upslyNIyM8F5KWttR64ZfER8ptUqAWyaxSgM
2NB6V7LrjYwMLECw8KOHQ+UOZ5pzptAnVRfIAv+sNGaGgYogqp2TJY1/qPPLro+z
c857ohBOBghYj/wyRBUFSEJLuoCrl4oGv46dfn/NebfjlV8cWbv4Fz8pQvIgOvuN
GITmCK1PUC4QyV3NBBJWIbYZV2kub92yXUTyFKJXGWj3l8zSbJZuVDFX7Ymy1ADC
rSH9Q7FqfaIr6VvfTAoCZjMK4g02RCU10DPs6cMVVL+dUcuCU0uqQnhPxC+d/FIG
WhMOw4TAiKUlAh3E06uEgRJr05DjWbqwlG9iqJ97H7bdRicITCGdijE/UDm/HoDf
LcJjVWN3o6JwBKrQa+v23QodYR7DtFQ1rCBFWp2dMinWw3ClXK+J/JzQEzXLwpnL
w15wP1lFkhQ+6H4F5MptE8t7qqDSKH3uvSJwS14PIcoG4J9eg7ULUi7DeGhHzU9X
IYLFmDh8zMVO/a1wMj6N6ly06L7JCD4hsKePfvH9YM+OpgvD3Uzvgj7eE8JDGfW+
AJtpRAEDvuPtKFWbIv4q4QcSmOmGF7IAT1mADSVqd6O/IP10rKkq6OpLvZKfUh1G
cLZ4wHWWBZGP7eWGorv5q4DdRYWZmZIynWj4icurVBIXu9Je3iHu4q20Ila6pet5
jQlTsZ25Z2f/Xam7ml4IreVL3HbX5S6zg2ya/HtrqMx2+Xj6hL+Yn7Td8PF1Eq0H
4KRC5C/d+D7817GVrY3qET+fT2BW/2VnKVjnb9b1CLCQwp0fbsi0M+XWthoVjW2c
PR1Q1AVcw3IdFVp01q3YbIpnf2nzd6M3EuAtSNNpiQ2efGd3jajklWMtjJs+eCWH
deTNE/11qlWkyxLdM2a7xkCj3IeQWChBWRv8EtqJSOwG8Yd+zsLNClp6hA+P0BaB
dH8LroTCRYwY6ZYZfhUDBC9EGzc0vHTcSrX6cjgHw3GtxSYIFjms+NBcuquG6HT6
q4e3Wp3n66SQX+Umza1UNyBK2agP/M88jCtfGbO8o3Z+wv1g2NmjzjW/qKTrvue5
aygwxaXGwTEOXaJMR831ZZB/Sk3jUn72XgyH44uIGy7WcpBJuizbl9zzQBMw9M1u
jl434Et+9McEUpg/DonjyEdUINecwhrChDPOHKLEfP/DC9AMlxMg4T1WRPhaKWkf
MtvT1zOlVy7sLyI2FygcB8zq1r3Dm/H2W/rLZa8sH6OoIHgU8zO2EplSo17ZNiKc
ezBZl3X5Jnl63YINJePXF37zUZLmSOyukIxQ6sb1tSjFO5W3dm6ZKkCSgIunH55l
dqnzidybyelwAy9RKxdu4nDQ7+wyMl9wen5QCE56g86QwEKez342qtk4wfIiqKdL
GJTD3SgrPNEQgZSjq+fOIOePogd7uoHW95niRgfZJge/FinSH6J9JTfu33tS7/pr
6yE2Vk01W7h38FlpwbMjvpB6BSId5/owLkf6zW7PcG88CNfY9NYl1pVKjnFL7XzV
KJlUa36u3aVMX80P6FabD8T9ctmbM8oPW1yngf0J2rgbKSQisVbZKvvrCqRannyn
HQveS/EFpXNtTm0pvFt/rl7Kuu4LB9GDMn2EZ2obcUvcmmzm+CMTcguyA0sU/LWz
RsRPqYm6O6haghrLMPnBE8huYO/6mcpYlvY39Le8CRJ4Fo8A6UkZNY1vnE1GWWrA
8N18F/Tf63DAEQj1jxbHBG0pIlCYh90Ojn2th8L5Hai38Z5EuxPsoC/XIeLn5WCS
Id1IQTbL8NHp7twg1HMOhqqtXn5BedSsMLjOyKZBBdeK0zEyD5wHTss7idgZ1SDh
lcxXHZo9UUrouj324FaxNPR4sqwK5O8SYKWOPm6FiyczTRrpA1LTQMEKGFM2LF66
twZdPwkbLF3quhKKcrZLbWldjctSJz/jhAXLsfsVN8P12mUZV8dujzb6HzwlTBfI
2RDZyhLZsVjLZwfyAy6Dqla4DIpt9ddncWVS2YX+FRjPwTVbfPyL1ogu8PWb1pbu
1cb4s2q9BCiIUKv4J1geKeB9gX1fcZZxDxdwN2rsS8w4HVJMbN4miFTmi3E3dZH5
dlIaU+UdPyto/h46zaVuX9XXU0k/jjrt9tuKh/yVv8iu6Yh5tKEdPq92fd6T/Vth
abKNLN81tDy6r7lPs86aZ7R7BwlnZ0H7a6clwqVu+TpuEx6+dgN87K6poOLRd2z/
d6tAbnOMzlLif8DyG6LxjsbTgKcVzIsLmdGNb4jbCqTiCWEK6IW8lro0qcZfWUSS
8QRXyttK22HQUwsOXbDJb5I2H6iycjp39NL5RJo5fyOF05z7P/furK+qCMfoMn7W
UeYF+3+KMtNuKAwtO5y3Mlvwg1fs3x87E9yjFiMsWTWTf+uuhyqKY3+iwpcr8QvF
upPLP1+CrXiM/iKbp4YCDhzp8HKKlvTv6asAn18VubAuNi6jBNndYNnPUcbIgpHZ
/TzwLTjyR6y1ERfYhF0TcRiNM+lIZCZnC4cbKyKWaEhDqG08O56q3IGhtrUCuuVV
WLHL0f4h2TlPpOqc39YMqfZl6uQPfE0jby3XJUPan/BaRQNBsD/otZtX1VYqH/zR
F7YinvMd6WoHsrghrIswgaKt+wHToVUYHUQ4ZWsoPg+3amUw6FeIo2960p+YHoTH
E0/G9HI5+J9AIhMhvITva/3sKhtPda4pXQdXg4XErBysVFRRntCRbr0V4Kupx33u
cVnzhRmhZBX0D3Lbq69zab9TnfbDGvPHO0mySKFJGCdGCPnG47mhti/z5SJ6v5Xb
ijyacpExflDDyBYyPX3zWVk+FQUHKZ9ZPjuFnZtYoJ7FkwjBODfvOng/iM4U0RN5
gJ+eSeJfQ6Wsg9HdXg1jaAhq4vQjLOlbizaGJLc0obegVmYV5gglPi0fX5dbQ1Fv
QZgw/X62rWJ3kVzJhvD7qk2sOlnw5NpqowV20mLX83VzRum3P1RtUtA8AJBd5L79
NLJ0JCvtYDgm7vm8TJOur7dNyp9mpyKTP5GugwMxo0Zcnkb0YFAuHK3R7bUV2VRZ
0PCUTCCtLn+cu04xo3RJdzzIDZn4eqHb9joPd/heKW5/JhKM/gNFVIlKaJe7zPH1
PEecbFUWO5Z8JTOIGTvH+bR0TlWmyOEGsCN3DvCpz63W8BC0M/QUgzVl5Qg5dprr
UnPf6LOYQSXcydJ77B/bUvOv+nDmn/n5TMhvjaOvqgN/Oe8Znm0jyF4s1XMucU35
tJQbFHTO7CNZKS4tsNyu9sXfPerke3+UvnreKNKqR4LGBu5WqpkCG3yEoKoS86xF
5wEccpi9Utz29h/nIcyT40BkQ0YQBuBWORTfot+jVOYnBw/hTMdS98o6eviwzan/
SqYxSUPvz7PsM1uXeyFqE2iSDDtDFX1Z30UHCeOUOJNwSr6hgDfjv58FK4NkMYYF
h+CJ7e6tmX5kRB9f6Cy0lpOTVwf9oH1TWw8/2C1PcMYO2V+h9aW9gpooRSkK7pIy
kAuCmNb141OYlphVCtOHWcw3rEswX67L3DUEKG6VfcaYOKb5om9T1Suvcvqy9MRm
aYZJo1b1+IkmIFX9+kHeXOyC/9KQw3T/aicaVCnqaVeTUzivhHfg3pRX+STG9zzM
OJYYnY4mJeaFr+OD8KOEOEgosgC1W9rPfq7vNR9eipocAcHZCV9WjIazZ4XTiv4X
OQURApNfRfkG2wS8zIVpedilwrXPZn+v3PispbZkNrvDbkYeRWoUQ5i12Jxc3S2H
jeYitN94QJ/PTyg87rhwoyF8lrFZIUaQPhpvnGobW3Ifw/MmoB08DbYdhyhE+Tsz
tubAJyQMMBFYcnCI++WzsmC3MOnjFgj8sSRB4XA8yHzuM3iRAl+UkgRUwRl/IEcj
mIz3i1UhOVrVmKUan6iHteJflU1PIERdSdCx5Nyj/xNcLMrXPBzXpJvusjGmtu34
FE9lfxAUF9aeq52s9f6OY3QuUSxMbVbULc3V+hEedfRirlZfx6vQdqnD72ObmxEG
kfTlIYpA2Cios4DaRaeWKImOZVHnZN8SiteQXXMJULHiCS7PeO1fauTmh+uVu5oM
9Z1Kv4jJp0XyW7l31JeFr7UbASHU8aHEE/0kBQq7n7M+pyY3hScRA1i+QV+1lY2Z
ozGRgJYGpARc9iAIA1apK6r9PLBoDxIKvzeB5H9hm7xdFgIW+uC2zIQv5GKOgoWP
khrbAo3kpeK/3XNiswWnRCNGYM2hgw6EZRj6gUvlDPcwL9GLrLg0pZThRoi80HLh
0G/c8crbpU0XmKX3xtfUv5Qp1nzqchoWF/cHRnCKbkQftm+dyYprajm6vdRDoook
vDBUrE96INYZ4A8tLKuqJUSjhIPUfaFW1d/Gh8lq6ArY0XMiGELSXgBUfmVu/ZjA
fUysbA5HfNcH9WIPV+EVbYdi2pE13mYtSiSmhG5jydV/CZI07/1D9lhcCgO+A65x
GlDcmTzTrUi+XvHIHUEpdF9JGcHKTECfunWwpcDKUty7KFnWZrLQyf6jbl0wp3yd
n1T/uKmLTLTLplHJymcflKQAwPkxjPY+EpIPKAzVatxDBaB/qedqMMGjgHBzERgW
furGevR1OaOlnbRwIhV3Xqz+39kwGFqHwfzX+7thTXML3TlR9/zwj5ypdJrwsq2Q
UIEgaeb/BK+1qCiBf62eDfw5EMILQ3+jy+eYFpvLEzXxKpeiTJXMOcgzfUllC8km
mRrYbfel1hhp1ezXWs4siphtVsjKe3IZCIYg33gM3qo/YTA340cBr+5hji4oHpGi
X3vLkHu6Pcd3ElB5SCjYCzv0mU86WsJPtDa4KcqelESGHy8bfaN47jyXe6N3olkS
ZQK0f3cfOJCRPZGtTTjsYhvozIKa4sSK0Ulgm7gCf9r17+lemBwgpQ7e9lvH1AbU
K0798YSsMPFgWGqS+8BjNpIjjjWs3teY9FUCsKW7QXvyI1PHmj9xdz7uO1Fc3Rch
EQgSWQtEZmyBUV2esW3NS7ygBqXx9f+Bk5I55Uhsp8MY0b1cvbsUWwHS3s1b/2WZ
2zt9R3lFiiv3SgcV1jTlqx5uNLZmUAOS4uAEl/sJIpPzvCqTLvxr4mEtJeHk+W+8
KQOTOawgkgIriLlQHKt6ueQg9Uw/x2NwekTGdgLd/dcqwLHJrxEkt5ZY6ejV2W3b
EpUgPrUWuWIJZ/fQIuS0qzBrlJqwwgkRTW3BpBDkcQKQOXWYg8GG0uCsxtjenJTY
OUL5j81CAlfYrM45QhIPBOTP+D65PlNUnV6e4HMeEFTxnDc15P+qq2r6ty7UyDb9
wkN49Cf921jv7JNHzjdc4k/1YHFWzQGbUvgS8ga2qsL5S0EFrn5Mb0zt21oaNW9d
Lpq44nL4RFXjw0mDh6PHZ1Mpnx6bDAs/ddU7ASU5ADSqFCL90cV4rnvgKwn/5Mx4
cgXNZnxlPrK7PIy5LZjxxkiT47Dz5+Wd6FVWqSL61QtPxAiItKn2oZyh92KZlOMD
0HM+25n43mACfmkRbeErBOcQO89CZwrlnnMAHg7Z5hlP8bHVmrAKxkHYNC52KWD9
GylAHf5kst82D4OYwJq0TsPHfpPLLioZQCJUCfxnQ8KUayXX4QOh6PN6rpWJDw5I
a7IPC6qUDXTOmJORYfzqis/4c1d8QBCzDNW4g+d4Fv8TCxqLUFPwvFj9ucRLzm5H
pyJbdGSdak74ywVgnkP1E7sJ4sdpCTSKvhEOUq/Hxv21RZLt5BuG9C38vVYaAmcR
e24VWMJkZEGS/erZ7RlEui+9rt5hLAe/v15SsjPe1ENCcZZpjLaw0XKkNWjZ+ZRi
Vrpr5REZ5KBOe8ibnr3HHZirBCe64ZSwJ4lNqSZnIK5UmwZhIKU+Tq3ydTPK/RPO
E2KY7pQG3dE3rcliSMBeCm2B1hG6sxsvkeNboGIHUiu78Rc4Rt/0pwlga7or1n1u
aEXYRdh/R8icaTOBh1j3Xk9p/wSZPWEAf2S1a9G2kSy+C8y6lWJjE7MV6NvMOLmJ
TdVeyQWEDZawKGb7v+HZVvh6o0uNaG3T3SMPMjDlOwyff1gD01N0bdO+mFqk8Gb0
c6fFMMM7JRbiFM31fdsp9DlfRqueE6G5Z9d41maGGma1VklHCCvzWYTK2pIf+7gt
kP5HsF27OUlCDkhyaHHw4QLt+TIgW/2hWiY03Epi46E6yrxsAnI8UF4lX/mixV08
XqTnQUYWHObEu5+92c5DpZEh2danyp6UzyT4eTkK05Edkbdc/VV20bxoW/FeC1AB
ciEZbGxn0D1fqW4F+q6WR8ZGXBRhp47ZAwSOKapR0AHQT0R1zyKfSgNznOOxHhbF
9Mfs8uU0+iwPuuIgcHiT+usJVKfy9USpE0FBOHo6CDYL0OmVMirz1B7Xp21MuQPV
VZ1KR1ibXoXaeAsEsp/nn8NDNYQ9w8w2M5lq7AZdw0NY22Zk39Y/z3DicomM6fl4
vpX8XuHgNYQI12WA5vW6Pd6o8aLNSlrE3AzzM3O6Q3sfu1wvhYVSWmghXt/Qsl7o
ZLFZZpjHWlGUGnQf+Ks74TJXK+1SZKICCByh1dVBdjBJe2yn6hXhTMt5OFX90uml
YD1zg+ksPJYdAsWk9Zt6+wak3tJXDMndDECwQIBl/OPPy/mqGxiKaLsnii+lD+kV
M5SF/gq0hn/Qjy69ZPsU2z7Qm2pnfcjI+nIY3IrQUXIXgXE7wow/uHWP8/KVPdfF
W4E10SQEoYs0D+rP3jbO5W19b+UULSQIwDYE+UXmEH0fIboSczefmb8kPhiWIiGM
FW4XSuhMDU37bWAxvWWEH7ItFgBKT3Y6D6XAiJCAK6Ii1n6Kx+MmpYf3XxUe2q+C
4UgbudjkoyP8xPDxo45BnT4PipC7E4b8vpcwMrOpaY6SqPXYToLZQUqQGk3ymdKS
8/0mmjXJODJWyE/JZeNTJ5uKrr2Dx+USnTrPdsRMXYFDiZeIydZbZLkhoHEch307
Unkbsfpv4oErhx/i5euRhYaW/SwIbt61qOzmjkz3n0ND9xCUNhksRxu0BY5IML3V
tFVPbETqL9b3S8ltaZ+bUFnlkb50pseLI7FHi/bGmYGg721KZo+kcZQa2bg+Q9TT
c8j/28lN/gSOUNaHAHD0RkWMihWoOpZOEEvwXjQs9qDeXH4Tl01aMtuxdTNHLUbw
2c64mPGx9xYbG1VxK8HxMLc8rXX0ShXU7h45PwrO1RqyzP5FMDXbC2qFg1R5DiH4
BUVdcVPjJXDRgvJtXMFTKO6YtEVXr23UKctDElbayYEk4RkhKIQT8c3Z17Wp3sU2
7Ih8WWbSHifksR3TrT42c6THFVM+O5uvWmNecq0QSPoXPaIw4+Ji1vzLphlSuoOo
Hi1weiSw8eDvAIT+MbN429OF1TUNJSnDykMCY2gis+TZphzqK6LJszGjcWD6ifV0
LK2lR/JHOE+HWWC85UD5bBIorMbxG8VKx+JutF9bdkrBUoFlRW+ExkY2U8Pp2FsC
VqAp7IkF/dx29tndZxYLJJaez4mY50fJywPPh+hqOReeWjYvnTFHorVM4YMKhjdH
m4ta5BSFyKNTXLD7x2L12FCIXUnFmeKhHswtq3vGn4C7OwuaeHPS50wujYTtel+o
zjr9UJOCXxaF1kUCbxpQwemWueyfZjeGJXd1yrHSXN8Gy1nEcBrp+LjQFwJwlvfh
EKv1bA2V2siT6GCx6SqTXHgtuRUUsUM8br3y0PGasBwmfR3WHIznOWIh0UyWw24U
/vsBfib/6AzXJS38JYuI7DZhqIvzKgIr5ijJ2DoSAzhxxDZm01+Uw1UHBGbvamBo
pBZFubSF0VyC8AveviHLH0b//6oiRoaNAiQsW5UZGf1A12RBRHooRU8HX4v6Orcz
vM5kR1sIJXR+I8Oiyk31auYQ3ic19iVMkkk+/yoYtD6tJujzH4qyzmXqD/SZWBGV
ZL/1zipYcP+T5FGEnv8vdiNmDd/rehuJFkmalloSqOIcoN7ZIdzmXfgQ+waR9rRT
SMVpcgvVriKhv2Rkv+PP31TUqGVi+jp/cCWG/oA7PIlVy5TxaS+UyiCKBU8ApNQQ
JXwVVnxxi3PRM0oAqDUYTouGcb7T/F8LjKYvWL19ML2gjVN3TKUzsTF1B7CVFhbX
RtNxBJwh/0MNPa2Js+fzC7VgcjJCJWUvVN2nY9mlsDu4S1rgokpDi41qi/spdPwS
1fovs5hOoTrqyCttnUxKxjFbt/H0tLMSPtcP/A5nZzczjvpM8QlRLL2yXI3V43Wb
KelezUV3J3VskVh0LyMWWi4VZYblPZ3piRNB0gfNtw6YeffbjOdQdc0hVgPIR0J6
4tyK4B1CcY3UQplRN9p66rhGalSCZrYAInCeEw+6Yc8a9hITdFtrxSp6NNf5M/Bh
cxh3klncOGKCgp4ZJkKXLLlmjN8q10lnxe2UsFRzFXExwBRT84yO5YABPjgL8GDg
7tAyOPvm3MpjbHVixFhUKY+UeW3kAhGWWVblnSrs6uzRTPsoe4CPypffuTRMSqf9
EkBqfj+79ffpoQZO+LXRjt8HmVzebN91jhDvWPB/HydAH1vcPYiZONhCQkGLUukH
4CItHrRr7lXR2+G8EyDN3y9GMNQUi8QVkHmf5PZQFfWhVQb1CFTVfbq/czbE4bzj
yOgaf06OgPkbWOm4LSQNGiVGEzDVhbu8GThxMmdaHAXDfG9Sm6g949Ia84DdLJpf
wZtRNlaVB1g69C+X6fiOkTuvQQBIm0JsUQZfUdy4I0WmP/AQ5GXzYGQSOgownAxF
3A//c61mtj5v9ocAphppa5mi1OXqyWrcwWVp3i3w+CwPJN9bR4wfi471FXK8FCnp
0GA62q20JZmvGnasjpHYWsV+IS2N/b9Hk7N48c1qQoTd8oUm75wvwHS3GbiBiXoJ
wSxQeMczDBLnWpD6/+dWLioMX1vM9nElfk0uXojLotXE3rKQN7t8ifn5XyhtG2qa
xrmXck4Pa6QQg8R36y/EmO25He/EvK3a2VUWpdLPN9t1XtrOGws737I+GnUn18JM
UmjdxPt2xyPbtNndaNPD1bqZJhtDdlJ0OQQiK39591jZZB8rgh4bCNdxahEpJ1Cz
XOR/RpMwtBUEx9MtqmSgDRgW2gSfuQBLTchmONVRNnLPMD9d0smLqXrVqi82iaAB
cEGVzba1h0B1ZV2/6f4uWlPYBbWakcJ7g9s4iaYlAjjSr+FQDJQ6Ibr9FuqFKtrD
tOmvvntSRTEsVaHbmtdfwd9g613vDMEFjrat3q+1miKOPUiv0EPNHNNSQ7uHDXbY
ZXlBiZM2vxUOriww0h/SDljKo/RgIon3FaveVQrr+YFnL/tPA6EqqhUfQ45oHVTq
h1+aO7xDS85Bub/5raWNVTKNk+xDtETBsQhOrmqshSpASGonxLikvBhZzTOYPdq4
sf4BHh+kdoAohWhmC7clXzXyUwrT4div8wpIpverMLFfC4RgWGCryfHpTqdYZZkA
mB3gKq4BEgZy6Ce2++BvzmC+e55aTQOvkCl/JrWNEl83Ny9rg13n3rRYX/STZb9F
g80OWxCh+EA3Hdi4ukBOFnof1+u0mM3eQwIaAXy0LkDa60Q4TTWydqreXEdFdTbL
kzGrWourB7vUdVD6w75VaKY3sP9G5FMF7cfx0xe3ah6IXhUXNt33tFmcZy639jHa
Rd8Nlvhqd16KMzV2Alw0zdbo8NLPYVhAvg1l7nruN/H9BX1PStJDtiVmk+o9gpjy
j5oR6xMSk4FPg0++UH1YCXVVjKdJimGsBZ16bkv5y2uFzgJZZnuu7DXla0/gNToJ
URRXXdtVFlfeZgjSkDcXvNf21D6ekwiOGJpuUwE71cqDBh8E34hYPe9u+F1ElzIu
C1u7xxma2Lm3LpriyND7bCg3wBfc1FtX9M/nWdgxdEyTr9FbWRJhV2HWVM8jdpod
vW7yL+iRQRj+BDVxkoHL0QtNf+d89ZHuoRYtXksERT/rzLYPjMPgBPdNi/KangxZ
jIypPvOF1r6NZ5TWnw+L7YQzwtbkGr6n0hKAQsaxWVDQkkD/DItMuvUsQYldHYyg
3umpYQasCg0SpdqP8/SL/SAkKxbhJICy9h4B//0Rlz+6oCwS/E4vn7XdYcZ3xU6b
l3iBmhULfdWgtNWMxGXX2ObTFNOIgr4qKKjP3nsXdu5WYwsJiBctpA4lzxJF5J5z
rhAKKp6vEGGAP325j9yxxdk2iSM3EFUXFhL43IBYRLdvVw8IFuRRHgzF/H7VEGwN
fzPcpuv6sMVIBlja357lY2OivwyLXvaYFiSc0FfaAzBXR9bZhbMpP4pkPXmmRgf6
aJPawnwjiBHLauzsEov2TkoE6CfA6NXFFUQ87lpOKd/inmlSyUjqOeRYUME9/zXB
qogYk9+LmUVTfwoGqTP1jpZBP5m/2+dpdZLURgSnWbvumTmDRsn4/q/jrT78++K+
n88sqhTEFnaA/xAVwW805Tke5ltsaRdef/hiPGjW1/rSbJwbGWy3jL77su4pVEwL
vf0iqqSoqsA6eD4pjedvD74AXzNqDNxKWfclg9vzYN0R1Z6/L5+0mEeTdVC7e6bi
pz2SpKPVK/nO10w/9QKO+Td7kaP6pGzMutS5yQW+zYaNtFZzPXL/hjbHtN0impTU
DSDEYLkDCmW3X4QFSwO5UpYtnovp1aLERYaxcKdbGtKPMIpc5Rtg+cYG1kDe4p9r
P8MUvWLe1tY5B5xjvYzu4YEhYTMD9lMCWPQIbEuwzMAvR3wYpwpMPq3klHAhUmv5
cSvwOB1UJ4xrhF+cxlglsfNxYSKuPVdEvhQMQBM2oD0n26s0wM7yhgziG0EyC4Zv
5g0bDo/zAmh0doBz/d0PkWNJyu/D1l2xYIAP2ERO5/xBF+N1vzjapTKW+3g2wUDk
H/TA+0DoCZLYBOl6c39uMKHjLF55aEZzMte/c6SYuV/f3c/YiG2f/vcjONcGyFgN
Y2XzwJfXWffWMoWvykrapcXy/nGPKF6eHoqmcYW6K+lfj+gALFsEGcnO/fV8A9b/
IXqKaON7mIjNMsfEN/Cp60d7EWcW7iGm5Pd+gpJtLbuxee1rYDuS5R/pMtzrHxFL
qbNYn5WTXmR5GwviVcZwuaUEuYyl7PDUI1vV6/XdIFFbpjiIkHEFmUjV0eO+NU+N
/fsQ1tQ5ejIgZ8QU3s/TgaNk7/2DKxWkphGb971IvYg42HB1SJLinN9UCZok6UHM
D3NoKTBgf91RJnfH+ho3+WRYopdiKcnZo47yWwqeQGRygyu97wHoAMgxKWVfjoXy
pIJ63/oJH97AKPgzj6ZCa1LBDXP8CzwzIMmlQzDy6UoHeBrrJPtnZgQ4stGM+G8q
gnnkFcyTDzKge4ZDg7WpX77LPS/XW+qlOxdQC0UV+to8raWGEPoRH4r/hgT04dT6
7jXJnBkQkl/3Jm9lPJhJJhqtewG2Krbdf+Lve1LJ31PtJEZ3P494s14mHIq3r8MM
UEwQXSvulLNxl1SNBMdK9LxoJU7JJfBTpSBCPsP20ApfwauzPjS4mIGgTIU3cEYI
cy/SIQW+LfFu995C091l7pamEuOq9rfKvFMEl/EPb8g38D6OR91MGuRMHdOd0k1R
DotBE+WjvhT5LUky76qT4Q3ruVkg4abq8i9iSAU8bwaQ6lyZKHhT2lZWmQbz4SiF
SNVw2+5TARB1WBC1VE4Nz7wIhBjm1Yjrbvfsnf6esgtML/gDiob4I8SFtya3u62v
oqS4/q5q6WQ97CIruD3V3hZ2z3aa4umA1Hrvf7ePbSyr4wY0agOGT1lFLRPiu0TY
QiVJdUgEYUcc1VXN0JuckvVMyreXTH7u8FgfXng/SgzaTe5WtDE39sRh27AxHjDt
WGUcb5RgqCAV8ToQ7RWFvyFl2ypHLjEJ+xWmcOB4Tv+LJFphsCglo9MdMrUj/PO6
u+5+KxtpCMcrvTZ++G75gPEJAWLytKRgf0BKdoE1XqpBEMVdV+R0Etb6m+gmjSZH
ZObiBoz/YX4WyFLg/+oDEquzzISE9y792EfFybAfc3YyjWaP4kfK4ciq1rvd1DSX
kWAT1s/QotRyy3hivP5PL5MZc+n/RA6dCew3Khpd5HxhQAU+nffMjwvkmE7D2TkG
4JxrGoJKu/4hV92fzkN1VP/nsw7RPwpXbdhy0MRprMM0YUCymkOOMJ0GzazFDPJl
sgq7ks+hN3LcZeUeXTHfPLEEoxcWDom1EIlnvCE2zg5l4HXUWFqlknj/jWV/EKJv
TeC1Ovr+khJb10DHf0Rl74pmA+UNXCLU8sjJiD/PtTTAF3cB/tC3a//6SKQo0kUq
jkdveED8b8yrb1DN91WeElMqLzNEPCd/FVItXs5qs0Y4D5LypLChzL3du8At2aFa
MSKYa6SZBxgpbh7bBgB/+sujMq2G2caBG3p4eJZXmsiydqxlaqyro3YlHpsQiQHc
BSR2MRVJJMJ28RecRQx6v9SOh30KEpVxIY1rsrpuT6J+YA784xPfjGYrN/q+mWkG
b/YKMfiLgMeBDaURbSBERWGAFt1wNqnpmJeo1ERfqfWBh7zwn8nteb4CtLxHY4sA
RFoSpJLNYAFEXgWa1WjgGZjCRxGoU1ecZ7KLzSvIBhRJVrnDWilNp2+SgDAcVNmo
YlfqkR4ztpUNqXhJM9/kF31nrv9IwSY9/rKwnYjGsr51HYJBQrqZ8CpecFQtJwjN
ZhJLWwx5sr+YnLADkhdlvXkG0u5frelabKNsLlFlZ7yGz7Dvc7K/VP4gQHCGkCdl
pvuKnM79mA/3WGN6Hl+bVf9xRHVuhPu+eXfmkTs1/iINTtU2QGuejAk6V4JwPXLO
hGi+MprbaoeLWJzCKryCQkDLREqXIUmeod9G9nJWG74uTJnne54Qa+wFT2wS1wE3
S7u3n5PqDZq4uCbsG2GpHt/QlYqzDEU+TPv6LRcTTO/Hw2NOwiERERNtuVkNx/Ry
76N+sM0JhZCuo/3WpsiTDcei8btS14ecigl4HVmjlKdSyrmSaYiJG5bFPLAUjGwu
zYjBT3WEJsBmpdqXqPKuSctOC0+axjpcKHfO+N9Z/8zG+kpF9UEt8A6y3wCir7AU
jR75YsMMJEQwCBgz0yKTg6l9J1sxG5GRIJDzkXGrAJXnIL5p67Q+sh2jYx0Ms57z
I8vVLad+GEtarnJIRKvjlG9ff9d6RS4sowXkh+vhjCPZE1C64D2F+vV3WU6jqUVC
kfx/l4zGQeulHFVuXhFr6nKlWPMTBanImOpVynCctV78MNg3F33Ayhxt7uYj4D2c
9gl3/3fiyR/fjYZy3lAry/VWbBPMJ8upPHcJkpBs5yTGIRaKB7xej90TW9xEo3E0
m1DAahmqh1KGoLkFXLeMVAVL3WI1k8izzYYUCUYsH9MEUH2+sKZedxeNDUPZfvII
sb99ANQPkDjwr8zxdVIuvPj68lJjVIgUP8Iyk5PMVmNgosCpXEL0CD0pXit1iEE/
YdsdSpoQw56B724SYS6VZ06ouyfoXAxwettngNmHjGd0bd7f+jNvIesNchNqahg0
Eva2gbXA6ZWfxv65Zvd9cU/lzV4uL6yOu7d2HC4Z+eGoI7VkxricgYN63RSPrWiC
Hhp9YjguoVEiN7wYkt0+budFVrFNHArbQ6b5XEDfC/chbvswu832pZVvbIzk/bYU
p6Xn/k0vH1GmALRlguArDER548VjGTLwxmqb4QyM0D+5cO2ec0bb4cWTDsOsIEKR
uS29iGBUwlbG8oDOCnsGs2BmBvdhAC/5/L/HweqdYiCMMF06ZmvjcUG/BPJnLsnO
8k35bLxEAN5FioXJt6Yi2kuTeCXKhxK/+OTVqMZ+r3dYecUmfsPl7LKfI6MbWk6l
QKL9YfR9BTbe2xXLp97ZZmiolMLypyDeGWR8RF5fS1JBmg9sDu5EEKNXezBvS9Ad
ENxS9hp3qwnescFTLQ8zeqZxCbWlvSZLxCLuOjioRyYIeBcwrzqnrTVp8mCBLxMx
PQM+PuY2pO3tux76uuqKbK/CL+HKJoiE0uwpbH19dEO7t8pwqgzK+XKEhCHTHINE
lqbJbDudjQdkCN4V/VQub8ccIyGhNNMJMtQkJr/411UhahRDMLZwnDuA3uJhTvzn
kTIX2h8jG5C+LB0PBoVdzBg/h0THmHhsHlLAnicvouBCEqdYHuiDYMB/umvuCGCw
Yt1J/JAZY8zDc+1ORwu7ff+nAqhh+qDHTTmtfGLga/JlJhh/iGb7Gwhy2DDkIKJf
JVB90lnPCJAbqvUf+zYPcaMIGqdp6mUYYbAXtvA3cEnTyO6NHaWxJhMaaa7YxG46
3fDTfNAiG7Y3vnHjhoFjl9UDafXjmzjTM0YZvEy3kZn8PpiRtQrmhozRBu9XRPT7
paKvz18PXcvOf0Nw3kacPL23qkJTtZzbplpAEyHAJOMA1O86oZo0cOCcWANutpaq
Y/VdGiv93LHeDpcdEpoKCJfycf0MLO+oqSU/LCFixHsVE6/CoIdr6rOzB2NHPNhT
M7mp6qDVT/0kEfwX3KTJtx9JwaUAnCW6QG89PuPo6qV6J7v+lgAl9WYtR/rfjIpy
R9g/KhC6QRKGvI47NuYgoKZPM7U7qOFK8F+j4oYeTCzL9qExV+EyH1XtrXpTqNQG
AuAfu1EuRQ4QhdpOjsFW22FoGduQIbX1tNIUQfpFXJplPMvLBu49ksSzJV9jN4rF
BdgAVCvovOmSGWKJb42FGx6PuhNGHzcTqirh6hLTt1X93p+gQxcSrCOlkKUwDXic
XbS/DLUuEUlc2DcZVpj0JUx50PALliLWZyjDS7gIWYsWdQMnXJsBUWkIU6ZVnXU7
QI1ymEWBfAfgztPPdKnyW0SRo3VCNWyvyPvsbMQW4LsLtZeiKKIH3JQyhnedwbau
g1Hy1IsdCffhzmLuyZzoiQqcJR9OwAJsr9MHXx75n7+VoybtbGP4zgpbaiAiokko
3uVuPlUUWntDPGigksWTyDgYF8Hl4n0p582zN12/sCCEGACnyvr86h0/VW/kTL1l
4uxnnevXVsBWK5IRIvxT/VFv43o5ie384tD2xXo7mEBix6Gk79jLFNQ28Y3OUhfA
k365sQpKokWy9cHFZGwmvu+TCyjDd8o1HD8js5y118XDUw7weoyGCC/NpmOkUpCU
g2BqgT597bAoiv0BmIEh5t8OQLR41H+xFYXPIXTc01B3hgfmtbHr27Ii/Yf3iUWk
wDfjAieQrUKtlDx7XhY2RqeWx0xtync0SM1bJKJfj8ky60YdnW3j3NJkcb5QXATY
X1VZjHwcGpvXDUjmwL2hu60JRfPw6q2RS02QzoitwlUdGr5kJMH1avfcN4lFlHGz
227IZTiDvPgRvQkqVqh5EbAAP1yv6aV1ruZTT2HWl4tVJ2vGfWswczdC8xjwOxgR
4eWbEP0EcbHtzCAdGMM7avDThetouKM83RHEf4jJhuY1czBnA8vSNgLqgNxEwWJr
866JQYAO4aNLtB4LZd/YrsIe3e2pfdz35WhkPML/307rJgOetILCYF2+rFArHqtn
5G8wky7pB1PaUvfjbpKykbzVnHFdfzYRHQvxJ4Gy/k6bH3hD06EhQGm0SnNLFX8b
ajK/ey8HGwi9xy9iHWELfC+9qsWWtpeUz/s6BGr3tC4jvMqA7shGfWo4p0Jfa+kS
UZaekC6jHcx2bvYWgm2DbfNR7jQKsJM/XzOB0mWZni9KeHFzfmxh48kOuTGvebfd
iwIvwZOjGxpsb8OvWxE+K+PPWrgor6WvMxdCNdakb5S4V9xM+Buk8FnDFcuhAxv4
MRnfirz8ResAfSxNOsFne36Ty6CHZDE1hzT6iTBP7VsW38CL//a2UCzeiFuYsnFM
JNLefwJ477iS4+Uqh+nAvbq8VoCzpr2T89XU55f7eb7ux2ByyJJS9e6ap7XqLXDt
8HVeW0pHUvMu+pjXhC0+zQgkjBBmJ8xTt1Jo4wHPxxGnR3M5IoOUHERWNlSvbgC0
bJrHluXsUGdTdGXoM0tCdmvfZHfOyciKoy3jYA8ntHOgZ/tiNqEB9TsfvP5n6VOX
U478BgWdXiv/eFMA9BlzJ1j3O8YSFaH/qQsfDt3qXINOnq+Kikwtnv/3IKPpxfnL
aWlBXU3izWnBcgEGapMW4pX8ryWPOOPTNALMD/rbDfEDK8hG7hQJgLThzNxm3rVJ
gDuBZVEATdDLgr4IHtrQAnaSa6FkjPvAP/jg0ufNsOj4Zfi+AnKADwRY5IrkbE9l
HZyYFzK0lpOWy/ijhXAgg+KI99couc05UKllaRJ5jntxoqqCGmg0xbnzX8RGii1b
F66UK+ytGkTGlac1lfTLg2ilNRztFrVagDCpI9C099uhjC8LxaAAid67oRxLS7fc
BWqjWtRBmzkonU8yIot+cJL3Eu0qPZ9ocYuSEAToCUoRJyY4suMEdwcjRebIBdJq
tDHwF9Vt3WBkZw0f7aRh0j2QJom+wuFzRatjMYATapYI+Qag6OVPvJCKqAY7lSG9
ejzXhaURyBkzS+3ejd2i/a4S/N7W29q8M9ZTEsDn5OX3xa2FOiu9N9K072RXO5jT
WinBVLswlKxt+4e6/ya3dAxrZN/lh8N3YuueoJgmuTvbe/S24Q88WGbVUc2xjOWk
OGpGnl34/Vo/c11IrY6TtFY5ExQkLSvFh5F28pNW3XHIEFgvM0Ubf42/apV6sNUg
+6UrR3DzsU3furbARH8n2ChsMfp/WmdFIft4OLLM4q1cgtOPTIz0vODEQ/Sfi6jG
kodY/T6R2wIT+NMX2Fy52GNTaibA37jPirSXzllr51mXrb2rTbgKmMfn9mVKUtO+
nqFmkKAMCU7a3+3TVNgQVLSM01ueK1Wdm94quVypc8n287mYslczMpD3pqFq9glV
680n9HsmHAP8i/+dRAVOYABbPv7dc52tgo8D7zMxWdVlGkWdVBfBaTnXicQrXImY
VbJaG/Um8y6BPItoAZHT/DrvsHWhfMYCutwA8Ij7XMzBr0GUkXEdOcav9rYrzF12
MIRW9y6Fx+m62dvxZWLvcQEAqChWYi52wogdUtHfLL/WAp+m0XUT9KM+fpHB5HYX
aMG0cD2C54Ks/Z7CjpnrE4evcY+pZI5QgZn2wUdProo8MvJMKPGNeoZI1WXeLjCc
O+s/bsRVFBJBF+TVjV0nVgEorBWwR/xWgCV4DHBVOMvTiNHC9O+hJKqRAwljcxYT
QYNZpkpRUDJs30qb4GvAhHAuoPAIeoMHs4T80+DkU4dXw0Bss8eiRhkHh6J0LGZ3
qrR5XyCYAUxMUNXnx2/svyU1i2UByBmN556tsbsjjJQVmabZUmfMS+kkmmpYNgJ4
mCMdvjE37lYHPbmmslud55w4exnpzbM/cf/f+Eh7yKaljrNxmQuoG7jTN9wziTZ7
PwIoKWVbIVPCtBCTEi8aI9qmuMDCROOA63LPdGlIbrp2XTtf+zqQGdpqCY8cY0N8
lkFJtUPQJnLbzOmxtkzQzYwSC9eUX/prVQ1ecnkvgdLkDp+V+sF2edg1wRIiwMM0
KAHB4rUDy0VomvQcnQ4oIbt4vj1AH4khTad3NVNMe+BXlLyrsonixnXIrFu/HIDn
ZcHQw75QcJvDQIj/TDpgTcjuawdIWx6KoXqQnsb9VniAQsd6KAVzXN0EWhQC1L9s
YLsnMFKCfo+Z/bNP9Tc+0ancnsHhRLXi3Eit9H0I9M1sIXo3GhyqLWftEUcBNBsl
b7EmgnJOwFOxSGOB1069ZX+f2jn+z3qkeWrf6RUqf2U6VeDVH7wCgxSEBUXTjpab
0rDTC7CBItF+1cuUNiiJLHhOUUZZbZJPNVdj1OtgVmDOhiyMOsU7Yo0MBDDe0KZZ
c2xR72bVcVjKszo2uVEg8zk2hdOS8BqAT3CoPfjg9GwPtMq6bGmlLzCrjdbhpr9J
iWf5PjdQ8HyEmS5vHtMOTjIndTkHCoKlUIFVyBC58KYH9l5Nxsa4ra8GyYaXzK8x
dQWC41y3pk3jXQfql5vHmtkxnGsk3bjBUvuKOU6lO2evMRcZFT0XzyUdyI4skMdT
qs/+i2tU79bYmLWi2oPg0nzJT8wlaCsLSn4iaQ2CMEBPVQr1H8+g4mgdc4gk7T45
5MOB62r4LROUCkUfX1HZyvUBAYoptuGz+jT+GtavyfySxM6uAAFjrnMV7nKat7+c
XhulJp70o1LY9c2J1BkhnJcazCviYowNxtiCxrboJS4DmV0vVa31P89VZC8mXB+c
+iCJSDGSkjP4kns1Vxu3Z9yQ6JeOPykaH6KQPhq+sAM2KaUQLJh9RLhG/QpyHb/V
ZFMM7Au8U9YThWeKxnOvVvZvAYcK+AzTxcnBaHbVVa7fdBQO6bVZaFGlrY51gLMY
uyJT1/kWj3LZsdycrnijpXzurZ1xnS8dzovYbf26vZaoic7ZEivcCMK73a6RW87d
9M3wI1EGzKN1JRw2Wz56PolF7M04sOWKBg4mFwvGeRBsD2+cuma7bjJLrQaDgIIY
lKfknzR7i81OsT6uSwaUmJ4RZmkFV53oJaGvJDMA+fIcicLWJSG04I6dJppXe7QC
p0er+b47F30eAdIjpr6VyAZJwTDj8uPhFFJ88SJst0I1kj0SkNVbx3fR3Q9Ys3+Q
wk7xzB63T5yAYU+kwg7cCR4siR3lTCFFcUCZE7pWkb3xYzwBinLQWXPtlSPIVrpI
j0Fqs8nmCy5IcFD5jCeOvUcrcuVRuXmZ8Ekl0lzYakiAb4e3vZSyl1DCu0056aWq
FEXF79pTI98DqQfFFtO97GlGtLyRLzyiHkZ6KcxZeeQnl4rZU+CpCEADITi6Y4pm
N6KwCWF9iM6GCiAtueLo/sWNQmYhEtVxYUPFwTX56kNwIp1J3eK8PbLQqKbnsrHu
UHUsL+cd0rIhpBPuZuU4a5cunsQU0XAKDQHH7P/hy27wQQk9+jW2oosFrcgFdhkN
Ozkdn33yOhlrVgeIo73Y42SW9G1Z+dtHSR1BKFZqQNHiE+/RDnsPj/ZvUfoet5GD
LXdU6tIySc22vqAJs28qCQ4fG4X54nhbgbeU9pEBgHi37oWudCZGwq05zhpmpwT1
nEQvsA4vLPQ9dv96sW7S2F87C649zssy2nQqfpKdyYOF64La9Oq7CIp8IiAy13Li
vnqc8z8XuuMuc+ue7VUqpym2oqKNYy1OPoxy+5I8eHrLjBQmNUEiATj/4b+2KAU/
eze5CuKjhhp/BDPqQqGKsn/hMaU2wmabpo/CycxVJvL+inxlPWCS2+0vXSf1FCGi
7jravW1kyq6xbtaxxgyvmF2flt7YUQpJ7THzDlHeWEwKSHhLiPnjNqBGesTkLLTi
UKhUR65NKmdLpYny4JhFHLLwnDcHORfJuCOd8vNFPO5CqcUNDSRV8o/J5uVuVaIr
g1J1AwmGB7Oia976fskjQ4EabcdfPUSpREtzW8Ale8I36loThw0tsZd8wst54FmG
O4wb1yLdyw+FMHCI7ug4VCL++zL/zzdvSUqcbkQVviiaKn8KCqjX+DtgpW3vl6po
Cgb+AWlI203UbG8V4W7ADqIaOWwtwFTxDkRXX9SC+5sG6RxpiqXJZRrBwF/g/DkT
a6hRlyB2t4LsYGr4ENn5Mk9k0ADpaO3d45hv0Qoz/5CSsDgxkUcwv39HIpokmSMa
Uy8U+GXxRw0oBu/Yzw/z+jXLpSnUxDAjOkirhgOJdippQfYlgw+lQOKqvJycMBvW
kyIGPJyQ53Ezb+mJMUoOFzoU/vtj9oweFnm1iXtm4CIoeoQDo3hOJItvFw4ALINn
/+64wBY0pwniWQn/J5E6e97K8NeyUiL4BewjAO9YkceBXDZMXACmQcV8Y4MaM14v
t9pNgI8bePwoNz1z28V36niC2NfkjRU5XAMo6bbzjFIzYtlhPLFq2+FmTpSSA5Ys
mHC34/4N72WXXg3k2rvd2KtQnf+Hpr8ST+lghsh4TNGHfgRq2xXNtXUvL55aWXLJ
znMaXkXkEcLmXaJ+Breg9rNWX1fKQUZTvmDTiAOfd1xTVgQj8BMj0s+gizrosSuh
uUcSqIP4mJajhk0l3QdVExs1DWqYDPJAxjI1/QoZIEwXR1ALG0sZBNCz67UUIRR4
iLlnJgogYqWtWok2au9Rq/Ise71tUHLuq1cvgHpqmaPiMSu61bprZfFyV3aUi+HO
avEx3vY+DE5jWLyT0dCIljDNEypEEYcvwBNJHQWii/62x3AJBUJGu1C2eEIk58gK
TRp2oXzE1nSNtrgt1pOTmQ5Ka7N2v/A50amQFzjZvx1zfqM/b9zv32dZZDhgL1Im
bLAZrhN5Dh/X87FBStsYIb5+VLxyCLUnqh5sOjbIyVEqortD2+MDB42MFjdVK+Av
PkVJO0t0KF7aF41/FDLaztZ0Sfrch+CsAgtftSksFaKcSQAEjYqYIEWUjHLSnwCM
oEIhglsEX9k/NeTioPmQ0GpWGZ5JfYKxuzqJd0g3BctniAk8iBtcu64dKYeYjYB3
EuzoXHovplLRHaYN6DBQSzV6gbQ0M+9iro4KPpsvc5JRv1c8GyGKIu7ykDMzZYaz
i9kwt6LIyJoptPPlPXc5djEmz7FVz51WsTq5qsMmxVS6QnEzr7VRvnF03FNBGwkv
XK8qaCp9dd9erdXcKyukdihPaz4RfmVcM7vPK1qaF3Tj0ZsrfCMmsJWWvZIeNJkp
l6O77GMcHncvch/Vm4TXAPlYKStTadNk2SUk65Q/AgIFGgR/i54OqIYQbVnCGxJW
/d2ByYkfpIGsNfCNIKb0Zvji+N2mUPJUMs8fDdNAGkN8ODp/liBKfORFgstPJjcP
2vMimnw6JF3MNS8dZQzCGK/FS93cGcYSNdFkzkBWoWSrqEZyKHqkEhd1ecDTuYCQ
pXKwdwpLsmy7iQ89G+iCMKiycrnZyzR3pM99SGL/mgfUJflHDycZABpKrUWm7epB
kCUUgp+CXQkff/hxgS8fLJnHtci/kUVrzzln2h0Z2au2CdXWyqXwTtz2WHAy0gqq
uvj8RPgSBF3KQFD4UHS1a4jHb3xBK2qe0z2nBNt1XJ1DMTcyttcGXf3d7MCTNdNP
R09MbxMeAVWM9bv+0/6lLkxnsHsIaWHsTmqN+j98G0VjRFP3yuN7WcVVzg6/E1dx
34lfDTdE8XUtDHp3L4vrxHH82Ovyd9mpqf6o4lcaB9/zFNZVh2U/D5d+QCRYr3BG
4KcV3+h6AM/2aW0tOpmcrRJ3jBuQkE35Vg+hBAlW5tcXRjTZwPGCOZaKxb57xMFy
OnD7/Nsn3P/q6aQGc/3CaSv25Bq0vySNGk4vqGb9jaEH9iCFaBG0VGaeCMCu8qjo
kIiGEAGu4tpwiRUXfTtoWp3W83KcS8rgliXfrIzi3qLustOM3+jEMu6FL9KMuSRi
S76FZQEb24H7ozSEa1PY33S4Rf/fWvVGFKPBQ9NHP2Rv+qtt6+67vpmegsHfsiWJ
8VpHUjLCAEmrpWUfWz+UuEyDkruCH15+qfKoTnzERx7ESCIsG0LSLQblq7UiNZl4
y0faWTw5hpnAgP0GAtzd0YLXXuJgsBphdM3QGQczyu6lhcg5MIx0UgYtGUYx2sd/
nu+Cu6LP7geug6flulqU5wHJwqsLQcHe+EK/gdifSomQNIgJPsIgp2v6sHd9sizh
OnK1N2bA6YXKrUxlO7+nISF3YWD6uYl47u9CqXXiCQEEVomphx4QHKTAt05b4by2
ViLhJRG9H46rXtwXWqYgYKGIiQdbBau++l9NwLXwvmbmwIgWsui6bW7qRff1tXia
yCFEdL4kM37+PvfwknIUoSkuQlbhbZMhmY2sebaJIIjQQm+cAt+vG9FG2pmRmU33
xo1uf6LlTA2s/K9BqnP+/RWDC+A4YpgPC1pOvp2x1CWbYgOxD3FuAYKTi8a7y4sa
bwwwg98N1F0I7Y0wgtRiQH7aD5i37WiQPdzwdZs9c3znN4EPWjLpg+YfCyaKgSza
cA459dsXMdO/bBysycifpr4V0WQHqu3Jo7MQfk/QpVPX/g9N88hoqjOq612u07lY
jxQZGj6BfSVf1P0JLLKs+J18XtPML0eyHY9ekIDAeN4eVtzyFvCt0DqSYFQfiE7Q
QavjpK+7LSrLyiNaCMQggVTVx86cdmE7Jp3M6JcGqsnzt9lBh+pqpz5G+rz0kAkV
dHsoq19Uz4cZeEp/O2Hgbm7w5qFtt5kDiahgqY5QkbNocAsl7qjeyHbYjtLWJpT5
zAqDQpzd0jdMErxWzl64Dnjrk0y+VY3+4bSnFQmDW4+uY/bpxh3joTniDDHiSUsd
TqESGMnW+1ysxpqLvNj9q22e+hvnHfEmAk+FODfdW2FPqCmdnMOOaevlFv27MoK2
x867OV/rPA2K/ly2WWOVYIJK2wky6LRpgW107Nwtd7P81psnHO6CGHDEo+fCj6/k
39NE5dXUnrWgf4/YfawxjN8CSTvG/tH5JrYG4z168OkpO1Q7JQNC3PN0S5h19SxK
4KJYsEIJOw/j1RFLRd5KWblFgAUL8/OjUtNB1+ElhMyx13rbL/OmABkIzSPf6jj6
BrIpjmtcz1YWmh8D7H/aevcCTN+qX6tQ9uS2GTsNRH1lWiotjI7j+jBx13cXLXs+
vU1EysqbHnXjsRXnG369+YnKrMnYoC5RLFBqkv2TO4DYVv9VFEkXn4jzsXjqA3QN
UCjSz5vzBHmyuMZcLpaypf9WQYbyhXfIQjj8GBDN8Qy8y2jM/l/f/0Tsx7FvWthx
XuB+ftNFj03Ch4T5pjEsGtcbYewf5BLACNJPYAoh1iPrea7mlrrx7f0FiqmvskFk
h/Gn0RtoPDWcFvTpB2dw/rDkD2ZpPyVFLTkQknlXH8OBu22e/7wgf87pNLrXTUiq
CHbIzuD6IkjDMpFeUQ9awLcQmmf+pTE91oVHLClun68dxHvctx3RYtN7rhFAX6HV
0QDYmW+8AMF7YWCFRJlXauKSpROhMyFaAw/1AqAzbOj9fcAPYoHC7Ipk4tpTICoD
+/WUjTfY2jb9JuiNOWnppdf1LxKRAuhgKgq7FeUYai1QSaITcgqDPzJkciNdIhWM
rBAWZW9qA5vUKPcXdiEc6B4s5DVZ7VNAUZrMUGtS4/7jP2Nfa9zfy0kTvXZ6qx2A
PPl2PnTrtEh4mxrdoODUr8Bkr38rcgxhabpeptZBhnbylMGRz2axbAOvZHe0LJxG
EGgDwXI3kUkYbMvzj1CmDJGSp6/w4mIw3cCgWG2hrF5BmU+AnPCiVxq43Yy+yKv8
DezfS1LeHHk2odV3jVJ2Z76rtvuwDrQw2Wa8l22AHAiq+q4ERVMLMC8RuF/4lsJf
jmLyJ0bJreoVYHM0vOvejRhcZ+aRWsor6slBX5wmmI/GvsTswM2wZFP89eo5kHB1
EEww2oOjW8uOSUXT0hPGpjxraJDord1gp9u22ul3KqTZqdKk5czx2DpWw8r5Dnu/
n4jUm3HtdexQlXDuhz1UETpAgc1dSsHYnYU8hAKQlT1JacOQCmIz/KD2doIDGdQY
fdFttztUmMynpk7KdGMIUrHweay2UYgN0niXHFTxFl4aOelYzd56hl+WLOjBxX6M
d5Qj/Tw3cEe7o3UHsycmCARUVtj1z6Z9ITFpAcLyd3JBkJ0hAhyjxz/LKhlE8VZy
bMcSMuqGJZTwLf56yRmHivwF+5mV8WcV2v6D+rfOW/Lcs+FvKsPF8uAt3dgZOeew
LHi4/JNb4o+ooeOCFa2oHjIXEKdirJR+ub7JwMwUO4o3duJ2BjLEah/XynEvO4Ul
2PIC6wTC3IqB+yd0hHPwF9hDjURgMHXwTZO59+TgG//YZd+TVBvnrD87UY41/1r2
BWB8gjoKpFRL8B+OGQBgigNfIV6zfWjNOo6f31fDvxuwR3aqjFotfuNUBgC+w7NY
wUdcN/FMRZUJJLq1Svw4lcGbixFob5oqEFul0frJ+6T+3t0yCobUZAftp1UAoWU8
KyJZ31j6Em5nU5wh4lgyHhmOSZ8RT4Lz3ULIDlFfnBvOf2v2jU8ba1Tq2sxjnuCX
oICrdxbke7ZQyLul2LV8FWtQ5N1BGG3hp+ThnAkx4WcM+xLO+ARmZSg5d8ybbUBX
ESEh1j4ZlPebCVf/qlNi6nTvs9MaBmFXogn8fHZd7VpvYHQWHO5NLsfNhCIC/z3v
aDQhRZiiRxqrKNDtN0WaYJXfixP6gs7/fs+LkZFjmP94/BmXicA5WtM53qy/n+13
zMBvtlWdJvJiverC/N5YFETAN6S3eW11ss1yr4vwkSPqHmDRVFLpYNSrFNUaPhkh
Ay9kvbclvhJTzoCLgId9RepJYTM1GJZbA4kTSvu5DrTslT6+Qns++S2MFvFd07eT
212YX7W3Ityw9jvNAPmUrOLA0PrRHwB+LUv8DFfTuKvya+SD5BOBznEVGiaQGt0c
28dF7/VJCQdxRHgAvJpaW3LcHIXgZRk6l7HWPiiN5UDHOduMHGTG4zEgqEp3X9ew
nMoXqh5Bji5MgXyHvtPhHYHFWNJPAsdiqhKpzBw28Yjo9jlYiITJRTbBDx4lpjHY
hPrMrTcI5Kotsqn08FVy5Q8UXJss3uwxlq7NBJM7mfAeQnwwR0VUEIlv0jV7eqqU
CpC0L6lSUoKfCgUjpj4+C+P5oLE4oYjx1yCGMbTTZvNutiXa+EhaL/LXqZyyslSl
y29VrYiFcx6lj+dsXHC3FsNKvqJ8P4x77MeF6/Tsei4SvHT7oxA0x3KeOwWRawpH
5HjS15PxaQitU6CBUSmgy5ElmkwmU0+xAKYiseFxRbbJfb58sQ4Oy7lF5LtXrLHo
VKKJ+VxcX4qCUquk2OoBsEjlwl9tm5D5NeObKk2d8WiVucskfwqqsKf5KkE/EJUk
B4Z2mHEGDqWtgaP5UU0CNfA+Y4TCYn4hYNv53JquT4x1L4cTshJUR4lxYAHuEtJA
JCkIFmHhHOV6gNbh5JWEfLH+IqJVefZ8UvGzK9JlWy0u54yvwkEL8I8PRGD3oNhf
dNyxvxfKwI1lvCb9adh7XvPe05KRHYRn/afFBUSd81gjsDU/5Pugv+p+zqriX5EM
iWJ6WduOqYGVNRCre13O12zTS82TTeAzeLP1v8UfR70ylyGdsFaI1jcDAeEan5FN
22JDOVwWkkpyRf7av3Z+yI+vnO9qvpyBVnK6pF2jhaIRj9qn4GeEN5FwRQ5LR5uw
2HfUgqXLAqGd3f0hFR6472/bcMkX+3nYQBlp3V2bXfKeaUQbWWA8oIwLQiMhFu2f
XzcMmdNekwCGsq95ppzZTPqVK7aP0HKCGGKjqmsHyIzIsjPNa9U25Kxu1qQfdcZl
drHcEA3L5aFqUPUnP2g9xdSQYIoe+FspHVkQtbndHxYiPp0hUz18mnywlj0Ry/J3
rtbzMGMk5eTf8PZGJgX9C0NyyRTSncMIdfhBrg0uTTCLssyPYBx1ehXLWADg3mCJ
6II0c3eLgmb2mCdhQcZzeDMYaxML8scrqJel1Mxxj3RgT0IHtLQYse434/Hky17e
WpwF7jsS0wgqgba1Axc8sfyVa6H4E2m4dKjxGJnBEWA3wQppWnjir79W6L59Pdpi
Hl7SZ6MBXCs9IueiCeywqa8whLhRCTRmorZknHJ0omGIPh7qyZmdKjfPgrdcvED7
+0PoU+V8IDH8MDxdNjs7TMj5Kl41lYuIMn4S7cEp1P5HjY5hZVKA5Pj98jRxSObr
9Ni0L8BDUfO/NEB5oQ5QW6HwpbDEgcs55tfOv7cvdnaQsEbWE8lu2Xlo48N0oIBr
KzJo36rEMeVALSDZ6jAj5FPz6iEnDOFna1LPVaHJS6aHyLh8KVCXNCnhwTSgjklf
ecsVDZv0wqCT5+MxdMIJfQcLt+WWksy8T0r+72Pm6iCjYuhAem90MfWJXQ81HUN9
yPjQqKKziROzxZvWjsnMahbl7MyCLG2A83DlMJVV9odWroIbzuaxOxtwpiFUSWEI
K4GSySPn1kPsj55zdj2JW/d0tuw86AJDTTGzO6ICvjxPIfh+gEQzTDQX+fRB+Aen
sM37jGrmrwOJrGIhb5bLGddhKu+vJeW5IgnGjLauJUkUBSn+MbIwXE6P5WyIka7h
QP8qb58SU7HK45smdeP/ZjWRMrbkKDdvXEhhaxoXAGXsQPqa8zLm1+bmB7wQ+Klb
ud90jRnUdZJWA1uGvC+GK+n3duChHjzgOvsxUW6N9xxxfBveIC5jFjvE027JPzeA
ACTfTNpzZwlP+vMIs8zuh8Tqh0tzmP+KYJUpPf8r5GmW5bjE32NQ37/l8qbmbjAK
v8w1juL1Pi4p7P9KuX6I4/HZP+r//J9X3nF49TA/jOQzlZQJFY/CTXiFq5qfZFFL
jXMPa55ExTJbNB+M+k7Hno35GdAhQgcAclvNcwyiilxr6/PQj2fOyTN6Dw7EGV/X
flitzxIEB6VX6M94wuMvzXp9bkCAs9hYX/vaxML3N2YWkLp1iqgFccflfrSqk5cc
GaeLxuRuOQ+vhxj5M7AXjSKa3AgSCV+5HGtojGQB70musGT6/mhYtB7v3RuPB5o4
2eIs6bbi4mm9szqOqavCbNnlsK8s1/Ugu9kEkbF5Rl2zI0pQ2eyhl2LOSPIac4Z0
2/moOj3UMiLB/skHZmws4xmw+ZkpHZsBe66pLwvc/+HCGAzZ8HNjU3eSplLtpGhb
04Uo0dB5hmGk+he4LZWcipfFKqOXD1ffL0NhEvkc8scj6yiHFXsUFjA0WBSR587q
nW49sa1UHWgxuGbtI7vp4QVPb57XdonLfpG2+ZV8o/45pPsq9cU/nlwp/Rrefetk
n+f5IgNmu8icDVbmMnICIuYUXoSa01fngDFpWmMp3gry4aOqn84xEXfe4UNberl5
vypCi1Z8dw90PPnRqT16q1jBEdheTkXrM4SR0UuMpPnD/ySRYLbqBOuXK/tku7iJ
R0D53Z6PsoOa2xPCPRf9rwBXxWsPbaNzcXYnAc4NbJaAU0sJgKgi3ULQRUlAMM5c
gWaJwoebhI5sGC8Edmu8tKGIqH9tOCfYYO/u8uABCKHLk7ZZ83wKFxjPmnSnn8le
UekUdlNql+GAu1mWdBK/AjxFubI91x8XsRYW2nQ2v0rC5p4dHnpIn37PPtnDSerG
WZXEZTTWy+Zv+ad3uVFQtAgEJpk77QA/vP1p8OcN1ijaVjWudQqLjKjWZYf9YnCd
hUA7z6GUwsBzu2L4BuQWhmuzCfD9QQQoF2z0pc+n7Z82PwScxX2gva3aKUHcx43C
+5hl5MwRh92nQcjCn3MOfWBuPR2tVS6WPEsMTk6hiLGqg2RHsMx/y3nkAS5kCbtu
JaztVIQ99QeFAiCmjmH2tT9JSEfKo5Js3UpQC2v8t1T9PH7ePIzU5YxU9H5KfmT0
YFKbXSDE3l6yBwGVM1B+EZ8xO9FJu4282z5bDIZ6192WwnvxUN4q3SsG3Uzo5GHa
zMhogjGFIB5EvIu37AulkxFZEvoK8wuN2Wqh8O+/P/Xx9ILcKEQlNqjAGavkHFeQ
PzH64Dpc4A6R7K2EzX7aYRCrkyRXzxmurKuzgIRfrTltFXDVWx5EndylskeLszDs
mRN11aFLI6HoIuBZRjpkm/U2tu6JTk1maUxco6o4/zntiZrLgxH3Z8BFU3cwRtHV
2mnpOWEcyTrnn8HXs4O3RM/MwchBqReFIyyl9ZUKBoWPJr2FSrTCdc3g8SAD1ewt
6GF1Mp9wpdhq3BXZqsRWl/3lCeyHAs0goQ/CAUsWLoqTU5Z4Yl10fP7twNc8rWAI
zK7K2zUWYSfeb1tzCU4/LRaFl3RXA1UM7F9Fce+d3e0Zl1mSHi8hbnvJw/Ce9sVe
ddnfZkMonu7u7m90yV0Cr6uSg05/fPjxMAcc3xND8OA6OZfieFZXWmoYFdQfsg4P
bTTs7THSEvIBW6fzgJ697yynq7wSUya0ngdNaFw5Tc1ZpOQdT9Lp31kUPvWmFxJ+
hNSjd0a9IFbRHhZuDbhsa3T2ORgeC/RTHTrm6G2WVgV6AnNq/qH3uLUfKpTS5K0G
bdBva2TnUVukfxQIxvni4TC4H+hnrRrDDrdJ5pceHDSsrxlqO+mwMS4C890nQ7NU
rIrG8c8FblyF1Qvsc6xVjjU0yrJuxlIFiCLjjy/xPCaNH++EH9NjCKWjSDyMn4tI
hSRpRxTgtDssHQT1jkfP8AqLBFQ7lbVlqRmb2HknvNJj1spQ/eZ1kVN2uyRTcl9s
YcjbwC6QQIQs4cBD+o0aWYxLEpnFDdMkZKBrAhTCE+Gxxf3TTNm5usNZFTB/eydV
NM0wFev2/NkFgPemyeObLBo2Wf6TIKfSaejG9cDZPrQml+OTBlnJxJFsseUKNakO
6/EPrbdGKc/sd2XK4Xx4T4nUG0E4e3i/GN5bNKjjDTzuMS1eDyuPS6cQAiADxjnH
2AUZRD55pEduKs2iNW2Ac/mxZYWoAh0RadH8J5Avv571D0v+/Ly6ojcMU/tUuEmt
tiN/u5fNM2sr4jmp7nm8xL/4RqBpJsWoV0OvkoXilqqdSNrziieXxtQatxfPPw0q
okATIlUNjdDlkmoUhLn2DGGT/EnSUmbNlo1Ulu1k47n9ny7GHuB0mBG5dk1qAQI/
/nJdQcBhdygFH05B266JxS8A2L/1ZhalT1A7iYLcG+FAAC8NaV7Wxj1Rk0OkCrSS
Rku1IFIBDRqFDdm2D0ZVtxB9bFencI2ByJyiY8kqI4NbUpezu1Cn31sdkzOtcdwc
a22pxtzS2R6nhFYlKPz9yDDaZPg3SOGBPRv+2WM+56eiznh1j/koaav0Zz5foSLm
DjEXMmx0ispiXrAYuPetPtk7+oNoP2nEBCc2Ld9M1/66fH1yjGKrcCG59nWdcZz8
xxMkXvr6RyB0UTV/DkM18dnc7lkQPhLcCKYX4KAFqZyQ5RWVW65fYj7jntowGVCM
6wwQmfseJwQjijRVhGLqkwWNGV8VEOxTmRmNP9jwCwgul5SO+LXWzAvQNpGVRn3w
V1R3781g4JalSF6NoHLCpew8aVrnoQBZJKSuxtFl5gNG+26WFX0XhQkdfOaMKhqk
Q7gGtIWeCL1qf1VCtA7/QUNxE5znnlZO+GZuhzKM07CiJ4eHtyvyfXMzWJ2APxtm
Qg2/LgKcNs/okct6uX5/cSY+b+C0UmMdEDza0RZbnLr5op6qECJonw55xSxPcu/j
gCWc3a5BLUs8DOl9+9oZS/RM+TRxH3NkyTUk3YNbxac7Y9XfkN9BPsIckd2rFDl7
za2eyIiBOIBsv1mNsl0veZM4g0DsVSBaf31lrdpiwEyX/Loq20AO5rsHym0ATLV9
FLdGLFcoUIXgP1w4QGnN8FzBf0Zpr4Cdl3Nr005VSLmlKmEOYfv+wjldtVoV03Dr
bSHSYK2C3hEJdpsYVYX+aEOqg7xV4msQ5q7uprqA6j9JUeud9fR1jJElJPRNjIvV
hJtoLfS9mxUM5/XLOyVr837zG/lYO4axjWv/D0C6iG9sCmcAp9sU+/bXupsVfs2D
Vvd9pe6lcAyhhFRt+X664S4rAeW4sb0OKV2Cn9suG+c1CQChuLM+gOKzIYyGKcwx
APlLbJU45HqzVBqQizstzOOJkBT9JIb1uNEp0XeKT3scVHwts53rW9Qfw3WSBfZ3
iJPsiIm6q4ODt92h3W2tKdOUiw7PN6kDe/kfKwMtNQrd0TA6KsKdkwLjSvryk84X
b09tmOFd8Yc0hom+Xq4e4t7uGjOlVvbJi8nYqhE2ZBZqIulwPt0f8cDP09LvfuYj
XMK3ftORf/unyXGaRc/A92x/sn9rUHCKQGngq70iUmbs4aGN06eJkaBei6fR8iR5
I6rNvUD4C1+BzysLsyQnKwRU2nySCGFQSn5YBb8kDeuPQ7ubY9CEuauo2Fpck0JR
gbAvOvcx4PIY1XhKN+MwP58urYzjVDk1zvSEyqUeZwgOy3Bk7KBIIVeTpyZJ8v4u
BUvk/nwDOC0X9/x18MrZfJM4YOt9DkN8yChdbMRWYU4fJv7GHXQOTXVhNxdn9M2O
5i/XfG+BavIAmerePWFQKE4PUFuAxg1GIzyzz3M6UO5Z+figaPh63tH4i2kX7g7i
bR+ACIAB1Q508XUYuiKmxSq+mEsyA1C27TXXn/eXVwRzPhIKScJs80ZPTEoaCT8M
MhCRT1Tw7vJh+PenbE987yJOpcUYW5CtQb05lp1nMVRi72BMqLog+UPb+IeP8e1i
mvppY7RBZd0DCQBpkaR/tjN5r9fE5dkbw/l0VmMzFfE9RHwh1SLUx5N+V5xEqQH9
agxdEidpuQW4ZdvGDr9lms/mNuAnO1nIOhmSe3AdsoGm0odklMRRgrb/inPsJkZL
7ulBRazEyzn/arkc33UACpT/IT5t9d46WudfW5gO5iD1QfvFFmR9Eo1EC9rLbURj
gLv5/jo1cNFh3hQTJp7GLtxt0u021VfkwNHqRZ4yXQy/5uKDDl74BLn7A4wougXs
2HPEUx89UbWPGzzqp3yt2iun/Vxt/DItGOVoYERYNA27CZRAkscVxMkpHGtvPkfX
aEbPX9WzXZNG4hvuvPEQQz0mgJTxGO/VewJVYKqI2B0Wx67wKSAm/sfywcuDN5HN
XeN4hMhKsxIagpuPtmtIhJFfFg8smb5CS07g6O7S03OEefVkOAVKn4Z9yDteZxkI
xSvUrvL4AoNThESt299/bDvAcJyKl5Gm8ELH6dit4jrwpfzJwWIosro9bYtuF7on
fEbi/NC8HSNI/+kz/RMRQ3xfVDuaJuvqP22R054EbACwkUSj9gszJPxMbeqyRDbM
eGrbK+aO/iNlw3+bnLaO8kGQ3zEn5aE+NYMHqKcPtytAHe80aY+M6UzUxAhtijY5
tjZhK9Aasj0hkyK4K6Lu99K551D8iHLbRCsk37fVjKlLzaoDZlr0UoFyy7olKwrJ
Z6/BgF0mLun3Q5wSLSPvYWBgw4tjIkZPDpoUrLX9FFW36/YfXKirYw19feEkd47J
bug8kFMJTyAmWQfBZaek56FsBVJ9Md9bVNXwGF5ZGNUv/Z5EdGz9GdIbbWLW5tmU
19hzHzpWhUuucBOcbuLHJ5mtzloWdz2DDOaqqQfZfpQC18LcbRL2M4GtINDTWUVC
xd8+7NbjgJSCbdZ9JL0mfjz6MPIRkVHs8Xw1Vp8l/HphyEdENW5fOvA8RVJ6WYx6
tLF8ScmwVn6BAK6F5+6WiIpSBjgmpDAoIt+i9AYFDs1A5NbJZZxARUgYMkgdB10o
7IUutJD0a+Tq0UbI6ybUQkRDAKk3eRY9QlCIOt8bYaQJcJaKI6EV3JbKLXairLL2
TzJED2hRmZR+Kgf1QJyhG1fk6jpxVBXLxBxFvhKpNuXQ+hK49w/SdtvJSJM/FyGc
Yh5BvdZjiEX8SI93ZXho5dodbnwmYJmbx/wF+c509Wc7O4lTHJsCx+e+//Om/onp
WIt/tWgTZ5RiHha+O5LVi4RXvQWEVhohAUn1VNjlTZi1+3tF2dvbFAMJPlkgayEy
/XI9hIrOMsYUIj8zQh0DOENgMFkFAMPYCvusQofn2oRgUxScugkRuIkJPSbCwafp
1ioaDQS6XbXTyXII0U6DT03VbXsR98JDFo183ZaCb+95iONERPG7jtil2I9W9R1V
0oJNDOzBeaE3IcR143jo8QDfUlcqXSHciUUxBo8OL4vRfyOEqPUYiEHKzbg82Ggu
XmSBEploR/xXgcJh58pEdoAHTQnMN8z7KHeaqRFP9nwMYA1SfYrV+jDGztgeSsG1
1oC8/Js2fAKr3wMID1B9INvLN4tAAiIptqmbhRtPFAxHQ6wFno8cs3vRwEli9EyV
YGuhs6tef14jvPu/DlYCr18NNkUSfnEnutUFKWzBb+6TQiemOLTlMuQcMEdVCM07
HjaM8gVGMJ+lp+gA3X4C7qDcvkw8hd5Nj0AQpx4dMVprcTaiGSplgJHAZ6C/QybS
6tdoV8SUPVbhqI6nzbU+NsVzRwoE+3Xde3kAtlWfZWgm4iz4qS16RzLlouGCokT6
jSGlKMIUaT01USeTfunuM+x/BQ5UMovUW3aBSBJMDgUll86mbZEtvFoaeD1wwWqN
v8A3zhBXmbERnnr8HfUjHXKeU/jJO1rm+6poQ4TzFEmHr9QTefLg5VBiHuvkwe7b
ZewdgEspN5qPwcIQbQgMIIasWvu8+PwwDt2E4vujAQu/QctZmjjLhXgSYUSk/0h4
yeYPtvsd/yFa/IATsB+HbsG7kvVW8aUywMcRacSi0QApIGIfhatNfp8qVaU6VfCF
1N8ONeCuJI/L2v3BlZzp5uR9+2vPBFHthJ9rhA7JOje1bbCm7Ttb1g6e/TDp0JpT
ii16IgAcQhDPrjm/d+SkYH7hK5r5qQ1Zu6XnBBja3XXyZyedqU318SJ2ji2m+y2y
8yIuAGsfZYOy6quza3BrGez0M66NHuPNZ3CXy5LWnqs0AwzN/EfiYQ/5A45pkwHU
2+I/81VQ0C7VdNBYkY54kIlvssZiPyZ9nYVGcmS1UaPXRR5C1cndZQXLTb7vwjq1
0jwsPAoKSIEzldYg9w/6jge0IujshhljJWFaxQjKbWosZ35LRykFXwFY7dudLWux
jHUVvWn1UG5361fPZUOsbpd9pajg0ZulMXX+W26pc+H7DM1fsbQr4ojLtXWVJsW8
F4Dl+dDPkMvr3sty7IKfq4F4V+N8qWIP4QAu2+8qj5ftq84N4kRrFlwD9BZ0HJ3d
W7elkGgnI1F/YWRPsisKApWw1IJ+VVVYNDTAax/0naw+MKa8JeAMOol+cl2tDXL0
lfAD4jodhto6Nd9PA3cHWjcQSA6sctrDvqv+fdM5T0j602rQ+dz+Ln8asrfAw8jC
IWssp7JVnlcKd0O93nceWmrmalKrOAUxHCC4Vi4T7UYzKqUK7Eh4Tc5SZXxqUXFb
57kEE3+sFwxomlBUcs1FogIF470VMjImYMIv1rNyk8ZMoMyjESUuB2htQDds7LGp
LBpEXw2MjO6vrrkxlEwF/LieJG2TQ33IPjKGJcDhZxWxqLzaCP7FNg8FYpxP/Xey
qrbsfTt/4+1UmXhl0+5AUbUZs7t4fNGh892RqujOwSaVi/VM0LxBo4qHHpnRiVqN
lZJMzblqHZ1lwCnJv2G+4WvNNJYJzaOs5sNJkefOIdW7bpogJg2pisC8irvLGZ2h
3AGOdCPVwSK3JAb4hqz6eDzt3ky9LbIVg3yW2o8d69ndFaARyZ0HNXk/Mg/T6m4W
i2SE7lBcNIlvuliusp8WqgukLFbLwf5qiIRcHrI/llufAHwBZKcnxtIe5smCnwvF
ocXG9LdSKg/3s+CUmXCqBKKLQUVG+7Z2kKfqoYQiX5sN89MY8ASq6RdPl8sEk8wV
QkimJU7PcFUxa7b6h+h2wB9AV8ccW3qslAy7oSCusltFPy4Pq22ZNHwGIMfSornj
nMk9+VaalZ6lOLxFnBWl4z0Fhv6QlJGEJO4lwzl1rZ3SDdgqGHBDe0zwRfgzJe4N
wftE1+4lAUtVjAY3RU5APKo0c76p4Csom1iVRB2uB/W8i7sSWGkIHKC3s8XmK5sv
MPSqJKC3aEV4NwdvOpCCa5fFzaysk+ulQuXKETYiIXJvRMYf95z3/e+ivkVcuBIU
ctb7SV+a7cWLcXjOe5arfVXPN4SdSO82mNmsGbKGmy9rInqsATwaHlZezd5oWc3N
wYUv/8/iZGWXIYTikHSN1qgEMp4DZ7C7CnCcnQQUiD/Bz9dgR8OL9t/EQKzMjoIH
4Ex1DPUykS9Vz4qXxJM50ILmFFjh+0Pu1Cj3P/we+cVyJY9BLP7kQiMyiOMH+jYj
ykOWis6mfzCBXbCF9uwPI1lzwFF1S563sss0f8FpoSDU0nYYtjun6vi+7xJYOJHF
/sBiiXekULtN7u2+be6R8bVrtTG97aNzGEQzcWtas04lqjtkhQkWz3yh5I3h99UR
qAN3w+bCU40c6/7RXM+rZVS9dnZPPZ+yTwNKpRGHbYGRhVltNZMhRqfEy7Cz4HRL
INNq9n2txqrQB7F8zIB6tpAYhxT8M8ZJoerdtNUQ8cf5BvqHeDEGuKi6N1CQMpLg
+n1nVSuSqSck0kaJrfq83tu5ocqgnnpef9kHUPS0cg/8NUokLa+3N7ErQKA5syD9
oDp4qzI7T/0vib0UN1f0QTEFHa0vh8OWjqxchha/Rc/pUSwRRyHlEDvOvYGYJpLK
XuG06hTZjWZKQt1erlQ4L5bM03fDhcuO0+CApJLQ0FGfBzAf60uPplLzavzpRhQJ
ebvtmMD+3LksxRzIKkgmTa3bb9ejR6rwB/Z6ZaqUz5OPkvRZLraFhoIZXhu16xkg
0nYLelAjRyps2TyuotbGhaez8OuCpqif+Q4UhU9Y1rM/4SD+9N9jPm3eyIh8cP9H
QOn1c8NdX7PsgnAsGUdn/73jzAZyTW06msod3EMfYV3AK2DqMpt8TgHDk6n4er9W
Z55lzavHYnkV/NlIFa5ZLRnnCeD70N9wOq6wUZ6/RPWOWI+TEPH0PTfxxX74Am+y
2+rNAkHvLVMpPsdcYPLPCfEWDEg8NFMYQV9vyL6sJWHbxyPN4emOirDbFMWu29VV
5UrqCdv844eHFSU7BzqwxsaF6ZarDkJ6AOf/1b/o+W8t30W0vSyW8VVFm8Pbc4Kp
OelHdGGG5Hmo51Q+BsqbA9hSf6drePb81zX5AR2wFV6nMH5j+1AW1NY7vkT/lhne
5Yz2jo8niZMMDV5z2wmGzLStlOGj39JoDnTC9RXGjtKr7JIY04LGGTIjT3OWXc80
XfRFIXqsrJCrsD6RjwzgeP3xzrzps2wbLaKtEYNbbB3ORQ5x6MIAkLjj1LNRDs31
8gMCBI0xGialReKOGfUlPSknA11RGp4p30uKUYL/S/kEdGrl0H2/uB/DS4D/juue
GhqsKOcawNQSCOq0K9o+zzr0jhBaPQs0GNwsKNVzlMepES0430yNASxXekcq/9+0
HUw2fo1gonGFb6BUMNGpbeqACihYDDOZLjpPF3dohvRqpdqG0kJMnrrBGf+6XUkZ
BA8/tXNtlYGzTdJE4LDM7KUzAlZ7WHoJNSLC4gAXWYknKfne/71L+If/BdjdgNzC
GT6Xl3F39nOyUFNcvOcDEp7FmAagmPxwtr8cWnNHJN9+P9raaxW8bYNpQ8ZPSEXB
mzRNn4lUkJNr5R9om5RzwBLAgYWaf8NzpxiLfghifU/oVopaQUaRHmagMfY0Ey5M
u2P+Kcw/7aUMekZNYidNPWN5AJWvnhXmtd446ImYoSNywHPdPnfABrGP8u1iF+/C
5PRHPObpw78L44kMmKlPkM4J19ZlX7HbymYt5d+qKGwwM0YTBaS2OXIRP3izM1/m
odCDFpfSls86r03ZuBH4sRB+DbZKezBmYG24xORpJL8w4AaG7fUUhyEE/dnLqvQX
9YLVKuOTJFUYvtv0I/Qti4DCGLNZrH5SUBWQaGgHxlHvSofNBAZEegWLoNlmIPD+
CFZQ8K33UoHWb7QbGkg0kMfKjlCDShVDj6TMjGp5o7K5mLAmDMYPOdAfi1FTTQuL
aFM99xtZiHNqvcB+Cq6lfaZ7Org/IeEH9XZX6+BxRrKUXr0FL06mlHSts1k94p5X
m6kSZuk1HQT/kSZg+jntFi3uWjbpZ2zJbDBUCrF6W33jzkVPZfgIraW6p2tszMfX
iO9dD3+v++m10G3xEVIZS4AE2pJp27iCWEDbJuZhJ5eM2RAuDjdwBa6XoocLOcAm
idbHTy3WeNQQVKDPj0qKXmUVgAoAiUNggcCLBi2Hjt7WsbQiQ0dfzAqk7UFZhcRv
drYdeY+h+a0iS2SlfEwbqXYJtURqVq7rS9juUnfEwurjgJpIMbJthIr8+yhDPfq1
5zjY8jRpoBhfuztCHbfsKennKNZQEykZrFxC9HSdWlfEPw76g4QbI6Tac/6URu9U
aaCTQRlT3+1VnktfyNYaIXy3zwv2fPAdxLFvZYZhBo9RXoasQ9XQKvC6cwrbENlc
DAAL2SY2mjMk9gN0rQrvW6LQ5plDbAhhl/V7q8IF1fAdFQTyUtM3QSFbQ/JPsrKR
sJbEVxEQ6JwL2BrvN/rsLxRRAIVZn0KpFqLaE45TmeRsIwlU2HOfQVyyOhJN8XwV
z6g856euDujxksYQFmcjYkkuqnTx/u0oBK/e4L4CSEd2rZ3oXVGWWyHGfF6ctCTi
kOrPtXJuLvh11VLgpy+S6IYuHBlxF+sky5/0m7OUwX3zPauvf4LhxHKiO1pfLYwE
yMbyakpRT46C8IWvaQx1bBAqyRxdvgZ+OeDQdUQCZ979xnYPiw8gwlJJWfBXg/3V
IND3MgqD/dggov4r2Eh55Cc+saJt+KspkFWLA+wu7liY6Tvp4zho5CS+xe0ZNDFD
rhAHrE1hC4DHLwFyjpFFbXaE3+wdKxgJdumUt1vVwqA7U+hr5AsKjuh9VScWHnUD
yOjriu9ZLLW+vz90a2MV5oN5AMeEMZVQf2SlrTcnwtMWgpnFeNajQi/KO3mbRM1F
R3YoqM4G4nEGu1rQKS9Q4xj9TEl9ZysGHmC3AnUgCUaJzakqS3jkobTgjIBmpE1S
5qZQ6qm2f75QYgvooWS4rUuqYz9Krgg7LptxNvREwKQj162KcFht7e2PJjj1F6z2
wTQMpcloSXBLGGkqdOi0X/vLrxzQHizWwEvowLWU70UCn8+exz6IpXkEgtC3BLxK
thDLxzISEtGxnuTpJCNTacQtvtk5yCj8bqRn3vMXW97BngdEu+9NPZZKKD51e/Dt
r1617uKyOQPo2z7v2baqPCFy0lz9PELNWUyhTmjMtY/XoFvnPeg1ngMYJQEn7vIF
2uWHbGAMU0x1AxAzGdtnXsP3Nr/eGk6S3lwsosEOus2tAUhyRGWF4feaPO4U2lS3
LyaBQXMbCXtMookAWhp7WraRSl6+F0NvdZxqRi202Ej2KjOCok4WDEVDOwGUlnDm
GGRDTZhBth2gABJy1c3woLsNk96MD1ewyxPr9YIWc2H7I1B3nKXPcDvaK68v3xIa
eJk39olN3CV15yW6SX4mSv1eP8MvYgcXkj+nd9IW4rgN2WnaeHdRTRrAXXdQZTCf
OJq4yQnAty50SzZIY9qly88CS021RsZeHQY8NBqa0aA38D9OsXZxEhlkS2BBzf+A
s4okEUONsuN9JwObbUea1eqZKzm7PhPHvHohQztbcfJGflsqtuROzF+DhjkfDKW7
PD2fgf+ens8GK6/Q2lJR1UMKnEavHnaJYsF4jvPr9ozBE2urtQ8oYirQ9UybpBi+
+osa3wO0pgli7T9k9RJ9oHjyFRXP0Fm7HseCGF8+DSUve1HY1uFVuvD9+pgyKbim
ZefLqLkGHiVyB9+N9zhMP1kjwh1Y+eLOsE+q2Qb6u6WEFSVu/2n63mui7rfK6AM5
yclERWgeJA5bgzhdywb1xEXOnQKLxxy82goaeOa9TGCaaSNgx0XRIl1+EqSpSwek
/rXw8y4OQfXfGgPWlpBkb4Q6qih2EpepYB0DneU5ZvOgt5BkXqxhtKo3sjcyQkmZ
FTkbv0F/MKz21f/65uYNTq4/UAzlS9ox1xYnOouSwFpQj33HHMJgP2WzKi8miFYA
RBfv0zswUX9ZCt/RnDbqX+hBALNRnLpfzZKyGfhdT7cAvVUi6Z9EcnzM0FE6MvzE
qHtPfI6kKZItkIvvMR7Ut9QRASkUSEDQuQTaJgL7e8NWKjY4xcFwOKy3gGFm5GkB
Fx95r7ynbALmCaEOM0oCIRFPdxPge85Jg41QZCJj+/4HHjGQklYZu50THjEJp58i
fQFDDof0CgRp31UPAfKfXmeKelqM0HpfgTQS+58TZwPoxnxiDsvx93aA8bDCrQML
dzSvgFhAPofcm/53nwWu24p7AFZz8h0D2OsbKmkgZgGiziga+Ybyrg+VM/CFFSju
cKquXu04SZUtjAAQS9AXH5RV53Ww8+nDaBZDZbl4jAa4LUg7IoTcC7+5h43UMiHK
vhrjcmxU8x0DUWtM1sVzFxF38HR7zdYgLiQJdUxjcQt6O3vl2xI46gaAQzzZPtlw
G6BP5PLltI+k1DDIcIvlxyFQ6KadmVsI3fvoGnAAlovlbtmOKSuXfGiQRaa5DhL4
8wk+Z2hZzueSnFaKvsqOIG9gi2qPhSwA5+vAnteFfbzKekmO4doQaNA2I7Yk3iln
sUUfrReDpNzxr7zUJN9x+dh6KOeulexK9CRnF9XORJk0FcD1fawX3HB9QJ7wKdGj
32e9MF4C56xF0ziwGMaEQMYKuYlaC5NDPP71Mued9t4j9+M4lYoE2HK50glq+0NM
/0xO/gxZHTys5IdrOoCdXAEtOXRgWAnjmrkckkYPslIp0rfZD7nJxkms5DivFaQM
SiqTQaoxHk4RDCNOSFX26rY2VZc4Pjz/oqxwSPasVm6Iv0Y5R+BkliqX6/gOg3n5
vo/KaYwiicq1BPe4UghGTYG3KJM9Qh6i6WdHBsPtV++us1MbJlp50ybaiU2X6kGt
W3Ix4Q34IR7tNH6jGGNc+/HkyjXOH3C9aRf70L1q4x+pT64isnz5JfX/yF0PFn7X
WsZhsoH9hVvoj+DRKDVZ5XamTlBSVO+ch3iOzWoaoFrI2rtS13OfPIGzYyjtyxtZ
Mq9rLV2OgXTyXD96JhIuTmmRMRlk4Lyp3SVB0ruoLOHIZJYKfjzp8Z2SFfFYJVJN
20IntCNgAlStxzjZCcmFkcjkuATXtcvTP/c1ecC5VklnpQAUesaXF4z0Py8hIb2/
cQ2GtMac9qquB0t3M9gTdoO3+EIgA9sNLiheHsCeD+Ol3uf/B+eCKbWiVbVY0OrE
+enlW3O/RscJ1Cm4okwJ0gNzSdzmPRFkTnSn0I4Aft1FV8tZnULzEFKd2+P+HVgl
umIS6+MGPkpAFI6Sxld25FQvRKrirYNrrs3t1HVAjqYEO7+q+JLHq6cTpzneu62e
JGxCV7CLQPKAUQ7gmRRj7x0fm37YcDtvndiQUUqyR+0gnkVak8JvbPP2VHlGbbx3
gSaCqKUNlBcpO6XGXs9+leTsK2BcHnmjlrZa0a+zjfsV60Ji0VKXpZmJSwfKoBFL
tsuB2BleMarxqXhAGzkJ75wXQsaSN7wpfhILQaIbY0NMVI2xHVC08Ks5nJLE/Jbv
lwW5aBFAnqI26ST5nESEDsfL3lwwKGdbV8PfuTHCBp2pcyNs6Wcc3/jcA6OTQvoe
DAXpTBOcEF4lD2BFJHWDAEqk9Qiv4zDVE7vhtl7wBPmewSohB2Ej3wq4Ssa2iFWj
QyFv4lpB8aXN7R0b+aXth6mKSLV/JB9diInFoRGOacpOtRDLUliwEZgUECurBdV5
m26JU8sZtOl9LJxR3edkCGQiaDJ+NEdVqa8a7L7mgnklM0YgiALxxA+DCHfpIPdk
Uxn30WCTw5FjfKvQmPLQFySH92fqrxHecHAhBYDmXGddnK4ex8DsEJFvVxknpB2z
NKQm8j77NRJS2k8fJuebeT7jY3cuYpQu60AE7zveF6o7BaiusO5dcQwr7kFEpC7A
X28tQi1M1QK4ZgQpFZ/IeMQX5autrNvZMcAcaBB2/DIBaGzoJ8+AlqJLFX5I+oKC
/HI7pDQ5REZd0zybS3H4E/NdsomYm5XZwbuTsBxPVYzyr/5a8LHedH44v73Q4SHQ
jCgtIujnaNPDYoQ0JZYLH/mjaWsBsdFLSmIBO9BWKxQwt6wnhOrTvJGcU6N7rSNb
pcOZ47XJnyyqWft38D23d1eZjtU3/giVMB7ZxL+unH2t6nmlQTLFTI1e0MhmmnNJ
/P3QPtAc+QfVhdtikKAG+cFdgGPc0TOXfYUaKq77HTWxB4DbEs89JVWhI763gtL0
kwyo/aG6N2ZY61t/glGLcKINh8N5GlzA+1Fcc4hNNR3OrNPY2FlA7RHD1HDUbA2A
EiWeE0EUiOzM4sM7Vr1ejDFDL+u87OOA4niIypK3dOTiYiv/VL38lss0RgktMABa
HQpkhzvZG5f7/vX6zxk3v/HgtRSBTo6xwwLviQwJ+3pZdy6Rt8ifp/vhv18wdqdT
etUWpOdnFLcr+TJVMRiZn+nuVmsGI/P2qCnPHu+idZGw91i51Bz4igDDS0fCqbxY
b+bkuuSMpTU9ZB+d/KrVMxPGdviNf/EsqixbxQBRCHozeo5/92UfA8Hi3f+7jam3
b50XRwjwt9HW4CNxJp51odKLfaBYVXOZew45956bZqUD2/m7Ofyj7pZvgc5Fad3X
IWj2nKcf9dUPULVssRaeduI6BfBOFi+nvYopwQq1X+08KwBXZ5en5FiO2VuhABF7
wcsckDFjZhHiIci7a9KdeD5kJvekdTg4ftLBAwwPcIZ9A+xhS8RR8+aD3HSPsEXQ
PJgwQAAxCiezNs5eb/pAZ10ScQNE0mFPPX7fjgffNjIQfaRJX35kEQh0+syRXHoo
unm7+bZ4P3HGbncwquQg/qIdibdEqC3AWNoYf7trHl4ua+SnVjfev0hJyvCWEJR+
NaoHArjE1zzuZPqcv1xiQbFiCnoXOw8Q2ToBEHODNIDoqhNTW2gMdU8zxhoYwjqG
k+0aEiO0fp5qkAvusYne5/YXvDUq/cBDy0B2Tbugps/uqOc88TLC3xYrlezsaflX
xKwWTrZrljopbFFz6OAZaQlBYbM2dNFRe2+MFh4bSYGiejrxkKs7oeKhUd96Mcgf
1QuHb48JV9WD64QLDSy/oHq/QlKRvd9XndSKhYfKJ4CxZUGED820wjjj/xvXx9Gi
Anu3XzbvBUuEP/rSIv9kwPxTFkZJydmPq9JC1rQRLq1G2dMXxj32PQJkrrA1W+iP
77eTiMYkO5IpDhesVtRh4hemQfPy6130p7NJ0yZrLOQY4AZqGICEUw8wwqpwH/Tj
skRzVnrHe8SVC6BUtZ1rMP3lge3o/ekd3zjnBw051pia1ygG4tPeJXl9IHN62uy3
VaGLsWSokyRfP/005/4GqrvP3gQgRQov6LUpego64lBATAVlA68yS1y4hirRWHr9
i9HjuOt3DShvRCncPsjm+rr0Jk0UQSLPcvkSyxbd70ZcP3I2EtbOb2VSPWEqTLiT
usyshFSUb8m+UXH2f5kHknb/RbdgLIykvSD/n6q9yCIJP/I0J6RhiTCTRjxhNSmz
4aySXh0XwNqIJBih3qhht+CCbey8pD3XA2UIhe2ZSsE0shUe6GfrGzaWdkPVBxWQ
xQz2tetq3dth1pF4vHRn+pKjgrmJIcfFLhGBtu0wJ7vFc6We2zyBUM4R27sdNF70
AZFHQi9RC0nJ28auH3x4S+VuwNlaJR3bjiSAdMzCo5YJVEqU8YVtBSPYaw83wRX3
B/V+voBAmu+E51Aj15Txgq17WMTC6XUbvVTUv5sY3hMexkEH2XnPOhb4kl5B222i
0+0yajuJrVUwUPqoYJwp58TbyA78KFgC4mGZX3tloAOxwlPxqBcEhfEiYeRhk2Si
pwSlk4s2uRvtZNB8eQDUABjpgmg3vcg1HZTKQTil72V/DnsG8/Rpk3hY9GEPzuDb
wIG7FwdkL+DA0yKloT4H/HzHVRphNxZgZUVPADCbmt54vZtrompyDEoLOe4BdBf6
ys/46TN8B/J3cmhNEq8eTLgpArZKAreUtsJLJcjCLYS6CAfczH2oFWOfVJZ/Ydh/
r2eb0j9AuRtu0sgbcKzxfoNOUAkViV1G3G1dKRklt4RIdLeaQSKs+FE12qXKViGu
ic1nKTXsmjxWJDJlS9Btc6kzFXLQcL5n13c5Dtbl/eKwiPqtVSUdHu5KMVOteZeH
8bMes8LSTUMQoPwG0bH7GtFsoh92llMfqjLt9/mCppe5yLKEuu8mYrM0Y3EK5sCO
8wQ/zYtqqy+CsC+LIj7h3aqWS/YnDGSR95Zj0UR+NrL0Lcgj1JgtSZbzLmuHDcjw
LP3GhFhT9r6z+L0qiE9VDK2n1ixQAgFdV+1ZByeo5guUMEeUSxRIUb4M8CjJ50dk
iwNbRYNGQa9Y83R3LKtJySXS7AXrx0QYjL/C1SMfnQ4Tg+FGWiPvMeQ7CkkwBoJn
DQSq0pbCaA7btNM6B8prypo0CaItPfbr+wFfwduKujqoH0jPcBIFC447drRVz3BZ
GhtY0Ze5xB0E4Ci9yoH3GTglJKagdw8eSzmUa13KE65TazIMUDIrDZw3xsXCgu+o
m/ajdObq5Ajtme9mpe0lzxebxUeSFmI3Wln6Jr+9XLdINr6/DUYiytKCfO0mdzoZ
Aal5TMajyeCus7mE6EsB4aAyg6sZw3NNUZxBAPUBhDoWM7KMkkUV2KzB33/p5K15
8zD3rKEgbszepctk/4H1o0F2DUdQ9JaQkke+KpnJ4eTXuC39saQk3MkxV/lVRjPE
8WdJSqK2zxOx0t0FGLHNZTDsoCEv9lhFKWXZb40iw9sHXvG1/Hx6dBNuyr4nooi1
AztLdN4Lf1qgJAb798foy3DkUvnuXGxbVNTaKU3Y+tILl/1jgX1IEP7ZgiV03VH+
SjpgS/dilDdf78jNDf2KhzK7JzAXfQEwYxZ3AE8UNvM+9yT6OYMv2otegDEmC11Y
1BCv+r6pSVp1CMuKeVZVR/x9gbcX9to/aWIsb9zC8zJORKjE2BLAcemsm1HFfUS1
RQKOJObKSAKN8aRBDUFKT4MQyEkOrQ4n9PtR6t/t0jgotzljJFNxKHkGg7lf+kDc
ygFK012DYOOdEOdWXq4yZbw9sK6pJHdQATkhU/+bb6THjm+FmuLvA8aPaFQIYkzp
fQitl2Z9NLQfY8I1rXGTMgUnBnWkSEUBDinIrZFaOXPCUzfvkm4zuPsWfyOjqqPO
ZdsYyXELQUp2A+GqgpWb8s1kddvzGFoBalYDqEqE8X2nMJmtj4yneWWHtk594wnq
9zpaN1hDYNy5Hcm3Orzzv2UIVJV/MlFtWYrnkHohqLLC6Z7QjJRHe2NpFmzYtGR8
el3NET2T4P2P8n0NtJXlb/GDNHW3iA8JChpF+JzcdMGwEo34cjMAKAt7IBfghbJw
B6Vwea49Vk9lFsqmqxfEJzgDo5BWp16cV2POs68LE4VYNY5/EI+wvoQBssJZt0rQ
iAXHjdG9aM9jTzL1vGe7xsJs9Ll1S37m8uRdCX25GEJ5vrqofFVra+xopGRd269M
VmmTbbDYAxcCZfdcrks/Nd4UUXso/+uK/q781ud/tcZ8t+F9N3KksjdOgbQAr+Eq
KC2ApSrvEZcsqIAqTy/XFqKpPb418xumkYO/L6qP58L26+Wn0d3thLEQ1VLXVx2k
o8ANuwxYAimThBwrrwWW739nr/RmL2K8N8t29Ja6vCjAbIKX4wzYtwvnMdXveHgF
FhmUQf2KPYXstLJgzCWZpaD4eH0J0ka6yh6LEkj7/JBNtpNpimPDXhLU1qfDCGTa
qXQP9pa8cojM0LFY0jvdNoZ2p7CuRBAvWOyVZ6IUMjaihfb3O2bBzDm/4l7RyiI4
m9ox0saAa9bD2iAFfTkxJSxRRlUo0i5/Vva0Kq1SsWjyGUdlfFAFon6AIf4nEHMs
CHpBAgJBVUFPdrETjY9xyyt2vUYrWq+sxC9V9mwP9ED+ZtCCLyiJRC98izieFj9E
gwzka/an1OhkiUlKFxx44lBeJ9A7Ph1cUNT/ggocRwnpEVW4o8tsyOFUU3iBdvtI
c4Fdypq0ZWR68pJmci451JQqw0DaIPZHQV1iSmKnwLS+rT4WAyilX4d24WA4kuwC
aqM29yeCnbVNYMPfHbxJMjKz5L4A+GBSaXSxIyPV/AgQNF6is15QgsSYKnogX3h+
tCObkivF9RnlHaqWZbvkAR8LhzxSpkXeArToNUqgLqQsuAbq1zopsSrZgkmAxrau
UzIxkKQ1LbSKIZiD0CUVW8FdsN97ALYypDIE5A75yupsQzY5461o7euk/h2Z1+HG
ZHL0h+1LUzRoHqJnyoJce7Cnge1dywm56JafK7oZPEo4fTbtdTqo9lJu46sQ6EMj
MA7mXFZtdlaRAcLf8BJuRwd8YJg80xUSiTVj2IDuhOnilp7GDt87rk60PqpVw4HR
oCQJDBd4HxDioLGsf/G09jGZMYmFESpOa4i3V2uWTYQTjCjEHx86a1gyTMcc502L
2u1tmI7224gicuxoCj2Dsfb1Y6Y4F6anmQTMY29Nzn7kd9qgT6egB8EKAtu3MRMx
d6mm9mqU0MRnJdR3IPaPIoQSTtfuw5jlkaAF1hr1SkpPMoQelVQlIEQ6wT5siZhP
FDlm4pqyDJps4kWMvPekaNbzUmgZfWVrhA/gPPOdNviI8wzaZcX74iWI50ZuF2dT
8kO1dxWzYEqm7nMJo63sVH0bwQBoad0rTx+f1qZ47O/Edc4DpleyXSvAhaJM77jH
qc4n9nC9IRWD0yHZE3ORco9pPIz4RIIUrxoanN0NSkAr6BCU/Eu0nb6heUIcdk6h
GltgFiYTsZFHhR5YPA4kfUA6jBzzmvY+x7px43H2ma5luUnCxdHDZ918vu+3q1o5
P4cDUhqDBNa+pph4ZjRHC24kybMmNtK0l0FIMirYuuBaw1O5TjvZe2qEU68NmRw2
d1erTUcuTBXGrIboS9wXtpO3emNxqY/+ePycQc4rQpvHMQI4F0WoupmqYmI2iHxP
K5FJfnFRRpRzWbrwOs1eAD1P4vPsjqxr0Z25KGem27PX8n0ZQGa/SG31Zfmi687G
KyHCAkU+7Jeh3ijPWwx2fKj+XoiJZIbEGgDrXYcRCu6K/e7Zb8AeHtRFnJCI0nN+
iU8DG8ile8UdFlkZBvYexAHCvTzcvNSl/eTo0TGnBAJcRgrV01p6Aiy9of5VJmyu
40Ns/CRFEurUPhgEKd9THoRCcmI0ZTUHrFg5RhWIB0NRXWQdpmeCu0wovDG7k3zi
utub7ClFZ5uJQ9waZSHrjBr4DvT4Bdq7ChsaaYaZm5SV1aagJLxePQiJq+MEk6Xg
Jn5smSxIwcDHeqgM4UjhnIA3Ko6oxxq+gl0ewfATm/vlcvonuduFTd4zAwbiNKCY
FTSkIt8lqTSG3t3p6AvSEW3N790m2At+/v0K4uLtkflx70MYeSwnCwkOvRF15rbP
roAt1nFJilJmFS9I/DZu6ho3c/bx0um97XlIcMIP9BgiAVem1OIl7PlgDnePujF7
J5Am9S9SmpaoxKI+xU4/3aO2pIRvUvqNInSMr/7HvfBhxtx99QrCx5a1mLkJkPGv
lawj9pJd+AYBY7YosI878hHYvaMAOTFaYguPglxMk9nzM8AvilVr/4vOSqJCMEGD
8CwK/B5i4Q1wbs7h9zqWnQAl+RUoqevOuRnChsBPu3Cd4iFLg9XYG7LSq9DqcnCG
ZAC24n+P9npxbHyYkx9zceQb7nHJkwUxtsJHgzq4ihE5nnkRpP1jlMWFj0rxspYN
UnQAmTFscJJd2B4Gz4doxhZxk1XVlAmO5biPxO4gXE21FElk5A/cBpQKJ4fUupaX
dcCya6OwXyyp723uMX1kz2Zg3JR4e66ZoFozRWU1mMvI2tL+qxSFhaXB3TpVWw7v
b9dHx2I3z98z8inG0o0rWHMb82zUeh5Jz2vmiAtKTeD7TwO+1IIA3ku40ZQISf9f
UzqK6P5cMUvROgO2gWjEZxUifn7ZSJh+4eBw90BM55WKiqW0SeuqX24neFD67GEA
nMoByUFfgq6l87oX6aXK52yhoEYQd/mru6TeDQRvwpAqT7+VR3HsiwkJ0WYwywei
jJJlKTnTXfYb/GBcIB8U53zsXeB1nAWqMJRMD+oUDRovBNovM1jhv7ZyfTkU+13Q
xlov7E3D8grToCy52/Ielm6cf6MtOgCl+R6KSREUxE5jCnd8pnFkfZz84QnmBcgW
1ubeN9PI/m5Ttu81B4Mwts8VMNFnBxmkBoFgzHIjBY7OXipNb5wrQfVECDiEYglJ
nccgWNpyqvz2zHO8Rylr2b2D4mtSwydWTnkerteHoxzRfTxxVnM5ERNuZLJRfGgx
pOa9V6g+K1q/vzBUMZKL6Y2kRvq4g5lp0AX1kILUSmlM3EDrKg+v3ZAltp4xY1e0
X65sXgsa+14r+z8oNjWG5yc7AP8ql8EHGXtO/InVecz2NVTjpr4mqgzDjCEuRjWc
JC12MyEWjV4TZDV6htD+eqfBXNDKzuATZeBjusjQnWTJpw9VFQyIqoLKyrGmnmB0
U84ThNcqlsx7TTo+pt1EaAb/3Y/4fh2peAXfM9L5YV5x+oSKxNZ2mUnWstzdbukd
jTKHC+oQuyfx7FWczqsWD6QnA9U/VCeBg1cjGsxu90O07qJiVBMbEjU9Q2lS6L7y
L2MOVKf993T16tCmUiwaruZLz+ltzFuiYlKepDJsMceDOcDzsrPRn/EalsUHLiU0
UZqWST3T+sPBBokYexTCQOGDDDZuReZnSjPw9oMsBIb+o3li7O/LuvwhQiIR6VT6
lQUCLnHDFmjBRjnktSoXbeXL0l7pdcIA+ujotJ2fflLftNyOr6CSgO4g9O6qOQcz
ap4yjSqGCaqIebHlaqsAQK9hovWJM0IpgMpKycTLPYgwxJymJuMpKq8htjWAzgYL
Dv0KSRYSZjSqUusC9liSX26Mt6fLVBhY+65+IC56Vvu0jEJdwhK3axEbWK6zoCcV
H42SUJog9nX2p/RwbCQY2Uj3GUp+PLYo8cb6AExkLLLMf11qGJmpdkICUfQcF8Gw
DHOAWFt4Ig4iZCfVklWyi5n7HFfHxiuIC0v/VtmwfAfZrRG2hEyNYWBpuzgpRu/B
fXEX/c9pEwM/ZH2Un1M8GhkUiGGps7aI+swLziPrm56aTE6qDvwJjxHczr62EIh7
WX6U8Jviv4UgI6agV0JaVh1OPaR30E+5WCQcvzWfBUbR8CcHdsuRgPNdNac3I+OM
dCIBMafoTeg/DJwN0+lQh4xstHrqj9LMOFNoH0XE0nnKxqnnW5O2m+t1zTAlk8y0
1CSE/DplhPvzrpUXK8ZB6datswu5lTDjF9Sw7FW3TJBakV7PUPKGnexBkuTEjXr1
l7OwRPOGNxGa3+w9zE6Xs+DR7MZFp5bV/okgYbFw9/Z28O66jCQElEp5UjMLOqBy
zDt77ofKnjSK1WdihYu/cW40Kv4QeUBBAaXmrlE1zT9G0sGcIwhbMGJ5oJnVHENh
OyCPkd5/Pgsgv9aDB16/0Ua4TRlDghfxsLIjdwJbnQLUpFJ+3Tq/4I4s9u8zSrL5
/NQOBE3tK8Rmi0mYYQQ4fpBYfJNXolX5Nf5f8kNLc/QSpii6WtaUcA4MZAUJm2W9
n5eUH60MxQIrTkL5mUluPg6C+IPwbjQY3WkkJGwZaym4gWHtMmFgRUIqKFiVBYZ9
ham7il1ZYUx7EUd1OKosT0Sq89h9jgSP3hFupxUkT2FA/jCiLm65jfq1MzkSYBCe
oZWUVMAzvYisbfUA0JQZQSi9XhVqkkuc/5UFluOsZqfo2UypHEwek1FRse4bczoP
4c7tBC8berVZojw70E566eRNjGArdhiz9U8kk0TtbM8GfZMFU9UZplpMaF43u7Tz
AHEnotkDa0jx5uehaAARuFpkmnb3nfq4DGF/AVj2+PSM32bv6S6EZYzr8v47Ry+A
tBY2seGesbdTRxajLjrBQ99RxP1CeD1f4+YziWVg1l/kqAWheENIoxK5MwmpFY0m
hN/j9/GNW1gk1jI6RM5k+02UDTFhmQHv+/4fuBkbcKEDAiuS5Vtec6NVR1wieOkj
fLpjq7PWJf5Se3t+SAOM89VedBYg6hBz/yLTjoRV5mYNxvcH++15HyNYbdHQ9BSn
ctRCZPQbTf8B44z5/MnN/ePOhFRuLVkvFDvBXm0p601hXI5wu1V/CEk9vPFMlC98
rI1YMpM3sHN980mQ/HjZSDRgdGt/+iy8saNE7vFrrDDGxO5dfELqetbqazAUw2gY
4a+4CuLPWyjSKzrlYTCcINHk7JSkn8zt97ntDaJUEELe+TFgTR0bHi860tzgW61K
w+8mQ+alrBgqoB6VjpwuJunDQ/XLc2A9kjIb/Yi5T+2Br7xBiEEuO/O4kaZOBO4q
fjI3GJtlG0jUEnZ0sr7/Q1TQMzEK9eaWJEnCAOXwxeyxMK95T86I76FhEq/dDHtJ
mt6yuvS/8rrZ5I9QuvFeX0ziOLZaGtUdl1GwA7W1vOJXP+rT6JRZ1cOhWTCi6/v9
fBRv6KtVk8bGECnOCy/ZPTwAkAnluko05of6RD8/h1e1hJ4MgHoh/7LU1rd9iOxE
o2G9PTCekUsaQUn4DLXSnPMU28ScrauxFkUQSFQ7unq3lvWAhbI8hLvF7eDEZvN0
TEmzvJAINpFp1M6t340/wxo9VIk4s0SbnliOsJISVH/uZbRuvfJINGLTBYEupQ+S
DT7SMw8AG51Sa/01Pb0W3H2k8Ed1HpRKi8NLRhEbwlhwxZwfwCohxFU69jU/Mz7g
sReop2/GYglwpjy5opbto397E8bmaY00sofnalPkW8M6HTWVu/vXLihRNHhZES1U
eR3RVEfEqjo8EbGR+ujJkvBhZSNTmMixiWPMr5RWvsebxWJ6CvbE5ob+6HMmnwT3
cmfl/deK7QttZ86q6lxxyDxJYK2riKYx04s6mraM9sS7Jhl4DLt4Rx6qmvPQwVbQ
XGv7x5wSnNdzWJgv+EKchKxUV2wFuzugVCqpIF6DOmx+2Avstikw9qMPM98e3VIH
jdqWwOGf1H/yZiUsa5GUvFseME6TrBvaGxKPFzlutxCaajOS6FItnfJIFf8R9wNG
owlSdpMQ3ueRNOb+9l0IEivlHBxlKzil4nKu32SlXwFb7HqI4ZdRR3ktRxylaMtb
zBpoXxkLp1PYi+7i8EdA46xvoSYAejS8PpxrMuD2EGXwmBIbd+3i0fOZRFXh+Azz
ccSlV/bcQVdCLNDvMFkUabmIln1e8hZPF69irnvbbxnkQponctCZ2urviumpz/yt
ZJvqiBLowGcM34cmdxAgjzV40Lg3/bSL736eCyUtHVjhi39NhWPg5vheCzal/AC1
lw5wWfl6E/zMg3F58HHqT8TLd+xzy6SuxaXSyN7WYyf5cAbOQxqRp12w9GE2nSHD
LllNhlELm4YRBbbc+r82RJU3nNedEDxIGkmSxRYKX4+Tm8imStXz28aWPr8urxIt
1IUtoADcUJVvzt/AThru5gIJ89+qo4803noZ/hsia6ql6cFlKhJVWa6DYKWrgBx4
J8JBFTxZzobtyslN/2woG8Na25e4iKdjZHNrZPJldqOsslhNfKvRdsWQY+K4d6B9
GzRKh+rFZfU/viUdj0KuE8iwji8apBaHmolK3X6TJsxxf+jANAM37J7cN8O4gxXA
JxiGQoDYST2S3cSBP54BoVvPojN4i1/Mif2yZvAhN8TpTTCw5zsSAekuxzJIRuXz
h4/+QjorkLgUwU+4HqU4uJWZVennbrs7K52tIxqSpdFLcwIOd8GYsQLFkwoTeYue
n54ZW5Cmv/OUq6gQiDsTLRSHLXCjWUHus4UDhcsLAH+cS8SGLmkBe0ub2+a3DkJD
b3Rwcp264T6pjwJ3oeXPgduZecs5Zh34Uk1ynyNCmv4sk9HHLtOHaltAurrUDD8R
468ZtpYM+vmZ4DS5bhZOjEdAw5lX/vJMwXG3+guRCwRCXLbLi0ed0NSgz1WzbDrv
Uf/W+N6W6lMdUKPKNl/CmR4RGbAfuS+zl74+GSlp8hmZzIn4DjlSxBkZtYB9VOdO
0GzFso3Z4zhLaieI/k+OVKj/pJMdDwlEOR0E2NeBDuvMX/ORnZvVyw1CMEd5OQWB
WDb6qRZ69cT7s5p6Wo8E85pD/XN5OX0UJFEd2FkQgXCUjGOp9nN+cv9gBnjgr0VK
RvA4F0zgtCg8wm9l8gKUQl7S2q6JC309Wm6eS3mOGgAzJi2EQAyPPS5RFcrfKTPh
gTSH7O42+biSdvDn3Csb7yhkP5FNjtNaofqMKWhmXEtq+x18eAqJhBIL6iRynNKM
d/jAcbZi+DEdHqIjfqHJMZPDb/3jnwirPL+UWt6MqcDM1IR0G6DdlsSyNGcFALSk
J1XD308o0aRBJ1P/l2CPmpp4FwMe/8bFCNjQsP1rA2/GUUGuZDraLd4KHsRw7aOJ
1TVGyYwda7tLRHiPBLzPFF3ObLGTizd7wtuVY1yPa0hrRY9/tUBShOqHMpdcoSAb
IuVixvsw8n3ZjS2mkfjjSNCBl0z3fhu/FaAXkNTBdZTCYyPIA8U1vuLZSYs/IVED
pcA3ZA5UJ580o6qzWgauA4vM0FX6hcJfz2Twqv07li2FExzo4wd7ArrDMgnCULnx
arfdANspEp403Be0yz5X8iyhyu0L0Nb8rpdJBiZVY4CHgDcj9n6aM4aaB2Gt1CHp
5FpBQBG4ahHjlLZFxY83vtkERTOu16vV2ZH+Z0J33aEEU7ehUlY158GYBeDL+sC1
rLEVsEhKtBd3OmOCs4oQBqjbGd5D3EMNfabbo+pGOk0An9NI6cP0HBESH9xUY6mZ
rcgs3ENcdUn6e8cOiDjQzXTJdAzA74wv1tSpulLXPi2bKzXlebiH60x00C6qMuDa
Z5P3935Ond7YW5U4zslRHuCKg2KfsPbcNI+SDXJXsX+qcLSlILwehvhxZO3RNO16
DK8AK+VlNdwnDF3SExb9SCmZIrFMo68Xrb/EZ0agfqB0j8V526ImOeJOCTRyBVwh
Cn4SCfNFngRxgdFoBojsv9AwrJd/LpMjJWbWstaejLanHxlu0lUwjeVHFGBNuzpj
Y3JPu1IuCUUI3qGxindyK30z8pmkLaDpUxiRGknZ5QLy+belVEN0hz3cKF8bXzsD
jYm2UkO0DPV7C8d8tq4KiteOEzl0OixMr53tGrry3DetINO6jkbRje/CrogOlUvV
7Vc4CskRgqMVXx6Zj+EGnLKvYSyNsc505vntR7TMSX/WX/Dj+ZWREZwudgw3dGq7
QWAeTE5CvCEpBrpFixPQpXo0fCILgvqVgu2TBqTxFlygoEKENP+hspbDNxHuLEc3
VhfVej5O5bnPL6aJ4Ub8/cBsyTSmdPPEyw0hucoYHrLD3kdbZa1da73TbbNQucIq
d0PJcH5R4Lc4OIWAFqHkhwgh7HtWD9X6lHxyrdXXoV8PkhbzLefFqrbYlqDYvKe7
dlMchPcpY6I6znMj0b9r9oBU6bSHS9jyDiMqleVVN6hN4mbu36sbs6aV7o8LnopB
i2kxHThu/xEeRIQ3fvZ5zShM1YFgKUs/7gga5S1v1xm1FwgPzCrCvoMAKVhY7pZU
+3kcAW6pbMkSNKmjnXGknaKevBZB9P8v9YYgs/YqOjw4wYozeRKAPwkIK46xaW5n
Fm0In7F4sr8PQGHVovEOt2lI9F2HhYYw2o4JUo3mkN+iKerYKu/Qj1mcZY+qqOaO
9TcTU1dnXNLBdQzjEW7Qz23y8/QWswlsj4l7fYXPRkdQN6AhE82Hhm0FS6Fs5snD
L5zLx8erMRtgA9qvvtdSf4lS02nK3HtUXCFCgv9YteoyG8hxPfjGARz+n4iQ+3nF
l1XXggH+y8KfJn9fuSTKuAEVX4QSQjIG7xYlSVSFbPcZYzo2jGssh3GrVlGlvhst
nF962GPOe8SoL7FjL7VErYVAfuvRERiOWaywuTx8lABMqasLc6CgnT7Cd0cSiwDS
mxsrTY8A+B7VneADjmxELjYEsJfPYwfQCotvG9Y8qo5x+MFZTgYS8NHp1JtODcVQ
nIS4Xa7FYrviB72AxYNQpjKSnq2SCbx6uhyGaXCbaFFluNpCjMji7lhfUuE8ERED
zvHU9eHcvH3nrq+3i+23wnDX0pAZByEYuSnMgsVz9YbIG1kFUZbCwKa64KSKeTO6
8jfHSVGwheHZVHglPTO1Etcv7XC6XOW3a/YmV36HkmuuFOZr8DvKIh4TGA9Ri5Bc
5334Us4jhhpk0lgXm9JwKWMTs/n9Rkoo3ZBCsrtfjdH1x9UqfM2v+WrmvqVckDLE
6osRBKUO8EtitAXHIjWmPMdjnJ1LTG2mzoRdU1XKxDz6TxC0c0ETouq+LiUAZMbf
ADr9gUdtbzxFXXVmTn0UNy1vyq5tpxNlK+FC1MgJsmMmB9URa9IKwCrfqsf7pNXJ
Q5ABENNgGhjuyvW/cL6RXhgbS2En5rbTj4E/GgJKZ+pozxTZEI1keSs7JfAhgW/e
bcBvSg28kKL+b07rAyfF18ROlvC2w6FGg5LGjquERwjSBKHcE8DBQCHqo1pEpxkd
nB8qGQ3/9MvxlSFRvo85PmSLinZAjY+LkRnH9LJSifl1y97K2TQq1MS87Eq9fFAr
Wt/6AZ+/pqZec32TILpW+6V3c51xDVuFjyX8L6BQCwJaIX9SQqEhwcZNvkieSp0h
TLJ8qG3VXpzfI1Zfu4H+9XQ9zzuR9KO2Q6R9AyVz2oQkamgcxkkNXdf9w6tzdNRT
QP7L3LwvCLPbfSAuLgmRA4soXoMQO0TktEhqK4NsPzZ8lN5WJu9puOg2YT1Q3PFc
qnNbKuybQXjZg6zD1QqlsC1UL5qrUKhLsD+j7kEHlFdtzqWRrII1mU0RwVJfTSLH
HRPhIiNROKnM5FjXz5lqzkgT9CkqDl6i4TCV6Razo/USTpguFYb756zB21qzc49e
KirnaZIfhdgCIHW3h/oE+cDnH8ilUW2hQuiOX9T6NfauZv01YMtLrd60RVMlJ24G
LyAsHWxXXikbQ8IOceopCT542LavraRVQs8Isk+IJXr7SEgkI0xrk8Qt4GyySm/s
82e5b5wa5sfwYFAK5OYrDImtW2VCmnOdb1LvDncmEzR10MKofbTK30/CC2dsgSSh
zAOs9B7NkDwL/4qIbG1jj1BWNExTuNSi0pzoZ3A1gX0JVh2VMKbAyiEj5SjR8YHy
TNbdonmOKDPlQDkb4zva4gznVGeRE1KKdeH3btyPswq+7i3RED6yMW7Ph6i6mvRO
oIe4T8JI41IqOgD9rdRz142cXycfqbREaJrSygairEvVf7hns6vKV4FNKp2H279S
POzd3rqP8BDpY6+y8tMZBagwtlMzia6Jr8BE64fmXJ9tmW/Sj98JHck7Z+gmb4GS
EVdKYp1d6nWRRhDgf3Vg9PufqB6bc5zc88XrQzoNhA0VnKLTYy36M/o56PqjV779
Oz46qRUNP4Yw3Z88ODtwNeVM9e1ZzEG1pQclelkUMzuBe9aLQjyATWkmkgaaVdO2
jnqgkUUaFD8cOIzzl6mksapZPrQFJ8Qpgwde5O3FZKoWebhIO9Zk+muqDvibSx49
s/Qg8VQAvoFCbfbCYztCGqlds466twHPY48sMUYq0vgqzqJ2k0RCw2w79vpyZbFw
NRNt8ui1M6pwxpQdCZsk8RARia+S0EAqW5E3EYrc1jdQvp5pAWA9djORAlK4BQvX
zSdP3Uijv5NsEjECk1xwIR/TYxtu/qKSonqb0WXfy3FBmj76qp+jJ7+MGZvDYACU
QeSj3NdJcLRdEj1ca3xHfEFtHdZmRA0PLGGFkj7Y+8ayVszO3CaZgUxfOfnmb61n
k/u8bzIGK8Irkq4P0368WjTy4+5RwNvG+1vY9eTRrzkZBW3nz18wb6sJy59tC7yX
lISVfeCakLL29R8NxkxZVnxxGahkHYKXux/5uFKnz+f4qhM6X2cT8xOB+RDRSPTj
JXVG5bim1gfpkAReenSCiqx4wcLbUCgE3M6cztW1qb2Q+ox/Ydd2InC20ugQHSvY
rWpxfP/gzDOl6jpId5yJvaDcPQVeD9zgAU1zlP3JvnhLLNkdPSraVIS52ybZVhn3
tiFidGkSmW2TEtk2JOCJ2KxywFZj+w0aevSs+GfV89VTALF8Zso9TyZUebBTz44z
rwSl+gyxQ50dzXlaNdRYRC1ZNIqgAyPTdXgCT6jh4ZVlAWPMjtgztOwQj33jMa0+
jHwzInRWPHCgYAi/eLfcZ9Ua5yOTR6zbCJ+MlsA4XEKqImQGo55HVUtNlk7zXqdP
F+1sS+BX7ulGuiqD3vkslPvV/s0Ynzl5xU4K44oDT1rf+WcVIb8JU1Lh7jfd5iA+
jMLDJvxPECksr4rXEUSLi4W75DDN9mxczXD/ARe/RnLl5I63gxhwcf6i8Emnkh88
oIYu0luxmn/60XS1ysj8/Qp/eNWfJ82W3XncY0E9+59AKfOJCNHQSwxnUWPr2Owm
4Mp7bY6Q8SRgoifugabzEcm/xDILBK/Htgxf65UqWsZuh4SfNmApQ/yTrnzTWT6U
OmQFo9kf3ZjI3E86v4adVHoz2mjEkpMMaVqnQ0T50ccTRp8+PsXqDfRfa6idUatW
LdMDgMP3JONwB10BJ30VIhj1//pA6V5Wf+DzXl/MbgFU2SGRR1wmn2TUotdmR8Mh
OWqj74Z0KdC1rOHyA3ymwOhkYNnZJ+X8aRVadoyM8kIzPJMrHXBQaCsED6BI5d4i
okt4a0JfbOcrvl967R0dKIx9A16PmpCEn4h+FfVxv5QmULLDly2C0TwxLnNAnW8y
iAqOL9MYNm50jxEzqFWHpMxs+L1wZ9C2TJp0h8FewV7t5/6amSJMfwC/0O5jR5q4
h6rI5j0bq5WiUvp5NoQvsM+lbU2k1evPY0t82T7q3gB5vizK2cf0jSTI/xguHg2D
5U/1h7UySIulUqEyATEOAVw3dZd3MOSzBtcKZHmQYwfiotVU462thECgfEO/3AJc
3XO+T0c6h8Ht8rAylAziSf0rjwOk1HkEFMZXCCNiVyjrNEJm8FEqZGZo0oSXX41Y
quVazAiHHzi8T/N6Omdn/DJzzRiPZt0/gfJYkXQQyLi7IAaPliq25gT8iAmwZdcp
IN9TNQmay5I7Ua9MpmcDBpjKTMO2kINvXxhQi98TeqCLpoI3QgLaeGGDN9Rc1/Ib
6MLyRmkmw2mQXEpg5t5gOaUBOGOIVVhiP6H0yp6QK08jPjPSR4PQxHQnKvTM6dcX
h6/XFjgEEj4AdUDnI0vxLSNUHOwZ0xb6WfndbCVq0eev9zuCrHxUdnSEMssCu0Dk
dark9FPq8sWlAJ530xJgYzfjCjFEpKKIaHITPSTnShhvGps64jTSXyIcyC7AT8Fz
+hKcvUZLwSVdlKxUh4HSs/+ENTVWjOBMrpN9pkDP+PpLfgfh+WfZA7DpXqo3Dv6G
8zZZJwG7pdmRr2OyWHbAf3FvDKVinF8UqXz1y6Ogtj/QSZTOd8tnQ2pB3VZgylMa
8S3xQc56zIsS65zK8+4HW6SVEKx24FNwwJQZF8v1M4mPk5zhTWEinuHBpsERJywc
UPWY7DVmfJ2ZS7eB4iUbMrALj42ISZ9xph67J01If6yZaZE97K3oOQrTuf0uxTKI
qTBbIAC9SCdDioXtmPv3spt3gnfsXYFIzweBDF8t4d0Z1BXpfyhlKQ7zM+SI4r0q
o0pr7bF+E3EAV5NxdxRhuxQd/15V4gAFr2egS83Tsx97KHs6YmOrf8Hh7ioaMzF7
GduOQJLLnckZXcMej6zwgsPhfdJBTYbABWJ9BP6nP6nwB94JvBlmjfu6u62e4qdl
XfombxWzVHryt3hCnEs+iELo276MbHonNw0JbnQqqSRen/JSa0SvRtNLk8bssyj4
Op3z1zoyaPmx+NS5RGSZN566CBTnUnk7EjKpKQqLKah0q0Fb1pr3WT2TdKB6eadu
Okemzrrh3p41DHT65ZjzSYzp1OR151qpdd4Z7zb3bI4ZghIDO/qNu2hOFbKZfsbW
m2IuSSUZTRhReXg3xHZ9XRyzjS6vvfRl3jvAjMcHZWLKyrdxwqvZDICxYhsN8R7L
NTfyjBa1TepV+5v73pl1LG0lP7D8TPPpW2IoRbMeuvbn0fVBjPTvhrfbDURqVmBt
mNj9NbQyJuG1N6gom5swcSKpiLtTVRWg6UFWS82R4mJBmDAiiCWfJW5t/8aMplwn
Bep+oMCVupHXkvnpSfiN/C2H77CcaMdMZBZCpNykIkb9NHZV2BYWNsWqQikp27Gh
uTth9RRpYmhJNzc+nOnldc0DsXp7ihJgSQ5smsCs9fndtV9Enc/xS+CaZOiIT707
hiMfo6C6xLUs6AVynFMMb7/jyeyb/zF+iaox+OCrureAgPnPrtBOOw2eI5pbUSaa
WZvI95ipo0kYHtOybbaXf/AL9ISgkwiiet5Hr/moao3+eyKNJSdTYlg+60g0hRNY
MgVGIfBpHUcZSaEN70QhqcXsPGrefSR4D5gRohM/UkWDBoG7z3hJCYZY9oxU0C+D
yb/a+bb9YMdd3ZqnV4S3mHsY4Kt8aycNK/xtzOsfi2ZJVcAgFn/7f0mlRz47nfAL
iyTUpkNoDYII0tBdgU4uuEEY4SZUZ508eWjrUKovhIOgbWF+ZYU93mJYsYZeexWU
flcY7rTInmR0SG5HkV4Q4GbEdWk8Y6Sxnf3rNoMAU+huLrI8wWfsvmDWTMsrGAIU
atekvJaE3ga6Kbg8N6XQJ3GMIhBWaWFkCXhEBbr3Zhen8vIZjghc+r+X6BhlwwiL
E46lhpW0Do3BvI+/3jX+lKvsn3zFEcJY655KqglZIMdTnJqULdorebLUBVpHthLy
gKesNKqW3PHkn/jv96/qY2q4C1w1CYNVj8oUSCdvtMyhfAt16oApRBzKh5su/iOd
/VwungMIoF5allQmfwR9I1G2jk1RLlBklcM8XNg91+4no3yaAXVzEf0QaNYL7FDg
1GP1uNnp29d/bT/qEnF62qsS32S5VGBg77S0GsAVnEbQ9S3/b2CILEOMsZzz0eA5
iOExTpA33Oq2UNWGZKADlyjPjokJ7wcfOY+BszKULN94DHlM/2oX3CxLp/yG4tf0
54UkcfodDtEA3joadjW0sbvMzwW8Opbjcyk1U7IehlI6g/370lMpicEgFRwOd8rG
PhooKjw3eEXFZPdL/wfdLYX5tJjjFJNvKP6fuPlUo6xGcT7EaNkfo7HSijReA9IY
B9kdlQgYWKIlIt/fZiPx5qj2ZMMqwcwc73Wd6BHI3WcfRh3WdGgGX7ugpJc6Kbbn
fQnsoi0Bo2x4PlY0Z4QLcE2s6UAGVcFm4CK5PwSZ0S1GEvkOP8948E96Esi2galQ
sWG9qr5eD4rivvzsL6Jbu2nBzZd8SnV1F9GpsyRNfp1Lorc8A0RjVmRO7qHqWEjh
j3GAvUcNrV7ECMg0Ys4FW0leEiBJkz8qY6ymNabjPXaPOUVadFHUVIUS7vLvp7UM
bgVTSRXrr9QxNW40jM/lbNUCY4pIIbIdV3g7r3sx71Fs3G/a5yUjiHbddz30vxzo
K8WxCtkfUcbkRzF8LWJqYdB53TjeEsAfjqDK3Wp2V9NDsmPvAK+23Gv9m3+dDD2Z
/D+LTf1/ODdoK45qp9B5xC2PEDUNzrFxSJbOat3DgifPZauKWqVYNXRpOexi3Vot
MgA305kv6NqtXuUcM29yOaltDebBCcBf55jFbFRSIBNSsBxdG1/mhh+6kqRW6EOf
54t2k2plz3yqrK96UM8bo0YBTBzSv56h6M50t0CYcwO+cWggMaOrMHvqvYshbCYx
XUzzCf93oGu/lgv9rF3rxSM4EZ6/q7jKEePemzKK2pUN39yTSW37go63sVgzQoUL
/YeW0X9cZZnPMU2KWesvNzte9rEjkwR9rDnmZfOVlcKo8GlS3D/DdrsZcVJBTs96
SNMGOx62AwxNTG07JVpmaeG/qATq3qfapVCixIvtuIdoGAkHjzh+bs83O8DycoV9
HTDKIRjmrlMlGgbAF15nL1qzxkVUaHpsZIfN+bJSbWCCck8CPOvPkaYt5H+FmVjW
RzZRApsjer+PVeDpyvzk/EBewNaFN63cVllWSl/NtPpsVSIN1vOQNndlsaAWI2V3
WEXRwe/GNVdvHaG2np7WxCN1dk1t8ichIz3QPo6+lmldGvhShsKljI97E/LsNc91
O9fy6OP3iX0Ba0UDK5/nsP//FpqmSQOvhlBIgoAuwFzwA7VV/CV7uXTe1v4bPWeI
SgUnqg9ulao0dMxYXpGF84IumI+khdruvpxDYTNg8MsdJyJ7tlUqQCAf9CWc+6Ci
a0AluB+t9bxHABv9ZiQCo4bNpRlBVBekCnlpYcPt0jV6bcBchhYh10zHuu1BPGrU
pYXfAA777YxEbRcc8Y1oqSyUwWG4VyKJpiy0fKFCvwYUybi0saoE29WUzrFIbamx
+uPnUcDyp6l5MjEVUxNm3Gmx90UWNWiZO4mzSFIlmyqwpJWnKsO6t5/CL50ms2Eg
gfwPoh8BZMML5MiKCAS6DsUZVc6oyAIs0yXCdbf8N/GeSghjOpXHGyt2cJDnXiul
sHJ1KgiIJ4PK+1WO0KrrxNNCPtBlbG1rbU74ivWy62rS1Vr4pShJDscJgQBgOLmw
6XfjDUITsPstkZwcVtZ/DLLOI4MPqrLPF4cCk2P1y9dEoBi4eQTMjIGcJlTZPL63
SQsAqORFmvuDmFk9TuMK9XanNI9TlBdnIi+UwczTie3u6alYI3m2NGh0FzQjXu8M
gMVKX3LhPjACS47VNydoikzpjzqk4CZQb7k7UhbvMgLqjUt2+SoXb0lYUc4S2EcD
44mmbfGIIoEp8SljMH5R7gtC9NMg3tlfVC2yUzKVfvFOJXyHkus+OJyFlKOq+Nk4
OM0LWQy2oZGYYkGgp3+tUdROd5X0Lhoj/nNLFj8kEo3tX9s64EI6Lir1NshilYwP
NJ2gnmOjr9aNDuJ7VjqARS5QAriXs4aKePRleMCmDbyB1i9SYr3q1cxd0M9FhQhV
9FF/D6UqSPT1AsVDTwKgGuFO7aT4iaVz3n/Q2uvkOOXFmCl2aCDpEvy8X41NHQtJ
mMHDbzRaBnHdmxWxONbhnVC9wAfU8Y9i7/9EhMi56R/3bEeh0a0MhwVlqlv/bzfR
E9Y/NBWvfMh5aldSgAEon9gCSarxLZtc8Dyv/tCUdsTzLD6DZ4r1INgwLXu9gs9C
rR6IXSudWu+M1bEL/eAsYk9Wo9794XhsPaC1TvSy7C5faXr1eKkhOk8Vk4IdNfHv
pxpgeD2TlLbykeTJkPcPurB2CjNgco1W8BGmOqkk/9lUmaI9TfgHNXGgrIdwpuas
iRUVQfer9lpcHuHIUujs2bd6G071zL2mwmhJpNMsRWiy1BWudMxxFAE1jZ0u6igV
yfBbd+CHFhMsPYOp/N16JRljIuxHjQDblb4Z6pTvDmCs71UDtSFrpDdJohCB7rKt
YbUxVWZFXM83LoYAr8Q2u8epryo27J1mKnkEtDiF0QsVYo60XXO+kqQaGZkbu7QT
9qp2Dp5tAnekZMC156ocuP4G8n0Ld1awhAJICCf7czjGPESfVOw/MEvjNn0/Zz7I
CDET58qAQVikcpAZJAOfc/yPsBDfcFExnzZp5FvjPBjkz0jaJer1npO76v9DPEru
iNDg9XOa9Pt2gcXypHpbhOVaDJJg03I/TgQb9UMpbJObUSoRf+wz6Yrs64VjcTm5
RRmVfXssSdt7GSkQ+3pyi9Ig4wEVa3U+nK9nws6x1+q/WkLoYFEdSsQQJ43epYOn
zaCcmMQQX+XNPdZ080YmfhE2HXU6ilQaxwg9zM6N9iVXTsYGS4GdW9Ub+fRoVfrD
8GV8R5BbIRCXXH5KbhoCcC2p5b/BrXNNwndzsj7rR9q/SDgl2xgNg2690nKsmfdX
zN5EDDvj1Edw4JhN0DmIjtFefDEkjqOjfo+iLK0liqoZldQJH41l+MTr4klzTCk3
ovVIH1mP/DwqkHJMYbblkE/2xDO/6RRb3Ex64tYe6TcKlZdg/XvduaF2jWe1mfBZ
2VPe6EfkwMzBWBu1UbtLDUpXVCOOduSK0cqXISZBusGfNUjIJ5zB3tMQwkUWuzft
MZwMw25eG1xmNrcWAvoVpCeW/atsjA7DL2y0Fin1h2OxitZp3MXKa+9SSblOhqor
Lj3y0qClgu3zctRv6jjcAXm775j62TBzeZbcSpjzcqJwDzDv3/ioO57czV/MZqG0
tfil13WbhHEi1WnxKYsUshilzycqUjW6dACac4vSuWXD9v1JELyG9jwy3H9iqOlP
Gfjz0Q++IREI6jXP6rmC17KQlhiOazKcVjUe0/bpGEjyePO4cdH9wkwZCQymWv7b
G3d3X1QeAoFOhLZoPwF3XTmOd2IcdYdYoIM3eyJlfxJQYLD1nDm+HLfEE0orQldI
4aXcz/6s+px6weetk5QYRnxltsNbQs11riIsne2pU9YNCqn0CdHWNL2JemQnyKhz
A7A2RNXYeV1EhmICmNql7rAKlfxK6QeucbJtONL8VnxZWu2AjSBpgKrWLd6VT4L6
X/wEH47DC8gZye48crW4ZaRIm6KXkILNUVgj6QxvI6I/Py36um7tCFm98RbKtz9z
z5/53jLHDFFeSdMNsBuVAXP95+qAv2zfo+b5OypcMvrDTdw9tE95ySWlhLlXKXNb
yGTNRUU2JpxQTr/M12VDNDnHeJl7ykKP9FgDLW0HtktWr+t87yKkUD+uz8Ga5zFf
jW+VwGDd66XI/g6rXrMQHj4KCrTFZL/LS/VVvansEO0VcSHe3xYuMcLpTO5X82gv
cbf4/6/kXt5f4R9AcgrRbZSkfhpzF3ZI552Rhmj5puSxSH1XoEFo8OjbgxBzk1HG
yvECObPWvN/INGTMTZ+M8fjKcgKfEJBA5s9WllDEqsRyFZ0ZkhokoY/hsyM/dhtp
0dasUeXkgDJec/VIckiaGjDeh5/ohvHuU1sGW5SFhSW1SyXIefpY6ALJNbZaoxcc
gsBkiYqu4xG+Rtbe4BS8lCPEsQ8+v8ij30UnIIrEG7wItxA7M+2viWvLsPA1OepU
jyt98z51IcKvH9SqQ6o9Ajhv57krCg4ICs8cJoaXtG3lqf0zuJcLYP2OOAS1AoU+
OUdQDVZPhygu3cafntTb4P2YZQTD0Kcj771AVN1gfS62Oy4Y4FXUItsina+8QYf+
kRLJL53fSLhGlvV+AoJBA072J7mhjHjXV1P+NX6BGIunjgnlQB2l2oGtl6eBcsKS
T+Dm1PoLKPLfbeUWX/IaQ9HagBoa1Fi0DP+TVjF+40jycS36/uEJJ8T25wopXN1r
j4nWTnO07QZuPyk5ioa+F8Ek8DVrLzjjAXKuVFpiLzJrwg0M40acCKbQpr2XtXND
WDJWGV7gNqH/s1jKUJOh5NtVGjyumbDguKWR/dvPMCUELCqz6s9BV9Q7/A7A7bjI
hiVvkxgUV2osTWQJanqhVmpb0gnJAVBInNyu++tFdZv+e/0PO/3BPSyA0CyNEX4X
qQygEi+TSMwYwKBp7VLzh5t1n4hOS5vut3RDefhaeNaPsakIEbcZ3+qRQvk6jcha
iFRlZzE/2s1c/cSGZqzhFfV5PTPXY4vfLyrID6iXYCULLp4BqtVunX3d2VIWW/0g
wyjiYRTDD2IgKOI1oufAQxQpLw/rQ1zkT/9F60vDpp1e6zHLSmJOGQ8UGiAJtd7L
xesK4f7O/10BGi8+PX8w/qW3qHV6l9TxkSgBqF4AgwNE6j4IP1feTImSGGF/J66O
yU1v6mgOYiRQmRWvahrkApTLTJh31IM2hBmdU0K6q/HuZeJEXWluLR5sylCsQcwK
ZkFr+LVwzrcq6P+cwQ6sY+k3Cq6bkIl1aOJDp0vhs/cFFGQoYYxy/1y8egqGuWq6
JFFmATTPg/RBpuCj8Jaan9UDJLXekYueqQm+k5OXvvkaJXazqiWJ8/UquSUYs7gp
cTqqQNFbWABPGVjcfcDoP3QhaXF1KduLsdfrTQ5Z/j0OKv/8nbts39YDql+qwQI7
irIEDLR7ivJr9DR+3uzWo8Uetd70MkCbZIyE7a9h7IJkSU/ei+YUTPkKcnkTZ+Ji
dQM9QfAOagHpG4WkWuuAh5R3stFf10l0XG9hSktXMHK2ZSpV8gyYu7DZegZ05bnY
e9Qy0jLpNxjuKiKXRNJUGS5WTOXPsp8DAxQbcwraqVXa4rZkaBPE2cYY59HzcdiV
3XgUlgFD2WGaEwq6PH97HFuzr/sVZC3UQCViAE3RUHEkQ8FiYMLmKW8GmWC/sSJj
jGFfqtNBGnhJY8Tg2KsVDKB4NMIGAeTpDiTcaZD+/w9ATBcE+x4lMcqiGq8RfGmY
iukqCxJAt3kfcdF7fIR7toKVrDtXvTuUgJue103nbjxKN6JYIbuSNjafTyWMAURn
rVi820pD4WITCpj/OcKreMrXFq3KryBa77kDC8Cz8AVLaLLXricI/mPCzM62vngO
ugycWxM7NrLei7uBgRWtWmK3iCYGwk3+aV4l26cNQj/VQNAYp07YGmFe15ldkfpH
eRBV9Vs+7IpzUUXdqDNwJTbAPUN0wM+X3Qvr/X5DxQ0VcX5DixKXo3RA59fbMrIZ
ExWd9DIA6paF3OlD1RYEpthpw4LCctuGyl/CXD6OZfmsYGRalcemkNYwATgxSuiR
QAOB1ZpHq6/G+IiVoiymcyCyyLK1rCQ2gaI7NFOhtr2/NY3PvDV8iWEy4ER+indd
nG7WdQh+eYXhryghegsuLlKoteYmTH7dVpbgUtR1tCU7fzVf1F3IeJIjTjYTvNNt
Io1vorm+3cKyGH6Ajl35YV7JxqV5xQwkZdX+3Yx3kQ9/m/s7UXhPBZOVigQYrqvu
+t3zgiErtQOjK+4BBslUTCRcj1ix140geZPTaTCPDVfhbFj+2kWIq035v0k4qb5x
irnsG0YyynJALQ9oQF/MRZPYVLJdKs/TmpVQaIFNN9hKr11V5wWwg0ZVSiAiD4hJ
1mvh/5eUpH1lEjhne4ZZY90vPOnnR5jg+8hlRlGyxXtLkrggwmbDYIX3fdFtOI5a
/+Go4yruaDR2v7yMIxXuCeILEosrqzu8YtdHgd+EjLOCRx44rPyXxdNk4EwcStrS
o6a9hNi0fPZCxDxPe3sa5EP6oWope3GAqOn09T+q+voz1ANXs2w9i17qwagkb/6L
pATJyUjBHQB+vBrsA/CmnpZH8KCio+gDslFmOmU1mi4wVgLRUvq4OSg93G1UXL9k
WCf6GM1pv2j7nvxtIxX4EiyI/scz1gLfR3aKeIU9nkoyZyyWY+MExs7X4KZmTkNe
m+RcxQRL61dHSu1/87YQVUvcH/VVXodSCzF0rXprcuWVFl8l9PMav9YpJi7kDVMn
vn2aBVtBnyzD8OuG7yNda6ZEcL5LEvLsA07chD7nrhBQRAZr36A1trPBbi5DCkvU
vg0DPZ63iqQSbgNcd79skGCx9N6jaVlkjaD5zw8T+txYAn+0x9jhH4YkAWMt2rL6
rv1iVGFy0hfgOPzsNT7u/Sg7voSQ7JjJAJYeAfKMZw6IsFLB02sY5MdGofqoAazi
SIkQnBpRSQKxFKu/KK9rc6czKCgg4eI6rIQ1YrILNMmTqHcCBsuuMSMMGzNZBwbt
K+wwXLnRvVwJaN11Ph3n0PaSAOARYGC45WgbwKglEX1M1CdSfbjV15JCCI3qgTM8
LMg04UG1UFd7Bk5C4/q+NT/xhfGYmGYxKBAGkoW+lWU1QHIA9KP/w3Qqxk+UvlEu
hEzmIs2Q5ubYh7bfzKHt623abl3Q1iYgmTkcaURhYRk6TvwL/5QYx5D7PKkd4XR5
28ezz/9t8zZQS0mAFRjh8N2zX1K7eSSOextBVILQRUJR29iG8Vivz4ZNTKmi4CDE
rj1g8aNJkDUae3dydJzkjG4mk2hpk8YgWinZBKT4MoAaNZpblaZq/4wxs7vL5+YL
MVo+yrIIT1X1s9jHPBCYfpo/J7JZMHOPlvd7dP07DOY+qHqxhw7SW6jy1oK3R6r9
qRGYJDMHbj5DxgECXhtcexnD7SfEzSOuUeZzMVB8TlLEdQA88uChCnPq8Dys07Nh
2/JWVZcmfpL3NNEacjDmLXdUeUNL/zmt3A5Na4faDvD6Aj4jDp0xwOWzzl4unsSg
ZzcC6e3YX1+ufhaPfEk0aJ7PsH2XXV2+xLvqXa6/p2eMiOYRxYik3RTLjyHTgmZF
0jJ6/V9XsY3k04TzNku/4Tp/+dRI6m3zlq/zwd7o4889pkBxmFWOC7uwJ1lGx4pz
ZMllhMNU/P0ZHlxfVPwSrMMlUfPkhKZEwxJr+pxIyWrrO+s/cqpdeNlEB4vG/VjI
x4oEqBXDSYopKhGDYwtx7sqGS9EzL4FTZVKnm0xnhSjwC4/LdeNuu7aplbVF69xT
jIazeNvtUP9pMtQUwafqgOEU2QJs6TxWSR8igzmLkezL8X4RfZcPu2AYoY4c+/yp
4SItPsH6Q5cyq97kKqjZh9lFojIi5mvXMZPJySmeCApKhMB3fa6XKTu2YBDdsa+U
/cbDwdR7Ne+yE7mG6jgco9lk1suINSv3jP+1e/N6sd4VCtX5bzffZDJJxN2yoeDo
GkdT9kU30STeEQDMcRTSHXfQdHDYWAAFlj+bQC6ytN22Bx84fVlg9TNhc0Zwfv2Y
PGouSKhQ9G3YL6socZMgM1Gs2IB3dQJM7c2TJjBKqJ35E5TnGBR/uTs97Fgokq7Q
YtVNnzr886bhtlzxcsML8MWWG4L3ILppW4f6loADzHyz3dzLPuG+yAycordMVx9e
lpSHAUbhoiiKIMrcpttLMenJrhYc1jwQy0T8LnjN/0T/H/qj398CW5uMwTjdbWnl
i8JymB+AzaxtT0Akj09ewZVOKwwVB+SwzWetQBcsny9D7IRufBnOq1nVOsVdyCeH
OpJocK2uYeXQsl4mS7TyJTG6uG2ivtgEKY87f+s/XhjjGxZPtXZ60Jk9HeY9pZ+Q
8hfccmvHgZ/VxKfTl14NgYxYEuk4Vyqt41LlMXgDRv+GLlIcyB1+Bw52j5DCdyIB
+cKLVPXVBCZgmqFFD3t2KOrF6eU+UjnoRsSx/R8jtuU9U21UxDUy8tmNwPBuA4VC
3FX2vjuRRCSQN7uDLoCgPAev/FBhhkoNopp8+k6jPm+RGNJ7y/y5VfYUy7BPNB+u
6a6ZlUzcHIZbFVF3G/UtbRa6UE3aZJI9/wI/PjMab4Q5YSwu9ac+/54uZXp1CaZs
LM+AKxmkM9SDTpiEWa25w2Ga6ovojkdxrA5Bk3epb6sYXzB0Zl5i8pYnQU0LjIn6
OaqCjZ8m4pkH2lPtHbzuCLSwQwM1iSN52GHv6AIex/3am1ErF9j4EUV/Ooph+uSI
pcXF71JfAE6iRjX5RDDFKjHNGOqaCroi660Hjj4PLokFxd4HvUh5Sj4/jaW/Z9J1
b4RuYeETxivQDh+LMKLOH7nsfrQh1v+iFelnnqxkib7qcqddyAFw5j4dJnQDxFcC
xYzrhF6Ds6DWAvRX2wp9NdwAJ6hSO4QcRtznW+7F29xD9t20m1LBWan3sc1A1m65
qiPW5fb1xrQ8zL012rNad9pYT9Th3vRGB4vRaQ1FF2MZUWKgXaGPfAvONPlmd0/G
2CXc6rvhKshmMPeN6sZ63QvDlc33UpZilE04M+LDwO06nCTXc7S6ljF798j4N/VZ
p46vW7I2LbJLIaY9Uojgfr/bksbXy0Q7EONvHt0jkT9G0+2Ng152h/TrbR+EaFnY
HlXp3y0ueuKUkcmvOTm8xSDuvkaruMnHvUkAtWmEcxZlVvIw6BH7sAmeUeSYk15/
icGKUWNQMbOOKQ3X7SlNF4eB1IBVMUYKkl4rEOy8UMexJ2j6PeWjOUDr9cp7W72M
L2eoY+WoBMlX6SQLkEPwBs8GsjyZBLJYqrYyp6AUgYS2/7OLGO/Lz4dJq/vprS5U
p7Q4WcGsiSlyQyihYmRcJMuCL7HDxNuJIxdzm0drQfVEmNUUxjSKCsm6IGvvvus2
1VpsljlVxqd91Z1UJEIJIK7KRwxTr2p+I6pnlBNYHDh6h/yRgWLzy1deglSeucFL
lL+rbaUFaRAp1eey3gZeMNCKXgEM0gudtPqrgc22PxxhXTlWWtJ99QpQsPhCnbWJ
rQXcC5SOPF0yfoUbS6HnV1FIbHOXf1Fpvevwr6MuITE0uMI8zuXstSJuticFVKF6
GEzz50MEzleirNwHnogSRS9fai28JmfzWVqZToRaH3z636pyDZL/4rCzHKiZsll4
45M/zHCemMMCMQi55VfiJ5nimmb7qWXgEzT/8FyaP1jVA4H61L0mzqZxmxBj4ePy
XiIejWGBE8B4+sJFIDCRCVZuoPVkJLKaYLr0sMvrrpHk52cG9H0J+un9//awHF3c
owqr+4fDFYd1txq0uZO9CHxGuRganmkdvPNXlKbk4rOz1wqAxySNdx311+vT/GZS
l/P8iNgfvWLE+4oiTHv4UpPwfix+6Bm54SGcNAh1oLCZFiEuaEmZa9N7sQylzmqm
mnEa0wm1aFz54P0DmnjHZV/wnuM/+ziV+dW408JvC/M7NksXqwLRRHCzdDPT3YDj
xeYp9Hyklm1euJl0C4goqLti3oQMbCw93lSyumAHoigw/d2Z+qKzIoh9+4Zgmy0k
Ze9iF0D4rx5SUfHYE52MUGZVtScUB1YdQQyuqoVhuYpmGoIvkkeb8x1M/8Pdpf4z
6mU3OH0GvWHYkujBiFz3CwKHUnZnXg64qAkKZxdpn+p/S0v+qdDyhC3C3luybdEc
pi+kMYgpeWy8Z1sfxMzvqNYV5M5776uQuaeeWz6+4VsI1d8WjAOXciJugdQfC90W
s2PxhxmcIq9o+06PLQWoIUqaf7x3G+IJvFwpdUM539cUNAAXoPsS9B/qYuscMZDF
XHHg75+azuYHEawRjPoJDUuBJ0ewNIEP9CzkW6J5VkhHWkmiDXYgDylT19jAWMJZ
YzfI6hcIGFRvDnboPAJLn5n6ylnikqTnxT5PDXESwRm+edXteD5v9blN8Q2XOJEE
+S55y7AKyB62DB3v1rJ0am4DlMAmwYRGKT1wQsN4vTt6xjeCt0U1a7xFwgaW4IDY
aWMoZXapaWEq0C2Niu8I7NW3MJ4RK5ol6T8a4+EK2JJMO/Zfacbm3ipLjBLo3aAP
eV9D+8U26kDyTQn7cj6pSsCo9EtemmlRy5CL0Zr6lCZ2uYfCBpDekedOwIgMMbwA
eAwliQvyhqx89tmOiNexWkUsj+f+axOa4JpHYc+lDn26sdjjekK9G5Lq76flZTaY
rRqC5ISJwNKTXvy92+rD86iF+QCZgRLcgabjonQh3egKV4GHLghIYb2MHm5BBkUq
cE0pgVvJaBqfwfS96nllEZIIFGHQE90p3a6v4VD9CWsA1w3z4WUy7IWakgsZmt1P
qmYEQD48tCm1owx6PMBrSoa2XTZbN34l8ZunSBVKLnNub3FVLGZ4LBqljFdC2i8m
msyLIAyPDnTAvWEMV3K4vQoPulbAW258awtIfnXZ6vrWMV32sMay95Hcsk5XvMsy
CYKjSjiE5xps61lH246zpsJPo5yFZcP8bpz0lVHbTS00kCYoIb62IJI8PWUlQKrJ
ln0sDo6Sd9GkUCyxk1XNtCLXk5gKiARRTRgbXl+FIn+A9ufDR7wB4DCzqmgAFBHx
C5MVZ2OGzyJmdbT5NjsV8iYeKQpUQLEkomSSBmK5t6UJn0k+/GjfSgJj9HewVas9
KCg/bx5OW5f31UkmYZKZxD7FE+sWw6WmufHbPlANqr79uFu2kqOSmqkR+ud5/u6P
hdzXi7bOPsNpNKfg9EoIolfOPDozgholXatWm/60+i9VjjScz4Wa4Zqf48TTFX8L
Ri0K+KCM1tJK+QPYDZS7ZxQ5BlBHo0quPuwVcxCtwXMT9j7IiFOszyHNoXLboFLS
SGhESZPLKI4HJeg7zPmPZTAzxtATsZgnPs0+UtPJQpRzVUHDk0IrLzNja0zLoiOs
Zy+XtVNnLuRwgGpOaKeZECHui70l05dqr8QG2HainY42b7RVYBtnNMAauZ0XSXlV
13wnPMY2bi/6+K2FnvvQ8cyo5RW9UDINnuW/UR0Ppas865PswXm//+PLY7yO9VJA
BJ3qYOB0esJk/pTVza6dAiMWJnqovnevix4raxmQG4wYnXWtgOzTDVxzznV3tYJw
mjw4TEGt51yBxUvKLAZsqudAf5m4zxVDftmrXGPy5Xo7GeMMlEZfGW4aQVSgqeep
S/p+TJJRMOdniD1JMjWiJcz6WAKGlTvsakR6sVTWeQedeEle5Ie5Ed23+a5+vdah
nUlFtdi+r8Mvwo4nC7QaWyJ3ahRJ/N5dQCrYt8ChXz6TaLrdABQKV6eei3SHgsPY
ptZOPmLj0DWvdhhevPaTb5z56pwdUABTiGvLmI/u8PyGhKktC0Mve2zbyiJYg5Cc
uPmwkAZu6OJLuuUHDkv6An2OrZr+74OY0ZPxKxzAOb1FvtXRvLCIdupzyi/Xs8nF
6yjagG9H+bEoC5w4oqJsaXCph84Tc0WuNJVDFiWINiiQ6tLn7zdcKp60cvt3xl72
JqCW0mB/hSOEgsvzuqiRnjqQvem6kVlM20EjwL4n5grOXEa7L57PyYFq1ektGSB9
C/Zspoc4pPo8Giqbfo//Sb/4EhFZmu28pvMZG4ivhUdn5fvbjL42mlbgfP8B0tij
i1B72mmEVMWdIDcNUM3WmcSYhmHLlm1BNBKT/k1nBCNpoMrBgXSYj82kx4oGXdhu
FjGpPcAfqKClbwbZ1/SsF/zF3/qWUwP7IdMdD3BPUPw4Q0hwQkkXtERaSIZz2ENU
5VGRb9EyB/1+KIxf69eUnifnLyxXOPuRMS/6BfO04sPiFE0eFJyVlEaibNUU9xld
7DVyxbrfFCAcziJC4Z6CHIOyqfb60KEYL0B4WMVijVcSaTQ1OSKXkh7wag80TA0f
KnJIZIXHNUaGH9GQnQXO0SSBQizHwCrG/D5gDcEYWIfvqG2lAzMKgTZeHLTNoi7H
QX2Yq1dTCjmpKzV3n4ShTWWxj/35ixUUP6kP5dzOE3LcBmt15VDoVuG0JsFwmVpP
HigaxbGp1ZQ941QIViFfcIEbnNZ8/IShyhkPR2i9KwGfSVu/cEv/XZhoB9Lg9Bcr
uHxGL3JzgTXuLrBpA1KAeBpKxi107bi6WajLYNOYDXleVmRdAFZCw6bDhXALkNGx
XppyhKttmdjpzrdlzVN0yImcHR3uiBsy2rNfrjgCS7wC5Mkel3yPM1abG3ld9o6i
nPTDQ2kiBN/YPjQdaEj21FWte6c8T1cxroFRuYSHfxfbBqVAu8zIfUKOEbVpH89I
xShI2cxevGt6AnkDVT5WiW3wzO8g1zpAwfMaXlr2WcZu1J9ogGW9j7A6oDtf802a
wgyoFJjBv+/rKzCdRV7/Awliwa1GM6wKhyr8tgNoflp9HRtKCLhqp/rmPK1un68H
EFbATlm2J+8vmrlOcBsX8P35lqXIt+QiOVoTbkPFo10DeuEKyel3AFGmXe+ryyXK
F41Nc0zrkfj//pS8LeNt/vJHHHLTfkKSCovsjGJAqcS3valJezWo0iiOB3v1tMSm
oXWQrKhCJoI8Itp7XAtDk9PeqTZhss45aSf8YdlC7KIIHvYv84LmVOwmqSS5+FBy
xv5Oh/EyTjTb6KUzH5x10Q13o7WPozUtevTqu6XhOHJ2rNv/yp5kb+Qr7ckt1bMl
GvUYeGDRkxmRtevoKWfCjYdVi1leVcsla/MUntC7NVydHEoO83OrmFEXHDLnpKR0
7H8YNFinjLhfNdyY+s3O+3oHGRWJ8aq9IAlbR1HAdD1+qpEwxBIUVbXv6fCnsT0I
4clqJKzhEomCj546eAZ4ptQP1wW2s59ygPpws79+Ok+gbBvUQJbq3rbK8YKrGdz7
/oGEv3DPAyL/i+mGQwUqIb8uqnQ2PS0blfKxu1LlL1HoYH6V94KQ7iBYZvHVeYtv
8NmWWXXuP0xLD0aCvTLk0s7G8eh5TmSOszEQ2Es62yN+N+HHVPiCazEZwBXyeK0n
5XKHRCmpuVNc03wscIwnKOR7IJw9uHK//WhzpmdV3PJtXYimi5Wit/GTqQa+cvKU
iNIt7+bT0aCHNoDE+XiFEfUVf3FRe1Tj289a3+oykHfgEloWVo2zQOCxMBM5cfRb
B2tsl0nS3pgWPtUUex7/C8GbDS25GZSGXr5B/IZRDFTR/yfEiBs95nVxbXbmxFg8
N6sTsukwB9i5cBCYgOboVtGRQ8QSMY5iMcur67k75sI998zaHvp6ps6Fsj8PDCj9
ALhVDeOM5WnPYvR2JlQ2nC5TLCDx42raJe13PBd7cg7+fJm+LLs5EOL/iv1amWT1
g95A09XRbGWyNuWXV2Ilp0uVy7uI5xpxnUw+Yr1ZiKqjFc+IAnjOnnKG4GgcgsiF
onMg00LaxHPR7a2MmUYeI8b59V2yZ/QfNmREJvryeRiia7FahbsnuboRzta06Vm4
k9crZDxoR8e68gVjcLPb10bde1e/N9kH4P+z3zW8E1tPaqGbniMDKXs/uCkR09/Q
F7FUAzePs+iEeGfLnH97eVvVZUtiiL3C92ajhthU1IkLlykPqk0X6qDgCf+z1NVE
aWE8Vuur9yVpui+LQ8fm/eTzNVNkpot96cUiHsTsKm7f6gGTKPOhJPQe1jwj436p
DiQNmA9XTUn+cFtp7M5IQxXdsfvLmCZS+9HD/z6SAfEW6PInvoTWlOE0QVgREhEP
SOFSBquobxYc/5xS7kIXiGsoFCL5eS//LDss5tuoNbG7eNH0ac5KfneABPUOfjFA
JjukKqFLsVPS150E12Ku/oVJI6yEFl8aJ7eU+qS+yLyM/Kt+3nsBagas7QDjrAmY
UQyzxzDPD5UamsnlGdLL/NEIFh6/FDbr12LtaeNenPCHRbyLQk3dOW5CQCGYZ3Q0
MCXCRucdtOFjomsSgGrLYnkjXQiBRSH7MCO7e8cVD6CrSn31Q75XQ+bvv0hRh5pc
8+pUlujV4r8340arHeYNUfox1N3t23s9Ximi4I2L6l85P37HCxJ0gJ85i12Q6nc8
wsHEIQ8hYb5HRI8GjnHQiwZlS1GP3e24Vq1dQSc7/h66Vjz4ecJJvPZhoJnkMoxi
lp4mLTjAdSwwletvj2dqxE7m9P7S0g47vPb1hFTZholXn9ZE8SVEjKZwbZUcGxpS
RcRk661fTRmP6+JLLTDnWFDnQDxrQEYmuBmRg1KulEAy9Ful95brDn+qmQOYcP4s
FpEv2KWcH70p2GkrEA1ZtCH9Pezg5gw9oVMZXP34khYcOvsOJ/jXyaanOl62Igpr
wGyNH79tm/mxn6/Xe+L1nJKaMPMvv9agRJvl4qbb92cgHiY/DDxgCM/VTmmiV5h9
tJVbJ+/c18N+NK6dRtSVzBm7pzBRv4R2lm2gGx9G41YE8QRCNtPbiID6y6vKjjxn
13LdI0bfpfgr9Fos+SBwMRCmLJ/7WyWkeJGKKk95JIm8G6gNN3erYkcF66Khviz0
8FIz8mmpUNVPAn478ZbYeQzrlNJDp3x7RFQ25u8QWNwg6/+lxFaWFIWTpAX+n/7K
p7/6YniItk01oNv9BRyAvnjkmzklPjwc3FOkVehAHj2737UUzOYONV3iaeVWHeWl
yJTpQfSD33gBnD5ZHBl3l36F9op+ixTRafpndKlnv+QihgtfrFrsoVFHSnFqa8bQ
x98YZhPUeYGKPT9Ce9rALbkrYST5Qw0Da1ysDh3JBCXMcp4rwbIrSwBbkrd5RcET
oPbo1sIBQj+YH+Z+LFMVxAcWfoy8mBs1gMjHCIV0y7PUSHxKu3Xi6Y/lFfZo05v6
XXXVSSia/KhWWbYR51YgxP86zhOgtPrEsnZooNk/VvXeg29gwqMmh8xaQvK3WiIf
pRn2gjaHNNWHXRf7kvFfYV9AS7zkBuQloZmujsOiJOn5Hvz9vj+YVsIVTDaw0zLE
91FHLo2GASz7Xf7wFFNQ5Sa0pTNO34FNBeHuWLXuVL1N/ol8OLcxFNOGBWlSwgBw
Ozj19KS9kqd3JSKhUBBXyWu65IglE8RBjnZMDv8VpJqMs7LwXR3Vwcxtiq8Qdahm
zGLhYZN5MmW8Y6aTXNQLJBz+/zGIsDdNQ8pMtmdwd2QaMn9RzO4LmmzoZrZjGMkw
at3mX1jWgmWRsEMFxUYyEuHer7FMPwsriQPCZINmOzcxeOomeUiv7YzUHOPfkL7p
8V+WuGrBMdKSANoWv/yhMs19firFSdsCrFEQkJNQHRXUFhR9GBg+DBCcsLzgIm5F
sm/7EOKLokm/DCt/O2IwstGRd57A1DlTOLqdZUktI3HXmDHdeE+x2G3BEK+MNlB2
0qMx7BdkIS4UUOJV7cf9aOudiZOFkMIPw7C2gZrtSGnu/9mbSlMkSsud00P5k8uR
hPEv+8IBKPvgs5gHEC+ega1vjS6MG3KJvvubOsKB4/Fa0s7xbtYFNro2NCqLNrsQ
29tPJgO05i0S0K3JXSxTXgzMrqIGWwtA8opyWRVi7Cvn+uGgu6mvu6gFMlElZ8HH
ciypc5MEUYY1yE4dJ6oj+o2JVrEchtt+j1v9d2m8Lj5zXG4K9yp4ZRXzLxxVGx9a
3WTKnaYMCTL1KaRRTSSjD1GDvGF8STbKAf08hc1yRQRVjeJqWg8bfG1XZ2mgoNSj
FyY3oTJxQF4S1ZRmmXXjuC9kaHfDliVK0acdPOfgoMtWkBiUwvyAwnUrq1+AHvOH
YlWpMHYUOVANtUovK1x6NeBVgPD3W4FCPRBPyByFTIkfCYs+hTY20oCJU0be7mQZ
vRDmmXKQaxA3sazCXZ7XsYzOyQwqyuPDE1V1C7Db90f2rHkIlGa0oaU5S7uoyxAz
8j1bsKQd8Z0cMLi5QQFaRsgrtPGjXQQfk0TnMZWVWo8RrNGW3SMFu8ZqlXUM4gsU
UPm56AOiZMSAksIR8e6pE4UAvD4X/z04OdJXvZgPumqCHSgbaTjG5OiZeX4hC4N1
+SAUlJlIqBsT5wNYpIZjoTkR4wBfxheIu95zd7M299cL1LhcpYto7XJiA9PMvEb8
BuSw3CDsjIRcj6TK8L5CyanSjQr1slhHbWiiKPx3a8a7cz9NQGWutYniZfGd9enx
MlPCmNbkpXmTgPGSm+sd9f2o3R5AKKvKGdkbIN+9It4XLT5SsN+jtVLrb3PoCB6U
dd4xOxbomfGaPVCIsrr4/ZYZzTyfYd9K/E3cN8QVNhEFFn5mEDNCzf52hv5ePTfH
YN0kXslRoRvBp0hxlMhqaiJu6xim+H+fQip4wSf6DPLT285NYpR/ZL24a4OUgStX
2WkHEbNrhWi/Zs+vPBaqu8Rd97i0ZoWFNfDFGDGKyZK8CNs9uwzV52T/ZnvYw7UH
XZ9vgEfkz9ll+F4wjFPKxH6Dt+nI9KyLwGnt1aIXgk7gxBEBxrd7AZ79kOzudLTR
Ce7qe9lmEcnLBte6iVL9ndfUKq7VHAMznkoU4XZs6IiJ2/2je0nk991Q4SQRqS8c
ZtcRzEhAhv8f2Ob4YgGFu7kWC9nVwaipjLHV6xcZE2EOdcHz1yIygpoaroZYidQ9
JE6Vg/wu98B1dyeJ1cCoTCTgXnzhByEqx3WSn5X3fRQJ84bRYIv8LmBa3LFybglf
K+xR2+PZfjQBCxpHr1zUMbwOdTKQhONC73GCusVtN0gd0R3zCwWI9hf0ewOAHUAw
kDP1vbkbyIz/lGOa5F94L4YP72vo4LQ1UxcgFbJ+fIV7j3ARZAuxPwyHK1IF8cI+
VJxOMjjCEFsheZAX3W8j+fn35o4So2h3McpI6ZrSSG3Ak2OQWfWk+N9c0frDi1Rc
buFuH9kWN8UmFYxjlr+/xWMt1ZYaxjWoUNX4a/H0BGk4FdUPIkYhY7zXKBFp1PK2
9VuvdnwQIFRBO+XVUY1EEcRow3CSFEzSPpMF8lZ7b8o3mOqUcbeNkDOsY/jFeLaD
io/ydV/4jXcsgHwYqBaVyXc5HBvJnw0UL/05fLpAbWyV7qXR8FhgR2a3Ui/VzxEY
2VaTd8MyI5Q7Rsfim33+oHo0+rjlTCm6sGWiC6fsliTwsnU7PyXoHKkBpeqkvOWL
8N7yGFg68+dPHV1wPFFVrpgwDg1WCuAt3cwObE4+5FFiDZKX1okdhZIZrizqc5l2
VRcrJGwFdmqLbcHXqBqeKm+uRTfZToInxbwg3rkttQ+LYsq0/8lBzUJi0DxH18U2
QIr4nf4CF9WLs+Ccnt+cbJKvvU36LurqiW62tYCwLNLrSFIR96GshsOew+k7H8+t
4nRAiDwEGL2rzMZf7/udTZt5D7muKYrPQFsnRKoBjQcLAXn6rbsIqo1Z1oUgDxjF
XnAaReihkjl2G+z9yZTBcy5eQj46GsDr3Lpxz/7E41w8fSlwg1ateM8+nVzyyHdI
Jo94V6ZWM1DSFah+IAm+BGKqQKPEXRwmD2WisIDbhYW6xiG7jS8/DUSLBGdHgsM0
ddT3Q9X7LAoXXi93UYaKD5SwMoUgLstXkOdEnONWVdUIE9tBCFPQHZG2BGv1tcbl
8zym2oXWj/RXrFXNLsQ73msTfcU9ZqWeAG9u6ewOv0OsRHvG745um4Qf+jbUUhgc
JzDFgkEBWkCg2TZZa6DyS6CdDbxu7a7t4vB0R/NZF2Wvry2Y+BQiXPOoZAOkAH35
zRq8qjs+h0Ep7lqNq0szrCChLhRYPjLDgfpnBxFs/hZUo378iAeApFXGd0BiZDVV
7anaP2tsCfdN0izBqu9Bh2zYJhi7uHA/UVrVEi3YA04hB6q1U/PdTPB0LA1POi5R
BFwUUgaleIIMx1CX8wmMpM5Xgx2G1MW3KCGt1647ZhCj/YDTFwyVjapt4fos/MbJ
04pilOelBaFXUul3iT7SgdZr1vU1gcuTzlDfml/tzQi5G3Hu7wTRUOFBkvAdltp3
0naFfizc4O0ZXrrUz/GH7XKXkZ4/OXcbI2gQfSS5dO0rl9PslBcTqjulBGZPdf/B
CLvbA7LLz5Kuc1+C+WBtAzNOiKYaJSPApsMwfPbdl60RpfSNtSFQztkdDVSCepBE
V5rFM8102qp5CWNwz7qevoEFaM9MS3mimD3EGE0NvpWFwWBE/M7Tvjz/54A/iCFw
Fau8l04TZ1PFXlZ0DDXnoKiA7WmUbV8ohuoz97FS0Rb68WkJiREPCR6ZiR4fFXyv
h8SwffoBNnp2jS20OOwedNDkM637/8moVVbgV0EfU+fhzfC2EJormRfC1QLKs9py
OVULDXP6ZO6YL9mjw0uV4M8vxYBPFue62TmR37w2o/fyvta11g35Ox9K55zAHPDm
EpK8Is4MI1PS+93M4JtPBlMyEJnKLnOuIiFKZISL4X5kv3Di6UaU7Q2SZgXPm1bL
IYs7dD3l1BRMPwGepzkTDRVJCuG9u+LEOBLnPISJoavcaJ9Ix8f+BC1dIIpxI4h7
JQN1VpaUgNJ5TUHxEeK5p+ivk6ni6rmATOT84yBPWVgY0HNIRhUGX5d02Ggu+rBZ
6d59Vb+mkboEpsu9NTylka02DHRwfXYGY+P1qSwLxtj8+zo5PRjW7/j9X6gYQTqs
ZRIG3shnDebU/L/W2xxvftXaRGMdMsi9RgJbV/JJxXW6tfZ6RgmHtF3AsXFW5Rig
772h0QL7njW7p+H2o4S00zwn/wBI0TSc9SF2kfjfpWXWs21Q5yw6oVY/hy0E5Yu8
ymT7w/IkAkQFClZ/1+tbAtxkwgv/PDWIOM6vbfmajfKh2cDRdQ0kkjSatrqnfG/s
tgdcMiQC/9OU+Ypy+Z1XWVC/uZhOd2z0hQJS2jAk+fqpn9odyYcp3+Lg0IIG3DD6
c/MYPn2YLkFHMIdLHKeMcE+xBTSvLvrK2ULclh5Rnn69n6QykuikfrqXPDD0HYV4
Omwc7fQwWzbiHaqcugGdFwcYZPXtldMi6AAwkff7LerERrgEIIUjlDHtvB8JumRI
2hIQnphlSRtGSRSVWZrFHbZ29wabGXw9+mtAsoIO49gbDqE2RiH9VmQTGSxvv7rf
ht0zmWf4kbL00fNm+DZsj3cip0HRG93XBOKBL/ke8CRU6OkzpbUyd6Gfnm5A3+QM
yLPMFUjN/9Ui3z5uVvPN/BnPRoWNKx6mj6FfBf1WzLmpJjMIvwyw4oNII+uNLUIg
QXH/L6gw/IofNStP8zjIMyzIkEk58gTc0C0qIU9piasxUiL0JresRmRmP5uu7SJW
wxPIcxyAHjfiYymPr/1tCXCQLTsKFhUY3WxvABe5m3vHaQ2V/JyUPdXqv87CU/Hr
/V/cGAQ7f5ePtJBG25o6JwcR5+590WpjdWRjEMpWjaeWsc7i1OEo7VjOUubld7k4
LEulk5GlfAR8+PwD+E23foCJT739UI8ZdBoczcg5py8uWJYBK79aAUUJ48x6/CIn
RKYpxnlRS/3w8uI2zSL11bKI71qGzvRhySmbgQG4C4LKTmYZx2jJAS7Z8qI0QbK5
IVCdMtcOOauwNT+Ksj256o143MNOvJn33R/EjTF6ElnFD7CIzjSmxUcBlqB+H5Jp
KnTiZC0cwr48RGMcGC11QF86/BAcJtzkaQI4nwAZAq2dzEQAsJSFFHu1NEiQcMrj
acq0ANk20zx+ivfnmSiiGNygfC6qzmBJRyxvVmTghfQ4RS65PrmrSy0mE4ETUIlX
sabxPhnhVnmg1bgHOE7OR7jFeTDEJ1EcoqMB807qf4xfMCJB3iC/LGTwb+CIyWLE
WELr1IZKtiebDOlO+0o0QQj49rkWou2cJaEexM3c2v95XHqRnTZY480fg4DX7Zdj
EmPXC4L29DWPxpsIuLN70e/aYTcQ2eih3ZCgmPfx9kl0WveaFteJqy69W0lBJUyT
CQeRohHVtopOeV5MMELxBHcARxh7r7LDpwQ6B0JokiTr+zPdHk0h/vM8YzHK69oe
BMYZyedMNdFC3THYAd6+etzXehLI++aYbd5u2s6sAaLoI3stOm4qWfle1L2gAG00
ddTqnlVR5yWmXJGlB7uqCK1p8D22c9+jIOLXXfh81NBP9eYwxIZ6bDcE9SbOzPV1
WC/rFEU1BXC+kdHHzdCEPQnyFvw06Ki2wtvsih50XXnX5HPaJLesdP7SaWY7lpoi
o1+uWCkwOL9NS3lVTLABgkw9UUd6qIQoiCt/ySML1/skRqRNk9zXDyaLvGDR28cB
SaNFo+UuNFhTqZsvjSVLIp0hmwEFnLFPxoyguoq8xCCT7aNJDrL3GO1uEHaS1mZ8
W+ijebWBe8jxR+n0e6nn4EHV5D/narJsrOwTOYa2/kHiVy0eMBuH7womWrzERB/5
B47Wfvbt8Mqj40T++O5gSd5NYAoC0y/xDgmFmrjQzCvDZv7ycCmBRWQsO7xJ0WU4
ao2fM6X0dR4H+Uqlww2Ef9y60BVp4IXkh6KGsWNrHWPtPkYkjCtEILlVVEfysk9F
QTGhPXhEIisYoLww5kwBcJSVlm4Dj1PWO+BNEYHwT77/skutqC44C9KSvWPyegxL
vsOUas4RFgEJFTspSzHQyUGalXYK6XbaRtmzesZrSYZK6gjkIuWRqFt2W+xAYK6z
JTlTaCtOsfNj8+ztJeGNkkzH+UlaRswCYi9AwrufMEfUemxKaocTir9dkfxJ6Wrt
aQZM+ufP9u/+8cQuqyZdjWK3bVQMZ2vdLH6vkJzaauChmJIRQ5jqaTnUQRscr4kw
KeYuAkwfMYtu1QTXt2MS2QH8H4PQ0xWoFYeHmOsoI6Sqk5Cf5DA528vUhnrKfb/3
/0T6Chy1J1ZumTIzMt1f3xnK1k+I1kJXQpP/H14+0p7I9QWE/OcMdZAwCPpZlqG7
odgnf6aC+5tBBGP/hw+/UNSpqq8KhpDQZZB9QdvcnU4TQvrOaeGFWeb91uyJogNa
j6jJNRiYPgCfcreALpCuTWXAxQlINoYgTOtqgwNHmmIgiQrLfdlRzcyHUC8ApvKD
jQ4w+71N6D6wxmmzFk2KQVVsLi6iW/tZSw85cAyQedzXCbATNg1Z15cIQvXUfsaA
0WqMmvp0cckM7xtrTnzWHrVZq9b1PgJ32SjLfZLZimkOwy1p/YO4Ib/OWwlj6Y5h
pinfzPSQO7syBcAuRwe1oO4ecEn2NxfwVVj4FaSX4yxTTzcX8SuYeCbNwmSpqoXH
fs02pRh4vGx3w2YfiRm3tOPaqZkvP71dmrdLjCWB8Ncamju1Dktk5kBedayARvwR
ICTJwdL6llUjJ/Tu0FttLKJI52gpplpvp78hm68ZvmUr7wJPJIZ/B0B9h5eYk8Be
3moTVAQoesJHg63k1TcIO4L5W8hWkccJbzLT3q7amNoi1Pa8CzgH5+BzTlRFF00t
8cpbEhqgQSE/4vRNTDkgxmoW5iDfh9syzPI7J0mU5q5Q9n2b13yUJb+gXTVTExW6
bJXSGIDhlUjaRloAeYh9fLMawJw6tP7pO8WhkvHOAexT2ZQKY/jPfEFLAm3aDf8Z
7bFhmlv1w5vv/bTLUxeLUjeVl54ygrCtrXRJwHYDBwLI/wVcbvq+rx6+4WZW8gLF
3j9UMsY5tKJ6j2hpN2VVVUONDpp+ujId16GrkAow8LEgoz/FkUh+jVFxTn7BKaXz
2SZm62GyufxW2RpREDKtkqq2Dd6HkK1CWQFv0Jd0NFR01ZigXfeRGKU0x5zl0tqQ
Q4puIr6RSPHtxFGeL26grIHMUNylYETcTJcWzujN01uzYrTvGWSdo3Fw2UZ0mknH
wcEOkxTM6MRKAsb0gsty8WXWH26ARx7H4NkRCcE02HGikbg341AyotvtuWuSzqF8
2sO5EILeh8X75L5EDIe4wz6mxzbWhViHSLxISO+Bioy876ckG+/zMjVbojERFBH2
60YofvaBxxmrBblFQz2lcFiIn0m8+zFQo6cgYjEbmcRN/SI8st2LcrD52duNvUmT
No4ZF6wDMHFjrM2Rypv2nkOvzMvmSy+SPNnpG46mx0qwFCbt+deZjQ7pbb27kp2q
nu9TpjOBEWBNILciHKT6YrEzXj2MEbS64ob/JdgU31ernYBz51qvm61Ax4yUG8JC
weW5Lbou7Mfbj7QFfF6IXDCEgGVQ51oF4qmoFZGuhU+7gECacUGEnnT8WYkCcaxs
VUcjm6WZmPQTsQ1bJehZwW5d5f3O7+yPoG2nA/ZKh6NrI8s3vN9qzJDsdnzKZLSW
dKN4hqliD2FsB8KYJtz3o6rT79lVUVgMLFfUlqXCYhmPjjsv/cga1NdrvNcg43Y0
XkZXu3BDbHXNyxGYE5Kl2foyMxCUfUmLOacZcMFVI+zCyKy3gTw7EWljZQFEXlPl
42kT9iuPCQ090smfPYoQ7zG7zhI4DsG4xcjpJ7GC6kvSvf9F+VZHIx2mVjyjfZIM
UYZkPSW/MOXP5WuMWj0KwdM7539T/bJCCqHlObnTB/HrMTwJ3fCf5bP3IxabtGsw
1SX1m2ZOiab8PapC81CqqLAmXKqC1RmnmmWvuUeT7bDkYB5INEgMfe50/lSnaOVx
Po1VloJewLoqREl0vCouVMMrm5aPHzuuNW4zZAvXQCd8El/4EwhsajYk94HUw4Gy
giT8TxTdCkzy3NsYSY0a8CvetEGZGbsJrAogWVvpe1CMu6iZjEDyZY6gGVR7uxWz
QJOn4emw4Q0FlcUdHh3eDyQqdD+rmyz7lArrBGa/IOvq43BHzk1zVlZHSKHNfr9z
cm42b4wPwueywkr8oBuuKeezO6UZnz0AYyLr6RtOLIEWzSbe6nNoorI+IVMsNILk
S9tmWZRuFJiT9BWWf2E/3BtdvY/tXLsK71gyJqn8fqlLuszO1SldE/+FX/Bg7Se6
DpxG3Wv3V3Z9Hs9VPCOPhOG5XkPK5XUzj/FpmOAfFYY3uFAUq05KTJzWAyozdCSv
lSgOEQcKMmeU5PBvQ3OEr3YHrebDeOppqno993ERhgEW+I5AIkEkTjj3m8Vccw7U
dBr+OSCRB8qzimRBavPul3g8nPpjyJBjs0ZOFswRp8hWxXgEQDd8L4xy/bAgu99t
RbTWf/hLof7sSnBvSjmHvnhwTNHLbO6TvLlKGPauGX/1P1xdSvimJPCDY4PE53jY
GWJcdXxNLjTFyjrtjkpJc2W3OblOXyV+aj+LABPW4rw9r/siZ3OW9b7XFLFRCg8m
euWDuVBLfE83Gu0jKJHVqI9yB6EW1sO3qBk9x/UPInrHcrMN0gghTTHt9/MLWHf7
GKBsPuwMxoa5eY6nWN9jsYCOi33BBHqxJPYDG/+QzdqrHcrlQNpbRUSfsh0SZW55
O7m9hKVuqEyi8oHnCp3Fvg+/MltPNgB8kClGHDa7cn6jEINI8+lAUswEptQpNPFL
ICcb+IXPePM5YzH48EJq2eUEYnGe/PNWazdPXoe3Sffi6UWiL+A3wTx2AV4HwJ7M
HBb3AgJR5lCrP1hmWCIvf3ezcBZG2pYJJGqlzfGXkrql4ksdMkb8+fQ9lBFMg+01
Kl7fuXbpnr6k3MM39tsQojUeauWfOflAwIWnp6bHku6f1CouiRdQUaxRG3cJA2Ug
MYYH80sJ5ujTYIElQk1rmtlMsTZnzYXOAX77cPhBnya831WkVRz3m8xIfbJ5ugFp
EMXVBXTvAr4VxGb+OBHB/ZFmXhOpHB3kIvFwA0lSgiGFcRUKXXfMpJdWf5fbTvT4
XSBYoofgSFlsQm4MzWpYNWY6M14jSHzmNn26czdQLGw1ciTHd7utNPnTR/+zuPC5
BxoXFdpn55WcQwswwj/Dm/QmKuFJJmCPaHauypNpWe7eB8eBiY06CHuIaJcVS51c
Dj4aX2b/EVJKRFSZPgNQEJIeZzKNHktenZUrNwGqW+W2ZU8hbIRQprCnxH10LeWa
s/hHgjlnUwnzu9L6iK/3dxarmgss6oQqTGjxn2BZ3ttw4MBBfdj/d3edtDIdEgSD
jNEZtNh44wT6L4CGq+Y+8QWIPDtQo4LSlXOiGYFG4BiBd2o+WkSorlLcq/jzO7IL
k9s3tQpCk9FOnFnCYlUkoR5j7gDCa8YguCyXUuOEvoLGJJwWT9YVSzDw4dMpK3+/
ywEyZelyMHRAkTMu2LnwUs4vSXW4IYwCWORETB89LZ05gW5n8XgbgGhIHy1AViHi
7ehIr1PCZPSMHLjyA7PgCV86kAIiU8w0knjaoWnpnFV2c/DlLmBmsYUolG8m526r
gjgvSedPLOxQ4B0UKHWNQU/WIB8GwZqnuTlb6teI8oyu5dzhHOnDru3f9k3qMRce
asRB48vKY4LwACNtAmo/MdbN5bafF9mjxYoKbLvW9OcNBLkwD6RBay9iE5VcZM3C
OBZRohavdeWdF5pfPbB79rzte6EPa8pf2ToYoMae6peZG7mZQ1eTtowksBwPwZLJ
F3lv61r8QUnz8f+F1mpwd4/3kFHl3bh4wnkIF1WKGD1mZED48AdbW3v8By9SQJNx
uptOdMmG3PYjTFnd5QoX3eQP7n1xj5ddk7doD1E+Hb/+bMeIvqf4vbnFU+aamvBL
sRL0LTi37ndrUMqURinXKRKsSrBUU5f3fC/CMnkmVpl3kf3T8+ygKe1BAHKzXILs
DM/21jRAS4dCBckmss3yXfmFu+tXYNOlq3gdVuv5lZUgGS0H7XDWnBQBcizOaqUa
HUB+VJeU8kqxFIPpBDmlMP4XhqhvTxq9cg5Z135CWrBXBxBRItTpON0xBVrIj4YL
XFw4hg3zk3T034lA2bCu/4/CjUHDNCj4d8ofT9ApvggbCw7uGQ4oWK4gMgvucFc9
Jjv7ZhraqxrjbKBHtlcxwut5xaXpdCUnhk99JKqMSDoCpIjTfPv92GUDCzVuF6f4
cRuxBaA4T4r/SM/5b3/QVKBgatlEwUy3lY9c1xb6z5ZN7cUPTnk0BroPrx0dMuKA
dLPcA/Y7dypskitLwJo8NI5exdcsZKOpkD/6yK5j15Ad1pBqFeMx4j7VB0JDUPma
IgeNVtqeBHKqCwv5W28zqnXlLMNUByy6WtaA+GDVsvwXiu1y2yj8bgI+B3aj3u4L
Mu38pjqt5lVOM5hE5OMgny4LUx46TvOEGxi2J16jZRRDSaZ5Ps10lXhBIMCA8liC
aJMglb4c5Vxy2tVleut9oBWTiyaSTY3BJNwVQ5IKwjJyYWhkwd3nJFv4AI1KaMs1
lUrSTdKSnzEMjSduNvToof4aimDa4IzykwMscmvHyTlm041aFjauNT3bw8xtfweT
XTKI58E2ZAA8Rww/xHfUBMeb20w3F6zS1DsvLZm0GkenrRTdtuG9ROXFGeNf0gxY
v2Qhi+6EmJehABtkQ7T40pJ5GJl9IxEjJTs3WJk8g1A5X1rFL0IZK/sljaIYVlSA
3RQ8c8LMrm+xB9JwrLUQJ4heyVpuVsec9RBTbbmmL7z8CFYR6LwerB8uCoBNct9+
QMDg0RLp+XPuRfsBNTjGmP86L8JcmL+tSTRl18kTwcamspy97G2p6lJEtCYdu94b
7bYtuskoUlfhf4srUIZ706nKbmLKa5/TP1XBQ5g5DMNGlJ0LaO3B+ZMexxfEj6mj
wOyc/sFmqV/PuFzuFJUIshMer/NBuZWf1GSdtujSwswYFCVMrxS50w065UlSjPYr
HLGzf2v5U+nPvHvI9PxhyjrVawjY8qKQbMAJNMHipkLUx8uX+Rk+u7p951Dke2Py
cTSXYLU+p5LfqQAf+0fQpZG6yQyddT9ywMTLOX8EJutIOxebiBL4cXXiKFlI2qcC
fU7Ul7lbTh9Pf6QDN47FM0LC6Xm45PQfpQLx0JVcIHjl8LKC08filYILTLLxGECy
UZwc19DwvgNIHa0QUNesUW1uBwA08BJuzCrdYAkWZ2jbIoGgy40k0i3tEOIVn3lL
yAx+DsTknlZZZizzkFYzvud4iviAQgRQUtYOu5Tfs33TPzjvqoJfcCA7Zvj7+XdN
O4Bdx47I3cZPDvHzTjGnmN1ka68azzOpOkt7TD7Yc1zR8cOB7P+ESGi71LOWo8ym
zHcIv2FhzaoJkSBo5ErxG5D8sNLkz5BsyV3lPWMF1cTJehAEnqnpUESx1If73hCI
sM8yyRCJ1oIvE10ZkcN1vlvBXDsrDH+dI0BUhKIXnoQ6S26vA5WtwTiMDz//Icsf
fVPhcSyvgceoTGP3JuotHUWEoRymz+FFXiB9XWj0YT5fwa6a1WqXRMFTfz1Bp+Qi
3fz2Ftj/0f7X8ygX4EDRIkd6VvKw1t/D0oiq6aYitLrgTXx4DzAfqC1HLuWqO1Ib
szO0M8LOrCi9CX6PaGmAB6lIEntyTtyaefcUKqE07dm4XP9qyZEqSVie94B4mFVM
fO4N4MoRSkDcFTuGSWFrd0DR/f19B9/5ccOrx2dT2spkPz/nCfuK44Y3rTBTkKnk
ejY0Og4EvuKRPDUw8p5NXFDhoXXq+GsVqhWJJnC4jo4YZa5DD58tB16dM2XmE6zg
hReZTj1yeFcGRPqJtHbg07Z0nbr6PlUCQ1e7GjHMtxKtSDs+9xdvSOndMZTHEW/K
nh+s/tDJKFpc5WXJ5aUNqFZu4wDe0HkSV+BlZ8X+c1R+f+vKJ1Q6IIsN+OgVRYDt
6Bd2w5MERBJvsHps+dfkRJDooO9Y0z3PnJzJjVSwMJ1hhhHZeAcQf4Zathx/D/Wp
Q1WaPQE1scF0ZTLwwF/OScIoLmawYwdun8EbZePaqVsB9m+uQ0THCkXQ7FOwa4d8
N7fHXcwAjnF6XEq9mDp91MezOK26UmRck1H6GXLVLxeUDf05/FZy9RYU6znUlQOo
LrJlq7y8NBXspnVFD7QjPnFr07xIq3HddxrQcPNzrsfUKhrAWb0m0fl6grAU+cEH
WcVjuPlS28xkBL7zyyZ1o6cTgdWR/d+jSBHg3znWLLFByffLKpT0j5NzgbWAe68T
HJxjOHMBP/eeUeNOCLdrRzDtAxr48sRtIhwNOz1ZIOILtBDpXxUXBwBb7TZ76qPK
hCxD7q1WRN5Alj8WnWidq+xVk2eID8dNq6uQ+43riyVdorlYHvoPDzdQBHnTCNgT
jCWz2L/r8SYjmzBdexwDoSx4EiunsJsBOlChD+3ZBJycOBvLbgQBcT0RBQdpZog8
ssJT7ChZqAOyvUH5U/P2I3FSLyet0xZRt2xQmard+++goK0O+j55h2qe08eyHCkF
SNhdrIqnYNjdUTPhoo98BeMJ1S8aPr6gZTvxYYN0kjoqzDfMFcaEoPiHoWPgfkk5
71Di7rqQ1DdP/itqz3Cn9Nw7aqsDN82Vh2WkbPZxtPwJ+0OH/1GSCSJYQ6LraMJ3
KUvVlR6q1G0fMsPS492AVjfVDaoBRrlOQU5GWzgpUbbgKHi77Z17Z8OgtUTaIF9k
YLUvpUbyb6h2TF32pETj27aeYB+eFuzcFJxovttjiW+nnDdjEGWh1dXz8USKE7NN
z/azX/+jajMGL0eQiK9UW2TV9+dDWPfA3s2jPvhcPjk3OwmrVzSoXukvPpCoKiSg
fGSqEW/JyOklRvwlf9XdTGI0i6e1LbIvM3Wny4GHQ4quQGT68PO6FrDjuH0oN9lz
kCYJpsmotAyUG+EdZS4oRiSzNxPromNdYA/de3j0AkBFvq5Uu9pHHGOqAgz8a0YF
vx8uIemTVSUuZE7CEkU63pKDd74z+O1maolOtt1+K/XFGWxbt1p2xAsRp5S45DMq
SnBS8Flxft+WPjHVSw0ZIWVaPQwqEFWvJbeB2bqrJBt4OyghovY1ggKNGT3PLdU7
krojwIalpIccdcPqBb+IWoTN8SYlEQkEmVE3UFMllGoVE5dT2M5kvzUutrI2z9/P
/LzkAnmcfduWW0xJ2ffGvyZiyiMujZ4hD8XCZracc58xkx1DZa6DOmBYkm0cfAXz
N5lfWpvmHawmMDcewsKUwSqOGFWXoCscHVAz8w5/S6vsizNeRiuGnOk1hPGnaIjo
IBf2Ean70E7TiXQusxr5xjOLBsizLigA0vdWK9Si8G166eg31i+RJ52hUHVCjJPR
vxUJTpWVCf4Mbc6dTzutIxD7D2210Aj2x6OQWzbQNKBVSjz0jIcDuJ9TLUDR4mQS
lTbz/qS5B5Bg6a+Dnepn2BHQgNJcvmFI+ogo3vilz2MUJkc/UFlfNI9y0foTlGiA
yVexCyKLpFZxMo4U3fhiW98nYBnYz90z/H37hAqDG3a3KPYsXOPONRDONGWOU64Y
go2QwIfAr3p3dneF7BOJrUJ7dV9bzeVJ8poithnh6uF8Uofzoj62MN6AGfnr8AXd
S42o7td+TsrmNz42/JkitajnUYQ8XrqMBhku1KSOYHBgq5Ls+Y7mGhTMiO53uouk
13zAlWg4S1hRUa30EO3eX/kz/YNZtSch/6S1BNLAYQs9yC+/Cn2u0r7UFNaYH9uF
yZ+7j6oz83n+IMzP6857mMeHQkaqbrm+VzFAkRe9c79ANbaq0jSgQwjp82q7zTaG
nz4lTB4gkTAnL1FaoLeESsV+5yrQHxNgkCg+/sY2NR3ppzIM7Y8mrJlZ4s3RrO+r
KosTXPShJNTey3LDrQOgg+NDwTvp93KDMJxBie6m87MO5LwgfgUe2PaZ3YW4tEHo
BjZDz9ai+ZlHJ8mehxuHCQiWYf+vUB4lZB00qJxTIu9d8nAHqQSL8MH33DKNji6a
rJR2eHnSpapHh1f4AHt4A/eOypEwgOhnz8a0vS6bTvckQg+HnsHjMp5uvbyrcQi7
9mCd8vAdRP23zn27Q5UAwDIXdZp/UDbpU/Vh3iME1qIcSJoZNX5tHTcTR2qtHvJ1
aLUAvJDAG6h1baue0/fF7wy0Xy/aWPcbaYnuAIv/wS7adkNoVO8N9K5hshVrtXMO
c8xqFpv5FwcnDb39/H4P2+RkSQJSR90qkUSnPIvVJn+jbYJZt1cdf1fE+HeZnfk7
mRxyu//KU0UqJdZep2D7twiNcbwtSYe2y1pO62F3KUEw1LAILa2drM+Br3ZZw02N
BQCKKuXNjfjOVZ3Zi/6waJUSNA32sDz42GV+7MftjMxGmd478tcb1CqS+5WWFGOk
UPrMQx8sM1lcyNugBqJyhoCL81D/T4MBNKk2LHzEN9/iNiuiuBces8d3FStk7+N5
2+iU1+5wWdoMT58QBb7P+9prZMzRoemVEOGz9cQ2poBCQVP8BcAmehdEuuFBfyqg
LxpN0uTxqPURh91E8dxljPmVBNw3pJQihrMO9otMM7+azooamJhmZwIKMALgBbQo
V+uRFWXSO5+C461+EmXJGOuspBgtNZrYaiUAyCbvE+2mteJBXZVrVo+uuof2Y3jy
QALfeaICMUr74cSIYIUUq73EODshlkz6J2IucfIUm4jwD8RMCHa/IcgzqOfNqyj8
mnLCx4LFdE1vONGGsovKZ2CdYZBE6ugpfODOvnFayWsGq5ojMsKowQQRcPzBOIcl
xCa7aPC6UnUONByWaPc66Y8aXATUwKBMDnmeJLEvhOSxvGPI47PXFExUkmmb2l/s
GP1XWzdXLnMLmcSDpk1xywDJ1zLPv7LCmrsO6bUlHQShJ7OKP0Z8u3MdwKZjMO2o
hiDoY7sklJUilVL3kS9EcP4D9XHXqElsnewvMWKQ2caDsztny+W2kMPnU5JUfXXl
x7g/AHOUv4u2YKQYRD5fQdpBPMjiZnUUpWa7QRQOzLa4st8P8iEcvWsdtYR2G2pb
oafi4akMomxSTFQsnAYzDLFGcEeriIV0U3FNe49AQ6C3Y8nSUexY9MVKKQKMZnNM
4VkTj3r/0e1NI7REVhuDnr741FQRVQ0m2clb2XeWC1ZAdt1A1jlgJh6nbh+9F7Yh
oVBDdySjxn44pwDR73V3SNwjiOvz5e8S4xW9uLJXtL/uAK4wVHlT8xnL/dtF7kmf
YLZw01JzUlUQfgeYio4wX5Hyc/mfjb+/X8+aZe+JyMwT5tosHAiX9brYxn9tjk4A
SsgxAJUJhu9wW47fI7WJ9BHtRxy5RxDGeP1pmYmGV7ea+tdMPv9WZjQyhDYdUSfV
9YwqaHr9a5JHJ9FHy91phjgQbYCTQWA34gwOAmIfQFZHlgD9BiSk2epEIo92Ghds
Qyp8FaHVWKQTCfjtepn9g/JnTY841UzqzAwnDL7SJtkeELCRMghjJox2ZFdI1KcZ
GnfPMi+vRswnhIhWeOZiYQzoFlEY8eG82+smfWytuH0bEb+eucG2UOvHaT7XbUU5
iOkfzoSywLGt5aF0rlHkUvB9Vjp7VlNls0SNwnx9fYACQuOx6ObXpPDDstwi9zgF
VjLTD65RVy3LURt7KCPi0rEy5giTLquYTcspExmGE7dnRhoxgOQ9j2DWwFkwauWr
kcQ4cF5OzT/Wbxc62IqrMt1/5kbCLpcR/4Mv+NtRfRYoy6b+ahgAOShEjadSVQZ1
nNwU7wcxwW9mhIHlk3AkdIlgBKfnFatX1l3UaLTOEX3LkpcuFH2bEN5GEm64+6Ef
FLCSsNrSt+XyOQgq6h4zTecRZ9YYye1G3sA66S5JbIw7Ta0sk+rtzEQxiteYzfl+
JkFpQYF7bh1zwqmCO9UwGNxrnYPvxKSeW1o2tZxrA5JvTxqHOD5ipU5Om1XsBL2n
YBjKNyb9FNMk3HIfeIzEAyemOl/Oq6zdFeM+gnyWYSICO1qrRdXEGUeguecqntFT
x2+0p2lxY2VQnNAnDc2jhpf1fqMbf/i6t21+uXfQKVcHvunoI7BEbGgPiQ6+YWVR
kUVbtVnQxpZ6qwGOAp98X/AtqLGBxaPb/dwF0n1O9DjkxjX9GkaDqmt3dWgBKW8h
1lP+chynTRcnvXGmCH/FJlwc91LtcUaiS1qEoquUdQkugiWcC7J4v3dBuXrFB+uD
LXCbh7tvJSG6OWU9S4l7jIcEjxkIpf7WvyG16Hw7lKGTMC+ymiad8QBUPuOITiTP
VAGmgHCSR49pXgJ3EOmodsw7LTqWmYHn60mHJDfu6V6eqwE8GwRSugkyE/UPD1k+
vjYJSu3Nqey3vRPvrfC+qK4JmDYSYeh9IHa0896+x2LFVMQVAO2KoF/I5+B/XP5K
orR3GgMnBbPNttCUOyJZIJKpVazOEf+KbWHiP76Xon350XEZ3r7zf1EhmRgDQrWi
HHwKSjTl/djONtHT8nhfgVGoTFV9s5oyuATkk/6V78NZzkkaljtMh/mdOackkI9e
/lbQ9EYRP7DZw8qcrGlCCREK4FowP3OJ07rUWeR9gME8TmCZCVqiLd2SmvdyZLrB
De3GvMjWoafcRCEjxnQQow8thA+zeS/13LwIC/bS6HkZw8ZuF8C6gLD1FbfaO3bV
Jh8DjIFalmgeayEPG7kF/vRc44oTNxOYhGAi4aygNSSF3PfHxLvgFXYQ4qbjpeaF
JcqUzWIfen07Rr+ZVJ9IVWQJeUdfUki2yLhns6aMznPNoj7+v+xOTxeVUWFvhCTW
9mhC2SKfzC67YYqlrmnxf4LHD6gF4QWRd7+LPE+HorQ9/HZcRGJsSCWzniq/AGgz
TjHB32xrAp4lF6h2pqFl7wwlQthAJMA+KwaCMFofS8mCaQS/94DloM1er6/ky3WP
THqc3/y9ZNwhkVL8pq5qFlcmsLNqBki2iMFIhMnFljNTOWR+ifDKBKdkeZnhtaA8
V6avjSbfos4a38M3UZqQ0u+Ufj/axtKq9xJuUx0aCbfCp3JSAJhhlCo8D3/dw14M
QIwpqYVrIwJ8Ib6+dX3CBcTMPZ8CLxFMYiNvKk4dQuuS3UoXd62HRDsdQwIrKZzd
E8dmTN9Rr/7GkY0AHgas1uvm9xYqJx3qvPuAypFV4+TQE6kxb9WFhS6MFLKfU16G
E2txhyG+Li4XD9uDmUKVhGwj7a/6Gmb/sJrOvZW7y8ZW0bcgdrXoaDajzGzk3WWd
5RhJ6us9cELDxKbVED6gLlYi0BNwDwqNHUaaxTqfXnyyLyrIkX0q8PpfxYNo4Ixg
48K5zTmzogTBrAKX8e7E+UB3nneG7dTv8D2iOYo7rMyH/aC7cRnNgZzUEKJNqpdK
UJkiVIGSPT4Ngr1fY52TRB51HmajWjxE2/fGFosGcSWtLRr6z8lRyFB/Lyzyt7ss
bXzMyCXya8YYaTDFIVx51l8V9khIXY+PCOxXEdznYVCa+huRRtJrfoi7oMQG6CyB
SjgEZP4Lcd4FMBoVAiSXAZoRM/7ymuqirD5yKdehb7w9jX4GqyFxyJDw5vcNEQzz
fckDIyK1BpC58xc4mWQOm+z0iJVeR3VZcNKw5MqWo/i1jQ8+IY+ZdAuIAlmD/l4R
1HF/82/XCPEIi2J5nK67ONzN3UYPEUhOtCIXysWap5sZLucQfbvv54jLUg8d3owh
Js4Ax9qZOsXnCwPP6M9NZBkVuTWQuLGQSFQPlmPcH4thJ8KqGKUWLVFQfk4n/vj5
SROzgtcG4XcindETtZKiqYdQsjSozHcC+8b/1hd0W5SmGt3D3oR9AKaykw6JIPBa
Mjm+tnvqFPPjNBSAcSfy5TOkPJF6v3l+7kXFeytFQIhnzSosoyLPuRkCQLsFWRCv
qRpxsV/83M//61jb8jliUI6GjWlQ5A2zB1zqWxt7KfCuWOH0m4qTyKjRSLSFqBXy
zovwhxIulTv9jR/iyVqAft7Tw0eFwlg9F/ZZ2NZrTOyuIjwxZPTdJ2cPJOlVFBNK
5kUlQjU+hfWUSJisTxllIqhRTKfLf55LdMsLf54+37CcJyvO6THi/PDibFqoM6HV
+QFUXVeBaihf/yqrZ58CmTLpOalmDk1pk8qfeg4nO5Mx4EEZa1LafbmLp4C7OZO0
j16PMi+96u35fHp0BuolFkHSPa9uMP6PKMA1PN8XA0IGSl5FK/mFzWWrcH7pMo4S
paUJAwHP/q5W8RU6h7tqsbi5OYWkT06W03NzXmp0rJNxN75xfRz4wymVR7+5upQL
WHR0jOop7a9Z3kKimxP9kqY22I4SqCeOOnjYW4lvxgsPWf4VwZ/vXsMAp1L7Owiz
e9xwZsydsthXtltFVVjVg7vjzRfI6ttmM5kpBiNzuWXw9Vvfdrhn9FCk/8O6RNTC
ooKmj4+/oXe3XpJ4pyDk/Yn46XkRPMXyoOF+5sASSCzk768oMm8YNhgLq4YhjBgI
vmBwmyJ68GNGHHTpLcjcpHRKhVs/gZhlenhvRCKRa0OhG0BZYgF5bPYRsCautD91
Yz/C2NSdUK21GZLuLHvIM6s5UOLKPN9/K2oCXpbK5eeCveRKNAtdtcBx3aBXgHPO
X7b/fnGerE2ooqmw5M0o8wK777gvBiP/7RV/kz4f8qlgoLws1Vyy/e4kLu5NQWMf
PRMQgbIQHtGwWk24yH9bh4/Sb60zdCdI5pNDv0qW4+QdKkr8UyGX8arvc8Dnyda9
+RCP3D5e7y3wEg+FM4EYYltfqLKMSl/4fNAbC84SnsNyhiUZCOofMISe7Fk17yd8
ScwLtqazPPKhCjadjK7u7cF7u/feJEhiIUOdgoc0Q7ZnZLGfVqvs+U+9QrnSZf05
DvgatSUSd7yI0ceDayjs/N02XmFGsBIQhhvWpyBI3s7ul8yK2Uxq6Cks1/BsLolU
aXNGdomkDqIBUjv1W5DgsDoOpEwUI1nC7swPOzjljjWLSJstV/33eaBRv/vVVlPI
Qtn44DN17aJOc3x+LYnaWrWb7Ieg3uQYQT6523LAh/CCHohG6ByJkyz63pRCxJ7H
8DttEW1P6pWa+7yc34sATxf1frkR0VHZ/Snn6LmIaQsGIU4at4R8Os/X9muI/S4+
bpz8bWaicJKfQL7TWTFpI5WKcVrxhox8bQIKLg/dhHTUJzU5mrKe5X1jfnZDRXT9
TuT4JKdL3izbAXAHHzYYFnCz4enMnG9ltasInXB+TGkNR3pYovO9Fp7DTdR6JLsn
hBqJOpDj5ZNGJDUTcIfkEui6osoY3hptu2tApAbRP8dV0hLhAIYCKaUq3J2bwesT
ESA3BP8NeXZMkTSgSEqKJa4x+bFphcnsn3iVhh57MUZZQp7IVJQ1UzDIvdw3Un9A
Q3s0HgrjqkBrLE9hLIx/314TiLzfSs4tIzMYKkLufgfNnhLcCr6V8KPyu95H0h9z
DDt2gRCTjEynFkCrc4MUOVS+As5sTH0dM/BZeYWCazDm5hh6QBInQxjwu4vGAOAb
b2gS8AU+TW4v2ohyItoflremMeqjNKutKQ2EEOIixSG7nNY+M7+fE4K1UJLPHlwZ
J0CE1J8S/RCJjzYk0Wxs077WIEInBYx6QAtUFal5PEnfVl1C5AuLVUNRoa2gRkE1
+D+tkmvmOBIvARSnKF/8lJiVowyWTrGp9hXcGbWi9vpoFrOQeABUkZEQ6Ip10h/Y
Yyp62+9TafDnPXHj4Tc+Hh5xbcEVfwrwtXas0567/Z5IYXpqW77lX4Rdit3c8u6Q
J0/EsYB5qogEMGS0GVuRDEd5XnL/AlcW/fOMp6gY+pM/+SyRI341dOySYrk2ebVl
rZmUf0yKiLyo3Fa1wyeCphtFYXhpNhFKDC4RbYylLZDK46iL0E7Kh7+Me1cRyZXE
c6aA1C9SPPFNRsq+CDCdRovhRDOW4M/D7EDrEyipSvJ8GP7YbXaZjEw4FjWM6AQX
iXO3Ml0HqmMCrI1PYvr+mEtqW3a7VmJh7PrHjtAwcMMBWLO2nsNtVWp542aRhGy1
JbaSAmV5TlNHuiecqw3SZ8pRArzuq/oeRCk7dVGIOEXFwgBdbaFJ1sWeygBniizH
3iHdCoPC9SnduVY3tjo9zs8kVkYTJ7uJ/PLZX31/+5L2PMjNa9g094xFzZRCIPRn
HFYyyMvuOyRLQTMrjmHS9RuL9PWSBke8+E34Lhn63k7Ng2HVPM/+n+Ab5PLpaz+U
fqE8E3TaaHnoXshrkdKH63pHBvUyYEJvnphKk+jDDy2dorQv0mW9rRFXiBncadN9
oH+0008pzuzJrYCMBZI2mFfdki7hW2PU/OCJONMp+b9OGrfAKteatXF9DABNBeZN
I/51Q789NxwZgPa7bmqBeSZ258dBYErAkl3zvanTfKa6h78WPc0u0Af2ra2+tzXB
Kbl9WOkvWIlE6/+OznjXHrbdezRQjDAs3SmP1hOSsZkZplXUFoeyJE6zEPW8/9hb
eUO7AHAfe/Bb/sGKeq2GCwHzZGXtamxV3EE2lYblVyVkxLgelEPlBxcklj2Cpbph
dzX/IpbP7ShocgfL4xZfAfeuHNUQ0JZBPLNY3YWefg/UW6cMjWCBtTdP5bme/gMI
sXYLxb/eVTuIZD1nQxdTfO7IlxnvucAVgUywoSp7Y6vih1mycVBNY2iVhf1JUIxD
9XwXs7pOoTiyqb5+HgAi5C5J8ph8clTyykvSkthDblJBeK7Q6EF+owjALcGAaXor
qdnckcgY5kBXkIJUa47PCMcwFDzZ+FpCTBP5WKogBJZyfxK3ywX7YZypXHv1Wn4r
+sH0RTpMc5/ayufpKykZdyAuMDOgPFFdr8WtQhr4RdYngGS6VH4SL8TILoSi1Ep0
j5YjHKGRmGbXrew4ehSP26VvvK46SImGNOXyE4j5eYByLabUQ/iroBOyk3P0lWTA
CRf2D0NZ8o6X4KNGUvPqzmwE5CHITvDp0+cOfUnTQ9qZZJ/vZfurmsWXeQma35Ic
YwGZrqdQW9S7NAu7ynuQYmFlGWnzFnxeK3vsGfVA4rbeh0tA5tgy1FOPWDSVkhpy
HjV9ZOrhsblYvdLX2/ibgem7KomgJIf/C8D8myISsPkrfscR588hUhaEnxJwYkR+
23hJtS7jpSGpRqtktvGcyKwLPBjUK6ZnwJIf8PPK73A4p/dTXzfdNxC1VKSQgHMi
efpKNzcXBWSON3YYO8fsJISlqf+gLdBwEP9WVCEo1sI/mEAwrzSTalDL53Dyd5od
Q+i/yRNANQ65AOFKGS0ub9F8Hx010Cx442PlVJyiRcoZO6YQ0QdmHF5b9qcMIbzt
0pkpFlU5TjrScaE5mMRxeDWQQHbkZ5eB2KUpW5g+dwDt3kQaHlLb0XFtxyEQHlt8
YJKBf+PCCeD+23YWsiy6lVqYZ4Xzx/ikvX/oBxZURjTmooNHY/jSOHAsjr3GSpD1
Q0y6BVhFmK4oYfX7f55vQZfAoG2wiMhKmPKZe1oUGw3HpHTFs/cyEeg7Aj8eHXmj
Yy9IOrl9yC5udKuEhulb0D6nLDUN69rDeFQLxpJQGzdhtfABLdB6zn5eExV6T77D
Dn/+amOHgGxy5uttcBadCOnDfAQnhyAD+/5V+o6AXYyQm8A5zpBUX2jr6rNlHY3v
ZD2qEs68+xpv1VT5A9w7LDoG73Eup4GNL1nu/tc71rwl6EndIxFhMKzmzm2Rquyl
N3a+FsL/2MozUflSkCBnSqMXRqKP80zIJrfIpnLqAr7QDU9sf9MlaVcEH2TE7PBh
752KC+B3eWQ5LGWrkh3nbObL7J6FVTxuTS3wjPjoJH8Fajp0J9iRa1FML7qUgr8h
WMqh4asXF10owfuUMMuv2+Rzwd567B3I/RFJS31vA1ACG+UWp8ZfalMT5GcYV9QN
VeZ+oCY8afiivAc8YG9xeL2d3OIn4JCbLPs7ETRwgYwTd4yatKfGLyD8gR3R5s6x
c3Tju9mcR8Hxy6I6U3HqUyHPF8391/6CIXAc0nOeW7zlSa4W5OoDI8+wHk6RBEV7
FZrJ9EXzhBEW2ApInKWPi0UxAMOWWuwTgzBfkZOOivqfYCczoo4h0KTBOdi7CnsF
9SFFgtVRzcEqyyEUDJ6juGOdqdePvwxjmwNByy9uhAsBvjLRSMErvFEL6+gN0jnt
gDmpXL4Uw63rJlkPRg2KmdWXvm70W8eJxySPdhMesoq20Z5uDG4t1L8KQvusdnJo
4GUHca+1lpuYSh9Ws5OlJf9FhHXrU4QlYMpHOl136VJ1c0QbnBpIQ3ZrW2UaCyMR
33Rz/L1kDxrqo95Sasif4wAbClTESDKnYSM6wKbmjlktfEQyXraAkUkc8UTuqzp+
UWSrXH+hmFL9+lksbF2bAh1/3wE8e+MUiRn5hAsNEZeihgATjBpUdr4K5P8g8cqV
FMvQlA/LFf/lbOX1FzkTm5psdrlXNuTWAlux9gkpdMynqAL3x7bEcShqse4Vq+8p
4N1blpM/RV3I3VWq88t0Rr6K+sFHPgSWCvut39TCPstAHyqCRy56HwhgySDnkHmK
cWANbGiwVZt8a8lhxmeQKxsmySSXo1fPGTjEtiLtqTUvbil0xLyYXfK+SYDhJARS
x431Hxl6+ybj89z9Obtd4acRJdO07l5nLCbY5a4VnRHiiRjuuujLW7pXc3UPghUZ
FymMURUioq9zRDER2Q9EzeVPg3QITk13U6M2n4j/dKSHI88ttfYZYadKZN/+RZZO
Ho7UUPPzFSmQFk5LB3LiKLEhTYKrtd8pbRPFllVlOJVJwjogLMCpSgKuI64Dd1li
Y02ID1TubbYCA3cd5dsfvCmuMoVo4dyVwhVFVngX8GIN0Ig1Avp8Gz13eP2CORgg
WoKncQr/zDw6ty1U88tiK8TQ9HVbzasGlftwcInCC/0RSQ+5yuCp5YLjaqVYE+YJ
2f+DhlSibMddl+FkcAT57P7QpKEOIBpigwOrrSfjj9qMwlbo6HKg13kKoe3fuy/e
k48w8uKy3J8h96aA0XnSlYH9WRYcFTyHbu0rrjKJEB/2BFfO/L4QgD5Y38eTjRZF
ac84Wy/8BFYWUXwQcYnmkh0jAKbpnxouu14l3XHH+TkrwKWGUILOjT3qBJqObLGk
h1zpAERBRxroR3k8K7+2gPpdMOte/DgogZ3ZcK20PmeDoZhEES+I1P1jloHIsgRA
5rBqYaGXNMTYeC3AR1ksbf6OpcMCX+u0YbcxhZlXZAngsjpKIclX79gEaH0s7tlF
fAvJu2K1GEbabbFK0WBEdJQr1RDbINaNIynXu2t3HyQBeY7rzOrz2ELOywg0jM/G
ft8xWKXvToK5NsRE9qzezazf+rzGmGkxrHPofCPlrut0FGN2H3mz5MVB2T9EbMJG
BCGUr4jYNxTXFUeGKdOYak3AyeWh7pQdbsBG/UEIf+OPgsldc+EJFueTE8Kv5Sj3
ewZBt4QGd8rWDyDlaKz1RT66zFNx+VznJaVR05ivTxmgDwhOTF67NzvdUCTEnBev
6ni0vxY4UKq+sUm3uuIZ9G6KoxNcLZcee0plgv3MZeJQm9sC0NP1sWws2kxNr7jd
IfD5eKJOOjWSlIlJmh6al0LHgqv0G6EroYnVjFA/W18FlXLbU4YZJ2OI5y4aR0K4
qmx91R//lI3EFCVTOsyfnSjMFe6fUXp6ILFSYpn/k2KZV8hlpaOJH+Cco4PiilqX
jVa3DcLRsjBQhsUjQHydkh4dGjT4Zsn6SBTMTp6JItN0/yEoQz1GuixdGT/ktXNo
njgpMzceqMxEGxnQQtfjcRJ4abu5k4ezZ3cl/vsowt/NHXTRayl3YChqOHFr9jzo
YmYGV/K7lFYKnIJB/rtEsR+lMCFjh/AbrStoRQOY+kFogt3eWYT7o9Xp8mo0hDoH
/wm3x1bsEpCLSGGCSRKhRkweLxUk84LT3su3nwu7kQVIpUjma1pC3pRZHwsvv4Ty
8n6q7hYiB1XzUJy6i4of8CKxo3Jrrs6uQzVC5o11l8L8xfM20vwIVk83m8pDAA8/
nujv2ybm/y/yZXcYy4XB5eN3SWtpeMfc+yfZAa9yCOiSv0g7annvl5ZbYGFv/k29
fyOnR2Hj1w8PYN4vNouWi45d9I0gLkpoj4UUwILyptbR4dAQfxsWO0noL+6k2CJe
eOmoxMUE6ZwQAzjL1n7ktmzCvRfrZI4umJZSe5jTboDXWbekb0C3x6BQXeudOsuA
Q3IyZ7oUqXuREh7vUgMByxSZeOhuVRk4Y3FCb7d+4fAMZfTtUrLJEWehhd+Z2N/i
sBmUGNyGtWYAUEJc8Y1U97L5hi142gwON4ka3yTyvF6Zc13qY1yTIa/kt4i3y5O5
j1DP+ySHEdCmzWHBxntkZ0m+g+EY3rSrQfYrBlheYm6FQfKBZDL3kvsDlxDoieHW
Pi5Erog7G3kdayjD3G4GZbj3hjf1jFv22+WVF6A+U1cb0QrBFRXDwe+kCNbrqltO
iX9m3gqLlPupMj5tjoqOgbSEYychESF/amE2Dak2Y+INgN3HGxZq5jojGJUNP18S
JRxJWVlv5QUZU8F3ufpeB/MIJYi/ci5KyU2lHQCSBPqiXbBvQCuU3KQLzMszsISt
4xtsOCnyFoDs9uzPugjczIDaSe40Kkef9tDxbaLSdV6nDdppamAGdFlqtjTz+BlK
hf91q56nk812ItlZNa8uf7vQLq7mLWJSr7UCxoJz1ASokTnCdSvQy5RLPO3CoqKg
JOt32ek3NG9A54IYjYNHf5SpdBtZFKbUz3nWonFfGYcBfc+uUmtN0aivqMlj96ja
CLxPCuE0EUAt1Wo3a+9YFK8vMMe5TkbNcB1djP4fto36w4r7YYawYQXT6a+StZRx
fP7Vc/hkhHracnXpd5ILWM2F5ew6fg/Vk+tc+V1c/T8erd5ADYfIff0bq2lf6xKb
Ogu3DfG17AT+4/lxwlJXd04PDKkD3GU1RXjJG9mypzie10k+q0KhFuFbmI7YoScz
yftORphutTtW0GXLmvSfMxnQq9bsQIk3SljU78JkT7OzY5IpspkQnAHsUsrzTMOn
kstiOnyoQlu3ZRsn5i7iwLWlS/X6nT2/HTc3xHqsDynjNsE4d8LMO2V7UKprYzrv
4OqQ5vvMmBQ2oEAO9Hldg5wCCUC0epCXWu6utulN5cFxPElfVhbTpdtqXL3xTdRd
yvyJzy1Ss35xbX3lVAalI3TpaCPJwGbwYfvc8s1o8lQzBRuyq12xbHCqiwXsUfXX
3ugHkssVODl7jRbuKzAYrkiLjcsK3crbTa8tX4IY/q2k/EedDECdS+XEZtuKoQ7p
XVTwARsMRaM+UkKa3dg6GNo6qN682dUqAWZP8ZL3sJn5WrKlFJbH6n6AjkjWWd+S
rvyo7qjKmkhNkuIBJ9MNt6/pT+LvW4Hu3/QzSHkKrjf54olvukIxcJxVNvtghrpg
1oibcA9It93IXTtspH5v6MKSHBZBQltCiYiVaiC/sA7kn8E2kR6NPYb9ietoSEbm
jWuoim6cD+iBTjh3uWlm1derul7kKS9npYHwBTvI3mapE/yHWNeATaVzZyU2YUpH
bVF6JgqqRy7Q1Q1PDbjdrRiOCAu3grhZwibrRCY5DxZmR+vC98ssDFAqZrEFRvxn
fj+s+TQX2tC54VIrKtfbhkPD5W/0r1FM/vVeVklFRPDViWnupLC6Y0YmtON+imZN
aJECcLZgXb08Xot8S3zBnV2aCWviQXKrl3bOPyXkTTqQDbD0n4AtmhCHgNLK2/TR
qu+1XhuCm+QeRR7MEylHfIw8hTrS14PPi8Lu+yemAbmKzvsyNQ+4y9f/dIDhX5qf
f9WXKcxn62uVLyh1geiIDjZeWYA+BQb+iAf9WDHGdGsFDrCHQi2iLDheQEwClLAO
l2VxApSicIZqEHyC67VFOBYEPosq1LHQFpynXVCiFN/BZwPg+NBIKhR5QAReVRpJ
hk/66EMC8sBPR2I6OC1ncPMmlbvwk2EHYXfRhaNC+etPI17sBF+Q8J3Qup9BZcUI
Lh6wWVl5qhkOGAn7lDIU4OAd+0GW3Q2gobYNrgDgGcvd+UVP8Ty964DeLJ8v3Xa9
qmDU2ElZXN0p/vJKmQCVhwlM05BPkVQcTXvqiCy6ASZ8QzJLu2Jhlf/LKoplDArj
vO3sUI6k01S6mp14++3o4KNomqadbU9aY2V1rx+N3ipYC4HugQQY7JquM2dDjRW7
RX0QHKIzgwcOr62YlIwNCU6MSv5pQKyCh+qSloI+Wd+XcQq4acFf7Cgu71O1/Qb+
FU0k07IU/xomjr7sF8Yr+9CwrMM8I6JtA0K+ildZ7BkgT2zQSurD44b9ntgan8xJ
YzBpBZXv82zVAlY7KzN4xhuEGLeU+HUN5nglHFGYUQCNdhRQh7id2S9eYAsdeRlO
Dvq+aT7/7AS1PBAz1vvI39cln2FSq2dIoB7xOiWLZZpBrrYYEU8wIrbgYrGNzKdT
0FEfwzis9D8CuEV1FO6NZjYnm5QOyQErCZGITZxlBDQ2y6eeBXGgP7Wquxn6Ksve
G/Hfhsmo4XWD7Fgfz0rqcNcyCVYvbxTwmLONecv8NPgTHNE0QWJ9w1h9MU8GYnP+
w14IIqh4uYwrtGLjj9y8M9sC3k8wG5jlOQD7wsilffUF8mPyHxoH+GfZLgJzQ5tv
wjaA7wBc2eZs3kmZIQw4eNk+AxKlhroKTB0Nd7Qv7IMWkobkfc7baCyFptMaWQAR
g1pr2wmAY8x2bBcw7wIlT+eiiAHP4aIFU7vYd0M7nGROCZlCKAQsZ3CnXI7STgEu
XHOkohBoZwAkm9JfPrl7C1kuRLTDKvwToCg+JXROLLWWlZWQCtkJkH5GQr7+jeEk
K5q/2f6589Aoo8IbnJt5aU1OqAiQkckG7gkLXwkmBGlxldruMOr134kaHsvxGOwf
/m46qf07tOIOmciBFvDUFa5wEgMlSe+V0zyGuz0p3x7Qpcbuj2d7Y2+y5Z3a5NWk
vIHNidIlEgOYkqnU5XqrqrH22+W469gsOKlAuQXS9+rCoRwrMknO/a9WCQoS11z+
ryhfxIC67+jARJ44KPHQaS3ZI786pgOXgCEoCkgceAeIELzQH0F0+awA2eBgZG44
xDhjAYGuzeqdSRFlyZuPpfoJtywvRTh2vD32XKQ4dY+DNfhpD6Vq3c57wumWlyGL
ctfNICvXLCZJxPzyPcdfP02uKsNtKmu0ZpLzv7v4D7B8ymTv3P2YIw0UCo8QPMzZ
4in4r4vDxxGH4tcMsu7FS3qg8LBfcmgQ8ULIBNrWKJRfWnsjFPBkrx8s/TwciT6g
t8c7xMzMJCwADK1Fbr68Mz1TZT0JlMvEVcMrkswQu6dvhkVY8D2TZK9NXfwgIg8Q
XCWJAnHjAGiziSypDnYNNNCqSU+sneyknyh3Ll1LycqA894wPwhg2uiIa7RG+s9W
Ia62rLTKeRbupzykKhTcQXzHQkQY3j+IE0Fmv3GM4Ze61fSoWkZOMcp225Wdwxqg
n+mtxIWgXnHh3qmyXO0AI/WMfp4K71JV8GNewFB5NH2mOXGCz+3EfCcSLmqlDhcA
27t6i0Nm8j4DS/PFxfK8xe9JHcSOywe2QS3VhKLnzk9zzOjjEW/aNnnE/5ov8s9w
OMFkHUyDiYZ0C+MwNtdttBJqd9mtuORcJfoP7DE32fjziq48r39rwYpalDccz8s3
2GYZD2ifZKtt9JRS4puFvBI1WVmCX0vMATID7ObpbsShScRETrYfr9+Sx71km5e9
rjrgfugn8J79qaOXj0e6YStj8Zafl2+uioH6aP5x5pffe/aECHH9TlNO9U3FY3Z5
xPSlF7CDPXLvQpkzoVkfHdbb6FhBzdKAX1XNbSaHW7TSftAHesY5/GJDNi5U92LF
BZiSDADgSniXgoKpxeWLKqN93yEkSbEGY8z0lIfw+D4Eq+hs9ST9iMzIHfkNWA1Z
N+C20acdk3+pYztujfn6gWiZlqWkPzdvn6O9HzdSILTNygFIcaUO954gIFbdEloY
E6oEr23WVfiGxKAYOcmQbOABtirHBKcEOF6VvheTJ0abjJ7jtuFhYezps6bMVy1K
hO1s9Z7C+V6co/gGFAsqoF9IvuwMHQqiYmOZ8YVcoz4aQILauJ80mOj5flZPtgmU
oUF/9Ycq1t+tj+Gc4v5KakW7sjKbt8Ao1tp7N5xe+U3aP6ePOo++f59q8EKm6JuW
eGLdjsbyR7arhyDucHo2Y0qPbfWQgMicNeOc0b6HgN3VpnPni7FTmrGj0ox9znTf
pKrNtd9dtipX1ikblBvX1YHodCwzsBP6vzVDWGdo5JG7H1BuLE4aNsv2ZmqsDicw
Ref6Jp7nNYhaw/iNPU1dAFb0fgjbQpUCqEdH/TFx6xQe2UPPZYQdpA/f2orNCONj
T5kzcVq1gi77OJcv6U5zv7no5A56WR87Iu/U5ZUqxbZyKbkNEJ/D+IStj23d5Yrt
jIyAUw7Ci3dmPYvZbcKJytQNmXGC5I1dDTwK8VU/6lwKrG7+aZofECahQOsbL4XY
Skp3CWC3whGarwT3WCh/QWxE1tvvTVG+ilpK7o7T0zC0SIBNDRFB8QF1icg2pIu0
MuikzeWBWTeAIVAqTdARKzHD+K3Ux2ErrAYj6m17emqUHVx433HzQTXs/KB8zshY
YjjP+wq38ywVGrSphzPrrmglOhvwhWkfX1/gxy7drjUeXSjm39EjOF8rfsgvau8w
aSO+geny0QLC088qvFWlw8i2tVBxLDVExJ/1cHDV392OrHweBAKwnTdGhFby4kkx
+ygOVdTACVa31I20kVFb/wXhMj9rci1aEj2y5kcRc0kKlVKg3uWl/lCdNfLJdYsR
fec932UeniowzOK6I44OJdRZIMhB9judxybX2y/90wDps2G0zfRo/Fph+zRfowXc
1Ggy1jaqoU4Ij86NfWFKEviqEYs2hdcUnSXzf/cQ/gulcifJhjqGc0Ud0FsMaCV6
YSaAvj5gSKxBpfeYw8YaWnCdbc4VpzjtUYnhTWgxmz225c0CiktS7psdhfgG+tgA
uoPyHXnNpjd7LdIdAwELx/K+06IzHhoY3aUYjQRgE2KM+hiXt17FFwNM3bdRy/Qf
N0KRgUAHN80DMd5NBAe/87NqhM8ELaLMq+9gXhCm+LRiQB3SfgYJDOSWGvtW6OgU
npju7V6wZSSFNcayfaNYxSs+uan1S2MJA7QSeaxHG5r5onG3mu7uOqnEhPBO0oLD
ZeakTVKROlOiV3pf+nBJ5aJnwUnBlqCpmxAQkbzH+c8QBr95NgVJ0ilOQe8B+zk0
82t2oIef5rT7GW+XHCkLqG5AUTOkiNKxa9FMTguX0AFTj0gIPaNEBEz7/ltXFRhM
T3OnhSc17kkpSPTYl2x8obgAbb0mL8YEgGqntNr8lSEsvJWofU3DHjJ8ErXA7P3g
+AQiZDmn9RvhD4Ohd+7WGb3ZINLzRRK0dq1HsYcdc9JbENvuymvjGkaKhT3c0QwC
3XrU6LAuURgwTUKrPiD+VNY969QM+CKfjn0qlCmCxgym9t+j8tg+ZcP3MifXK88y
FAt6vjk34W70odSxJosk+UNrztvqXXvk6lhGm9knmPT/c7eixNNTi1J8D2XyYG+T
/4Y611juhuJ5e5wI5JXAZ2JFz/3uxRxQdkOF+RJUMTVmuUfqFpj/6BtXY1IBu1tO
tzHaAkIccUHiUCnYz2FkhIMclg5X++7fue+e7PYbZvhWQqywa+RUjny45SlDkDxu
g8KOpicv/ycPtqn35ikxNOkl2YhDz6pv4VBxZX9irlp7FV10gYnDXuUetxmw56YE
LDln0M4eTIRxrsn/ertxcI1kFVBSTt8/uPj2zMZh5u0LDQamw8N2E3I1a/KUm/XB
BiAagDPyHltCRU2GN8LN7ojPvOEndg/LPc2JTt3ezrPn+8AUaBHAPPZfigpyJbcN
TZDmX49QIqzslG/On+Z9bNISyogyldactZit0ueIWmUQPM+43MK6zoXzPedoMwjH
iEFTD89zEy+jBJ7rzDAL6w0IdlNE4jcqOKKWvxGKup6YKVnZQ4JVEgCCemaInLKW
fo+mLRe+lnvl+dBOtoUVeS+Y/xFHqd9xQxp13SI7h9DAPm8pBRKy1zQbN5tFU4EO
UoeQhG8wyzC+JQ6x+g5BZy6ES2cxQdJAne2aTjyd9k/Sli+2GQqwCgIMykaAthBT
e+ZrIxONnqU7pWlGYM1G+DyilQwBW3zioQmksuM8k4hcBkipBT5yNd/xSaEynq7V
JNgXyMLoE7WggkDrpnSv3mG+ZyaGAkfQqPfhlKof112dhHB+wHX3NG/dm9y1fFSY
mJLC248qtbNBE8q5Oc1VXzSh5EWYoyVYe5myGMDHldxYlIfBbxBFJhEVHMuGtaWF
fFTFikCO+oYMSStooIAhr4WzgsLIzVnMEO5KcQYYsrfJOItXqZvXu5cIXfdO4Ibw
sF22GHF0X0wnTrnrQove5Wp1F3yVoHx2M6KUBFUSHo5C6UxYuUkt2iU3yxFTN+SR
PMqijVlxk1G+DXqTMIOOo6rH48bK1XPeSfJEYtAco1kLrqzlaXu309qN3gu+Hl7N
YXgBD2fc8+fS3oAfQG04EGdNWAZAH4kKXdcKiQskiHQNNZKfk3XMKMUsFK1pa5px
EE9413Ayh38dCvTqF+D/9D8BEYgcoxUZud8XPo/EUViR1PxTTFwfD4iim6/9VaIe
Dkc60n/RLhC7pDwBL6CCBqr1LwcrFO8uzk6+rrIN8kj/tn+FPdU8CdTZCvYnBqUC
gWvNXd0EU6DfnjQFh8MSvoAdk7ZRsdJ1bv1GmfRf4Kf8Igl11gsDRgKEnMs6uEQq
/P/AxrDgFdnMOd/yfmCjxlUIaSqYElOP7ycn55TgeAbFYQDYPRDiuU6ccVoUDw0K
uHd6qvsnqw2RKYNUPUJT+dADgAoyUMueH1ZWzPzapNOVTpcMXquAwisvlSICwNNZ
nnWqxz3wHP31jvvqmOXVm+DhalMJcyOCyFfwY3f5xR1v09L8wIqIY2YjNq8PNETh
x0GNGiQ1pXa+bnrzvKDsrpG1XfjH1EgS4o7Rd5c+HgMSljWPk0Mo9puQ7kdrxJCz
WHUgf2YGdyc6w9Gy88pP8YOqYXGoN+vMTBZ6AxAmIk7mnbY52DtNGLWswHHrHbC2
M7E36b1gA+Ov9OkJD6jACL4+u+3vYp2fUho/saJ36GHSJfmvW6FY13WC02DdeWtF
PnrzWefLbyEAsk49Nkoud+Pfl2HjvWTaYRhIVhNCppZtuinFV8uiZ3771OOcY4sc
W86/fYLDDiNdU3yZum5kJk6XnDqpJb4mx8LBlI1P5E7i0Sa77DpNFPR3XeQBeWyp
Dc86xnV3pjninas8HmkOkPAr5g3CweIP5PxJvUCTGpsCwp5gq0pzVNgEWhmqi03M
vdvK4GwSKmDQW3MImikvY4EWdsNDcbxT7rApOBnQkiqkJ5DtOBGcg2jZ4oUgXQVd
QEi2y5M13jLpR0qs50s9XRaBqgdnLTqKbqwX4eu80hc5hEQoxc4nzWoHJFJcJ+wJ
iWysoONMv+O64oQnyq3shxlLzRaDB42QhGnNCP78v+/1+pMU8AhyO3Rf23T4Ennm
F0/jFiYnrpFjwvr0m2QHcU+mvIuW4UACiHp/T3itGBR7pak3NF+61b1cAAkDywk+
1wCWWLJPAXO25QTzyJyPKWxgGYOq+pc4IrpSNhESi329mYjjRtJ5l/+q/3OfXRyS
MOptxG2DuLTo1CFVq0VZ1007hxWS1yifdCNdwWbLZd0GmuVk2ANRw84R8dAHxXbb
sJGU6nDymMunpbTPGH13x4sSiGsz3ea6D0EsNnGhMcdw82ho8bfIs1smYPZR4KXU
uqsOesnZjp+BRrzxtEc0B8hGRqIU4fA32BhwZi+iFOGkEAvXqOrkEuWTnkaIQWPj
MV40v8C2oMsxqafGQSpmBZbH6uniEWGQGJVeG+aUf9LUKkBHPtVRRRd3ciwt0bbB
BDwTtFVZaHMzULd8nJ3y9sf6p+xY+qqLGaLYsN3xy4/QfrCDwlVKtGzVn+5coO8f
p4Xsa64CWNoHOBWkN4+MEJ0rw3MCxPVVpW6KOOjpox1UxWbDt1P9viBI6TnXSQ3+
3EWeNGLF6R24T3mGDwR5V+BRchnLAGC0IzphQMyPSYyd8aCZXypMh252PgChUPS2
BgazevctI1H4qwGRcKzpurZp2Ink9N9Wub+5D1e3GswU07Yl2OOgGFgqJGInU2GI
4EeHlkUmJw2wKiyJkNrylLpo9B2Td/pVlK9T6c0Jga/qsXmWhk+dKh5P+QPXQUca
a1at/IQ9yMriExGM7yGk8LwOjQdQokown7j450B1TMTEhd6cY7KYmSZQ4pAeLCQm
0CdOoXqXmJsM9oQPhBxT6rMhEYGezf7NEF2Nd2OzJWqW45ONEVUPaIajgVqYk8Ew
ue7E529ocJnII3IN/HeVYGxTzAQPHPa8YEV7M9Dz2R3VjUKp7heHsSIdg17shAYL
T6ZSv6Ru3W79SSdLssi+2nIaAXBfsRa4XPUL6XaKb+rYBddDZgGBYjz/tIA//K+i
xXKvdoqriP4H/zxZEU0NXgNDs/b88Q+rsxO0UU2U7/nN98ymyLMX3bdtvjtamG3r
pl2bsS0wT77KZTEad6z9MrZxji+5fqj+c2ZwcIwEyTgz0SkefbnV/rzDhIh+cafj
VlHLKna0BjEkGdvmxZ0ajCWRqR2rtf+bmI4mTDYyaNwO3ZkkF+0X2uJu4sz4t947
BwNbcaohzviW8EprSUailnOmhhVPZ2v1rDCB1e2lIsUUShU6As2GmsZHdzKjCPKx
bB1mPvGaidRVPfW5PXDwEEeJGE3sjedzbptePVftm7j2Ir/Wq4XTcSJVlbV+UDnW
wIYIZ5Co0DBVmMi4aBVLoMVFa6tnBco9DVgRRPlC6CaZAL7RrvO9qK5ZpdsmWlAw
kUaODcCMfAjYvhjYHHLpWQUKIlSO+BUMhEgi/WqjxvOZ3eEMgWaj4Ya8KC6wlwoU
hqRoG1nYRWKzZUPPegGmpj9tw51YQ6/Pu/9REUDCVbuhlwKtQrqvAKi5QjvNXvaF
FHWMtkINQF2vMHj1eJvb2DsO4tLAipfUe6QPcPbX6+cQ9Jr1K/bypM2yv+9nTRQM
pG225qt3iC0CJBWa5tA7JZ5E2MtAWyS/RF8pVifV2pCP7zM92iRkzn5JoKwN3Srn
zXZs3FAtpkSSViS7qmS7+72kbeEQx6fJDf6RR5Y5D+3hlHyq2N6vaOLSwkcR2dXN
SxHMqNGwQU33aHWnEU9/FiX84Vq5ZZlRAbRd5+g1WeOf6VyQ1ITXzHw1ImvC52km
JkfeDIm/gTkwoEX364lzZsFfv58UibbizXjARhLjGLpsb37ZzCE32i55vANY5gth
drNXtE4wkBURTb00lX66KYBGlfXNO0lrRCE/oBLqHmbsDgCFzmFYTm446wKzTkm/
RQ8iUM5lZlNaXBuMnWgOXqtWfk6Uc8gJcnYSYLAowCax0RWnjpxC1M1LoVZYP0fX
B52NrB54qaynd2GqoL0BbF6Mi6rrzejb/34xB9bRfOb728dKH9LLU3Uzg1yXB7cl
kyNBAsKnitpPpye0ZCI16t+ac7OoS4PczAelctErJyXCflxu0WIsYQVuABsmiCoW
cMACnu7sdT3+1yW00hKxCeiFDVjGkbYtSnln45+xGrH71JheNRKd6Jv1tiN+HfRM
T5OQp/KP1mDaRUCT56NFN2WpBtISHL1idFTD65XbUM/iWP3v9GsSyYgS5D/6LJSx
g0igU5ER7LMXHt88t1LnYqwELG5YGdL1YiFllEY6ZO5qBkCb26q1NCf1oskvjHWK
/K/cWWN44SIRREb9iOpBvJuXAPRQBjjcBMKAc7ihS7ykIRUCl2GhwEDEYTa9mY5R
Ywdx4jgkkH8M/Fuii+qdjwkt5s1YMq/ASKv1tLSBsJPkA+mp6szWXASmYBtCd8Hq
gzvLZ/nY+HF1KfAStvPApPsu4xlDePUV30gBMxElGfXGLRBYlG2/kjxGI/FumwuK
UERUB2kh5naWvsiJH7LoxEZFuO7rEzxSQTYqe+j6RBeCzg+l1vVExNwcYPXQHuAv
VPo1h+SQfdxoG/hkOOTFRMLv8ymijrxIx//oQNaMJQygt+kSlK1nxWbY8WAq1XfT
d5Z2CRr0jBQa0/X5lLThZdlagBQHB7NrgUchmHglRDsqAa+YEGKfEjEazh0XGpMl
ttiT6eYk9+vcaTQ/4U7mbaTQ5M6Ai2g0IYUclABH1GdUXT6wWVwvO9ms/X7QZ14m
Epya603u4RpknRWXfAXsSsC5ZdrEAAs6JBFaIp4jUJ62bgJR9Uz7yA1ZSqu/eqyP
NDjzmbSA1VeN+iGMzUAczyvTJ6sRTwwXTHyakrfSec+wJ0wUp83C4g4fIvY53qWr
3hn4JBTfxUaqgV4QQAKGIiMe/WdFugqnypFLTovWFZkSbJ5QtNtxNTdFYKnHxrYJ
lSqpEpnQmY/zV2ht/mML+k8kIDxp26+q1/n7Apvd2SeI4TQ3SPM/OSV0QN5D5T/8
Y3LLEff8oeolDnieESKsL74ruAyhHzjSkYvbpucltaq7oRIWTv7rnP2eXs5UbLlB
2tf2YBQpI4SF8iSLA8VDhlUShB9EELqxXNb3H7vlXVCTuLShveFrN9lToCe3rJwS
RvzIhUmMWIAoedjXmZ94frLxAB5jYSolusjSRgEFsGzQefaeRnWDQUP32IgPEQXm
Ivo0sGym8UtaC5C9OkmFRnkoc2P0nqfivamQfEVLEOGqNLCqgtM0md2os78cBsZL
5H+Fzt9/tpAHZhW4ZAdiqp0Mr7QkmPdhdNtS3qDnnxUvOYeofDCnqmMSMXvIXXkq
q1lH6Ggu/8oj4GhxbJVvUIcDDC1M+CqmZyojKLi4F6hAKlIxunh2g3LrujMUeah/
inPk0e56rKVIwwhmPPKt+Vta1BPf0mS/X1zw5Q37W/EuZho9EDCwCTbIlLe/4+Km
k1NyPGxFjE7S8TPYKlGRU1hXHgzD2fzydbNgchhpjVp/eaWSUWT13tgSYWQUeUQn
Zvez7Nn5npEuzSUFakDpECQedznU5qxQVeRY0kvlt2PpVgYtGuWA5G25qqUGyeJ9
fBi08Fj8QHW7V1gaPACC/eVr7hm1/qrfnkSPVOaTHaTw7hUjh8a414VFF2Ue839K
KVOQAj2nU4FfRbhbx+Z+DodtWJ0aHhCcz8S6i6IE82WqLG58ChVliJC2GZUZ3LTs
jqn3014ufxnqJmz+o33O3YfFxXWRbOhVIeOzeYLmOVlpcgNlO3A79zRVpXooe6aB
dXZ6W/au8gTHaj5Ow5s1j/rJtP8x6ktmFFQMdbaMVxL+buHh4COgCHjjDwiOpUcS
sam5cOH8lUrsu5VRsoa+qdBbdy5BtEYxSbEGMoSQoDKPXNO1U6bkHAzWzvBiAr44
yeqFVJGhwu9Gr+Sbyx7JQKvtqJefj4C4fMPhucQznfqEcSxL5f5xCWaNQFcyKKmg
A59IE/vV137Baw39dq48JBvlXRsznLdAfg0xdSMREjlCvhYEmaywiwJoQuHWyJWf
+wSfsdSEYQb9utCGbpEwOxUyJgJAsk2B+kgcQaqccnYpoNN7sBGGleAFamXABsl7
KwuIEFq4TcTA06HmYu233ke4Q2X9NvuSA5mR5pPwaAJpAMJerPeOuV9tKDsg0T18
tzra8o2x5IJgDpxsGsPbwtppFsHKXzHEddrcqHIGuHPPf/FsFYs59Zei9yKMgFYk
PxrYGGJTX5Om0QCOZiE5YaaQg6peks1UkjvUapvklUs6t9ST1GzEJwfS3zaZ4n+Y
pqqlEEiBBb3e76yqSDSOpAbgH65iz3J0ieg5guJLTxChwhs1SsS/kkCOSAvCHokh
jIQghul+wWag+/5CS2Gpg8bFMaBY2PmW5CCUapohAZtaGz5OXy01q2h5lQOGcVgV
BNiI4s1jYFK1+XfjLXEcdxc0E3CWT6ShaHTjWpDicMb0OqwEc3mr7TjztTS/JzSO
KvFgQ96aSYmlkz8th/g20cqtblJMuQW2mFnCtw+p/rpI407xCJMQjmzzVVf02ebR
O9O4uTzaM3Mbgdn7EIPN3XW83JdAQt1cvb2hmRQTvdhZ5AYqUhvsr+Br1mw9CBXR
1F1CJp09nXq+jgR80wkcm34Ni7Y3U1empCsgu4SB6IQqAMocGFr121zKYGXe94JA
Gc/ydMpTgQNHPcTIRMjRa9zmhP1+p4YMpyKUC1Zt6LzFa1tAM9bgISFTT1hgBZIn
W62LgCLJrufC/DcAq7dvWlGoB5Po3YGSBs7/um92Nhf/U/1xPraAYof4nCxO4wek
knMNnAivC6FARItjHLTMCoRfvZhxIgULP1BhMuBdYKo2ZgiFb0/PYulPMOO4s2QV
H6E43jW6pU8u5ZWtCGnp1I2U1OJe58xhiChIXhFk3zsXQE3Yge036laBtAX4J52v
IW3BjhK/JAE9TsbxHlE0DWhci9nLJR/2zGTTuV6dHZmicbGwty29jAspoElyq5/8
z603WOMAwT4yjsYZVO+oFdNV4HG07zmu4f1OYqq8WmYDKYA8IWQ4W/oqPElHMnUJ
lqJk6GTLIFipS//t6Z4symrEtKwlyIlWaN+v3/jygurvIUxvF+eUs4HaCLyYwOIf
yOpRLJCWR1bFCI+N1GkDIGwNWbfEPhJ5E/jcoZNMlFX57vOkhWIvti2y1Z0hnaeG
V30ZMfcwPyKQ9wIThdYD3eWk8RjJ9IkTZsnI9uSA94phNxPegjMCIHWIIfLjTUKT
ZKhwJe3oayAzhvA9BTNt7MKELbpO2Hpy+igZjBb/G7KtQg+Fm6Y+Zd/X9v1fa+iH
J1l/7dELj6VRdjibC44wx5QOFcrM8P0Zsm2dQjltXehOPbaPxP/gieeMhD0s1bSL
3QRNUKMKV8aReh3+Kqw0PKSUVkk26AHa10ESeWiUrCW4JP50i28w5iBg3EFZA+7+
Pxi1c3tV6ciAdG/B2y9bcn1WzUJy3x/r3APzw7nqEN/0mDupfD01SLg5UIXty9QS
anEIyZ8jAy8Stalm/A4+oTOZ8hPxIvybfkXmhfkzKJtusc8hf31F25BoBygMnPV/
QjjRnAe2YmtTB1cPPeRL92X0kdA+kmPe+IAUOotuLtIBmoBGfIbAW60JifsUXOuK
NPZsAbpe/EXBwLe+xBV9GXm6WLD7UoV5l6NCPRJYm3VC3D8Qh5hgzRWuXmMBl6Rb
qwjVx6DaaiM7X+3HPcYgTTHWb6dMPTV97g7Q9Y7Kwq3RQLDZt6Yznjt1JK08ytoy
t9B1T168YdAWhlDA64C/pLQf1Uyb1PlROOiizOA0oanlzGU9fxDxj/orTN6G3sgp
eQUBKJS4phG5UjLj7PkIPzbpL3RI2Ss+hitHrUyJaQ/FDQD2miAkZaVAM/mN67Ti
kYihR5xreGUMS1JADIyHS8FrOxHPC3/0fSbYwKNi+XBjBqu2etqfJU7ambqL081T
Q+4tKlQw7jfSH8hOPEcs/TxoLWvCrGF7FmY0IMYABRkps/j8tjNC4BIqPS365aN0
REpbQwX9x4J6E2Kt6Q+exeLfzP8qTpNDaiR7WpsS2ibkZNnrGeZP7CIty8Oc7s38
JVSi97I2xBpeN2RhfJugitbYz/OGOTIdUVlxegq3Jwv09s9jwDwd/hw3JwzOM1my
SnlmkEhWeOlKSVMUiTw9PVqy9UgqbZsT5UeUe9iLJC5zHy1W4pFWkN8sckxqCrkI
WoMt+FvM+HWEHdBGLUu4QA+bLNi4CnrLGqnSZy8F5Qr0cLzSoXxb/kNckzkU+Nmu
9RIEdwUBUgPGPBFLhxmirY8iQ47FZ5KGXL7UnWGfloF7ifP0yRFvsNva9ww3XxGj
enfPuCO4Y/W4uslAwl8tDQv8XSW3S/u8QHjZZmm6QwCQM/uVrqx+T876bn75pKHZ
FUC2S1Un6/DROKS0uNvPJOBwTn5NLbw18BFtU7SGgkiD9z97pe81ITx2x12gmCjY
K3CVIEYV514G0/2/WusA9+WD7w99WhfHDp1wfNnkmFWYzAu70DA5d6jgBHOkslW3
pf4ra8gKjCs7WqQzrLTwPt3t3qFgOcjVV4nMJnVEDI3P4d3Qt69IjJxTC4dFX/UA
45FWodDIg4Sjg6ScMSaunYScq53zGAlry3D6l7MtYQr9wvkWff2TeXWFQvrxO52U
XaSxpmecrR0JxGLT6bKf9hdvjQqZkj+JjuaVXlNBHuqWDh4de5TOLGXd26ICum6l
L47T37ZfUtSvOEOFezJydlloen3yd38Dlc1gV3i8702Zj9oX8c1G2GN+xXJ5Z3SJ
vsy7ZCfNLxfdfafFfTqPrvnjV/eBKrGUu7F+0zu+wa9wz4PJMw4uf6SSkUIxtGHc
1kPlZpeY3RtMWAvV4WwUPeDqtUoDzek5heR+Pt1AFR9a0K8cXJcpeqNkwF+cGndD
CWwz9sc1r/8Vf8S46d7f2F69hFQNoJU9UoIds6BuwZO8tXypRgtFgNoWts1o6D5T
AjisbEroYR3FmNIv5wi0x69QIMM3iaRd5P8NTmlBflQToBpYR9mTUj/K9+AqWqf+
FsUwwGBD2ZdLeLgCPsbwWYc7QvFKssDKLgVxI+2Xzd2YrFygJV7mhlyHSctUrx08
6luBfeiKu7FbSfatVSpUT1XReqLBSx0P87YszS09A4M4qVq91cHBq5D9X4EDdJOj
ivK9psh+21dOsdtpQNPkLKFXk54KkwLqe8m8kkQ1CiE7XxScXzG4MKX/3ZBdJkau
JMZbwyYxBSxeBmawdFw+EdlpdYDjjOZQh7oOZE/3FdPu3H3BviD3T4T4ayY6smBt
mEg5X7BnfPgzejqFeppwNVavpUdPwS1kS7j/KquS66WiXxTnmZEk3lREBdc4gt2Q
+S04Xq70H/MejQ2BR9gI/Y2doirOpbzLinVcxyIO91R1BK7fEnazdRBcBwo+ki83
uh8ZD6nTxASLY4RlV4P9nek8pQwhuj9damXdIr+cUcXRI6hxps8Bcj+9f06kVwDJ
FJiSWUyuPWDF3GICYWVWcu4o4eWYHAHNoNg7vjE/GvQ6ABWDoZXC3/06NdxgXHqi
s3mCR4EWIxzb6v8YTxmCD0gsb/SGUSudgwbIO7oNuFp/ZB18iPtXi479BhPqRdfR
0QD2GQISb3Y2MfstC9KGwWNYvLPCauAE1UyIvIYV2Wd+zJLInqRRF33rkSEouUtE
GwU6AInOw3dg1wM3KjdAM99PTFUu2Ciczuhgzz01/mSO6oAZ3Pb5zMcng2mfVLN0
mpBgvZv0GSO8EkCyIm+NlYno/mxOepOFLh/GXxL/MvR/DRP1ralCTGIJUfLt1r1o
s6OG9LXli5qKOdp4IFYfFe3Lku2W+LVVeQZee3iMScAyYI3rzbZzdCFbxigjr6/S
0/8gyLy558jesUFLlAQSS424PFCCJpLc9fw5BBPliFxbwWMN1jnIaFcNUOxcb4si
4oVK8m3wwWHH325ndQ9tkYgxeqgXFLiAr4rALV00DKt6KaPVZNAWln8HsRS4RYxx
qMWZf5MfKMdrnIaTVl+IWLEO3NQyEOYkoHcfmrpAydqy0syA8SL70AGHHL2JSZiu
o4Q5A/2Tw0Ta4CIuqOgaJHpDH6L5ZM6fZysoF1IkLQbDWAY8peUbRw96cXI8g/tq
Hvd0bx0AdJ60Is0j/8hR8Okw08Bs1Xe1BpJd12iO4z4TwpqZHIhHRdjvLHXteSkB
vjiyw4SYOrIvJONZYhzWA4brmDQOwYs5Mkyr6TJsTqYqGrfcwPiLVZYgaIc5Lw7Q
gcg8vjBv8ywXWLWIkBJP+1FEdTueo2otvkB/NQhvPsYC7oMQFLoQWrSLh1bna97z
CFt7PbMeLM1/23Aa/pWb0FUeM53kPuOz8vPdmNClccczC3mheh6JYtaYl7Pwy2XO
+h1oC5Eid2LXlc5oQIEauEd+yWTTV4UJjV9VbAjpDK49XENrW1IyisfEVYUGfedi
18TSv3DxMIMNJeO5MKLHT1y5p9owDfRAsrbjqFmtj/EKa4KpuUjov8YQfSOB3lxq
zExjCfrJFkGCoZvFfcn+snw+H9ney7geBKIcz/PmZAPq6/yP4ZUtew5I4YwDGEjh
gN5JC1UP4GXiDgF1JcKtZxt+PMAVKp3Uilgkg9514gnsADt1WQ0VZBeOXcGDjbYy
9Ihonw4rJ/5VK6ai+t8MKivnl5LZWJIOoDfSMpd+4yLoFHXvVIMQlLmNIQ5FnjHi
srKSuWuiyHWMih810pjYJY9lwEXaKtgbFG/auMcCJFsR6Gqi/i+X/S3Mc8M2icpt
2cJvw+apJDsScpVVxAE/p03yY1+J5O38gkuo5oieVyXUQm1VL/6J/qcAPsGMn1Yt
+8TUU8MG2fru9xW1TWmK2pTDt4ODId3JDeopVU5V48K6lCtKanSpsU9c99sRx/st
zxagjO6tP8xTQhu35Nop2oL8LU6UGIAyoyyXd8j6y6YeS2/lyX34o97mWgGvC4Ro
0BkvJ3rghfBvwGuQ1cdRGPgkY7wB2O8RP6G2EDo78pZutiwbLPna0uXdnY/bms72
ddpsg9FRSgRIawh5NY5Vhwt99f30Jl0aYY/EispuherENXi2JlQXorzFM+ngJmze
GgsSA1b+hfV7Op+0zwmdFOwOdtOq2cbrmO4mnGCGyLN3zKsVL0+Vhn30nE8gYi58
kbIQ8IlFJFVa5yhHn1KSre0l+9EbLKfUGTHZrsAmRVvlUzzcq9h3PWeV3fmiu6fK
2y09vCxiJE8/k12XDdnyhW3ZSLVRdpC00CccJY8UM51yoN8szZibqx2qx8CgCCcT
ysmKJofNPtd47ENLgIr5ZXcW0HYXnqh9S83BC8+8QgYIZxYClMSalWv0iSImyL5W
V2Kgwrw6ISsfEohOQEOEPS/vtNDYZwfc4TZsqJNPEUf6/gvZ5dRS9psD3iLbho/I
ACFeH+GKoq01I/TohdXNeTiJX2IgeqHb1YV04f3osozfS7q7L8YGKr0TTd5yjqvC
cB+tUzBL+n2n9kil5ZJPzj6blzF+khtw6nqeR4b13Sdl5saJVIIdx+xCBicuqVe3
BuvAhdHoXACk+bwaqRagrjK6h3lMejpCeMJvpScDvHB7z1WiimEPcenQitwLzs/p
TqTzdg/KP1siCTDBWhCJdJ+o/Ms9YScM2M/JkVN7uz8nJgUwQauUsZKm9mhvIMIh
jDPwM1s3VHf4mcDA2Pi2ABP8TSbsPLLt1ySOB7gCdeUQbuRCyH4a5wgaVITb1dzk
1xsNXV2rGyf99ZfKFESMarb/eZZPyCr7QzfoMoyMUp1GqhvNT8IAVKM7ChWA5oeU
krKpw018sA8FeYRqFX3bShdqF9IRbnEKEbhaDb5tQlHIe8P1xsUgnuz+gQPcMM44
7oVPL1d3fhY8ylR1lM5Pab6nqxv7K2o5bN6ABsVrsPoKbNWxKufwGhOEmQD7TSQu
bphADY8bcUDo9naudFz1USVhLz3wvmANATlheP4ow9HAz971YStK6Og06BEhK3Yq
oGfMHnHjoD2B0hwm+Dr+VIjhxmDzE9N7IvPkv7HobFhuPYpSlanlvj9BILgF2IIi
V0rq4I35+45tA3cfQvuUVOHVZ4hmesLWkfqoI1Lt1AYyYRdmCPqOs2gXR+jIDqUS
MzguapwOl9ECyqaA/K5axW7YBL5O7edrBYrwV5f1l8KpvtqxeBNVpMekw7F2k2lX
R496KAeXHoZAxEDwSGKK9ruFka8JCSZRcXzN3/doX/poW2XWFtpd3vEN71V70FWm
kp+8P6zXTciKVoTHHw5NswFyH5kqQmvCpr9rUjslAUvcIsFntDuXApWGPdxZrdo/
Lf6284FMoQLVtM14WPzSDSu7n4WVAmm2QLppHUfB+UeEFMp07aU81KfbEQFdBdvf
cyM8kBdAnWTSJFe7BBFqtTYiakEEaza7xB9rkFLOuBLrND8mgyTi4HmvWZ9K2bsD
xtcw6F5MRKcTyoXoDzYLDeb3/wHJ2ATZEMIWcnLpXUCnk+zy4byOtDZItWQBzSZ/
9FLpMyxTgzmez+Y0Zz78qBntKPM/GqAxxMNIT8iekeU52lFi6V0hjN0mthj6YR+S
uAtSA2wzbaDzh7entI9VuzGBvockgCuXePpRIVCzd2bmbbHRAkrcNc76IBfoo7CJ
jIcaJKez3UJ5sMJBuLUsIEv5gOaFJfvbOfRqdV9hQwDS5Q8adE0+qFWGIO+07NGC
BeJsOuumpHLM0Mg6A+RbBXMOOEdn+h5E4EYl8nR3fFzDBjs3KO4oVT9LS1WvdnGM
GiwV4/aynH0v4AM3Ms2WKkCLZRLB1qRY7pdusiKCbSZroaAgUb5nZgHN8PQ9i9pT
XwEF7gKogKmaiazV1k1Oa0wb0ynIfTLP6M9dXtWY7aeKqF+4EWRe0GBpBQMcWKUn
XmgKFTJXJyElB5K5a7l/4ZINbfwleutTecEaaMSW9ooXdu9pQaBQC+ovO/EpfAUX
nGTYL963ZHf0/yjefP73G4YqEfK8f7lz613EL0VGKfTU9SrVvsGjOFBf20F5VFYs
MCSW4p5mlteQjKfBRbJSXyJ6iS0aLZaGxQ+Va4wKVY8/H82ZbhtfBAQYIMu2mETs
ikFBI5bzF44k9wuB1d/1dR40KMBzPvspVq3dlPJ9T+UqN7ab6MhWLYXhCubmQa2t
XSuqmL0PK/LGkzjHbLyf6k1xjrime1etumgrci7QmALLZziXpr5skoDvlRB/BjVK
Do/n5zYSg2yb1BjLeLBw2Bk7YkNddZuYNiuxC1aqv2MAsA8Ex+IE5e/yW4ATm9pR
XG38ovK2cRcFsphTaTBbDQ2Xze2qmSkkLFs/Ik5YvBn34K9uWcLkcP4hGXu9t5Fg
3FKTsFIccf+aiZbecmlPVGxP8zRUDng/hK4+tL6BCtn0+v7+BuXv+DfDA6dOFydS
WA5yFjuhv8W0a5A3DdsV0KHh90uzmOTrllmFx8DJc6UYOFuG8YXkYdMK9CqzYQQn
dDWir4c4ClLxORxB6/KgcWx1DALm7ARKp/aIt1soVLFUI2Kzgl0X8uVXsOBDlgP6
Q9Lt8MFrHyg5Qcl1TdFMNf3snfxJFcMQ8g3k5niWRy1u2IhLvgMV+mNhhhswiK4T
vuo6JEvVD/llKyFT+IxJi8G0vQM8z+aEtEdIJtIVTZNmrlTXyNEiVEpoD9lDpMVF
YtyctXkrnbXEr+ZWHj+o5v7l+Y2yb+dnx3TfSdSYDmBrYtu7TTvbhFmq7HYNvsiO
f2s4jiyUnOBXFdv6qJu2AYdOlOyCrxP0mBQsM+szWqF2983sckI/dCZV2Od+qFMK
KJaI+1IAlfXRGBHgRDIMEVb2kv4jCTkeJYAXJhfbL2s+jW4x6QBTym6Rs8q/VtD5
OW4PQWNDB8gTcj13k2jIz6v1fJnMG3bnNP0GEPhqJOHBz5gWsr3sov+kqfVlLkKJ
G1GTV4/H8lpdwh1pzw3ulz+OOBUyunns4mcOBixhdfHpXe4U8xV26tqHulwQBPxn
BbT54HSJ3RvCr3xo9Rx46AtHCcO81ibdnm5As31rHZXFgQDYWS8aVxYvMwoiY4km
wWeeH2mBQMg3znxjHO73TquPOCJBYmRzic+E0+PnDb31wfNVXPmxMnZCtgKqel9/
aCMJTMhgl4oMTPEc5rynfXKA1ifG44aiMIPXwV/XZpY7Ydmty5EvaK1lawF7g1NG
t/d6ITaTTDSwMTocShSMxma5eocQB1tXXJaRyjyJwq2SA6JXeIlBtN/As5rDU5yR
6Gx1mteDubEhO7weBjke7fnLEl9Li2LIGV5R3Ua5uZXL9cHeHRSWkwKw0WdBA3su
LqLDQ8tFjudMr83lp0hqFEr6ZRD9x8lH5/dnMH641T+qNOMtBqWjMpB+U7pUx/Bg
7nhoK4zKfC3cPbOVov88K+y/E16U495u9jQssjwi0X3zDBmbicR5FRwrezouUqrh
9+XJ6LyPlJGGT+FxiXvNg4i2AeniyEXP68vxDpvoLjhp7bjFz8RjMx44R69S4MUF
rcfttmfOZ43HNfe+7rgttp+Vv5v0qhEVvLCa9cceEBdxQLYqUMbKiowSnikNDp7A
ZhaMfwPg9QowMi3Q0ltFo3/xqCysJWVKKi88ATJYG+s9qLZF8bVZxYgX+GG+oRBg
tTxPu4IxyQNVw748G8997Mr4eHElWbnRLKN8LBoHn6++f3yov3oQNNoeU6edW5ZN
MjcEPUXlR58JM9ysu9NLF4JJKx6edMkEOoGn+RveeYY1VIaE1NBy1wFQIUkjjZxW
klAMhoV/7CjbcfwfUs0CT9BwgHVXSxy9CYNatgsN0f2XWMqksAOO+B3bMH+Le4D2
/Nqq4elebNSVKtuuvK+B55gN1micyU45R+jMqmLsJf+it2Wf0rAHXrwMTBdtsJdj
OVh5a3eU/txjPgqrSERu6R3GZIqY3DlM3PZO7a5p1X2YiVfn7PjBfZu3SF91FPdm
Oaro32oQkHTJdsPP6gcpdJLjYP3r2uOx38IlnfSiytJgb6lfbDpUN5955QIoVBiz
tB7e6FA19FMC1/HWw18Dx7gHomlFSQzbmAuhlZUa968tbZqfCiMYjEEDR93rWS1i
ipwm0JZqeyqHuYcwp976V/sRlvkX5Mg7JuKjBLiBR2d1hdxHmApfQX/TfwNeERhc
m+BY9eG/XHWsnt8KzuEYhWXhPBwHnUbAqhwNlbpHOPzfrinBPyVqrdnGJk3rKNc4
y8ALcTXYgsxlf8gRJIH6IsEhR3GA3Jbj9WV29WeamowDV9W6Bc6n7AHT0fVBjDfJ
UirtyM9Yj5dMh93mmArMsm6QyQUtheQLOmqFacNGVekjLKXcHCgEbiMBY7yYYoa4
VCsBOSCcYcO75cpeQJnBKOcf9Aft92m71Phy/DEO6EH0Aaxy5WdrafdYGaaIabQS
l1oI+NmJ0fddFjgk3yP23KZfKQMwNrrMSL6zrsCdQQzyCRZBX88211WjdTt5oGDg
OGMkx5C55biAsVg0jOD84InDPDdJLBNsatW/WnCDfBcrc9YApHBdtya+dOqS5ByS
jdHvep6HiFJFX9KnSlYZxpwhiHxu09e82APNpq2i3v1m+Fjgrb9V+cx2gQPPFgOv
3mX1jC3ndwL4zMKfx5abtq8bZEC8g1cEKv2C0gTX8F4Z0Wvc2ogVlnDFwcM9huy4
ecLew9r7ddoEKd760gDzaeXbwiTT1hEJmukcIFsfnvDhZlvUzfFbJsQAIctNRZrz
qfT9BTtAyomQ4xNCZh5zdYSxQXgZWRsCR7TBEgWmdvWICfJsHgf6MDHlV1YzFM/w
Yd4mQNkXl3bz2ZmmKizQQ5reARYZCkhv2aEEm+P1AWRDE3iVxPwzn3su0cvs+POh
xH2X7g8gKDY9XUdjiLFfUzqWvu3PDDvXKDm+OSWTr10zTA7kTy6UbarSHtjXSRMc
nhXfIBpZis20GqFZ/ArXsRslPbNVGKj1jQkUv4QY1tDuNgnFnYxw0IwdmYvbGCio
AVKzVNs8KRcRyokQcWpJQw7WfSrzWlEhOq6J3eQ3i/bf+oJcKSaA1gNdpsCu5WfJ
Ezj/CJJ7E11TQxwY2mpfTKF4kpe98P9x6hNiw/qD5ZLwIbdt4cnniEVmxpy2WIlp
VE24HtlGH8bSldS4tKwS2bbR60WcYWgTle1YPBv/bQOhE797clutCCc6uuwXRZ8y
Nb9ROetbt905WLI2PVIf3KzthmqtAZPfX8aLMqPdp+i2vVlJFkEmTgr/g3BHGNI0
uLbSTg61YNNtMolkfjSkFlFPjimX8R4p+bQf1ttgt/ReatXQGyV9ekruwQJVxen+
GOjLUGIObDkg+HwDt6yOcj+g8SRCiwf3y2yQ8Su0VmVu9dfCzWt8u71fB9qtPLeN
5b67tG6a6RTU2KHaBGQQ8BInMfQq9VjkTpDTPqo1fkIBrtqf2Wotp2Aykh01jEsZ
cxot0/1aeKsn8Y9jfiyZrWe9Hku9mJFWHW5MyYLF9ZlfM7I5Q0h7RPsObx9nwQ43
f8BAf6EHrlHFSnE1fu5axmKir1dYRP/HtfmeUwhws8CHZ9UVQM2jlsebnfNLvdyn
giugqEptZbatbU0J5mForntwPrHFMq5YVcB1ojO1fwY1T2JhHeOVtgHluE2nEVHk
J0kTdJqP+2O2ov9+KHUBmhjm5ISjZ24g5+BIsm/ngx+E6TKlm5+KoZsSvT6wjYtj
0VZvZ8ieZACd9uYQs4DrqqtFc8lJg+yfb4X7Fc12BTVUySwjvLQJPdNtHvFxu97f
vXUYVqXhrV8HyNyZCTOiGI+LoXgdYfoCKF44Awya2l5teI9t0pfeanPaPCKnao2I
n43KFr1srmeMp9kaNngUaL5hPxKmWP6Xzpcl0Mn4VqI5zhHNBre5XPmOKidLGen3
wrXWZ4E3MDOx1kuGBBCv2FAg2gFWlGXvBDHNDXeLXZ0DTL7iVZanBY+8pbQMQTM9
trZPXG0CzivNtEDIj3ZlJ04KWv7QL46G5XNFvtrI5+q7yllocrTHR1lMLm32aYcz
gIzhO/dWq+N0p6nxRdwWP5GPw8fyeImws8e+2tBGJHznl8o266doG9reoBcc1jX0
vqhiz3yfdD0a5aoNRJ8KYQ45fGNqe7EaTE/sQqloOO7SOdnxDPKs78Nvy35+SJGJ
ffyrm1K62wT8WaxyP8EGfKiiv8MMctsZT3qBbmh7kBrlGjEE5R0URMlwSnO7bORj
pz/kvs4umqQ2/vw/38FH7Ny6mpFR74mXWiyIE5WR+Jbk9CzsYG7BTdFE1NkP/clA
eDgi3jZ325TokBnb4mHCq4wcxSBrFPzkXvPh+4wfj9DiiOs5bVKh3jzxmWUHJaT6
q1DiiniDjMyEtUSBpCmcOzSwhYM3+H9Qh5VFRSO/L2B8dzGsv9nOFjhOVrQqsswk
hhmnBNtT+k07hfA5diJBHEhxHqBK8due6MsF2xKei9JSdzaugiXK0PIdWnibL2HS
x8i+ieVHtEotTNOWzWaEL3IQrlAfT/GNrMNZneKjj1yh2TwkDXHmXLZPmLquhwib
pREXa9Jbx+/euuf/NDqMi/jE3lZ1XO7N7ztA2gR2juQr5hYurvRAX/fe87ZRxl8y
dJ/KPYY1a4xFNHWpUi6ckbhwBB95Z7UJ6iwlFsDR0R04k3nXw+eOO0hX1bcgFswF
krQDAP5RmoyAq1MVAOjC0fFxcEZl2jyjAAlsewjo9YvSXO0XJNWblSSYXJV+lWRW
ppsYP/PKHdfAF2lOVBkksmetiup457M+xpOMMTS/2yG7OIdVsNkyFZsQnjY/40hz
XLbfaneR37K3vVFs1DRdarzt/kUXhHGMTEDV5UPmvlrkltova00IY0o5jWm00VYT
OkEeV/hQWqs6yXRf1rY9mmWExy3h8O9tgNGOK1e4znd2lU0JzFBPXhUnWZtN+6+y
cRPwSQHyxCusQrPWWFygzLarPkcApIYPXQWM3JuUZukg8ufQ6ktnw5/004zIvc/Y
8ucKcHQTHKn4VUCUjWxCkEF1srmvSVUJ3TEVGjemlG6MFLzYynncaue9Xb/x4ePB
CTYNmwmAvQ3WlN67gIAQwXzJKVmCQSFF3l2nX5i5Rdk9+dYtYnVxWpghzKDakHFT
GXMvrabN+qFEKhRlQd/JOncxnQc3gt3/0KgVLJ6welQ9x/aWkq2RWWuS6X2oYOg7
WUtrq8GteLDMwOiCATSoSjbkFxzLir7nNF+0JegjQgjN7NRxRjuJdk4VT3o+C7D3
qYVV0XbLEWdayv2rVuxzafdEA3wKkjbe6QBemI9TesI7b7FLa8bZFaTA+zcfMZqk
NfcswQW7vgjePfoiul1SVAMZuZdm1OjIyUbzJMrTZD4DS/QW7/vp83ObObXuGZka
yKxwpsLgMXs+nBtkKTMkOEFPO3C7z72kzf6l9Yy0LkN9a7aOsKKz8DMkEx5oEfqd
oDu0+FRbddyHbyrjIU4IlM988VBDDK85GEiXTx3BHxVqNQAxduaur1krEYVYJyq3
dT5a8GLsHdq7/PGNNw4BZPwLdT2e7oqYmql2ewQH970lgi1L7dFI6ZDSfS4pjKG1
2lTvR4NaK12P+CdAaWkEhZZP9Q8j6kW14+5ljRdtU4FhtbpsvDs2soDIt6QSEQK0
oKsDmbqMXzYKqnTjCxFjzQzz/sIU1r3bUFiKeV+T1JPGUBXVDrQ977Z4nVSzT11V
DRs1UXQWG98H1VmDmGySI/mKgjC3VZEumkp/nWzd+HgrmtQRLGEKt+HDx8D27EFo
pO7MvPR/6XQd4+544zwUrbYyH/aaWSR4IUrXYkWmlFQzeK48CVdV50X4K79oxFSu
mhMd8vw4CjNH26Ay9tYfcKkQOOt1klxJYnkdFRyq5ZeWBCB0/UvBrLp+MqxrMAdo
v3U9InzOeWX+nhSkmFzEpAa7Mi/cwXOgP5VQHGMvyNPRUNFRdDfjcj18TMkwp8+o
1MixZKDHcqLYTZA9ZCqS4HzYos32KWw9o/9UK+iJIFIu/IiLYd0586qWLjWuASU8
qZqjo/dv6su22f5rjkld1LbiyOL3JFzqXNk5Tp8VnBIXktQON0IZQCgckpbMCvwy
Ummc3x/q3fj8QbG4hStuRVY2nCjqXDFF3TWgLdZQ5nuzzbgQA0r4tYvjaPASmOjX
sUjILIgpriJO8elAsu5aBnwxc8AOo1YBv+Btyi1Jimn6McqT0hG+jm4ljOs7Knx0
wwJjrMzmTOe8AXuTT5QSpvKZVk/9h2A9veQ1HZwFEIafU1AuOXFmlhcW3hHAFShN
NJpAPxDXjbezBgfd8Kgv+Z1P8hwa467Tvw3/sUVx+me4FD1uoov1gO5oE/wjvIw+
OsAdmFa4hW5XfW2MqedmyvD+Ygm6UKKK2DbglIDH7md+2/wSublP8ArOGRcb+RUI
zLtl0XMMszsgGUPZLhUT3VPSEVdU1ynrOm+3Q/e697f5PRGLgeLMBK5WBuzr3GLc
jRX/0Ud/2W1okvofRPaqK1ez8TqSReGoxQBwUbJd83hQsNgCL4W140QSDV7qA/tv
KP7+Uk9qW+KRzk5gSZ3q0YxvQvaFU4zANTaILCr514baEAagdSuJxSS2ThJcv0LL
+PN4vngzu7b7oyQppoX6yOyRpeDeX6J76MFBYXMO1l8oLE8Fietg4q8wxuj4Gwqv
RT8HRmrfaetDVvZUH8Lj7nsns4bjQxmzgATiwAgqIn8g8+UV0IUIA3npUmc+9ego
UQYFsgnLwB3SG/+MNW96CkdSQ/BRK7oj7xVyTdS+XYZCAWArvDk5RdD9VvXaAsA2
NZje/0ttYMcY6SXnkK+pfXmI7mat5TeYHw0Js/UELv8aA30jj3/e2sFvcT9/Bi8t
IE1c0rjxdEFhZidCQsmcBclQtbCfBFkrlVR8gC1LkkJTHp4OXtRsHGhWUJkEEK4Y
bPsZPfebBLJ7WOrFI8L6GcEepuTOguZXzEF2AuX2Cyb2mXCFZS83R5MQkzFp09qK
EC5xoJCV780LSzrrjIaIUjiBAxF8sNQ6Grcp+7mb65dNsv12suEBSi3V9CzpPifs
U9SMM7U01+drv4rPhdSqZ/6BCrQsZr3klCOhzavUP3n3ybBCH8AwcySJxn1ueHYA
7yOer4PwK28jq8SykaeNsXtDWbmbNNjhPC+zwS88sN6hvK+YFz/ZG57WJy5ujUJt
8AXk+ws5iYGSRDFj1V7K554YsM7LP70jJ/Xk6nh2D/EL6V/Y7diMpJU5+mcRtXmW
pgVO0EAUyEDHnKNvWtZBx2We6657psTdHoJuTp20z29tBZcl1ytVq/0Y8rHZ4pr9
ApXRv9FvBKq2N8AedZA6pG2CR1dlT/YBYoPP8iIxSGweQEoPJqZFZ6E549K1qsNg
rnwqfF3TqxWGdHorzEl1htSzvBDB7e5ADYToCOwDbZgWW5fjOAjHKuk/hcPPEdnv
yR7iQdd65wqNuoLOYNEtz6VUlLMUem3YL/SUmXF99qc9T4dDwH+sK495+bFed+uc
iP9V8Q7wc0krY/x2ZPkY2yJHjZ2gSREX4wdGNHbPeKETJNsMvF+lXICsOxhyr3XC
Uwo+0J8ECCyNqgwngJqB42ww3R5dvGJVp1L1Mz/Xan1JMlYYMnBWg9h9TNloaFAq
8ZAXIdpQWQRS27yVHy2D4CtakWTsrxAhPDUNegCu86ozsWfjwnNMTqJUE5FxR1v4
o5sorJp56fJIskeg3eoRp5YItyvVgF/6pcBSQUuxyGPALJTCoKlDx2K0nGXJ+/bk
nUJfbUygurw1cIqiQdq1uZ0pzfzICSyzobCGp9hrzso5uVqeHuWDKQntJtzIT4rc
QhS04NBSPQ94TWGPAyUI+wTAsp7vgBTNca5ajLLbDv8yTnVEAvOZR+UhK9M98aDZ
c4qAvSOEbGrdIzizTZfZc3LfbJrz4e2j+mTpcIStnCPwknvHY/0K0tfwIRFyYa9D
HD+Tbbisr/zD44SaLEpeRAq1C4ocDY18Qp18/wCmrC+K1gfwT6NGMwL419thfKFr
b5kYCDn/4CUCs55eCLcUDfXb0Xx2KrdvdrgLJRtKiumcVuGlsA04oUIUQ0sheWew
RPCzK6CAqW1I491BEoGYZK2Ey11STu4nn6OZrlFLKFZPS77jLZQe5e4CzqpDNDvG
p8x5OesdUuXFuWDNNfH3vle1GXbibUTl04N33sG//2hAFmaHcz/u91wBnfk2J7wI
vQCXoH+zZPt1NQrWrLaAz0muYzen0rdeTij1FgwJlCK7P173YZsULIKb+qFrvJ1y
eHt7RyIwYx14F38w8mqfYmbj/rqEvDEDxIXLoVMvvvMwqhTXISvkC7yOeGc7PgoW
tkXPVILgxDdxXoWNbZaok+NdlYLfOEXKtZrA5KYMfOqJE8vYQQZ3xsG76JP0xvq1
PKjNQyD8hgBhmtn1EdzYONKtLbPDebpwSeTBL14PBkTb6T/iKciYnBfBfcgbURf6
nDTbhiaBBf0Xs51xuJUvu4pkSTpZNVuOK0RFG/NzTpl6KE5dIhucYaT4Ls+NaLpm
oNqsrHI6lK6nkxZDeHZ0KIfRYvmzdzVw2q/PTzzSvwBh7Zdck9tK8UYEymbriz03
LSwS/srkkg9+4fbpbv/bw88f6OppXvQcK2sH3ZF+QgZgSAee/bBMv06O0PKXBOyd
BWF8CHSkAhfxqE893RvJR5tSG1HV209FVIUVeijBwHZ+r2G651LIXCBHwOYgho93
FZx09ip4oIDq4tFtYWBUhZBhL577FYFw6b9/w22W20sIxT/+drOhZsAEHHj680M0
qYB9k0+8KKNTBOlcaQ9/w+zZomW2xk87Rb+L49T2fvLQc/2bTPx8MrXfRIuEpuJH
pWkfQO+KZZ0RgFVTsnn8atBsgZyae9AGm+p/n5kBYii4ls1RdobWF3JfW0dLcKhd
kYHHsENcIYvR1EYJfLKCBVFPHrsEuzlHgI7PIqrndWr1M+zMPEfLywVrPH5UnIYF
+vAFXcwhNJSQ5efqXuYIt7TQFGGiNkhFQ1e5cfddrjwNHlDnkV8l+VPLM3Zxs7Vp
7UB/2d7O7aP9YKrcYHPGix191Hv2+yAk2ZydBi4p6b3kPgjTM4+kcKNJNBHf9WfS
foVSoevH1P7t5MZEaE2pbTgLkNl4v1xMtFt8qVKSWT5q951kzuQSnpGuGPUdZLgA
c4fr2+ZfyZI0MYW1KTA3PV9uGBdo4eOadfy3Z6loYPtU3Who/ztSA+26Ai/E+pdO
0qTFdJadqs5K5vjlq6p7NF8Kczy5E4VwoVonZwM5mmxG/8hkHkQp3TeVa1QUwwO6
2s/5OnR4q+zJaKexyHmDY/j61v2hxvCspXg3g38dWhUOAEVNgsoT2VN2Ygzu4SHt
BeUiKSwG7Myz7zU8b0R9UQFz3FjS9gps5Ivy63ns/Amk+i0cY/T0orDd6wdm4M8Z
jNJIjvTrqcIM2Nc0Wqvn88FGZwpj+i/zDVoVl6fpOzVmjevtz8Zl9GMuEEOotshp
bJCZLQx/fAMEuz30pY+LX7qVX2TiLIL/DQunADLXVO/2KPRjzFyakbI3Kz1io35X
diry+1SBWKn2iyPkVK5ewyDvIX+SSvgc5yIGZBbEdiPVuPC7srTRoWW3lJZef7EN
mLNIFbHCRLrSu4NwFnLKPrsR3L/VBbxnOMMrKWJSgmVOVeLIpzR3Rv6WZdqQB0xA
n67cG5LJAPLN0SfljShPjYtfESYxIby+LsmjCpoUuJGtISgm8+PWvWmEvpVmpaAV
M7IaUSH4yW6ei2OzjA3Y/8N2mOJ+u/TaKKsJ+Bf9bN9bVItpXxWxIELcGgOxDde1
aLFwn3yMkwM2o68Tiw5KNqFhd+tUlJk5MTzur54G8hGeTPSQMfACLwnKOCOUq91X
d6sb/oCg8Ef90CmTb/JXIGNAX/8RZetP69o0HlBV9iGiNJppjiOalyJxHpXyevje
DWFty9sSCjqHcecOVe0drXx7mz4wlfTeLlTIyWF87LPGlo0yfB8GwcEHcX0UAQxr
02F9IAHvcqzPmRbYWZyVDpYv5Uf9QFEN+vIljy35SDtQ0EkTaOczOIiul/iBXR+h
PyrPi3YCH2FokmyTjmdU5aS9XM/Pvr/5u0sO8Ax23wU5a/IVRLxwNoegxgnwjrn1
rRVyoPxYzUIqx1tQREasQq3Y3NcmjLckqYtH5ibsz9KBcXSgXr1QYjPN2rNh0xYp
BgZFDHqDE59LYiDUO48zNPXMn7h+20yti1SpNbowVpuv6GfpnQDih7xc8Ti3bGP3
3KlUx2fjTFd2t7o6b2FGgUbUpm6icwvuLREx9qH4kPzWIzs85Yip9Gep+JodnBGd
TZ0fn84PoArkHXXuhworr7UO8GKpMe68uPiGguPptkFW3G7sMs/tEoRI2CxS+N7I
Ij9brOTrApqr74DxsLdypeBAjjI746GNtxQdHAjqTEPXSbI8PKgsXrShfd03nbAg
IIRV5OboIn2PYSzgM+Bg14agTDCECt7rloNGzvJWUoDZx+xoWwLfy9HPUIvJtH8G
hLH+vBb08lD2L5MWcKHmhvKRY5qbwn35BcpCEqZhPK6khwkaIBI8i5qexONu7KVI
tr5kR+UNREN4cgewvR6hjKUWcgk/Ex8SAnhQ82bNvR5uEOjjnariBzVJ8TYD4Zxv
HclNKrI+3KCVJmq5uNrYftK/Zf85PR0uMZTgUZpdon6VTAH7fTfXtpVE8Er3I1wt
/neSnNGlPMFm9eG2EEtEfhFU5nKrzaKVS5+5MZgUWOopSq2RV8grqOOSkKZXgh+N
0cQAU0MXdon/eYxu+OEz4Mo/hlELsbAy0JnfZwzy5rkMu0HGVIKIwvqfRfJwbu8G
efsTaGWl5slmpHdH6Selmrru2yJIVr3wsjSgkPGMFR9XzbtiW9sAedV7bqOrVHlX
+U2ZLA0DZm9M6c39m/DcoCf+Jldh00RclHAY7lQsNkC3Bd52UudS1s/LOJScUjd1
48W5nYmW5Zm6OWPyaNOJkssoGHzThCNlmPWuj8KAOPa6mSzguj5ZvwkdwGDfSpOJ
nPXlntLkdFK4ylKm6RSVwdeaLVEzvy7GDCW3u0SCrky0JBRX0qfcpHffMcTQvV3G
O3rv3GqGp73Rsi4st/1u7XMCN4kdh9dUDY7mEqYP0Ecldy3qf7ht2i1JBissbBjK
WdUAOicIMqOctBMOXC6oLzx0boyjj5hgdLnizX/3U5R5QTXB/DuFkKmznXcAj3tk
ipGLHNU9K/iZDKIV/63t90NXDGhWEo57i8prpSMyTAf9BIqJOOd++LTxnbjCoGls
iTsAXkVxe1REuGsqWruOgoMRbf1D4v7JNHp8BeEE+FCpWeR6J4zpNBQVYA/9YhDd
4GIeK8RXjzsulfO9qVnjP/Plmttq1Efgyr1Sked8/anRao4lLpfKgiGseXbG9ixu
uz8mIcGEcd8aRSNToG/Zzw0ZHFic6OFg1TDW/Y3XI8/qHLSu1q1EORuuoAKRCGsP
TLv9ZjX5snMBfB9BnU50Si016qXj5IU+efyEPKjxSy4K5fb90T2LR7IJsUVQzCFI
VWKPXkIb7sxPrFziNoXlWot9NNd0Lj0BZP1NgU+8mkUTw3uIAQbjQg4v9UEGvh3M
X94iWxYQ8SWVJbHb63X+TLJWbvzBP5X4zzx2t7b5dr0zvt5OU1M9khdqJ5Cqyq69
ozH+a/fPKeIZtArMvkUhP6XqQvAsW8uNA8EdbyvJFFRv09cvXbFr/95+eni3ra2l
qz79WuN6pgk7PUGTQNgRO96cSpxE6k7VPailF7luOAPTZKTC10nD/c+HA1WDZ5FK
ZEGHBeAGTQZWlOMid2joHEa1t668eUfemAjC40brU8XvgGwfUSfDdut6zw/8DUVq
b+mX/+EkRomyhrpyDSKU4LjAQdidhp/mNsgJUWgN8H8YX8kSMqAnp9NQMVg+wpwk
j2R8BYrWVvwhNCHxUQ3tzYBS+is56NSA1KReiVjDl8eDhJxlayQu5BzSkZ/oL4XG
0faarPwUNz3PmJDGCKs7W1nox1O+GSZStJ6JY1lJzoicaUDN6wO6IAHHnw+KTHzA
lWzMSYAgr59BM9EZuVjkL+Fihs6gOIiOQySJGIMk7bYbIWSPWJE9LsWy+st5/xea
FNAio3ATdYEkODKRkiiUDDzhnA4UAnpG7wdqWOev8348zFvLaV3B/LyZKToiknNx
uvrzzUDtvp9B86OSkNDuJ86sWpSeQvkvvKe6skqzG1/MBW1TFUWpfKsby5GFFR+H
2K0adWxzrPEAvxrKXL3UmT0DFpML4+9k+HBhaJakNZpwc8+QMbtQMtc6eAFi6kIp
xN6SEUaSTdmDrCabOd04UBUibZgykoV22G4mZqgdx/E8akynDkacEAMZ/VPd+ERm
3guU4ir4UgNtPO4muK0p48Yxx6eBytn+c7JuvqA6bY+fcU10Vs1h+LMkHhoUws3I
wlVyY5uXf3LEMuN0YeptsxSpOJEHxgJYUNYc+mJ8QM9TiJBApt8xKUI4lBB7a/Br
OxRSsxOzXuFLySv26S7X1sSucHo65tMgrROkM2+c+DUY8c9eZBEriVKFWa3I2mPe
5/SpR2g4xylnPgWEnuxeSi90oPZrosDTmJh4w3FVlqT84f4q7uduy/i7sg1JYWBW
h37Qyfq2JFW5MNoPzATpXLTqy16mPGTLtKO3tN5aGyztcI5wt1yQ1p9D/WfDg0x6
mpIEBzMO1L/4NI++cECWe+wqqQ9xuQTuJIWVnyh99pfBMdwFaa4AD7Pxn2vi+18z
70U68pU2K7xfk1kpNhcrSya5fBBc08RLl8yeNwHjAIDrEESDyDs4AD/8uXQ3Wecf
7HfCC+GsZdPoWeOBwB1XqLGIsv40GkXXCKnVgGaHeBvI/HYyUE9YSLTtqu6SynAf
7IUFZsrm3W7gLAN1jVXXjAKVje7dd7fmS9t7N8hWYEqJWV7msERd/ngLCptiT4Vo
ZOgci/ywlsSjZx6/8gzu8UE6/BKddQtjfy4Lf+1jrYgjnhJ6IpkERTJxSXNeh9xC
piJTYIOmOomFzqPiDLWq64dEBdc3PTP3X1kLGgaO0hC7cYrbYpn6u2+f5KY0cly/
gd8Z9NJpnqZAeB8NH8JKJKKqWS+f1lTGYz2dDU5HfpzORS64vac27vL3JLbtj7jb
sv/3b4EFoOmitTAUCecv11FlIqei9pzHIWuA4a1ZSTlKZjuIqj6vKcg5ULkil79g
v0V1TEtEeJFdXxPKXNCtrnKnwIZzS09kx+9ZPowITuRtxyjVC7nrs5iUxKSuCJ2x
iackNHYKThlsFfSoKINPql7Tujco5WTYhgJDXHEfrPIvoywDLBYeI/rbPjtMAC+T
rGNGhSSfCc0uCk3/34ZSEq1cT0VILvkudJF+TDF1Ke9yGUgk14CjrStmyDwX3OsF
VqcEv1OFR7WLs54rHubAdbS/YMbsmXdauLO7WIrf+BZKMe55YErzFopGu9kSVj8v
TpxTEnb8+d3wpRi92isGPF2TaQYjqDcr1LAXjkd5EpnBHF0XUSEWk3QRQY3gpUb+
1f4lisVbs6YuaNx9igYGb347guvOR4vBZXstRjg1dH1b/nFgNUJPH4wH8t29Z5p6
gcsHpH4xNPYcEfMaEL9yxRas1OI7Zs/gtsVggs1w8mO4b7SHAcQmt8sORUhsMTDv
Yk1NdYzeLD8HABNYHp5QR+iTc+4XH/XvKwn0eLH2BTY2PUf3bv1Db35YC6n+o3LX
OGyklgAxymf7FYyyuyVOZr9ND+AlMOxEIN8QqWYrZEvnnJmi+TRUjsbSvhcxWp1P
sMvGg28xxczacY/sIfZueHGitQeYTfdzJ8+NWrjEt+LL/yLBJdxg1Ievkmj0Vlqq
59TTE4Y2zvfPbJWxPR9wnYS8L/MJAx0mRAC5j7d5WlMsKjnTHKwRNp+O8Rx/x12L
2Xr3uBBrN+m0ZSu0Wbfxm2igSYkHR7WN4X/MD1uzO3FkrNGqQLhcsSkOi4iD8Wur
rW62sxuZOqTj9rDOUgBGRF8FIMUyUhuZJHI5ahoree7bJmEbTwXmtF1v3aM9CVp/
BIOBguY1STIaFUFJdjg9HekHUoEA3FT81+p1NBD9XPyEh6IPLjdLdDgGN0Kclklz
WNJz+MWukXaa6XEfjFB5da8AQBmYep6UdZAdDLkUruMdqDwDx4WyJrlIG/NnREG6
RBON1lsMlc4Xgg6i+6DVqD0pcqkgpub0MmmVsk1ax6zVHtwtX9c0uzm5cRg2+J90
dE7FV5yfuku9Ssi6ZRVF/IrH7bQixHU8U/lCORH9yz4z1ecCJAisc/REZO1O45kU
z5MSWVSSPJ6Pslv+tso4840u04gROF2yKnS0O9raus/WvdLp3MkBo1HOZzjTeF4x
XaCZvBKerOvuiZST8V8eoXnAThZdhXmz2F2TuOBzopvzVyHogHzJGNxk99PhSVLo
OHoVrf43q9FqyX3uNy+XsE45yTNDSGZcPQE/82gptPx4kVgK5wPkS35iD17Nldsq
wbLkAPdTn7YjWYkahAmQohyi8G+T9Q1QBz1Evri5k27OzCR3FqtMJsxHRGWWSUQ6
9R5q7zNOscfWxsZd8zUwRpsyIshE55YU+lD9YuKla6ZE/ycIcRzJbsnN2V0AEPrE
Omedck4k+3QcL5qKJbvW5Q++hC2O3HIw1sai/sckQo3RLkWFEtDjoqJQNTfR8eAZ
EyxWI8VvG2mfCOLohQoIQS3Jdp16c1Unnl/nPoVAT7/HtwYBi3+6Vpkd0KsGvhm5
h6eC4+D+AdBK0zgjtpDv1rnhIWIJY82qWFf+UW5PbQwBCOFbTMb2GMH7HclsPKEg
+eUos+4FEzA8fry6wRXOpGfg17s7negA2mZDpRXhMsxD7C2zjPKT2yPWWQWJFpTB
inDtI/IgSDMFzCEB1J6zobnSntDTGRe91/TzJzcvHRhvxCWUl1r8NSwjACv0RrTJ
8B90qHYAmND0B+TyQRJOA4PMzm5Kk6LHs37CSKVNpSPgC9/GLD77HdqVyuETUp1C
av4Ny8sAy3cvs3ArxEq5KDBRBnkv5HvEKh6+Z/oPXEHoOHdYb/BVddySpIIywfZc
Zdit1hkR0Uz9GjCGDbcqbWh7vkqTpi4CZB2qRWNTeklndRkSevCU3YksAmG9tPs4
kw+Wmuwa9YXyOUQBu0DMwMmS5U7d6Q8gppcWWpwTWYBEYgmFqciqXwSXBRmHfUL1
+CKGZuGtLkpzxl66ZuyUd6uqKRdg2YnXGg8qYZuN7LRg/wMwccDmm3AWoxIohBYE
viQmels0MYaWfxA975bJ7Mn41Kzr0dMKxvyy48HhSf8CzQjVIMwFv2P5DTCvQfaW
WkaKXYuvwb8qbahzv28vKf8l9u6lCXzpfXkTFYjo4rzA6h3icUE8bhmxC/CbeRdz
8LqIL8FevMQcEaM5lZveX6ennbP2QKcq1FKZ5dd5VknY4kq0Orqb5F6qGC+wJMk5
VUWi50vGSvW46x4V+prxWd4Q6EK0aBlziWHHoZXcv4kovF4KXR0sggjmoLwMwR+g
MyegnLroRApkMqeSwSvazQUcnJVS4Dar4BAgSL3tDN9aEq1SVpJGUoYa/QgMIuUZ
ZyYosGpNVuF15WWkPZvSZJsIQCCxvBOzz0+CJBGbI+IRAbSMJDA/QJ6DLemHISB1
mXfobY9mlLjGoeiTo/eWqAIuKqB5Y03XNW4SX59svzv2Mz85KrtCvJCkUSyMccID
g9B2LVtAMsioLiuGNKxxVPEGv3z5lQTE20E1Jjzv0tSFpQkh12twoEl5ZUDXNln2
1yg/NGeZl6WPsvzKD46OFvRpP40Sjy4c6UP27qbmrkXwPHjYUk1nSob8d3EbhBrX
AMkV6fBZ39q++WAuG1+rjsf9Y0+wHUyr9XJLM8C2PeSe06XWHsv8qbT2tIUiArnb
UgdUI33iEIOe6TISuAha6htsPSpOV8yjVY0qQLXwUirVmKrX8oLOpuuJKrioHZiY
PxUN5oXS5vzeXFo1ygxVo9Wk5MFjmpqy5hPHabm1HrwMDpUH2diOhQHHqUbcoHB9
EQ6wBPor0+K5WZViTycTXEPBE2IgLfIa0e506ITFX6fVGA5Ae+NlAlmQlHSJz2ck
T473CAcuwbGDzxXI8VWHBbn4AeFlY4orh44zL+2QLY00J51R4eNsPf9dAETxh0cU
5Unbh/CghdjwPnwCkApr10o0vkvxkgI8duleLHttLAStWGLJ/2Weg7PNnIrLVZd4
zYALiEALHG2IS/pPua5iiINE7/UoR6mVZXL12I5vLe1sqeV0KY5tzSYxStPcziaD
5D/HBr3Y7SfNTX93/Be/uSU1xrSA84EA0yTNadtRDAgm5ZWC1/FWVMMmgAkFi5GD
Ps3B96f0I2aIh+8mkUAMVockm8FoLNv99LWYJ2J2DHlXipvqu2DScKZDfXD/qdLV
fy4xEZwsTqti83A7d8/oZvosJ+gptgYFlCG+EfVG95/nj9sJO0+BuKm6GwDuM/Ze
ZLP6xwzCEPU9R0CjQbH1sy8CAPbQbkIii8EG9agzsrVZMtVPyWdBgJdQcVVjrWTx
PwO9msqaV0HHjkUlzm3xerV82SZRk6o8kxu2iSQQYvwMf54A2RasJ9NQHelsCwES
eVmmPfh/wTYtKhQZmCQYNMIB58D883iatTZ+ZeHym7NtkiFz2WcdwpJ2ViWMyhad
DNPaMm+V+L5/6o20YSregveSyTiPqt2jX5TuYrY9WALBSH9BMKA7jIGbYqpp4YyG
VdAmI3BJULt8LWKN+jW95Nv6xkwwHyKiqZ9uaKxadFFqUCPsQF8ZecBuzxp/HRDN
fexx1KKLRZbZLvZwQEnq9ni00UKUe5NkgIkLC+N/caU0bXDXcXgnkarcxTx9x23U
zVCFDNVDtTI/z2Gkw1g1r6FtRYwgE5HQqbHagWSdW6g6AceeH3jze9lXjHbLCfhe
x+StTih1WprHZA9CuMARkg8dh0bRBhROnPufmJK2GvMgSoTiLpk4h01gjrjiiHlG
7ILKpfI35NcHBfpBxTkPi4ZGZx3dBI23rAv+svuAjO/cqbD/DnbBS6NC9BKdsgsL
jw6hxfeWzba/SQdmx1ZNEmlm3axB+V4o9RZ+tCMoeTWf9YYTttwY6VX1tvLU5zqO
ytp5vP7CdeANd1Eeddr0AY7+9i/kg8jk1JoEDf653peHi/78YLDN9BC6zub4j2+m
x8roGGFRxrCooMqVONTebikIJ/DCxM8i1toudMG9REQZ2BjdeHKJr+LDYeXUJP6z
CY0/Ju6MWXH6Rb5aach/VQ/RIABbApcHB2CCAdIwXDE+/wSujNO442RPUc//xSuR
u/v3XTA2mqhSV7ZTGH18Ovs/9g0ITttWAurmA1m4sZ++KQsTUZJeNdt4Cw3GnnO7
U1ZikaQrgut/Mn0ZRbbVJsQnpa7uDMjvpaLU71i5D7V39QXHRbPtjyP4Rc/KjDCw
5M/upISDzecjAigGUjhmLIkxueFc5UcR11e+y5cZXNMEBgF04uv9wLsMRh9S7Jxi
jga48gIMMRm6U6pcLGHQVhDe53BL6Qve/eJNWHX23vuTq93nTz0YdHXUV9r6+Qyj
TWwFHKR0HLzBwvV9edDt5xtEvrAZFeJa0QVkQGWKcpmnj81FIS4wkIKkp/uyzwVt
g75d45JIjcy+OR9t+D/LgG2GDVy3akp21FGaRJQFAKgWMnCTiPz1mZvPA2iBY2V6
1AczWjlUs4RIvQvAOAB3xIOO3m4+HYB7Bm6B6aBRBY/xVZw6Yx11VQrcSZ5fA2/C
2mXPaXg5f+w3yN5Tqnvno2rfdskiXk4UeIaGpkEDHqnhHm27Fizf9eSLsnpHauMZ
jmel5/xMTkX5+roK4gZVZrQJZ9TBoAniXpeiucx/hjFYW/4n4DxYVpTAucqSUWyK
UZ/Ipx/+N8ZLbKzEBcBhTQDKAJ9VXYggIrvrmACz65JMPxIO9NUYANEpFvDPRZ0q
wb+i7XN/dAfe3PYCsWPyUe4FDF+zRQSZvc1mbZa/xhuSGfQz+eW7mYCw4WGrCCIo
DJzBAf9km8UqD+mrbmTlh4BABrdnEx15clNuwK5t3t/J5VLZ1ULAkDF40kYjHGMI
2VPyFlUkqxsTnsBGMgPFE5ND9n95Wg5VDz8h7laMjP1R+Gk24beIJaT7/m2IqPdn
JM+MTvrMI6032I/wr+qmAxtpKq29SzFZ8iANpY76Ypq3/Z/aPR6yXoDjF8a3eloL
JPssyim9Vsx8NgAMpSUHXxapbW6cO8hS4TvDLBC8NXbxtFULyYdYxowXBStvLFHN
JOOTvwWWJEYHbZv8gYN7xT5v4xWLsgUqy3z+zHEbmKpHG/c1mG3iG9LgcEuLEgZS
5E6rBNwgUu1zgIxHpPEszp1qukLjbmOjWVFRHN76Qzz1499Vm7zV4nJdCtYWULDy
3nChVYSJaRKIaoefjsDUO8dRrfuAL8tEBqMEg7IHaofggSgX6ZdhSHgXniVdJoCc
I/Ze4DX2IhM+eboNbY+w+0KUJla3CyoO/jW2+7j2+dETuxP2pawrvn2UlQKsLKkM
PU+NA7RI/FbqDM4M4fnsxFl8dhLaRpPQlCoYkEpfvV3nEs58vNJS8dBV4Bei+bVR
vDVQTZKndm6s+/XhuGt//S3Dp/Ndr4YPB+cDar7235xkRz1EE/1AqGtfAohwIsWZ
odbhfujh95iu7ENVGuQM157jRgTOEb40uGSzT+EJ/Tw8O3njt9wtVSIIuvODS/ox
hGYkerpuXRDw2j+ZppCG5ABLlf17RG5p5mUqNQX8i51kOOs1WLE2Hn3Svgm2SRRd
PqGWCZa1zhxkLsIf7PcbWsZvzv8ED7iljujwUagXw4Ux5DpEU8w8j4evxK5neCU4
sH3N62mrfg9QDs0SvledV0T0wazJUWCddj+SLr3s33iDUnF3JhMZGq0OdFlrquW1
CB1/J8+uAa1ii3fiORBz5VdgdSRjyAzqQVlYjtX0zP9vycnGZgq8LBGhGnhpQmKK
XRjCZBT1lFOnWGQ7fSC7L9KKTl9g+1ZBnnHdnS9iPZMDbp226et8qwV7tco0I72M
E0/acDi58/tl/D8nNFH57M+I3sitOtYhz4/GgelpspGlhfvOWSiwlAlvyBb80+K4
bZZCmlt9u6qSld2xuqCdE+jsTChdfhGUoAtUZ2WXEwN0q4E9QI2Aj2BcYBJeKGF+
8OBo1vVgjcuTFXafXMMfveeSOQysZ2U0YQ2KwcjCGK/FTr0UiHGsVgHU4Znlkd0X
y3y+q9H1i98znpYMq06TcICz95O//JMZ6iaYodfGOPnQYzYE0pTjAmCJqt/ZLO72
rON4s2Bfn/WswQ2qlfUiMNbr5YzrB58v+6sJHHE04fa7ZeFBCb9lYfXNWx61VWO0
P/LhW5cEsy1ZEsBEwUo3992AFgDh/uKpbRzfkbdH+AotAgM/4tI1k6ZGak8a2K0u
rf/ujBFo2WzGxjW1IFDdbKWlDm4PREnS1fx0EkMcoAE2vp+Fw8ZXMdJJ2RJ48Im0
y+vut6ujrQMIiR7i/nznQxl00sef95xDRiIoVmFbOiHHpLqPcr+S56C3nlEd5z/g
24WIHJhPOoF35/DyOAu00BOkyYTsCIOw9Zh521fnGz+uw3s3SmkdO/vunkGImZ7v
SZ6pBTxJRc3PN4J0JE6gY0I2NiaPEFT2xeSviTt5nTZBVbTPw8g4ABN3WY1onlwz
Hmx3WwWgYHwx6/MbmpUbto/ioR9sKpGHaju9JDxmXgK6VI2CU2oviznOdzBWajMQ
lv6wzFWAfDWkvg2lgubOdgTMF/CPvAKzMNJyvaKpf9DnHZAi6Mig5lgd+L8TOKJR
ON6YGNOPWkWJiJJKrkQz3VteE0QryUwIk70CO2VrVz+vUit6Gp5H7kRpGLzsAgJR
gcmBX0iCNXdQfIvjuE7aR6KdFPqUj4g3AJaZyQg4burR9IZl7At20oEvQE1bZyLw
nvaeLx1gV61CWsyKpLXBkJ9Kgi2CcEXcfbvOgoD3hx6KaBnjyFPqm0RTMAwQrMGl
97ySWfPbpx85llhNjYcNvEjAAAGGu4ZG/V0W3a+870iwtadT3Ueuqzq4Op3gyY7z
fChdPiYdlPlgBOCW/vWdJQjUiOvubWBnro6JTUrFfWcgCAO0vSHynVR9hgrRUUwG
b2UVciDRwuDEo9O72g3Y9NXQjMn/37W6fkykQuSEM43PXny+1y6FAvD49LJz3m4h
DUPGCQ7nMgVuWqVPiUrVwTu5zBTaN815C8022x3+wJunHwmA2HJgZH9JiylcnjNU
ABQBoJif1SL57CvmnXhB48jcfy8L/FCDUw+HAvgAFxrvESH8B/BjMeK9Z9F+8Ovb
nu0RUL1zI4NrbsSe2cDNguZcK9Y34/mEcAYba7P717Fqt9rjukKhHrqecFdy+Mkv
Q9KRoqNDPwSbCL33ayLT6zE6bEpLEgw5Hahi46VGzdODPeuL6MZz7qhoozGW60Mx
k4s7YbIOQKwZksPbk9SHTcB5R7plDQ5ji0ubTY6ab1+3igz5kjKw36BS8qftdgeB
4iFLAuxyseCTcOtK5n5o1DjLdhLSK8Z5JVKk9uqmrULeR57K2/PRvEGtnZjJ5gIk
n2QwlCT9zdy0rLLhjJFSQtT5CHj1QiWooD932/2OLpDMgpfP/TrFZ9WBO1jt9lfB
kNV1EYw81lP5cae3iyF+Qh0t1woyQFIqwYABY7EX2HElMHQWs2DKJOJerMtTCYj6
OVSF+9YJgHOFYKgbzTLoKycZi5evcdDSKKY7BCQtrBFrTxMOlLeCzX4uAT0uRDF0
AhNwRLtezzuUBhhK97DLEk/ceu79dnmLyJKCFZa5X7Za8qsCszWow4INL4g123wX
wftcTCQRoiVLsR2kwlMRZZUXv8JenQ5Lx5OYlbRNJKRm8xrCdMAbq3S6TkXy8yQZ
xcuv4IK5WRUutPio8kwLuHLIlUykJ/GkMLdtW6iGmaLyTETb15QGSz1tBH4YHL2E
G0qtjD9UAXGi89PzEeamggnpbP9mQYfx1gGZSVjnjbkTamYBgNIAFvYEO81OjAWB
RHHSTRFcC7MSyBBl5vsKenpuzw7bR9U3uf2LRMArL6iNDJ324k5gSGnuFTJm/n3K
ZPU0/iESRP3Vf5j4w0x8LxQyOVsaf7PJmngr9zXCFtP2AAZH96+gNaRg9e7cgEAf
vXNl6D/KGy4y2HM78jwSh0jmyu6hfaM5aoUwt34p90gISRz6h2kSzJ2I5ysGlpRZ
N1NIL/pALsRcValdnbCfRZV5OxQivG5B9XQKiMTlBUw1G32V+ZdywuN3Gbx0S7wB
DlptrPvVhr3YjmUOdhigLFQblrqq8J3LyV8WyvsKUqOgkCKVa+9EUYqUb7pDKguU
Z69mDkfprl+owaxFu5Z1rZpgxXiPjaYYaVqXmkHkYmx28k+z68ZEChf1tf0uXCTY
lng6a7sHTzL3TMXXFAGnBYCqZrvuKUUgcTA12ig7LlyOdWN73HTBPK06e4dDwPtG
xhYwrbiHwHCAfOWEQPT8dMiRLyC53kdvuc0Sx6qVYBCbC7YeSe85o5MIyjHiMg+t
uy3aoL5sHdF43uOUL2sjcTL3qsC3gL4/lOlSBB1A50O5uDBctVHJmfQeCwpGDoJZ
PLIyJWsgPp37MRhqm6lTlgjTD19qWI8LLUZ3fwLGUzz8sh5j7Vtes6cw7RE62Q6i
lfu42x6fV22lzRc8V5aoEPz+phht3d9+LOLrnsrlBt685gLHDdFzbnj69WbRFNFs
T2kQVwdt8lATwN8F589ii1j3QLE1J0avIXUXrSD9IJySYfLsDhp0zO/CYPAnjE/u
pX8aKUCd7vbpCEPm77lxHkYkOHOBblQ9iH/pDueu63VEA9+PWkx2T31i24sc0gP3
CLuAouc0zDkSYki5rLxo2hVxAbwlG8xvubeD+80E4H+OCNueYIuqMZVD+BkIIynX
KuWn4stSENvo8SDr8DiMAbl1CCz9De8EiZ2dRhAZIsHO2W3rajvO/sesKKX+C8Qe
NhvMr5jj13cyPbmL++fVt5cDNwTEyZckUMBJ1tV+z3vxZmbhE4zHQRwJA2odoFrq
47tUOj78lkTzfYbwrcKijePNnDpcYrT9gY2nLDnS54H9PEfQ0UPAsbFXpJno0hz4
RENQgK/XyirrQc37DbX1QNLaXXgBbjqnw5gfPEKQ6SI12e9KEbT+uy2ck6HC+q6G
EZsthVLiOt6OYnxAPJa2ob7SsWmr6TWLg7e3cKXBdNQxhI8f727FsYpUi220qUVE
KEPmXAZWSLpQxAonpHl1kvhajivRdqloUmcTu0wycy0zyAnZtUQTlHkJJ7ZmU5P1
z77TY88Dq0dczrya2uH3t1pdLkpgIHByvOYpuBr0de7YGtub16GSeNG63eqb1GMF
6QSy2w/KptRNwyv5DQZEykkDBpfvbdyQ9A0b1woEgH3nQR2YY2tx2CXtQtcT7N1o
wvTkBq6W/vCXtq0ofIIS0YoW4eGpOnK/Ktxc9/kiZsS347MYcbJgGseSIUrOIyin
FokEAwofExbrTxetzPW57rLtwPj8cXWUeSOwMsu+MR+cyk9kvSz4nfNQCoJhTC6y
9Ih+YhpJkNfaJxf+Nj0VDzqBOUMkS1fIM3H3UN0l9xOqTgmTWhAoW+GGjTVjqLvN
8ak1TqoVVzY2B99PHG7NYouHT5Qy2fG3n0xYo9G9VVeUZ8pscC+AwRmDzGPvh/w0
I6OQTqmD2aui8YDeB/yjIJUgVUuzXi3E59BhcDim9zu2LXhFfkzAFr6/2Il+LUN8
0uXiX98WZ/9QxQNT2sAbzCwQcfE+34xEVdNOqHR2PuNO4K4y7wDYFqc6wv9Mzb1X
9EKzfHY+nR8aT2Nkgj4MKtoIwXuMEb6Lgt96bJtlolhj96d+A2XKewYFc/aAblef
WCTvVNYB6Ox9y01tvK0CVxI+4qKoGl0d5HVMhnaEMLjQsm+FEiloGkDZLk1s2rJf
xPCMeGFgiSCDbTBhifTvHgv0esz1QI1cWLrdYKL0pZ8A8f+uejSxq03Ec4dRs15v
DteaxFZT9xo6IRoUVuZrOP/yekrNuNhzniM74avJXS0JVuzpPk/sBj1p+KSqKg1/
dsGznrIqg/5YjJTBnQ+8JpU/D/pJcl1pBtVksr1rvvmJ1yryx+S5JY4IoYED7dMZ
w5JzdZEDnnkKmaDbfkKEyhvRxHkeFJXdI3UUvWE6jZg2Kz48iSOYjp+LbBunET01
2EwzReLPdawenDT5qDvuMENEWXeAd//u0N+645N6RQBoLylvJUIU6KzbZuckJLgC
UFhh+LfAxB1YwYgo+z05Ylt2I2qPCGjLKpOo6+f5r88HLTdm4LsMQOkktaZZyyz7
9gg8v5sSx2mWknD7cxzlNYWPvLO9+9S5fwY5HWZNReFhRoDARbo+cHkid8yoSOxF
QiKOv1Grryw1aGS1Q7r00oX7ibSx/uGdrlYmjDZJNGznuquHQW/iCtczoWrCjDXF
RPDEAW4efy8Fzl+vPu63pTcdNagMJJFgEBPx+u13BF7QLRmso1pWmXfezlmMx/7U
yV4PRSAjhDAqvrR9Q8LIyl82m19uZPSrCyFq/NPAtpx2GsmZF+7ZN8u963RvFOFq
B4VxP2Vs4uHqEB+0A4phw0oLoSzAJ0cyCUlCQ60qfxMGvvwpka5IKjyDoTAcyeyQ
WBDhcpJG/kxtD9qrLlr5ugFk0AhiA7glyUGTC1oCmj4+DwxeEDG0eGdcvcri7MCr
1+EgL5sHY5j50ZpdWXOFWwMcNURsKAVqwjTCPrCe3viUH3s0cR40pa1jlQUDl6Y9
T9mHQdGU2/bP6qQGAX4lz2sANK+Yy1Q67mPZfHZvW/UeDBKH8EP5xaop4wcKJa0B
c1DH5jZBFKgGuN4bg+mz7joY+nLtil3oBgblVgms53Aq/Xt3S5TiuP0HlfmUaXLj
uAQrj90xT4TnE2wEvnNqkILZHYtqGQPG0k/1m2i5mtOsVZg/alXeCBd8Ys4upsLI
+o5KHl5Alt7riskZI8HU3K+nI0IzUzGEo9wwo11FlE/pU+GMsAF4FAYEQdIQGRd6
Rgy/ToeDjEAuYY6rP5tw8cwsBxyHUGVRnvPN0p5UDfgjxsTFZO7oAII0KrQbbQ+2
6sJ253EO4T6idFzaElGtkehsyoXRjhAiZaJmU/OMXp3NxWG3OacoUeHUxWrDoSxY
0z4GKAolkhOMCXYfmKIWmssB9RXeExKi9JUBPbB2i4qwUytPVKDztplg4hIBgDWA
O/iBasoZ+5cFM6JZm3ThmFplEyj9H4fIR6cPqUOs6rrc9uwUkBmFT+/Epqg8gAfs
iDEesxkLdQP7Wf07XOMCmERT0QCOFdtpcplgXgYBwHKRKxQSAHyaOxw6NX3vZAE/
1BiYTldAnsZYMKvgvOMRiEMUfUtkcMJENG37MrGSchDdsKO79+N2V22ObNEmwuZ2
8HtdNRduwTKIb47hl4BmhSok8XzITpFugGbYZGvNicBbP7Dsc1/5lEnnJfDeqhu4
jcgyiUoy/ya7dVj0OQ7vXPYwtlHm3zkL0yF74p71ts39A7Bw5RDa+z6ykbSdgJGM
ZX2e0+WB2UEeDus4pnq+1P2ohqEkqkO0jM9++qA2Phk3bPxN7niXtxN890arS5zS
XbHlUZu2R4CfWQ2rXzlR18k19KvK4g3EeVApnuzK8dcCuWMP0WDTI7opPNvAXf5h
T3w4U7H3GccTGkiYYpdTZ/BKMxPe6o/jMS4j+2+UCnXjRmMaIQ0BicLiI2zd1f/f
pJRB/IZt8aGR4cT6KE/6QP3nxzLGfY0edQlr6p46JlbrOwuOcUzQK8oycz8y/CA/
NUpFGYu60fw/5da+QUDq584gwaC8NSVr83CsQQZJVFN25nwYkQ2uv9fGwYSuEi46
KJ8IOlAFPtWRNs+Xy9URfee4zJ4eDtVH0EF/7BLLlyg2tW42w7xv/Q0SQozXVtT7
lMMpGCG36IkzPFB1CceCin6aeMf2KTc3O8W/4xACsU2i8I2GCXPfwmqz8p8SJ21f
9cnJ3bITnpf48sEbGJJSmDlA2c2T2kC6Laaja9+g3Iwub4pCmdidbNF0JFTl/9hG
ttua6r/oJLk0qfbOBnKHqkh8RVENvUTfbJvajXCFMJO5RB/zRtc0eqVj85UBLTgk
o127fONskUQTT0iJiQoXqxSzyxkOTrvDeTzEtsYYptu2vqlDNZZi6zmKo7Mf5JoW
cnyQK6HU+s/95Ww13nb4/sovHsH6Hwk5nSfZOawv1g9Pz6KjwAODlL2obvdCnnDj
xQQn7EOtUY5XMjlXXv+qdRYxe5yHsrjX12W5Sp9rGLcfQZqoHauTrfYw4NXefZKV
q1fLW7dMGFnLoqZRYB3RfF6TNHjf3sFaU2IlUE/AXh4K+RpHboxFONPKW1V0GmgT
NU+amwQ2XwroFyUpM4b71u/a8VFWQq75nqZzvY4jpfPIHGLfmwX2S5fWb9vQLQ5g
auZgj5xSVSf58juwkKqTm6VqiZZXkQazcH+WzU6ug79kRQ1an7J+f95qsV6dV+gc
XjfbRpq3gUJtVa78U0vNsbVCg0tz2LU4zENyQtIA6HamPklH07vzMkhn8D8Cun5Z
b/LPd5W8nYGYOPMRZaKg/cNQF9KYjjm5YkNu19ku6W6SFavP1PH1zvesyHHoQvOC
o7oF7reSURGwpJxA3XsBWEeJQ0LGSgJ7xkqW2PAgasmVlv9cAwR2GB0t0ucY6qsk
mUJyNjUAirdPosgYRaO3gprF1FkqPd555E8p+HcDd2Xl4TwkfhKp1SWyosFJZ9iL
F4DgE6QVyz6v8HB0ArnuBv1VHeqbVOSIiPG565mcQs3USbCPJlxB1gcm2hQjmfaO
k5i+s75IlFfqvekr/ac5X6vXzy4htrKOebA8NTWUgSA1l+CFNGyi1swnUgjqZTpx
qaTKvRCGHZEWM1nTe2rqikEFeNlvfueVH6CWiqJyzHN5fky1nbPh4uhqtzS6GuLw
xJRdq262Twz5suMYtFl4/29rdPQvhk0LmWd0XjIvh0nOIGgEnsJ7s0FONmLQzTEA
9WgeMz1F9F/yagqgPbiT0lf+nff+S6qLWvnIjKK2QYXtObMv2E97SoQz03QNkj64
SE0gXIfBGB5ArgrjAZfya7iNWBp/1dU81A9rPBZA+46btN73+fbFWalytYGD1mCS
VGdG2SQVl3y9QoVq56v0xGKZtiAjupEV+b34bkax8SWiJcvt2Y/YPu4zx4PCaOej
tltEI6pGADL0cYY6CT+rjtBYO+lnk545qRgoc/S4pd/h4uyBdw600bqlgRrSpKSP
4Pj3fywyEuer/lU2OuRkKMWe9n9ezgi7tZnk/M0ETBdm9hKk+EiUavxqyCwhASj7
ezyfKP+FenEZmt2JnRlKFd8WpyM+GJVjjTz33aaB9uBLQrDnJzibEPfTVNArZfVG
JyyKKC2qUCBqL3I9ovxTImzrJ7cPZyocxT19lhIsxo2/ygmUsiE1x7auFuwtSIlK
kYsYMMSs0radEdaCwDOae+ZTIrRR+vNFRZT/vcBzvRuDZnweBQEXrYZ5HP6G5U+P
5BCdZWo8njojftLwq4HWWdtynxvb4efjbpFCBXd5KO8sXnU3nEqvHgJ2woU64wOs
1PA95rWwRRI+VcZVAQIOoEUaMYgML+NVLbCmLpmNmI59zhBLYjWDshe3lv4lcRjY
IHvuE3u/85YN/svvGedcoPoKsQi2kKI/MMHVORf9bnA+EI2Eg5Ssf33LLMC4GWmn
YPWSYXK+or3QlgqgqM2ZaEbeoD/fbDKCpPzHi7n0u7mcus6vlV5xN+fo+HA26YOW
XKoGbcabcEdsaC3mFmt0ia33LF/gs2C+dDfZQPPLeONy3Sb+it4STSvXaL6beyQB
X9F4u87nbIqV1G+4d3ocnwOlDuLFqfZPxK5/PZRmMTdBKpTGd5ExmrLobMUPcz8n
5D+tssteqTL4xQLpeJdMIm8DS5UuvafDFyb12yfoXJnYLkKDW5XQT3gT7q0SZ+tx
bEl74V5SnQz+HXGGet19+Hnj1CD9kvuiviamvAwXZvxQmrx79SRAXAL2iY5udO1m
TGk7ImMfJo9sytD4ujg7QmOhDy5qKc0sOZXx9HbVPZ/uDXK2irl31xDhSKCAFJTU
PyuBhnDzC1R6jnZgZVTDirINLVanHsWr3wSKs1mPAmlvvaBudKSKXt9q9JfFJhn0
A5MkLLmmUna7HTXUy16ERL6Do76oRRhhBOimOf+X9s8ME3ZC48VgBCuiwYrnPr+n
smUM6KM0TqVPdQDNiEtacU++y0hqQHk3n1QDG/N7AqZ3f7Pb3LhJOThDYZwEkoxE
ukvqE99qe1wXOfDGrtPUxnGjVDlHsEUXKa3Rmjxl+mzaIeObSrIekAU1h76rU+g1
MB33wgNuqfVli38GaDrHQ6FbXfgaKRuSPoHOjKCzPnISggcoXFqBMO08ZECEwHRW
k/r1Ve/GbW0wsTShy7yqGnv90bw6WzrwXtMsdOjzn8njiYNwUR5SPU256W9xOAkt
izhkBFzHgZHRSxZ79fwY5WZojmflpb6Yxk4psT7a19h9Siwcm2oWJVf2GkoUpe1l
bYVjMEPBzccHeQNnVgaepJkCuo3tXwmL4x8sr33nEFugPuT96BpykzOkOVFRmaf3
4W7rpaMf4fLlxyesm2HoTLvMDTh+pyMQw20EEse3z7uOCNDncBNOsnP+X1GGzPAI
PxBdJmPf2SS+MPFD+zPObw8fUjYTKUqEOevJpbLlDseFtJM8Iw0Ha8f4hX4lVg7I
AD/VP68QPf7nVyTTdbDVAYsh2KTZdwhimcgO/cdcPvIhWsq8ehAIJ+EmnlPOxDEU
zO3CRNomVbh9hMjy7VDEX2GObMN2CWbUPULUFRlm0d4xwux5hIOgRnFfDfwnPncW
F1N2RoxalNCj+oUE/lzJs+ZQiVUhqIMO55Yg8+nzHi8fHWgYN5pBgjaHOONYOoLV
YZFQUJNV2zzYdknl79wASRd1UDx3Db4kcJi5D6BGZz+EPzeqhTW/uv16yYe7JFxG
VIBvXI/sGRS19JR3NJTRVxmDBYycQjfXx8jN4cXHN7uYmkcCUBcmHeU8KdAhWqcl
tV0nb8S3De+UGQO/Ox5xQOXzTIx3V1dvckj/rV/K1fKibroIs6zeJFs3QxV8S1O2
jRhpkSvc09DcTeD9/zDlqPUr0MiUtf2YED155yDD5Ep43UrYHv6iarPPuEy2Rmth
L/x2qdu64Rlei36pUt2j+dsx9r8IQdnlOov/0GPx16QHeWn5aIqnFhLtTT7GMpTt
fV3P0G9YC8yMOex2tC6W2j9YmTud56+xY6lCXRQ1w7ByCjAAxufRoBLYeuYB8x49
mCb662bJG/pMs5r8PTL9pzSGMKaVFYxApla+CuNsFTcB1edMQcBtXJucuA9hLCOt
tfxOlR7T7O8qAhbOu3c5WCidfi7f+fWquPvW5VAweHcHbaRy5qG6pUJhx1tZj+o8
472wEDCgWUjmux91wX/uLuEeITTLaztX9poY/03g+Ui+XhYidSsVWsswLc5SzhSI
sl8zjvPqgms2lG4xMbefW0EdqzsywY7D3/JN6oPQLRnqzUcJtF8G6Fs8ZlgwVMvs
jimSuMpUMaVoaaCH5h4h7spBgIXyu3cXcqw5CeMPeDdg8vLrbazUDKRqrv9rdmmD
YoaLaf5aAdA+ER2ZdNkgczNxobRzTzYaW5hnPBaKdVYo4xDilNxrxrIUkEoa8EW0
NA2RH5KUQgS2Pze/fndNsUkNztOAViIG0z5HdX1ZEzqVLNlUa5gAvxUD+EqDLL1m
klu23y/TEJY1MvYGLQs1osa9A+LLwmocQjv0RSlQbxhNjPIKPeAZK7Vr6dE31fK+
qtmRQKm87zdqI+y9ah089CkISyzc01VN0SzAlJOffHWs12obTj/OuK9p617pLsEu
uVYyLhO/WSVyiCbhA/QxlpnTADrJzQ01YIgJl6o8Twb+NQ4HDqlY34G8Iuf3qCqU
AeHc1zXjvf+j3u81zJ4bxrdUwd11v6RQ8uu9koVrSB+35aEMeySBSQ83CKSYqDFX
vp3xjI25NK/fSx60TZR6LoNfCtoXAxn2ipyLkeqiCqxCPdw8jRAqB7DcRBF6+SZU
72duHfEcQzfup9ZT62i1fcCSgDtYOKbr0ERz0ZQ9dDKl83+Y+4hQX/4GdvfZMpQk
GD6xsNhCehw9XXqJ/QuTrYNKAlSjai7AmtnXMNHqrww3NsbjZavqmNRGBC355jzD
dKLm/yUgNLcuryw/J6b/Vbgk/DKHuDqagMFcOXSQ1qnwfUoHeECkKsUceK7uxjJM
WA5Oom5ARTcT44+4ViDgjMopajIovqzAu5VoTBgmM0nsfYU8KBFivYRaj6KB7p5j
IWOYX1FLrD1mOHRaJr7OpvWj4BaHeqe7ctUH3QQeAq34l4m01h99ApqYp8S49jJf
+cfMKgIz/CfXH/6DWmJX1WRHdDmRFtYNtlQztW5867KEVKmRjS2LxxLb/zT2Xm+2
HOWldNDbmoo40FAL6KXbTngaRrzAnbZpO9blCLo68HQ6D0lti/xuU/fx35psXh00
AELAzZE0Z0NOTFkTFOZdtbsKDDpsrsp64+VEe8E2Ameyatz8UaksyjgbXWfibu+2
NpZjcWI7aWoDd0RNHUFJPsBcUhGgo+SG8mjpwr8uM/VV3rWm1L1+Tekgk4tGZV0F
FtvN3XN+1A2s2CDPUk6CSdESBMjsOqQs+bnCRF17o5GDI2fAn1GTXShLF7nHdJGg
m0PFpCqRc3pH5ZktSRNSHIsLSA7vlYM6W8loqqhPknBRYOjnLovd2oP+VgDWHWQz
4sF1WYgyDL0/C81m3m4OdHq5bFdscqMQJ4JoCQLOBlvFmfaVAQFohSL5CzD/fG3j
Wv8vBGqlhYQY+t7PIITMSGJES+zmN/4uWgj8iQM0Eco2Q+48ezVXlJF6WZPC0+46
/2eC7nKNFhB8i1Sp9TWFdcDnF2iWA06hy+c4vWyp61oH5NT9C7ZYaZhsBuzQKeVy
FtlhE9Wu5Yw+ivTAPcyn904IFpIi+v0z1/201aHmCESC20JIapbqpTMjBNg9byX9
5/q9jwavdy5V5HOiDUTnJ2/CfzCJ/bk4FNIajqhfm+ZRZR/rMNkMEBmAD0mJgt4+
aygZ3C7+mxx7rFhtj2yEJ1QrIcUD+uuhkd59ulc7oaXpFF1ayE1VRYUrIhqNZFcP
sL6MOwpTGlIaC75z/To+1jt9dajpJtg3K52sl9N6fopp/CPQVpGDheuxcyWDg3Gm
uZCXHW4JUmuqVNvEPjxkt/xdWfX8ZSskYXzpxBfjTt4My89s4nsiBoELGoKjiekf
9l4i3MGOLa/Sk8x0hw3MokKCEkzoH7c0CfWhwALVOSWxYGRGJCpsSpBxB/czcW9t
nJCJMTJ2vKbaBGCDevv9dYF+mFtQYLPqP24+mQvpiEBFyOUNCONX2lBmPlcrhAUe
Z0frRkzk+CQFBJYsvBKyfD2+XxxHFydW1rr6G7gpoB7PL+hR66VaTbgOq4V1L5p4
F4JYKZRHvFPemb52hr287YNh/XXbyurrKr4PoHg86YtCSIjJueAinffVDmZph49F
DV8gZOG7FM4Am6HQzlxHEY2skOwz29AYWe7ZW3vHq06bRFih1oTG4oMojT1m8wQQ
wLJDMrs1DPbDCjWBt4tD+/WrIzs4peVL/y+Aa0WqBS08/SDwcmzOsKUr27aZj6/y
j8ysAmGVYb1XSF63IYL1Suub7YL32LCHgV5Yi85oo5jasn3ZFcD41diD/hO1myuR
e0NQnA1PfzgnRTSiThoxppGwQ2MoAaH7Md7uoSR7xjyJw23jOt7h1ukjyeiSc1wp
sjXFnwjoS2ccJRqbdBTdBDQDKWPa/hgdcC/vdDK9WpKzpU67kFPS+APhHy6zC9X1
DwSWX4RFZUqJ/ZTy69Mad0M19ngGb28wMPkSQh3kYzBSoFF9nEnoCDESagYO9vhF
GTUnBLZhZXd3wO4B9MymCKmdhW0no+6uGzx6B7Yl6Mq84Bi3W8H1nbvJLp8CF477
w0I8myzQvhQ5H53f95KucBOEO9HS90d/z5f/XYbK6FGKygqEb19fWvzS7FfPoVkk
ZEc7HolD8JwMHRHx0rHMYjx64LK0gP/AGJ15k1WDBw+CZEesh6IwSjhJdriiEWtz
y948+X3xq1oTT5XkygQuveaEVGTz2TXGC90akVJ19oJ89sel4PuP0YIMd7P2DYZK
FvWpWRdaexQtWADa5ug0ZwnGBMniDtpxribnSCboxScmFzSs0PajAFohJrnnOviQ
46lrcoYbOuTpwlJHplDxwARDsixueEi9MPJMEV6D2IxH8kS++b+Puz3VDh43Zu67
R1dBHcBKD9zT0VQa9U6OlY8JwXgs1Nml7kKYbJqL1v8rMXLBF9SZv69J9UlMekqR
R6qPjYwv+iYl34sIGIgdK5f/sbX0TgRfbtCM2PT7gofEuAJlJP3DBjwBf+zrGbMb
FNo2qJb3+9z4tLhu0/G57qBcK7rS8EK6aCYRN6EnEbv/qpRzhUvPxE2S1XugweHr
2+XhmCClE5Dm6i0GSKQXiicLqJYFvcSKGRBwUzqmDlMwCbNEzjlpohZb6VaszTb2
QEG9vmHE75iCtA8Z0QsJR4lB6beO0R8ezLLKuKDaXen+jVZo5Yh32hihBeku4ljK
IjWfwLkP3HbhmtOLpcFAdeP/m9NRJRzLV2Pu2v7xMuIGOxXdYG7UQMo6KVw69rQR
xQdBxUC4zsFWN9D9r1VPmkr4swL8SdfUcjYbkdtwPJnGDUP1fFbnPpyqQP71ndXe
RzEgbpl5T0t0/iN6+uf8KMz8Jab78mdCi4z8A+L8Dhn14DTaGMPdJGj/f9wfHhEf
J6RplPmOTH8J4Yee2v/3USeBaz7bHqqMsFG/uXNEZGJ08XEtSqswDDhWp0WRVi9p
uv7wyzX9W8csx8qBfBJQ5mpQvTUNG9Kh9Qo3NVdi+Fyk5u2/Z7E1LTbjjKSBjkJa
DeJwCv2jMVoSn2NBHSyBZ4rcpRLOau5JhFVAFBqdTAt+cvFi2t91v6roLnD2XR3H
rpNAEZEs8XnifYYPYBa+x0ht4SnlUa7hpRE9wtIcZLTIQAgWLem37fe9dgqT5tIu
I5RNxCClzvstzWxb+KKu8zrHJz1OnwG1p/EysbqxnQBmshczHq2cNvVP4nviQD/m
LE49M+6HdzxBYdwtpd0M7bqZizzFCVF7ouR9m4MkjYMIpFwlwjaBdXTio3czaApM
zcKQdg83CY2n2XXZnHvcGDqKWjyen9EySDXXVipARl/PClYdCCVTYmIG80FecxOI
7FoDK6x8YgGyWpgxWL+W+3XOJtKpLgqrxGgOjKqM1nR56tigOUGkc9TQqV+WAvlW
YmTG8XTIczRDGoe/PxyOgywRDwxB0RKIN6DX7WX2CRLNhz36BqtTmb4l++f2uEXv
IeInp7ENnyVCtZqunUz6XNbufJv4qgGsMDTLDeLeJ9IAj8Nft8Q5V2wNza0z3SvO
yS2OaiSTY7ChAbp8faIM0gkzGXY3Pa2hg42OlsnHvvn2Kdq7RUDXL9z24jQwsf2B
1s+NzuCT4g/AIGcHuHenL2iAb0/LIkbge6Y+WLEhxVmjhnGeqiRiLAbkeInxQgXA
27TOLpsy4VQVbLwm3mgJk2AXNDRrEqSMW7ar1gkNA05fWEQOPv3Xtj1uBFG8bX+J
m4+iMlGfqrPf7fqSIjG6kLeoa6ij1deCX7uCLo+PttUhwaEXJfSKYx10ntnWZ792
sSSh3wImCPejANzghXuUL0P5K/GRDiLliABv+vD3RVYy0s9pfb91mXB1j7ZAbLGc
6a/RtsJYBOze2nfijDqWRtBjelXI+4G0ztqM+2Xh14n0xU4SQejnDsLMtM9mxNR7
/u7pRhtIvqA/MGlecxlrhj9vWE/nHwcfaAaQvctWqGWXB940KD/Ami+OXWU6kkX7
ieIKOTDzzyi4MXqXboe4JU6opriHQrSRkQ28HF7UgMvArGhy8xDiFKGFbnsG5JiF
5qLP5oyYlHvaAS8xZ6uMqo4jM7tMYgnFvGZ4CakVS3Mfa109acVMx/zH5WJEFm4Q
KTtXaPqenfma3iNuyxci3qoI4P5YMUIXjFWqdyfvxjRrlkxw4EAr4SIHmyp8jvKN
4HYDMSiHIMLiPLThgHuV0NshkFbySa6qpr9afkUWmXkmyl9nsprz4ceZYGo1eJXX
AeSwRCGAUdevpHEK+84WMLHyf0rkjhq0gbU2KBhNKuVFJrl2RNYbUxjNOobYhH7u
x+fuJPnaEYj1cUS3/a/qbK+LUi36jxkxSRsfwCkJjIlTNO+nAiuq8A5ARAhjF9oD
6/vq0H1jSzlRB8nGOG1r5vCsBSLowzo+2lcftvgntpQiamYzrfsLmDYSK4yECa+6
vYedudvj+2f9T0OPjv2u3dABL4TY7C5GdP1FMgv5PcmpGNwpiz2PLTL7ve+geBQg
yA/QTGdHZbP1bu2WyE/mWeBvzyfD61HgOikeUmL96x3ywhbG8XUuj4aJSHflCQiB
OLv5p8k3dJ6vJNUTiUp5za+dGygNxnMknMTE0rsQE9zoCyS4jTdQynRgBQGXJv5+
l99b28mi3MV1oKEzji3hyboAVEOL2Pf4KEJ/HYRHQvvqXSDotm3bgTah1EQOg/ls
8fcZUGYCzSRt5QdECfdQhmcUZKOejqjzj8P2s9W9QmGyaISb4X+JPrRH7jsvwod8
aCl4kHXU4lyoxr6O0OlHmeKgzaKnfPJY/s8sQM+lrf/qHOABISwPYJWL8GUGVJ7f
G4P23GjsJg3yQ9RYcj04n9HxaRlODK6VsB30EqQ0MugCYp6Ro5X2eIVaYsdVYc36
cdNDeubE/lDQbcGCUQKZ7maJq4gGACYg/9NePAc3TsY2OqyImmfDz4rxLAHYhw5K
y39/gZ4Fj3xAYIj2vkFV7F7XdJw26Az380aRQ5E4g08AXzebieITQ4ZUcnvFLzSR
w9VyMeHYZNOhiybefANQR3ZJdFpPDQWQXbaV1simnIWwQhUqKa9KvCUEkXg6NBn6
nEu3qvOYquUWTMeRtFuEJFWRiwJSvW9syDF4yTHETfovM7fjs44597a+wbjLlx41
41R0CS6q+NH0ZkIaXVJQBHzl33fGUGN0tfkaDZcnxlgeYf29xSDGIS69NcWTOaao
BF0KHL0wKrxm/wEaIMGOIHZoLTZayE5VqU2S8M5KKqR5bDoWi37OtYYqOhx5unwM
Gt0R4S6NrZbpnIJmaHq3rwj1muBaH5SHm6OAMBgJnygYZyGFDqKwGMFZetma1kvy
ULAqLyNPmDnu19vEn7J51s/52fl3a+LA2i//fXi3yKfO3Nq2QpudrCjz63FsxT79
/pLwYI0I6+T2Xt2QaJwmao8HFHd8u6QAukucmVwXkxt3BqYbgLZX5C43t2WQLrjU
FtGk5KkM1YTHgV/I6Xc6748tm2x3m2N9G3VBQjSHeBF+CpEs1V3bTZ0oQo4Iz05A
kVJGAzR32Jv+dGOM5guHD/J4WsshYFyvr9UNFZ2Hsb2XSz0EtOUOLsEzm83jug/j
kCH406kS4CU2X0hfDutZVCMZP7bpvQMI1edFrYmlDijJPANSBPA6GK7kvJsnikmg
wcLQvv2d43sQ1CbJ3KV65k4Jl5LXK0iHxTq4EWPD+qCJHwF+4iDUQUiI8mxG9SBH
QcX5cjjiVKY8s7mBLwmHIqfJ6QtEGSdgS1g5S8HLiv8499sw/D3j/PTHE6yIF9Yo
H1dFtYD1KbgPvv4PrUTYIp6hKl2lqsnt4Ux4xEVSIoapmmoYfgXrdAcrbn9QYIPQ
r60QxkmyAGp2EV89me9F+kdBe675fsWkDDPtAjgDYEAm9rR5V9kkm3aJjsmfPYsf
Yszd/Absx3gNO4cfJmeGuSADZ7Ep7BKJbPRKWpyljk7f4LOprTilG3vRmoVvGi5/
isPOVcuE+LoBRl23Tq8rHnL9pQC8okVG9bsm/ezyTwuCL6L5OH4rMpD2ExGBuKZA
Qf1amRbs4EcQvKnDDNxmEhbKqw5Xg76nFU9HZyKv63EyBU4PdMAWUVra1NktddhW
JNbJPTvYJuGactgTgQevAFcYe90//bqYJLidu59T1Cr54n4AEuGsZ9uQ20jXZCHX
fRAmTGtAC7R7agnJoXHRJWzrvE4XfcbbOXS7uqUqoBOCZ2qXDYwf01QFsmQhNOVG
coLwou/IePrcWA2yiptHus8qH03q0XKMzXLMy2uamp83/jbd00/0p5GSjsSabR7v
WPn5DiLz2yPU4Bb0OQlu5iz9Us1vjxMUWfqpJ217nkJCsUICkMOC4PhUCHb3JqYO
4VikHWoxV0QLNfxO/0bxeXAiCJ1yj3JdNCfsLQpgNSuhGiYozvcd3OJmorITzJfX
FfijK6xZq08etvy+nk+jtdjwVsBVZ+jJKk8lj6/d7m+MI2yJjLGKZkeOTvNKribN
1hPVmQfQV7oPU01Kc31OTFbEBdGqpUyUS08ZXjgaH4/CFnNaqdLZZi4gH6po3wQI
P4Nz7sINhVwwLU9kQKZZ808u9tdzu46U5ZfLNs7Jud4r15a9Ia8AG/0g/cclmH2T
bICnliRq7IO40wKN7A78kgkql3zGG7qsVWnY55+NYH6sb+IusnZfowsHYQva42Pg
x9/dabz8Smf9BNAsiA3cyIPLc+J/XSgYWzs/YrwqbTKNTdfBCvnava3P68ilO1nh
7q3T6gIxMb8WCHlKgeGoF6XnZWgo5Y9jS9pFYrVD23KzoWro1U36UINdQ7UnRTMg
HaP9fyinH6PVo5Wu9P4p2V5qgFyPkR4i7pFyipaIc61BHyh50zYBBpsme6Q7R4T+
PL4bNZ2wRInkVtSDPJFUYjOcDmsHlSO18HTJ7fdMYFGkrrGWXIilJr1PRF5S1wsV
WAJu/IGuJPF8+RpVHUYgI7ZRlS8uZlG6koLBmvZJCTE1gz388rfZfQovxkGMu42p
ZryWQjTVvEg3u8OxynrFg4ArLwE9G0/7B7hRlTI/QvolfuJX9Ise3AaMYvFImckP
vMYUUPnnnrzkbFumXAkZfGZP3sxxpszQnDklfQeXikqBFSyXonKh4ebgZFrztJPa
X9RCXaXCfeehXr1F2KRjvWYaX/FhFWc60G02gRg5B7Tl11GsTSPDYAltnzWnih++
f0MwHlkSVt8WjtiO96n1wk4cPtuULEqHXjhd38PwgaM3JIbvObF7L1KcknwSuL3w
tyyJzV5ynR1IKl+45uZ4ebMLG1xPpZ7oIzaX7/3FoQM6JoDlqrHfl+k+iv5c+zKb
fMAlyMGAWpK4wy2XEjvB/ncUw9WdU598SsNtVLOhpeHh1hO2xm1UHntt65FH8XWf
7+27ftszDqoxgLQbkqOPoRmtsYvAKvFJamIthWYvqQL3TLG2vbDE5+TOGZ3h4ePt
+TqXPibCX5+0V/e6RY4sBagMRyvOMTlO+EsyspBO1h3Yba5zW1UTYlonMtbse5oJ
7Wym73drs0kdCIAYTWXhtyFvKs6FeY2jHHQq/hv/54TC8UhWTT/7aP8woWE1O+SW
zieVW7XLoWowSShzwbqX/jWYkto0b/ni3SiVdn+3RYu6HfztIa8gh7d1+NV8Mksc
fISSLPBoYXZHWs3amIDBWH93cMwlvedhUwb4zzDlFigcHMaRK0dln5lYQ9g3Iu16
QhNYzhRu62uJ9sAX3NKfGXcLxwoxcnPk9QPF/olhxl9D5rU9ZI5P6S1tksGdw3Sm
4t9Q0aWoXNsdnDMOansPYet/mzg/eQsoixYQD+Uvyd+nkyDGTiVz6RnIPV9dSCCn
7bAS89qhbFwIrwikt+RtEAy2xd1UQUtRJTWh5YGQrQrgD+mQLE5Nycr5Hi2QeiaX
Fx7JBKEEAurJ0Zew4T7IAYJbEm3myZ9QWepDPTXmvVBJ8hVVYRcquhHNvNURM3AD
MrQvYwyUoVRxHVCE2juBWO5zNeZL0MbFki5GV2WoRhaenFm/OZKwnYXZloaVNw+m
l+QP/SOZ8iAoBZxn465JH5QSqwEC0BM0DzxAE95rQXyCfVjZXkxjSFB9Czv3VPEE
QxCkwpQYKu7D0sQp7/moPru88ETUltGGq8THbRkNGPCDD0gHGPcLtKala2u/UD/b
9ZHhquAC5OQPJqslnxrMgRwEbkPVmJqREzoxunEEegcuV2utZhdUEA6ovB/orgxx
PKenCJH8Oj98jsXtc7XuTg3J/aga4hYi3QcVbmxy0IBTXs4M1WGwxIzZZoVMAiIZ
mu3F8Yxou/wY2rttS/3eeq04xdFuAzlSdDpx4OtBtpwBNU6RtBoIL2WNwNefcJIB
5eOJJdOuBIGy3/0dQkrfPB/ghAFPriIK7PapAoKoFNKCi2sOxPjMUAww9/rReoTV
C9iWA8mkDTYK3FRf2nFBBw4fYDa3LBaWyAN6EkadIc5ZUBNddDyFSuAlr1Cxr60u
fPdBWhK1/ymgZfGaYhvOPfys0uu1UqAkzYEesoH9XbpnXU5fqvUny3Gdf0VTWTXJ
vqwgvdMVpXalSC5YZko6C4WdOfPB1uYm4KitJmGp/2kwxwtmsKsqzfV+GekhQ5Ph
Fc1fGP60a6TdF2U4gpt/uz+l4JP2xSKY+Y1ydSD6VkoM5JhgdgB+O+ypm978C2zN
6i3PHkdk9MIAvrWGRoCquuWjyk46lcovYEw1GmwxV/Se0YMdlXwBsBuRO7kfH1Hv
Sl/mUTI01kf0qbqXP7e8cux9tuHAU1p29g3HtxXOugyuLyZCFtvRT3qx+zFxn23e
rbZBz1F7gt7f+ix4xaSXTgg6WvTnCQ8Vl2ctnYDfNhIVYUD04ChGFacRE8jsOSlq
OWOslEfA8upuhEolmmWvx5kB8adT488b0OmprfuUfRfPwjb95QBLEIKjqzEPkEl6
W+XjZwjBz2qVpEMByBwm6KetbyONLKsbRiXzQ5yq296av9IqzMxOAI6oBG+frhiS
QBfrnT2eXR6vUc9+ZrcX7cp6DYDlcNSk7/Fkus7j/Hy/tMoNFjSMaDhePzalECZd
nkAwbYnvqS9G20mVDKseY0hSYCoTXpuYBZHwpf6thzZ/WeJcwQhYE87gml89Tc31
0WL/hodVJ8981FJ6Qa4a8gAnsp1W70PRC0jL3mk4ezzwQ5em8trGOK+Y688EXxbG
id0l9fSkSrcrbWfkb7LPe6t3P/SqAnqTWw/j8TJ/KcUVq3D2Qr6KGaV7c7T6hD5N
+pUvJuq629E/Is413SuAOJENtCy/0kTGgplB0+JLnMSLKfFeXIoEy5ZIYQMiAYSv
yxrJFY3tl/7mmCBfA40Mkr3Lg9bZk7AMpvTl24nR9AK3PwcB8DSpkvN8syfhZD+2
Fuu8F7+hFmTL5KPCflO1SEmn2zRsZZuo2nWK10BK6yH9wO4SdXto8bMbmEowvvUh
38+MzfOHKjJczOhnALqm/+4PtavkDoxXVGECIssWniL1mdfHFNbF1OL6d+mX7DTo
zq7WkT4xpzjl66sqm14FSQXn/rWaejYwkfEbsz70ExkeRYgZZvlxlXuO7KRq6Snk
xlrsnOrCC1V18/vZbO/+f4600/Qai3hLpSNBIGDAcOHU2QHV7SQwiA5b73US6eUf
dPHASIyA7zeRhxmZEty/J8X5nYHcTohOAqbUTu59+FwnZTu8zE/vIuGHQaRwmBOQ
DpWoi8x0F5tXmx09Lkq0SDuP243MhYfYR2xflCg1FATf5DLrj76MVVNBjwbi3B2b
yWfR1VjeYV2nKhbv26qDypzTIw731Pphz2e+r7vaIxyorgnOeduh44WEioIL0nIB
r2iEFL9iXLyEGdnRAcFKvweWDc2OkXg5/I/RgRLb2zaDQOyLmRaZ1xz5B6/Iy0x2
0wwDXRBoX9GBQi4JfMwozdxK7mMyD5ow+e8q4ERPYcV679e2hLidJT/rXNGgeohO
sORx1pXTBsFT3Ojc5gwOnEY5Evdhd89Z0ZVl5EtUr6vCqRHJ4gqh07ZiezmCot49
OC7gElo/CoCDAcYdMiyuAIlVKfeoLu6TNZqLO6sE0pExbstERTMo63BWhzP3Mgvs
FW5+538l0D/NdFr50QojHF+MRLyfrlVvlxVtQUwjBh9uX2gBNVYdXOsS+tjiG9JQ
ywwBkfY5rFLc6TTGEIM46WpgmpDMBajSy9v+HojreMvKg47XXciGb8fzznlnK2aB
NZ5FA2j0Dh68U82y//VUGIyeqVMKruSe/IvG81WL8T4hSkRek/VOv9eIB68ZGrMv
SbqAQmgkO5PKDsD7MBocfZAuFdID1qf85HKo3WSgXj4TEjLNWumR/pdhZ2sgfDyI
vdvfpvrWYrrN34hp6QIvR2t0Av8VTCf3lP8sXP+5c1JrwTs8s4t/tyEAvQN3pxer
YF34JHWv45FmkLBNSuarZXDbF/AgzJsF1qm+/Ke6gR+pP/cLMHU182DA3zvsE0pU
89iOWTdw0VVdcm8kv3jBjkNAq6ih4dCfLbDfbfRhjPdZ0x0Vwzy0SPBpDpxB88BH
tQkv/rHbTtZeet18E6rNl6NMa/4SrhWKj5JU1gwMQNDI/djObBunLVph7OdUIMsH
Bgy0iBn65uLMUUDf5Y4/68BEwcM+BX1uCIwh9GkiMP0H0PQ7LUxN8xecN2r3tzCo
JmqfgzJLIwIfkf5hVswSSx2m1jYksxw+gWPB46Bf+QTJZqWoyYglgsIQNwn+DLg7
fO1k11FMJYKxIit+7hs2jYQm91I1s7WgzVEjY7HTlbm0yOApGaARxncEM3O4ki2i
37itkTkcQlKfS/tnTosmfaRkaS+1CesHuzsv7zgnM/4kysX9cru7k+DcxIUh8xU8
KzWefCIB662JYFDG372RMOKmJspHNXF2zHx/WngqfCIgTAa1fMVCGE4bp/TEb7fA
LEPjF7v77COLoH1DR+6PNBv4Gro6Tf/QWWVHuGI8CEoUxAy5OphNYplwIxvvXv+8
66xZkuktkUyaHNAn7cl+yxivT2GoheIoW5XZ0Y8+V4f+RrHzVTRVj1XDD1kC5pBA
1EbBpwlgtMWUElr3BF9fYeX9bbeXmwfj2GmQTpMGx5X8ojnQJcRssdJ6A8V3qd0P
BH6GPS6aNjkbuxY5p+DWg/mHaZETzT12DyhpnKzAMYNw+ZMlHwZLd1PS8gXsdukK
+JDawYIpjRjqP+du2uiUbzQGC9h19KPTwamgRYske+Yvz1jzv9M9a6m6omJ2s5u4
gkkjn9PHXehVteqGEM14nxFE2+Ogs8UK0SB4ZvoYobcsQlhNpn9m7Qzh57Mr5vYe
fosYLY4uYDKI1JNuJ7CWTenFTuKF21i4kCf8TdwaZt3hW93tZs79Z3R5XF02Cd5v
M2Ced58KgblBCSRIpcwuzrKzaT/BWA1jhfVBXC0qRzgj6QTbHXCyIGVD2NICtlcy
VAFSjKy8VsAFXaFe3ckqKaTRvq29YhnrdAJISofZT6+fRTjCphJ20fL0dOfx9slC
ypixV4OgsUY1NLHjYuzD9Xpv/UJE1a1c7NojbO8xjiLt4Tm/G2VYthvpWCd1Wz6x
GMLdTRoAJewpdLX2P8fw0Y36vge5t05XxFc5kO78esxNEOasbrme/ca1My1ET99r
JIDy/o+XvyPVxcYknLCg95UNO1/ETW2BfcZZbpvMXkRqpTQ1au1TrzrXqu/6NYyd
PqBZ9Mc5rz+skPQP2hUdZ+Y0kYLUuZvS2ZLFniAZWP+/MFwZpgijOwMZpyHybAxJ
lIOoOSyKW8JoU8JvEc+mgmndfntM0hBaqNmdcIse7ef3G/aOyOhCh820oohDOfX0
V6Di32NLdmdaISQARAn3vt4sd+oXIxUcFRjht2ahgSGfVjgi97oQPl7kPqGg4yas
LVV7J3x/6oZyesQLkQJ+0Xh+a+j3VLrUzprSlm5loz7xMbUqlGGraf5FJUe7IwFc
/7cXRMKRAOOKNyc347JwTXHpd5PEmsUrs5pXGt+6ffvJLrsVl5sJB0ks7TVQ/HoW
XfcBlE73BSXrV9CkU8JuJc1egDJ71e1/NbtxJY7QNHvM8MkoHqk1qeqkSJmxzoMY
azaKss6I3n/CZUHVQHapOgz2KNKNn/5E7HGb9VBAXKb+Y53UdbWzlJPvcFn15v0o
VbEKSW33EfklZNPINHQoRBvQFPCuLFF349DSXMj7jnmYs/VfzthGxRY2NA148ZG5
qDwaleIMaapOBW4T1ugvHkOTHGP1JtTXw+i8qa4tDyU58Wa9mOUjRvnwo9FK9Lok
ob1s3YZUvlhebj5nBM38crhZSEUS2zSRabxswV5bFYjBNsF34BlBqLfGtRDsvBuX
uX6TVd0CdpeJ2ctNOfwTx5+opvC4rekLC3F8S5KlL8KJJe8JAzPaoFZzGTCXgNO7
azR4hmkaDV3hpOG20YmtoyJW6jwp9J4dBJu56/QiaNdubmeTepVNFzTLtAOSnZKJ
UE8cKthWMe7RxxfDK+wlkn/yWfrWnsQTEynTzDEhuj+IgRe9lUMGFdHaEWIvnTUF
8Y7yYLBkn9hkDVfI9bIZJ/yUMmf3tRC8KlGgtsBH5HsrE415qVmFDrpuoyv9MYDw
Sy69i5ONOd84+1aCCVEXouKx3tVh9AA6I6JA8eYnGuZGIinhtH+oI4YydX1j8LX7
4ZSdnacRU5oSEPF1Bf/IKRXecVSMR/88X1iSnE88seI2FXGjr69SCBL3tUyfUD4Q
qBFb1sTPTFFgZRA2kXKEHitq63tcr/GkjpBw9PLaDpRgt/CLGUOV1xNA5Z1IA/cx
XXiBPiv+E/Gw/PNKpZoGzv8X/YH+h4igOdatXY5QAE3moosVAUFl9h4QbOCfANLZ
gqfSVj2zxULm1HhB+Zh4H0COzVWJsZne0mznKuRzxrwBRn2WXEoUSccJ7580O/KW
WT8JFSoH55QeHP5kZ1tgjEhUFElplZJcv75q5PUo8qZeDyMGLd0hOcZTH7GA/p6u
EKtoWOyRPggV4b/tlzSew/9aa0syjH+wCDeXEcx/613avwhIAVPGaCbnUg3PNiEe
s3empGAFQmmVdwZCygFf2NXl6gvS08Ls5EDwHgBsXGRAmLVZU4UfR9hN6rZDEuq0
FxrID5WbMTyDjdSNTCZhNjanqCLr0+hIJahh20dXf3Jt0c67rVVXDB7YTsGQpQNc
D6gABEuAmfM3bh/gxU0lvRp69tTeFvQnuv9J9d+vk4C/3/b9oRAF393bsHNAInNO
7ItvBVdN5eTTdKiuASf88pMAAUYZ8SryxNsRgsT/rXA1/6HhjiZrpUXA53iYccKl
kHxk2xziyS6wozdQW6IBKRVe4NQs+cdkarqQp/GpZF5c6ACUHksVEy3NCpcXDBqB
wwucdLPksV9e+Hkecnq+isD6xcJvwv7wITnIuYWeq4s1g/rn3dj9tc67Jy6iejWZ
sIM4muXeUQd/YA7ZKdvNoHwcvsbtC+aQS8bJ7s8I5xyA/HXN9HInSRj8NmK+1gz9
A7nX3sDFmT7Pp92n4tw7wnPS5Wj4GhcxmOUbphxwLGKS69z/XXL+jBUjfHPl/ySD
ijX/albytguCW8xpELeW4o/+aha5dRrIffnCiauWzFSihwMov97sZYLrG+iwKoFv
KR4VyFpPNJwyY3qjRzOlMJYp3KpQBzKzkbdBx/l9jBW00TmbkXhMTTacnCTjkn7v
LP5tIPVnf85SbNAsHldl0peIz9l0uiqnKjv+l4vF3DWhg3/a3HkvRplGawC8Isyc
MAvAlSUzwAbGWSk7Kv2qi7y1ycOgiorM0Qra4T+kGkdKFN6euC9UXbZuVTZhOviN
+nBfXAsm4+xqBzKk5Y9YjRoUYRNQHB26ezgKVsa8t/lckPpxbah1WGuZjk9/Tf5B
WFpIWimzCtCTRWcEifnpvXCgWNI1l0jIp0IN5RAd9dr3HP/cAk9dVvgTNGDVOapK
mxyoCh62YEL5S8QVTGHBZRYTnuCougX0N+CNJ/6PZrn3vqMqGuvgSHC3rBvxgFvA
0EckQYEtq1//flDbPnBVsm7VWh3uyXTcQgbM7u4MPJX+o4KQDVs5xt2/Zj06Kkmu
uimINL3uhCRNEQFehDOgqOEFx4OwQVCS/IINU59bgCuV0XQBwbdqtCv077H30yvX
/A+c7zmSm+G22C+4/SnRQUFitIxC3NRGdOY/ILj/KlkS9N5+J1uL6M8/0ArgCo4d
1iO3dOQFVHT2aeBT0UlwIBn7yT2zLWuORmXB1uGiBdedidqSto0U+ELN0fJ1cznG
oIHOc10mowlwDiHhJEIFPZx0W2JReLO9kDZb+Qls76dl1z4wg3CYGmhEVY6ffcRx
tyboj+CG1KSN5eyjm1DpP/ggCQ4mAgqxhfqWkkzyyycAW4j1QXGSaC9y2UvpLsst
TkCZ8xxHZJyLJOfIyAL2ZgFLKWY4VErv132wL/McTtvo3VBXzCWFibOUwyiDy4vR
vb6B9VgPac1SrwTeBGhyOLqPOBv/Ea9ufdgP81c9bQNDv1dlFtSaRYQPjLyEnzve
MFLgJVcS7nVfC1o0hzGkVeEspKrYK3V7qs7KXjQ44yxNwBb+TEM6pohOCGlO+MFJ
inxA2nveLdtY7GIMDbFz8L2Wrg4AIDrgUS8v8uVqhH9ptI2iVIZ6WNCFRyAtZEoF
pDh2WUmMZSNZS6jBzA61duJCvgQsnFxEIKNPt1Aaqt6QjJ+yyj3/5ADUzLgiPKzN
rq9HlCSTMcBnN3DKdwhpxURjXH1JB4qctndx08Cvxe8SSnRBaCe8lPr5qAH8E+r0
9KRyq/128gItNFYytedAWWU5RnvBxYv73DQJLd8OiTrY6vmTM4JN0/g9AGLGKClK
2vpLa/xUoReU06SrBIvHMnhYf+PIpibiWZpHoajsW3hc+m3FhJ3F3wZTfYol/iGi
V2ZiMRhNds8RhBHd+HD1yLOILVHMf6N5QtvHrHYTTWpmioLz4zOXO8IEuGjuQuhL
BjH65qqijD8/z8hXJ3Y/Z6r8p0F3gZRjy5xxXRwhvIju9JPIk5oNrQBZeVUxW7ux
tt1M+pSR1z2NGy5UfvEBHmlIFaVdMxBX2po2ae6WNeCkXd98Vf1Vpis3mq4JJVgG
V6DPVRfVq/5RvUpLstVWl9QsFnzZny3CVskzfeo6pbIqEJ/j9klLUQUfwF43yqqf
xvsyfU3zFVzLDDa2uBAEmNzOwbQaao2E+V7Ybvwf1OhV2GgOi/tLGCwPkG3f8e8b
NceG0a7C3KxSS+f8pBwn0gqsB88eSFM0YnuxLK4h1RzO38cVr9nmZbbFlk7LEtxB
VtYWH3Twkgl+EJ/CDJNxl4RSf0mupngPFDInzTKId8y0J1Qw7hss/GLd5VW9MIkK
LHGP5w4hMt+2Z+KIYMWMLyCkINxfcMJhREPW2XxpnMjctiFI4z6BWg0OidHrhkMw
+yUnOf72e00/qA0jyWkJoYfrL3+qpnEYfovLqFNsfcGZpMGHDE6sNPmoEWZscMS8
H6PkCihc/MBs5lXSBRp3Qa5xXRbtd8TkBm2ynC+jcSrnaCbUVWhi+7bQaTNGBrd8
3kv3YEFVnMOJjF2nsANw3MxIGo9tWET1L2KvicJW2Ev8OEStdMztSVDemcE6c05Q
V9wom5O19Q09gX9dhiYLM9KtOgVWO6qA1MX44Ix6pxspPWPuvBaVBjraAwy0feC2
eU1FVMUshe7JEpVCVDrIb4BGe0b8p6Hc1Cc5MClj1kbYoLK8304MgdnTjO5YE80h
P4ndrnwG9BUZ0AKVjv+U6yCMQM+DRlYiji+pY+AW7XfFRhY97YJ1+Qzz5u07vw4l
HhqGsp6ls5FJd++ClFoRFDjPgoW5z7yh1hLYfay4IM75lcb+4+88152utVNiSiYt
EDB0vMYW+A9/osdJZ8/AyybcThW2l3jqYEsOY2e90pLD20NrXG/b57+KYAMNc0r+
9dPwq/VCROxJmep5IgzurOQX3UyqGc9GlYRpxvdbbIbtq3bsmyLG99Jtw9lHc1qq
F7kQIP1isekRZAODjGJhtk6ohRG4BdJzV2YvQvSaULhSI3d3/aAxm98uJSBCqImC
wdF/Ldxm6yl1iGnynEzT/UGVectfHT3KgWr0lZR5AvaraAMmCYs2uR9ViIh595+Y
oRzX3OZuNexuruAlwelBxG7+o70ZYGmh9GOquIien2kQBtffX21A0kQdjk0oUwW/
O16ehPuyj/iLSKZRMj+G7wvwQNvmTXJHTPQu0uvT7NB8OSWDZb/D58R307QnfEmq
DzOLEi5WbCk2fvD5PpUibizXmNbMPAo17blGFaqHnJFaHSWpz8BOZyIipYTTcV+f
0PQjxHNMZMIBMY/ETI1UVOHPGGgrSCW1qIlqq/H0h1YGeLc3BY1Zp45HjD4xShov
J4rJ6VCuarjFCop6h+UcoMqMH4DTvQk3sf182GqE3zbPWTBmhjoRasiXDwMAeD50
sgnPONZ6aUWbboPBz32zUqiWpPll6ed5pbEpydcb0QnNeOT9Q0QD7Zb5cz5ta/n4
l2sOPqxuQsw9gtPMddPWo9pslfBNCs7GPLrFMfEwkFnCXEgl9Jz9iI4uOPQQ1X5f
277QQad9Ir+FKGnKRfD4/nmiJ0Q2f7wMXy6bMttlRHeGwjkucZjC7bzWz3mMmL+2
IfaSfudTkJQxAmkQBVkPwVjDAHKe4EVBw5Vd9zOh92fyWcY8/uM8RqxDXB2W/kiE
ET3dis0PAR1rkc/werzjpg1+e6d80WlsTPJuyOnzSY/TQ2tDoC6au/0LHWLPFjsL
JEniGHsKSD/s4QBHnDEJgCSG6E44vbhSlAmfzjTm2NfidRCLM7oZajZfV3cVP1+1
ZJJCPLh2vpK5/0cDZOUbjbVtD0CBOkNsoV4ZjON36Ak4GZouUG64KGkMtKlvjr0G
cr7D4M0Wm1ZqDTlCHuBEaXcVPYXNWxzRvGqB94UsuOTUGPVmhKA/CsRScLyFW+H6
LEtzE7D2WIzwTAxTvuo9CAxzQS2rHiKTu0m0a+7fj6Jz5PkUMqbFJBsiH+Wdf/iK
xeERHeA6xZEni5JnTmDJxdfoSkMCrrnF4oy/8cdLHeC+lqjs08YeCW2cUn6WI7/j
CG3C6X+GXjHnSdgT3XOiY/jIwogJcIGkVeCx9vhfQkctOo0mdU7MXcniZonkdiFL
3N8oSErVd2OsGN30q5jkJ5mN3AOT8VZluju9l3eKEpf9tdM2UwttWBLgDMw5T/MF
IP02u89TIvd4WWgJtBCGCG9CqrU63feXAik9zqCeDSOb3SbHzIWUHLKZHpvpBD6k
UQykIMBZOIeuzDFpkHzP8ovkAHULdjGl6TW6mwCrUowPiTUGxAGk82N8B5ZF1y3B
VA6wl+LZ5TxMzmoFuEQJyaVgR3BH5pvcsga6q9ynDsXcaV5fMPCicUd9MgHFJUze
T6pWTTindLrX/lj0badJ9JcmPme6vmAJUiBRDZS1AaHPVVhtcglTKw6Zgq8l8Q29
2xd0Nufs9EUqiaL9pqhVXHvj+rxYQd/ARC3ElS0beKcLABWhK/HcAfB9pEvxi0na
P2zr2C/M312/lJYnhY/2AP4XTf+BZImJXMZu9tAMueOT23mygLjipzJARXkvd41l
L6pn56MAJ0I4cLLP37mU94MnblMjJybh3Gxel6xTSU8noIJLD9KOapOOMihOjwU9
P0lRHL1+B577slTb761Yrb3PjMWUBuz/foFKigS4hY+T63p+kd8RgkTiWhk5rQ61
ja8cEwhtlo6ZKrL/IZ/i4HEHyq6xdAWhR1pr73NlnTOrof6NCzFrl5LLrlvDOzaE
m0HEjvci0zTNCFzy+S6pV96QRWwnOHdf5aS3AJEL9GmpGyINBrveZxCYtQV/aKRS
MAvpX3CDB3NBpFN/McZNdYy2RqfvUq02jfCEY+WWxU11KKPJr3GpuSaM45urD9hv
5GuG4Xk/7BSO0qw28/sDel0ZWaDIpc7Mc+TwYanooAbCIPmgOYlcgNl75m+q8qUZ
ZdxjyRYaceQvihL/j+76o69vFE4EhgikmzV0wtATpiZ47mlcSxES/er2SYTYnlCp
IpvVIsuVmhsgEVqJwyKqISshPpSCUyp5YIHwo17ZAig7kHeYGS9ufc9o6E7OFncc
j0EvPNu9E/1o/BOqN26hQ00Woz9Fv22MLFFO8x0MR0+p8AT/P5MOA4GqrlSReSNe
y3oRPnruPf7AGfozqY+iTqC4E/HljRNP+7OXU4LdT8OZXacNAGJCnIDXTqjX7ZhV
L3TW+59/TcTok6/JNNB7BhF28p4ehcrZT9VvSC1iAVSR8B7aAUaIw2C01J21yTCd
bP/h4fINLMhsJD97SFD+PoN0ZQmYc8yf0iJREKsFa5Dx8aNAG9un+M+IuUznsRSk
YJHO3Ef1f9Wz0pcKjvpGCFs9fhxNSfXxfSdhujKv+EURYXsYj3n27TrsEc+H5U+1
Fwz5JkU6MTbVGWA5C7Qys4uRQ3VjgOUvpP3M8f4E3rl5IBaPYm1iUxktiZYE9kZh
WOepnhX7uuw+TGW/TuPZP+XqrSPIr5dUuwbjZlq2XqTzhH+1c9pwudppP3FzCb1T
PiEuxuHV0K2D4JEKmKvixu3etPyCAJT4yimGdzIKEyBHmi6S+rutYBUk4PuvbI5p
2+DLESq//J86el69PS2ECbYfNISpFlj6/kJ+VuxCZckxb0vJz+0FQGh4isqz8f2S
gSvvpk+vdBfbEgDcu8E8wOMjS8du+VlSlBZbvOUkbxFC9ytdFSzHQQ4onBB/SIQG
KQUUF9bIAtKDDoXcwscOohbu1WJds8Pzwbed+CkFO66KrSeu8hGZlHAqfj6BUHiP
557q0Lj1aiJbkyP3tCATaYXAY1D9vqe486KbXZIAgNnCzJA/ksCWH9EhdyLZ3ZaS
EZgtd095sGFyNywCv1l8202SJDf/Yx+fCkmR1fmE+49lsQIJKU3zNfsY3ULvNxWB
yL6lVJCuRVOpCTG12a4OGIxCChAXh6fAjMZnaYAm7oGw+0jWe8g/2CS88xw+/LLq
lBPk+rsHapXHgDIO6sbT3kqCIKXG1Toi4DXuMLCnrLdo+YWB1Rek68TORfSafgzY
3eFA+U1yl01nIdkKKFTU6HOMn9C2w+ANITOtQBSs/6xw3cUn4CW5h2i5l0cMJo9s
Nz9Rw4tfPMZtaw15sBcqG6E2bl9oDhaOcncQhuphIu4axYCBQ42Q8MW2PG4Xzkcm
GrY9aU5HDafNeARnS83NrBbhQTs+OZkQI1lJCd6sSQyZqgdaPvkoRGCoM8YdUCch
txwpB1rMfhKYY/sk1IeEjpKsCYHeeJ47DIM+gEcCS2Qk8nvngxVZlzpXuo14f3BL
UkspRQ8doGk4w2NmiaLZofJhnzx1ePE82ETOKxZVoHILi/vt8ZmnCb/0iyQ/bBa0
589MwAdS8/8dkxXGqpwhsWw17eomiQNBEvy0nKhsnkDEjChCC4Nats9AgA/2yUp3
chbdICnfcrbnbWPdr11+PkwTmI3589/qfr0q1Jmt9o8lhr3yp4Yf7BLD3wDTjxQ6
guqv5ZgQxz3HzlZQ7ptBqvXQBh8riZAGxJQBs7+j/kXF0M05LPhlcUUlPAlbTzEu
C8hawXr8xAlBYfH6wVndrxZrTnOmCYnjE6kVhmXw98w/dH8AFN3Re1h1QpZfCrpf
Mqbb/fLMpwYAlCaKEsEf46l647OhR0qPqJbZq0vndRP18XrOuZQO0elYD20tiIHD
wBxlbtnnNFhhc3tFmZ8zGE59Zk5trkl6T4CjSKI/bubj5u7BHGIEDdvfcnBKz7Vv
agNzEHftduvBGgEyJp8OqF2GQktzn2NfZW40KsbV0q+W9Jv/SLks1Jem8yEtemw3
j3Ng9tSaWEw10yGj8bAxkFYlu29GnmzC20WXe7SKjIhpmVs6+L67svJXm2QD4xRc
9yLtg35Axt+9m4HC1jjA6JuGlTLVkfY5LDEQcJSCirWe56/g9UChX16GlgeZNw1g
fv/M8w1QgtXHuFQ4QxK2ze+R+HtzhRdI8tOVM3s2pjgY3XxfG9QhO564LaQwZknn
jl28jTv65/FNvxQI5MrJhu5ISn9vOiA5ezxCDma4U11m/jtNoZlkUhiLNXw+i2VH
lhHmTR1yTNAca3WE60gSLydZKYP/8+HbRpi1ppAu1tkkzbA2pdzaarvKfS/UQwEI
K/KOMR6448JNTZveYLMJtCq71BS1y7R7VK84vYQ0eR3psF+wFs4/eaNeoGYdLqe2
wetZyWVPHO2rfKx8obpq7dbW6pEvWoMxeWYh4hL0saU9Bxrz7Qk5GJ1HTxVhLRVQ
L7q/oLBw6vDs2OZGodmz27ShBW9YDswjAdpawn4YNuJ/J2fLL45FULFD92puqmxR
7M9+JiN5wEfd+oCWtkNjYAOp2NErRLhz+jJKeDzPcT/HqWtPWYaYuDtQOwr6c/wH
vgt/i4071h+0WtFzgURfjgYyqucH1NmRpknUW3fB3kOyrY0NmYloIWbb3GJH+G4q
v1R7kwhjzkrc7EVDEMJ9PJ1bMtwPc/EkpkcEkBE4nkYcbyJ+GEka+ZHN2J4Q5BHh
qmIMZ9+OnIHQBkoNvS3ej1a3qGordP3c2mH7kEysL1PXtuOkRP4AXin0bkyaS3LX
G5DkpS2cuLg2g8WKCsRJ+JcKRJ5MPIPU8tIk5aJPuQUUXbPxPGD8NEe7PKxjuRGP
PekD6AjUJhRTHtimQe9yAZ4zgK/dv8bLlRK+LJHxwgiYKPl8pbFaMaZQcHPlVMbf
WpJKTROF6PxBLOhxsReKFj/I3XG7SEj13PE/1pbpImO4S8hkjt3+BMqf6MzZh+9i
Xb0ooJZWdfrgNHayS7zplkkoxAw49EgZtE1VWFniOBPGTy9gzmrzWH8LCvIgylIc
Qyc6Wg9knICLcrk7f5ZP9MRR9Y17pN7ZchGZtbFtMLRpJ6/24KH0AZYaERUHM3ZJ
4udabJq2RyKNjRjuao79NbBrEb7AozKW0fZG6KomnYObhmc+JSd22UPJNTAHo+t0
SrMKFEwkmOBQbtzhbaFib2Q6Gmo1C8gN80/+eFEodLruy3B78jO/tmUuWZLFWrev
zY1LFGE/ND/T3AJs2O5mPw9RmTWQr3m70eLwsRoESFxdm6dRR/GXwDe99ISzN0IU
tkLMLE0Agzxxm9zKxcynOiFHBmZ5H8UeTCisBOwGkJeF8o0jDucYT8TgObTM1h9C
nlLS1y+UNnbULxoFosIV99pUvVpTholaehyrtPB2gx2kEjj/NSkexr1eW7/CBUHh
lV1mSHk1hqc3W25oXo8kPYnqBdzdPilEZdMA7Cj/ZjGapBnzLG5e8sFCyJUrm01P
ugV+vZNnF9b5nE93S/zolfpxTBbwzhYiAacgm3W7b2N17Tit7TpXhKUnaqAZatp+
tOqWfxK+VjMSpUmhVnAdlp4P0jaWMgbM6NLrNLZHe68bSKJ50LPS0J4SWtknc0og
q85wFDk/uKRjDiHTKt+jI9d/TCqzg0ocJeF1l/UwRVz+Yk2ZWYxUkXvyR9meSlq2
8oALqYaKwECI0z+Dp7d4kwQYqQolMpIwSZc8Rw4S6tqSiZVPeNwu8T2KYeRCqyh1
VaIWC49BdMYWbr0BGsjkrmJgykuKAqVFZ3C5CllOZvTOdqlYtpDq5MLIIZOFYIVV
Ez0/lq688nlYDarguEJ5v7cFnFDPYx/BIfiK5/7JFy8sw94bXlYb/p8GtBvr1wbX
F9GXKUQPk9sycoBPCkol4evia6iR+xBaBQivQpgDBJ788P5zd0/pO9pBW70oYadn
PiA43XUX74XIBBmAI/BfGwF9FHA8SpJq8rUxo5aZbpp6/sQUGXCi6MT4yKO2JJZX
kTAGtYd1zWDZLdpLEgcNaLMdH2GKTjYdLAbLiP5Hsj/z2kjR0awjb4+4E8dpjpwl
r6bthAv53aJb73IN8MA1yN7OEZvIA9ybAvNff6Nh9f97MatQjExGG9Db23YMXvjY
Guqz0MW60+Gq05AQic9S4rvn12h9jw599pSosM3Bie+jT5FddgYbRLzdR9T30u8G
mJKkhPVZDsndAGZAIgZKVYDii3UHa7BhSkR+A6ynzANmgnsUth4WVrfL5qDqtMTo
rc9DpkKJOADZ/0iiQxovOfc6Lm71kz0ctMvQDJTc9R70Az2+xH3cP10iKG7wgUVI
uMZJglj1g7aTEe29Z5OpzyeQf1mMWk3o6So+2rilk2qnIQawWYA7ya/6lXJqn2fZ
azCWnG35z8GNYKwOH7KdV/y7glCoSII7AO1NLy/tOM1tGxJUM5hu86yNvDYgVIeX
O6Imbas4AWXsL+LixRtf4XaBVn6vtkMoujiAtsM3EeZ8Dpgvgo8VkXHIb7aMgDF4
kL8KfdjOZ3lD7gYH+eBnRq9zdZIWekhppM9u4s9diP6FVRpBzowx9sEjzdG3uA12
nouGex/CIHZbOFongzvm9y1p0sbhuRpLQvRGNrKcaxmdZwFHcqAZfquuprsW07ui
gDRVKgxA4K7hPo0xzDqyQflaIRL1icIFU1RHcCpcuVauGlrh/b27QY3FbpEflQtm
GRlc4VGy0M/1Q3o/wRnMYsEGiwd04BoI0tdh24uFrOuOC8By+VBtVBWcWFYwWip2
O3F1t/cVj/Thg2i3Niun5QNpB0f6bdqmbPlZluPfy3CXqZ3jD1buekNlgtg9lY9+
nLbVGMn5PHMa2HqANcrhO0EglrcimURWRKg6wTlVa/IGXu4Gc5gD/oWHuTkbh5uc
cZ4ddrLc6ob4yxWUa1AOH34ISrgly8qNPEVUa7zoEUnexiNODrmsmC0zADVQlsw3
O48wtNYgnU0QBoZpveJxH4dGZ9PErtmsOX1mIAA1z/MmYDj1Zec1bJMJoN3hbSBP
/axkcHJjSSzPBaztfQL0recs0ngZhL2T32QKIvs6MPyncukxBbG9A2P1adHHRQPx
yuT71i5bw3ORfEvlI9SBw3Y8yB/nObpTt0jGwk4bMMKmsYUmc7P0klGN24GGzmEf
XSTlyv/bGOn1Sv+OX+XzRT9Cezs5PjXZ1+6PpLLoVEYUcAs2JxtKIVL9/nTPx5PN
ONDHbCRLYP/6M5/JpmyKNDwlU8rd3yNrmQnQ5/yzIrjbPlkhfq6Lul6w+I0INwY7
c9WD3+XwMgjZG7MJlhIuicOTuWQty3LLIUCjeYGDJ7iFe48DG2DmorG6LOs++ofJ
G81LTSC857M7//owegLcMbkJhGBMl/cRCM/oMSs9B80C8WBFzznQaCUqUgvZSBjc
+Borpm4EKm9XUhQezeYeQ3WlOKBT6nhekMAafNUtL0O22TAVKWIewBRvjpzHzf/C
LX7efw8YSeGv99eIh3FFFZVQgszLWWMWQGRKl9/AM2+LAAeTR5jI697nFZ5OHtAb
n3srnP89G7OOjPgJShvjtTlba5UrQvpg1Gj450uJQTQEj4BBz9RFlcoOJrB8MZfv
1v8iMvUqnjvpELThRVMszvOA1R6t7Ovq8TVNRHKwwVJiPV9Gr+9WErU8tSntEXBO
sNoV5Pa+0HyPqOx4LUElOV0XkW6c+koSbjyMqNNTfoTn2iGZmsPd5Zdb/Xy0BdPV
hR5ywU6h2REg6N3prggpBHLaYkiiocDBu7MrcLVR5jG0GH/YZmjwJGePvfi5aTXv
Ty1iH61ng2NIthsoLj8QrqXsNljHISLqeUWVG6CaZeJFUYZ6QDYLJdyhrzvwqpOQ
YGWlL8En+qRpTXds+99++KnUhscnU3vvsU9RhE3G+rREjjFwGQ8s/qFb0eUFBEs1
DkXGs4us81Gc+YSk3Z8z5FF+QOFTn4IiBNC83+ch2ZYpykH9mM/mgrGpgRMJpOAm
PdOo3kStL/K69eXUEyD1p270qYtB3R+W1FxtrCeyGTU5TiihGgYcwisPiwg/eDBR
jPRucp9CDhM0S1M4q63r2RPqoNzu3HAEu50Pz9QlvdO/O4RfzvrOgaZRuUOrkuBI
3m+KzrMM/J9WpXcVQg+Bn1Wed7frLmOTuL4MaoZtU87rZ/IxSiUg3fRCmOcbHSyN
lY6yMdj3hzPn2DYy+jGwBsEeVa8seQO9i3SeHq0SWmYnx99Y0ChgXlhO8jg89xod
wmguy5VyHpC362tGnK60fxWHHKLQ6B3SIIqLUDhr1CFtGjwa7OHmhoXhBi/lR3Os
spNWviOALuDcRmkZojuiartFdPvCaPJEMgxQA8f2gGp50+isuO3F/6HAbJPmDqFX
AyAYwbbVtmgFrQKs0pX8uy4fjU1yJ5Rtwb8nW+90kFcDCf9LOM/MbTVudoPkFKYl
qLNW0yjC+hvo2Q3Sgq6TPeTZf8U99VL2uo9r92cLzSBih/m4lKjWUjS/l5GiHoVZ
xQeGPcB4plEaMzBjPE/82fKfDrj30MjgU+LTh0BPIMVbt+UhaTSBQ5ik70EanOf6
AWOZoYg7HzDdZbCL1dz4CrCVS0ErC+8WhqKGUME2k8v0a0MoX20GvhrnR7CjcWF6
4Rj9v5kqSxWMFtXxLN8FsW9ZS43vNdqX9cgBzXWzBjf9IfSDvXBVgoO1DDbsMymq
NqF1pQ2HDvgVX6p7lYMl0Rm0nBimB1tjTJ3IJgtoAGWZ7FIrnjcR5OkI1qC42dS+
vzeurvo47ppD0G+LycKYFXhXj624lKADVUb5gtGJkU2YaOopapEBJfu20QqRbMms
J6QRThqNOxRdDA8OZm6Hsf3SevgPuzGwiFKBoAx0rbQXAC+HTC0ncvFxEYZ5ssYj
A3GQkqbEzWclZBHo8bQfNzsWm5rgnraZNHA226qFmK7jonJmF/lz+oxdTE3NFGPC
E5SrASx9juld2qyjj4APPWS94YctDfhAjAeC754lxWjwfRbxx4q4+ywK3gZFz79e
NJJSq3IBbSA5Qg4s3ealQVZkSWPs0KNpwogDO9mdjn1Podv4CsqELtNmjEaLm0QK
aIWVs4v/iY9NMFVoe++KJhzMAVFPn5iLwrSl2g8j21+WKrorEIfrx1aqpdGLZUEG
8zx5HWlL0Xr4DnIkVrBlR+zEs6+KyTNJ3NiZBGqJVjZVX7ditsm8z36DpEZXZPx/
VuCryRfcpzpuP6aD1SEGVqWQO+0EMn0b8jqUGacIFpjPPt+kwGOCExyowU2aVwox
cdX1MO9pgLZn4pcH3UYOMREjI+ApLyMMgrJ32ukj37gt8Yvk/Lrh8bDznei3bD2u
HCTfqUUO4YuL1tkpaa2Uq5APkyOSP7aVO3PYGySy3XuNNnizoo4umeC8CWXMBIl7
yQknsczo2slk9NKRc6kjboM85Q1xqmfpBtl0BQjWd8wlfminruqiCVMsac2dXquG
VxExlTt/ao2t7XATEMc2f7HftDMDEsAiJoq59ZD8yXZymGfP5L9PXDOkgzOFQl5I
d2vAyaUhP8MYbq+dyPfnOuYaeiipmyyeZBeSdQKVzVx61XkFuctw+YjXYQCUeJ5w
ZuK8jxR139HRjX2uauRbdsRaafGmSBNkpCkPDBbKKuvLtLDoUXmnC1Fopj+tQgkY
BKiklVFNYjWQsyRO+phXnAvBXzNF6mJoXl/To6Ta25zwTd7cyTh6pezu4vKeRnxP
qvVNVB5aUSHcz+sWAxXjmynxeNxoSzlcvoWnCox8e0vdXSo5gGt6yEhs/lcsO8Yd
CSNMydjclKEgz7ufY4rbH/Kiqn13fTNEmXT8jVZ/VnsSRaNY2ATNXJO2n+11zfeq
IK/C1QfN6mfGg/7f9SYOtgZu8yzBRJsKXIChkIJYss3/IL4k4zPAaWE0uw5TqvA/
d30KdGLnF2ykqTmDtrMhufFxQSkbBbgaB/jGL3x6rKoAtV/mPMAcxUwghrzwiVXA
djzu/eCFo2iQxe2qsK+qeY17GOhBDjFhQrgR13Ms7EmntuhoEVCyNyGfn28eNHfG
hJnitFjpHPvNALgOhdGuWxZ0wFEp4xQvvrP2+Lz4KUj/+f5gTJK5tDZzqoKdV6pk
rKFTi7W3btJ4JphIT+0H0+o4neOmQgSGEKd/UB8UG0uIx/G4hzQVCye2JXkxg9s/
uX4QfuFL0xoVphU34ZS6AXYLGZakAf78HewVosPi2gm9CwW9JXUB2LNaueN50MH0
AjHpq1msVO2rK8MP6XUU++y1YumlTN7sZ2Fr/iOkoGnSkD1ZJ9dX4pzzYYuuL6hN
KFJq6mcMF8AQG0QvMmvtF1cexbWm2tey7UWKOmwa0QBKINMHWrQPpdhotva65y2g
9AYOq44XoCiBv/72pjkjhlKDOscW7usbM+tTIz7FuSDFcT5aS/q3TGWvXwRnUG7u
TeZW5oVaRA4Do/ja7Oxkd69EckvRkx3c/pU5taxGIzSG30rqum4BMale9hoYje1S
KRiIzR5J7Hy+sYZLEyVmZ5GCD+PmH+arN6cqNqarkAOAHgpids+ku+WNSXBCflFv
BSK5v/nVmAUn95q+eWOHs++nnb4Pb4auxmZOeb7siim+CA+CUtUHCV9B1dHOC91V
AmbqmD4AnOmP85O2ug+f8WAelwamdsiZz81d3YJKx8F+q3m6wF+3fX7B3QIOqirn
pxV985ErxgqR5u0yiG0q/6kx1ccz/idAZa7EEZk4udyFzlxijJVvN+KaEFoysNHR
RTy+4QY9PYvMZKNaBhOAbWK0QemUCLfPHxOtuT0bMqoq5gCbZ2uucZSESu4lgy/4
eKzCW2A8A1ErKz26f1OLFpp36mOrp/EPpvK/vpFFxV800Ew+osiVXoO92SPpcbOw
CYQjl8pLb1mxqBjmxYVRZcskPuHgPo6ht8etJtkynmYbGBv5wQuUWPRcsjg8ab+/
LBFAhiTAzOUhZopkGtv1yKWuwuV/rFHngKjqMg1hATdPS+vOAZFSMb/U3gwQebCn
makY7J35ATQ3DnzUTpcxXzuASXeE5GoXFbjlqYcXilxRzjK8CXPdJ936kGYoFFGj
MTtmZmg8ntvcr0ppxjvfpDvdA42Pmh7544vtZlLMc53dKYKFDtc4lsGD+Oq+BjpZ
RyRA/0xYou0V6/DrpEM9IxZd3UKmm7aQ+5SCuPS8cSXfbQM6qaUeKW6pWrO+f5r6
PWEUvbbEz+fDX+eZw9C2cW8Lp1qdIl1Ez3oU31TPScsHX1a2FkvI0MEiKhtltaD/
3JUnTPhoVDNLi2bQtKnz7MgyOypqIjaSP12fAFFvxKYvTH13FZbD36XsqkHT9PhC
x3o0oTeCV4oM+jEYMAAQGvM1AghYcUPpDJXdw+HhxbqWERk3krudPH2rqOqUKU8z
am632MQsSb0F3xLIF81V9Y4YS3zfugJ5g72L2bXI4BP7AGI2d4haQ6Znn5brc1zt
BbJVnrz6tFZkAuIjC1ZUb4iVqkpw3ny+Y8KL2j7/jAXcMpQx68jH0JFBx0Unz88y
U0SNvzliCTGUxACqZ6t3hgiu2HUvXVsC9DOiuNQvaXon8gVvMgPcfohoz19jDmNY
Lgo9RHujlc8L/njUCgdEqOngXG5Rb6P3BfWDwRAjIYnzkqcH4aA9LvKoGzMZy8aa
V3gRY2HkNtJxSd7AxC//9D6Jno0rLSaeDyaZJ6jb9fWteoAs3arvH/zj20/LbSYD
LY562A6VfzeMwu7MPie7H+aIucEDqUnkR8rVwy+dU3hoAPkkh4WFQTnuWObFRHtI
a1K4S2PtKNgi9eSyXXYyOwD252k08q6BM1TwdHaFDHnoIoP6xeWbJJLEP9IbgBgY
cElqdOkGuqWdesuz+jLxNbzzeEt5qIfQ9r4QJVUbPpp+NT1lVLhDKBcStGGJSPDZ
al1TMngYN6hA0U3z/cPlH3LiUlF1699bDH8XY77qt0WtqXF5gXvm0n7yJrQDAcR2
CP36+qiGQ43PPx5cdEeia0MDFo2v6byib5Z6T0020JeCQwImxbBlBiEfjJWEFgED
n+BUBCOMjoeSoQ6zE0dWNZuw7irudAQzDLNyUxQZOf9mi9HNK0gkBhbvxUjcXw0I
TlJjwggaxNW95O4qzubBdaZy8QaY12s4RzR1ZQAnLJ5vTKRltUdvexBd+Kl40rmJ
lLRlpILCRseiQvQb6h1w0BezAIPUVFwI7miDt+BE30EKrNEu3+qY8/cXMicYYhOv
5tBfQn6p4Y1jBXuoVqECi3BusZ5KwKDaYXIGia1rY3oeg0E09FnoirJvhiV9rkf4
YLFz279G2XFjLV5q3Njr9eSPRsFZAjT5e7ftUtzsmhiMsAKalVScIDMQ2kCTbLGe
JoGwaH2utLGmqkZK6vuVwm7EsoIsbSHK9Eds7wSVwCnxGjk3I9fgW8rICn5bhHbg
c76VR1/+jB96bfQKb+nZUteVdmANBefnCy/cYgidg9mwow3j+jroiukNImOQz5QR
+Tq+UtyZ6nXo91Xh9Eu5Anc1mUhHfbGe1jvVoHqBW+HthbEgAYQmVtlRemfx8kUE
QiYgAicINEtJCctmyG8mTpqAD6NASfvqFHC8W8+OxKGNinn+wi82DJZtF5ICETyH
1vRnn5Tn87fOuI8O+33Vrg9gTHGizBdljNxudrumzeozauQwjGj3qRCxyUcPBqG9
CjDJ1x7TkfwMQjbGuCHoeNDcmMxQ3SPNCRdrK8x/CYFJCGP1F7abrd3by64JLoUk
2oLTI2H9q7zQsNfTnTiaaB8Wk0UL5zzkhJJq5FRXpF5sP4DH2sCK3aHKealGvVRC
ffrXcpFvnlRQbLxbU7KZzHxjuo/PWLcWAk4zcEDAjq4Mk/KsMhbFUlPnyocHX0Ug
Hl5+38rb7ZvtEJr/XfH+VeVEcjPfFuvibScXYzJY580VPLOcX6wCK0cWgDDM57qY
EfatARcxk3HEKukIlQmfLjoswPc7oQ8PgW+quL7r9nXXweHa3KHKwH9ECaeGQuXo
75qhMO5/n9uhA9TL6fLjObLXYyfSSe71EH1Y186S20y9vwf9v5n1wiZAL6RfsR15
gi7+AtAD/3idNqmYziAcCcqWHHqGmn03RQ3BDubVSk7gwm5azHLu4OGttCZuN17B
a40UI4Qc9iNmFTgA+zgVCprvt4XkzhAfg375wq1udMcIYLPpED4hWD4Mk3NcXtTh
TvWqLwbiysjVv7jhsJ9ato0do95Q5iYspjabm1myVPzxdn2KJwwmzCLuqfbN04Kb
7h9nEadVc5+2SacKv7lBKpkAJtrQO0feibiw9MoMAipzaXbgJb8gLP+aRnQ/qidS
Hh55Km78n9V2E4/iTYYuF/kYiGJxhLR1A6UDgsjqzb2N9gEhZk8JZ1vx0rE8Zjc0
QsxdjbPyhKnIjqSr8Z7f6C8XZak0igvhJHdoQ8COE1dWTnHWZB4z9xh1Xr5KnJPj
H4VcWKSluy4yCCAG1vhbUpd0U7mownxgXzNtv/nZ0oJ3Y8fMFgX22CVeQ3F4OUee
naqU+baiar4wosICTVSbj0daUJtY5qOpouVOCOCPw/oOk3SrN32v9DpuSuVkrExN
9dAT4HVFmiizoGNlEFZqH5nzaVIkS2PCbieoyLlEZyDLMdT1EUCHxF2mDuCsA2x+
xGsfMU2EyEufzshKZuyypV9U6/1NKXgHvLithInBpQAWUSWfkIxnh8nPvr5nujOP
X01k1CLVSNBVeHwCCXQaqUB6pMfn7n9mdhxknbnJQWZ5TLi2zEEZtF2teV5dkf5B
EQ36LpwFuD+KeM9yDv1uRW1eI0r2Roykdpyucumx2eMhZ3x6CtBBCKWy5+A1Sygs
kR3OxY8XqcwED91LF6OdBHPO6scN2oCoovpnDjVYGHY93x9zVNKxTW7X+4Yah1Xy
joa+T61lRcV0TESySZfCLtEhZx3biuTp6Knyk+7SoCEveX0pcY3D4Zu5eX10OCRg
lMXJ6yQXl1mARXQXzpfTcuY32dcNCT7jNTALZTXvMwRqTOhppd2mHsAiiEpYOeG2
7dKcw/JRtWFIT9SWDatw4ViinD1bGEkNfa+ESGt5R40dsGdq4D/qXdZniXh87RGy
YxjEVFJVHeRpFZhdI+i9DuPStLikAsH61twdWrdvty+O+ewNN+1TGFH9TvRNpgRm
ZVzQtZA0FIR1VPiBJofnj+uGep/nWYnDpNkiS+1HD9OqzZX2SpzUkDGx64hy46zO
ZEdwnMPkRMfWfd8JH04sSu/uAQQR9t5EHnckZc7MZ6imRkMLwgeM2QgdLPpo7kyX
PR8TJfz5lWHNHh9XdHsWOLybUqgVqi0gSnP//I6T51PJGjrRvtXNoTWzX/oVJhGe
eKCRgx/DXqglsmUs6QURL2vEouYgcNOcBnTOkGFPW8dLlmKJFUbEF3OD5olMr2xb
AAIcMd0oL2uan/jQHPTQV7TKATFsLhna5zVF0qqMthWRz0pesAJyxoKWUCBfaGgC
1OuTThw439SR30U8Wc/cco3ICshm/SSdRje67mFPaBbpxZx8yCNpuIVKM5H91Ngd
ctT+CsvOXgX7BtoHlK6uXVl776EvluxHf/ovVLrm7mqacpBTf+sBZCerQuKoBPJu
MDYJ0NU6GdIvduSxyg/eQVyWfKe4pjVs/z3A10wUToWc33onjkyUesyo1C2JVSsS
bfaM0STP7Z1wAYamcxMDTqrs3YPgr2x7Du4BmOqctxuwy/oK1gRfWoKL5o2/ZwMu
eobUaLFxpWJxlYsy0yfJxps14tEWikwFl0rfbs190MZkM0ya/RkoxFcogb8rgIEG
Foe+nkDM7oMQpab+v0ivyazJiuMBfsX62Nm9RqY2S4Ow/ouCVMc8yXYneGo69iM1
czxB3I9PBnSvXbeZ/R8+4EEqB4dX5YbOnDgxMmFJ2gx31Rbx8DAnwYPBXIzdTRfH
+ttXLmMvcwW6LNquNlK5+yvUM8f1J16tU3PAs3ludaLWg2QqAddy4dzzjzy8CYEy
NWH/NbQwENNvYDQPxuRWECHJkaGH5F75I2DLrjIHTQykKKSWLtkYm2GvgC9XF1d2
jw1O9Md1oVsCFe4C4wN0JFJChIK0CynMTQ82z6W/h0h5+ZQIOKMs3jmhi0pgSM3U
bHhlkIbCTTsVv53laHgmetf0dH0nHM0DIpJligxR01nUtQbE560aZxrIPNoGdAsp
I0m/5FnDWevpv/ORpQCVC0wa9erF7LxGL5CSummc3HBRn9uIrsi1TsoemdlZEdsD
vCu9lhtKirvWYBrohXsdzmiN/7PrsODdfR7qmu1QKZESZxtHcAgUCEOEfWVs8yZV
hL39QedA/uDiSgVTDUkIoc3kaRQR0yYr7drOTk4fHva80UaaydW/eKI8BiPapCWS
QQM49k1EVdqXlThpxdgIfeOKbekv1+Gk47o9EberWzMCPWAsoHtkx9zBzkME5HdZ
IwtTpjOqF3lzdmEbB+Gx1QhLJMPYwKzjozp4TRpvmXdPbyrQI8cR/qdHVCbllVdV
TRaHZ2zJHX3TiKr4W+N9NBmfePPwKSdJP897tB1DrC3vLA3dsM3hpBqMepx/1qfJ
yqrovtI4LJuWe5RrHEyL3QSQ78VqhX/4LJ7Ms6jQpnktYGy47FmytIobuEZKlQE1
p1CPKkqp/qtxX2DYoRFWBizqsBoG1SbySSYiFve3wa9lCwmhW5iAnopdZm6ZKcUm
3rVqR59PZ2Vp1xe3KSXbhhrdD0eeQrt+NywqezYkZ+jgNBR8Sa6IA/kANcXKQUJY
kLKUOqFF9Sb5EgWAFfROWgYCT79mKjx1kQ293PNm5WxzcSx0Gfsf5Cwhe9BY87Q6
DPzZFAMQGuFcDpHi9vL7Jqplgjtwew+27gSxZivEELIyZj7PG3tm4eW2+6WRBgmB
JJGT779HbT0lwmfxwNkAzeAvmysV+b9JpYpB2bp7Lvy5+NbWETXcUkbChrAuJ+i9
9X57WcNYmmsldqoSY3Kb5s/lYkIWvONaEVy7MKLN9xyA92sufU3PPKDsISH7GeZx
Jf9dKx+3wCNsWfwkV64Cp9QYPW8hXwbBHlJHSHmPRJHDM9SoDpq6wgLJI7P+c86V
q/uelHT5/hsKVrSgmaYgHXOpABemsObBzGElksKz8+I4ZXNQ++OegxuGBYY9VeCp
Gbeg0vC4EWjfKoCkVzMbvrGMz525NmxEQ8SpWDph9a38SEkL114XMynVBJoU/RBi
nUYT5SqyZ+NP+5LCweqMlOpL1vPOZOrxC3kyw3vX3Fj7JLBsiPXZOuE0f+8Ftq0F
S/pM6qNyXKyyLHqzJ2w3Wjkhw3/Te79RqxtStTaNPhBaTO6Az3qXTewc7BUsaepB
TfVdQfZbVpL2WuwXPFN+7aHcvtXDGzIHZwsozUIVzaMQCBUS3K78FQqspYmDzlKa
xFX5IHQhSKy4nIzRmw23jj5Ak1T1yXr8VFax1lRsIQ+sn4tNQOVwjrCIhaVnGAC8
MpXbOrdOQJFbse0IzaDDOaXVdAGNkwXx27fN8+YLA6J7wQREmJzhVZYCS+ABbuOy
R15o6sOb+ZK3SEsA/dvQXFnUaRcr1881E2mPBVV1MKFWndiQXSpLY9C6f3y8Vzfq
Peef1LR7vXK+bgb5fn4fmKhMgWWi6HY0jGWElzxbd9JRcND+x7rgHmhz5mT5HRRd
l5vJHCpi1cNyYkjtVazhV6SY7eU4lepL/BvKIdNz+CbTwCA2bWroNnmUlNBQcUCF
Z7efI0fNorTdz/BALrkhTb+KOO/6cnH0JFobAWMTA16lXt9ZD/0/I2KWqc7uzyco
K/gZOEb2VSP6a4VY4GpOF/uiwHrv8dtmktSzU4xI6f+d6AF2npAQaFGKV6YQHfZy
H1N6Rlw7TPu2YBMBntG9rQVzHhgvK1W70t1RnmvjbI+WX2HsKYGTHwAwtsxmtAeX
/3zsNI3q5y5XjrP6ZivqGcK3kupBJDjMl5TSDKa0JsQnXwfys5iNL5uJfWmB/D3V
BGbGrtubwrp405tIP6BlEVcPoqz3IO0TVbE8+zB3ce4UcV+dkV6u8YumvljJblyv
BCqD0RgatRE9tyVD4d+01fPQpat6ZmNe8asHmOfClupPITBlmJeDNWdd3F76NjMh
FgC85wyxeOI5vZ+cgo3WomS0OPTxikSyX7ZNIsjSQwxAjyYJ0MNLQnMYjj1KHDTy
NeCUIqkmup154/t1XyrjbBLzLt8X0fUNiPz7h7l1fxV2Xq/z5VwaVt6Y/eoWt8SV
UUrtqBrjMIMb1yW7IWBZmuVDK1Q0Fi8U/4tK9yj9NE+uyStbISfQJxtZ0XrX6X3e
9LQ0fdkeZK8Q2EiSj2UJN4EDGNwQg3p2toDIkjaATAzF19wLDRo0PDdHg1q1REjk
nwp+akU1Xq+RIv6UNW32gYSoI+dfSku057anhu9Q6s5Q2QZfO1V/2JqRb/yEIF5e
+6uyYfH3IferR8/revJztB+Om9giEsKhxmstVH1H5zdsLF2phNBGDtbLJCSjHI4g
2l0aRbmZVeEwGw1uhafX1wB5g4kHTprs72SEyvkS3ugDS4YMwsVlhNiyZCo+D7rP
BJ6uRGjDAh7/m027NijCxhUXQ1mWKCqJ5vq745/AFxfQXWRz7SMKxZsOCTayi3FJ
JtbFQt0lq7YFgT2Tbv+6FxS8xd4WScePyLDccazG+8+Ha2JpP4pCP//aiSVsGgSt
EtP+fanB4t06A2+uxGbdvnONe122NAuTHnHf0AVDArC9HrLMUALzXcQFAAiv2x4y
9C5OFZbuxntWUuHcRuT/iuOKYJREUNwCsBuv+i++DZ4vamdeydAgpK7e/RlHze++
Q7Da2ymwMxvonGjEMkO8vBCjNObwqvkJXq+V6Cp43DvIG0FjNGQDnAEjpb15tRKI
BJb04Ge0iZaFygqKcETM4D7HBTON26pe3hloOhawijHZSbFa39g8B064PNo64kHp
moj8+wclcbcrNHT0JH7HRP9eVC+hT1Yd8UKuqgVrmUOBl9U5EWd0PUEsq+GRhUZ4
GjJZh2Od8TbHEBd3Kce1/thrK+uEC21ohOurUPRIGTIJChOeq/In8DsitwurgZQA
1uZ/18fibD/JJbn5zekRLzIZZIa2ecEEUX9P/RzeTbPE0ABtnzLBQyQpD43z/Q/k
Gh5v6pw0mnkqtHyU5YEIWzkfgVq/ue1wm5wcL59i1cmCFQUY95iVwNa2Ms1rcG7Z
U4xw3MuP4nPpG3l5RjOtB8StpyKPDWTubbh80QFvxVZhD8G/N7De+Q0YsMGR/MSR
thLY5P1Puq1K1lQfPOnJtAK9d0yQnORvXp59EPb0/dhp246ENUR+oORGyaDv8HLr
msPDzamVV/IfqkFz1gjM0Jy9jbmzdO4Jx4O/lrsdsz+mBXjsM1kyhlV+NSLP8yvx
jcPifDeG0HIELHtvD2332Ok+XQ0rqeBWmMiXPlaFp7fdzIXdaWh464NJWCL14JNq
c7+izDTUAlo1TMdI1CUY100ZmZMtGBuylBA1h/DdKF4Si/FAr0sQkQ9jU/rfAgvc
r3Ish8EWdYmN6dAnVBORNBThuwKULcWPZOSa29lutzoErVwFpZ/1rv4vx9hwUJb2
Gggav+2fNh0/ql+NrQaLHL9Yg48Kd0XjGrZ/AG6YI7avwAccTKcV/ym+e/rVAq7Y
fMH9Pac5uMY+1J+PgFdZA26jjTkZoKAmWmUVsQFVbBEFuucFL+dxQSYFEdux3Kkx
XUgaGmLxX+8lS02RK/iZ+VmsG8Bkte6tv3xVOVXGRpHFfYCL6/5axceL5ZNtfKCZ
/qA7Ws818Xfxw/sPzzlsPxAsUqQ9er+awiLFjMJsbIwLbCx9Lno0XYg+bGaAQisN
B8g9SF3ULkdekQROQpvL/rJHKdhP3MSfsrvmoywRzW5jbjxn9I8IdBAe6n6haWN8
gVU0nxH5MTVpvbbVJfpLB5629fKp3kGTDlsH7jAVbBGix9vuIjF/teF/FvCXhZlD
WsSg/sW4R0FfWB5s/2WX1nMfoZ+5yOg35NW9Vhu2b0wUg8cWeQqh9Q8k9xDPU/+N
BGTS3sGlbr6qktJ/YNeL7A0bAsR0D0UdIhENdYSloQLMrhLvXFiuls99p6hGI/9b
WaEsYJAnse18fEjEQbtXl6a05ZemDMbRbWJmeBZxycWHnN/IEKePdJka1RDk4+sn
T9aO18xC8YWE6OYtuyL1j94qfKhtQ2D2Diu0IGMhx0TSkKkZDDiT7VQpNqOXXL3N
KAsB5/50bTCbLG4et5LGCrx+CyFqmXDWvbdKcuXg1udWYwWwmFfNjGEEOY+h5Mwo
9eWSatUU+AhO6XXqPMzMfXYCewT9Gcv/Q8cMjNaGOOBdxxJ9xnEcgmVkZ0RhdvTH
zwZNVGRSMTTwBVdTd6T9AKTHXhYIbse4q86k1v+UNhYqqBPzpMqpRFOphzCa5BvW
CZlhAZGrZBGya7IwUxTiiCQrt1KJnrJnLZ3rSbgwkKfW+NHC7Zj0UnK3H0FBLlwV
w5RYgu3gtxMo1mmNG+fMKdplLbV43MutC8O0wCrMBcXi1/ZjeH630HFBdi2nz+So
pQThXX1ShVS/KSn3Kec0QvAal1FyFRYn/prmVK6dcZNiN0Fg2NEvycwAOgjeBmGx
h5WyUZ7AYzgzCzuJNBvdzRlF9K02/JEM0S6FhX6/yEMmHHW9t5/1ydpn6+1DbVkz
YyeWssNOw3DwYAoxq78HXUBQz9vrB3Gh09LSUxHcBUqSe0vme9GgVY1lpbX6jbze
spMpdUXGSvBo0vZV6B516YQfUnsORsZoNxttgujJV5FTEZNEpRY+n6NLaLAFAn7/
UifFlFxu28X9C2Z54gi0agkHMTa+PG3RS5fCKHnfoFQXbAubZwunVc5BperMdaQG
u4qbe18nGf/Pva9oRRb/4uKBP/IXQvDEou/2iZrLcLEl1D0IZd1sv6hHlLn3xCBD
tLvl1UNa3n0jC9SjLxEUDykLL6R1VkuiTCiSwVYHdZ+oxQdUQD5Anr8jr6v0B0Ev
mlMaPymo9U/byPXqNWTZq6SzA4dCjOHqVvW7y40QCsy103ZAEA+Iljfm49wENAnC
oU4Tkg+gzEjle2WG0JneqEXpHzQFrN/ByGd5M5G3UF9GQChFMmVaRng8SgJRczkx
rMUQtWle8IvET/KdDWV/QTPOdy7auEmnOh84R+WtG6G0V/g0qpadGtHaD21vrlp3
Gkltksov4NV0I0Cw3Z8EAsOWbZ9mFJzYN9yJBMStMuTiIn4WXhJLpfp1CxoJUuDc
1vvatEfvx5tLofnlo5dzxYxeIqcQPv8BTXVIH+eim7T6fNHt7Ld6q/u6H8rDQS5n
1MffZxzgNq/MwP8G/fdymvNdcaLVS5iY4INkBY+wjlGsTj01mLBCfYkkJKSO2Uv6
fO5PDSy5BkIib3CBBaKFaleYhEd9oLYTmBHDkhcFTgAr1+2b0gf1MkXydwQEOj74
7KQ1zm8E2FgSGKpmMXRO+/UJXcBj1AT6r8nog80dxCtMBsIjj7Tgk0c2ob44kRSq
ZkVXx02HA9eFI0nxhUjIqFAfA52qawvlH7IspEZPUEbsVGlWVqeoQ1c1puHRr21l
K0xqFfcB/3gsIyUN97czXRuMUoCAwow+RJw8zKmLMtb6unYjrL3oz1sGxYxAueWf
RXG4QDzu7LviZGtAXMJjOi1LRu2VIb3bdxc0d94COKWjWF39V0ybmxWC55Pr6pNM
S0uniism7KE0SsYOm2WkASAd/HSxVUzvxYQ6IrIyahAwkNN7EF7ABnntlk8nxxLU
6M59a0SFWb7Cpxyq4sgB4qynQYKWVBT5pc7UfaDiAb10Vy6g396ERHvhg2wBkz9+
JMpiEoqHRcUJ0sdVCxzIItyY9x9fCkmvJfzrbRxq1jRPGwZF/Am18Pcy1JHwIGSr
/3BSxUAwMNv1SNPCZHVjgdtSn314Pno0WKRo+Nn4wmBl5YRvvS0yYsO1iJe0T3dQ
PaW9p3iIc2IX9qexy72usif5E7mMp58SHbdLFj6LhwoMVbQkb4QI+zzhhulS5gpB
yKz7O0IdsAJkPaFYD0b05GZ2QXA00jILUleXawFET2dDzfP096yylcMkJpBEG2Mk
OLabw13/EXhOM9cBTQFG5dVBmuLhqjx+sPeLv1pBVTdL85tIIjkAbJt1bMUsKuCt
fr9qi7mU3HVniaWjx69yYoVK0t9WIH3Auq9XC5PlHsQgOM1MBHRcZeCG5zr+kZp3
MRLxrxTYPF5ZMjV2cdXO79QkK2jg/eLwgSjv17Es/kZlavlMcY7oSCYACQLCphUX
3EYykxl0kkh2RTfpVRRE0XEvr/+uNCOn31B/PO9XHsKw8D0mJ/nnfHPHzuM9wiMG
uLGuGVw4NGtP4LJVRKAU2skV4PuQHVzObCR0+WzxL1NH0qqUBYpiyBZjzFdUsZS2
1xGd7MgTlePz8mReAqsXf80UX/AVdEzSaDBippsXGZOIgla+evoVYcvDdU5U4AHV
grbRfvDaidn8BmG+Nyy7CQ5VWyG6XdFkmAa4hBD94540nLJfVwHhYIRLJhlbalIB
4e370QlmPyZx6z+Vn3lkBtR0eOKGkA9kvnIReJ/d4gx8q8SMdsfLWzlZ69SA2KAK
wn6airGTMnzJGxg9oVuA08kIp0D7Vxj993rW/5EPIUU9YtoRH/SlyyV6PMxqRvL8
qNQOfzxL9LBN0HA/aY5SswplPp5LUInQzODqwsORHGoU7Dq8STdXikMZwIrtkBZX
qyd1cv+nK9HmMO3slwlVLrDu4MMfTHsIitO6zSN3TebP4BiFwS/9nYbEuTl7f+b3
ncXCF7C8BG3qc/jjfqq00rugFn7aLHdqAXccGtKoAekMtrD1FWnZORWaSuN3ZkU/
BYX9RtXJuUJwRvdA/vN0nGNcgegA082X1FBSkE7vellBhuzOZCv6CJo64t1Li359
kPO/xhB4eMzETHSzxIqyjmQA9zMRbQnr5mlqSqz5MQ5r4ke5rdvBM5artUVf2b+/
8R+aFG13YZZ82RmihCFWzKaHaAFkaD0TrpeNWVgvqHCpUS8y/I1pjAX2XjsdcbRj
4dIYr2G03N+52aPG9BX8vAStYa5S0QOjM0tJxl8PoSEnjVa3QI0KyTPuddraoIDN
UYJXUpzuCcUUhHdPRyn7bb+OK5F0+/UdMjmmzzTV6hQmcWluOVUHAWWVTCpERDoD
TVI3BXYTk0PDtIyVfCq8Nw03yYSSlhDfmzGiKO3uqBESdJPixR6IQgXpZzDztA63
KkyM01mhJtGPfVBKgkeqvinp6wfltS9iF5uQgjv36QpJ5uIg4K7bgWbGQVGCquob
BgDc83yV8zq3Xbwzxhve62Qi1b+mBw8iz++uvRMMOTi+RSXxTLF9LFRt2U05V3KY
CjDv9fP0ka0ZNsyD0junYAwZLydO4+Y9KMgIsjpntAcM8W/yW7OaqV9onYA3hl1Y
jovG12425AdCUm+o8SZDFB7DEwJ7+/yGTBFVmkjSoWFGdYxfAQ1WQi7ym21mdAB3
emUrDl+0T1R/V7k8zwXUkG1veov/HzrCvm5eF8xnc/nAN1p0x8+Sm6INM5ROBgwF
FD6+YM17P2RCJHtrQSSqB6IrDnyyxflOAu5DbELK/VR/e5fqR9jVud9QOvlGrW7C
eacHTrXdNSKwhpeXsDUG0Hq6ZfT2OB47i7mMAMia7RgFaZy6zJua7QWe+4jUVQFN
PCyN7+9i7RjAKgmYNQbFZxkoOOKST/FQUso4hg/HfIiZYOKh+6+db19k7/MBFPe/
0Ra1tN1QdzskGIXm2O2SjIghGJiJcLnu+ljG2xH/7ZJkSUJRHh3FIibTb8lgDQ1U
U2zy9htMVpoLZTd4aG+fx2nqyBkY0NBp6oBUFTQiDAa65sWA7P7+8f0x89aqkM+c
UdLecZ2hSGOHWmO6CkYJ2KAND2t0LaQfqDh7MwXpfEYD/gVKbWednwjrb+E9sKi6
JCMVRM7BvLYj82LOXZpnLLNFZ1cNWn4kbAMbGu4WqSCUnUWPPAQDT09ayWLzBQPQ
HIQfx3ehRUWM6+Jiko93FeocS6LnSTKWSULYnLRaEX+hClmKisrbLgEV2iVyxS+E
Jw5AjM4UD4MdPDirBuY2I3RKM9f3gJe+3zkJvUeTdwR5G6H8B+jfZt/9R+DWXwVQ
1yssPtsLJA16+fJS+1qehanAluTPeUoyMmlDVDbBbeZbHbwnBkbTFbq9naYhBFiH
I5z+HpQSTmHJngTouO+J+h2MSj4IcAq6hxL/Xyxv2aTN9qcdPxFWtPMGzolkKvGE
zCl/YhK7f93fV/v4cmUZfeRRTxyu9M/DenrU8kX+sjFwr8skxmASJEkB44fbM707
lksmjaXYJ2bQlCuLnuuOfa/5srstqggua9ac3bkyc23xPJ9VuYJL61D4iOp/eP6Z
Vz2PcYRC/NSep5g8yqYIv+mFeLv4jRwI8o0Hsu4+VqnSN6LVU4xkIjZbluYNu3Op
yD0HkpvnfbkQCuQ24VO16HTW0tAC4xsJyBqglZCpgwcyMgoGmUzGGkcPr3mtEaeC
MHsAkxIvvtFwDlJ6XngIorsDIbXvTZuH11WoRXw6kkvLKkHe/DjB/G+vCSvVZQG8
zJyx7Owygc82j5NPvjgDpY2+llO5ArtAI8aR4MLoMCZCYt81q25eHKGbHxOmweom
3Eb56Beeo6dHRYHjGh1nElzXIIwpC7dIs2p4euZxLjRWaA4Y0Xm8PyQGInRth2ub
IVE9jRGSGuptHfjG7wuiez8m8S9E7Gpv1n8XBz4mY7NLbeioUw1CeFbWKOifxoM4
AMFNGDJ3iWrB8Ijggu1GtczYlkEZMU9cixzGmT7tf7NKj1PzrqOZr94w9x45CJ2L
OlRz9enlkM6GeD+52RKjXcLfxjq1V42/Rq5jag+6Ip+kDNX2ou5JODq3nZIb6T9k
JJOeAsvVcArlmM1uDPgJKt/yCYOSR/VoFytsiHpS8F8w31B4S2UcDyWxuacztbqN
6lF7bMobzQF/JIj9vmIGYNybofpLIlOnLeIE7LXjrhuYjUEl/KhzK6jmuX3+2HW7
1UfH6Zft69Pwch9ThMj+u6GwDXljYYYBW8Syks8hE+sybmc0/v+eoY17EQOpXNOS
T8d44V4MqTUInNJkAlC1CKiXd2DfyUJ/WuUlCmlZRwSJDCW2JWyd/U61/fDY8km6
gpVMsqcc0x1lsB4cTaJDlQZjKua3OJ/6QLYGKD8ZVMKdgLudQ3HETwzw3BUNsiYF
V80tFW5j908G9KWwH2Zxfl3/X9skJUhFRrXvPRu/2gCjFX3aAquTimr9Lqev4oC1
kCLjVrA5QGSvWN0OBc/MpLrjfZOJhrdiNOya4VcgO+TKgke2adCSMF3cGRryw63G
eMF7s5SsQCmYzvIXtKscRdUGzuUrF17DBktw8OW8MpwLiwRSpGgXG1BzLJlgr0qn
XqbkMcbj/VCLLSK2XIc8CiWB+lwzdJXcFWhxQqD2HF54jyQJJddBovWgYIDQ3DiC
AOEGE0BHbKzAZcZiZ4PvVn9xesV27IVM0AbOmTHzfd6WY1cXQZHPOuwAx5LxvIH9
b5oJ/nhkJqydTm3fOMpKaEOt1yrpfBkLAL0oRjVIwcY/1SDK1dTUxePIhBYPimcp
HSMoA19Nie+MHd/INkdxPvOKD8UDjtNRdO+FNTrVHALGWZsz7447Ms9wRIOoClu4
spN7vWnhngVEbWroXkFJ+Inty0DCnmPjhGDvmdvRn9CjvVd+Xs/JPR2EdaXotPDK
DVCGDMM5Ot6mC8Etc4MeLsDFliF/NTyx4oc+xkIKuGdvvbqjSdY6/uMjZ8DNYqOL
w9lCVtZAp8JZkevFd6lrNIyFRBsrD1Jtwd5v7ue0Ej45wvv4LKnaDtxi1T3p89Eb
4b1u7LLVU6fW0ah8AUsLV/XFEEcgiUEDnEoGyOyJBx8Xp1HcR2wnfXAg+CXAFSUw
ZWVa4tCU6+31bh3odvtIq5/IMBYN5XW/o7VfEArGpxpv9rffPg3lRjKMUC+Sk/Rf
TzMBvTOvxkDOQBOnitdoizb+jgQoNhkbbJYcQxMIJMX7+/mun/lHzcBz8lAX365M
PfXaxhG+TH7tz84mg6kuoE198FxAlFyazNhSrMAz+zIf0MuH1CUiS7FuMsRAZD0H
m8yIEn/VRqjmroIuFbZA2B1XNoMm1AO/eaL4g/ClhmJejOJU6d88utNctrz8cg46
MfWE8jgjeFqZgnMa88NwI9I7Drt9Ztie4tvqllYwHT5S1ClFeRyx/xCFhhwMTZDq
AxmnUgUHUOp8Vu09m7my4Uz/rTyJJsh9T0jpDJDc82M1H+zZXgN/gAU+6wNytD4S
Rc+LV90oJ+wTp8S5E8ALhbmVxUs1aJ/aankBrP5vrxla2qmiGo7FS2dpJCpc/XO7
gnXQwj51M/DsboVUjpqg255LHdo7oi1Kb7l1JMzgAY0gP2EZqMJmS2LByOcYw9OO
eljvFPFABDsC95RUqYB0kl23f/2Sn0QveTbox4fna6q278OSAkRk524aag/cjBJL
fBTIdZWtvyC4HOB+ZkeWfpezoOJd0QXLJ2GDL3xWiekwcV3l472GKcibqXrKYqG/
18JMVIuX8WbDp+w2JJ3oZelNog1aXxnHigj7jyF9D/R5HAmL83MA+u1lMX3S5Bac
nXPSd93DUt2mEQQ2ElP2VxxwbopoTij9Nl/TgYXyZ8LQkVrznECP38CdX2lGkMOo
deNgdd+7M7FBle4a/uiMBF+/vOZZa85yCA7pBrTVwtSu6vuvT4ENfWaHcUaDLv4c
q7tsartTE6rDj6EAE+tnltlbrOjh9Sh9STst4/C+ZpWzuvGPCajdC+AzeDy1UZ02
8InLF4Zjl2sgWcyh+OKw4f+oY7ets438n0LpkzDzk3suSwM09JDHLa9hLQn3CYnQ
oo2VNBS1Bz9gYxn09A3v9mu4pwWB3+SESfCYCrDa0blLXMD6ZWSBvxDH7lrQn3jK
eEbMeob+CXDLYXhGnrL2ynWlmIiMqgs+oMsyIrrMA8VS2lGqvtRtmLZrO7bxdmKw
k3Vunf+9wTQBiuDKtqwzKqa7xxefN08pvNbqQ1hhgMBHFPJw9/HLqKenVTaVk1yc
yMHHeKYbSmkDJt2nVJJJkIxhprW/A3qlm5SGc4cW3j0q1qXyUxsn1+GJie1axRXf
GUffdjOKq7Ab8s7B0Cu6EvtpaC3zb/sPCkENZpm4bXrQ4kUAQQJdILr2p/be95nP
Mt4jYbY9Hhf3w8igt5JYy5JFiWJEPS8VBudtCgARbomJIfm4Wk2e9ZnQX6aiaHoE
lZfu+N1UxorjtAUvos4yaCnfmrB0ChdF4Z5aY9Od8ppJhqMRMfA2do31A02n0E16
g0FBgmY2CGZw/LFTpwi6xlSyO02kRgR9ezChWn3SCf4b25Dgir8iv3hWCbGy07DO
xLTHtg+cCW6ObTrAP9g8KtIkc5HPHOz8SXZEZdIVoKoJJQlZ06ulYlkfgK8GG8Eq
VTehBG0wnGRCGIxy6M9y3Er6xFb4OZo2FI+Zl6qorNFyequByTmXjbZgYuojj4tY
dH3PHF2Jj8de7LHXLDTYgqzhLo26CKucgkVtqKgbyMUoMiTLKKZaucLv9JSCTtYR
ozORI9spMlPRVgehj8jMifyU5cppqPGg8RO18F2E144Ew924ogP2v4zUf1mmjkx5
Auv89dkXkkB4aGcF09N2YiJLPrPiC2rQqjkY1FtkBTzzWRJLDcx49E2xDNI9CxAN
NLKxbYZtkM+vwzIVCwruzXNA8O2dfwNw77ayRaP/rPpDgvJ9osK9STZQgNSTc8Dt
qbDWVLM4yZFlRm1MumbfarQ8+uzYp+4TJmv5+IhQ6puJYb5FL0kqiTf/Bxrbw+PZ
9+kPFycXq5YElMkjmQ0uptXRw3NfxvtvjIeG5adq9KWfrfBpymZ7OwXV/cKQbMTe
b69YoULA5qxXR/F8WYB78FHLtA3jf8/Ss7YH8Sx15F3OtHmIX2wO15AwGLR/+EFz
+08r2Cg25MnebeQyRoEejeeCSDRH0Pg+ghtuhX0s+J8BtnMu8zYHICnCPXCzD1p3
pNjjqiLIz53qNJwJT97mYIc9XQ8xCP2R2VY5PGO4L+4yCrhXVuebVexsyEqtqqAG
yxcw9G0myDXa0JF1BdydlcXV3FjvImJHVkFQmrVn/xHffeHm01bdWG3IR1P4Vmsi
0l2Zhjr49WQzH4W3xGRqlDzdfi+m4/clCMkR0GNChFC/aZHtvQsPNfkj+MncGWym
iHbM1p9/+R0JOitXfM3Npejvo040sHdStX6tkJsr54TQt7CLfOnYYvb8YC16c6JX
LqAlCiYo7FQnZ9X48PJUctNdFNCpPxz+Kmpn+bap9P+mtaah+luoO3CT3sJxTyJZ
Bi2S8h5l3SXbxPavEVyTiEFdw3KeWkqUKpjJHFuni9zF+OModlz04IjagU5mNbRy
M+dhC0bqWEsrx/teMM9cKd8zHc2LA0F2ggovFQ08V3C2ckruM9IiMZdEXkCs4Fnu
UQYUNA3ex6CfuXst8Pbqa3OaqeueN+0ooHVQbr5AMH1aJM3X2yctrq837eCVmt7V
eUtMNu1DjPJM9Yl69Ca5ptyH0h1GUQ7rOLDnOIgR/zG4VYQbbk9q9SxzExS0x0Cx
ImU2OPVSZk2eNEL28f0vR+hf5TcO0LHrh9ZlkdzpIY7U7Lxcf99SYKsf2y9bPc3r
qCAVAoQ4vJ58A7+hGH/CPtw1nKdy/kJH1Ggwe3pNqRwOtjNRQp1LnWmBImEFEFWX
ajbr3LGvcWLAgBi9ji4Hu9IlRJOYtr7p4CLVU4NZqk3I5sBaz8NC5OGaRq+ETgfJ
AyycS2LtZBABaisUo6at2iCBytmHHYX5MBStCwU/GgSCbai3cXuIR45mk5nJc1qD
eQ4SaHi2oGE35wqoJhRjRVOO7w4HRmtdaXLfGF9Yci5kBjqdnw2Z7tTbjE9fshw1
Ey/9adwpel7NE40oNjxjGwL90s2iLynOvcHWLLtJ9GFAJ7mwXWJrfENtTyox4Grs
EZKuQkCHJAJvNe8f7PY0wkS94mQbwS4sdFqxE5kY/JhigyvckjETft4XW7NkSrOg
h43eiduRNMC5Hr8VaGoh53ageQpJuP0+QxBva2HVxowlgMhI0NarOeLRsPXp7SIc
FJyVNuqiKe8btAz4W0BWThzOCygGEF1FjgU7uSKFI7S1FRwQn02hhdGmx1ISnorB
EvrAfCrh96z0mRBIHBVMB5PAvrGqhw4zX7be2/8VfuPUlP+b2gruPcCBfxQE0+L1
UE3Q1sK+G7mgK8rI2iMX7YVWznQz0N9FlbbdWSR8Bch/4doCaJlAHHCquEZzszHh
hSJnnwdGzgoYlx2YIh1X30AzpR9cfBxPqFAT+Fb2SXWkrlpE+GU+T8PH/N1pInk5
Qh25WaVL/9B37C11Z5sp+CrUlilx1DoQ8TyAvVV29Gl5DQhYBdODv4ozd0QR7gFt
DiRVCuo0kCBf/Pgrqdj263wM9lEnLDrnoJYNYxCVCczMtpqE+QnmdzfC8w5GENqH
XLdef+4pfu8WLGQgaw4B2y1Rh6OfSyJFYKH5uOBYUlC5wvDpgEvdK4vpb+1gBWR4
lK39LXnU/47vYYEOSg3aPfDopgJk8vaImV3nJ2bpyt7vw1aEfKH4Gu558gH7ZLby
nQqTwqg+g8jfR37VrML6Kp/7wpBVTvog7cD0GgtMBFPHlE8hJ1dX2uwhPonyn81p
agZ01vzBNnSxYagaus1ZKr3AmWJA6gIs4VXCX4Ux/EufSC+RFa3L2v2WBRj6EGa3
KJxJ0Uum2xz6+Rxp6P3f98PyAGzxHg3z0sp7jRIRepruOXbEkEr4C654HT6ZMN7F
124GE8LBddsd8MpShtnkdMNZtngwCulDSq3Jwe7/A86Te5RnT9i4t7LltV/9JiGe
pICRB0r7Nqs62HedEVwfpfxO4OYYSuLwfjJE4VBmJuI7idLvsjnorEpwd58b8NCP
qtLFtAMfsv9iQVelOMWldiVBKPK3mzlrWwI9Ytzs261Rm/+FWhL0R9gv2SmFn6Zn
NAKTdDbaz6EOUpa+FmCqK020Ll9ChwasFkJvDPBFDQIpdVqJU25UeIZ09U5t5hJm
IFckmU/tpudf0QDA4BRc1eYFIj87ASV5XURAIHaJ5TprcTcc5uT5Hik70xNFd7qb
sH3/lA72iVJU7loXU657HqZgmKuGl2HYh3AnY22l89EFhzWUsXTa1bnlrQeOO00h
67wDAqtI2HIVDe4YmUwxs80IJ5CB6a7e5dlLyX+CZAHerNoPRrzlDlfAAuiHsAJr
SSfC6PETcstXTqoxq6BfezmDeFC8tEUraplvRi2VJTUsLG5PDKqt4c2Omtqpi/VN
MK4PbjtitHoztwgKLWO6Y5EP5nan9WJNV7XhOPUIOajsuEd59+3X1YHzk7wwr4oP
cuWrb76rO6SgYIRuZEjEjqbwazivNIs0VTmP/8/LRcsPVaRt1TnFbNo/aCnXhmci
PqKBfp71UkdOwwLveyGM55EBmK7IWC+42WTYlOtWdk6vG8WqfquGtCG9fvRO3WB9
p12ZkErCii4PqtF2cH7duM77ZjW3Ajv0RrOB0GlC/G1jv0Qa4Alq41xao/rtBMds
BkNvyHN4qHsGId6I4RVeAOUtjswDqOyb3nCo288Ol8/LhIOdBnG5/S3mE5PnKUZM
wm5Blm2pYQap8hvblAKvLPfXzGyWp+umYTuet59N4KRZvlBsJKmxZ85C+yhcQloe
vAKUn/x6b3P+PaMNCcxIi0GIFYs5Y1LrGoQzPPfx0vW867YG3eqrbfJ95mJr5lQa
UIobqBz+eunJY6jGd/pHPZrE1IHPS81Ucpv1ZSoRFN93QGq510BP3yPU+s/nxxK/
YLBCJ6jdqsnYkj86xxz5e+mCVX/E1/UBWZVvkhXYktYKIwwuBos1dlNgT7xexeeO
OQ6nlJ+Kmz9VAVxtmLhKnNI3IEEHXXj21sUvJKGEsc4ue3Apxy7MEppLrzJcL0kl
rq3VKI4rFpUv8llM1X4lyCLFnF5S91fpd55punsIwuPgu2+c2pcIU0L54OhyXOl5
L4p3Aq3o52tNT9FfRTi9vJVXFzPNs0Y35Dpb+xeWSs5EZFb8pyJKGdXTXBGcLxWJ
99rU6O7fJUm0/M8BOf4AgdaJ6F71JA2dbHzUQsnhL89IYhkdxsMgxNnJMKvhy2KL
4jYoSTU2jN2EAanxm6uELkFEcsPqLRuufrY5MH3PQGZAmmNUwBikUtaWRak28dRU
VUs/JVyEYToSKDe+FiAnSz0/w/19QufrOXcEiIK1zh0ulTX3gzPVy2LOJcOQOXZD
KRqbl6lP+dtY6QbOlzDPw8f8zAgcdsyk2aLUq1jn+41tTaOSzfraxFyAmCbt1ENB
MLJXhIEpqsbDKu3dXgeA/+VKm02KNNrFl+BgRLDwIWWfwEy0Zv1OcZn9QwvcJc+Q
fF+q9bzvg0n8JIhXnmMWboqZqRBQmvjP3jV0w2mPw+20/v52NcW6ckXCw2y+Exw4
EmC4ZBS8TmOagYaCnISMChhsGhaAnjQ/gkA+kaSllcnLdpkONGlIYVm6JMSdhuLk
MjAIJMFVeqNrRbsdJforRZqmRTYHPBlNTSDYrk/vTp8cV9QuHathFE7NJ7MfhY7U
oYcXkz+JTire8oqOk/K0zb5GDOFOcsDkCvS7iANBi45aLPw4J9i5yQYRNi6JBrbG
UkkQBBOvohJdiXnBp5jMSTmwDNahWEZNSTEV4BNoSBpZHmTyjtAnituYIjpdN7oq
Sd1WGFovIfaYB6Z6g7qbIUt9xV1wltuWBoxEDQPTiT+AhTvBdkBETKquiGTWfAax
UmiqiOi+9XWIKcFGhNC5TkkngeXihpvHmcByXXhNQB7QVktomUsOoCl9gCmIIWE9
h+ud0r+QLoHWdDSC+tp8T8UNoYHV7j1gBw1+j662+vFYw3gANAZlyuK8cfhZ6Ar3
cr2bK2P+YBX0FpFfPZfSN4lHP7NjROjnkAtunIvKPwwI12AQ1e9xkXO4WvcAMsn2
cpuubGVrT4QwDKR4OxCL20vnPKh+jrbU4eFqaYuajTdxlWy9oiNskjDcbGA8Gyqa
jgSQdkBrcIafEG0j6tKtwliN+zIOfYK34Rvbqyl2vu6nN78rB4dAxnx/o/6Tj29a
fUxKXcVSRNhORPEux0l09ckp3icqD04SAM8NWGpKfOZmma3OBLmnvPbLkOL1TrOm
TTN5KTlLQQzfi49KJG+zjZ0gplDcY5MjEEXDgZZWv1NVk62enJC/8IZn4Nj9Ny5s
dy9LIBGQPxcaBxmUCcqRQFBV0actsW8SSHLn45Sh+F5Ne9nibv/+92oFqGNzxeRA
55jgxF2bOH4lbVDf5l9TTHzCg8V+wABuyhwDW4cSm9fxoxDRbO518SKKmHR23Uq7
nnrhqpuba9yZDohGMLPRBypFJFZCDIenKZmuIJ11cXCXr9uENu5j1sgKscMvcjR/
veUd+UxJ7ibMBSMRwxDwip1pzbM8mB9L5bghuRaCFjvZgPdqYrZ9bXLP3d54CKSW
TrLKFPwsMErA/TaOjepjx3fxwKF5L92B21Mf9y5Vb+4sJD7/g8YwmcIxNbm8mC3A
dr22FGiidEGuzz8P1DkWPtXKb/Wrsw4eXXSpZeBgubooU1hHAC8MmPScAtiVsHpD
MwgadpE4KR66FtrHBpywTeb+DIycauGVr3k0k0kNoKBHMU/T3r5QK0xS2mXoDRsm
fmJFxbz1VUK+tvuh3Tu9nQOSmwu9K5snSUb6EKtlz7VeJ+zziMh5RVgxFhmP48UD
7vqaMEbb/V4ERUa3uwvX7HCjFuer625fnwuynQKY+/w7pqDZpStAgpcSkNcGYdKS
uDIb5OS91KB7tWYb402Yaq9KAGCAHYNmT9ivOQCRMspgfp8LwGhcDCcgRsVjIYM3
l5BRsW5lTFW/WdA6aTOQWzQ6nyLwA+pcyjOK8tQmsxemYmSVe3rLOuao9b9mi6Af
fSPZKv9DmCZtTSw8wAbRBE6xKEIE4dIfkZ3CQFaJS07Fg/w2VMGZJt9B+Cfxn3aB
/rwdxEcXMa5DNBeLKf1JfnL9Sa/guF7mLrvpFmDuynLtNnZa0c2VXCRXPDpo1149
X0l0oQiJBG0vYmjZut3D9PMj6VPcUPjab9otyFj5YlKpnE0ZpNagvnVO+opfnCQu
KAym73k1YebTKFRUGzhrktjxUgRJOFjRWFgJmgztxViB4OHa7+t761IT5+0ase0G
loLHnyRAu1JfK4Xpw9SApgx38nskQ56MyU8J/N6buyN0qDJtbNDS4TQtxbqgQbFC
Cic8FrbGNCwZ+Wxh2OlvlkHiUhuxxdn0gATIcdF02AHtm61dFy92eMftHl2pwvqY
KlJaPKhJ551qoJ+ScPs8X65kLuZibn3Lc03sPeeVTAHB/vVwE+Xa8SPkpNU3HHts
efbR0myvgA/o8yxsiK6lo5fT3gD2sufUZM0ckntkmOqOJizBGEkuOLUkFotp+FDB
0CBGowU6Mv8UuCMByZZGvyKQ4Ik9IdX8CYmxCj7g5Q77KAf/JeRvvFUt6C9z8hQp
RqsUjSZVVmWD1kIOyAJbs5eqkDQZiqOp+bjB7JVmh4njAu2oWd0dGBYW8RR96OYX
vBbop9yKn7cB4fQOI6WwueJS687JOrzgxPRGt5P1/Y71ovWaE9khvb2BkqSKWGrA
vZdABrAQLvQnbf7F3svU4WkKmykIT6ucqKW08Wi6jkg8EqqNTaaqbnLMQFYTAFt4
s4zVRWcYoHOsfbDwGC1zrQY4H+YeQi/tUTim+PaNepqhz4BKwTGQ/bOVFM/vBgHX
EkilLq+ut+riiT/h2X1gOk5+OHVxTUEIs9VBx1Q3vwwYuzIRnIKxbY1QZWpHEnc8
xBKiyTDIKiMW9RWYjfSM47zRZzt1MVygbctNprf+dajX/rDqHxEPzfjdWOiRQIb9
m2i1WorB39unzZVIcg3cImxQJn/M22gJwCRLIT6/iQS6PqMoELxMkiyAVsOscj1b
2r+IE64fqdkyu0JWuCw0i1mSvlVZXltW4vGgVFR21Ktsw166LgiNMO11U3KKoxo2
VDqK32psAO+rkVWkhR+Eu219tEcR7tIAwlCZeE9/2hM5wH9rZpbUSlrsYoH8h405
HXQBmAHU8ws/VU8y1zKu5pocQT34irxIilIID4I6JdSGhheKrqzGMubvd0WmkUJH
ymb76Nf10TZymr96bBaHE08JInfTkfeZj3+0M2/pF+oC4xqmnSdKQhVWVg/x1Luq
5wClWbFBz61Z/lQyVnwZp4p9tSpscXM2uTmNoTKOv5xaubQLMjcA7/ICOTFAnIxf
g3KMSttQCzThv1krN4N8irh2WBnDelH43ZoOyysVQI0hSDGkEQdKjfJmFehNHHMj
z6f9463+sUA4nE+7up9bPKCHhWX+LFZ+aSFCuAe0sY8sE6Q90XQ7L7kjtUstrQ1+
v4o5RPpgpyQqE8lAHa1cM7lDGMmQxW94lJFgRCxY7hnG3LWq3apT12FTYUXgqtqG
3Dqoi+SGA45jkbwXV4otKEu1zXKteseBPIV1fRzzWTurm8ujRP9/A+vHVJCyph5/
7pZikxAVRM7XnYfoQAqNaNBivL90Z2uBPXqp5bumfpUUsvUxxVU884ZZFwxmNneU
HP573wIFVsOwi6K8cGzEPYiRNXj7t4fV+UtGEMDhYGwvSPPCd/akXLlS0SH5zkII
xdSyWpGg31VU0UrEjkqrHyutFBnwxn8NMrv+3hXAz9IllqfnjGcQg2hbl8BlO8hK
mHuwnXO+6sMO82MtLUnSzn7DniNeK9gH5NvwjbqBr6naLhpIa0gFwu1Lz1raWCGY
N6wL4hwwUGw2EKrAjy4m8DW+h22v0s48AU5xj89WzuYt1yPQiJrjpNxEWUnEm4cj
ip8cpyz4IXHl7qZb3z7MBar0A9YgFN2rjZPXpQN7gy5JVQSINYbI7/XKPpe81jtj
vHr2REIuiWDg63cf6z651xnrq1wK7tJhqNdJ+iSQc3h78xIKXmLHXsFmUMBd3x46
2pqrnGWIhdZQa11hLIn0dBb1b6DA0FtOMlNVqtJ1+ZRWddiWGoWbGPPnFKSUDdJE
uNUrLBNZV35aKbZbmI/PL2a/KjUbk8OWp3s5uzVWvJBwjjeVPneE7vfktNKfz7OA
Iiu6nr2IGVpeOKljHNknq5Msvi8SJd23DBwnsyjptLm2z38OpCDf+upFTGtH2x61
201/wGUrmm75Btpc+/5OIQ1p1EOAPCYtXcf8jd8qPGtOPHjTLUT1wrY7NIm72MDX
ZnxXsXRbZy9E5YOk8S0pQfG9IU5ohX0i1ahwTeg11fBZmMFamVGi75SWaKyWrIW6
DYzyIW2iUTbselxZmB3dNrPqPzUlW1LLnn3jt7Q6Xzhyk7C6pEGHiV4sCCsNuzYm
uwbo/11Xfp51TDNHNi/gfZUHgR/hMUAMI2hL+2q3L/OdvsM/kiz/2DJewrHJ7zWI
zkjhRonke4+bO7MdG0kOwk6NfTzobO/gGBH9sLuZ4jIZaLnXA/4nFENYKKgnIzTN
GYkG+5E+32yl70rPcyErcGttK0M1BfxzWnnSWPIyWuje5+F8E3QzNrYtwMOo99+y
i9p7nPLwRRlIqZiyt8lki6VWq6StoJI2MbpF2Knjktq2UHySUJMwFwSnTPBeFcz7
oRUQduWi34hgfiDR6Z8MJx16UH050DTG958q9pvsmQVMcJ4Ossj9vS5XMYfUcufm
0TdYnCZOSZWbA2LblJF0QnBHLWw+KY3IFPVKA29xvq8yn8oRu6zS1cP7taaBCcJ5
jhoEqUcW4jU+okifg8QAo2ziFt3La4R4+EcwgG8NqYwweBvpqU7UcfopCSukGgCh
9FjIpea0K2dM9TqP2KFi4cHoRgl7f+QNHIN3xkyZCb5DySMi0hpMgMIJjzvBN1Iy
B/04IW+cdcfRwGePA5p4o2G9ICKwmF6uSiWDmF0KBwHaWVWzIsEU56TSsm6VLyA3
i2DQzSTa5wKVYIMqFmQUSux82gaCdDZT2xLcjbujD4hNkK5jvxI8dl4SWtj/9bDa
xaEtNd6Mt+uFJM21eDKSIuyPIELRb7eNGQPVgG+AkMXJB6ygna/7KRlPwPiYZL+X
e7h6CIr1qDp+aJiHT47fWqHSBsSp/OIyD2epeXDE8Hc/uAIdo5EizAWD6F3MEjaW
uL4L9cdkQo3Cw1MGGxs88+bmhWyWunkZG9OhT1FcuOsEafXVRL/yFQ/VTSXa50WX
6EplxlVgut1GgC7SkGkC8op3EgL1CEdn6iZg6hsJDqbBzSLy+RsTvVUflhPdstS+
PSky7Y5yPfGPCHTpiiePtiwb/dZlPP0UFZxl18xOVO2ayeu2pz75+KsNz+EFXgQb
SM2vLlYIf4GZ3wKH7jYFdJIrRTktDE6ox9znlgvC+xUwZiIsvVtN/kN12dhpQmdW
+idBHJ536cRopVSEQlpHqaB9H3ORMtx/fPiG+vdtr6SRD9Cwxpsx2UGOY46U3QFU
szVOd1gtW/6SgSQV8BZuCGsUwEvIiJKpDmVkU0JWPGqeGdQYRvjitEEmqyMtbB8x
z3xfIsqWZj5ill4FJ1zDyMv69HI2Zz2KRiQSXXO0EHF+X3WdZeJ2PAv4Ybn1BWbM
TLoE12nOHmObDcOiJpNQgBdh6XBagiml3TNBMDwS4MoeNGcS/CRhE/sTboZs4vOX
fmW6UNCVqICedjcGugYNQ6ezXpicMRZhslYEY3q9C8d1pWdoUWLGzlA060+3Q9Re
qvRVSy3WI3Hg4O+5VA4ze1dSCW6/2Ra1JHzJOqU4tk0aaevExsQYhY325XpatbiS
shO4/fZk3vHfxOE73RiYzrqPZJxPn9uaHB8sd3ieS3zYs3JgAhyp2PHD2yPSjemB
sNTvzPz9j1eJCB747H0A0uJw4jFZHGsWEkwqNpEX8pzYNSexVKeYOkU2NNIu9aC4
yYBEma3AGXKu/fgb4kcv6Y8w6A2YQS6hVe8Jap55vX9xDlcEZQAqCG5+QReb84eR
7WERDZAoePQj25P8SDZwLdP9cag2cvNmHr2DPYFTUEcycDb9o7pHFNZmC4GnAfBx
wGFaFKUtE5mFuLuxztuORZEEmHJIINVwpLODEUhQJfAXl1/BPyvkE+mPfDEIOVAH
sP2hQxKDYLP/e86J96PovP/i2134Lmog3S/l2hdjEQ2cks0B8qhGEf/Wg4LsEXH2
JVy61XYYmtcMjUheA5LZ1MnlvNYJCshbbAQeDf9kKCkMC6rUteD68G8gBxigJf3a
yN2DKOclvBjBNLh7J2qtq+YBNFuD9BToQvN/S4lWcxXT8udhKR85FeA0h8c+O6Rp
tqjUn7vp7zycBfi6eNX19Km0l30jnGCmbSO4pWoxOpR8NJXLfve78fcRpyF9a/n/
g/NQZ/MJ8tpPG6Q38wTUedcRaC5Fjh8sst8hBzqfgS+WrfR7NIl4u2RvVBWWfRhc
7gnDRUm/QhXt0SHXui7zwH/t9PbzaVTSExNJifBjW7c/D06OTTdwzV3UKFF1eYhS
U03YFe1zCEIoksppqaNOIfplsHLoTBwUQQy75COAgM6Q2WV8TAj9gXFQCOFwF5aa
8diaS4AHc9huFIXaT55bo1aCAV1UqZliKohGRRUgLUMIYn2X3VweYH1jkYqN0BjM
eJV3cKp0r5JwQUinoi6+HeCBBh5NXyACaKLt537ED4a/ZBXN4AosC38EzYokgtO/
YLbsFbhkzv7/75Wo+LE/YjqvmaAQIx2T4YzuCc0mCqVrIrwwJAveBfmjHFImKvjH
ntu2a59G0bBWtNgF0Vs8pSIf3HtWSDpx6nLSxIwErFu2BUUjHfSA3OusXwcTi6Ny
8jGtAcL23CFBFFdlhTQOLMaInivONrqgUNLnVoudGl8ywO+4Ti4bZRGaeOPA4baD
rg/xbNmZ4RRE8Wjp161B8BEC1t1Zr89udxzPyZwN8aM7r8N9THRutUe4rKmYuMbg
raoTY4gMmrCl/8qJjF6iv30J5u7pTJPH1Yi5x/L0laTCCq6wWgpVomrU2KcrKra1
JIDPM2UiRw8Jk7V24VjTF7IrQYjsWqIcJrsB7Frk03YO6ldQkbgz/m3EogKSfvLA
GZnAOuqfCZKsavhk0SubM/tjMM/oKzWl9R/YsBCqOh6GHcsiE1dPvVZ+qV3b75mV
OUQiF9dNdgJoIK6LNVDWeE733KG1ye08wv5a9G5i8q/qibaOibBHVPdaVCw0VEKQ
1E+vhM927JdWdxXDLk1hSg24wDwJBAGkux+vJ/v99izpR14u2Z9uA8yXe8vtg/YQ
+9C91CBbvTd7ctMNyL6a4HoA14dafisKRFqvYgRJs1PTC7vXWCUI4m89LePLEBQj
dED9b39bcJKhDeZyJTYVMc9sDQsH05iEXe4VszW6EXHcdQB4ZNVFJezZnvKHg4WW
jUc5JOLni+yPvXXZYfJztDTjrteoSlmJTPFXCe8tsKCPmIQZ6lvZHiXN1J76LyLG
ycKcYXAW98tPBUuUlo4FHVZAE1dDySvgaMbduR5RHgA10q11Ig1srPBpxtdSneh7
7uf8sRmwMFuNJHFmgbuULTcudRjoTqU/kurzfP/tZ+wjKhG11oKBxx3iDeXHHRCf
+7BoleN25PJigjeijUU9nUQSFGKQ6w4Yp3p9xZCXvzAuzu8XMKTSmWQz2n2MVu0q
JFvdVqL0et5EOdVn3sFuwK1n4ILTHsXkRz0PLpStBmoYeeBMkZIdSPD0/Q+CrbK1
aZfAAdHgVUKidHOPAPuTK2g0KC7EeBRjUx4wvdBfFhV0emRBGR30Ic70/7WcRKhH
hqYkKRXKk+REZO3vGPGAJBwRwX3yDtq+8I86Voo+a77FABltknIqPLQ0jeIOZdp1
VT/P4elCx38ILiiw6b+fpQc3JHUktogLnHNKB6Cg3nIjHUfs9FtHl0NO6fzX/3w3
yswi4wRf51u6u/irg2VyqabYmhWYjbe1iCJ1dQVkW4nxZPtVD9AxOxUDv2pVfYs5
wMou5JW6M5p80JxkhHjSRyZtdJE/UkfUjTr0/bvBLdFx9fZZN36Q/JBJSDEE15hZ
B2cq5gt/IH7aSmN2QQHJ1Sowxa4k1nFuM3cyuoPZMWjWMmqM/VrTUM/HNbMhtzgz
r8057AF64qr6FIXsX+AUfRi5Ntmgd9mBkTUCmBcpAbh0w77Hgp4Zo0Dg7j2erEZz
E2rappYV302Fni88/1Ouy2LyxcfJXuKo/Q2XZybR4XAabDbm3IBFeflsUQnWRUiM
nzaI8HRMKxd+sc9EKeH3tgOne8heu1XOdKGHZ/Ofa0IOZv2RbFu2oyg+qb23Ap3K
ktHBE95uu0qh34tEneh1sBsp1mTYCP2L+sFMbYb85sxEt1kGvXaAGYR/BzC7Td1b
d/q0RQ+4quRtHRESmfNmpnY6DdxNv6Wcle8OVMPbyt8TdW/ZpWX8zurevOgNf5HJ
QdhJpI4pl0V4WYY77FMhyHAP7qIoYyHlYlPhrmuUuWMFPsoILDv90XIIkj3NlC7Y
vEFT4pO7HZ0nBbfe+7LisMtyoMsmFKT7XlMITi4ev/m+XQj24mixvTGBWHFZrLck
t2at8l+4pbMe9WGcBJxJUqmXAMJ0GRhTNGL7jMNyfFs9352bnf1tqlITnBdFQkdF
PsYL7QNC2vsZEDKbIYWHGkY6Dkc+lhq+7MNyPPhXjH/qK6r/7EquozKiQgOcD4BS
IlTkEn9HAuvlbqSBPXgA71U+8FAMw9vl7ElIzV1FrA+SfiOB7+gcXUpk1/+yQoUQ
kDK40p5g12l/zaDiMNcne2UpXJGPNuNhqAp/dGe2hbMg3qcymujLr0lCVYZf58n8
Ap4ZBjv/VJ9id9nKjgqH9fTHvvGjQC3sk99G28zWAOBqBHBVqYzMQybe1q0ZBdec
MgMngycJmjdCj2NMvr7oZxcnQNTyUAnJSSLxCOULetCG1fkzvXfUjeJrm/9mjbd9
vXSr45oRULa3aYEd0kDwEw3rzT5TSOQM6KFxNt98LP1yryI9WTNA1TphqoMC8huA
hWDoXo5fAWgxUJ6oQ6eZt4SywLIXSb/PolsKhTIHO1CYc0oXDL3BOJQFIuRb0imz
vpmLuvh6w5TqTZBbBFTZKvaYhw2BZmOgO6P3hdyVPQJPjZ+4VSeT5LFrszxgeiIX
LzDt10DRymvRBCVsaNSVf9qc2vjFpRykoVub5nE6URtZcYsFEEKPbpk0kOcw1BJk
pohsY+cIHIHYAMRw7zt9smbPtMzk3vSxV9B1QCDvHkOfOkYVYm1EyMHoXmOYGKkX
raoYHFEoAT4mSoq0k6Y67dAV8/loz+tnpgoGyuxHoCPKtZHboLXEa62BAaCrgfNs
mxCF1uhUdLh1AaPKB0ofBzQ7G+U8C8UXhCSPJFHMIodkYD07csSSjXzk/Rk4qJ3x
aXoT+WLby3vo+mKW/1fQRvQ3qCCwDLcd1Z7ugCbHfjFJixciLjMsd930iI40iMLk
9zLqhBM6SoUx1TqtQqLzOhf7WE20PRuhSmrFbkpp1GMrdjuDsdHKFf3MNhf4ES/0
P5sVVF3tixWVcKTrl7axnMf7Jl61fbdb4bnxtB68qBm+9t8As81cpx+prNByKRKY
Thgx+9HiLp38Avl6vBz9wPxDQigmh9kCt/BvVBrF6I3VYzLo8xQn6O5TcdDLKQAw
qYRH+ZPn8XSR7nuR56oa5PMNkBcwfJEobt0e7KX4WpRq15eZLG59rsQQSMu1D0rN
GicMH+PuwOs33GS0F6ZMwguD6QYybloxmv2gsUOdmN1Hn/n4bmZ4nroF6R0LQRqq
+gl7AjOTFWLbEFUvHRq9GzAE992fcc+9A8TRaITdn/QQF+qMQBxQ0OYUsSco9nn6
g4Q8khygjmt+mW5EbGlGuVxiPTHrP5psJopRav5Nwgz9jioAZpJoGno94M3B1Erd
FcKm5PJDHM3ZZ/bzGVG5KCLpgFqLJsjZ+zP9Jrz1WgxFOBZoQPMY5ZAhQdqvCpYQ
6cgEzUzJzTuo2OCNSZIe5sDZSYhAHLE7zRvDCEFMuAbcjP6CCUSHzTJ9fcLESLxq
II8S/PZMs8NTrzUdjVyxGHMewl5ig8MgixSkxmZSr+2s5r5M/W6a+LPij0RWAK2G
B0VwuWj1M9Zfq3Yx/8MpafnJmaSIaARzTMJFBY420XrbFIJ+8ilfeAh5YHkoqAZJ
zPMFirSdZcnarIbwMI5aIY93/koWZPr7E1JpXTedbaviVaJf/+MNPQdxiYyey6fN
I24u7PziAhp/yLQA0EYUJA6VZ3DmDRIu7ELjLOWlLR638VX/LF+3KwlHFM5bibIS
5WjnmtyMd6mCWcZSQYkYrCtqZClbVcZHtT2pHx8tYX2g2D+LV9tOwT/D8TtZukR2
v8SOBFwNYSdgONm7c/quLKwzWWAi8+QRAdroTu85bRdC22Y9/cks5oU0ebEziEg2
DXxSC5+RpxK450bXLxicMUKPSKiKCMuMz6Fq26eC+zoYT5rFIydc5jLAk/LWsFNc
0n8OAD1T6yq42PcGZpo9mGPos84ffm6juSLh5jEWReDdsuIQfXkZ2Vrha045ma6Y
Hh6x3eJYM3932JnYFAdHWWS0N+uScPieNX6zyAnSqLS+H5sLoeznjgWH7TZQHHXA
sN1dz0e140U/Rhp0XjVV/5Ep9UWNhGsK8fcffVOFwDHg/FXaIZwCmWnB8VlwPic0
hRd2zIaodtMVmPkSX0jQdq6qdggrYna5qXayRs3OIwt/iNP0gX/zbQXXcyBs617/
Eo5DOOHZUj/G6uWXHRi8hgRA56vtzVv9lOfbXhbEv6U+T9IzGt0ew4NCSka6fR+J
foVgl6dVeuGAuYsShbcf9ezL85EyTNQI4QNrkfEF/u/zC0azfKiLJZ4y/ZwDHL4D
ae+gCKcMjLJgS2uId6QbAJKQ2XkGuuKBQEYBiMWHeKAsxOanuI6VvNwX7EnhTgBa
NrmiqsWPm5nS6SkuOsD5+DobZ5Iwkk5P2iG7Td3dTler02pW7XXZRs4bSe6tIPwG
OQDouRhjrOEDR44hSiVn/uWj1KbrY7aG4ABj14XcbrWSiUM0NtMSmUuQ7+kxKHwa
hutBl8+yHN6GpN5tF8+nLagByWE3EciKBOiIFI1EQs5KiP2Cgj/8/YHqxlcTUqm7
wDb8IvN5OwljJm1//+twt0nktrstVOh1nFklsIXyR/FwxKl7Gh1PeD/Ng1siGLmA
ZjEOmkeBUIDPhUef+jHGC5BGGqXo8snWT3K8x7+5msm2cHA2tO02cZM7uutkViH3
KwhU6FXNVmXOMDJ0+Cz65xnr5mep2VORe+o9oAMwB2vHO+78/6wDFLDtScwC9Uyi
IWOOo+SkLJlAOi7r8P/aLw8/eMfiNmqdSjvMJOq31QoMjDkUbCIYztulADfbYCIf
GzJFDbnWiDYZPioo5rzoSgaw+4C1yenKwicIgQfP8mKNuanuNSaQrb8mc7FVcNoZ
+dHdvb45Z9oj8PA5QgWewxMnsPY8wyn41A57bi7q2+Exsz78a6E26SgA/YM4VFCH
OfNpEGCzOA7WebgYm+WNEfyqB5+fsdCekVjsSsmvK1PXcSAo9+NxV0acvpJrsyz7
WfhACClT3BbMCrhJs58pB/ChdjGj9oCH0cYlQ81IhTwBaQVkNX2XZpUVwy38ex7n
69uqTNhyqKYau+c/dXjQciAORAG5T2Qc7PA/CT/HszHtBZk5kVPYVFe4bFs+O27V
axpD6PjbUOWVzopalGgwcklMXh9EJN95pTiSoRzhWf3m4nPzO92P1iybXaMfWvA8
2AmQGugTxNl+5FqLBgFSH1qISFAD8wMxVTjumCgEsK6HS3RylpZ4g5Rq1WDfxFfh
Tbcs7dZOz3+VFySNZdI7bCjDu/uvaPfhL4Qh4ocXqyumWtoP0NSZL7d+4HcRYDbb
bwqbxAHqYh9rsQo5cUvMQrH6EXdpYnbchSEEu4hCgACghLa1dIS8LT4t5DRKw7qp
x1NywGL7U4vpFLzIw/qsmJI/6fLE4sg06GnC32EbyQTkYfeGK0tsKCsStEbNXb5i
1rqNEo0RH68PZ5a86wZQSoyAYW4E3CUb5KEYXWe4Nf8Nc1+dAtEpuwxDg+c9OKFu
7hNS2tlyrJ/6vQKT7a9Nr4lJqVSEREk+FNfpyNjoLhH+AELtNTauJGsomvkhjAc+
ZbtdWrUTORTqAec44OzzURE37Fq+E+lGAodvUVecW+nFys1iQGlJhpVDgz1HT+xV
6uDy1eW4E3daChnGmk1Q82b7QkgKTRwZBDMJ7T1EsCWWmsC8xie3MZKc/ANnFFrM
CqrOpG6OK/YQW8dkFyz27IvNogOOZneahRqhKnoy/kVha1pP+3z3w+yonwK53uYS
5ZO3GKG0f2CWEiJdWE7uCAwDiCrdZFHphvBe9T8TUv0uT7gj64p6H7EllcIHeJmf
63639JD10tzWJ52s7FjKvn5iTNT4f9F5Fd21BxGmBIBjofguz2837Z38w0f73nuV
CfSgrcg28ZMa0nNM8UFufn0uXfYLssnGAeuXKGvRUOnWjfpIx6qBliEyVhm3M0j9
WeiCn0GoQDCCkWdZngcjQmW7JNDWboGRu8fkAlbHvBz1SBmR24pHWVN0TDpPJAtJ
uaZiugRvoFtiyeHXpEevJuQ5Hbt7GqbZbe35KjAYjJfAtluB/YWXu05wpX5Mc5Mf
PN3Gzruor2qL2c3RE2eu/HRzVE5kCt5/TpFP05NiT7cUsrnj9X/mEvMoB/5me/qM
9JJwPMK8ksM3kCPfSxFnGol6gahPtx340C22bK2flCxEihjzn2+01+TClb2cjFIB
sCvMw4LXCs1zIUcS8hxRoxp+oHhj4oLHB6bdGQWeIXWrQ2e+AazTDxBxtyWCtFqn
8t96v1g/RNUJKFHmwMwnNIPOaba/f593oYFrKyvyfvdL953Xi50gUoSCrZ/uZSv4
ZTWMKOTfE/SES3VMnI5byaidbBy90uodOo0gQQigJ2Ptosj67Nmp8m9xrn43VY0b
KKjqHctIrMezp0EBCYL3cidcb7eHocTkE+uTj0AjaUCVSp80tU1r7ZH4IZ5qEeR1
Cav4fa1wXsSbtZTn1pN4GpjMuB53nJCMOfPXQM10R0pxyJHHNiB1eFkgaQG69aVf
GlUEPUYvcB17P7i7NiWc3K1blctRc6ZQz2iEFSYazqKzlV30rZYdRkyuOTCEJ5s3
Al7bVGzM2h4O2fu5rxKtl41GX048Ll0B3++nFmka1H4YBuHgLDTrSHfEt8/TNNag
Y4WdvQr22XapCLRzc8LvXzskhEMDaZfMq7ehFUxxv/k7NOtACaV6H3HzKKhYoP8k
3RuwPX5H3p+q3+7uFbbuOnWtgNY7oWWuipBsnhOBbB0nzlblnv9+akolz/y8p1Ze
2Axcyh8PsX8prEFpHOEFXAGBc9yRuZ96RtrVhut/Ujgqxg7RM9BOs7CLilbSy+Eh
BDlhUxPfY23VynlGEv8hzohy6I06uDXei7vLVo0BTxrlDNjhrJjzgkQY+S89btZB
maRZ5Zk1gKgq5Ln3DSnlx/3xJ+cDOBvJoeWneMT+HYfJz5vhusws7PfKQJGqwUOL
zCoRDTMJ6CcpwDJ5OKs13itb1PpeZpk5XBVtfWYFMSJyYe5USxx2867RFmon+ax8
+4LpgXN52H209wRnhACigkYXMzWMYsRSB4xeVZj8PPPTTUpgERtop074DFzY3ZRc
+KxywJuw64DLyNPHjFeKEnPn1Ye/OwLjKj+ZuDppP1bUD19q8OioCOReFNhhisx5
WfvMZWZqH4Wk+xTrShVkMiiLsEYFCkPwU3Uh4/OyrW18AcyiKReFRzq1CQv+j0x4
bxptjuX6AXDlFE66nxjBBH1upstzy4ix9h1qfDf9ExorE7/OBYXUGRpZivHpHaQr
uMqE7qnNhKT2f9jEB6qjLsvPfDoy33AVA8GzsVyVcgLzVarEc3hg81KbalPngBTe
4k97XGezXul1Ft7fEJvTDwCqBEI3FTozUXpSp+CGBpZhyQjlVAO3pCPwWMx9jCHp
ZKPIovDQa0vh0r4yqzxMtiOYsdov6lHKLcDBg+8GDVhvVwGsrYUyzUm2nOUvOjRX
ikLoPQ6Rj8O8c5ZP6OZ5TUgo5WmG4CwuAw7sV1nb57b5ocXFUSdfpMg6HqCMh8W5
Mbxczi7wHX8FtVCAZg8WjuQxf+Cev2M95Xh0YwsKmGqM1HODG6M6yG8tIKCHWhEe
PerX+s7j8BSWaQJ0mEtfjmEKv5IhMZ+dOaNDRYkrO6a4ewtGoadMX0Y1HT6BRJ1D
k5SKZbGsJf8duWHQo7TDu7T14OyYcwmKVltpVMiqRlI03irTUxOn2ZM6QlXt+P24
6Ll4yksjvUG+2hlNR6JaM7po07rUF+ApG1NvOCEA9JIAsIWa+BlGp41Lf0wpAQ94
bTA4h7BdvQnYXb47YK0IIMKP7KtTAcwJ558P4Zs4z1LPk4SwN0PTgvqZit+19EoH
QQjvFOXpRKusSOc8sX0J3xV2ixcsVlVH+SnmsGXe9anDFSmOtJjlVwpb+7TTOffm
HRGEtzymYK5bUVq8+wmPEsFTZZeusnyiJKcmKRXjsdPHRldVfA3GMQR3Auo+L8P0
OZwpVR3z2+N/Fr5sOw9oDVD4FarR/rakpAozyxA/mPo6OyLMO898atQiWUZvOuwQ
xirFncAnB3Tm9TW+c5BRh0jWWr9mlgxyluHmpS8MutGrgal9Agg6o5OkodjcSH7E
QdMWcjpOhM8y9YhOmnP40Y8QQ2H8WWxQnCZWz0ubRoGyc6Xo93C5YiN8d1X3WBoW
bmGF/BdULrxm3VWgLhUzyh+enZkF+RnXw+5egk4CwgH9U4usm8up91ddlcBSLD4g
8pL8M/2378liiheNhxqrnAlwo3BUcZ+JXWEnwDZWFSsDkmRuCt6ww6H0AxRnOmZ4
NhEgwH+zKx5n9gJh6JaSXWRTmh3hCwh5McH1dKVZl5JkGvN9XNnjzLP5YJrBZIXo
NBZHcfklTiZ60iLtqam8vGFk4Qt+qN70SC8RfO4tx+WiaK7uXZri+6Ql5PCQKkHW
b8JleHbyRiJSwvGEJhhvczkUNSvXvplsEfPrmbtTrBNuZhZyWY4W1QWb/QYTem+G
ayzDVwV4E0t2NuFTqaGi0S8njgZp9bdzA6BU6KRmbq7mSLUrudrPDM8UZ3JiDdtY
nxCbM3MsIZtRbpIWx5Bu24hOb1SZRJEMC0HAqhCxMEWrAsrFucNUxhFQC2/ZMcSf
7SLs2/6QCNsqCQvLIFEA14khM/oW9QIYr3IpmcIliN+rkY0XTOM9eThTT2f38Z16
cJuLaUOVFgAbQDPR890Kakudfqb34hJRm9/AW5F1MpPa4O0FpHfKa4wXB+OFCHEs
JX8XEF/X62uW3Xz9+Cl6rx2ljNbvDlH7q/hfe3p2Z9Nib1aF2hbl2Hb3yghUcX1Z
DtZDIwIc2t8FdgxEdkXNqPZdSYPKwMs+XUyktzMpEi6euN+iYtuCF813Dav9n14G
3Y9ybWVfgDkodfFl/tV59bxoP2AO/1Yl8MKJJZCQbdDSgS2TwXQbFBmIVvQOpNit
8tzWsdkph9PtaLv4QTCPu/Zzf5hIXkBKb/gWqDNcltRba5eVPU1GLKv+/m0pwE9x
UUph7FK6PyqjMqIiGRWuKzBe3pt1rblS/DdtyD5Jy4iXBOj9SScl95OTvr5XNE3E
KW3isuyQ6fTINqbqKNVzJUvu8VZ9f7HqWxw1RXERKPTLjPx5k+46v2TIDw7pGKR1
1XwkiYDH4/nHd9xsenzwOUSV4vS2W64ZaTDLqvslA6KlcHEi8DLAAOflEwITgUhz
5uw/p9w6R57WCm4SrNTu25aeHIAKogpjWNOuNLLISiAxeaVpPHzq1UIt0mYD02IP
4TE9Ruo6d3dSqyEktHdz376zzx02DGLr5B+OzV1POl3iu4rJDBeliwvPhrzrqlOX
a/Z9jFrgQCbXKnxkun76K4yBFzmUSYTGYfWvlaKsVrrJedjPSNQ2eqKW/yy6eOG7
Am/nHuRnmvtVPGAYXfu/SNHfLwbXpQ5cJ+4gioRPGWttVIfdBkOaIcu+LUYYMZGz
qF1OfMXZiApf43Poh8b4Fl0OhL9505O9fe+lGzbImc34Og5lP08R8U3HXSMVK2PW
z0F0TA5vM3ywRynFb6gjNNe+dut1l9C3uNp8gBzQQ1ib3fmX4FLcq6/9KBEjPsB1
RjdcXfm5XeTstOPEkW3z5bprSNNLd98kpbs7Pl0WFFkulAWj8s3qXB0DeW4+A8vv
VHzdFiBYTS4tpwoLYfvv0tzKd+hchnRe1GEIQOJ0cbvPfGxUagScftWuDAqORywF
lTMieQYaWTIiYm1EnkJPxIfaO5jMTO5/5my3ILpqEjx7xMJtk0dtps/uyh+jjsaH
eZJKWfB1x+8b498RcgskR3FL9KMPVuGLv5fSbFfJQ3mWDi9qb6aON9Zu8NAHlx4W
xeO3I04MilVzOM3sNEywG33QzVvVNM0rNfPrhY2wxyZAjG3QVOOUB0WFseYb/a0m
MxV95vqMNXSkipqbW5E1tnRDS1k2HchPnGLlooSJXRyzip/pVB5C6+KeG04cAR2p
CYhrR8JlF9bZORfjmDx+2J8PqeLOYdjYvidg7rHhhs6mB4inZXuEG1pQ9pN9zvuZ
Y8VC3s2LX1LwGOUCrA5dJy4mtUM00GS3k2uJqmSrr8PbwCBlQT6zMjg64/QzNF/l
vdLCDpiFy7M7mxuTBLqXPsfjT+hTz5S4BFMURJzHZQN/i2fYlKz2UhLy1wY4v1xV
NW7tRRuUgyO4VyMiSPVPYAkEUm2RTD61k1HFxECVVGkX6HF06BCkd6MiauxLi8TM
g6NqmASD7v7xeSw8G1z8lWFVUsqkliCfxQNahM5VIxpRG+pniEZFzDx7rqM4Fj7m
AfFKg6QqsTgt0169xMuxf23BXetzDSZfAQWQFxO3ieWUlbl13o3+FSHu8ZAUVy6s
pX3qWgOZIeapFdA5ZC8lfdpG1c75Bm1Su6C7HZ2hcnYmB3gCl2PzuM+C8VnJkidq
FTaR7DSAj06+8gGrLaWP/YjtllJ+tPFb5F9NEX7AG4JbSKDyrFqLfbjjs+2vqieJ
V2RyIcrlXaDsO9xRBzu84AQQEqAzIayvC9a8qi2Aeo7Iksj11Y8wJRgsNS5H90Nd
vBnKRm2gSui++PLL29RfqC53qco/zzKiFRlL4hXam9uMCXzub/iQm7n3K//FX1eX
InEt1mdbtE+hatQXI2MZ/e0MJ2p3i3706WzrjD5jbu92WUgTkj3Xio9ESdGZTAbW
6QL0ftTEt+a26Gin2T+XnXZ1nFSN4Sy7LAEi+M1IPaqqMTRud0MDtyCyvqJXKqYa
qTFBcWj11vDcggeSeWDSkOI2PpeVxFPaT9xDvNjLsb73UOyFsxMIH+TqI8wqz9+Z
trK9lf7pIGdljdTQ6L2kZ+TWfGGCZMCuFSadllTp+HibdcdZ4IW8lBZ8kEbye87m
ZxrppWwo393UXTDGRUuVID6TxmVrSYSSxXPV9H5gSjLwd+ouqfz468D9IqtSMMJY
b5u/pXFDXr/HrZok5DcchlqKsSvFRbntYF+eouL2jfPIXM/xvst6PdVj/aELuHPc
XihW01R/NA3uHdrrNtuMyBiAEo6WKaqMDM1HeJgXz6S3eZt8SxapE+MaSffGKqK4
7CvLwzYa3/HqmhTfKMVlnpDI4xLzVwgq9C25DPW9PKgyHGZ5fakruUqlGZ4Rzeuj
h535F0El4mDHZ2f4uB/5qtyGaNYMQEIPkQ3iZndhpgxqX4nMgvjcbckWFesw2GEc
/VNwTOptGz424jglcnBv81Go7v0476ffJ6auC+SAiVT7BiGTlkR0m1qXVKPrl5qu
pRKqpkYGOG11QMNWkBvU/JMLxSQOMP1EVe8s8yxEHHpX13TRpF2epqmSuKK7ThKx
nUOMqOlr4o9faGGFeXZFyXTW/v69DQGyXO9Mr4KOPgUbkmgybKUoDUtfg2sAK4lL
Scju+E8ruqBJ6hpNbvscXJhtKco8pHAWQ/F5cJD4ONFmyaI3Yvqg4Tm16/fioSmq
MaMq4etFJ7yWuYadl1op5UTWqEy/LoQrhlfUY1P3GjaKEtmfSbIXxKd/Z765Xnh+
xl5QsjQEi9ILb4wn782PvUGseDzt1cu0zrEbAAFVGF52WsWWixLelUW8MZK6RqYn
qlGpYhjhAvSpvHV3k4HMz9WZFRHbrE6+mWM3hW8ebsawSAlibR6HN2NyPoID5z+g
byfezoaHAbNGbaldGM9ozV1fHX+T5j039B2dbmOo2s0bwH6zZY0seKedBzv56+/e
LXu+w/TvBMhEXzsRFtRGS1nSURBsI06Mpw51DHWaeeoNylqTayUSlKptl2AE6ZsE
S3Qo124twXLU2ZUQpMtWDNWpd9q1jLwDNAQmyIn6OQ2+KeOsOs4vlya1c5D51Zwz
IcNbBX8Ni1WSpzQWCkwxkxK0KsZ+Q1Je0ypQlG0Lco+G//dSJYEQdSjomBgU0rM6
8OZwQsUbK5k6dpBxWZUriGj8Gql8wrIOHEphBVhS7bdpTkNq4nsaG5Vv6Ie7LHKD
Zx9k9XSA3WkFo9kvmchob7mNF6lutZhF6Xucu7WBX5qKUes7L2u208YNMRT8XoDb
DBV9/5SHzI0dEq1JARaIO4afcjxIS9l9nwUDgT0tZ6uuV9MwzGGvCe6LhkpUtJTx
0jzsN7ZsvBZrkJfCBqqoUAvegwbpkqeMnuiITw2cRoqnKy8SpDCCVswMhVRzGwy8
P1Lj+kR5OyWVrirLSCigEUjFwFZczt2lC2oGcGWW1AXn8a8ViQldGPM0W7Ko8yC5
0iPMHOXNCoJePyl+lpxSNVIjQGJI42d1pbdqop0uHDY/hh2izpuEuWX7pguZ3XJk
YWdLANLFu1S0LtniWQTJu0Jiy6XKh4k93MIf7XvKrgTRj5U6JXyJJpgvXcvzAA/4
8ajTxqWfwJmD2YpExNvX0Yax6EMnFZKD8nqqp2kWk7ZHdBh11VN+zN8OuHx5/TqF
yvnm+aIjS6KcNtuqme9pYCsiCVsMHkRdu7oTjT28DhNYklX3pKbq2wJE0TMndI1l
jG7uoCqQ2H5Fl1aCrmjk0n5ErLe+BHhzeDmLzkNf+iLrArUfOdiOjlmgLuy0YrGM
CKWgzh8bH6Gn19tEsHin+Z8W0vSPfWwyXT4Fzznp8w9NfxN/yz0kdoygMbQJ6F5u
/dRRLbMfXWnmWfUE2RiCcO/t+yU9MLFvETtVrPcDPY1To7xeEUCj0GEI23fvlujI
JiRAMm1nn6SpDCiujXCCro4VeyoYFhVPVzwguG/ZaHTzVfE826q9i39trizsDuxP
YrvdgRjbD2qUbqjbXn+0+mlsCj3LcovNyeUiNCdukmXX73f9T+zQeZV+uaZMf4P5
Xe/IUlECkUpZvo4uybkQRNb2CFY20ykTiLEo3daspbKP7wHmfP2wIa+h2Llv1tXD
MQbMJdHG7bqk9nEUCUG2iR0XZCokFDkefY5bD33FTFsQidayCSIdSNcdFPbDkDOi
NBi1RD6l1ZxlYWKMMO4LRn39imA1nnJZmisHUXx0VSt//pj7r0HcOeclnY9/EANu
K1GedH6bcJhV21EApKLXjeQkoIT6kViGAC0XtkzoIHzW5sVOexg0n4PKyvmGZDQU
IQ2MZthqGtBw4NoxiveqvOArrnA+zZsWEkuEa3YyPOl/oocIVfcM6Wga3Elx1zvd
hWrb3bNb8vSyf5cUTrih0i1J7PURSNHGGL0mNts672B/5QLYd4PTySlgu1G+L4RZ
bbNXvslAkMCDJ6x4Nu4EersSpO5gdShuoCMsxDR1X386eDOJ+nOEP1pFV64g10dq
KLVpqvmlleR/Dd6oEWyA+E8kvnhLwyFhuWRixku0mz6SK4QdUid3Vl4YGzLoF38y
pklHpKrxsuxRB60lAfgCJNecJF6Y6il58+YvvALDeb57J5pmswW21WQnXWzLk87R
7xtDZ1G/xdgsg+X/VX5L/+xxO/TwUhaDkMtMn9Ubv6HU4JD/kBK0tl/VZV5KdyUN
nUrnbMxFkaZ2l9OQFdpgooJ16z/AJiTOSzg9srDPlanRiGLE1KZVyKp+rpp7nVFC
CnNTSHUu0owDD5XHiAs+yCBgcKV8jDmNqj3bE3sKQMFf3lvvZO0MNQZAjxrtR8hZ
0nttu+Dueu9nvV0S++r+N4So0hdu3yVW0eywwpg/Kj7YzNvGw3jf8GuGZwV8VEq+
YJmoOzhtrmF6EH0YMkyQcQqPmpBAWlCDa2op1kbYHdUnDSTD2s1VAVsq4GKegExr
H+/WvoTBXPzleBQlV0cK/a720TOAcLMRwVXzcb2o2tpMuYM6QPkG9EKli+S50GXI
7rDGEzxp4tE1A8WQpQLdS0Yej2zxCeOaLozM54HqfeWB63RBMhrO7Q3+gJmeACvd
kl7SWY/ERrNcL7y243u7q0MezHBfBL8RmHuWPo7znxfWmKK0mdvhLmKwJSLWbe3f
lpWqVQq+uEfhQXQ7PEYjFv/bCDXApyDKIUioT3f8Bsx3snHH3GRqbfoPVYrVFksY
f9GkE/eveV2R1nUlvDRbENYYsCrL4W9OxiSCOpDWfThDC9idX22gwLZm4a9KI7MZ
hAVnZD9UgS53MuDAzFIgQa/7+k2Lz5LELgCYDaZ8pRyYjkMlAio9/i2+Jg5ssuBb
2PT/5XdcDxN/kHp0xdXCvloWI9ow65kbJewkoChqkSeCjtMLHmROYk+Bc3MQqAEm
uo7Doabguxe1AlpoHAM1gGxj+j1Eh1iaolkXDFyFC7/DmT0hdMS9mmqylutd1eki
TOJ3bzdX3ljd7aJdqELVkl4sPGMSCJs6uaPQ6QMWsezEFqN7wIvcdDh3W51fKq3I
FoIr6QPs5uV+dpliinYriNBXNGywVZKZDuMaMpSmGlusq/flBV3XPOwdqOA5Nho1
N6lcstY+fO+D1rSZfte7tvy4dQxxq8XIlgjJRbXpdlf6lYTL3T8nWAdHduN8RlSg
cuNOkSqwYIJlcw8vpMPgAmXtqNQe9G/3FeEf5sNqQm601Ll5E4chY2OXcjMGFFf3
t4fs4rPO5DUyrgcR/fJy5y51xPEQns3Oj5EUhbEui1PLBrOEjw+6R428zByIWUim
E/5XxFltui1w2Ya6Hl6MB8tGmD18IPetg8f+e5d2HeNY3j3ds2CA7cPe8AcIztPU
D1N/ba42JW0T+KKh0xhIyZ84DTZv8gg/WF/Fx1Qh5bwb8GZ4vD9kVDW+OYNPztkp
YfwPrFLxeqNr4qbF9dfgTsXy0rJ9A2vayUkjCUAg/WICaHa/wFKG7adWCrz7U4yQ
viryMmsAOQZABro/dB0uL/FA+qUw1HIekCZup0DM+TPWHcQz7ZOOMnUUrQkIJjE0
9+4lehEb6yDMRHGl2wjq+8WpMTCtXmluS9MvOAgg028GE8i2nMKd7uOxqzQNqkRX
eCjG5PFOullBOf/ESTZvJYCUKYv+DbQq7hHmwMmeaTvaLdZ9uikBOaTCiYUFu68e
A38mIZTBouYvsqho7WMflqKyDnwDe9MPbebk89ke4r9EyD5dM10aTdxXbgamL6O4
dUB5nsGaU8+WtFgH11aUsRdeGhQv9nxertX1xIXmFuo4P4/QWPhpajUUrCLByGqK
uVWwQPVy8zN3rKi5hGUnd7VoAYyJ6D6qqabsYgFFxLgdkc0w/LkA6FC5StCWhkfD
XEjizamQyXqENfjfKTOGwbZ2Q4Q+L4hlnuzbYaRfXY4CX4PaDB8FaeI/tJRp223l
FPzNqtzC9h9jVxrL+aoG5kk2zK9HVTZv9JvdgtoZa07cj141XToUmj98/i8nHUnR
4Ph36WZC7u9tADt8POvJlAE0M/L8rdNsNdMzqUsrF1r+w/t+vQE+QOKn3FUnNClF
pvX9AR8ms5GjM3AQX44cU6NYZ/FRNEF4+sArYawcD2aVv6PSM19PgMADcU4XsuvY
VOGMkD4Wboj+Mq4xTdUgwK81nicpsvmd2ycd6PtsgnmQsDWW9RFS19HLIqx1Wo1k
EZ1D4eDu8WD7UJWONlS+vRpg0WG/irkXDq3JbGz/7aqkONBQW5Mp0gazIuNSFQnw
u1mevFnJf0AudULcXcNnr2pnvqe92xCwdl+5zSj8EOv3Qh0txmIjfJJh2AT+kNoI
MvtKDQAt7fbQhkf7aQhGt9wTky4ThkKEiKtUM45dZhJ82cCid4chDv0kMONB/Kz5
EQexIi7Js5TrVWYvBNp8hD8UP/eQx565tndze7v34AJcrTTW8dN63juBumfa2mRE
mGqkgFkMS9Zx2UrHERcSHXMa+duafJ1vZqC7nMtVvBj+x0EEjvXrZKCJYoersgyZ
fvZRuLvPWVp7mkFMRSLymv4W8bdOxuyR2oGH0DfuLuNPN38mTGx5G+m+AsjDvCSU
Iue/0fVb6N6PGO9zu2EWx3AjGg7bXuhNj5dISSCStFwa/NjgRgmETI+qZpxRZrgX
PqP4Qz8uRZWteum6Ee241L2kgDSFSNsJ0pTOGoJ+nPvCLjUWVks93EPyxdsuCfUI
n24gSu4CdRbbJNFPsiinNfIk+UCdqMZWXMnHVU+NZS9f4sq/cN9OG1GqMbW8sSJZ
QywqZXDAGj8GKDeC6vStv5rqePV3BpWySuPQbu8iQTzyzoFqFEDN982VLvjDo71l
Xy1WvFH9cVRwx0DKmLtoJnvTxc/BcxCSLCS2WgLNDpUwsTkRHX0/S1PTqqnARyh7
zTca09i9keMByW4fNEcU6fCEMeWYpuApTnFVXCRAeb6srQQ8SemnizQBVbvghaDI
bKT5ICBuXxcJm/ROE5ga6JB8R8zqu/8B5tkY9Eegv9kgmlzgI/tNLzO08/osoXv4
UatBa9QQENzyr7FqU8ZVgrAL/IzgO6dZ83LXmSF9kAn+Eqn35wjGjoJjSYUKwnF/
iqxqvKVROFXjsPp8NRC17aP8pVl3rpVEKtrE22Fs3zornpl+2D1o0P+6HDqXqXcY
ik3RB9ac+Yl8aClm7HdoB0dlPxLuPkG/lwrdWNyJ1oLP5Kx28+OCRXbq3ec7qf50
WtA144qJLErawZTCm7qnsYkEsqBYzPUjMnekDU14kzhfC17e0QbAvXVQ8M12xw7X
i5z74FB6+DUntpzqgK/UbUoA0IPXgNb+EbF6Be+7RVmTBvSXLyrmNZeZlLAaqQUB
Cpx2mkipZgVMQBwUiNL9stj+W8cdfGsXZ4DtVkDPi3Shwvq6bt7QE2VLJQ9K4a1R
k3K+2vatjTEgveZNgkGWzEItalShLLFTVlXDpZGFFS/1fjMfv9xoOjRh1f5DZ5qT
glDg5ydbhzPbFBBJGZEePTfB5r99CiPRVAF8vldod5TowKNvo+1KB4b5g9ee/ZHt
xMg4TUvWlz1T6RzUifEyKR1QuwlF8yWGnyJe9xpSZazYNf54olyoTmVeYSfzCPvN
9OmaX3uZuhsKhFwSx2tYWXXc4SGgceP24NRhJvtoJcZjDP35zZcAokqDwnMPgWaE
24CQX5I++CSjU5K05oxQ12tHTcQH/bIV+pv88Y1wh4GjVNQozBXxrdFG8RLqEZ3B
7SNXmY4xtnbe8/ptq6XwoqfMNT0uJxfnEfLYUSssjyLlcakhDxf8DDjiBvfWhtA8
ExjtxSsidSEk92Z5s2ll8IE2CiQ8bYlfMt+iY8rNnd2VjoLv9nsSPbM9GEKBNg2P
iCTfTzRqy53nzMjuffcywmboUwlWMplR+03oapX6KkU2HW9WFGep5FauVU/ugzW2
/dwsM/MVt6DN24I4Ojfz4blW4DWoHji28v5+WfAU1WoWB35g6UatVNZVbkMWC/3l
QmNkvTOVSziQ0Khf+yZayJ71pyEz4ODgsChm+70bDHlolnekpU8v9Os6FFw9c0Kj
xFmREXTohM3xF48gT/eV5UISCyih8FqL9gq/Pdy3sfpEou6qEbWDXXRz7runAVaB
A+Z284ZH/CvordoDIPuuEkJlaqFsaM07oT72zEbylwQAdxX49rslFOciP8MIhDdZ
XEbB/bjvYEim+63NX6VONHcpTnHioJdcREmPkL79Kk/pUwzobBamnFL5TDda6mIH
7iAj0AMd5ZtYL4RviKemfbTCkePMzkJYD1gbfldF9V2fW3uFctTyOFabPI1akguG
AwMKi7JI28kCBgAuy3DoTXj/BbUhL54/uwztlbNz1mSgCNeQ6vq4hjiCezE4g7Fe
5YhRSVA8BhBNGiTOiV3xk0fUIbDBzd9bIAph+YPhlHrTchOBLB/ykX2ESZQ1SSgC
/42TkZKGIcTzL2UGIYEPN0mfQGFrdWEK3HVttOAW1HnpNiE9Vc7z9iomLx35buMx
i49Ki8kz44ZwkhDcBKd5ko9nKBlcnBkNX0r3aeqDgv20lyqOo0qy9Qx3MG/EhBkW
ODh/k9DnitgaAz2iIEw6dYQmyEPvmuc9g7bVOCRwRJYJJpk488F9RgnXcfDO39lJ
lW26eFf1z3lFhTOknHwIYMa55WxcQIOLH+SsWiDt1va/nkQI8QF/1MLOorPSVIAC
SFFnsXrUxQiMe3FxP4PZ7D/5FtJ+vhGJQ4ERZ8RD8Mhf+u9DE2LUiP49eNT4qwai
Tg3eiZVTn94kYWblS3Uy6zDx5xkHHNfhKzvwIpcPI9uJX5TbikCST+5BoJOUw+Wy
LUbH3OotEtWpw+FEa2YGC6RapS1MtPybf/a+GH1oKEdCEzLZulU/v6elyWXlOP+6
F5kumIpYaXRYt94tPEF/R2Q95jB5xWmwqz2ZckZVLU3M8zB7nc9cBSC4AVm4fG9T
NkC9ECHT2lcuWPA4g8ASxc3jm8k7luoHugqK4MmA3otZJ7/1fipXfRsrd55yD/fh
2lam6qUIZCSo89yv5b+QJTFiceU5JeM9ztvi8NDsTBN3euxfSXweZg7W8BPiWMfw
b98/zKbR7k/hl4oYPK6EN81X859uZ2YH6grVj7gDvpgs+UW7m+Yf9tCOI5PjbcXc
ZL0yeP+HYn/fsiLY4+CPjEnPR5IJJGfziJF2kT6nFERvcCShPzUo0bXs8IcjgBv+
9WYkb+1JkZfkJDPt5HAE84OwJa4cmLJ7I98HSjhsCcJNsHURxOu8aLO3oSu5be2C
4SryS3b4K9cSDeqUxpuoPkGfcMXuBwe4jTPzgfRU3SCSynz1JBGliYxKr0tMps7U
Osn72sSt7Xh89aT+WtG4bhDBvFm2RiPE47fKfFXo8CLK6W2HHVSc2zNAYEr/Dhdu
0TUYEcYsBDSREEttgmpeED4viS+GL8t9TwdW42ncXxKbQciuJ2Zu7mQdWXwLkYVw
TQP9RzFa1UpwuULbDNG15mh645bb9ssejeeKE1SciMNmRuWzID7lR9fa8PRZf8EA
T7hHxxEFeR9Ex9ou2VKHS2DZGGw0NeZ/yJTTmGHj7UW3ntsNAiJAXW0x5CBLrxTU
ypJbxJ0BQ3hFJb/relpQelPz6bE4EKZHhLsedPF9ei70CglpJQT6Pj/JOhaZyrh9
0/tlrqIdROWJ990QOMh2TCixU7LF7JVN6xmuqPP8ZF4id6jLyUFjGkJ6USIH6Cu/
KndV2wEp6GTd9nNnJyWl2FEV2swYtZK4W2m6gdU6EJkVxSr1HysICW8N7w7A8uu/
k3P04xvBmNWr5eRSSuFJaD9XmFh8O+UFRiE+XqcIer1aA90G0M7nhIdafeXHAEWm
+qr7A0KuDzATbEhOXYnM2YqAB3Z/O2WMC+149ZVKaYW7OIwSM/i5KFJV3SXR4a7X
5dDdGcHN0uihrOq0YSUeDQSl+9+tyb6zolYcAlx/nY81MwID8I7MyaTGVVDFfEGO
HYXsh0rk0bURyM6Vp9eu4r2IRgGjI8cy9iY8Qf5xUedZSZF1w6dAWowmi6Vma8em
RUnPqSrwnFe1fbDS+G3K7+Ej/AQmT4JkPJqTCua5rxKrxNKGsR6sJuIGeY061k5C
leycyRYX6gtVPhrL/gscLJ7EnNV9e7h0o9p5OzYKM72ADvlFsWWItQnx/MQlCJhc
BXsaiMCVLLfDp6tsBdohiQDnsqLAxDHafR+Hr45tHksdKm66DDDTtkS5y9YbKNI/
hDGzKpt1OlSmxPB7STg/qEi9IYHHdgWtF0Ie3qmtzZi875HJeb5E8qiX3lOsHOPH
a/imgO8FAWyU/b/1IdN63APbjawR6kngxcXA7mX2K1OPJISRrNnwdZVXB3+kj+Pw
340rCUxOGbCP++N0SyxorOA8g2f39+f22PP8bJFM1Hgg6yTY4n99FfhJ1Xvy0q0k
bVWSnhYteT/tY5Ud6QX7i/w1tW5LrPuIJZWlczDRhySspEdR4p+NrQg6q/V8E0kg
gq8j/EHookg8xekW/UYZhC9+MHbyHomu5ZUKB3osXt233AJWYUtyvreqZmM372L3
ihjpiPB9L1aYOpyAoMgYuY5DD6AygmSUDtghWO3CdIQAPUuxa/acaHjE1ARWuAat
wUxopFcS/slXUYDT0KlFH6XCHXoUvZJppKjscOViRFnwkxQoPCHxjZbkhyIL47BP
tRkzfeASaPFY7zU0Ty6qd4Z+edkG6h5BXEO4cocLjO1vtJMzbC+KvJOmZAe5rn4e
gdKDopCjTe3jThl2MsuYr6OORiCi6kZjWNYzjIjMeWsdm3B0/8fbSZNrJc/MNewb
lZFPn462iFOoNDOaaRwq8x288jhVOBPMPUkwG5xLHjgTimUvZEKaKL9RKkPtJ/ys
agfWCeA5VdLGV5xhyM8axtoBZDq4B2h1Hi1ZpDjfUOwkbsYbHH5bpVmMP4dsE7lL
jMosYNMlNiAljGtIPGWOyEoDlcZExBTVGS1ZDsD8efBLkX5UtVpTboIErRpdFr7D
ESIbHu53xP5w4QaIM0zslFGy9kQ9zl654WAdjgMsFarxE8DJiWNbXS89cdP1Raxs
kLY6bdOhLBKcLOkI+YzHwXEuJwDBsdAF4svgP3ZsyCyJanUxk6S/mZOHSjEKj4yW
KKa76va2+3b8RC8ZDShT2e+ZC/thf4I5/N0EsGQni2pKrVoFs7ESwjLWRaB8b0Fy
GEOgyuu5Frn/ngPdA3BaNJTSIWL52CXx/Emt7GIKTBFsbnWQ9qZ5/BkdDNcrO2a/
tbXKBXyEiD7+yJahvJ+MKlPrxh7IncoLQy0FFj0tMOL7m7q0ZpAfzY7jgXaz2c8w
DPeB+E47+1YVn+4r2KLRZgqZSXi2cwaUi72P6sIHOONvjmRXyGwQwtB0a+cni0UJ
CumcqEJ5Ew3S3FDGWSXua2bcs5zr+vOmGwBEtw0WKJ90sVKKKd5UJbVnzAIz+cY5
GZi+6GmVye30gpaHWOyU+PIh9ceWTtzgRpHp1rOPm8PuL0jn7CzADwlnw8xfODJQ
y8T3jUvquHKOFJn6yh3iXDx5bUWVxt1JbW9zDBDDuqZcGYfGC2Ask7Uk2/hvQWa7
MsR6f6ycyNMIpHg8GXi+Nj4NuzAEXwLIsjUESGKPrFJW9zy9X2IcWnhAUI30SKoy
4P5E4OYgvgK7lT1sM+0w3Rkn2eq3SR1gzxi5L859dpGpWxjaDjF4nYoZte4JyZC1
1ZbFKHXurVKbebqq9EG0cX8gTtf+ytE0KU84x2skIRipTj+5v2p477EhwYyxC/su
0zsuFTZbqiAAcnphZCvjGTEXmoPQYgVOqgj5IaijA9VjBVEfQS+WVeEXP+SBEqv1
kgHAuTRUAC3KnwlOXChbK7KkCgpqIQ5uZBpSjgfDFdHTxG7jyH5vWCjj0Lcw7NzY
HDVLS7V5n2DZwwm7jbz/aBGAtXfVXcwP5luSrBDOCMXjUVDoUsCqo2f7hgTxj383
HxQ+gBSkYhhW3ruwRWLBNNAtVS5JLU97wPnfQEu+F2FSF/2mTutr8kd4riVf489a
M4RaBVcE5it34V36QmN3UxlwA5ssmXLSKR3DEHtiqamE1UJd0UNEN06geEFWfnMg
+0h+cTmPz2XOPWVzJlKFTCsYhMBmieyAq87+CPlY//ukzBHqcxXx5aOoCURTBVGu
ocxpWWH0/eCPPfzK3+ntPVZVO6njUdDmdTO/v3SFRoAn3fde6+A/d7QOVFf34vQh
j7pAiyKQ5+OBKRCN5QoF5Te8Klk2+EjRlXrj7dw5YcXBBt/21VDed60JFROrdqyH
IZ0u5DnX32uBtMhdHSC5Co3QzB5Wc8zuEeDaSaWeGDi59NkZrVHzcHcyW7m9SEAh
0ng/wYy7zN7W9CtYDgfA5TDsH84ib24MrDm4NpWqsQko7nAw1R2bwZUxV2n+n2ET
0hdSyTGzlOvfCu62nw3RXkXpQRTO6cV4uJtNuACBk15F53TN7cBGHmgQujVRLvGO
GVvhaQAk5g4HVGvoKP9mI4Weo2+a67DTJ8Vys/3tZ0p8yDMlCUwVQhqRZ4bFFEHO
Ubi6Ys0tTbtVrscuPMxNAV2XUOHjmpNrMXgM1a7EOCvPBDoaqBFLf0WzuKVpSzyy
yEw5Ek22uF8g5sCteGtAUWe9WP8yH7V3Qs+g/eJ3lDxyLjOo7hwGrXXEqNMVt3jC
aMZMw575a9wp4Dd+vH3SWOaaXRYNj/WwFS3bPa9XnnHVzYbKbBqDyfLM9fW5XnnW
/Q9fzyA6UCA2Icq2+ZjxPVDqvuFA1wG/hGQhODMkodAJaN9YvM0xQ4sSboPoDd2B
5UGYHlyTRGa0xEzETM39ZX9nGZH1W+lwO+p8CEyTNY2X3w/9WYilzc+RXraCGP58
c0XdLetSgBbVkjjWgowviJDC6s7MuI+h8fyH8GqtErw8RDdZ9ZGAU800e4w3Juo+
g/23RtIQ/Pmy31s0ONMFYcZqeNGtT8QAfN6SB6NJEibGPE9dRPq6iyXyyJRK0c+O
FB+wg7B9Az6Re+aQa+CHU4iwAwr7jBoPSESSU12d/oE8aLu+fDl6FiG8CwadZDzr
2FWy0QZErRHMa/fmcPgUpYZRADjUUm5WCnd3b5nV06Myizs9iPwjCiUtV437Tl62
u98jdxgX1NsxQXAdGSvIWmihnlQIH0KOUM2L5hUdW+DvPQCEIk6GspJM/qNoDHja
9vnxUqtwvwtBiWn/8olENjGikIlwVRoLWDlZQ0r3Ov7ZZY4VmRlURJb2mpZ6wJNd
7m8BseAlfBUKykqfxNY4y1qA7iOWsukWwcH7fzdGhNyHZG9HFQ1iYoQz/+yNbXfI
oFOrmpLR5IhGYkeQsxLd3f5Lm4JMVeWwN+tjAy+YE3sbuBn8X0jQ3+Utg7rMh3N3
cRVKeyd9gZKczUtfg9yIK8HAbZVVCBxSYjKfob8PuUI2bRD6/LRNpDzLtdIIH2SX
kN9d/eeZAfJ9s77Ha2adE/2KdQdNZ5HSNTLzV5ZOsXSin3bCfX4epS+jg+NpCAz+
e/xL0tb3LgZVbBHCcCA+PTlUoVcAgWuWdk0oGhlivnrzENWKPTRb4OkRbfkdRNe0
IbIk4nI1/Ko24GPlmpNqDBWkHfyUytQoFPZpLbLyfRm9RAur0G/QN16fMMzYElML
+YJtn35pNnNk/tdnOifL8WP2Blk42HQeFM4N5v7/HNljwvX3CDk+CAmiEO5f/e+R
Dr7ScgHYeHghf2FvZFP9Q4fVM8/SPns7IKGQ0zBBDdjERUs5VwD/XXZwtPufku3c
pM6AHYLlm+B8OYMQJL6X3wDInYGOMqkNgs2f1nZZI1b1NKfYHVgjypt4ZOjgffBQ
ZJVAv7knCfKuW4dgpMTb/YQpfb7n0JOqQ+Gu7JDQ3I7cJXG47X1yYr4lZkpLKsO5
i31xQ7fp548Zwh8HaXf+T2Wj5TI6SSG0KsEFXGbSpEuj9x2o7QbcXTM3lGmG9Tch
wvLs70xMpw6Asy641TMru4rBOcmZXkDk2Xe3hdwudngfNjBRj0tYJt5uAm3CO0p2
rcTrk1fkdSg+PC7gk0t11I/AcpSCm/PH6fBrSGHSAIm84qqXgZJ/J5wfKvqpC9Gk
sv8mUX5fgBUK00Ejw+bHBJtzIOj/u6B3e4ovFsml554PBNU8K5b/1fJIN9uY4bjB
VeCa3KejsD8/Ny3U+2mGvZ1rlW0GbcpqO1mLtdXUbq50ZhjYflHK46oSY+W75EKG
Q6cIMMaAeCvJRFYv/6Zc0qf1rbl6pCrWXiyuZSGpXXZigpyuTIr2st+yIROanW2E
vUSEsgNdjxtXLSuJKUGwzY4vgwfSpRDqNeaGCNPhpHnv6F6Bn4qFPA0hCnlGW+l8
sIVXaCDHp3Xh1LR7jM1cs1tnvCSm7d4SgvJGiWnfyW39VEQbHQFu+ofJkG7Cdzn+
Xs3uXIJX1iKPeFrIRwOdsGS61wntY9d7EWaDXC+Jg1Y1v9itSdEw0FD7kNSYCQxf
sNgGgnhcS7zSL2CVL08+i4el45qVI3QGdsdVOsHTMdsxNBefeugo2Je+BK8tv3+T
WZ4LA7GbIK8RA2ckmSd9yzvfeE/CZEon72UA0cksIgu24tKktngu2Um759vzB97R
Pd3tBkOYgi4UVhlSMb6n3aVHruQ+kYk22T/xHhZ5BBVzcFCfhMEKcDQAb71Vbo11
qdwijkYV8LeA4fYA3PO7QX/7xv7g5VTVkXMcdHp01/9ebWokXjxyU1JZV/E79sEu
W+SyeLb4UbDeJoyteHjUDidwyD1joE75nBMMMqGcDUHLG9z44y/w3gA4ddwp5+GO
gLTmBvk5G6nQogS3F1kFYYqBfx1UfC/jIE+b5PhEECltZPaCO9gcbvaaaK6C7X02
5cAf2YlB8/rATcv6s+ciNvIwoxMyL2WJS/uGfo6ML7wknYjQME5/zrYBkoGriAnC
uolkEHHel1pASV+laWU8/4QiL5WoU08ate+otSqziscW+wfzh3qkE9eFrxY1RZtE
733UeHTKF9MnxmKAvdRAcC2fctKikzWt7wgY5xscCZY/ELmY252y7tv6ny+PL/Ta
GJSorYMLqB2dSHJRW7r8nkFmhjdvmb9eBn1gxp63eQMVn+88p0woNIPfGnz4Huer
uhwwN/9OBK+QFXmebwpBhzje+B+O0fUeKIuEXglBW7ilu0H3OTI+wRrvBZ919Y4V
gc7r4ZMKGmiAjiVB5FhKbSD8MfCam1u9FWB/uwQujeHtUlGYynkmaOg0GzJUnbRF
RH3lgUE0PwZ7wod55CUMOnNk1GSuPzNmXJIbCzPndAD7eHlM8WKxBemfyQKhsXfI
e171XJFeYT86sELOeLxQIvJvvmU9v631BfgvzxHxg7gCSEjOK+XXa09NuiDd/lMI
D6kQHW6QxoLwH0koeUj5FS2d/vO0/59TXy6tUL/Z0iIZSTFmR201LAWClaxv1ITO
gaTD5opJ8zti2GlMNhJdAf3AohoDHQJ0pmfJRM4au93vh9ONGNlhD43gIDPwmAmA
a+cfsIZ5e1qH7ZCvyW1EbkQeS0ViLfQy8JARTMlN7sbj39+teiKyz/9Wt7dR8cvU
DpKYdmxZWHfQnA+G7xD58vlVHR5rn7zGVS5mHtwklqAhmHmALAalCVYk8R9w0ZoX
rVlmPZVePtkyT2ks7hA5G01HwlTJB4Jej74XSIxE5rIoVILTRHLr98gPqL/auTgR
yRAsEAV7EE14Rl9RSXbfzEMw3q+vXs13HSAXfGmjBDrgGvSgpt6DfLzXHXHHF8Im
4Y/EYfN0Y/Pjmb1sdxaO0U7v6LSvro9Gx7EElfhzBdFd1tXLycfXlekLTEjQHvwj
qT1CWJTr+bpkrl4eMhuaLAsXnakhiQedvmUcRRtJVKEF/ZMV44N25fgkd0UBrg3R
lLoAXBxMaQKBr5G/iSIjSv4IOc4Mx2xjsbfoDJBiBWFt+AWEO+HhYwoo9g6oz07z
XMkLINFSK+UHjV6rHP6aGSBz6YcoWyNXf1WImpezQBipLnoCzK0dVtvGTtqK7DQQ
uySpy1unITtHn+MfFn0E/P9L/v+tgbsOy8iSTYc0gcqfyXzdikzeB9OCfraIKFKC
jn0g868bTQ11Zxki7yf6QL+2UWcrxGKSZV0tYj9tXwsz0Fvsq4n0HSrpQ1bdWfpy
Hf6piiaPeKPW8OdUjrkYICFNOqsDmIojS4ora9YOXnEO+d8OAf99iX51WKFWYd6h
lY36H3DEO6nP8qFBzuEzGu2HS/JI9NfEv4zP51PFHRkmQykG4cyVeU+pm/TR0Mo3
sZJe3UjVjUW+MUrCJTOVFkhNFk7L08KHfeUx+t8ox/2EyQobmB92V1tfMEUOPSVh
s/Oe4MtLKGbYa8LqdqCr5IhM0770pM+0xWm0CGXyWkSepQba4JGm1Ol5F6JieZ3E
4MdivFO1wEPtSK8wQn3yI6U2T4Iujo2aK2SXgDdwJboB9LAaFA8t9Po66qwtl17O
x0RZFqc5VviEZxP0sazorrqfk68qpn46dbpFIxoPIOiG03F9BGhKJR0bzK6CUex9
nBc7jalEbHOdD/JbDyDQlVB2ohFoFzcpDFKt3wlf3+ZbIeUoDUALkfFBu73gyHA9
WrxqViC3strehbkh3YStpg5m1yqgbijQrWTj7dtGW9dUTl+pPw2zdfHVvPVlIpaX
F2BuYtOleoBjnOyUBz4Ozp0HSdpMaUUtxL6p3/RAyjF5TQuqHCOWN1a2CDB/y0Cr
OsYONJRVPVZo/7ehTUUcHn9A2c+V+kbGqeCioGLb62I/W6++vtC8tlSyzv0VfnKl
kROAvYQ7TDLEJz9uW9hYqZt3w4lXGksJtUoqW5YZ74gkyOppJ6PlCF2jETApO8mK
91m8Z3vw1nZbIvKS6QsuF5vAeHQo6ar2c+vtvJ9jW+sR9io84bZeOVdJj7bZaAds
bh3Htg50y7EUM+qTzZy29oSEDJPA5VjD/nG9wVPO3vzdIBQRv2g9+bXCBFR3ZOw4
2Njm6Jm6spdilmI9+hGpbcI+trfoAQyCrivZyFqm8Eh7bL7jwJY1NfWZu7WmEwXt
KuM791y/2WnAx1kcQGuNyTQpe8gCY/ztMr7Bn8++VyDK3tLTQLsplA/DL29DpXwm
+RTOZGLMdTMliXdgJHW8AO2P/GgfdauTRHu8Rv0Fe4+9cs75KTFRalcHnxW2cJlQ
aojnlAqIGrGFPs7QuQwjc9//lELgqD7Yjk/M2ZfccqJo0LE99Pu3arEcDZaTLn+5
pGRosUf8C5Urxqz988G4rD7J0u9JSEiJzNgCiRG8ikO4qdMghXf1LxwHVPUqkY+k
2xxZ5BxNV053Aset+c1zRwTGIRmS5LobA8kTrNJxGY8KLOBEZafsslDAEf+9dzMG
2eLj4NioMejK2yGGtUocYRO5Sn4wggMl0AeDwEiWeb2T8jNMEliKFy3KTUqZwdQL
eFcyf5nwW7oNQ9revfM5AEzdia5KgqyPatkiesY2COEOz9cLL1rSKHsNNXoDmZZl
VMUU0lg7ZfpA+K/wIwyq8+SYEIndZmeeFN5lS6EKVLrzRfehXbr0IzNOIkM6TnzN
G4iKf07+57Mjdnuzvw7GgTgbXqQZzh8zxjC9STRI1y+Ek1LlgQgDUZNkZU1T+YKR
5c2CgXAcSieT0h2wNPClpl5SlCZ/sqeeFsJ02IhRzT1rk5BGMucMv2e+EHBqAoiQ
57amAaglsahQ9S/hHZgU+2hXNRjsQfUaW8PIjaT/6ZWmG+4Tl1LIaRDDmNwTSRs1
xk7dwdal4QLxlk6s0fO1h/43TiasJO4Le/nz6uxCTePrCuio1Ma/lEpQ/TIfmDYC
OBQZa+ahmRenPqzNj5cynwoO84ss5EvFfg5i63rCihsIcYUD998qiABF0+feYizX
X+UnY/mR7ZgD520aXYTf056xiLCKJdtAkAnsz2TyLxnF/5wTy8KpWv8Uk7ltRpKv
lBGGd6g43vMDLlA0X1cOTVwKnKwnHUCDDtGyMon9QpZy6tFhwGeBv9GIEcvYADfy
r2b7oyivDVU5lLMc/CTXufQ07LXornL2gRb9y6nhkh9heUdElqT1Vg/OWKlvG4sB
96ISjVHYhbnhKdsxkAPnLMHccRnN2qalIE51ae023WBBIK2iU9audC8s+LZbTGEa
M6ILWE/dijieJJvAAbY+vRIA2uOAQuwI9PrcsnDZDS41bgX71um2BK189r0SZyHU
QBxCJrHkyFPFgW6neeXrM6Ye4M++A52u0CVOaVBJXOe5hDAsLMBIbZNOG+8puihp
BpOl2Xl/wP7LmwZF+nIvw97Rb2IF8Tckxg5gEFHCDMUmEiEAuKTyFA/auGkJ92HX
j6QHFuZRqCF8Bo2rnF3RpWTBHGeyM1m/De3kVqUJl59pA6d0+xKWofimYMlrQWMa
1EUvk38o+C5pklf+hJk4nJyZa2PXl5X0mIgQjtnopX7yXpxAVc3+R5s5GLpX99r+
9A/37UkbcunvBl610fL/iKldPINS12sAziCSKU/AClkii5y4Aab908JLxg4+3rAu
IGVxS0MHKOPY5ZHfmEAmDrNQOofzZz5i5ZYfS8/C5COPcL3e9CJRWoA0IBZRf6EP
jxn9VW7BP1FHXw6ZmkFkPA3ojBKMDJ1ArKkc918JovJAf7O9MCVhQouWdSm/3LXM
eidJU8O8WDe+VCkHYUMH/yuHOGfbws1FJQzGN3zzJxxR1OJFdMKAZ9dyUrtxWhJW
TjXRGE0UDfavVpgmBsQgJ59z18yo4OhanI9IWFIyfH7XKFX9ohQ5EIbLjNodZIkN
/5Id00YJCoX91YOlZk7wncPxBbFYRgOMOAJ13+Nywzroa7CqxsJdMFtvxD8yy0Ga
bdaxIRxBy8VDo+DsjfmmZwxCOnA095/LlKJqhG9C3D7UUVe0TXO1I/3DiBoKZuCZ
8GnW4pZARoQkhfmjJAbYetkPqwt3PoMDlUMYF9sANhi011jWKjjU4aRqNUW4FLH3
NIhK3vFDz1db0sdykwMrK9FZ2pJxLVAY/W4yAGCPAVKxGirxlc9ZY68uMrqwELNG
QtMZdspgxa2HpY6YOL8XfQ/rWl6Arij2BLqkmTnZ/ZbhtY3a6lJrmQbkmyn0rVOQ
gbwhk3giwMCGjGSGHExgInwN6QN3je0WeUatQDwTXaIIBQwSi/YEVY9ucuAiTSH4
vbxAJwWLCVLQ7+jnFT6TPY8x/b/guKJFVBqBdYFF+Huqz7xI1O+c0f1cAnsKq7xX
LTUlBijZ/VpOkokeivuDn+cUoJzd6pO123jEOeV48z5BpnyCT86GFqCuMdaisD7O
Q7DNYPScMYLHeE2ud9fPW1vwTZ7OcXmuJRhcmSCLoEZGXVPf+KmRmNdr1ST/ya1c
CRap06DwNxFvBbsJ/9Hq/4zHJTyjNsZWtpsythRMxV0K4WLQTYy1GcLTHCKCYVT8
MIvpXsjQvOvFwZEnLBsKCzSlDJmetApASBpg9Qovg6M/v99CpLyvJM/Y955PfRa8
lkUFOsKFnaDv2b4On/FAKy+vI3Er1GfyzDSFLG0YXPqMKaTx1fbc4M1tkTnToJAW
LPs876RCM/geWvEvMcpJN0tVwYkSSgX2CAtGPkbJm3weFRx8N6+OfoPaw3nlV8pY
OojhstdH9J+PDObHjOY5LVdeKOjaPta/n6sDKlyvprUO+UVhPts6LW8eV45mFdkt
4yt/WKRkG+ZONLJigRsGId3TRfPPejgyzZ+C/0R2XmPVKRB73gpkCXln0t/4vbSU
iOdzaxW6hgHcDlCVMux2lgs081kHspdp6/nCsAnPd+AD4wRgJ0ErhIXj3WHH5QQ1
yg9C8Stm5hQ70BFP0o6vonhA5VtSLc6bvAqb1NOdsGbs8CO8lyq96+++n39LxOBj
H02U7dCIsg4dwOLYxLV+VrTknG+QC639nZnoqPU8BaEwVJOeG6jAWOdsZpc659Qq
CvgxJ0Bnc8vJ3rtDH+y6GCW4yYSR1ohpeSgkDKqgH2ALweFwK+Iikm+nItmjBr3y
3oe9pWk29ri8O0dVyCjEBSNfg0reCb1HRJ8QI20YVOSYvyvIG/UHiaEWU2geQcjM
XUVsV6IZ7yFgMUY6SV3IRu3hFtcJguwruDvNVIEPvYb6YEE2Y4hV+/flgrNCw/3e
g2iGeW2bNaug3a4AO93fE6h5m6pfYUV9MYZPhQr45D9yEqb7lLxcdzP+mm1sL6oA
wwt0W6aJIVILjBb7Sn5Q4rh694WpQKlvQJvKSaePLYKdE8yDX/5l38bPYFku5Z1V
sZ0TCWaty6nNPkliAEWTm4JlQgN7MkHwOZBx3muZ4x8nYu3AMsmz6LVpUqlcSvto
iSqczltFEO/qMlXMbyTq/U3JV+7DXaqYD69Fp+cfA0EJTr3SFHnb4iSQAEd+Siig
cGqoBmFoZ+fKXZXCoB6UVe692gund6bzB30Ab8Abbj/t2BlaqyfB51WGMyRavguz
U+QPkxuk+31RRpkL6ukStoivx8mGoSVchqh9fF4W3AsefUXEQODV8VisLNSHryDp
Yf5FrMQprghxQO3tujfC5lg6t+lQ32GYe1J7Pu9/vTkINNnvabs31iHabddB9LLT
d8xjsszyvB01UfUt8yFrfu1awpTfCdhKe/BAEGrh7hxDVpZqKLgNZJ8K/oZhg3kZ
5laf7MqaDXsgeKsOi51rENO5SCeYBQ9i7vNHG4TKBgA1F1lPmRHCVK2KJpgBpu/b
nEjq4cyRUeB3RPeCIlCtTjKP+f0ThSQ5RSwtTPyxM87qy+48/fg6em6gh3Ro8bZ5
0moenhnZ8GdAu7Xd1mXmcx8/hTzMQ2T5mBtxtBS/pxZLD3F+b8qMClmZl+V17Qru
bt1IkawsIVawHTpqDENUBxxIW8HYYXVLxgoulGDBz9yYdvA2bcXbpTr6dhMeUOaM
yiN5MlQeNoBu/U4kfKIDXkv5JRAUTL8EQWp4vAiX+VivcQEpmgzc4S7+4CUNCoAm
stfkQvv0ciSVj3LozdUZwVIc2fm1KEhYgPUmJcEhNZFt82BNLV6fEV4R7S+jGPYO
0m7JPlwpfYU6R0vhUWqwUXd3pmKGpsjyE2vyT/tFsSWPEiesaPClRKQNRAKrdvP4
WydRGFBTdt+SSzMgo2y96IXqQfUjzoidgZVUoajjG2FLPwLvQcqGHU4RzKPAb+BI
fR0Cp5MQjjC00o9gqEbiBTj8VnW01pvpJ/MqqqoDwq6+67LJ+LKp7SaFSeoYar2+
hToPULvliUfo9OmH7bYGJjnXJdem99dmOmZru+4om3JDgriZSiC0LKLgS9zN8oUU
StFPBOuvRqR3rLNZpfStluDxvowJ6Qjsy0vGfAWAWvQK5OTyFjK5vDvrKRkhMH2l
V8seGKRvmCLpij9mLDyM9fB8SOBxH6zCD5/gEuChIq8ZbIByxWbnsOfoZ/iV0mvS
k+byIvsN1IHt/NMHHM0pEQx0wP91+L7q2/OtOkIftDr1QGp8xVWI/46qP8XdMn7C
9FUrhVicAybJyyJNVzyYwRHcaTvI5hc3zZuY04r1HudmeOog5lULD/CM9G2WKnET
l8dC3yHqwvbi3d788pkeGZn6pmmLAIvhMBJi63HzFdSJ1fyqh/VXV+vAWdCyaeP1
J/hP2ypCJ/VVX3mqPaBqNHxdCh+XrKZHPXNUY+4/B07OGCoTVZmQVg3mJhciSrHW
UEbatoF3pf2XgJaoTQaKnZVmq0Mb8zUvBYtB0ng4bKbezvrfn0nQNKF4HaHDIGtW
ny5/geF32PeNWzDxJmLPJXp3bTh2gV8of/0nDE9tRpXy3JJhpUJb8LDLgB6bkWvE
yoRT6unX4M1UMIcwlA1TpP86ymN/7f1h8fxVCfE+dZo3AM5ocFv62WjvhaPQS9XH
D+VCqQ9qx8OtFTyzV+NYHQSo+ymKvDM9eRQZs0g2zht122OuDVUP+MInWMYC/G5Y
uPrJVtj4rgLBuI6SimG8xDqAl6sU7oHddfxZHV020Z/zumSbSeUJ5j81uzwPQxDc
Po7TUWV/BFSz1JcUO9PNt0QrhBJYt8aAJyV3DEatY9c1EeNS+9T/US418xiEnqN4
oV14ng5CXH4CIeQNBFEqFnfU3MrI0jggNPIKkm/i0JZJG+dbcm3MRPRkr2UbdWF1
mBdMsocV1VcoLiBiTYQ27xygYmckXlsNMvXTbsUSgSh7Pbmlpcmv0slOsyCgab6c
L+5gzLhekpoAI+moej0PJBI7Vd/FPI5LET9+pSgwaYROnKFoy84WcSMqNXvHKzYU
nU2KvWdoi4nQc+xFPU6GJbCX53CCgwrChCkU3jA0pjaUaYhzZG1cL4gMlLjBjxv3
TM9h2jT7LdV9V9Np8NSid7K5UND/c8bekNxNm6d51z6HFoflBGVuEEGV51Qe5I7f
GOzudG+TfVl4xbTaBNLJCP/VA9NGIFPQ9LhTuegRsG6UKOml1AsRAFjTAF78vom4
Qd64MhgyGyszodMsmvp6eOFf0lKLwtxQ0koWgR1XcIyRP5TU+NBpDc0/pChSRrVW
h21aMqXHdL+9+ty0u1qHeVBmFnjgt6Aer8XxWJRRsfmXqPuipunOFbtJ5eFNYaWb
FhEw9rbw4u5AreKGOVkrgF3TnkfsBNKTRRtj1FTgE4F14Ma5UH5cpFl34AZwDXb9
BHqDu+PSYYnW0IcsvsJaz1poQslh+InL8jsHVueL/eAl+asGoTwK1OvNDj9/FBRO
fVnIFy+B9kOWTlIZnIpT5YVnQvO4NVQkCKZMOpukCYQ6az12MPAoM1mhB0jSZkrF
eAnkH6lGUI62cTdB2hxQ7G+ig6oRQO5DSGgIFDDX/Ovpt+PwJ79CzfY6uBOyheLG
jdMIgvecC0OS0Wt1I+eP3mYt9ekC8gFjD27sT0lDskrb0ofjkzOwj/fdAvECN8lS
fxldFUxK2BgrUE4NNipmb9HPkhxO/Bex4yPcP1uh1AbXtRdf7MVJ4CQMgP9eMmv+
WdmrS3xhe7+ua5QHsDn4CyIbhcCXOwRz/4pPhTwgTSVz6m7DkDyIsJmRpAc6m9D0
H5qv9phX42Ll41M42V4yOKWP2SGwezHHBI7fDFV7O7n0IkxbGJpCCz0lPgmeAvhr
tlppiZKT2MQdEV1nYhAEn97sUiijNngaN20hGf3aVZw7w/kogPco5frDhlDEdDRz
fUw7dPVRf/QDOU8ZDyuCDBsAJaSFjlrNUxAGdxK11XEOn+hgnOTsFTSDa7a6lM8B
wGm2NAGOTIgXWp6wpnufC+cAw0ZDb6zstCfS/w8ow3hdnYRDcVsfBBP+mzTcDEOJ
68epBMmL4jT8Yz4NsFXMwzFFsadJdJigNGjKnK2ZN2CFRI4wL+JYoTRxP674GEqp
VXuvAe0ptwtsbKALS0Yc7oGRKgZyroUkNzPIkxGrwyonDuaQh9tRosgRGnn7x6x9
OU2xI/Igmms7f4G/guh+VMYUuLBlRqePloc5RroAQHmu2TqtbTsS9NbRcbKFBnMe
8DYQih3DWTy13wT7cD/2/ik9U1i6Gv4L/z0utLMqHQF4QEsIn2x93IhfdOHaHwDH
XUBvKqna59OIz33Md0QeRWGmDrz1wGNXWeRez0GC+hSMI3J28R4hU3ZP30fkhjuC
qwYj/FRbWSimEyLro/85P+Vs3fyrOg8o38zza4IUQWGjQWAjQlI0YYM6BoFeq1wz
h0ZrqKLIRk9BdTWkv1oJ4AVTkZta+aGRBIhnyZotJX0iCNIZ3zrlJ42ND62DqDSS
dtkd4AuDLJeNM0ZoeLYUDndX0f7q6LBvYnX6VYnIPQeidCeKpeiEm1dzoJxkIBfA
mi91jW9/xlt34uCNWNLOLyrQJSul/B4NUgGb7h8vEsfl+JJNCo5I3E3IGtqQLvuy
WCyOWK5TEBUdwBEe0A5TaLID17/0Tsp+XwebJa/u9Hc4cQMAGLq31P7AxlUVsmXk
ZUYO52ztBUUXUCSdmQ7/gyPMGPwJrCk0302Wn7MwJ6EYoq9HFyZDe2XldXL0u0/p
RpFRjuug09Y6hQtI+t7XhhBuhrXt/2hHiX7fY9sl+b2BfqA1ziJzBOwGRQM/k/Uv
7cOdN8wS3V1t81ZI7J77Ij3yu6/i2g9Q6clZNRGvOH5t8HzysqzeA4c3EY8hjd3V
TWSsrHKSkQZeCGITcDcmFip2LIZkJ8AGqCWzlqk5fzKfPw5cnOXwlcNRZWXKlIBO
oFztDIdcQ2sSbr4t070EPe0PHLvi4wyADPAZj0XeIaAyCakUxNqxwZmIptv1zCFi
w7OtLMwL90J+qNyV4Sb8v1VIEJxuJcdece/9KrFxPTQoUlNZ1G7xrRs94uwMMhIN
wgVSHdQ0QOX7FFMLpve/X+UlFE9FhNoar2h79jdI0Zkkbgfowccwd08icAKXQCUM
2DEhZN9cK8LjCD/aY9DQcGAt8xxJQlCyAZWI+G5Dg38GByXyLofx2uGprZKAQNsN
MaIVKs+0CJQ/XX/ieX0MESQ3li3kX/8QJMQxS1FXCk61WmvOiV5bIYKzX+MGFdWB
R5BvRCN98Y9advxbOu0hY2Ww3Wzi55W+W94bkcIJ+D6rEVM+Qncp3yELZ6WMKt7N
iEA0dYCEHh98CoPfpo+PMMUewyWehGyTZ6JA/uKpjH/KGgJmFxe4IoM8621SJaCS
gnJ23Z7ghVv7GPCNckwdyCsiIIwP4is2VMufFHstfNBPaB12zskn3M5ouYqTePmb
wyN1zHNASettNWCJcYCD6ajzLcGYmarG8pyP+u8a9YsB+7BRzm21s7Yd99J+QG80
ntMLCsPOqomMOl4o4hiaHG2LCET5fnlxc+YnE+ndKAoq93fUaMkl71cNjqm4xBx+
23zJ98hQU8b05HvpVQcN0f/15xnAUmGbNE7u7n8w9ItMaGqW4TPmO5AP1DnYJpBw
CkJ3r/iqBA1fIB5Grk+ZkzBe7CwWTsAQz2lWGAfZJARUEmOWaOfYVnnkwvTOkCN8
t4Wi5kVyKrA1V2OgAQ87y8BQMmDRUOjo/Q82SggE3GeIYT9aiJlgqH7NFxkFipEI
ftWLpL/n1b7Rs/5v+FFET4kgMgor0dXuBcFqtbJrsQmtO0XZ4Irb91Va/r3DA0jA
nlOjBz8ngT+ap9x0vDMbkJplbJbh9kLu8CjARZSmsgl9Vk4Xa0tSY8rbPm0QDKcg
J7yKLcDDIPTVeYicYTCG4VFSUuisvEXB5IdwEph6FWXNWz7ukN/FDgLnF08W7guu
120a+ERF8H9gYDZYnnb/jNr2Fji8wP7h13Nk1sqwAB98AQ1gITNWknv2RowXGgFm
TlWKt8/UA9YndSu2iplupiwTqvMVAtXu1sGNAOHN41xufc1M1B9y7Ea+dJgfqJ0L
F9Ry0F31QVuc32BWtax/dFLxoA7KQYFMkWgb50L1mr2NDN6sfmM/RYjLYBYd6Unb
4Gpx17nGbtxwL/4DPHIKX/TdRXj+psaLEskEYPIEqql1cN4RnkcK8EB/07JyalXr
zSf7hbsEBoN4juaLtvLq4aF5A02b72sBDU+VkSL4IOO7nVOff1qZsQ4Rm64+91vR
VM8eHfhVi0Q8MwA1HScrWpOUcYIEghaJ23CATZkFIleDu4bMf8Pg7rzOFANBP+Y1
mozyRNlwmdllBShM8cs9kzUIwZiWLKc5YhNLQ7TecUCOWrocB60DK6TiapsZEnxd
TlPldoJm+ePXIwHSLqE1lJf6Zg9twgeHx4wf5V81HL9BfIggyyEia/UyB4oyOsyl
eR/9hFGvPd9dMsIcQxQepk4d0PahkGJJikY1ilPDkCzmGVdNhNSJgud/yeyM6n1Q
vrM+rR2CKzZu4JFYpG02CqymfIQ4nuLsL8mKkjXbim5BCw/yocTpcHoN9x/oexrH
IfWm3PZxcW5ymHokazGt59CM+koSnBe8NLUt4dxPf8KJiDufoNgBXlxE5P9V3JWI
cYwf1kWvNB+13wyT5/R93iwSg9QS7q8MsGxC6SbE9bbPc271K2b6olGoF1Io0hn3
X9GMo4gYLVqjWLW44MsgOTvVxBrL/88nK7qBg85iD9lOCTH6auogkcnFMG2xh+h7
LlY4qOrFJj/NEyiVMrfAZjeNy5sV+TcY92mB3B0agsvlhWmsR0YFa+CtvzvfTyDP
cewAzTAxNwYXnQw/wrNZd1m5xogAStvmTSOp0LeIbdp+V/4j+4jCekUiKnB8WnRZ
9gydQ0YJQIkKYixa0ZPXKtnZVuGBOwf/WZ0hIeGmrUYbU2gDabIRMHLwmrajcSkt
MYz5aUVWRem78J6PGGNpLl/UOqDASG96bGqG+OsoH5HoH7Buid143hIcf8m94Z8I
6CFNnFBBRDSN4Fx+xtXWDj6y7s2FmZNLoLOj2GC+WAu8Bf7rOZVZuQNTvtJy4B0c
fXHtdO7h0slUKpRLSuxM8e2axFWZzv6HsBI/r2RLU8y2uY9sCzTkmP89MqMpaqvw
RM12UaBtwFSGLKG5qbrCbs+EtrjfagvEXNZOWslQGvASMhigCD8pwc35InMLd2OL
Y/NPetFe+jl3jDMSvgmF8zbX1WPZpMgtUuOTKZ1LsVYEtCANwi70GwdKU0/Am+xB
vHCTLHMS6cIYB1aMRGDOQE7td8payCZio72YUOk22mU4VaUlX1xhWJ6Euy8KXcgh
dadK3ACvVymLSCJ5nOeJlncIOnn7MdXurAsJXQ6x1rQQwudYuS8/8doE9TwKVKoX
FMdSthUHczJUpQuBKVuxMQz/QWqd0nnq1B7saD725Xsa/S1BuHXWrnZF1l4HZimy
FlnbxXNqk07Q+twjzQ3ScOSb16+TXxy8vA2s2BbQmrzDKs4T7jHXQPBGkXuOwR7D
SfaWvX0ivilllctYHVSXBUQNwzGCd9ahGLnssbT+qG2bHfL9xbXqGi1AWajsLD+p
GpeItmK3LAvYLr3a5HSmdLP3qSy22m48SEFgXgq7cl1xFAteEaHwA7S5Tt4rJqlt
OJQVO3W+jHS5zkeIUAGM3gTBKzxEUZukJjy/MC6I+KkFzAW13CdLsGKW0dmH8uyH
z+eoo4FKZGz43bt9buApVwVV1HKQo9wLcYLO1LTQ3Bx2UbVqA3DpNs4zxBWw84Lo
m6rlhO8MsBmOHew6sXuUzai89Piv/2GszWE+zUu9FgrW9DwnxEjXoAGSnbGA7IXS
XjkZgoKpg/UDXgCfZ55l5SmrAZy2dJcrzYCLNn40wuAO20hcgUVjGpeIwSBZICQo
tok+GIvtIRSaCYfrdOT/0yW6ZzRHIVk1VuM02ZEtoDAY/iK2YxTv8pSXXOxjJ8D1
PhzVmFDNEcuQ+bxjLry4fHNkpHEkagPIayyVyhu1uHvXaEQ1cVK40AWg6uauGNU6
943YvMZdFvSTBvbffzFEAbKTvIJFLEDP3EJzRUsDWX0cWeFjqFthFCHCTeQ0jw2H
Yjjjmfsqm7bvj0mYmi36KMjQ8AZhkMjTnwvra2QHqWIaaa23l1gfQHA74W4Zj4DV
JukGf1k3M+E9wOtCYekh6JAmENLgXPkDbCpExP+1MqMWU2dNBSvwhwmtvYL2EPpS
StFOjOmDK+z3Pyn268Di5K0kzHEhOTyGFwz5QwNu/gRKpkUuB5ZD0lgErG3p17xj
Gd9apQiJI5g/IEAjcaX8hdBQlcyzGA13nYRpW68wB6a8jdj/wjJx1zXBc+z3VbAa
v2RSzBnBcISm3CNrFERib/mARcx5gZXtnyTlqKqYb7avhg1dC8dzrRHzl7LlrXXM
TtDUMt4iTn4jBNYdZpV+V9ZFiUJ26SPGZLhBvInNecp9tHHqsiXAnVcG5GDadb8q
TRhccAlMnMx2iuiz4lwhbWih1mLSTmxyiFJQBPn4ysDpBrp68K0bgtqljXv/zm/e
zGjqZ/GSjp4ykd4Na0TAj6e/9PTeLQ3ETezzk1d1EP3xztPPYWNo3xOLPh58+8yy
shOp5VuPH5QFNV+KSJbtE0OXu8CCLOviOs7GcbNZXKZDWLO4EIMWmZ/plW1XPg32
GF2IJJT8UQkNbswWsj8C/MnKj/me4r33bOCLVKDR+Hsf+SZA7ErU9zFQ9f0Rqagp
e0kDulZqAHwQWNVE8W9GdCxUC6oraKbBkfgnTlam4krLE65xkVscrq2lOh/2+Qu9
/RR+48AFmdBwTDMCrc2wpbf2lZmpxYaBAahpD2Rh5R+CWN751EnEEM4ZbSKVsk/r
qND/brl2ccKP8ORFmah/+pS7u7WN0b2gUaiDF5/mXwVxLMRfHlYC0qNvMDkvRRoj
UqVh5Fe1qbc+leXUoQ8hwdhZaMEmV75GyPDnR4qRAQXgcIN0CCntJT8DuzWryxqV
PNGHVtVclajEConwMky/fKF7i3yrTFw9rR1AnFS/1wRPfrZfW39FSKQcB74Qh7bp
OV0yr+dB2gzKRQVH6u55T/alrfbPnF6+f1dq8DQtDzn8dhFhjoaEj3mTLWtE5lcx
bOWrpwCmRYsSaHxv4Zmo4fxhejBobHlAbMTVbFg0RcLpgXGfTc1LA7f2LXrrSwd3
LVwg8H/lCHhaFzuXZG3vBvoxBV0FExrl3qNjhmHxdP26n4OOxzPG2exMvuTPXniv
lw4YvZjxfzEJ8VwYZqsAv8spN1BvHJlQJYJVHhAtSgmGiBGgR56hoQ5oDOlbINfe
JhIXNVjpD5TV6c4WRr4IHaxkRxuGTk9A6+kbn/TWD1KuLbkgMjRdZb0VTMxMnjUc
FmrQ6l34MZjbQW7B2dFAEHxJrehjJPt674hOXk2kQtlD3T40ZD9QFYN/Bn+IqAhi
B9pbkCNp1JNYkiqSwsOw7lSJPPPWuFfsEkeI83epirGbUIvEJ3TKs0vmgbYK2HBV
W1HuocD6uiyjfSAj1+XYHrBLzbAT6KLZYK7KI180ulmI8K350b9S/QGyYVpnCvXx
59sOOIx+HWkLVEofUbbyvXHK6J4Kw2cZrgHa7gk3KQYz/1Mde+k+DK/zhfMi/RYT
GfaXGkJ3erRe5ww02gXIv/kY1AkFgPvVKv3ekSAshTHvu4oBlgHjUT5ISj+IjTog
lkVnOQUsgDnP3xgXZG0SCcJFqiUqKrBzrj8au7jx7fXNtxcgJPhKD3dzQK6YfNvu
bAWZd+PA/FuA10DRfoTNfnXOhp0d4uYn/ih2Ay8eoJpdUq57OutWOL9NRJZaYbNJ
qp5FvMzhRILdjTB3vN+RcjI5qarBG3UzjKdtqpuQ4x6IwSnB4TRxWMPx7ZnwKnW5
+QzeNbyGMwmVEFv7zBjfJf5YYCPkFk/001kFaYT/b6cqsbUsqCnFZl7fuYT8es6h
1Xj+lxWarNZkTq5hae/i6/bG5Arc3VKFbIrsKpidtXekkuufRxRVEvUK9C+v3iQs
PpebnteTZuGucxcF+0BTEvoINvkW9u7IrSOB4Z/kN+eFX3J7dugxbBFEgfMqKITn
zBfod1XwMTbR6t0oDbcLGrR+j0ZuHx3Uh0ktjBnfU+HRoMpf9jIaoA1yOvweMwoY
28vEKeFEhlobO0Hqw8W6oLfzkgGjsZLCiH2IuyU4QtVTs61fCKX92ykvSELxyFcR
dxnMqibGiGGA5E/YOEGdKPAWpPmgdLiUY0HksCousVyv5vhAhUmnRXjGo0tJUskL
pEc0Lbfgm82B3XCY/qcMw/kYtDcv5Q4NrGZN3Y3lZqGh5eh1/xhcEUcnRIIv60Fd
Jh3CNwYR8CrNyuE0RGg93DW6xJDzdNBuZEUkUZEHrr6uzcfnMypHZok9eUUxLoUN
O62wN75UzXlaJQqxbUkPyewcMSCkioTyU3+PAOwO2SQPb8/+4jyI28LVRBvvF4cT
2WFzQ41sHfcngwfTjaKvbl/FvxckabRwiEJtuHRRYga+D6s6gdZ5Vce5u05J62Dm
3xLZCCgKT9978yeUpi8h7i8wnK8nN+tXUQWhzWyDgK9oyX2yjzTd9tyrCYfiT97N
dmqa0DssE/QIEyhaw8oH8ZT1S96qMKkAfaXaV7cmjnFghRPVt0LIvYJnyA65FGFa
GWIqpcBSya12supmdOGM0qAaIwqbj561helX0XvxElv6GRw2+7HKvQZabU07QXKg
9xpC6gfXzEgCLX9seJmCjkwcODYghRkVVkAMX715GuDoMVsG7CEhPaPE8BVs0dWu
xcGHuiCVFSpjNlGD7jO4sactHKDdy0wZaQLzEM6QpTckjBZMmwBOmf1qKitlUPxx
SbC92prtNZ86uXXPVMBLCv9rGJNxA4Opc3xmUjLSbbyUWF3YK89QTfg0tEqMdfMo
Vs5xzHGBbpfNYSL6ftvDdX0D1zGgneTzBMzF7SjZmOyl7e2FTStqzDIVt9xcpfXM
sgD3vx+SaJsCHpCGkoACg78HXt7u9fi/uNzQ/LdL0wymsp5TFSa5NT6jqbnjZXTF
sFnyystvCNIPxLVuXOESBhBebuBUm5v+QFOVmD9kfjMtfr+zoT5l0xmushdL9RhP
NhinHLafLB1lKuxn8HtisHlfutCFU83dLD7PPROs6iRq6iDAsF4Ar6kUwSI6iyIA
Z+ZAp62guu5828gDbWv/MqSwgrqDBiP9HO2uYDP5AU2Zk8QxiBOz2Cx1RUn28iNN
whfVuWZsdIHcndFmp+SM6LLreSlOiJ1wQujrN3Mcpl11o9cgDYECm3bg3W5GjOoK
QnYseaQHtNrfTEbZkNxRg2gcUHTPg3fH390FX//habmAdJYQuFhaooekGl1Lpssg
ZzySM8CQCmpJNKocTEPceWeEFwLeraFZypLKQXgYW2o9zXvHcE0COQTn7srhImLe
eSVjFIqxELHPX2CymdDWXDjD/owHXif0OAcipxjqvkgkZqgX+F3SIAnwTulAFioQ
R84l1EPg+Y/p4CHAY1Q/OdOfxr6jKGsz0aJLHebyi6LowMwoP3ej9rI5DWnrcxUo
GXllaqs70kljZ6x+jEgKNi8v/X1nsoAWAvIer52lY+bUsdB2Qc1NvFVghHgNP2Ar
V2WXWZJ3AqQol7IHqyvkHy26gTmWuze9zqHsuTwGTxNTz0CbWlAzRJiAOJQ+XIju
nfKc5PLLoV1tRxgfvT1zb66puQoHj88kDYISTBWH+pLv4HVCaz2GnEdrvSSZVtZm
vLr0mT65C+HQ6u8fHy5qUB4HXvutSsoHVd5wF7i3fcRvY2kq4j0hQld1cnsxuY9d
YT22/YaUYwbYTXyh6KS3k2QEcsjo69g+qekOXX+iqzwH/KqJkvlKvC5rWSfDjir6
BF2Ii+f8bD+3KaEjzNeAooJvFlck1Go8M+nnShBSwwc1dWdze7t3PBpJ8DWYk8bw
LCmezL9cK/9ra0zimcvrtR8ogWPyHxug0zwmzkH+hqmZ1RXnRSPD9XzxTuwlk+RA
p1VB49KSj5KJ8sDjAF5RAzaGI3Y7KT3SLXixfdXF+RqcsYKstdTED3yOvqyZvThk
WXn/RiAlhG+kgEweGG+WOHE6JMMg0rMKZ/AgEE55xgXw8elNeZUnrllrRX5NpdOc
pMVRyU3smpKgu5eYeabzypmewniyCRK7hY3B7R03DA+3JlVHa7refJFo9o6oFC4j
l5YP1QSqbhNBAyH38PcZNd+PEGWxTqaTGPI3EzPe14CO5On54v0WwlswdGEWQQmD
Ot+GfN+yb5en2BIC1ZeFzBff1WNFuBAzXw/bF2OKDwsJ0TfOAA2irMioyxNArn8b
DDPxX82QsOYfOnEBX38mK35jmtJD9nyE+CHa1Mllapn6C7SEdaHyKQCLjm2sXL73
/FJBnDR1WkZOeAmHg/JOKNRK1LN+uG7lFmcwO7sgDmnwCn+5SdXoWpThDk0D6srV
z9flRDcVovJtEDDchnGXMeaUoiaOjDVc8Iln+s6gwN2VKIkgWzAWs/mCfyaCNN+T
4X36c8Q7QVlmjzr/S72SOA7D3KvW/Kw1a91y7kOb7fGhghZcVckbn5NXQNc02lH0
1oT4TKOL5AlfYuG4m0OVMtZ1yk439xVaWSblteyIxCSuaMokb6r3bUcrSG4HdgQ4
nv3c9rc1FjG97MII8YK5+AvRC9leCeZdIXxGjWzZ2AzNguYs+81uYHsyOz5hJ9SH
122vn2EYlLZn89+mW9QLcGx/JOg9FnKH5mlKWCc4eV3VXwf4waje54+1VbUA9/wS
iAaNht+/Fsf2e/OQXEUy2T5Sfvsedii8BdkaghNfXTP4qi+/1gAXJrHMKcEDuyvz
T6JnsHo9c1te/w0YaYZzPP6dD++m6J3oS5ky1ZHcsBxULlwvSjNF78djESMULMUt
TFNPEhc+TwfH4+ibW5r+qfoTCSg9zI4zDsddJYq7hEigJkrfaxCsL4U7gcgK1g/e
xgyzMiE/Zqq/kw2vaRufCm1HfeqArdU+4+R5xinpB/DDyn180iqk+gfxm+mNZxm6
lnc3VepzSzYWobm4CnRmAfnB1OZvR9r77LwinftRAcgOuCgbQAnAgtNcDnwJFkQe
bKiI3Sp33SyNaqBKpi4c9F6ZXihzxLfnc5Qj5VY99ndeBjB5K/GuM/O8SMMOFn1F
gzjyjikLjFl91anWLPSQ5VGsJq04JgWzmDJicIgCfVcIwavAZdx6/TFVVEr2u5p2
PCqxfdjjPPW/yG3anwx4MVKRLOsZCyno9tbyPphy28vfFW108NNZc59zs9n+TXVM
iFIIffTvWM/quOyKYev/GbYZqztHej7NoyPKafCc7PV3y1amGHdAMjccbsjaOyL9
YYRpsXhjROs5FGQUDJqaOV1y6iRUCfZR4IyiMYEchsIFTDWg4gMkQSQtMF11gH0K
UKxVyX31pU1siFV6vlNFvAAhssiQqSdzDQWOW2pQbI4t8gGoT4FAnXemnuhVhSi3
n35lldze2kiuushc/Rsl2Fps0sBlse8YcAHx1J4f5ZNUUk4/192jZvLDU05kr5wK
bAZafxYXjAZjiEb7039chESN7DIfxPnOa3tN0eFCTFSXMis2WA6THi1OtgcJXMCX
2CfVLePOqJESStwqjall4V9verJpADDgtnP5C4NoR6sF91Gk1bG/cudgkGxATXea
VoLyQz8MBKIafLIwj+YCdcR6WPF1i6PUCyukSWFa+EPQLDSbYXS+wNgHdmZXhPw0
ikKGrlT7PBj6dtr5g57yJNEWvB2u/sbY2vfvCcMcrUMzW/aobsO6nUNa8GqidVCD
eBoyrAjTPN7FlqICjFav4dTc+v89c6izbCGD7B9pnOz8FIDh2WE9nQL5EyEVBZGI
/86zB2In1BF5Vj1u7Ljh5jFf2D/zdn88gQKZmAzFZ/mPYnHYcQSHewyfdE7YzmTl
3AzlYINq5dMO0th/AJnOV0B30ebeCDXbrfewNyfSFH+DipmAyi2wJVHwC/n0NDJh
rat/rp59/+jEMDIs9GtFeo518ECu/NDcsLyk1Y9hA+ZEwE0IFoWSHTj6HqxlMIiY
N+5ohGZgEmJgNOUVskqDzEGUe7eElzz5EbDRN0aRMPSCavVs1CunszFzhQE8y9Ke
3sgUFgrvLPn/JmA9IJw39sGbRd8sySyA3WQBSyH/c9LQo2lLLaODNk2oN7DF4HJJ
4V3nRbePlkeAaqG84ORtDd+Z1YHV/r/ASk+zicNf81WhO5FvwmeaR09IBxKlX0CY
juMtN8glfeNK7n4Kk5V4KDBO2PpAygSQtCiK5VMqm5nESOJXQH4PXBbV17GryZ6T
pcL3QEuUigugCC9xF5n3tHVnlXKjDpC+59Xj/iVoF6WgFCykyotNhiNblnqQBE4W
rJ+W8XWYfxl2FJFHrOw0eF3D6pCNel8hHKhsECZ017kUsURkyWvdILZkIYp0d/gH
pKwU/OYrAgiDotF0T5vcfLV+GcVCn5qGQJ4igSbipZBVxggo5Jb4Nnsmb0S0Qji1
h6yVhH4cdyW+4sCm00OPR6Dv4CNcSs0tpaHFhgyrAerwRblbGHfyqIo0WPeIx/U3
/jn5ceu681QmACRvk+8aejCE3cXl4B33S8EnQKluaBhdzG1FZuHneSTugspjZoME
3t8A3eg9/x6S9d1bD5kjO2+4oHrJuBKcvdbGWLuvT2efRjJHDzS1Nzo1Mj7h+eoj
7MwVT103cFZS/fqc557Gy76PgMUc/iP5VVzE0t+4UKJOwgciMNzlJW5nNdRj7GJL
YBL+Uc7d8OKne3rG1ToKdQccqJj3W1LnMGf+qkqDczAcLfsTkYGeVWec5DU3xgKA
pX842/MrJcin1stqYXf0VMA+X3AOFb1Hb28I2Num1TXM4nWj7uutaGTKk0uiN1RG
396fHTFVotY1S2F1psOWXf9LWsI4i7rL6ZIUW8IxJbCrD3D9emR6/DusZ3841eIW
odbqFgN4azqfmalnCfjpGwTXFNT1Mnve7dXXL1cm8LrPqa8GjD/yivOECi7+dyXX
Rqf38iwE9HYXYtCzMNskq0dCxbHejMcgwO23ixw5jHJCI4tsJ+Ns3GE9IUHydOxG
n8FzEm7zyAwdqheuYzVazUkJudxDmj/0+yhG/MQANm2I6Co7rg9wiA3XD/lmByvz
x4lNcRqZqxcpCpYHD+6GT8Zfd3XxXm589RSXD26mZ6ZZyjt1GRsU4QHkBheFQtFv
RIVy8SwlAzTNntSffmDamBSkGEbXhGxtR/OGBSiPG0PnzKkUd9iCkAEUiDSn/lFg
wV/px6T4dX4lpswzpdW8vYr1RevuxsM4brnTkR54AloQf8g24XzR2a2HSknpg3uN
hNr1e1a62Y1wGicyFZS0FzjsOfYFvHlvED35HtrJH/SgENt8aZfyFCT4GSGGYfKK
fbY448q9GV57D0FvzNEZSONmDL+hMGcSXUJ6xyN0s480qPXnUBGgo6Xu1/wYQseT
XQ4OS9Ihm1/V20fhPIfKxVb7IFHTZYx8gpdYW4R7CfLnrhvDtqIyvSwht8NmMDzv
S11XVLIGQKMH1dkcslDPoXAUDbMmUXkHgPoX6IHLOStcI+A6/f2WzEw8zv3pR5yO
2FFKZZosPysnicwrHLp9/UTSjbeA2OmX+Uz14HIK6VlrqSx9YsS9dg4tiUKgVw6Q
f4JCKoO3wW7bPZSHb2xwds9nR/Cl70AYd5TGZSEJNIfsU8+lTthF1JR1YLPYvDbt
vAI522Qo9A/jACdBrrmhetMLyw2qQ/q38NKLECkH651HMrhpANrgg0QQh0t9idOb
yyMrJsR3N5khefbNiYk2X2gQqOTLJxPUJTG8YDF6UMECtwQ53OVyx0zbUdwbk8EC
FRgKI9/v5TO78fjOuNZTrlAmAJmW+G3lgUfuULfoJzOiCJ+JFRheEt6Ihzr4TTKe
/vtwOTQyjtG+DUhtiGRlfAPQRU7304j2KaXBWitp6xARXMdRWztnmfaP2MEBcj+a
CM54AdVzB87XB4UR1s/BQvSUCc5AKbfOnT3oWPUGk8nA6Qb58p7VgCU306UrqCzg
SPifo4Lion4qF5nR309E6Vcy+aHJbEQj2BA/eoCoHNa8JV4z+d1qZOHNi4PTP4D+
t6klGyNA06DJKStJ4wNHDuwLgcskEpeoSo+vYco0GbFPnsYZY/ZWGnfft6Vpp1qE
a95PgOctfMeiZtmi77w2Ea5GCHJT+OCIJ9a6YZG+R1Tf8O1DFR3vUQw6eStBQoXe
CP1OfPA7KPwTPz/dmlBDyMnKuSnQ6CE7nGn/Qpq1lUGAsxCQOSMT5EsB/3oiwRO0
i//wXvLEb0zIQCcnsTXc7lxs8EQNInq5GcZw0+GtQe7sCXxOyYBzRvnLJEvcfDbb
gjoBKoOfFX8CtB76CK+uKmym046k9J5f+rlC8/bekkbLKwkwTaonVEYVbsFsymxE
8Ub+fuiNiILMlW0SwHXF0UYS94swq+pOdlLGSa3CvLxsnhjbJJR0fRWQ0Ek5P5G6
bAjSEbCMUPPL/IPEqD1ZHlS42QJDMF4Y45WWdfSx2NZBIo4xduwElUYh8oIIxv+U
52GLTouuuV6a5JGdptsI9r9ldwxjFuBFeq3JHMBnBswgXxY7+G+aDxM7ycexR3tr
vxftGmGYzeyIxdBCq/eg2TYL0ZzE3YxYUAc9dyqXbu580Mh7sqfnu+vZkt0BVxou
5szs3rE0Uve+oOCJj+CZvw0Rheiaa7cD1wz8B2oufn1b/ndh2gmpcsQF3hz6+NvU
42U7JsQ+r7/fgwrq1+H1L4FqeVIyHmdIIupSrCk8XKKzVscCHxYW0oiGUBcRNRgL
vYOJk3kdbkkkYBbNBla1vzDmaKToe4ZPNNG36nOpG3Caf4Fq7ofOOb/K0pY3b0of
cyPBsPwtN/j02tR9s8V/R0YXfeFw7oVfWEXtGg5cvTTgRVQ9hYexZUG4ASK+Edm0
ps5vGZx11asmhXv7JM+GaDUyje2BKpxxT1ElINltdbiRY2R3UaJ4sw3/VmG1MhNg
w7E1971mNfHoy761f36w0W7MDaKCbsK7UUI9UCmKpQbYTlR9Gshf3ZTVley1+S5s
gWAMXwcTMpKUpZyoZq9sNncObqg9wou1N6I5O83pnb7T2SLI5sAgMi1mGFLwqj+e
tFzC0972CbG1WKhxodZDQ6ulA/NEoBBZSh3WlyW0r3A85MQBWnj1ds1VvQ3IKfTW
PHmJjPkpAeq/o6ZGfuCmtZaZnLw6cmqD1xbtSGlDT4TS6jB1hn95OXzjSA3UtT7o
ZMVFdpEd15D17vkHr20N79msNVE4UIwGy2cwRsQsLxp1tSBKHwUM+Oa+6AiDqLra
OMbYB7ckSSIlmDHxDbR3el0ujjsATIU2lHmsV7PVLNzYkj/1EVuPaLVa30Oavk0Z
tYzvdrPVFMK/TdkZz2SiGLJR+nt42mrhwZfSRRgBPwseX3zBTZCL17EdaDVQFhNZ
+/dXeSuROdsCXjAHAM5Mp2sz2qGe3mLmDoP4wyh9JtgRNsBq/yMBRj7tOGh+9ka+
tERNoMtvfakuu9kyGlnKScveoSjphXny2/fOH74pGpXVeHxCW3ZyI+73lzJIzRAz
BfkwKi/cDQhfsQfOcRe2AV9U0OnGjy4F/gYxQZo+itUxJUhqg2oD3kjf1xtOENzF
w86j6HmhywFiwdTnTFxmIUZQlYU/veXrVyVFLmQJ2MM+94crJ0T4LHy4ueTH78cS
RmdShlu90Wj04InzXAMXkDa7047KwzHAoKVMdUaOojsIobVeZAA5GfDxpMCiFXD8
jTKq6OZSQu+K31HqoxhKHAKnFKo/oko6IZ6Lb54f+k1eoQA68OaUO1ymRUbpfDte
9jAW/lLsGev8cCxnTxVo8HtkP+GKxJsWX6wwWoQH7e2FUlqFYwS9RVKvYO0iDW2p
loAFWBV3r3z8agidMzvtDJ0Kps4+VrVpdghcSIBSKXsUqjYonRCVvxuNBwvwFNuN
t19R2F3A6nX6/PEzNGYl71kVV9xH8NONkf9HURubprxsTBChLAqVHytc3WEjObWl
eWdcTfdET66G9KrxtslbC3igJBkxZ49V7lgd2b9a2Cj6L3OSIWqQ5Hs0h0RM3KDD
+Db+BSXbnuixVOc8qD0rIl1W8vdEa1aZ17pNSDI2UyxHIwcoklvyuK5r2PfEe7fV
TjOyN67E2lcgcEr4XR7C3FzSPSThFDJXYtPlVODrPJzKFrBg7qJPjE+pztBZptHz
SptJoDzjiBjDXMBQRUhfDYKG7AUBnItAXoctPI3rkBa+6QhX5VC2CBg4/kz1SfyW
CSOCS83ne+x7bOTBlm4URvvpUeafSTJrWXeD8dr92ez2Vtz2pM7koCz4neCbkdkv
/R6Z1yuRngO25Lh5kwOwo8jxllUVrpi9PnLPaCwIZl2Wn+Hx9e8RSRxh6AQd8gT8
iO2LQfhc+Pnb1+2YqRiAsNBavKLp+4AazQ4h3RTcjuZ9GRp8JrMa/rDRxvfWhXa8
WdmphqfE1z4Q/HlSJiGHzU+rjIB2gdnXORl5HvWuRTS/a6ROTBKGHomquOpjADgU
vbVSCK/Drdg/ekg9y02BOuw3D97TjahrpVomks6Mrw49FTHEm1L739sXE53aNoWe
FxxvYMKQvOEyTFfQmRphhdgjNuT5v3pe/ht4QkSDpJ9TQZoQZW1wuuggWVGBCzmX
ZzXlZX7hWbjKkNHECia/yklcPg2dc1XLmcjtxMzaghpRuRi4AGH+Wp2lT+MO9CXT
nrjnxTFYHEp8ERXvcxqYhHzbj+kZwBADc7ff0D0V2eIZ84lDpJXEdjs1TPOPw43G
ql0s6p9DGBQ+MjtzLo3uCLN8/aOqjj46MWzP9RBuodsLiU+iKXhLZ9PIEdEYeGOc
4+mFQmxk6rGIkSI0mvWTLLNTP0P3/r2mJZ5chdCMqYMfwmrZFxtmi4m2jiSKkA1g
RaU3fS2+0Wj8eZU9+6Ue7Muvkr8/id0OEzNGODOjD99KHzBwRebvBqpACOorw07Y
YXD61fDAs8GtBi6HJ+DJQcGBseiqZE7b4qNb2Wa3RIrwCWE9mZd4PnxxOsvQujFq
Clh95MBx1TBPx+eT8x96V0eK2BT66PdBSfSiUtIzzcfQNvM0Rla+ORg/7AARmvvT
TRmb3SxQisZyxfRshdW/hIAvPh8tzwFSkVtdl+PYQ73yWeNvf1j7uz4ld4l+ZPpy
8fzsBcC370UM5pcNIjpvsXwETD5M2+1sHkGA8CEbLTjeGKvW+9MT+NI5h4VeVBTs
zHtD6xEU9UGbMNQdWamgxm4hg7OjU31ihup0lppMfIi9WEnPdcb3r9CVoEKHXCmC
6coX0v8kym3zDGA20GJIHC8Ul7jxER1wi5NBQ4QqKCivBIArW/XNAxFRowjqkbHU
fDmB7MxgiVAkB8ELMIso6Z+eFpYTllHVS/XfXSWaTDLaCCCNlofwXw7qyb5un9jQ
14tVIdTCSZ+0YoRF1ReY3DQkQBHmkCw+wnvJHjusQ8U0oj2EsjS9YQigpDtJwDgN
WqWdDe28lSJBG6WYxa6NlgacXqp0XEX2iEjhXFZCOKm/hAYTWviijrrhUh5rzfAB
xP9yBdsCEPpyehpvaDotAfCR0cAk3CXWkUsN7RRoymWs86IWDOsC5IfenFPHqhcj
ptpAxGwWKglgp5+qi8N6AlLI7M46mRdJsylFaJlzK6N59ciUJnWu70zlCuvPAR2Z
iQ6Ci9HfPf5/uw9LNKs69jU46LzuBWsEXMOb4/r8afeE33LTlrM5FV5iA8kz2qYl
jdxe/0BdDDwSu6KHuTcJy+rwiWWruSbV7PcfBn7nL7KXGQRvYb7dQSb91nD3QdoN
2qxNBsEcTNZMLfPh5aoxoAisgsLJva4uJ/3fTlFpXO0+HDsrks53Wh+YinBiAt9L
oVq7LJPb8vP4Q0ZislPQVafOOyd/wXDfPCJ+/sc3oYSfEbdgw2bsAfWzf71azreJ
euSckOCd8YlM+7ziVPn5jjgbLHFV4rbLakcTO1n26VKbpcRMQaU+lVFPvBmOGBly
fDYGrqadvJGPtLzTtacZj0HhsuPaPma3SdCvVOUh0muR8Cxu7I/vK/jWpJgyABU3
EqasAzQShgGvItYLaYhAlimYcuA9WNArjhaZROehfh5Nx9+LV6oFy4Lxx3Aa4Lfw
GDxVuQ+IhaFE9f8+Ak40YdRLvYmeJw83LtPf2QxYZbCJZwg+Ig+nY5K4C3bDNev+
cBEVTTdnxx8tm/I1UuAzmc9sSn5wL9vQ3lRkzYHLBj8loMShKYfeCMsBnChfakoJ
M1ki3/XLm1ERPRQcabZVYMbf+ZWuQsClIohI9eErah0WgMeEWGWB9d7VJoPYAY+i
Vet3pCIp8lireATBOLS2g3EhDVEgBNOnBbqSnFfW1KVRiAuZwEFJ1NHu3onm7o3q
L6lAml6JhfjjbfS4ag9k8uDz6eiGT5guEkRktr/8kJgrq9Ugj5ELcYSP9ngAfu/I
nxaU6ri2DbIleeNcUcUxWSSMxAPcTm00AzKjH+BtdghwlVpXj8XKc79LIWkuYpmt
C5SsjEdPRDTv5gP7tYO5U5AALAee4+n5fLl6AwewKppA4WibF30umtup7vYVPpQ9
k9ZtxcwF4uv2rMBrBIRbA/S4zd2lopzxk4kE3iHK+YwdBYwwmX+XmgN8nenubQaC
J6PvEQCMu20LcO+yYtxgmztez6Tgkl4ikYvuj3uMia2GF9nZ+v9Wniy/0jjPGE7r
L5HqYJ3o0xqUdq03lKCOx36O1W6M92p2atZKWqtHTyatxJbA4r6VsJPLCrqF4bJc
jUfqFl8CVEh29e06ZGkLCu8hVj49ze5uFC2q8a+ZTzZ7wY3+Fkdy0W7YencDEarI
94tObzYyE9LyP0mKZkrkUjv6ZRbeykJ1q2RvOcm06/cvV8A7FcAjwmiuRxIF6IQ7
8OzrDXdfavZxA979XFhhGrmtf+EiGLi/PuKHExcQyPAkJTrFrV3tv/ilfs+b+Le5
wFtcR54W/MBuzHQcfezGHZkqgCih+fRyQhivm+yDMUusS8UFwgLCo6jPaVQLV+yg
lB8t0ZMSBfrcZRHDDfElL1U9I/QWzYy6Y0v9PY0Lh+Tt+h9Y2GNa4tfe0bUGrSj9
vtrO0HoQrf2p+AqU6jdJsUhqipEVK/ak/eopKXTVv7hA0Ky5dJy1b01ViSMnqQ4f
OyFe6tOHyKCOUC+913NA2/2sG0hvQ5LIB2YIZCcXlL4slbnHUNKcNIvdCkwtM+FY
SoLvK/3znaVyQ5VblMXHrVAEatlneXzU1I+UphbdUCw27VAbU2kvaKUN47tzddv/
G67Vkeoo6vihoUvsOZg0Qb/FviDK9Y/MWwGup1WdWbDUwC++J2jTEoCCPLdPhJu2
xh8k+VU8nOt30DTVCSswzcLdVAvlegDIdQpm1579BiXIJgisk18eICr7hWqeWxA1
7OubRwHjxsm1lPoVvyesaUxjWc0Z4RgEPJxCMhIDi6nBifu6N4p2mviITP5LkqF8
tIYCTw5KVJSzGIdIszbBf7MircySa1DCN+dX5VtF9SWNUJOGmtDWi6Fm9BtVRxjN
t6LipcgLW39grDe95ZK1Ni47JSTRpvkIgg632uFnRD36nmFL2RiwLymLqeUQwmYW
ovwp0xlXCDwVLRxfGWQY5gnpwSHjL5V78vWLdPIUzVSSvftDyP4Mbl+2Gc7NiKUd
pj17/1M1uGHEOHwlQ1HnsdnXrSUdaAANB7y9ryQjC7v7uPg97F6tcnQKgWKIec30
Z7cnkfYgGHlcCKznRYWhwGqfHbYQNpur7TZFJcZhgWW5HP41BEmGAsXMB1sXM2DM
7468qORBGeYxY1h9f1ju+Tz7xwFCpHUgimKSJGoScCmL1WsABgtXPWW1cFPN+cJ0
iSZURYrFWF+lSeY2qRRv+lkRTMzSzuF52+lQ/L7lgI3UsUHkXSHrJifI1agPN5GF
kHIuSuJKSVcO+rVjemUgqAlCrHu4EV3SbmcAZAuqfiHPCPGSLgbV919gqwNja/AR
3sQ6I77HY811SPeZJIbOZn9bZ2Gvm9F7A/lRUCMvZ/I/0isDYNcSftJTozIE3nj6
blFNoV6PMXApjo+vLCTYaa4RMyAMcX/d13hr13VdyO1Ay41/oXU9boTBQGuDy+7a
joVDlR0bJSrv7BSVecXMTuxxtmC0k2st0Z1INe+8RYJw+gX24SriTNGEVB7WUUsr
PrNEOrt1gWhNPWKWB7sm33wug3vzJAQ9fvxIhp7ahnCV1ypMis1fPL7H97EXv2SG
w2v6/uWIBHgTLjCq0X/R5seGQQKb4fCjpP73WfwhnaBP6MGwaicE71EaORDtUIFa
tK0ymi3OMtFFNRh55xIU2b+A7M2bx+4p429ZHNEqkdyVFdOL/rTTL1NgAyTwweFJ
7GmtdXbnDF0Kp9a43+s1DjRLwCIK2V0JJNrTS78PGA47CcD4wF0IfAxQVLnkzDlE
0KbX5coEZK5CSd/TUkxAexGTn2gDP81GTo51YQ6k7qF+C5wWXpLZYflDP81ZDXuW
zHFh7wfeQeeNrEgGasa7SULV6RT2+K2T69tcbtYIELheepiPE0uU3YtG8mal5xdr
INVaFAVcvK5Wk3lYYphmR/76STZQKS21C/rdCWQB1RwJybKtxNRuwGKYAnq4A9QN
TepA2UzwHyNN7wQi2oqAdbyPrkwY/uqpcgBKuuv3uN4Ma6pN8Ri2iwFYCvr9YwwK
ymbBzu/BS0JFDKevnPX43pPYJl3w2cCX3mFTgaI53nCkoZyG/YGxHbXtueCZ4Dto
B7xB5S/EfHQ9bC2Nfg+m2nYueEhai3T1H+Pw0RYq/YlnK+nSV3HH0bOPbg+S/IUZ
LGMglB++bWgtoVqjsM8JD76d5CLtgdpxXMjldz/kxiPU2s2w4RfNiUZRNb+cRKVq
mwLIoUeQjBfQExUsg7HcHtGZ9UVuIqGGsHUN31ikNQF4EGPZLwaMLzK0g9arTE5Q
yt6+hEQHEWVAf+ve6khZl0GdwMkasb721N0eMEe5vWytzXzVDFOfO6n+ah8UDwmq
QEeuKWWdEIZl8Eb5Vr6IoduMdR2hUNisujQ9lbuP1tUdv+lOSwykrjm375AUF2qS
Qi9xzthxCNw92HHORhxHO/2WdJgjeCmA/8E/fVUDPhWEAhEhtCR44sTDtwgqNrIC
8OOYrG8/1jfRLEQTuYDnoPBgrYEERdYi2kmZQ4aaz8BZ0naAkv2jrbi+sAPsNWzT
zszJsMdt9xSvbetFB4rMmDJCqPKCnZPYu7cBSpIbwkTGKH2sWeEiFnQ6NXwsW1Sq
/BQw5VchEQQVkbolS8oc5WTvbBQfNqmoksjK78kB1OAH2NjWGLsvg4qHoHo6KYSq
f6bU6EAZj3ZV4Vx0bEoFpqOcJoIdRaYrmJ5+PrMyogYZ8ffgrpIxElL6GpUrc+vg
7EG00aHshSSkaXB6oYA1sMxB+WxmBiTwvp9IlL8I2Tk7jigMxotfDSJ3KK0HSRAE
atCQD++h8EcO1X+QLvLcY7TgFYpXjdwqU4lSyhZjV6nJB13eRE6NBeLRZ29a+7xU
E0XfO1Ix+9q2UnZUdQ+DNFmGymy3Ga1In4/xfNMUR9x4V/lXG6L1DeE0qLafWe56
qnxbJQQtHfctfuYCgpK1zvYO53PTpYORAFe3dDQHy7tFBwuRUTSemGlpXaBVbxUp
owqJVmk9KZNxY6dBtQ4aLUq1o4qko5mMthzW+kVrgs9wy6KM37QvdArzt/KhOhxg
lTeO6ZhmfoRLlwuYWqFKnNj5P31B7Y+XIcBZ9QsnKZQn23UjJXPFjbTFW9jAjdC/
CpzJAmmUZ8itTk6JSysGoUmwktqq2mHFq/9S1OuNINe1FNGPjFaumTQngFPMx2wY
suCj8VZwQbH2dn+ELJL2JKy58jzXwKYlO5mnHpb3bMvxfkHYl/KP7GCyeH+BamNq
FTuHqxh0rryl8G1NIs2wy74oK7Ys/483Iv5uwacBdnsXnHSjLLnOcYDFK82Rql+b
+srLH0Vgt/p+VvmexGwR/W+vna1QJapraAK8xc2KQgHMqQcs8z6jCdaURTwdKVRw
LE48kqBKLBRg8ThqGH449dpnjQ29gXaj/UcfakajU+iXVRx8Q0PvDzHmioM8qsm4
sqCc6jZrVYPlWbH7timt4+DSNpKCTSbuT+ECtt2Umb9pHWaJ+AVwNZTxO+E5yVVE
Q7Wsx7fOD3msl/HPLGyeNeisKEuXzY/UdiTPY7A+cLpNua3ypPkhjlgYGk3b/i15
bXZeZRQQMlK6E6a5TQoHZeVQNVWyPTMCJNnI7I45+jm1QVLAp8xcu57Qe/IXGwK5
SZOQf+cF25FYhSmqYIFOgVUV6exnkX4EwW+w71iv00xJeGg8liPL6CTMIkmlM9G+
X72KvTdPcFyrvYu8aGamBOXWMpYMSQQUVmc/XvCkxpCajLZAkEszuzrrQX7FXJWF
q4lIBKijOhS9YOu0i+l/JVeg9SFTNvBGD1E8q8hkhYXxqHVzrPm4lJH2Uga1pWX8
EqOVf1BrT+FIwCcSq1KCrFMWrA1ez8nc58rFL1QIVHAWOxRdcb+STQGBSaGpL6Pe
fnjQPqL3OoOM6BlzfqD3S2QvBtMDcsZT8ZlErBzIYWYcxnbjVr/4mgYpnVc6dgKa
7z252+eClJ7ygeGnrH4wxy2sTzyYDXaBEmZknW0cwvORT5wkuplOn3c0FsGoVP1F
E1g2oa1paGkgRbUp/D7/12KUeVJoS6IfaP8ud605lPp0nBbYMJCCo22CGfUsddAf
3skL3nk7Ufi2yty7goYSfTx1mq5gX2e2Y1oD+oen5p/XCG+STcHxMJDRNucbCaR4
6cx1LcokIYXMw5o2sqpuoIHIv0XTPNJiRo9u75I486+rodqz+4yB7/7pcb7hO92D
bADU0LMcrjGnHToxdzdOyIGzemKgeKMUJAhhgn6S4gUSaoRab0ciVxFRGQcVaa08
lpmi94o61NQuJPEWoXVNM1XbiVHDe7WidETQcIv4LkdBBONsXJk5yJ1Kor6rLucD
FgAJqucLmFxpNUu+Fumd0GopTr6zZuvjgheZzwyxSaPL+RD6lNyx3bV+KwDEDcyu
SAbrf1cHZpcBsOxOkXYP/zrkyrorx47X1V1Ohcz7VEPXG1IXigVOeyH9uBCi29wv
M8HO63T881Av7+3v0oExhA2QTZ1A9UfkvnF1j7KOceTXgzeSXNeuAB2rprc1sOEP
TepQJeoLI6SgphBRaqY2yLaWLjjYxqCrYyLxVTJt/yYMUk0+AzjMsZG/iNAJsZY3
dtjZSimsz39phyIHeg/2kZn3oSvAPDJyqhv0Glkws6TCb6uvXtMFzaqOjpfRGv+O
5OnaawNXE0p0fnd+PDixFbgwmo+ThK8XIta5BRNy5Q5HoEsn93Pc8S8w0JFYPGC5
I3WfHWSS1Wc6syLoE5/yfo0XxjGUdCIGkkSuu/8BSEE0WEuLsrDYJe8p1cjBEnKs
X7z4aou77jHrBoRvUZz/ZxGR3hexjqKfcbFFG5qmfPmBqrpm3mH6JZz1N/Tuiuyx
5PN8PmwaxWRaAdKcYhmq3a11y6MAB0TTPbu4nGqtcmA1bH0iW4xMn78fzyuMklZX
eX8PA94aM58j/QrLOTMeFs2xHhDD8/dVsKXaIKTJSZgVSSaBMGmvdy2WrmnxtrLd
4UDMtb0pENJfpbMFzSSMt1Qxy8MBJZBGhFdEhUnxK9tPngJUs17y3FvngmKTOiAP
dwTfvCt+hjRUnX0zZ2Q8WNGmd0LTH306IUKhl0O1rj/EvpQ74McRNAhFqk32JeXU
MfgYniNx73IHMmHMTwR70DEiV1alITEG1dbGTyRLNFmbPz5ZxsewAFRqaNxjYkNT
UMSHd8jAxXnt1UaI/co+m34/nXvoQIvf0gfQhVRic2LX5QBX0bqk3OiJKqKgK+a6
gZmx7qoZUa/I8U2bb3/yvvJYUu7vRne8GAJmt90ez330VCJ8VpzeW0CWiG6CaM7c
h8yjGapNDaXdICYdchNf9p1eWLnLWRqxw+Zp+WKfXF8ET35Z1bI99CH/V/Os5TDg
2nLcV9Vv+Di9oMBsOLkTLfRvfenPtoib9EKn2W0lYjud+DJbLtfYo4GECjrC89bG
NCu2TqXMTZXcP4L6LJcWVpj3ZlVQcqvnc7SPbvqHnLvAD1CPi36Q0d5B63eDnsdc
0AM8lSphnXbGsGMBKw4EuPBYEwqKhVwJg5pFheavhYoGaZ981kSpased12jHi4Ra
uXzEMKMKUTk30FRMn94CwaSDQ6Ylj+TWO9ChoQNdwcM8qxJYxqfi7aUQs0oiOKtC
F3kNxA0jMHNi12f3IWx8cXXYeNs9Lj4jpR2aCcnoCkSCTlnGBis+DWV1u1aFPhpv
hlQBXldPcohlDsqnvIB7QV82gdGjiSVOftu//dYp7YndgdqbotcBPVzom0CP9kxu
pvyLWE2yXWS0EGMOH4t4eKUaj+hKaotL09OqPwaT4wFJo+kyDcKi//GMphayZyrW
cj6f0LN+NGw5ntVk9HldkDseAzjIjI+uz3nfS+eGcbs+3g9U2r2DhNGlkYMA6C95
tbFnIHz/l4R7cQzGCbNQJAEsftXrH2VLW7BGemwCH1dUZ9MYZpzmkHMXwuEznFgH
McRH2P0fVx/Ruz/RHX1Ur9z5jjXKD1UND7rvKVPbiqT7eM4GZqJsWZnQbmL4LyRw
XWbqFlEb0v7Peu7xkC110nj364jYTTt7ta4p6jITQsmLuZQ/gaDMr1DoOEoYOfGz
kGziy+ACFoEG1XHi6VdP9GGW2KXDWTuolMpNUBUiDWpJ53kvyvdm+YoPbaGRDbmd
U+3aUcwkZmmg7Q3ObLAsQrBawCVQtvyFU+/zosD9jmkS1WSAnm9CqEjnKkZgsfCl
gE8aQmlgoL62dhzf8hhKpbn+9CAQbUdC/IV0rXtzmQbaxxMJPLorOSaYrEJOzZWD
l5idiXdClwfZlSZgW4VtfcSWhhx1jWTDMM7HwofQMv4dana1v9RZ1oZbWR2WE68B
J8tOiCzZC8YL2PxDzyerVnAo+d+NNxKqGwO//bHB7aHPAw4gR4RIbSTzWR4gccFJ
C1H3nDK3aPxIQVwXyYxc6rNnsOPwF/H/EVykv4mz/zEtl4degQuw7f8gVKU4NVRH
SP6bTC5CRUulSn2tBnO5k1CaioNnje/LgCkwlyNN7xB/zREBjMQOnnbnB797OFNC
fMhcXoZFnZpnAYvJ0B4UbJA0hXQT/euyXLlLdn94nELA4adT3BOe6LqNAn9pgO0M
eXFGNIt81vhTVEPK/ueab5Z4oC2tfrLfdE/cGohZfU79ELfFOhchG0yLwirz5UYe
GaOcQULPiYui9j1jPcZZ6e/BO16YXhXD74l5VcOMaHAe7Gq5kY3t5Pv3uDmbBUiV
bFB7vK3fM0qIt+mjMmpMjjBsEwy3/+KYwz1NbThRGUnYsqmLRI6DRlKE2I9wCPuR
L4Oz5KOi1RNMHbjak+77KjtGadeOcl721TEXH18Y0R1BNOY/+/VZueoZKjeJbOo+
GMdkdQ8GV9ymiMUpaV8ToY2ALEaRH+iSGo/KM75dXoHTR9PuuQ3vIuiQ+BE7Hyer
DyPQ4Zm5K/RnVVOC9UGY37D8u9orVJrlEXRxDsL5QkDXRXUOzS1+me5joebrC0H/
1lpdp5dW1jB55hYIsxYtygL1b55ZpZiOPutMdx/CvBbvsNTLktIJ8V9Po6FHQP32
AuPiLHF6/n8MY4BIk51RD088nwX7/Vx1jJgfhzMiRuA4QilPVJjVz0lvnIriixf0
T3aSY8A0TIbHP49XpkN0F/OQcBPAtPSs6gOddGm+sl1mlVIr0S6Wh/ZPI5t7qOOP
pEHom1fbKv2vWMpUheEB0YzXRHks3GEFfZ/yK6QV9jCuwfPssjPEPpvyrblzoPM4
ag1hupxljd4jmc/Vmye+0KhTaHVI2j10T3N32uiBXxW3vKoyBLPC2p2EWrPRGjvb
MaVxcosXEjVqKkTLyo7YnFxdJaJh/1ce1pa2tWZs73eScQ6ml0iSWxuZ0JP1qhIz
/NqX19NlAd4S2R+KN8w3RC9b/7RY74rZzlReVvg8fyNinrHDmTIAOrMKiqQqrhLJ
uwF3vOG1JGXNkBmR/dWzMggjNOkpTXOw+bzEBeDtxPSChSKBQvHYhCPBPVrsuSSW
mjExRbFby6oYVrLBugczDdVg2jXqcN9JOvfKMIrdEtQ5fUsejGxyrcTpggLuaNTl
iYS5+kjQzihWgz/i7YNBmdL9ISHwita1xaaMVHFvDky8r5F4Ty/6swD+P4v+mpN/
jI6XqNuN4yaQ+V+dGAJdQi/qs5A5VpEhLf7N2qjjXXM5vDCdZ5zPrS8MqEzJAumF
fCqog1/fkvQgy64/WH37sjhXis7VTagmIC7qtA7qcesHCdJbcZ+5ZN1P/tVSt1X/
pZWWDNVf//yIMroKJczB2bwJNZdTzUATkcV810ZAxiFGc3VXGBrX2vYcqaUXbn+S
O5jTee+Xoj6kwmBMgiolFZlxlJqzyQdBU3w1L2hOpDn9GDhO43ZtrqYyseQhOHhR
8aeA0uoCcVgebd4md5fHaPijGxvF5opT6Jl7NnY7HPvyoJ6h0kORjK/n3N9ogROQ
jM1FBUwPze63ZzOa/NCkSb8nahwBsRECEWwLQBWVBJU2jhDkbkaZfJSIXOJIYeWO
ND8YMq4uTAbkEoEI1Q83AEeCxOYAvRC2tPLd6TAGHxcVUMNvExFF97KWm86TOWR2
xoQulGzV+FmTVIyZUqWXBcl7xjpgZm9jQCZbIiKpDov93OjHdr+nKRn59LHCkrij
vIxW30jrEWR670HJahOrGTbqys8a6IcF5oRkTXLAPC7vQOQqSXk8nplEvv9j5Yzu
pNLcOmL7UbQKt53mQ7YNtEMRp/Dlay4/Qwc9TiivwVDjucJdU8jKp8c5T8SBRycj
cf6BsnsLCVVlQeWtimJVyeaXhmm2o8eOxwjj3vJYLHQBsdZg3pIo1ndscK+25IMP
rA06IxwEIEc2pB6mfNJdsgrh7JeMF6ist0YxWvrKkWNWBvhe6nm+KX7fWMoQB8wa
s/tJ0+N5X4Ui9KJr84+b7YgYIBOfk8V43glIsBS5XuUOL5INohc/WmfrI9gF2ZpR
ZQPLFFZLBPvn4xmQla91rtRdRZwhzAUtvYtXgFlfjLn8yEPi9sppzebJql+KMsMh
X3ScmmJ+ohMoELLlKztU6SR7aT6AZHJ7o1BENsTJfs6RSpdOZfMqCJVHbh6IGrhR
qoVas2Yb4VoChBpfqEsbZMtJqCVIseHQODXtJumOj+dplUL8Ru3Fss3HOGr5ajX4
nrYQ0Vw7hdiK95gui6Jn3m47hHmZWtvL8HRgej8vHaSL4km70cZE9YyCqgAPvis2
uUKyEbubjFpQOaVAGZN8GXbcwFl9FLorjudyQVeLwZ4u06VOPM5WNzBZuaxg1d56
+BVNLmP6PTC+ncCEora+BiDVeL7+orDkcUzJRf+JjNib4BXSiaharjhuGlZ61KYD
VbnTOWAdC68kYTZOMMe2bQKTvspkC6Xy5N389B1frkrxQUxaByU5E9kmRBao6ZwT
Lr0gAiCSBQNCAqyLRb27Y2htw0TtJuUChJcnogrN6jCeZvB2jCaTl+C/Y7ayUmR3
zCHqS/PA/xAAtjZFTh7mS1jxDtG9R1ukrX02fdz7yzxhmiV2/LmYfxf2xBPEMnIA
yZv/yELaA41OjMiBg9XsR4wQkiQQreptBuW+GhssJ30bbLR1P07dBCHyRz9KsB9U
rieYgysbufjAMP/3FaabyK47QhbZCToSQLr2jr4bWCcZpoSlnxTe4zDZ7xN/CAch
bjy8umnQcbL+rpgVgboIxJWrq3QY8k4jtN6rTRaekdsqwGCNFwadYczhJ24kRsIv
oO/Y/Zv7nv3m8xtsXlxXMM7SSuS3YiG3Oh4IO7G55yb42mlBLykezxkKvC4UnrLp
HIdl0FHQFW8Kc1l/6BcYlL5kpWJ5t1sefROVxDtxkNQyqO1oO/rHAI7mfUYZukFO
W/3mZK6zVOvIHi23O3IrZ7qiMt3O7IXVriPT76i6X/PesCiu9NURRQCbNDtzZFyL
qi+1AgisueQCroPr34mAQk6oX4Sk+Z8a/dZJfq3+uFDMk3xuzC31R5tHlus7ffOi
2DJPenZHnT+WS7MLZ7iLeD/fdCIpwgD8D55UzaDOXvfejPO4FbDduuRYVavXeDGZ
voxfZreLCzddcKdaA6Fri6BeAjc9JjAbpI5GaiCXxXnq6pCs0Ki89i3IKmd1Fy/S
R5cXvgat2MeGLHAcgaxuxqlA1JfackqrxhPcjA2gZ3RZOewYSph+WiMl9ojjHnaG
dZCuQ9EZs2VWWAKf6HhkYSLrn98sVL9m29Nmkif2K9Yxa2I3tBSacadg0HmWu+nk
dPah6KHi013f1YyYzo4EZ2EUyB96aO7OAhSFSG2ZGM7oIMq6b1lSueuqgbi7LhlF
/VAyNvEs95ePTKdb2GWx43R+6WesYa+Cj0OCURyUm5pO2pwvLE2EgMoTQeSh+Ez6
AptVUAUmu9kJ2sQ8A/0d0Wlveyuwh5zabW/NcMDnqlIECmF4ACSXvhwRufaQQp2O
mIEFDWWX5MDj3/qfu5czDbsQOygMBMtHN9wqm8WnWp/GQNKDW5jUNdP6gRi8HcSd
kQeaBMDcjXd6pmzCSvkp+b003/7D9tNQC5o3pnqUb8ok5FNF5mdjFjekyFU3qkAt
WZ0YMdjqXF2b0TvjaryMFJ1yID9c5v8UGPXlqXsReQbJvseDelDOEkTv1jSOmkfU
aPL/RL6y/6v8IT1JXvgUhvYxM0vTYC9y2mamr2UGMUKwa+0iZZAaaPr3Mr+PPFmC
08B7Z5nNwumWpaD3YU2hxUifkChXwBsCv4V/XfhGRmuWcNK0VMRoCFPe0uj4DTJQ
67uK1lm/PZXNjpcApgtEYCzZ6gZAeTFJETN6TLPQRPF4GrWUXMUFqWFrMQG6EIQg
cvZUh4uuAPR/L6RPg6AabHJ2k5OpNf5MgaehE+eF71QMuOrMHCIubeg0Ov5JPrd2
HATqLmVugmQ3gPLnNKEHYep8ApKhAw01njyifFTjJ8hW7h/k6OsAeLLQcRhrr4fu
j4FybtuB3JkiYKgMpz5mg1WRbEQGnJmbj3Pht0NcwLkuOWLkz1cmq5TL1z4VANRH
eSrhjuF0YvoyYYadPTV3xu556jOdHoooede7KUuyWxKFfYWqNHqFiTXbMIKk6rE2
vNLHrdQ9o/fyXQmMoiQhfLkqSjVQrxeX1tEVdpB4U87yK5LQLrx+ZQw6O93FyIwi
nzYaLjwbpPKL7H6io3T/1d0pi/7uGP7GIC4gNQKLyHVRRDyqkDWF0uF/nzTcRtM1
jY1yzxS1RV6vU+Gc1iDbgy4RNCtGmc+Yqhxr74r9Sk7JQTTOriIwhAWDox9cM+YC
l8XsEF8lRoudID0IpWYgM+QLVVZUOsaF4uOtTHccws7dCj3+BODQj9K0ntU3gWWx
EzmgYOnANRqs7z4wR0pqxRwvvuuow4Z5R7x/csR35dhEAU2oPMDQfxXcECZ+Yq+W
jPkAzo2EP9Bqya1gCChCOqHos8/fFEjDq3R/5o1Lh1EhViAMfDVSOvPzC2h2GUvW
6IS/7Nai/PNNLWHSSEGkB02WwzPJjjkBD30/dBZzrZut+R+Ftu6BQMdl1azsBwfL
ZxtmQJTI8F8hLbKvwbJKIrqLPUE5L0RSuj6gABawFVg8KtqRr9KZQ1ffmo9Jz3eR
lk8RHj+lIPCLhyYRmWOYwPnMrovIJCf1AdaQ/Z7svojIEY2PHdvG+4JsSWu1jbf6
JMXRSfoIir1pNBcnB7BXhfDud4ak4HimCG0W9hJ3q51pkt2Tis44pO3sCmrjiALd
gzGrVEnFfsmmxNpkwXdFcaFqD1o8NxYpGDwmtuGXXpD9mx30F4Mgf/PnKtd1reL3
pY5Dgq/wEiuXgPw0KpGLFQmoDrGVW4rzl7abmJ+JpA+Vud8N8xboVTWDlvUGww1S
rjFtNU5zbg1wXwGrrD06ofqCzPK6ANboITR0P0TuvY322y8gEBS0wixJVwk0EI9L
m11k43yDRNHKR0sS38H/WyeWeh575aa5EV7R0qnQbYyf+ZZkKe00Tffh8zgbvotB
y9sc4P3NG8q5torjI6QZQrXIdfL9qO6bYPGISlDVvJLQkdXF//jyknX3oWGQpBye
3jHFuuNMtEeXtrZr7jvkx0hW3/nO2chU3Eah8f1dOYNl3x6tvwMHgti8UoP7vt+C
SC4uSFhAXg0WWMYHaTSqgraKqqAWEmxuhZqECsaglCm35B4wiAZGiGaPorMLA1m9
jxmgT+hWiqCbJD+6Vkd7PLUhO5+gE3LWyt1+OPmD6knW5TJSdKVdTidRn28tpK2p
tIfTCMjgPYjQ7Ty7EgUZd9Nhbb+LiUHMRM9FnZMxyWWdlsNPNBtfbJctsErp3YvA
9PHhoQ+JEgsU8lgL54W/xlt+duf3Q0Q2Jp8yE5noNc5HPXPWf0GDL4ahsYFAgNx6
p39wzVfiBFf7q66spPWxlRAmGv9PzBMijfyLLjW8afbeAny7TUKV5sWJrX1328VE
UHaTEO5v/fTBv0pzzgPISHilYxsUL4RhH3LdR4ECJv9G7yCabBQ7QxeW/dTb+p9y
nrdpuwVxbg15i5goMqR4+7XUx05DhCQ17Tkg3OfTVOtQ3plvjDNFLU7KdoXP0YG3
MeoOtZBrhSm5NaOSGGJE7wvI3+wkFPXP5rNJym6Q28Ubf7ii6/STDOBZaMA1Btd9
2OBFivFwI0R7WuHdLkChRe8fsIbR5BLAzzKd5FJpt4s4Zmp1OMiSSz7uXS1+Ij+y
gc0pa5upjt4juyfammf4mdlsQY/Zq72Vp+LarGPiyfdWRV2/y2zZ1HvGl1SMVjn5
SI+NcoP3c6Zm8gwmc+yRpLdDwKiiD7dLJgR52lrq/F4QySGWwff8dFO04vuMrpPy
gRb8BevmEycwYPgBpSKV4jfxyxbS8/KQmdpoF8QTjf0fTXxtd3GYhFEJXb1xKNw5
HGj5ddxQLWYUzIgqyqyf5ap7VLnQ9EK+lWUsazSVhJv1Ib2gtbGoVcLp8lBd9mTX
iLYqh2f/bAKWLjnU7twh/qRpSWd4xOuNvmECgHIjOKwB7c2ydPKpkgGaIolR1Ozv
baM8d/5jV7FiIQUmuMdCuZ7QIQJ77FkzwyPGWc8VGtv1ioNy2w52OGCDWQI52eGO
skP0Jwbah9CKa7nBsxjR84J2eg1yj7BszrOs6zQe2htJniCCVXzGgu+XqL+rqLxE
s9X0FUbwOyjjC28E5fOjwi7aHq6EnkTnFBLXPxCM/o+0m4pR6Seg/0C3C1CR4jZx
gyP9q6Lg0RcKQ1TdespuyBz9ikb6Y2FbW++7DHXFUDY7ZLzhLqDFrt3829gK8SgV
KFSzPow3PfaTnJfLMvZQ9Itk1E9Yt26TgbkxMDCvK2i71KRZmT8AUqyx2xkMcHqp
Hol+WFnq8qikmto33Y0fHMvBtrsbipab+jYoNZ4HcyNoyeAWkHL/gwciAf1On9OH
ze99rDjQWxaimV8YnyBnnYFxOMGJiVZ0G/JuRocPmDm8NZ6jP+p2OM2ClnB4nzZY
85mT8IZBtW44enff7xDH/g2zK3QmSsAazNdcMh9El2oJyW5ONnJWnDDbT6ySi2sv
w1BcxbaGOkhz6DSo6wtbxi8zjKkUeTds40mALzPeD+ALW28i49jHX79LLNXKQJ26
0VoXwJcw09X0wEJKBbYpHXug7/8Y8x2OztIdoZjfn2w8/6TcmVh2/MFvb5P97+kC
uj4ZAtZ01MOLf2oNxcXgGm+AwFoEtZR7+sEuCbMBcjQd9VDLNv141uIbxhcpC3Zv
f5vPbFn8I8NtD1dlOqrf1Dwg05IqLgJxq+TnjBl3f/lkU4O/lqcJvStxUG4chH45
4ySAMeQvNoC/UP6QTCI/Q1pwQgUkWYxZwn0MQH/NidIJKYHu6vQg++HtjLaL5EIN
1ZRmX1biBkkoTfnWOnCSG+qVD6YfDdqh3wicjhFTfbGt4cIKARAy3w6waq5hwBa1
5/Umx5GwWEVD7dXgnXfjCuxGh8jDNUr1BIC/n/xZDPHyL5BgSXQOJFc6guPU6p4s
rP5zctakIqtWu6QaPWIzz1aHvW0WFvOvY3NlBJj/r/Mn41yQk4D7+KRcZopmvhzS
/iQjvBZISL3r62gJWWolopbwYF8CH+11lRf/Fbcw2aHCEEVzYqxKwGGGf8caxu4a
0WlCtUeH1AvmpdGvDmDsRRX/tFOt+PmpaaaqmbFeZy0RSiMoSgCf9Xhby9jnSuIl
D8WMs37zNGucbM6/cZ5zyw85/vZf2XCoFWdG69uPMYGBw6zxok4GIhScP4yX2nvH
8Q0WARSQlLz4PUqK6XaIaE+wQPbJIB18H3ws2DmNOT0OI8O3f7JoyRrEMAdwDQjY
yY6D4+YIhJRTPl34h9rvZCsmYLqYBFUwpnoMQsbeTKPsOLc+VF8y1DX4kRzVxYtL
8YABPnDYzyA1pOVucoDBpBpxaOGoGHMSLx9ikIEYIKnelP+87CcglE2p639Pi9er
gbS/15aJf3vYZglRFBUGPDhNzNFeRLlESKzdKo2kSStqNpvwZvTJjXz4jdtatOmZ
xeMHZb85bAw2ztw70ySoV2hDSd1e1EF7G3D8iDDdsJLcMVf1mPBAoq9aUZKPy9w1
7YN5KgG1b6n5RaMb90I2WH9HSAUDGVw2tWLExJcNhnhropxQl2/mvXp6OeKLLE1R
OjJkqNeVMwr/5Y+DeEOoWSbj0eREy3vwuw0AGazFqwIjGUj0aJ6UXl/kPt1pcVHF
fCbyTizE/yD3DFz9xcQUnJ4MevweCHHwygn/0KP0k5Q02CKEsHV5NAvoKk8U8OaV
Yioow2m72namQhvxoDyivE46KBHTHZ2uTPlm7J3Dw5waHwUf9FFBtfACLaw9tni0
3o2ZUZiSp12NWCVkWOWDaFy/Tg1nXC1Axm29DUK81t+/CtlScBvHItWNTB25pvVs
PO57jk7BqgYN12/O7QDU/doIjMfjBsqeKqdJJzHt9D+Ex2c3LXoPN7oka5RI1qAs
6RDIVVRTNZ3OMZR1+7xgFtWFkQMIUM16qvBiJEGKwdZQFeM56tYmrQEQOqWutzS9
f+NuXV6sG0DB0xslMxH1kVKIEJKEJMsPrKepRSk9oe83IWDkDBLkK9t1YHh4asBj
KC7RbgfPr0nNwJWVD5ZQVssV9L7oBuXE8g/FMzOB9EUX61B/KdpTsd9hX5Fht4ik
k/yhX2No2HnR5ePJKJG1INn0e3++3J1BCSEfDmVfXNCFcVh3CjjmeKY3QYGQMT9z
b0n9oN17+ymu9Ug/v8puT0YOC1W3wJ+2vgBW9QRmTr+2Nu5JMycsne9z6B4OHls9
OUePtYNVu7kBQ9y8sCZ4umg6Ic1lZi/v7zHahMtQVfZ6E63c8dnxZe2F4prGmaKL
ABrGDCw13SJAW8LxGGnAynmKrc0TUyxmMjsQASNa9gAYjT0H6cJRys7cBhvfQ1jj
X+NyfP2e/oT+tUDpjy90oYlcItQOC1v8DtDRoWleKcpCGmEsgGGqLWukSHXzr3rZ
NyTPKiFoF8DhTF6mdTes+2UcX7QE0X97l9YvaBDcJLqz9bhv3H/Ml9xz8SbetPQa
JAJp8qc0E7mpg62GKfb4TXRBQ9uu9wPOw+FtxL55qDmm5QdpZ/NcEwWCkTkqns1I
psRHewYHf92sbIK3EpI/egaAHJzAGnFUS4awQYE7HhwrRgbxfSrcXV5cB8SQEVad
chZ1Fi9yaCkm2Zy3Srn9L3t4VMPFQYSXSetd8S+nJNdMvmJeQYdb6CVwuTRsYTfJ
wJOfh90ClBSv5HhN5z2ZImjc6bfbN6KIDo68Lzne5B5HgpDmDeVNeA68Pv2/XMXG
vOHV3UoMTZ0C9n7Wz6x42mgwRAP9Xi7cl4ZPduHisAZoKvEkkxKH6QS+0TA7vKmq
gFDECkcoraQt+n7/5WgRGG24R8Pn+nXA0rjcD1XQIom5DFD3Q2C9LmOsiJo8l3fk
NCCByHvB58GJVRyTKGTsV0/mqlu1/Q7WXpkL8uSnR+PPH7rZNAjAIjv2XdHiQTXt
rdu1tDqQ2q+gnlq+jF4Fq+fQ35iUu92HCbpZ4z8WUGIa2u9qYBaEl6DnslTe3OmF
AB1psF5GjDIKeOFuDwNvchz/5GKDhEqtt/QeOw2yHmMMO493F3TXpwJBobdubfN2
t4Cihzde1Incuz0tsVDrmw6pqAenSjYM+x8bgtBB3WZ2kEQuU9I8hqZ0dxBx7G32
F0ODJb2thh7MuCYCrwZEF8/aUR87aCY4dpQg/PgiY0tQiZRCzC6XkhxgErBhloMp
ntdOwhoSk8naYrFX3PK/K3CYmL7fFLvTtt5wKJTtNkDNdufKCjb7N/Pv8B4juE04
r4yhRO2eVRBPaxeWmALxw6DCSEv90Jnkwlh5eeHUFpW14YbFkCabes7WZcHnUuUl
wrzEVX9dMpoLkQ7KqHr/ylkcDfU+8QjnGMjWjDpwYS3BYNL+gGHihAcEbekf3u2s
Be1jonXku6Ymj6LGOXpe33DL/irI6z2MeY1QOJNeGShpkA/o5EKgeZNCI4ZEwVGt
QmgdWyqYQenKpKTaafj5Ns5mr7b+AskYeb/1w0fpN/NOdKklJ6aNZKV6cQSNjGjQ
LZfhrFTTFAfA2+5Urey4ckA5ocgzcxkuIvKMxFN2vE1FlDi83wTLDNx19is7b+TY
1A1LLddr5i1Awgdr4Htq3YhIvUAPfevXoccNJJMLv2F0CHZQOjB3IFkI8Xy6MEJZ
u0MX5o7Nkcz4/Mjc79MmkSwD6u7mtzlmezFAtqFn9jeWIeP6ssS0rAkQuN7ushoL
f50Y9e58GHSf1250VVpqtZTYHwMAOfTr/v7w+tIQ53pCU4dpBtgDhGlxhVfFq0v6
Fz0TgaGVC4T6FrtQJrLgag4s6ig+SiF616WEA2cgjAczcdU3FoIHKBsZMSxS3UAt
J1C31cka9x3M4/Ni5r1QjCRxpUGveo1qRa7oscviVUgh/Vh/s/hUVJA+Fb1gT4UQ
8J2vBwPj647ff3cQj9MopyTwSgN81stkJN5kAUaXY3hNn03pMjnJzw7V09PiZXT7
gv+fSI8hfC3GvY/pd/qZ/fBpbpboMdQ+1TSSJh5uPt2+BSPLjRlmENg1Wnl0I/pq
dFr8lsXpI7x9+UcLvMoAy7rTyaDiqo4UuMjC5sy+ENYHz7Fy7c4AuhkAVWh/4fvM
2J0IVaOPF5bXPsVWsNbxm19YoPFZrBe9YeIMKbHuXv3f5oBJPqNH6OIAkjcW7TKk
5b2eHRlX1pgAVU+oM4OPxfydAdWFjruTbBuemDwdb/J0TBp9nnHSrmbk19ySoa+T
lJJDXQ0uN72tK/OO/9RipusL9kXAXKPGmfwmvLN90v+8Mz60F/ELyIlrZ1CcOjkj
gobiOKGDx5J1m4TPTmH5csOtSpie3AfRQbZHf1q6FR/Kh+zQEK6Gt57Jk2bbalCE
dBXYGDUsDzTXwiCAdTbkMGchSGS2e2aMlLJ5Tjgv2+vHLqgREtkYZh7/ZnN+6z9m
7QiidBGxx69LsC6VzjnJFSE6ZPmpTFwZBZwCMjc7ExRlbkc3hUIkSccFTYzpl9fE
Qf9xc1dTKpgxRp/zDQ0XpCWpOb1z8EGyxWbwtJGHlVMhgG/v3MOJzKs5NuxiPtj3
2f4+6SytAdnIi3hOBcgAszi2GUH+82nLEtHHUYcCp87U/Co+soviEI47pDUx+yOC
mfsYqbfQTgEayS9UQ6RJV+Ek1D+Cwf1N9he7aRBzrrCyEG6nXMSk1Dg1vclm5NPu
dFhtxmvQGOJo/968M8q9gtqEcywee0YyocU5bApMNip39Qo2UTeJ7nzL23WsZ8cE
p9ajBWWsNl6Z1tEAc27YnvjlpT2gYJ8DDML9u5q2CxgU+6grwjBwvQSRgKUv9TQL
fO7EtbgNXEvpQY89+L5g7Ox6FhSgvpOEATVK8Lnytbuer4yGt02beEMs+ahjpdPS
tapo0Guqii+fQobR3z5aNYQqqriQhoobtm8qcr2AoewAPb4yKjBx1FBY/s7YgYGS
iIHtOOmpp0/KjbEDPAeHjmv/mffhUyZaBAtOBuYcD21Rpk2mZ3BOFFjJlBh5UvCR
tCwCiwXvmsah4+rJD7SWvSQJuhWMlYDhbIqZjUWPb3j6PxO9sXBpBMJ5+7o3Rncy
1ii0OJ6viPCWzgy5sDok6oAqiOuAKu6ysZpfbx/P376sjNlUB26Q0+uWpXoKG7Nl
3W261Zpv/FePrXTTCmup06Zbsj3SryJY5tBwM+xDyCdC3/HyAfrGfM03m0MXwiSn
S411VyUKZ67pkOFtF7D5rNbSPvNRZQDjsLFYwwpyHGqxdJ0YK7L0NEqlqjlpVi1v
dCrkpGMti9oFm0IvtkHaV0OeFRwON/+PnU1Jz3IqV5YTW/1ofduEv4MCS6u08Oth
93ZDve4769U5WVQTcnlgq6Qq2xkN/5o6DmUAP89qQGtrb2dzDBbawkAZidyrjzW6
8Pd1uVp9O7ZfK/Kgl4d5VoN93Omy5wgM6Ezes9E3Kuv5YVTd1FmKUTOqid0q5Zu4
KnRSRoqK7ly+T4SpTYbuN8JbtSbWDdQzjemHMjAbTqJUkd6QFT5v3BNSnh+XeDLI
x1jdSHtdJiniG4253OWTAJ88gHx6tOgCms5oCJVHq5Gp+pcRl9vHWO/76aa8rLhG
J6zta7pg4qN6luE8+UnfDXAq6jtpOFVd4MpLUJa9Fw39gUkoOmFmjzHLvnsU6lgh
MRq0qs7fHEx3USn92WxbtfSaBxrnHvgecC/Ly5ZBftSB/05Mz4E4d+5xf+WiuIy9
RQ5qeSlEZd0CJIpJinV/1DnQLwdO0kk76GjfFaMntnlL5qo60M9xHXVvJpFK7dgL
f5MWP3AgkV24sjiaOkhdnrrYRGQMoud/8ZPC8PmXFR4DNZUljFyLCMBamkJyJ53q
73f6y1ZWnsUwMyApKSY5bGU/0Ft+o8vjqf5IiMr78+R1uAKc6MYDx6rgo5/sx5FD
//eWJkUbW0IUlgttDmkpjiSFhqVWX4Hlqn74nUuSBL5zNAC/rUFBfinY6nkB+RWv
hJHz5qNer5GTZ4+6uJkdJXR8eR28tasj5co79q/LWxrfjXWqXm4iHKa9/rpIEn8S
gXvhCJ6soXZI1zZ/FBfU9bYPmqcPJrzaDNollm5RfCxngC6rqtG9MlhMsN1eNK+n
nihgL8Y9Pv+lu6yFPn/CXz/OWe439WX7i7nKTQx70ReWCm9AoRL8dvWa/M7WQxBX
eMqstC2lhfmdW2lAba4g+kE9r5/Y1J5JCkb2VQ2Vp1QsqCbZ2l5ijAu1CIEPh8+R
w/7/X8VcFoa9C3IFqkrJF6qqVWqxen3X08OiwSr02X+lEyWZOL4KT/b7dY9NQNmF
Fi8GCxIhlx+djs3bCGD+h6tnl2qvQsY0CBjLYXgSAGYcy29HD0Q4EeC3rjlZVR9n
2/ckt3uKbf16x0jMlWeRAMU+xwHRz8SBKO4XryxSNJMKrBE3SMVcqeXJb6wvxugL
czRGGQc/+53nTaHpcFDua7iLx6Dqw/Qm6v+YHGpFET/MBSP6L2lpDbZInUOq9Dbi
/B2NqXzwm0P14hzek5uIQ/8aXGtWmSiUDF5XF+d0M8UQrtAsR6jLLvzmhFlAGEP7
vpqmKGSU+hTwuTF9iIxsgYj/ZH4k/mjfwk2Iqi1OfRr81BLmP2li5qXvUqiPDGPP
25I1ciAq02bybpDIMjti1vTp+tSz84gHH4TPNdbN+Vtr9DVYUb+UmOCYVBNjVYr9
AGBQx8xfHbplJK92ePq+3xV9Q8Z5/F48QyYK5YiesQStVyXQa75LcGqz5zZIWmnd
1QiLh67SoLKNpEyPB1+ePJUPA8iDWatzDMSr/aRbwvH/TRAh1H6QPp06vhPbe/qB
QF47jQGRJkjQQP+e90OLeZGRvKI/RbLAkevQpdnedcW/SmQolOziQdzs/8eSbySZ
aZXtaQDau1+E33MgDOqL1vAZnZ0capLYP2gQMcm+HZsRcxgICpxg9zjX5mNcHnY4
8I9HNgFjh2OI81EpeBAuy0v/I8F8ItJbwEtIDfrSiBAkQ3iHBQkwlx4DqvohnHjX
1KcZSPwer5UsXSL0vNURLMTeaojXzHpLllmj3Dm/SINAUdU8q4TQGoinXykR9Tuz
8LoMKknKgpbmz1SxmqdRSD2EMlrnAQHitWIiB4dGriOtw5LGmVomaUSOL7pKsrK7
WYeeS2LsYafFBdCkjBt0hCz+s093k2hFvgUlSX2raWjzJtzj6847rQsT/srxT0Gq
aZo8sKChSDyFCy0z0kuoG9vnoMsZjX/h/hUR7IU9laA5o5L+kJUNps3epCrdp6NY
ysnPSntBsssKN+bUIy+YlblWd4qtrqZF4zY0CL+ds2aTfdSSGKGIJGhRH16LMV6y
9L+CaKm/nlVyaxCuLAtiP5+YgClNMiBTT4lChBdoB4ImFH1zWwE2DsUJMWNQgtkY
ULNslRrg/8oPh9sJEQwS/xOQL2BnjwlD9LFT51O+rTrU4RMpLMg3i8OsV0wpno1i
Z2utCSFiA9N7QzWo+jDZnm1wGzJXlB6mMzQQxv7QXXwhIPCLPBQyidVpsbGhRp03
xJV3FcRPaRyjEfRKmlbNnoEislvkBapagcHojC9eVkTZfJejKpUjsClQy3QRrU8a
u+e8xoyYGTwXGnZum7iHP+aG+qffMZ1ALneimGJrxW9V8ZasAWR/nOyO0T/0SYAo
5/wtMTCtU4T/j23fpJLjUCk9fUEz0fFjgCAabxbcprSi+dUOH43MZ1Nw8ZW2NHiS
tPopmSpRyLWxgTzwa0DA7BtLg8zE+cfUJi85N4bp4KTIUiycqV/rKfDcUnqZ5rOg
ZfUSr6mea0N4+ka6Ms6VL5EuHizTAAfWynvbO9RxXY/GShWoRlJhpohtolVUu0Aq
CRl9TdjsKJPgyEtVuXpdoOOcnCAGrZ3rnjDlnZjPBs+fwFm8o9Y5hafw7GJep9/g
lqFmk6Gygq/fIgk+2zySlc7itAUC/9dFA57XYOoA2/gyluh2RljKxc6n5cONlIYG
SaTDfH4bylWaR0DPs7hJLgLjTXzOKLYQK0RaTEJzoQp7rhhahIsR5Aw4pqa9shuF
Wud+SCKpDZD7aMBjVBjNh0HloPqjYqBIMSXMGA8ggxJ4C7/+12gpR2/0+GeQLaG9
xzw9/Nq4mPxGEeScOje2CsWCABJwQFCzIahPdk4Cm5l12GBr4x/JskiSen+J9tlz
30yJJn9J1gnDvUwkA3tdpAnFdvhvPPzlO3o9omMoJVyiwoUo4uZFomXUx366IjrD
SkijIeTHSwH/oFaWAI1Wum3BzNS+gNxdH7il7JaLKHyWl0qYHoXtCN8llacwkEXa
EsFe9q//ZJdR0aXzGsAnz7Q1SOku3HCXCK22WdlBFNUUk2149kvsvQjy+HdwI+EJ
0fVDZMD0hN+7avVC7vptCqzRBWF1j5rtag+ZA5KP5fr3s8IcarKJX48Osu/fB5K1
Gu7SLUGMc1IvXWEuBtWKTGZ2kh5RGTf8nR/fMYfEOhbFKvkCq3ZGV+F44EWOnJJi
Rec34EHchTMOdWe/jCdXxW86IIsY56bSWzxaUb4oaeOEgyjm1o45PXUu5eNQ0U+1
xyMhgknTpktLfdNGpIbPE5Fsr3QYMB03YXzBJCjbflspMKm4WJ1C95c/2KzbUEar
aVOsalTMqYALYLgfvdjZ1SdZDSyeA4qOlhgQMHjaQ26IRrrax9xbheaSQZBELK/l
bwdbevS6uKx6fi/q1Hnop5+/44BpfrGNUEBs/fZikSgI6PIPAYBJKLEcm+v8e6+t
wEp993wtDRS0L1LeenEGvB4wt7yhzGThMRUjptyWc8hTT8ka2e/MN/U2vT44ztat
H7kCNKz1GV1fXVpMDD9IRXGtNUjwT66lFfx6fGVe9nWjdcm+h89EmifIKDRMxm0l
MeKBCRWMtzmEro0GPtBjFj3UxjyOqM8vChYt8/Y4DvR93S5ECih7+vywtwG+BdfA
FcPDbgEUYPEJGl3Kj5GGI7bn9L3HPI6ntDxYJk/yahexr5U7NuYWAIockMYz7uNT
SzotwExWa67/sMuicGH71nB/6vbJukGA20+gg0sAbABK07LAeQqzfHuPKaiBRBjH
7zEWh1QBS6d28pe194CIWRD9XRpV5pcfZRXXqi289b8r7nbxmnRqGTi0xg0Im+Li
VXX4VAmh8UoYWdbhTIMdGzUTAImCHrJvHARiKlHb5L0URdZijjNT0EovNWA8cVlU
nVtEJt6W2XwJoN9Gz1hzexeW71sJ+nLV8Cse+4rKq8kJPJoOdtYhP/Mm8+L9Pg/t
Kml+T5fNDvttJ1mpyZ1DFaarnZ1dKzpc153CyOY0FqIlCAbAxIftzQLB1bo1qosb
WzQQpUVy4+ayYBYnQaDHq83/MSoPujwIoNOiLIh2/UPdncsYczEGY5vQIWzg5x9b
Mvoo4gRjZwKV0pitn49hC6b2gqHlm/FcrU3r6ibTD/umt8er6mgZkepZIpYkHsTd
a5qdhO4q1eIPz9txHxVADSS+ECEvn8TGZSu+uyv677SrCabbDiJOBnSP4Nll8GQr
bneANh7KId+1ld09xrbL5zqb8aJhdoT3OvBrKjarrZs0wPt8jWt5pG/ZSZ18Dlc3
bHQJZrPQErxKtgYqUO9oOqIRiwAvS4yXIsU2E45ADqRjLVgAk0sSzggKvvcMsLIK
znWSLQd5yWJ4km1ifkTYhqjY8fI4I6XsTrerOzdjBoJho1vF6ZWZ1ZSkFk3r/ktM
nyg0aXqJIMxTCwfeROWBeKnXUiO40F3iKdI82eZS4QJnVGhSegxmYhzJ3G2niDqh
p2vtFG7CtsqfRe92ZwjEmaB2AGnCw9NjOKlD22K1WLWs0zWpmw6FH5MoHq0OhB50
dZfj+iUZwaJD60z4UYjWlNTAU0jCdDpkW+c963fgoXuZqny8hSQniL8LciIOXaiX
55jyufX6BVpcDVrVo0aEfF+hXBpzzpDZcRlTf8bjz3w5CTO2T4FVaufYYBB1JOLr
GKJkeZLmvDlf5rkeGYSk2UKp9GnoXQgNCdd+csw3S2zrvzscbh8Xx/WjrKkhLEXQ
GOyTXZ5dnXmYjvsVDaY8aJtH3DJfNIlqQG7/+zmrpaUHTsKZiT0bcewpqvQH1cfa
0sEGLGuwfzXGKb5N6aZj9Ond4Tq76GIktnp5XTNY7pHZPqfp0DJ5e3566nTiD8Pl
/Fnv2I6I1iOt2opXoNi726JNo/mAdA/nahUAOUEchymeVVc3uuu0V4NPMKw/jijm
E9K+TXrVJzq20tpcMIOe1PqK+HzZ5Y2JE3Q8i94CwD7kfYqXvxBCGbW8ydeeXPa4
UBurJpigmlURPh31KcUveVP1XJloi515sEL9E9b4nd+E7WGrY+eDtOC994g5SQGi
p+45aMppeRLPsFzJuTLTR0FmVfkwMG8Rl/V11meP3YWNbAyeMqxvQKZKsFrxtSCs
sdUyRtjdnwaIk+9afleL8v1FOyGgn1Y8Iv0RVBhsVSeQd+C1V3FP11OliBYbHjAu
vuo0OcZYOwW+KE4UooiVaiqRjWLEuBWEBFwoc7GPR1Blti9BcCmdxKdzjvlGSY+K
4VTslwVdGUbW5q3+1AzWsaf/UQxpOllP8+9bMFjE94uY3bGFi+bVN4kvQJI7Hra9
O3OQf08cAjrinFmk/xoL58K8Izg11aslnDOps8+Lnz7GrtsKYaJeQFGfQOno8X2F
eBmShiT75MSFVDC0/iUadpdzbEHUAvyG8Vsk4i1Q53S8ueUgm8iRLczMhpCF5jW5
U3xd3QT2YJyCgPbK+n6klm+6O19OvgG1pXY6m7BbQqK/tFTr4UVslNY5qWuoRR3e
ARU6Hz+q4G3kg+tnHkvv62t+XOUaxGyRyMA4+8CKAgt574jP8RKCt1F3XJbzBKAb
NgpHI5aN09qfuCiRrSnubipPu1M9IHpiKOnW6TNMDAQFggnUw/KTiLh3EB8IjqDu
eTirpi9+6vim2pPC0TJMb8d8u8msBklFraMi8z+Am7Lhm98j15x3rl6SXt5LubNh
RKBzx/lUWsI1oi9v27cTG/SyZPnnKoWcI7JUebTBl03bNTcspIwixG/4ei0w3+z3
diZjNPHXqAb70fVTDbWcfFhVFHD/D/YPbK1cbfOyDYjcOdY1zt+2UYE6MW7qgGCx
WfyDBFaLiao6a0jFiYkyD1TjJRNw/e77KKxHQ0uVd2qqkFrhDXzT13KuekxTS7OL
bps60NjnQMtUv2Hv7O7uH9Hks31ox17E9BQCbkZQXptkyBB9Z9n2zK5ez3yo8IMM
KyZKG9CVrNwEpQPp+Th0YVSTtXiPoRfRkQwwMv4Pq/L/8/8SgOgLV4Q1vd0FbUIs
YzrwQOVbF5PqYt4OpHVIvptOpfR4y1owh88JLUB6DHtvWC+HzvBhVrpo55jhbdVd
qbDw9wqmtPK6zy+c0dndhFQmySki8jXp3FLy8GEGpSBPzkEO1oOpqywfcIfHRqij
HxcqmrthwhHQ1c8t7Ol8n9duegE+7EaxNWuQvaXNZe9NwZMgWKK6Wv4pU3pqsiG/
1q6P6qvc40V2tCEjda1VwrK33CWNzeGpMM1rSuijLpsTaEwH+6eBKiIhwqBH2KuN
EhCC6+PD5GLc0jzJHzZotmNRYOVCK9GQQv92Daw6MJQu2R3L4mQZVGqRKOlHj7ut
oSXuBex/X1b90icuO65dKIa2h7dCOQHoRfhODvHnN5ZI1PLyJmr7Urx9X8VJkb75
qL7GIiXQmwFS+van6ejKAgIQx1Ns4qk2he1KfXsGLYdwliLUKaxEDVk6MT3Mgeez
vrY7H6yzit8GKxtbRMC+3je4GOv065/yrw0iD1JI7BEsdIip5fCaL5IoVjQVpyh1
K5l5JWKbRCtZ89gxbhvcg/S70vTmlC5lKXyjTPNmOK1FGjQRxy0NZs6z5MeaJ7HS
lQyjVuz1bz8YHFSZzTqiT5cjOw2nW9jWWKYlTLH2uY0J2EYbEwRckz+lc6oV4514
3tfu7YJqED4aXPd/czmaHoNcWInKFnx61pVz6G+ii1mC/cSBq1AJCncIzyKHUFiQ
8OYFvfq9uLoaF1F9ZU2gNIL2+HehzeXd32Kjs4DJchSFXPsDLLdn5ZoBSUxdAS/G
zrWUI1b9P//NIwZWSJy9Ckqw1VPccHTcHb5CvcXbCPXce4YW+DJK/IFwbfJgATHC
2+SLaJmPd7sCILIUXqZeR0UPgtYkVmHX2vVk8RMYYUY1XFLv+K/Kii+zPwn1yIR9
jYIBh3wZg8z0vl3V7+6Klwvo9hkG2TvGmBGqMYWKWXPGsR2AoqAxtCvDglQLfvY7
WR0X6QYulkChiqTpf3CkHp1smPaoSzvVqvFDSJNYRvkFVMqsLJraxfCJdMAqLK5j
LgqJ0tTKOil3krlA6oPArOWdijJXBrp6+NWDWhiCdHGwz3kVKpEJiBL4d6zeX8se
B7NguIdYQDl9pnsfPwx7c0qIpilKkHu24O9zgupJggCOJ7dwD/+cY+l6cODkMutV
LY+EcbKO7MknfLnHvY9iSNjvZjZQump+T1SHgC5fuPtxy19PFOKml/dLNlQp2wxI
sUpT6jTMxp7AdadwAEmnzXpJ2KqkNo9fZXqw2R0D3xiBavbFDxN9z2bVJ50ugTL7
CLLFpRditLlHZ+p+joGV20yEuN4rTDZKpLw03+FYPNUvHQZkdqSAgPVf2TZifgcH
cl+/YhqM/eeiSW22NL0+pHspIasF5MaE79cp7PWoI4i2cW18KzQDH4koeslxcjnA
afEqMko+tEJ/vvWA/xsRpHibjDhn4DukTRntKw3HCtF0GAfhCZKznHbA0ZMSyirY
6Zk2EMShQ4vncGNgt/Gsx2d2Z49ul9ivfSnIRK1IGLJckzZsvJY9PLoH16B9MmVk
HvQXTmDhOJ2v8InjDekd2utbUUhPUjyacEwo0JPOZNV5/LDTI4rZKrO9Mc+qDCb4
kqQPArm+GRJAfwmA7vCWX67RLfSWcsGUGWlxHTd6BJNB8SlTEeAEnd1XwZW7q+Wi
qn+2p1kXBA/76VVkYIZ50Sl1MB9rgGr/kfkTq8dK+Mu8FfEpa4H1QELjb855sn8C
Z0P9eHrcEZNh/REPF9+QCYz3fIs9T50xksYhvZMxOS61HILH2h+MUYlihXRxzNhz
iqfKwex8ezYHxtE8tOLnHywjJvAxljYMPrRQfBLxick9SwM19GjHfAK1n4KAkEVh
F0VSdD7//lG+i2woNqKXPBW4cHM3RJmSXyrWgNLbaSq88ORQiqglp6YA3ci1Isop
LccE13GbK9y/Ay+rD3FlxCGosvsrNUn82uEvdXeEqPWw7X2e2PQeFNH43oEVO2+2
LahZxUT+NhywE8zCEYz40qV6pljR75/+XmVyepZWe2Er1AZBmXVzOIINTOXmfEZb
CuoWF3epYgoskuc0SiVJliyKgJdY6uzMDk5/SiwT69zKRSxtog1avfO1bGX6kJ1a
h1pDYt40Q1bz9YnQujyH/Hfzjt/XcxP3voo8o/EHWKOMANMT8253AhXbSvO1SFIn
6g+uvWbyxm6TZzjxLztuHj8gme1tiWUQ6HJBQ4arzkQzbRgCtCO1wonwAKukmD8q
3Rn0WEIT5LXxNRWz0hWAhRANyEDpJbedUjAFQcDeS+/rd/MNcyLdnhcIzc7sXfG+
NMzbxKlHarhtpL16AwAcsAYL3AJChbawURbFvRlyIbF/WLeInDGFnI+5fzfCLFol
txFkhvevd/PJbO9xZA1LTk1NO7f/t+l1pVJ2w6XhnFqqy/8Q7Dqje19Ft8MTd8q5
gzuxDNiwSCb8+dfLmAUqEunCqEUHBYVzllfw2ZiOCPeeRJXaRN1UNo1naKHtfUA1
CuNVL1dDpxGh5LmOJao8+vXWYSRyDynjL2rf3OmK7+HeFFJI2RAjri/PtMkUhnjs
+FBiSQO5PVR4t9phfuRU2IkKqQTvOKJUyUVsFpRSprPou/OThnPAxHBLKTsgyPyO
zEmleusqN9Jh1uyw905iwsEjiqqcwJYs+XTuXorHe/wGEUQCxtg+Mp90AWdfq97l
XX9j2zV24Frts8qf8GG3Ow9RHvsLdhGytuFdIF5F1pMAGX/LBpSH4bsi0iiyxP9Z
zhyh+3AFP3s1ZUNvPnJYoHX9EoLb+DMFYvNkxZxWzW/gp7R8nfS47i3r1XaSiH1f
9ulaCVcgOPIhCqn5xB9CBHEGfs3PS+kGCQN8qFwTEFLh5inbyFqP0uELCfX8HHFQ
StsEzcvO4rmmqarIDbd4+Q19qk7wxwJ54ASi18JRpQf8PL4OAMtZVB4p+IqAl4XT
bHkx+7ZPkxcG6pX5IIeyHlc+36kXGTuBtZJTICpbE3+BVdVz0yVVsupvoIN1BP0L
ndnpEPFw/g8lHcrMnnX88Ywga4C9qqxnfvgPggSKS9GcOwpItYAYu58AQOyrVcA8
PzsRR4oCLx9vGi1VvKcjobUCY3TkkfAs+s7mu2/vXykxhKdVjcxF6+9Yjc0tf8+h
/cjL07YeeAYiljifmRAA1PCHxGvxzIjv69dgnHZkMCps7Q3+/D9Aob9/Q2ngP4Gm
kWpx0ikp7fAnKQ4G61Z8kKVncwREoH9wewc+3IGAQ2e93FmQLB9nOTr/5OdfYm2S
mkbKCQVT4QSCOEl3brqb69brToJp5Ryqh/Y38eDBDT4t7WL9kj5Tn/JHdx8hZeOU
nlkJ/Q75aJ6KIubDKwpg9IYiht7drp2WqLw52zGt/v8msdq+rGuxhCLH5fF3I8ZQ
q8CelWbAyBrKpJPaQxmOtG641K3mcu4OROwjF0O8Er/DzfR8OOOlnN6O+LbW3Fw6
xwlRwPeHWv+NC5qLkMtnB3qeTSItJxFwpysUGPGlWcT6GWLeY6ZZdFAvvmdg7Lw7
h/UICyzccVLcVc1EPmzeHGCokJhHYstQrHhzUiBf42Be7pmjQK+OhfvaJv4Bq31T
QKXHcE8a4BRAbZMxn1Fs2KQ33IjHb8aru+1py0/xD/OSj8V4apjlVIq+S/lu8MSi
sKAv7s7TUtoAmh8dzgebVjw7WHDGsMkDafmldSU4FCS2m4g2KTZ3+TJR18Yy5Mw2
2CqtaUuwG8e4IPphF00bMqfhdw3kd2gTO09UXR1ZrX3wRJCJBygWfxiO4GMTeLZX
zCbQpathsmrJEdn7/pHrMYIUrsVpl4Inty5nVMA1M7c8OiGNDEgKGsavfvWuB2cR
ujMgmv8x4lbLx/KgCci5AEMOYoUcg3rUtLwXxyCKndRYhw5upF/2x61nfzAiLhSp
DIFbnzSWIsakwnp+xPn9WzVVky5o7DXCMg4aA9Q/k7peyTD3FCsqrKQS+lPHaqRp
2lHRDSmAmYEiaLquNmDLUhT0K4QglOeVNJgnpVFRP9b3aDoOgwRMrEm6CbxC5/6E
Yb36jmmTX1PUCpsxtJj2gDpUnTVrC4vLd4ItB0Pt+TqPcYCXDY8+J5qVljQStoXC
ZqaeRraPQVRqEyQTp1acm9PVhfNWp1USCQAhYUmIlt1aObtvR+s+J2OiMDwgZDwX
L+SuvpRdpwW+u1MpfuJRWTqg1soZxbMXqul79akGkEQ1aYQPoM6+Z5xO1fQ3bhRl
K9M51dejSoqh+XOPwrfixXCuwtT0FfZo9OHk2FdxpuE66yY/eZ5rbXJudcz1BLVP
e+ZrROQLeri+9WEbwckzGzJzL1MEj23dvYhJNrX9hi470ShSfagStusDRVI+5W4e
00UXiGJr2RYFsjEjEfwMWVsjnrAn8tKByESNbkfjGhwctqr531tnpMWr5PWDzou/
Lav+ohcUB/dkT4ZZV9pdUBAzaQDg9YQ3To7dwHPtVI5c/KFo52Af/n2eot7qRMxA
nA3lSET98r5UixTSESGMwh8hCPVDFNFBa1Fs5NoCRYrGK7nO64fNJsiLIgC4U4q2
+BCUu1loogLlh/bI2pMx4imDq7NsZEYa+zU8kOxNGmK715OLUCw+BS+1u3cjCXgE
qtMFrFTYHywX6Dh23qI/jEMlozQprEuWl2AtfRh21TwB6xJGHjraP0dU2rw1FTS+
h7ZAh2FiZfezSIq9zioKNlCMmiBbuu9jnLUgwOC+/j6lZKaF8L4UNZOjCaliJrfH
MYCV0RnluR2dFwOyeWBTWBkaAJPCKbotnpF9SPWib1Fg1LeytkTDd+pBxzcyPtbK
vJtxY8+X+pqoE1l8kvW21CANzwcpk7MQQHFDckiHMxgjrdhYr4mVgSiUNM4vdYvi
1rxSWc87WWLqCkuEBm6B7QFyMPF/2qvYTtnm51TYrE6Ax5oB+Y9oR3RfLIrLCvMc
+I3fYk1SxPXCa+x1NPB41CnCN4g/wuUG+dJ8V8keG/n3PkGOVpMZqpT5lsDOUHxf
ukkYcmg+W2su+dAXbDYwXmLDzjsydxLM7a0u05Ag5Q0xYm1i+h6iN1rX8vmVzAon
gcqNlMQIz/YMKmweW3BC+5RW3O+hXTcP1I8JChf5r69NjsV0jVkUawBjoaDrFIkn
OyJZQM2T7UNsdYZHuK7PPE0niiQdeLVaziaah56+9Kx/+nTVdpTGJ1Y0udas4LvA
GC6cEcCsfAp54QI9fY9myfd24DNXeu1QeSKTfjWROWLTcrLqjTPTzyULyU803jup
CwIoxoEpLmsDpnzGtD+mVvb1FmTql9OPlKrphaU9UGiY/WQGK8NESNIh2I1qZjFe
fvEq/CGc07bLvUiR+5rGaYbn8HQug6ZrAHDcGxM39TB6/Lq/BkbVHNGDBFRFYlOi
6XJ+boVDjekVgTzGZv9lVn1ikm4PS32T6nC/PJczyhWfZ8QpVJRASJDmH3jyyLt5
PAhNi9RXWtstkZbYqtsW35piZXF3O83VSax7xSWjKQHw4suNKjPpqEv39y4q2s9m
iqlbOF3XRCKKOgwqF8ymG3M6S7LXu73rhV4r6IbCm0nQpoF8kB7im7EOuDDNKFDp
gCrYJnnjU0xX4VfRZN16mcNB9KLMlOyeweSJxMTrJc+qSdPqAW8eAPhJl/f6c5su
En4MpMJRPZLA1dR/ZlBWlCkuIPit2KGnff11jWH9vJXNH64Gts5IfGZQc/fWDLfD
rTojJ7c5t2OohefAhHbcFmssd0rP1apMoSqqWfg5AcaxuQ0yXqUPfNh0H4KBKtkR
J6AIBwTNU6PWwtOqyQLW2TZuejN9Ls4HucaieHTu4R3P3X56J6EYtcsXFU1mc1gB
DdjdkvJRyIuG5uztdYbuNpGnj1hVilJTgZAGbzR93jb3xNNWDSXl7QRVR+ZtKn8o
AdccADjsF7ummIUo8g9AN6KTSrL0FypWwd7bZjv9WBq48lAMMntencRr9qAJ1BAF
eM+Uf07l1p6FTlgKvyZg+Rp9AoftAbZ5UgnnFAWKacQe49tVlw4Em9PeuX3E1F0T
2yHqDTZELW7QwUfupuSKCJcozi8/v2ti8LfbDtFA7wkNofMeHlTs5VG/1ckF4Vxf
lki34F/uHuDf9aUy5u+B51C+idtZJ7Q/mXWiVohE+1vHjxsxuDpFHWrdPyxGOrNL
yN3X3uyIl9wZTwmeb1J6ql+6MrKW0lCd1GBIaPh10JVc7jYg/mKs30hGjgGlyRoZ
7I31zjH5Fma5zIaXFdj76zVb0QZ85z0rvoQWNMNmLfv1gGsMnpWXXRhMnWiaz9hQ
Rq90Bna1mL4q0WnFcWZlkGX6/CT47dwWCm8ulMvf48AU/dheUthV3ojfXrzaMrtU
Fj6ztPzhVPH6+CXLtF6Ir+xcl3bieQQEim9Ye1Rr+nYy2BVBCfDKTArUl5uk1XXH
ZLwcMilv3JtJ0PCvN0I4wL7ZndkPzxorzCBDD6LMgRphdPg/hwKPKe1dsJkY6x/1
5w94FdwO7Y/VxxcD78dXdzBicWrppQ7OXC2IsjtyK0GBDNz9oND3pi57axU5GDFg
yK2LFL+4o6EVS7lGSNcrpuZyeBW/pSa0RvHaI7qu48RHMXADT+vDCHOYrCvdlrfS
H6TWT4Sg1htJuwJpE30/ysgis6N4dgrBgNdFtUN2wDid5dmGlmvb4D6bJb88CZ7s
KilfiLfPk8jMr36Pbfs55UtMU26HItRQDp0X8xZ1PcAI5g/Xj+zgsTBkc7rcxdT9
IHNcorEfg2hzTFEvS+TGjnxXNi5fkSG6u59zRkmWLTpG2JmsRWzouQsgPpozExWv
42UHEZLHkRR9qS6NQ5879f010bdB0M+sOsibrbiyxLgJsv1S8XOKF3PtB89u3RRs
kUx/OuuaB9BK10MZ4sU1QuRrFfd4iyM6HiL5jisx/9QI72JBWFynz2XXKj4M3Im8
mgVwv0i1RUrUbGEuE+QwjfjU+zYG+4RpqO0xjv+GJ+88Ysvec3b2n0cG7ntEZ0tm
jCkVxc3Q4ZZJR1GLvDn/WYExweQH2vchaVUgx1jRr7KusT9S8QzQlD1coeIIdoMB
rMPF0xa3SJakBm+uW6dwntHptsad8rzcgLHlG2doDMza+Q/iiBTYUw+qlUPSgORo
cggl0abxNrI1zESgyIuQ8yfT+n/Ubi7/c3qZ9qHwTkU9S8isvAy0jbT0Fz1j/q/V
MZ3YITNjwz780Y5kAzCqIt3dXbmEHeSDQOQApYeVppVmkmOqnVHbzGYk2eRB5xW4
hoRg7fOTDijsAy05XNQwLTPFdh1Ut1uFfT6/359OQTgzPkzu9bbK69NGTK5O5eOS
PrOsETZhlZT7xV2yEHpMpPL2lv6AV9x2BtW5fK8Sxfb5evqiSPc1OjSBrNFYybAU
MterozNtMS+Gwa+jgIMQqsMNs0u0Ghfi5O87h9Bq7fhSGW4Tv5ZXzQyRzXodHiLT
ZpfAqeWwlZWJPkXNZtB5twTxQMmwgBeOemO+PTagBDKOh40h7DQJmlrKKpjMgkmT
DsqebMD1xm97EDZOk0MPQ+xq4dX4q4p9PwTEFCofiRqCBp5gJTqvpryCTH59k+h7
m16LEUxs/hoKjLSkQK2Db4zBsVUeOmPGjvOgIk7LYxNwbNYPck9uTKjwq0oye7hM
9UEArnjNUcBuyVV7MqkzOB97XO1GB9Wy1Tz42CtMPJ2spV3VK6FvN5EWpx07P8RL
CuseY0QbBHw5E1xvODkia0z7Fdy0gFn2jq8ZaFCiKulZqIkrEXH261BorPj8cVZu
Rplze7Qb0jgST56AtnA9MBiK+sZ3QeKYhyZRVXS+lNATVUCHxJwZXolQkiPO4gQc
IT9MZXsaj52zxJCMr68b9//hUj0F2f3rO9m+miZY7hPEKte8caSLaNUDepQHXP8V
rkSF0co37+Q22lNuVxKBLaQJnE6kKKzXWEPKK83mGQ14xGBAfReA1knmxJMWQeXp
IL8dDaenfInNsXTzC7gSBRMfC1tWogeoJSWvqlg68dWh11WPOcjgzS8Zb6NEI6JL
RE66HhDCrCeLxwwI+F6BcP7lsmsAYVEEp3BznVSwDC6Mz2CWm2pMcPGkxiNZ1iGs
BBWERnlSfx/qhZMKdv89GvZzGvxbiMTv674ejWh9YkEQvQSV8oo4vQvYQE/s6RUQ
M/HYc3GtY82+DBEC8nmX3Z9uOOTVm2j6YS0RVoMNkfOfGPPUQOEHn3rTCXHkh0nD
xrH6SUJGaJigqOl3mpJvqwiwKL4XRBeZzBgbXlhbYiQ7wezvAZBif40DTZ9LLLhX
rASaH8o4i25S4RTYez/2ZGyZ/vm/9J3Wl2yKMBeiCJ3lTWNFAO3xrWoadu1gHdyE
DXbggt9tbs2E8OWXpuNha6ViqLE2pmjnzbGSQyK5jBqS95g1EDOg3O5MPl9Ezey5
gQk8k6WJ9aMIzrP51osb39MnhQ0jNBs1xSjt2OcrKao0D5jbOmGL3jdWj0zn5hiB
18lzZE1Nko7ZVRA43yPWf25epBbDNpWPSDCtlScjPO4XFuy8wbfG//uG0JjToEW3
JPZZUO7GDwEyjwo+Hjyqo+ztwS08Oq4pHTWH8/u68y2Gt8uYTjNUdpdI7kmfC8eU
2QgzJaxNszw8jlg925Ex3LUVD1pWUfu+oQOzXu8QGfVrJPWR/x2r6tc2ABvypOyY
JQA+WWEuWXydUtGWlZi6i1cVuSEbysBtIwCwfgs6SbmitNRIzQFUIyAdqbPkzUEh
wjOwqkCCT/KauIJKpPDuWEmwEdFtU04tswrtZqqDhK1CEujLE2yU3nS0i8NYf3yA
nqt0FCpvkEpPYDNKV6fZ2R2B6TEKcZfSYsau7Z3O87f48XdYQi4GSdRTGmPdINLH
SbMpd/uvz+MTTe2xiH2EveYucO0kItYK5oxKCnwSfKoV+ZLv8asbMXMT2Chhaauw
tIi4qky6bB5y7lSJLMlhQUjVJvwx928skTQ286xFRYfB0PM0qKZ6rr0kF4xPlZSk
pd9rOfZgZUy3w9W/WIaNiFTlDMgBlg3zEM9Yi8Bdk0A70F7yH2ahPD7clwFLJsO6
EDkl8Dam+sKr7jDLTNU754iGwZa5ZFs3R/qDM+4RkXWAeEvGZygwY4Z2VPOktwrd
uDbovB4NnbXpDpM+9qkgJByGGc8Xc+IvgZuo4bQINYhOmACmnmTp0Wdg0xAIWnlL
PFYnqKiYgAj/OrsTtAwJ+aCcyslXw3nqMf0JsJZrYrI4nzzLFwf8WMnyI91dbdhM
vwNFlgEpU6xCSAPiaID/VWeTryEdDzEJngPZ7vG31CiILkY9ITLQt1mQ65v819WG
AfyeZg+D02Ufhp2orLaZlKXC/WBlvwu6pqKfc6UyceiCNjWzW9MkXd4zSYznm8Lw
TRPZQoA3Uuwnc4OLpPqtl1pbnDL5+MDolcKOgsWQO13RgtUFaUgqPYnn9Ecuw5Rp
eGIIojK3SHKEXzHQ3SsxGmv+3jgnDH4grvvc4SCUQO3+qN4iND6sbZgbJvXq4IG5
lszU/fbBiys9pBgVBkG5qd1jcUWhZ/jIBiIW61rrlhEV3c8jWPHXmgn0MlF8pAWB
ESO2pE30eTQZoalCgIN2bnX2n7AZfpKEoqu/GWFnvpLKyT7pNCe2l+NkPPUWKsGz
lneAcSulD6yMso0qHARTQ1X9Qhm1ET94yORKoKebjc6xNkLY0b0SE+tmmkFrDU+l
SvfTKO8ILwEUBkKubi+KbLJeIsXmEhlTHbRx8O5EX4whBWJ94tg6aEoK8LGwkZue
F948iD9vJRg4eetVbtQec4GY8/ekiih91HWIN17aOF7RjXM6LE8AMlz/bSozG4Ow
SNHyq0HzrDDBDm+Maw1YLItgBM7JErOeEWPopOygBl2I547Le68/hmHZvw+PR7FO
ouaIu01Df0HcO7OXzbtqwBPF/3ZMLPuGiF59+J4jw3wC3qhy/WW29S1ckvmZIbkd
1G2Q1gBuvcwIHgHE3Cy3VcaGknjgYXhatwxCuGM7SPLZOkoOkXZP2H7lMkDpFdRt
u4/GUw96o3unCNWHtRJpzhUI7+XpdSMEi7pDpxJRwJSJMjeOGPYGZJ/+lKyvCoU4
4qx3RCUAfRp4hJm0TFaF0cavksT2smAzdS2wVpfgapoOV/prHpgAUs9Fl28e7cXN
bNt6tI9m4n+UQMdol98PLUoh2PQopESn2WOzR1TJTw6vxRjhIRgu94/aTdGDc5Dl
aIs8w8VluBgY5VxOh322XkzrZviu9JHAfSNkqBY9Ky61NaYhPXPv1pZqRrZr2607
4AuynDPl7fLo34pwYitcn4apBeL+OMDX1jzIFq9/Rqyi6armN1PVQdDVcE8nv0lh
okK5Opmb55EJj0pdoiFmMjJPEupZGH+6SKLc14SmBn/mJwgthhtZ5iWeOXGJC0mr
9unPYRwzo97tqLI6R0ZFY8Fqr0cBsLZXqHsObqkgDPzMVU6QBKDhI/eO4WASWpsA
orz1I57l6mU83HjNyQVXTV1/mNHcclxNm+FM6Is7CYSslpmW1HIWAq5FIs6w2mcr
p9AU562XUlBijkIq77Ng5rd8hDZ8LnyuluerBJCgUwiYX5wpftURNvx4/SvzTGla
/f8bRPUpsHkuJabtThVH13zPBht4SGhYzEskNiC6hj9QJxij1twWm8UgJ6BUTg6P
Ej0+ZW5083IwFojDtOlK2z0WihpfniaEVt2D9h4GBoPDklYNYutH1XJcme35EzjP
0chrla3W8pb44NqLN8pPQTD1BhsWngANQ3JrM/ck3PH4stwT9XRkaBlBAB5VgEgr
plziRZnxwLV+8aCxlCWO3z/B37Q8/vstyHtxAF0Pqn4gaOafOz+K9WVXYAnK/BXm
ufDGqEeDpTNT7opGqGkKUGCf/5GJBsVx7Mvr42HTejMmrnXfFY57c3c9n9Xs7wNF
5akOMAZr74qfMnfSiVc7lVZupX+ADap9X4KfglD1yPdH0LMOx/m9VNvsEi/6qDCL
n5C3NSAhgFUnlc0J+6zpjw26wbL5X8CFij9inHRhYRYxSI6Rho2/ydOXRW9NJzpR
KD0o8EQpf1CJD8YgtRnuWGo/3ygsb7A27wr+biH8XFKPYWPhWdW48RqDaHE1cyNk
XstZ84fqSs0WLa0YDdg5ZhsYdtBwAGQkrXN8donlivM4cuvECnND9jVgpcfWBHSh
ekLThRqXSiSFmBwCm8bBskhTRnzw0ktY3tYJOB9lMXeZY79pmQl3QU0u70SqoxtD
LrEG5naph4UxfYsuiIBAvzIE0u4MVhuIG4vj1uva/k+jZ4dGRGRvfGACjz9JEQX3
HAQ+2GNoVYY0GDdHnNCqp0HU/EmfTDv3msepAfoqjTtuKUneXCQw0Teh2BVXgeuX
aZ2LGwL8ZWAqvYuZMh12X/fMJnIMkHq6VY8TnIQlSjdIOT30LmJVN+usweeVp7dw
s3f43RXMvqEipvdaQhx8Lf28gEskUrCH8x9sJ2HqIKRsTRBVOAKZRtY/azmxGK1L
LBWj/2Dfna2Vl3SX9L8GJ8UzXetXhwQOaYre/ChwtY3IRTbrval2+pDk4/4xnjmH
TVIu6T3FEXVSjtUNE3pNE69SwLJgbI1O+h9YWKh1BREqrnXeccgkr8l3v6fsjOTj
wYrq9JnMxF/ezyV/CYSmy88Xf+0Gf9wwVnkpx1vJsaH+hvU7gQZJIkEEPeNz4SgZ
Jr3yQKrOTHh/dm6VbeYLR5zRx8a/b4XS4QySSUxoFuU+Bmqaa3PKzIHHkq/kwjp5
zxJn7UPHxzzRCN7BQkxshHvoIP4XfWLXmv1zXztnTDuWPsDrD80oP14FzlsB2/6J
MFLNZFFuivtybzUlSSa0tUTnblhfm4qLqaKnQIgnOAOzGj9IIKjtjFHnvQ0xQi8L
5HB0nLJ5UljrrbOMBQV30NzleUtIfIbkjnwILURslVFN9yWrEV8C2Gy+nM0QRXq9
Hv05ahWwSYmbc4Eutsx3ny7bRRp/vQZ0mQXGcwdp39JhnHZzly+qKnrSXGuFG0IL
e0XgLD7UFqqFTc7hTmogzLvAPGAQeMDTCHF/9PYN7lK8+OpLROXJKRneg5A0oyIs
AR+gKG9Jr5DdOD/qRzMZ35zYZpIR46J5evvpBvXO6qk+WozkCj2fRAQBBi1l/+On
rTCgyAwLIeKJLHEHo2YS+f6dHCrKYQrDHdvi4tm7TeAqhypa9VjA0S2FAcdZT4tK
JLpnVY0KCWWH317mNebKD0uZ8kZ50vLGIMLkRkqcOHznAHGiKQT23dCJLcKYc6Ko
dx3gnc0cHvG3rTRq7CHKsydV9koCGDJ1USFNpVZRLh3m+W1VrNDjkX4+mNZS3A4C
+0yCQWVViEjG1HXm6dunDRi4Q41PbtY2keFtsKD0xaSsy0qm3z2KIisLwuDao812
rsZ7rkQ+RYqzsZvYqrWx6jmz/SOyIPNhJGwvk1X58dVUifuMYoJT35e+3ggYOsKC
PP7L5RoOEX9ADbv1CDU6QDLPEpxPP7EYXWJ+F2t22C4Bf8g8KLvqvLaeZLbZMTu2
hoWglvfFYPdWK9o2s3LuwAF0M7sc9GPhMceg2tjDtFOXHUQFzRfn31mzeRiIIKul
KqxjNsZS+MtV9j/HMZOLaZx7CTgKzrso0hWYBljB3jBzluBd7HT07ermAJEeM648
JnEgoQ19xebOk5Sna9y5ma0kULgbpKJqLM3GgHO2zgDTmQCy7lBL9h919Ra5Xljc
jsBjo/fE4h6DCvs/JuJE5sOFUZiKqqHDhLf9Qssmj9hv/P644tv7xuVI9nEmzQtO
S1ltfbu4uIvGT+965AYyJ8cVx5YAHNRNmanLTCPoXKEVmZdX4zr99LS+zltig1We
ygJ0nmfnwRFU+IRU/S6MELnvSV6tRRW+ZoeMpxQKvo4VSxEoeYTnlie30eBp8z+5
8e4lOdIziuS4nM7swToODgYzw3aFkfHCsc7UiueNVzTO+PmIU0dKXIXA+NjgPsuH
cHjxzX/hiTNaN1SGspRhi+e51dnLyyWJ6pzL+/scu7wWkO9iApOCzTuSw5441t7m
jAZ7l7vM2fJwTxt7hg0MiOrxHIJpmn1kSKfbj2Z8Lm6YFDmSPbzFKxyH9Iu3O7UB
cotlgFwAqjAW885TdsX2FaEbh+zKKL2Chn8AwZjv8x6JjgfymhKlOlYgm9QcccEy
vmGo0fwu33AGvEcBZNBsF3WscDDV45bHT5bhYMA16dckOHPJfh7lL7HMA6VRLxB1
kI5Lzl1zmNmlBcL22vERpohO97M9LtnxmG0Q/BjxlAePsGQUtl3vk6q9Hzq2mmEl
jGUyWSeW4uPXYOaMelJv8RFW96AWeIGEanUcbgb/PDjAYjywUuQs+c5fooUPiTmi
LfbGyIOXP03B64A2wqZ+LiRZv9NmkiQ6zi4J7PGLinGGEgXjHAjfFXYMkCKM7uzr
dTmFCjFtN1qFkJMWNfZGPsej1TfCHmRJMQhOXyKDq65424hLL/0T3BhS10K1P+oe
2HX/rxEbPESxLqGirPAdKhfsz3fXyi5Xf9FrfrhVk8tejS0mAbyNSXtQH2J+f1kM
xf9VyqmLrMnDx4+Xe2UA2tPGYgORpVCjTgBj4O+QC/4i9Mlc6dns9Q+Pv1dv0ANl
5/P2SScoNVog709N03UNiJAryVWikmiuOu8jDhhri1zhalpwiFIrQ02D4QZQRAGq
H04H2rHyKsXtaW7TBp2cVedik8IBZJxh5kNhPuIRK2+WhWM4rGU13VbCTrfNKZAc
vKrAe3w0uDO7XiU4aT0r25tVxJdcEyCr5yckA6bls1YHILc2R+rPZjwQQvwzT/jK
BQbd+kZetE65tMrQwwcCWmzqeraB9V4ksfw9yscTDphyqzFrfe7WJrDU49IFE37X
pQvxLyOBK9Mbt//cYPix1xNbJVQIV0IH6POSlYfugWXkdIMeMtnSHtS0CvuWM+xB
9uYyGz7fOyNenLZmUTV+0LD9JIYWoSeS/ymZLOcQYh6ILey+Bg22sdJbv7jDZqoC
7L4qma3LqxSro16qzcDWPsvTBG6bSzP9rTOF0v3joUXLHd0XH3FjqdoLjTBtdVHG
SaMtDMtlZ3MVg53tg0/iT6NhWnwFzzIN7SJ3tsx+iqsFOWRkSa/iK5DhlSksMzWt
qbzjbdSvDN5F+qJxuT6ntjTCSlxxaIti3VK9T/LXt7L7/fBq9RLBVyWxKW90lXey
Vtx8U+SR/DqqVPybGSJg1ntivWKNXBt5F3RWDsNhG0+kid3jaB1utXmNDYtfRTm7
lFcoZ7goD2qVDh7kYmODOMNDbbTGtNTFchwPHkK0CBz6CAtSiY9V44FP5WFby8SX
DufehBronx2Bz8dD8t6njkRa6YWZ92ZTQQKsn4psjGi+hZPrzGjnvhEtEGZ8Zfxn
BVdFgROsTGknOKQ23XXc2GH1hMGPaVtLwGmX3polfOevwCNQAyEnrWNYtblsN3rp
DpRhijYdrkrKTtVmqYDp8MaBMOSL7ljAhl3SehuBFSM0QFllvAdDaGW6q5tpLPvY
VLOZarnrjhpd622lrd3T8mCG6ot24cHQ6dWvBmNlxLpr7VppZu5ZIg6jFnwAy/vy
8WdGCvat47oF8dxs7vrHK/elynh9x//iNiqtSUcSWDKzLySIVZ+jBOSOkes9WZLx
KNw/0or6n399slrGYtTxulu3uWHK5HwljfmzPLHfLZN/d1iuha1gn5JsJVqHVkGv
xpgT9YHM2iQX8K8LOi/BPA3aSOqT6L0MlPOgKqBeXM2sAjTnlBGJXxmU43fdxi4G
a58pcqmBOP/3DrfTkdm1upoSzT7C/U0paTJftB8+JOsNycU+7G1anIk4GHIdZr5Q
BdM/mheRXZYSZnKW6NoX3Z0qO0RBhgJSSJursl3+HaeBZjeGFAl66Qnunma0vKsW
WSEiB0keX8knVZmeLP49pZVfSJdEa2y5WV5EhAZUt5hgOZ0b9Q7aZ9UJ4lMKnGCL
dx3bOUDUmB2aO1IjM2S6p4Sh1TnvXHwovKpBEq95682r88vX5kHvxkotaDR1Mafd
ENScwhyCkCby7z+Klrgy+GbUUfOAlChW6FTE7EFfzw/CiegyVeMlU1ox+o3rFoSl
3UG68J5WrGyDKa9MsJS5nUEUT7fzG1oLEnIqtCBS+5u8K1lXXOszldgV6EFx2P1p
yzU1f+Z6JwHdwBnI98qu7Jao0rLs15/Ymd3gFgSKMP5ica5l5WFhtDqic0KrXWAi
oQEVRjJemcyziPAXBjJofdQVzgp7g0jjAIMgTy85541Y5pRDWZZYrEY7puOoLNgZ
J4X9/FIjYzbQnPjxPSO4+1GpFlHVyg6+Ts9mQwgvuRR/BxMkEZYwd7WtYqxruEiQ
/+R3tD0eaLBuzjjiS5OPc5lAAMB+cT6GakmGAMuoJaexJ0d8dQmy9pg/rYbXEK3j
hIEWtvLlOAdRA6ck5MWArIEszsscRpUBNbr0gr65PmDLw7x7iS8nJ4P+GsJQS0It
Dbpx7N4eq5WOlZtofpCU34SalplS99f76m7fK6rVWTrIYK6TJfhU+STC6xCOGXYb
pYBgTgm2T3Mb7iPDv6ZNeyVBBnlJcSqnZ2wUyeHf7KF/5S50MAsLuQPkASi/Xadb
/4wi1UcDY2xRomM6eXyg1X0subhUER1ebUmkLgGcd8CzVo1/j4DzRcoKjNICVUsm
N0miijR4vogdhtlCwgiHhPVhDRmxXSbwJE9PvM1mKuTSu8WAuNbCBc+XFU+mbGHp
j/B+OunatGxJT1STgFwQQwArp8+0Axz70wuZsNaG4ChxacksJcpWspxjwWDr58KY
xZlN5oEqYn+FucYnDzO7yHPpPUxZ8a53OgnhS8/PXET2nJtamVD5rtfli138FI2m
cWCanIgUO5a9uYuMmgEDQVmLI+KFZuY6PWUgZj/ZJ+zkB3L9FBAMzNs7wUBjuF7h
muVshI6sWMWx2k3xFXK3Oo9GpBvtSUHpQfmINBksLw6DnNCJPSOAq9fY3aERfzNV
9KNp5919DXDApC2jINefAi8hQvO6OQupgVO6ILLTMDyRFKsKchbwSJZN+Yh0OP2X
vi/tprYQ3JEQXFFZH08VpQ3M6fwOgcBPyNKvTbq2PbvxfyZqNmqTZ+CdnB+EUyu7
5jfw6KyyMQfSsggcazNoxB0LjC24mTRu2Fk4bGUDMxiidfxA67ewB+e5ejw8+xLr
tizuK9BuBEmATTg89pVWutALyGzDvn9GaleM6GHGP4mmNAdOXUyYUiYy7vN5UMm4
Ig+498pJrIZle82mZZexgtGW54n7JrL2u1mMO0jWqtTCPqFWss/DDdRq8b078AbY
dribaxSr/3ncsNOK6iMtucYiN3wDUcWtNxbL1/gufCJ5YNRLfla7gmnsaZe/qi8W
dguHzKhZoLcKcwgSIsVZZZ9kcTwI3QqRTMXh2bdnY6fWN78kHvgrfpbTEVTwBEf1
3MdL1e1aGwhKOr1ODyYR4bGIT0JQa8abeGZvulHOsL+kEGKTOHjFiNDupNahTnbX
tcpn4s4UZ5QSP7Ksc3I3iKb9E5QbCOnN1Ws1YNGuTbSK7RPafDgbh81pbNKbhBAa
J0RbHwy7hiUGoZJjcrWbE3C042ytdhU3wdcIfzXFEplF0ZOXhatsBjRMaNZw9DJY
Y0fYytam9IZw3RXoibarLEEP8vCDPOBzs7JLcC1CTgwxRTxQ626lG2MfhZ1w9OM3
EI7ZRYj52yIS9CKLuhPzHDURztDwett+45A4IDS1B7JU6G95nARlPqRhgU1HV+TW
c2YJVgYg+/fOITB2p6fr9NOjk9jV2Sx/hs+JkRb+RG269EUuAamQFexz6kbNHuSU
DxZS/OoBuEqUflmEsbypcUgnxiw+cPdzRW1SSwwjx1l58w6UiRHuZJJAfjJYxfeZ
Dip9/5SAnGp8KlQbtBFzpzYz2oseX9VCUrKd+GzxvxLiSgW8gTgHoYo/y3KLm9AJ
GzPklndt32+Auz9iqtXcpiwrQMSqdavK+h5tQvavGUOMRVDLC7FMXJpmNTp27QcU
Ns09qWzPyiSZSKk9jDaqYp4qKZq3wO4unVhqYl7B5yAY3rt3gMhsaCAp1FsYkfJ/
rPvS5+0dZ4P/8IrkNWKGS/iqYErSHf++IDk12TV43GWasLMjhWbdaLTcKLmX3G9/
ohO7DZk/Kz9J71N+voz1VbCc35z/ohdgFxOVYQSLxaMvUOzidINES5y8/vVo4bjL
dEnTBBgi4nr/CH5U5vXg/OFAz/XONGbdAfnVS23zwSmY/8a6frESmYQaeJEHCbAn
wN/PHtaIQU7493lgJgYuufbTPrXGkSaAk2MTO3s2cL3TAKUyY0XZKTz2m4PE3vW4
gTvUgOsNqTO8NfORLOy0ASyUFw4avaWH5V18igbKKWo2qaHWspGRxuT/gQI8qm1B
RfBi3moCYSAXmcJLYLBDqE67O8JWWtNmxRd5mkMiksqDPVUd3vLLYlggvj8Xzuqp
2BdNYb0U5QAmGN565HyQq28g5oOmGPO45SyEPKjpR4BRxXFBBbYjRAQk+cQlAYVI
fvQohmLLC/z7004Ch+gtV+nZxMdts5vHUlxny7jRNFsLZNjhmiqNM2rsk+t56Ki0
ZesbHpif6dr35Lm0ZcsV8pgJKKENQ00XDjYKe6t7EoY9W9cUVAFcKugEIFLok36a
iXwaCTEnWYtWDZQ2hqy+PEsPQaHKi+TfzgEnRG03zZH1TsOvgFX0jH9KsyK66wjG
J3eiAEckNTWbwc8jmJcOFHX7Yl0KtsjdFWPCMdQ7krfHF8S5/A0z+Jhdvi/aj+4Y
Wuo6DnH+4ZUQxg0EUqLqUMADeBy/es/D86K74m41mWd4GKINMJwPP0kQWuuHJT7W
UXqRZTDHSdxbir1/EjrUuDqV/cgzeVd6z4kSeoUo/jo7Te55LEPeOovA0u5xyZ5b
ggbXl2gffgwJZIBnJS8LmTB0kaX7MYDvAsT6E3qkQ2oFVqnUuUkQK+XqiRypiqVt
br/zgzI5gdlXlQTTxcmOo/SKugGZLXDg/Py8qp1PkE+JMvQJUm8ElGbLkb+mTwHh
Zpa1EiPBHjWaN+g4Lf2iWZ2HvyuTbLNm/oPF6IGEFf5LakKsbSoGCygA6plQnMej
Q0Hj0uJ9hDWLIJ9k+Wm9zJVaAjF8zsBQTp2iogLMuDbOGzU9kiA98I+M94zNAzfo
3R7zkN86DrIzn7lH/WsIvPwAS4oJhBt1d691SQIYUD0jRzbHgVsxvnB3q3kBlSLS
PnS6185Bh+0rajMAWNiLvYzaBy5Vq6XFlfzJzMzXfdrw2QB7vAp9T5iCxZcHZV/E
YFRVDM+jHLc8ulQG+DDWqSoZSnUJB+j7UH3iQ+YJ6Xtwp7YNfcgz+4yhA3wccSwc
UpMfBf50wYdHpNtDVsDr8XHGnatqim6dnoqzLepUdp7soLdvWjEskIobtln/9sLE
Aoo59lt6u4mkqKoKYp3jo4FAI7hbsYrSHomPzEDk6O1VnkqnoAkr118QYB9MIhG5
Fi7GXir08DA4Ig2gKyb5vCCQE7SF0fUUN+xiJyHcWCXfr6j5bzAnTQD1Dk7eHFWr
WrU4q4C0CRJVMrex7v9LU2I2d+yd/0cJpl32zyEAViqy+xrqcN2DPze6WEde56An
eb727apmJSX/FrMg0Ss0jsHWUSwuQXK/dtEQWxoYPNFqu06C5qKv2D69k6cKXUuf
wItIOJE57tFLU++HsNVMzbPj5X1W5FcMFuiD28dKJzbtiHKKX83v1wqL4MQbzHIc
Tddz5OzQIp3Bctc1Oo1/r1dDsgJ8hE+M2mRpncdG27cbFzlkmKRbPfLRxjIqqEKj
yhARp++CIBEillWWu7E2RcN9Jvo80/8xTdCf+3vTJfK4QaXD6DtYBAUGgbAetIxi
VxHFe7IbAiygARTjqdDMUKx6dKoVvpDtQ5+83kpd5dCgsJ7SqXspePy1sdi9+/Ff
Ko+lR4YvLPY1k2nm2M1B38pd79t5vM8qCttTmdVoNgvMHiReRb5Z9jar1CguCWze
BQTmRCCdviuICd61oHtvOcS1FvpwmJrWAcOtiW9Y1Dli1APeM8dHdzv1L1E6TEej
n6z3G9GMLAlEui3LQBL227I4fOMRDM3iTM6Tq4xPo7AQ5aOMYIGKcelfsXg+BgG1
+4cwan15KFg9jutummmff3Xm7SuuY9AB7wODO1yaByeIM+pO1nMe5L6EgwgiDhgE
tYtFhYI2lOsaArg1lZN/yO3NezRPR0fQthVwUlbZZksG0/Uve6AXvwEkG55z1kjx
pxNST0UDx7G2T7YpHvtZ9GNIN6UFVbEOs1dKmG/m7tE3wbfOWvGA6ZwqejOrmcQ4
AfM13z0hh4DX0AWZZmMR6Sr6KWxzd+LHhgZjBMYZuzgZZB6Yf7AE9eR41nRkUrNv
4uc8iVjKiS8kktupYl2JFwP1RfVIBzMiuxqilk7KxVkvBeZlTI5zbUcz0ekrBOyE
/hHLTf/SLcb0E+7ifkRtxAthhT4E1DKCccWIG8oLlUQuW5IYFqQcVFVVhQzMf8YR
3LLNivyW6oQl+DhsbPcHr2ut0KxAJrwO0rOuNc9XBYgzS2mzkfhVwA/0MSrsROYq
QtjzV0m1+ddsaQqYAfLR/Rc0Wf6AOFUEdnWMo9F3uc9tNUMk6M1vzc2W2wukHCAW
6O6mXDrMtRm3Bjgy2YGXUSkaAS+/Y6whpSfj722OoGT/7g/uuStkAn13cTQb+T77
vDDmGPHiT1vj/4KxNMoz0m41oe8i2cVnwcJoQtrbwTWdvq7TFLY6t2tl2TNnErTB
g7K3Gy8lbXxyYxjlyoWxtjzrT1AkLQ3uXckezBA1Kv3FrDm92tOSTuTS9MX1buBN
Kft+96+Sdfz9UW4nzdYgYPs762BltJkPy/2aMyThRZqwTj0l3WR3+wepAopUi30v
NZylfdqaKyaH6+VH/0+8KtTigSaQLXRQ8irQUH8jX+JFLNYu9Amvl3fFUxmD3cfM
p3yUSwmUrYRrR88b0KL+/WmmWD34me8O/XGHWI8v/k7qqGSwClCKnWJ7+YSn6T9k
J1Fu8vtNiGii4Pj+U3cmC1Adz0phW1oaOn9D3v7H4sNnB/71sY3vgxTSeSfnUNyG
36eDqSW3GrXhkvTpz59eU8FXWepktgDfbYVZGvi3OCb98p7bV3xLWlIOSkhRNwee
/K/LmhSzcKD/cT9e/8hWVbc8gG1Nk2N8hn6rZDwMzCQDjqKpHWIJ5DqNwCLCYDAN
ZuYNLM3XC1c7l0uQYXNiWzQOMRuX0qTLt3AYTyqSHHlxPiQxTQ+NKUM5+mN4QSsi
Nz6rtuel4clVWJFCkxDf3Mt8robY562m4mimBYCLhA57KlpH3BbAaMPD1RQRi7ku
DMrTNYXfBN+5QKL9VCCms2AjwzrJHOWbJsdIo9XvbFSYkzMf+45+xf9iwv+iZxsR
GOtY/WK0A9httDFYY4OhPUF0p7kpOE1bI4/Fb9390cvU0SUF0IGDb7uMdXR9tlja
e6alP3WAcx4ksDHfx2bxIbuOqcLPRBpf+H2LEDn1VmpB/1pn/eCqjXpBvLEur5Cb
N1kP9wywH7rVIDG3KWdEjolJ12YiYpHFLAQf5I1jUcEVXHUga5z2kfeYj2wTyNji
trNjMN6WPgMMUHoY7ViMTGu5O65n6EUagbGcWwHtDzzFqhy2flIeMdpItHDn6dIz
PQgm4K3PBuz+Kxy47Nr0EBYEwb+hLoW8k8dt69Ke7CeZwLPW6jd4Yam3EGQ2I78G
sgykl93bWxAdhbnl4L96GEmbJEITlUqfQjADqWdTPmtX31rXCFLx4hPthp7GVj9r
jk6Oh952SXGGp7NhEzEf+sRWhphsgvqtPrU+U4nkrxfCyLhAdzNntT53o/OCx8lb
R+StN0AwZpRPi4/vNeEb4dRlI7H9F9hBZrHbtTICJY2Lda+s/g5YLxXG3AUELlvh
6+6vEwH2iF4JAdlgP5Gd/MMWoM85+bTregEXL4NsASQXw1qPsbQPbfSo8ncRbaht
ZFuOQhuilxyY6or3R9dusvHBNFkXIFjRaZm+ub0xhPXR1DjgJF6bg/0GAZntG1p7
HQHK6HblU7asMCV0eD/OJPhSlI0rnEhvHhfBX9H/nwvPvgY5EqJej9tHYTqndnCs
h1ukSZLcgyRP9ZT7PHTrWygWD5DJGnJGq0yrWS6fGuPNDcwkR8dBpPmhXb6Py+8h
QpRebptW5zBUmWsw28RzGWws+JOXje+UCcBi1grSL7+DThmFSCClV25zWP0TJ/20
pbvLQXSJVVsvIztZ4l8S+zj95tEkhP5bieokPZ/F4yySZLoejcWMslpp41J8gDPK
FM0FaFLYVMcjIGOydLk9ZOjASf2oMi5o1BQHoYVxGiYfQSFjzwKZmzdBSlijMxUG
Vh5utDqc7fEmRWIN3nhAveoR4cdtAWtc2HzCHzMGqh9WSJ57zoqOmwaraffcv+Xm
lpjtpinBO0i8cfNmA1giE+sLhW8jwCIC10na/1YPEkil3gtAR/N1NMTh0B1bUFfD
phXBmo0x9VFRT6fhayIN21cwPzzsp3oq7QhJmyvE1bKGC4n5dcf05m8w9YzJpPU1
HYMG8gscaFJozf+f2Wmcr8ReywhQV2LXcYtSewTE71bZeeeQaibb9ZAPSNh644jU
9wtAJ1iAg14wvBOhDxvfqb+vskSICtZ/lTITuiGVjcteGhJCNpPLMzwL+Da9bLlj
Uz7imaBtEcA1tyLGs1GU9nQ/sXMb19a+sbGL6qrGjEPpUt8RSPGO2RV8qY547NEF
CV3sQ25AeCN2KH+XjX6fLStC5c9e/pC1V7ZzI164LpzgZyDiI6ZQsdHX6slCZODl
52yne2PFZbHqvya1wWRLI0L4AEcpnQ8QefLf5iSOgNYhEfmKjcvHMNXUy7u+jGYi
iaS3QcR8Vztm6iLASDmdlfgMlCe05ju0vbOd2LieIpHB1lm0mNoD8FiKjBy6Ujg6
mOvMYN+1ch8mLppav1QOP4avSYwvsDsMoIbRqGuKK5f1o+bb8D8T0Xaf7t3HQsJo
KZxnsgeoSaLuSl1cGK8rAcM5fWYT4ph3mFedyeJvgmRjLjZDAueh+iaQ+Taxrvuy
LsiO8BESK81UBgm92542Qs0pZ/XKDK3LgFh+lwMghb+R9ax0a8mkWAq/jf/GFWdM
wiIbFnKi2yy9PCTrONemBN5Oo2VDTyArmNQxiUinSXQuXfZ26MnthCu/odKFiU/s
kvbxx4C10BbZpBVlbHgg1PkupdJ2YWSECGJciY4ViSGRfbmyPT6op7z3MA/sbJxZ
fFZsLOz+cdMZgYybUmCvd/AVhEMUZmGr4rIiqVovWOQ92SHJWNjADddCCuPyY/6Q
G6f8IsAhVHwyKF1id6PdUhcw4kUQsAUADygDr88lt9zNTrsOnWqkivRpREqDatoG
JwG9eHa2yalH1j+1o4qllvnf2MMuNtzwA461xn8G/htWssg4p28jzp7twMJnmn/d
KlJz+/9VtK1M9JfiinUpfpHqEqJNOg8pETlq+sahvMX4x6I3ye1DRYTCumxNm70h
6GfxLtp4kGmMYAYch2n7B+KRpD3ZNfNpO5Yeo0cjlw07Cd8Vcer7IrnNWqs9h2Y7
aBH094MWYrv4MKOIdcv1HWK0oUN5OPLuLh0A3prRMbvp1/EN2p7kCRJOUYdTo8CV
2zABP7UEmwbGTh8iR/W/R0Me/4YxFP1Qmh65wzLvOMuzUY/J87R0kJFlcjw60qAY
31Atsy1u3OKGK1OS27MO9hQ0D8+OgvQcekSAX/kbE3SrsCSAfickzbIyi4PGCeBr
5QMK5B4cGq6S/6//bz/3VYeiHLcaeaxc6koKLuLOhwY+3ZpbM7JQrb7CiMLWhycr
Gv/d3F9zLB1v1Le1liy06KJu8qWkt/MlZEMfIMbTpyuQSR5SmKYKYtQhJj3+kmtA
YXik1CHW0ydDuZ2gJt8Ht4Byo9AuD/X0eqAMyfp/aYQTNc+ReOVINEJrariDORSV
/aKGoiHsXL7WKGgdR9X+FmqA9n9bD7exreNINr/s4UCi8WTyNKWKTq6xoh5qkAie
R0P3yRjq8Z3w7+gz7X6BtdF4iDF/HSvwuNlAB5ywXCsuLBcsqcYJMQ2pHpRHzBbS
+uiYszb3JyGPgUCOaOh+WE1d0w9u8StIe/kzXTtvMJ4a2dFiEIYaVt91TEqCKM9H
eTRVJpwZzNfhiSJ1xOqtagZzMe0/eFamJWfvZTw+5TDFEuks5UPSAs/eyC+Qb5Zy
hgdJzevyu2pgKAysfK0i2JI+pvUUfl7loy65wFCspwgnrjXlt8VZv0vUn2vcQ3IQ
mgstKfXWPWcye6A0aIBWXCk9LY9gZYqWLbrlZoS3Ky2Z71b1tVpCtfMk2UETLUcp
tsyO+GN7EdSMwwWOp0nDCvAX+ZMkmGCTHiTLNHzpHSiiXmwFHfMoXCD4l6tDuoPb
3RVXKfjMlozNiSP/2I8kil3qu6aqviYAagaJ3EHftvNO0XCaVou04e9BkjxAZLaG
4bgbfgrS6JUYkBbKJwoteWkMZcbVRtfGV/N8IyRzZnmvgDplI+EDbzFIGgS0RQ+P
VtqJhTmFraV8FbQf6XquJD3s+mDedBK8DTAyPQnwip1ZNcq10JnSo1uL/WItv6vs
c1+x5RFb2wzUkw53ZKGzyXFxReCIojfww4Pl0AJR+q7glzs6S3RmKACxfYUl7jG+
164FoYbUEW2vDuK1ZOh/u2IV2NeDFG2E/OVVFtg6p9GEg/bdUvKDqlrJvDyZ5txn
8a1T3CCesKUIsJsW6Ashvh1HpNM0eFOsI/Zhg5QfnyMnT+y+Ze0hM8B4czOhAyjC
KvZb5u/sFPf7ll2Olhcm09PggH/4e+x37nRi/shRQi96/ICeQjE1N7Jwnj4Ah7fW
1rFdhzyjBaEvp/iCtYj651z+YQCvWiQtEKScSq4S3L1hsXs9bytnc1+WpMOWcj8J
Q3Cq9lVFzrHaivn1+YIJKaZ9JEnLAvHaXsdhFhya8NS/B5t46Xp6MYWPVOZsi/rg
cX0VPfp342QfhVsk73KDZxDXoieDjMDPY+Rvl7xBHbWmniLOnLG2mB+5u1NX6Cst
mePGSDhxUj/PdlRmL08Sh6tMHAjB5M9+kYGttkD1H7Xh11HuT0t8sKn0LMq/hIEN
2CxbvyY8PXJoW+UNlIB1doXtp9KDveFLyjqgloor6IflvT5xVxoAps1iDKvn8Xjv
43v/Ig/ZTgBdxcPQDXYQygopaVcWpJZqrGgCrB7o9JGZyV4Wj4MofMBmpiEPTvJ3
kMKYryvSMFpRKfvXtQ/D9a3nlTHAJmEhATyhGQNEusXYAc2XUZCiyPHXjdIOf5NO
fDxoA928Xtrl1OJWTT6nJKHIF7P5OERjuUVkO7FrtbAZGUwi8kJ7IC40qJ6EsNsv
72dydz7vz+Z04Xct3cawnaYaytweU5cnVJG1VuPAYGKbN8ZZKplBmJPA87T5YBYL
oNqUKWBmIkQWu02UgR5Wi6T5UqM66aWkbCKvDEkai4cDO+6kPep1R2kDzoNhVxxS
+3mpegdoKmw0MdZr1PUo9eSMt6fWXhXRadPVuWE+W7aY6okNLQdKWPkzP2gVvUbQ
mY6HCx6lzCqt66WvpUl2CMofimyev838gDYbevzN2TWv1eF49sjdoEyrYPZ8q4tN
VW1iWuwUMdQwbNyc0ycwnJ456SMZE5CRPzY1QX/5OkiwJNGbc3ki+08PCzO50bK8
WN6t8HO4odB+wn8QTy5SN4L1NcCsg69RQleesTBhs0WZ4qOYPPy2cbEl5ky2ecb3
QMH4WxKa9LmJCiJH9pW7xh2X2pZxEKbjk1rpr6trKLX8iIAxJx/3pWHA24Z0E5Sm
xtAa5c+ki5KkTlKYUR35N9/n1eLmqhmwVQASuCi3nVsZ3xRvCm0GJ4UbsPy4zk+O
5Fa/2lG/jlxHIHU2583nyB+pg8mUd38jCRy+6PM4MieGB+qjOV4F7431KC5Zcvlr
0GnAadOwwanlCjNyP1aQhh94GSduWgMMpju1O9dCuYCodve4WTcufTLZ0pVCa/md
yHh8kevs4UYMptGHrGCoNJN4WghjAQGvbvsw13ls/V6fIDuu77AcxltNLghKH0kd
8yQFdZSDHfa45nSeSDhl6wvHqWPiu4MrjxCDq/biEUNNQo2EWdpzDGJnG70XnDgq
meVVlytJ5IknopFIp+VCwkI7L6Q6vWPk3caajIXsRLLnQOWVFMOnn+6a45tzoSZG
IY0qWXjxr/AxJIDRuh66mxMwBPlJNvl2UMCN8KNQDe6rSczsCS/BtKCFs5m4G27w
ca3An7g5zpsiJ0jTQ4wgAnwyi30clEyZ7Zp4BDkxtpfHS0/EC8sONZHxGXFbp624
ZFne9sOem1bEib8bS/vhknzCpFW28EZNWgmAeE0eaGavUptdP7HeEl09PWw0OZ+x
KuD6KCTSkSAeSEqPT2C/T2eNg5lUkMdzB3blrhU6+BAC5XDFCzIwmAqeb7KBhgHu
9GyWAsdC1Mk119AI9nrNoXpEOYKI5w8MgipyuQy50BVen7TGHiikjz8rnBUdL3Wx
HWvQ+Iq9/Vw5wYbAkUxGnhNl3Hx1OtCfHhZMhORiNcDui6RYcDgSI6gnLtEx56qF
LhvY71Lk2//gIyOT/23/c8tWECQvlec6xrkXxNWF6MNiK8u/gWodgClCcGk3XCdI
YGgcudJlj6M5NEBCL4nArQneFA5OrZ075kYCs1DEwz+CM70PgwaPv4aDNgJGouYz
a1y7sZkhRa1ooq/4d98jp1WxETH8BxBiM9JuYq5T5bvKVL+U/AXXp5cESduqbllc
YaDDOY9f00Xn9HsGaIYUhmPO1vBtsne0STxvhVeUMLBX8+/MlDqvx0ZlbDHm5dF7
b+R3guu0Hmocoovtx+enOSSTMtXP+yp5zxPiaQiQ7b0JMLEgEPbaabVRp8MkFyNu
/rolIrZ3/iSI0q6merHCYt6WRTfeGdCWka0CrPzMVtukcwhfmOjqwuCCX6YH2HrQ
gIX8OBGMFcEs65hHklure399XxmSySl+qSQJVe024PhqqarBJ1qJ+nb8kBb9tXoG
5VMH8VVqenLiHk0aJpeIxtcX2qZKfQQHl9bhf5GEPowNXYVK1OdzDBy/5z8mN0hI
f9dn/WeG/SL7LU4p4qAoHoZ4L3Brq4XzvtGUTDdyQ2PpH9l73gopzNiwlLLxdAaR
TofeChxSNRtlv6TsS70OZZ/I3havPR7gZC8VkA2QV3f9JQVBvbxel3m98/5IY3qu
laCV0C+OGOyDNdcZD4yulw44WWcDTeJLtaVUfOESSZ0q9j7412CIgHgwlNMbx9lQ
vgilEkE7uyhdlCKIueJ8eX+71isHIsS2WaLsW2Lc/g+/AAc3AgeRL87ac6sfX8p7
Sf3u0ZzrEkdtlE0P8xTaXUqF787vuFt/yWRDC9Y9EYtj87Rvtz/4JK5XLowMYWJV
5uqca0QGjypY0kOJpDgmLcbAiX/Xts+SGy/2D6wcj+aEE5v5W3pLbk1/F34dyaBg
M3XewHiUF2mhkymF6bjhFFbcaD+SYt/tLE4bv1urmtqRSWmkFLiaul1SDnEDArrj
VxHD50WYlRR+RWzSYF8kWFNPVeM4RMhpqy/dO6uBbF1Tcu0xUGsDOzu77c8BDCVD
+0nLKBlW3LcY0Zoa/fcDSjVzr5woLONvNEIpL/zxTS8eFyyD8K/yktc0X+fDi2ja
iEwPNNjsWchutFhpscHCJYV00upmIyYY9fKn6ZCDriPCL53++PpJBfj3u/+vSL8X
Yg+0QrIE1NWzCMpIEzRUeJp/SDKJKymuh0qffrWuPZc2Fk+rSJ6TpA7BxokP0who
TShiIHWpIobCSUh1iSvLipZHKVcAYpx5HcCKWaawOlJfSyQ2CxMaryjWOLKiVlYu
qhsg/k3vc9p/eM+m9qihQPH249NpzD+0Og/dySvy58NcV63V7MkVn43PeO7IUiTB
V/dlXf8GIS/JC0mN1umliEPB+Ty/bh5hfwZpJ3RNYCtEOYghGNcy5haqALt7xlkl
s55rK7YNLdK0c6xn7mW42Sciz5hWAF2BsBVl+fRYrXktzuaayO4J5FO4Jx2xL6hY
lyBn7Nm+iPr3OoTqCRlbramZ/AijbXmrGAG4oOXbTNTP9y5FQGjfEIhPHuIXT6VB
/HtX3uUnx/kcUO7UuwuNLC92+RJrW2VfNNRwQqJ6R0yA015AvmdDdnn698ognmm7
8iahIpcTDfJjs6tfrcc8ZEEV3ZEe+KpcryPxE9H5dKUWE6mUynYvg641WDMWihP3
LuegxNN+vV0DfN9m/FOKXlgmPDKxkK8bgxXwR2k5W09feTTRnI/YlzXfISLiwmks
jvNf/4NaUGxP7Cm5GWq9uC20lLTBnAZiAkXXaxWrNU16NftuCRPtSDawNnaNOL56
xOHFrvtzZWYST/LdJfjM/hH6m3DPWSikH2gkeDGM5zK4soEdx9ljcNYcFWUSBlkl
SWgVUwiPCwC0b5Kv4dpDrKHuFyB9T3YRE3VNx3LENJ9gYTPPnwhyTZORUm7F3F/i
IL/+Sv9o8DCpMIk3OJg4r26TG5wO9Ua4Y8DiDato37bff5Kj7tECzywU4pAnxUB0
fTDaz7qhfZrhUFV5P+66qH4PdCtp6DT64UCYc2oDQPfz0oSExavYRjg5OKakUlsW
LzDmINaBpAeIgEeW8VxOrJmpGrmG+cNubHKeDJMVN2WuKPUrAnrIKvDHNdiqrX4q
UoV5YoZt8QA9lJilNQW65mKc+0fakN4pffgBTkOl6ylweFRRfb60jvGKBGyK9jxY
78Rna+EKYq81QgJUuzbzkVKYXwJXOx8fEeeSjrM2DK3R+1Z2U8+ewcW4UfXKfsZw
us90LtdSgeaYaiWiVRCXRG0H0xPThVck3pl5LF53/X1R6ZCcsJmbbRcpFKNpqRsc
FKQPbNMQemNcfdMVzjMj4MD70lgBDGpN7STGbgwEwI7mmtdVVQa+dRmTyekJFWwL
j70J/KWVjmMkWF4YDoCg+6NOLp9Zxs9xlwDZNE2APHikuGiC3xi8Z1cvodoTi8Qc
FeAt+9LaA1zK7XuLRYwAvrMkRQOWJ6LMl7CEcDZDPoXEyaA5tx4pipc4KxRoOFRt
wQzeKf6OzHJgXJolk1B55xQsruRPKccbk7G0Hf2mpnllgsY6ccsKw5EXNzvO7/My
QSPFxqLMbyg9azYHAUueLFPhbs5NA0EqweB40B5Va00d+eAibmy4Qu4ayq2PzGD2
kX1IF+57+Z7rHDlhmpWN4qFPAyZ7RGbYBtIlrfelt9Mf2SLrQK5jGxYDLQw6XO6y
/Fmt1aKU21n1oXBOKO3Mzf/8dkuUdDEBM+7IN1BY3NN8OAmg3wma5lGYDJeJUE15
80oOwahSJy8ljkUIQBSNAHTEhZ6rxnD0kws/WMmtpFfddAfZlf+q7cyg5PkOkXS+
1WckOzV4K8lxl8t68D0RVgfdtgWvc2h2TwKlQTpcxAU3nhdzT2kwmyhx6olhJdxM
mn9PKZgowYHq8b3WEH6fhor+4o/Yk8byrTRlrWCFDJ05HhHPNIF3Tm+e8tAwQZ+V
XTvdTCwYGGWKWvJG+G5l18vr4Q9yWfyvUpWU9CPM4bygCwJL6iEit8oj6fx/8iJ2
2mohROyciBOTeLZZh3vZslS0byRkXDBLOiexAhsgHid5MYEOafmM01IAxdhwGkgc
Uu/uhUGNwOMOoZjC9BY7HeN95JqOQP+VJ/CtCl5KC/yDo+QgfQHoi/ntqyyACm91
YBg08FP/es8Z7Mzxw+DQIg0VPjNUf7jP+FN/PK8FHkvDNOnRoA/C3It0HWD50d+M
0jkG8Mlpni2IzizN0qJLwhpLJQSzei9Zfoc/3hzXrWHIjbaWJF94UdFjIuYv3/C0
7hToSLm01lYZQYjfDFmZM2Zyxpyr1LXCu/DSOoLgcgiaFzacCwsw1R36Q4EdBLNr
LraiWdR5YSzC10JC/NnD0k+7qhe6H2PWY8d3TWnPOHo+H7sEUBEqFDxeEKGf974h
84gQPeiysNY73lNDk9bn0b4F5KzK3KGysheXug+MZOIumdg/tUQ9+j0A6TggHVQk
4bNpE92hrg3fCkgTvbjsZQbx45YpYHTLv4dSjliP/X6hXYN6m02onO9i8iM1qzWK
1E39ShmL/eyTG4Vl4hjcV9xMfstUbEkNHSSglT+4hK/HKEZ4pg3VE3FoN8nkhdHW
IGd4Kp9ZwVinjZKqKxaVk3Tff5PpHOTi5iJk8fCEcIr390wM8RncMf8IQ3JOwJhG
AcH/PbEw2zDsf7WQbq7y1nJxIfNkBGUh2oupaL16z/UbGYzweAemdeUrp3eAzGcS
f357py4lktkDmJsMeLwCqT6YxkhXs5Bz/OSeUTrPrc+ACWHjtWsHNDQfg4jxbZoS
GU7mx3sy3enai9nLzXPv8vIk50DwTa8BLD8uMZHki+C6mAfSHw2XtNMU2OyUV8iC
VQBxedd2Vh93Lbxx1IZ9e5AVwrPTMxbhEp8lmKf7b4+DrIQiW/6X2GHYIlI/y6+3
or6wH4C1oj7Bjgf0/c+KJuyCNnUbDmIBM6g+7LymroVxXaogQqFDg8QIkdtiNKSy
Mj7mPgltJFZWXrRcZjeMQHRq9Xwgk+W7gXoX+VKRSuUHKUJH8pZktam/KB8B/nK0
I3DCkcP951ary++OrK60n33IBFrjwJ7wQffuS4giK7OldheddFynk6GfcSgEZJ79
0BdKeo1DJUU/xenFYT3CEmlomRFaEr0whl/7Lnr0vIPJFvXLb2IhcFb0/FjS9A8c
StxoL9yVyHwkYlZz9/wk9dygAII4FZggs7lfaYG2zSQZ6m5pTchiJsR9qZZ4nPeS
hl2Uhnpeep6O57wfuVHZqfATFJpozLuXP5luJbG0tPjEQBIbWVZOmc1n/gGTU4Tq
31pA/2YUElF6qlrtzL6qA9BUUrKd3UVZrup5szbbfaxPUhtbLUJz2SdghrrF0zZD
TWaXKE1oG8N8WdEfbeMu8gWA3IuN6ryY0qkJ5Tn4bR6C/PnFzk6KD1kZYlH5bOo5
t0Bu9cr1V39OrRNvNxSGTnwEIb8OWbiT2cIjTU+ge1iO90Qv8lkrIwehlf7d9EK7
JhBkUv96e5ILYLJmN5GoaHD4apfprwyCSNI82mqBwUAhtIhxW2B/kerxlJNc+VB4
9CUGImyYVj9HcTVB78qWN3tsXwIErHZPs8MzSPCOE9AuxLHkVmfJjp+XlqhfwWh6
BYHFWtDt+Z1uJV1CN+i8Erc37tHqd770AHO3yvUqa7iyxf/ieFd5Q85dnhOymUQF
G3NhFwla1VKApdJwSrozc2cBHjujQL4ZqItWjjzx+chozI3Ha2/g7G7Rm0IA9G8x
GCdicZW/piTHpb4SSuI8kwpw+/5BBz+q/osth5Ihv7bZKN6O37X0CwUHsyMOGa2O
OB1E4g7a3fjj4tQzOTDWUe1nw49AV9hTWcop/76PadxHxAgzzDvZl+7t65/KIDus
kUYyPVhktaMvhPD8aHgi5WxtqIHJVdmDrfWYGo/S+yP+SHi0r/iOl09UHcRdRCYX
H0BPMFJD6OZdkBgxSRjqWa9Xh4gTJXG4s+j++wNRUT1YpgN8CA+sSQ3g9hPAloms
DabObyG0mtNpBhMDXRL1Z47mdGf/CychTEzmOuLonmnlkEIWcPBSBjqztR3sJuFZ
2kMc+YESCHe65uAz1hoU/QauP6JuSE6XP7murym1+wMAuhUEggofVXbsUwG3y88l
/9JHZNDcgBdtjN9ysvRZEODuaFlRPK1Ar0edg+0vxx7YHjI0XheHvvq9Q+n4xQyA
gPl7MghxYpeKlSvU+Kobwf7rQmvg2slmAqfMPCnDzE7AXv8SvAumbt8cHzZoPcSr
oHCipRHD1XMC/5BKF7EYnXG9u8uj7kewDkNBhhCrtx+5qcbWrEqwklrnnjBEW/b2
wCdJg/+BCF7oTZ/8fBQ0XsMfyBmeM2Vb71VaXWSD7akQ3PgdXHVXj42+LAfrblEB
qTp8Ry9SuS8wuRAHbdXO6FbnDq/t8qqVbAN1Dk+egVCBifzuRbZ4c3YchohtRapl
hsgsXe10VpnSLjUyEXDbZkojuqZsxHUxzG5rnI5PQZ5Yj1+3maXo+Sk0op8XlXaC
gOUFsLG77lY6b1mf7SO4jMfrqErk0tnC3FWqYoVBS7VyHroQug8axUZ6VCrlhiFy
CYTnu7VvO5pr4bKPthTTls0l3tN68IGwWO7AxOqVD0l1qyz+mmDSuWO1B4hr2rBC
wxPB5XNYKVQg3+lhn2ECEEUnjDX2MImXfqhqmlhgz6kNzWp6SMsG4wVdjwk0dW9N
SoSNqCeYxDtpPdBm2jaYWl5bqNjmTzwpq6NDeWNf1AbcCOZRsZwyr2iwwfWtEl2I
2VYJSn5y/0wkQ1dSy9pl8dgnRE3zzvbDoPOpY0GwPU35Tjk2Mc/cAqQJVnAoxIyg
yRnyejy7U+6RUQ2ThgWnik3SAWUlL4p1gIVypNECZlgrDNnpAGP4PtGAdCTR+q2W
c5D3SbkHL/yl7XMn9SW+S9NHVGjCLM1+5QOZlSrFf9PNp+Jyj9OfBTOl9admMNzd
5rMKm5KFf61h8tNDHnlVr3KvnsyUJjUOtuhcyO4Q5w0mBqgYrxoUsV2sZHp17AYL
9YgxlNc4/rhEAptVOOPq3JVqFDmBAZJ9IyO9kgClYvMy+eyxmFTo6PRidizfJAdU
o9RFGaxmwCyQ8YXuPQsy63dS7gES2t6jT2wfI7PPMV3hqQk+qOU4P5ibVGe9123c
VlPtxCjsYGHqk1QJiJEZno0cDTi3REYzlkKBO9aCPVWSBk41+RBYIqLObGIJUCQQ
kz1/YgKYS1ANET+CdwjhQPfRXCD/RlzrYddlpxN/k4wq4HHBdn+UaDTnbVUUAGRp
MazoQx+A4u/ZYpIsKQkuJFk0iSlwLGt7kqAnUrbGJ7J2upiQnU2jNHBZxim2XElm
vRgFfzk4I8LteVAiIgoGhHxkJQyMukUAV7JKK2U/zXQMsO+fCWePKM5sWWGExfl8
mg0dROWsYaU16citHEe687/y4kecIswyBoX25OVRCZCfzqpvCdRSvytE2sW9FfZa
T915/xxFycIAaNekdn/R6t9nHrWwySxf2TuvBsjmGqMrpO6gu+HaYtFwAGIhvU7W
1J1g6zDIiwXYKHwQK2JyNZ83UzOn99TPP0HzvJrW6xGhWMBO6k9H+6l/22fVhH/0
vFDaH7ROaPWG4xGDBIYtEv+VEeXMH6CVM3hcFUQ4aLRtvGInVRF7WbL6IomaqdF+
pNWTlLTDEsMBuutqT8IkTYE/4r6Z8ckIdam8fFRuncS6hbxWCyugkTB8bZ/Cp+1x
wrN5Y8V1yKujMsdzp+PS5PnAeIy62vFqmsGsv7sqjcNQlPOSnvG5fMMNqNB7TI8k
9i3AGqwWoFeNqWKintMgrRxKVC26ZJKyaXNRrDYOI1+jZwTeeBB40eXdIO2cwzOi
VD9fODQMA0zk0aDpC9jgRPfT03aF3AKrSukJg74rOObWUFivwNwNi3qedzvCauyR
GF143FuzwX6tIg18flgIsmgodJ6NFTS/UwkTnKI1Vj7PaFqN4jCOp8SHG184+ATB
7CFLfAq6trCQHGMTe9lsghHJ+ORaEXNnj7LNAvKO8igWa7IjnpYrTaKdq9w4rKng
uhtl3WnQhz6zcHTEDLSyBCr9xgHsCIwzdsQRKqISDSPgldq+yrX9Mq7ydh0OsPht
QF2ZSLuii1/EHBpGWMFegPZ4jcq+N3EKzX1rHb58D21rN5596E9TG19fgFaDxAxk
9cy2yOmoUgdqVFnw/Kyz0Vsdo41jE0wg5j9Ku4HAoVqD5VlCNqxH0hRd0q86jc88
WyhTw0fetAR3fIkBNshUmdJ+wuIahe7LxHR/m31k7iUQtRkFAdQHQ7ralIPRsyED
iAvpKxyklfFBwx/oPuSdW+NtKGFwQt+T5p9ph4ypjm2biKKuksAREnsviq34PTpj
nXDE2n+jgS5UOCYOyK3c20sHi4tMyvBv9vXi8OV6/EOdN4M62douX9qGnKA3FipS
vwrf4R42zlUSCb0cgoobpBR9qWZlH87zE/I2zBABUNYB51vBhELEqGIt+AH+c+lM
VROdz+GtwjuCQYEY1y+5uzPCxOSOwENpkjBxa2UoMPucI6kd2u822l5x2Is3hG15
rdd/rziNj4qW20Ru42ywUmOASdxv2j81RgLpDUCbw1kPjQPAE+8XBkL7fCYREyN1
XyGGzo7oI+Zy9AglhsN0S86y23f+eAuEyvZMrWYYNJOVZdDfelZFy+3Ws8WVVqPn
aMQKzl/jT/PyqXgIB0WjnJOLkmHxHglJVynbf+xahZOaf8IrjV3FTDDyJDboWdtw
ZEZP6cxbDfmv5We3ctJdhvp9CCMs8EqgHmD1TZs5Nn3Jkqz3/c9RURaRb52lQsaT
0FJGIhZ52kufsL9Q79Df4gGEiUsdOhxonD8hzLw0Jdaj9PNdG6ewoavr+xAWO8IB
3o0PN8kV/baRML8ar1j2pWEvqMFB1DJbl5noaEzvbWLOI1uz9vfRfdruLHdmfDAJ
/ff915aUSzyQePQ2XZEkeWMKBo2VkAMUecicHskOcljRSnFB8OMnGMf0067QDwE7
c6W6OXFE0Oc3LC7xPt9VNXMJV1qiKmhFrkdceOr3T+Fo0IbNh+gPBt5esOp5oVgd
rEalBp1k1X/OTFU5GWtuaUZ+kQ3SfSka8kjh8XtfOR3frLA2j8AsPiWPUidcox/h
Pb7UZXdpbCbD6xi0dPFGP5ehaMB/ctOz/asDTTW61PPjDWCuX/hF9zRnxe1tUsmt
U039wFrUHC4lpn1bbt8lOqVLDSdBEnaq+WyN/x1DMj9NCbFP95UHn4SlQ1ekL/IO
JwdILzOzFgSBfDW5SU4Iy45VcKy6/mPNiZGgHAw9vbZDAZCo3uv4ZMt2YK1Rw6vV
xWCtX2ArobJMTyxww6+evnnm9Sr4IvhSY8+GlBmrGojRSsqi4bmY32uGDVwFO6a3
Nsw5l28N7IsgSWzPwRrv2JoVyz9BLaoQA6/2GUpBRRvtA/3nje3rvBhHXL7I4VyE
4DusO1ajW/lgBj203dHdr9N1MXX2tp5ygOE+B0U9tVuEwabciTMs9SHpmoviH8pF
rTwBUHR+X5mqWVXV+ho14IuTJ06aj6ocySxeW7SwaaoBRINKT74QIjEYg6bDEpp9
eoR7wzfJarGcEtdgmikN2kqEMEgHWS5iLJ6ieaXcaNTOpfTA6gdk6rvfs8QqfHw6
ArpSq/O3CJ3d1uT/Mj10eqjHeeznQXCgzDlV3eOdoVzZeibRFdDSlRbkXEAjnnGr
hUx7+os3ADwkZmpi/rxJKojNjwwvettMYDkRfm53oiQFrLzcAvvFIxOjocbOlP9P
xzc5K9zXFZHhCyePfXg+gZEXErisDZO08zIrrC6oujGeYttISAltdduZ8SUzywCn
EaojM6dfv+wrNpZo0K0529+VzUmLTC0TVcOskEDJV8Ij6ponjDXKH7hV+W0+Duyg
Vmk0aY6gYMb1+OpEXbIr5K6Y9IPkjnVHbSZFP5ROU4+ALpi11WaJIDRIK73BOcEh
PPE/Cpxp3XAyrnNU9wZvxxlu1IEGOysb2CycAA2tGenJa+HFa+WJu3zA94KIYFnK
QPLUQaFwG3E096RWVk9Oyxo/EVQ6t/rBsqsdqVSP2vAhb3t7GGnurceEwZEB2IiX
m7R8QHKYqrJsySrRh1tGmx8rOA4+d6siEhCqYzBknKZVeuL/Oc6SH0zEW6s/6l5/
S0lA8WTBV7NumP4gyH3MSZ1NlEnigwvORj1CD9xRxHV/IuiFRdNXHvqzy9Rk+3Sl
0iqkZKetn2uog6jBKa86lX4snQ/0WZkE5mBAVtK0igH41FXpeRyPJdZyzWQqdkqX
hsutsGhDVNxoyXCyh4kIDUGSUTyCsAz6kWTUK/3RJtd1oLl5ziZx/CBXLc6RkVXN
D88eSo6Dlph+WQykG5fYo1gcJjsluJB3HhWaioze23t2qFGutQvQ5ANIVyGZ61Ml
CJ5VoKW12+S0iLbCPf507/61m3IzfGOG50Jxur0pNaUYAmIJemF6ctMIPYquDVLn
umgetXSUe9ccCt+/Z03JaSAQCdRnsoDR2FaPRyygLgCm/vARh+UVxbr3qQ0jLlyV
K2ljE4jy5s6wiDqkA+By6sAS0khHgFtAgrtNXHYMssvHHI6IaI5uXkkrZe1stS93
N78HbzUDIxVBQTm7m47Vg6+V29+4v5OkceFANrfnpda6MF3Al+CZgNEq5Xaw/pjI
FWuFwy6oO3CUtoQA+hvF0PQ5T02ALYmhndd5zNIz9vc6y6ELmEwISwUx9RayKEql
rOpYA7D0tgMkWZHAX2j7hI016RHROuziG6wD0cg5dd1eYvsiepURVa/LRul8bUuT
DOjl+n1DHM8xmMqgzFDiEq1enTzcCdEeDKB7KG2R+4Atk2EUpG93uxF6ejXjP/8t
JE1l02kuWa8shm93bOAr2GPjanqQZw5jRWEPDenVEtQ/3D6P0YwYNkxIeStGQzem
1tC4TWmENwR1mDwA3WxbGjjmwvKJezuQXUdZJdUQiZgHDwNuj8lredxrOazt9l0l
Cqlwc7bcZf4eem5sThE1xH6rH6xhUt5jn+/F3EvnlX/OtAgqHQUqGikIIyegvsSc
mGHbwwCRk7JBst92S0M6bEVRGzlfpeMlnkT/iLp13mRkDN2fQdJlzEO0G9BSfG0q
wl5SG3IrMPLsdgAHs6mrgySkAMe2Han0mpzc5zCVAR0H9s1tqqYD8D+3sU+Mmtlk
1FAPWLwD3G9OIBLydoviwU2q+/IgniTabW2P5uTlH4Klpyqk3OwA/4/s/zypRieW
6KSrbPvCuqwycy/FH5Mei48BqSiwXqtiRsYlMnAQ+VZlM6gHPjmCEh63j0cJ7kIM
dRyK86S8PraFhO0YsaCM1h6u7N5ETWkldUGUwGU0T8JIEgnkjc9m2+HzSR2ZyyJj
GFvxAhsouyJclMA6atCICxkZZtrqWfEeBFW7lAW6hgsbPhHMkqLSatQRk9wMswlR
i3UENMiDijMIhewGqQzIrk/QSEq1j/S/asHW2R1+3MpdpmW4kbCWJHyCbTVw/U5B
HRCdrVKaTYla0G6fu2dzCJNvs90F5KQvJwfrGTnv2OMj5Z1V5vHjg+zQsLh6UrtC
sP5LwrV1UsQaU4Tid1O9YAM4ZFZtsDUxgJqLMUkgWcUd17b6wc+2iWioJyl36lwD
Ng5NkeCNPjFV8YsBb/ocDBYFAbF/taBVSihaPWcLcBp7et0T3DnsOn1EQ8484wzP
MPqYmm0gqCPpL9Yo1CYVAybqO9ffxakNRFsEUj2PiJGsdIAt8BWO0ZtCYdowz6lx
B05MXsWiJ+fGjyMOlUQunMpNEFjDWM5Ig4EWMIcgWaOTh4GwiVrpjWzvUUY8zzlD
0XZijukanaQ/ks9sz0b9m6qNjdwnK+kn9beWVfy4xkHnKqSPtmTKeouXJopOQgdw
XJbP9ztI3I6kAUGg/XnJHUF0vjGq9JQztrEpsIirUJCcPjRrZnNPWDs4do9SoHoe
5OgR/MUJnvuRLkm1eyQK/Vruykc36JuEtv8qqR+ghSc2f/dLTPxs8stuyKbtYLmD
hCMVI7JtSWKAAFwIa8hKrk8SlVm+/aJcOr3vBnR72y3lR2LQSx1TK23InukFHGs/
dCiBbJDAhUXoKZnnDOf7Ckx+7knhwnK+DhUz9DFDsGdKjSc6xVqlrOTiehFcQNVe
rfJhzmzYKT+oZnaDeRCsM4DCduqvwwyvzdmmL2VLSfR+5nKUXGp2K71KoUoSaN9T
trtFNoUmw7U+SvesLur8xgrU7UAk7tFtcFGHpiG7Cmgi+9IwD/CbdUkuNfqHphHo
Y3NVhvJRFVqNaeLlmIvgIcNYDLlmg3njfamvN2hfIKMzXMIpNAA31olWWZxBsL03
E8iKesClD0VNpr0VwHjHlUbK8aM2rQ8Zh3oQoahoTxKIV9SHESGX5lem78avlU9v
SC9gRc6Xq4LmLTzp1vhViaNQtG9dXjjFrk/Ks9gkN4oKF2fCgCLEz8fdOWC5OGSm
qEP6EuSOdx32xHTiFtg16sCM3VROHoXDKJE+1ZXQgA+n4lC6grmKBbgx/97/++0y
pjtmTKXjPglAy9H0R5Pq+PGHN2hduTwnQ4e8gkL/bc41I7FLsH/oCmv3wbWASHRC
od5QY1cE9xTU8oxrk7vEA3jsNhk4uGGvmbdQoE4Tl2JtPdG/WZTp7PwRbnjBGOxT
i5pZ9b3pDkMS8fpLP7ZxvbrgEM3sv/+3RR07PttfksTaouxzj4g0X34MJPizdFD8
+Q4SeB4YadrSwXODuHFv8ak/gB6JiF+zWjhKPZPS85gVaNtfGqS73Dmlo088QRc7
pBlua6jfW0aVPiO+HegQVSqJqZOxsJEnifAa01QHoUSknTmhJTB+9jx+wtjtwn4i
LUAtBg5obmokOJRHbUjvPcGSGq34RQYgLf3fT/eBQlZTa8OFvdnIAsQxGNkAjscf
ZCAKI7tdJStsxQyGW9Mrnn+4be78HvokzzdPliiSAjeZsecmsJsWj+Nja9sLeBeu
OeWYyJ+vLcxmu9jPY9y2GiVXQCyBi/RfEENjY7w5qivW38+fQ8GayJ9EaDV9M+nN
Dyg180kCTpvizl26RZFpqQB7e0GBHDi/TMxRK232IuIRyjGTiT2+nMIInddH/QqP
Jyg3t59z+60A7zefPvieg1HPWl0Yv3RqKjdAX5wJoYEZo+KLXlEzZugK5ABAEfzR
rv53VndtYJ0XN+T6WUO1vBh2MIlpI3/Wvi9Nc1BdkQABHHmj8zXBHInrWt23rvDN
SbSHekZ6fF+SCFO3PzqKhYp2nUnisrJITG6ithS0yLPD4BDDwzsU3FfalRyAon8s
jkxZYhP7ZY3Sspq1CeSmsWCeZ3SIosBjQTEkA5EqYH9K5usWufohHtabsGNgsbzX
mT3CPEB7AxjDGAwEEnsY47YE5rl9QO9bfW4xRbIQpacZWMWzK4G3jnNepy1tq74h
DkuwXaWkY+fH0DshT9zYIjSwIvZTwFDssyq86BUvP9JRb9p5f/I68anfRTHZTT60
lw+uf8DFs+wHFB3LaUupmqvzuzDmldXAhaBJlQwokZ/7JFOx+5ktw9/z7CMxkHg7
8YsE5qIAnx/8zCAWSZvnkC6yyMFaWecUNeYhqPvGfTV3VAfLfnwWrxDwM0cPQOCj
QdqeRbrPRNVzVCJjnFxrstMYKLEmiCoKnS/1qiSWIced49oi//p1Rl31OqnaBxYu
uxNC/b+xgp8P6z2vo5cz+A/dRbYOV+uONSrI7dOj0MF9dvVw9K8K0IAIb0nxNfS0
N0QCBdK0Nnk7wNHdaK4Kvnxux87sFNIzHvomNTGb2TKzIplj3aH+Z0XWkvU1vpDU
bV1QBasum3xmUDOv9aXUwJfFpZmfitJDrqwhSYoO3fus3IQ67BMlaNshSOXl7p8S
4lzu74iUwvwfntLDojedZoC6cfcx6rjWAYitoc4HZE9pA22ypbzEg/81BAGpP9c9
mbt/2fbh+mGVs3a9yZ1/9xN6xXx2+mQKxiJWh20JJyblSi5ZGtIcoM5HefUVKPfF
l/Jc52kh6EnNe1N7pOhJnb7EicJ2ZspzUKZmsRwmx4sRwoDCu7KX66j0PFEbAZot
cQuQokjCYkogXaBmHHIh3TRw956kr3EA0U8+knSjsRNtmaggMWSAB+AMEJwq64Yn
3I44FlIVv4a6joVmR59xJzdi6+G9OA4WvIwvwDKATT8BLwHFCbRB43t9FjsoW9yj
97+fEV92BUpthUcAehHSgrVXQZ972WtP1AZ4Z+lmY3lczWvtheQxBYwDgyjmXgXB
7ahJKdnAAnE+r0FG156qjp6xGPeDEvYqXdxBM+husaxe44r8vclqVvC9Ga5UFpc5
sV4pCQyT0CsSsHbtR7uMRRpNjj2DOxxepDvEZzDQXJAQBkCbX03TavE67cgVnwjV
0Ps2r+x+b1g+u9uPvM4gDnx+GtD93fCabZbXumxF7nEjmP82BqLmkw2i7xklFZIP
G65k7KmArsV/8dVr6Ee/JFcHeZKesEW6FDjinAWk+9ELRdqcpKxJRvcNIVNmyy7a
kztM7uYPMrQhO1V4/utATvV0dpa3QO9mxQ9kAsT1w1t3GMubIzor3Spx1LVbLxfi
ioj58QYyq7T1aSKBrE0boOQCgYQSDQgls9WZ01DmwRNcTMsoBw5SaAbDi2eqTfQt
jw1PKn45k+VrQvHGyc+68ZJbhPVEjN1cmfHllyKy+5i3B60X3vD2FtSyAQGbYcVj
T1LkbMd9xFG0i2+vq1aQNNCC8G66I/jnOm2xzl+APaQQs6G/1t8F58GPd7SaAwIU
JnwT8T80A+4JDVs6wxOqUIdMjEfXpmbkizx0JRS5AwgT8DPWnvW3JModGX7eCf5H
YVAN2xwiNDfTKkwI3O8b2CG31ec2KoccBbyb04u61TpbOzePFeN+GcTFwZ3Tioc5
ZdMdWQDusHubxrUAHliBR2aJNW0cMKFxmobz/7/CRmg9aAmdU6tYbnB5/jABA3Df
RNvb61D7FQDgZgdiq3xiW/YBy0PYNq7oJcXTm9Oq/X1XBTIEXL0kvsUBNiL+EEvn
s7jNqkZwgVYOo2QDNizhkzsUGJjfUXg7csNVJ/sQwqjz4lgBvCTRPsFK2oFfUfVj
CahTYOwNoG8iWhdIm44aBBRiWAasSW/yFF/tjq+0WTQtFaWgZZij6oVaAIuAd8TD
onlcaGFxgODzPLasyxtjahzrVMxTTqjEcxhqSfKLk51CWECTyoSYfwUwces1of3b
sH5VW8VXZKGZ6BaZlBPqz1LDN4fRBu2l5PQcFUlmU545Tj2QVkeblcSTsVGclnTV
3TY6xsl98J8YHC50ljzVJKpzXvBSAaN7BK0OvDrBqRTpNPJWo4RsO5raivd5Qa2M
siHDO3L4KnRissED/zOQ1ZI2FBeuEWbBQlNPhCUFVEkhlrUZK4sNsTlOgVJHP3MV
YERKslj2jMOfrO+xhrhU2zEjuR0B7BSu1vcClj/Sa1ZCNnUUx0UC/SDHZF+KRw/5
V88ZmLOZ/9LHmHgKHx7TnDvh6A0rM9FyNHVLrt0lkWdALJWMEQcfvek5KY0puz1u
ZXMZaOjAz+oJIxLvzQongguJFIJ30/pmoh1OD9KfuA3AgwIFbTmlFLioe52cC7qw
xxclZkFXREBNo5p67afWzUIBJ3UBOv1116csHLiZJKz6e/Yl8P5Wo7iTImzlU1TE
hhyYydNGFnMXQHn26hzqGpoLObDaGGU8DoTSKPMz9PkplZ/aKtR/QEp5N1g/BCmk
OSgoQS5Qd8LX6dLd39Jlt1b9B2gbjo1qpbGDIcy88gujvSx6jECAmcb5vxJK2Jvx
yx9OxtH+yYo5wBr2BYoZB+KjO8Z5wO+pK8bT8AsgP5DkpwpMhbBBMEdmrd6ouoJy
NSTVPPkqh/nT6a0dlPZMmLqduhvLeZbTd1ekt2BmnCx/CdV34fAqysIV/YVkLPCj
RLVo+FMBRqcfCPQUjrGI9Lv6GRD/MteWLBPuMWxCzCK1prWL2bZ3iMFGWxNV7NRL
KEIToeWgGmZ6b8f/1PmdL9ktLZrgfHvxvYuzX8Nm4Jfl1nPbYMBJ51H3rwVWlI7Y
t62YOSFg915qzaGdnMJACmW+k/+5H2bn566ApiWrfTxnhl1b9Li0H2FGF7uW5bEG
x6yV59Ky5BiLTBRLMx668umqFxmLpCaPdEh4YYl8rBMgfPOr3lm8cjYwPJLZb+o0
1Yp8pnxPbr41MYzpnT+U6naY1+SjXXaQy1tx0rCAmhcGeCEfdctCxzUFxCppWEbA
5Nsj0ShJ9Fz9224IU3xd4jZ2Ev7qMuBaFrvIWuK9YWHkSJwj9PfBpfG2OhSo1A+n
Nuo6R8oB261ue56KYPwbJvNzAx521jaECQ2EP2tKpdOJ51SoAcAxX5JujmtAS7Zh
RszbCerxNk2svVEAdkfHwajHqmP0SaPjN7Q6mT6BFgq19WxGhfh5DOul8OGhiAFJ
M8HTcuuwErlN7QwlsYUzGgmJUX5mvu6oGA0K4D7XMhFOJ9g1RyZxvrVzWTzhMhoe
H+IFGkGj860/TQwdZrOOPDMt1BVzrtQMzt3pnkUnIix9lsF9ZdAH1oUZuxRVsP0V
0Uky2d2uWymEPN4BqjJBbRCVW+zP28krZYfyfRDmzc58vvZ+1+ECWpRru/biEBoQ
f4MBeqfEs4fDcKdP/Xci9lsv4USox0UjcHarMK9BeQFMmHJUhBC+f9ZrwxgqYY3c
nhesjSLnn+OTJzsAdyMzfdABTm1VRDY1tj0vBFK3yHk8smolLvc3kDGqPvrzeWB6
3KGZjoAKBas2j6ad2Xca4RIR/Fgjbu2pOfu4HWfmttrcLr/6wA+4+fUzwF22Zu4e
HqUthD6o37CHvFrBd73SQVbg7m1Lz36UxipUZwGiKSkw2gLnCbQXuS6ROaWvDLOA
4QGY1Zv465ixvxCOV24rA6aal8ufhBC6xx4sbqTHDGwcBRVkxVTRcItHSSYP3TV9
B0XygOWqh71hgiyfzsSPhDMAbigPICUJpxsK07LQKGNCqbw60yCNff9QSKsTkbz5
XPMO2N45ZX2o4Gc4sm9w7A3RFGUI5g9P9ADY7CVyOo0AZ29coZ7+riemE2XP9Rdo
udfhiXdQxC+tCYWOYd1+F+jWeeqNODfCAEabofIszwtcI+tW17XJeAYUe8dAuEyv
f+Utxoul/EMftZd/W5y1ATwRNw8itq5rxGO3e0PpheY1tWD9bCZKOUhOsT9zyZYo
+RLwcmeUGVFYFJZZpM8QXNMbBUrZ5yLKNaFMcafRrDQumv6FnkhKJvQXKw3tBCy4
Q0XHH04OVxZM8AOvllVG2Eol7rkVcDAT8y8b0Npx69EPffkU0BTllxj0IfMTkF4b
kDWZjozx4Cp6Tb9bQhfCqYpmspx8HbA7Lkvm7Um+GsYIfcVbJX5bIWcShjcFrJUY
SFTqKeyTGjH/mZ7jE0HFq/M001vMVbgjrWj5djkEFnT/bGt+gKmDGWPsXqqlZa6y
9FFJC/nh6XPDkx63IRdkaufiOt422g/8xe8EBBFqMY2pVUL7EW3bMSz4g62SkhcQ
2goDEo3mOfb3rGtyuZ3rVhTGUieQb6xYGJjUTSqY60cKAEB6FaHyqvpd9iA9rcfU
8lDbG5bFECfecffy4n6BMPM/vclHGEgFRDbCgXjP7IMzuLYnJJdEbqzk6iOCX2Vk
VB5osxVFRUekHSTCBtD87GetjnCjgJZWAZhibDkALQLmYo0pfsbwHdPeGSD/wPxr
hic5HenKRi0KbJAAkldDkFQXYBXMqd1iprgt9DGtvP2LkpguZcXFb+AZgaY3DxLi
1FTIQKdIoh9lOFxpGxFYV+DvNyoqQHTYw0WeNpKUJ6aFPBHxzycvku7gCaEB+kRV
OzfkpLr/nhL7c5TyFtDs6ueLjngITSe5G869D0qr/hPz7UuUWfddPzvMBwMN3eIY
3Bfnz2vTn+s+VirVdwqV0fBS2iem5VlEWDIGP5wuMfVR9IW5+UCTUqcsw7Zcy29z
UBFBhHwALcqOgy3Hc+6mzXZ64Uo+ED3b2IC92wOtHYu51Zdn0NCJG1ckw3PZkKYv
WCHAJ7UBiWHi9d4X6DAAxY+Ko1vpR3g8Oc4KdpYbq47a6p17n2mblp4/9Wz7rXm6
zv6PADtHbf7TYX8tO0TKcJ2a7iJQmO5kzRNI0G/0fwKBzKK8WHp/s+HD8EUtBmmO
CIIhQlAiwA2D1vw9vOJCJpp0ukXn7HBgWUJGupWKn5NakXVdhIk7B+WDU0XPTQ3R
aDzwbfeMX9HkmFUtouoSncrWIfnJryjhuVO1+vQDLCiQrLN1yNkK508PumIFZ4zw
6BoyEJgTF9yu+85T0eBrIqUhEkSfsx2hpM9m7U2zT2ws+Gyzn1WFiCY8Dz/9ZZw8
DXPaTZ7Dn0zFw8hyIcBmszA8f5fPwAYIYmhD2FIZ0XbxS5y7RmkTeg44sW+5hS3N
joAZecttzdfqXgUxyCv8X4dC014tQ5D93yvEHdOewXycKCmNzFpV8nqMTmMJkTPa
KN4CdGmTcCJ5606+WqDMso/D7OdZFwCCXCvb8pp7l9LKUZRbKKtz5sbjO5WkBJVR
aNIczlfrk17MRexstz8IbYMXwv8buYjGLaxxROnUHyGw0RMPtTmsvPfto7xWpbjb
XLxTRVMe6Fqp9QN3Q6Knm7nDbY5PY7DOjOeeeE8wJWNEzdKV2FiRwZS5PDt254rK
UOoeBQX9A1NF1Br9rts4FKmLWoh0I+ktniAfyrPfislEP/IPFKk6FxqG9n4/ueO4
zgJBHWoOqrZ25PNj84loqVb7BMgLVSgbo2U2K9EBCO929wIT3QdAlJGCfVrQutVt
1m1idLzW+zKUqVfzrhlQxw7RDkNfHFNH2vUM1rF2Yy8fsuk5Hn/vqqBsNy4fvpv3
N2Ju21MJVIsgNyZUSTzFXU0yvmYuiGzQmPctpgSSOcoSc8nxYHEN/KprpavRF3YC
jdsW13Nts3UTCGa1aO9H5fXqPxPGSY4DbgdUIGNOhQlWV2jNkyHpaczc/ZH/webj
w32ssnY4vjdxBfjIcJteX1OEMBgkme7+BeTtiWVqz11KMlHesUflDaz19lSp0wJh
N1NBerFPEk5WOXu9Y9EPQg3oSEUu7T8tFRAY/vmLQTz0AEzsNNf7BooKiXIrxtj9
QOruLkvgrTBUrxi7H8thBRpJuDKX5/m+XXBqnx7JX268FWpieB1vqiPxTnXy5h+E
ygOSFfYkvlyM0Za/GomV1x6qEx1f/T0+Ai/uuPywj+wWSHcrbDaZlN2LmPFotF06
WncLpJfKoLnhd8mKF2ffrjcaHZ13v+1RXwd1FBlKl8SFMehNN/lxMTgL1Z88wFNY
eMXeUAUgqW88glRZVqM0PNKNgtPXwRTrzXsPv8zTCkitC7wL1cdt8Dal4/5MSh4I
Cz2tTPrHVGi0KAUVJk+6CmivIHcQ7BPCQvgynEcPrlKngyeb3qpN9lU4vA1R8J3C
VZO2Jm9eh7DQAttmEkea3sR2Obl005Hn2884ofBDbVUhpFW+mPREEXVe/WvE0t/M
tARfpOLHlrw1O2AcfoaJ/TGzRhaLrRxztlozuUr61IKPolUiilapbZQ3sF4b0imc
u+gK/bqj5SL4CYafbw9/FRxZ4r8KEzPvk0mtY7aZWzpTUziPbTpYGgfYTM/QaSrB
aFCZR75jVVnlGxx+daY1BhLRbpeipJNsBdHbMN5uiDti5UQUhqU85ySkbtO4ZgEX
K+QGEhPBVhgO1RQQycDx4YOjW2jkTf7Dku1z603i8EJWc1qwy46+xa99uwlczNdS
OhpZyNo0GunRL/OIXTC75N/Ru51VJ0T1GsDJwOXQjYHSKEQNtr2VQ42yqqVmZzaJ
f3lg4C5EWEQwRSL6f90I95G1OwlXjfxk/gUiDmZHLJakPZ6rfbyOAKAekPNZ0f5P
sPdMF5TAmJa6TjhloVqTR75jBcTjm6MS0+n45U3Hp9OjewbUA5qyjd/3avF+QC0j
KqdbjF2YuF1NjSL5V7Tt2oi8vtPVpmHmMF5bxUpco8IGK7cnE6JgjUgTW7F/WM8G
b72dL96IXYPGH+wbrvkoVGg5neUQMEJP2FrSgPrchex2adPzucgHtxqxvrK119Ib
HdQlS2BszoevlDqoKRT3+kDzScgjSneKWdVzfb8ZRpaAV6LhneE7HorhqtccQACs
2tKuoq4QL51tHreopWMtqTMTNO6D4miHfY1FCeyTcmH99JQjTzTpWaNXSoBUciC5
YmniS+44IMSiLE9prxii+D+6LG0exSK0OofIuE/ZGurZ4ntg4au27baVNH1Km+M+
SjP3YPX2vAzoL+Hs4Po7Iu/GmEkVcJ3q6pA3hq1xTK4zOrRBaxdp+3awa8ZnFQ2f
gsbfpl+In548n+UzKFErV285d5k1MMLCi+T0jxlAeb65DvaxO0pVnGOkWHx2i83W
qgbXTpRENvxBdVFR7sgom6KhaaiIndOcHUHDrq+G8Q9mUxwC5VIw9LyBKCeNXG3M
QeEqbeHWk1fk5dvwkcITl+f7FjmI6CN4WrVj3SV7ARF73BtdnCllWPXSF3QND25I
RzI4LTNua9OSZdhPw/+k73LSaY5+im/XCwG8o6rx2HOA2kKBWG6mwvx95yvfHd02
EizLFQBQRdp9Ncta2jWhrVyT084hGCAD+/yLo3jj/t7HXn4LcZtvanT8AJH1Cfzj
u8WDlFPFmrWy9wq2BtwgqZ20D8JEI6cQb+5zoobMOlQoCNWsUvyJA3XDbZzxbzOz
M9zHuHb7OJHbROR+fpIDmFNWq+2RsdpIhfxj50LhZLqbYHyoo496DGrh7zcULaJ5
YzdvzHCYMFwtwvd3g4Ys71MFFdszzXvie3nxaz0cvh9VRx6jGr59cTOadXwqfrV0
X+ShwHo6hLFynF8CGdAGIeR8a6ampEq9fKfecoSlbWivnWm1YCqbJtHvJQS0QJ6U
dLasO6r4yulL1wWklbIiW0Qkql79pT1bue46WHjUoOzqojC/pHIT1y8kw9iXek4X
DBR8hpJ1fQNjQIoRLHp5tQ2a8zbtBKfDfeLcgw9KOpWv4XbSJ9I4lRGvs06rL/mO
MIXwQ+aknhRDYGv+Q+aasURpX6BS+2F+ryVmhLG8wD7jMP4oFkKhikEIP1AP2SVp
fuvhn8/AsH92UKNmOynTAq986KCY2xUOSZKv2n1SToxNoEq3KH/ESlljWQKZfVp1
9EDvwZe5fclKJeUNCpBv/G2s3vQJQagorWawY8zC0f0FKiqpa3eXxB/vfLHVwciE
zh39mkN7RNvxqM0OG1yfQt/ph5+4aXZajtlc8Z2fqE2Dixy2ip0Wtxlpjbd6kG06
AC7AGRSarvJ+CYzCoUxbIFbE+04T4EJfaToI8n2n6zp95b5ma39LeIW492OpnCjP
WNK+VhZtU9AKq+3mltI26XBvpe02eMZ7sD5WLInAKEO29acAPf+VgqZh0Fe5Ks9/
YEgTCS/OVDV2iO6ATR7xUCsOCTALo6ppUDJ5tNRF6WvAgqKnoMy+hRikJCSZVb6K
ahW5gY7jc+et06uZRGax3A9kNWGySn0b1+TLZj6/scDJMvtohhj44yvsEln5IkwE
VCX1b2+giMZKYHXhFg5Crjb7st02sC2Nj+oyFKeuaBJrhuxe4BIfflUpjGzQqgLm
MJZkfXo9MfUs/suIb66Wz5c5/+W/2rIIVxTq2UwcTw2NbHxnVwO5NtLndLWxjcsm
fwwNAakO4L/Srajqny7/1TxLBe1Wd59m5FRZV0I5fQzh0oEdiJx0y5Gh2xG5lK3u
oiCix7s2C2M8b8PJHNwdyvB9tlhwk101w0stpV9bet6b2pM0mGPpevDg7vimYqdz
5Xf1l84SkwS9mmA+xARCrHj1rIdH3yzNCDyyHup0tBJulnx5e8wJ1K2w1RhGXBxJ
LbxvLjUI6qgBIKm8jK12mCxmr/rRPJHA3kkY4yBVALbZwcm+/TZiAxeqk2OxZGm9
ZEX5jFC4E6jLnUweM8wwTybwySQxliKlTXid2pIoB0CeN1+eXMSy/wuygiVRmPuZ
mSYNQ8/E8DZs1sjCtNwAkfFYP8XkI6XbUNdf//w4t0wCUivQGejrSinlyaN4zKDW
4oFQnvUOkeUGfOu990iDNPHJ7pfK7Pzq4Tkit/j6vBmecnmMvdzu+O5b2/bIgc9b
LwQOCi1rgWHk9+bCuiQ+9fGW0QFzag11iFI+j+fpOBoQ5GeexXgW3A6lcN7cIn1r
ChwTVMgHVgX1dg/uKZUbCBEGytxzayg2it/UD2302X8kxn3MG5TIoLRO02BKLV6c
w3hAps8g5UmPTQ1vCyP+sUU9lv7novCIEnb1Sc2p2A6xaXyHtHpTaNpaO/7smaRf
bIY+m++EEGwLJeWZCUVHBm7VsA62NW3/4FLSOhcxcF67MghsNlJcwLIJdcNM2hIA
c1Q4A51V5HHjHJcBcyAA/28vivwMqxfHyti7Fm6V/PMx9MJ41Mt5ryZ0nI/Ty4lz
MMWvjGayHFfAtcxrm2y2xA+qdslLi/eeaGIZfNS7H5QHzW02F2zF0cI6aX821j0r
QBWW/FjUPnVVqHRxKw8csZjfZchcYzj0QQnSzfslqg1BkaPP/myWux1TnJgo7vcd
gUPHy1PRgpG6/tbHdlZYLHiu1QJnaBCIUo/4S21n1Ai71jgoaQLoehbKKWX6IQim
JYbz5K3soysd1nviZfI1tr4ek4a4xzWcG/k9SmkSfL+xUyeDtOM6HxY27cC44V1s
L94gbMbuBznSgLSarJdvM2CvexaVeA40KNXv2DBRoitU4hyD5gpyfX6XiklwZQDK
pfVPokktDf89xUA6EyHauDKHjhsuWVXuY1fvj9UiM0EWWQBkupUUEYwtj+yGckZz
PlkKAI0V/CCt9DqoCfS7sClZhHatHj0d6oKNAsNmsdmkfm1I3epk/yQSTjOESKS6
ZGmLkBl8vDeXZaH4rLYhhrJOTtXv2btlQz4e3fHzx453BCxZnIUeAjbXQqU9FRYL
nZ0RoygBlM3r6UVGhdcbD15Db+3oPFVO9jKS8rKS28kZdgeoWVuV3SIDByNSLqDh
Bg5CXU5huQPyoQ66SAwupK8sfz3L1XeeZGEwZSQsnVMX6kjeorjgK5ljkxnF5QqU
yGoVIi+UxdcwzBiNVebIW5d8/4IHeXR8VmIIBcnJdBQYRyd9TjJ7OuqH8E8wFRh/
3p72q+OETS77M+VSn3Vc/bNPNh5mo6QdllqqEo1KlSH7248HAZOuYY8kIqCn9f0V
fD0gD5jbAUDB7ueMLRp+2Tf2Gf/Eq1N+7Aub0/+atL70LP8Ge5dignQH40DnZo1S
jPisa23hHPsRG7ZB6VlmwO/FAN7EN6nL+8Qt7pHPBvxi5NgCGjDevzkAvbv/NXqR
M/adOhTs8zNRfx0wGexm2I4MGb28WuZ0dL6+ZgSR6Y5cUBN3qkIqBN0sjdDtr2gL
zKFSKVEk8TjjIk6S3H5/ING2NhKNROWSOad/PYfkFAEZBmXgq5GfbJBotEt0CI3/
2+BEYJEEhQkwR8AhuSwC3swn0nvslhaHmTuFo79IHZIstTVrYcuATq7Ub0E4aDHi
s6f49Exmy6jVGn268z7UCNtKkeILGz8A7XaWSkzb4TRTcIhV9yVM4R6VSj3WxTz0
Qy8utyaktkH7htqXmNO62LyiHd3zj3SqYWs4mRFTXjlEhS2PvWymulypQdCDCLhx
ZL+ibctNS7WpTqyUR3zRWPEERYUGvsDmZpg01oxAgt9MDXfo1fiAO7i5jR27FMWS
uuWULWXEOh2amE4s3dkGsgBP7Dq+SCjDorUGpUxSXrt0sDirDwnV/ULvkObZ0Pfc
bjELQ5ecC14dwQhhy1fyZuFvnRrwiuqxLuYMIVjoAqOh+wNSNYwJc/oqpbRIluk/
K4IleFvsqVde8c6vX4+8Hj+EiUaDji8hax77k5DwJqAvFelG4dHoL///yGvRth0Z
LSAGGnO3CKE0XOHfpovPbB0+JigaOQJgAHj7A5pJ506f5zxd2o1lynE5+pfAppYB
5rTBRx4uD7Yu6asp37SYBpHx9ei50VYakeICuPG8l1T+aeOLAIYly9FJXo5ydxOp
KxKZc3UeigvDfvIycQY1w7lezSi5mhiBwUCx9c3jqQc6NpuNC9N0SlNjdJekL4fl
JQ31fEdvlBmYFqIZGDPOsFxVj4OZIBE+iek7S8cQPOymW4m5sE/4WRRtxeSKBg/s
KyqhHgtwYyqSXycPEmDGUKb1561aHbsDNoSLTgRJ2S3lp4BZGA12CK+9bBpmmx3E
GvlsDd9j7PRu1gbYSk8P0R0txcRisXNataSrZ6oxmqHOwFY4fHIHjc+N3cHk6u57
DIEfElhnYwg0lr4hSAh0ec8HBXH3/SI2RRbtWHtM1hcwp71/vdzltQYh++vdUArD
SrtsYJkc77Ay4sTXXaTPmneSxjDo8zwsCP34OeiDNCfRuIjog9VjbtENlokqabDJ
gdLuOKUDPIrH4ofh69Wjhj9aq0yLzsJmW+OQhfamj35VGqX/WGUEMMbrOr8VMuwh
XhSA8+Q8Fu9bw67R61VUufpu2/DO6DEAboJqSH2a/ysl6mcz7F6ONgL3obqNB3L7
Ix83aPlNWihkEZc4fMsQQsN8mHUbDmd5ZpssbfcbLgz+Z31UmvFzasytPz7e5iVC
3+uMpssMBjERHl3ZxkOuRZ0mzywvUs8Ey86Su0x1puFfHFAnEFk0HvkQDSj/F/im
SETXqrApXdov09aCHQqzuoFvK/OIXAxYpubsy6HP0POfTsl55nE8K9BYnJY6fu6Z
+AEFikqxhEBMNY6+XRUDaNNujkiZyfHn/bmBPDWk69ycDD3H3HZrQ5WPiLUiIxCg
xtY+vhIqjyB3bNmYasP0nGge6+ppkD8vDlY2bSQ7Iffuh+Pv0NSSDYGOZUASYFUm
dDy2xeD8Cn56iJIzwnu4MRqa2CoKPOHdabQBZ2Gz7C5ZBHT0NfGIdnhZ5qjBac+M
bON4hhM/zS9hlHK6bwVbV1rcAyuB0wmGSri4n1Sv1zvaTs3JkqBqledh/YTjksT0
jmApyhXM9fsZ1v4WMrla1zuIP47lLSRT10sc/tm3Gec6JAAJSWeCzFWR+NjGHOYr
Y/oBOVcZ79a7DeRmTDUp2l8qZ3wAidOYBGjTSXOjQA5LTRKeB/2LI8ppCKgeE2SW
f6UYI9wny/OxdQmB8krcX3ST/KedtJDMGwNYNXzS8dSWPCX1ZztMcC34QfiWDcO9
IhgUnyaLzQZfemp3o93CQ2rK1sN6T6IWNtoxrJxc7ccaciX9skp2dBATF47yWALC
DinoPkYeWTaMUNV7dt3TMNYUodJ2rhJjKJcikHU7FBokPAwAyi/nI2u2Jh4Zc6Xf
5UByHbwjf9dYQQNVWg/wXhVkV/fN2Y6Js9dUemnThz3uFkEwiIiYdG0dr9pLxN3A
C8K5bnkRwF6Ck0HS4KnJJ9wbog9k4jCBHH7UytT8Zmz7IkkQCwxmpt7OMLJavok+
k0uPYnYW+cePa5BRvZ8JC/35ZnmiY9T3aXfkVhv1F4DKeztzGXgryCMiMT3aZFrq
p2i6Etb+JqXN8VEwqJrE+CFe6GCJV74bqaqF2r8S23oBERgZZszio7N7qBhC1WAv
zhpjsUhuVIurRfIO/N41HAq5Zjc1rlhfhljVPXuqResXzhQkS3mWWLWJGdrB3EgM
Enjc8Ana2TB/7FkSjreIG2FG25ktuAQs5aXxyiqwINP241u9Ig+FEIKknVRQ6+8K
I5TfS6M7Y0kkEetp2UAEVrJtumxH9eS4cHRvYvPgjuZjRKny4zmVCm+p14G4FlCh
vophkJUj+peeUaBRIgUhVmtDS4MaoOyMituiUgswPoD8IZ9/BUIgy/dZKNTSHV14
sqn56naJaDPvwhJjXrqzQQIAOcKVZEEl2ez0XOyS92z9JSfG/xSFz9qpxLFWadjo
sxjZekXRoKJzipAfFhzEP8k559HmoGFnwhm3IJLbRxoxeRiAI/CYH2yQ/0B3OO6o
8wq4uHZUIn0dySvrQa07p/SRAqgs2wBo/5BUzrODRZZNUDfMc2+30gCIdF1SVlqY
lOlYMIAEVcuyio/cYAaKriFcLo/WoP9Sn+nk5lKSmzGehGWYVngScYqspJStEW0v
HT8cGgdurQ0f6beNk/rHbC9/4f93W2pQXFlRwKkY8GBnK2LGjuROLGXvAGnTLCSt
owDJYMrPLcKMe4zcvhimNDKxyOp5GTR0PxDb38PkSQUtCCenxxyuwFMsrirvZx8M
nGqrfPtTWdZC7V+GO7oQBKPuCQPg0AlVXiXPHI8SjYCinZiO9n05whOIR0hzTa+h
5A9d2j05lVoQ4me8UeCoV6HpMtwNZMZW4SjhFCbDUm5gTcDBoFhlzVy01okSnvDV
rc8DpqPQ0GTgQTA8cN/HVHTfW82iQZfHUbOHgoNPf9FcfgkY6vjdz6yGiz3clan8
c4Yj9yekWA2ekPSNBenng2UqEMQcoz/lh8kMRi4RbQRSAQE1usLJd5pHw2YvB/2B
6rhn+QysXZr+T3ANdBGLXasJ6QNL46WOL/AIx3JlREwFRiEPyuiq6xAnJ7CBIlA7
0JjrSpRk/rTqAUx2VuIcbzTeJfRDcri3fhffy+Y0Mfx/S61s/AwhzNBQ2Ravst0n
i0swU2neSa2tvCf9jRyhZpk9UTikV/lRuCluBJ1CpdNuRuVzMMCvFHQ7rKyrJZo0
ZpYT14e6KoAMaQqCAHgT9IoKevEWYgtWehSjW2e4r7MZynFnxTuan0d5sqErlYfd
aHhTXiqJdeKxblxcS1n+Y5VRfT+jlzN3TlGKlxhkEWOipQFHebc3LfDdqbMIG8kf
8LqscLq7daiB9HZRagS5hMgcIiJlAiBTlNvRF1gPhH2cWgt3g0sIIF3oRIdcgOAy
t4YCLUW4ctW1VlrMbDH0aA70SjnX8riEWVUsdlj4B+C50d8tiG+1bKRKF5jGOvCV
iL2OqRNJHEl4JXcefCiao5VJoDvopQw4BRj4Yt6HI0mB+FvMQKu//R/dOsgaSg3G
s9iD+hiepTsuDHwwTEVs017E2pa9Kzdd04hRihCqDxRxKw+pVFZusbqoXBNeGCDu
AjLjWh4kUJ1ofDaNR53SH7y+kK2wXkcYVqs+4tle7FeltQJrDYN5lhhqA9HESgFU
qnevDb3SrcGJBLwYgNbCnrvkIM/4XthfLbipf4AbzO/ggl7VJCtRMA8g4ZjG8vgj
VHylWij5BSNoqDGsLtvwAjU/1aVJTOC6O7LMA9x5Oaq5VyLPLvmgfTDMim5ur5Ae
MAmc2hLU49lFE5cEqbasaF+QRZjigF0UGw8SCAOF0ILYIZCKxeWElpPnMgAANBHh
sFwhXigWN8Sf9u+7aNzZP5BCu9V7ZZGaP2bzvnkEdysY3quYa8Z9tfsvjQ38euwC
X1JYeoM5JjWZuIyN7iub/Vrmm5SjUGGg1xW2rjAYVUIRH37Bw7czrcYzrmNktAEN
cfb1pBc+6ouyD1OdIi6DKXaAWE+T2U7eTAId/GtxexvC5awYEZPx6LCnGfsuccds
p2oJ2KwLsboiLo46zJhWmtmzMNHltiZRzUqxnop4nSRgoZkwxIX3I0hOv7urQBZt
4klgg3UyJ1EN1gIaiyaibTYou0IL36fpylZSf09Rbjuptt/8EFe7hqzzYHoNNFkw
7+ALLpywA2ZiFK7QdJ7hQRniPFIpfroBRS0TMGi18S4QFK1TwrZhCu6VDUu/HQJM
CsiIfauL2McwzEbC5jYMOORsxdMFryT/NHBu14TCT206EmBLGGbm5dC4bkEtFhmm
2UYMxCwMdRRTQyrUQl6YPxEOqOZE7SwN4B3HsDDcVWWumMWLbypZLuC21bq3leJ6
4QUHNKkbuAZ+lPrHmFEVQ4eAlr79J8CRS7eXLgp/EKxw6mG0vl6YEurtayYaTjJy
x6AdXbKQABJbRi/1H/VacBlPKCbKnSN9xsc4Tt4jZxZyqYVINrcv0HKEupZtf2OA
HXna4qZbHVY3Y3Z2JyEKziaNUC6pT9m121ZkN6v/eEBIRbZfKMmreGR2Yr4PzbKy
WjPWISrTEZAsWkyv1ZLRy9X+kossZAOaQwjfX8vZWxrpkbzj3KfUf+KWpJYjaxId
HElOXzrKzOze2+gYDNiIwwfxJGgQZ/XVzBYOeLuizXXee6D8ZK607cOWD4u5oJZw
rgFAbUkZGrIkNwv9j1IimR9b/Hp9qmtcLbmKpKLgvLLbc0mmBNGtdJCYDFvGa1nh
X9jN6c4buWie3nmbgWuRIYiWCsC9hIRioHSvoWyhhjem2Gab+fOa2GeU0KolY1xY
AS5nw8cFQp17F7F3ffLXWFFZmGokujODNhTuyKwLMVYJqTw5XFw4BUgy1+zncqoy
lY+zRCxo8tS6zZHfeYvrcfSzlL4ByOchJ7N4iDuJ0Z7ZOXVJb5JeKqeJB4YBi+yM
3kk9U/iY1p1ViYDZ+FZkCkKHMLYjrGGKG9Mtw7RKdDfxC+dka+TS6/gD6yqq9Bd5
N0Ikn7eG6y8oGunv/W7FlYzI0wAp3gSDqlHpRxO0yNfMhnueO5vqHEJt//J00Z94
lME8Ib3380AshI41jE83lnMvBkEy4wRHWGa+wpWh2i24qRo4sk1FdR5DWdG3cLcd
Vq34hb6jbNc6uUz5+3fh8kiSsk42Jq+MP1ZxDpCwD46jG2APRLMf4I477c9DJ8TU
kLl4AfXOJ/qwxqBLM0Wq8emOYOSB07kcZH8WMLuPXhc1/6bP0nOwmh6HS8r50bUg
UzBE0PQOK10e4FE0M4Q5rNXSXZ3Jvz0UIDPyhtq3EEe+Mr4eUO/wmw2FBIbj7M0J
a/uddJhwdQ5ajQhmbufNShisN8GrhM8Zz5bTHMSuRo40/V8DEQspYuel8lzAAyxO
tGoqHPfrLF5t2SpwJscwd2AQx9xL2icG3T53qQd4pK+pjosDt0RAU0oeuCkFLQZv
92iYITP2eS37SmABmwy7VYhxoLa25KQIsb7O167InNYuvt+G7vWJrQWyah777BNI
x8Z5zsvtcqzrHl4Day8xl/JbdG0nKersnjtmdmF+iRogfMsDmcSTlFLg+Fi4rfmJ
7wr6RzhQEbxAulckXqXn/j/Au26bHPOos2bfd6fgLm8oeLx8tYreJSlQWDUN5TIL
78lXIUlh8YwYHadp2cDp01F1wVkpP5PKzyjeafSVXxR6e3oCGi1ZgDD+/jL9NYl8
7ILXO2EHv/tJPr67kF9BTTMQUaXB/Nrt007AW6DU/xJVA0D0/bs+Kbhqn4SH9M0r
+hzrIWNkeOmxMUI4bm4pDTVraqm1bSRyW3tdmtn/EgOFYoY812vcwuVSBTHjju5c
Q5F9yUEx8x+jXNqigiCultfbTrQ+LapPPVEOHkP2zsymUF0xiAAp468L9+DeQn0D
8SEjUejvPjxi4EKDl0LDkhMkKAPbBRSZVOpexVeJr0thDR2xthRy4i4pYysNiind
xMK2j0n3oGweOl5x5BlGVx4EMUmCF8NLMxcO7Crh2zR3ukjbSGHEgoDtMFq5u034
NwkrRrI54T8xah4JX5oYxD1UWBiGulE6edPszNLH97iq2eJSBN2pKDTp3ljOk9on
qRpUuxTltbXp+Smi8VAo1TM+w3mKAk5JtuxXT9HxXvP8tIwdG3w+e1Helwm4esaZ
bXcKf6NiVRMKwHlCvQ6Wrvx9pF39DutQytzrWjHQlggZdIBAOyWEm15mRTaM+/r4
3lo9RKt6o1J5eNw/C+6x4jN2CdI1ngXD5Y8tTxb+MQHUSbrFHe8G6iMrJbeUpR6A
2s51eHFgqLNqsESV0b+2vHT24/5dMI89+dOSSQjJHtC/BczK47jcAIsnyMsNSdei
xi5QR6TJisFMqLye09+5RGi0gTtzipQ9Cta06BjeEziY/f94hKjmw9kbebIW9+2F
DGYg7/JjxwbHtSWOds6gKXuQpzAK6P1gSZsIUrwayozAvZmVkGbdebnSq1EZDGYL
scUmxQoWLL/nv8e/aLxDqkUnR0cmV7rccB40r6LXqIaT1Y+WgRgEEymx1EoyroZ1
hPSIK9Dqonqgw09bkR8b0LtpB+36jCy1RYbMfKW1MB6Dr/2Y4Q1WZbVSLBBCXdy5
nsUMREvMvZti/OPM7MTE9Keo2KrJxeFtRcjAM/9WOwr1tEViI9GHODADvELHnmxB
nnUihsAaUtKVuJpO+K9x7SQHcFE/mQDUbscIyLQinTzTzKPHyo6k3rWFi3NYBbMV
vQ44ZJVWEHLjqUEvAhSw3ZFxNPeHUqDry+elXC4MoeM8MhDum5Iib865oWGkl3dS
waV2Kjl7J/6+mT8d1sfJ8Yyh1loOox6JBWO0xThBqaM72dKHkNh3QlNQXSAvTMrH
nDt1YeyDIKOSVonjCP1R/qsj6jNCvbyFFIqynlKdiby/n9IdNvyh0hO5ORsg2Tss
qgzx3H6t0He1UVaDn9mhyvdgi4h7s5THAQi4XkrspRkGCSwbLhhJ34sbaWeXwxmj
/U6fH1V9jFX1Ua+EfnVdfmOfuDI55exZ9aAlecXK0eL/gATMTATJdkem+1xd9F7B
dqFnYTpQRf75AyjKYeEGCt/ivMko2rNRZK1DUFW2eZGhuH941JA4EbudakedGIZe
08G+O1L6P3ElbwD961A6b4DBFJckM1ZFyjqueaGX6LuxZ7HzAOfvAsmJYquM+foI
nZleVS17GOHHWnyWW5frYDhELxOVms757t27oM4HIcHd1aXiHMS1crrjPCIirK3i
0C2qYBOlOVi6ZPjswXkZDshQlJFMavZvwp4NZVzM0cenEjOBYgRYG4ag/mcfm69d
/pPxUjoZ6oP+NVhhweld3buRMomFHe+3JfgXyqQyKv0oJgpRbHCVa4qA0V47T1u4
l3Dx4IJPBTYGXQa1VEEMdI02uCSFu/M4lQrLlrKlCVz6IfM8KuAAfhp70+HcKzIY
2qTSJyEJcuNtrRiAMC08IWsKdfjakQ11Qei3eiqihzaDKoQ8he6//iG7IxgQGKD+
9qDhKu80TnNq0xUjW/w20PaxUWwUP0vHnBP2mLjNm+g7dqmFV1yS+jalbmjYyMqd
ps5VWn2mSTq9kKVqQS9Tzf9ANBUso2k2Tjl8IsM3euGXOuaBFddlHMmlkMAMWcYb
rk9ck4BKbvhEid8c/V4+AvynMeyJL0g+zPOohEgTiXx1uGdKeMT7+S8761spkeKq
iKU24kbcWzWNLaiUqM9h80nRH/H3SosKbvWcVz+aQ2e3uA5BjQ7N0o3tReHX9sRH
1QS3EOC621zEWZhZmOmKDlctYWjL3EzjDMDkRdt2417ZZrh2dgT5/0QtQJxVcyWf
bZoDg3LZJ5DSw5qXU243SGCObbugGJPaB7PuJzW+x79L8o9B6sj7JNaTtUO87iya
j2RQ9XKVFFGoXgzWbUQysbCaLxxV2RYR/j6qyjhuWKPPieuv5102kZACp/MInc73
lN2662BP5+LtC3B74Egd852FGKsy7BwrGia2aapRAl69Gak/5l1GqEV0LC6iTjGg
IPKEaaR627epfJn//nAW04jNlF89d3KzuBp40lmbI8lAV6Q4ypAB+3eo5Wn8tM0N
iJX3rH0J6aKM5Rx86qHOAC53dz1K65i1cGNZIpELvCAK2H1Ja2VJZcvWhXRwKa4K
BonIgm0SzZgrsp/q5O40qdousmw9ZP7ktj+1N9jIp+R7FeAcnH3phiOiSlcrkR3r
PzPmU6QqFuwjJVI62PuBjvRHviAZGQymq244nDRZOZKT+IpWKoD1o+bkquwn5YAo
Xjv4ztdLpFxqZxSEDIl2GsgBJHFuZcEw3dHRswigsr1JTJzcegE/LhR/dpefaS3/
5U0CRBX/tCjpnOmbEEIyueqVJC62y+obR0XfE84/WYSwvEAOrWomT69tf3/1zGye
rUXF8OOH16clarw8C/JtE2s+hya7MAtsVIog1/CgQQZNMMhggSb0ObWPRNcO9hOV
2OLgVe2f0J5cZzOmrV6LQrSYmnzljgxCxqDXcXAKGc8WxpoMuYPJN0X1XZDeZDj3
DP3jcmu5MnrwP9y+VlfBIYD2lOfn1j0e2Kbn1v73Rmy526tKvT8azP2irPepdI2P
3KQBTSRkFvBcVjRettroygnGBlM+0j8hulfqH+zPZuOC9Qi/u8Ii6QsLkXqwAdJW
fOG7XtiNeC12PDHBIwurAKWrGmO66BezwpiIliZWvTFv0XZM/WjKq5wcS7c9hSYb
Em9fuK2OHUJD8IusaABOpgE2qA5UMJ6xAKCR2ETfyC8b5HJ0xfNoCTSSiWyHu0L/
B1cLGm1tpO9G1lfYt5CCYEbiNJBzhImz/wgMbbgcKpgqO+fuRSPqtjNxS0LVU4BT
jtgWAGtSX/MO0dw2UJGiZhF5eJ0bB618KhV04RGurU3Y0gEUfkMTkJM7eN58RSla
h7efCNHnFlffZdbQ+34BJSQtMsqHJNfNiHT50/MDukSLXggJO+QhcEC2KovG0hIX
8eaA7Mb1FWeCuCZrAZuLWSiJSmhUWzCtPrLjCvQKTl3sMdCmNRD3H2OsSiUWuVT6
+gomH4Z+rCYSZZ/nUvP5arTXKW4ZgEJNF29RHvc/5YAxFGvkA2dYm/o9XlHoKnw6
oUpDYkZU1e1vKe4YLcrTU7+5/JO+jaEpWBphQP7vnbj28mte3fRBLGlkHCDNVVgw
dbWfkeAc3W/vf99HyvLKOxDOvduU3TgZ91zKB3nlv9hqF4u8eEsj147cYZo+FNsu
bz2BwbseemX+wpmDE8yVsNhDaHF4e0NdszrrhIifHCzLenropG8rmLAS/QBtAVfy
o3CkERex/1pOEGYvhg+9esOQc3JLZ5+32JpeIdIuCWtGlC1WCooBBs+Or3Qyni2E
TTDjCAzJs7x1f6ln0HqqbMeGmYPfaTQsV3df/cbuGZwT7BSG2kuhMoetAurerYJh
YklBB3+ML1qXWuiikTD0h/EEOJoIcMns5iW9c1/yzRV+pmQ56ANcHKe2oOo9Sv09
PvLxImcS2beOKTrxo726MtxWCZ/Xlqu7zGAZYmMTXjf3qXBEHpS1M0+KGUyqy78i
g39wplkusKgBmceQr5W7TBqa80OPVoJbrpj3XLyf5KgBfbW2hXHb7SBiIUt6HmJf
zTXtRw5RCL4h10e1ayeqOKo8EEiNXa5K3njqlc4yK9T3HRZ42X20Jz/yJQpozj0O
EPsb5uwc+vCJDqhW0CPTv34mtrfFMU+MEFY9HPCS9GEAap4NoeRRQtn5RplJTcNX
E0JFbt5SVxCpYLoo8FlrHxWwTeGXtQWCjzHEb1jqJrgjrU+7AtByAxyAgyrvdLSU
tumnTp6IOW3KhfLaKVgLjVI74P2a3BoFCzBlt+kpR5eQtvAxZTiTB85E0E/ExDIO
qRkWvCnQUfc0mFX6IQQmj0x9oM1vlH0ZCXD4tWJYFLLu4Mh6raCmIu9RFXer5fVB
pbTWMf+ldORelk/JPXUH9+tCkYMqEkfxk8lN8S4AcvkpD5NtzGePpbmo3zDAoFDd
lZXFCCJQ0SvRMxdNTNypSwoaccRDWXiXbu4QYPfeUQ/cxHCuigVPcgaWcrB8jvMM
1OE4kPCF8dJXRt2CLC3KgMk6iYLmhv+vnggUHvTBO1THBwjNO5RdbZLaoEm39u4/
4T0to34IeXcw4gs7KCrfYabW9E6Oru+rtkN9A+9+3O24fB7atcGVBFXMS/57XY3Y
i7DUE4kyRTbcAmHtCnNsLluqnFNdlW8j4Q61ewXye2j/t6ZI8q8r4kDJJaJIdWtG
ey7AUcDoR48D/hFZiC5t9hVrb24gsPybZtzViMlEJNS/k5ZqUYZUGj/dO9svta9f
ckGPnXc8DadH+9D5I+iWTejrIAenOYVlYMa7jfU2j9pYApRRdbCF84cbrChNQoM2
Kt4UBcUv70lrAvqUH76cI6I/dn6Y/7MP7AfXIVF8cwoep8x5xn7dSEDUqkCkFiv3
Pn/7VraL3l6yeVlRU0c/d9cvnXh7twg/CGNP3EkeSWxKxW+nCTcZVtr4szZ7ysd/
vpNMMO0tgbjvFbScTEUXsl0ujbwGcmSuFViIsSrBTECn+wY82LU0jPPGjjNPNn4e
Eq2sfGjjzFGAkN5MI1otA7ZHwmG/y+0utyHDNM5ecO7TdFICtn10YP84XjOIUfY+
khhD0BCplkmpXXZYayvu8tHCAzIzfxnq8isq9Ookh4N5PTcpKnjmkqmVkPRhogtH
Bs6RB3u8pte2whaY/JYy6XPEcz96Ui1YuOAOR1IRWALHEPMkDQCEw6+CP1Yb4Viv
p17We6/nmKx8o0YJNOPoemJSyu/BTvLALO9ETb9/u4AGYXmyu26bldW6omwhVtzV
nd8SAEnHJY4AjORnvKho9q6QAQYF70MkL0PhcNTg908R+zxwrFvh8aAfgWnsFm3Q
guuw2pKosa85s/c6IDFXRbuCps/iH9P0fB9EZWAEbzFKhX+Zj7kIi2v7wKA806qw
RgaFbFgYIWJ5tWUYXE5qn7PhTtkvRcz0kJ/trAQIJfOSyAlyccJvtcPTzqzrhMSh
DXXuHxlenytagjrF9gLbr0Dz5soaVcpbNW9m6rI6AW+as+bPh+h4XqPtboftqIzG
XJkmnMOo23SrBVcmgtod/C4MsOkZuCkVZTgdrR239ZANphN8p+FlEHMQJAxpI9IB
OBGz9yDG+WO4fR1/e6KT4VpgRXOwsf3zcK60I1jno7kX6nixoqPVLDYnhcGOqlLH
nEurwEeCSqtK2vUxC6RPjPHIob1khcONUKT9/ZusWjFzVuE0e3vbyUdcqex+VE2h
KMpFOZ70gIQ8fqHZSEJ7uwMgY5pF2tADuC0jVy35PYbN9hXG92oFTO/b5kSVDoSS
r3sbrBKFu0U3zKf1mOwlEPgeZ980Cttv0rbYD/qNNBihg2ULYWiIYT8QuMvE0PLQ
9cstTf8Qs7cJ8ud87/uBSk06RDK6eF/F46oC9h/5WkDE/3gnNaWju8bzevIxzszD
uHgUaG48r4mOY+i12STbUdw9YDmUPNygwOOSRTcZP2we+jXWBXK13hQsQf10F4kw
DoB66Tixbc0DKbL9Ed0LY4D5t6hSui+zZXImWHvPzuMz9ysUZe468Qsk9hMypmk7
xWJE03wUtR/jA8XWyDtvZ5wYeloOIosJ6u4DiBiX3bb72akjB8SpgXG7WJBmBEGu
l2TsdTpz1Xg35Lmvve7lStWiFOqwz+Zpn7NNcQ1vRzfFi/jjd8F6vVUMQ6LGYrNw
xPVpaWtK2j2WtUrgVcQcqaByol5I1zgb7zjq00TFLaF2bO5PMGWvSzV5iSJ5CsCq
jiWN8WJGchrsM6oKDY/CC5FUdboPJD/f+T8jilBr77lDFFOHTQMupRNxg1hbZjiG
c7y9ETJJjW+Tnakguj0c+WTiOdDFyexp+zZwczcnbfRzN+0zxDoH3PJgOA8sryLf
LTKhXfP2Zkl2Q5w4aZR9TCJo7hn5E/E8dervK86o3+eyN8X4PWH+0xmclk4JP9x5
3QZAHaWFq0tjnza4ofBYIVx4cZ38FOuhx+M4DydXn1tuk28pmP39jwnD4YaGlLUa
DY4ATvTV+Gp4HoHlNk61NQvA1qmcCj5wc4csOpUIRivCrirqKw1LUUzGtBKL/ofn
p51H+mPNJH3ewDWPuvguFxgXWKDXBtnliQWxeILvreu01DeNZWnVKjn9nc1czU87
5GHANUPy7gudZLxKXZPDZzwkztpZ7d9LZ7L4zVRGoszWA+klja5KoLMQrSZovOev
ibVu6+EPXvUysfZ9RmSbJTHk//OrsVWZOkxt67UCROKXAi26vMb3ROb6O/ZfZddo
u8yJ586kMDG/acE9lTWNn1gGDeFJs9AN4k8Qq6vyWoSxhWOGPy6/0no/LPhbjaik
ki0itHEjq0ETdHBoud/2Mp34o7mBHwIQSmy8RoExgEGRlew9qU4eiBYlD/muSWUj
UfyvDzAvFRLcdNFQqsPDBiyE/P1bj/EXvVKwlWQdH3x1C+jxGDsMaIsEox1OuxXA
8emOY7vek319cEYXNT7vny7bYgjIX0cd8CRdZpqT00eQv9p0ENNo103Tdo47DZc7
9yKPiEQiKi9B+VgyFuafPue1q58G+ZURYQq1FsK0ZYSzDZ+FndGSiRDClJdgQYS0
3y/E3bgV2ME44T3JJIwioxeYw3PvgsoiYjsRGzdXlimAguvc9FrszzwIYmBOErTn
oVICuTn0CMroHVo23R2TocwG2gg6GiEaFfK7TMtFrfmn/s71wIsHdZe+KFBUhwYd
uvCWLg377LpHVEJv3STSVTSHrDYSuY3iqzbtNuRCJZs7/YAXtnK570m5dJNOiJF8
/mu2RDExBT4gd0vGXSk60WKt5o2BGDcEIfsGQbyIYQCg2Rnu9lqFZ0v3ac2UBWV9
QlwgiJaqIvZqjFgndCl8n7gcPhUoXvgXrDEMHAfwaM2yc8je2orrJDf6VEAWe2SY
wmhTTL9erBWGaapsye9L15MMnZ4dB6t2637Z1EZlPpPSqpTR8PYfQgkFtGOULS73
JdycEeUX/SocXiv80r2OnbudV5IwR7RXfpWFqq0IL3PXIdTNCWuXAzOg2a2JvLlK
jyXKUgKVdsLpI+m2C54smVfd3pmt9OI2KiHaiY/Q8zwnYm1GhjNxOqbqY4bdnCeL
qvH9WDoRIdmIGac0O2XalWPbtLc/r2GOl+bVyK/ViVPZX7psfr7KK8qfMow3bOse
UghVv1eZ4DptbcQBspdAhkr36/2NPkslh+EYW0q4qiP8/XupwFjp5mTGtSJ80SMm
+IhAm+EEX8fqKV+PALbfeFIyfEZg9eMHaeZRUQ58/OFOOYMJDFOINjvyWrDKQEPt
dXXT3jKEum2sGf1fv2gPA24DAeTtn2uz887j7e/2eoOtKAiyzR8Ith9zN9O+UhHQ
B7/OFPr/h6bUGmOMKmm2bXupFhiu6E0YfkyTQvCEz6XdE/wfDJLAfpvckxMyu8uo
ARhO4kMSt47xFLQ70wXmuPN3WGXNX3h2jNoNsWhrI5oA+J7C6PqIAP8sVACU5/w5
/5H0Kn+d/+Y+bB7AXKT+Ih2BX/mUe5kikUNDp8/0MkwSDz+mia6/IpITd6H9TYjh
QtPoGRv/Br9YwC3aiE8KnwKBHqAn/Y8TrMQPYtGOSSjhsvqqiBjYFS2dlyBc+s9W
GDXtYZrl7SSRYL7D5pNFlFJWIsN61RPjJMfQxa1ce8bryspei/mmi8pFQGSxGpSZ
oWS+NVKyeFLsdadAQ+JPjP7t6eCF+qcU5/SK3XxwU8zYhmEVPg4+gDnxUx3R2gtR
wZME6OJQKM38MzNX6K8dzhGbYxvJnvVgiwXnDC7IHcpicVgdB+YXhheKOyXpdEUj
7P8gSfPJ6pMGaF/gPdI+1gzenIMw468oUfySaGbhlfig+zzxfeCm16x8qsNF+iOj
g8MvHcWOYAQoBvGDP7EgpsVtB/qGRqL5n+ZhWdd7xQTk9K3jRCWddE55wNhvs490
o/9kLVr5h/82FUKGyDe3/eUSDS9jGQapkKjsyQ7J7/Loj/DyD+vDy/T9bB2eUIHD
Ab/UF032X0bqGV5rf0wm3t1PkVmgJ2aANSzfs1/FNe7z/SQ9yI2R2Fu5ZRq4KcQj
iY7pfQw3nkoICBrPADDaIva8YfZCO06dzZah+zFeNGg73o9tyM6xEhc4bh8z5fSE
8k93wSHIcQQg/V2yG2JzHbPXB7U2VeXfcfUSD7HexdI+mQ3butI99UYOWYyQuKo4
pA4DhnPN1BzuhQBUsAoheeS47j7edKVgO9FysCLV/6F4yQ903b71HWUo9cPAQc/Z
ldNG/F9ef3JloEYwvXwku+EgyEejE558WpnMkHBhFj/HaMtAQ+hjzElzyJReQrkV
QbHYAHCuhYi6K27Fk09Ab4IZB4YHAjKhqgOR1LOpv4qj9ovwBlsAYhkzfGK+gtzG
grRfYCeYmfzyuSlJk0xKY6/TIAR9+5yKZSzd7HgISIm+wIIaf2Yxk6AwVKrN0gLn
CHDRlJN3wP0oE5fSOgeLOjx97NwQjGrfjOHZvqbs2Amyz/v7UBMgff+kbp2hMikX
uJ3M7LpnZJQW4uoZA175NzKvyJzgWXOQwL5pxwoMy3aOaVDBquiP9NmIzNQRnJ+M
685qf7LjiCXbH47S9yqBDpcd3aRi0/JvsWTihbCr1lwtJ7JZB0i9sPKn8GaGSZew
fklERUKTMMFWCcOa2s9iF8Y571vmKXW83ObNi2pNpFAsulX941bhAxNRnN4AuzS+
PFMD761PucS3hqd/8ZzvPYkE086eJU+D8uHdhPYx/YR82XL5jHxq6uNcYiQFxRq7
7fJUtFJZfIKwyww34aYDRo2WIP7n1py5jUyK2cjM/Za6Vo/eYtM27nOjibxlTKIB
yepbp0F66BJGziq6cwk2dtsDz+TMvNIxwPZx6F7R7LuKoDhRfKUX6up9N8ZcQZ4W
GuRmMRrB+omTfhk/6OFvcijJLHpKCCdREpk+xx/L2orcqqzyqNL2tGzZdrINsNUh
aY9fYmdJo1Aj4zzlmFv2xi0k3sQKA1C+uoQLxclCUsb19YJ4U5oMTcpdZjfvFoA2
FMzW3yXlPe0uVCx9hwqgcN7PKXuTbct8p0OtWYMKDTyRqKeggx+BClbOMoJajoiH
X878ktnXOfgj9ixQGRF53RpOs/U5dlvVpzkTrqj6l23f03bEIhD5PJsR51CPfmZv
kDlrJe5NDrGVqj7ECuZoXusxEQWWuAOu1Yj4RiEc1KpXD7O3EfX3owo0CG87bi3/
dQwV+RxRt0lGVDmlEDpq2QLLI/hH+2k3gAIpTcJWitZcHpEoK/kjDPTKttAaoDi0
rjL96SlfQniRVsi1CLjUaXhQTD/cGml91q2c2ugOoXNdHs1hCFRLHfwwkrBQ1sbC
mknhs865Om2wezZZDncBjfcgQSOFaf3eA51DpHPBOiILeqjczrad18MkaSye/ngn
1pxkSRrcf84idiHHXNYsEmTvQnrB0x+9UU2fzOiscC2iUhr7jcsmBbMeq1IsreeJ
Y7Qu3WHPTk3+zuTR7KJdZHXty+kcmbJwidRKg9Q8taTGBVbMmd04j69Y/YQZ6nEE
RVNg+6W5uPdvrPFvk2Zk3e1qpkodLJzO/ZbUrjboghua6MWbSPp9NdA/YYM7Pd1E
gApw64E2WlaRrV1svprUvqFWDzi5uMUuiaKx58PyDOw6d0dho3ZDfVTHVdgJpGkZ
dRRz+VCTvByLDhgns/TwuAXOlT6FIiL+20ExASvi2asM72oE9YTFkfcMlkAcMMak
5HOj7QdOAFMKCju0rjhTQishuEawiXHhXLs+ejvSOy3xCs3dyumI0vL/o36WYpQV
OGFhU/lN2I0gbGdoClUuxoU921v7a/XrFbS76R2m3Ygy56Oa+l/ePlYZzG4t+Wow
cInNVBf7VmnyUjHcjmDbqO7O2lrrnneBXQEg/HhBimypSAtD5pFeouqVVoxk4vGE
PIZBUYwokbTWrz64fe03SxojfhbMHSV2jiRdZGelLzU2uVyP6WgM5XBVc3yxD+Ov
+WNOxDvURXkEVal/THMiVK7NAkaM4kGAEXYUmmeVB+axSXOju9r7/8SN+byRogOv
S1FL4HOhg0vWiFdjytHd8p8Etvjfw0oRPavsvKWc4ENSHcslJWDYQgwBnGKI/UDJ
qvpZVFiOBYlJvOfgDhrlv8Tl84MDSu0187O4gw0nXIFPzDYdiHqZHs9epZg9Tozu
Yf3RocR+KAsXW7XHlVWp9kE08ZCOtozXParQED2kq+s4nTyEABV29GtCOV6jJn+a
M3tIHOqk66PBd/P/+z7oUbxVDSrsflZjb9H3621rdmVfg+6bIJffCs9H1syyo91G
3foYd79xYSLxLbEXeKsJspErpCHIQ942E4URE52WfDP9YbJQ5S0zDJJmrS2Vda9+
HFwcd4uMY5Db4sMNVAF0uZz52IjN5GropgBVBq1q9vE0uo7E6qlWSeAtM94u4gx8
a6KtTrQAMK3A4qnOCfoqeekkvv7zrF24mkmHIOUlgih5OKoZjGYcu9dqj6yNwkzA
6zxTLlfnHrabjPHofjqiID3G3FXsV6coWizX4LdJegsZGDKi8OzIwj9lrERJTWtd
CWs/reFj6qklK14xoo+3O0d9e738QIVEO5r8WSQ1YEDEHhl+9Ir7CuSzQut4mcXT
ZQ6FyyYNg6gpA92fsxlteC/I/Dceyp6kaGIwwyDZzU0h8I4WGr2G995dVnotq6Hp
GUKa8P/nJBfDealp3K4JlyXfgBdjG/ZgHyg4+YxyhLjfRtawKtGgmuvD7QnQrZ6F
u/M6Lnm9xyJtDLerTQCI2mh5Q/CBhV5m6jHjUXo7MJHM7XYDWq87UlH3mCJKKyfL
jVotohltl0VFx7aBMYXgtuUtEt3ZvlhUtnbvUAe4hLGu7c2a10Iia74ds5A7W+Dq
qu3CBnge8Xw27pPCzCTAfP7Is9GE/anGqmGz3YAWLUPIapb8rAo26E5N62KBMSHz
LeAdXw2q8nw6B8j4g+0hRBr7Voj7FCKazN68XxDHQa1yE0FreKIZmFoOR1ppUrF3
1DJwQcwbPLXSrt51K7ifUwIhHr0xsD7bTHETkfNyuAzvEIenZJDpXnjE5i9eKie9
hHyi6QDr0HQZTOtvaJ2Oz5GBdsjFTumwPFNM/gJTAXRdchCjT4oRcGDZWcJV0v+I
nwkdPJMD/vYGOIfFYMf+AksN9v4DGNqq71Apj46EidaGkOdNLFmoimslGgqxyt6/
WLfAonkGOD80ikW7klCPDaEDgzwqlB2yBpDYNCIXGWp529JfFWEjpQ/CJEnqpjhU
t2Lx9qRYOFzh2IInbxy6LRIC3MruwfLycYiiTR2a5jzm5mHB0+QuviDvfmI6ye5a
FIPfWqvJe/V6PP533GuERWezGBs4u7oSoPlzywJ2weRmnRvFdFh94NM9jv4LIUsO
KqRFGR0VtCTreBy/DE9MfAtUmjOFlvlIrGbK3DN7BZ7paznBp768vet+kIobCMSI
KjQeMeeulThUWl/wGQxtuCY8DrL69CBh85pe+TbCvk3NUS76TlmUn4Ahx5iSCwtt
kHVYqM9m/8R/hMBggpIRmLeYxyBTWk+Cp1zXukZCOXvNSxtL5377OMuK+7u34g6z
G0l4/xh16yVFhGEyO4T96PHJdKfcwq64jzvK5EUfc3cgn27RNW3tasXlQfOHMuca
87BNQFr4fu6u6IKccveji9SilAlXypj0XF8qsB7QDB2jUkclN++oEc18JI+QqoyQ
U6NkGTnetDbsnxgEtFhst7+4m/U/pvZ1hdgzO7ym6Pc0yY0iwwj9elf0IU9dK7QL
II2ncDa/vfFhj/rOZtN5ElOKWdv21sW5uKubY2CziisD7mEMSVe4qdoMGVLSFPcm
HM30i12LhZXH2GO8f7gndc4127GzLugSKmt509FuKscIVekYT9rig29xAZ5HzHl4
2YWX3dL5ZoRiGOnuqqxbCjQ4GsXagHCoTXWFoMmUxwZ0+UinfDrt4vDavYkbpOmV
XD31TZsHoi2yn+UWADkUXiHqkpaNc98nk/1rHSMuVv1H2m2pRcCcP3R/Sbe7AaBW
LoacKlZ9DA6eQ5kzI2zWXvNiTwele9+3QoR5K+dGK01jsj94pAxQW7ge1yP+me00
QsHvuu3ZMLTHD5h4O459I9K3S0Yj357uDWzQcJoqZg1vFSlUvPn6fq0oqdvMKoXU
MlczuymLt3tr1xoFOeN38a7oP+i9vmMUuB9lXtImTl5iQl9yKM3M0Stk408DU2DB
iG2Zcd+t217bzC8FSoaxJEXCsmzJcSUz2R/I+tyBHlMkHiZ/bRNJeACiUFm/qjii
4u7Ek2947JgAIDdAfdDa1GvBAnmEES3XnbobbBOJMG9xgV2Ei13SpkkjP7r7QF0F
aGybebpTKfqCrkszd9VCi5iB8/h49yCeDzb9+JAfOzZVkTYzqh45hJiQIfyHT/h5
7Iy2WGzxyvjgEoHK0SwYJKyBDhSXHXwIgaG0QIGdx9BJr6tfvDKLm2jJCzqDMQS+
UtTd3quCPSjERREdYvohaA5r/pxXKZRIDxYZU8nQ//Kbek7wMfBFx8BZt2CTI5K3
krgqu/vy3xTRx0i5nPQFXJK88URPhcteDK9/SW9EvK+YWWL/2Efkzfy3amiMKZrR
86FarxlqsumDBL9Jna0juZAqubND4wF/k6bzgXD9DPHbvai/nFNzl1er/zSy/phY
GF8lURg0TIXuONifwzF4pepWBUsTBoxsKnxRg3E3DKWhlrBpKhM7J36g+pOwZZwp
LjmZg18uKFhA7B31oVJifgU9NWWnc+MTPSPYul0Jg4YCk9PwMfhFFYrAFk5e4EHO
7pfxhb9M4skN40I/V0drCEBkvxYn4u0ETKATr2ld0wUbFzFmQrTEF5A9d+UVI1CV
9Gpeo1pbZJl9cYFmMcNDEpus4rYXyhOOpLm0XgNYjyFooq0lsglRLtP/JNaZQHY6
aZI/rG3QsOu4hwiTFVKdjHgZDXo7H9W4H3WFqxSwLNCVwqwlYbs2hkHTEz4hI/a/
Hs1HR/QJWAhDS+H0M1G1IXh0uOuDMF4LJdrxSDqFwgKpD5/857ehb8fsgXIrDWaL
AH0yZFstu2mlBFU9ElfAaZmq4Q9rnuRfr9CV+lx+eS7W1a0iDBFuQbxCPenMQZof
cVHFWsehcOCdrMDatKnQXFlM+4Xgv9lb/iw9Wb5CIUOQf9Aiw6024nqBc0rNvEWF
InKblLcWKBSNqpH1OSGZpRDCS51Egc+qyL4nz5UqyIPPDJ85nJZguWC/HiACqE/v
AJHpgMfP+o32MX3Ehq923QL2RiX9pFF3X+XrkT/zTCHwhIstHt+ZJTb9n2ZGmvBH
5lPkUPNs6krC7ej6Oltgy2sjDpeNWFIk1RRMv8+9yzqW1x1OB3qjxTdQoJyMfDH2
E7QK5swlMPrCTMxafR4Qx7Ip/iwDOPzFtzj1PEcOR0dMGrdiGlRzFIQgxZ9nOyOw
l/JF+VHGCb5jq00uSRZiXlA8Pe+S6EP979pdhqB5a+7AqYjyroLTy2P/bhFnAUI6
v0vtf9yFCfGtnH4YbD6ovVM+znsTNbvhizjUrJuB57F0agCn5L5eip6gIqZCOUZM
xaBunfAFl5/ZZHKqEFlfrdRJc0HKITIVo71iZovtGwbe5gZZ5u59fJVs5LmoxynZ
PutLv/56sxE2bmZgtCMPYf+xVEb6/ZKB+qRufIO1gbXuDtVWaY8FS8hZkLE2tjSt
vip8SvcTpv7JtyUeTA8hqZFDgKECRENkZWPYR8fOf7NgjI6MeVMPQ68EI9bSyuCm
uhbKnkTaQxl/q+tVPZUHGeYQ8/eTwFHMr2BaQVX7Y10GLYWNgY8h63p8bTFjRGL0
XCtPdWdJ6x0rpxk4lgywDS4+38cFuS8aY8o0fUkCJQnsaevpnRkdLgPD6+upd4p4
CA3T22YDY6A3/Jb0JpvONHfIXSQFLKkXwsSODEka2CkmrbXRC1wamJHe7dafdUn6
2i/Z1C/BlCpkDjqq01D+vD/YZJGpKXDwKH0Y9K4NegIFe1uYPqM6yMBBCXHrlcRO
yuCX/tTEHBAMhfBDIqjxrtvDvTWAsSa5WpmyNmaA3aB9N0zYGJWIHTbHMidMBeuK
7UULDDeFdY1GtjPwRszY7Y7xEoCYM1HkhEV3sEX1xY3xwdDkOxUHOfLb+ZcxKFBE
/FK3H/wGLyIOJpWsBqU3RNncfd3tOtQj8cnwTDzrSX4nw1fKpSmuKuf88jaAM3aL
meM4l1/uH0fzcaizxyux+dN4S9GfXfXGpAJEsVsmsjZuizNekp+saPbIaxLk4fOp
x66HRNR950s1JN16fJYdX++A0lI2wfMWYJtmx0gE7FbOdntChNqA9iczAd8PGBRI
Dj2DF+R+T4DdF2J0WfbM35WkV5xfXtFgQeGRpmdyqEv/K5D/igdQdYHpdslfpPfC
JpQrOZQzx2rXPvkgOrca8DtCSTA5oy5Zuxz+wHZvIpk55tVl/C6Si/XQTwNwX6L7
y7DHFaHzLPvpbwyl9FUIuXMOzKppPoPefFzb1UDhpfTYmqZOLoSomapwK9GIc4OZ
qxDiEolZ9ygf36MJUj4FyA8CldTjn1y7OgdfmS+7bjHdwn0TiXpZ3pw0FePvXuPD
sKFD6QBwaUlzxusY8b1pweppdO2QsPivsvnsmH59EPKeSZmYRi2wZQzdQK6+i4Jc
AknTugUh5JVqNAx+X7LYJqTvgdHrQfA5rCAQawrCbXkV+wuazXn25xM6b2CaDRTF
uKcKiUOcbxvSG20WFUE7/6PGJb8LsQ5NGE204VSPq96HjfyureBNg64A4nz2FESj
IOmOoDAD1IMdIasM1mIJ8as3vG4QFbdUH0X4AajaapcLXtApUBVG1RMMj+pyOiwN
JOC/qKN5M56iw6KHXx86NL+fZ9IYFnWNZApKKpDdodqcekzX9dqPTIcyPnldv5RO
A3CkKFzlV5/0wbbJPrxlV8zJxFxeriLwc5zSfM+QmROxadumwZbi7vWNDJxxzmhO
4V2N5xh5CaFHiNLAJT+BYPuPeD7ESTNFYT1Juy48DHQ1/gRZM3JyM1tExnbGoUf1
v0fDhBBtG9qpY4EbYtYP+RVwjDCIvOYfZdLBydUgNuIgXyYRk7pgtTXF9jBwoIHR
XCLVQMswOT5sdKIK0U9ZLaMEOspB96F5DNgQ45o7mi+qjXSh63DkpChu1fKYiy7w
w6Rz10R6H60ybKcunWsS7NXJlBrcCyz7UyGksNnWVSmu/NdFBllynyI/WEfSZOu5
evhVcXh8GgXKmhXqF7MPmZdreG3jK0hzn+PWA4nnDhk8j3UDgytQZVhyf+cpEtlv
dHxmNUMd8tH8KvA/VysB8iLPaW5VYR/WP+azkGAC5U6L6efk8FUxxiD7LNTRI/vh
wqbqN0YxeCx8xsM8z1iWRIFvs/z2NEthvFQZr1lAxfZMRE8LY40/G1ay/rZssb/D
qgakUR1eCrVEK8sAUrmuMfs7iI5Wov9GBh3xKQbcw+4/5+XpfCsbPsE23dauMxTI
EtKvA449dOpFKR1J6LrAv0FG6cPar2aO8/rk0BMnd0fKFjHHyN724eu5hqYuvyI1
Q/Hyy8bXSJw8WeLfyWM6vwu7oPr50OKhYOYzt3uPADgg7FzyDQRWiyAGhlBtDkCH
TbWnlhYJgAXN9TPf1ABipJ7wj/qqqzxdHgc2wSPY2LLqy39j9yg++ALINu6Nq1a0
iKCNsyvOc45smAoT/l79yfOcyK3NALYLWKWGlRthEU3Yuuv0PgUkKu2HWLIgwjfr
Yb7AcMQgN5maPKEIqQUsY58c3yFE3KxlNwulHw0J7C4gi5GJdKJan0qxdbVyOfpr
hsdTUxiG293Z7YJALlqdw1ES6KyGkb1j52Y0ui96yGw5OYD+emDOxoZlsR2o0B55
lujLjdNkJFWnBmGpznYh8cry90YkUjR7OCPKhrxXoJnIoiywHq9S3RhUlhUN4FH+
aZ0RN8jUtSYA75yZq9TnQ+EaX0ndaSjXQPfvuTHrCVqyM2XOd3hI/uLg/Vt1AX7S
Sxg1llJ/Br1HwqfzUIiexKcKI28pYdFKgsngTs8wxG+XLe7yE0884zlkeKc9rpga
zUAttr31AWHxOyX+GXNKxBava8X37EglB5397k+WCRG/unra0aVMOWUxL0x1OUg1
c/FLUXX1fYvDmRZzqM9bQbD+vwH5jpW9I67uVykCMF8av+hTJCDw+IfINouCakTT
v8daA+Bx4M1c4Q6k3XfOFF7xiPiWSXfqiS4uPI1swBpt5iRl5dI3rXPLDqH/Xriq
BYzqN5TP5DYQPnu/c51Gld7tGKuVDcsABkHuVOmB4bEdXf0Tuu7888j8c7SedkWq
Fzx3UZ2HhzY/MXybtGewUZQRSnaIbR/SSKZR6eZX+y5K3FAuInupkXbkp0PVBfGK
Jp3P0wDDKA3UePBNo73HuqP+1AESUgjIgFZJ3nC0PON5rRak3Pv4AmwMRsGI5MOv
RqKha6kXHZl9BbeJ5zQC98etnp8HWXhyXAkxxlNMcDZNXBGsMguEXnooF2duPOpz
Q+R80mTSuq66XlPNaAPNUF3u1Wu+o9GbyNI/MA6BhdDU5x5fLnOUX+S6wK3vsfqn
R5GMbap9spDFoTAhWB9u/T4/IeQvJOtXT7LQVUS6VXiObKpLMehVnQhqxe6dFn0R
kMUBe/34jyUB7UsY/ykmbUaSjpQ4UjHH8YaPoLqC33AQiBzEguSOW+uH9puFSIu5
cFPayiVHREP2coz0GoGsBdbZf9CFqtW+Dha93Q242OBDSxYCWBJlDb9uFvhoQWNS
30VmxhM90oqRf9yphZBU8kVd7A+ovFF80pqRZ/MX97dWywP+ebAI8uluY/pW7TS6
10eLXtde/Rb/X8w6CBLiJt/mr0mOa0tUHzxEy9LYZ5RReWkomr1w+KCnvlM+Q7xZ
ai+FVSRKdBDqduydVT4UQb6q4ZfZ/CaIhvWxZKl0CqzxuN67/muBcyOLb4opYYpM
9/Anob7V9V6dCXCZ4UoQKeN4xgnXhIRGsGVGzTqsB6ZrxOjN9kE78+o4BbWzUExA
O5vxwVZyd6Ti7izfC6jrj+uu47A5IgbN5MW50VqKIYFsRE3VaMM/7rd6qxTlEfD9
wDUCuPlRviuiPYwEi6I+X5hyguzus3uQ0gNFn9AjGU25ydZd/aiPbnVWPGuT9MkB
Xn8ZDBYZvbO4KdE8+YKxE1atPXT0VTdGeFS7p11D2QdujFtvYK+gfLMNsrylYBcp
EL7AvCcRS20XCkgwYIOQSPO4PVHytGVF+gl/1qXDSTFxg2NI5uWOOYrW+eZvR7qO
1D9h3y0DmHQUA0WFUhMEF8OTI6/zbBiC2kvBP60UwHsKzfysql0AVD9opfdeWGsu
N6Alt36/WVdmhZfUdBnjthewC+9511T+qOgx4swjhbTxAyy+8raWfDumrUu0QI91
ol80PCAcpRzEvSW2NXgVkCELLfEV21gNXP7d+gKVdzFc8IG4WeGFO4DhL7qziIOQ
VgYaTeNUgtwvN2iYoYJ6yrlCyn5xemcjwq0/SxissMneXTGwwIwyIX+Levl69Jir
6Wl71M5xG5Jp+KW0WuDlt0Ik20UBTOgBTM1ijfenbbbf5L2VEYBv2CCmyRJ5g8Qd
Fo/+SYdZ3vtiW/n9qtOYgEktDk883a9NFy3ptcjknH652HX8P7YbxHf5TKsQEe9I
4U72FumxpwPVG1Bfcva31wcLt4FJmr5d+dCILp44thIYfpqXCnzGFPg3ump9Eq+v
HycVZckWVzD4lLDW2wdk4+cuKUPI4Bpj8MvumBzIwyWFXorjvjCzCATDHhi0y0Fd
qILtzOjt5n57o9gyw90W3xznpGL2aRZcK4vVPkMEObb2yiGKaCqYuYsSMNvONUhH
89+gYszjYCgK7yFvuKZGE77U1xJ9/8LI1NP1ETCiCfGvWuqndYjBbAvGqW660OaH
LtiUeSwqI7BK1HnQ/Cl1z9lEu6XSoiOay1vhXJ/aHuoM9Pf7CiIP8702LSPGSO7X
lyGggxvr2X3GWFiDrny97tPiJ75bt8kE+Xc/47rdfObBmLmho8pH27WPp4Qz8cxm
OLfUH1rqSYgFl4GkzE2w9n+KYK78gPMQ4sXNslEiJghOwkdDtTkdFwqlOiE5yYP/
c3WxsHNiljhdf4Z/Llxj5DaM7jH1k0rr0p6iAffVwfofoayaS59LCF0MaBTMXDD7
igsJ1IUj3FboOe4AR8QYo6cnoPpsKblZSOAMJZjwNOxSzEQYDXjDo9JEU97CPchJ
Z+olNl8QWPTdIJhn+OCAwL23NI+d84M2cK3Ts9Mgq/jxR/IW6DtzXcFDFPhxYorp
YpaxcP6jTRuu1GBF4VIFYVyY0jfVfalg3B5Egvk8ii8fZQfdqhcFmGynLYGGOA//
U67s+QsEsjCc5+FAwgd2mShdmh5eQ3Z321/E7Wjsj81pc/gNdHBEn5G7bh29cq8w
I6NY2ICGKkZA5lhzWLLn8rZoQ+izFQTllxBITkWJvEVUXsLsPXaQ1nKaeAIIkgrl
2qOY6dwNnqITdd66OZ6VSgpz4WpZYHszGugk5cYl/kBy0YpM+YHFa0CRW5qvQpvd
PynKdNCcWvRtsXgd8rKrciicHLbsO20UrhcKsQoGOIo9+GXSM+U2cBWm8Evxhqgv
+4wXe+77jp7RMxctBMd862AXst8IuieJWYU4l/JUobRpIyoPH3AwQyvkCWIPkGIt
kNMcUwXCWbfsNJRTpKqnoCgVMZI10pwMBeeqC290I7/onqBdsS5K7dxdztE7+0ib
NwNtrmBw5+m+PExmAgBaMuy0H5yKEMjnEywsIalKpdHL5ri1mD+LWSGr3yxdQdmw
TQ6iT5HsJlvdfAfXrzP3B7y6NUoQBvEaoi5jkwbTTTp6oavZIRMyt87YExPPM8Iq
BZGbqZRWLLArwNNlFG4Y3WeF+ZRvstF+KgnzD6Coet1mjH0WuxJRYiwRf5Lw/q5N
UY3fcvYWl54fioUTe27I2GkGg5SCwDrBsp2rZqPRYXIpYpTr+3ChMH1FxCL7hVVu
g73Sz1GhP74rHyeZZMsS0i+RFTSyhg+wa002QFxEEaZNo8peQBjYqUbWe7CY6Lk3
02fQYCt9m6NRKHqJLDuv49iAFxeZ5cpkzbQuiqaYLkC0qsTzkvFRHmZ41hcSmxoa
c2wHHOtzobEUoc04i3Na6orUA4ZFcJOppmNKbtuKhKpSKuT0d+UBPtlfVr+6WbiV
+hA5BXVpmdSZeBY03tkzYNxrRppYZ9PuQ9AJZTHfk+npXIpCBusnAgGaj568meQh
ZyVpSGUsNpyG6Dg6xcFviaq+zcltElJfiyOX1Kvps0eTLlCGwEI/cjNUHoYzbF5i
Q8l6X7+0IvMDvtBRRy9/uVOAwq3y9nleJVDmCxu8RowbteOS3BGHHdpYG4/TW7mP
/eedY9DzT4MCXMO+BHXP1pNn/5qB8jNEGaYi//jFdKeippriDixjRuWBDYKW95px
kcCM4gsj1oQo9o0SyZPwmv8hkkH8/FT7QC5z4OTRZtkorRVW1uYFBmuOIJy0Vg1S
xSNXRZd4NBSo1IQR7xi8qOFMacWSjoS09VgNtH001QpRffsABIjAiIVZq1xyUnPd
hux/dLGSp+e2P4OBedsJaolR7SzV0iZm0ixEasEdrSiyQgdBn17pM20FZe+ZGccb
eQTYhHW2RbiAtfrNQH6LeRyZoGCUumUGxiTTamJSXEiEgMmN1vqo0sB3NtKUHq2z
OU5dWji+7HbYiLGHCkBykfHPJTTQeoWHeuYamREdrEWYb+PrUR46jOMlhy/DNYnp
pLo9R/DUwZBeMS8aspmvHTxcbaY7N1oZ+3w31j97gIOMML1SqsyztOU3ihdq5uUJ
qrOEPINk0NK4cD37uXjPSIVmxYmhqS/isdNgV4eIoLmt/E9TvOnNuKt7yYhzNgfI
dXHjAqaAG1Jk408DqwwPwpHRYxoCsM2G80j1bU69C1ivj3PJsh45T8ImVynOx+XY
2/HDD71hjtQR5lardJkMts6J++rk6sgsTVeJxtVLzTaYFnBQKs6hxW7CHieUfefD
txvbjGGHUwogc0JWljc75CljFst+yPopiBn1AT2AMJNuuuyluD9zQF0Q7eq4uFws
BLio0GYX+ojpMUzH7oD8/ak51o53aOAAsNKxfhDou4HKavv0XCE2uHfijlQhTMT6
aNYRxxZsykBRIFgVsTUuWMAQORTRlgQeSVun5kTX0lw3otlwgF/A38nPk+kpXotZ
hGZYyuiwdJOHpmT0mOpE+DIBGm2ak2KSMiUAIx5VXfUuENcNjYnJidkBWm6392FK
1IifhVdnI5GJLgHEFi7wtJUl6jp/bCylvs0Ks3dtQTFU4MTEsqPtM3k91SdlrnuZ
g+7aRKcNh1IupyriUa8NaSw1wQPGYRVrSmh/yJq8bJWq4SSmzAmiTiRm1CF51xeh
zZAkFJO3Df3+WxE++QmQPVAhGXFJ6ekdi1ZciJMw/XATVD+uEtziAifxSY18zv1p
MLiSMm+I1ra7FbDGc3bp77+qGUxs+PE0gJU2kHokMmKtx0JZQD1TOnTdVw0BMsPJ
atEyBOHCOWkcIvOeqxi2FVjZ8yH3Ns76bSWCFRc6FlGXJugwN8BPhLNaw0Qnrijg
62uEzqMtjdm3HJRsNMXqE1DybNw6YI50JW7MhCbpUA+ma+HwPO4WIUZMfA2MILZ9
caEjaM1LHmjtG641UkIf0dOwzgh6u2jYomefE/wAE3KRiKqi462bD4lSIhNWMiT6
h5aVp9mxKY8KovduVuIzr/yjHnLOyMPHzaU9Va+G+LCcWll0oG6pgFYc7p9vGolr
O2JN3UYIsVhw4KT77txEbyfo9SojyD/DBCL/LGdrZuLwlq6zQ/v24PbN3+I3yuia
Sxbz9YljguHeQyJtUmG0bnhwrE3+d9cXN19f/W6q5t8oMD/AsW/8EKvTMk4FA8O3
8S6z54TUCgacJGPjMDFPcn0T5svgYFKOks3Q7YRtuQR7ZIb70S6fEmqO2CoLc2Rw
asER5RE8+vJEsheDOJFZz44yHA3Yv4ynrTiJWJ0FoXyz+tyDlS+Xf6p5RARRizjO
WuFC8O/30crPhzuB2dLBsELofcMuRP5EQN+yDVfAbmEslXON1hwsb2ndkGp1gGeK
xUq08U2WQWR3PauxB+80zxvRT4tKXaGOIxpHA6JBhuEfijeEwj6Wuzw7kkCcZD/a
J+VuGJH4oNFy0rn8Q9zlCoRHoYS5+rcTvIY1aQRZK4ppKC31J7f7oIX2oM17IwnH
ypavfUgEGl3eJcyll5DEPuP5mQYwNcrXOzO3DffnnaiKp5HKgr/ep5f3ca2XhUZO
GVQ8p6iajO++sicMX3ohU2a7ZG97C9+YqRaqjIVoxS22HEjhzl1ckRH0iEoh5mgM
wLS24N2BZ/as/XJnaX5AD9veMWMsnAxH6zOYKDE5I+xP6zFEzQmpuzkeM12npCTt
rLwxyYoL0CfsXftpgkQnkBg+0rFi+UvT+JrVnT0j3uw0hGJuxj1N+WBacPhVIQ+U
8kTieR+VRiUNvbY+uAQ1/5AP+7y6XV2HUH1CDCphqh/X8NwW1/OKNkJxqBTv63We
dtlLrqaNE+qQJcWGJlq5hvsclqJzbZTZMUP22FOakcBJtw6/P7uT78s4pLTZnXqj
dosA3vaHsM8Wvl8eA62UgtIhj+YICxeqIep+Q/HriHO7puDdVjbBJxX/ayH56+uA
TmK0j6MI4y12HsZxERlzfvd/goFIT/4HXs+tPZQp3qebcPALnY3myFmPdz3fsJO7
Q4RZj09iFkmpodQLQ65UO2ew57kqHHGPKLTOhvZkLFi7MEmQGdj2/jo961G3BH8W
Zoh8E8UYrYYtCLMMahl4bSgAJJ0RNIf9Pv1VcDeNl1/hIIGuXFfHmLqD7IoMJ59Y
AQa0O2AixPf9np4tlxExbzpG4ak4Si6OyTl5EJVjQrZE+eX7LwmnwSpIZCBXEcck
6f8xBVc42Vs564JSn0vIbWOM0A7CU6yffmVo56VQ0JMWAvWw3tcz1NgX53BJYpHM
PFB9mcopnJe+6DMcc3AcwaeBnyMTfTbUjZoCntL68idKt47DzGpb4NvoyCY/qQYl
g5sCufvTiWOy8K4pRMyfjAFJor2qQEhgOdpfMWprcurwCIBSomyVDYipFTOf3Fwi
7/nKzom0ocnpejXxvAHJ+NBD/u7bCuvp8WSi+oXpQS0n9sEtt9oAhci/JsZnDZGD
QUNU4p1ON2F3E8r/TQSuFFhHL5rkLl7xgL1TElKjEuA4XOLdAb0PSyH63HCUm8cu
RvyYB21Q96YF3mcYUOGCUKv9GkM0H16lMBHLpcQlI4e4meIMeACVmPRcmR53+13c
Rd4qvzbIo7pKp5BemCSS5jHaFnlNrbeeMV7psiYsp9lbQtHmufvOb8bwgzLl6ZM4
unRMHR1cQsPzPIA5NVyWSliIQnzWS3AT17ILcc6l0x16M+zHn4EOgyqDsp2BJEFk
NTFwuNsxCzETBKUffQL+83rEyEVRsvvvnUoLoH7/7odYDpDI0B2tYP9GyiVycUKU
yInQLfPWU66JVOhF8/weSD6DHViCYSGM7ICVnoaXv/FdQOU7gOLYCJaA13xM5DZe
yA2Tz6eqQpxLfEsOp2QihWKCUSDBn/FbfYKtKNBGLbOdwitgaigPWQXouM8OeetP
Ri+rHwDXqI/7YqokEGxbJ1Vd2JBaatAef0p4+jVvTI+blAQuY928iUYGeOw6SlXC
N9AZBE94q4JjjN/6ezAseKr41iIjC/JYrPQU4rCd3Qh7Sja+ByDsap1DZBKZqI6K
GEWaaOJTGDczdGAjc33FBufepN/e1dkphUlFBwztSqwDvNEtMl36iFskx1ahVS2f
vOmJMrwSl4njyFoSYCXuRviwjefsoNFhvCx6nPoJR3DvwQebxyuNn14CjV2OAqZZ
C+PDb0aRANk4GBl9Db2+RUbO0THip8gqficdLf7fbTUbGMGgW421KgfV9TqCj0LQ
22oiFmLGllDkLfTryEdaoyOaNaQ07tGyle3zDj8aNongCAy92a3arJiCEXJLR4bg
EocSCJjMR46OMMeyZBYNX2XwxTJWgCPJe+EMcSLtuZ4Q0oQMHEqqaVRAwrHUTaGn
vxL+C2J0mdgcs5oiogWKcVGHPOSw2AMqANGrwqOEElpkUrHt6IBTuZ4J3PFMoXY/
hynU39BDNu+uDCi6hf/+Yzc0AIrYzBbOIZgNtoy+cfcr+mGoa7OkO/9andhscBPd
41lSXggfNW5o2whelLCpJv+pRyJsB/XH6HZ1mSTBhnFW4NZQ2xuy5ArpOXk3Go3f
YS6JwBMB4qJ3iKDEA0D9y2Do47hLaYlVXS0vqT4TyFUcy/38mG+/GCFtqWZa3a6j
gNarZ+Lq8KtTeox3EKxtL3+KbBlhcS00aCSI4ybrjKkFq1HZthkIKXy66k0HWvC4
FZ0xERkauyBEVBVbY1o6vnyocoYf8DCneCp3i4VenxYe9IN5zT+aij9xybm3ISOR
NGa5vOUKjgUTBUSXB5ld/25BXykjoqoErYuNfBCPO1RuEJh4IhFLTOf4oO4IiQEi
3fn/v1ZxcBrEQ/IVhBQqhe2LptprmF8PunHxWyhy8VNaspdFHAfygH3d2g2CgFJ4
AhHRq90SJGs5J7aaqE2ox6YL+FctfYQPnIjAvuNAGBQqwkpyzq7wfqdsJsBf2jPJ
XagNC3EgJJAyYo/KxdDdMhCOyiBGS4hGS42vBmGZf9PqP0jLCH0D73pnBgYvyTMZ
uX+9gROXLPqbYos+vmsbPQdoKe1+7zsXQAWngDfeS3YPMWm0WJ8V/BnEEuEaVNyR
SkRaFIIw9upITruFpV/1vnyPATqulKUN+ttiVbHwwJx9IQmQnnG+O46rSQquRJLW
uIi7RLFjQo0UQBCTPTE9iwxYvLv42lqNq+BxfoB9TvNVFAMLcg0kL0sNo3qKyiMM
xbwRU+Qgsm0ElBlEKy+DB5QbhE8rGZ5fqTtmwAmqcsVXmAOLLQL2iDd2RmnBNF85
eSE2eoONPAWim8I3njNj0XfNa7GRmUssNCWeY5R0NTGdiWq0F39LvhIcM4IKDiCM
WS4BykQeZrJwjsDHXHZ4St5EJOIbrExytTJM7q5aqX73g/lwbuLRopFurxsow2TB
OkQptg3tXe5ioGabhfZ+y6ts2QhLiS2T8oPOxd/rp7VXCBTLUTOODJpF8QN5z8gJ
IzOSUKixiAWs6X/3ZCJwDR4nsRZ9C9SoePVY2lht29TnxFFBaJAr8ITuopsKGkiu
JHeITPCcqj0xaKsuTQkkPWspfDdWkBdc1c87WDds5sDkojpmpfb+qCcTSa7u4Kuj
ZSEd+sRg9vvsszCKFzx8ZGjAFBq1hVCYaVzaWaLeGaSIC2KssDW4L7gHD4CEcb6a
o51mK+PGhqLQQdJn9x/0g95/yL5lQKq6qEHZYNbcPDuekw9fH9Cpvs1QlGI8UUrY
vPeJh96FVf0vZ29LJ+tz/hkpP2SiHCS3B2sWP0Sao5JnUYT1098zMYfgsZKDr1YD
HDEBTBr6qd5C3ZC/jvA6ka9EAQLk3a83kkvFIrvzz/NXV8XJgxS0OrJNft9C4jSn
tk0UwlUNWZg8vMN3GbCW5hV+F7t8fxWXlRQHFrSvTkNMv+zQFquf5txk+Rfw74xv
6exMPS1UToP5lFRz2j9Ba4+e2omOh9F2wXdDQho5rB2qkX/l8wKYcrtASigt4LNI
7ckjUydoj+dhfHao5tqFCfYbK54vAzodnxyDPv6GeofR3EYx/Cycqdn91tIs0VDm
r3hwb8sOB1y0KZPyG4hEB8cPyqbqYrgACaqw3bTzNq2uoTYDVlqRUYj5NJ+2TlGo
VixGtBrvSX7kd23i3etef3yIn/k6lNSqgqNHGyYXFqbJDknssMKGDIfwnroywvTk
X0TOwv4IiUcEi852jSfhdheMQiAYBbOln0XIoLXJ0+VoukElnoa1673zJcXqiHwM
qH6+3zfQFztGt69+4UI24dxwOSjqOK1ry6uTSLnyWgDN+rhP5RO6eHTX68l9ZBY0
OWX/SF+2bLcWGOWB2Xfn6b5BHk98RC4sgHZMFOA2MGHkFp2Q/xPMZQ+Rk1Jmjgpi
LwePUZvot4y5a7npDS0PIXyCZEiEZfjjrjnTpL18VAUfEgIuwfK0qFotUxqavwPS
+u6Uz8b/G5n1jJqWot8ewTtFRcD5GL+JJLzqJR9uNlDKRXhkxMo3yiRap8iaOJf9
t+ouSIxjKFY6rqCExmZdh224UDMX16LZF/6G1N78Pleqb5E2roWNo/qvYXuxoCcm
5CRPGT1N5dzd/TvMckV3Zar7GY3279o5DPQCHfWNwdWfN6r4yVCKZLa3jvJxiXwK
vqqiajGsw41S99/dBpIcLY4P/8DYAx6x4dcMhP0K+Rg24kirWHBz/mBCFA339VJl
zCIsKHSPO+8I6Iaq/T4LBaVzcuLrINCb6VkpvXG1/Mh7FjZzyAXGTC+i+SAdghih
pvkc3WK4Ki/XlSIpvQ4gnzYKXkjsPnRAKVRGq1Vb/IW3Zdw24P5nGhjq22QN2NHw
XVcQG0RgV2DyoNkCgnnmaPHTbyuYYvFH+uwTYDZheiPI41mNEu9KdT8xT5+rmMA1
GfQVyqRAudduI6t1xyERLzgPamIGJYvAQLBh03kzDH9nXPRhrufqFM0RwnfypqDE
RuANwVoSre0Czk5VYpI1cqvb//uL/g9n3DyU59IjMif+p1R4/OZAE2Ls8q3y1tlf
Uij983gWQ19MbybWIfBI2g4hoC1jQtnwhXTq5W5ustt7UjftXr8f+1Jz4b5cMvQw
trirusdchpXlGKm+/qOcgfJcrJMuntM44Ld1yfXlUJ7Xp/PWTiFSWZ/hV27FfZVD
ET80oZVMABPQpsbHpkPzmbLUXwrCxDK5QGdUP7FIZ9XCRxJnCeT+I95jDMO4WuJi
BqntCTTZD/u65VfFqy/JWRRPZyu37JzRL8ru6e6q5qkR2vhydMg8p2o1YCP2j1ZJ
Zj49x+3aGUAiI3zkJjDTxKknRnAsyVOteVm9k/4ebuJjzhNKDi0ig6I0wviYKQms
Rel6LWbZMLDjoVcxuXLDb0+QE/i76w9/DyUyn1oWONTcmbgqGBzxKJ2BW/uerTnF
iW90VQMgRYHc0K0qhBzlOCLpFcfP8ht3i8C4tG34KMaXqYdiT7zrsX/XWxfkxya2
BOqFkgGMsXg93RYUM7D6AlKEI7NhTVAieFxT/mx8E9OHl6SNZTdVNE3MuWyLrG0g
VpYI0VvZmr0U/b3uxOhJJuXS2XePdxHZdx8KLvlp+ugS9spgkuEd2F9wCxYo8Mo2
ob7UbnXEiZlKPcAdAllOHcQe9oomedoXKCqvlPU6igrK5w/lSfroNXGGLjjC6gDN
H2ROPDe6MMs1N8iRC6sPXnfhh+YQXcZvSV83oLLTW+FbYVIPJ/SrMcCEps/v9Bd3
Vkr/jiDmbAl++DuME/YpVsqUhtnSelelhbcRtCszvSBMrg5nqcyZcatPurq43+J3
zhixehR6b8apgOPgchguRxYAFW6vpXPtNYZmWBTN2Y7mvBgCcKHk2pBF8pSG7S6G
q642Jg1Ll3hrQXidihndedSlyk2mF4Pe2hoAdRy8hzztwJ6WeoTAvzpzu93Gzzw6
hZy1lzGLekXkDwrDlXPnF+dfd8O9c3ZMOstMFwl+Dxu0GrFywjoavsDHj3P6e1lJ
yDZ0CtziyoedVxgZrdhftu8lhGo9O2nwauvfWTJv7SnCtRRt0nPHEOZgxu2MZhH4
WLoZskJtqPGU8fVSGR5/CMzWKZ/PnA6AMYkfR7O0yQjH6ZWYaXZ6VrskHUd20UuS
LqxOoidxsZvZz6LHqRGyrUObmIrZ0e4ROyy0hNTVmGd04uc3setnUtxUR28m85Ib
iDAGRBsZwibFzXXK9bR2OZjrLPkjH7VeSkAsc7ViZt/hwKMaQicSke60aJuY1BxR
acA6xQcpvXqV45xuTapTaKhHuqZ1dHL0O5mDmOeFmCMLqSijpIlDyGS6FhPap0aV
OsvCLnzq3/tMsNagBC6lPID8j6i56rwr2sW/hTwy44vBp4xtEuZOmiNTppWdeIs7
dIyxSMGylW6WwaXPLQFgA/q8rgkQwKrb9BkRfEELN6sD9F8YodxGYxh2IooMgz+c
SkEP+gIsIHaWcn2uq1MFOAGaU3VT06pWB6tUS3aj6BDQrk6B1gfIKorK5eH6HUN4
QF57+zkqg8KAo0I044N77gJljmn4MJIzFDP9wve0ZcxoZndOvMi9/7tRENri+VXn
wo3OegPWmelXWB0FBF42Wnti6rrKdSENoVDDOHmZ3UGNGQ1T/Dc1HYsoTv5HDANR
S6B0+re+7MBiIFWgCHqWS6cog3p4jDZAajOVTgabxDQZLtJ7rPUsm9OX+LVJ+hKI
tthUvTW4lQBc/QLV6k7YkxYbk3Vac7IpRhRwl4sQe4eKf5WUMfMdlspxc8JpAgQj
zsHm0nQjXTiOKNTOZYZssR2jjv9d9EfLl8+egvq+Yl+t/mc4N8TMkWX8vjN2H6Pw
PXWbLo+BEX30J5HpME1qDjU/bAC0lNdWw91d8kqZLCB5ao/yyZc5jtw4xkz7CjtN
MJAoHfnun2vIMGQTTH/decIlaCtnoY1fABVluDrzttHVGhvbvR/kebmS7gisBJsh
3WHWof4PP+R80EPjf4bvQkMhsEJKSIWIDNgatkkQFmBlNwtMD1vuZwiUGJ/kgCXd
8oSP/SGxChH4M5OVQiNV4pcW75BC4c6a+k26eXSwhcSelltMIqg53wi64X6pn/3G
6NrcOGDqP5LkWeDj4HsE+q+CEQsXqexz340dlsEZUKLLKU2vVBwFlkNlXEbMSnr7
4KNWR7OcQb+73T/nlF9aawQ0fultokb2QYXNnlV4b1nifOISptn83nw/SSaLIsDD
ak7JdfaEEsDBvIBmYliyemLmEqj5amj2i3V0sq5DPeMtEvoA5IJ+2CXT/xmveyqK
M0z5tQOyxGj/bo1WApf5AW2SNCWaXT6tA5hJh3iLBZ76wU/DGHLeH5A9UqI3IBax
/pLI9JiVIhDKlBPfaOHm1qLs+vHtlYJB73IQBWRGubN+1QyZ9Ivz90stJaO+W3J2
b/kh2YfsQgD/iX9uJtGDzhSMa9U2VzgjkxBScOJhT4hLGc+ew/59CgzmShK2lwig
ppwwKOvbLmMBY40vmbmWAdw35pSG+j2LM1c7DEzkREEzgnj2SXzZmG8okOnT1DiQ
erXMtGeRHTOw+6Cimyncemy6IuzLQI79kiXTjassV9ELVFSeNtKTdqmnjlvldAVM
FlLqB4kJQ9rannd90zncRKzIIDm59u9ba2XYokw1o8czPk+5IMnywsLzcDSlRsIu
drmvWehmScoNljoy74cc4Pt+VfPHdn7/mhSdIsZ1B71ejNXe0Np/WGDj8exGZfEm
YmofTNeGb3+/wW4pYMkUxY+dVhJlpVt7JQ3GIBU9xQ85iEkvvoexqc8dVrhaVUtA
yRQZbUF4YoFGaGwnhvIG//yUBfZN0f9u+z7PYARBB9AbDUpHrIscFnK3EY+ReFvG
yaIJVNtzxmisTQZtMM9mTxaU4OmCVuzBuz944TE9IN9EExBLwdBRGK+X3YuvLx4G
M8AoQanlawbhiKEIEgcX3e7oP503G3Pov8odtzIvZohNk6jv7B/H5zsAyncM9wG6
OhOJ7VllDqi30w/LCzpOwa03uTUCMqUuYbTFGWCFYWVLolXqVMEdmELdO7G6epj1
cAk8w1M3kr2Nun3O2CI0r08hCuZcfZNVTtsqMkGhLDddtvD6hOt27dEKmwvSEB+p
UQVJcbsaXfGDkAlNYCy22O16J8jtSZtf7ontoFuB9P7HzA9BBQjFG8clnXPajIyU
kkSFu3rkEvyRJ/nXXO+ubS9qccPKIMLoTuPKOp0Kurbmf/Zblb2U/ue9QFDeC20A
+60gDP9L9gSf7iL6TM3rEQ1BrB9fv2CPZwmBJKcW6SZI+8O/tp8wrmhBB/sIfASR
N4MaJVHJmftAhc7aM2gd3yaVugvGTfhtN44IPGMezLH0jJ2sNiCwBg/AGA58J8Do
OVygsUHCzO9Y2pKsWivFAEIBCItADdu2Du4u4xvuYzOv9ZFFjs5IrqagXHVyNw0w
qW7716bIBrxpbUBUdpcDJOakG2/S3Ftp1/rMwuDTtS7nGEJiE6565pL1r7CxWIPd
naea1b5wOAPHueVKWsujzi2AfXlkpHuo0WaBCoEbyRlrpVHeEwv3NigJfTHAUAMK
Ip6bKJMlUlCsGQTJGu0pEe01SLaiSIk6OLOGaBnV2zZ00rj1RDwUGeqdtZNTOElr
utGGdvJi9wTtyr52i++2dMHLq/NcSNzxl41HrVwudZ4ErglB6KyvuzkhzH4udhvQ
gyYQSh5Y6ZQF8vwgY8vvFgwDWRp/OkezPdyq9r4gj2iGMwgKKg/YslG4Vvs/zqhp
ps4jhL6c2obJQkuEAWmh2ObRqBcfi/aK/r0/HjOv+DZwmYLgeVHMgZk053RWC+Nt
E/7OL9T3eFhGnnq1DSGG4q7rc3wWEwh02u2FrP8xppXvRkxWO7RIyV/vtagV5noE
UL3lI+Ldw5QV2OpslZ0vZEPu3RZOUPcEYSWQ/EtupjJs9apKLEneUHorRIBudLQJ
FvW0N8/ZyQN+Fzy74BhLHMsj2kBNzXEkgd+MuAAGHBYTtGGVT4zzR3UuHHjwnBz2
Gw+mR94PvDQIs5xqY8lHsOr1MFu3kHXBO6o1WQjMAbq1xmX4cXo5y+k38R6ECocf
KOlHwTTQCiLJZRugwBw0rmWlbzuOEDbfmkDBoFej+/pMeHulfa2syR029NBoseqH
BGKF8IqeCJg9PHgwCtXfXAgAl8/uHQDfsNFuowSNTAPNLVM6D0JnsZoHb0ItZhAC
mmcEqlQGLuhEtBuq0KnnYv4+EsTOKSd1qlXUr0QEmHm/H2wYrIocTzhV3LP2LDuS
MxrNa8lprq3soqpB+TeuELZrs33Cv3T3wI1GRVOXxoNnywNZZ/i2JC7sSfbQeO9Y
WTNKt7u7rd7Pc5SF1u2LWmBxI5dAYQJScJXTtR+J06usSbYunE/BrXHoclBPBAqU
9f9MA8kX8dgNcaJq8mYWKmuI5dSDBGfRLwYdysC6+h8En3AGWrg8ZO5zEG6zj6Hh
qnGs7u6MfGfoWCxY42NXihaY78tdcnD6DP+xb6uY0OcNwyt49ihxVKLgFn9KSBB7
COlIO/WGLR53zQ9ixzm7KCkeet6fnH3+8ulCqq0CL3B1FcLM8Y5I86MVOKx5ckgn
LPDfngJ+ifrUZ2C5f29520ePVWx/0Juxsopv9t65EQOX4I2/arW0VFlGCEhST33p
azvbaQoy59qVve/qyj0VmuiG+NSiFpgV7qBUWXIVMlRAOq7z+hD//8ZB2aekzFvl
jak88YC6K+YQ+DtYsi9dAdY2gwgZOiV4JvGUvo+bAIF121Z4jLJDDqqtu7u7wkfu
xTMAt0CICSaQ10IOjN78SkUYV/NHXTmRkyYQa9uPXYH5jtfy19vmiwt06raTnrtl
QiEpo6r9Efn29fyIO6Nbj7Pp2B5OxbevSRS8bAfRpXk7R7nsa/d5QbQpfAqaGOkO
RHsS0N7FiMhgTWvFr0pzXJpzYAwKY2stocIsgw9vlVBy3wOhb665QgzJBPpIrk81
mZz3jjcFBDT6TbZPwmqaDcPJs1mkJq/8BT0bfZWi9e3Tls2kRIBSjm8ZE5A0edMs
xjyxwHmp9F3VrnqNh3TM1YEkZ9OzdZCWDlyVtJGO0DZ0qYAzo1eKtx1SVC7ovgpI
6WUiX9v9x+pUEKVoGN0TE4aI+cZwHL9+mFzB7jJwoY9uD00JM709iYMxBHezjOjs
US2e6bd2lDDi3P8fZmW3j7ZxBSfs0Gns3jVPVr6kFdvuZZj9Kv0ov4oFTsICsBTT
6yCG+C7UVLGAtL9KUPHhgLvxc5qtKZXlAnS9H0fgU1c+zn9xHlCkFE/c2tOO7WK+
tUQaSJcmV2GBii/xrWV9CrRx1lQk1S8PXFECpOuhS1S0oHwBBPb0+qicojUnDITj
FVAqiTfCOz6Rw+RtcG+IOnoX15a/nSmQ1gg3OxKxOVlmwdI8yj7g2jnw5CQOHLKb
SNN83ecIq7WZm4YhvNmafXxbGgtmMpzKSl2nc+ILP2bPlSHOX+k1AHg2VTjDm3t/
EMzYnZrM7fox+0HxTc0LIkZz11nN1Kk6xquxhaHZzVShRYdBGMp5e5XLqFYOpsPl
RZ0AorETUFV2CK+4PvVZ0olYLOcAhqcCF7+Xa8BVtC2Whgcg+AuLCDniAyPJGJlZ
0bAAwPt+KioGHhV6EeFv6YlRrKaz4/6siPsQGwUADxVIDB/5zgr1KeTTqtNwebyU
iU6zsylRXfKFL5yo0s5RxvpgOJl/8tBFLBSBKY5XULfFbmGpqDdS3En572meZBXK
w648cbzP7omACDRM/oEGUrnHoragWZkAezf/D9brqRvJAfheIIBFluMNO5KnIQcB
J90dFx/6eT3lZsn7i7gS7hpLQRLrbyhrvy8SOz9/177MS5ubD3ETKk+SG0PLbKFZ
6cW/o13rNjI3k/VYmnLV9AAaKFeHyGt3ebBZ+AhQj2m6Ld6Fs8xnm8PTkS1IHMml
1IiTImmXGClROt5hVPF0gAT+jZoxRO71PpIpbM8QcWOsVaCCr6Es2yT5KcrSo27V
6Q7ObzhTOSm9NY9zR9XBSAXjQyg21Q2Yc4PYlTqOElGh7Mw52cDNNI0hNmJzdWaS
xZ9LIC2N61xR9mWu+XjWNA/FSMKTSondSgq7B2rdcHj1H+0nqnWtlrtEjPFRoHmk
KdPb2I5L2kQxZIj6DaAnHmp1WxzFqXG/BC9C36QVr329nHkjDW0xDTKP8WXcG22m
mIg7fogZ7sBWGlgkdvbTbxBw4wISNnxVfuy+2e1ZQ5NNvZ07smErgve44etd8pDy
wpOGjQxzhD6wlRwEhdF4ZMrMptZ8p5atsO5fg+4L1QH9pEy4n+6PZ4GYcG+kXVff
Wy2Ck/FSJYwF+C0LJZf+9y2tMtnlY1q1cP06fzOsoJregMOZodnZlsDIh35I7A5H
oOrEdfGCZnIcarVKHQhRXbB26GJD0eUWttaDtoEzWL3k6qpX+3roVK80xT5wV5Yq
pv6t/1puryC7twd4zX7mhoJ1k4v1KkB0wIBfHrO//b2QLf5rOIT24U/CfvSdy1rb
K9F3ntBQ7Od3O8JDvH1uNLSR0Hx9F0iMMqGSW1mLk//xCZNpDYpRurqpAlXEANeI
NR81GrO0a6/NMelYkgpbQO5GnQUiYNlbk8RVmLGTAy0hFrFv3HqjT2+U/7bNlttg
2KP/jx6PG10llDnRvplM+BmBbyfHg3srqnE61+ddN9MEtBjuMjek/gtqccJiCzl6
ccBFIKVkTXRJuuEhtTzTtvnJBAZdvwJPi5C16w68GxmhGPJYfkD7GARDewmxHNpv
KcbSOOD0ztNV958KDeq5NBfxkhffbMXQ1uu4CuGIrCbCMJrh95pTJcaA85EkkjjT
HP7gifZT2AyfUwx94mbaBHROiPsROld6s5cPc7j/mGNkRM5L6cysvFItYtI+Tjsc
hqbyzhMnsh8Dt+Hfqpwef7awb/hV6WdtcsNlC1rkamX37G8X+WknpvYe3LNkTi/Q
QpyUecWWgaFec0cHIEKc3TL7LxlKqoZIJP1yq5QMrIps7jV07zzU3aAUEr2D+P4V
FGV6k/PaVd6ya1OvtSPHfz/34q5LhtHmsOf6RxB/ZXnnhWHJZKEnvCtVvWL5dqAF
8HR2Rahj6IUwJEroAfZAs50DoRPABRTwepLzCsbNfkW9b9DxM7wD5En37rVGftgR
32M6RNeDRSIL0M9Trp66jmUsanKp+SgPhkHSrFSDmmFlj5Fn3J4E7kifNb+nFbEv
hjufBVVLrphX3XH+3FNq9zUqJX46E5y3T4urCorN3XJhF1E5UTBQmQTUlUbP/4QF
uqHVAC8D/n9fjYpDQvlrHKZRb+lIEjSwATu/LDNFM7Wd9zFSzRYsOnA6u7I6Kpqf
G0qfCw8/h7Ry2O7pnF0dgHAwp5g04xi3AODelgKo6x1emg95pIY5Qz3Qi11ypOfB
Kcq5gHodQH/F4l3o6Ftb8TXTvaS5zZiqUHZuDkGVCU/a96VWg7IeY0MwpT7yxmb3
czR7YY9k8hNTD1J010/Pv8yDu8z7jcuwl0jY8d2pfa7ddRbNlHouceCo24XCCjTT
1uhj4WSL1qz9dlWYmiTtO8xsggJ/W/02RYzTF9TCzkO7aYvBs9IdtDtLqKg/wEVs
0RdOoumy/2Sg1GyromskGaU4H6bZiPFyk0cdM2o5XlAYaCMEqAITmOAQbbvnUkd6
DVk/J54tGJuRkxGzZdPBLkwdoJWyPBA9k2zvcM1SIWX6Tojry5L09pS1l04NFt+M
81W2w4CNEhu1njD4cASpfM20G+doKiCxB7QzWKKUBM+cVKauk6CCyM5bcjdKq/cq
DOfraaAqgu6qPGmITQ6aSYbsRv7JWruUXIxcg+dS3WeDWUDKMXxRh9dmVI6BbXvq
gKDjEzL9pBGYFoBg3uC2bKSuowHe3WxpZDnyhFRL4ifJ2hakiW372J2CkTiqSSa/
jJQwa7sB+GOyzmjnXweQ1AMeGhOkAKTLlEBxN4Ii/jNfXpm/zPaUWmktb1iwgQs+
+PwsM1vm4jxdWaC2omoano6XysL23oLOaLPO7JLTWGyL4fAtRRTXWVln7p9zXYa4
NDD31siVWgRmR4E3LwBF/zztN3Pz1pqrbYsPkrXvr3+rrZ7idp4rWzjhg0WA0SSP
9mq7tgQmqQAs6OFvvPrkXkTDRSBbhnWDQSmioJm9XERGchDKJUFr3HLyT1Z++gml
qgcAH6xI3TRYCTJJw/RaFB+qj8jW1ZBLANcnzFJUG6uB2vRN00SPt/8QKdcMhZyV
OyDQAz7zWizcu2Jl4rjwALZUCfUlHRhETOK7208Kx7Gx+SjC9suEuJDBvt4zHkDv
Wu33cRsD/LwDkFn8jJEwLLyXkrB6rAtdtYi139Cn6AdyF29O/Nc0uP0tH2qyHbaE
WesnO/L7n9oTp13JUd6AvexT9wYjRZTkLM+3Ldo62eS34S7tslSfE7Ow1fVN6Ecm
5zfrGwsldBh6af0KDnS7uZ7sHnHvCrC4lHw6pHfbTPbf2trTuSYFEBmNBrIZtKpg
+PnqbtkH5P33PyHIRiV4oMUsYfo4K+B/9IHav3ysLVj6ZnAUlUaF4lwHrOSmuxqH
iG42l4CXdezF5H0igZMYp0FxtJSOY9PU2g5PxkCURd8McilkJrDtwCI41Yc1KTet
6HrSVQR4HBWsAjx79u0Kn2AG0+hIudaZfhU8zHbMUqNvqs3g4FDxGkXKvxN19ssz
zFfSYkiaUcd2UGar8JxbWKKFR4n7Ets8ijvF516SWqEfLvomdDDUZpbwOAGs6n3O
HYWS/aOH8vQFSRcf4ruReMvEYVUC4FXEd9rXx0mZaToSCZ+1wZuCNVmD/eHphuW/
k0dNFitNDFKFLww6IwQiYT6lnwe6yK9pKv0+enrVZp6zP/bBZ6mcPcbp7qA18l3m
oVn9Aay6cZHSt+OgVlThZVgA43iWiroGEvk4W88fXWh8ELyv7qXr1ysT/iFpyyjh
/4ZKhh8uLw5HaaDeCqC8EujGsF53JtvS26Hle2zEY/GZIjbcNC7c9GvIp9ZdSbIL
qCTX+5/y4A2qHoz8liocyPcUvO0z9zOLK0ZxLzkbsvtIK0FjFhoKmSfYqK/YyQuL
yJDcl4H0D4eAUZVk/tudmp1U8EB+uboRjw0RAjfk7xGpLdu+Hk9aVjUJSxtxK6wR
WJtxuU8xIhKPmvrnvuj6FGVbMt/a4c67KK1kj7goT7o2uHmWWTxW2YOhXJUJJn0q
2MvIPS9O4UQPWr1SN60Ys4uUH89CgSLvCFcsCr/I/z9Lr5w7BIrzI+4rCQvLeVlq
Sw/O6DqH+fClK18xWHGGlX25e42oDccPvE5/q9DIGjLPDoH6McuyqiYHBHnIp1NS
G8zwc8xN/1K/8+vN3qQOwyHbSjwSGzNaGy47Az+wBLEOr7Fxq38WTJLVD8Pyuglv
eFWETOcrVSOJX10rMeX/Llwjt8h2DOzdb5gcQ4jx5zd/b5pBXmQZ5J2kwxQla0ek
FrGInwbrgiRsBX0dJmmna4Br4QW2HoysA7OTcEgQZfCCM3rEGVT2PI88+8b1kdMc
CFtO5cPbeMrJpcRtbTBGpiRqIIcv2R2h2liulr65su7zdAx7ub8Q+0IVbKHGOdl6
E9b/x8gtmJPpS1Sz3as5O9Iav22sb9bJ3Qdl5vLrqOW27FJL8h/e2TymKl8R7jdo
S9cJCqwEdmXenLj5plxFm/vYyKcjkIl+7Ll9gNJiSAimvUYXWtspX86X/7FGg7hD
lb3aVhyVLSGWUI4iRF08LnisG0m4KkzakHtmy2Q83yiw5g43Kyosa3sm6nEge6TI
LhsWD+GVot49Xq/AmmQvirrLlTFlVwUMk7t8FyoIfBoxuU+d5JaMpstLtHKc6A6L
7gmrABACrplJQrT7eoIKiyCRN26DSpUvAX9bLT7DC5LRrBmVnpcJ8V6vvp2FHwuE
tAwCcSEZUA7xaMK9lH3LavUw44V/DUIoxZZuDdeRTvkjKOm4esS/6yODuHP5vpve
qm0yBloy5TFZJq1IFxbTF6jfP4WCRhJfQhIYpKFvEFTtONIDD3hK5AavPgzkTgFV
MyEHFzhAui7znbEeZdjQt72jtXhAGJqaTqsa1+j79gSMBxfnMpCyuf2HB2BCpljB
ecSsWf2HxnQvQ8OJbuv6Vx1gqYbKWujWxGVYgH+5mDTZ9yfGVcqU4QzPSf7PAoEs
ch2RbjLZWd2TdrdLYWHwc96PNsBYhXQro4dBglyGk90ywKtwCDj5P5YMm4QDxmhx
7urGqt1Tcw1KdtCl8ClwRudCp8oR1Mxg8gkAiKoBLLGVecBCYlcdHKFOht7rQsbN
S36GT2orS4TnC+F3CTvyzHjx4lmiZkOtkR2l3Ax6kOZZk02+J5BLJQuEr/wrTk4n
7/tKpsHihfObSXUmWAv3zqMIRW1mgfqznkf96Oc2ioVT1ax3iwUAKfTdCiNlNiij
Y3cRWw2KkKR3zwmJYQjEpcuf3RdIPchJKBUre1h9f0YnXONedv67kUPdLVumaofN
KMrsxIzvZID0/cu0wR+8AozzZ5zEgmV9pA+LYZaj3UfyuslfeSMydwfRPc2t3Zfy
yeh4liVgJX+5FxEgrd6SBiROLW3G1G0E5yNcAK4GuQIuzu72qVMUBNcPay7wuwhU
lXz1ViG9FBrsWNYSV1m0LhxngA7zmf+FWA4M9uJ63cTf57Fx1PTeiHGNDNZ9yi+N
YPEfqJp+w/xtx+0BhlSsMF6Uaxh4HjMkUdxPOef8Bkqfbw0Yi+vlVdB6DL6FOUwg
FWvi8j/LK+J5D72aHFt6hioWo0KYih6R9rGgcWaJV4o6lO1XOjCsgaBuC13lRfMI
khNZJ7ty6LkRr4R7KKV/qlawzulTkZ+hwEDuFZe2mp15/WlaSKwMyL2T8/a2VlFA
Xk6PBSCS3eihe7WQAXjb6NkzAu0MaDA5lpIAQoTjMMcIwqtXYOOLYuOcDV6UAyw5
wb7IdbbWWc7XBg4I+dytLA1DDjMmBt/Lw/uLywjqS3GypBU5Tf5ze1vGijbSQGNL
cDM/ustahoAmXKsiM5VpvpIHR9m8wQ/9tKp8gNPD8f/IHZvNd9+ZH+1ihUE/7GZD
qJKfApSurLi2D1Cw+iU82Y7IJDX1+zANhxI18IBA0lZfPRhZADTzFIhPguflj5sw
HH1xGBEsGSBsRcF3xZ17USPVriWENTmSkZZICP509rLv2DGcu2sHS/n68jjR9tHc
xp4B96cbAPNzUS+7rr9SVz7XPRm4rkFgwxSccxcO2jVVUi4SSOqU1ZtDAn1wlVSn
Cb9CT/rpwdZtIDh1Ow/OwSdgXBgaK7HSY8S9jzPsKXkaeO+cNLWt6Qb+1CF3JYWX
IdpGDBQLjTpyiBDk6f4U0xacbg31TespXN/o9/dE2DyEPUI+YltDln+llYNVveaF
S/qX0sRLzPHQUtdpKzLLp+2g0ogh8ZIsl64G7lPFA06S2TNSyS+Sy843U+2my0eX
etXgGBKCmv98CRrl0Y6eWHzo7JHPkmC8M9sPBehfLInpJfBKGemsfIWnNMQ5L7Jw
hNu0h8TEi6+F5+IH54QcJxK2BMv2A7tJkOpSNCp2crEgLV2mcuLb4fK3iCbhNnxN
cS9uvWjjzqwUYuJsXUTL6KJyAeSdTs4e7ugnyhj4IFlLHtV3Cc1G9PRyUhELetjc
xrHdOTpGh1P/V8BPAH2lx7flZ/gGFmNTxTHyrVxw/xbl0qRczgG2tP7JyXpk3ieH
m+137++gmcAZGZbfR8aMeNz3c6I5SD7BAb7gwEy5qEKVWR+3lbFyQXvf7JleMA+3
RCJA/SP+WP0rBDkTGZNpbpQRQbKkd3qH+PFn+vdTRHjgjTysNrNg6QtlAN5jN2xL
HoDtC0RFcPLl2YV00zCVjai+U4yq4szLTcclv1TDOp+i3oh52ntavFIzD2NidVUu
GMQOpu5IfjMBFCJti44VeO2NourwPHkLuOxhlcZEShl4lX1zG4M8ClWIS9rWpCbB
+O78JiKINCUxuIO1hndbMYXVvewdJwnZJ39UruzJTWTBry2J5+ru3YAmLIj500vn
OxWqwhEwJnAawY1n9aW5bCMsiecAyuIJyxVy85RH0gXFcuVNMcK0XA8lvHgkKwfX
DSPd9vFeqtHNAh1nxfT30ycMgGJ3isP7M76VpgNdvzMY1kWuEnjYk6ObJ+EPggWY
h02jkAJSLUaPXcdm+XY7h7zTdxSG4kJ44IuLyT/sqtLuJ8JEFwfZtlBK7lkh9PTE
/dlqlooiW4apLARX4ESdoG41XVniTfXjtFp14wGNDtaDWRGQcaQ0RRkpLeuqQAXo
UE85777OTBwUoQV+QSYKW2SzZE+6bORmOxxVpPvtnr9ApdhstFFMguYhgnAYD9JM
/oKfzjsJ1N2a9eQ5kjgg3PDqq3p0dzRSLrXV/Dw7BeNq5lq/Z7RNcD8b6UWw5uFO
6PFMBcoUmT1bX6uHGHWza7vb1bd19mxkXz41JhAr/Gjm0mp/zWAs/xVGGgnnhdB9
jCTR4C4mc7Q0wQDoJGpHahicSGENSS8eFW8Gksfatfu0qNI2p7DV1+bPnR28FUZz
MPLkAsRMeRGBGtsL1J99VtV4BmdVFvHKkTMjLx5v77KoWCA+1nNfBfJax+8/+VJf
jGBgiB7723ahkxEA3ysRh9hug0FKxwm3dVBQVoz99u5StH3eMMW6cLdhJC7NgcYA
V68Vy6KOYAx4C24w4FpPp6sEkL3gwH5MqnYhuBt/rpQfeVtNUwtWnHeSzxQ5VP54
EDSzzxg29T8OL6JOV8cciKRqAnZ2js4zhq0so2Ba5YdDcrVf+177O6MmJ5OI0Uuo
ZCPIWN8nk9qlLwr9W75XTw0Za9bepIGCyJs1cd3oFWBmLnb+e1sjVSLJ/LXxGnUL
YblOGJAsxp8PBSV2PDGWHG1aep3rFq1qsoq0gTMBbwnPI3RRJXz34vI/jIgArpbi
WHaoOHDhAEnRl+MRZ7OfT1XgbeYeGe2d3vTc+kw0BsdsCwYYAVOCE1g0ZrScabxs
JXphz3MU9G6MM39rYqF2inwgznhmICTYIWMWpwlb/C7FWjo31tjEP1rbJu8GH47i
hwKrt0O5e97z21LVlR0oqXLVXGZVTkrJrRAin6HDGrKZ+rSgmUypBEo5L4Ty5lV6
VyQZSw+K27n6KjB4j1xXNvPWgxF+XYhhA/zsGMv6PwvjPIzNMMMSvXqA9CFIKOZP
G0cyFOYnXKCdzTnjM7e1DqjAGb5QwRRF9Rq7w70xPbEdDBc7Ww5SGQEOnyJidDKh
vNq5o+s8cSynRVfqJNqh74cMz27WrN9+IYhYyOLhz8wDIU/6pMtiSTwY6ZHlqNab
DCq33sekC7ACedykiOUGbpBeNbaeSxJbcZV8IJ65dba59mmUjgsHMlLowUS+LZ3X
EzPDKN2ASXtF0NGTGUJgW43IBAOmHySJISxDe4D7NxJI4qnl7Vtu13CtJnpfpaEi
ihPnShIS8HWCTvC40DjNoIHwjAWqNeZS3LvQlvlwWhccDXsqeld+CA8oKmSMSl8z
RDF7bUOGun/YduNaCnRAMQwb0VeZW3s65ZXaP06sV5zNSon8TcL33A6A/cBHJT31
dEo+VRiEYH6N2F/voAfgNQJnsxozt5aXrGkCoOEoJdlTDSC4fYqsOQyav52qJxAb
7n+8sAY9ELsFBZfq/D9hWrQCceNYvfZi+C+ofuEeyhSO/nAB+pSUE4OMB48Ppa3c
gG0QDNlGMkigDizSx3AdaLJu+mzrAwirXIwHuZ0nF/Obseoa2q5AqdLjnBgDJRS3
4nQXAhmmSBv8xY9sjVrymOQNQkKR29Zc10etq86ugxzU3elwa9gn6LCIOyn5q56w
RCgILGTGfLVEVo49CgbkExcDV7x9LTe5SNcdY5G2Hht6l5fiZ/nzAIDEXuHnPQ+H
y/Mf/wjOPGdDdZafODPL1mMiGknqY4k6JbwoTrblsq9YNDMDhNgwdOBDFbuw73SB
lhk8ZbdLHKv2jT0LibEuQVYVBpuH98coM6T9Bgx/jxkP3pbJPUGIY2olI3Q+iscA
Qf+HtwS1OU2w/37GLe/KlJMCmmhlClgM4O0hDYF00ZTdqJnEdHFmvPqXZLsRbT8L
Ft30EQCidRULu/FD4HILT8PMI+URe8UwwLLu0wnmHPQCsQ0r7nqcM3Ad5pxlZOl1
x6Yn8naIt5fFrseBN1eRJlRAZWjhNEb/XiFogx2Bxs7KKq2qtkJnnXPjEn83D8n6
PZoCThNBW1yYTYu09jzjgMTxxVotYAuR2m12xtqGapcHtJdkyle15LQAEMGlKuhb
v8sDcxjI3yG35V7nQLOxlJFRuPQQeIxmaUbAzB1Cd1WmniWHzOmWD45i2dQ1nYEo
Tu3hHOQBhnP2Yxr0LvbrvnToGsn40mrvOhOPSO38JtZjsy4lkiQtoK5rJ+aGpg+j
HEVYEhqApDCy5WvGQ9qSQGwSxd0Jrx9tVLny61pqb6t8jw1Wnuw9ztrEnDv3wUuo
wUlBAwtaQpZj4qWybGxoTGke7/TEkhQbBbKZMDMWh9EYdO+5KqukQvdgSgZec6pl
2SF4mH8H6jvJ8LYw0uLFt9gc1twT+lC5C1eC1Y9eTJFVhstQj2r4piUzbblRwwL4
wSHMmu7DOSmjWzxbQ3JDp8INg6vDWh+04HXYzxuasAQjvSRwARxLebj5KO0xnCil
oJJ3Fmoy9zpAiL9NNALFqjdnJlM9p16avneLWDXZ9kr2o9+9r14GlCx7PlaKn/7p
Wej8efNwPuc+CKd3usN6lu8a0EelyJrjGe4UiYInItOhXU5P/CoCQtuertBRa+nz
zT5o9pLsvK0UllMsREllo8N9XBW8KSXqCJqpVEKupJZQTaaCLtbUJM1Dejta9lIY
BaMBNpwOH7g9+B/3FuPwVDtuxI0GbOIdM/gTSo8VfS3F+qq911SG71Fo4XQDUaUC
mlAPQoqwNPWxfYQYcdfYxdV/npbEwQ8VWnMp+PsDyYWhGlpcEVyukJzztcuIct/W
QsbMIDrX+i55iSa8xOdLMcygCUvOb71Vs+Q6p0SRjRMkRWd/wh6gpVBqWQr9hbA/
VmUnplNpzZkEKj4cEXetQaNQXu8R1g96CsxVnZoFKEvP80p3nVztQzB99+Szf0RV
OcQq1NeePIP4xUvJ+3nj/EFPyYFg8uRFZMQI0meynatb49EWQAWg2WLMndFVORVj
OAzFAVZg6d6xpmU+22e+q3O89J8tY+AHfcHeq5nW3exHSKNlPqKwRcKnLxhvrOb+
0vLFgqzs2uKRf+gViAKjWy9coAquhN5ByTpPP9Kezo1Xfv7uivUiIMOXKWEErL6o
Ptt8gqEY5hqaPpqY/gXAvwbl1zDPLlrogaZx6sOPrRLeZszUFBjJaxCvxICyOrNr
7E76qcuGVEumln3dFZG7uYCR3VOUJTVrc0G0VLH27sOd/UoK14DUrFCHzErs1uqr
VU44068TuePJnw2HWO7sRcg9HlaSY7498FUaoQsV9yBHfx1shIacPll82i8+2fGd
UUyuTuUQoMsT35cclED8bS2omCj3f1TyGMSAj70oq3YB5T4u7Sk52r6ktn6i7AlU
TKGuwuP86m3UtNVKv2mPvc7DP2STUoDIMkvmvNNlwJMASkIVbeXXCeHNsUw539rl
gu/42Xo5X11otNmYYlxqabDKifKhpBHLyA1d8eKEFFdFc1zTlpS2IPDbD2ZUfWM/
D+CRnR/Dba/I7m83GsrGAlrw3p1hFNM6ykKj/vBiyEYuiAjShOIOPv+p7gXUY36E
g26r2zKs3TrdA5fwTy8R3ynzvkZzGcCSlVOx13M5merXvMkpRYadUlWzRszvm05k
Px+XeVrREn5JnsfI+AKfYvYSdc8tVM66lqB+gNuanvvnCmgmeVSm0fC1GeQ4exJG
8faNnz7YqHy1+JmGv0O81QscAtNU4oEALU0ZGf2pWp0ZrZ9IGO2XIUAdlRNky3Nz
SmGWeaK2lbxHiqwGpsUNJVETmBwutSot8yNPUNgK4nxaEZ8HSI8IhWo0lDIYB8P8
rZEUTpZmjpBuPTbRz39JOnrW8w057gGpitaFxVxwMcd7sjDCUMi1FZMM7MZ+3gje
XpWRyNzKrMzeveFg4mMsAPwhHKANvB1OUinzerDkcDMefTgEf0wN1KQY2YQ6Enl0
3jjTejG3lmEZrtsK04gl+utJC9MMycUX8WuQo9Y2XfaHKgu20Omro1IL77BRTdwy
xf2xKJTEy/bn7mMVS0hDfQ0xJrfq/VX8YXtxN6nIp798vxFPeFcu/BVzihFNeC9y
9yoxrXyIy6g/7hm6OOquvgCpAAnLsS1utnGMiyfBdbHX0aryQxmVsdvNvVrENqY3
2YaTkmn2JZP9gdadt3tKj/7VRS9+RUKn+yYU/PvqGafPR3NZaaJ5HqakLguueacs
xB87esOs3naYuMhjU3Nb6OXedaTkXBbEpYUSjUS6GT83wUze7EuytWtNiGRaQMXi
zhJt4myYlJSqu4FKHKIKP95t/76Wx6Lx26fBvUSmsbu8OHAoei085u49xDtwywMA
QBswntSuApAFW2KF1brYZyACJFuah/f9FXPoHJfuZOvnWlTgfNc8ZzDbvdr4+z4x
tQamGpm+r6FMZBAb8ZNKhg+YfnS/IuxiIWucFALzwAlZvhFCrPjzIFTnE9PzA107
UP5HEvA9bAQO5VIeRa93WcPKHSkzDfgBQVW5Inv///d/k+unsvE3QhW2p4AN56ps
oE02/OCFpzIGkZMuGqPMfh8xPomdecqRkbFykPYSp0DtDSGnBFrPzMyVyKI+eZtr
9p6LkJI6F4pWAh2bhTpJx9uiyPnp3W7Nug2MTq5qgYB1HxpLEpfVAR3mktTWfEXh
HU8tx1vpEkA8DpSSu9PWY+KjBfdjLEP+ktWCn6T3lj5ELwAPRtKxNgXiUWbFXsav
uw6Hx3OhScnlISqXj/YMbvvTqh5gHZLaOjWjgosDmXQBQrDB8YbAHW2fnaGplEjc
r2mgxyDgbn0FqGhXQ9E6wvlLAQrJx3z+255JUuf6lG7s0lZ+VCGYwDtm/yYRn1mq
GsAq6mLXbWq8uuQcRQc1Gb/z85yzMXDPMfh3jJlu1r9bWQu1QJme69Xn5ym93G2O
wY8+cOa3foXBSOknROaTJeU3h4ZpYHOsSN2xioP9zyoA+vIXmdfWoqSHNTfHNVWf
Od2ar4BoKyFBMyfUWjl9x6sv4EbRdj/Z0oXJTnD8iFa81KOhqbmkRqg0ivDnDXls
U7p9yuagQ1sSg/RECzt9MIXiI/cdQoRfTW4iZZvXEOR5YfoQfrPTD4zqHDBiK9bg
33HRPmXTcpHEbiInRWBu4HXFWobssKx2gWpGB1X9yhl8zbK/tIw1tTf9MPrUwcA7
773fMM/Bc+mRPFhdBQQN2/W/GVL5n4TDCh9oDkRiaSkxuxujXMGqHfa8mOyXoJjv
86QO++jF9WLn9TimH5K85/I65wYnutHoCuvN3J7x3g1TfXvUw95B/tamqv4eBqnK
+n/kHixkzWuV5CJmJu6jcahYCcjUeXg0KqoepJVKTvII5QQ1v8P9d/92h/hx4TQ4
8+3GSZZm3if1E4roquNwdF2vitVu7uKTqPN38gXrMdJpF/oMOTk5WBG0EbXSDalQ
FN+VVRp9eyRVAQaggH8rJHgq/NLTkEEIXAGnVMK9mHtLjkq1cCRE8diLOdulxfCH
mdaR7r2u7vinxd+vzMaKJ5dHWGFaNYt3q0GM6fMN1CU1c7okWjfhEA5q8f1aCqGZ
s496Bh3vqVHSKH6oxZDpaafiDqB+EshaWrj9SvK0wiIBr5NnSew95sZgHRNq/zbW
jkBbgDsWIjdFA8ZpjvUzUQHWL3VFPm36u0+IoHf7fOntDGj+QXwP6pw4atCsII9H
4K5ZoaKubwu/4S/e9kIKK8viihrv5NpPZMAOb57YWsGCd0iH6CiRVCjBMAdU3KoV
Q1jH6GMrE4tgTQzZ+/HTjMRjC89xHd9Smxns8pBLWeLk2jqxm9xn/4HOZLTztU9+
TSxCazArN2UPSk/aScHDSUWBxV8MauWEQTKho25SGeeLiOdP9zP5sE/pEhfdGaT2
Q69nFSCgK3G5wG4Wa+MnNMACssfqh4Md1fZ0RjaRAr+07syD/fqJdS2va/vUoByn
qprL3ZsXjmKG9iOyw/CjBpk0y9aENJGrSNFwoUncEPqONuXEaY4TXbsiLH6pgI7N
kzKBWbP727yJvHzrX8ZPOa7Dtp3PNlBMd/oTWvWfq9zZuBoxDzfhpgdI5Lrubqqt
CtCXz7LMx06hZw28ez6UhdWPAYEG+hm0t0XNPpHyhTgUhO72ghDqjJLFN7ON2jtT
BmKtltmpY5eNHFBVV0E4UrZSZxZRPooljIY61x547MqrYh//sVsTs4FDvZRivXVU
jWy3FhVLyH+Xs0DqJi6fy4bMQvV1kUyqitW5GpNK0j04WK+N62BOkfzk8UAcg9iZ
V/aZsucqRqF4w2CjhSAUhooHZOS5HX2XY/h6VcrfOkA4ia4QNunnA/UeYZfhbRdW
sGd4xcPl6W3Jk7qsLYYCRza00fOUDWemvL9gdrLi846i8nv9e1Zj9M6hJDiIbKAD
VOiNpmtG+7TPpzqYORwbv6bDSQxsQoDA1ijEs7QV9Lqy084Ab/MPjUWBRi0exJdw
FesyN0bjsNXVOwAQGeWlz4xW9CVPxNN04iAl2Ibsd3QCF9YRwKb95ocH316rbxW+
osYfsW1+HUpaZSUaeNdPKUfXUx3zFx+AAT1r13udzvbYedaxN7MJXnndDfxvboO/
gOoUXWIui2iQjSAKXXjg45QpHKhrM+EutmIfLZaRj8NYBXEf6ZAtCdqMrlQWg7G7
aN3qxABkcpucs5DWTHEHojdCCrSS/2moH+HKrC+7UKp5E/+7ScIPWf5OvlypR04y
+VNqA2/wA9sY9ox5964VKIdcEal0doyuCyrE61csnXMCUxDYrarUTxars79IKsj4
eambI2puntUVhhLXTSqiz5KHwOWztKGaASrGRjjV9tWrLlxVOkZsK3Q5mV2C/6cG
+YqwtkY8fig7SFeufss+ztts7CgN0tndmR1HUt1YcClnyIoXi2plpppPS5aYGpPO
KClqy9wXYf0QC8WXArEw24tCl9/p9YKME7CtmaYe0jOrHVMxPCVWkRBJCiDomaxi
l1vn0u2GioRDBk1bfYsGnn2nVyEHV2GM0/KFWN6LpKZcKB8zonlAjkw46+p3xVSj
WSiQkWVFSpgYnkWFAyiZbCoOQHqnc5AuW5La5L3Llpzk6hw5jEHrRN5Vn39tfzHp
E7XyUcI9ruy5tfZxexTSz6fcM3UCiMXiakk2ogyE3eHGTzarqjbLWsgu+oXadXGP
40O/7yGOIukf+mHMz5dwoWoAGczBvw93SinDp55jJlFRVPyS/A9IPIkDMOfviO6K
GYBFaGckpSP+OWumB9bko1jbiEIMgF+aCFgHk2zHbV6j2pfkK9NNEM7PEghbf5Yz
THz2HhHbZYO4nlK/XI2ZT+/U4Ak0FZpTLhBV3nk3/RtwLCZlzf5aj8FEv4u2RxUX
PCqLfHU0zXbavaJEjRXbAsoILGJPgXZg0OyyV0PNifH1hQeW+Bdbtmle1nw4iifM
TWBND4y2zM/XEI3+v7dngHJGjqV2n6TAGu+ojnVPbyAUU+/iaFUFRjivLp/gR1lT
UZRqwxCiYflxlRCILhaeDMWM4LjU4V2gEOY+IDhumTc/A1kL7M0tMRQMToDZ5jRC
WXwreWjFqqLRAmDK2/SyhjzjFCsT3J5a8Ygy/DrPneZbJ89Zx3Ngv5haL12GYdyH
kJf46lkpiMpSCaJOOvvkNNXSi2Wrhtr88fKM1jncrPy1W8HS7/8gWJ7qu9rNbc83
TnT4gouAhyNkZEvhigqYNpK5fwAQ9CQZC01wDCJuiAs3QK5tfEhfBjC5BfGhZHw+
p6Xi7VVjj8F9Uta6J1aXtPgnZHbAycrm5ZYSSjavYjEGpDUpxvs1Sp6XWLJd3zEF
/a5GWFUmMjf/UOSwac5QCp8tYWhiGgEZy8R3L7ndBUEGQkmnn+pd4w/qAvHtgftR
pEtsr0X5J61vKHWWulvkMLFefycJdvhMpmliVpip6Q67o2+IcQuRyS67tuUvVQyO
mHob/vZcjNgGXmioHv5KOaLu/jqIxWKCLFJj+ObQnEtbP+AZecavYvTnjB6hDVP/
V1gpkL8PFZbHdiQKQIZZovb7vabR/ZKVC4rHBQ7TwL+/ImlD6V6DjH1SqgB0vN89
tk6MVTgS76WGZ+5TxaML3KU1xcoRlZOeaJvSXDvQwNqS1eCvHVZcOc7CFNMfAUby
liS2jsAspllXNpUZTnpMG80hnhwfnDGEezxwJrjojPiorDsmFcblobgGhB90BFbj
Qq+EZQ2gnFXXqQ24hBCRwWl6v8AEkWvPUSprEuEhdhJs3BIOwSm+7SQuIVVn7M4f
Q/NBXaNZ5LNbVArjxW8pKLfzu8P8MSio2tZPcd678alQjvaug4PweG3EiJ6y8jxm
8nNG0NQY0gep0rnNdlRUHw6BpqrXqlt1h6gJcuhY5WEBuof2svWd5ky3VM8eB6im
FGea9/JPHW51FHlLD7u1i9UAyOewt03FF6ONUD4J1w5DrGB7oebGraKkwi8nJaK/
7+kgMbJkrdJxMCgpS0Y2xWdbP9bT67P0Nz6kBlyqxM71GIb9SBHI68ChuVjFbczo
VH2/U4OdDxZrsRjjmDhdJnrj8SPtX/Irq+KB2ppoOBvZH6JcNO3HlOpBTGuQoirM
8wB4DZP1QKXoWNnu9zLGAjoB/kGuJbu1t6mks1b9o5bmkTlIWZE1NNxF9vd4zwql
SJSgoTjJ7DagjH0ZkFexv/LZ9SE05e7IwqnsDNOQdJBR1aLLf4P83zpxtcAv16qk
VVcVrttyLiMJz5MCfeubzyXzKe9QaFuj1Vn/xqFgvM2G5Ds4MSrQtYp9Qt4aguiB
rJwXcncXtBAnREC5IaBWR2XOFF6gN7QcLjUBfXobYd2oYLeYMEM7p7/Id6bHAyb9
BAvHCy3wTmeg6Gr4v1A0Brfu9v0BrW729QVOttSa/DSICrdHXrww0u6APYPhX3ML
k/fGDlcp9YZvfHrqVi3/b4FKxvNKgHZiIlDDLn31R9hoWb3m8aXHEbBiVQ954Xk5
Rowo9cHyZpXYnfCLyUJqeBxlm/8r3bkpkhWQHJ+TT8aaAra4GtNvM4cTitM593yC
plvIcHU/59yFuhW4AyFJgrYeGXxY8oi7IEHHBunw0diETNJga3gLkYYZPgDWraf9
ZaGRqCytgFwPuODHLlrPlo+A2kR0PruSbR1BdFi200Kam2wXZV77ahWRqnmENm8L
5xjKk2yleyiY79GnXeOZF5Y3bEzO5G4I2/2SZhv+8JuO1DN/a9B2pc+3vs9vMUIw
S8R/ADtuABs2LQbGJvF6LvzjTJcJxqxMHF32H03KnlRQMHABP5rDBb3H96MOPwqZ
PFl2rW4/F9xW1peabPz7gBH/rSHbBl1Vrkq3OYeyS1rZ2PnpFiK73z9pfL1lHNxX
JIHi/w919CbKOvphvf5AvY1bN+SyWpVnIoS8bwNbCxMDBvaaDCVFnd3CPDTrNSC2
aaUgMG276TRzuceJE/IQXveOyske7CVxo8WrAXS3VWLENwLoQTOhlUc0CxD9enr1
MrWtrGFFvDEzhyD9IjegTAbxHlBTQUuTV6asIqNaM84aLbMbCtxPL6C0P+LROFWh
+gBEIBYzZaoc1BCpH2UAV7tMU4xYukRCMl9DeJYNtQlwdDwBBGQcpgnUjJk+ZdSb
LdkuvE16WwX9jAVOX3mjUUJif1c7/kaO3bdx8eXR9/rTUtD/R4JiRIKAPleFjM6H
nQEc8kLSbYtfeZBkY9p5A/g7ZL0PXH8dnFBW+hNvt5zEFfehFRgi1QExSu3m+OK1
nXeHF+veW28mRl+SHWCwdYeJNrFHzp8OiYEgNWxuPCfrltaTsNPs30jiQt1HSFTF
4lAhN6v3/08dq4nM6stVPY7Gs45iJWprY8Qr2foIoGF80/xbjWjROo0VhGKPMa9V
fMZ/h4qfjVAHyUZrfw5HNnbBwrtRMy1FHcHG1kUR1A/4XhCvuY6ekUgKh1n10VUh
morO8VEhAVAxhgIgZWmTue7eSxggtuXOtZgDqhFBNtgA2VanCklPPspvbyAWxgqQ
sMABxMOjyc5OcDqplKze/pKoXp8U7dqs59gHWetLf/MCJrjKaiiqRI7Vs5E02c73
bylmSAbyXXv6cDbMMgo0fsjR3swU/ziweyETtvE8ZmSep7EK+/mcdHxZgjwQWtHY
na2tqOUWPzPWExHb2ro+2I+UneXS13Gi8AlDlAoBfPb4Kmvm28VVaeLygCoTsopJ
BXBTXNzsl3tbseqaWuPYKNiK+oWlisMt9v1zEfvUt/vdPxRUG/xex00Hdr4b803i
fooFA/F+b5YqYMSORBplY4uK1GpI2CTHFmEgrBAcGZGt48yF37PFKWmKPVRjrygS
8GZRdsl0VQlLN3eRStqQt3dKDisl2UB9FXlGS5NF0HHFo7A6FIAAtglh/XnohzHO
SuSPJYCh45SaZ0z4bRQeRvui767iw+IvXw3phrnzEBurtsgWmTD8ICydNJf67QZE
RsP+0jexgIQuiVDZrR9EZT4wP0mnh9YC1YgC+5DN1q72+9v0VDrzXOK98WSAUM0h
K9jEoDgxVC9uYoXMSsCSRayeRHdR+q7CUqvVZoatZiiZTkMthM2znCsqEN/GLPv+
fNLZKgF8qxcVl0m8xA9nDkmqD2gG5Ubh2DAUcZ5LcBoNK9lXS2z0tUAiCjK/YKix
skkH4ZepMKg8lZD92gC4Pcg7/KsFhUQWBRl+3M2ozS1vg0tmqrSHlLneC3dQudxY
+yjjwdj6t/GZiyCWbZvDuFK09SYHsD2TrsLlKQFM7Yh9xV0qxl1OGWZdgR5snB71
7G9bpBWqsLpQPbVir1ZwpS8jNFDOD5TVD84Z7tJw1g8Gli0I06M1Wl3r8wOiYCKH
SpFGSwOE9l7Nne/JQHrAp2DeIO5zy1aNPQHua2avt8unqm+kH9mpcd/4gNuP0baj
VU3YVGdGdn3kAkRfW6zu1eee//jSgTvAcfPlJQ/X9UhblhfsjflSNJijX+Jn8POy
XAGsJ9xHNqdYAQAIZKWYdYR/cBJfAhu2A0eRWPDIKCNoHRcDfXlExk1y+d2saN6k
tLdL7XJ4Ay4hscsl79KNy6hlnuSyG9qmoQ+m9K797J+dsp4/MOuH1FjE14D028qw
wJXHVoLQmOpgppbkB9rEFHvs2+BUHGJK+FNWXJZWbnNzmSS2bhQrN5q6G80sdmFP
ooS4Cbrl4otHdIAUAEfrDe81C9boUoTjilHwY+RFfZJb9/HaGKn+keAKcBHlEd1V
ge/of3mP9lR8X3y/Q/ze9QDGqnIryeqsfDO0AW0VB9r3K5FVzTfyCuPQ1M79v2qZ
0wvilh+r+mxME5MCqcuplLjK8WPKLLCUA9Bet3NzDp+ZoPi5aaUjC7eVAcWnJ4mH
WNPVSnCicpJZqPc+wixIIlXy8tQXkL77am4JRaMAJjFLNOSrHpoFeaObDzp2J6Dg
R1N/mx+jti1UzF+2mdyWkxslh5kJ4EI/DaZgiSx9+KMvy4Klixz3WTHigS+kcZ4P
MK5DAqXkwDffROK25ydqnLpb7ogAkvsmzQiIcgABtffjgsDNceOcEKDyLPR5faid
JK9n77bTjQgQ3jEpK1pGy96c2qKL8YiTyuD+4nodj5xaQi/axCTS1tf/zAcUYnXW
u89laVMI616a77454/wJqIlSyesftBEJNGGx9HdF93KOX95iKSWq7JfeQYRksNwq
w7GXuknfit9vLeK+YC4X4gNxLk06hg6xzE35nB8MEi/mMFgKDYRJSmyBGXLEYDDo
ttzUBuxzxZyAld2WX1PuWeS55SIHgayaiZCkbK5IePgNmO8DG4alu3rgrYWMKLVK
QDO5aiICQkUW7Y2BljYFUtujbFC5WTRklkRPZelryWcxLA3KWKc1PKvq9dZam1UB
FEoOTr8Up8nBwfKo3N4XG2nMi6OtI8VlyaK+JMRJGyp28Fku29KFPFSfOHznS1Mi
W8CLSclfZ0zsGYuzDc9MVgq61yGCU5GHr/0rPKYBEdiEjq7+3y2y26iFbX1z0NPK
iq2K6Id6OYkLiq6OcEkgoEkfh8zUuXt4abrsedf6yGqFaOmgElYjk9zX7+I0W+oa
5YByiZllmSssiSMpXWD8qNTT6Y7w4dlAMA73sEDj9Zbjg1k5R6LHwVxc8+ETgvlN
WwogONsSci/XXvE59GB1BjdnUb0USXwbcZuTd2JkyBXDoWhWkwhhoxybQMDqbttP
3/wpSD/vxkOMIWtaWHyo3sj9BiKwfm98jVkfqMcKTPN2IaEfncDH5EPryLsgWs6a
WEF/NCxYCZbPxMfqoymaFVjo2ih0i/CPQ8egkz8HTxGGNOxCsfEwhzJb2rJmx7zG
7dDoxXVMgMGPpXZ4pSynIxFJBURlJefH5PMVZCZwcXMdX5vYy/5AvL0FxgylIVzF
orO3glcP/AHe2DpCuiXfi+TZDCNz0G9PV67FfjONrnq631gZ8AZ9JGveBcxlATxr
X82Lgu0Mh1QdR7yGDLTck74NGEKhuepuWaRLrMQHp/dLDSiVzghjSLs0+sDUwgPU
py44OGn+VOry9W0sjPpo9pHnmoCQ9aQr5XrDOatxOJgZPzm5sLdzgX9PySFFpQZ8
oXyNHhWN74JfefM6X4dmwzTemDFeNwO36lKLq4aLFfXs2e8v4vCaKU7sOLnAvLry
0UFBabZdiGxOVaxJ8HU9WaVzaMjkENAvN2a3VCZNeKk2T3zXP0k0Tyju0PgvCSNH
VeJS7+6/fvO7B7yBMyE9wmyYSSdkDGGu6iyIl4tg9rzY+/La6VoNzoW46jZ8kbXp
Np1g9V+RY1gEVqubxFuJBgz4fVoFL+BDQxRJhcNHDAMO+MmrHnT21Kw62A+Xexxv
eegFcbvpUvZZHljC3FS4oe4FiRxQ04xq/SL5vp7gVOlCmcQVqIu1aJgF0zZ+IRs5
JTY5Bhegl7NKbGH/lGYyDEklxp9OsGD6YzFVRV8JFYi9Kk03vB4eckyI0W0+78xl
onHsDJC8g1KkB8P0mvIXiga7vNT0rLOLTzfJO6GBilE09oLYTSUCz1T57UeEKGjK
r9vE8PKWpYU3cGJA3kXEkzExbqW0bO2qJLFdY9q0ji2kUTk/PoxUvhA8gHe/D7jS
WHzz8EkiyjuwusDD/56FYcWlisyD9vhJSfllRnFpYqp3PLGf4p7DK+MSINDrBFDd
yhX221bDZ8ft7XGQISezOV1YWAW53O60KKbf0zseGoIPO479aD1BFYlkmjitvnfr
4te+PTjMBTEqSkpi7sH7uGFbzaXRGOM6WYv6O1cPoS2p13bROSaQ9E8gv6/stEPC
SjUvTUBZuQUJkWJ4NV9/YV5dRV9ckdeD2kC0sPoeskyzZ/O8HCSrtk+tOSAAyQLj
3VazLut7S7Z36+aZTZ1S+jmdPInb0EhPkETG4kPchuFkTN+lgfinb4eHBUft7YE7
OIER3B2wVZdMaGSTmlMLD7MCEGumq2a9Ygib4xgLFV40vj5sYFBgWYxqrtbOVS/K
yVUwN66kfFO0eouVylHDsuNl+rC1uTYirB8tDrm7qQWOgjeCZkFxvkmdZpACLhiQ
pFEm/FPAASng8tjy6/jhX1tiqCR+E3leVTwGxUy8bKDaQEMqxa4GiXWsEH230bw5
pnGVozgDlpyWlqoFxQ6TQhRYtm4CZ3ebzs14aiWhoKbBWUFcOY33pUq+7zpF1C2H
sYC3iJisgpQk8OS+0qgdCOdSWV6J04YLBzIHVWD3i3EjwzzDgvlr7WT0v2Hzk62b
J9G2rnpDt/W1uNcj/hM0bFSG/xhAQQYp2y9UvtDwEQjfx/wTDVeXuUGr5RtC8+/T
IcyXSwJR8EYDCvcdPz/cn3PHNNB347P9FWjNR1DOBbwCcgqQk2A1wGBDtFyUUkTJ
E9p6Q25Lg/GCQ1M1Y6ao9a0DmKDbSB4o5hNkdEeKXMu8E2wx31VHT8IGVmeResw+
YZx5LZp7uKGaXQEofYX7a69krez/5dSmIw/0CYoBTBuJYz+dgTD1Au+Ftu8slSTa
CrqYgivhovxSJkuAkQQgS2/qJaXNLpizeVAtBw1B+C3vYCKQrSO/qr3VspFU2sty
IyshNSc7IgENTvU/sIK0IrNiyG5yT9awMjBYn9zOu609Tpv+aaSH3WJTcmezdNPD
QTUzYASB5Gd+C1Qiw1eno3U1DijevrreLJHVUMZTzuPlkcshM7HJNpGGBP7j+2ym
HCpM/k8I86oBDWiARwVGUBFjhKLY5de9y0sO5BGfD32DH9Neu6XO13QjB1JdUr8L
p39NGGCZifLkjLt4up5VrOsRxen+16LDiZyqHBwhWEbIYEYeCuvFyUU4y/7YOEHr
TqF9VQcDZsNDrI2LZ3U/D9Os23miXJK9kkEe4ejNO0sFhjqVqfGUxVVFJtXnKH50
kuQHvy89HuVGbPFmcpDipnnRpX0a4s9CgVSEUtQWZsybLq6RQkxdSSPZVCT35jba
T8MknNmHkIgCMzINJQeTwsg6YmAayHQ2LjFEZ0u17oSfZJOZM06PdoxFN+jV1K/T
MJYDR9oKziCxAk2hhpRKKAW0GbFaqZY4yQfWdXuxaoIYqYUFFnVWm9M98pC6rEZY
CJ+hZqG6MTY343VDd8Kae2jr4ibb+E5x1wcwYV+1GU3Tg8FS2E5W9GeTHiyYODN+
+GaSYTYxECZvmV+AGnYbvNwf0g164UljQR9zKdmbxIMEcwmfrSor3a2+DcfZFDar
35u+lk/n0R33qdBz1glwmnkqJEIdYTXyrGFP6f44QRPdNlj54y9hBRK0BM3yiNVi
D9iAS/0EMfXlwIrLJl9NsMMFUTVoQTasBmOVLNXxFvudTBBDW95QSfXEyi6rQKAS
OL9dOwEJ7kWUdwqBmOcLxByKKJOenkoNA0fWyd2y5ummm64vJMRP3UxLHw8qyCTC
pH0w5z35hwD6T8je6hcduEz4Ol2QRbXjFGKqgn2EounX7J5AVMHi9cucs3fF78EL
QdO+B9HMyZVTPuDDrsZXFwRCQS/ZqSQFiR5NaU7DL9sAV2alONAkQr/IJ70P3OD2
RIHaGqtdAZ3ZPQg602WWypvdSghgROYLeobKRGWqyfN9YTrxVnjGjpzTDdPvVHq+
CDToQXS12ZeaSBFGtCloHv0bwTTXljG2rAy7r/t+BEIzPd44AQczEl0UWWeoZk0P
AWmnLiNs+aS5yduBZMK/+Vx4Kp59Yhrz19vxxFFk5ddccjhg15RwxQc+5kKeJU28
RUpzLX0tuiqkDUzwjMT11SubhysPbIr2AhUVNY3WpzklIeEOnJAsj0QuBhdXFpsv
t9TYHNKcOs528JiO3UfncOXFNVsyrYm6t5bYkQK45Yu5P0IzpmjmzV32h26NiisG
J86sygTaSlwQxErVqHBN1ztle7h48beohBjadB1r/+J2tgQoyeg8Ow0pwtxUMiDb
BTOV5BbHxju/vjOFbpcNrf5WV5kYSlHx6P8OxfFAoq1yjZR/jTSDVOe3NUi1r4kT
OWMl3A215iaMGyUrzVhofDKMyPhFZ1VMw5XxYTtROy9JgFdJ174OTpdJgt46lgBU
9YtwEYpzcTaBWce58wCmEATR6GvhprcCchsYNQTYO1bOzPP1T25e9huJB22Rkpjo
+F7aZK4GXN7u8QjiNI1+PC0hGefoBNV+X0JLb8JGtdPp7eYRqld3NsY0g6ZcimDF
6lKcfyaTWqYCUZvRcjGO4QPEPvurEoker+h+rNgC3Q23+GENm9shBPOCu8istY93
l96ZIfDtzmntfKR/zMUQlGpKTPHHBQoAh1SlZwfTB/ucWyTnDk3KpBVJ5JOxlKg4
DHYufkCEhEqb29SyYEO3ikL/BWsOnFlMqnQXqjgWnnCnpb9rIkZ5mT8uIbHcp+fp
rR10E6TyoFShCiIw/9tAhkAtEVOt1uv0n4U2KmAy7iGXdnYwKuwThSN0d9UGJ+e3
euVRz6bI9sJftEv6ig6/N1qwOCTPq2y+9+cVHLWa30e++xByrAbMG8SRkhxQcSJF
VAYVhlMQgTTs9ieO+2+yI7Xq3io8GGY2KVQvcbMcI0fgZvbe7MDQfviqAe6Bu5mF
wmbq4/VQvz63rHTXG+NJRZf8Cl+DZHz53KDDaYn+EYgpQNINIzfHSRcRpa91a1sp
riDIfKMeinA7oRr78BYgj5VanDQxCY7vLvkE61/3P/i+aGvkWU7XpUrAshx4gBtW
LUnxXrgETXBZ1Xg/fH48WLZexeQYEQirwE7WmQWxo8axwTzSn7iTS+jwMLxvC6/l
IvVIJj2SZrJgvUE+Zb24TUyI3KnQa2zpo5T5XstAnLicCUsLeG7Y7tFhPRnwSnEw
Z+oNnznwp39h2dES128eoj1go1hccaTmYMNmbGLd1JAmiAs3NZGHShQFmwHb1x9Q
nVW5v0iaxJ/Ix+LWSGMaxwtekaSKonLcqfN7Jg+jPOm2K4bi77JRAYvj86k87rqO
2U6STNX1CACUcutneb19vSFOZ8UBvut11nSKUGvEynHnaZj96hUCfnRhh+4ye2E6
YE8UhtQczwPo0rMr3m6WRfwz1gmF8XwmqZYzGfrlEMsMmKYa9B610Jo+Z3iddynx
lBPf0JOBwRT99z7leeqaHwHRu05zMPFLZzvSi+eLNbQK1qRFPKYh/sMGFDMJ2zeg
vGjzXK+U2m4fyG/JAjcg8/ua2MGvuHrNyQNNuSikd5G9aE4j+HZcpBRl9x9NVMHb
o5v/RPnolz7kGyC4Uy2R4orjNPEAyTPZ173dammFSTfTeU+Ys++tJg+1KUMUPCrO
/5ymoTqGLSw0Zxg/jjJnfxPRyieZQpkgVjniWefA4MJb1rsX6vHifW+Lm9yKZgw6
CA/ber+C7k4SM0y3lJV1yc8W+NKqIqV3GVtj8fLrd0KfmReAC10TEn0LIOIk8xoT
BvxPWm8XxRhsRXLjUcsFFKmiQkNyJaUVk4QZLTlNiEOrL8YqkCrgMMVqnxf/iXWD
60nrReGb8zrTvwuEfUvJY9bmp2vsflh0FFyUuR9R8S9mjB250hwGW1gIxmAFkhcJ
XfKk2obu22wOzUahkWZC1t79BYvCP6EmlW01UH5mQLZ/Nr/Dw1JrrvHaEPShcZaT
1TuvMmMNTDqciqQfU5okDQqVbJiHs6rArQ5RFxmNa3pF+K8aalzB0jEpqpGzt3Os
6M/VlSrOI+38F8RE3gD+V+WUVmHJzpR7YDH3VGQ2DNxVVS3yffvalatW8NOYHGks
5Btcry+lwTwAqEqq4ub1ydVKhYh8YFx8HfmAzC7VsQArgdTils4m20y0/h4CB7IQ
8HFSZcHheo8BMyxAVQPK9zORg99wIMBnNQPWXK6S5Jk1N+LJG8M/hUCFiHteK5un
fsmLl5DA4A9G/awsVLYOJXRQwM48yDNDeD6UnVz0Z0aWW7rcTUT6GMceePKtoO0W
5e7tEnShlg8eqJLCMHs5/E+CH47gJW8tic1xIJZr+GyF3BXbaUnIzCmaiodfnuD1
1raSotfXKHtJgzrtBEDOvTcceuwXHVusuMhEQHTou9QYbuIWcWMrY3gmCGEkmYQp
oYdXVpbqEhyP67NZ7P+jMuxXhdEQ4heRdupRTxxMe5Ees6fWRn9YOISrQYI4Mino
4lDsnhdeW0+UoLKdb6/DJJTjR+3wVL6SVoiX0knBRX1AesuiouuD6zd05mO00iTf
AKC6/BYp3WFCod3bkTr59ipZrs1CuqiE3lLgms3NUPEhRWdUG5g4ApyMTTVB+Oiy
R8q3UfA3RVoPqcP8k5oGvq384wInI4Vd4ub5KX61RQ/Ee2AeKossRDTM938YNGdU
4Zqne8TORoUF9WcipWVqdGHq1vTCeweuxY5dVNnzOsUBTHkl5APxofhuoHaiYFFk
Y33bu0/kY62DUMXyoJZBuZAT1YbdCOC2MlvcRID8ydYpK6knxIIakHJAWt663Nun
tyQCiB/R0NX317Osy6R0DoS3iUX5xsVPN/AzoRThMzyZJUPFxuTrHCk4T22Oe1f+
pF8Fl5NbvxcmIA1Wv2ylJ5jpbE2+u57zh3R+vlho2bNaKzeXaN/cirSbHCyFd2Zk
HmNoFo02XqHfBgSQ3eVJNLrwI8/OHvRTNwUDH3AD6/bWdOzVspW40j21xuOuwB+e
fZi7RJY0OBifDZ6dd9n68Y2bB/vxBNOaT3wgxUrUsOvy0o323ndVK6mze8ZAURox
HtrAXRjre+x0+kcL00vNiJoQsqTDz5RtbtyT+Q5g/6A+be5mb1qtOg/c9SRBa8vW
srcYyyhs38I17+aLDnWGMdJsrM5RhhjnqfIHL2sdP7HRBcRCiMgsAspVB1Lgu0Gg
VLbMYFiuCbasW+978zNapd7bB44xu7vxKdFzdQvr/6pUVL+1RS87iOWWzisscKch
yIPLrziSITZQfZj7IEEDJsPCNTXM75QN/MEvHzscoplmNgbYWCEaegoGbn65LNII
wtG30rGWE5CkptOTZO9BBVsVo8LOTCWT/pxH8Q2W0XHIkSe4lHidKuH11+KoJ5IM
X5Z+advJ1wDPDsCjYomkRZY86giHYtO50lEXM+Aa6JMwqEprOV6A6t7WP7d1KuMD
2KqKbtHwU/bMoavdSe2xu7YWKbMyYUYtljmgtxiBE5EgkxQSIdMIrPSUZbn1a1R7
X4Jp7eM3G2ZGJW479DL/xe+aTq3WlZFEQ9v1zlasburkjxvsEnxa0EtfyiQ+G+Qd
3nDggiKE9bPDBuua5eS44hntfPn9yWdB3ZzHKYjOUEnKWDP0pGStNWj1cb55XPM/
zfcx4Ne7oSex3nObp5VVQvN9Xke0pOWZ8a0MMcP2KVXiYvruhRly3/A+2SbhoZVm
3nbuJ11OoJiHwujY4uuvp3y/6/6QKXhZtEa2XkEzTTn+n+JnVciYfH+otgSPXR2a
y1YiTQeFSq6rnhDgPw2B/u9VET1Pq+6PzYeC8MNpMo2ybLwQvqyKXIsRHJ1ScLhr
VkHCZ5A3vvPd5iiALONBDdxXgwaPQkEpjZIp/mbEMTbi9GwzmS8FY1I2cHxU6vb1
r5LI2o1NLAwoP0o3EmTSgNdJTQtEQHCnY3vVBoj8yrwT3cE/XT/Q5X5Vj6m+VU0R
35F6+iTHN2mWH7BNpQVDmubGPcYAP+EDf6/5CM0RTHdoUNIcs7ItYF1ODikjplua
Fe+/7zNDuh4BNfVgH9UDYENBmEuTrLQBo8HGI5ZTcwTLpvHYRhzrh9cHWSlBcAXM
v4fjWqI491PzQqKBCdjBJd7OtDZIFlNPNKA0wYX51osrs8pJ0F83Fg71wcj/RYFU
+3LiBpv/ezAVWdnkeNEnUPvCCGCCXS8a5rA8UAscrBT92fQ5IScZZbK1zanq/gh4
LRt6CspTX72Cs2S+Z06aVIkNnSAVTkTah8p2tESqkhApw6WjqvNxvll3IxozoaFd
XfBwDaBE4O3Qcj8brxHuvfVb9YaJ26XWcNloFrmbk7GZoCJNoznFJVgcOfKqwt5r
aMkX6Q0Ey2EJFZKGQl/k6SlK3IdZRoUn9VP40N3ZQB0/p6dlMHjdecKd9SCV1i9E
6y++TZop5UHKeG5GoumAge0nlcJ4Q+eAdq9E1mPN7Q/tzH8E0ndVDLfMp50KqRog
w1QL2fj9f9w4xMEMePFpDJe+VTW8UQ+nRaF/ZL3cBF600W8+4jOcjb0LeaUXdimS
/MW9y1HHwkv5Zifnlh7cJwabVZjD+EG1bT+Crsk7NWBa8vtKXPLX4XQrFooXrtda
x3/YGEHCxFyvg+fhsbhjJYrPkAJeD8qmcRnIwNZy4RDyiLmNtOJMeKzIy21pJhFI
rnFNbMfH0w1zDsvd/yhGTgczpZSGAAKMyA49b6XKzyu6CKjYC8VwU5VhMRy7f4NV
SqkdZumNoUdogt6MyTrd+TMb9bbEvHg/vEnytW6rpYL0Y3ax80TOnryuTsMFnzpJ
i6KB6SBnt+LwD8+b8oj9vvdPArJLo7AnKYzs2SzT0wNEpYYxKmyQ9KA/JcYiGu2F
gwyvZ7D8EZXEg0NPBA8gaoCeKVFDAED3z0goaA2M4tJo/rMfFjqt5jYk+SeBWCzW
RLLdlsrZz8AQterXeF8R9sCyhR4dJoiV+yDO7pubVP/w0GD5pnfCRr8fCcVTjo4M
WMZuDMBtp6V1bPDFpXDc+dd8bIXj3wpVbXuSo7rHYVqduPBrF28X2JQ6IvkXx15A
PK12ClzGM38tbi3wzzG6EzjIWQujttwiPHVX9Z2nsBA7+u1oK66XDHmFHwkWV45f
mjb3m/QteYR+NxhTMbK4cD7l4QU/gISMjD6TXquR5gphO78y+U8biozq3DL1oAk4
oIQYaLFRXp2ZB2xi23qMuLafSeuPOv4AgGpFagU1fbKKroq0RHcQnsfvM3ByAOp7
25b8rB86nvQDks4U2klAbyvs6SVlgN6HHErHfvBs23BstEtmuSWh7MMAOkofPUxL
zT8IHqglOAzd+exeTsirGRwbqBA1YQKSQnfjwlNT8RoJ3kCmYMY18RSbCmQYFITi
4/8L9xWesDfE2p+E7QYKTZvVLlF9iS82dN5vY3uHKGommB43K3ULA8io79M28HnJ
2tX4se+Dl3WpMVppDZAZ3KWb+93lUnjD+fCDQDymYn1QtskVcU08UhdOTO9SiOxp
hX1feH6tCTGuWVhBZ0+XgeS4aXfgjasweo+Q+w9qma/s/iImsFuRvtb2SO1kC/95
CFymQwT/Tm+0j3rV8+D06efkzFrB14NS9P6HXKv8HS96+jEm4c37Tr3o5l1sI4V5
CzS46tfNK8Kiy7CEeu9bPBZvuQIO54bw1z3ZIJh25O23DzJMa8qBnisBUrAdGrd+
tcUqqPtVZGFhLSoqPv1wNNDM37zkNEmqbiuhSOzEz7tZ4BWVhvL4y4LoT0fduk3o
NijEImLdvgRlCWcUIPZWBQQT1O1VTb1nO8w2VZ/1mSmOCgbltbRAzfTA6rNf31PZ
vKVc1SpJvN1XNFM+CZCoJkondc3bLXYV/pFtuX4/X9cPqFe0x2mau6ANoqcNcKXp
JtTzEM2OtVN5Qx7zvK9urJLlytiaM3SbsaAysn5R3KfnmU5m2Zp+i/RdJufxhKt8
dkn5B0R776HgcEUlZ8OcCvQRPqaQ7PbLZ7Oc/iEQhTAJS+e9vKK8L71QEiisd8Vd
BNuOjEURcc+YVFZsWEjVlbzxTFOab4ZxXUukcVPOi7dpVnnHnV1niULuE5GsgVp5
7hp4F5brmmHkC3NUaFV6YZIKMNK41GxInXTNy/1CT0BONxLNTNNuiOy+djEgz0cA
sU7mCGkRsgIt9fS4adp/mvA8Wvk1pNIFuBw7X/WSNngIGrjl6MQrSUvje0lx1NQV
Mloc2H0s5yxh4O8tneemhkQQ/rSVYNRemJMUXZJzgAGpvSeD2oP2uK9U2k3GQs1+
11SoRmcdr7rVujs1eA2/oSMhAEIEXeye5SjJX42QvZdnFAjIOnMYSU4FxQv528DL
haruWFYi4yefoRU3AbYSD9b3BbYttLt6DM6wVSnfQgZ040zGEOFA4HmueVWvQ7rC
4Yfspr7/dnwpHP1Kne7HkEsgRjIOHNLlVW+sVGwBXz+BKQCHZ77KdcVDf7MK67rR
Vc2j5YZ8+wdfGVY4GRVy0VLK47ONg5YaMGxA4W2TQiN4bzJiIylSSbw19JBHOeAb
ux8q5nGCqTnI7p2Kj+oc0jyrm6D0BaLSHy3qVE6y6VTeZmc+FrPxPz1Lu4BTYocK
lJG3EeQkfRNZAbzLp6k5B1QaRXu+0kGPgQDyWMjc/9rXU9sdswkRRG/whR/IBDaA
UnTZwOYs9Goq4UHQ9kPbm0Ldlytsrbw8gu/VbZq3gUmC2V66HaChtEgRmeyGD6FE
IdXMe6pKGle4b7KF1oiLRZ5tEOpEvpJVeCbNsNP7xFFoVlQHYKlcRbexcegfa4a6
V4v3ZuVf/1Z/yVRV3Vsehn1NR81k79zpkIrUyKxFp78EkIenFOOHYR3sVboD0dde
ljMPZ6b6EqDpCG+Dvriu/LeBs2KxFGxq0lLlZAAJv48eadwo554nQYorxH4hx6H8
tWzwgtn11LGgZ1rVsAQjurKWCkV3ux8xuA7fp57Sud0FWovCfYCRv+6MPTCMMgoC
mAS7enh+YF5ljMO4Q5HCx0mpQ4pLA7A5rdq6aeWzFf+DVoN5C/docd5BgrRkYCT3
6jM4Y4BBp6FrobW3C5lnTBdR6Y49K1yuaUWyi96dM61qfa3kGXKcXkU2aHsOXWlY
IYJ0E4D7Zu918NuiH6zZA8+iUKvyfNy8LNzgTOhDAJKIWAYQ82KiC3Lg/Ud1VKM5
TiX+dwHt969FwjBLqOMsZlcGsaTH3WO2GmwAVkgI3pthMLCq+JJsMKgdDi0ksdu3
7aic0Lia/fuHD+Tyc9EYYkcJEeKRPoj4rAdp5kZYTYXO8kdNAHjZLGJKaCL78Y4t
HlugtYvS97Sj/QCQChEh6TI6lc3icy76rCbPii/kBh+rkdq/Oyy6B99FckzXaFpo
CcgVsOrbrz/brgVkQaYSl50SkSs/W6mt1B+/VxnxBeSCMOo1OGcWXnQLC/TtQ7NI
xadcgox0tSADCmM0c5qzxo0V89Ev3z6Ssy8YktKa7z5DjWnQd8/VViLFvDMnxIbe
D1RoNw52oLg2EWRLP6pqIZ4I/3K1MWQPqPmOQwE60MmdLp2fFPZiu6LdpAXgQyyf
JGnaEH1M0V11kMx4f+ctbAENM5K8LRDEUkh4Ql5j88lrpDK/a8NBC8YkFXfsyOUr
Ol8LICeNv8hOasNu8ANJcYkStHRNwN0/+iFY2gwuMtzAtKqzbW/TjFShQ4Jhgs2R
zMoezVFeoZpKYhU+IsHy+ezXK1TFmQZWYsU4qPedep2/VTO3uzNy6sofVET1j0Mo
/a0MQezMqRlJGy80gEpklw57wkjR7pSQjRIBcMhniPjRYoJ8C5bMnlJyowvZrF74
n7Im3ilCnR5xJccEYXKPgZzZxJ0631JhNAn98ZovDHtMkU5MZD0gql8blGyY9vmg
z/6IHWdt5RXvhnfP5Vv5v3iQWS+71GyKER2XiLgp2Vxn6x+b/sALmf7Req/0XzVy
eXjb0WpznIQRJt/gHYazTrJyXiQRebQlr49sU4UEdfh2Asx+B1TPE77M2UOwGzqU
hu3cOIEMfqzBDaoxrqMVadjSFpyvDchXq9s7N9ze5n1sg5rmSQLb9+A2dhQ1H3R7
4zW2+nUIE5UL8AscxqexyhAWo7YfTnFtiV+rc2K3wnx8aDKVUaHzYSdrO+r/rdMb
M8pSPyEWElxgY+qb6X6KIiGBUGmTG0ZB0C1q48AHReVA13luGUKJK8Zk56NC/ZOp
F0K6aD17tX33Z1q29jinnyOrz3ywf+DxeSJlmdsgIxmsb2Nq1mlF2wCN528m70By
tqggBrL0e5KF5WS3F+mVqwZsoTeTyvhLdZuSDVwCwa4vp0waNl9PK8kj1P499Bx7
cd4yfLfUNypy+nvOCDAMNqF/OfuJgP/xaEFH5jXb7hAHGdudFcIS5yi/93DeJ1SQ
EU1FSb2PEJ1q/34nlaZwM7aMpGZRv5ZFBuQEUeLTC0tywXPx1FQCfJ4PnYZXRGlk
kg9SyS7/GYKcBYhGpKqtbkKsW/HQGVOHV6DMthEo+dGgsZ8ryDDHXvqaD/wSrgtm
H5UVUT6+GDlpLCNxoG+cCSlanN6XqHFuhBdLpi2dYJB99yX4+rCysjmpUA1MhAuJ
NR4+itZ+eV7dIVQR9RgzNX1bqoroUWldrPxEEFyv0gRSqsmeNSRjfckEAE7J4eYq
cHVGhIkc03WO+rKr6WHWf7vDuQJrTpHFpJQvJpibkSXfIM4E7BD17ar6Ax22odar
gTg07hH83yFXKBdlU4AyE05wO76fGbhxrC9nOY6+hFmrEeRsgViMrFngS9vDsLz4
XBlDFfQeqdgBwhiNSM3pNYtoof7t1WllTg1O4AJtnk2kzJhBaZkJjw+JfxpvE/kw
K27OCJCIVfY0yVi4Lf4nCLHx4NHzZTOz8qLkwtiia0lI6tUiPmYgEppo5IA+omWr
Kx2Nc/k9hw6oPTt83HNfErvSt1bGqXG1DKmFKbn+aKWKGW2RjPk70y+5V5zoMluR
gv+V7RS/YNvDIl1Z9sZnJi+S73XKPHJoE1xjKROcOpYMnaxlVWrXNA2shBVCf2IM
08kd/SA7y3hYBIbQO5vXatb/4+txPsCTE42JUGTTG42imgZqICyN8VX621UQa1gO
SCwzbUmZy9GzH/MKK7xLHadLOPvJ7B7577VHVPfpa+M0ImOgnndUDAxUI7Mmf3Js
6EpP0iL8pBzCG/Zg4NW8IrRrbk1YLwZvGnHMLhdi3s3GC2lqVxPwG3fU1mJ79A+5
YqrxlDiXYZaOnXVRDcjh8shjR+8wsy6dTM8lOhrgiYA3ifZ3Ullt0miLtdSVYxEX
gwECs94PIoPzznv9ucd7t3iT0VLHUqTANxziSaqwL5rqQRUjLLszg4RgeyDwJDrY
N8uBMlU6vrXyIXzPNKOkv6/Ijm6c0cRvP2NLd5wEongA5Z5bSeNj2K3AtvVnrMWG
muBBOxLjO8HP9HfrAAmEQ3FlxA4e7TcSkgD9V2QNB4YaCPzJZQmRJc97bPSOXqhk
Y1DvPAL0QFa4Di3x+BaLUXy05v3Y0239gFXVySgs3JGXUaQ6UU96sCogX9nxDo5b
Hh904RqdVnIMCvZ9wp/PlfCN+3YSXHHpGROmaOg6s5V5l30r0pXdh9ShBvzlYo+3
71Y95UfXO5Mn3ZOW7Ej2OQcEunT8AcdoSmeDR7SwaDdP5jB1PitEJn5Y4RYnGnQf
gLGFJFRaAwPckHuf+Df0ZZYcpTqkXsew2dUv3eSv3dpZ8biw8yIolKITdWmOg6zQ
MoVp1L1cj9pOD8+LZneDL8t2GTVkfhYdSbssoGh4FO8Rb6f6k39JotYJ+1ahjE4v
G6FDZbfgx+jRlaRQfNJhOuk6BnqZK9BbUKNfZYIy9pl6ap4OIW3cBK+fPEUUIqg+
bQ3KPGu0GE56IPiLc57eRMSJC21ftpAid1BkMrArv7gOaTX9ZQGqWCgfrqkdka41
32FBhpLf/XRwFybO8vxPk5HzHnG2ugSrdj4LMhzsLHH/Ietne/rpQeci2AELEE9E
dXAErerI+UCxq5V7E9XiRQs9dz9Xiy41jTecGr76oBmQd4DCxtrYSiBsNuq/yaOQ
zbwJPsEvlV+SY9C3h9cYeh5pJpDs9X0PJKGneoevwDdlTOwPV1k+Lv92QBbJ6duq
1JciTBxvA2nKoYk2c92NRquADHuwgr/G3Q+Z+fI70/7YscPnUBiomsTDtumhhhH2
2GTB3bW1hlS6N7TTQp9x30OdBXTjSXZudhA/PKzIrDrb7D0Ufv+yREg+HTi6fl8s
PaTTBepdhzyts00aTjmSkgi+JyZBT/jxzhaKlQAT2mDwYvpyWUtr/1G44jmNmwcj
+4zj7/RHs5t8gDnYTdkF3S6Z5wNtAhv+IkqsBIo4xSwD09eS1Lz/fLg2IXN50qg5
Hv6DfxaI7/vOKpA3QsLTuIIIm1p52iOBnBj89xAZdjss1Gzd+5ozM5+HKaJ4VytK
izTPLxryOU6M/Uz3VY+4yuzqDihFFubjeF4LUBVyqDz+I0+sH32+n8QEG1hcMFd3
0CmENd8mbyGu+jvaMb3HYSf0B5OWOMgzR0HKTj2cSRSRcu4z/0KjmLJAuh9MUgG5
wJS68np1uW+fFpnyS9Yx610J0dRKj8XVBnoE3XgJb6HnPZkefRvc64iXxY9QDpvV
/LvO9QxHxmJpnNxtuxswDCb/1zmqdYW/UMM+eg8uFP+ADg76H6sGkMEH1rpOperO
yPYeCEVfHr9YB+z3tPU9/9MdRb8EmIfBdnFE80HZNg2VV2xZFw9mkpPfYcI3R/4/
GgctjQA1b1DTu2jXs5mWGBhkj9jTd+vH4AhDzHwGWveylcQ5SvisIsSxREIOi8Kn
8wp/DGfiZdshLbtYiJtIM+7JnfuFMICatNJtDCCLEgsMONbt/ghCAnQAe2BabxR0
/R/0HZKWAhf+ecKOjCaooNrhzpPk1TOLFQoUloSr3lwPfwIfVFnU+qGFu9D+U5UZ
AbwZ18FwilOGk2oO06IybwI7hUENG9Z0q7DuQ6lKsya7FXpLeii/PbyvMcQLR6xM
SX5+39/z+ry5u8rXVhV8LVp81U/uVqBcH3BldxMfHXh8fMIY5mTjYjvUZnoa08fe
VkrpmDHll7XJ2mL94561Xw8TNXliKZdoVqSR7cXzLOMfVZ3VlyVF8VI5F1JUJxEX
kQtGLNHykD92Xw5i6PSE8nolzX5fzabJMV6V3AxHu51LEOF0vqLiWLFn3f8v6OL6
+m3zrLZKwEfqPYHKbMLS1a1P8JGz+a6r9JvSbKU5Fo5GPHfCKgIBZUhZ7g0mDlda
ebPmHe7fpGmL29rrzmuRtZnXM7qYnPjC4gKSPnOzZdiLAmPvJ3j7CQ73ERId3i5T
ARsHukoB2AGT/lAjVGD9i2AMjq7Sg3+aovPgTPZFhvIoMOI05SeMRkWOKPLpn3TS
tWOYhF3vbaYxGhaWpzdg4NrD3TBAMVqbhjGY0QxAxc3tAZn3GMnNu8uyJvHW7S++
b1XcXSH19FvyC6lrA3i3JU0UFO+djXGTMaQIjSFqleq4KyfwJNaNQZ9z4mWqa/UP
wERaF19NpnM5SPB3YqJ8yAdUtR6TotufU2z/+QWxRFgDr3RQ+RDrM5+MR0Gb866k
12BkcXcFj5eQLFtxnq8Qz0h9iOMZXG/AB8hGTa43a+7KGXPR+4jmGUqaQ4fzcO9p
6R0qTrbiSP4H+U/x+75znM3oBsfCyFJ70HqW2FJ8iHDCFzjQrt7jacF1UofuueeA
ogWYHkGX1NyKJ2rBvk6KAg2LcWjBsU6tGA2qQY2L1pqDqaabKQ5c8nZLlZwZlIVh
FQB4MebXQALACGPknwJtgE6AeMDBvsauZrC0/ecVocsjX8+vCCsDaL/v0J15jaZu
nXJTBzMy98sW74ijKf07XigkavnN4jIkjmdq4WzSZg6UwoHlpN5RIO7qTohD2Zjb
qTUJ58sPxuFDlFPE6dw9988oDX7vRg8Ujyn3ffl7pFz2Je6gcvc/mJG8HUrWWVEZ
t7uBFR3Y1mzat5DBsHRyJLLRO1IUES4xIF8Q6lgxHy3LRfBD3TUGZSFcz6L2RmC1
xatOf8DlaFTbI0uAsn5/ggw6SpG2zptZo+g6QeE2yesQVwzzkmp9v+VKv3PLMsX/
Z0QyyebzfR7r+HqG2sb2QsBs8LU/nQxVpdYzvejsKDK68Qr5tc/csY5Ob+HmLwSN
0Vou3ccrO/AftN4FSQ3yK8x25NYgLbB5yPFl/ia6yAaQVFk93kNYC+eBMPro2Owg
0jix7GQ3P/SgRP5h3mJheY9n6ydW/9JhtATg5Xmn7HHrCboM4DEqhcTj3wVdaHOz
VcTRaW7mUTgvYWlm2m7ijniclov3XaziHsa3QatxDJPlhpthSQ2dZqYQlul0Apuz
N0/ydkEvKG7ovgiIU7VnBtAuMDTp00Jl9CL9T7Vgyz7kL4mNt9BrEumMZ623ZtPW
KiuIo/eJ1NSQOvtJHk1re9KDABxUd0V6vvxO7J2gj9T/pUzlQ3W1RjEAdEDFqUzt
OHFCkRrFSYiqDLrdAYr6xsJjQ6UJcT7QlhzXPIJlLa7WZXGMLweI4+4Ack3wA+SA
pYzrLLtHbBnI7fY4N7PfvGg0uJIAIBu3mSLbN7WeMw8/99VtDiLChWD2oylu2Lb2
5FjyNrOYD+YJD4P0BGNiQLEemY+u3+yVTNH9eKzPkLFvLc8jIxW7H71l+JeLZAJ2
XaIonUXpl00fcjWQbUEV6bJVW8C8G55waLLG7U5JVGnb1fPBJCtYVwT1CF2waKlY
XgnEdJa6XxWwxEq6hQi8wj72H93cY1PKvzoFANsVXYYzcbuyK+OP6ueKluvXXRci
gPrde+DCmmfgvX9VIvMYccBj7kBdfNL5FhTpKQnTtnYHIefLa7qwTDv/9w5wIwBV
3ZzYoWdTCMg90ZmfHBsLQmVr9AhrJy2xLI/rL46qBvnV32w6tn6JQ1baR4nxQJRe
tuus02o619Bo2RdXrEmsx2OSJMffcgixni78PQ3W0DzdaUuH1ykHO+qRqZKi+nkB
Z2r7Dcmyg6+zOq0MhR+X0XC4TkprEbtJ6vOh0zw/SmIpibxE4vowU0FPFzMFtTFr
b62LClmaAYfOiJjhUAWlS8KpsDbq9onKxs/dUmumn1i85iAGzDwpgM1nc2q1eQy9
4OjpZhm7DDtykLNmrbfRYb5nXW8MM+wr5bnhM9Xxri7VFkDzBa9Q8pHrKW3sMyAM
QsTNQmu6V/RgpEnRAp1elzxVWsOIpXWKChcNUQggpvl1jp6ID6J4dCMoQwDTxGlZ
jAEZIkpSmSqxFFaxqnRdDHvZso+j3v0yMT7436iAqCSWFedD25j8E7HGCIN/A673
My0ZFWIyhsLIaEXwQZqxrQLebQAvxHL21bOnQTx1ak1UhHDWSMjIDax/ooRLxgZf
ei8sR/GCz2DFW4J33tukFafJouqz9Os9XyUMetuVsMI0ArgA/TPwAd8fCScbrJf3
JEGCIODxQATE6Ww9p3Q8S3z7mKlKTY9gDj0x+arZDp3XDFTcFS8PN5wSUXBoI6rS
0byUYhptSp5xFz5Qe/ld7T44Cl1PvSL1Z9dgd6iM2YbZCJZw1qetdSi0ntcO4kxv
1f5GSHIqVFUKa/u19aaGwNmCCEyyeCkSNnfcTr64f4gLN5ygtMnZmh51k4rujt8I
EpDmHJJPT1KSkakUCXecbX2sQ1Bfht2UpmarZxRBMrPOIdKNjbSAWEmPXN4yQ4Rh
KNKtwX/TTl+9G6kmYgUQFc1ZtEX5QHxOGHrPrKKl73BicnMjD3rO/4psk7cv72j4
D5MK7VyqN1k+it0iuoQOKKtxHWJjUqxkjDG6LnMTwkIwgS63+xEGi8IbaS4YlU1O
+zrUvl1jbMA4rrZGekh4tr+JYjBlnrGdHOZ7kb5duMfmRj7+Sfy1euYmvCtvwLFX
efwcWBArvjX+zbQJZ0xwQNzjhQguE7a2/0lRJHOraBrQ2CfFRYycyXs1yXisbPPe
1F34Z64tZt3J9YnL8aep3TLEvtEXiGtncelTU79CRN02XV+hDVAJCAQPxyxeTDvL
nUO+ghPOwycKzO3L2dyr/3xnG3wiZ0EJimS07h9SEXmwMzPvIY+7pSf91dg5Lj/H
xRPG46GVTxBsiIYf19dhVC8G4a/KDzauo58xY8Bla5eeQ1Iw+YU0MAABiiKt9+xI
IDRybbdz6ITK3YBgnpiaIqcgDML+guiYfxr2V098dwMPt5o35PAqXcjB7fO3jMNL
UiHH/qdNbj8eOfXT36j94b9dZPq/xinLJ+pyt9agT0UK65Jr3AVAi5qFlNmNy0an
H/nXIJ2U0Ui4M6oVp24JgQPazlVDJpq+0yqJr5LtWPBF+4B8ohtUloXBlWX4EKEZ
rI5YKKnwAmi5JOxzg0cRyKrYCAEmR9Rhug92fzFtLbmFj+EWi+97vkBdYcaSMMx5
jwt3tP8vpGob36ygB/s4QWbQP+UGCENBbHJLC0lRVtR81tUPNS3MEosOJ5fcy8yA
MCU1GGzxGtQfnqpHFLJ0m1Ozb5BznKZ//T8IFA9TQnKXcDhNNTmhbWYvCI7Ak647
MhJDqxwI0WfIiAO+hcUHOV5bzb56hVEHFxuzJNv+canisbSHUuYba1VrNvPCwno2
kXFescVkgBV2JfX2wLI9UYS3gW17zKiZmJeQ5sr5CQ/3Gr1gY7XQIV93hEmub2ZH
kUA6C/qhVZHH04GJa0qUtSfO3CQFWUAhIyQJk5tnH1E8cWOGFacpInFx8Mg2QcD6
29A78uczgkdYwh5SRRfeGEVC+RDMEwJCYYKXpS6WQamGi2yBFddaooe+qBB8A6ze
Q0Bl0H71u6ZYm8/6URzzB438uaj78iI4T2bcFvOM5tHDm0CBax30RB8LPwBh6S65
TgqkkeW5UOQq+TZH4E/yNK33nUyDGOvUGVfdr0gl2V42BaKMNr1squzZ6bO4NOgU
NWJNnp4QsRDMRSreje5C5wq5jiEbjhEpwakXlw5wCKpzYZE3fakI2DdGqBmyRwzS
ZM3KEwhBj5cPJGhI9mEyW6zz9I9uwK8K7+w0Op0cMQGjzQkfruFWVsoSKT8zS5Xy
OpOtCHEjQ1Lp56Q6wAhIfZO3WPmLCMe8Vk8V9JBBgcEwkRnDm0Lc2qTkUb3bDqnx
6+x32HT577CgBIjpADeHzwTfETZKl9acNqDNDn6Ci4KdDZLw8LucsX6cea+W8rAi
xmPJwLJqmT+8lAqX815RMYgIr/rWm3x4+GoKgizvGTX/Pp2dbbAQwhQn4Q8FGo9e
J9We1pI+mwe/J/+vdc9RFdkb1vL2LIL32t85RgCK0ZpqzZRETcvoTDOaxM6ibUW5
NPTbsUskFWiXmCX3PZItRQmfa2/oY0jUH9d13hj1+7fdZuuKRbksAGJZ0OtKv+op
b2dpeXIHehsWr8ONfRqX1R6d+jbFZ0dAA2AtjnBCECl8IIspTbqlXWr684nSzK58
sC7KzimlCiwCyPATg1O/HAzTKxfRPjCZaBAxmfZ48qXJZuJZhG+8YZks9efESCss
FXh8vvgb5h3mhHti5on+Kp4sD848mHla0FaotQEZJ0gQX8/A6OARhdxOLd9PPFRW
8sioCiJAqgZprpw2Mxiz00iMeFzREhpHA+qd2AU/BZmnG6szuUP8Q6cNo4nBt/fp
cA6k8T+EMSf+PDWOvL064wsC/kNjJ36DVn6y+R/TZLwOXdkGZeP2Z+QzZgSCBIIe
G0c06wS1CL7sd3KOu9hazLJS8PvjpINADPMI6OtSU14kiv0g7OKAKbB9gYnlHV6x
EfOw4VGJPz8he/eEfO/+HMygL644D5FkDtRP47jZ9dSA9Gf+nUVoDC6LKAEQe/hy
Lx3cqUsiLsEXlXnm5A3NWTAVswSAZORV3eWd3MhtLSPn88PSS5++Kv+FIllH6wiY
4CoXmgkDo/bqhA814NX956aEPZBWr8lJT4jsZqjWGSIQqL/U8i1tHE0/TeCE7kVv
eWxAaj3i03esXbMhSz/NIYaNISfCXILvRYU4W5ffIoRs7liD2Ap2FUWBvg9bOv5v
Aq95LbJXSVgOXlH2wHaR8pSK6/TxOE+lIQmXXJxxg7DUMPbeFxJ2T9hDP3WzFfbg
LREent9ptlM7twrLqC+kAFOp3R8AEJ6o2HXNRVaCmE7raISP5cdifXsOg9U4wxXB
w1P8Toq/gpRVuty77GNw2Vlq0NdwnnyiC9wbPIeQsoGG9bKcxXiF7X4zs6P9mmR1
jCenYF8NPIB2GD5Sy7IhCEo8irR91e/s2u0h/3Kri150p1AdXSz8SCS9jK5BKFkI
BlrGQ7tlimKRCH9gZBbIzbt7Wgw8Z9GwcY9bZ+tB5Iwx3aVloWv0TUsbC5+zj92X
VPtpVKqhRgeHJy/4usSDjPXAxyiU4YWgLS/Vq7HFv92jMVOouGXIUrkBNN/jYV1E
FVsLJRRayQCpe2+CXhVV/09JLnNr5TWywwc7gz7gkTxaafrPQrEn8kkxZbj+B5M/
o0SnuTvaGILugNfJboC83LfA/JeTnv012Rpwtb1kMp+VqM8UlPflWCysfJrnNPEq
AnK/QZWexvgUSbAbIkNM6goN7G/+6EY4gbuyLJAs/lPG9SeJuXTKlBXcpFfSwAUB
55CZY0sX0e36ftAB+tIFvWhHPdlrRv0oASRDqyCeOz8EAtnVHIXs68uwUHV1Equg
e8AC2jF8J3xtjWNFPwZekYPDgqEBeqbHateVJawjpaGZQB0pI6dBCwITj9GwYoUk
1IbTyJd0o55kTYQKP0/98eB1qNplkRdrfNavYczSRl7bdZu2XMZxcy1PtU3B3S8s
xmTD+8LZcr9o/6DrtgiYkyOrisYdFQaddN0VTOLGWed3up3FqPgfz9Fsnbj3i29c
lwDbbOY2MwYx1Jnkzkv11r0bt0D7dk5YWwm/r/aMxnPuEIjs26JkKfrS/XD3TF7y
S2NQ52eZXm1lewCXZaf/uWO1LT/gzGPF24pPPv0/Jn5MRPX60fsQTB1tl8yvb/aV
OMEf+02T07Da5hleGfUQhnSE0ivckCRboRBEFGTeA9LZ2vGqXg7xOrWWjbKPpq4O
gcD41AseNioNtImO2edgPhnNS40dTIEWxtddgPpOtnDUV6R2EvnDmUBv5bdzirIH
b7ClA/9EZ9NrQ8zF/J6z0S4zcHS9ypP3rj6RwuYhOSCgXCTi+KP4tFqGg0AC5lPk
kXsQtG7Hmm5LF4hDzJv3Mb6guFlqRfUzs8Y6P2oFi+u6YRpOoi0segkjKU/0z7xa
TDqhS481YThmH4zDR4zO8BWQY6Hw1LE1TwlR2pqYPi9QjTNGWtceIM93h1m5+xQS
G46RWfwLJn2AJS1y+h+E1YECC1D+pKk1ytf0E2YU/ZIA52afKvVHWA4SML3wBD5+
tmp+3BTIC3lC6sKTkk5oJh2IpPjD/Kz/cWJjJZIOBxmDLjnZl4Xsxu8D9hf6aKC5
TY6d4mgB+y8rugk2s4ypr4HkAH9tEyvf43WGZOvxuGplrccUMv69B2qt0uToVcaV
GOGStibatF5bIuQhI3bp7ZmqWNc2KtopJy5soQgJuoZDKxMKkuDYaTi27+PhwOCl
WCkKdC2p9KrLHoeGflwbHBLiZoal2NJEid+uZlhyRAr+MVTPersWNZxCe8AsYtm2
UU0q14hqBF7F6mg/1GccpaQcqq76iQ5Po3NjO1CzTdQG504q92z+68BQgVJlkhFn
lFBEdyu78QUxB0bukc/IJyZirIKn25ODDJaXYgtu3YwXviUDBRjwK98MfLrvjXrL
GHIomNCBbc/v/aC3+aWzfGBjTsY7AwYqz3FaiFIDE6VeZmSkbUR+qqcHaVFeyejp
2UszFNO6l5jpU7iJDkabi7YYG/cQ5xyp3waK3ZjbYZocwMtAqZLmzvDHinnwPqxD
6+x/oF9eaJ3cv5O55LDfxyaIsu35pcV5Jgn2xg/1BakMYujwwFjyDYzMsPQdf68B
Q/XpAA1RE7mIykeRwEbcmbNM7sibpEVUoe3wdh0mgXg0/Uu+f468c55bI2ELWm72
v/xLCl+MeiZOx1zCoq9PQmBJDcU9/aBxaLFSeE6kqxFlDMygtVVTJVMhPi4SmOGx
LaguH7G5D7JaOGiRwh9y+/qvLhCSDqLXxAkfOqyW1GzgBVcMtQndxSD4lGD3wrMU
Ans8GYPTacwQkrpAxUtNR8yAoekIs0pGwd9EWRF/SDk5U9UH/lIH554r6K5nsGd8
qW7d3EnfPJWNTKG+Jmd/XqrqXpKlStfeacVk+2YvTzHFMHRyF7rtM0OMjprgggvt
whKkdaT4EtZW5c/fxOoJiVqhYMH6bT3TqA7PlY/QNXfejhfsNcyz8sbicexQT4N0
cBVyLQdlKTYNWk6Ok/3kjCKVqADZ+FFaTB4Kte/6TwlPOgsyc+KLU36eXbVOwHhR
Bixn4qswRB4/A/Ap8/kZbZ3sTg+UhcrJEisUAy4ZRfDI35xUMPGHDqYEG2F08OZd
ztytyxwWnTGKkCelb9ObZeqfqHVx9AVeU67v72pXaCdhdgAbXo8Q4058+GiNrSG9
ruVKP+CUbUqSyHG9dEiGdwW0tRP8f4+Aq4RUsaw4rbObsfu5we+b4n53dpZoRskm
i6hyhTkwQgpyWvEjXcBoB8dOgkjFUNkctq0fsLWc/6XIsJf6ZP4eAizTN4er49Dw
395hE6FQjAaYxppA2xfB5dN/ulMZZUh86Aex18aP0IK43j1uvImZJlhS9Z4F3eba
w9UzPxdhAmgNehet83EzcuGELyvhy2TBw92jXYmpIIDg+b5GwNBezyP4FjMfAPSw
BuQy4PwP6FHzavT2SLTjjhc8gISJxgarguDSmB1S+QD6a7PpOTrzX44uc/LvA8oz
fbJDQDweuJKjwVH0h9aE7WoXVdtBYfq4kmF3vHjgOEZ8Vv4rgXWU4VjjuMFgy3T9
szZd5HVGUuHWGrYmhSmJ9kkTeyvEQuwL3b7Z7FUnjJJEiyB1g2J5CErWpuFKZhqc
EJpmInNOehfeENYL7WrIdBUJ68TK0QmdRMlmACEwYeBu1pAaLW5yauFkNVN1T83w
xWKchThIAJ1xAJloXHO6X6cchCBUd/XdkxzI7RrxOw/3kZqy3MGfd/eu6eBKk7or
JYof0lpiujVapcQLhgL/d+jKDGd7xlNF5/zoSG0QyQWqk8rOWif6T3OP7eeLXjIi
/DMJ/JsCr9pFJFpTULFXoagT8F1/V1an0gr6yDQiXwP3w9paPqYMq2My0HPoCv4t
KUh4YGsbhehUaDyJWfBMeGGg06UeJZdHzG8pP4YIjJlnWq0mPX30j9iLUITebPaS
8/Wm5ySvmWw7QfulJtg0ezZo4BiNtMawRksI2e4CDN4/wYU0Op1jq4d1pdxFOhHO
NMvP70SqAE1xEqSOjI9e/RhLBrj5hwd+5OOAcjX9eWZZePBJKcFtQzw+j6MmgkJH
P/kyVEE0u73BtAf0T5gBRRFayMPMXqs6PsU6IwckQaygEoe16/8IDfKFCxbf5P86
hPpRvyZlEFqSA2gd+7Lwipxsy3vq1s2frrPEX8HWNH77rBPVhbrwGejMY5Renz6X
taz9XXmK+Z84GHCx1T5KScm4y0d1SbtvnTj5nVXTFMb/a/jtBUfu6qGLRW9SWk0x
OBoEtfPT48l3nhklU3BQpXNuRTxTXtZYPEew/+FsQCzyYiQ0QwbsOl887NiG6RBV
gGfClNDJOS3XBpwWeD+EhCk1w1ibjZDS3IWxcRo9mrpjokDiaeE8FvHcR2FYxAgO
vRFGBb3iMAomuvwDujg/29fEA800XS1/PeeQ11TLagMJP1l92sl8Dt9WHrpepGrW
ncHwJbkTXRMn9bxvLYiOLbu+eV2eoEmHkpoRqOJNqil2i2VKVOF9mA8TX0h3Tfm2
NV7Ao9c8m3SLuqVQsXCBrBg7Pn4TytBnKoCD2+7dmH+JnSggPa+5tvq3GkHlnH7y
yb4EHYNtoB1r4afpM3BOl+vkKxBGCSV77tvoToKL8R003V5nqcT8p+tlcZMwBFhx
mf0S79sMLIU0UVWvra0IEpLM+EM7l823w9WIRd3lg62dknSbBSC46XLbm7Eg4nEN
p//eKlC2MP6yhtIdoAzS2N4/69bJtCsMipcAGxEm/9QRcdN5QqLJvUvQAqVVQ6mq
04/lkFQpaZDzd8L9IChMFebg22GeiAhNEGcSzH/AdBXkfjPZdKq2/dFKm95pD9MM
PitztkdX/mjdDBZBNShCaSloHcySTgu5i0fiNuaa9V/NoeQIinyEc2xZre6AvOeF
G67aoxMMaZ0Y9uVpLItvvbI2ClY07jC+MyTI8ikyDzmd7X+bYqNoFvXhOMichB0d
zDcgw5Z6cT50qwcYaSraRlBMBUrayldGO5Y+xxV4e22oH/q8OCqXORZii/AIM7Ta
pPqY4I53HKP/7KcsPap7PB2cYP/v69M60iyvxzcbg4aHdBMlbadPWWG/uiQTtT23
Hh6z3RKBwE3se6UFP2vvfMoxeZgrojeyBs+dMzYZ89idH01d39XnMiUsf28y+lXd
ThBSIIPn4Zs5A1i8/ZX5/CO6YjGNELSNQMpZYEPmEZon9X8fCjHhtsS0PWnK2Pqp
HH80RrWO8t412YYSqy4g9EPCqHtgcjujiq+maiiVf0sP3+HNXtGjinjEK0gvXTCe
DI8snNou2noE2HhvcCBpnn7uAKC+Af6e85RCQ0nVr5GKb8KwFJCz/FuDpYKhjtgF
S+CiNQB5VxQ/359reN84Q3ApZUaipq6se9rwDkMQVdMTqMtkhGflvqN7K3/kISa7
zykCvkwjypa6Tmex1ZnMuiOZNNPoh1GkqTfNEm9Gr97cGLdUy5EeUjXXjyJkR/QN
bLC6VmkStVRSseB8x9vwwGDqitM4JLHY8cFL9pEjDRrHlGqQf5yUUrcQ+FKhd+kT
X6Bvr7NZQFiO5Blo/YBnHXYCAJT9TdeN7ATvvTUaQ57EzmEXkUpCupy8l4anIqz2
vWtEDaX59xlBCZ6K1WuPikc86Vfa+nh6V6PUdS7gBdvPgz7NsTmdvAhg7wL8UpVw
L8gZrZuUE6kXzFwvU4NtIuX3wLqVBBIr1U/7lz7iRStjm7TlI7PPPvPq5VpXrYSQ
uo0GhRNHifvrMsbrsfTf2/ZWJwWfx95qtpjLK4mRHeRTB0k39779MLQKKpahvaTj
5fJMb1kM1W95nIooI8G4l1hsvO0I24zrN1Lh2urELJrzQKjQHbVfZ045cFMMLt9a
d+2cNBt079rojZVedntUv9by0BRMvM/gZ3RkJg88FfW81p4oWZH5krBp4KMOCibs
rh9B3VkvexCT+zkOayMIn+1SAgoikHm3su7G50zFzfkuuUBVI2av0/IE1kUSuIbt
6SeFH+u6R9smc6wdy4CvFKlXiWtDdadI5Ah0yJ/jAwlMMytMt08QBhi45y+f3sCr
8Getmgs6ArPSDTePZQvgZ4jGXZTyFLZj9SGHM8tUEv8ADfjNqzyZHTwWKQ5JiWdo
SAT1JLZtbqj5DEWhVYy6/+Lmxg1f3VdFGXWm6rHKEdFLRNA7+bFSjtbYSTID72jJ
pxWqZ0Ds4XJZwuAGe+hAkTRQYsSS8Q6nL84P469jXOlS29Cz2apkci1ljGc79yWn
AmFgnUe/MOlED0x8HkWo3ILmK46iTNMcCExXaKXt0+5NKF/o3X9gyqdtPlVkJzo6
a/OJYlfAYJkLLsxvpVc5fsnwxdG6xE4bcKIQX0bbUOwQAOjplRVEsHmYK+cUtJyC
3Va32Zff6h/5pxTdS13Zo5cZo6AKkxv1+x+7rGmxz131y6Ow27QZ/Gd4Z4Ic0+YV
nktPXA0j2b6EkJ/CbBFXVkPTQSLgsr1HvgVU8cr+REfqmYVTUXqM+pRalqXDkY8e
5fXaDveX0gFGyVojP4qZCsII+Ehl5OW0fcWrRc64WA6oesb71WhICSEaMyfx+0vF
IswrCRI3WkQk/tqjD+O+zE7xDOp+5HFyuFhQb2Q4/3bfuPDFMBGlUtDt5B20CfYW
yFh8KkK6TU4HV8M0zXGVQUioQtCCQ+dnqsFkwGHzp8Ryq1u8I4Rpd42yiZv9IrfT
EiKrLgMtXd/fn9CnsfdbBjeeG5Uu6PtHkK8+DZjs5M9xYRtkZcCyLzmyUCfBpuhc
mQ/+YwPx4QW945oYXxexZxUjukDFdSPXjfkqi0P6Z0fTmTp5Q0PkzsJTsJX+i+yT
v5VC45wKLmLKZo14yApnG3UHb0Lj38JQhTeq9BIcwdwLZ/o8L06kO8sjqYC2HPph
onlflmV4PU/lPvjH/2uGcStoeYDSb5NpfdFMQrrYPkf12w0HFtoMzpFjBlVIoMrH
SSHwH3kVfbn1VZchpVP6Z2GLxhzdSFAwBmo+5qkf/lf1MDr3fsyw9ln1Un6fvqzB
MWzhWtTCk6I2PWlZwNpGbiQDo550EYSZ4aNoo+/t+gZhZUx7yHj5xqGS8sWy9n8p
62y+fIE2nET/jXP/n/zn6mV+hUgje9GtA6RE7EHnEMyep53Oz60vXN+JlqAKfWeH
m2wm394IT9YYOO2RYXDAveoLnwVhg9rPR+LxCf36VH0jtBG0s9ieUkKLlmsNfrhS
BSga2Ik/FK/Vqkesqd3pWyp1W2MdZ8EPScyjkX5w14JM0yojMqWzh1nwa4oGM0g2
0ACU6/3Xma3HC0n9Aqqn85weEVbvNYpA1xASyOeGsbDewc5Wgkg3JpzVyVeA/2sH
qK2SPyAJE0O+DI1aeZ5pmOpW3zOtzBv0Su3IfWH0EdPH1MH7LEact6s4fmdwE2qq
Zw6vlIilqQ7FMCsGgq+kMHZQsBecUmr5oFqDTD2ga7KfV0uyvc1XzWtGIEQXa6Ca
Ri7dL+1nxkNgog7ANOkvTxLZJuQV7B5c+ioRjzITVPboeS+2ckoJg37aAMqmoQtr
ucgYm+mGYitlZQajTCEtjTCECIUvhP1uXunXkcpYo3f+qoQ8BWrXXqFYFKT0JJHJ
lhNvFsQuJMK5ln+kDUbEQqo0LYM6j+p2R1Zkc4Xq9ujoxMcHDqmqpBNVUkDcS5V4
2aGOqelKwkcQC6RK0LLYq2XLkSLXJ1/EYzpnMTDCj4OZ2QUODAnZfguG9Y3+bO17
3ii2ZMmqRAev/SIbB6+AfoaDYRXkDksot98P4ODOBmHFvQohf40WgOOaaRoSVLWP
dURvmp+zX+3aEmB6Trk4G32pnvbqhJMQnDionxQ1satm6kIaLTpsysz9s/DlCRfE
DZ5sYGAx4zj0Qa3wnq1rUF2M/Lnop7dxnJuBCPFNPSPx0mmXVlc+d//HRBiXqihR
pxwQlmkTLFClrjnwqn8BkgfH5qMe9qM+zRtEkYOLI8iMs1zqmQOxYwMgxT+1BIRl
QXD3gMDgeECjy97z1a1gzAvmWhFFCNSp037YE+GpP0YfbJCtQHJhoSo9corDEbZ6
CErCZ39JYNWXV/I+tX+drSopQtYzjE4EWrjiXXKYTXMYMMRXGLvGGZqNGPn0oYTO
M2rEn2jzmGqt84UT48wN2jZx+s//Ln+szoVRUOTZnWIp1T3F7NGFHmIm9pQvR4Sx
sXCGRegvY1w0uQVda1mB3ruTjaDnKJlh6RSnJUPAFBC6NmeGGWAFWQxAblEexEDz
dZtimTbmVHt7WMChHrP0aERrjy3rIug2ATJl6XcYs1syHTIZw5SJeAiueGSFFIOw
rbvIHDwOWq+9TTQ63LYbtd4Cg4ReKP1HuF2Z428y3z9ZXgqxnTpUVe7c/tKFqflJ
JwE9n8wBUFHcWPIu2t6MN6go3hLKRKhcFxz9lOs/cG3efWk0NaB/HeAnrgxnt04L
46SjNz8COW5jCOyJUm6porjmxs/0N0WVdIkCDx/00f6UxhSh0LwCqQwU4T4iNw3i
oeu84dtiP26oquF7VMaCfJqfT4o7tx+7ezVQfDe3yCsYIKhSZWT+ftJslbPslY5z
NsGab3wFz/s1+hQztAWzIU4UmztCuziMZqWNsJEKzXAK8xf9Ozq2HK8jrJpic4n6
0c1mgek+2flnGBnzXELBN4otMXcO42qDlwLDWJ5PmQN1wo1muU+j0xLSiebP3k5L
1dc09AwnHgrk0W7re5i9gg3iZxMm5W12ijf4pAWFDHNsRQvM5mro+HDF7gwt6epK
IRFDJjPHJVUP5ekFrz1djJmw9k/UbcZP6+hWgFrbpfi2J2zU1Dvx6vXtcsb24nB4
tw7EjREPjDIKZKieVJkmNDAGehN6KsFEmbi0kD1ifkFNqY8jxOPQn1Wu7jukFxX2
J9NeQNDKDWFphD3yEQmlSvhqmbNIYgZQ9LfCIj7WUV98luUDueWZbLm1Na1jUbeQ
Nu4mz82B/9kQt7Zh/Nc5cexPIevva5vH21N5jP+RvxrBYv3dzbGvRpStmsc8VBk/
1n/F0uW2YjkdApGL5mGjp0M2U9dbeAemrTmKJpEkdm5TqfPLSmHIdbM4KFodNCPM
ZszSfzbD9Igoz4A/Sfdu/+pWeIe1G9JefHt/4t1cTwEo2XXuCmxZpsMWiago401P
AlWhD+DOWrhdGR0Tyk+IA97VUWsehCA1E6KE6Q6BGmh1Rimqap7GJVNtEOK9Oe6x
gQDC7hlWEV/NgJA2hu9PX6zfBkNexQp0A95NdRw3PHi/XNTlDy6oYSguH4gogeNY
575TfrtI48lugOOhO1HJ+jKxlNhP2cxJCjvvVhaN0i7GaQxKuYJJqBY30d97jtr1
IQwMPgvtSnG3GKFQydbTedeJwLkJbyXjn9xwseRlQmEHkTB5KtBSrPFbo6lBQc2F
UR3EfxQjxKtYZQXL69XaSKdPilyERCIzd7K5exOQ75KsGgQAM976jBb725LCMDzX
/dpmbiFiwgFwY/65sJhsUnzMUMJJbXQ9HjglAcByjAoAG7/WUWZCd1HDPGeYJtFq
Z1QuV2h35CWBkOWFEor5ncNpJU1GYY0RBlGBsagD1Fu5sT11DCvmdEyN64hoUspv
45Ex7DUwn/2Zt+YquV8T/gC53vsYnTca9kk/B9++tYdcaYSWUX9CPsDobWWEQBs8
Zjo8mb331NBSEnQGfiL+7lTGw/KSYKstMT5iMpoY9ZRNdyqWA8cMVy09i2444WXz
ewiXf30Nt+PZnWSFZyHWONuCa69UAprSQB3s/HBnI0metJwaeLk/zKnxe/i5/573
yLaE6D6HUO8lI/jBCVS0960IlmcAxslFXDsYwlzjXNBDp6DhlIGjPtxkCSpUQuOh
i+DgZISa/P65RPn7G9hALt/rQTqR6CUFlVmg7LCFODcqAjTohcvPYvKpJtOoCqvb
DX1hMpyjFYsJDrV/A/Ulw1Z6aQulmsXBd92ZZQuctRb3k7hAdKqpzV9pL8+xu3Re
k69/DSjKaq0I+ZYUTREhH3wMsNFrqtN9go0uESL3Ux4ChVip4ZgLf4nZ8RpD/UBJ
2jO0hKx5nEwF8WyZ5S7z2I7ZwLFnNtSvT7iuguE9N2zmNmwN1bqyU+YhNV38c4M2
wMT5dytRCFJgbImJ1pUROs44JHafJvyT/dpWKhbK4UNch07Wtq1YVSpbBQPcwtcY
NU5ZEFn8LGHgCIuQ6EjN786CNBpL3wr9W+mf06tF2DrPSgvCsQHdVpIGZJfSGKMn
TfOrkWGb1p4OBKfgVUsQsy8dAGPReoucc4LVYfx1s+A2nQfDK39EZCp/ujhk5c/e
0mZLhFtRK1GhqqLnRtxoT5ax5GCsHvlv2LH8pe/PhEUWupQHVSAeJzx8v5UTDNKD
gBVoCgTweQHIUytl6QMDZB/1kwAaymbxvtJzPuGyCmTDxYR0rnaE982sWIimCLsC
JKEKVTIl+N/9+TxJDr0BVCmfuIgTimT4CZIY0DzLqux40IHbBRCuUAcAsR0vGugw
O/9tCasdk/fMEs3FSpt/D2vqW7fuoDi8Ye4Y+IFcDdeUj0XsupB+2VoZoIf3q1Xu
pJQVuJA/kQqHpQlL7Hd05j3QMgqLE6V7ws+gJyVANbMWMfvYY+1gyDdknZRei+5R
Y77wQQxEnzkaH1j8mmIvfHXTlivJbIXzkzsMepPDijPR3Yl/TMM8plSZ/Xg3nkGF
xbgfKB3Tp862eqFD/mn4nQpme8D0Qi9Uhtn/CSpCuuJyAie8frZGmJByoM8quSvp
Cx0NzW0YXfsddX+nyvZqa9Vq4owQitx5rULTSym4bgPSf3IbseCZSSo6muFENbFy
168daRfug6Fzy6NzNEtqOnzx2qIj27OdCDr9niory6WoNKJAQrLO0fmjqbZVR7zg
EeNo57X04i36KzcPRm7ftxAiarDTOerWaDWCTxVYXQN78Pxa2yQBHFa9scyDFWpj
rCbLr5k4IX/8CCwTL2g0kJSmFAbNaeHJ5h9pxFxrmBEL+i2iAB2WUd33hPG+Gdkm
E4/A7ivsZBibVns/aeTb8vzlJJbBJ8br2ClQXWqfBqE0bIG+0utf7dWbaDaweDr+
8HgGi5NqxG+JSoz855U4rcg+picRazjbgqwBM1ZY6sOzABwOA2jhkKMp8u7IYSdO
CQ/HujC0qo92ytUbxVflQ7BQLKsLh9Dxw95Ms9ZhlMSHZF3L9EncHRyMH2kktIBJ
pqDhWUE3CJV8xWYWcIUI9fducvrtNncY275wCLIOBcq5BABNSK2dqDEQ2ajFlSCj
66XRp3AC3fhK6ugYKHcsDe7+gZ3c7J9/hA+KMWk1WUi5QmToGaz485PxsexuFD/l
2mRn6ocbH3m7FNMhp0kgq6JXnFsFtIi5qupa2ywVKvECEK75RJHklOdzRVhgEMKf
bsZL5JK5kQqnGC+cQRmG8BOj4KLBwgeASuwkCJ8Uf3Y2lt0pyHO0DY7AbuOqtHem
bqmnFR9eJJSKSX/hjnZkNJv6kRnGBgB0WSms3gJcP7lj63zXwOR01Ncy+H46/jru
g6okJLbXCKjB7vjvlJ4FWCbenieXHcocqcTa4P9/QgPCuMBe/Tuw36IT6yEfTXzD
hx5hbueZiNQg3LnZBIN79mFdQ9M8zGLYBBsUrTdH9u1bBgXlhjbBcUClqaAoJhjw
AOWxgy/OD3JFLCrXWCSh1gUg9svHSmHxZA+VW+/cCTAqQ9GwzvlouOBRoKCFzVc1
bS7SkUsCEzk8wF/Ui72ZLUFsroqUqAb7Wf0fVnd2Bfqn6YAoR3hzvt/oAwNoU3pX
uJs6ew/8BW52rfe2Jd/zJANRwOVYIVdtvoYZ8FdDeDNNy1SidKlUUvwrdOtdWv4d
lF2AXV3vY++GzX0AgEUTK3qowGpHoW539YqCa9aJKQRRt1MiuUDL8bDYDvnPVCiy
8JvPmdnNN/9zb6+OgnvefrDIeaW5ER+pYTdfS2sgvTrU5pv1tS/CzsWYlyXHK7TR
X1Z+yVjaYif1nOEn8M3faj8KSU78HJeb2YRwkOYjveaoCLdYheUPxyICAf3w4LkA
zwyPg4IKl8eZUULYMtwGEScevwDbqM/kXSFFMMOXxqtY9d8B6A5QKhmIOxT7QY6X
fB2+QAvqfYsJ3ffQow1VSv2tP87usJ2SqqHhMlLv78T6TUc987XkyPstpqcj6BNn
xRvNP888lA9ui4nCwnAevXFiEuPjIVGH9IgkuuW1ow4+1E3aVR+tGFeDonP6lw7i
/lTFSeOlu2xDmYuggkTXkQd8uC/0RpKc4ekO0moZEnwWMSS7b97wuTSqqP4CBTI4
Xi3ziMkLOOOBTiqjWGvxeBeLIzyuGB1Ap0sR+ojbIzZie99ClMxKRt1u3KtO5OYL
1A9t8h58Rp7DLrdQN+CibCjU6W9II9/HHWmqAt4JBgMLN+y3is/Tz2K93tuP1qDf
MUef4++rjBnOb950L0Bzzs6M6UZC6XM/HlCMG4PGNCEQsJUgJV6DA1W2M+7zK6JJ
30a92SHLH6TNKVNg4kmpU9SlGUK5fUro99jxskweC/KPjYqAjh5C8ak7sHxbz2kf
foXA1yrKvPsQiKqb/ny3Z/yPf7t7eaLi/hjhFOeaXbw3kkuIO8baak+zeiFzof+6
fQXecfETx9aD7vmKHKTzNwJm88lhRn4d0jtXeBfEtZTxYjyKdIvBDIdjIYV1Pgja
R21fttikp25v1XoVXrCYB8HYl/BLyPVbfYs/13xhkX0p9fRtwkW+Tjm3DH4V//VL
Jq+Xfhcw6HexbjIhGMv9VRscWfCz7TZbJjT0+9vnmljJrSUhiVwWJT6y3Icf0GkS
M9MtfyNOKJimWT0uIvVuK5s7Ja9is1fkBkMIXalT4fwTM+3T6pPfItvuF69y2xKp
7TAta8S/3EKKbym7uVnHaUDFaRSyp+fZ0go0W7ciDoBwvUWjGcERh36/17UMmgYD
XPEbmmdIQo9FurmlVJvowNAFfr3lCaZCiHtW327roqgBQznfBn2R+CQjVhYk3Xjj
le4YnE19h9z7ek/U8JxnY8ka6lfalnCrim0D8lhGvlqFl/oJKV9Yfx8QKnh+57sn
nIeH3vF8MMjf2d6g1TKLrq3QrRlM8qstUnipyYCwm1uKQQUox8U+xPaS41uPyZ5p
bQatSOiqX00dduW0q+AN86F6jomswHYJS4k7njKuDgW8ECKQuRMOv0dsZaz/8AEK
7UYfTl6eH/os1xrwxM5ZndDEGLgBBkroaUZ6LRcltcbNbL2YOS+TyfcLMUvF32M9
JX0JB9XrXJ1XGsmXk1sa88t4aHaBR/yX5hhPgdsHNvfb3eSjESqKHhIKSd3vyUwc
BZhEIm0Ckr4ZgIO4jYcnIpI5LCKVSVxeWVxZH/C0AvhE6Y8IA4I6Us4vSTX8EqaO
r7jvyhYh9Dk4BUhh85tdcVpwTNE0oHY5Cy+uHLh1ljA+uoaddg73QOHK+u5xMjJZ
v2tSYgS1hB2Coka1Ui7fH3K2jSDPlSDnSlOBuwYA1GS72QfrXiTnlH/j9FbSe0ju
anAafnMamn9B3eBTZgRdxsvDuvfD19OSZWvHubkGj4wjTK2+R1PdCvCwvKgEZdUH
xx4GiZt5DuoF7MUMtgAeb1xai6qG1y4yew1D0ClBOEctlbBIMrxwdKaHAocPE0rC
DBtZubRBT5WVyvLZIvDYg9uX8xtVkOB/fQNfVYUD2jBhZ2r55awn49tteAQZsrjV
+2bMfrQ5EDD85zcft0uT7dg0KaZ05h4P1oyDR+aX3HHg5I3uBrJz5UDa+bViLON9
hbuYX0UOacaCP5BEeEXMnTuF9olG6I5zgJXAU98jBFcd1yPG5orqhVyQmngwxiyU
NZmfFICos6ZM6DMP0GgnwCgoDE8JkjeUbwovvW6VJcjaMkOHxAveIDPS9ECzzN2S
C+wSzNbnqRBIgEMPyXxfyW06RRXOjdlxJr+imViH8GMnlcuh4BW0Qsa5nHeKXsqD
hUYwTmPLdE3xvagIBE1RXl13iWlNDjPOi9L77uTdiretIgqVdw1ox379C9hRjbFW
KSgGJSjNnvEmMJLEU6XB0KHDlt61QFcmWg3Z7iv5wK/fbScBq/Zr8Wa28QJOVtjV
DriWnfL+j19vDPVwl8AyYutjMQp3Pw+fcgIDYa4gVssmvLOaYS9i/YDMTwxlj278
G6U3jks4lzPpbzY8QJFQULRhKj0d7pCdhcI94GMfJ24kfb/7hYIpIX4CYeu8nayU
tRnggrVZpEEeWmYSi9VEmdWpwUvA0WPOOmw+SQTTDn8mlTDlN5+XYDZ9GNZbYcmo
G2QRt0ND+Dsev3ozOHuwzDtbAKp9sLY6t1zQvV/fxS36ixcHB1kCRhcQpTYRPuos
SLQczpmnylOFR6cehxvSVBx+Qo1DxTKWo+iRXe6j3RdG7GJ+lYvvuiD3jDjhrjvU
Sf6yuYHp1yItDSS86Re6dLzI2hSCtLh6buiRF1T8S7WpeGqwjGga3flPzsHm7vEt
1ofNNwDzvdS1YmVEr2PLQcwSdagGJ6K5925niG7GQgsdc04FHRQPQSWml0J1B0Ms
K65z2PCXJ9CftuG9V5BWGWNUWC0/uoAKvlurU1ogW8N8oQH4jAmPid5XezZMUWoh
X6Nm+bRSZOanRwDE2yHTOkBOMwku1tRaWQv0NtVaxedx3SNUP9at8RRbHBhE/XaF
yH9lIrNJJDAX164EE8F2hxpFdRZLZIMpefZZ2e50KFq/2QIuNFc80FuPfI4h2mRu
UMDodL+M1nfwk68+O0Sl2g3gkyiUjxkWpvFhYoksW4fDGUU+eWxSeQDkYGDYeYxK
2F95DeMrCFL5hzpI759Fu10dHN643BGGsn85H5apRkBZL3LLTxAjWqSHVh7OZ2i8
Zj7Ulyt1AzZ3cedxI6zHXftBs7DvWoDLugVdQBc8F+MsvG/h9AAmh4xyu7NuACRs
oflu7HK1lIY3zXCOOnEkl6z/sdP1PMazwauvnIdnvarXsj64GQkO4ooLmvFVlBAK
tUefEIrCcQurc1Gn7gcQa023kVu4EAX3tq5+GB1OJ8+u8rv26XD609FoQSnDMWkZ
A8ZE7VGCUX1kq48pm61xIs97DZgtzibuplGCPk1jSj7zNz+0SEf26+ewZYU0C+bj
KsqatI6l53B+PAWZ+3tzWCPt7BhI9v5ZUIQYHKlMyCC3E8gzRbEuUHm2dKxV9sNY
5SxlYdxnH6nyFXljYCuwB2wT8g6c0h2rXgCa+cJaTlrX3jSSuXPZ46jr8NYpRn6u
SgsCsIM++ln0II5jDQ+JRc9OL3Y5WAvtzZnr6DEOWanaXxu8MQAosMm/3qOxbO5P
Sr9ELirNmJuTi8sCsvkv3V97uqe5YEFgIPd+OzK8ABY3QpZztBmanERO4KNowMW1
eb5udnrWB5BBYofInsb/2YuZkurBMMWZFMGF0Z4L2sGrC2m5gx5JbZuKQaHs0B5E
VEGVHPfkWwSxriRShVI4riGbVH0BVUDYmemUDdBTd/gfhXq4ylIcnXI7QmXW3Ay/
b1IwQwzdwfx8WodLlukmiEZbRF+vXZ9cBy1w4A846mJB+C+QJrPX4bFeiwDzTtw1
j/RKNbaZS0rwaFIUGSbNmPqYr2/2Axm/tPE7I5r42u8q6xMSfTofFuE7HH+ChzVp
8w+Shez/lM2BDe1y76U+DLirbGZ/+xQbypvrNSO5ZfceKASwvl1/t8/CBFanQjPb
PvVss+1/uWx2hS180Wfctsvl2otLBGl82RS9bQ2RVB8u+3ly/kC2DBXa9PtPb9Zk
LFzETtXoxhV4DVwwQcIkh+LYi7wVtp4VBdyvHeUSDSiPpg0BL7U53Okx4IZrzdrQ
d4TQeySuyysd09MB6NyEDIUd1lW/JXraRvRjxz+Zz32EI4UTDzh9Cd6Ye1+qbBUK
qWDf3y2DAwgmC7vFpQ2S+4sjbu/s7bnryah1lA/86b8j0Hau29UXhnH0FeADydmZ
9XesGQQkiPz51g8zC2oYScQTmQq/WE0Fn6FD6WFTN1jRewruZNDH0Inepxspi6pV
SFwKjO48VjLS07yDSm+K+CMkcjxymnd/74L98k3eRxpg93ZmchShl4/VTNCgb/5g
abj52wHr4q/A+xKMOmjM2rIMuLAL7fOBbhLf5RbbFHKgqYwn/aQQa7oG+DrYR4n/
+6jSF9eSzRcpgMmFkIYRH4CIb1g99OWNsWn7pVXsRYEo7k6YYoET7cC2L7Vg8Nl5
0l7SSHzVmEXoo9+pI8MGCesU4N9tDZLw6xkkKVDEShkGcFwZRg5WINHYEQ/ssbJK
S3dEECACdK0J8rSp0C9xYDjSQ3HwWYDKritC+rS6FBmASZZkpIWTDlV5ohK/VMdb
SIwDaN/xCe6kEps/Jexb6E8FBBllKrHQ7wJ8J8iCGPjkzMCVwUqrOkZvyLJpsD81
RwGLj1kkG0xVjSIAtS/eiBiKJ59ol92++LmEGMuTzqzQ0M3kDLtcVguuLj0rEd1f
JySuZAKUc8KpnKrfcuBrIhECOljfFILMxnN+bP7tGAx2LN3wSe3jfV5Ugn20yEaQ
To3BZLUKrywAxCO/H/Vffn4JplXWxHYAuNt6o1w+yJP6b+dvjUkdFjcUpjfIAClP
eZU/NACho9P/4Z2b140Vx8kT3LI6ipLnroEiTG1EBlSXudq5bJzuD1SCtyg+3W1f
4EGcL+XIpeIR3hd89Z93Bpm7VT8XVz0DuyPvaOEin7nv8oNvD50u5+XMP/V+qH/V
CQwchTQcS+LcUEudU/iAFexOCeqXjbh3Hurp+NdK3pfKwDSE6mOrhwE6Wg/wcaRS
Zee8EAvZ7I2ALYnbvOQRPhEpanrJ9COaXvXf7qkhNfJpcnGH5rAB0otGJ8FCN9S0
jv1F0VzMaDziQFjUzCSEh87D93snlKFbZIiNjcUxKmmlSKP7gThr7ESkESC48pii
/nflAVNmdsKMIOGIAd0e4du9v/48HMQy0/H2Avnslak00UHIeoqBUzoRxShWtCVm
GO8Ti3ijg/5YsAwj8MRe1RhRDI9O3Yl9DrnwOfJv3gjhOVDJMlpGidrWLOsdMEiM
gOD+vaKysICMukmcfRSxBLefJWsXZEaZ4GW4gvep8adM9z6OeRRaWgTytrFuW9Nh
mJso/hsZagibcEqyXCnlwthFp0hR5rBs5i12HSAO6gY0sXaeHfqOAONGyr+evuMr
UQEHP+frgiXUmTmZ6kI1MzZ5xmgkYPObw6UDzG5slgzxFNosH/udJHjt3gThflwO
METhd3Wgd/MiLEBDT++2ate1a5X89S2J0jtA66to4lxwPvW7H3teuzO36oRoI1j+
GleDqkzpR2CnZjLCr+rTI3Es7XR1qVimMczG1deDv0IwYIlFzn0e3a4m52zsuwEh
rpgc9LA5U480aFlY6DUCxTbDkdsNWwgp5QPF0ITB32uBBzaUMyjD7FA9mrKJoTmM
0Ql652XeWYpb6YRSQBiWavq2OJcX0xQo248/SsuJalcgdIm4EAQRN8Uw+LhayX4+
GZhKm/f9fT0PdoeYLP7ZUaYGjqsC77a2cDv25oDckbdtC3G3jmL7rIADJZazy5li
ZAJjZVZL3igy2boss8Ol+1Kp42VhRl0ppdM+CfiRxCIcT6yo9lj191eCEgUFPH2p
OAdtjG+rY55fH+2N7FE6mA3ns/NwH0r5+ZOixmuOXvda7/lfmI1kiEKekMtQHIOu
hpmMwIhfcsGU5JJCahhZlxk0befIen4HihfXR7VxSpB6oe3BVoYyx0a72ss/Di8L
ENZ2GO6FtJRVY5tyC76UvErEqYVUm0m4gtQH6qYE2TafYmgoUHFsBF/pVvP2rakw
2TDfRNnE/JCH+BQB/hrP3l7jp21Jzh1gqX6/E1ShgcgwB36PBaUS50zuogAwg8SH
jPo63si9Y2Aw/rvTX2lrnJ+QZtp0tbf2ben4HwfSISGU17Qy1uekCsEXjkpE8h9R
mjWAOOo4aAWZG1C9qTD8dePvXmDrB8Ht+ZwxDhHfxBGdZHYacq9liHStv79+eF/t
s1yQJmFw/fBNu2zN2FfqQNkjSknV5zxJ7/4Jy0MmfACBSwX3pVVOrPKKruCqtW7V
7R1u4huL/Qh+9gtKPfuBp0UumdMhSeebKafss/KNQWROwN2UejsP1SQAGtmOet7R
Ji2xO04E113yeS07UH9HaA7HzuhUe7XaaqNntNfcQIFEkC5auJ8fdS04VHuh0xFq
hR+Eo+fpj2j26wIlbh0e0FjlkJD9cNoWvwVwMLvBo3kRrPwKDvykQV83/XkA7k+i
p8/WbOcW/6TFEw7qn6xABbtRvkv6aYzdHATvY2fUwgz5p1R5pmEEqPiGDck0duau
JomVokAy05UQ+FLBCD1tODUVlmD3VQYMZEqr3JmmrH/+W8dcYXBJwaF80aJ9uQ+/
lIVpDOAOdQouiVqvHct4213icf488ZlTGuP43TLxmgdvOLAO7thujt7bGUVj16/A
SlEOM8Ma8BCNncPjQMp7sei7975euDUIzpv1kTFJEhQ8mOfMMQYqKUrVq5kq8dzg
G0eT6bCcNkEjUW9pmOdlwunQBoOjcgYbNCuteZObAFDFKiLjMr8Ag6qTS5oX59dS
gyMRTNbMt8H1kZ5h4CTTQejvBkGG/PgZUBkA7Bh5/siLee0VMbd3/DwCzn6u9P9l
edP1UY5rxqhARwoXLl5K9k45fT6mgG8iTpBM5grcCiSKHJtI8mNpm8Gme7FWMV2v
apYef1rSm+D8bjK8WyZzDvQ3m8tZ4Wfss7CAR33Rs+lLQUpvwAs6HIqyI8XGPZM9
tu84qz/S1Ek3rlk8PsYb+uqZO+EZJnXBFzcPgGWVCuhGGf6I+8MruhH/PHdroOth
2IvHUt/9CCJ5g7UHVc2ECyjhh8QR+Rhbojih8CM9mK9ju0h3Ggn/8aa2Df1NRZDD
Jmte+ZRUi5O51E+9t0H4bNXZbntiyrHvVGECv+CYTzNtXgp1SyEHyJpkV2Z8M9lh
ow4kJQJHHWRMwG6zhes4BYx1VMm4NcLriSxE/A8yuhppVDTf0cA3BPCnMuy9MJ9z
+F1u+reg65H0i4ped/M9LcvwzCrpIcZ3ee39FEEJXKv0pLOSGJMzGwHg8yNQwp0d
lZChRccuT3at0jaNIxovEKcsxly7rYtBrwW8eZ5OQV1jXJnGo+CaDsx6twTpLUic
KZbEarrf4bSn34vwyqNyFTEw3QI34dVV+C0xppA3eEzWJsBJe9v3l3hbcgq5D3K7
JGlvF1WI6irZHQcTafmLCJ86giHwJLF38dsB+cmDMTAT+1o+p0to7vUa9pT8yuJh
Tdgywo6KW5O89jyM3XuFrjxncmLN7cKMoNSGgCN9/IYfZFdjocK0ARh7AS1KExnR
kD72VVNxmDcuwbYbKcJLEw6Dq25B0M2APEvYn/neIzvJb323aCcN+dMh8xmcKrcd
+Ai3Ab+ocOtiD4XFEJgKAJj9lk0HQ6ZR6uLHt8oDAshmQ8A6rYv7NZzb/7W90zqe
nLdhwIuTvUVJXTbOopKN9p0BWVB59UKJUUSTiPrHMY25wI0r+ygK6larHFVjpg55
hEeYYW389ftOBIdAUHTYyQaZ8GdZUMr7JUlTp4LPEJK06hua7JPP6to4hw9PjSu/
hFkRvO2mll8MoRS0mf1EIke6dEGjkXm1zFZm8wcqKN2R5xkGBrds52QMloPb+EXi
YEOOG85+VZ0G2FAAWZPZelFw7M742uMdt245jatClen/eDz3RoKC8xLHHDnwIFhQ
OZWmtNV70rau/3IKDkYCkDYo7cAa/LxaYSGXUrX6xgCInk1gM8kwy3SYFiAFnIBM
rRf7s+GriDsx3PaIfdtgbAm+esFyIT1IoCgJlOJ+HR+pE3OR52f0ZHGUu+vi0TM0
ao/EtD4CBKZ4hySBdtLu0iNPK0j0mLMqf7giaQlWBrhLsESt4MnKtMyR+rVh3nUp
mu8Zz6aj2OtQx2eQD81IUHSho/Ff9EyOxKGI7vuiK0yW2H55gvVPl86xP0gR4bm+
/6xOONz550H8589mtfiS13UNRpGP2SG/uA1+0l2MzQW6yvPecRMzatdgcg4RoKhR
WZ51UZWW09ZwTd7bZVm61xMOOSlTDeyZynPw74aO352ZtHX1wsvRO+6PRG3d1nWZ
c9dYuHYVe3DJxACZZnETeugDG0but4KyOGbqG7sTFP7gK+TLpTbIqHvmeyIRI3bI
Ua1hEW7Yqjx/o2Sf9idu+QVg1TawRfifp6cknZH4Af7hu9hojW9wmpkBo8N2W3rY
cfMNAgmIkG+vDwrwRTGhRN1iz3l+5t5vlE8mv7/mOuM/2+KrhlIqDe96as0ToNAG
SkwPa5QzCkn18dVbdFY5caJMAjiYZ3OdwlUBFv3yg8F5jrS4qt4n4sk6r1a/5YzV
Y1OOJLcYdR9jizDE8/Q2gTqN8jcE2DtlmPlckfJQpMaqfR0ic+6DzmKitE8NSFmp
Rg8L/7B8kRQOlKMaZa8t0P4mtoDQzAVaLMn1rqkOiMNo9S5T/lgjKpOdEGzAfuoL
MVb6K78u7CPcHNjMLMcfwOQ00MsFcUURTaoUpKdPQ/ZVSezMA3dr9eted8JTrM0l
24MKDmOjkY4mIebpB0JLKBp0HT9v3fTpXyxrseRaBocGx1UwWRjuGs06y3pr8cXE
PVCFpKkz7DIhsrYNPejcFVEsva4C5Uoun9DihOVqtmzebaucRWsZdaGHkaGck8tG
y/x42h29ut1Mb7+tsz9kNLzvb5iySkN4rzqV4pOFftGQKuiB8GmvQmZbaV975XeG
5MH2NR3zED4Dy84CMPA7WCtYoO/gRtbT1o5nkm+PVl7pdWlrG0jpR6zEVGhwOcXR
RiJRzinJYPvDgMu1TDms4wzHOUi3eCr8hQLa+Y5XPE373D3Vk8DgQEeIG405KGQ/
kaYlIx1h94E8Zk1tkNwcdR7HaKXAdpe73Mdx7VAmH6Ghn2+sY7WA+/fPr39z69jx
tcf9Q8TpqZjET0JSRIOFVdszIgqrYbLr3YZM9aKqNpVFlpNyyulXoAFA9GhTF2N6
NrX6qmewFML6vcIW91yl7C85kIG69pDLw+5AQmoBKH8XLzvyiHKTi7rl9hP0ZpsZ
d/5e2sAGIb0jh6+7keo0g27O/S+tiEm1sZAFHApVY7Q9by6jdXYLxLdCbE8SIoIs
6FxQZd0C4Kt8vFw+Xf5iqyAEejmattpKqgu3J22+LRmccCMrdJP1w+yr+QrfQlfp
yemwLZNATMQMBH1iagQZKqOISVj7PiTWHX06XziMpNLf0C/2xkh0TI2iVbPqbJz1
jW6UTNTPPDj4ctQxMJB31TtnfUIw5sHQY0FAG+iVU0S+WEiAKdmNcTHWg94C2v1G
2QyDhupMXD67LtGdhDb+mYmsY38Iiz/cjQCH0WnMZZLUNSW9NgYOr91vqXpIjq1O
qiQlpL9cixQslM1kh+8wcLghg15rU63DNUSy+2ZiSMBIHDnnXt92IOfHjXYvh8LI
5720lrbXMu7CcsP22nq/nOUL2OYqX924C7qmAQRhDFMeg9QCvJUajtNpwdleM9hW
2gpSmgtnfwiNI17pDHn6wksKs4hBw7BplQVWekyEW7aNDDPf8C2SWo3y1q2YeiCX
uG/FaP51KFir/C3G2gOY081cL6TihH9SPgiFJ+pZigQeNJwgcmv4gF172PRUE2cg
N8jRyeH91KvWBxV1aLAx5w5hyOFT3qwOod6mH93Fxx8ymhEXVuO0yPZLEGXLNcgh
aSnIEw7/PC+8WdSHD+vFloCHwV9prErF3cbm6u1WOhJGCo8Z0iuENQQUXkn/zTpq
SYJIF3eDeiojcSlRMtynbvnNClSAzhnrtAsup0h8OcuH/M9ogyDcH77f1Tqcv/HW
m5o3C9PaFql1jtIjfYW+kKX4rf80R7O2as16nibWQfG7fmo2VTpKDx4Nd79U0Jy0
OWZ2WoVsozxIu2DreES0LQsUsx5bxX2SLr1NzeUMiGK0TgiYJdVnNIgxY7tw9qcx
TkRp8l0JbSvK8lFWAOclNVcUIhvCZLE6tUkj/GQpiOyIOH84hyZxGFnoIdY8H6SB
a3bPWoM2XDenorkA9uLTsAfWEo5EVhS3IlKfouiwotyW3TFwKcuWd5jQDk4YdpN5
FyeUCmpLLC3i9O700g15hiygaTSrnpkDlKEAjYbT6eyFzF/Un7iRm5a2KwReLo6c
3c4eztze+uzMpl8oqderqKiiS4bvGg8yzXvV/tNthWputwu9vO/sBx3scmoEgX0q
jALhnEX2a68I7J7mWCHqG3Htz31ifKW4wU2Jnh8SC8MDc6SJz+d1F3fR/iq7vKtN
hEKTV7o8wT5+a1mtQ8217R0jIR3B0lgOpSQFyZksL4dQ6QV4i06NkwV3IvuvQxVa
xQbEPUxGz0E2nj00j9CFz56HGt9/zE1cKilF+9UbGSjkr1f/Hi9fk1h91cMdecUN
TCy1oigPxHiod1/GsUa4+G6Efus4Mtid5sH5hZOuaisAci/UbfmFU1f75IjbN3AF
uk7ucJYOONvfVfQBi6k7NNsFcHkD4qW/qpE3nbYcSg9ltGMAxOU39COHtta7b3Dg
VroH6PEfHR1a76YsrSUqtpIo5AWS13BQMslNAacYUReQH4F/VpVKNOeVNtr8VxZc
309tmnZBhfwxiJtlzP8SVMGH0gfCKkxz8nXP2b9ZwtQ4OdBstSD5gZma+QViT4zg
2z9ZFzyaoMAI9RLC4L8lApwRuKtetQBetsY8OTmLBj56OYEVu/bA8czMBhWp0sZG
nVEFOp6G4IEuW7IE9+1yM7ra4kSyGXm7JYYL3VfvGHrU7612sc2d6A4pxBIFhixI
+FNWWqjJNY3zd6NL/scbe2lHDaqpV24hNzrzFS+jR7rRL0TSAuhhOc0fqigV+p/m
hfRAc6NNsU2mIVngBrDDhl/VUua1ZNLzFFi294cb79koNjwM4wPu2chjY151mDrp
yMgyYiHJoc/ki8u/sJSjHjEUD8ufLl/ZtdUT+gXGuEQMufdC6YXmaD4N03pGCFEE
y1jrHfVgPa4iF9mgPmDgdzCoMWhDFGu62Eh/JDgrFbjAYRTkkVyQbHj1xk/pXbsB
riGHdClwgbg2J/sRHV6iCcLBr8M8dd+JgopUk6ti3ujtz+qvGBQ7wCJYY824rZNv
FgifiWj9UOrvikbYyeI1DYDUeKkEnz3r/Ci7tDQ+whCgUYtnFibUiHgv5rcuVO1A
Ts6QVqn1syG3r5PblfrXh1iyIajyNT/13jLlxRozpOqMZlItMKARBPT9qMjtJt4d
svmmcm9Icnzle7Wrqco/kt4sjvfjvnCOGpP4LA3QNDw8IKcNhNjQuTor2bmE0Y60
3Y1fusUcay7yFDXI4snxGKRrwL3r1z1Nww9ZwVmtt6MxXSRtBwkEEv44tnfvqaHR
o78sA7m+RYfiAoBW1NoWW7454IEVEBuGcEjF1rq9BpBQdmOaPWSCFU/peaOsiqz8
1n6DQjJ8zOTZBJG2SkwLC5XAyjTSvFu1GL+Wt6I/izlgKmzA79J832YFJpzELpa2
ewPk6sgcy1DGvg+ujirmxdc6jn6UsqyJCcj4a58UgdptFi50hxVS2tMGJiXKJQe3
h4cudS43KLp5sDJJD00xDyCCETCYzexF5DUM2X/7cxaCYspT7a+f3Y2+dPwk/tOd
kVHlfwV2fF9KpMG1O6NIQeWwvcntSEgyaZWa4qgKj2ahlmBqqE8pI4AuZjYJ1i2E
dWHhK0wKAre6x6nk4QnyIe4MuNJzUUeo/WAtXLIrQQPEjCisQECG2VW/t52wo/sg
OaTMsB9TVnV/bXIoLVG5fN0JE0hNrYJur0NjsX9et4MejS8GLOY+4YZ47oIVuYri
CSez3kos7Pl2gpIyxBkbDNrwI/ny0JK5yUjlYTgF/IdLDU22aXqP+W31pKKMcj77
AxZpVIgoArspWAlMtaVMuja6NIBiqceA6BgcKC4H9fDH+5NReEBdPH0+zIuk4uoL
yUIF5mm+xrGwhq/ojnKpiepzKGuyTXBzgdWXVXPbGhWfQ08Vi0uuyyiur0YNIcze
jWaPDsUWRjdkFqWhJOuirTKNOKHIX9VsYBlVxlMJXkQ841L3xkWmLSiAW9/yuQW7
XIpMQGuYouiWvGnMq/HfYkfqVMCuraejCr4KZgJOpHjdR1eYpQQOY4+ibht9iraT
XJttt7wsbPPJqMAM9zPGtR61jtyk1AkAXwX4vn++UPGOMLWE/c71K47hKIKF4qqa
BVbh86uAWP9HkEGJBpXGTIMHKKQhFYVPfx0gaUNPcPRqTvCgTIVLe7pOZNdVvC7q
WgWnqLi4ovASpI/+XNC2Tf4g9dP4dIzaCRqZLDqKVKOEk8ZZjctQ6s2na4U0HdLY
4Lr3oKTGclWT+KICE8Dqh1eoSZccPbM/3QPEXujN05fOuOrUlN9A6xzLlVhUmaEe
z64xJ9XLn8oS6ujAxmukYTrJMLj/JEWnzVoDSgE+YeOidoeDTcgmYbfoCiUcHsSd
Zen44zYnsGUxTWjTi8KJF+wEWtCfwc/hoCPRuYmXH3bh5Hm7fcxMa9EzXI9nlv+k
fultw2QZOLAIX0hmQWFNzcza8AsRRJMSA+Xh/0OiaGzYRAZW+dZstXL2nzQY8lKm
ELIMg9nRA+Cqhso2KLAJZOZAqvaO1mpaBgYDK2wGVU+ew3w+i0zXGjzlfumxVrJ+
iKvBWIr/mCFv0quRV7fq3FQ4yA5klYTqwBb4pNAHCegSESOpbigDmhEOwdr+54AZ
qgCYgcVe+Vj+Gj9ARKzFCMISQsMOZ6v8Imb5ie6IiKFk0Qg0O/PvmcAw8OYssd1u
/hEgb5wO65QEWDVH4lC9RAw5FRZXDlfsLGYXf+Gf35Mcd0mXqKy0bnxm7LD5EnlM
CVW/WaaMKcMigVq3JXhjVwH1VmC/4Lnr/GvCmUIXNnWQABxhXwM7JOEFXQJNtmOi
ieUeJPnd/RUvP33xTyT25CJEuPJW3SxvVEeBAzO60vALV4Byo+fa7Qqq2B4JbQwT
V06bvLi/QXq+/fn8UYhNVtjzHd0GnM7/OlDPCxpWDtooe0pnhBySNNEEtK7DOnSY
5frsweFhGZhVs20OF8U/4/8Pa0Iy1XVkn5+2z6Y+JlAg5emCH2m6RR06kyJATqjW
g6Id/7F/SyTphTVtU0xB91ejWs1O5XvhPsQg1zh0G6gcIQ5MPZ1gdOT0EidmDgNO
pskTEfLJcuPM+dYXUP/17wacUC/uw9pn1WX+AHLdusUSKNu6eShw0VVObFyPjz2k
3BLWttgbT24+5XCN9gz5BWMMIm4CelXfB2Igg/L8wTj3Xryus2UAAbwCX5Kk39uD
Q1qH7QNUWz1qGqu4P6hTMJsfF0Za+OwrYXDlUMXFQBRhGCkIGAoxk7gc0omPUNS/
M/K6bR5cN53AO16bMefxCXF0GM6amgp4Da9otoKzUQsxyn0zqKbclWVvDEns1C3y
IGgxpFmDLqXxZrmXPn9CRpX/gsM3O4SXZEEOuyCiXPz1Ub+y2x9qNDNdNsCT01VD
5b2SoDH4Qd2LhqhVebAbha0I2IhhATH61sNc7/98/QIKt6TdGT58jwTtQ5bbHtHd
RODnqUSS9NsIg1BRR8IxjIOUmDIOrnT0yANCiNW1vD8s5R+3JHXDU8llFvvwpiam
VVv9+QtntCMimToi4ozY/GTcpmfG2t2Dpk2MKNMc5CwVONIrD3kb44NYFJAJE5oD
AHWZzxZ//XQTeI3Yl9FOGuOq+8gup+ukR979ilRWJ0ZKZFArsps2sOEqfyuYhzyc
BT1uJ32VLnxyIoDqSKXlR9/QeM7w49Nv4Js5ZFMbho45pdZsWrlTQTwfCKLOprc2
mDjFAv8u/ArIuUNMvkH6kjR587fUmNoqN5KGWuK1NPB4R2hSm18iKknLigGRMcn7
oY11EM5VHOQJqMJUhrxgkjclMP+ANJIP0gnvmscHTvEIrkdieZUNfJF/6PFV77iB
TMh8ymbIVGqz6An310IYlWJf28ZrLo2JXVsBP2WBn4rDKWpT0HHh2jyzfBTxXxdO
lLVjL823CJEsjoiu6iCu2mVjctSZifEDPQYJpbxuOjjiWKGB4LD/SR9nJnXBHpUq
Tk6ac1jKcqVUbMg+R4Zjf920aVQ7rNZJ/lQh0hccc+GuSCJlAe2AjQtTxRQkJ9i5
oqXoIOl2g/h+w1KBesg90gfTMasD72NfohV5ou7vsarEtP/Gfs9HTy9i+BsiEWJT
zpaHemNVOaDCjR0zinHRQJQXcvtJlz/lYedONVjGniNhPFuJHKpqqjoEsR//SQ8e
TAI1xNPfSaGa6YOyvW8NRxJK+aTgGMWl2bDRXR25rQCufjbk+ZE+xedClwNSi/fr
1Gr4lQC8VwaPkqypDpQVT/OixGefMnCn9/hVVqHubf17eXepioTwhMQJAIGupKcT
PwCEEuXUthScw+Z2590LaJ7DthsxY3E7LwM3RvVZ8mz1rQ7GZH4my4kHTnfE1qvF
DmeLQ63ynvoFEOvi+vQ5joAIEkiOu8B3pyt6/WHrqDWISEJPbpYVxXaZtuVIWEUM
gUj16XLh397YDQ7I1dpfKvhrOUTQPxsO0i5DnPZxKz932uhH4qJ0m+WLbxL1CAHk
0vBoWMuZlP1dVmo4LT7m+6ld6LKsCn5kbDaWhBpFgRTIB+BU8490zttnpslolAjJ
N23ARGmuH2qiQAvDiTeSA8iZi5/UKM0TzBxejvd100wr+tmWxGOONKZ1enmICql3
NhOZSyYZW86oinGhrcn7yqRXTn40lgUc85sfB/Rv88scYiRZ0rGwLVQFYt3KCmrr
SlERlJuN4FkY0DMXzDW2fWy7k3vsJKSHlIT9mzqBq9Uy2ToMmfQq7UZ11SG8DGDH
A3bQw6/cHKFHTuOLPx6yxemPvpz0CdAwfSRQ3BZ0V0hy/74o3LV/yBR98glx1igY
mxLaeITqXnjlfrUZRg4xn7FaX/gSEYw3iKPitwaWoNI+k6Jsp1FjWk+9wJxFxtQq
6Nb+K58pRhDt17pV+0LA/mEn0/AM6Xf68FBjeNZGwbbVTaQ/g0HDTJngiOs7hs95
ZRkinxBsE+K0+1CHpb0cpvLyu7DYSAcCknp1O8R5sc9nBRB7WODb/X6b8wzl5WEl
ZdeVWf3I8we+ANRokm4mot38xbjZkE0CmHOS8Sj2qBj6X23BnHNMN2Utgkpy9vV5
jXdwqmBmpZRTsAt+tWa0n6B18YotvJwXahk5vQiqcsYKstV2Nv3aWk1xt1gbvXya
dCvTBC1/8MjL20Up03kDRRLYjZfMpD3zpM/mB+akTLJT/JdfflgRKfucbB++yJvr
FyRo7TfONG6c7EZOAG8CKDfmOKLOo5OlI4QDkj8DK7jV+XoVFeIdOHScKeNLe2jd
THqEB2bJd4LqXjbXtwE+IWq6TrgfATvBIArOK4UdLamwcrhq8tSibDPHi5gkc0c1
rjjNYuiixCux1EmEhrdv779C+R+YCmU4mnGZefVO0aNX4Tand5Q0v36QywA4i55D
pu3ZPsylVKa7e6MPTz5iGDx+UFNNC/EK0y19RFS6A7YxeFQIOvudfypurerO1nD3
1KgM4WI1Yzx5rjsvjot0WiCTJxEnzlbp+na1ifpXT1RWh089Tnc43ROL15nXDlS/
72/SNE9xRTLSkKciL5+RptYtspBhPjrjJsXmDGhQlC8xAC5OkC6/mwpwzSxwFhQ3
MzJei+rip1W8j6aXReCkuMru+FbPwyjt5BCnZBQ0/Qo2R2bAkI1JJX1Go5EU68OM
gtM+RZTSQ3iq3eOczQ7uamalpwvBN2MgDGuw5I0bX5u8R7NwbVkkZoAEMoseqhBy
KHQCoqkgPgHDPqO67G7ZYq1PDZr1Qn2RVBebKDboBWhSydmykatsZ89Uy6dVUZBU
D8+Pj0Ddt1lVLLXehRNFyUGUQlbGsN2eCEJu8ViCvk/dSeyf3SkJd39qQYGR0ykF
l4hU1n9BuwQUEWCEixwrC0AFWdu7txJPV/LxxsYk2HLmsZsmX9BXTZ72MFfKK4gE
ISIdURoADCn/oJu6qh2w2zB70sXZi+7QC+ydmjyewt0oUyWT090WQ6+RxjA4LSH2
H4nZoy8DusE8ljVL3vOMVnCBDwdsyg0ru2c2l2OYzgDDgqQkuY1f7A+fzIRIkYA/
UwgBBy6Iggm66xQPHWRhVlE4Qc6ca1bDZYuwoFiDtNlVrPF94puhKjKQGJ1daJMa
ML2AUJckhCWjo/QajzUY1Q/hbiGff744U8kSDAAKfnq6ruK6OICZifvMImNK912v
5dxxe7bqeFv07Zm+lKQFjpSH0JNeyhP9coyknjCbo1qK5R1/b4HfrX5QOi/BTtXd
EPS80z1L2yhf5DaV+tXdPAwA4UlxfOY/5r59Qm2TAVEw4zwfaoa2i0PUvUUMIZ1n
yrpA8/XNN9g75nODJep3T8DKGov/+zIIK4mRDTh944LBwMeXe8azUuUOoGaR4Zha
0RTwvvq/WwzVyLwZLu4ubRsjz/47CfZc8qTN0+jmN+ti47CxuoTsD/AHWWWwbsQM
ayDDwEFu2Ya92W6WHtYQCogFNCz63MHH3eFwCaaZgejHEVAP6jexIJDNHZCjTWwi
3UtUkyG7PRx2fbiMu8dvX2M0lgJxzmi0lHG3KBlYfr9ILS7vvWlsc90WJ+BXQ2Ps
n5LJOJHlbJNL7bS19RAcBe2c/t71KONOXgMt1CplivzYFTzevwQNf3DLnLBaKlvc
l0zvLSi2NVOY5O6W9um7kWHBdQJc8IR23rYB+2lMWtGXiV5ogytJePJrVTaYF7M/
csNgewyJBaLzbGkDl83/E2L6LzvrqndJn93WjuuDxufTGhEL3zHiE2WvEOuE1cAN
KR0acPi6E4ptDZHSm5jZtmYuHtVyr9PkPJkQyBg2O8A7jRzzEPVf9py96oEO5BtX
FUORjgTdw7S6I04umN2Skq+kVijJPh18HQO1usmk1YvqU23OGwzJoaSvpxPMqgtO
NAyGc5N3aIg2iTrvONF4r8P2xo8F3kqg91uahyZ02zgdcVazSoghi0dNukcCm6Tf
oVIOfMcgwDwiMVUHLneWFCAvw28M/A6TBGjgLPct2gPveEeo5zeDkbGtWWQwuKY1
smFLWNlhZ9oMe3v2gKuasKKpskGDYpZ/FyuYsY5S/YKZapRbjCt9g4WRMhbg/9nR
9MesiKl5eLtuH+q0KAOtf+fYTP8yMaG+4reVyuS9vNAsmvHsAc+wx3B1Va09yC6V
RlbJ+7ObSknw0C8GZ7lNvYTUdsOu4fi7jatLhT0nK+LtBGonss4xPt6vRqkY3vPO
yCKaQBFDywRgktrjfHHSi3ag2dBoRBAzR+eLfdAnWrOwAfxU59uI/Rd1pPFmz9jT
epDOUnQdSApjo+3RpLsyO9qddzkd4aXDt5N3u/xoDDUbVmMGe5dlt7vA+oa1iW5F
J3WY5OIRXH705DTcEjvIWp/AIn2GNmXRTNrtaERsXd4KoUSyv2XLIaT5ytKASrVE
/iRiAlAGeF3fs4Efrf+ePYSDzYwCx4xEjg5gyxaxq18vHj/BOdIpMfQa/yarrLiX
Z+H12qub8K+tk7c9hwkIiAyIoUucp/Km5r16raxhKAeQRA6Hhzw/UcpGInSAbgtF
N/EGDDzIypZsTbHyJcjFA0qzrk+rJISGethSWClIzxxon/di9tKQuM93UB6rDrJB
HAoBaXRZub2M1TaEU+ZUHVdbE/JdG1zK3xEdDD5CjxNUGGToZgXRymObDQDk2eLG
cbK0R0LFm/94R/gXgTDdsCOxGcW5nn+hNLrNEc85A/u+rTu5UXLIhpV9iJPNXsME
S0HvogwlR/Ri535Ry875MKOIGrRAf6IbDZrb1eZK5ixZp8HUpycykIuNV41p0C4y
ICFoWJO3g9lipPEahgDWr8+c3wATZrqs+ffqlntU9ShVMwQEFAH04WKPCj0v8Gs9
J4/81DwzqEmZ7DIkaCrWlTQo+dCTC6N1MiBReBtYlusXaqd5bGBIQkwiY4z2XhXB
qj9kZ2Y0UAg3JBcM6iixOQmPOQMNuenBMOd1XKe+eHUEFcfMYIA4UgMWTMnmzX2V
F3ZeSBmavJonkd4A2wsV0vvS55THYrf1DrSTXXJufxKMX5RljA+evnXe0J866E+W
u9DVKyonNKqIn/cNFSE1aWpGshO/kHIPzCQOAc/X/EXP1uyNYrO82MdrpRIutu7V
/Qw9LFMbRRBgHWL2tGciXMP+NYjIkbR1rQ7HpoRvgTwjGOj1pZD8++IHh7emM+Yp
yKa/B0XrKZePDcwValgXQ+HtfXUQ+be5mFjZcmu61nTuoYxrWgInj8Jt/7UFKn4o
YEgibZbC+NRVvumGCKtFREJLrodHI32piFvz0L/mJNbxcIhM0TzBUF9y4TLmi3t0
1f67UvEwJ7jSoMUjzlIr1eYYx9UCJHH0dpGplohaPOF3+1gS0P8+NX6sopJn/6yV
FipejufrAanwRivQF6VOPWhMpsYZIpMVhDtNmIRcDbh0KQCf9TF+bIFFrmpXBnsP
9HlDlAdF1FO+fjbBA/5tWoxhGlHvRC49lQeRNeKGNgphBC/CXCYRJBxqiUFhKqlF
UNaa1cSBlQ0p/3y7aowcAgLL9zZFS4JWVjyAbkOC7He+5Yg1yG66wRvIAwImVdq+
yFzjdaSK2sf57K3g0pEtYRMtWyZDMIH+Va2MTkEnkpmKgMW5Rv+z5Ce7XgB8G6y0
f3QaidR53+ISXdfSl8ToXG278Hkrq1sFZYVFWZ6ZsxOHosb+NB8J9IeTotGR/svi
LFzNbV7bgRZh4K43jICnpBozHDR5FbDxe6bTTqOQdh6mDtRbMsghM84/Sr3u3KWx
aaM16MWT3cd2Vjvop7YJTzLqX4FEo92LsMxVuuykCZKMwMiQtHSLwSTSSV1f7Prr
YcqiAjhFKis4ofJxV/85QFrhlUT7+QwuaLp40OQ3ivQKyBUjwZz2wRdP4VT2wEn8
NZyPNUZoNK0B2ehj3l58M1KzGeLC/B94CMXaXQgwlQN/tUftPmFx58Fpqroxk6NZ
69UZKYGI5kxoFwiCIfT+WQRvW8YDDBt3GN0k3FZWDF2FYq7SXEEpuICblGfYxqSM
tBkCirO4botpd/+OuJAq6oWFTep8bewPPUgUCaaa+YXrNo8MC67ctwlBpgQhNX44
DAAnMHW+HzZEfSNWqYwppACMJyk9vKidhHUsG91Hmto44435CehaSwtPAd8xLA3a
ezeHC7/IiycB15oQdfOIg1m2ilihh/dnX/AlJpanbL/RMepPAjvsQ/dfConXEHTa
e07VpMEsTW6dU/m549rq7ScJth4Ct+9RCU8bwL9AVxvtNl31I39BcCXy5icHnuzb
WJZaqwBiemiHL+48amROCWfPOHKxCqY2btHyX/qg/RfFLRZ+XQVr27vDgKakzvTc
KUF6Clwvs66AGlolg0VQrqrvNdqA1xZfWH/gn10Xq+Z91sxLnRZJ/GDcxaW6XWP7
c2gCXjDBEY4AZ69Jn5PGfNKPBy/Ky0JwNv9dWA/XOopWlM7GN90SOOCKO28DUtG3
/YSGSh6D4CaiJv4TAKwnJQh3xrIkT2sdJr0n1UZhAyhszQr9baKsjXr8VA3WAxL2
JCU8boj7gef5XWCgsUX2kiuBAXSwBSTxsAKK1WYIQRU/CsuU3z0XjVKIRa8XnXg3
/Vys1RnCXGLBaw+vm8AI8BW2vdQJ1GfAGJ1LjXj4vzMBzdChff/D4Xi4beFUEhRn
JmJ0KaIVM3XGi2jLA9ot28uVNAX5oiIKN0pi9ywE4D+LhODv0zw4UzEfMq6TdUwH
A+1YVn7vbTzv63ZgfDF16qVYqrGT7/sSf9dwT7EKuTLBktR+y/qWrNLc38uBkBpQ
VdEoj+9Yb6zfEKa0jMgjwQob/TXf1GxEkXvpB6F9kMM61HvgVqPb5hkolUmHnwHG
5jsmHq1aOLpa+bxcSg8TrtE6RRPbB/fmi3Mc+Bt3pUTCUV8qhjwyTnMoXCRqtuH9
xv0OX/8QH7Q4K0Y5uszdueQgbws5CsBTdsYk5w7lQMJILijB6t4t6J8SxTY8Gnhc
jjD3t5vKpXBjL7HRWh7z5ZLIRhzf2Miag6wV3/iooeCRUKTUDTXRFT9INsgfiGDe
BQfbZaZHr9Eh6eKJ0hAfjHPx+f2a/GqoXQHgAZ+UhQ2s8Drxh8OlBIjZCADwTRu1
Uf4Ws8tYaDcs98te/WapGeYr6fIldIPZfAcdU+h+hUAyG3g2x/9JCcoaGu7b+oE/
sJQhwdTY6Kgzo6KpMKTU4ZxghJv00MiYwXsiPuwBjsvldi/rAbwTanQCsmPHKK9z
wDsJ9+PiCc024rm21MeJYDO/q4vjFBIiYeS+0DkIj3kTE+n8YMpTdhXrat40fnWu
ybFYldie7MPRMyXrc04yeXIE+bGOGJVRquKANS1SqdNNsBW4UILlJOyGyy6ASWVu
KvALKpc4axIV80iWMnCYfPWT4JacJTt1Xdv+RRvF46vElqbb0l9v/p0FSlEKE5iz
RaskZ/+Jk5ucARDHCY7Qru1zEHxS86hMGnWKK+fgVxtg80bSCA1zNM/uj0aMMhf9
tSrub+cIZbuKNJb/HfDnvb9nsXFLJ/hDuX2mPsBWbYlGs0OOVOiBErrMlH5f2m4d
1TjTQmNFknWUk+Q4YdHVgKA0N3imF0p5DQJeVCqgslL/57XzpvlhIRKk4xgr/OFe
IXSuj0Tj8TEHHsrM6lJH0MwE3qJYiFN3dNNXg8m5F8LNpU8shzqfqxWUdgM9z3L5
/kNsqvtl/uTUS6RCHOhtoVUek4YFLwwiWIPTnxq/ak3p5dP7N9pjK3r0zZIeF/Ct
d6eG0bJfbFpm4t1Xdtm0IWTE3qzooQjdzrXa0KrzKVgBUzAV0gOj1zP5+ho3LaOe
FSCXlRHbtFoNpxbbnWFKLJgt3y0TLOuqqz7dgOTqzUg5koJOllFn1CUQmscyC7Ve
m6TVWBZPdoYizXH2Wi6T46JlgZe+kd2O0YM5Fp690R4x3hKCCEu2kFftILJO/RRl
2MP7G1rbmLbjFJUcNFFukXFl/nMGbiZNC2MaIUp830ZGoGEbnQ7vS1PM5MJsM5SJ
OQvUloltqhZAOaDrYGzHfAkm3Cjd2GbOfX5wyxrBRUgKFPdZXChSCLm/m1IDKx5u
yNVx2aYY5BNLSOFJyRDpUVfiCtP8fCgI3SHXpGkODLYo6zTtws2o3o0tHd3pwKFl
QxH7wlH6XObUeSOkKj3bPm+3FtPZAPbwfUpWWX7absUBpb5vrKxpU3iBtHcGHj2j
rOPCJoW8e2Foh8wPmpbhvUPGbix4KQH/+kOXwWpqmcRHDHZktgVem2fY66gLJ09u
uzAFFqkIFLM1ellt/TaIWfejr2TevJIo5d0kt8HmTfE2GcuNq+DJszObGBlBX/M3
sOuFXfM9Ve/C7nWRwVa7aUrir1bcJPPeVAgQZQ0ipRle74w2kvXxYTQswDFQw2wM
yy+jj9EYhEcYmd1makt2RWVcKt594i3MBmFB4EDDRJXTBshtPq0nApcuKfrDwVCO
pzX1iOQZE09UfNQCnapA3ca3onYNdn0Xd5jLOrV89BKX4FyQPYQUc9t7uKVD4/dS
Y8Tgu8Z8M1Id/ogqOWCphCQE9L464l3UwzO+xA/8CsjWIco3FjGVfE7Kw+rKvhh3
o8b+RIxzbFog+fYV0+Wk4tc0pj4gseC/G3+T0hCSeCAve1xtHHX903puRFW8veri
VLPaOdh0sKIeunPx45eOVdDQra4h74gKhVycfoMNLqx2x6kCm+1ECxzIa/PshJFb
Ym3trCSNMNWGnSw8SB6eRx2coqQlFKbu6zSz7AnKKxq839wBThK2yeZKqRhtSs7s
zewcoWMds6sNmFm1P2gVnzKRtkR6dM5Dv3R6QkGQEwmBU7smp2f5O1wjZjaL8Bog
Y1H39H6BhuLSKNRV2TzC5bYzZAVQ92lSEHgp3tan6LSAFNePB/XAffol+U1DD9ug
9fDAzf9UpTXihXpA1TlZ/OxepWWpkzSuG3RAVduNVz4DgsdsyaLjyTIUTVS+aIcz
H6egeUOs6MK8iprsWcyhUGCmWL7HsGPIdFayCurZeeCUDXb7QC6ya6FueqISjiuX
PG5LzwrTF/8TVPEAYnVx+AjaOxBj3k9NFTP9f9fpIu5Mkk4k/+5ERiZxYvxcfKul
aWfhmtlPtfuxP9WJuTkxE/4KdC/ceqFH5wc/p7VJ2Qj+7RAfQOXQlWSmjMyHHhlY
wPs5egP0ov5ZHyCLx3B6MXrbpxpWODBGSU5ul5YHR80CxrE8y3PN7bSeG/b3kGD9
YIpxkqoIEELvg1gvdHcFyjHL0iJpcSPpdlyMbdDyTtGUSAbgm1fiMpUkU35culai
2J9dmjoEHGF7ujM/PgtLrx5af4ZkAummWVTWquoOjt10IHzXTm/a1PEh4xlqMK+0
OwsOQNiHd1lEl1Yk9T0914xauoPzWQMysTuLw7Pg21kFeLceexXnoJ7UQ7HZnlpx
BRjAusqf/CIsIgvruc98t1fULfWxcTC9DSKsJ/8chxYZNs8qOeM7otbPa7pXG3cT
wBKXXFGvFRUXEY5SWCg4v+Dei0abM9XIZaGRv9QBVJsVVSTmmsqchCRi0Y5mcvTb
nARAoaJBMEznWkS13HPT6XfXIr9zOnkuz5jTLWegQXIruOPd7m/vX/OAINstRO4H
Aj+0kTGRJBjSvXUIbtyYsqoJQx5vrohI62X4Jsb3YU49TXqJotjbhRlUP/wGSqVa
OjTkmMCSvZmzoNs3ztVtJA6+nApNry/Nw8JEJ5ejKIC5KHqj/KWSjfRNqrc0MQR9
6X3TYQw6PC3iFFhLaLDabweELRKBaLGTOkEUnZ1cBJyzTRUw7Q1wcOftlretZC4d
+ZFjr/K3UcZ+2RpxBrUfp/t2T8wMzHOL4XqE95UBdHUv9nj0QlH5K0UpvrKfM3Xl
jMbV79ritTMbP5IjY5XWXfdhzl/ZCZ9YBaIicAaqOMvB6+MYsoXXI5xjh+I5c3qx
/RfcE8QOMEZJ/2A4VJ3qB3t0+lPodpMXsMBcec0NlNIPKloQUpAIneRBpllFxC93
X0VAQ4+vKPVYsDthulecY8dQeSD4Tl/s1blSD5ftabBRoj2zwkLxdEx8soWVKWO2
X1/2E4BNt1LkWNZ+NLAtbI0Na6fcPNHtM6QOFGQ89iASHkFqHdpK2jIyMkbcXbCv
GxVLrr5QkZUjrBPW2NxlHJRJClcvPc6I+pyeW6xyBsbONTWNJiHPujV/l8CvnbDM
piTSAEYFZlRprZVcq4YSOXF0vc3hThfE+Pc687kKahKsOePAUXSGWwAuOpDr3+A1
n7IkctDJ2wI5Bbthu5RYVeAy23T70EnYoWzwGQ9yN6xZf+NeTJn6L/h/3Qk44Jf4
WsvloOqK7w63OVMk01GxR+l3AbHvBvEgHVjeAh3NIR3YYlY1Q7CDzKnMQjpCDqfh
jLGc8DkmQv6n1YqgKWJHC+6o/6ZjaotvrNI2s5p67rDUjpEvZG5FlUfrEem1ZlmU
P8DS9j6sBlkQllYWPFhbvIUp90muo0uLJjsXcl9e0rdx0A801hbgqgsSUGC9lOP4
jDyKXHFQv9/ll6Jw+mo19XlcMdA1EzI688UCvGW5EWSgYY7wplkf3z7mMq4vy65g
gaGCpupj2OVfaJhWjgy/uDYhosi0Zct8meIMJWysCMrK8G/xPYIoeEpnpLTJa7lv
VfALsdaA9Yic5IH9qMVcfSP3RVC+GP+MxgrcylqyPK81+Pqaqdh2I/3Oqf9FrciV
2TgAIkI5QAubvHdVAw30nifzx+55gHxJwmjvfJLZAwcbGQC8ftTl9z2jI26S+A1H
CWdtyaaQGxCNq8nXcwHui0CkpAZQMPkB+wGeay8BKAkDpeUQ145vCF7KawU22r6p
99ME++PTqTSlYZai4YbCzm4Js7L4rEJAk1jWCaw/tlLioKH2O8Y7CpRuPTKeXgSd
TG0WxfwhBKsVuuwEVZiWPwvKWd205oz6uPC/vCTDL25fZxmRWALVw9BxK8KQzNlV
TvkVkQ6o6u/CdhcM6ohXOeKWuztMDn222IVTRq11YzvEIa5IhGUo4zd1n3XcxpXB
kKqWNjDhvYseiWkjMqBiX7nuEiiAfGhPgI/ULGNWl1M0lVuNRnRa47FrTkbhzKix
A9IuZnlNQxdKssjYSq4vlWDkUqOhuqLSkFjKreaXJ8WQo7q7QSILeJsEQCLXz8Kg
hqXAp4lWLJmgEzEhrqfleIFSI0skScKHiufAkrlqyD35HiAimSehopmlcO7A48BI
zG/fIdk2rx9a+eHMfkpJzRZb7isEM/Ac/gzGaDdeXMpTh7+dgccx0uv3W+17UfS5
tDIKLc/bIPShHr8g96Zmis2+j8szTmH1jdrDDB7FOCodXPVnrjhRX2XtTbCLSoNX
vn36L/Jng7HLUPHFEJVu3hNLTWdMssANLFxzjd1w+FSo3xlKTSGDCxwjRPZFwYJ8
eM/A7fwrqcsp0gZGHoiourXddbh5V6U0I+M0aQUzD816B9aBmx1kVjiGkGQW8ybd
8F8mPSb6ccugaxeK6KfJHZjWYIz3i/9kQ4+1ExTD1616NdZnY7Q6pWHgOHDGyINg
BG/Gbu2nfpbx0yykhiU9kOb/QLcBMU8PgV5NhmOwV0We4fTo0c9+m5XRUWip366P
AdXDpy2YNJ+NCamYwHJ1PkMifzjLcGkN5xcxWvDig6Y/na7I5/klQyFZQpKFhaps
khuwI3KlUxtQOhKjkbx6C1mplq35sCer7PpdUfj5B5b1INzeKzC2CvzPGSpbXS4z
NaBzWB18wEHcy5jA/aqUFf9qQIxt+ED1uIwUEE33J8xf7b4d8wRlmCGf/GsltNp5
5G3wpBzjTCq28OIZbugq1+5EpqM3O3GLBaTW3JFdJesvQyk2mMLnFg65RlgJo2n4
eJy1dzXuvsbfRAh22cNcQmWTm1aC+egS43uWZ0O7Sx5q7S6ukEWi+5gP0E3aqlkE
olowMxyIWEoqXZJrY4FiojKMWio2tPURzhlo+ArQTxsA88kbFP6F/hCetUkBgiL8
FiGQnVces+faALqdO3aOgsXMLYzBdx3zB0AcrWnC94Uq1e3gAsSMGyCSVpxhRURz
j5k+3aIiFywRnOmhRKhYN0oNU4WCtEHQHt7vZcFvmoBY7Cb9sZoOQ6CL+U1sqx9B
wLv4I/11DB/zqaiQJ0iR8aLGgMJrAnGLuVsqhLsfEorSTjAanpHA1F5igEqXHq8S
Rqefk/ccERinLyCN+cLMlw7WcVn5ktEUiu7Wsh1ymKCY391weL5/qodSnzeLGfA8
D9kZ8fkl06UrvlvlcZ4P+iLvvfwzK5DSWBqEIt3kFuKksN96v4qb0CxPFmTVEN8X
PMs+uUOmkzKmfsvHpE0i8i6HPl6YmfnEuqfyefW/ungwCHWQ1Orlj7OppMTtL1qp
jUIUrvL9iI8nbEDheWExsO/fivGYov/OnKaqDFj+ZTcXg76SkO2kL/VKW1VB/+iS
jP7nXJkt/kHUiK1Ty47vHK+n7hE+b6NMaDOriVIJhGDKZSSpl8f4ELYWTKqWcYDJ
5np6SUUNwbsR6R3B/rEVgDardGv7BtoE9p3au871t+3RvTl7qqZVSy7LQ2Tnd/Ds
KX7jhLvPDPZpD222Nf9s0mBGFYVwE9ayw1DRyLJ4JV5pxHsApKTT0aHK3xWOva9+
uzC+Ux8tzanOTl0Mzpf/N86PpAJYO3mHAG1Yq3ljuxEVGwkkHY18ICTJCUISRsAv
NErWZ1FXoJvliQKdvaYa1rHxEOXQzDQcrmHljY8FPkyOo6TM+Rw4IBLuhZclFxHG
V6RZuKGHcTfRk/d9nAlXgIyw+EzNGJAoCf8GrlqhrS2dOGijqremFlrces0XOTLB
DoXAUxeiwc4YFgvjPBejfELVi8xpNihh2i8UDhNNKZKMcqbwA0IxYt5bGm4k7AJq
LqkhCvwkKchXdKI2xuG5QJVog/t3lNq7KGkOyqrg8OPEiW/ZhUi5NrBBFVC2vMgu
UgPQBow5Qx2Rb/ZMMmXyJQZmoMGmw2zhmAfilI3uLddB6N27G/kd9X5r8L8QS2Td
Kml1xAqOSC1tPMtgBI2c6rfHSD9wI8pnfB1zpFr1G/6CvGAuVhUF4ewtYOIxC6/H
dHOVWgFnNAHuFe8rd9ks0p7FoT/3vt+uqVUSN6NPEOtvBr67GTtkuPak8BoB5fTG
U1FZ9a2+Q2fMTvO1S4e9fkazJ2xhXbh9ykYXi62NjOxXWPEjWd0RipVDmTRO9R7n
mqsQOIGP27SpK9/8pPKl/Kn0py1jDND4UvBuOn1BY5MsOCQNw90N+ykOczyyHnJ7
vZqakuySbeGVDlgl3rFHbTE52EA4dIQHMNX2SFTToBIUz6eaLN5so1GYPdo5sjF0
QjlbSOnAH3pVsHLZYbGpEWc541a1UCVzB8/V8EUp5CakPmR3TD3mcWbHqAgrIehG
i+7rLVjvMZ+/bTVaGXEwSWQaeBW/XA8+eVH7lGzfgPM4MrtLHsTQxmCmXCcKzM+t
sT3YgPY/BMCWtGsZ+rXqcO2un7HxnTXO5EFx+MTrRN1dt91lTM5j2/+Zq9f0hXM8
4XoWOrArOBJah2qQuRq4sGvPB3cUlYZ6vdqViDQj/sdZC2uvnRWdddCUJGSZQ4pA
x11UuU/vZ1D1GNGYmZvOaLXxNgiLF97nkEKoJeYzeKjOuE2piRrNoT3WXLS652mu
zapRMDQtgnf8PnectBq16sPXarV0A3ouHAOQJhKTSx/xTph4gNRoi+B1jBJ8YEb4
lA7opKrzSTYgt7hCzZaF7CFOIZBJZK1zpkxouzlLBLfPaNNC4p8lsoUcIe7BO2RG
aiencGO1uARLxaktSC7foJvmbPv6LdMZ/if1lYbfLosmsyHVvvPDovAhdmt44DGa
eNDD2rht2c3Nhn3SnvWEKPDWZ1pPRhiRKCrsNIp7IvhioUYA0Ib4I08m/uNR4Qr6
JBJ1M/SKAWDZro06dpg9445YY5OfQX+8whM+OsiSkP57opilnOAsu/bEBnxC8v4K
5W8wEwwuKuvDbgLVmBnhBALsC1Rj4MtOv0agejP8NLeaTXyhecc5prNboVNsF6dY
lQan9LszG8I3ffF2/6ymuv8Dot5VcQtp6zPNRSa4ziMV0JPn4MgIKD3VPLg/rkm9
7K8pFJ5AceLhkJT9Q9c6JjOpNlRIP5tk0XhRJE3ITjkPf6vXe5gnnCk+G9GI2hbo
Js9JV7tzSoRupCgCCJy7TRBN/R/RP+8JopI7kgSf1hfsSuDK0T/nOXQzQvh3hD4B
NvtAcvpH9y/cOhdArccN+cV0hyzQwTiFB4oAW+QMeNSLq1FduFOvi4fAb/3hHHO5
D9646YMpGI9xNuTBO2Z5wSVRsD/8Q+nJKm8JtyolJDJhfTbFCr7kyuH0GsVP/Zsz
91HO+3xsPYVEHyce4GfSwnV+Sh24vjED5PKOziC5lskKF4sMN+95IOL2RRrh8ndk
wJzo7JEtnYXE1jNR+d2giInntdlV0t9Dfi6tKMMBiETC/suEujRSWLzWyPD8tzUF
EmLp92sIhqoFU2cI/nKIsRcExEVdF/L+L6cbV1fvaAl0ARfllOxaO7ctYN4zWF5+
WwS83B3LnVcxdPZ/fI0+yEIUjxszdJkPtKgtgajZMd+dWMHi9nZtNkY5yIB8Xoj/
pHGeMKMbV/PcOMXhYf57i3jNNoGrbo6PS4sDsQuaAjKsgAV9AW6jYF46I0ybK8H2
urH3YPWC14YwGSzn/VUoqiON7vpAVmbgMFIl1hWbI3birHOWlmiTSb2GUTAy0fRS
xaYGx4WcNm3C1i4E3u+8SRgKKwSrk6cRbbBF6RH/KJYrDQMHTrg8qz/EV31K4WMS
NBkFVreaIN1zOgIHte8te+q5lDC0kvzw3MAC/EPsAaGlX6HH63Uc+LhFAI3Zyz1F
WW7beXBov6Stj/QluFuRpb9bbog2rH8g7xfxdvLku41+jfGSrahvqtg7Cvlcwh38
mGD1QvviOh2ItpXXB9q8MSgx5RZx5NoGkBg/C1S3rzjMl5MxMgyCHAGCAurNXjto
PVfGVweboxb6NLR0aE7HDXamDV7eWReL/5eCtIYB++97UW2MTj4bY44aE1sM1BhI
sQGaJWuYVzG3xS0JY3n1F3Ya5F+gTp2ei/otJZnXorMiido9i6uYH+i8iJ88fWRF
TtOZZlwCcl8g+3TtXxli3115nqvYD8BNSelKuwc5glDE2cqs9kwBZIhhYwl3+wcb
RCOVKtPVJug3PzRGgyFKyQS6QSEzQM7rz6Rc7s+EzPKZOKgdu/qtbyk4S4TRI0IR
JKICShdrzcQy2n9imdsp1xI192enF59jP4nCyD68/GLLEZZRUlT9u7JqTxpscq4m
xd3TCKuApqobJdQdasSPuQAFe9JXAUi+737cM/mGMoTfUJGRCXTuZYuw3oZhHmek
V+WtDjOr0u4BfbFMlhQgINSlgm3dXK6Q+EOdKLknMEWCasosQkwDRPtPvhSoMzVr
+I3uiqxZsQA0LcPM8VIRwhGcHCE11IUF5H/oBadFWyvRvX+8Stq2Uglv39aDqngT
4Qb79VQ/qQ+eug32zeWvyPv3ictD6FPvApEFkDECUgOl6ngEJlhnNy5KHDY1MFcQ
PfsJIYyJgyv4T2dKvHkmdGg0h91mbWdZu7U5p3LbCsRJiOOa584WCWCConvNPe8V
ODkerqGsRUd9xOo2bFqA6BxWXnEaYFSzXA74N9qtECnMXJtLSZeuVO0RxaGPdsIR
5DOAKUhZW3aWHPLg6dipheFhQFzrMD13DdhPhXhfIn9R5VgnKkh+NNIzsam5lcLn
I1KyvA4jJIMspqCQ2ZwjlTX+xfn2tkUg2WqK1kL3uw6wOrZi6iTOG1GHZI/Djccg
UdeS0c6m4QeSptbN5uJX2e9SAHbwtAPC0GXN/KF6lf1cK9jS3cmyhhJZFVZPZx+g
pIXW3sw8/qgBa2596UGVbkwSC1LIZiiO4TxaEVJDRI3pYA80DpDn8dPl07vmCAQ7
S87Ma4r9IjoIdhlqXNp/LS1QlegnphwD8MVQCk6vc4tVNlUYxmDtfX1TyyCoF3nb
IZ/1cPG/k4xEAFoEGBhfMhONO3YBH1h5SpeAz+OE7lEICRCqkYVjMXtzQIwfpwXq
jx63PMT9A4r6nknQI3a8A/cmcgUUGqWA3XmG7uk2LnT671OqryhzQ/ptu7vmnAtQ
/1W+VYk+6FIvrulAw8dY/ckLdMdiz3UhJ5EMF0ZfXB86iqXAxjsKcDy7fqCtb3eG
giJkMJDKUZrWF+6CKZrVv/PxXXCs6zhVnwQmwkTfLbAb3aA6cZJpeMr6dN/rDHNe
aaKvatCjsOFgbRe6Aje4oKQHjF6SsPt8wvvCt41d6DJ0YfnjEHarevubBKXsLMuv
6x6JwPXstJXHlAxatxTDEQf1dy7HukCw/tF/VC2ug6hO6/NpDQDgDYtrCIkuuKhF
2586pROotY+boa57oEqTwoXtPSy3WxX4bfACTDlU96uCWZ4z72Ve+68e1ywBOMlM
WwddVAZOE6pA0IJHoiDeHMvsH6/1jDFEIzKPvXYX4+l0kqqjH/gLUkZ2fCo4LY4S
cEa+BGDsUl2srGORZyfpA0Nj1AHf0ZhEvsJ/7CZIW6hmPjJSt8KhGCVU3vIOF+4X
1X+6xu1vglwNc+fpi449gYIXlIeAP/b4w1pFlHs1julngTMF0gf0M7LSTQJLtEYK
oAhVloRDdetnp/ixjVn7yVtDTQo655kALNkl8vq8z0DZDj3zDWmzJNKZM9CKmTFG
siGnc3tehIaQc3sBioJ+P0RAgJLwXKG60dKPN9i5jogvIppYAvxfzS1IcGmdkGHJ
ll36brKULgSzEQqFsomKbaZ2WFY2UjMJox2Gstz+X4I/nPL1g6Llz6OxYo33wFlk
DORoWdblOsACQdlwuqcCQ6DmOVRt18GKuUWzHc5rax3q4eT2hWWebEyDw/Q5bIFX
/IgwVnntdA1wgiOl/KVKnK/zm1Pt6g09NsUDBxxKuRYq3wBicReSqV4KdCmO6al1
0WtSZqHOY17s0jtVzbq/kfShue97G8ABlwqPHBE+5PgwqntKApo8GDpMxENJasc9
ojn2r8osv5klnkTy3i3/qdTWl1Z+a4PHxFLAFpZJGFRffMJnYRxNfbnaL3kn7+Ko
+41dbToevx3AnLDcECeFwvlNx/c4zeZPGnmzicUKwEPFqK6P/WNcp5bhOFHLeXqz
3Oe7wdmglZX2/jNwzIuUR1rtmzXP33BQN2pY/bjuXFRNKuksYOKCLPvcnPtMgLbF
+mlIAY5v3IPvn7dH7GR+Iggy9LC66omvxxjWnV6BgEmPLQF8et4CKl25THXBjIwt
OCSChEy+xDTFwPMUuTZXMiOROIqVKUwzhoG/zrpPs3y2JrKRw0DT9s9lW3I1KEDZ
hJEBarMJqz8ezz4Cd/2qJthP4I7IkfjwFT18BfWybLgXTVESnwcREJ8rT6WJE+JK
1cB+K3dazRKePPh1UaV/GuHzqCkDjXQyvNwAc04c1wW8II5NUchJUROShIAezDmW
U7VpVeNskeo7djJaE5vBpQLBro5Up8VYG8PuTVYzxUuWgRcy8c6P9wSttFoFlqQN
US3jBiv9gxv/pD/HCRe+rS+IpuqJdBO9ylkAnkXPKO8rvyqYLnoalyEhQ7Oqp4YE
kgo7s6tPkmJE/ZWn8CEyvxpW4OaZSjeuU/EnmewFoYfophWorBNSAmDiCofM0GeE
ENfxqSLxTrrkBNO0d5yROfJSG5Jc15sk6rp2f2L1c//HoZ2pf+ze9b83swdPLwjf
422aFsXgrHSotj0NuSdTfLWlTqnoasWGq4tjkgrqa8+rMkp770IdIRR6BPgeeD2V
GDrd0ane/RXqr2vyDup+PsNqFsmVMBKfhFyisXugI+Elt0aQZNLzydMrKkPlFpFa
NFnyFc+uaL451S9XQVOJw6soMRF7ue3LqntXmsknAQvE1V9BQ9Y95FLnF5Heoa94
epxpRUCYqt1AUQaK2F1VnQOtYgv+Y0zOeIyhakMV7KdGEHA+FPedEvfrbz/mk9ke
hPqappb66ERl/uPDtD8K39lqSK7bIOr1YyiIfcyGQXcAC8syZaiMimkYQvK0ZuzL
qyrQg06DcitGq1eKc1eFhkpRRkKjJxwt/P1n2zwmEwRpOjkIR1YA4fIzMba+XqdI
lllx/v4nXsg+P6ClacgkG6hlgxUinafWCTqZVPxHVdDuuVbYl0Wt5rm9wklas0vj
r8OE2wD/9AWC890VWwU9c2p21TuFsFL0iLVYpJdfg1YUa/Eog4RWuS2BVVuFL7a5
Ytgs4mv9Y4zYdMyzfS9vlH8MtPngcD0OXUdpZDG0zTMCR8yX69YpvAAI/GCHmKPy
JVsWpjfRycrvhMYLAnTzwo0nSbABB74YJ9wwngn4AxC9XfuDL0MWhkmjk+3Ozsro
it9yLTANaE9GxbbYcgCRhzfEYQB3bu8fLEqAckcQ+eyhH/kVzMVF4lVcKY9WYpWu
QldYUR0kcKRIQw74ZIW0GTP/sCNseEoFUW8wOEzh1zbWbTMpnlWU4zZhPvXlb+IE
wwLabt4mimUclcQXty9HWbKRKTy5BGRT71YK8FMXyiF8geuqZ3F+mv0cbsD9rrnv
0fWNKs3LXGMgICrwfZ+YbaoAtK/TRS0VhoMrWgmjIRnDW9qF4rZrgBXyqWlIHbIJ
54fKndENrqJ7DY+lkHRcVzs3H6Kj8raNkoncs4mwOfzalYBtpCPAjw80lOCTCy4e
X2KPVu/0BD8d+EuOLctak1g23JktLPDEu5OMDXTG5+jzaymHllVkVxOApRUupyBJ
cELk3qYhlrVPHhJCEowJMlK7KEmGXig7xqrTlcV72DnBDjJiKuGOQR2eCNQvVh8k
tcLjheytF7+1OJwFhwJtMAthowtSyHB7AI9rVENQlS69m+ZAADmRvOGMH/JrX+cF
rRtGQfZdPH0rMuNpcBpiWJmClc5GrJZ0XhwCyr46STXKAVLuiOrYUCO7R1TZoCTq
HDn0LegK5gOmkPi/5K/NrlP2pgmv6VPUJIXKx7Pxd8rI+ReVPED3w4AW0MJttoPH
++CjoVDLwduiyRlKfttHZGfDn9W2nhtsFVBCHg4ZnvKf+KYF8McevNFkxF+CkDfR
s1DMaXCfdEz1KRbbs08QNAi4i1awUqvOe0lJnF1fTd/6+n2aKC6xE/5H23t5Xyde
L6pLf0qAhb3G/HG0dh/FGygAguFhX2BifL1p4qfhTntJWGP/HNjGww3ZgTgfCvJY
Wrph61fUZmBJbFQS2kNQyU9hp96JKg30mXkTEIhkN5Uiuf4w9yqo1c559NA9W1X4
NHt6e1D79CQMwCxpFeapn8GEq2WibTNlupmucap6uRRoGzI21Ysf2uz9gofRxpFI
BYAa+RV0nlCvKCY6uS99WVR/Bu80jusim67uLqPamMBv/irpfKGESINxc3moREIy
Ss1W4GDJNdCZ3DzcXquBRoo6MiAdpuKUsSJAC5pSfxP8Y1o2A87FN5kOWfxQuj3j
k6L2T2KShth08n/e/62gIo+Glr1mtV27vbAOmq4nTp0ek+uuA680GtYAEYddk9TO
Mz209Av5lvdxtFela9RO+05pdINL6Je16Kl+r3NTvSiULnHnC5faa04m5YpU7CTo
VyFrqkW7xUe8hO8+S942bkDAQuSeCAQ6v8N+5O6VDjLpOu6mYaL/86MpJiZBzphz
yC6ZTHRiY7f1J9fsJvsqqnA9zFJIN32A69hfTqwxzD2JbgHIxoBp0TLJB4vbfX7r
j7lz85uPOV5IBkjEvpDjnrVYl/V9bmtAGn2pPbmDVRZt1RDzQtPgEdSId31GVq8J
82rwdxZk70UK8hIrY5xJ7hftAWmbgZ7NNpkPxAbtuX3q4IrmXFydiUNALRrc/6MA
OJLpn/7hC4rKWdIJnl2I0dlg/8LPhGwew7JQda+9YHOpRj2cXZMzhZxNEFSQFeyo
HxUx+ew0+EpuYzX5enpjFlw9pbavqiGvz+Hn7PSxPneGcE7ETJCkrfTNQfbh54gT
dy5TBgvhkIU4b/neW643mfWEhsEewDHqKZSVHFjQW70TVuR/ehgJCA0yRmxHSkUz
EoZ/wceaZ6Nbsore0Wvy0GnQOwTv0MAA7jzH3ZzsC4PS8IOXfyB0VMNHnZeUvT4U
KX6H3bB8+Bu360JIt76JmAT8v/opFSKmjBaxn3g9Dq3hoFXwhNGwRsk1TMeNOfBY
3TP24SnbIza4Vs2oNn19mm41pEJLFIUxzemyj+1EpzsWe9nXiNaPac3kJ4aTBCxd
qDIP0f5XLilVko3X7pEPJ7W7mIbG4jJxQXY49l7YrQwVD4RYt+dRmuJINmrEOwXX
b6TfjZ841MojJhSs5Yn+Tebev1MijSu+68P4VFbWEsWLmRksSU22VcJJ8owG3YWG
VmuVXHVp+cKZZCbr+AVJCcRMF4iawRbXS/w2JTNFLCAggHVI5T8/u9JSnJkb9w64
Uj7SAvRAg8CVSYVdD/4D+NzqEzgfdeoXaFQD+pcDHUg2tpCnIJebfOD1lFQvE89h
hFwiGgzLvxESYKOQ+J8j0DhHRDmqC2Pw69N52hnh7jCSgWHho6cJ4tVAxnxgNoPl
Mg2knPO46XYRArX3oCNVE46VrtvF6rBfnCdhV0xLqbS5O4K+BiHXVYlYC+KSwc3G
ynJghC2SM1Rd1s3mnGSR69KmiNOjzsNaEmhUDg68wU36GvSymTUJgq76NVyWXSSN
DZCjfhpAN4/g2RfckYzt0AlTrZLaY180Q3PUq5iCVNWJFBp0niGiM4ht42a7fH3u
7aoqZy2BLkWp002Xw1RX+4+VuTwFcQF91OLoz7fnRoTpXmutrOb8OJYBAcQTeM2a
z/YXWBHR+xTiyEUx6AFHPrys7p9CnBUVUKWvFJNUydYHhG77iPgsXDrJbyBzVAkM
mmbqY0EC2PsKn1oWonSRJ0kzz3uGJryEKXxclQFkNOl+Iql7uGxAY7uHBX0mq4w4
qjJ+lVq22mZ7DpfNYp7zOb+y52ubWTst2x3VXJun0wC7nPtiUPdnMBTOgZg9c9Kc
aRDhV12+2wKG7XEVjmsfYMeHHLbbWGwsJMErelVvO1OiIVZysYN59WRN2abL/RQz
oFhEztMf0jbLCtkTsPYRBAzU1CqeuztH+pkG/5vObyi5H+H4jCUE9WvQfTRA4Phv
fGHLPXpNz6NkwgdvxrhZNwSTipO7uWITFeQwBFw1zHZ6eLYIeDv7YkxFFeILz9Pt
o+vsrkVLfbADnI8SMmZqBocusi/Or/FJTwrC9zHnC3KSn7rEj/NmKu6yM5GUa1+x
W1523rUXmboNSPclgxCgOxcKFI9U+9jRQL0WlTHbA40iIW5zLHJ5kAe3xPbAUVsN
PY+rLJUy206dBeMiEplckxfcMHsHga3cW+D82HLmp3p+ISjgmoxEsISpF+loqN1K
rCfTcZMrjBnMTuWPwF3epQ1jGVhPIWHTMLN+XJOrXbMo42xMWw+8xZy2fQ7lTkZ7
HIGqf5FxvI/5FUjaLG5nznkpC2VRmWtjdSYTPPjqWTv75QzMzzpsKxJCrOfAsgry
5RISv6cuEcmoL/RRpvcHrpHYLwmjCGBznZbahpbYe8zmW7CUbfdJz7MmlJllHbmX
rtmFBQco9uKMBO0DgpGSFPrfaTcKFq7+a5yy0vuUn8oP8DotZwsg8Il0Y+78yqYc
87RSsudIW6IQAKD13CLwLNemq/7UXwGTzvAM9ihqkoF4irUc2kC1huox4vGDyX24
LanDFGPRNcIPEHPxd/+/eISQf31odqtQoKiD4jcbihnchZcOE800LVJoGnL0vDwf
fExdrlNQ6/58gxb6iaQomn+H9TXYDzKDfAuKx4uDpu6t+uNezNe3CyeLG2zcVlVy
3PWdEPYZg6MMxfzAvabWJSfcYP1IJCKOKHrFsCJ1JjvxppgpUsVGuhvxCua0vroa
dFKFbjwx7BM5znR4gzT6XENBMs3gqgcSWABKMpnQJqFam/S+q7TZSxKNaK9vnDZA
l0p1blhF5LW1LnEvrZwXLZ5nBp3810fqd6Ekc/5800nt06J/IRbzeAmbUTSTq8AH
LQFxcfVqpGVjvmIPlZdp76YMknQcv7ED01IVZ9eeIyV+PvilDLvotE2m4OQF/Lpj
ReLZoEsBfIBQ7HeODoee6u21WBPNJDhPsshYiiPx0rf5pOxG5HoznNR5oaorYTUy
iqTyUOvM0o7SAZY5n4dkMud0aDDMXqC2BK4vLFPbYmuf5AyA/qsFZsCu+rzaIfej
o0vY60n5BrNLTh4jNeJyHOsTxdzAldn4JyYZm2TOBKv/oKNg/0aXk0xaXp14iE7a
Wndosg3C4YGvLJQjW9bBcj9S9p7z1WTC3fK3bK+/jEUDTVy6FFxy0Iht3hWxQL5s
wZG8mr3n3lWtsdNXlJGIeKulCImblUAViVTg0HejNW3eysM5Pww2aN78Xs7t9rdm
+w5gzTL9+ReyV6XtaNUJDcbtAXSdYe8Q3zJIQ9Lfg3wniRbhf+EVhGLCWedSypwb
hoVVKTDGF4fPiiP7W1QDbx0mGT2dj3cEYEtA2Zcbjlgf7/TCS8Q1Xn7ui5XXx17o
USmsrKEw9Q6EZMU1fFK+VUnFwuEaC5VdseOG+xT5EcOwtt177DG9tZ63Ur1lXRac
PUvwWA+k0KFGXrJRBeDJaRd0IHGxzUmh9F24YkojfXIMVJ+MJSy0A4HFsb2UmeQE
B6BGGAWpRB+iSv6aGJJv55uLDeX6XWfLJnucyvB32mVdJxATAUIuNGAXO6JkLlAT
eIvSn3uOMuoJ9Ufzg9lD0SLrH/rBwvXVfmbIko5oN2KeZ8NztYlFwTFa1uUh5zVg
XjIchRRX/mvfJrQg5SQNt38WWO9cf4/CnCviQgIaNQoZ05FR1l8yey0okFKcobea
EvGqWWCrYnKKJK9n0C4dVWqBpB7+GJx2stvnM6+HqIu02qWvH2qDdfiCKT762Dij
QvoJG21p84foutd13uSAY8A+aHxFDRI7z1bQtdnelJ+aZn+vrZYP38bugV4nMbHb
A27epdz91UGMnViba3HgPMxR+0P+TRyYBo/6FzqJ4Uh3F0GMe9ieTor5PNh8Gp0r
Ef4OiHot7yCn/HK3E8mVr7bFJ8X7r9Lgk+K6Hepmeu8hUATIgqwXJ51by6QT/DS+
TPt/2okLCljE2h839zazhzFNXnXSA1lS19BSAj65/RzfGQgw4EXJ6RGEG1GeBl6+
6vTFPDPVY5wMsb2XQODLOqzHjhjQJx/QMNU5AWohttPrX/GcY7GGXoILj1U9HxmR
zMEknXQ0ANnxMiCk1vb0BNw4NarDIlg59OUurqUxcNF/WuQ0buqguhQnpdkJsZ85
/24iq7eKdeyOg1KiOXHH3FJ9hOZcRwx7ePapVbny9XPRLhYSmyCQlNbnRu52HgSG
2Qq+SFoLoOLBij0Qj4Q+vMuvET5x/65opxS59WxfvfIiF6hghnbYN1vEwj/xEUyD
0GIEsI7qNz8grFsz4qYLRcR0WndVQIM9PU8Fa+E4XPK+45QTcUhf4HupOiTtJhKw
2SY8sfuScLkO+J7vUSg2/S28ST6ApVJk9bZFXp3uoqT8mcc9lMoGAHc846/zfKt9
h8qJaW74+vuaveDkjGEdkZTvCb69xZoFrQ4T5husGI05X21fhizvscsznO9mw70g
jn14jGncFTNgh1svdNwtN5KQa9Ct8P2zRX3qVaU1YPUXCcwFiA3DR2//y+f37gIv
Xb+Z5sYR95f9KF+2sNBa6zZIpAXI0b0Y+/FugykCiTFGN3Xkg5xgotqzRq5piRJa
NKcU6qys+g96HuRUL3j5fIGyEiYxtQLkCQ0s5LzwLKNWKczZPInNaZ5xVN0wSAhb
yRg0Hd4LUDvwZ2blLQaY6SfDCSki/YKaXF5+YgswHGiEZ2ZO11bEtEHpJhRkywVw
1ZcCJ/UjCkKlFq2/z4rlKW91lf2e5K+9eVBU2bCTzuFr4dQ0b4iExSJXIp9YDaQY
3gQn23YHkKoYGRabDEhb39BfC7JPf6A9iCbini3x3flujO+sTzTlU9r0/emxoQ/0
oHkq3ggBteAtX8VawUtgYd2tuFtSY60/y8YxFg20NSXYhq4xXacv1qVTik2RBD9C
lpRSg1VNsyU75TeuZVU6AqaFxhNzKTECivHz+1UKMZEusj4+YYiw3Ss8yDxjeoUJ
BDW9MTxE1hpqEVaXfKIMGFJwIQA/em92/KwO0VrtosuU+oNwhIFvaJU/SQ8U+j1+
hNyEt6bPtTqnUv1ALk1RW/w1IRYfIFv7Epkf1t8NhvIKoNOLZ2IV44YVtltiAb3r
1QszJkrQT6l+05mObQ5nc/c39KLUritEd5lq8v5XyQ0bg2O4+cLHIW3DnmQq2k4C
EIdmO6hrJoq/88X8xORsFvbA39NVuXYv4RqsKtweadaNpsszl6r5EvE1jmSYu42z
S7cRdi7Bjl3DF0AcE5CvZlfr/Qc05+7gKJ7I1VQt5RPOpiIicMcRVCcuwXZ7NxXu
PraFCeBeotxhlUwTQB7CZ75K/9mlDGXw3K6khMSADIM12Fi5ikKC5hs8XKARRsFp
/5lrCRVHEo11pHRsZgvdFPDwrj2MGsp7rUiEYp88uuwMLUjdA+auIGaK4sGe6Vth
hYiPaAyHwcmbcsPWEe1jI/EncFiGvofQyS7i5IWjJg3lR+qmz7HkkAFJAd/1gtG4
Ih/APx/nu59IP/FTVrh95Uery8MIW/pRYm35FJCHo/nc4fNE69azuWgTNz/jIAcx
BhE0GWn4/VRHI5mU1lGCKZldtLq995qZDe76Bi+s8qI1kQ694fyHy7X9zSs+b7dV
xHs59l3hBd7buoMAbLs1vd9e783+DfU3BzoH45f1gGDIawLuhpjFavOoz89OkJWA
dv7EatoV83aSaFogVuyA58PAUt78UVn6zsJQr+3urguZb8PByOaYfvMFlzLuBxQz
YJGMoQLvYsSsxjPpcbikNj6AQlZbyRdd4qo89ka2XtwP5Q9/dXaq53BWpV5g/mrP
MIgE5JR9CvhOd2252VBfI6wOvCPThuCvwE8dzn3H5Fqpbo7tOmXAWjil/KtbLBhE
AROgfVuI+tyk/Tw22kD1gdChIr39gvkRr3ZLRyxR36UbqWY3VOQ+/o3qWG2DVgNu
uBvwVpTP0oSGD1uxhKzX3ebh0lv2Rmp80bYkXcB0/Gn3izUa8SAY6eiPOhuMLF2/
7G5gkN8ls2tXn2X1ymQdoSDwy1azp4uAXskkaohs8y4swdYPlAV5eX3RDqHOJ9v7
cHoQQ5Cr/6MMcxk/zeueGqhV4I1CwP523lpunDDWbqCx93wO2yUvB1hBgZlx00zc
lCQ3pFO2VMQNyCB6shEziaArbbbt56gouEUDuX41pl3WGaXY173+CCYupOxMVv8c
MmpE/R3jPlPN0HOyd7rEIY8b/Uc0nX6CN1Y6tm/1FoNOUHXlHD1aTz02UEoa/ENh
CTaEcdx+OjIAhnxFpcuVNEtFMphcVvQEtObbCEnNUyyheVAupWoCvAB2ieNClfii
IIDO0WgMW0PTgvqn1/osdKYl0LuZygY9k5XcpdJcDMqQBrWoIhex/AWQUhpUbzYc
SmNmVsjV5XXlzH1Kb55iPKmBkIULq2/5EeHzi529AU4UBuNEZqj9g9XCdvMgOLn0
Zj+cHZqU/tTLXmm86NiPMMm2xSk0yRbMfVXfm1zcZ19s/pQZEErCWFeYXpkvWflF
XlNpFM6YVBxwKFFul5p9KOCUmeUkcElf2QpYsEIpUiVirJlxtp3JWLb01so8uECQ
IUVyy4cPrTJG2BjGuBCUNz0P1A5vjUqUWjK8xsmfZay32wdM9Cbe9285wSKOXZx8
+x1FiCzct4+53DyzXbje9dALIaXjx+G3mdO0qi3KlP42PVPgftM7ReoL+QQEwP/7
o9f/BJWL+rJXpZoZMMmSQHcJ9r57tFlJ1SSKuZZMWDT56IgZo0SLxYaK4qXkgQVb
6PMPUFxtOeuNw2ikec7OZXcw9XvyehTlitOXbkkMRv4jbil70U8pHIsw6ZuE6p+J
ILb3N7KggxCh9nGHf73qc2y7IfRstoVUXJcqjg+xgbR7P7l2dl9ijILonbC6VR8A
FvOQhPsIToZ473AWB6JHJquuhHpt/ynTbrL6Z5OlIyQXo5x3jsbTmhKqp/BzdyyD
Bg2X7LT8/wnDWTehTIvrdO5JopzIXLCZacpYrIQhaEHBloVh8DKZPO86x9QAaJ3r
MDwOvgDsmLGkenWY7QegonT1TqxCjOG9N/Cijrk3lZHRLm6gSjzGUBran92PAL6+
MnsrWP5/x+zi6qYmA38z+aPRVBkvh0H47338JhrK1aNi0ROMDndE5IugzeKSZzTF
rR6nLbN22EQ+4eWqsAs0bxHBaFBgXKfsDhF0tuhXKtvgLDmMboZR4Uk5O4qiI7hb
Xg3QGlwbn2y6jX8D7YVwapNDG6fQphxFbboF4YhqYMpY7tsvvGfNnDotFIofmWlw
mZMZ32s0+3mCmF/AyFglyvzV8wlDX/OBaPgAzkgQ1hwpCbEprbMJKu8tSUqly2+3
/03V02NrG5rP9Wv7noanISjeGMao2xgLfoj+8QZ4LkdKkHFQcrTMLYf+ArmHs2bE
VMOQ1JbnrPhAZTVznKls0mv+yYCB37Nc3QQKGyI/T3E24ZhX+fQHHng5hZuJk/Du
Ca0XYMO3FK/OXwr/ogFcoUmtGAZU1dvkLlUK9BXjrL4cl4ry+q8tHVfvhZemX56J
o1LtdpjhoNthHDZWCCYYqPTmwkZIozUY8uyjQGpAQblTMf037OHmVgVSgpaFKtYC
AkTi7obbja8nM1JHuF6sk6SfFXgvGYV9+a1Cmiog9npXcTzJEV+cIEfzLVyxZXN+
50A9iIrB5/QNti/lCtqopP+NCIAzQOYmjFNQ86bUvCExFYD/nCDW1wUDBXsH4Rho
5el135t9jZwSCcnsufCTrtRMkyZ0PUTq8ixSg/uOvczHdmOOD4esdGsmb+bUpdE5
PVczDg1ITyqGrghDzFtAe9dptTPy+j/OFLgjiflPGe3E5wav55s/AcT8cXED5Tlw
s/0HSIqxh8CjfUGoc+2xZlQqVLN0lVsvfS1S6anptS4wPOif6UB6WpXwXv9Fhjhh
EcHfGDeM9NlxczDrL4faLst7V91Gbs4Y/i8HfGTzFTCKpgOA6UZWa52Off+HcOyC
1cJNIhVY0nrB56kr7DlA/+lCmM9z/UBLrZS7Gz7d/3WxFBZuuANGPxSYcyyIq/9S
TlXNKRCYjL22lKwtGrneus3Pi+Xf8ldVe88xEMpFirKTyGsBpx2gvFePiLVni2qZ
HZiUKIH+gAK9ARYa4h3Vcg1OTV967IRDUn1V8OeRfa5aAP5usXY9Hgjbsg2W7Wr2
MwHmXeemelvyaxeOdMWbPUNIQ1iYxBUDTXi+r9cMDFe0Fu5549aVNjo+6L/4VQaT
+pBMJcpzbTQcxJ+sYqaiVopv56zVANHv6YY/PDtyxyDl/GlU8rjT1svuCClaBHVi
zM333RLNRSeGZXmM4mUNrSOyhsOmcnjHSeGIpKQo32SWjrNlXxiYQccfvIHKQG+7
uaMN1g1NoOJKN5gnjvFwuF3jW4KmJN+DQt9uvR9tdOKnFMNve0MVonnY7tRipmq7
yvVDfqrtgl4hs18VXwHD/4zaWEDpjVU0TgwR6MB3L0j8hzqEU8NLv5Vpe9IyUEmP
w7QcQkAKSj483ZbODRwO76JVaPhRjZs4ZRl+vZfhEsuRzhw4GATYLvlZIiGabpGe
xocMphtOlFml3kwMWqWgCiwL3x3OhN+4/zj2aZLGaNWFI0x9DFZkhAqDNipYjm7x
CydnmBCcSDGorrpgpq5GZa/irm4yehSje51d4IKPy31xvJXrkerXaNXB4vkpykF6
S0Wz7DwjKeX1OuprxosCdwUjJOAfG2RHIvXStqoMYCRU1IcsfDFGcxnPyRfLIcQb
Z14/3I9fnToDAayzPA/Al6zlzfkaESfBj/2w7XdFRcLK0iOonIj17R0szKrG8XYi
+5ebTYXemdo1rV3IMVht2UmZTpyfaFF38j1knZfHLa1DDKcFYJO+TRq6IHkVMeqw
oaO7wRxn9ovHVOzmwY57MKTaX/P4Ib6TRI9fUNA4Af3SaqXABNeBtYAALUHLTX4k
rEdCdqbZ3VB2TRNzDg9jGFBRDIExt9R2o1zZIdoiGv8HxJYMXTQFcWstLjv7XgPz
sXu8f3WSd0G8yr58ZIxkm8U1EVYz9MsKbmT2qPgxccpA7zJ3ru3EbsewnG3X7Qqv
dBYKAtBIJIoBKBr2ao5c5vIgbFCwXgxoeeTUUwLRwhXOTs+hEWbTQmKZ6c82R4C/
xC+S+DHN9wYSzbqVUTStDvy0yoXgpzZSI5iqJ0WFXApOjSnDe7x8+hqTPvePwAaa
VXVGsLmJJsOCv/fY/7isRm0sBKuqWgdJHydJH392A9lXoO91xBh++n6XsFpmbUsg
BF+ipDlN+JygJVK3KbpB0q2U7LFLI1h/rccFVU/LX7DNRp7Bgu0wByWo7P/0Q/Oy
g/JiwzXUBmhr8Bi+WINrYDXXE0A7kcWpgeRRYSRjpsKui9pkqQJQ4gQdzuyIYYKj
n/3PJA/e0cLUEy8Y4xDB+Z3J9/cKGkcxfcDCf6uZtdJAkvtL6W8ou9hu4NuxuADP
E3SbA8g5XCgAif4m20VagGM8HtvGFOFi4L1IBQBrcQBCbOM4vOec0K0MtlbInmxL
n4/pnBaXHKUSX9KgHR08sGT9cWmL5woucCnL1iozQrofW8BtlMKNRV/Y6/H3ATdl
hyN0eyyWZ86GnewkEPN/dEOvrYorEOqKyXsA9nxQw+RGrUP1hiKmuVPx4orsFArS
ECDW5ShcNXKH0jsRdnIZczOmR7Cic41qRRgvcm6HtZoU5EKuJ6aWLBN6SPEhIP9D
RPbCGAHWjkEtEKaWjbtiWSXKDt5yfHHyN4mtd3DKKWdrg0TLZXHeQQHAgkbbzBTe
1DEdtVmGIpsmosFWftml3bHsHN4yf4mW94rjH6Jh1lYQrAbxKmjeuvIj5eQ/N/+W
P4rnJ6lrIIRFyq7e/YzMkHiPmp72sNbMBOyh8NT8l8TKpBY7PxPW/RH65xNBeVfo
eCrbWHwptTH2m+GlNCL9a+KflAY+S88XovOp5a3wOoEClYNEzeAhTRh8OYQUFbQQ
7I8Gu+UDiLYB1xF7WATk98ERQq/tGENOb22aSzCQkbz/huRlgkMmIKRzQoslrt+t
lLHvH93/my3+8qL5wSdPQr/BY5CJUzKOh4Rf/r+cTWM55vCNCbe2CKZfuiyrkrzg
/lIRaCOI+67dbEtD0CzXzxJyKdetAVYn+VaMjX2vKk3cS7k/IwMLflkGQe1UAYD9
U4ThJ3mHhnFqLuj/+syU1+M3ACHCM42kWbDUmwOYGA15TDwQ7RYpXcIGalcdnW5v
oVAiSx0obma4tdy7pALaHWN8amXurCKxFTpU8D4J9zMBH+6XrzBjAYTB/oIm2F2J
KfzYmHgyouEYRSGyeDQDvJ9daF6FiyQJD/7jgX0Iwsjr8UKscDJoQ6CIquDxojVg
Ijo/fkR5h3/+SQ/7ZanfYwcTF/xDSftd6WJBZYe2tKvY/yV6CEdEf0dRuU8pZm1O
lykZJMpxhnc6Ngb4pVE9WvZqwT8zI/MkxGMH0XhslnPTEDFeqoDjF1XBkoiYHy+X
VQmXTyL+J4PSYJeLjw2cKt3zi9SZRA1wzbVnlgNAUgOeevODcDgXVrP4Y7HWiBQX
/p0/eqiDP5nhuunKh6RzGikVJcbgY9vENwWXrbqrLyvUq2vWvFI53YdgDQBREuGd
7JHe1h6IrDmiFR6QeQF8vYzZQChTltXP9+aWDjvglJOBQ42Aw6UnYAPeJmtBALpK
wz9DTBn2t8jK/zs54T8ZQ6rf42cNV5QbPu+YXDTy4vXoE4OYiWhewP7Wdx9iV/q0
8PRjNsMQmP3xaoWLUckAjrO2tpw0CY7s/rgtLXNA6vtIEb5PCfnFbfeZwaAY+GyG
66TcFcZ4d0w9AC3Yjxz9OPftfAJ3s0ihn6JzB4mtSBnc2FgNjBCUdMVes09mZr3q
sUuJNm0wNPSEUEzek3XU3rhZEWjCiHo19Ibbho4LvNbLRMa1admW1L4DgNwFi5K3
LixAOpL2Sj9US/u+hF7XigV3FwXSrDraKo4nLCIlm0NydJmU2hQxCZdmxWNcRTnN
RtfbKc0ZOHGpSFtbIssFDhvYa6xPfSRxShzH0dxOx1QjpUa2IsoqI3R9cMfl+WJj
sDlJbwYBVVFm46WHMqiczDnLlwxNmRzV0X8RIZqj5OYRuPKil7q6aWTciSs5cH2K
1V/k+AWntkgThxfIvKvwOXWTaebuL8TNmT643aHTHrNU2NmxdudRMl0BHwt9wU84
7z2FLURrB68Q9q3yxiWHQrG+YlStWE8alrWzHjSKVTUElXvwgjvfYvSbA7InFCc5
Ocli5xJQValnIkIoNwg18f5iy3GaaUYZnk7JkL0LXIZI45Xlm8kKazQZ/5SehErt
SYEBTrGUTaKju37mvqqP0lZphPJGqsLz6AdjkD6Dm3jfiSCKrmJFQyYeNOZlolFp
gOW79Zq+Gp1iUs1HEc0RjrJiO8vqtxRZkDD1WqJ2UaalU+G56ZzX8sOSDkmOlZ60
OjEjSSIAmsXgkSUCyg4JHMocafNlLzL0EO1WBMyJTOkFHX3JWTjsqbcgKNnPqOej
Qil4I+Sxyw/jxCoNhNIEcxHmww3Gcuumcv3rrV6VgL9j6Ur2BVB+w8OQPjDvpbiz
l/1nOVASjROnVe8fvfD8bsKeMn3YgzACI8VsrTse4EZCRynb5Zes9vBLRURl4gHA
3mkZ0IGFIdigL9Du3iv2IyFaH0eN3EdnQvomT20D8qG17TpZJ0QVoZzt8zp/oQaz
W9iY1ApWdZGhSwdESybZGaAJwZ9pgi9CPX/HfX+cWlI037OR1CPk39b5ThS1ty9P
318fHkARiGd8AXR3HRWKnvb2bWiq24dqtGfibyhTE0/vlaZ7/R+aGHjEKKCBNZS7
qX1Ndc0kT17z4oig6Zh7Hs8ZuvLbiZszD2nJQ6REnv5uIgjo1O78b5M2eLDy7nby
zmnA6ZqSg3tdXNcI/yLAgVMpX0sEoTyNOM4KeQ+CqhvgPnKD9Ee1Ykh9X2L8uXG8
hrzl1Z+Zcl88nqjplvpqrKwRX4/YboLKLOoK3OHIsG+NGF0jOTzA8Peasc0a63AC
6Rz23hCTg0v5bjMUPK1yHQJ8gdDPB/to9a+3L97wlvJkU0W9k8u06gMHnjMSzyrI
7FnnaWS3E6NFz/W1NoBBHOnLyIHG4nmSaIbDZTxJZAQjJYTDRIQabc4dBNxg+vnW
ZHpkdcPttJSckrh8J5k5i9hqWlvZsHwQrQj1HbR4ZvcHWzoN1N93Wwhh4zLs5MfS
ADz6Ip7yYpKypE7veF2mEX8aOjd1eSDEFZnjzbQbpBLj1VBMDj7XWhevKO4lAS2+
pEVNsHrnpCKcRvZmNuuO6MpEmrGyVDUy/Dz0EQkpTyLnaf8TacTBQHN5JTXgm0jI
aYZqwRusJOm04auzE3yjdF8q/2z4U1piYOhIspFxhkzDzsaXBphSSO4AtUNLQ25H
pHi6vb/0yR/gGC/rnywt2Lr8DiP3jNp4NvhccJmMudTlnzUKG2EoLLNkQS477ddR
W3YlfZGI41RGna5rifTbi8Ft8kjmg+v/Ga7luNCV2CmdiIi/5v98kseeScyUrELL
z1coTG41CUUHtxRg+5+8DenkThmWCnl4ftDPE9xIfKsxdmGlXSbfV1EqO7x23gqZ
EqCSeurCproFM/vc3FnD7Pg9x+g5Wxv/Gql1bBx8Q+okX8VIF7O9qFRW3niAOBb+
anrkWG1hYifKZ//v+zvRP2PhCWdbzpzsdzUN1JnnGw5G78fYjcSdSqcGSOvM4WKy
CyJV4P8obcaHnzlYUrNdv4icb7zApjG3sYQQHeKmgM6PAX5avefI4veYFPsivqSl
Qfdhla7gzHSrJ49XQsN8f+nm9OGeDOqn6gK/7vwPnJq2W6bihAIeqMXW/zJGR782
MUzIkX9dyKyRFCvg/DylgfCVUczkG4zR/orSNheioxMcCFlo0FhiXfxg5fyBfE2x
sYm+UUnkgArVgWcME8AAJQPJvMDoxLLGrqz+hqBevR/DRlTlKcwsq1YhZDmBP+dx
iAV1SJ2RRNVX532MNRaWt8PFAGVej0e4+PuSEH5sxaqaapAyTdqW5TOEcGgSuHKP
fSAmizvl69h02+pfs/3Mp6A8EvsWLl5aD8lrgoguTyH3YtojRILAzR6OJ+7OF1fj
PcngcbsVTUpjLbXbhBspGPJSd0zgdYtXCoAOiBf6oky5zgHTkRieGXJPz/tnw02U
JRVWMbdbHqwU8hLzBvmVAzvbecAgUWToifBvpn9lwrYvr65QWw+5RnRdrKhi4M/T
2YKSsOzSAKG3GdtyiVX7rWGuK1A5cjO4rMh2fu+7s+QA8/sFXc6fbeWR8/N6jZRe
MVOCirpXRTmjFAbAzvUKmbmWNqjnbayTuWsValH+diZDzLIgguPJB3gt2vukU09R
cXy2kMTcDdpTQFQ2e27EqLwvemhisK2dc+ZEvap+qs3CXR0rt7c6H6SWW7+Op1g9
pHGZgsg1ijTls+Gi7CT8KksCwc3/SRqAGrBscJY7+9kIsxhoe30fTTxw+A6MkQ0m
eKgZCufjNeQ5QIOfPvmPsVdZDHVodbS7EkkmeBpoXPbbn7c3gIp12+fMrVGGVYCo
lBMQD6p/0GYyqg0JkuyH7dUE7lyNiyOnuWMwJzCkRigu0VllgBofHNov5QTkFDAi
V84zDqrUTQsRPFtLH6dURz7zU8Nr7p/e1QyTHsfKhgrQ/xH8qbVkF83st9Wrpq05
fB3AME1m5J5i4b3L1sLhdMUcbbygElm9Z1+aTDAWM9SWdIF7Xv+L4bF25xyhUTkP
8rHv5wUu7TD+zxALf1ILdaBUrX2ZS8O5+7b5/msd2ozTtWjCUmr9iqhAF9dEgnsL
mgX5SDSKgVV9aKbL9uMfBHOtbUWf+PFsAgZ3H+hwI9vACt243Uo4FVLgOqOo2Bt6
FUN8JPl1vIYAH0iohDiT7t56/tSR3JP8f+yDttOP2ejoQawODJYrA0FSs7V6iKtF
NMklTemrhnKwWaEe9D7NcVaBRIO7LNqT/kMI01FzOLVT/Tak853jwe8orNPIACwJ
SL/c6MBDjU1hq9BEOWvbba28FRvVhck4i0+dWiwVz8hmwbyW/ukXMMLlZ2NH8Rzn
E7BYHu4oX+yLrtiXONzsUPvau4tD92EliEE4Rfi01/K2o0tkxFw9Z6fM70BOJTal
F/EDFLn5nJxiRsD2Zj6I3GtgsOO9FHa9MJRXU5GBg9/Ko9dufaz0uVRRr2Fja3d9
L7Y7JNCJYPDNtoNHK6OlwfF1JNLfUALLrhx6dH4Pwu3YCY8GsYZzxToWRsaeYAqr
16hyT7ScxAu7uqivjmjALKWjyam2Xa9Ezd/xL/cypJNwGY15YUf1w0bzjhI+WsrT
KCs8gzn7TtmFdyzD1RTXJvYtH8Bwm9ohQ8n7KiVZz9NzXQAtdQuKVy4w+2D+x8TN
k5ocwNHunmKyhCM4JfdJl4xvGW1cxV0rHwgKJEMhoDJBVaMcHKXp0eJceN4eYfCf
fW/0Nb+Ds2YAgI1MivX6t7vPwjlA/n9W8tjFaeKwGVhttPyRMvNNI2qI2ql1WfR2
doZ97DKod32taltDr/y3CFAHZgLNOrQc3HMzI0ZCSQq/oN84bGkREgBjzSglYcar
ZIReQ2l4MvD4xxVUL6UowF1qOLZBs0wgD7zXlcnaim+ap9vm121b8R2uCX6hD56n
gy4Gd0HgWW2pPKsIgoe+VgLW4nlSKRKLJQJISx69rS886fyouTcRkL4tQySbFGtQ
IgreX9mwrN7NfOBhpcXh6TCxheZduTUivpXhote7VJC6Gk20NsObrDdsh6QyawUp
nwLMPNGT0PT38R4JukkxwVNTxoSVJeGCGmQsQv1S62sna5oDrWcMT654N7Ie1rSf
YLL5o/e8sFuMHVovhUkMDFRxt3vOO/LHAm9yrVYcLpHOl2ESDo+Ynn3SDDCMseWU
3jf1Fa8rrpbDPDByZLvUdf1Bb73E7pg2XZLqwIVfXX9KIwjoJvc02s7HbPaLmxJp
N8nEIEiYX10rrd38s0eAHSNl/IOp32DuoppDPzuLnGY8DMFKIQBM3qJjeyMS97aJ
Wq+V+SWyGWlhdo8XrzVepJJ6FkPK/fjxxMJBDHFjwp2ivPifKjtVbZPq7xkodWFi
M1vMGu/agXVsPa/YdcqRajF8kpluoQQVsFeu/s/xHEyD+2nzoac/QfOz0CDpXdjC
oVatgvI5hCjvPvfLZOSxJeg3FLEkSCakVN00zU5dWevsYcvAeJ/Z33aCbLBeVhJO
XxCgk/wTL18Vs7vQ2g6y9I08chMzojmXt5gFfIcUhyRPdgtUB9CaYdaUW2jpkNzi
eiCrhqQ1ZHX2VE4FQ73BCHfW0TgGDHiMw8eNDtple/uw/biY4GlUjAzVQmAJj9aM
ECRqOnUAvN0J7HFZyxPpWZP+3uf3GEU3lTQ7zLa2SCyMT8Tw7Erc8hiQlbaIE7co
Rsf2qsKKjHK1Y9IeYGtynZezVtAWges/AQZVSUsnLu0k5SBupiq9Ohc8HCJUgyPE
ubjDn5lx/qXGJ6wVGl01vl5zMmTLrik2Z65kQSQd4soC0PlC+fKCO7FjtSuo2jZ1
ATWYp0YqpfvWgqYXvbn8Iph1b7/vCXUp/j7BbFHzn2KurBEjMmro8pSEhbnmmfF7
YRKRqXdGHVSURGuuyjpwbFAD4P+JZUbjxhWyUTKl9quMujjqgc4PJwTeVSXY73mT
eD+WtJLMZMUpcujIv+ECMaLoOaAe/1o1Ybnx277mJJM/OY8CIR15iQUldTRiUIgp
qWG5HMyYHYn/MxEBLBZ3FLkhyeIGP3iVNwRyfg9ajYeCwpje21Y4UsCts1wKzlaT
eNCXmPL3gDWv+GhV3sjQlwweABA4MHcxhd2rbWWysZgUCbxdOPTLHM5jENzkJiip
SP8d0Dll+gEecauoJDL8CaCGOWNRtsidlPL33ehArHUOCAWb70sJyJ95oxoba6Ql
+e1Ha9AhXQam6h/d04MikbXnnkOexShPfRon5qNops7hd6JuZ4nkxUq2Tnw4yvo3
XRO5zHinf29G5i2B7DQSpgagrQ2+EZiDf1UcH9GzBy/nscAGxRLCzSzovjes6Twh
iMgjNs759zuMC9jOz3DfRVsVVPg8mPxQANrJNjLQdvZXEqHnLHR4mLX/zt3wm1f6
HRyqnr6J+K3/tR/sHwpKJh4a8vWwChz5hKOYm5mEay9r16NHU499MfnJaRNiZyOT
mD28+AnzISWNh4YjIKlY3m1zaxaBikpHwpviCbH4/sk3/nUyc6Izajjkh/Dlbsw/
y0KnPFgkB+MHvsN1WO9OpMP/pkDbbYRt2IdABP3P5RSwediNGyz8FR8g/dlUAN+a
H6q4ddjo+2tuRG7naTelo5opXPuT5Hnvh2QikWB/6yCEyBuQ4Y76QC3dhreug5ha
FzmxqITD36f0sJWU1Kto6ORBpBLvtfGQk3B2d3lwQLsFYRy5a/Pjacecypk/CTUn
zVOfJWSRkqcvxfviQ6zvUXGw6Vtbn8nerwm3MViozcfq8YeQpaMOZq9XOf7hXy73
lZ8adhcgS3zEYStCJM/lOqF7ajVwGa9KjQKZmtsg/ag1EjMvrwuo8BweRYkOEYAU
fhGc3+g3qVwallKsTsIM7YhPtLvwV2pIj0R80dgSKKWGFSWF0bilN1kraABLsbou
P01EvftBcr9y7v1tbbYzoQlmNSipXo9oZcZWdBOOhKDly6VC0iODIxABtGs2Il/9
O+NxI7znKd8eLzwlCu6imUN8RS3qo04rTAJ82jboOTog6jk+NwQfMEyMF1VMXJ5q
BzYJ3E27zkATtjaEl/ZaZrvR92yIZZErO0QPHjPcKlEOk5C/RppBZ+WmSpkaCnIg
Db70d70g+4CXeaNMpnnA/qIYhvXpsF8zExi1b4r6ixxQHv0TY6hn6rdS/N50/3bA
4IVQd3KanAHeXyko7OjNysMo3tMDShWa0cDhHeAsEBYAl339rrQ6+DF+89q0f3A4
nXOAW8YPPcBQPqEIvbjAlb38mtoSsPgc7gBTyZjsebuktSR1WyYlLlL6IRWFZpW0
SbiGnIqv5GqpYKpfuTGveGSyoM/aK2qmiwX32OKpVXInm4tI9t+Hj1HW7rY849jl
pAPamjZJIGaYOA1XZwPIgXNf+Q2TIhpY76DALFFbvfwDaISJqG1oWGEbP5PCnepo
t7GlXVkT+cbBfW7q5RC/dsEOGrEadsW8EZ+TycjvVIG4XVvifv9MB0+/T/xUkTpb
7v5R+azfx5OJj2tRODLhvZBbqcPeqo4pWl97tTIl3u+0fjGkqexhs52L0QDwNnAL
iqjIYsdG/SAHpVG/+TVvHHl/N3KUOd9aewJ1A9X7C3Knrv1LbMpKCB6fiSGGOWR/
X9DoL7fEglPmQULAOvdSEfkWmSeCR18aF4bqwXJi7W6XAPHGrudQL3rHbGY9z/D8
hsvbzmfdIzow+HnaQKnu3leD9PSMA5sw3l+7jgkgJA1aNdPq1wQrJr36yEN8UMk6
4SeidblxKPqHjufR/b0KMte58AAQl/+lCkfbV4k7xTjJFNXjNEoT/NvEaMuYQ76o
8lyGhBy2b5wB6WQcDXwbET7j/ysHs/aoaVcCvI6h21WvffWNmMrlYVwtT5nw9TUn
og2AL53q7hPjfTnVXxxJIeHr8EwA9YeZUfjmhVQA5tvgrtXDwoTUnnm1QL6HX9lj
dvwk9PbihFhyZ58/r62v5Mc8Z4z3AvZVPkEdMG7mrbmO7XVeVZUBmFg4chdjrHdt
T+jBgDscTFuLglqR3Ei9s4ksbKT/JOhqu0X08wJJeKkC/os+5Hmw0k5nIyph+Jmj
gdeBqmZn3MGcGoB0S/yOgPZzs2Pk2GX6pEllb7t5rB8PRm9uCodpIXlZ3Rhuo9FS
jGjfJkVIXB+O4v1KA9Jg4LHXCRpPcOlYHp7B0oIvFPrST3wYvs5DXUYx3HEB1XRh
8+aERxVVnHKeSJW6kFrvPNpTcYiuAK8QGSRNApJrWUHDmlv4eyYjLJOukFeKYwWg
cdlHrZrp/47pOoz5/AbER2IUx3zeRL33q+NQHjLnQgppZX2JwzDTNk9swtzljDgZ
qORup9BAzdrYVtRIe0ktEeBnZ32iI8p2a6kXQeGWrbB9tvMtoPdedeIEuDNJuXmn
2gfhjeS+FLx32Ta0xjAbIGBrvNxiZTrdpJOLwEB50CgepC9x31e70kkfs7hRsgK8
SXnJ1dCssaG6ftohrH9KWZgyzWiSseNL2zn+Ay4rKtNtG7w7V7oU+/5UAdDqzIlG
GDstRqGse+ZtZGzxk56jL/Vp6NDs2l/qyMXGikXcnWJRz11frk9wbQa9kqSXKPle
0C8SkLc2mv4GUVNa/DKykx3HcJTpvPpHCHixHJY19ylOK4mioBAKfkOfCIYMyacL
hKtDNstkCam2uWpflb8ZfNFiAtrHMU+P4boesIdU6AQ4DP7uB/8Op34JtoX1FsRW
uDg8txwGwZH59nnTbSXWr+w7DDDJKv/5aT8heenBS/ZomL033dNTDWS+RjZeStdI
TgyA8y5OAKwCjaXwmYrkyW3rghodeN/CJ+EVLy+CGfqirCf63DP+QqAYgqbbtVDJ
J2gRFWxbEwVIwaMMxJlEpQzHoEIuSkZNm42sR4MvuIHOPEirNAUuYdRxR239ynP1
uauvD7B+2F2LT50oUurjp6euTGQwkhC0SCwSwEMlzabvpNGLyblMQXe6gETZH1L5
qsI4e2wzbpB53tBhnedRSDDuw/rV9hgS9eQZmxFOYFVjdayTIbrnnHLnSOhJyTxd
2CVlF3SspJHrw2JUqDMaym/v5GOV5KN8c42eE70jJej36dw9wjKJ5a/IN0UCeT9e
cDl6krPN3KMCP9Joa82x6oLa6+xGVGkbGE0eXlhK5UeLtdSdqTQ6owZZLBo+T3oZ
vaQ+NUh1FbvUSSVP3KqnUdbSkpmSQwJIPbSHhvmnV0FKXwcBga8LE/W3TUtNYkJZ
LGvUJpQX+771CmvQcvoZm3x9YQzlhp1RUWHyU193CCayOUrFwVEE5ubxpgRLXwe1
DRpZOTM4lslcJJQcjyZux8P+gfcy9sSQ1ZyEhn3rXfVwQ0jRpFWzgyuLpGnMfOEP
mf2PbmgxIbCd48Ej53cDQpuCQ3lxu2n6J/dB7Yr2/wywgSHJToVnKefoitBBVTkY
npEc12OuPNlRCtqtwj9gaQkZOaOIde6utor0IRxWmnWg0nxJvLAEQQTO+ktPwBxz
MX2PUh+0lxK5XIjL7lRV9/BKE8nzKrdlKUB+JGl6Y5vroWPe7ru1W/LC80A0PTE7
bdZI7qXsXB7qrOXENpZJVIagh7XtUmZeDqQGerdr0BhYYP4t2I/qzbO6KpCB4a+s
f32PLlRGvDhb+6H34UwInroIyhXTq4Uls9X+9UVi+nhuq3jOQtcCotlgha9MQ2i6
bKOQJ67qW0uxHRjqzG/UzchQNLtZsST5DMYz5bjoXt2zIeUb6p1TDIKdNQqWN/QP
CIHStDMbKu6L/idE6bACtLY66b7hFSMLOBd1uSRFsCLkh6WqlMdP0z6EHZ5zRfq4
k/Z/Ly4h69pbDA1XiXjt+8tS1DHcDkNILz3L4r+iltW03U4/nUoaWAXMytz9i1qd
cKXa8nMyKHx6A9sgsIzBQVC1LRmfOhGIAAOc5bQk5KEJvIhDsvE7CYxoh2uz2dQA
J5FGjqwEFnAw+dUyEd+JI0wNCTHaluWwNJ4iI9c86BShAc/I3HMi031p0IIlKL1E
fpXELZE21ABGdZm/k6PEkANTM/X8EvphqPUYRueaWUku3Q771Iwxq1qcvOCLg7SE
sSII/4vvaK2mJsTuhUESDvdUIM5CQOTW5zYYnqHYJw14OxWhma1eehY974IddBIe
OF2+EbYU6uVGnwrX3Dya0nwIach8qvz3aqJHHxb0cF9QCIacGNo50fBxSRfdH1Ht
Eu6VCDb2WqNY7+KLN6XskeXnvSMe4Nj1DCQc9uMPiwls6egjeUmCfPOQyO2bbhbo
qzscMC56PCQMu5UfNllGLT/85EBseeTMMHC3JJqsVXJIY7AthsET6VQMtIYs2Ocq
FTbhDNRIs+EVOg4IuM5ciC+ic8GFiB73+3nJceoPeRNkBk6pc9UZ7cGe7r7eT8mZ
090iFzFwH08jQGzE7OvEz8o94xo9+WldaaRD0eyt6hRLIBjS5eQNFUi7cOrA2Dou
TkaJ1Fe3rj8/rEN4JIBARFHG8epLMKI6mSDmYFJ4l3wyI50LvsbLu7rAapG59hZN
F76kOBkdDVX2y24aDWrzOM119GoiVyOpiGyK2+WsjKadybQoUJ/L7fHNKL8ftvTT
nsKOzirQAHC8IBCjWITdIm1mZ83w80KDSaAcNMk2oqi/GO1cN6lT47nJGDgVtMt/
ctrz0fjle3LJhBBT8bvNcsPFar+a7qK14bCqVmOPJes5sRMxoT9I/06EjtjZOOm1
gR2hbMR+TjiHaO23c0/bW8SYgDli0+MMxCDD97H4eLM/8f1K9gz+9K8Cxzc36Yov
lIAd83Ozp96CvV6bfD3j+OZX16sERL5w+G7WIYHg+LfHhM4WHJDbgI4FvPxxzB3s
EREkTMXlxE2rFH+jC9Qj/jOipyQEFkEAx2nN64oORSyK19pizjkAFM8NFJdMSxGP
eD3AdPjFXzWbZmw3aQcAlGV9JN6bvqEiHnkrZ3zW7hZLA1CGhIz9haLkhCg+3vqz
wI/jwY4oOn1MH78F3iPdSjqj9JPGtFo1GOc8KgsrNKJCiR9G/OYxabb8gc6O1ldH
My3hsxKovunjYS+9ImxD5BTcMwwlPwxB2jhwaXTLVoUDM+MErFtwFhZXQZXJrWNv
3zuo6s1gROzsGNynkQe3679MRUdJPTqn8A0TveBzh/5EmhMkRKRadk/r2RfGudVg
06hu3uAkLdfo8EcEoDu7ShBaVPKx8ZoXJMbNhjdXQGrrZ+2HTc+V86jfYYJzfMCq
q1JToHs4KhKRhWZ3DD8EezwB5hg3QyARiVVUAx3pVR6FNK5s+7SBqY8g8pmU1V0C
tYAkTs44PdRt93+zpS6wK3biLG7VmDOtt4u0wrTtAOemWQTQMJXH7YGm0AGj8b0F
MZ3xLytuH1NWiDh4rUWMsBacelLmQjgXOTme6X9MpmVJa7hNmLNshS3RsGD0H1Nj
DXXUfvzr31PR5BJHYWXE06tJCA7BCaOzwdfkZqLjyvbXu+jfFrr9yD8tIzQLa2SD
XbuxhMeekoWYm805zq8rBpoMqoQ7ImZmMAAb7sEBhvYiMlV9VXMDsgDxXTdfQ0l6
X62Stfzm2FR7da9Ur8Nr/7Ixf66PuuQ6AvCjGW97MC7p6CKGLnLLjd38LmWxoX1d
7erm6c0twmPHLjVJE3bxDP9LCIHJoA8grCYEJEYjAXSdkfw0sLBi6ofdzSynCOzk
5/30Osf1jC+Ha5ixpQmehR31XlCkyWdsobd0lLMrgsfoMQM0mn6c059eBpU01/Yr
tp4cTTc4OlAQI2V5l2RIkhG96JyzlvaRTrLB1go/fYxzo2VtwG2Fwa78zeRAqqFQ
ojFwbdjZrgFoqA68bS52De1M2ehl8C+/XZ7vxgQbd+xlAFQk6NGxPmWcV1tj9s7+
135CfzHiAoLGZ9NlCDNR6wxMKeqMPVu/FGs5RqeQKh7imWvDd6iuaWFAZYGvFNAr
pqJXYc9W+LWsLB1ciC2+zU8x8b11sgqFQqHhApi+ZZhzR3YSkNDEDxkQp+r2pqv6
PgxBTZPBjWERabjwmTHAC5suxHCBVYAiv/o6oHFRU4lgIUW1SkY4HP0esPBZX4Rk
mN+g6/VrPRE1obQ5xSSdsk3FcUqg3RPhuAq/rS/icPceMphZ/gLNrAf1ScCJO+i4
PzExhdSMFHb6hHhRa0I+y1O5PXZ3kTup4wdSoH7xa7srIHstKUg3ypAPdg/iHCUG
tMEDf4KYZQ/adA2YSZr2Sq/mLholcQG7OCwsbpve+9nWGDpg3/pRmFmGQ9vhG5vp
XCIjbUFmxr9IzLnPNXBBNEfTnGpiGmxAmeYz+EfvAhLFD9Ueiscad845A+E3M9NS
/uddCDUwjtOoUtJByJsfbPbdITAzh8gVGfJvMcePuHe40D0k/C5WXB8mvaKBINOM
FTZ50BWlNGDmQfeZi1l0pi0AHbVCm74sVAIaPlgeisXxVdDyBikaHUi0I/0hjTrM
UrI9nMMDETcalC0Y3SGg0H/DCOeTj9JVY1OmCp6ERhs/A+VWpDvHr9r5PokdvKQ+
WCzlve3Z7fUayFE/SzAfBTu+L6TjVmtK1BWX4jnGHb9XaQjy7HbW6XXNnTvuoTF5
c4GE7/LefUtqBLwVYyuzwdv5P6Mos01r8hx6HDVR7wHkPY/wsXCVRrtve4YdJMep
PTdGAvjHw8la4JDkm5xk0GX+giJG3CcffFTs0dTmfaMhh+e+71Kh9W1vA2Kk/FYT
5OQwB1ftOrxpH8Fp4NwxJRGQ1LqOP3sWVBNRqDHrY4DZ1+4TSf2tOIVmrk5iRD/G
k9Qx3ZFdconR30pk+soRnVODfeiC8PVonwZHbboKrcht0BrHjcuKwIgPXScfHyng
dN1XzXl8ktYPYbGUuiisjRJXX1SFICr6d7hWpXxxrSK47yGEG6Uxx4HEmgyH2ZWt
6oEdAB7d1XO7gTvETQQK83fE/pl3T8A1RhKQ5M81L5VpSjjuI8Ez/9xm0/wQpNJR
vooPlxnqZaGcEvHABVFtjEn3hpYuC7xDXuyP0a0Qj5/0NF4WtBYckOe7quwppztd
A7F/JY8JVIYb5Sla8EaL7doWL8WXIbCAIoKu+OEYvSjHC74TBF8C18Boi53he/0x
kSvngDgHzxdaofrzyCpU4Zk9XutAlwQWMrsUeFlNA7fvGlZMI0kKzx/NNK7UW33O
Mve6AKedCh4fu0WLKE0LbeCKixV+8kiZwEqBbpseyGBcKnrOX0DaA5Qi9luhZU3R
4BiNIul89IzbYn+hr3AbrCueGUwJdYXg8pk5PkcJnZE4teN4F2NffJRAbBu/EryN
vQMlosTr6kb9PpLkIdsEa/P7ayjhod9XqhpOv3x4qGBmIyBohhBMrfgILZAC84fk
sHBiSwXHns7K6mT2Th7Yr/Sh+kn5RgheSrvcvqOROx9UMCt6K8rbX0H+pYKgExM8
b4vCdqFCwwWihzh/J8UT2HWoVAOo9dgXjw3VxU+ax58I7mND+kvFFz26GXsZKvlx
LnvV8JHULRg7XV/1n2AdqPMhuqq6TZqEDfTni6UIFg5euNuwjpJg13xC7E48S7Uy
HXoy2IhU4vrfaQW6Qf66zNHCzgVyDsIfuh1z5+bgX1bSz0ghOet+/yiX0Fp7VfQO
9t0H9LlZI1HE0tmyxyJoup7RHd6eLygeULL1pQWMJKeOiWnx9VssaG+BNKyGfGFT
V38USk87qudslNRyfMtadnfM1VtmdvkFOdc+BphEdA4grxYdlEyDKZfsnlCl19Lf
kBYSDBlwIFKNXZ3iGwMeQw4MQlJR0gqKL5y7c+N5RQZeyDJlTvlWemI76PU81xyW
CfHY7PxjhivprzFsj7xqV2I+YK9KYmGtaf8G9wus5jlUUXpEmuS7Pr64CHe7/ksd
V4jjGVjHbPNP81UssGzUyY5BWL1Wp98Oy0e1oHNIAA/cOUjL0X0JjlNNeVVsljsj
wsnIg4OZioqSGzIb+BEI5W1PCS3Mpdvt1Q2bjr8oIheyqlbI2p2UL0yxNA4fV/HM
02U+3zR3Zk9Br5ulO0ryO4TxuBOJOEcUq0/lm7K+wko2gNJ1ETH/0UC86y0HtTdo
NBg1PX3DmMzoOMxQLGpsYOdl02qyNh2PM6e6aT19OZu8EFHFXD3uaUPP2i4W2xt+
i7KzsikhxaziDMeKQ3m61LOVWKV59mUvccgmvvwT81BJTtm7LDHxsGBtotRJKk9K
XyNa+ZPAF6Buxbv433rZUI7TNrtJ4hegA448BAopkyz/dA0qUEXevP99VwTPW3/r
lTAQ4eUI20mTSTfWa/FGhBBUGYOw8PmIjgAX1SCfQE5fGYbr7tXqiestCYyOGaGS
iKDdSEv9yEouTW++0+sh1rxkV9ar/0fE1uFeUjtBUeZ0uE75o+HX15Ia9cpXODRO
GYkdIkxatuwIuwF/QKoUS08tGdwhPzo4uXXznqRa2UuCKdr024d9lVldUxC0ig0Z
+peE6xfHpi/J+LHK8MbkzDINR+NUqvZ7m7tAXTvLjbTEvNEkAIBx/axavtj+ld5F
V+cEcOlLycUMy3hYllpqu3e8myFaIodyqALhwGbZaldLA6v4dhWUVwncdHrDiyQt
lBA3DIaktS1mxtSdBZNIUxYwEX2JUyqW0Nk9Ib8oj3hzx/VWpRVlBCh1PKbLr3Wo
UwIdoUBntGdG5pkBtV0VcoMQzCGnPR6MXLumlG0z1k2apJRAlD210Iu0jIEg2gnZ
POsv5aUU5Qnr1d+DlEOadQckbchfWLo9qO1uqOsFvNYxMC1zDsRYqJosiQgPMCIa
ANHIH3JdqPjf2zwsSXT427RmBYrhVoPPiykfQBOsRhUit6WifbXFooDj8LimxAic
k1EckjjnPcSOoWCV9ZrfzY7YaolAivaDk6qJt/80cyGkWSE2A5eLG+Xb+Ny48NST
W2wXefpQ6fwMv9YpuOEiqASzK94jqmkOIKMVB0+TLZNpOSSCBAUobxRtwHrRH7xZ
aalgLqslZZdREH3pU5bo9L5dVQa8kLTM97AGXGEFIUwYSO/rH25eHVZEzYHcm4pH
FmtQl47m3eAD7K3ABzUVERGNtKv977UJjmin7O84PiDyT7vzgAzmJbtLrNIITT9k
cF/GaPTSjEX51m2ZarH/s24Sprwuk6mG7wwZCg9uunwq8t9uFmD3Af+6ryEoAqZu
cPuH+q9cRtO+Qu9jDPmtvN3o/C3KYDfgKMAexqV0rasMYxPDSqOBOKD27I0SdtW8
yYZmIETyjb2jWktptSQoSwh1GswJ64BwWJFW/Is5GRTPk9cRTQL1YH9JGdyzU9qw
MtKe+GmpZbM1uzwnHSE0PNgrDZYaZpGpgnWj07MlHaIswTVn0zXe/bTA8cnhpgrg
4oD74i+eIWqT+DaeUqD00N0wwIB+zL4YgoDwvxUN8P/9qW0OrPgoJepXuujkeA9a
ajSRSG63ts3omBBuEskx1T0Q9OHbBhp3xAhSIsG3Hv+3tbN3gZz9ovM5FUkZ/ITH
UCEob+/r/ieo8qbWXmHXYQ9SZNILGreqqk0pCNA2WBnyjOs4b46oJBx4YQSetWjs
MjZ8rodyWFZW6kEboI1Xn7vjcGACmX3X4g88cAfdyadYDX5X52G5/1yhhhzDgkJl
e9ByV+uWkG+t74AF8661nc7Sm1qPAF1cEG4aCSohT6BgavQf9TLW1mO87ZRsQX5n
knsvM6EZql2U9L5rHI9Z6z1V4m7GC8OAsd+QLxlq+SDth9Wj8cW4GCvnXov7qpWa
NOoPC+cyEPkFk3/4DnxWwTyQyy64G7YIQYCuEMPOe44fpVHf4zoDB3bzNtCct3AV
Sr/PiubqwL2fRx87GjW2vvgbMWf77q06y4MS9DPKv9MaNgiSGB9tCEviuQ9em0uJ
N+8a8H5aAjur1nUcL7CJCFBO33A8mlWE99gYE5H+A7gHXhPXT12rnQ+QVqgcdtxm
bLb/cGsMgqZtP+Y9m4NzehFw1cWvN+cGiQbRNPy58CfDYOQeTlsNN7uaME96uAkG
fUESFHgODAFZphjVdAX4Zv7LNewCkqj2cZ4IduE1p5nHHBsWH0FvMxkl483IRCn+
9UMhNyT7SYz8jj3PsDlZZ3OCiOrb1wVKK1P45DlUL/8x+tm/5mc6FX0Gv3IZDkSs
3viNsgHg2yLC2wwgPAuJrcDBVIQAZm+mFHD3lUpqs1kW+zS++YMzwugdCfOftf16
tmJh3vg4BaLi1pV6JCg/Kx3WxBCzIAGl0MjTrw+g63VhmAZtMvAJMVQO0kesyqpE
aPrSA3YAZZez98km4AOaa0WwuDWhUjLbcaON+EHM8dV+MiHe2YBANB7WLmR7YQ/P
l3orhxhDPfTqS++9cfsj9LqYHdRjhwD3nsEMTtyuHBYJctQ9qTxNdxHv7Qx+oZFP
yJBZKlQNdocoh3d2PD5GxbSgED/d2/CCniaf5jiSm7QjjCtUXmf3dj+dmnj0TejN
Si7BJycDvSkSfbhT2nvSB1BF4E85q0tJlmo0ZsW6ARXTjwb3GG2PN1r95QmOjGDg
pDN8YA1M7kRTRqV0sfpgLur+nyN5457AbvHz/KZBz9m/KRlmuK/ikvF8uzXSKsqj
FPeAWyjHjYXv0zZHx84y2pPmAMjeeBzmQhoiZdQYbjloNSiEj3akvt3mThMoGpiR
BUmou72JeXfZ3kQgMYPacshHineqA/+B1rG2zHoJLCGtdh92zFmhz+Ht0i4WPE3p
Jl+5RXUy91xYlMrRvDLYMFZQWW7OeQ4kDgu/Vw4BlXL1hA0YdLVec5ueKaCsoHeK
zPsMutVkbCgn+lT8dXRbQ4o1thgq4pFwnhyuvGjejtGg/oG3Gbjcr40RkcaR3lRV
cmtaohQNH6iyqJthZ7QmHaRcoq6nje03gISa8vuG9fDkRSnnq1NCPw7hmV/K9x7T
CDqhBctQSxi3+JL6s2qCvefcnHqfrNnU9LNFxDhm0mwhMPHT0PCGNr1MZITCfcyu
V0dAqp0EaVDVl03m09cl9hMTBC5Lt3IFWJDqUnrZrD/n94vG7Ftv1qv5w78IVpEF
IMXhW5P+c295bhIU1aCYuewIj9Bat8gMRbNX9pAGvIU+3vuhWRXDeR1izJWLmHUY
/Fl445/MVCSNvkyH/qFAAJemlT0DImqXur81Geb5kdHW7YR9BvWxgl5pVAWwO0eg
8DCEtRZ5AdfDdiXh2e2fOdLL3Ed4rnbykPjyZTVBeM9wKnluM6VDat9RXZjYFI/W
ehfFbQMg/fmu3SvsRV1xA4JzaMqGcHLm0TYe0ZCzTSASAR8e6iN/4RsSVynpEGQa
on311+VG7auuDqVh1ltCsPs2S3AsZxUOFINzHIvYumPADXCo4iOyelDOpNMclinU
/T1eJ+8DgdHCa2K2vBdmeRZJwTFZHWqyTcUmCklWD37/KzbgbkiEJyBCNKlXOhXv
TEQCCNhe28zFNK6EaRuclnWf26RBtPwtgRHKJjMvREEGuc8fTAQ8khLLYs8z0Iz/
cs81tkiYqFKXNBaHKnbre8XZr0oZDQe0f4+lUxCOqCUMcOD2uZHiyXfMrhG3eWaC
Ne3gW5z0MV2CSC6Qf+be7QnxDhmiF5ZqckvqEQWOCfWsJYMFM5hiNF0HbLJJxT39
hcxzNxU23VYlNA2cFCVty+RY2IU+2yLW0AR0EAkoLViAt0M/Ac0TocPNuetKMrSi
jL3W0Y1jhybI2bjlx9vIMgl04rhXfrkruU9iLOSvCBNRX1F4Z4GluBdtJ/plNQD8
4SFrdZGL4w1KeEOXXCdSE6qpvAoH489zg4QcyvvXY39MqZpNMhdmdkI2h7Q25mIt
aW3FzHxUEupyFdCJTyUSJqJgU+kq2em2XeL3EnOeI2vcAKY/QwFalObOmCZXjDKM
k7WoqrJrg/FesBj7x6YJOK/L6Lk005W0SsUqN7fJ3CJMrrfIC+Si8tLPVVmYtBg4
G7TjIJlQRZJAmmqVW7l6sDTLFeJAMQc58vqvFxrLnSwld8WR8zKMryOaojtJKZtg
6jhYR2hMDHvUIqJ2Z1M4//Zc0sTwxL5QkkUCC8Km8Rxusk9LHObhpiYKsHLTAqA9
bZxtoX6wX2TbkqC9/UmxcAyW9lsZyf8TRkqlDztHk4lyre2tUywgBWQ75asLTToT
nVVz6FZeI9I+5iybxOJ/0/d3KyC+GNy/aXWJYvW/lIX3ZqVaNV7IviDZJL36+7j4
hRI9nWj+EAR6kBR3fjkZjDTwKhk1qkBDNhHG4TBYRWrps5PRC7vbI/Xkc2zPvO7b
JkBywIuMRRH2rsKFw6Bgf0yTprGZaPp0aWMNajcwFz0wPlRUyCsg9UkEVrTX92G5
v3rpOkH9RSjfRZ17NHLqVcH60uVNTOs/7MTtGR9hejhuxpIZyEIoAsTI1w6XEasV
zV4airEZlXS+WwT5+HQYzWEBOFYJrSuTFSCaY9V7PAU0c92QLQTqfzMBagA9+f6q
Vnj/Vu1MuqfFvzhsPhphAAwqPh83tbE11C5yVwAC3HImRUYEW6qNyJCYnba0X8da
RP4+l4CxwBg3gqAjAfsBRxD4rqxF27JulK9qszRaFy1CFErUXFY8axo3wH+JK2IN
GepeLWsG2Nx0Rheitg04AAlKtjcEVI5f6bwMeRGHWtlUbrxrKE6v7/MRdIcyPM8p
5pssXW90+aSqiR9AGnEUev3IIc54/n96VOHhew3atEIzLpfHoJRVQvRtIs60NlPc
g+U9phkaYhajVkd7fxRsil0pA+lM0EOASWT2WwOb4gN6NIwihX0/55JgEx6SPPnN
rkcHwl6H3tHdz4gnFZ9UQ3tLTf4IbQCl4jCSBYpD7zxjixQzT0lpiBlRIqMCNCk4
L6GPXbD5Z4IluGSC2RSkEE4htL3BVI9LDyZatbWldNJOTICfnLecKubEqdwn7Dsr
I8OXcMWgi2LmPa2f8Cn6SPHB3Bkkr0Ytbw68F45nRVlRJyyVK2akWEMPLwZUg7y5
xvgvFoLFIhCvt7f/NXNUgHIXw4HbuCLFzsf77rGXVLXzgurMy1uz+bMOvZWqMK9R
4D87njtXY5dxqmKTuUE4bfwhWvhEMAEDV1ldeSF4X7FLNbnia64J9JiUdhtDe9jq
CHmQK02NmzXMsGdbKQd/DfTyx1YUWHFKucIPgWlY8AvQBw3OX/OYk0SwHI7Crx33
u9u23OCfKyFT2MOFS5tOqGnedIEu3NQccaulgsRZatQv1lV4zZ4+TeTa6MlqO22x
Xrpk/ZgdzL6xhxUqEEOXhDFNWOQ4aqpuE5Zp/LQRHEpVV9udSKZqcWRjp/PITz0q
DXFwK/8aLm7JGkP9fiw3arpFb/G4WLmeKDO6xXS9Zh8CXwdk6Iv8bt72Ej56Ywus
JYCCMJgO6rIb3GabJANAVDu4K4buDhGTN4Py/EZ0u7FMg9xQlcJozwFWiBNFwl/7
vX8IefjmDyh38+JFpfXDACH3WsKf58gTGRnCo6lVM5OhdFide+0d5wS16MxYs10b
oO4YS90F7LcJclvxsmwHIfGVZVlc9cE8fPW0MIpebaJBys3PiCH6AaEfIR+dhN9A
2fOE63gzjUxcV62/Ugo5p3FzY7nJ9AmN2wlFDLy25NOXPxQ9OUn41zB4kkjRNCNx
9+MEKfZciGoYVCMxzzhyR50RDtG8sIEzolUD69AACaKs4WXDLro4PB2VSLudDsUc
mrf49wreNbtHI8zNBaC7p+jeD7qOk66osO9NhhvGIwGJj60gdzseNby44hK4l7L0
27ykWLAT4dqsEuWIGV89aqxgBk9nD6xB/eKsksbabrt0goY9blsw3D7JbUYevBnk
RpFrrQeuKnn7eBCp4tU3dmECit2L5wwR+G36o6BTUx4vToyAZKrvGrsdf1zcM7Ze
TLGtkf4uBunJ3JOhEdY2a3uEImzY1O7lYmPtMx7rmMbhUsqkdyG/yuXwbS8NoNVZ
sM3ya1gIsZYDsT7X8sUOAHz2HQgEqvYpo2AcmkRZQ9uiRbvOr0+ZrqLyoO3XbPtx
vfJXO6RhEyvBkgYnKx7BvCTxy2k7yWQSBO0X9LLAl062/XELensMLa5iBCHcShJ+
5lPTBRjXxAJHMDSOYrHKs4NOEXtlt8W9N7D00Xs9EPbbE/00TdqRnwpdL+C3g1ct
yNfCxsduL3Hv5WLYWsl5eBRQ00vaEukiY7FV9W2+NptyftxNuVaDZxDrKVlEs51G
4ogLma9K5lyWMgDjPDKN8fV5VpZoy7IF6j9bfzlFen0nzcsrVBMBV0I5JpdFkWvi
oZAPfOorSHwWrfxkcyGmP87ocF7GBu5sQpo1dY3HhrEUKsfg38FFS3bcpChrZyWo
oziaqWFG/+O8ieTgEqEHbtad+K0xe3D3mXBMX7q5/BttNTsOHF9siYw00rOknhy+
DRwkVjemDc6Pyxg9BnYpfFSy9fbHmWR37v2lPwtzKvBPg5uOhSL2AfGuRhv4IdhR
GdGT0hGv+/AyPP2f5UXI6rBVaBXln/2wkxd5uBfWjqUR7+Hxn05Il41Xa46fbwyB
aEUP+JwhLH/wXyIJwCRzfV/FCW/Z130dA06lvyoyQsufcWvNegWbC2lF7v0EVCBi
NY3GNjXmvSDONxbo7L0VuTcpbj2UzN6RuIiupLVE7XWnkNA0w7ZbzEXZN0I1axlk
E8gmQPUthfEWUuJaU+lIrGYA1BwVH0j/T5OvNPLVZFR6nhWBLZMyS/gY3ZQiVFtz
EnkIbXPtUIiMTwIZMON47NZQBtkG9G9B6I4Xzekp/8GANeFmvBa8Dcly9DQIOJs6
xIoLjtd9osgU2wkM32+323QWfPdhyGEyRpcgudD+Mya0uAML6uMBm8MvDB+OJSEd
ivnMfjiMyhBfTXaq0ei3yA4YDV6iFZKqsx3Gqe+EH3CETz+9cLfCqlSkQwITlM29
vfBbgM0OMy3kmzAXLuQuLnbwb0awB+u1DP7mDnJidKjHZ5sdgNIb6cuGXIOzvlN4
WfseEdq8nq+qsbyMVh5Yv9n6Is3xWRVR7WBFGa2AgFj48wX2ECpeqDyUv1KHo4RF
+cEBwOpumSpTTre29AeTuUNS8dKzevAuyJ/pCAFTt1rqcclw/3C6X3apawpkG+MT
ghS/3tDoUQFZ92CnXVvwlNEwspIEoLXL98uqqrltN4qdQ4zxvqgeey/ySLklW4yq
cBy300zNkIN60g0K9IDqNwjQIAi0xwIj77GSyQjYD81T5LakFnsaScOCzoQI+A1S
YdooaUm//unqki84pzzxotaif5E7xipGxQz3oljCT6MoVXDSeY5SlWXAjMxH4fxJ
3iOaR3Bkv1EbZpYcDk6E3z+kqUpVBeVmJgQqjNpyD8ypcaPokdY1waft9eiNzVxq
w8n6EshFlvIq6v1Gz0zNS9szPmgbCcfN52ttER9p+9Sl4aFjCGXK8Rh3l4J7yRYd
HjHK5hlbG1omJEXxz62Xx6GQQFcks93AqPey3Yn6p+NRwP3ugzQkB5aI2T1OZrVG
NSYxtCjmiUZ0mUDvmslyyKCVkAwNr3ZuSOLmG7yuHfVTB5Y+2FyF8uv4uAVFirnv
WGMvvhUmtuGYJSu38Ti4QxR09WeXGSGbVNkdZBQYgixRJvkhc6CUqxgHTFe2BAmA
LxlqkXytkDy3Cw5xLoJ98/GWFuC+WRAokxD7b8TcaZ4TEwGFHSRnYR04kP3IYLEc
boNPzI+fLYrSc4VgWgCLkOGddSx3Ihz+lvmYCisho160pGqlKXLbpk4XTn48iC/Y
uALPiSj2YwaLogxcNLiMCMnTh3Qcb6tIToW+Nqdo9AbI5cuitVeymQrDP0acCxot
LcWq3dJ/letglt7y8G1iwBOrpUYUlq+W+49NFxXFkg6yYKatj2EfeazkfKdJ8Upb
15b9SiSqCmF80q9Xv1SZ7zlTXkK/UfnNckmilw/Bfl0mz2P7+CRMfm2QUH4tuo7n
APvniU/hNYJ5ED8GJdfq4xlv4EKPF+lub6f8vDRnt7Mizu9h43TDNSpv3f5wZtAS
GdmJp3aTBrPm3dA0Owdn0Er/nDzWYVOX2EkO1WK/dh1+js0c5oEr5y9OMvyPq2rz
Ri8XMQ0h40CeuFIj1O30VCG6snt9X78PaJiBkDh4ZZWmuHLH9Ioxa6wFFJUZIbnq
06nwb7tAg7rp52D7LbXjwAZGsYToPez3qfSw/ioVLz8ki5gvyX6UHECoE7GcSc8C
4R7q8fKCD1ynEYBdJnW2m19h7Mm+zmklXuZNa8SVrIaxqZPoYqtTj6PlwifxRSLO
heBcxx8mEZWdgE+vYME04s5gTgURomeI1Lu6fpePOJH3OxuwTxSL3LsUbl+av5Zz
a5kdxZBdkxVy+wYv9A8+kzEZMVo8EWbM8uBNncNAY+Ljc9AepVrImXyQe4aCVrmr
SwF64O273E47vEV6GdB1wxB8OBpb2yfTiFwl4mGiSH3zJfLiX065PLV3rNc4Zp5S
i0gYs3H72QmJw8qdP3XYyHIg27nu3h04wG5r0nRjjSm1cXVLJj9Yixq0fWk57z0H
LrJQwUJjogO75m2L+hKdrux6/pO1Sdaou9ehTJ3BujMCWM2ALJcU1DKciJ6nunDC
hN1frMYqsvL8Uab/kTCCd6MM1x001D9Yc6OZoUswU+mHgN7BOtx9ITMpuqqzS/tD
sa8GVyr5KvzEbN0g+Fo6jHCVGZyAnR8c/f+CKFq6HLghgR0d6jwf69SSDgt8jFKu
aXV1527k3+rVhrskfzGIo9bH3kvkXYSybj93MmRV8NG2FORwcPq+LXbcc4ROymNk
BZU6lFBCa0YMec6xsNMgWf/Fpirx841YnTXq2fmTKuHby+5He2R2rGHCtWrsHr1h
546AXzFmdMzyO0gUvCXeVFDg/Yf/aO2O3zJcqxrsl42GUd6AsJ862tzhL2WMKGrX
GwPyteQm/+ri79VGzYRWEi6+03lz2ZLKQuAFfh5xHtEXo22w1AZohzhiyfWNCoUf
l4EkZcneM7mRRaZfUig7To//lFZf+CyB1WLbDRRFf2BiqYypoTMnhcLUVF5eETV2
lx/dZ9leBkXcMN6ky+2ograY960Z76y0R3KJ6j7ABDVIl4nYzcMlg/bg1uhbsovr
n1ePcIO+GS2JrDpUu11VoL+VQBVk0YkcaZcLy9KQtLkpS6bSh6itEHivsxt5w1RY
p3k06Cqyt5U8o+cP2doGfgdS7QAISn4EYKk/34J3oE/zrc66M6ZB64i/e6qkRJOw
wAQ499HQA7uW0y7vFNmwbndfZblel6b0IvPpls4KdpxeuD13dZjWQ7TjiP4bhkfi
PcMT3FUxY3NCBuBD6BxcbAy9CAImVJaJqB1UZ6833/Wd7nw1mCpEUV2MMsR+e7eF
34pKcs0D8/Vh0v9fDaev7kQdnlWJEdW0y5Q4ZAnbS0LtkngejG6RraCo5+JxDjVb
W1OcGW+bpwtNXsy4Q/Q7Y1ywKl65f3UF91IJBDq28Idkui8Wgqs64Jo9a3DM31SN
u55blo6hWms4mcWxioVKv1fjhVUNfjrmQDMpTMvTIEQ/QmwJdS9JLwt1+HVftQbU
JF7fxMoK3zyTSdLTMfSzjS7nvKx1XHQ4JfQDjIP2ZUDAxIz7buGsqHbyk3si+r1G
vj5eIas2tVmy1Cd0L2XPhcUbwVvyul+HAs8ZDS4pV9Ch0nchBLMusdgRnmAdNohz
fKE887kgNbvSAev46BQ0EnIoYOrZrLEOASdbedcQl14va0hWbkooxp6vc1igjLhr
Sfw5EGaL/pkndiVn/PgzZHEGG91Kp0tFs893iztcfNX09F6V4hIH9FLXk5+p/mEg
qWWGQWoen/5659mIsWo6AgFdip7g6ipnzU7Odlo8ykqs2tN3qNq4u88OXLTHHOCl
HuZdHSqwdCxd8/WYbTIBpcLRCGJq6GIMDCkx5s0XVC28d5Bn/MHDKqPRsdVI0lfj
iDoC1Pnus9z9nQ0ZFMaXRg5T9W3Z1IA4LGDMP5JtiCiPl6Yxz4KglWxFc6oxPxFd
A9wIjfSkA5ytHD8Dhg+BXp2/mTRdGIfiIZL+hG5mCZEsrS7z5yFVIvSF+EdRtTB5
1Dwd4znapDwBt3C8iTEG6cIZOosgs86hEDYhBSMCbz/WX4rHtXmbPcFS2ElkyiP5
6wrvpN83zq3NVw46r1lzfdUcChvhdaYxNJe1yaVGle4PZhFHSEFSOy4nIlKdfxCH
4s2l+PX+9rQ+UmdrXjDA8Ta6vTuR33f/2Aa6lfLPpFEl7wGDh4cQM8occc1x/MNN
aquYl1JGTEi0JQsDNUrFy0uA/2hGUsQrZ1frmyZh1d/MFktcvfDGQMc4XUHsPjhz
KuOOWBwxadLl/QbWc+/1Oy7s8ONPid1jPXBBBX24TrvPYIFodao6yMMT7UTN0T5H
eYMqYxSmDUmShQUnsT0bPMTGaelMlj7W8EpfX9jD1przeyfEY32p8VumOky2U+Qy
dpoBnMSKkp1dK1nm+Z5LF21rY4DUK2/+ZeSgw61kUmC7OGvoid6A3YxBRHMmWuQf
xvoTeMUCo+V52SkQ/aT5w9ks83JrE7iq2Xl0GzjolJmugRPCG7cIwUanJ9OOSrqS
/BZrI6zYgcu0VGqwzhWEJ+hLCpygErSEt5TeKflXY1S0vE071KJYQ0eauInVOIcZ
+UVdzMs8xed9THhcoeyOV6Sddm7b41E+je2CmKboo5DHFsXO9Q8AYmMzCqDeeL8N
O+iPwpeMsrsfBgrgXqHoDPc/R632JwhLMIS9BGbKnDEGLaMj09QgIYGr7Ll5fv7J
hXh4XOnbN0ahS35n6J//uUheZ5krk0Bb3SBHt0EE6ssqHlrOI/w3xVpAu8ltJwxd
amgC9ez1NpnL+ltWMFhDpxAK30TJL9iKZLLtUXNA6CDGgXMRAb4N88egEqyyfOck
Fj5o24ZcaGt4uaxDQtOCoTCbnJrDbxCiB+7htr5Sjg7GJhxuxo685CglZ0pCy4TO
1l7FHlbiY2BAPTPBqVZ9NOqHAF0i0IM3UnQvPSJ94wDBcDW9nXynfa/ezr371BIV
X1TBuvY52mTJPnSucD4pXSOpkwr46tYhk71TqoF7QZ3l8KQy1KPWMDV7d0Lcnno3
t2XIqxxgvUK0z3arJD7EwSmZJMG4jUO2cq5+/uVQeFX7WneY2hcdmJ2ciqqVwQhI
j+zfUSDFr3qcZ22eOoYhzcupIGdHMFJx0a49uFc/3z+nn1s8U/lqve2MerzDZZoi
jF7O0cHoBaiB57hQdK4dTq+KBw0pBYghSFeEEBG1LkwTN1Zf0eHvzBVdPosHU7Gy
lnpSyyVsjZZI8sv8lwmVGObs/UMHIK3E4PEd4dFyDxo0Bq2nEtQOkWUw06nAVaAf
zhH8H/569xz4yGlJyvRPqM9DVr1hIPbGha5BhM6pjCO/O/fhA7UXKUh3wWNbClcI
Z20FBeW/kDN+EJpvhXSkwqhG5Ylc2WVJ4dq31Afq6mx2tD/QsEfOr9sZ+6TMbRZ4
iDuBh2RE1C+A6CkHS13PXYmOijFGKBlH9aUG7cVLO0aCq74c56YMclFMMW37G5VQ
1RZVmj2DHTcxWgVXsg+8fHPUSQ2Umd799BSbyQef1AyiZIKqZDxxMas2LUmVJpcF
NyC83+RKCkId2owOYuPv5kNmSi8rQtBB4648nu5AUi4Q6RGN7ewkMtkPd1L0sAxB
txE97KhnSJH8cvV+FUVToAPy4R7Uw3p3XESwk6Sw1BPKbT7q3ffTYXKBK2aPwwJB
Ibg57GwCcgMIp5j6SH2IsX/AZIiwKCgBAWV9Di6WzgSOn/8fUuY3fsGbCPT2tGm0
eYRyIa2ySbEbjW/UBeIf7yYfVHRRE7kBxxKaF/Sb5yZ1WY4oNadWaKAcYhwqXWmB
iWLLjnKpNxXkfKqdMAb+gLh8TiaP8axRrYsu62yG7kgQb7KmXv5OJy+c82cJyvJe
FfV+3Oqx9hdVP2gdFWvXmkcCpOS4MsxirDZvjFEKzZsu+uKr87o5ybSc2LejwbC9
j6jbZfvFh/QNt/lrf5w4Tfba2KWVWRONGgOOJ9left4+srA4LeSAxZcS/IVdxmyp
m0VMmMaMkV2/TEG42/eIoPL39LhcNsZU9Zsx00seyWQ84awAsFnxMNeU3bUvvAbu
H/yMJ5OA5fg25M+ibugfr3Tb5O/F72mGYzV7UrCTvTWGP0zyDH7ozPaQA0GF8cTU
KOqiCS+u0GzzYxm4xB2LlLf5aAzSLywRxNx8Q/CN5xzpVRgyIWNSsjRlHngTz/eT
1GO923i30wYGGydDv2Sq80W5vzR6jw9aXFsqj8z6EaLjqxb+G7q7WaP/mu+uGzJZ
uhXxOw1yk1uHU+UEQ2fOGU78Z48Ugm9X8qqPyLBAXGatSlpgjew1ycOG0jHOZlOz
gqPoRyxeeXwmryanszydebRyilo9lGIeYzb729W7QwFB2q4/qDRPmxZlg1GxREBn
1dE2C8y43Ca7U16IGTjd/ayTRZ6bUSlK9pjL4heXY3SOWGBEp+FtkEWanLwqe6gu
B/05zekaSyhfQGaj9Lcspl4ie4Amw1/lnFB3PrrcfyXBs3n3EvZHPGPrB5o+5fIV
iup4I39sgkGIhrv6CQVGPKPl7nMOL7+Yeh7/ups71JYzDRQTj6NrVDiepF2ywWLs
fBsWbRFMFVBv6Szszkte7ome6r6na5zr7pP5EfF7LYMg9GPlTQ2jbsOaQY49d6nf
uq5j6qyB92lJ38GqLvnr3qMu6gbn05A7qrmWaeCOw+nnOLoCMfRrWNbNd7uFC604
2hR26bhwNP0O5wwOTIyO088FqtQOeq/9rFYF/Iw5T1TMeYDBzDeGy2NUvUSLOMj+
Y/fbEAWs5SqDdU6mT5CFj9VieikKbq6quve1CkA5ZqCW9FvmShKAxF23qk7TbqXr
76QcSJn98mN/oP6XhVjWGZZHHuuSUPMVXxF7r8IVHnFGaDv6nXCF4ZOuldAt9SGZ
JtcDyThqLu928oy5O7e8mgUjOsvTzXJCx5DEkv2Xvae3vmsDW8FZNphUCU/009ct
uc/6Durrvc92D+M+K+UXU+Vih/wOAjzeVe6k0fupwUt7E1Mo5Kar2IXI5mjwIDAM
CiasxatQIVvAGfovd8Z8sAdrahJQkK3zWMVF/RzCpdn3QDkIfVXHQGS9tlM2L8vb
vcoDstxog5xAIqJC3IN4G07JjTV43M19UK/td2/MVOqkg/YQYYWN3iWLVFyhzxfQ
8ovcsJVEY7pnbh44LLILB+K5+ticNwNobhUOvRKn4UzuFJK9R4b4l5fpzdTgLUuI
GC8x9bV3xgNCTnmfjIiXpjRMXtuidpnl34Gz1XYRUeRDJOVR35B46puc8Pj+aaB0
nCmNKBlwjLYO4e8OptMFIw/YVijve0VfkHjxIQUbx9QVFJg0EBsgEgH72+JrtcFx
8eNFNeX9m9DMTr31C/b5whhFA/T/3Cf20hopQMAV0avNDLooRX0RT4KubCRxrzAj
ey6i9+SO1P59KXiQmr2VttRtMw3P2gWQhUfkSLTtwaTLIBews65hntk4DOcOt8rB
exnoFO6uBxHJbEZZMU+iO/OTbqfkZ3DL8JUmDczE5uSMRWzY2MUSVxowR0T2xV/w
qp1cYUOo0th0AcRflp4o+yyGjEICY7lqZo9ZMC7DigGwa5K9oovNYXe947I/Qb0E
911qaFbzegY2CTxqVN5FSd7Qbh28s9uf/0wYvK+e9uEA3b9SDN5y+4vhcT9ZZBM6
enMpUnc1yToJYRkwDXM64+3SZiOuELWvRRo+Sr8PfPFPHZ/t4kesLi7Jol9yQ9zj
AtTXqDY6pNLifurexMhJF4gALnoB4XoUW9RNKh1YWAJln9ivgyEYcmOTz7MUs/Uk
mpZs8J3EaBjCGHxDRzJJt3UXexVa+9w/ejpHBjSh302xNT/5a2Aa/jtbQa96r/xH
umw5ZqJ+NnUu+yIGPB7N0fK13/Qcg+k6HA/Jn/df65eFJzOnDk8vvy8l+OBlezwX
7Qm1cQdF9AjW0GoLQPGc8FF7XisxK4yCHSrXfpE9IbO3pHxD6vVI0Ujh2BV967BG
rQ6LD3oPFtxstZWZ+Vujv07C6cjfD4/fraeKWoCA0rWhVsv2UENc+IBwAAaAUuB+
ggeMa26JyzesAIJB0ahLmKSikyBFPu9/sqcK1rf6pSFjUEH0CCAM4B/oEInUvg2b
iHvfU6rq+H5nSDPJ5HgCQsJwBoa2O/48Oj1MTjqIVh/zffHD0xsKAwPQDAi5nKNY
O3ssrlrbzlOWGk2QYSkHL9tjr6GD/Xg0RTAxCoePjxMkRGJwAv06WAJ7muIXrDlw
tOQlERjKS0wyp/8i7uvWDv7dUA1LVmVXqbhVHjjN3K364jRoffo/d2GrbCdg3lHN
gov9LuFWF9CddHt+tQJ9WPGVYGn5PayRaM5dGRK2p8+oSVg0WgHoOFgLaIE/cKxy
G5r1H2UmIoeTxEB6FdA5/bK6X/a8Z0F9gbg0yFy/CzcSzaH8Ze2NJfvvrxSBvBnW
EbrQzJhoaORRVQIeOvgUMgDE1pix4Hdb7pBVbhOWkpbyYV84vd3X8O+VHiXo8UMu
A+HWN/81ve2rq2XSW/QTHx++eEZIULRvOtjRe/U6BeLvrVLn6EdKcHpWLcnEQR4A
2xI01wnMvzGYO5zyZ3yfj+QD/k43faqDE35LT0vPOzuGwdw0Mzt/8leC++YhBdCT
6b7Cq74/n5T5Owyd5ymiR0pyNkIJE9Btsv7iDlm9bp9gLcd1lyLAXUpvC9ApIghp
wwWsYJtb9snE5KcprkIUX0a+ME0hiQD+jvSJfaZbSi3F8hbMxJUAgxhyQOEmkL4q
F8nzEFIroWoBKloRNrSdTFj7D9WBIb3wSdpthGJUowUi+ExdtqW190/RGEptNv6l
B0CPZIiu2tXaWWlf5f6JaEfkfH6zdV3kFtabYHUqCsY/Knxpi4RRDd8nP0iTb2DM
yr9BjZvmYPibfq792uBWHUJkQUi2IJyYTFc8Fgx6QB4I3A51ElrbMJotHcTFE82V
4NrW4uDRpcq/L+fF5OagYct2AbzXRu5UedeTfqOfsENC+h69aou8QKNeG990odFs
zJo7C5ya9XoZx7zI7gXP6+1Kz/tw7/g1m8LpLi8+T9K6F5+xZ777Rg1UdSQ5FGU9
nzV8e2XqEPQrIajm4XFLqsvKZImlgKtZDQSas/SZhF3Vb0HgwDCJ4Yd26jTr4GvG
mE8SeHBFc/1Tr58ux918sbnDav31ko1atNCnxEKCkfwEaXvTuNXZYPBZSx7jNVzt
1pS5+ayyl6JrzVUgcQ592bKU46/PNffwnywVBGlVb9ybEDKNmCpWhB6I7pq+ssUU
UOpWk7u8TNT/s+RrCaG8yEj1CyVuvttciKXUScR0exxdn8vDdp/gzNM7bis0e8a6
doTMzFYkYMhgUMP+KXjeJktD4e2803X6kqrcTowe3WbYvJRgu037CX9/4QyDojKz
QIRoJfnrR8tk0eI88N4nh83MfXEtNuvpQsfoNaDtXq+M1lRAZNMlW2kT8ElFkY+x
yh9JhCAAD4TJ2r6Sv/LUcP8dEPsh395/IAEyBCq+k1dJI3yjR/O3Y+xe/seo8hQl
BeGgYTMHtQlfHGchBaIPMF8/sV19dVfxceBL43ZR8pglIBUVJoZY6GPUDbv/GunO
xIKAuNp1yeh0qz3+8xeTiwsfGdWxG4288YHFKMu69khn3oUTSPe9A/R+aF5FpyWB
KOvioCzE8v8H0i0crI1GSE7KoWFPI7coe/9yRWa/jBZ0fjmYsTLLKwTfpFl7rzzQ
oiuxpaqHw53hn9ydMn2iIBUIDSsv1FMq+G5SWunTge1p4Ni3ObxlFgxrQ59HmKLJ
xqtWkVS0TKMjjbITOXgi2SNgN2EaUVqIeafe1+WEMBcd76EjSnDu1aSmoZ7O2PkD
pY99l1yFnjGLgVN6n/sSYWIf/2Ox9lIs/P29Ysjmr3BWWaYUJek05lWDoz0x6P8a
lhgVXNyZCJUZLQotSiKHJblZanplgrIuX2lMLw/5k82StATVEPyq6BIc5BUSvUtd
8FfMLS25ht+DGtkFSmKUkcr5H/bMWRV7T44ZVkYWKpvirXSYti3ll9neADgaRaPm
naWCq8pyXMacXIitrk3R/Sk+huvo4BBWt3wBKIJQtjmyHcaJsa7GGXAxIhPEqVGV
jpxRiSeGcVqqQ385XrWP1B5fVn4kL58HMXWqa0dpijaE6jrXYnz9LqygUwQNg+U/
Wdurk20MbXnyRUmuvY8e7Yc2hHqrpNV1B/PCcLUMcN3Mhs835LkecAq0jKXpJ5Qp
vxH8xk4j+ELcFgnqV6HaqtTFn/fCQEP1LBZVv9WOmzmtE8B3kvlPjs5v8mCiKumy
80ItTj+yEVHOsjmjh3DA3WVWpJ1ESxkUz96L+vh38EocEaGAxnIVYEIcLDmzqZzR
hZHBtYJxjeu/6HNHPPBNQewq3HsEeDhvdqHLw1oVf6+9tIfXc429QYyB9NIzsKFH
lEa+MxAAyFKo1WlHDaCCVSyBfvMxWhzJNtHbYk+YjydLpNbrggTJMo8HlXYB2K0E
YOyjSoaG9CVcSLnVMWPbSfkh94iENrHaE0GrrD59VrMUIphAJHyOED1c2ITTcr8d
cTwin6AyPQ20Q4QzS1gUSC609yzfwLPJkvJvhFwBcOvfN1wG2/hbBH4l+yxUU6qv
RoreQPT2ggjwja8azrjNZLfKpKVkXda0kKHe3KY4wCkARIe4t1pazcRSV+RTXaRw
KZ5MqpqTxNyhUPsBZWNAWUVUpptRsh287A+RwkzcOtSCzF8TwiiGXOVLpTg/92rb
g9u8iXuKbq9RJwMUAsA5GS7bxQi82D+140xwX+bKFwXag5c+W6Aai3mRkIn+6yXT
tgpczQMzCGmeNN5s8CnS7FhRxhx9i5QhAlaOGNAgpTirQUAz6ntjbvYHIYoEJbOx
JRKJhlcyj0jhytqfcQ/EtcK3R+U5ZRTRXoFUjE9TEtVIyqBnSPWAdjYFkxOzpPnW
elmFJKP953cdqvDPaakXIaeC8GLMzya9t4ch479HmZ0iPHnwFPndhtyuHYhlpw42
dCyh9GZvAdNsjUHyzPLhcYbDFYWkPZZipkQeaZddy7wWQSw7I1SZfb5hf8Gbjk71
STU4+VCEf8vulpH1qDFRCAEFxkBz2xkJo1igDvY8eEUPAUpakEoi0MRHYhoLrM07
kmUnp5IzN4I1Z2KGb0ht0S5tPCvpuDDIo5No18NaQwfD1XwdYHUDtN97CRlDjA9c
ZRMzc/zXikDLKpEv158CbROOoIZqaTHSW221BTpS3P4CUR90vPsQ+uQp3Ufnyj/J
ruv7wqTnBjZ/TqDKF8k8qMEIy6/0p2+A+vUWy96TEV+dFjgsihwGnfwJzM282ip/
OW0ATPy0DtuVEoZOXhoAIBb6+a94irrhM8V2BQ1oJRL+74xSCmWjyBfst2iSWf7G
GDRyAa+GrESLolFx+iad/0PyPByyYGdwOyM7uJzjJ5bQjYIkdvBf9ibuEGR5RmoK
cl2Ed5zwGliHNFNnd4iVmBJi8urLOZUqgQEjJB9X+bNuw5zQ653Wq3OOT1uV6LPK
g2QF5JS+DgJBY5LNCdvQli814kAfCIulc7vJKHKcOCG3Ew5LhJqznmxPtazXJaHJ
KjnLij3WTo82/H1v5sBXKV8/Ns1aLiGMVsBAjMyX+9ZSJsRqKsJPOyUMppz9OWnb
aEsF4AAhn5RwOOQEfLLAu3oTnfjdTpGvFSdrYLHB58fIPc/o1CWVBsyc2PVZtd/q
PaPOD3DiCqMXegWRGbRbKBK4tibkIBCI5fo1ps+K9CPpro0S+hZakKappS6kDtUA
/46OpsEuFe0Hpvrzy6dA5MsWRN7sIJo4cTc9CBtrkAZSQ073AqCWjhOQc99tP9Nk
cbmOe9XKTjjnamX0k6+IuxOKjGUHi/UT2YExr0kQAU+hdHYxDb4OPKKBbqd5HwBY
bFhJvA+5e4y4CktA9GpqpF2F/4Rp1LHIw4Fmyp2wQSH7A2ZFlOK4EZCEuP1xmdCd
Yikozl04IFON28/2awNBY7pujHwZgqTsuajSEriJAg2l13HM9EKM9t7+L4LRCEgt
G5JAV5lVwi9hsQumdTjvk7l2pmfn0iTgPvxhdtlG7T5tGq+qhD2cEpZ0dNmYBKZe
VG0Idc1nyWMMHeqFmnfjjnA2vvBMQujjSLCvhppxvSdIpMJrDfBS1kA43HbvPG/E
GzSU2rzWKH0+KV8ArGJXi1TsU1DU9+gjej656jHNN5hbnD7WYQQviNJ0ZAcI5tZC
NSFSiSDgUtqANCwUJ2yPIj6h1dC3sAH8P9Sk8SE87QycUdVCAQYWZvfgW1xbDuEG
YTOnbUP2/4PylA/UlSyO7eOnUJ3r923xymUgc2BefAHkKz8XcLdZHoTuUbAxhQVD
AmS1uLTRKUSFNmsn38Tw0A851655+1vSWfpIeju21M1c2T8dvP7aZE/vxpwfdec0
Mficq/JE/bXxR8WOWHDUbHmGcorga1+AEbxyhUfUIHCdX8vlGV0Q9gqWJeaQKJm+
efUKUOOxORazO6qD9zIocylYOCEP4oneiTcUFd4KqYCv8j7FdLX4yN5qWZgGf6k4
RUavsOk0mqDytv63Fo5TMqhQjxBnAWy/dGJnJAKaCW3OUYGGhWG8lkdSJufHIHYk
Nr7ahWWiCHT+s46iHeoCHJk0VHdGGTJ4Uhrjy3PZvvhSdwRwQEQuLy8Xwk4A+ivW
Wa0lE/g0llUpRQSDLFRRcgfBrQ9DwcI58FpMccf8gVjTN91dwx8t5gdqzpsjSYLh
D5kGbb3Y+23TGPTvdvmR78zVPruC7GqUEZ5UY1cQ0BpzLJi+XlTvXITWrGBMOcYP
qsVc1eDqpap6y4gejhgIrvqVJmIuuxonw9n3RnQukLL7XU2N6sE9kY38HJPJq/x0
yQFcGUv6DgfHwxRQI7rDHc0ia1C4zXn2wkXPNglvh1/mgHtVBKSNbQuOf6/IXNSL
As9WyIAN4GdyB3b0uXDBXyKYBWR7Z78ejHe2KXlfbnYJtMkXI+/eTn3d4hVYuNkn
g0A4bhygISe3VB9wgKI/Fg4zvNQpNyBNKvG77e63TSEmERdIRdxRM0tDef68pB5l
HFnzeWSefL1PFv+yprfk4cjjAKoTrTHNrpAg6YaPx0ReQSHSy1317KsgPaCavN2a
e6/EOWtovBRBwdNpkWj2Ghv/m+N+0I82L5JUY1ph/Ea+YgjlbfFXyBBtwB97YLoZ
gHJJU9JImfX0p1yqVEbKwLzJV9L9+vMPGvWc340zSGdfBqSw9G7EIcIXjwgn29bc
uQh3/WnjrW6t3GPAF9Y4Gpr7Aq/lzJxIsoLzSrf3sTijiKoFN8UiRiSplbbHFWC9
3tQkKElQKSbyITPys8KwD1xOOsaxGzeqSpLf0iJFiEd2/G/kcIrBn5CHkEt3/s1o
9W/tPSCbeH51ZTyvyNKu45x2/b9+1ShKeNzQI1olorYGY21WGSOPFIHJDBgftNvW
/wictXfmghbaKPLuBuUtqCRcjzfPgbU7E7DYd+8AY9m91Vb9GkdC37FcLRGUUvVP
MfGL63ay53O8etQP5sPIcizKNx4CN4niMLpfB7TDpJUWqSfh3TPf3R3U0X/LBUQ+
kUt8vKYwjveceOHNz+JvZdgBq4f6lFn0ayMASu0AqQT/QXykyd0XNaFwLBaizDyB
7nh3cZFCLmGhRimn7hHE/dCxZRY92QKnYJjS9uDDf1p2hic9r29/TyUVceW1SAXH
uihbc4qVlz90SwhohVVch+8/APEYhwlr8L28zIejj9phRhwwRfiaEIK+xVmFQ6Y7
p0nCjzpwZfi2/epdsjcntR0iboqpiSctSzcgabMRNmGaTsXj7gZ5Wpug53JeLctj
f/i9TgnTmAaFb5yfT0HoP3PcULTPBwsNRh1MdwMPInUD96pIW8F7VDLHPIK9s4wH
nntb9G2vUoVnxM5w+3y/p+V1usHXprLlNy0BVXu6CtrRtNXqgVYRLvYOe1Rz46BF
veCzBHQmGj+OJ+MEL3bz/O6ekJ+GU8CcvkB8JB7S8cWAWbLnnZexkZNfxVydoPIe
I8PJ7KSO7+ACoFLDXGhsg9kgtvBe637bFzLdUm3/3AXfjmiXWET/ylfhRBsw2S/5
JSjSC2XSvv+1c74BIE7pFx/sysRvNQ6MK4o8Q38Be2+4Di3vnpyL28vaQccmB4lZ
EJZS0nLCHk/f44FSzTTO10YW0LAo/cJRZLrWYId5zUOvcKSisCsvjiUiX0wbVc1f
ZnYsaAkTs1xNJwRE0Omq/OUQoVmwL8stTwNFMtYPyizOaIceeYpkWuFlLJ+3123I
ES90sVGufzZH4tDNfkqU4tcQv9yGNulDI0FLogyU1HJegtUi8e7zRG3rEK0fuAsp
srqrx0xOHM+4MtMQqM0elkjfv07qRw0FiceCv8w5B4ZRQxGz74QYuh70RKz81w75
uqSUVRTr4ZbkhO1k1RcOn2JXav6Q9Epw7ZPCWkpwCxMkThWfgc1blWsKm5yGV2pk
nnu4j0zu/FyrHyvGQBVdVhimFWbAsNweCDfwOl3Q2NIDge/n57Ua78aIWMOidLba
3QaJqL01B0BHB9a/+F/k3b0+3yhsTTi2D+hSm+Mp73xaM73jYOdgZ2h+mvvUEO53
/VRq8TDYitP+ATKigwxTZyRSDRJ5xma4qsNS8si6fiS/xdzN6YEvjNfPO79hT69e
U7p4xR4fRvzSgMpSww7oxJj/6JLmZKFz0tgrHbH3umLO/N0OHpS303PAv7+S+pz1
mUPEYokEsmSUHwq82lz81poEwwP7DsnYiTY1oCcsRyvLfaHHaIC8m2Junasn1cba
n2AKR2xg4f6NYfkUzD1yCOTe3SnCj27T9/v4jA3+piCM2IBRIDvpzI22Mcz6vtHM
XFcOvLB1x7Wkriot2xyfGV88WmSILdiuB5bAXbT+IZkWRxv/jPne8JsRD8n+3SjK
wKTeiljJ6aoPjN8HqgnFWDEAEYTY2YXf+fPhPWaK2f4a9WWVO17Vj7W9Hy0RofBe
948ig+wIg9F76egImrFRggaS6xHjnDRaIGtRB0QxVgA4SbOFyfwN/ZgEFqT/jygf
fdHUopqMmHhUB1TTYe9VHqRG87ejTQ388eNRdDV6Lkje34fVTo26tdTcLT511glO
1JyN5lu9adRhMSslY9KP5mtVS3ZZ/z4FkDLhXGPtiGBNmOHQwQx3B+7SlKIePWcu
WTn5GNPW7aqG+vFRZcJx2EKH0YpB/v4hcThDfK0MwArF7942thsI4RsVD8u/kvsX
6R4PE2+rePKyQtPsiFDsZ04vltgYPJoEtVoZpsU5I6sG4GmpoNMI1wFTLZzzbN2s
QZMP1llU56aX2KkNHsC9Pwcvr7AuwUN/bbfpulZsGS4NO1lRvdAldnPa7QtApN/g
/bijeO36GJaDcaJnRkOK4V0ZjXZobuAX0M6+60fBrE13FaO9imTLgvGc1HPk47+S
SHrLxyq6maqfKtCTW8m/dS/Czktgm5aseVcg1P2GEQbGOQD7Ab5/sZQYswsdyJCr
aXNyPIDOqS3oHbHXzRzzWgTyqG0fK1FzfEg1XAySHkpMHNAqWFfLiri1FkgqfHat
ugF0s4JDrXfcpRbGCE5BBOeE5lBnNhhfRSVBsHFOuvEKrF5wB64On646WwJ/ygyq
6WmQ8Xfo572kAdCv/RNSLgWRPmwB3xOyj8lIVqhgPZFM8jdJXOC3SvWFiH5RJosh
cjSjAAtF8b7kqs0ROkz4mokKupSeY6M2sB3LHCAtG3Xg/DHGmvttPPoUv14fbWfi
u0XyWxLLihANeg7JvKNM37QKw+HV653oCyEXDJIXpmQcF5wcxtSFQWVJvjtL2vRo
uPT/9fPC6UFFCTgJqsG3bU6c5U3rz4XeLBdE4DBiU6Bud1d8FHc7hMhhPeYpvUrV
y7nEIjwPTXGs02u9j+BWJcy+lIQg9WiAnq/f6/xQQyUYDbUjYDOio46T0VijfSi7
Ufgab8DOffNZH7us6iI7eXJP9kt3wcAH47vvU0/DaywxtAaxWGKIAt1yCcq+EaK5
nNb8kaDInZzRNYUV7fxtm5FSIhlF8ds0BaFFXdM5XkaeLzQDWIO+iBthg70ec3GE
t5FgPlmpcD3OZphrc6wO1aCAJnZzOozI2OGbvKhjU+mvzYzJFgu7x+y3WPsW1pby
wLoISus6kQM7gQXjZ99nfoxZ+d2EQNRRG+w7rWp008rsIt+Mz5QiwJPB5NMlQkYa
kFMj5R1jUhKlVYl+RPgubjeqBIRMq2glzCrpKswu0M1ohkfOLtnQxC5JsOtWRcYq
fBRyAzzhcXoYXhdyQgTCzTjyPEt/Ro5Wdq8EgxScaUA9ves1n58dra/XadZx8m1W
RdHn5PYW2DaaPzzNRYmvly/5hH5uYgLEOn0Vdj3IsFwPV+fd/wAM9MJdxDZrYcDZ
9Tgxy2ZklutUwN1ZDLzwHiDRHM8EqdCbgF6fC6bXD4eJTudwDODta6inq0BGvf3Q
SbQitCsR8l7Oao+t2rvlubLPA5Hk8O0QBBxJYUkXuGte5L71jQxXSM1DDqot0dV8
X8Kn50ntAEvJhfqj4URRacZllVVOYB2k2vsAkatFPepJ/vDywxfs2jjzhIwq3Dfc
OveuOXT9mv9UetfWTjQ0q2HKSXKZscGOszs4tGv21qz5nBkjJVYiXdyG99sE6ASE
zxvb9NwzUt9ECcIhM/oxLSVNfv2pvLb+jyIlb5BtXdwYGtN8fS1o2C4+UiRN7uEU
fo/rwtQwuPDUAfbFLbO5pyeWOctsJli9QorxJe/ykUpzbmA7SQAIJeVtCX0BafAQ
QmielEVEvubFcGL3qqF6+jmixU4YeSGIR/NHZzshr3PC338NuNnlaYBKy+Bo7zi6
gwjvinfKGnyo4AnWmk8xdm91EyuAxojP0RHWQe1nIWSPLLhQcJg3zAJQLlS0Dz2S
NFX59JVCtXi6IyMPMsKbVUaatiKix8YUvcXtvjL7sQxIxEYhm9Sn1i3M6j5vC0DJ
yn+Hm4+HGpz63kQa7ZwP4wCu5D9h4Vq/BX+PWdA9Vg/3r4x8RYidAxR1I0xum1dg
xGehekkrfWMYDsKmTSKU5H9TJMwd2oImUeR2R9qnx5fZGljqFIboMqBjVksOq/+L
a563IU8YcvJlSDXW94nSLaQZvtiusOKZhQI5vz73Gt5Rq4SEV/sMrOB9i0cAvg1z
NSf8J7fzVmnCJbG9Qv9scvI5UoPt1D95azyJ6q5L3SIK4xm9K7Wsbsq5SEDYn3LW
otgLNZAb20vaQ0ycd2VL4N8xB802aJQtIJddN+CrAl54nRwd7uPktvKjW6wjUyS/
Lvza8m+dN8X2+rEezGVVGyQ4B2N6Cao0upIeAKv4Y/KL35QrIjcE3fSuBxrD/62N
FgFNge4uzXEhJLwmQN1PAZnA4rQ7+pakrqnzokkLotrXdIK2jyOY4vJRNCuFfbZ9
gZgtpryV40azRSEiG2dbcwb+JvpoQIXGq2EanfPK31/3AVlcPfii8tFZc54K7o/S
mPqTOd2xJ+t44GB3aDLuJwYTlTL2iomXZj+5RzKtsLckBIYqSBd5q52tMhOO7cQk
nW+KkQACkAQAywO97zy/xkwYZKnhpufNv20jy+plTNRu4AEslJyJ4drRl6sStYTp
Z+6rvP5gdiq23r44QA8wb8EbK/7g/uolOoOQcebbsawwXJU1l0wS2LjcMvYPW8Vz
zJSzcEBEk9dlff0RAEiVaaT9e6ie4SZ9z2KSlAjMuUNcDCXm+x0PMkL4vcouxvy+
VwEAPA/tjfxOs72CD/zpKabp0B3NMEaqQM2cu3rMgihHEjkRtGMEufIZCYHtVvKb
s/uUBI79RKcWIcvDXt65rKPEvc9tpc6euIbIMHs97RINWQZo+AewZic13yHDvCwS
foZaHsE6WElSW+LyZmWppUZINsCdEDANop4aVKtd4cc+YLevsJwpfZxUw487MFPP
QeBmC0gHptlGE4HIuLZM5moCJ4K53ThrsPWYVInOzEKCzkiIgPKMRS26VDEv920o
8JE3TxtBY9+JqqmeDuuV7ZfltnlNpjz3xONQx59ERKb1Jig1c7vkKDESdvGGXsFd
eOynBu/PNpwVaIe4CNnXFxU29sHTeVa3JXoZBSEvxC5HuQRIKzZSH9EsWZrhY7WT
Bt8eATulj26KWlKH/ALmmo08vFIXM7FP+3nGwwiF6o1xEpGJIm5Xwy3KEY05UJw2
++sWYwBm+8UYiz8wZyiENHS7qx+P9p7uMDCWhCraQjAZBzEtq2F1bULUDFghzqBq
68mL9jE1uise5KcpDyTxAnJ6kn1Dn/9RJ5qdY1oH15Dr3fbF9Dj763sv7arYgBk8
iYIBGZH9xUMRLQ7MOu9Sa6sUZwszSukJEIaJSIzxVfruNGnlI081koDpXGBXu9cW
qynnHkcgtBorFvHqQh8y8m9QUrnphOt4YRHln5Q+W9t3qSgglVye+4KmLCwScjR0
0VK7bgWEO0pOuIK4viXTXoQawJds1WGbcJiuZ1XNf6AoCXgdcgtAonItc2a80QRV
GLX2PKKQ1ZXHibr+6fC+X5YBr5fWpcyPR8CDlY+ggUG8YJc875CavU7Hx4XxyAuC
FXEqM+soY17ZovDXLmpC/D1s/GPHGcPuYHdn39Ih9qpyoDod048x2DFpZHbohKwB
3BHSNhAkajh3AYYau5rPgh62zho7YSx8fWDorSl4kKal/Ossla6iM8kqwBBk3/rX
H4LYFN4DpmPRemUTyd7PeXAql7JayRTIQ/XGPH1djz2dd+AkZ7xa76ZW0NFKW17s
FjwxrGvtXwk1V5CoZhJOenmDLayg0ZE7CkC6ri+32T3WCmwPhRW3x8SX3TGmgg78
7KFqffZ4xYbkzs+CbZJcfDXGqfjO21dF1h2aida5dkPJU2oUgHzDg7KtkjdMgKH1
mwZgBqIuGkOBfJggE5zWPOIjlakmsC6d11OGpJaSFmO5BBbg068oajLHxA2O5TA9
j1fOeLF4AxJJhUfNniLcu+0A5AMoXaQ++FAEv6PHJPAu6z6mZ0aAMvK2AQyNgCgH
eHq73903oggFPD3RLHaptupZcoqPSWURake06JSMBb3OnuFUOAWyevL8mfOnnx99
t1eu4oJKbn5NIXpIoZzbLx7PpeBzw7C3oliDDJCp1lQLDHD3bV/g9HsQjRibPNJQ
+H1CU7PONZFRFr6L8lRrUQHcez4/BRfed0UQmh1Ad/BK956LK4QtXZ5/MzLivUq0
mK2TcvvT87bWyfURcCC4yZAPFSwgQ3enEGwxCHS+Aa1YFLxbt4U5Vs9KqWSUBBWn
xmQ2umFIB4MxW6Mn8rO+mquQ2sMMZhB1Vz1y4Pj+9TqSMetcybeAPf+Kej5OAhqA
KYwf2KWbQ9cHKwXpTJQlWnlQVY0D2bkl1xcDhJDXtG6WuWV8PjkVvyFR8LpRXmY1
9kMh0YAPCtr+86Pd8X+PgwZ9qQAY7nncG4XQQyh/2FShk6qwxduG9xx98yvK5+SB
qS9oqjbQ/bSK9XxG/rf6sji6adwtqh0dAHToun0M5k+NAT9/uvMd0nO5jgC44KNK
obsQ/vVPAcUu/0XNUP7+vveWWfDG5LHJpHYkrQcuxThN6H1mHiuZ8VEf6jBz0psQ
8L0Tb7rMJ6Qvsu8natKkiws9fl0MQD2TVAGS2cYKErnqFNXgKYsJ2gTnVoI4zX6z
PzLXoWFdUCu8vfpXTBEmF0bXo66InXujYhZa0jlS1cxuwt7TxSuuo/kksqpTMthE
TPSorrtYCi3fpQESMRoQTJHEUG/aNdvzS9wdvC8tKQAk/4B8b3EB0ZUryHxQ2Z0I
h1gyaHBIJqwP8G5tYYyK9R5PPhvVWaUCwjRQEmBBQhJYIclJONTovVSKfXT2FHaf
ZFShqIJVrhkfuAf9Yn8N6Rkd87BfnKHHOmpLlwzKNd81vmleARF5tcq7e69simO0
OHQMZqZyGwDaS9VZdTGVaoZi2Zcr7rINUKptWQh1M6brWdjcjnHvxLJ9grPGsqTM
kUK2abtVXYRRx+nNzT07dHaW3WYsQzTCIqkY+A+ZwzziaHQZ2ly3UanTKhBw36vT
F+OMwrCiwnfmdgNOcvS4xvotjjSCuMdvpfRgkT3t1zyYpUUWEso/JR6tZ9fkiZIG
hPaeFPxU5nl3UP8IVMqJk2rNBKSIlYBuVWYp4wz5OKuCvnTjf3D5LnaGtM9b5CnJ
G1vRbSCDKymrKofWQIKiiBLKKBaqxByUJnCNAMEh1zYepKextu5fxSavGM8IvYUz
kLRbrYWXLylDOWD/R9knVpqwBAOeZQaa19Y/me3AlEDi2WwPFy5j7QP6LqtydKGu
fApNYOIQfw61f876yW1gZ/GNryi2RhPLUtWn1lcoQtcv1aqW+2aSNSEri6y2S0Uy
YTLvPoxef7aEw9rE79eddToKqYYXVvXVaqYZCuc+prIP/hSBEqHuZ7+6UuKj/nbV
mZimH0eZaGK9mQ6e+cT3RPRWN9Gsj2U+lQ/XhYN6xx6IFOLxUjuEBTklujv9g7gL
mze/xSso1EPGWt8gkdWQWfLxEyIxrtC6W/4Q7Oypwy9Hppg5Bve5T5d5jzgsn9H1
QZjXIjfn5wkuZILj2KbSp0e0KPn/NUjjrLxp/NgscVon0FLAfvDmPrfbIfI0fjjc
vBU83E7J8TYUxNXSMAWXBlheRw6HFJIEJXWfaMZkbdpStgqgeiZDSfF4qh1ydk73
mp530Z1MbR69jZNRzfv4ptnSJ6S/O/In+Vmj090O2LZ0sbH1tb5UpOtMfHoK/iTb
tXr5q9HCeiYV+bn/pJuPq5kpZNJNXVv6ocPOm0PutcVq6WlSPhEdL/C0ctRKcErU
CeAXjjo4M0fQs1iRGCK9WCBfGF2PHdcHqufJa51CbwHZZV/GVy2wQxwQSyh0Fsen
5MoGRFs33ncJveN2kZa7aNeEZGdoyHN76MQ/a4ytIzmOCLKEKrJ2Jyd9cXkTz8VD
KGr5fHr/5FEjbgAokitsOh6slWhz8AiYGP6O6MR5gUM3SW2uur1uu2v5gHDjGMNt
S9DcbigVJdqvxxi1BPHH0347tFtY34yfX08BMYH9h7sMoLUCuVcJdd01suVdRBrt
AfJcCiJPqBE9x5OuOuIwrqlPUGySRKMrQEByQS3fruugB3+ti70Ej1V2eRLFaXqA
kmbICNv++8pQEz8qIm84B7vyvvwzeO2wJHxYX2YUpB1gzBUwhyz5Vwn15lBzfGC2
AE/PprCbLQ+oRJDXLRchFyWtDhlgEh7+clWgs8yDmhdibkZpQ1dfQkL9DrxlOkel
fKG3REq6ysMnygsDYs6D7F+vDTLbYaGnbp34CmNR6k7JR15htbBH6O6vrHY5+CR1
iijj2brceBoVDhu+A4SE6E36EigXgBr3zu0HEORErRR6Kp4l/rrxTl2SJZVDjO7f
39alSJYxmZ+TuKkRhX5IwajnSbbgwDIqpGl+HO/Dbzgz9YXaOMoumk7qMi3uGg/U
rpZ2IugNCRbI0jy1T8RQPVJs9MyZOufFxqkkwxpiM4tBUoQn5A0jTGQ5zzya4c2Z
bPWDsQeGmgbO3cj31utYjJxunkT8vTcXgJNF4o729/HZ03qF9lNmNhDSl92zabob
1b0AJrXban3hRxfl2Lb9GC/xGlJezLsnHtxrKMfILF8NhtLdeuMt0noM8Vauostj
FtozcKxFMx3cJ6pTsMgkn7AJ8N6BMF2KoCoxXfggPKuW0bP0alZvBQVAFgFz4a4t
efCUM4ntwe41+FQVYG1haDvrNKW9gmB1Cs/Eduy4odfxExwYx+watvNXkUz/axCl
AlId/gGMHqsx0VHgxRARbgfWb+5SrqZk/C0BzVF8tpJt/19NrKfRj78meeUaVvkh
YAmuVSyCBghi0om4IZ1/WhVLt0sAywLTCDFShHFn8kFvyIF92+TLl/3yMQWFmvcD
NC9OcD7MLKYamCRW1HsvZ2kipdbVDBLBBrnLeF9WBXV/4oZGE1rdSkRZwXopwjaL
CNUKJas/G38X0r3mimU3lOd4Y9A2jXffY1VWT2HHPOanUSBlNfL0eVgJCioCZGbQ
IehNRDETyIXBPoY0CZ5ZUrtd/MXPbRl8WGR7lg3q9pL+HVMKhhIwhedM2gCjKzPd
tEZ1udUKf9BeU+yHY8zZvl6z42LnlrWuyssIiUmsx4jbmom9bFxr3l3b1xUyjey8
BGYkjsT72btkIc3xpalV8qJ8cuY8VXZ5tgwLUrXCexFWdwfkMY45vcP5EVgMErcc
gMa8+umE8d434YUy47F0bZyMP4aVlj3qPih9c69xrVZva5UBL9ddyiCUnxSdXG9l
mHfpxEOhXBJTaf0pPVQ0KqAkphUKtz5G0W+qtMRgQHc+wkRk5S8NYIASydAJytJm
6BKCM5PxwCYadfo0+NL/c0Op64WRjB62kvA8Nb2rme62N5UEbklGE/FX1xeuBfTw
FZtW5PkHAT7ebUa8UlIHfL+7JI3/NeURnysRzOH9v6izmF72jXX+LjHmx4mHWSDj
YbOt695g8O1OOkUGPHYQrZdaKsco3vsdjuq7Q+2cizqH+YX0g/pKfv4E8V/qo8L5
mD/jdjXhyVmpHftL4uBoXZLFHzHECBp7D6TP7p8BxyDQH4y/Qp49UwwaQQ2AvQRm
0dQPXlId5HWg1oEvvmBZafQGl4Pk86ZJKBqBxZXo0zQH2m0Lx8OKtLJd+CEhnS96
m3WgddOVfAUOcYyZLU+CVYO9w96fNXtyhiG1yN9VUaUhPlh4rs6+TxPzvnrapZjx
lcbwvv1+9kj2Ps8C9dmr8y4H3iCt2hln2NhhC+sVFEHPwq2Kog/I4oO+zvMWk1OI
H14S87jewfYedF7C6Oj0UZzxO3hAj2TCFSUgP4bPEHhpBvaPQygZR+C7gzJH/8g0
iaN2t1XoBozMex6OVSaTXlnDmpa9z6BYssBkkSftcF7Qho0ozZQtb55rYT6hGUhP
M9cMHAHjD7dHMLDrjNsIMxPOEBQnCZrwwWjmdaAm+MTxxMitq2LydwhShMUVW3hd
+EDufnEj4ZzHqIYkd3r+eKV5vhWE3I4JsuLZ4hiJS0885ACeeBIKdOQhCNK8SEVw
NxgVzwyzubgk4x+0UaD45Q7hGfnSEtPuopUJbQtZo9gAzZLZcW6YfU7hvCtUl5dq
8x34Nqcv1t8Ck+KG+trUXLbo1GinItoegJnISnUm6V+NByTF1nWq9uw3PG1pm7/W
ou0u7X9LTLZ5WgMUa1CHWvh1SK/u0Kf7mBS84c+LcgpAX2+qUNx26lj2+nhPKuEW
NO9diKBvzRGwxyHiZzZxBm7HFBSRPHbr989V5c+Ga+FrlMJyV1RJAOmynCeMT9nM
UntZpivZTyYHkRcz7CQKxvc3smnaYwo1xQVok9nf0rO7Hd1M2k+yUKgJRFPDgt1F
AjN32+/NOA2HQnKv4gSBwVjv3+c/ZTHgcqmdOYpBb9tqdiz3+/N95FGQ3TxGOE95
z3jWJ9SZGP4VKS4aIemgeC8BZCvtIfGGdCPNN/13Zws0VTMBI13WOgziLOfQ9Uk4
cuZm2qd/KiO10GGetAdOc2EYF7sz9qEPCf/5Mgf40jH/dkdQyzud/dyValocGYhB
tUUh2OqGgt0Na9R39Mm/8EbG21SSqrH2394y0nXT3T6DKmIB2Vdlvy28ufqb7lh0
SGIW968TXVNK2z0Rfpq8A4AlySU7vPyAJP9t1dXqqyJigeeOhnpFVJpuJm4kExkS
huDfy6v1Wpf9E7fMCtCBamz+MimAEg6VINVninRSYha8NuoJ1D/fMGQjvLkVitmP
agKCVXrS8sPkwN9sM37Am7CUDGAInww8H85A22GC8qfLu/hl7tx0yPpbbcwinXM3
T4Crn5VlcrkvHcpdQkbEQOK4NnTSRkXQ/UpjFVDfgOmRBg+YlXDtxUOkaZee7yjf
MjIPC1kzNt1Cao+6rBWTwf8TyiFOdc2ALrKiBKrPbICXcCcDiSrWjVd0rsv0MUid
zF22pLoXNxb/oIs+hwwdkjwIhdQTlQFNrgRvx6cQMhEvKDU6wq1OiBvUAebQSFI5
jbzCsXwqF4A4hB3u0R7iHo+2TbOu88j2/nr3du6bBX3QpRCF0p20K97x/xohkrAl
yFJw8nncy3iy6zb9VbNLJSDJG87QAwZNopg28ExCd4vb4owYYtedA0VJhVihDIcN
kOgfungPFdaeL/srC7vU+mlkhMFY2tXZkfzeMtn/xmrmApbInSJZXfooJGjwd8Ek
oUkMT1baRtYFXqsjsb7eKW9AppTqfucPJcrqY2L5jtazwWYSWI5bk6Iq4bbyQBy9
HEJWG77Mc+FyYBlFjTNN7SUjGChNOCp/xkHSALcaOab+K6s0jqEmyJUSNba6Jl7u
WKrgr/tOjQyUjNw58q/F26/Sei/Bhu8n/6mFu77b5VmTQRcLB/4Am5qyOaYEZgZE
IJnP+3gLbaaqa1tDHm606SWlmhRd/R6Qudddi3QwzhWnspB18uKNr6M4/1hLHJf3
Bkp0qzPllIBMoBzIAvLVufiqexM61g86lQYtt2g4UvSYIL8tfG4d8FXBuEbGs1zJ
bwl19r0rEUoUjio855BLUN4Vl+G96qAqVSe8Lh1WyjCPAdk4EMGD1Ypqdg+bMzgs
0L64SJgHRkpR+EAKhcIniMEaH/7riZwOcoPzBrGXiizinyTx9Dic2iCpI7rmBK1q
6bra85gycFcCnvzqK2VarBvIUo88mHJtsCQHCqgbcDL5A1dMpCNQm2yVvXcCZNFe
fq+/Z8Sn8DtNHiSbZ5HoPCmPWUEsDzmHlVQm0rCLgJudiwsq5NyXsK8+khsDYGF9
xLEIyceZhbWMdJ4jVojnfkztkT/vNM+EKhIoG7E2Hu+7lX5Q7rnkCMZj19m3yGwB
DsaBU3fLdg96qYHlpBLOqdHWNDrYHelg1jdAxUkgqgq9unWv0J1bBpzrAXYvp/Wy
oEyqPM15UdEWjHPnVNxhX0819+br7h9K2Z5jgnD9QyvXzaucMfeITHoZlhPwtohT
DlGJSyELiNMaSDfl94cvYxzC4+d/7aT9DEipxmdv5bGs9dc+RubJxQw3mX3rYa2B
48nPtepZXd+IcjCPIiZGVdM8yQVD+2O7j/4PZJ35UJn52SonsfusELyH6iZFtfZy
ZPJ+Qo177oSrWC4VZENQ1He4SJAKDXH5OS8DPaL8gTc9Kv7yzg7egBOCNtVXs2kL
wZZkxzui4PgMTu/uURpAQlnBOvsti6JTYMBZYao0MYkWz+j4ss8cyXc+rDQoiVwJ
sErrYWjzRipEbul6GKzjgZ6nUuojwp44zXOCDYzNQxpo+zPZcfuWO8bqgw0GX5+Q
fABX9KDhb7lPwHHzPz4NyL7MMDn8T5jN6/U030OxF28nJHcLJzPFfiW+d9E5sxnT
6bQRRhweCn3z59fa0kJ62BsZ3p6BsTyIThBODbRSLOMhifoFi21EXTP57nO+D9It
dpr5vDcgIomdsTUk1QREG5MCsovWlsg+nstwx0ygzZH4FSTHxF9/1ARCfcwuWcFm
92T+Bvpe3Ea6LbZ9pyg+FD09ymC0rPRUoyEnuSFXFiSYUPj/yCk7EpzYWPFMdb0l
VlhFj4Zp56bF7TZnpCxRUTkfU0X0mt2GrCi33ZEailQmlndYcYhuk3Oon1ZOghkT
mboNTjeXNs81HL25l50Hp0F++I1LntXBeV6fLLKhTI2gpwpKa9Ezy2ucasC6uFTa
1IE8GX2udfK7FgympKqeSTVLDwUXvENx+5GiiAEF84HOSD3HXpSMUUjV5zzFawc0
GiFnEHEs6ej61+5GUcNUd/jRIZeVd0MfHnn0l656h3xB8jgGFNDasDJQTckzs7mQ
fGh4zS5PZ1ZCEOq3Ik0D3zxnFyGKRnhVAa1j5OSwpZDGJJB2289JiiRrxlkTqHp1
OtDCEIfhlr3iVnSSbG4Oh7m6fAM/sw5MW7ZRJgE53FyJUsD0vFciVgVfeP4ma6d/
NVFPkAmqivorC2G/y2hJ97AsBH2nxyyTCcMVocdlFZM+7Y9mF2y8MEaLdc33ymq8
/76yf0D/eyyF376LKDu7nAnGKf9U8E5koC78PQFw9zT8fG+Xbcfv516P4k1Ku3T/
IIIFdSELTAPsqJQXS/g2FmF/jf+vwoGXAKvczYU0ew9pMK3Ed/2ZtvSe0cuFi2mL
q0w+yrV7Cqc8gIdMnKI1ycxe3eZoMr1ZfFHY1Xc71/SzlIfpf9RchQ2X0L1GYvEt
4Enn77z6MM2NUYCN/wgX2flTeVRSaf6RZ27qn0D+dZgPgIUzpPbtTRgZOOLa4n5s
S9xcEo4z1cIJtBJBGrt3iyiGZyRwMFyUuqH40r2o3GHclQd/n9w2hcOIDAXTLE/f
SHM7DZ6zHZhb1NDYDIkDmNg5BqBwM6/flGZKXU0zxQ32PHhQRkMqjAWFj4nBhhOH
F7+7s9u+F1wlG5TvMCuIqnZWtTza9Uw+lHAuiwvyih87GvM/49Qs5dQ9jVLYdFHn
maxaKARHG0UQRVwZWCwRGJLhatZ56mV6JvWCq7AATg9tK8V4wFaQvnQiEhl+BSH8
tpTIGi2gmsoJolZR81Og6ztM84Bnv8Pc7wMUaYPFMWvu8Z5BvLpmymt0m1OlXkYD
/m+gP5n47650QvDDPM7UDxcUMwft/k1K0PWwge1bwWFv3BkaXDKzabsdmm314HOo
MqBIgvQyIj7Q47addEd16W68OMSwKzt2R5P0hYChP3PsZbV1sS5RsB6xipuesxBA
oP3mQrkdC/BAniry5Vcic4bXhHSP+uQBB3J0PPpKMKL+GzuGpH3m3aIwZLZaTrK1
vcO28A06175ClVQKmWkvdOH2TGgB8dQrm+7hpVjK+hnWFrh0aoO38MKemGFndnpV
BzSo5Pv+s8JW2w72+CgJDT+BiHSGSchY7qZkRvSTtzQq8mAVDhKHt4SeEqNRVN8O
18VEyTIbl2VsCTWxE77Jkl6RSUV5LieXwgtl99KU5in05kNqMobn18plg1NpFcad
9NVxHxE8ctcC2q3LePfAulEEZ6B/yXgSLPhXoSOaASGCHXzLK7yIzCKk69HIUZai
BBgnx7sgzm3LWjFL7DrSngDkzrcEOIEQNqgiVlWDCE5A+2MnvKNLpAT9SASJTTR7
X8hPqhYjDXUoUQNGVs1RX4WCAq5JwlYsF5i2cc0IZJm5Fc0xQyNd9ZAL61Zeween
kchANQDvYOpzon0kH7ChDjJO10kZgfhj9Imd8aftHLVyDygfN9TvfEtrVF/TEVOZ
CxdP51r0CLvZJDTsngssQ4syig2bcru+ktlLjz9Uxb5sdiK3EBeZWEnqmeL9xt0f
ARhh3RSwxiUZvi2A/3N9wQiPwnzcmsZfEMUK3lqzacYoyUTr9y9DWMPqr/uqNmZf
7P3A2M8PL3Yd6rX49mRQFQ+wd792UfaomN8tJQYO+qsrYX5jNWOhcgSidlc5IYVV
Mmyux6QDkG4ThB0IgN95/WncTJWlbI96lj5AcLeVuKR0FywSLVVtlU6Chhkwvhgl
AMPP8Nti7FFmX8jVxg7KCnYH+vEmcbk+6d9Xcfkxq1dmwVm3EkuYDUjb6bwN/xOI
WwxQDlf5Rn+LRV2wZZIQjLySaSrrfvu+IYuC7wTVvrAX/tqYpRYRh9KtBWfjJr4S
GfyKWePSoBbh0kJxDcxwGz0qufJ85EN690PLduzk89D+SvJOfZkEwhecsEfXfUW7
AJ/KcDXF4MN/p6oEougp9vgMex4nDnSHz3pqadbXREgaDLrCxtz07aVaKLSfyHV/
IXnxy6Ws5j9XFCXD/SIhZEa2lVsVp6JI9I84RVh5vdLIPjh+hhU/sbamyqrHJ9pM
knjzqMHaovzBHVslpMGgYZjVaelPXn7PcBhN9UTOaMHPG4c8RMWQ+RDC10rdNbMv
bCue3BAwVDYfSsQw3nJPDf9G7rPq5oon/XBjfN/dxhOiMl9GomI2V1EP/KPN2Rwm
VB1kiLGCBgOJ8FPCy1OUGrEC2fTjgf8JLIU/yuqhBMe5nLME3U145Y6W60e2fC+8
JdO/Y9a0WKGPFgzXj7Khw7jrXNDh0PQ0lIUq7KgBwdaBi3sBgVcKxcnZed72ZocQ
IH1Sz5LyM9mRiRMOAnK0KpIURrsoCPm5ojuqQ/hbdJuAwgieRU+mzJW2CjDbez2o
azNGxd3wo7/yZHYk+pLzhJVJilWmcxZhLgL7lFAsp1+/fIa5BZXQuMp5VMkdYzQT
4AonDeo4J8AkD/pEQ4DIQYR8RNciGvWJApWX/JQ9LY3zBDBdByVSbBCOvXGqr0TG
Nk9jS7HB6Jx22VVFfWvINXlf8YX4lZnC/kvtWbPuqHd+XtTfvU70/Bkn5iUFHjjx
JwEog5tZk+DyE8CGvmB6FN4HL59s8Dk6SHFvmdoZDv/sHFmaIcTsnugZ2tqKZRjn
IU7h00Qj26d/gwMfR2qmIg/TJ1niB3NCvCH90mZjETNqgnE20oW4xjK9IDp4Buvd
1vdxCtYlByai1s58CgoyR4pGb7nYPKe6zFffTFo8W7va1taxAa22pmhRVtgU7HWz
Pr0cs7n92yhWyW+GDPaNumIrWbyVelyj4IKbMqtTrE7YZeLitX4R1utzhp/SwSVB
ojooxsue/Kyn7+N5eYBg9SPXtTyq66JTEoHGRZwapGRS6qtzZm6d+RckWGjC36Hb
QuL57y3/KXdI4MYmYX6XB9ijm9hfP6mK53qEGdaVca6fNQcon5+TxdyeJOf97BRf
/FcusO4HDM/6DGsM+xPsertQYcg3RrSHKqOvPKhsXDPunVYa1pMtimQyRZSNCSsX
k/YPhLyYAjud1r7dkXS78Zgh39TunIC3wTHiw57gW/4Yf8RKClB2C+apzmLWQ4eH
68m3cHdewwm5hS6pOtEvDSJJGqr/AOKfjDKoDJ862fCBvpubEETF2MdNOFJ7MKGS
dAhKJUaAngtVJ8xWXx9SRmicbo73DB7UKtsJRlq3JcEGX0BUYq6PgMOnWePzdcSa
5tCc+Hn65/2qcOclfCr3WahN/XyqMNUuE3LkI2Sd//T12OMHVrQhfyGaXSZmzrzC
VZcS3rlTHzAUVeJGZBLnZRCndxci/TheSvV6gOsWgz+PjONwvuvuBy2r2N+Xff6X
iwebBtdmXVIjTS2dEqqzkJv/wVJFEaHIMQz/iMtSEENelO88/4ftu2ysZhm0wVlM
+CBju0hhKDLcDAHPONVHap2mJKueTYPnhfPAAtrKrzxUw1/E+noeZONDfCaD9PDT
ZZgBfjGKXBZ4fqgSsjIYsEewGBUIGXn1EHGYqb6iqI72jGGhWY7QqZzmuFljDQ4U
LYDWj700tZQn482aprsBygSLrOEQ1N9GDptphIrWVpDuV/Hy1bURNtHJqYMz4dIr
3Zgj09edmz0y7UEjYlK/9mjlYQVVXA6lzl7JqeeYKTuaZvRMHz+zuIh5xvF1Gif8
UlWka4yFlRMjFdy4RRYYbC8ZfkFzmBtAdnRZfWD1I2udFbLPPQkIcuVM0h+PYHUZ
YJNrgFhLQFKo2hIxvHHQ2pVS+hmddC6et7jF+1m15OXW9DFLeIKyS3PTiWWt2NDy
WVcQk1QQnvJ+bvqQga7pcZTMTMr51TKGkk7I/zDIF5X7/CZqH5Vdc1d9GhUbP3wl
+ref9BrAspc+EYLfJJ34fSOqrSf/t44IPsz+nkfaT7JFdZjG3PilHmblIad7zTQj
HjLGAiVkLwP/4qFQ1ZI6cYkO06fUqyT9AJP2yQxa7GC37yN25yJ30eyNPyQ839XV
0ITTfkIJ9B5UZYRQSqsyskBdP8V9LJIv9GTYwM9JKXemchbmHBpxHUww0acyI3Gn
KspRgKrYfkZCz00c9xgtlXO3+XhB69M90PA/n4Ia4l06WY2mMig5sG81y2h6TuAc
cuscRaJigMNqudB5K/Bv1eMCp/sw4l8YIV7Tvb0HoBw86Rd3MCFvhSOb78A8DNy7
t7wErDv/KU1mTnwC/q61AR8KWRDLNAm2yEjyvktukatfsSB+2csrQ2OsRG7OUuCe
ZY2DMafZ0cy74khyiU8z1sJeJWTw0YuxhI0mx/WlD9CzaYX7+4RjglETnTWow36J
IhSNeaANOIOyBIfVnUCFgH46CHuzfQUzup80fb4FPVwixW6w02avaIwjxn0i+pUx
3IWTUYkZL5imWBJg2ANtMoELeQEGPDibkxtxDq9MU4QBf4UkfMrdlFwLVfqbeiEZ
nqHOFBpxaJauADLjeCy3qCbsIF8ekjmZsrE/DMjAqic4O8khKJKSZ6/yK3vmB/Pp
sc9s6AbOqipwQOaHbq7gQIFQ7ImKtd+cst6upU7PBjFS0ABmxD0lSnTQNPTx4zpW
p2U+hdhMaLwum3k/KvDHre7BL5Q28oz/evPXl1kN/D8oe0vrK2fqlECj1XngZnEA
FzRGD8ph9RIMikxkQzXSvXj2yHKP+JtBJcmZDPYrLR+l1j2czIuVL3+7+idTIe6o
/AexfwfGONa5kZ7YHGPVSZ5ay6e8NNBNGQR7Y95W4baaGI08fFXig9I5N08s+3at
BXiS2kLGMPvtMU5T2Liy0WxPZ5IAsvWbXMM8rCYW5aajC7SkneMkt5CIYP9N5b7y
lQJVh+CRG7ofnyyRTShEOt+1QwjnhriQVNsZBsJ3OmgS33EwCVTlbYoAXosVn4DC
JunJ6HdFDlBPXSf/CtOH3m/dWbLLFN90O+dO2zaWcJ+cbI8y0zjBVms9ilK66b0k
eR5Obi8ONqvNPMcncvOclGAy6G8v7yy81/fNGYeHoFCrVz6XfpiNpALYHo4h/77x
Z2D96RD3bmMaKzpT8iFx2jDyGbGNBnWlNUFtbWShxCmjR/NThGPdQzkX9MaRVKvE
GAdvFKSYAI6S56yVI5GZZN7GhMRjz5XMj+Fl+wrjHnsBLFQPCVm6kde/YOoPsfdP
oXMaRlDidbLVN3f2n8ICXA7rM7v2l0o1NNonRbBQOHHwEdxn5UDiB+XAuuW/0GW8
5LEcgnJmM/YhdEg+FLmt2cRLdPyvJCCzKFRTtVVtBd7z/PlEwoVprxaZwTNrhkyN
5APjWzXjNytsx0D0X9RXCd2/vaO4H5BlNLET9MI9wDJ5e4s9fekvfD/YpQD21/CT
ZmO0kDVNdGaO+2R6nzBG6LcSFrht6gagjkqjZXlcNLTXMvliolPmjzpGTRRUvzqq
wJxPVT6DPoaMEkB4856UjOj3OcBY/EsE5tpSN2S63Tp/JxulJLJ2NUkPFbIL6thT
oDJTAVgVR5W6FlSZSKQ1xbhsqIBfwI1uuCKMzuLnzn/HekEAcVnafJbRz2KIbUW7
uu7ASlCvEt5LrPCOdbs07wj9zQjBjRUeSeugUvi606Ns+vgT0/u22DDMqpX7/61g
5yhwRIFM5twsh1WpKQhPi4GwS4m3XIGVDrayq57tBoGnqiW2F0dc37COHdsW42Jx
ytUypKdKfn3b8EwN2QP3lUUPERpCHwpQRI98m7tPNKfxAH62Hp4I+pe3/E427Pv/
c0UpvUjNcnjWIdYWXmMPrbifm3M3J6c9qyGsD+c3P0lh2ab2XX4C7bLTPfTxJ3P6
s/qWMSClioFbj1ngjhJzKL1exKctlCN2XlBU+eXqUNkOpI1Ux4R63puTF/4ee+Qb
Cc3gxwoMy+jXHgFcRi/jyWaZzMbE37Hsn2LYCQ/WHg3xXkJCNvjLVtquiIlJNiPI
OjcFHMmUtO/gOglRhzgKt9731vKdwnfMZuvLbhQ+AAMvH8uQ2jPujlKdk8MTxZXI
To4jPWMatNEczV+L8u90xZz9yIhBLeoMlzTmfj7uYn8qArQmjxY0aUlP0OpcRGMy
MtZeKtt3Ao78nc+VCVSzNRKhrCXmL602W+Eo9UUAhhoRuIw1tog57c5qlQcZbVjz
w+h1qWO8+Ot56lEP7YhMCPmjw567pFfcON00MqEQrI8FGw6R+fd5H0nj47xks4S2
eXUmuyL0If9qFm0HQ3ow9u81tunzzNPRxC1dXV97XrWW9/jALgRBT8dsk1kEGs9c
zEyRiqoKVVYjhphoos0IFMXt2No7sexj3xxNT3hvBzrwKaGgA8auC8i6iGKgJmVl
uj0B1kn2d8szHtzxnBvMDk8ytx6OlhPRkrBB9EtZpynqtRrT6lfxXA6HtXwp+HgB
PlmYif5kwczpzHANRh2zobHou0dNvoFGxN16waflY5c4NodthNOJMzgD5CCW2ctx
smbf8brUUIqDW3yHukoqUfvk6fEQz17CDDu68rImMHNfSw1CS/VruhvfYFTNQ3xu
yjYqZ2+4BZtNvz9JSN7aNdcsnqsqMYNo9LmKoC2VY0sKJXCQfMJE/uBeKfT99pLO
pErpMkAVX+x0sH5Nmp5MD0+NwmluAhcyM2ExycdKCyFbIgLzccZnbIHNgQtK3E/k
Fgqg9aZS6TI71evZ+tkSUg1z6BiUX1ccEx/dooOdTUAtuzVTLD8oe7EnkTn448mq
0tUXp8HSGdPNYlvBVgGzJjK9Sj7g9NxP6UPClszwcwK/c2Lpu9/Sf8FpkFlJ59Oc
t/wTXBNUydOc7nB2U2+pnkLDaXSqRuFtb+VN6WnmU/qSEFkNR+fJG+UcOVBPljiP
DCIVVIUvFhrnOF43JGkb5xo1XiN744VGnWtguqMgkhtasrS0N08aT6+ZbrEIRRuD
EZMnGQky2zKxmH0t4YLThq63Ob1hsyjXGuXj3ZnyJAkmwy0kstXmh+vN89Vzbxu0
KIa0t0uhvmblTBs+zA4xMGp4DuYcZfzDX2y7mIxmyf2C3HxnR1CbvZ4+2g9G5v1z
+OworDH/lrBQ0TTqH1KW4TswyJoU+ali/zMl6QcAUZ0OFoDMatbzmNK/EfoelwQK
HA9irtXmTBjWTBCSKGmc9dQkkzL/T1grz384pLEc6jTBiRp/iTLwgm04Xi1CfB19
hOO35dOdoujTEPK+KMqwmV+Jf/InuL8nRLxDJ2wGsOhxegE7nBNQNRZ2j2CqmP3b
sN41WHGhERzv1tU+64IH0ozsoutwqGRcqoQvIAlfSd3HWCX9OYWolBPOeVYGm86B
1Fmzc1oGG2Bz/PFPrIkC9sBrPmdgadECHjKVENCVU/C5M8JnoYWxpk1JiqEcYD+z
PEjHsbDywcrk8BkaH+UCj22J1D7eoVEKVdHmo65G40ZbwEoQA02hIVhZpzCMeodk
/nQs+Yf2c43Ba8zfHL3SE5lSGcRHx/zQZmHSueRP8VzXysqCOyYz+YPiUE3baO7c
H2jN0GwM3L5mb23ax3JB/rErSFftrgUXPoI0rjMXYiuaWzhV6Ng7ip8QCoYQ+wPm
OX46s94le2KzAps0nI7WH/IM9hiTHGHfNhIt4d4ZDoZvhNE9L6V7c4+svcZzbSRq
DWYMToU0R9lTfA1Hr3aSJkCNZTBL/z/FyMKt5RE2JYcnGaD4xd3ue9dzRxhc+BDj
gK63Vrhmik0ANF8uqCVaKxyPyN6pRlPcJhqvl4Z/8O8pE20F9aZouuRgu23R2eG7
WHS8l7tD2igR1yDcRQ2AZtddaK2bx/wcTVDOaTuIx42X+Hy/0IFQTXqb/0gYZ/jE
rex+duaxz4v5JDWI8UCXP7xtMc+xuNHvOKmq6ZfRYtAInvIqO2hMMLNNMrz1fbnj
cIvhg1/eDd5lbYsAzMIfucd+rzPvLd84wU+5M3LJ/Ogw5N2mrYpRxs8VY0sTGkmh
GFfWZVIWzpToheWiBQsGAT71veqpzdmzcmpXg5hMopxhq3UsHy5xEyeVzJi6kyIy
6Qv3u0MK0SsDloK16AcWxrGsfpUMTA9grO6xmaxxrfJ+teRcpinq+xEE9YRd4I7K
YohNNsaxxO/Qmq8gIuhU6w/tafEe196dVWQWK2mQoisBpZSPyoPVhuePdpvxWad5
gG41LBuqjngKNk5Rlv6Aod3K3pP7qLiE09ZKSXKYmwF/R1yvHdPAxR3c6GwlH9OO
07mOANW4sS9pZhClPg3S0XjJ5yto6wFfx1iiMYXfkWZWr/IB5wuZrWELLa0MCbpe
hAIr/WaxXusTmxOs9c0/lglgrUpu+lsps/Rj3USBxo5CQbmRNkR7KSPwtas6Tgpe
8uDKrFCQCIlRVj9y8gsh0MT3RryOwIjBnampUNaCKen/clA2QMUDsEWQ//lx1/bF
BsHaq5RqhOsogEHBpYTrVYbRn96Ub8gf6ov+T7jLebnPAHnItagmANFYL/njU20x
gJDjJ6Y8LRba58v5hS26RDuUY96EgMSQSTA6HnF00+gMuE45tEYbDcfgEi0hkEBQ
J9kh1pM8dBxm/UzEFnhKpOnNj4sYH5R6LU71Iiz+4mEd6V5O/dQPCkOXkzuuRq7F
CjuC1xl100tkqE09In7Jnwvx9NIwyptkOHvLJAGy3LQ3wy5VZHIaR74cmJ0CD6CB
nsJiq/bBgyMYXZXftVDieg5iuP8fMcaxNE+ouZYYw+tWzU8S4DEmhz3bqY0v+sUt
HCe8LpfpDfiFX5+KVCM15/HHdQS71SVmE++kSsP0iJTK5gbWng6nncSlrIOPCVEL
q7DLSOY53R/fulbKReA4Nh9cy9oevtGaM1NNIf5P5Xv0OCaB355FdU5DumF05+Ac
3AXFZR1TI2AiXlph1AUKXSSFYH8kCdznJRPdM0G+2zPQjmXqykdcspG5SqW9q9KK
OwNqKnmD8tFXX0zXF/Zldj50p0PrYwpppDnn/Y5/d16AQZKhouzgcfZ7Bk/FNDSC
KYPny5Xxwheyf47wsoyXX0mgIAtubCXrQAlY1z6sxM/ynjMOkqPR4GgqzPjz/wrN
kAM4yNpy1cReCInz0+gfkO9z/fCrz+g3vN34c9jW+iORgsBsD/2GQUlnlhHfcbXM
JrPiCjxibd+nCODDcHSp8AARMcxyZMf8GY+xUwEkK+xcfGhagJ1y1aKcEYjqvcuf
3Cr04fDKvoP+KOIsvAhea8pV6ZOXUkM3oOdr4zDRcheiFIzZNmbncw/GNbQH3fRC
Uexjfu5RlgHhMEuyhrgIDle3gIu17G7AeMQY+B/ZFzfJvftTc4GHlYTrLjo1eL+M
iKQr6HO6PB839JSADFc6wtHbDROttMllgRNwya/bfYcb478xRP59yXOR/ejir1Wg
x2NSUZjbkB5KU202xAOuNl6PjpyF76NpQwCADo02JvaHVYR5QwFg6NivGSLC9tHe
h89YD3OodeN67lrsVzUHHMasPdB2jKwWm5ehONc3VtEgUiqykuj7J/BM3A8zGGsa
gSxrKMKbMpNjq7BIg56dmq8zXXIq9sSETWi25HB082BV5MOTje86UVaBdkxh521A
UrBAf+awtP0UtmwMXxFCyopCvW0w4D9RLXbEKjexv5TzxDtERQRqabFMV+gC7MPH
kel/0dBnfxXVsgeN/cbMBD62gYfzvRiKHKacxQpdbF2kMWdMuS4vXxpnToCRT7OI
WlbN6ccyhaFx9DmVDg7m4WNN2VWCzUvV7sZ7DtISIvoq3aAQQKgjebyi3IJ1vRfP
GuZWzvW7LfV+NdU/xNgNz+Ku9QKu177Sp5N00E5uRXH6CSirCaIUDO7y2NmqTAhp
WBYmx0zqFs2C9Es2dPG8Cr0Bv0xE9eIzkC04KyA914UN/XhAL4zC16hm0IZiH8Lp
PCZXR+N1Txl7Vvw+Htb30BO+mv+Fc7JZx1p62aM8/nR47kKp9FuwWQjrdqcMQ8Ak
YjwSPjB9lBO49YXcoQeZEkgtZF3/dtvQ8KeqLrMBXQ+AqmbDig4v0X30LtkBRNC3
y/R5XP2O7yh4VUn3vKRpA+ubHVWhr+2s6//WVuIFb4O90B4dbcyQCPlp9jKAsz0y
9OO4l5x3m1WFg011f3s+8Dl38bwsLNyfqZB36fO6HdwOBdCRjsAMcY9WN4lunn19
i/wQGveaZTlcTnsquzm+wLh+yqrXYYgiT3RIIRtgOsmjn46d5XZbNAjg2PFFMk4G
p44w58IZ6IM4k8hd+RgBg/r6yXOKTCclipmlTCkH1L2Uaj+u/h+4GPVRBgMVZ39g
zWWghhAcjjSOgRhsm1BpLcxWVW5rgTzZMfpnbgCLrMvdny4yhJYhh8Ij9+g9/73T
Z/m4hAUdnrG5niImK8ezoWXevAIlomCjpoHimtEzi5GTgDBeCeowxbTei9bnhwiX
6RdFP0NlvwQ6F1HB2AMoDwRjo4Uo/pt+WGz+YhZuze2ngza66n+paz327IljkPXK
epKSDuIYHYuHXCeJvfXuGa8sXB5Jk3iZxLlTfKw2qwv1UB0AIM6RGjbO3r0Y32RW
IzsErPQQsNgPK6W3UK5NcDmdc1Bj9pv8TEsT+3N7t3kxVHDGAcGj+e31brce+HmN
eKfbXFwmm3xNVg6BX1GpGCAQHrnZtoXk5ImKVIz+GMys+IqGMQyxBl1l2EqYrxTi
qrRrHmrZCuvIhoJnIf3Ay4O0nVGGsT+tI+go6t10SzDztYB3S+jSVwQyj3HYV6Ii
0qNkJKirbMnRDjrunvpCYdPpx1+EAVLp1/MygeibMCz2B7WmM0Ec0UhD2TScJ8TA
H8axI5fgsQoBkJqLhbNeT8091govu9p7KiLMdqo1d18gRdXAWCPYq12UaulbeUPm
0gMmOrmw2MlulNnkvEfAg2rNMg7m0UANBzbZkzGDgbwfG47jCt+jSjP/G5p3pepr
kMUgexh4NmJ6sezlIqTBXxxcjfLe0OXJGrEyp58+34vPj5ybHUSZP+srjkpSHO5t
W6+yVqYxdc8UDy7C8HQdPNab0ILuW/odGSZqLTqfx3nL++dVTJLRtFLyqB3Tx8Y1
MIRyUcDAoIu2PPgO8nigul6KAGipio1iKnSClXMOhKAUSgLz/a4RDoHd3fwWGBmq
O6Lyvd2UWneP0COli62FuupbCG874dd+S92vbKkBwMh97VR8V11kKCf+Bfb8I8bJ
YUWJ6JvM72Hk6gqboHvyL2yYlgQMABzmz7z6cQAUeLlUInxkmtc2RvFZb0hJuQOP
WHc61/jyWsnSolc7Yen3rUJw+bo4hWEjy4oi2e8SWkb56LAxX8lanzp73U7l9LNy
iZj1KQsYM5pZaQXl7WIjSbNX4PIqFqnuiyGGV23eoME9pXIDC3/s/jV5L1mgiUoM
F2yWB3J7aVJ1mM4hiWMlVKQlzofD/nSuCqyi0QVwqmxiacgdveFCrPaONI6iQklu
sWW0sKzVCRtOhTWPrW1Pi73OUxbKNyl2J2xaZ4U27q3Gu7ep2z5Up4Om25Uk5tDR
W6NUd9ICknOUowIRaX3n8vKYDSK0DtNVdkY4hPeRYQcAxUnVkxrPXiEdsqMINsR5
a8iglFBVJ3XM3oPdgurR9p/0Tw9UQEmBeS7wrbx6VX6tLvRshJY+egPPXrIlCcV9
6/BXes3h3mh46TIeZAI3vWroj2mrJJ5TDZG2A9PjzqmCDfi6IoAkgz0FhqDnFuaX
ttzsIKna7kwIOD+OWLZTBLnhQMYU/6Dk34+2CbUcwUNvHJwNxDM3QNvxHMv848Tx
uDXC5E5V+982OcHwEfB4psbX7gj+o785CC4tLB29n/bUvvp08gxKhJ1PS/qT3ooY
gYDK5/ceh44XuPaiej8fGgnhQ5jFevg2SCweHkKdSlFojjKtWAKeEtaRbbWRlXJ7
UewYAGtlfzHq/1EcePNpsiVG/+nUX9/YMLbBE+5xW+PufM3xwwrE59w1i776RfyC
oNupm4WqRSwD2rEVv2wo9qw2LkvBAfkRTrKHpKcOqfO5cp+3Ko+7nKgKVELqRlLx
6LvnOwaf2a8VLUxM0cLJu3xVgelntU/kuxoxrWUQZNuvLAPm2ar4C/MQ24G4UeEQ
vv66Y/NPN3r7jx5bZN8Hmk2C4n3lmPcvpXkV+5VWy2ubmy5Gtyj21HoM3+kuNC+t
idWyo2N90tkAhd1O+Zy/k6otMEeXQbeOu9/itvpvfHypP2+eVh3tSY85G0b52l83
ZqeQSiWJtXtxe9fG4A9sPfaWieq2jcOO2rLcyq6lfXRnjKVK9e2mzfcWBvssvcst
GBoVp1GgAYzdAwE9rPo6oVb6SLtre+7KOSiaaXR/qWA3KJ5xFeUvL+IZChEHhSTb
LBNW0BW1pbQQEQYGo2h8asaUnJWDFA2Bxj/uPF99Dsd/nuPNuR0DuIuWvKlKpU9u
71UZKq/igKxDl0Up//xj6BzwY4UuIZtGnq1CCnC974KCq6zVYTdl8ivyDXgdGJOc
sIKCYt/9CG7R+leU6W0nUmskaNWTalT5NwvvUEZiOiMJ/UF5z+LSHFbCbvatCPMu
w4gRYPXaLbvZQNAGgexYqV2EhQ8l5b2itzpE2YXcE3vLYuuXzVcyutOvXC8dSa3h
yvrKfAYG2RJ3Qfvef4/XX78h6jcGnySTakLlWdS08zGKsSGMYirEEBw9JmruoFcy
miyaOx+01GNIbyXBt9kqPcG7L640FrU4qhSfGkw+ZqbEU8qpNhCpCeqKhzbCDzhx
2zPxQSG6n/DpWbgWB2f+0QNDf7pNzFf0dBV4uG3ZZIGgAxci9RDEsMXBt6NxpdMG
SFVdDZ8XAabSZxN07eLC2SAtS4zkWXxGZKrpDf+tnVHwDO3xoZaddl1zUp12uL7Z
7pILSpPnJoBzwFEnHOrf/WELnovkir76729TURO+DnvdwGg3UKzfsd1VJbWH4hbZ
bDRnvxkfj9k2gVVXNL9H81SK3oQuQBo7rSd0nNuUiQm8OgP6tGNdGGbV1tGdeIOX
JF/BzxHb82V3MwWYP+D1Hma+Z95hm4743vJf/E5QS0KG2g18VjNASzd/4EgD4llY
oSUbT5x238Q/XcuQQQgMlycWrA6M6BiOYABXMdGTVU1pU+NXpfS0Bbai5y4uEWYR
ugMdDhIReD89FJG4q+6r51M4+kCmSnMbAMLhHktpreiHgRnL6dqGToFeRMkBKko7
AVUvY+t10m+Gut5OaI7iyZxASNyYDkJsgFkQn/dwVbyVsr4ZEkUp4po43GtbXTCF
/iUp3FcCo1Az9Trk2oyoNrQ7QZXL1GR919co+QSo7/VdJoRcXnSZyHpsO9OZF7Gd
Pt5MYr4l09t8GltL5KDwg/iqLFrYhPlyZGtB0rWUn7eTqrhIt+5AT5oCCJh3DF2d
FZld0FuhdpTALu0zXrfddW9XJtpiOdXK4BPEWPnI4DfBpC933Fu7bSP+bzMk7N15
fJtldr+0E62v6WwhGeDWh/mHWjcjhmAms8xVBsaW5ugI99M35XtPzrvF7pmiJjvN
dIMOMHmuttx9z+rP0PPbCl6lWwA4R3GM435FMFHCwfkHSoaGxR5IK8AETcePTFoB
LMe+pFAjFX6RRivtz9fhNPinZ6X6In7Fh9lhG4a4+jO7p3Yxz02PzyinOStq1SMg
/K8j6TDTVDXKJNXFw/AuWmXqNWPzKaZfUVLQ8eU4tb39wUIOadDsIAQFifhee1ks
E8IBdaE4A1lLWs7e2Vqg/9NDOIaryDN91e9nHqop8Kiy30BnFaFqDFRr6qH4TN3T
TRBLGcRTdaZufgmW+BfuwbjrA8FdFnrtpM9KjQcjuCft4FTTr1BpsIGWuUPg/xYA
N5QY9TnJYcH5EB+ETKhuziFJvkwxhI8s9FEPTkChbaQAJG6WzZSlkPZuyebr583v
j4XWW69o0DEb+6ODsAXsa43tajsHGGORB2LMWho7olqugYH7Oyw88YPP3ouHVXnr
fBLtgoa+fqNZzACJNTLiffHx5XPXDC3932BTz0uVQT4HIeYX2NaidH0AoE2vXn5M
Co8Cdo4aJLnuhvMOFFKEncSx+to7qqR8d8ASE4dz0V+bOs9N28YqTv7kwTLDhg5q
HNyV2Dtm9dT9N3Yc/ZZUeHACBp5/J4VA612Kwzudwa7ak/0RId96EZAmojXQMdbl
QIjm/bwYfbO1FDdd03j5zXC3gerBOC/QxAgjCbVKnRAIIRBek/uKydqubRoUFyRU
dMSp9sHr0QomQoWyRSIBDIsmfaHIS+mJ0TIC0UKMWAtwNcgGsbkqeDsv+eH6q0KH
Il9zfVH/wLJPDyoGVn/OBX/Ihm5uU3ZxONboZJw5ei2mJZ6kDKjgPdGvq+594bnX
yIP6M2bYlYKqrGrQRIBqXpMajPfyUmRzJXJMDbR1BBKZKs1AxUhR7vSXWRSwSF92
rnh3lfjW6D5VfGAlJN1vMrmj1VGcKdxAFO0rHc5bkMwxrpWQgnfm/HLhMdUD5Hh1
g1jNHImK0gMUAnywoLdSCsGiuIiP2faEuGZt9QiBpH43M6B9GCfKipXKRV91eBEr
O8+10WKBrVmouW68O2AD2UDvzFXgsNtnzAdmKAAHiED/CDLvXf7HQiobF2sohfxg
Xv8iuVxbZT1LkSM1ZhfTi/rgHScUAJAU7e2laV+3QZA0A6ddfxXXkVhswqNaQYjk
UKJinL4U0OT+VyTfccO6ZmLqYATSlKJG2MuvLNwh/bRtArN37mS6yYy5O1R6QX3P
V0X+qFF/QlILX5b+CMY3hRY2q5gGUwyomFGa30H9W67L/BfWR+yJ7YuX/kb4cbJR
rTYtj+oPYMNvUqLJ+h4Y3v0bXvanidQk8nrR3J9xLI6SfEaWgVnW2ceeGMKuzYZh
Pb5/0BbLg/7DMuaHhVaB8vFc+hxaHXLW5HZUGzio1L4/m20efCIejQ7Zs8SZk1UY
03zuGcfMoT9iZPcZvfdoEwxMRfrhtel/8JmL5Y7JnYt/BdBNQ1b7VJgw2aoEeBWm
ZPgzTXVlgwZHSy3csL5NUtQWtwo/QfPru1k7EyYmxU5pqybNuedaKsX5yN0oSVuG
6owvj+bfCxPix9sCl3SnSM5gv5Bd91yZUweMFfjBfxvbQjb1fAGO7ybkbCDoL9Y6
k6dRJ9SJCYQFazZLiiHpexZAPhb/PdWBQp/XUJuP+rv7YsyGgKUqir2RliEzRALT
EydCgMsfZ9Kf3b+F0cZBpa9WHWqmMXEFX4cx8Y2gDNLZukQfAr0AdK4qadcJ0mgo
fRAJCEAAv/o+ZG5manSNYrf6Dnnx5lg5gIVFPEFBVt+IvVe23b2idZZAwuebzLLO
BN56SV9nKbaIPgBHKNunuWTBooiWjMv70tpL6jyiBc9rB5VdYt/4gLdknpTmD8XP
jgF28BWRy4Jd9Nj7Wa+mxPQsd/hcSS6goDi6v/O18aYoSpYh6H98t9tJdqTrc1VD
Vz3H8Drn/e93OIWYebyoZh9AnRer8Pp9HFZLO1xe16Opb5qjwburNlCWizLJOFSH
r6iPmqk5Ru4cR6diS6hTsoJwXsErS8VkvaJmUQ6ssvL9BaWIM3tquLR8ecxEjIZH
rDqBGY79Rhube1P0K1EW+TgFIQ7RGj9ZBCIzP0UpmBEVVYVlN6wkGSSvJINal0qu
z6MCyJBFE+InkRRh10nt/TuFPXTfSF383ZnECFcNDjD854x9xMzFHV20fB+nwzTb
1xhjXNLSIIcy28oWMue4DSiKPB+gw+lv0dizL7qZuTN++unIo/gR0oB8k51B6wBk
IArpzUxJFy15+gqXfBsCC+yVoWjoiqtooharVLZpKYXvu/LM9PeGZ6M6NZT+fOZw
Hhg08Ngl88xBpZsHfg9/707r76V6PR8xFmWO96Y4mx3tpGHXuBn3oEV3nr5OgZRz
RsJR7WHMLvtRv15xOnDU059SqnDvOZs3554ldn2nAO0BfhoqA3MS/Ga8+QqHzDSd
mPlZ2lR6KD7SN1UI0XSIuNTKnbiDsCrPfjcnq2VQGfw4XRz6jaPA3lgRe5TCKTeh
T6Vki0J+KWir5VJ06NJ8sGGXfGd+9SFGvmgo1i3IkMOiNYSOwXXuynBHU3DEK7kA
alMm6qcOh9BoIJNomY4Uk0Kc2JyLbJzo8PcOufo86xl3HI1ymiVF3bKstJaoD+YM
jluvO5ZvUz44JzaWPmtTr3wCwLjjPX/KyLFJBO4GedCMnHv0+pP2eYMBNq4BjTKT
V2jC3po8Pyn/R9o9IPC7u/BidWWFXaxzAg9KILzfF/spTwbmGgEmF2j9solfdE97
sc970nt30/xlkfPVLGjW1Zjl4PK7mhzUijq9rL2mIZDU7fsOTfsX3yBzTvKZPp5v
7BGdU6gZxkxsSAAMTMGHUXAXNXbyN2FTRRcslir5W8QaeDJq3AdbIR9dtK67N9Nn
zzcOJjfXJp2VtPP5NtINxSZ0sXQKdXlgPBCNSSqZ2wlV4IHmKaGiu49To8gQq9b/
ifsxxjUTZZYB0bc4h3hZwvW7LhPOcjrCmRPwxWEvHVq3SbK/WSSo0XY59e0Ba1cN
oYbozoOho8ySm4mCgYnudS8vYWbTR2rbaePpR3ICKIW7J4W29nHY1wvqN37cMomQ
N8DIqY0XejtGfx2EeZZtI/XefV6MLKSj/Y/OH0+mt7UUA+aAmuYwkvN6ZlAmqj2E
Pax6xMqKwmwl83koNtPW9yNq3lnIQVnwoQm8uWCvKk14cOfy8Fol/h5onk0PH5QZ
VYssQaa9K5Gph3K1Lsp3cAmA8jIYTJIGC63OB1lJFp+N/D9br1ib+B4exaTAwH+j
mVioxxRwm2p1GC3QsoYmCJyY1kkee1lja8O+3lhCRpa0rfmWL84QpeOWf5ZoZZ3s
BPbDRfmKYfxlWKy1D9ZQjedaXVmOafBQDBnAAvNCaFM+FBz6OZKVVJDgv/jQDsCT
Fe/q8HgTOa+xsKWJBo58IvJ96IBuHZ+cOL/GUe8/OKplaxFZ6AooBbcv9RNbm/1H
Noi9D1/YjbNDulvwAmypxPdtumXUKd/eBhMnDIWX+HTgTXZfjFOlc2K1xHbCndfp
n4R3m+B/qXAIhmexm8Ie1kKNs41f7URvcWLTjkE+LO7tBYRZzron2UWIJKVqpg93
PUZfC38XzpZCl+EAf0TWhPGKNKy2jaZu69g54/3Pt21c2eGNHa3tf8kzsAt3K1G6
EqF8Z/riBSNmBRcHuIbrNYlfa0q7RMN82M5tZpGZG9RfAGGuMrS/mYJPL66GaW6W
OOebAGMei5YYCozKnXoKD5IJtIJG4vtKSBHTpdwmVY7NluTmiEKF731z3/XNyAoU
TcYZA4YOyWUcYoaZAkmTggXfopvn5k6e2u4QeVQxTaGJlN0m+lmAaCqsKVXuMGxw
v9WE+f4mwhUxAgkEZTFN4Xlk2Kv21E6YufipIXt15Kf1LWxpuLDtEhTsX8uCej1C
5jgczic4Zdb4L47MFAYHC/ltnyhtyIKCd53O8jU2BKQQ0Lh1EtytbVQ211QotNuq
es15sjMeiM9EDYGzvbY95Au0vyCfoN/iWlIhTpzD41PipUu1z+uWLl/u4otO9BCM
xa7ABUH2QOyllvR+Rmf8Z0jnQwoQ33mna6CDNl/q7+Ryd6SAYiDYPa+n4K+uKOYg
FgY2BsCLRaUiqxWzNr0yWvUCz8pjKjlA0D0vZagKB/+ugrr/+kdVivtrSZt6XO0u
Jurf26de1K5ktL03Ei0NdMJD+migVPZQXPbCsgekqLAjKroCsncT1ejsYEMNroNf
HlOyZgRuficsGFUATIiTC9JUTHGGAs+NJKKz2k3WKxoFZ2ojJIf5Nf55p2BCs0kY
hsB/AfConazepfIP9pfkCeMYh5acuXV3JUbVursZP3iNQv8WF8MbJ34mO1I0xvSq
CbAIFEaaNMl7PNltAZQ3KsG4bnC62aoAP6RpxIrbFVBUyq6syoz+AIhMprOMroZB
14GsHbTr8NXUzvegucVgWlQ8Jo2m3nIDUkJ7R5zpHmyk+ZLq4ZSzkm6qlhCaGQpr
iNJzSAYMkr6icslex96tq77A4ARWny3Nrk95okkC2jDyb9uF1RgTueiSapZRTKxo
tTa12MCG22GeKabNcV/5+INbqwHtMkmXVNCic14UO3D6TBErn0sBL9VumcNkzP3f
wD48MFKwQ50sdes8iOc8iJmLcYexWXBUAX1mlrnbFwSbuOyQ31pjrVioZprtDvqR
dyejl4HnmvtAsHa+L3H4tAdmqctC+E+vVdP5oBiYzlGkmhWqehZaISI/+2qKx1jK
H5B6jHj5G0Pk3JaaSPp4MfkKxq1SqeFJM38kE5BeGed3GKbx4Y+6sLOz5YNPcpii
Kb4VngO+fzv2rlP3tvo0+Q34gIYgFdyB/cVsVsWn7uwVD5HLfa2sxg2nhVNeVzRS
gfYDjod+n403Ep1YCqt3qbdyEdjzJxJt8yIpfN1c4eEQ1vOrvsRLnx/fHSVtkQY4
TbcRgMNAV2DCB7ZuBa9lhZ8pqvwiAM3k+OaJFnibEVxWwuiH5YDPQaMvDdo4yURD
qDa3s8Lo5aBP7A90VQ7u31AAuagIC7RauOnp6x/XFPwxP2CBAc2nuj/xbruQorIL
9vyxbX6U6G3GZ64fCsEXe6auWwPqc6JiurQI0z4RKRWr14X43/Fvmh3kF4anFXS/
PfBcty/rq5yop4scK+qy79p+0OhDJbbWlUXRFuW/210Lg53D6F5plQFndLdVTMpf
+AkLBV5lNXkra+GizEQej+QjWH4eEmkN+T1pydbhIOxRglWYPrHgwyhft5qGxhjR
HGgx0/arwNnhQSOJxnAsRlkxQejeXVoPSaELYqBh6k/O4plX8HMt5IJ/sTJp0vSz
WO9e8npGBS7E/Yn4qOxpkUmc3hiooO7it64SC/deSnUYuQ7MT09iEFQ408l0gkd+
Yx69AY0qpiQ8DHS6Qwf8WmTh+N9tvSLiyWH3Wpc7jYS3XJPdFROcqdefNYiVjJyw
inG/UZRcyQD2E0VAiaMkfe1PUicUUEmlLmfsJhG5Kmy8oud0wljyBYJnzZA7py4B
1wXPfPZFHSj/vG+oqglTmcfyEOEBLKI2WbyJBx+vXYUBX30E+RUNOcj039bAfUNv
c8GFNeLlRQF0VeGjf1ddQD1Y0f+QU/I+nRxhQz+XJF4vjWCgEOF7VJLFBLEoU9IY
a01Q5o22BtHXJKEgZQHGJzSNK+BzfvREQ0oMw5F+RjHqv8dXQWbAvCDuqGYDQMfE
0hSp8i+v0H1OTL5JJCrV1BcaHWGJtVi+2lqVrrgPLX1hZuwrYJFQNT/z30ehT4En
bNqNGxCNYEq15M8RMTxZZmWutmVB0d/HqBBqAMAwhzqqUd2gbpmK2PjRRtuUsGqk
oTQK8F2PonXn/ZdnzKtXR9Nhupcr2LTFYfJ+iibgZiKM1IXgisVjmHZqNUhFLh5S
sVbaL+Wx31d2s6NtGOnjhVmoioryN2ssKz9XIYnZRYrx4GXQ89Q2SrlYw3XcDo5e
Z7aZ/tW1ACCFJk6B9ZSiLfdAYAEkV5Wzt/W0xVUEpwT8KJ2b78zu48bGk1vmPJ3B
UwWq3elowZoiteoK83NimDYT1UELy95R16YfZ5QjRJxlm6vWVHgRNuAKK32LZDgj
24PtYZ/wVlXogHC6BzJWqqAsiTA1FUGZQ3/geOiWuV9Kxmsputloax0UprqbTFjl
8kukJvGG5um5IB7kHWE7jiBXH+eU75PsN7beNzPzMdC9Gu4kyWLFppyD3espYpaf
4xJWLZ4eNUmknmP0g1b1Ru4jgUAJZ0aNF47rIVGgTX5GB7oz5ypPzNn4A30GibrV
BvctXcctyEUA51biNWfWZrd/VVLFhMus84fYhrvEVyWc76ZVrTa+BjL+PqklrGPR
C7XgcNIQbs8G9M70n/sUKkzPrLhunPKRvLtetFkdZN4lwr8v+Vz+9J0EPQsxZc5D
b5gHGmWDUu5gRvP+3zb8JThIEeE4o5GJsXagqK20mQvzeWYffDGQAHJEAjq1Z8lI
ShbZHZh9dtwi12gjeMsJe8yUUbYUgqE3VMzhyY1JsVgqsCoebMK5YycOCR8jfgPi
7gxm7M1xUa1d6sL3mADnkHmgON5371NaL+9UkFygje3ONQ1AqRYkUkS2+rzS4P8J
YPCkjsPNxtSTKzmLkj0BhYVJkPt6y+1u8B6qmDmUgiRw9HVFaHMhooqpppNJvyTY
+2EGplCBT8QosjSASRu1A8tEKWSTnVPtx1E8/vj4YCi8dXacRkarbWn8+sGBu9G+
7sAtuo+68cUv44GxxwDVANNnTEh4tkl+sJHO8xxPneJDCeHjcc3GWhKqkMn7TRB9
eJGYwECOrklk3POGmsKN2uH9Pt2P5tKZNsTPmtD2gyk2Dhzt0me61P/cz+p1nMYg
5KOygSVK1LXhBI7poXxib3Mj505yzLEL6os76MrRBdfa+hfP15OZYeLVhW5BkBe2
BxGhlNr1rx6YPkUNaa6qCyuI1jkoye/UeZbUodVJWMkj4H9yPjy6zRp42f4wo6Ds
FPbvMAdaQsKe8CKcYKTEiJNE+M7DwCJhfcA5cotWEnUSnqOL+qPUqoJF/7+OWFuE
jbZUCVA/RHFYMN533iHa5SVTqyl91HCUJJpRpvVgawoduAlzU5iy3VdAIMUunX/L
FFFSPPoj1apNjU/6HP6rZQTp2FsTooWDPAaLhVDzrkGn1GxL9pdMVlR0OLUMwGVJ
agtMXEfJYsg5TKPMJQiFHamFrK3j2dBSUNJTyItrSh70yqAFXeKIDDC9ADO3s8+j
q4jy19CUQVATsoODnCBJvdeH+lBQ1Q3GlAikYfuJZMTXhxeQwWiTEaFCXulZ4L1D
8vgwcOleDVDxF4tuKt986djDyPBjYOe4dBch6PB27By6ktRlO+uksMMVoK8d5MT8
4mRe7O1w+bpEHGsZk/e7apaELapNi1c+P6wNgXxfXRAl4KVvAZ3BLYKQlZ3PpnAX
amwf0hxYuzXIFoD1xOF0TmmlGx7ZhUZf6VDD4RLDBL6B1ey+1s78T6pTkq1wB3yr
48ow0qEdIOyVwrxAN3NxMSetyglvcj9iqw90b/IBp8w4eSsHaikFOxgjA/s08Vl9
YiduSPUhrCJLfwN2tihKD4BlR6cJINTPfD+KqWquK5AHfWGKP69XB5WhQ79iU455
k4TgpNUpr3d9vJDbcxZmVYCscH2X71BRtBj1CpJofYLp/jlUo5/l4QHVYaQuLhhX
Opv29dLO6v+tjU+Q62u05R41ZYlakELEBaYTb7N35sRACHkc8os3Rei9eEiu1HBx
gr5MsMG3W/Xbt1rWItn3rcp14iPCGrZ5x9A+qQy5onSLtYFozpHdHh4t8YSHB5pI
ntNRxCdBydH12a16VIcU9sLoALIvIbcf6sRiQlAl5Ob87ZKCpkB4gB0pbhhf7bPt
d+3gwC0YxCA/z8Rov/G1qkmRGKRgyEumoakCiLRGEFS+tErayWpIwTiwNbip447d
oqizL0J6jqXr86PesAeSvqIX5zm2MNUH2swI11AsCqj61xHzJfgWm8jM8MIHoP6F
u5D5hE5kaiQKkOqL8pq5q2OE2omYe64z0xRQ/BY+hrfpZa+VLF6zWpf6NlNItv7m
5Ylho8WbEmRFPWQZDadwPmyiDqormls0dOzWIt2bn4kKbGDbggR41BP6HNi3GLm0
dzWiN94H5zHqlpaOCPXKj0Mx/UIN5uOrLZ27iuLskfw6zbJH+WGASD7g1u0vtTnk
oIuyYL2cFlusfaR76zM1e6gGdQupEmERHXEdnv1EUq9AIS1IZbm9sJU/s0notBJe
33ipmUZXKtSjspauY+GQ2MX+URVQSuY2dD1EkavDrd2AJWpCy7SldGdM/+atK/hU
L8yUQ4cia9NYSz9Jq/xRPXQdRVCqQv65/EmiRa8U85WimYI9KljowvHhMvjiMZVu
oq1REj3/yiqVt/LTXNIVTDCKWJBhYmfcdwOMIwPXOn4C+fCA/B3acHVQNXYVGc0n
78fOuGzIhsW6IlQSdV6v7I/kmm67EOH81lS6WGmrwld9ma032H+Sr75iXn4NHD7B
0aR2aZSWRwh+mOpIquLe/LB4Fs03NAP2VUnollI6g3UiIAuSHRu+gcdUluon+sZ9
Vu9LqjPI9yU2BA8B/ZCocjqy1hkDsDB3pdg0MB97vlFtaldqmHljX4g2tJL/zp7P
7m1WhOM/PMJw9TJgIMyD9CIVGuQ7Z2dXMzlfJbsfSWQDz+Gn03jawAO5U6Nqr49x
QvVNO+HJCphXv+i3liobxa9H7hmk22/9BPOvVo0MbHMtXOTiX+HBsiDJ6DSiZorS
9XygG+vVlMgExP5zIqIhBurbAP3sttCWeLALluoWzyqrBUr6sEk8oJGw/+Cku8Fm
ZhTu1A2Hl/f9MKk+tAeQzg6saNi1d9/aKIdXxxtyzv0/Hza3i6Jk/X3o50q5YT+6
0XtsSdbJDDUNNvGDoCU6viZKprKjcNVgmzM6oIt3Nm6hsj0lKFC1SoaiOln42YPQ
BHUjjA1XMC9ghr4I8STZj3uAOJxNnZgER7MJ4uLTyPECdiTiFzN5tf5B2hSf9rj3
/UuQfKwrKjFHd+x9iCYPYSL6/WClK/AJmQOFbmhaK9l84TIH+0RimkM9owp+Qa+0
JvHgo5rubSjZ62WcNq1OZ4/SrqJwgsUHw2tBkSBUnrEojOAxv7uC3X29rrFddIzu
YKEKFz/PIh8GzsTXEfIEvZxMG/qynj07eSExBYb79ON1vinOlXQdjwHVjmhKjasw
oIX27s4NevTvybigrl4lP4g8W+b2RgH3GZjD9H2mgVikA//LoULljykiTJQ31qIV
59w19Kh3asnhDU5ASxzVNANWPAvCNRTVDl4x+NIHnRTrkgteXGprnT0Z/IzHfR0l
Ib9ncTE0cqiJ+7pwBz9n63qR32UPhr3xecpDmwaJg5oMQjt85BFpb/qPmy/7RQfR
V/aoZO4b8zesG2BZet1SZ5pBcBfh8XlqiByktzh3N+q6vhhX2VT96eYEe04lwf1N
zPAiz28ZH5l5X17wVDe8u1sXmjbKeLvbSRbUnlA3gdswFGa69uhezeTb7wOANh9H
7e6eEWiLVDe4zwnTAefQLFhF5DksDv1SRrta/bcF4LylxnFB54dY1QBVAtsMEDaw
dEDH5Ru5TJh+bF+FBF2fOqaqFqpYU8E4L36G0i1ISOI4aoJKIoBDLovoqwdokFgY
a7FV319ngigcc9yamPRQr89b8bxdKg8LIOFCBCjCmmwkNglfxtrXMHgk4E52gblB
eW5/1WKnqKGs5nWe0uMhpUqqtFHC7z3ah4kh8lF3Y0KgkIKAfN7vwX1OLvzgtA7f
yTkKeuyBXXM6VmMfhHeAxcxMXSfXWj3WpWNTl1aL85Bohg6FXZ+7t0k/rlYkCDlI
vD0s3mNZecdZY+DnjC3eaL4EE6CvoIcbki2Hnyxa8T8JvYKW2sGQnqWu8Gazua8T
UpmE94d8L/KY+Pz0XuHEhp5qyvrPhAL3cu2fAMaP95u4sVWR3M5EPIz/kY6LOTME
1mqEsGPpIrv5miCy/29BetJCgJyLQMN1sN/duYlkLdXvoDe9Fyjnmb9lEoC8oAJt
/SVi2sXqQWTMkdPFjz1Jn5zX7j+9xPNrOYvWvVY60REwrol6DsujX5nowxCgl14e
WLyz3UCWWkj0O+9BY+lYo65nd0cFpl5o2uQJukj5FOB9iX1fK3mjR17MVSOoTyWD
0qYnWnW618lo0cwPqrZo49o/wkVIrq+3Zo4uG9TtsgDX3etmaC0mn2e/DrMDBSSJ
jnX+knlgysaH7EDwSHV/yfOE9Wfz8lGPCgzlMrtEeUAZ+8PXbE/zFKvTKfmB1t5W
XwiX1vO6hA9PoyxOmds9fjHWoI1btxnYQkOupx/OLcxilblyRhpCuUU+SIjN4IqF
qztL7tEpFj1DlO2bTScnlQNfJIjmsnEoLJs0YN1n9aqwtVrg9tTjqOog7H0L7lQ8
HPe+rSA3C/xm32v+VoI4pyfiEhJ7hfRVFs3irKTyZZ7DWPX/XonLA9ABQUs0Isx1
bW2jjJL+3u2KDwxJ9dqysgsuhN0SvpRPjxuEPAuYzoFa5Lp66/RGdneE9yMsQW7L
+f+iTBEYsryXLqEvHmvdQlauDXMGVvel6A6w9Vki2v6E0hd67wuo7VgcWlFEWgo4
ZOpiA1s7vVBSnzBpFUAUntSs8aH/tuJdJbXD+Lpfv1EgomLWFT3kqSXXpyGR6/Si
9/mkcNqdx+e8y76R9+TP2e50KJ9g1US8gPIa8ZykxbPEKHDwMbm+Y6jm52SMUEGR
pUb0YcZfdM0bg+C8zUsd6d+6kYacS0j9h8L4GbTaXDx+DSFoSWBEP9xcVGqU+3sR
kc+zz9yfrxwQioTvd5WhBEhQQomOOc+/OJ6DdrsNnyra+9gxKNT1qwUjnth4R20n
96G1Wo0irPrN1Vbsa/uIUk4o3y+LPXTMfP71sJRkvTL2Lwc78S78Lq7Th4OktpvF
8d7B6f/r0jCeGfZJEA9IWfkI+5eFvjEQiFCsKVqsscWvUKqPpKucRHWD4ZQknOr8
riu/kihe6OTxUhfbD22eAbdyEpLtWrtCLEY+RrmkqZ38vDYBQkB6YUjDm2078Z98
7lCJsRW1exPO2HKaTzS/z1ZCmvSCHlLa8wNwcu0iAHFbNmRSJiWCnAvOxD/OkCpr
bsC75Rw8IRZgyVEkFjRfAkmuy47GwIf48h5kXOrkwZWk3CaD0Lw6+Gjm7rFw+Uoj
bU+mTn1KQ/ZK9FvJXWtpcRisiNAvKPXQqfHLAAxffbYniZ0U2hm8FywJo66ZGjmI
pObM5K7fO2NlDF7yGN5p/lBt7Ue0DTEt5ykzbv+25Pp1Sjr97/dqU6LVglSMEQs3
Djhy/MQmUQ4nH8P66xJYD2la5iES0H/1Vx5SWFPEzHI+0hmwX1KPki/jyCaTQ6zN
DDU0xebD6U2dLx/CKfKtu859ePi+qtH2mrxJoggZbqiwgQm+2G8swoqcjHHLOvXv
jyfkW76pXGXTCOOx4yUFg13r/hBOKJSQ83+mapBiMegpLCTuSgr3kox037M5MImh
pzOoGAropkEZIz58zydPOgLq0CIeyNtVOZbnxvmIAj27BjIcr/IgRjY3iCL+/MRl
puocvJhFa/fUGU894tRCHki6NN7g9w8mSnkeXeBmVOCEZwZPmF8sB5qErQ81kZCg
O5syQNKUvMh5ywJWOh22P9Z4mhyIOwqAYTMnGd4I4h2ij6fwrPzdONWw+30DnjeH
JwJ8XZ/lKewSQT7psw9JaGcpmGbwfMOfUMhsza/hArOhO2MbHiN5mlC8s+XDdd2D
8f6D3CN5SnFZaBAPeoTD5KooM1lzh0WSt1ugVPQT4fBFOh5L5D5Tzt60g7D7lWF6
2oly6J6eO6fo+3dG8ZYhQAnyA4/IzVMkT0fL/CJwqBb7mak+180IDIf8k4ek+prj
6mVpo9rvhu1edbTf+x9UNG6b0Lqb2PI7bF78CDsnP3l8kWhjY/16P/6Q0bOuCRrn
gj/ZxKlNAOARh3sIighHXthXHxMLnMG8LQlt5YarbJvOGJjYCXZc8WJM4/iyQCP9
Fmri9Na6m4IZHy+LWscgleDIXw+Nj14+n7zrI3ieRtDNmwnIFlpcQvuWya0xLXdr
sNYMsTe+a3QwfQm/tZDLqmGRhK7grO/E+01SlbEKh6tdnqJUmWPEO3MU53xfNoGs
kMuWOIkPrdt5JfLNGzTwSbmDyYx+wm+F3Uv+xcywabUqsgP64mU7g1oBw9bc8zOQ
pMgEHdBZuEkImNawu24ylHMB1bCrnBODlzvvKobvYER/57fdyZhtks4mqTVGvFOL
4vy/gPdsTbOpRlu1b/7g5wT0nvcuMoVLMNcfHsZOjbpyQ0zZ42FsYbDVyeN9CPI3
fkwBmN6QDKJOrurNImp4Jhdmz9QrrEMlg+1aGvf76c7i2e8FmrOhYGgw50qVjhna
qbZ35vzuvEOLxxOvpnFnVnTNrZY2ChxstgeShumg2hhCJYm+l0UK3IAl8qaTeDab
CyK5BYeoeQ11uqteFPKLIdFYmeCb1m4a1Gnb2EwOXYhVAIDg79eBCiIdpJdzYign
FMGQqDusYJKbJoGXzzHQ+Izuyzc/Y7AVhGHtRz/EGeksovhDQYFxb6fD1CApeIiS
RtDmBbcT3IM4DojdHh6ykXcfgqH0yumMIJWvsG051GcGRxZQo9tyqVFOJnPOUxmN
0z5MbXYDq8UyWfGMxUxGazJ2cSLKNOrF19DwGCLroVCbMtwGC2W5dNu8Ehk8MrEd
3KKXEfQaRubWf22KMnl0PD9mOHZBoyQLJjASFmmih5YJup9zU3jNbI5r+LoR66l+
akc/9XQI4dJAr3++TGQ/wHwufsmh3JxgWY3w+s1/+ZP+8WeRMy1MioGF2EMV34RR
3Zqd1brfdE9BFbXr8ncQLUG4IwEFvUFpyelAC2GIZeKZph13zZKWs7hQYjMFuh+1
DauIzP1axkum4+Kk6Oa2NvjGTAsF67xflCQiARMaPjYDZnxSSvGlz9MW+DqqUHev
DtZg2VU0atG8QtMfxOLafO0DfcEr+5Qy4Lp3og+ZzKa7gygjGwa+5j7wSWTWHPgK
LNUpgLiiKcThPYlm86VJTKS+kBQ781T5OZhlAjoZpuYiypusMB2RuJhm9va/szVr
pf0I3MJNg8U2f0Xn9cCBGYAdbnyB8E5GMiYP1feB3l+UY/VfUkOVIA2DE4HkQpTA
JnVDQIKZuNGL3sZY4S2RzHZB1FI8OdvvI2bPr3ieuJ0AXArwCK+HadVOp7U5rKk+
uP3109K4k1ohv7/APTms0dERl1z+ed17ut98sVosHid7W2moKtJM8UjCzTGKqIhd
7ARrwXkQNqllsUMGF6dujt7uTTxLLjiSMDdPxOBpgnjqVFi4alyH+7UqeLHmEuig
J3pdDHsLGIM0S8w7XW5D7syu4NtAOlar3nHzVDvzpM77CF55Fp0E9YEpcCln/oUx
eQdVSi6RQFHFDA12Z3Syy5GMuj1la+zKq0MS8Lb6DdM7l++0SkzIWfKSNKsgT3d3
D/dcAilirnba3jYB23io1GDIqCDbVHsKeVadcnLk4F59WXYLuQbadGWF1ghwgs9N
4lu+o8jvtLBnHKSoQU3nNG07tqy8GsNy3ZaRWvbDRNhW3Dw1MLgJ3BKR97nKMGUi
54u1VFfFCBLNBZ07jn/aaD5xLrVPn5Up31xGuAiLV6HyO/9x2i+qrtJ3mM3H0ge4
LISNx2QoQcr65KHWxt0rfh83IxNb3iJndkj3F0lhNOZAsNLKkQNPec9v25OgkCex
WjVOZnfagoJHg+Tv6H2fQ04EfgnS4658xmxqoVXRcdc25LO+s3XsGAC8zjHQkKvu
FUtPsJs4+pdl3h4Q6VNxo2hGnHCjfpnq6CQo91NVchjfEIhMkR0UoSQMiGyju3xW
iBQqq63Y7lV38SHaEcmuREtBrFYSdggtErYDgAv3HGJPL+V9cINTdVNQudb6LyyC
X2IQS3DscW3jITFbfRxDlMzaF/1BsqH41KOguXvDCP4WPVlNHwd/uWgPB1Xg0Tgi
XyrVebXb2q7n5qs94PHzUA2d2H7AYJ+LsVthdjfdhj0b0DHDdFSu+kKiA2bORFE3
tXQcFc0ZAfBNR33JA4igmwbfzMDjy/6/b+FkEPO4mbWsdnYk09XpaT/UUbaW3mRo
Syzo5ON0xEIszTe5f+vsBTPGUQ4zuzcIFAylj2qEVUpyh7w/Cq05H+8bnl2H/695
zRpA8msBRo+rtvmWZvW6uyP3PldBLhZAIaVqWoPDSx5jlV+rseefjKwozaOWu16E
4bcGvd7XSXsa195cFenZe8W5/DINwhhYubWob5flD7bnfnKasFqCpZ0a//0RWTD8
6hS/yYC6UEVTT67jfw1rKQ/X0h9eabpR4Xnvtap9KaiynPOIE5eSqrgTL+/VWgok
u0kDYMQMs82ZmihKbQGIKEcHF8nCsU3jgEBkPYckRmwH38+CEDM7/XgQ+DO5cZhU
OKXfX5XaYHYFVOKjpEFosmiioUYJT0Z9HqB0HHZfRKVtTRwYiXEzTrpn5zcZ4nkY
LQOWa3DZFNWuP485KoPpGlGwO+/p5qJ63q/Zc5/SL5mNziycg6DmF1+q3CYULwAg
/R3tCDxNj6aeLEFnjqgB9jNofjfp3Gm4rdrrms3RRbXUgK6ZAS41/XXe8skdllr8
IyE6O1g+cr6ST6Vafr95kWLaBgvm6OXoKt/cHb13jWis+cTangFFCMv8QosGcQQJ
bJnp+gysnqFFdGY5YxrkVOvRBKeTbLEzSn/X2a48SeYcB2O0MkcauecHXptzobLf
Myq06DR3L4oiYhHna7Cjp+G3IOSvCJyDsjJaTrTQ/yh/U6BbHm5wjxIJ3X0xSd1C
kShfSfMIg0YWDuwz5EiRk3l+maA869ahtlJVi4Nn6g6Wqe8eOEEHbobAJN8CaoyO
6ewJvKEYzlgVWt4sAvbewWOOrGr4rXW9chVAnJsRAFHmttj3QCQdw/lAr9K2ov2q
9SjKj/ykYmYjjWBhnbCFIodpPD0DwdjPrhvmBAVGOvSKjw5UZYtmkezqIll+S6kc
cVkgLQw7l2ZarcnZyKqTgrhkHS7oxDU+tw24/6Z88je2tKfAAWbZJSvadboOcEBc
rmudBoTP/x/dMv2l5hU7MoEmVSkkno4CMmZapfSapLHlUHcLBhDj8f1mdexP4mK6
OVWSzyt+uy+1EGmcynSP9aEdSW49Kuv2hOE78CLKKg2wa59q9thIiTpx0ZW5mQaY
FF6p2chSSkR/bpAm6aGJh2BM4jET/YpdEAJOJpR6WZq5t9Q/xBP5uVP+UJFJ12k3
k4Rkg1JfkLVZ4Hv9t22xsW5bhnIPaM9q0gdyCVVs04kOn5qnhQUf+xou4HJRU1LX
EXggNjly9TX+bkLYURVdtPRlEOEr6a4uYCcLC/yZ8Now1ZXkfTfMBj+p5w3FZ4jB
ERrhElNq2Sdk3RKyKz7Z1i9Y5sx7uiedYvZpbaVfp77pZs94VGh8hcKr3hBmMVJA
xWFYlPVm/47HL56h0WTc42qxm/HnleHr1bROCM4bMvarQuw48PKAAdTGL54Rbtx6
hdujHxwJMn3S0RmquqBrTT0S5u16ZGbDAyfj903YufSOJY8EFSbM73PtE1/EIE/P
aSPM68WS26JTeJl/z9rg87WRuEdPGkR4cse/CczhuSHNOHNhXA3YNDVCtyWH+/+3
VwmghZiehmcDJUbu2ymFJq9qi1FXJqlGyQyVf9VmF6UC1MBqvyxCvtyrCqqo8X1b
wHbjL46wfQQzACk5kulkf5/7nNFx/8cn7HGkR5280PMI7vqS1Xnz3yqPXxuTiAhU
3u6/rN7lxS7It0UOqqEGs2Zn6JPKeetNj+aiPnH6/h3G3JF/IBRbntKyplKPxjjL
c3H9IVAP/+JKNqAoqHdmZ4UjLC7Q+L7xGPgfNMshwmR4SqZbv1nY3cmzKo5lfxVP
N2BN/amQ6e1nWo9aZz4MmGMO9owFzY4z/pJ+NSe624kxYhllqVql2x+tjPwB6Xir
o71g6gagaSTOXBYzDxtDUD/pli6jgyMpWK4ztltn8m51v/HOA/g3otpI5FCAEzPr
ttyS95fvjyPNJ9lDY3U8zN/qTgNiJzZgVyq8AskFYUJ+rJiMUSjILvsERXAhrjil
WY+omz0rpJMrnypQTmvCzbHeY9TvQjNcLlk48W5stSNkvUV7MVL1nzPHgMucfREO
sEpan97xacUbRCxg4QvAD4e7Oz9QvvLS8taqJoB0ltAzUqN+EBUMoiLCl1lGJa19
lKmLKVlyauD1XDTU3Bmyu9e7YLmhLK1Fun3qNynLAQiwytQGb599UOPeTXCFywAh
BWvtX49Yi2evztJHrPoixpKQmyP1QEjQ7Q3ewgccTiLkcd8eiga1lpndbNerdJNd
pYedmX91AgmJBst7SYiJAmjMv9IY68fVP0HirwuSi3FUuISSzQyp992H91lotzFX
UOHxb2x+pPW5a6IozzEyEi/uKskz0OQPN8tyDy/RXeGaOb2tki1zr/OWAEnGYJd2
GjYDESnPhM8bv2BRqipEfl66YkQJhg4LgnIAVYHrOS2aiZfmQnD0uB2ROPQXwgF/
lZqACnrTNuFJVY9NSEm8a9HjwKQrGZNeLr1LfAiFyBUo8wQnh8rdmXSirnDUwRws
reRa6CyoFCBZXJPxEGKOSEM04hhjX9Qu3eu7hhHWtggrROUH68khqhqbQRnxb0ui
MO7lRBrp9TXsV/oxDPNhEu8J4cbQ0t+50ECS9DwaaAMe0UOhnckIXNs6PPYHYbIl
YFZQquHrLWVo3VLn8LWJNL33q5lBqssjax6W8j9oNVxcy7IB9cvQH9wW0j4G3NIj
vCcHzrctOqXnyPsf8lRnk6K0Xn2Wb7XYl6IboiDNliNJ0b05qzttCsIFZwjXve+D
SVyRRf3N9QrsXGSSoHTPolE5eZzvgDCuH2qsP2e2ckhxhH9j+KauAEcDVI8Oprr6
AVezsUUSaarnV2/U6wHN7zGa0fQZXlkjknIEbw48P7jGKLeId3MVwdxq9brdWnNX
C98j3jWrV7fnraBlui2A2/u9ov4UK6QuySI3qm8VXdULkgNjXpWDH/dZ6emmJo0Y
HWruzTLw20RdOAwbPLTZ2IjTgjzjVi3sC8z9GGRFxs5qBAym5KLzKlLG6CDCju4n
q7+FqiyIl4APZnynX6M1JhTT2SnnLreqY7tuI7pQUWQuFFWkEvx6kuefvfmbpoZN
zkTsUgQQwHmlGJUaXcu6ZoFnprKFhhutmVwGu3muIcjHky64VIhaDsmqrL53PdTT
7IoWoCBvZB6fgvVmPRcE7Kyf+Oca4JwdfC6b5za16rAEHCCWMvkqo4iZ1pAzxuv2
sPlvCGmx5Mtp6ycTiGVHxkVT7TB5pIKQRctjN+WKL3Bt4sVp8bY8xYNfR5E6QjNp
o8buhOrFUvo/yAVh/1d/eQMegXMZSx4FikSLcmfBRvGZiLYJpyXcCrXH5zf1t15x
9WwmxDwTHynoZ9Lu1InAhtPVe562JiW5wl79TOwtJ/35WO7up4Tqv0lqwff1q5n5
FB4muWXY3+h2drbflKVI0YERm0T85+gDPbrxzIC757tZVNSR2oOEmle4gjmhC1mZ
W1zQk3EKFHI96rSmSD0QvE6dTrvo96n6CHBe1hcbAsWF714BMTDOhK3P06LokFVB
CZCmwYCg21QkW4Uw3iNq/Bu2EvXLX3UIVwZiB6ubmLX6r3QvdnmJMUjRF8KWLgJn
m8QN4vpTzv3Vf1gBYLjLOGY+bCqSu4UN2/HIsPsEvEr23aeivH0QD9767IjXpsZc
Bvo9zjz5OWq8kKXARjNQn3HEHgQl/QDh+50E65CyTr+qHKCI4kqetBw8S3Y4qGTS
NZFZEBDMxRGLGYzp12WeQE48WY+AxsBY/D8N4AmW3xFQeKkCuZ3eoU/anD5+jvJj
euTZq7m4ufkmaAGJfUh5aeR/CtJQOZPjMswt4uLai+weiC9HD7Y1HkZv/J8bjNZf
gaMkfBhJgK87vVMp7IJumo9huzF46yfiPV5WAsLyixYnToHpJJQKRriIio0371MQ
nrd8QkI7tyXTo7yslytbVFJoWq+0EfYNlyhU5aU4AzXAMZAZTL+FEnCulz5q5PEn
ogEI6TjG6Y5iwx+kt5wRpL24CXrjId7uJVpquTGr2q5LKVUdBMK+AJxbT3oS4jIr
WtbrmZbdk2L9WSbcZGSDoCyPJImm3Tl5XZEnZVoT3LCSBlZ2Rc8Xb+mh75n43MNw
TCz9sLFudYHBEUAHlY8FxkbKKcXJKFSZClC/lsYtfoTVLvaB03DJaSeuHeh35BM8
x6uHoFCxwJiKLxB3uZxL6dhAdAwgkvyiPXG3Wp2uwzxxLx3nAAqUg8el+HXYA8Av
ZA8iTmo8mlO/ZD0PA9vRfmNXMa+rK2f7ELGbvtaKoOG+AKru+31w9JTZb9OT5ZP9
sS1tg6E4qTx/cd0/qqMGa5CGeZnWeH5gtOj/FzbToeV+2G9Fyli3AWfY+1kPx1j4
jPK5KyGQR5KSp2Eh6lbzrQwZ8qnbz397zmF8BCIFdI051ePDNMUe7LaQciRsUaVY
oi1nTmnjdG9/kAfzmEuWah6ZctOGjh6xCPX9cQbHiHhQfx/AuZwKpmlXeviAzujJ
/zQAFJMJ+DIODb4I8pq4mqSU9ITZVH9MgPGDWdFtCqtRb96h1yJux5twLlOync7B
kmgwrRmaJinuDb5erC+Kx01R1wTCQLO/lW1peDcRqxYSaxw12UfYd2AEsMiejaeq
WU9TTi2yebWjxb0rqQreOrT0SzGTjwErDYI1YH+dq/2QQkAJKD8eXmML8jnFiK7p
TTB4+c+UYTbdfs/OoHQkxLaMiZH+aNmiDAJD2pkk3O9AxvDlmYCY3clumNHklX+c
DQ9B7UtK2/2ytuohYsden87dxL1uj3xAbXzH+zXuvCZcQzJ7YgSBVogO420eiTFS
lsSfBVINC8pshp3JJ7mBVFciwMML+p6323MJlR7WLhpCvh5u9gE6He729x+qnEQJ
2YE3G2i8T0+mBY09t8a/DgkQS1nk4yaqvMvQi395rVd6R3UJ02DIaNvyWLeU4bUr
lwIravxug/DYJuc3ONX6vc9ELxvrn22TodiS/5RSz+Q6dp126GCPqzsbTRgoSQGK
jC8klXAb4LrEbW/3lioX9F+GPjqHvruFPfLMEDkr2dzf+dS53BjyDcvtKF+TfsrD
ZFpanoeMw8pH9+AlKjX0m3HpKVMTPzBkkH+ICgCOmqZobQB7lC5C26vv/8H4neYD
ONZTHjaHDdMJRT/4L8NVoQUT5SrqTUjwtwMc/Zs+gGkytVQZJLlD1h9IKxQDvX6/
AEXwy1EEk17f5XAtOIxx3On4ScouFM6Wg7ar+3SyMmiQz/wbGOw9fyJPB0RbCw04
CvpuMoxwIqxVT/beIUFjxkpCqMaaPWgeuKuDeVXCk6Ba5q17IIH3BUAOxgUHu83f
nzu8NGLmpO2SUnRkZVnKa9jl/fB9IIr+PntHjPqq4FxUFFj+eyInt+zxCQVGUGUL
yn1BnEaSvz2mzD+UPOwspoEJGFeBcID9NTSde/6I5wLNG62XpGdkll4Sx5D8LFmR
072DFH5Z6wIajorU5FzS/GgVdweEyDrbWEpxlWjj5LppoI1WhKG66A0PlwLaxSuz
bfLm8ecnY6dwgfvhySjNY76T5g/6lYw3S4oCa8jK8TbraEkNZAm0ADz4bZXuaUDK
IOwIIZORRzkptzBf1LPF4cro1Cbfzs2ZhSrGOR6X4WPloB4XKcIqSDP4D3TBBsZu
Mie10ByWNB+kwO/RFkysO4jl4tsBmrQay48RhA/+M5PF8c4U8rl+YBwCM7RyDhE7
GSeOdsP+d0I7QKPlYRIK/Mz9D0lo9ZGFpj+gfbqjONSgPau4ZkNLJSIQ85yFt2CU
kSC6Tf8UI3rLO+taIDszORaVW/thDbOpZ+WT+5N98xLbXNy40y4uTxMYe5MS1cS8
PjsUkw3KkcMN4dzWylGgFSmgPIuUYFrCiopbWNTxg3ZIhyX6fK6yB88mPDqylu6S
FL/udzh54fUBawBoJm3XxAcf763BgVE0G7rup4NnyPZdFo8JqZuxDzayhvWtY9UC
FDB+m5DygNhMTnzHS+PEmqD4b1aAlA7tUiBSK43R+/UC6JFn6k2E3Ht8+uy++JRq
v4Q1UpoPzutZtY8KMHXFmojHe2vvFC6XIAUB4/mlgmzfD5lXJx7+ZNBq8AkX45LC
RefclajWkqNK6unxNu5jS/ySwcfy2tIOmJXeoF6zDpCskvXUO8kmLLU1gFgdHowm
uD4zeqsv1l+6WBf+C6nFpKbrOXbnTDtdvZdMWqaI1D9BAPzo4g/a+IVhuxOjoe/T
LcYTkupv60ldAKG0nQtHpnePKdNu15YEIUCaHEa6o6EbxEWrTgbBgttg6VrBKtxJ
gicwrlBn8uZtp7pF3IU0gNBMyB2NXSWrBIxfTBpv/KYXH8ReRadl7lj1eF4Eos14
uvpAsSP33wYvhiezzobvea0HpW9QUiWrjzoroXZO0MCWdfM4YimKfW6s1m7nSAgX
BROQqRDEBN9aVvQLGhgrMCMZ8QaoOe03mw/Wr1xDO6oxBnqnrpOOuQwkoo2mBIYH
jAt2IDMUFy7Yo02ksjSgpnd45afaQ0MtE2xWxRjciD5TiEazvej3/lUoLaNKxmpa
wrejwyxb4/KduVCD9bUv3CZ5SXFvjuFHdIsmEDu2i3sD8I7Ch6ZGg90FjxibLAh8
41mfDL5ahammm6jBDU4XFeAPRffSI9+o4LikVsZn4djACxZUJFACncJtYVieAy1/
Xe1h/weUcB0mTk/FfNktFDXmmJaMp8R4tTZJZlnfktX+rNQLoUm/OpJ+5XtdbxhI
WymnJvZuxNs8+RcM5owDN3N1tnMrdYgYAzIWsyudcK+dSbTx8RNnCaj7Ci98JRuN
vuzgr+CBpml6LYLC7Rns+vH2S8WfFB1avyijS+IhzfuJM3QPz7zMuJHb6fh6OQmk
ELWBmn5Yly0FPKIEg+JNqkn/Qx05qYJHZqoFUvJ4iOxevaNXU2KnVfkPFUwwGhDv
s09hNAnuis7xos+NIvWoqGah4z0ArZ+lUNupSUSqiF5yxMT2tJJKKkYxkJklkCZL
IrH2QbARR82hdO+2mk0FlN7t4zBWK4bMYr38jMyD+7XGBChlfTfv8uPmS8gPtNag
z8J/OUSBvV7b6aSWvEQs4NO+kssA9ZSvByTBQuWZdsFRLv5M7E7cAK5cIOeY1HGC
jwCLQEwhqoiP9zDAY5mW8uJy3aesfbzudRvuf7z42XNriwX0R7zLKcm462nriQG+
zndadzimZPR62lOvYgYLUOhsiNeDzGoccXYUuXZrCPyvFRYQj+gOpTbRP4w8N5qa
MkTxS75xv5DpYshzQ0mVdFWkUph1xzkobPX0kWa+hsq/ejpHKTXlm6jSvRjSqpC/
8uQMc+aeOWqUbw1xe+mppGNI1hn3Kdi1VH+bkxvfs0MAyg+TL6Wpk/NGZsRvS2Xr
pC0BTCWXBK0jGGFltcbbd8iGS/TXCfxVThqHDlbrXAEGWiDupHVYv/RiM0PoCCGa
eymfk5RFjgWYfCb/Eh0RAtqhumlwR4w/QtX+GDGuX1oI+f3TuX422mtIKhLdZkVm
VbvtytkCRPVZgYlLwYD+YlWN54ky+5Gba0qRHyK6tqgV90sUJq4Z94mMxwb1zle0
GoevKU26fe6/wFnEkcDbqFk42sttcy6lcPElSrlNRQuTbxqX6T5oAOAkUYaMhwN+
xT9gXoI9LKkbUjd8JhyM4hAW+F7kb60jBxm0mYMUPGWAuqZW0sEPFJsk7UFjbO/u
IRyAw9RTg2WRR1rdH//aZcf7fmMPL31m5odM6SRCOuBckLDbiGJ0b+6MA8Dlt9md
xF6g5IvWl3Va9sBWmYYdRjC4wKxNVIXIdGJh4+e+eOGyT9v5O6rkk0EZlhLnJtCl
QcRFUodLp9T2U9F7uyo6/s4hzPrjvMaoXrEkrTjeUV7JxDkqxObcsfM3UYhl3X4b
J6PbP3OagcLzfH3E+IURdWj3EBphAxPkOE8ajNaqyd2HqXPXjayhHdPJGMy0G9bB
ZSuuFFGlN89aV7cJDYLidom3ENwYTm7aBLkfPQAvKiOsHb7Dels8AXveYFJ7zmdj
jbfazUc/hWuPajC5Gvcqi9BmtOEiQEI+S8DcFgtlRa4jUB8k8lvrHusohJo2uo4s
+YCDdcFdgQtwAOv23s/xGBXwAjpORd1+M98iywjpynx5G7EyQJOZHOQ3O0uT1Oon
c9Atseh7s3nELMNr8ylOMMn3BmXFbr4rMfS2TUkA9mmExBuw0cFqmEWE4Uw5WUgc
oNsGU0y5zj0PHjN+pbk8C9+ThcD2clMMcrl3NxfDF1DnrK5BGwFw5nczYW4kLkBC
RQq1p8CdPUJu+3I4bijOdVy9wNhZgmCPSQawZxmncPAxLgoe0JEyQ/POTFpo/X0s
WaBIrm7RPUmQEqMqcGEGASzXWHKPlIt9xmOg96VM+4tEBJLn5aLV8bXUXb0/ixxx
+JmwDzq7yVgwe3f9nf4UY8EHdN7jlSZga0Uw4M8+ur8IVbIHFRtYcDCQcnqC6QPS
2mfPn96kQkCOnFoNwRTp3mEQ9SdbyGSrlTYwdMa6di8OMTboDHaY16O4Az16P2gh
syTM5vHQZLoJk4nOWNYSKDFSivER/bz4BnKo2ILvZQ7RKwUX+svSJWGxAcVrRhr5
hmnAl0G/iICDrTdmiaV8/4po+nQfhO70M4UCo6fJ4m95uzjcEfG7gL+mkvwECuvW
sMf9OL5BhzNEuO+iGJj0y95cyvpFHi5+Hu+IGF9uD96l4MXhXm9p6nlv/oh42C3u
TwrHCQ0ntPYzVNUmOuzNXtk4Mr5DsdAORlDnuwJpr5akRctx7v6g7p4KR5gmUIqX
QESyLrXbDhYwdkl/gTn9G4lBfJ+v3KUQ+k0ZXqHdbnFypa5TlzrLAdjIPNWAtaL4
QYqs2w9S98nF+CH6kP3zepccNN8RCfkJP09qsndG4yokrVCXWYYWr5/MuFEUSHZU
E/8RmwiiMQWjZd4aFOUoMcYCqP9XNHURGUr5I4LYbW+TrAzukA70RiJVD2JAd+1a
XXDbydYXuOdMaxM90pJumyahGXiPLZWEDesgheLhJ7FbsnZsw2OOHyA3Jgspf3fO
oeY6Aj4l/6sFIQ5PB6P8KbCKo2Kd50hu/1Gly1W0ESlrcX9v73KzQs0rzbkW0Slw
/pTzXofDNUNUnCC39ksQH8sRU3eLfPXDWAiSh5i/ucFRLPr4QSqqqv6oceJKVeWZ
bycwMTZnbdT5V2y57uxxZNVNz2KVBWRaIVQ1M3LANEEt94e3H2eicN4AV0nVTO0Q
SKzuLIhyIf77naQpQnHo8W58EsoGJBPj636YwxS4q4nwgXT8EAw5HexIMaPH5I4A
EjEcMhYQaxbd5/CKRq5vXdOg+vi8AJL1WYbtIUoa1AO6BnCIdxcgx9fnjXExb1JR
mSYUOQBJW/+HJt+4DzzoCCUQariV/Huy+tdeNJIzuM76y7NGFiuORessIBz1Sfyd
osQOISEQG71IPwi7sxw/OXca0IS4VFwdJgC0mrSQp43DLPuP3aHwXF6/7hNmUVL0
OghHzuwxPZrA462Gf7bhuyT1eiVcldgsJgWJsNdCvQrgMlAAPkWnpvj/mXEwbxIG
9w2gBt6hjxe4R0uiIGkzQuPdeGGZCeYA2aBNtbQ+AjgzwknrIkWspKvl0MssKrCJ
qyvHK3JgQiIjdPaXczPvc90+VMxz+gTzo+Bm5KMeu3jvThNI1xCedXCJKPWEQ4qd
iueFAgp+1gYrXXlZm8EWYZvi3yJbIZwpuddYZMhH0lA+LB7vbovE7u5d4P+spEDg
uX06a5PejgGhFkDca++DLZgLNPzOewRJCfKnvHcyssiVNN9iW2pnfSnULqvLIY4R
T8I90CtZQuA8fkQOBvcH4G+IvJG98Qomj//Kmmsx2RMVvj/cw8DYtKAJNyaoe4h5
C+MpOTYWdWvfQACg+FT5I+y5AuzFNXPVAoiPFv6MaRCxSKwWVNv2Tiyn/TpRMjRV
Kf9MNnC6Ebn5QlIMXA/kDA9cu4qxePXWMdlvS5sGiv9HzfUeUOB2KO5RStb0X98S
exOuB39QS4QA4o8jYrH4pFulae5lTQMG56eHLGzHOLYkEEHfV0LyUwn4Vc5hbp9R
oVoBcqLhd8k1IucNDBrXXYbOMmD93QmiABQOaNgVSl/ZtOiRR3rL/Z/lmRKrmxSt
KdwN0TXJo8slw7NmSLITwV0jJiqORF+4xg73nR78A0Gjs46eHDVzvejUAQccs8Bd
dWHIeia7e4jEqldhxwmdX+kgLC7Utlv+fYtsJp3RAmy4039DGJQ8KIW2GmZfbpJZ
MokjyH+BvJ6taR0Acq/9wLAsFGKa6YoWH/VLkzCj65EXZgH0NJtMMltof21yDIot
6YTRQygm4U1/hnFHs7/adoUNIHfkXJJOe8qTCI7amFSrx/w859l4YVmOur0b0xOH
s9GAsPn0xH+72vwRoO3/o6YKP232D/MR3YpilvBrtqyuXk/urSsyVuP8IhHq+cXu
Yc6Ab5XOn4elkWOZWWT7ehKczIzbQkmuZ6kn4qHzfs9/5pKmf8itroWaoh9WpjwU
lr6ELqgSOFBy5ztdbfzvlAtLwPs9uEUbNDT04++SrPmEajVpAIiAajH7UIfSW8qZ
LANZEn0NnMrGCZ/dLHwQxJ8iq3LwR/heFs/FgQJrKB6X9UMxGdQa7YojuXP/JTFR
PWXgfxgzBPezg4pfCkfY5duMbazh26A2Pt/c0xigSXH7dtqRD6l2GndssMWKBU3B
GZdmQSRtZI4UOjumZQIwtkZxuMJhEmH9RBQPyOdt0hE49uCB2oU7A9KavDjRugnu
vHPKzIZvSBwKdBf13zVTPqV+FDL09F8uHbmv6AgPWD+RhFl5yc1n029Vq974RIQ4
RQH21oCVTPfoA5yoWIIoi4+23A6Jx7+r6mF9Uhqo71RQefc+qVbI2696nxVywssF
O2zTqiaC+EELsjA8l2GmODW/V4/hIWsbOeO5gBQWMHZGbHFm9yRvSSNNyiNIDjEj
kuZbiQJQkHngjrxYbUx2DR3FIkGbzbh+ujLMkJUEgh49I37noABoselcTKfeikYb
XW4pSMlREld7TDAe/zF1WuaxVNsoROY0MzXBICaVJ6fDK/BJUQlECELuPZjkWvHh
tu0SuMqSqwTuNlI2ihxgDoQJgM5DpXPnMHutLqagnhA/iqZFA6akP52uE3EiPDlo
cciN+ZREeYst5iK2esqFbRQpPpBIO3PTHJtATklpyT3lFzf9tMWASesF+0Tlpwp2
ji7sXvE3N3lorIpeghOJZXXk5Xk3+IuYBxhKeJmQM0WwfgYDRpbhmpCzpdq9fbae
OFPzM3Wxt8aZSNArZzdSS003QvwJmMhyzYR1Eaq8FKMOkWGA8hOhTxAYRhzpzxHw
ahdjzKl75a5BXQm3APXcYlhXUAlR3Jqa85Ezoymoz6+RrCeeY77DHTNWmKv8H+0G
L/PGmkpZ9LbwjWPgnu2oNXi+iECLZyKvIWXLx8nW2zhe6i58LgMJpjqu9x+XY0LD
HQUvTkKI+mbf1iirEJZhMnqbzIo5hz7UVIKpuS36PbsbO5GAbO6LbktYYS3lrniQ
1sY6+fIFru88hjej9u7fjebmU6Lvsx8hqQ8xR+4LtwjM8yOgQEPJVrQcU8rdwmia
yonBCMWIOjzLTI1Zs9pvfY/xw2had1szrancTXUw6HhUsU8urmdy+gtimZzjS5Ak
kcRkwNfYGe1wMi6598azWRR+OOmRV9c3OTrMUbb6rqKbe4gV02AHITKf6Ft8Velq
FdmIzPgWVrDM51WjtkJp/1qaY8NkQXtX7KdNx7G5prdkJwpKpUwRh113RlwtbE8L
QlsVZpn1EsoEBuqbg5D/9aPLyWodJdMlV2qcMSUW7Z32OIMXA3NPiwJO0Jw6CUrs
638/Jj4wrvyikRym8Ztr7csCibHQDXtQoQqavI2maaDy9cD+sgaSOct66ncaaahn
Tst1RCH2dF0DWH5LyvLuDH9mQID6PetE8aWftKeN/esvU0RtdCFkjVnQSf63DP/3
Nnhz8M5R73Swq7VNa0/uvOuwr0jKUKHas4O/ud2tpgi1QCVOXkvPCj4Nw2RooxCs
1H9F8ZyEYt5Bj3R8D/C6bNWPyXRfzLgSzm4Qb34m+MGPQ1jHL4MiUNEUO/ZM78JV
SSoUZ+BojOXmTeqvEsW8z5/d4DiwI1LJQWrq0oDdEN68jmyCSFMmBEaCDbIkwzZK
L40pm6Y+EXuS3EouOku2xeq1BE5wo7LP1NohhIM1U5dW5mgvKUKTMo8WjAbaeLno
FJOqFbgLUQ1+zmbXIxBoSd2VpXWbTevaRuuEpS4TKopKTo51irbnG87/T4u0PpFE
4bGHgCb9j1BPhCf7PUolbJ0pwySlJ5MVPhZZxh4rhj38bRC3aS/5CV5tPqsxMnur
4aN/pgTIzIt4IEWMwUujIZUN1cItLLeZFZoXI0VkLXMYCxpK2eebDI2dlwmD+hLr
oA+BYUn1QaVeQlcoZhpwT+87IGHZtxR9qBYymEGsAOrj+yzmWfQcbYMdAW0Lyc//
wIyZlO8lWXW5uxNky/aBc30EjDesshPw0/2kwG3vu2asGP+ARadl2htgNc5gB2b3
gamIo/sa7PHKFNLUnkbx+1A3B+0pZHju98wrN5mR1e1PT0ZtPd04sMTYax/ZBAiP
klEVYkyJQy0lIeVrtNRcE/Q1jRysohheWfWMEamLFR3VSu90DWoYAILt/iPKRZ7v
UwU6jnozXQppQebH+fnsMlnISmjnQjL4auS/Poy5VHRnsnhj//2u9L1Pv7M539bY
8L1qNcvTEQqKqAy83o8jo7zTcxJs17DJ3LDjoFoG98y2cXpOG0oUcB6S4xy9kmLy
aAl7884guVY1bKx32loxqeMTj0zpYsmTEOnIpKqqHXpmwBg2JIFKt2wYkxqK+JWh
ZEX/Ourdu77HJ4kaFu6ZKHcoFLrCT2DkMC8YW1QCCXLHxsqA8KPS6VpwvkBr00HJ
V7tWuaFbDYC8hb1VImNAkx34fzzW7eSWMPBpyXE3b5tWW+yH2vO9CQZgwZf/Kxyx
Fz+VbNce1VDFjuhip39P38skdA3H4AkpKEwd0ZML6baVTEu0i2toGyHhRcz2vU0E
XODmSqWvT+ZQ4EPLGT2jxTqNa2SjZ5HLtCDLkJn+u5bvAdQh6UwwJItyv8s+fKqH
DPt8IWakNVivBMomAIPiYEj01Kdc+ymb/t+Qkr6WOb/zWgKxedyzjH8GDBluM1Ga
rhSvV4e7dTp0FLoiW430GSJUj34ausDTT4X5TInpZKYD5vuR/RHJDx8/aExptkwj
KjQjZ0fYnSC9s1eoYgKoRwuP5t5qXk8zo/QNaNqB7oyNO0NQ1gqwAcXHFhlUt+2r
PcgP3yZymsDhKb7GhdxUzSidyjrxCCZroRy+FigeGvnOr4C7v451kAP6TyxVtJK1
S5ACC1DeY2mcdQpK3gpGFvNi+PXHGFDQ2xvOTFCwY3i3W4tiNobwt9BXRZ9qKj30
6iNB+2MNxCWFduMvl7ovyPPTX8r0VmggbEG1gLb1HKKky9EEGn6IATyehb1QOYve
czUHKmCxQ+QhcOTPC7J2d84APiK7m+b3iqidUtLLdnNrE0FgqaMfGS97enjRqyBN
y7D4j3X+vecvlLoSOSmEvp/s5fuiRT6jXLMGY6520rPTtgE+c+12p1Gkce3FSnAb
vcSSYv9d9EpxUNxWH/T6b6EHVP5Ej19gUR0aJv6tP68j3wKtQGKsfpu/fGV1518Y
VZRU3opN9UR2OMCLK+6MPhlZdMKre9B4j6/msEfixhuXeDLoh46Wp4T6hJEXFMN5
UsjsizSbJl12NeVii9FvGitmo7bADIkDY0GjIeqNNA7XqxnIqeqbjIFXTRJxEnSK
vYE+3Bzq3oig/i1fUCJueMr5z4o4uKA0sS++Y6wfUsbl0WY3eRQPAxCwzqnROCzE
7EZ/6Lkpn0X3pXsLVXLH5D8frjan+5CISz2hzfEzCRnZAg1+Zuhi7IwnHwte9mD8
5bXp89xbb6wCwa0mgNhCszSKUH344LramBo9yCwjd0LqbAq7qpHyV5cUWn1ZLTWA
Zuj9JCpPN/BxoMjNmUO9aNvh025I35SMj1TEe/uIyI5BPr6zooO+sx9TG9XMmArG
8EFFdi9NyXAUHXCzaMzpYP1Khr/t+Bs1FKk0OSkZbd0Hwa/74qtluBhX4hiZMgwE
cp6M36QVaENVin9vhEcoOd3pNXeRk1EQaPzs4gaHAtn7F+uzeTd4HkjEf2Q8oRNH
Hyz6UJaag8l6q8RNS4c1NV9rEoNHI0RhBe2nOFmd3cf2mMuZ9A/7mjs6+VUXKFwp
PmMHgD5V9ZAS1oI0TOgsrjxZLI2kNn22SYwCoeX1LQPozlxQz8VFkCdhjVpu2c7M
Tn+AuoPJex8HDOQv8YGrD2yk4px7CekHAQ+8ES0FARBo9ExARnXXKU6rAzUJOYTW
2M6CvomvFiYWYZGBvzbrh6nytV84wNzm83rwKZJ/v9lDxypntQI2JA8SkmxJY7+G
bFZ6pbLDFZxwZ8bGOlWCg5VmuQCPP2G0oRRV/ToAVRK1wanclU60x9Sk/8fAfIkt
HjOS6yIkXUPcvCdPlqnyrpCIevy/0awTEzQRQKHYhoJSH8VSMNi5Iz9VHL2ggiWC
h9drQ3yS7LpblbUC39mMVGeiB9ZnX1ub5oAjetaY0tQq2P3nopqdaEL5wK1cPjli
mRa8SKrB8iCJbHaBun9EniVWvDZnTJNORfUqeWkK86JofHpiis3n2JgufBtmf6da
jPyutdF6r7dm3o7CuVa1sCiCY4yi2ekvEtdJV6sit0QrFjeFoeGlzqdmX0V7a4JJ
Yegpx3QbUB6UV2PGY+v6f66qxgBsENclOi6OxRaYf9UZXsL2G8C4+wIcNKbTSTwz
Dh3ihm71VHRME8QrVp/QeQl5xyURv7HTdVmLvJq58IvunK61EHVgcTfnPpPdzUH2
GlA9KSvCEY6l3mNgA1clS12WN1MIh6YYLre6RzKwy71M1jSZf4OKaM60cmIRR18g
VO4XKlPhA/Hwp1YE17HPpGtRzN30K3rnF0kpnWoNDM3EDtR4wKuNy9FMnoscadiL
2ysH8wQFskklDwHifytdx55Ny0ZgY+ki6aQy2jQzJAK5T7fpfcNw8EJy3Uif/WYV
doDziylLDnqpXp1+xp6f4BhOpLHi06/BeKEvkoh/CUlYjJsNXqvrNspgxmND5aGG
ffIJC1VofV057kAGce1NKf14S3DIZv/Y3yWAg8AWleMVJjmT9RdJ4WMT6tuY00+o
ifSbaM2tJN2zamnkPE2qxpn4CC/MI1CJkqF6EpeNSywzPB19x1VhSNyMPoFwNQ+1
JXiu0X1CvoHktaUP+3/LXTqkH3tCUmSvRZbIZf1jRxw6mc8AdqQ7xNlF/AsTiKLh
kwhxqqOxGaRUO0GI+sHKMEZFzXMTdAJBKLhIF7L1E7TlyW+x+8xEy4jo7wiY+IKC
ZNH1Ji11zQIjP1R+Uz0YtqqlHK2q8xXGY9I7gZd6LnJdXsA4R3ZsD6eXHHREVWea
7arVyb4M14gb+INrXlJ13bTYkPVcc9PksrCI9judkkHI1PsH5IltulGUV/BEiRnD
WkohfiUJiERM8QN/7gUejjbvQo/7VVWBGvy3Bti27Obf8qfP5o8b8ZYNkbhd+B+w
/+vOCpay79/itSgxamfKJQuYbspiy/bjXasCwJnUq85VXBKPn1aBjrIHEJ1CbI3K
N33N3PpwSt+uuTCn54L2POYH0w2ACUlEk8WZ9PgF9+CgM/TYhOXmChPFviR7v+dH
N5DSp4Iy9HTQgdGR6k6sfcZzpNwZASOAqhov/DAm3y8tqozYibdDen9qxOymzcMw
4AWz3wmmYLMfyFBhSSVzZFLd45MFoYttTDRE1I7BcTU8HHfRh4UH2tl8Y8s3Cx9P
7Z0ey15O+xOqDJZmjCnrRI4dDTabYOf1Rm6EZq8xdyxX2mtLHLoK3B5osUcvR7pe
uo8LpSlDh3f12FoJPZemRvK0HxPBk3priee8ZlwigwLTacP6ShbbeSeDx0YaaB/t
Kx8K3lPYme0CZp/K819mJ8slVojCYrL4pirFiwjNNpGExuS4PIt1TzQceq556LTA
IDySdV8pZmWX6ssoY6JgQ3+Ss2DhoZQn/B81e3hlGCZl5sat966o38ap7ki7HfXo
PZeASbTVN1wsNlyK05DjFH3w/TvJTXlJwgCRMAAkoWp8GVY7sQdDqlT4xGlC1Mve
+8Ip8rvkLb143haV3n0hbXKjfLWgEB642LPbk2rtdGq2HqyhOXdwmoCtV9gjHq1O
ArnvtJRLkBUMh1hPTszIx5xfzZ31GJypFh+gQk6b4j4vFmmrVj3jwdAqYg6yHMNb
vpW/opa0mJxF4TmWH/TgjV3+tCl0WNLTG5x7OcCMlLKYYwfBFBwUfvhR0HWQqvIH
XBofQSNy8rPmRSplx7VfkH/+yoNRuVqWGhqK8eKCJBWGooiYXvQNqoRqOD/k5JCK
OnBuTP4DtS9+H7hLJZSssG9r64w7rJ7vaoxpFRLvanEA5DwsJrfL6aitxqoYBG/y
jaRZatijuDnxfQuOF+jT+tBMh3tk7XxtVF2GnUwRQ8v+BzmjI5mF6FmwM3fBFXVI
O8I6mw8rqBohtVrMB2To5Fi+gl9Hnixyvj+roYyuOotJmI3EOOatPs8rVrv2TFRf
qW3hkwTSOMeX3r00IhxJik96zjjAtJnsSrF4VxZS7iF1p7xVvx5JBAzZJz4aWluu
utFFpV93MwFz9/mhZfg8D8iWJamwkzN60qAtR4CCkb+MeD3QPS1wf2s4ml7xLqB4
eK9NS0f5a38okkvwzt8NM67NvXV+P6+wc15GkrBXgbSg4B2RM5TutYQUk0BERFN5
S0HMIfMAW8HJ46HCTG/JBr056C17DfjnL3/8U23c5pwzEA9sWxuOnn3TfLi2yBgx
LiP4fPErTKAgiHBeKlfl724ytpYEDfX4D2vZ+figyR/LcOushcQM6CXIGXokf9Qi
wUSPhVR/9+qc2Hn6eLo2iW3H6LjtXNYwi2NMdbWDMrHtmFQ5FsbH4hYnJJO4BrKr
4p9vbDfVhgnEv+4HM4UnGLYfx4myLJjmrxxBQltZYCA7nNwUmUzsmBBCAcKHngNN
0gkFD3mn4O93ptmwUFlJySUZ5YlHafN8f7hi7Z/4Lq8fcwp/99e046oEmY23Lr+q
4snODZ3quAlOUjhzSVVHSbQZoMCCEeyD6Nquh+fZfsfO5vOWQoQ7noKl85sa8tIa
69dGOUrQ6CUABy/lINl9qAxdAug9ZXPAEN4a40q6eKi44N4EG7jCZxYXNsfCyEWA
P+hSRKU241Q6rb0bzcPTX6kjVoQbf9lEzpxZCct5FwPaKVKk2r4cb47gWGbYOQYP
RHYLsFQVLNPV+ZKjsxadP8VNXuNVlm7t6H/75KT4GCc5WPzzQboaBt4Aph2Utw2Z
eZgU4eDT5O8qMmmMcvFbPzbiKUqf8s11Cq1fwhlvJ84Jdr+3D/vjeNNrSypD78yG
v7MVhClz7B2QlFg6D7/+rwfOIkUG30UpjMm6FuC45n+yNKmBILR5mkHH3ioaPDZ7
CIbggmZzFk5Uiz3Yo04vszOUYGgF97lj3I+fsu6Xy++6tiNW3R6dSMuZwDHzNho5
uQGh+dQoiYPp3s5cgPzvi3O6SS9Qw6UuETcbN9dkzdEfoDnAJV07T0CKSKbKeMEe
5J5DgluORcI/C9G77MPOsupoZ5beH/MZ1Scu9ZAzOhmf6ylmKyxdrSMVBtu2iw5J
7Nt1tOWIENz2rZ+7ohZUGRf6VSWbYdORF7kbebWxnKadth8GXNKMqjZKVimoDm6R
VCZv5l2veFfJl3wBTl7BQBABYrMqGLpVjyz3dc7qmG1kp02GrrlJrYAtMy+BD55R
EGcOtZHXPY5I8l54ahG38EJzXSRlkn+BzLXHvcyOBXD9qybkyBRrWbXT0nWuDsfs
Pw6+sKHFu5aJZPwKTGKotK8+yHGBiKAM+4sRHmROZ9QPhgJtSpryE9bGS1NcFBDq
zfoxd7wkzpprnJHdfXPvl2hVmtOCw6YBrGNiVNpNT9TdyiXg6Wb+gbIMT9+6FyIK
Xwhkr/MpfeXE/TDzDx8dtr70akQYVuUZ6rjXJnfKkme3M8WLHNHAm3QRtiLrXuKY
JlMm0vbMvBhNK2ZPHMFCGYSpQkSoruAiv1jk8U78y8sAG1tk7qF4ESuJz6kK09Cv
aSmEAlepWWW11IW0K+AkBs75hcxFeyB35CegiEESfpNGKL8fVlDaWfPTsLpaWojo
FMRqVd/B/8FMcX6o4BHAIitE4HEJD2L3sEVJi6/JR4UhE9VjmY94aKZ/BQAwgM+q
y3ag9b6MpIbYMsQABoZhjfrT94I4X8ZR3SAEIXW3oMr4Wi64i75ZoROlJkXSNUPK
H7hN+kPTQeNTjuR82hUgA9Wiq84Txwd1N0SyMCaMgr7crkvDHJkHvRvO5nFBp2Oy
BS+3Xm46kBzXeqkfcHuGO8Q59/L3ycSeShByZYw9dW3uv5tcl5g2otigf+xPsugv
Ey1rt+r7E2uiGyC8G0ev68KiYmuyiBICw2bPFOgDapDA992xK+Vt9VPyKizSV+PQ
8HdYeT/t+NChmYqLHxvJ7uAxdkNHxv5G1cqJozWU4sTxBdd574Z1aqNuE5M6JPhr
9zFtOSm+Wqb11unraULTsc6HImQgWImsL2qHk7oycq08qXjhL82sFAJKKIN9Cm83
J5itmyAD8FpKw3DBKmqpHYK0wcDk59fTpkWvTmuk4gC3WhRZQH9az980TAJg8OZH
fDLnBROVs2mSbzRGyNidXYPuqPQ9WeVtEC16GUL6+akzkdrN5D7nuyhCMhW6l1G6
8X8lTlyNQAusBo0rFAdCA/2Y8+zH4qXex6vK/0zRx6JY8oNnX/FtF+JOV1WJCcR2
WEQ5FerZC/1hJ8ZQBqmgvHRVsC7KyDLe2CxMyzaymt7QuPIQBijOU7CxVDvx2ul/
QbZ4AOiA1Ivk421F5+s8hqCH/kcRCj2gcQ/0i8Ybj1ljLz6SNgHv1jYk/1WZyeW+
fo0mMR3/HDKeIdemPf8uoFO4W5Ay02DUEjwRIkVv7Z9hGdCbm/E9jz7lx9uMjSP5
cqmA7ieD8U4BXB7dANFSfjcv9CGCZ/0L7Rm44Oe2Q5IBTYKnM9JVUw8+Lo6tHJPF
tKBXqXo8iCoLm3X9M/FuYSsswuc0iw6VhbWx0mcJQdBAL4luqwE0X3w7HfHk2bEI
w/Mmgm6XJXfEpQW01Y0ZCgTP8XOroo7mjFBHjP1QADqRrc+FLOoy1gaUPOfRzXUe
6dRY/sXpy299J5gHx4rmH3bx4c6/YPGO51BJtA9MWeww/ZwKAfjw9E0+Q/mNY69y
QDxSIMv15MTSPYMTNy+QvFE2zWrlXCsE0rhs8XBDNJ7FR5YVqypvaxQtcsMh6Qfa
mfX/zruXb07AFqzpDNLpxMe1/JAz319zQcLF5kqrADpy23xGh3es9eyvmDW//aXF
jfc3k9zwtc44K7XnPlYIwspyn3TnrsR2017zbFtt50fCIG4h3E6wD9R4D7yDLoAy
aC0yPYZxqqVjFgvpEhdEF6ImPBBhBxN1k76/YXc1mhHjGDEID91EKeErX425VEc6
9J2XIoeG6VseJcqLyXM3L/tMYzILAVCpu5lrE0D5Dp0MPtzyIW/x77Z+JhiuSPkB
34r7trk7zViaQrT1+HioiSUFPxx6handIUQZxN97b9sl+1XDFwPGuuN25v4/Ejnk
s/z3XZp/yHCklxWI12of5gA6hsvPDmc6Olc6PhqvZOjvUyozDldLhGj00Lv3JQzX
uKQe5UhK/XS8rJvFyn2rK5YFUFyYdU8DJPK0MA3saxMLPlezECH3r3uPVCFlNY4S
3C5r8VQ21xUhjgTTO4NJPCA2Waqdc3OGbHVW9OKxI+Abmp1DLU5z32/rGyKa3iNy
lFcRUuNDVA+qkDFhkVnpscpRj8rhVs0xoF/SOjw4OUuS+TQTsttMSX3ibfCjAHND
/Uok2ze6e5L8zk1HU7aO3MR/BznKzR9qhP/8pFr2OUlvnRwWk9k00qN5IWOj5Q8K
R/AexZb7fS4E5ixcEchf9WdSSpv7znfPSZ1diDiT4DVy+xMplVIz2VdjSwgvlVe2
6hXjLs6fexC7PSSRUEOcfW54phtnoCNN4/ikOFaC8F+7APewlpFVRf2N0dI8381G
Sud/cdV6tTg+Y6+HyoqxSzNqwiSdRap+aQBKmwSvRLfmK0H5emVQNPNm1i8kUJ8T
jCrCqQmSqCo0n8W92m/j8R0ECXcspyykFDXN6jHqmTI5TcYIsMMUzGDvi0cLyY0F
EM+JQB1nI3SS+c9koMENlTmUzGii1T91uL7nmCvwqnNPo7520k21Mh8rOsORpXXH
OYjR2Z+NxUHdodOTHngpBU3bY2LEr69UxCacCKOP6jRv98caQi9TKIy7P5d7gra6
tn70Q0lsCj7qlcqvqPBcI18n+JaZqTuoJJoc9Kg2nILiX3nFePJIj6vl/jOh1nQ2
IVMLPg+hgl3oWTvK+uIcpa6EuCJ/3edLj+8lLHmxuzTUQWY/4At+XBLARp/noeyJ
Tgru/z1iLUKw6/FwHcc/ZxMEfsQz2T9RQUpBqDfu/8NfhQLVPosMBmT03xgnRAJl
PmCFkOZOmPSELVAhLJOKalNxUkU5edxre7PvsOZt+5uid2KfvfKOL7VXgXWPxdwC
9swuY7M3MsPK1kinCFewDQRkY5SIg6T2TKexPE7jXwvtYj3Hb9DqR6SoFw6H1GQq
U+L0AYLUV8WBzfnas3ZWDYNEaK9ja7o/KEe/E7mLDs9Hm9SqFM3Jt1T2D4GU7/EN
5WgjuiRWfBJ+JK1NLv6fagNCw8qBOyCpfFe2Uc+QtWgAyQiLeO6HUcus53Mrqu+V
KEb0pA/l/FBiLpx6Wu4WomqiBu7meheCF9OFeRoqziYsK9xMiqa/mNyKpAxesoM9
4ch3WXrDY7YxRoF4bGIzh5RMyCIm2Aj+pvnY8dn49e/Dz42YFEAHF0GishuNmbCg
EX9Uoz2LnwiHstKseBf1kyuM9OIL/hVJnA8PRo9diM4TA2p6Xi6IY3Abxgt+zYOL
CzW4REWXAq9qIwvsoLJK/MFtp2vELx2XsJAuHn71J7OBEZWzGB0oGGm6Ktz3hUo5
N7dIUnCqD0tDgbakC6JkXS8dJyF6AgBEa0Y8NztDtCAL1Dlf40g77xrhzCzG7Gf9
ChQc3ASJcXw8JukKsbzOyU7Lo4Vni8b++7qbDKOiOzNHILHW1IIbfYCuRJALpF3E
inoZeQ2CQJBCxJW6BLvP/tdg05VDmbrDf8jPlkP9Xtlg3g9DxwzEFewZSCClzsaY
zhSyhe0/ievkxmU5yPLDCwGI3XKUbdJKSiIXnzRbail079o+F2dysETopsFFRD4Y
kH4WSt3kWhq/DvoRQRSY5QTiw2FUTr4nED+RxrnAvS4Sa4vIXZxIigj0lEPGXjuQ
JKlmGFiYy1EeEQ+OlwdbItS0FHl8BR6y0wgih770Xukwsr0x16XbtC+WZVy0aoKz
ar6HqxU2L3kMzFd6ArzdvIcUXgi8oU1kYyXYjc5SGDKTlwEtUTu3xfSw6qYerdyC
uitnpcpiTjBBpBZBQJ8iM0TkNDUt0a79GZYsmpE3L1BmlXFI+R5RTqi/MNeEBQHC
srXXN6uVRHwO3gtfZonJp0uiTn4tAXghTTYdxafuTKw+xhxD2dsV9Kpl9Bt3cINS
/NVE2azE0J0o+Zj2/FvGrnBnkV0Duj29S/0EKa1SepatCHbRqE85GjZMd/f9/SZo
ppYw6qemoS+GiODyYCMHsrnpoLprGDCjk9YosH2WlaNDNwG5NqOtIgw8QJ5zFmn+
GTO2Qf6BR/hjN98vMNcRZCKR7Gzu3wrpp0zIYLhcEvEPOsnbggJDYFOnIRo3O2No
PuwvLn2rr+sDNLNIBOaU9hjlxKqBAFkwcKjAeXwps9l7aeW1gvXO9iewEDBevjjq
0PliPu3vDQODDaDlWoIFRCL7fNGdOG1iLo434ykKHv4vOCQPORfPDNEI7IH6N0nZ
tCd2tgfieY0M0/6Skwyl+axb/dj+qGKA36xmX65+5m9qyFi5yqXOfQMcujzE0Yhh
ODCk/uPAm6izNitfJlNb/mGZHV4gk9GwG/PYa1nSgmehYLcX/VWQ0WntmG3yJV/R
bNfYSKFk3xYbaDAkPkyLAdg286Caj5ViH16BE/bKXZWeWfuMNOcxDAT22w8bkx0L
d66KeuMWppo87EKwVNOthmXnu8klpPuyO1V1545Fopwc5x8T82E8Dh7ZH+IlQ91Q
ObLgPycTzdQEZcIvtkqf6Xtr2jI+LvuPEiAmnoRtftCIrADIsBkneHETAJqknlfn
TmFTG7TMlfMw2tGdXC6Mn/irdOYDvs6BNLKwGraQSWgoMyKGROB1lDXcNwEpnMbM
xbKu2BmjvbaDD6CYMNpzZ3KBTSsfrjCIc4U/l0xXkGkGWayQkTMez2J3Zwl388R5
jB6Of/axYmSOkDP+1mYgQaBBW6Socw2ibPZL43t36zfOdveDEN37w6X5BXBh0cRE
HOaJHbvsylRSWnSmpsdLKSr1d437yXWdHkhIUJ1LLpbnQxnux40/wh2Q7TisjL++
D5gMzh47gpvWehkkegbyCmYKedJ+3zFnEfwN3m3fEK7InlZQR+INbmYsMvFeHYpp
r0sgk1MFWbUkQAFYA7vFfe9rq3DXbQQfptHGwEcR/j26LpbmkEq3kbhv/uaYnmbb
2ucn1M+GMG1F0HHVDC8lBUGYbLN/uDp/S8e+dMs2xn7RPNGGfHqm01jGbD7zVabe
bIwMXI9X5IOLg0JDHsHqshTk7217AESd/T5z7DP0qkstB0AUVDkWMKw9XyKfHDwM
umxfIvS7eM8ZPuNyjs9WwomPoBZ77n9kKO7bWdTfh+kUZXDVNfQIp6/AhQQ1A6KW
Pa5jjitJI7u3Ks/JrRVYSYsPcFgyh9HJL5NNYsgBckK06LEY7VlzurP4/kGcBhkZ
E2qt3HkRQqllucS1dlPJN6jen9B5HeD4bREwLVbkuiSNEagz52zHfC0hVsLzJOjG
IYXEyfXywzRPSuqcjRf83TSFz7VoTAsKbt4HsUa6iVBXrYAAo4neKTzoZi9eux4n
Cs1rWKPfQHJeiAhXqdzbSPJtmgAZ32G5wJXYCZ0W/DkqVbTa3PbCQTLmSxZrsDuH
yBiap7pCOI6h1GXfgHol08O2u5wQYyQcfe2qOGpE6Iwpq7P5kB/J2n307a83o9FY
g+1zNNnFek5gb6xGJfhcSEbllt4JAser26MuNhyu5dykkxXyInrXf10+EbTm/WqY
9Fw2EhrsJVYmGk3pD1yfoh+19+qKeVSqe+X7/6NpG5DoQ1KWNvFLvLSlIm12gHa0
q5sq27lkqhrz0GEd+ARWXA3DJCDdARs5gOBQPtE9etMNNaa/rwoPxhPKe4pYp6Iz
yrI77et1xdSCcL+PxmV5hYD0uxI+niT8kSseTdekyJbngW7YkRUXoJWGfJS3YVgP
WBoer8a1aeaWXYse/r+da2XHNGMSOs5fBIbtAMxqfM0rbgHgVVQxeIkqxlhAeK0x
BvgN2RYYLu+Z3owhppi10GZ6wUs8aBK3CDfYtPIgvOnvb773rFvgaMkjD0UC8VL2
koijtuJwWnN7nI+BilHaEJOepR8v+iX4A+4nJg5llKxrpBbbRpuye/xG1GNHKwnu
6JMuzooScAeRwKePRt5dXFMHKT7lRGSTU9B6/XnPTRkmmRfhIJmjgE+U/3gDQsM+
Cn+rboyykm/wruniAfBR8uZnqma7dyd4tfyFTN/7XivYr4DuTJV71XZ1EV3Mwxj9
c0mWcVWodqj+QU9gdreYcUH84O2ugINoqYpWczUB91+v30jQE8EfOEZQmKf8DE2V
TGVCE/gEhYOp7kXhjHBtW+/zBuuYtAa9/y4toO4BKDRthhvP0e/hEUh8hFEQ4LrJ
plPatxYu0RKiF/IURS7Ulq3d0k2869jToX1WNXs7taOjzmRCmI5RTBjMW4Hs4hji
zIHgP7GU5lqucm68eelBgb4AU26YtPQ2D5sF+yPwGim7Oy9icNN/kNglxzm2nhh3
kyuYy8MUepqPJNp6G2soJLW6HollrJPqn9bXqZh0YDCvUvG0WclLqicf/tUmtUL/
BBITyLYaWTr83dOaHzwCk1tl+X3RfiKZLbQqE1C3kGv15h5bOAOmmfsC0LomMd4e
+IbBuzGl2Dk1maCbIFBbtJniHH+SMM7f/7hBikYuTJVBIs5Be+L8n/e8XvZ+KOC6
xmPXkbVE2xn/y5uNfRT+OHPrRy1dDsrS0JcpwSQB6ETbvpFfBBT+89PdyWTKyb+B
pE6YWvBoUQwiPsyAOEul/RdQIAUskVUhhuzqoEAWg0ypxeGDeujOBRo1Ovcs5qBb
zc0K+nlTI811itmNmiPjt/Y9/Cefy94/BGt0v3iwsleLa8H5zIQpg/PWnEtlLi06
WM4DjZu1D4JOVe8JvfHpzS+79nRE7yXW+eksteQKX0agZthOLr2OXSkyvwV1O7iw
xLaQnGMuOPZIxtq1xjO9oYHotRKgIm20rz7HQgyIyd5NsV6kyZxwNpPdcHNxR1XB
pOCnN9JJSImNiS9uQq/VBeyZJ10+plUqLNBixwIAGmpvyhxbyK85vcIkgb9k70HG
he+myJPBVeD4E8KgoQ12ZiI9/9HdAvv1Ee+9UyZGMGWrV2P/Wgj4HyRVhMRodrz6
OQ4UkA8tuvmcig1BjFjlIun9I2/LsPx1xEGB9sagk2HPXR/fVGXFBjy7T9wPCnqX
jx6oXbqNCagRLY5xhPmN9GchLTEHNtR0VGka3sgyKLZZM1ELbYtpVO//iZNOsGMy
3OM7q7tapTNn8VM8/u6/ifG+698N5y5yH47dKzSsdC13oLwzn5sQUrnFQCwB0i40
JQ6JmQRjehQbD/YpkPBv/JZu9yerklEiXVOtIK5i9VaPP91N9GKrJSWgTV7zoj1N
LKdYsOLYGlXfCa7MlhlmPtUVENjykn983c5Cq/XuS+aWityHd6clqYkk2DQk4xwW
VZPiU4EkEwkiHDBRJQgBcN8I2RhjnI6AK7BzsKtk3Pf8pZKuXwrPrlPVPvlqMmLz
RE83o1qeQ02HXyJaEZibT0Qyqe1E0XmATbxtIpxPbKJFvsS+79c4X5eQMmANmcl3
Ic0fyXYdQ85T8AXu1L7XLzZ0DAaSkLKzXd5t0J5ELlBnSDhzgCfsl4dKZ+fVPdtb
Xwa7w/1DYsElmb8omml7u77zRtoKPob2hvS4irqZv6tjlSNv9ZACyknsz/wKp8jj
e3t4R8QNsWlWJ73krleG0b3NWa1o0twJGYpvsZ91p7MXAywxIXvo1uaFFozOsipS
e79kUxUwK6XA3Dhsa0BHsHGMDYhr3imhEnrwTeXR6SVPr9fPhCyqIhlYYwXIkO6H
KlJ2oczOud+2nqAljocHSP5w4urrHL9YDv81NYDd2kBh9BEDXj+n/Dw/szMCAd3Q
AruIAGkEBs2mIL+XLHmOwIvU0Ipd17rmwbNW1QT5b6gSWTkRSUwKoVCBrTpo2x0W
0Rso9PvFryOtn+177tcZXJXndj242Aw84n0/piQqknmNRvli8/+jZQxN9NhCvlCh
JBAxnHeY9IOd+yRKoa6IqscW0fRLFiHeQJSPI+VmcZwsyDiE+XHMXma0oYCVWBLf
kdmRvI/JAZq5ANRRQhIVGmBpBMJaqOVPptADzBCdoVsvGE7tyUf2b7DLW3yGNShB
TZQglUutlOGxJvrs1AKTrYw7y5oXe15qEF9lPHIdhdDFS4Sz70a3zHM+ZLRd8vQ9
gkuSLRmIrpTpDchlLOaBxMGeYCyUBXF5Z8PIi4279XITy/pBPK8AZNTdOznkyYp3
OZoNk0Fl4gIg8Y9/uLQ4EN35CaLCJ5KYTO4P+y7TYirIPtOf/vUinEh/MEPmwvxW
49lJIYqj8U5WMVWOE4ujZOhPB8EeUq6Cagi8XJiD8z/QDbrkuR98JzDQRdla16Fu
vJEj9K7SlAUnfBDBaoOcrfc/uUXjNuLyEL0NMet9Z0guxRzonZ0U0G/G4Sqy5qKq
TaRU9yGelJ58csxe85Fr24atXCrCtEUUyIUMuj8si88cryfYQiOuUNzZSOSdN6xQ
Eppud7En5mJXjnbyB20ZrUXZ0/87sNMajAJZPVbyjJc37KlBKZKQvBnt2HXz7vpF
5l9QdBDygfyRVpzhXrDFKm7mhj5uL2NmLQ40IONaa0BOh+jTgfJHIJVpO2KV8JRs
qjx25hsLCbOh9H4KVdKlhHly+LN/d8rUeQhevxp7QHbXw33x4wfvONDWQ10I+iqy
eOH9NFT+KeEP4tFBgvWKEZWpSVsWiULnt9BUKM55+DEb9SwhVqyMnVAm40aG4n4W
0/VxWdlh9/n97oJBlN7j1t4+De/HFi08xhX7fGQSSF1/4AR2PztqGEtX/QUoERVe
0z66dzlG6Ot4H24yuu0sZr3wynB26Q1vF1hCdtDHlJt/84bQQpPEfyyK92faIEBc
aZtQlbvNg2kV5W5hxUw1kwnv+U38pg+thMxTtTSO5ZGPeYLevQYXdrvYPXZCApfv
3BtIJA49rCXrK2hA+R5h2mBeqC0Lmu4lIeuxT+Awn9kL4RkYEAfextx7lhxMhSq+
6N7BeVCpPHZR1u6A3Oy98i7IaCOdCgIZo4VmLYGfAWWhbeuFGTWJ6AYgrI5KSKQQ
TOoBvAsXZF1V57AZl1XoJW/Q4gGS/M76VAwHWalB8Cuif72DgxsUzUtn0xqZVbxC
ZkZfafCT+aFoEU49ZgkgM6X+AK0YMuRXeQCZVaB4I8rsP/k+si75/6cKA3FS+nfN
gD/Mu9atcON9HvfanbEnYnpkXzML4Aio8XuaOAiy35YyGbnvtKRdL6h6lWtjK5aW
lcz/HEIE8nWso18xEMwzfAL77jEkzgwlfRcm8nQ+ogB4pXGMMoNc33F9JSBrjnsn
lCPXR+tvxHQ+Btc6Wc/jABHx5ybyUavj0/LI9XKMcmehD/anr9RVBy1A+NBRFkWb
k4V2pwKtQZjaA1enc6YcZqx7P/TuobifYymT/oUy8E6q6INQMkwUBNqaCzQHOwkv
/MxB1vp91hRzZZXShkj8wXNwRomm7ue9VRGeXkpQ8GiOBxHtFbHaDhUk7EcT91M5
6WVWJcbBRqTT5Un/SAuvxRjVMcgD6lKYqv0ob/we0OptjONh+5pAzt9z3Fimg5mg
egNkZWct0lku4JY+uCOd+2+M5HrjVJwYum4AAF2c5l80lZaaFwljbSgQhU09Z93C
StBCY+1psLsxwMdfzPZV57ZMM38SQuRwDoaiXRjD29sZIjd9Ko3tqsp0IBnqWRp8
x81dXBrtH4OqZlgPQFsaCxoa8Wz96LUljxopoB9ZYJaxDU5db0GuPxq82FvCXhN1
HcpZx+8TV+k3S/ZHQ5fv3wwO+AfEczulYcsLxZMCjMgjKGEO5a/hQyImPAk9+bih
lZL+9LA/ewBKkNr4DoAO9rV29gm2FG+aGfKFdKWOe2T14qA1GrzLIYERU9/uGMqY
WsJfReLH0Ze6sxaxxMJw3czNgBnufBDco1R0fwLmoGUFVySk9CqYE2szLjJ/dfJO
H9FqM7Dx4BH17wD/AyH8jfeuW7ZsLm/MhOcGNmMIgx01KANjYexj187DqbWOH/Yw
OCg1cwm2Ao36vlwBn8jH8t+M9dMSa1PFVQdzHveZovSRwYvVjVyIhLJxZB337CNe
vk/Zcd16BUKJw+UcVWDGy1896P8vxt/azTU4J32L7WdmtvqExSdBiWVHVoD81Ly+
uRagqIcQ69P+t3tekacB3Xemt4fO7uP4aT0eVHr7v8U+46e3XyYc1VAnaif3gCIX
7BcXsp5yq3IEdgaZy80pRDuZ+VFGA2KBhP4f67yVFfYa3xUB/acP+B0cSHguiUl7
D741pkH+Aa2sOhUGMIfGIVJgrgXQTClX09IAt5VU6NMA0fmKLhjdYlRtoMLusfiG
t+FmPz69VmBWA1fACYTGo8pnHVCoEZ+4VQV/RFLQ81m4QNZlsp1gVLFo83DlaSbZ
OkcA6szOLDiAxGp8wo7deSJN65ZVaqwncPUtk5LhO0SIqkjBE/2SZA6wMBtjve17
bHTpuRRootxdqMjm9KZY5dTBCEzkgHKoEXRlDh5WBM1w3fZSuMan3u+GCVKKyS5j
PBDjr1iON5lclu5t0DxyoVXyRzHNd+ZdeMmyx5WIDdw0tZdQE83KwDsFALtBHg2P
FOOeFXovV4UHJVMV/leQlnyO2Gkkvb8ucHtumb9Hx6tRCKL2t9bH4IyG4n0TXNxO
shVHn8ZX7nmQ9dwEii61Udb9kJGhtCNVEeL6tjtG0nWd2e3k5neiFWLLsiSv6CDg
U4ZG2FvUKpU6o8C4a2SKaUJpTlwxnuiU0RZ/1skWa2ffxSYS3U5ClQWBGk5/WjgC
whO6AMX+bdi8x+22z6PPxrzKJD7RMbWTe214/gD/cj0KxnJxNQFk3WmMOhLrQfAz
Wc76oshsejsaVKrZD/iyRXzz93ZH1D4QdIYJthlcUGqvHTnD5kSSNJKfb8NrhVIn
eszF9CPotliwyPm81GI2PoZBUfchVB4tOXaOhWPcqCaGFJ9wWEKIa7/JsfsdyqsX
88jt4dELFOGYg4O2EEUUVsC3cAU23VTOdKoutThZzPunt/YVTC6Iplmi31m3AiBY
IORdSYlwt6E6AXMLqHAcD5mza4QS84i0vJrdhye8vVyknplPypfzP9B2QNTjDQmR
rU6XryBvg/KSZBedeP6b6Wq//o0MB9ZcRB5LxrL9erdcP9pjKJxkyXQXKRhLSBXF
/LWNny2wuAcrp4NO9JuM//kAWD2NI+74AfD9820+T/aC5Iy95r17L8radwZ26W+P
SwTVCT+mlqnitR8hPS022ZaeXcpyz6P6A3bgKsnpiBFP3taI+19N41/UgEZPVDkQ
tyJ7Lium1w4p169oGlF2cv9UjIAbRE88i/VSE7YFVlBdNl4VgLEL6YmoyzoCIxr7
d31zyNgSlZT6oZkYqezR0Ru84+gHF/Y69+AMgEbaLEUMs1PL60K1mUoqN4d9ZsHQ
3pX53hLVZ708i3qlvs1UrZesR/xMUcn3y9QW78Df1WeTgZJyULC2GfTEZGbFcb4P
ywuNI0Az8jmGhjmKqm17zIq7NOziQnaND8RY/UG5H/401/4xGoBU4udtBQAdrVOf
yK42bdoL6xHyhmcq5/MmaNgPu9KUZruIpEN51NMpNG9dIN3tUTzJ1Z3jApWQofsr
7/8qCjWQvdLvr24AU0tnxMMmadCdz1ay0xnSo28xvqLQN1cmt+cCtosT8odVvv2M
0O802x8GmfmalnljVEOkaFwjgBiz2WInj1Ohueh+tLxFrguDOr0ZeDbxpGD/w/lB
skK0BvJBDFE4KaoAGBTq2APWHlf5plZVE4+vz19b562dRQFFtDlLKFpH/3UH7m21
ZwHZokqLXO4rBa/PMiCXwyh6wCyS5c+fLx9A5+DRsT+dDMucKSusZmC2anAS0Upr
o41o5aVLf2/2gdQaOtMmnqS744GTPDuUoEnseWa6TfEGVNSQ6EQjgozSou1Xbnb3
mXwWvbiokEKGljtUjPKFfRXIMPtIMxEH0sSzTWuiFy7M82GRHtZzfLjx3yCGH62c
qvoxNMfl8smClHPxh7IrrrZHLfGw4PM4yNSQVcQ/rxguCQH6DDPs7NVxg79Qtmaj
sDAtZNUbwOj26UxlAAmkqODrGyr3aHDUfusB3RFPWLWTK7AmuvzUfbV7/FNgcZ/9
KAiueIObYJcTxqce90a3pRH4zwFB/e8qVUmpJ1UTTgBquFw73fFYoyxYyBCaD94D
bJidFhpsCQne7irqdf2KqrOSCASMsxTXdxUv+AVegQBKO0HnYs2r+TjyRzmLfiRK
UlQm12PlHTrU6zTcnSh/i+7iF1kY3LVDR8tdKtVGIouvICdgBOVQ8GmFxLdTYify
wj8YlERA1hHupKmxemzuBvQ1ytiRMn7IOIPvBmL6IkJWZWZIjLyKWlGS73/Mfzrf
6gMWMlDKMPZl+CAQzXGhaAt4/WdYnmyiAkYDsJuslrm8PwRHj5tCtsRP9gBiekgM
p/G1vUnDGF2Yn96Cr98UN5CQEqg3xA3ojKDxG1xnzYfqVkdQCKtHMIJp2IdffkTj
dlBPtLCKXPmK4x2eQRyjupRg16ZIcnI8eahCLFlwtlHOK4KX5jcKXbwPm0puvVgY
DC5Z0STN71xNG6y6dF/tYi70pXPIsfdbf7LXKosFr3t4LadcP/twVUCuM+LD7J7w
mAJcfOVSMfUiBepTLzDVm6b5pnUG2iGOVaNMXRtzkXtfVkJ7Jt1Qkb3c/81IXWI0
auab6oTgiBf27zD8ZeIexGeN8A5suSmYZfI6zDAxqIptJNgPz0/OGlqOaRn6DXEj
7pw4D3IDO8332wrl4RUk3xRONKYzaVfmjMYKzC3Ma1qyzX3+fnrpb1kaUV1rU3lk
M3uXf6blC5KvJJmDAliiYdpXiHDOO0+G0KlnEGvJC+/TR897QNoWXx92yaGpG6kA
77WGEQZUJuvuMWzkkr2ShqUzgkaXCzEe+pob3Q+VCOKcUxIgf8Jxts55uGZsi4Ht
6thJrto7EeO/37YJioNpGcFNQcZ7EjdkIS9ws5o/cKFPOKT8HeTDzMh9pU6sh032
RO1ju1c3mTDFifSDO7ncvDNgnt711P89rpDnOQhpdtZZpM7wzgpLf3QTSS+Onmlv
U+B9bIt4QWBWMbiKv0SlLVsmzz9PaSmQ9HPyrkae118a7ORrVBYSyhcMUo+THGHb
bO4KPVCtGQTLBYuP8Jzcm4dKo1znW6YglAortfqHHArlPXuchBpl1Q2KNzFBOg0f
v57Nl7UR+XrpFDlMzsKQcBFSI2zvRQ1puE3jA7t3u4zb7wbawBTuVCwf2K5WrZ4/
vwKMZ7JfPR+NHDL4e4XU8pV3OAeom01rYLl4bO3lZBifXuTnhgLNMlEyJ1Kxz8+p
BFaorvH9HhU/P3X9JcusPdDPqYA6B99Rpzbjkvz+TedgS+J/XebLyHduBf2S1y+F
GVAuhdpjLo+AiKx2VhJkfCZBuR5KUJV7YBzdm4JIw+5Tcy2RdJYA7No4+AkpAaXR
t+CVBM0ePvgIrDHHZJZZy9K9SoGyREvVYV5Ee4lolwNJseZZ+EmuPC3BcyoTLgKD
xEi9mB1jkldwIuG4WJkRwynVnprK5vjpn1lKF+H9j8dK0e8KAMYjPIz/jJrlSRcr
xecChGVGw6kz+sqxnj4RJov9OwWXNvKIWq9WsegQx3uVjvo03npPaFkh0tXtpjHv
Sx17fHofh2ZWMJOsABrEcO66cC7VPifX7hOy0IqHanxYu3KG1mw5/wGCyY/gAi3R
AvuL33mkvB/4/IT5XXY3oWDKnPNdrtXzpIj9dpEMa1qbn7rfLnzMZkI7QKssFIZO
0jrpMpeV82Vg72lZEksIczIcAHyemBwayyrDHBkrj2wDdo0veZPuKMUMlx+O7cY1
GeVZL3t6aDAH0tLE1Ch7jsvXVmLhegs+H59/wTiwijbiHeYrO+kBIINoIIe/1Hhf
nsBIEhnmwR9L5uCDDCUJSBgvVgPQkKQ6bCkfCfBKCuAaninnTsLEUdfkMYZ8egxN
iJRyGz9j0Uj3/uGIBEFVmoOe2fuXvMzS7aHtCxNZG0aqii27zj13jbbQtTtuMVLm
D/AyeShsjmklJ56wYTiJ+Mn814XpJQzT1j3my7Z77jRfNAYKHMD5lVXzrW15cZTU
DziWBBw9N3j87xmWZAxua7dKCO4upO0LDEb+oc2K2ngF72R7RBow7y3vR/vKRM4a
gTJciHEUvbQNth47B4hpS27LM3Z47yLyqnyHT/A/JfD4NW3VBZLVI3taJCHiOx2r
Hc94IQjokLl30vkr84szIhDwOWzZ7IZqglR9R5huZFqE3soDYCalTW4eJMpoCP4E
hjXp7A07+ibIbRH0weme0sKC78pFF/4Fh7XXDBcwFgbhAIMF3tD1YOIkyCWTeIL3
eECmaLImiT0wb0bSmYGNU0h+/Sbbv03JDdBSs8Wdmz72bYE8tpIn9k1y6xFsPGbS
yuZ358o6IAY6dBeu/1TSpyZFfLCDFGJe6KU4CcfnMPNyjYbXNHogJdWPZ93RHGQq
6gG+IYSNCxk7MIEwZEMwV45x2M+yKmfKZZO8vyVImimK0QD/6kWYYw85HFg3tfv5
U6+9gykZo4chem05XodAnBOux4viRT9ZqwlQb0kNVA7lIdjpxSXSfFvbSYrMDkhr
DuGnRTTixfQFc8aS/excc2bhZHaY4aIcavV9T2HDzq5p55JIxHlYcXjitMKG+ZPb
q5R4+X0e26EyXmCsB+LQaxlqr5pd4Vrn5YAX1LH1pvYOzo0QZDwLfDC6jf/EzbFt
nh5e5VKLsFwnZuvJ1ntNAGGBI0ELBTaAKLI9B9ABVLtfF/TauplOaGRTjjrNLyeO
qs8xbxl0V6GCzC8r6nXxw0EVQcRzEKoyws6tJSEnVEOy1eQP3CcXfBKToV/L+QrB
c3NATErMB3iplnsgBbZvTfxaf39JSOGfXr1qBpLDaE6t1PPCGSf6MF2C6OPKCH/z
BIub579gcMMmhPDN/jG7VkDOsldpDyxiX4zEoBZQmBVWOJl9LyON7kKycO3yjiAX
WiZShGdtmAWBSu2x+e4rAvnu8vSpbiCudchBuMooMgCXPplajhEgEvjPqSV9SgEW
T+0lUWg8pkJ0i88IDVCzuvogdyoIScrtEpslkcEyNw39V0X/Y4yJaLjiwnsnqQQt
8eh7erzZ561/8t1Zz+gSJa3pJ6MaOQaqoeLW4Av7nYy8vSqYen6qKXsyHAbkKsIK
Z8ziky0/YEQcLt7c3bELf8gtHnqy9XWwi9jOrdm9ChYRHYi/n/DyQROrVZXiVLbX
uxfNDuzXY/G487Ja1ddRX7xpmYDbJPyJu7w4W0H/RbC06e60ZrSwb8RFhIK/Pt4f
rD1K0MZUjZvcKszrd8isCeFGhNHlvQR8e30NZKE5t3eGpHNKYmtxwMnsApfdUmM3
I5CpG8scNtSj5UrEOAPsr2DNryMrUoU4bIVnnCza4SjgmpNjFNQkvtP0z3j/0U8I
9FCblYl4oDFhOt4JZJNOaN6KremysRHp+f/zQvqHnb8yKKEWbPrTNLFZGT69LJUS
YmEQQGKpl1KVCi0pMOTuEQq8RshMPMV8Mxb0Eil08g9xj7A4Ur9005PWO6nWarTe
ii3ewv1mmAic6GqFi0fLxT+gxDr4zF3IVLr3Axcn1BmNQJ5zSMr2UVVGbWoMwG8y
Ip155jJGOoSSq+nfbidkzayHIW5x+lQoj8Epukx2UrLmZsDJydcsZjZ8Mzrc7ZgS
LagUSRRa/fF0LlO4HADODztbs2s5ZKYRsT4G0n2TVbhmz3V3VzVfpkiU3aCGlxkR
iYqqqdUQiTL+hOxw4qGRBLTFDg2D4H6gWMnUjZiz1DD590CZQ76kFFuoC5P2eT/c
mcCzhlWwUyW3RVF4hthrabz/iMfKxHtdbSFcxjLv54IdooSf9rgeusdR6wNHZ2tR
SG2QGhYS7F3SXR8/dZXMMnD3rZlfXC7eWOP1T1g4BKJTuNDbbyasj0U4g40cVsnh
ZK5QKR/8aAQglm6ZwP2MnnOe18vjDZM4hGo1JTovviuP0bUk7AoxLRueKzB+2N9y
xJ91iXh/mzOVU8HtfG92NaHKKSrtxyRKTypxzBHNl/a9+VVnV1799bbwrl1eRluh
2bWgpONo2Hi1Yi7ymXCMIdSTolAnLPVuEDSBCidngaiPcUrn+xdNFQ/t3irY8nlO
inieELcztOd6RgTgGimwZ0OX2vk1iKD5FRJ59Wh9JhPS0fLxws5CSrX3HlwDDRsA
Ojq/LKT4mh9VYxjM0lzvBBRLTIx9moUOFKmvdiZDY9JlrIcDGBr9nglI49nHlMF0
YtEiP7KZ67sR8JGZwecnro3jQYdFryVAy3hcTna8mRk7eSejhivGfkq89gbjjLAc
5f38qySKDaMxaUJCQDrJdjOO+lIomcHcIR9f8wzw/6QeQCOlNRdKvOjr9OGHcMOo
cXT1XmbxgRIwxFMHJyR3u0VzopVeBZba2CgLXS3bFjVC9KzW5oCasKsv9TzSDS+n
aqpvG/AxoNEOxahvQKgjQa2wTAXsG+eowKpW+x/uvbH/oCtEDTmXJZHuNHyasdMp
CWyglz+kJb0cFFJjC32XwdLktlzUpoBxf2i+5vj7yiVgix3mxzP/GNjw5hzOjLz7
vRekpITqa7CMCfVXPslgae+cr6gGNruJ4H7vy33vdRBtln7h3THDACwFVC3duib3
tAu0IK75e0JMUptGJX/aWWdX3tweCeiv9f4EoHsqQlJRt3tHK7r6CGQ2v7pQlHgJ
Pg6A9krv3rsYVthW8evjajzft1B3o8UzrQgdWg+F26nQoD1SL85CdUpX1OLRJclv
6nnk7Q7qW94RlC+cmJw4O198BDkvxj31RbgZAXJAOQSWCk2WjfCTimhLtSepLiGf
PS78LFp6d4nsWBIP31u9Yt5xY61e1TYlBMgfaECyljgVMMxSWxeN8LJsAaFZHAON
AIFQMtUV0R8i6Mk48IQ+iH5FW/6VvgQcUiHqZo6X2AkHfPP/Nlb49X0NShpPdeyB
YuCqodmP8o1H06xWZRycUnR/eON0nxZDwKjKX1ikV1rpufdZm/U8VKPGtDS2MUyh
JaBFigVG7qRab44QE4V2E0uBODyVJcJmxRUwZ7ERQ72x/Q5Yd3+k/rQJ5QwtwQo6
EykNxkjjVn01ZVR4wRk2CHiajuA6ZrlVhxfEqdvy3tGBf175lY5YVJivklx6YTMV
KGIuME9NHpwmF3O6pnA4AYDw/w2dDTkqe1ci0DVGspSn/2G/oNDkKiAaVXLpzTWm
MmtZxfKBm3bYqvRVvzZ7Ihw1XavPWd25ff0GlWZ/46eqG1nCun8ESUE+kfEx/H6M
qzLj1+rTDxxmk3nGrzV9f+IuVD0eTyV9Xep+6uMOLlF8RFiQDsiMaD1Ov/9WRzd1
xLZSS5HawatkvDu/oVbQUkDBbUKXAHywZHXM2XH43OTds2CtWbCc+7Qkf1SvWG59
ZE/UwhK5l8yieKAFtuXTsnan5dySQb3V+smMRxk3irNt1/BJ72ZM7BJr6dENZCqs
OtUH8EfpNBmaB7umMPWJIoaIejYzO30vrU9R017V1URvVFM7O8lOjaH4r2yuNiZe
jnOWL9LTCZRatNCbHA95+EHfYIjItqCClBpuDDwq5B4JzYh+kxlDe55/5ohIxUJQ
GX/963CJrIWQiALecYEVyFcfS2F78agTAjydKHiRVjT7wkHBDejxhDXQy4R0dn4l
Bqte5WbbCa6/pf6EQC2rFJPRfgOvxa/H/yymLPILiF4PQiQV/X0awEWErHTA0H6X
sJi2IbWJRgSP0yzrlV8SntcgXwN3BDrO3RqiYgrCwoj9jU49yrcXw6zBTUTKrE/b
yijJJZiRPV0KAsxGF21tYEa+OIoJy/zs5f9DPoSMb11oy9/Gz5UU9T9TZo06bfM8
uD4VFJr0Pa/8JB4nYotTh36c03foYqwl3ySdGZn95RD1KUqzBO/X2HC+zsa/4OO7
rB5Qj/zv87B1q6gQ4fxVTjMCnvg9Kv8hEiuOGNEzn0nS+JXIvvsY5aOl5VPmajDb
hy3nJdYt3wZf//RnEF8GqMzia5AbVoWYXrAO9F0g++BqAWwF2IXY8SO6Qv7ebmY5
Pzp0M/CQuXb6QD7JG+VzK+QbSnCrDWRU/UN8x+SFZrrcAOPBpQ1wfqi7vJp4K15A
v8YMYvzuCX+LkLhLPMC+Ylqqmlj8Os01pFSRU6nvYCHCxeubgsXd4yrMN2Bh4LUX
luLS60Iag7VTYNduAjddrT3RZjpE4ssZu/T5vORrJO0x+ymkyN/zlkk90vCeqK48
2ebdkHoUfD9bFFRS3eQavaCnx5bTFT/yFHaLScGtbV8PluIcJ79Q0XnPhjzeY3LW
r9bQfwPBfsUDDGmW3or8IBIyoRv5Nov8RmGjhRk8KR8CERkXVeyypyp37aGECmR8
gFvgMisq5TdQhGH30bTPMFs1/LdWZJjljzgfl8XgsKncKraAcuqEz/4V/jiYIQC8
SKV/uDzBjIkGz6JFLxeWnInw7mieN/r9uCFTwrJ3Yf3Bzq1+KnOPqVf0nfCWE+du
VfOJPXNc/wAoVK03mbC6T8n0SSPfLnkHv3BcuirrLCge+c3UfPp46tWT9zFK8CkU
PQqbhE5Ht7Kew7jW08ARHEE+6iffLVKLGOGmd3UYpDgGTIVLyz0YWhg2wIoADaeK
JfH6qG9z8nQvu48U+20tTY80lLr4vxzk609EHsXECsRyguWo7UnHHbHECpGJQzQO
a9/HDeTwr70OJD3CkB2wwRsmkSmIIuqERGacClZhrqxlUAqEKw/4JcWl/q7+MzUT
7Q7+uG9ierHQJ3RbAoKeF66X69g87ru+plq4cSPVTpI21/2MIMCku3Ku10eEY09p
zuyDZYkj6U9cROeb/pY6cm5VXSe2oGjh0oetrGrPFAkrYrYCXBz/ngni/QWaeSMX
dkteZyoK6hAFCKQkWxEM8ff66wv1STvt0WuRRa2WUwuFr7CDLzrvse3gxeNeCxgJ
+k9J1Runk35aotvvKRHUB9Mipkj/AJKGPoQSbEYCnS3pvsaoEU7ZFByGqqfDeAJ3
NnkObNfnLlpiRYXZbiA/L8dKyz+9Hdq9CONWNrqIS5MT9B9m0legIega6ZMDTBYC
rkqLLUpGliR3P11BK+U0NC0fkDPDwBwQYJfBZoelw4Yj12hl+KcdVYGdWTO9oQtE
166nXzBZLuE5UNf7QuuSO1O25pl4DdYOGwtUkEqVTVvx3NFSeq/VvVIeTXJMdzB4
dwdMx7jSCqm0zZMH8i5mhEJCeJ+A9GatvKF88VDZkf39qL//mp6BNuXBt0WQxD0a
jBQ/BxDdwYtuP6ZC2f47jJVynptAVA4zmCYbb5du4p84u7EmXBfp83Eh2gakSojC
E0as2nceHJS/6F+JCQ2i39jmknJjcJ3UIuBG6foAlyegGT6/uMnsvUKtHCJiigj1
7mdrsi0ahWw7MOJKLSdDIrXklsMdV/kz6MDNcqOHVihMQKvYLlGS7Fuh2KM3vm5Z
VXc+H9Y5KAkoVNZPsUJRQlRpCJtefFiSxW7H30iAm+SExIrbBt6HeYu19CWor0qd
sxJrLZdaq2tVxG62Yzm+9SUL/UfKEOOHrIbsjIknY++ydaYmThQYOARQo8uM8Z8u
N1aXmTAeeu6AnhcZ7bI2UVDGHWWlVg+s8CAFJlK5eMeNLefICkRz01hcLynDrsRp
6j8F5xdLM7ERDS8eYfTgj4CoFmthNJCM9mB2P26XtAu4M/dUln/iwk8Lv6g80znx
vq87vcfMqRiduwip+Oq8Br9R1Sd2cM3LLbyalOVAgmrtLXJtFBtTD60Zdxjy81xc
lUbyKzYS040fzRDwwC8Bq8+efsYX0/PoxD7EpPRychcA2WZBu9YcPMdWRiygVo+T
PiL+030FICppCdTa1pJ+mAMvXFKcTjIbKryh/x062Hv00v6J+RaLmYfbKQ0rpXbr
5nLwknM24Q9nsEzUxk1077XwW4cHxAAExYzySLff0ow9J8LC6CzNDmXDxGBC9am2
37vxHmbjt+gPH2vwTKNpwGNfq64nsZ/hvzazbiAQEA44acNXUkqZjxhFfma+h8++
tfNBhUH4+OGoPJUcklNsxP6Db7/3UkwzFLA4vEpNoDdnONTM4lDWxm674iRkRCLu
TUyAjLo2bq10pNdP8EM/Sa9oU/jm73HQ/7B/JCxOM4PI2Ku53mj3O4a/XjFR+nKB
igho/OBpi/VNV2bbLzZrSLD4N2VMEG64NeP1UB0J/EL9CDl9z8cz4V5e/5UPZo37
jitWs18yo3T3VwYrPTZ3kL0aACG5hFQ7ljHLd+kiPLtTHxUK8H/3eai/5ijxtVcG
x6uwVgW9uo0XSPJNecOicCx4feJkBrkw/jla4xZ7NppKIKE1A41vNFYoBw7sF1S9
RhNtCin+qOaCTc29LJJObpHF4D1UUBWZLEDgj3Xs7SKMBq4waWm48t1htX5ZS6Uc
s2pPo9PYq1ILUbwx0inf2FNbyXCb3xRE85bM5Oscwi5ogEqt7BrJG0WzjsPxiK50
d5kbPnNVzqA+L1OqQBrNg+aVlQoGunVbTjJS0ZNz0LAm5aJN41vT8qBuHL8LL0uA
tuj/SIOfAbQQ8l7PS36EgumYUGmCDtNc6Nj7TBzFFxQwfFdsDOB8ADjNLHXa160e
72axrt8+yHn38EoIgeDd2BYWsC+0Cj5nhsuum2tkpvZaxc6UsOjecDyo0XuJq8PH
RUbslPZcjO7Nevi5+ElxzRtyJcm6sT/w8yhThLqF6VngljYUp3s5QyE9SshOCHFG
MZBVk9F+nQaLfxf9HDV8UdauqEmf8map/neL9/xQWHmZc2SRXHIj/nf8oBXgrWcy
uwFYaLnWf2NlcT+fx6Ve2ktl/Lh0F1Td3LN2YS/yCs/ZVB5EpGEbyPdB4Pi1NFJQ
wKUbe0vO3RoFBxObfPRvrX7R8r8icrbzLXPFm96KG34UOXcmcOCSfJM4HH3SHsFl
462fe/51RJGUGdorWWQbLYd2+U6qZ5Ew6e4H73JsBcfEQdxkNaPcrvL4MSSpw7kH
5KjJpYS77dOMcFyBbJKWoTNG7BR8HjA7Jrourr2CQ7xoJcWCpyZABpuUMJZgh46v
I51Bf7IQKKXSj1IfoohsztmcX1v1sMnmENphP9F3F18KgkpFAHMCU2zn203lNr3N
57hxXgfUzFaIJAsGY2vy1pdQnfrZ/Ns6ns9lagj5gi6shoAUuSXUGaG/lak5v9Nr
atIFTKIBd7gXaDkvZ+DV30Du61SgsCYFEdKZEaqxQk3vKAWn+c7MwnBVQ+QBV+28
bojDPIkOvRp95k7k25w4nucNU7JFTKBPipob+GzhuXmoX8aLFirpPKE/XABNmDf6
5GRL7O0ueMU1tsSGW/eyvSqQNFm7+bAcSsTa3b8z0VfNThM/dzbOIVOHcmvuW6qh
/jBnX5vKzhtnrM/olqZYe80+sBKiak12XX9fWYWQZqvbzx9PJxpdbcM3kBpdBVWz
AF9jKJMJx08iFtDoEtE6sbfaHxE0aAe/IgXgbIsLHgTC+QKZ3q0YaWhnfvvhvi7f
/E8a0WjD3RT7H5OJx5HvgQvq0su6IUvLdFrMORObjkXl9duB4Hux2tQ0FV1isyc4
QFa+7AJ/T9GN4F1hGEwSZYNrUyCmztAUmpMYdG88H8Sifk1BGI55Zd42gthqLoWZ
fUW3NVvE3NZ5hPeWEZRtnN4l9+iOwoKOMyLkFHRR1hgLsqyMRVYNWpSeZ8jZOt78
tKQoe2ZpqpkcGWMbKt6n1FzW28g/V3Qh/bxIP+E1MmFOSXTQNLDMB7LODNXg7znP
79GvHFL/FGQwAM7UTuT0lHVWeNn4clT94VQ0YRl2CAs/JP8xKALpL8RPpctybiX4
w9hY4HBL5t0cHeX+GJw8xR4T+Z2SDncsoYSsLAXbtfqY1IHfbg9fmCcXxMnKy20N
xGQED9/8as322Q3DNBdtmISxNNbK+zz/MzPf3W2lb50bhb4xOkL5WimP1F/T+F7Q
VcggHGy7BFhAJPl5jgc3CsRihP4ZDmXH0H238nzlN9hj4P117OUlWBggyt/C4Ayd
KvheJPipvZlfYQcL52KmZs3+WmobXQx3CXN51tenP0DXblQ2uyqZWLSiMhvaJF/w
uqKjgr8pOd4QleGiyh2APylTpTjSeJc9F8CUJtn6Bm2EagHCzQFMgNBY9Kxe65ez
JZSfRy4J+p2gSjvuUWQtMwYG5qgBvxz2uTrtBC6CG/5NSzhmxBYzsWc0BXOeF9oJ
JiPHl/iiziRI9kZipjWI8L99z54Emqa9h7eBsNUFpFhuefqyG9r+7+agEiepmfMs
qrhMF/iu6bxTvzclSY/kZnKSbL4vr+vKaw1vInmcnlN3I79ZNZXvHopAg57NijLi
j8d3TgovjagLUPjVVtZ1KiZPpRTf0PbhEYN+biJihMntr8S5C8TtBhhjrc7VsDjm
kubW/soQlnOQCyDH4a4gC744eIBG+kuSPYedT4CYKoAmyAE8aC3WgHD4dRBuWcPm
qCF8hB04Zkjm0KI7IPNFifbs5gjkIhykpPJ2g+f0XqwQBx8FTuIVmklY7QfHTodM
BX65GMnY4BRX6S3sJsvMseggk/GE+UyQslI/nYLkmzvbPnuR8odg/T57O2LWl4bX
BphC/hJ+8ugE8l/uC3JB4PCEHr+uhBJRMPARrM9/a7V+1snLstjZhIJsL19NRTCa
Ut/+IMP8qO/3/z8HwZVc4o269hfHrl20VTpL11d+aPex0QxUskOnMja3b/SA5AN3
BA7NV1t191Y5pYzHUno/NWeHUjKVnSiJ2/4BUGhvnReBf2BFDFVMMhn9lk7RNYN7
5MnEXbkQyyzbeVwxXuLB+wbym6kqxb+dNAt/0ri3req6gFgSh0DiItaWp1XUjVpo
+YRu3C6+HiD9v3l00NKS5DrJqksQ3R4RwTctq64tKB0TrAxmpSsCNlilTe7qwTS3
c+HyrN2f1Z6W4e6KAMlj2yEOoRN+sRVytLrLabB7bDMM5xR2/DILPMwmhy/dBdoN
UfA0ynUv3bxD1sMl3yXZn7t3/ddi2DMtCh1F7AD3k7f2fvE7oz7ExnuSSUAHryy2
fn4pXwWJ3AD/4XKV68JYpvdSzU8OhAIfmGen4mRnEWw4hrBlykvzNdFqsZktEJ7T
whsE82YaW/0ksaE8PnCjuVPMUJ9AVC+uQKA7DyMuZti/f/nlm4yfZnjvPI4Fmxai
boU2BH/2xcuxmvZRpksLXkU3F8kXMHhiifXs0nK0NRH1mtjc6fKiZANS3QZalM3Y
Fs5HjwuGdk6IxzUBzR2Z54zH1r7qJFZhKarYpC8L/TIk3w7Vk0TZ7fwsAY8a1r6f
XG1SDS+YAhb1OUfTSEBwe3WZhF1qa+wqhK9nWG8C4uPCnfPTtP2X7rbWsH05s9lT
ROP4FYtWqwgBkQK7836j14+RI/0uoNC5KfBY/tX5NY+ESnWBBemOzOPA4wqOepws
ahC3KvuSkyjMlnHLCGTOp7+CdfzEhd80KqKBxifMb7fsHkNWxi9TWjLNCSyXmQVO
+jOVDDqtkmseN4ZDk2aZ5knHqaHMSqlHeh2Z3q7Qbn70rd1c78c16iXUDjVi6Nku
4RuESbttyuO2lZnGp8eXsxcDo/qc5cV3sqDeU3x/iR/3eL+NIcN1CgOCK8G6zY4W
Rf2zYw5LCgHGdTgCg0yOLCp7qZNU0BRuAg7PQ1IIzv8cvROgGXaL7iZ9b/SPThaB
Qt4nllgxT0T6wU4hjx5jRWtcmpri1U3zRe9d8XVfyMoHBLEFRcpxEqFWdiTH5mlF
iObMsSI0jIHpLUYzBvBacRoeauc8dANRtrqZN4/qVg1UlPCEWBiBoxSxJoF+qVUC
h6FzsLPM2cuLzkIB7OPL4BMIp6pbK3umaMVcsNVHEuMqBtj4uqENMFrqtcaSLTLE
WS6rrPV3tvPvtb5o3p9QXPCD3CdYPw9GplcGTTt4rUQd1Xz3rGy/HMh+t9834cQJ
FfFNkI+FVjt2H5tv+crGyo6tWWNnl+Xl/TnEFjY3F2JCGX9LNAAWEHCygniNmeAb
E2RZFPSK35M3WvEpdD1LGCy8YhTpHOXYeHdMvJQrMUb8M+shTgqM1cK7vAO13g96
vxGbJpaK1ATI/+7622P2fq73dwxVXYAyZPnSr5OTKFvsBImb+z0Typ0SPtjDJafP
2yyZmlooifMarm05cCLXtDk8jGhx8Ro9K8jmZBLAIFwwtajq2AVFp/eH8CFrgEAa
xjl2FPu8FQ929/TdDETtXjonfxJ7FSRmK6AgZxUM56RMRxQJG89thrh9fo6Q4Uns
9RS3MBde8pyvo7MrvStmmSIpdUUMRhINUlZ9pwCSaB9UAnoXMdonjnDJY/1Xm+E4
SFoFlzA59mb5SbjKag/N4yu5YY7UDg9jfkvwiglpy3iYvZKM/k6Rv3ngCrIgpwiO
tCVFKQsTolEWiQO07VQDfeoWRhVzm5jeLWJQqMWVhQaFqqs+4+2LluhFH3kqT5XO
eu147LALlWPL5QVMx/VZjMpx6sFkxa+G9D/DcbgfMxDTtCClQLefgvl3roVsTeEX
Yy+R2zGqaozDQIqkOuxEZHZX4yAl73IXwZ2oaFHRpBITV653c8VtQZ+TRsvZoTNT
OJY9f8ZFRtuuMQNlnmg1QVMkHXiRjZtUEyv7lbqKblLDD7bj8+5pTwdI95k6cOAj
Jf7feerQGP9vsHertaZAgGi50OWVvdqOZt+/s38lIOYtghQm/N/x2Vk26tZrSLbn
0ixfcqpbSMiDWeqNpj+GBKN7+WiRrv8kBEKBv294OOWFrd6q0v7fucmSrqcPffYv
3+PIRt6qKLpUstG//ZwqOTW3IJSVo6y6O5OtAGmfyg6SGHjvs6uPyyk6ytkz03Cy
i7R8CN4lCwMigFZMUbmlU3/kgAYDiuiMen0+g/oMc+XBsfQu3NtifeQDAEWVaX/U
M3+69JEwMTdDxZGM7RHjxhFCAK1dDvNn+kP5qJro6O0lew+iLDRzdAjy8xU0XokG
hp7t/r8E6vpGRANJJ9LhtKqwXYKx+7jm23LDrWldYRq31FYymxPGoMYroXB+VHRG
cfNYKBJFQ6QyMlkQxrDs1+bfdSpMtPU2Jy7ZwBY3HDuAvF8PJcQmhp6K6y9qec4z
IN3F/kOrS+Lzoaadxa8Al9JcF3TyqTSWj0bBlMLXv9Zq12H9iVRowzzmbYaIjeP2
X4oVf3Tzcp7fFwWIvahiZaa8mw5iROzt8P6AxU36SXQqHb7wTSZ7qNQLkYZiBa2y
QYE+zZjut+HC8qqgqizyJ0JXjFOkx6Vz5rmcznnZcDy8r38jEGfPnUHYmY9K8/+d
Ll1DfosKN1GwzyfM7+1cTQvjxyeLysJvWmc3wFyPsOaZi8/EqGP3K5bqNYrK8CxE
qutaPca7GdyLrE/beXAJEJOaAoyjw5GbQ4Wj4IsOUSyKTA/EIwRgtgE517N8XsMz
XAGdegnJWRpl/ANpzV60dIzNnuVjHsj/Ne3uu5grffrgSJof7yVXw2v3EW/+wxuF
RYeh6YCm1F+EklGYcIjzD2YBmjnEENadziLXpL4KwlhqBNwHTu+EJETVEIW+xDLW
hzw94ICe3O1DK3Og+q7P+e/FqufQoqfo8P61QHUY3TL/C+TVoAfyAExl30XIxdgC
kKgDB2Tx1RTJlgh95HWsA65xeYkiBBCERwnhYJT3+rIrRNxxSvBH/SLYYigPiDaH
6LfYcN4gasgWmLRJKG1UOIVnVv+rvvKBOK35NySN+qUQnDTmLA+A2Ff3adopf3Wt
sw8V1FEFNE87HAFW1SVrOgv/1DOwiOIHwzLzU0wGL3P88yWPDMK7teLTgTZhnvUd
D7BzqHrOBcRebMjTdOCzUxlQlKmLLHHv/jKCwtLw/6NHWrecuHQnYjlhJlRAZEah
bDYDYWI4nzefb/M/tbfeLiEUhaN87fFFHAF1Zd4SZFlgIwbMakQ1rFKR0oOIAcFH
Z/12MXhH9Sv8iePxyOLwiBTtJ8zAPbk+Zqy4zXss6cRp+18H+1sewxsjZrgtdYeU
A67hsxz1dLzvoauA5nKZ6lOgcPNiNK69G5mcX2CuQHeH/tL/opcX9AFYTDz60tHY
PaVSRqk65+WIXXqNkZIpg5A0s3HeuFft4SaMn26ElP6LDH8zJn6xPTRhxF5BHZD8
TDV9pGsC/Aj5HupDZcT+fme8TY1oLVgrJSEa6PKZv8MDoYEZ2wn8rPt5DRW2gXJy
oFzJ+ajACUmLv10W78jgGDdfuCtB3LaQamTUwBDpZzexAe+giCTae4m2V7S0emov
prVAu+Jmwk75ghB0AhBLro76KG4d0dmtkiOf9bL4fg6Uab3Jtw/QmyY47DTaofBh
SrtAr2d2P90G+YBM4dMNcawy9lUMotJCbCB9PbGygpt7m/3UEnyVd4eHTUDQSfG1
0dWh3ambIFXaClIJKYGJeyOJRo7z4jub9WbnvuS2qpt/wAVOJ1GOnMhm/6gkneZn
Wv5AQyNcJ8zdzB/mRHcxWxlCtD8BQciVshl53kIMlt6uT3qfAWm306dLhDQQSZ5E
DqlIzHALUIw3lF27pJU2tDxdBaz361kjmiHl++LHmQKA6D59GCKvvvo7ueTowZ1A
SWKrSxyr97+qx6pFAptSvxNr34WyfNhcBl3dEGPlWm2z+9RiSovX1Ti0V1894xbV
FQI+Ms03MWilgwC4rJS+U5zsu1CIBXtr7KbyPH+ww3sIIFxF4J0DVakVarVVqZn6
XS5AAN10VuWrwASV3iPrR7YT350lgb7tEzcOvFlbrucrU+qa6RU/PDZztdLgVJfL
OEbzZsK2vGNxMwq3jtCF8t9jLcz4DmQp2mraPo1oT5J/eLPF0QkAnbbOHXiAG2sH
M9GhALokJ/ct35m61bM4sow2aIMlSLh9Cfy48IrvOHFDbkzFnaxwkA593n+SZk92
Dl5mYG/upOIiKa2Oce5k74oieupKJSWbmOjXb6Y456rYFHJQu0rz/AGssQscfpLc
+Ujxby8QiC1mkA7RR2uiimeG0af7SXZAZtva2L8PA6DpI2YxouyVLv5DgxujhpPM
WtMeYAdLX9LYVCn/Wgy6RVdezNAoh9iX6PC2DLQsFIuWxou9TR0iVubfH1FsXrTM
TY58QvuIzgNvGUW938shZKQHQeSX5HVe0bZFobF7zwO1/tp9DR3fAcS4zhhpO2yr
ukQI3t+7g0GRD+gZYgfq+678rBPVizLfNZxLj32/PqQ0DtZqc5+ESwuKf3HOTatk
TswnMA3j1wgf/hRfPEWKEXFbvwTxq2Iukk0xRuXkCJrTqscShQ9B6+wlpqDbyCdD
DaubdsY260gI5UVplW3b8MKzSjB46sHoVbIHzosJQzPlZO34/yt0vs7zwcCN1kne
2ruv/tN9N90A1uZcjY0/erjunn+gCfYoH0s3gKCkVbs17UCQJVEKX3btaQSn9gZ1
q37gJv39x1jk6NrAmJyCZ0xJ5Kfl3Pwu5Jlva9zucnsCFZv1pZQHs21EETkopyUQ
n6BuHNLTYaLjC74oiHNmBM3ReGLts4HIb50roBedoj0jd4FyhWiXB0tZ9uAz33pL
Xt4TmW+WDN2ewAlUNYZ7OYaZ0i//yUv5AJmJ7GX4W+Nk9Gaaw+feu0sRdvRr5xxh
s9649F/CZL/fq+ssHkcfIJo3HF+2P9cM2yfTBgd3DtJrwnBb20rCWCrtJP/4bcfo
hGZ2+94eXkZUu6BO0BFYHCLHlMNvmPYyWJ3/W6p+aFuOp6M0EtQZKZ5f9HwzEZ39
ZqmbhZ5Wb7daYMapCw8YBTiKR+v/duxlv6te47QdAHdwVg5FF50AGnF+v7SeZAG9
IJ+fWpWA8Q0LUdg2uRgRkUSnh0g1QFeYmpC/r/r2tUkD7Ve1b9uWZVWhuD94WYBD
Sv2BvFhlrhmm7ndrMLDJFEXGOdv111yQBHznuqkT0Lum3IGCiXYSxVo3gx1LDYIf
rTRhyJyVBwKstPkxFAoOyOKvHrYtv8FK6LYHRadLRdOu2wAXwJYDVGI9VIHYjtMD
e3RXAg4winsRYP6avXtlIXIvrdAD7LPuq4JYveKRB7zwvdzcJTP9yQ0imfNJNtVS
2AoC4Xc38TM0DsNjj/Y5DOKMjg1q1Hnh+18HZfgLfkOUmIJbltXZ9TeV+nGRHxSS
D6BLUl1duzNYgbp8RLnjoF1DrQWGaZtp/oQqCR6o8pqOad+Fvf60iveBwBeEicLv
HnVzBOKNRTYrTr7peBhLRKi2b8/ZGbyUXlFV6t3rPW5SVhDUbDIFaj+hb0YkWQF1
HTp1u5qzhXOX7hbx37lw7QO7dmdKSmowW7KDOp0b795i3oouYKTgVtJDq5JTS+MV
FXm/ElKB+WRYfK3O3POA2TNn/Knx07+AB4zYpMH+kUhObDlwO5zVeu07iKoPaWwh
HDoMHrUh+seTMVHN21g44RCPhcaoyAXKsnG3xXeami3Iy1dxjCxp7hZaN/0BtdEu
LudVhZ8LMx0fhzvwNUPATMJ3xjM3DYVU1e3pL2xmsO+v53xg1yrYT+PBbtohvWx9
ezVAuKn/4WvxhOESoBBcuNlF1XeZ20oCyKc4oTxYv4WNXXIeaPzQtusA24XfIdtS
s4mUNB/uLwHA4TUb8O5+Dl6dWwCMcvTO5qFaOQ/zsi7ET/f/v0OUCokzKgceeoj1
g88Az4Pub8uFTw0TezVtt7Dj7ifydJT233nqWBGtG8eL4+X1ioRhMiBrIyHPrNvt
Dx7ECVBQXXSInJTVHiTj3u+CVjXTtMfMmJvhTS4LpgM2/7QP5/zYFfES+m0dIPy7
XPhZe8U9CTdgOK8maQx/tdDMqofmObKeS48AxWnR4GUe/i82MF7X4Fab4b4olB3c
2aENNBlXSnScwvTBYC27xkSFb2stgtGxwbxX28BcH/l/kbhB4qaf5LMEWQP06TPw
D+0eJe6Qx09fbw9pj1+VNEYMbjF04CMfR8kVsw0htnh7FSrIYvaIaP2KQWL13XxR
X/n0zriXZ+DzvTQslrE7bugKcul8CGKSDqeZLLm3VenC3exV5NkcwKTGN9yUJ8dr
ayWS9wmiHfnPxntqISFj3CPlgbV49FA3lYKgVo6oa6O6yviaCq4JLBO9XNkvGJVN
uYjCubbZYmcyANLdfkYPQbdkoXrgRhXg8vo/Ldy+uXVyYHer2QOsTU+3tx85qE0/
Y9lOg16HYlxXi57fXS6WxrJmm0S/kZC0UdJPfqDMMQX8QBUYW7YEFnC7u0Vm5Nxv
F5pVjlzAyOa+e616+wLwoW0UsaSv3Izh9Vj2h7DxT4mxxgZp4vhlBDGJPjlTM9uN
BVr6aZy8YvNuysZaD1vXGngnFWooUr09F47fUuMS3jxUgTBuTC26xra7CFzzKks9
hjHp83io8jJGEOu+BQlpByb4I4/cTspYUORArF2l1YwGe/DDPPF3cXbJ3BewNFAD
EeGT7Iu6pfx6RIcA7GfXg3i9t8RWzdlIX8ZdgaksddMNpD0gZ56sBKk6aw5ZOiLc
U7JBu5DhA/CGkBOhj0WBPfnu0bRk2Oxt7ztVqgQVORljA95DKKTxz2m4gJemvAHs
NMiq5veErwzIyV9D+eorOzHY6ZxxlAG1OtHA21DlIAMbK7VwmHFl9S9/2aYeXzLK
l8k8QsDVrb4YVgWvSO3Gpdzlw6jKUVN8LjR5nXzqdZmpLGE25yeGeEqxbi5yQzz6
V8t8cda+u3kLlN7zt5RAbArRhgXffipfVGJ9QHMS4ejVuYLdTXIuGDi1V8w/9KYV
oLbcAmBxgUO+kMblOhic7aLFjLm5CSTFAWTAr1l69nGowO5Ejt3LzVWiRTiOrZFX
uCHjyKxVamQIf7mPlXK1N74m8UoJI0bJtYRTtqdSBYkfX2FXoh5pEZen325vyNVD
QgIh7lc+jXu77KBYbGK6co2IOX/fwa2jQ0X50kp1pRnKZoNZ6NughjRaU7xTgWAf
O2qmyKw4XceGJcERFsnWbWNGt+cawUig9q5r7hOdwW9Zkpe+a4GIFza5NSNTUMw5
9RerCfHeCoCg8aUQhpze8iV6PcZ7Ye9NlPISa/CuYIqAd1jyVNWahPCCTPn/SbNp
NGl010aVvm4WTVvX4hm0kYjaylS+nZKs5OQUcQammsyWfFeLnIbcjmrCVdp5jguf
/qBLal07/IUp2VHL1L5tTFq1jNAJ5WGqdLcKyWo5+MjwEhICHClCi9Z5Z0GsPhcw
nJwXE36owpdxlZEJFJicEIxi+v2sFivOvQQEStVjrYGlnZ3G9NDRfCZOzKAq+sSG
yBgyYCtMjC5GwuXVAxCOfT6nEbM6fVwQCamG8sP5pv3w25bC8RUibKH2DnydIJwo
y8z7J28rVn5IMQNX4YXhOJbD10FexwDbgTpfJvOC/5scqxSIIIdxXGFDLTSgUNxb
qFISDEQMa64JjK9Hf0VUZHLQQ0+dyp4duoUkZQomMf2xFHp+PpWG1UKxP/Ne/ftO
eRxqO8bAry1tsy2NMdIxqFd7pvJIL9hcZebpEDlRstU5jPPLg9N2MO1ihVhnjh5x
OausLybSUYuGdxZ+RW1MYdioADgm3Y6eNtqj4/s59bUO6x61Xul5T+k7VA1DeTOe
IW4WBAtve9msu+4zABede4YRXwX3iPxuOeLgIt6mKJe4ohg+qc3UUGQ0ZxSJW9+n
g4185lb8r4k+YuSbMRsf1MnIozhmzbcNjCxJAuwik5lQrDk5e7RXCQpe2atj8FQR
UDAzANeKHHvHE6ULhCn1tmI8WqFRGFFDQ5k+egm/05ggmukgE/cuL/XJNi/O05Y7
L5xDnnpF82X+BRfgXNDfEedB72cvAO9Ox3dzp2hohgXlXKNx9MJFD2p8yy7N4UTA
gphSMbirlInC1gOKkF4eob7hrHdjs2aO3PX32O/oO4vzAWdrwWlnGT4hoPGxpKXM
0k7fCEdlKgu4kwbpB6A63oYx1cwWMqdWy0zuP+sbjdM0S8C1kw6xq6Hl7T3F0LDk
i3Tt4oRXRmxwrB4P1v8w8bLE/iphcxI9ycENnT8vK+mKOD8xMJyEVqJrA7gIU2A3
IfZWV9fJ2UM/gfq7q5anSS+tmxXd+dZeuIkk0WLeNBATqg3OkrczeFPJwf2Zj+bc
8P+AWpC17Y4AG3So8J3zmfknXnzF5SZKQusmSV55IsPWwg72o5aqIflXhd/YUU9z
V5jqp24LXr5hvxJfbJ9sc4K202E9UYMimzTe9mIX+EoaUTemv9CS9Q393mEv/YUo
wVXISe8YhoXvrg/mS2O27pAjwaHPo7NLl9adnm/b4Qonko/j8Gy5I1FvrTJ9Jtk+
RC3Hxv0mXHwk/pMkdse57PoSdwX0C4uyd5dipeY8AhaRViBSPs4pBt6lZhZ34C1p
+Is+5d2v9AUvgF5gvsVeyNaDgMFmhyKP8EpZe0ckyFp/yDxWzm9ZnYRQWMVq++nJ
GpXkwlfiLVlQhLnk6xZ64Jj+X/fmIkgJW3TFU0f040LKbVmjRmPrcsFUpVKio7vG
qdVF60Ju2Ke81fCHDYwscCpO3CzeDyZlVhB1AkR0GaCDCvbSxcyd8ak+KOGXkR2z
9RDUHAkKiKfE+XA8m5kCdgl6a906zWx9bZI39kBYwnjBz8Yqq1EoAmgqquyYLIc5
nONbmVm60q1sulhec+93BRmI4dhChQfTSkoHEdmmz/57neIJ+XpzAXNpm943GNiD
sxT7zcW3zkAEdisjbg8IGunx20Xga4asiBcbphhVwIrJ9KRKRbRq7B52EpB5uWXe
BxwRO5kn+0vw7orK+eKN8GQcF/d+xlQtRDxx5ArNGyM7XxNsSszYBeynfqA4xrJm
sookWf9XrPKEf1Krri3Oi0A9C9lJLyh5jC9yxOzdx1lXPVKS7Iw6FvflZUEEE7MA
r9htb3pcACpnLimzBAM0hR2gvQ4Pi7PWm1UbUI96tGG94apOrq+qVgk1lpd2Cz2u
8iAJl+EgoZaAnzSMmXPAsY5QMMq3ltr79VIHqJQUlMB4oWJ6Vo1T0jPWN7GVCEoS
OUQ1hKxKoRGXq+Ox9Xh74hTBaEYLx8AyjgixOmTl59pe7WWADtOsdi+aJHkCpwk+
HXGssDbmYGCTpPNHP5WF/pLIBtef8B3AlRlZ0JJkCZgLSdXMZlPF8aNZGqbgaTqX
W6J7zAOLwA3+w/eUb9QiKC00DpsApt393xddvFsTZCDpaiylFhDA7LWRySf1Xc9L
m3AvQKE+nfEwbEKebsW0mZWzkuVAdBitK5tQrJpNHiNDkBYEOR45+xQ5WrTV3RYX
Qo0DQhWyGVBG62urBg+wdu2v1JcwfAcQ/HWRbQ6N6SjsY0cows5BDJPYXpXCTl5b
3GtFpuIDENlwW1kBlTIgJmOST45tlWh56TVh7F6k82odTKs1ecU7SFC/Y8/cjby7
YcIOIbqM/Rna8x/y5ynPWxD98GAGbRmTMYxjJ+OyzRes77TPK1+HoSJ4E98maJMV
HgfFcx1hQQvkbTBZI2w5xB502f6ppDhNL/jGgkUvnycq6i23BFupa627wFSABl4R
W6JvNdJyeJkYru1/MsPoS8edkov270zmX4iw2u+33UGjy6156rJ6QFvP1bCWe1yB
RTd1ocssLjNjbjYIhVNzRtw+X64bqgq+l/9pPq+/qdtpnRWX8edVSRL771r/dlWi
1M60hnlOvn/Ybduq8IGluLQJSpEI2+nL6c4CMdhtTUUx3Z4nUphWy1lQ+wSiA/1i
U3eh2Cp739vIbMH5YKM8vYuv4ZnmmhRXeLgqm8BvRCJ8FJ1Wlr9m7eYf1Y2Ju8zQ
W4n/kVG4qc4+Ho3VqZBp5VFHVOWOiTwkAPJ8QFam1ZjJTAMBxFSX82RrAfLvFRaG
ta8h5PqhjameKebuJdJ9Zw2qVaIAwCQHkGJwZ72V4IQkwOrv+ZBgasWnB5CAcybB
WVEgqb25GxwhsFoSNOMDRAs1LwWXjil+aC/uy5nrEilMVpEO2CDY38JC0wU0c2UH
tIg4HeZcVcBR+7+ofqpclD9DK6egKyk+58s2fPRIwYk+y96+HGv1mSTQB0RpVJX4
D7FMq3DSc7hLnmu3B6e4m8Fiut+qwKB7XqK6hsXBBQ+rJ0aPk2ax0Yt+1hcscR+Q
B54KyWl4fxKtBMK0o+4FRP6ESSA5gFQ70urH9a0L+i+PF6pjAlMN+E3ALccefQ12
8rwDZOOpVzD8cjksrRQSnjN8jtDbir4xqdX3OI6Lr3XVBsybIeZv20CXvbUPxvGd
2wBbrFuHi5pkdwcsobmF3hxjgM4ovL05EqXKYCpIk7/UhNGLWQbK6KEvY0LwLPfv
+ZB/JxDOGz0j3PWugis9ONJ5qWgauilED3yabXTNilSFxX6iuzIa2Zl/dXkfQ8dG
9/FSi1V00JEvYfZmwK1+KFItpc/ib0NTrpbKFtktXMJ5sNJMy4dPBro+ksfeKTQL
f3fVm0AmzEPxxRcdPBgE+HY3JAZ01ZC31yBossdwkX8zFDK3ZttWNPmCYvy+nnyw
6j+eYw+cU672imNPAHKGNDptkFUkV4M/SOz27AP6TBcvIlK27KDw4kr7b3Oubd5S
zl4Rx8wtZA11LEssgUfU7jru/7tqReT0qo2cUxQIQodGABJtlWbCMcgGkCB03Fte
S9Ni0JwGp4IkoyBG3bsTncZo8Fpzdxe16kSTsnt3624EE/ZfGqn6EZ/KYfCfcs1v
ezrENKcF0dZYnWjdgjkQCTKJA119D9xcx1bevZTvCxp8ylLxco1vTWR+pZDqIoRx
PkNcpQ36IrEpuFh19CV1Gf/Lbuds2/Ow0nTJk6p7HGHi5ZMrlFXdcJYY7eGkjGxl
1Hlfa6/5Pyc6/bVQNq+KvieesWCQhXAKxMI86z+J806qHNsUlvjscSaJ5pJLSyUk
1pQAf16K+6sb/VDARaEYR69hpglrsNtcuQHv01UETrkFk3otxrhm2xG6Q8PmTNks
3Q+7VqUzx4CW5Isxq7BqmfmjKYVrh/8K5PZDpfj1jrQYzmNVZ0nDZPY2ZJD4IwJl
+61P2Y+Y8QwRBJLd4cmkvVmHgsENAjBJjC6TiRvu/6u9tXsgJKXDgLmAJvqK9Bw6
3YoSsS0ieQt7Ad8jkmkoF28J69TwEANK5/j/iOqZR5Dd7gtLA9OxPyriMepFhbUO
snWyGCqwc32P1tqKEpKZ2aNlTQ9qlisFInGSGAV1xhw3RmZ0wnaDVMYhjwFeOFP7
nCy3VhRNbty4u2R3w3loZ0SoPCvX5zSxh442hhVw0HirGX+ZKftihNDlq12hpdNw
ic4lGdE4wcLfUecfcfEmitdq0NFN8Wr85C3iTdynyMDgMaLT1K4qPg7rTL225mye
3BYRQOnMmS5B7uue/mEzXDzskPWRxLnIWyz3fBb07iP3tvzXiOy96JClJQbZ5NkW
MqxtD6nwKg+X0QLtayl11Yl5GGXRaRFP13sMGpVHtsdIVOoHrFI51jpJs23/bD+n
bzqTSFDec42vyPpRuXbrYB5OOnhHs4vSO8rnwa5LD7RhZUUdIglLTBhhs0btmW6M
NVN3kti1Y8N1WrZnNYdzsLoAR5w11fQIV8dEEKy4pl2+91ic+RH8KcDVIEPpj4sy
kP1oghs6RN7kJ0wRXsIzbgaa4tRm24b6ePEwHSxBd7UIxJIDPclkW9j8RmuXRJ0g
zF0OggQIgJQHNsqc/1n+etVBGagb3GiZMXfLEwJXbvy2tNyQv6Ys/tR3PzwRH/5V
voHqBNXPXOm/k/JQDYfYg5nv7GjxiRtKDAyp0DJUVZdVsPGlwVRNr1q5gLibv8HI
rvhpHqyigPFyLCUOZqWXVCgQZaPxLB+hmyzWnmFJDPMpj+C5nYYrK4QQZrK3PJOk
Z2KYdlyYnQd2Qco6h44RJocR3S/5jNZphi32a6pfWTVE/Z8tvGrMoY8Yoc/Bxl/e
DPniGLdn0JKhdTjKxvNQsDVwp+zoOvrcRJTk9TrCmwB7aVOPvrUfK6gsH9IL8fXM
KMTtSwa5p0Xc9CEpkt8pxl6M1/CNmTcVi2FiUuuFB1QYdKG9zPbS8D9AUN1EkCiW
r2FVwWX4//QcqY27yXVzTlcE5qNhHak0rI8Vbo3aNfQJcIKIzIwvnufZD/ZfiHZB
kAjNgL5B/Bs2/KLAnMr8UHA6hulfUpeKNSYwUy+nuMCQVWSoJGfkaENKFvJ+PvRT
yrOo88hke1wM2TNPH6uSAqKSIXOYPGwQZ7HVLhEPl0kWLlgvTKQqEMMFK2oaSzAS
6lWc+HFLd//rz/DcT4X1PkOCJk6QMhEa2qa1DeYmbzEEw7m7dk70mBrUGWmwwcYb
xJyC1ZrrjDsierB6oc/IZY5LhXemz0UXkwnz/7a37B5f+3Vg2lw62J6q2QoAwLuz
dHDQP+zpHJWnwLDKReWYvq15IlJHMjA91W2ISNcf0LpBZorPLPteYI2eb6UyXOH4
dSF/6Khc02cS6XMfZ1R5XFVUdkmfEn5lXD9utDdBNXrrd5qld0bHjH0yCOlMcf+Z
1JsmsnYda5v8vw5KyeX5p1O58v2weom1bf5FMZzRirweqXdsxsbWZ6HEBTMYtlVz
rlB3tc0VMcgCrAE3/p/unRWY6FjhVdqJKU7TTEDwwctdf9RNn5JIOV3BaSODeqpc
1oAddDlR0FdyZobjhwSpkGSCpMBhAUmDxadIXQq5ucfzrlC4lMwAE5IJoq/yfozc
qDkXwsVw+CgPttRrCILppqezB68gK3Q2m1fgPIAlPdxnEUWimddv14e1+YXpegpR
H07gIdzQHMUbd9lNoDlafuBZUWhYDxA34gOE6YLkLs6ulQNdcWLFRdTys7mKNBa+
9+KttCDZBC5WtVg8/gIKADMLuBHF4zMEnU7QVyoOkyrWcZZAJB5PBuq0OgrIBoyq
PD0L34zSAECDhiEHxkSau4HgVexU1wB8xoIoWx3r1Y/W16SMjnF3hToQAT7izIoQ
+CPR9SGQn0bkDp5LhtaOukuuffepA6whKva1rwS7pG/anHru6bDbh6zsDfoiZJYf
p144UTosDPP9fNRUOW16zw2ApcCwv2scFe209RNGVhW4n/e8ZHZAtKWb+YS8JpEj
atrwo/sLwmaqbHhegMQcLSv5fj0dDBOfy+DWFpzInJ37UvnDTB2E9TzsOyDE56EF
t467RpDwqnpnBY0PaPJ71K8PNm+TEJdP07QULWNr0hPEfyD166FVKY8YJxdOJ3S/
jRdoz3O9pEocVB72Mx5QVZMSEl3f7gSpYYQO/8Q28EAqhWLMhNnSRJQ2/I8SZ+N+
b7khERG1+hvM3zGzikOzY5mYAO5giBiIytR0eg08WQQViAjlxy33f5AFhrxwErHd
IORRn246O3lUWPoSk2F2QNBIiXolfJgiJben9jj8OOLfVecYmb0RxB7VBQZclNfs
y+JRxPzi1x7LZUw067S4h7NKCrJ0PWIO66Omodd+Sw8/S6CRfZOoxTt4YilWKgLl
O5/C7N+SoKogqj/SFYngNEPJJhx2BqcSkimSJEIE8o3aNhEONpbfNuBEIiMPMqUy
hUu/lpjjFn1nnt1c+MatHEjwC/71GXfVY+C6I6LAPD7OBKrdRYWy0nTdGdpmKdxv
vEZ3STEtVsspnFKAvL6+Zpdvfp3utiCE8hRsy7o5OQ3uCK1UH6ej83PkRoGWTP1J
JW/xJbn+GA7ZWfaUuAW05By0nDTkA+gq7YmL/48PXdPxfNsW8UFYOaVCFMOAyw7Q
KCTsND1gZbD86aykuLNDyhGCbyu1ttmq5moZpUp4v9G2kudqBcNlQ9YQMjGB5ml3
bK8joNW8IiQIfjC9bo6SqxaLA24O90QKFrYrsWZYHjLBP1fhIRdDzBDQUnhC+22r
M2Yqw6A04EUNgFk0pvYFPfJfvElTXPSSbJVOj3AFURnyE/Q4MYR7PeIUR/8suqgn
aU+ypVWX4uHoGV/j8Ib91BzayAJ4wsXR3BeOoHwLCTna+S5UpsH3xZlLo5jBbt7O
fnq3GbtQU1FWAqMFCGK+5bcQP+ETRzYaL2xAVLH/8ARvPTBXEParKQwEAKUOas4R
o3ag116gK25gW0qrF+1OoDbYiB98TvOyc9kgAJOqPP0W2Os3ZHSc6FiypAng+u1h
peFCeCZAXydljrMHCw5W82qZdL7yRuzl4+v25PMwEV2rG9SsodnrEjHtEk6APFWd
gNhjHhJx5Xv34ChEe4wVR5ie715orAoGmgd3dJtt9xGXnIvb5JhFLvOPfW9k7dxC
lWNVLjJLSRby/zmIPJzAcDi6yVMSG8tiMmF+kCvOjlyYAweJ56JhJfHyEP+9bCt0
vYQDTxMMP0RCntdL6O5sKkRK1ZpiP9CxwNWfamQouUGQt6GZ5ZVMjRtPAuotxXsC
2uBPwzwx+wKdSsehlAa44r27Y3BSfxKCbf3MQBtOM3p/EkSaQeOdhxeJVr7Qyvde
e8y6yCDKSC8a5s6gtg/rogp6mFXiWKpJwOVIYs8fUrNqVcVWMPa3b8M1hdMI31Xx
BtVloHb+bm9bULZrqV+bZkWQRBmJtdP4ufjdEsQHpelCP9BLuYJ7RZIiPAZHsQUX
y9OgnPH1AoXSrvRFQ8HzoncDcLe25aeBpU/2cvaKg6A5rciew2PXXC8nFld1N6TS
+/4y/PApfHrUTDosOjk6hDzSdT2+cdM2gOue32Fn6MoUz0aKbnvIz2Mg533KxsP1
Qn2tCF9lH4A68afNrxOUeHjzulsWKYjJo2PY8hDrSdAWbVZGpPgU1Cv+6/rx7jW2
ojuVIATtwb87WhYveUsabU5aK5WeYm/FMcP0AlQ2sKKYiiSvVrUygwxzzvII5R9D
MwxyWw2bzCmFpi/O0Xn7FZ3TZUT/ruf1Uzinq0m+4q+Snvw3PXhMJ8Kj2r/QHGS9
PchwGCe90C+HmKd8X5jdP3MrQp3g/rvspDANVvu8JI/P849CaV9toGElZ62o7SRi
hFKHcwjdkh1OM8fo9ToR+RUNfQMMCLxJsQW7Wo2mJ+/O0BN6dhlECAwqDAzXag5V
ZDcQ+w/JpgPnEgkbUCQv0WmDPEZM2vVYUNdkQn+L9H5MbYnj3cVOUHYiqYM1TQfN
LG5S5K6WdZOlJoU27WsEcUV15Ay/ZZKASxJfedVcvSowWU4Q1DhmNgkLp8SS9dPB
CTgSjDsX7OOcMiv9PZNezNfBs99HbFLQGW0yvnfLEvW0KL2ijL6ufbaScZl41r+D
XbkYJ8/zLdDpIjTJterdUWLAhE+wyy+xz00Ya7Z82q3lhsFqv2c0hezHpIpEG/h+
+RVbhWUKr9b/DwElIP7EOUvKYm8DwTLWf7TjcSX8wnocoKXVVAysdhlrEYQMHoE+
EjIYxbD6lUXkE57guisy769Z5mqjwJUAIzCz68+rhyleJjbDRBYXIDKBC32YGyyn
0TN7Za9+nM5hp+hQK4MP627AUXtg7G/NFtEnA1WlwdiKL4Ec2XM8DkehbQQh/nEv
7pWVesXINKmbYBEnkFvKOYf7GI4p1Wik+yMOhRjX+KEavYV907eUL83tcrXDR6dQ
ZA+jSOzlLcl6/2RDzqfsaQIFgBMfUQAAti08oqQjS4/fYBkWDy0w49CSK+Grn7eE
LT9dZn63+REs3VXmNiHjVJIwnor+/epGKeEUC3f1zbbKKB5exETtgD74Q2rd0Hcb
D3uvvBPi6IBKysoaO2VeWTBQvB9zoaaRLCF6vg4miuSFzIoYufRGvuGzI2zP7+Kj
jz+3fnsEDj1GeTVZVHwfgR279lvvDTZOWVWRqo6UKMB7tkJyIhnQ3bzC5cGA+bGA
KUtdskUdIwcZfzefvxRh+AIcpf+7WcLW5fAMgj4XqueYa8eSjZwTa0IQUDeZPzHD
TFiGfo1OGXYuf/nB6j2rByr5Rt1bFBGkKsy/GE0aONT57fl8kj/7uSyMvVl9GQ6W
Aoc8m6kK9TmpEPjosqvR42kkT1NG6D2Vs3ToR7CJgP3DSeEA3fv9EecIwDOREks3
xq2aGRnaw8TDP5GYtj4bA1xWgVTHL4GV4VbvKDJfMLNo43vyNXMoCPJIOMPqU6Oa
d18RBRGwPi6QM3BN5Aogof/0aLe1ESF+EUvN6N2BBX4FONoVMwrdCdacku7VezsX
7WsaUet1V8eB2DUb0DlWP4AbDUIOhvYW1NigeA6G4SVYkW3Bff0GtJSmNNSW0ikM
ZUNpP+npF8xtgjCriTCl1+sxIh1aD/lAs78Xv+Bm8SMOSSup4L7F5+887Ogka0qZ
PEVsBMMd1FZw8dlmRl36iDywRzVHQz3DEa2hn0zhHDmObPI4Q3T0tIz+84KQ/GVx
1mtUMR/nAVvpBY/+r6XO5jMpbotHFJXMxCg6wvL8Y5jT5r29P2FtJs9vsEmaGMgz
zHTK9G/IRK0uaD0VcsosSpWmEskupbGDpeTyh1lLezMmN3NaW2xXKgWz6qVAkyBB
cUoYVfAAxwO8MUln1RGJ6hIP4GE5AXgGWXOgAmkuuEG/TZWl6SG+KBCUPrl8xWPP
dGFIYRZ9mOCtNz/yCqnfpVoSCUXQl/5jT4iQsDQOgixBqJWkE1jrvEED54oV5Cz8
M4NNaAJ4vfT1Pqe7Mhdgf8t8yrHYib1JI8QG2qgWyhegcX0bHHZusRy18J1BAcZD
CcRZ21amQgbbX5dmQgB537w6AMygxU0CNamuzbpSldbZI3IeCEHdCMsymZmsuheg
N6au5ndaTrjpLO7RX/9FWF8x3MfKEBSZpQbM2+qqMvWx1tOp8xlwrPlLRlIhwtD4
y/aj+GDgF0/781LKxXkzhhlKQSBxBfI8N646m52jQQ58CwFJbZguVo65+FK5VZI1
CRcoWmq2DLZmCnwNCZNJFZnYioVZTvUncJUG87CjWA3Q55baZdMYYkKWkSjPzaUA
wvMqEg6PVtXJhSohdrCLzgW8Q3Nlx70GssSIEW9N+92FEzN45wiEc4Yzi+h8ip1t
FpSPCZs7OZfizvU52P2dJb6VfqIgVHbG6+tntgpQr8Ge++lBn1oyCQDAAf5pm64m
9kHGJ1z4VvgM0dvO+VTZmUrLxAlz6NZlqL1X8OyMfH5PHVo+TFBqDRPb1vcgNPHN
XiN5c8K1nn77PoADqKGW4r255MrN0/RjQhnUXSTHqpdkX1j2s9vhcTIaQkJQyWkE
tcQ6q76uiN5lTIwvzD7MIeCF25wQb2QRwR1nEGuuKYrBmx/NLz8un/TN2pOwdV4a
1xJ7+uiQJWq9RSpKaSbPgS7mZ5L2p5XgA027Gb0qPrQMUDTREWSK6aI56EoY3My1
gaue0voz2uUHX/q94/PXP9gyq+29A0CkF3qmfk/tCZ0r6ZYrEhafTlvrMkLuwIVu
vgomtGNpYLYeAJa2dP8S//TwAh9MsNhLMQjUkteBf6X60pxNYgKUDA0yZYyZZ/mB
GvD1/VavmJfFp3b/7t06meuDWL8TDpYLRTf8mD1Z+DWtrymstPQSGMyGj9LmHcKt
zd823Cs+hpPfaA6cEARgVLDwK1gLfqV/pm1KLCDHbycBj2qE2Dxs4FnCw3vxRi26
4BdCNTID6j+d4PF5OnmLEQ5jUDurRv2vYI+As931kKZuGgaNSVyvZV3sdQcuO0mU
X00hl/X/l4cXCOMaFnfXRp/DfLFAFKYTm0AoxYYzGgOWOdJyF0G16WPG+RXEd+/G
wot1FsgGMNZTbHmsF4PepCDN774fvF06Wa/CQtEHSpxfSq2Q4/2BPYQdWvTTn/ix
d5tswRpQodbQoof9lt7x3CY0/JJhyn6rMTLFxQB2jnt8IlHu+BOkj0UfDWvo27EX
QR5yKRTfl7Wsjnl224WTzxrc5WSpL8YdRkHyFBqSCLQIPwck3skJ+QnKbZDFu2mt
6ynq2d06DJDnZILIYJhviPk/u6CaKqjzSOL11BzXEV33hjXZJxK9Grq9Hex45sIr
/UAkteoI4OCsZ9huYCT0oUa0fz0VsOHAgd1Dfuo/cnyutoFyzBHAdX0j4dV9UBgu
cM8lhCOE4YP20HCijAha0ADhrR4NV5sTYqpdjQuetUwWLnrer1vLKGbn0PRaQnZ1
ODoO3xwfD+6JudHAQmtsxDnWkjrAG6KNZHpSZWWSsoTjDYAfwRAjG3YHpteVczkC
fBgaUjcBJ5anI+8Kc3su48uan1nJyPvZxvQ6f1t3saQSvD3aVgOk6JThNZA6gKry
OaXov+pLTY3R6wQAofqK43rGe0YINSZSo/jzDTigVSW6RhDRR8+gZXNSR/PhZD66
RLmdvyBXOi3emaqG6tqFDM03MX7xFFfhG0JzipEMLBZFC114DxHYTvLKSE8zdAR5
Yr4qEFEmRGPSMg3FWtpEUatRwELfxMOuul3wNYhQXdbjLsMA7vhaJBhJVY1wkaqJ
v2C486ko0OY8OFMRZzo8VFnTdhpefVfa1/nv43M7N45/ahnRWGCas7BRjbkIgkLC
iiZ939mwVA9jwdrv9wF/6f5ZUByoTRsCZlJaeq1OOb4XUNhZytqg2NNVMASH3R51
lvpAJvfJ/DDRvoMiRMnzY0yih+cl7v+kszr2f/67jMGtJMi5+pWywXNL/74JvVQq
fhHbO6M8FLDVQ7EhUm/PoorWSjgSp9qzzicwxXprVLYJtndJ2qS9bOH+2MeDyBIF
jQ8S1wONuBe4mJOJ+NwM59VMZUSzY4+lgfvh4nR7qnhTBOyK6moBHtMZTMarUFuO
Opbs6WDUJPGSJlnWPqu0nNp+TlMqEb9TNZK0WuV0xnuVBq2qibKxc5nEIflV5cfn
T9Xl7PO0a1U/y9EkcrEApmaJKGBCVL3D3azOvRUTD9+Xah7uFui+5kfwZRoOsMuQ
F1HxvlEBfLQvP7JRYxFZH86+aHeoESirU46dGwxpX4fUwT548gWjl8MKt5wgzsr6
n9yCl00EfK/k7FOTw++sB7MzjjYkDnoPgJmkDvsLqGBCDUWAaYkpMujmMvuKPB/5
V+VnuGFW0pIlucuhTzVmFgFmw91jYvRBq/sLCtcqlx7T8Sv0Ee8Blic4C6U9UWQf
lGTZOlwqXbB/3+kiNZ6T34F0lR5Q+pTwto8V7iBexY+2GNSIYptMhXymrM7PSzy7
vUf09cUfYcGURglS5WGHcRqrZVnzdZ7XDn4qyUlMMzm6AvbFXj6m4mS1+p+epIPy
+akML22eS9FjlckbIAxxWr4lBSKir6axa3LxB6goNZsrzpiVLKltltWtXhbpilZ8
FSysskvY6y5YiQYjw8ktVdhLkG8WjNGolQfESNV00yEBiCvhdLHFU2CKn3aVV3Mq
z4O6PoLWLkgKUDNndWXJv2qgkC+YPbWBECh7DqUq3B4ykca2dyjNfrirVf5BPzDw
gOPP21j62lw3JDOFIOVR5G6XM+MFrKw6YC1medgCgoP91VHGMe1cxj3ogJvo6Axf
gHsKg4ti5fxhurRId9LtrJhRezhE74+usvEXNrFPjAA5TS9DcjDMT7tEms/a7767
kCPfNePANYa2QXDRSVkINQgkIS/7sBRTTvlPH2yrJUnH5+1uU5pTsCSjg6MVPmxr
w/Qcl+3VePJBtkZ2YJ1SGzXsRqVlOKuXzDvkwOLJC4pol7LA7akOrkA8kctrFaDe
0YfvQGoijFtjZRUoO3vVsX43lpTbQ6sOSqOLWcU8QIfZ3UaSIr089XYm5xbixLVv
gMft+ceWkqoNG9+bpyVPMAu1WxuTgYacW8Lr+cSjxELj5aCy7eYKljks5ziaczfK
mosZIfJ4pA9FG+tBoAGKfJbYAAgaSLquzoWa1VizRBdGEC/6u9AYaCmWykgodms9
KME5u5Lh8ShEeuu7AinUKcybWXDV7u0q4lnkKqOHfrWeGfzqj0OJmwWbn5q66a2l
nUfElTskC09Zule5NY0+hfd0UnkmaB/GIqhSjFY1hh+XPkRZPZIGr++a+dbnG1og
FHMjXBc27/nReG5SKdD1QlPjWKQRmFEUATqS7nhwhOozGzhjLeenJ8gjEHeIgAYn
xdIHdVcw4kv7TkPdtYMBA50tsN0ifo64ZU/KNY8wqFyO+sWSSEotgO4xr3OesSTH
uQIdN3ExDBuj5ec/kAyixrxr+rQ8nQjj8FEgUiXu+z0LfNukj2pr2SnY9gplu/hI
tZ0Bo/86ke5uG74ZyuhkpVkX7zLi1f2b/9afgb5lWhKcgT1WKFABv3RJXGHlI+sg
YKWRBpMSLX6R5RHQXmgvB62kvc7R01qljcTRcDipRdql29TusrAjzp3gqIzc3ZUu
Xd7kDchL8SOnOrb/ZHxQta2+0O3bgIlxPTpefjXDcufnsvc7Fh3XN+fwggICz+TE
czE+GqDkzmVIdcA2D0M4ZIGK5rq5lFwaGV2IyKdrJ1ng3U384DLngVe7xpgpSegj
RP+jx9GjIqxxcAcjRmPV70a7MjwYkqPSTiO67yHh0tCFAaI0jMItVf7JtDTxpV4v
3q8ro5bMmA7j9MOiiUg46xFHI56P5xZ72awB7OTaRS5K5v/rJmyJ9O3r8A5Bzf0Q
8B79Dk8GSUTRR7SolBfaEUTdRK/yi1NKF7GqN1jxhkKNlvoNt/Pvo/a/d5u05JzX
5x76ePQleOFEwVGLuHAgyBqHC8q9k1LmljHCt3b67RLP+nbu65TRxaF0U2YWsxQg
kgZ6vO6acj21Jf9bpDmb8UycyBzVvXM/fo9cZF2nbl+vnX86792ZHBASM3y4jhi0
TBqV7flZtZ38ND5xB68pGtaALnjuTB8mEsmWGnbrKYYxCuRWvNPNFBtN4g80qUd9
4jXewYn0uiprUw4DPqfJ0ihJv77ZUoSkHUbd3MLfj6mJ2uZLYH+HbpRRFfC1+3/o
tj37RSSq/4GL8hl8wmDd7ZRkwV4R+jmoRNS03wLHnzWbYOTCSwH7BLZ0cee80/xe
SV/Kfv1nBMpcLHD1ejQmRVEgvIX3fZCElNOotQaZqmPTeDOkhq+HncMN7acq7PuY
B6UGxZJy9o/iveiIC1hMsBA83rxLaRzobU9g8NgKYqoHqp0pGrCse60eVIteZlsF
QL5kLt+25Ezf6gQLSD1ssGdfnPN9p6OwgVlnhfA6Ab43XS4fhmssIBYlJtyhgnq/
kbQjOiuAXWEulEfeJH2iwdyMHfjpG5fUEJtm+c2AHwvnOP1OO2nhmAQFM2erbriz
2UQaQuTwLPFB5ZLp983Nagfsv0w7cH3D953jeApIYllJPx+5t+KCtno1ajuJjW5w
aUAx3Uux/3jGJzZL8zlGVtMwKfFSoyF/ymfx3rLE2UPXX23JYUaARgGRgRh2jwyJ
Kj9SOnWxgEdPNsvHGWORnd7TyzxVBc/tFtu91+fa/A4qJBlwC6BireEKiOVAlllY
4vtQDOhZJ7qkolRcub8fpexouJSLwgrqMkxdbpaOi/ntO1a6GaskPhFAu3zzOkle
p8KbaHFN+CzXMDVDIIkae/siZ0zhf6mrP/d3NaLvgBlndLoeEfmAnSN/Tuf9R/Up
X26loudssgj/+AzAw26xvbvI/bIwWpLJOpm3kz7elOV4hk9wRk4MoVwDwJveNAz/
LTG7OZNGQKogweWrSSE+hI7hAJ2W1JmsqWxErrH8FQ2Bwhm2kxQpyx36JzT76Buq
JH7SJVzmo40HaVx1WXkY+ii4tUNWALsRDFxFagPx8WKaGFe/S2RbTWWloaRDLAnx
wNkteoYzMkSUD0FeHWzcZrhagLSS57wikro6MEhMwRNpF5ewB/6vxQvjP0L3Enuw
7gl3Yu9APJCfHSDKFd8gagRsRS9xiRGVRAAiWAAClJGgCepN+UAqm8q/nz8wBmX/
nUZcDB+kUr337hxCGLm1NMW0Y5VC8lbzTG+NIIdsafqzBqgJDcPJ+245NltclO1t
SlKteah4Qf0vautkNiMjmZMVvc6HqUgEHL4O91XQGB76hv83zcObz2fEt0tG0nHR
fKcTaXAU3GsoSU/oCfGIA1Ii9PmAYOslfvfNQBa7R5suShjAv5TXLlyhzlm8cvpQ
lOr4KiN1J5JAn/jNyI8+9We1jDAD3GHMnXrTbet3RDuBA7eEwrOWkUKeh4NdiDot
CYxZHGf6xf52+D1Oe0Fv68dRM/G/5R8HOpxOiwl53WdIpefvwPHNFJUo9ab0oFI1
6U7FefWqI7UaYn8UNBt4++mwZAw6BS2zeXXSOeDRAPFhDJhITxziFKZmOoBQPSnx
760RKGciDlpC44jNti3ZKzQ1qsr0gEz08cKD1mev7VNS8w7+J0vT3fLCGDXxNXPI
d9ojEFpRBNavGZh6O2LKcDVIlB1yz/C8eeZ9CULyMCbVubkYpz2vrxOFy7VzRqJR
gO/uni44mY9lG+7lwd0Yz1SRrBOB9FLJcdTcUK0FYH3cES/xf1LBsZ5gdvsdTEc9
Fr2rO+19WbSq4tES3lVJ21DJUDPlA8u+llCHVJiAHkm/IRh6W/iTWpzP5OJ3/SyS
l+hBij2HM3l1QXxDDG3qrn+Ts94+bJ4vBxtT50LnhGnZvxr8TByT1wPlYnUvTqnW
mGOC23ihJWl4dfNsCuJ9nM/ZckmpqBp4D3FhLHLTL3OM15SHQx6jJ4YIlgSmSpDT
kHxBitrP1DbFsJ5xLdqTIHKL8cfJouvKP9AbAdWnh9aIgt6ExLG9V5UshtoFlfxx
YfYmgEYBLJ4ZnIKO6GUzWAVSrxKMBxl2R2gmI/2qpEjn1KEk3prnJwJAxHuEeoy1
neo5XMUAJai6mqzY8Dxu99Rgi4wl4rZoirilNCm4DcZhiEz5BmcEMvfZzR9RxbME
iEy3CPlPS2ru1Zqjt/13eO9EPZ82nt8jbiMZnv7vwbE1lDKGk2bS3AY7VRVfiVyR
2+NhWxfF3ygNDbGy+b++XdKYRAkXuShho6taiLLy862kvhC1VEQkJq65DMo0LhMd
hEIeoyHtWij9rBXxipfNwdJs49/fmXcvS9FFPeP/SW2ZB+953ucSEOMiGYg8tYQF
Kc5OIyV0OipNyLpO29aLhM6rPwxR/1EwOITo4A3rTI0R26hBSb/8CmNcYN0Eu88R
65UvolVx4TLE9bR5A9K5malS5Ar/eQmLQNpC7AH05MdhV8Ek4S1VBA+hEtOzzjn9
UsvzAlOkDEcG/R2VYk9XSgEW7OQpctsfSV237zsGIlqje5Yuhzr5PhFn7ZF6YEeK
uuVSnT2n8cB7iGc0p+g9Q7CgXCOc5t7nrXUES/DPmvsTXKCzDwREZ5FfCxI4U1Sk
LndSYoOHMAHi/xB47vyD9enRsgk5x2b/rvbZ/q3gZa45W524wKQy5YylE6bgdIUX
Fn/J505gKeTiJQSsKNlKu1AlU2kr+Y9HLyILEaSB+hnS82AgDqim2jGSOFeBYaiX
wVe88/UXxzG9Tla80QLDwNSe7Q3bye1ZIXqr+ob8RiM5yLPjn+W6dz+C3E1ucl+1
Om0j7EuWfXvjR6oAd60PWumMi3VIRr/MpwqnjeYpeY4vMO+Jj+YSFrUec7NHSVkP
ZcqDGlcDlmQNaUZzTtH0+a8Z4w/rsaAndFHZ+Q/34SHbgXcsqNnPgQZCErRbBolb
byMo2FhdWkHv+c8L3w4ooEcUZZ845Y/VYEboQbsnPsFzaJrXtf6IF7C1+HSYo3GA
y9s0wzB69FPDh2k91UDc0o8o8jGozN7hJN2mcyWrRR+q6OehIJgZZZxCuh0ZGTu3
Fj/xQQ5ShwODM06lwOJMELH5Qrrs13gYqQyYe32QxkKrVhOBVx+LZNWyzUDpPH1P
0HVSqmoLfo8Hwx0pChX4N8pSMuXsyD1bE1A5wmx8xnRvTufGhaOq2+rAZeDnyrMg
jeu4HOmiCERE4+ssGKv32ZAl7Zih9FdoeSBoBWDNfIF8icZDPiEuEot419eflbKq
tPA6kY+KABLPZJjejAK49+MbTMfr7Jd/76S0ITCkDlBKDhue/C2kVTRN+cbDzeC5
oiQ5NJjkX5GzHT87YhyeXEAZoHUqXZvXwAvlXu/jdfBqfufveDoPU5/R7kmm43vT
PejTHNb8MLec3g/LG4C+Xir8OUSLpMor59JAkRtk5inuhLfGpmacnwcI24j3nA3A
Y0hFoB9HuqdwBZvh+ji3qxVsXD94wGfQF6a9jPKtzx3MPES1l33x3AcXqDD6vvGn
clYCPTQOcfL9PhgvhFrLjdm2Hmq1OgpWbv12jzKJqRv9EblpdLl2txRodAtFbpxi
/z+0amLvzZjBjYf7V5K9zanAodgl44OipWR1bBS4TchPOOyZTarqhHNpqmaIv1bU
8BaH6I7GifSuWyFevVaurrsVoxqbYWBPpbBw3hiJk/qA8P0v3PPaMsnDTlLP6CtR
DPZLi1PWhDxIBCDig6+48wL/yLZmuw03urtd5hPc5fqF7LbxT8hplGPv7qiXvj60
T69zb1IUR6x4jYcE1sFOEH6fsD6vauh9zaXodK6inWrT648qnc5n+hWkpTrxd7A/
j2JK9wtQ1yQjF1DxKxpNEP544vVCzyAeieS/JZZMADT33L9pHOIqu/JYh1dJwRbE
XlEHw2ESfV9UjfjRX7AUKZx7L/C9dJG/OcQQyboLVAcbFeDoVwlmGHjGHp1jIwBT
unH2EZbKzbTgKj22Oq2Neu/KgQdggCAeMaa2bIsUbpYMiz3J6ZPQFYn+nVBzJynD
Y3yjeraoE1HDo8goKPGMPrwR0vnG89sguEXsk67hZSE2AL7vK6dra9erTj78MNep
mb3bpxEGTt8OOIqMtVHxnKCEewa6l/iKeR6eqS9AtYmqoP1jBEBAVpnCyNlbzSr0
CFd0k6GshG3ZrnJFwT8oSoKj6iOuNYsWCaBiTlrCCrisCkZ7iJ84JF0TDfnKyYof
GH2iFw/ipSoBAyscVCvFthM6qPMCmbnyysc1rUUJEQU7W4syYueNW5AyN9o8lBC1
qM6tmjGflZLOL+ifQr8fTLtHo43CwYgDyovzLBp/QKhEbXg+XX0PeEMhtlsFKgJy
cyK7ZU9oWwINaovD7kjw6MTbTqDD9eyUGDIBpi1nihUVuLeH3d8pNlpGekTowEHv
7+3z/rYdrSetkb4YVmm3zJot+70myOzkGUfrpzCnBBnXAvX1cr5MMq+WNJ6wpBFY
OlUHyP5hLue2ZXzoK+ApUmPE1EAryDiJZL8bFEU7npGU2uA8ww9V23QmeonBeyA7
d1jS2ET2tMRw+IUUTR9+bf4sjuEOK8lnzJ8KSQB0qxzQMSSJp1kPgBZG63V8SPK+
bvRg9uS0iSOQLTGgGHqUODzdDTF4JXSieonmkB4CabIZcaVR+ovHAOQvxr4Dhci8
UR/P9hzgsAAev9i0vd/qZGCgqvvJb3IkwK3iWWz4+HdU8xe8q/jXtl4CjH+KFneQ
nfRzEUG4e0Pa0oHgak7f8IWwMlDoKDE+jCTwd60p2SXcQQSQqTPGOXrPepGznueI
v9Ly0RQeA73webdYLesmNDaSK6aONJZyUTO/a0ZC4GYZCApJJ16ODqpwIwrdFqLY
3aKFWZWBvKq/w2Wb5V+qWmd0hImjNMake1IJr4ag00qlwcbKkjjxZ17IGiIcRzZq
SinXZ9JmCw7V8Sw3P6fHePL8yWd16uc+/ofIsdrD+N28DYTVTEz9l5ov+ar/oFwT
mNqfk2ah+cCFHo18HsTGL/5P+1M8at8REZV7u2PH6Rz4supj8Ga4MEQPVgb7oHhX
LU3TSX9ffYbnhTPxCywYCArm/rhYhi70CYF7IfzZNi7BANDmeqg6/TRJTVc8ut1w
MYCr4QtxSBVOgCj2hK5Ln+hCYtSTsGqtEMfAL+XN2WLz3dCTGP+CuUeKjfjUr+gA
qlywDTs9NUbM89HURMSR1Af6g+bXd3rzaYETesHsSxGl3YI/Jfr8RNWr/70h0EOO
lqcObezSU+VaTRlLBraYNXb1a4LvuULFSAVwiYLat0yVGdM7f2tUyOpv3kJ8oZ5m
yLfkzGJ2+QH6SWAfGqL7Pr7kGgnaaiWVl4K+ltfPBSTjFLfoq05k271Ye/Sxkl00
483Zwz1vIadtKxjkZYS/7TsYD8xJZ6JbZEpeVYsR/604siMbH/qQuWTTRiFFh5eb
o1UcB5/BA3izzamB/rI+qASfLs8sbCU6d1180sBs6TKXnmJVNnjbCpiyypqu+QrZ
C65Ba7e9NBjUUED2iaQXtdzChwmK0enx/jdQoNYmu94cHn01WN1OU2BdzbjagFVQ
IX2VOzThbdWi77jNLUod4R2IRjstpdUP+VnX4z36eT2Z+5OjqB270shtNPeBv41x
4ncQO6icPor/OyZGgtR2NcAM8muM85YufVHWvGmlIL1xfrZh85w9sL1sl9jos0DV
c9gn9610Gqhs8N+goVmMJTpLAGCxQEtZWh8Ci7ouHqnnP/OdLmTqAWv1GYtiI5qA
Q+SSgtq/k7k6yIuwKcsb4D9PHW8minrR++1bz/bld3wfaoVNazXTpIbwvC6C5/4z
Jl6ZelvSAVkiqyOuzQB5DdhYRkDJQFIU0VDiWG+XdvCa64OvbABWr2xRQwZxwscB
t79f5L/2+iaAydiZ/Mrhwg7EljHQvUJPaDjVVNN37mk5+ahMimaD4G/eLO8XygPe
LVAUK42cqX5DntzXpvtYqzjhypbFWN1VsJ/d5vACtlXfMaEOXfjKAw0EhvRvyl/V
Lc9O02idlTPEjdZBDWtFRYhdtZMh7qahJy6tffT0vyPTTgAHD4qVwiNlRAvHcMFW
5XJUTsZf1HNdGklqgcFaLBazNLWe4/0bEGcnT7oTqdISAu0C9lEbKelu4T4RAfSe
TW/5AkLcTdtKTfoE1Z9SD6jPS6afm4zn8B4l4xi4l2gMza0b1fcVVvRLSu52bVzu
1dqF6SVfo0C1b7Yvd4+VtdSUbCyDJ43RBCZLRvUCOWWrHrtZSVp+b7wyD3RHU89T
kaEF1fFI9k4MDSojY7zX+RCUPvnGnqDm0Rj3qUMDkYtQrgWdHzRDkT5pFntOR9y6
Cw927p18bi5yQkIExFbBZTxGYHLGwtryH9pj0D2epdlaiAYQLsTmCkn6U7QmiWIN
oNiPrB9SWgskE2Mwbdrhlb3riOYhP2cKb7ibNAP0CQAgDVV78muR6XOE34upxmf/
5eg7SBl4pF0odQaL8ExlFNSvKGTTR8TeZYxfyJ4Q2o7Szxn1daCq1TaQoaNJCfk6
QEiD4tBUGysFclPlnqWyaIx+CURYPotngAYbus1LuMLzM+x5CftLtZ+3vi4V73+2
htrW4qdNzZvrfSGOREHQNUxPWCJZCvztuZp52I9dFik57ibSObbLjgbSuhfnXdAO
HE9owjHROTINi8eHLw0UcqTrsCUz44Qo/02bRFDhvtNfGTdkWcoMVDv8Ik04RLRW
3UpqUYh/SW0nFBJPgxX6B2YFqO9PmPWu9l9d7obtO3ge9v8BuzUOzQG09iaAMGPw
oHSB7jlnNdw/4noFKHJto5wBiChfXghq6WtD1ZpWzg2Xr8z5z5GbXu6oQmsrp1y3
xPzqtgKMqT4k2z+QjBs/7X8FNngF0Ophalz94U+xr6n1X1SlOfGYpYTYZqzwzTT7
PFQTqE3kI5d1cj4ZIZTHt260UkxTgcqqaTm3zcH/P0DnYE0YLo4lX3PXhWP0GRPm
rd+nFeBHs6QzrQqQZ4QoZYlWJyb4f2IY7GBqCeIJapLZvREKe1V/6AWMskMf2rRc
Tt3Vcp3BNrRCMUNOHpR/0JWITKr/OyBQ+y8i1EtkWhOjJwXweeJlCPsNaU55lyKy
HNlS242vCpL0oHKlgMskzOz0V2yLSptay9NpWCGvtuGE8V2FNu/RAi25Yn0SCITg
yAURGaV/4t3xHXFCvzp4JnrWGeeERY513XBoS75xmmW75j+rSRp+AutXwneTfaEk
+kXYXf8UbiEMAR73pG0+VVV4XltDqVcmkpuIWax2z0V+xnfnpzqwFq/ZqEWg2u4y
NOw6cIQY+FX6KQhOyQ18Xk3DQ8lfbgX7wSkqA41m+u5V8CiKfNRQ0qklpbfrk1T6
BRfMwIwtouoBhi+9unc3WrJrefDGX0Bj/Ouc/MtvaM6WEeDlOJZNT7JJ1svQtA+p
YffWfF3S8kbNRX7E780PxXVJJORQ/CXxdisr5zd9q64QBv8b+FxNP8ldevocDi6e
qV4dzLd0EhE4LEDWxZIHHUt3gocWRhYoXD1QhiwnOGH5Z5Snh+3b4WybHwilsjvP
K3lCecLdxsX4vjVLqfz6LJrDoNpbBEnazuq7uVd6Tyl03SA15/EWj05IMjhUe6ti
uq7+tYzKJY/1Sk66QjnJaALVCzaFTuOT24vZrCStubVdDJlwny7EoUg8o7gP1U/f
nimr4UgjlTFHozLSBvn//w9pY5agxZa0xQwszjhKedtMcyASVWT0btmWXXnavKPS
mlD58KTSfrMWMTkKb84eRguve4kx4+YiU3kJ5hosVL3j4I8b4z+SlDjsXsLzJscS
855o3/RspVaaLYFPznSv6uRL92huiDdbdYdqc0np2/7s7WGNUb3VXKLk2u8xMrMi
ZOHo8sSCjobdXCsroyxpWE1tLnI67sEdSl9naYamYmYiVm0m9sAvrtNRb7rz/cGF
kKvg8PEcMN1ne8DG5Imt4V1DMs/zT1FjEiBo+t7Pe9A5vmJIfhracWcZchQ7vH86
lIXuFbHWUpJLtzWzjvNa7KAP39VYxrUBp1hcrszy3VjhP4v/MWK9WJ0fBuF9SHmF
QJlTMANMBOsMIq2n4ZbI/IZ3oKHQFKB0Ca350lv41DQD4vR00M03Jia5K0p8r+CT
V3zMqsmsw8yM7kgBI8BlYdTWYMtlqWqHgg2lVoT/h5BwVVNxzIUXmzgle/95qwKh
Gekk58r4W8dio6fucVnhW4XacFPn2hdgwt378YRkeN3WCpFRaC9RwKxIoIEqntiD
DX0Vxqc4M6m0o9W6EcPQ5PYnZpp9lqq2zhjmXvGQwwZxlxq+GHQkvX7OhJA9XRJJ
xN+4wd9Ctw5aFWA3m+n1gewUQtxHiqA+8h87PBUAdnfnh6IOFIQqKY+mJhw3MgkR
cdX/MqH8iswih1JrMyy8IDHj4n6LXo/qCpHZzlLG1Nbt+yrLG6gSY2XlH+h6RD0d
zbVWwjOFNEI9quwxWsMgrY9nPpCD3TCScODqLTUUCdV/Sx7y4GT8ihdPorU/C5PF
+kEfMPCmOegh10+CAjwv9Zrm28u97o6tKUAD3RcR+yiJGHiB5EK1LOZ8Evti+1td
0HtbxktuxYiBRSKPAR6SfbylTZIgMaIKnGNssVm18Fb/APe6kNqC0K5+eAcPBwYx
8+m+huyItpBjE7tyNLjsbTgqIPemC/LtqeM4abygcM7hkG6Xp/pPpCQCTb8OTGvE
aSFx0/kyZDRBtLbfLpKIWc68sW8BG2wnTwghtkw0LarCjcr79BVkYah2lX+bXff7
U6stae2yHk6YD81+knIk+Pldtn1XeuwpZ7DprYnu6e8zO99HXT2ZhIZJumhr1ByW
AgTsTYQLaxsT+gSI/tINxSYMq/85j8U3ot+7Hh8kpL3uPj0mWiii30zYpeAeDkzE
YNoef67iHeY0mD377KBWI1mRaA8FcOYOqvDcySC7R03phWk3wznYiBEBRK89/Jww
F2O1YQRMwFW0t4OvPR2ojqTAIAOBRWWnWCKpngMnLMbNbCjK4C3mh+nl3UD34AZb
z6vP6HRz8fIRuW9m+0IGRQ4IvVNk5bILnLJhy8TbEwTTuGljIvWLdVPYIEISw10e
ayHP+PEAq/SoGRU0amNPwgPnh6j7qEuofv2W3b5Ci8+aAAzbgkPp3qGRKLmVlmFv
H9lTeTBrhWpeRdEhV94s5EFf6dV7wpcA2V/Rez4N0eRKkn3sNWqwnf1F2VITWUeM
KO5eRhIcqyPB1mSThJQVpLqecQwgBVROD36p1bpHM0O+DEucYmYhbFkq61JlQ0d1
BQ6AxMbMumKPmsiyfDi7dCEK5adfmf9u1wRexWLFKzJdYekmcFs5bqXtbwT1mKQX
7OiZIQPj8gMGm/AStAebPrOZrmTiMzppJnVGh8PNkyNW36j9ciaY2EMaz1PfSOfZ
xWwmLymiQ8UdWBABYlsRRxXzoAOPVGxgLvDMLhRo/OBHOeDvR96wD1m9fB3ASa59
qAipQwxHw+qS4RifSJwslk+tqIkw/PH0zOoan9PFr5a1xvHI9ii9vO8la6nmNNIQ
C1zH25wx3XFVuu/IeWBxhfAg87+3B1LGWwVpGLfydP2kIpwCPHY4btpQrz0i4WUv
TxGvYNnOIu8CzFF5sgv6oaE6hlFAGRAkaMdU9YElLz6uIy+bLP8R2+2iUhnqmyTX
ao5Ri0IlPDdhpaa5GNlcizX3zQM2XdPexOQwUcrz7HYqhd0Q8+E+Vbquib3OmjzX
WTgj6lBlhl0v/HlmTSC9xzQFTiYAsBHiUuiw8T1W3uiOutAFSHQg6HyS91aH45kQ
unPYyi0o3lODT4s1FLoComGKNQf/l+Dk6p7gIm8zGvcBCfrtzkBvGHR1M1tssQW1
yJPsgQ0sof5Jv7gpVCxihZSm0EmllSIINGdgIssERRylxw4SOxRn7DSV9QnBRFbI
tCFeHTUOBBWH20TxfJLZfrafDM8K+UasEPRGbh4Ad43Gyw0G/fQGoxMDR0Gr+/wS
FOi2jANanori/SbEVuJsxzplO+eCzAI8/Sl2kVPmqVUudfj+/zEOMjNApKFSRqdL
b7fGqfj/0qZoO0MK2g2gBKE2lnPwDAgzjGbdw0r5xXjeMvgSSvHzflpkfXD97uPV
z7Ps5fOJHjyKL9IN0khAVDpUpFytgPyieOBzf5Pj1MXaxcrGuPN/51366x3WpSJe
IWsilRB3S0mmt2c0tQEP/835llMH7Uap6iwOmZdYW8IEOvuhjMrnQyW6acyxJ4ow
1U1u9GuCkdoDl0cdhk/RPlVYmkryhq7/KhglQNJ4fVPpn8Mq/eTLjA6iBLFQUnbx
zr8tVoNSZwEC1JS4YNCR7DrXMwOaOAQkGb2rA+wNNhnK6kaKFLtlhe7oYPBwawCS
0RMj/aQZqAmqvbR5P1U0Cw+xglrqntNMJwU0G+J8mMyOMmD1frnty0g49ydNcYgD
AhVzqbVEAr93PNHJ66FeoEriK1zPUbVS6F2HRsh7QZrnqdg+7uFqfXGuzZSsiAOe
Q2CnjtV0EMC7eaUkKVg6hUibHWLJ6u8OIXxPw31R4oYajYjoT7oaEC2kITe09E+h
VWB4rc1ignyTCczBiuywgNeS62oVPISk5PZ/TXiw0l3o898fS5cHMcQNu242aG0l
H+1ue1udD3o5bkNoDqDqXtnxaHxbrrGfzW4K0n7sftEqhnzGASBQtcXuhICyOMoF
N+qP92J9QhzIPHr8LeIW7BvHJa2kiTvGr1scDab0rLXl8HkVDU74HN9Vl7NYsMZw
OHiGMkcYgnPjRmmeqMsyQ1Xssv1Lhn4h8FrRg6Ts3rWFCBIIhLr0oCoaVZNmqx2B
GQyrSVcXDHTgH0cNXt/eOuRfL61eWRxebHPJbRWj8/MuXSCgAhr+oXWeqkfoZyTP
L31ETalVTFjr1pbqoJVLjjPTXreQRBY2EuwamYLzp1x8r33JBXSgGdXq6hLzQ3qv
dZm71rjO+IicioXgOBxTMqC4EJxB+RtJCit3zrd7CNYjnG3C6ZgscOYbR26zzI0T
oRvgbTEm5fFv1yN8rgdDbUbKugavjAGip/2kE+/3pPbAhlWK9kvWVdoeO2iiBHFo
MWA5CTlBUUxEPA9bU9rY3ayz6i5zzOV3AW0YtsVntAz0Ld5txDMoLtw63qHhFuyY
OF2Nh6+rs7O8mUUQw+GFYG4ReFyOY5BYljxhBNmAgW7Jqx+ygvJeGAn6vt5b9PZT
fcH2dvp4OJW6yjRkKz1pavNLAo5v9zsID+pnJ/2AYaOIa+IP/7OJr11CtQahRpy0
yHuHtbUWZTzYkorK2tSftkYauW3fGqYQ3KiNjPfA2utS1HJrdCwDewscbWlXhrxU
5e4T7Gw8vCwCPJ1P8Ee+Saiq0Y4TbwnVs+j6eQBhPcQIs5HDj6vv7XznMjPV0bXs
gQySoSIpNS7sToCQZswBBEnMzv1mYkPQay3rjYaeX+KuPPXTXvUtO+F8tY5qiDP2
CN2ZgE3FhvvPxQYLgtCNDlTBTIyYRYlZRjgfngZiETv9asyk1X7CMXPT2kmJJPdP
bBFeFC8chVlNqprRVDUvdqsrbZz13pG+rXCSK2Re4CAnwC4cn+vlWlgesZvbulID
A0Dzf7E+YJk/MPrJty3wvnDps/Z9OqKd2ADGSwwyrYnwW37pvjk5aDN8VuZ3e+vf
9AAvXu1lzz1XNz6U6gSb5AjX7DZ/xhKnukzYiS4tv3arLf8jd157EL71Y6FxZ5tn
I+Aim6ZfHyCbUd6R8TEC/hdPOcNCE6lM4rVW3UINYpsOR/seH/KNt0V0eVIClf4w
Q89GN23tsBTABq2Z6krghMuiUqvXuANc6ZjIWur0cZHH0GoALV107xH1oHe5D5Od
6SJIOvTLzqdEKHOPn5GfeS0fM25W0lngRGWAhA316+CChA/uZkiv/hlTuje9C6lk
Th+g0lEkkvcM1GLZ8VR9LNRCOd8W84AVhpnD7bu2Ru43SBA4IeC+4jJJRr9QYEc6
hvuO3nh3pFF9/nrLXWbl8jwHfVrka+q8aPLq7niILiIwSHGbJxDrjwF7oFwUG+2v
evOQlG96RSozXSbxpFmfPY5pfAYYGQQNpgDY7ptn/1ink3lr+lK8xzmZqTDWOPya
UWm7GMXnoP+iiIbWYEs0v2GW4L1IvTjNHEynM3Rx9msHW7a1Aqf8zLqvhnLo3rVW
JzHIj/fGyB4uyorbW0AAM8kl6nbMvBzmn9UFPv/s3tNOFQp2w3Yy45nSe7q2wfJN
M72c/Z00S6bPB/60ENvONc4eySLj6bmD+DCZmCPRYzMesCgLZYmKTxeEA3ucLWsE
ZUzeDZ7aO8pRAO1i2I48xwItstY2MsoNLi9WfUJ1yNEhGBtOYkw+qEhaGG/FwTmx
dwowdEkPZKZXpIlxBRbP7IsZRcab69nBtD2ToTDOTlvF3q1us5xNIQKjwSdt+tK/
QFuZL2ZH1iQtXpNf7R8KyNqmFaN5S0S/TMBDprRRXHn0uShnEhYtnQTmHjljtWk1
n+kX40oGsqi4FFi8MgdxLd4Aj7zaBbPiH5UqDm7RJ24qchZBEaakVsv+kZDHO/Ff
zBvK+y1Y0EfLWjFOvlA4iyJX7R69TIAGZH+Uk5wjTFDCkEwzTYGKf4ZkVCX0XXJW
xkM/lAb646yKziFHeRUsOGoh5UER+DA3MpjoSCjrSXAr0pucshMPAzlpaBc8zcdB
/1dnPzV3BnpjXktBJ5psGZO4fyIxCHjn78MZokz3Vo8b97TQjpsCFEawyOHy7um/
a0WjL2Ir/LSNG0Q6lbEkJAsvJDp2G0Q1mBDmHD+Wz03m2b05uHgMQU+E9ljXVWRu
o4Vb6/rGhNd0dQm2MaOU9qre1MZGip14BWERS1C3DEQy+M2FxUbOpvdZ93um9pZW
3nfTvNhniJmtr50++W0T7zA7Z65/Iaef4XCfWJcvEAUUGJ+hMoVgh5yrz7vRUie9
wMMTyChUd4MKDVzyCjDsaHveCXG4eTNOF1DviqN7hX/A6piy+H+r4zQNSsjugoar
5Y4Hh+MVVnTEHLgByIIkL2AS1PzOtdCgsLNhleADvXWf3IhxtCQAwh+14mbnTAVa
q1snFAw5pI+DMWZn4sF14owQ2ooLYVzTyso15TnanHX/fcFmte7ssF9xllpq2fwR
vp23SNQQ/COV9H22MpbFqqPzfNx9CgJBGayi48DoZ9rakbHDFR0VklCLXb2215Or
s8assOh5TxX9x6/35rJ+cwWeLcfllIxoHu12UVfqvTyPCK3FpjOvVFFEksdshq1M
lVdml6PWa+CSdJO/2mYF89SjKikj5j4WiL6M/IPBkAipYJZr8X2Anwb/ZhjlxId4
yaMqWTdJ8h12WV6+sJzCsWqoHwgkNl9EBDvF7tvR99LtnMR9DVMKGcXU1dzBu/i+
OhtKb9A+wtCVmFr1ASg64IZYlgtv38KUbTFaNKtE9Tv/p9AN1//MpCiCwaSPl0p6
hwpuc6rmjV1EeFhnz+NdwUnfw9CwkkBXT11lJPnT7/JmBD1J39TZARjVP1ldsFJd
8GIzaAcXFUtUPo43TbQJY6LIMw31+EdN04sZv1oKwqabXd1BJFR83l+VXC2vxnJf
zgY/sjfn4t4RcGDge5Ja0O/xpIGymT3WmsjeRr4PpUrNXlxHDQi4S2d96XObkmgd
jUItiB5tVJICcTEYM1ZYAGSNfGyI6UYR97v2NH4mVyXxRAXUdFz4hw2tOlaWQHXh
RuJurHIrFvOCbhmBD6G6VclG5iOPS0iDwYudUTUS17TO6AjK9EM9FZsS54lz69fA
Vqz9cdJ52+Eh8le8WS11G8u7bDBFRswPjBmINo2KDgUT2yVFParrtXeBc/sbxXKh
W5aBhes0g2fT1KIMc2gMED9x+DXuUj8owxtUb3o7gLOPdSto0eGukv6XI1bj2NyR
hREtZtA1WSOI8v1vV0pYvUvcWHV28JL3v+niRRy59AUXiwr8RcxK39vKLK3W3UQg
RUwZ5Laujm7iBVR44ceSeO/T70OqZ9jS5NFZ4ah2bYKd3Wor6KsDB6audF5nUiLg
l6km9TU2u2YYFgwjSmFgu6HId0PHHbfeg2BgXR6a11pMgNHlnWq+LFfs3d+dYiqp
lAKsfsE6VWti6XGOe3+ftsUMPEnQ2O3R7M0DoukuERbDLMBR2mIvSROu28E81jQT
RmBenPo8/rgsrwRop0lBMay/Jvchov0SpEF9eMj75z9V025nTk7l9elLxCpzUy/Y
Q2tDMfapi9yFtpGHGUKFzYQ/lzbTmDKau1PHyRE9YfkpBZESjogfNRL9b9x0TnSU
X4h4c8qWp/M6cRQx0EFH6uNwIe6i3ah+YIuCALTuklOVH6vSdTEypJ4J1FrDMJUD
GHmSaspi+ZfRhKIsg3ieNtc+QlTvdTaTIxyZvt0WG6cl8kW8nddq55hlqR3gbX2A
WbZsaZLaJNkOL1NBd81KGuaULU2scDRuqy40Qi7DCtzV6fyI0HfK3xBKHAMjwGZq
PiVlKShBYz3ZcxWueLZ/ai3CdiklwT4C3BUao3dLLnKOBkM/QVaEPQQ60uK7+Rz1
TeEQ7ot5jVHh9NGP+cSeRYm7i9SBKdH7vkCdxvm12Q3XHABd//+G/ZeToZKSfe1p
yjTlgOT1sWAT2P8YMAUPUPmRrOfKERFwkWNeobe2VFG3fdVtCCV7u+75A/DdXEXL
KJcG8sspNgrDP2azKho20WCD5/dFKqTGwCbVOWpxoyoNWvW5LN3gUsRV5AhVBVqA
q1WI6LBFdVdvkqEcZZeVsSh2sWRSSpS6u6wtw2eS25wxm0iBsUxX3VqVtwecM0Jb
lwGYpXHKSb5CGw3hAuPK3JAUWNzzWqDzajjLSTpaupiCcx3KNUeNsRnRd+6HePCp
Mt8w8urVvE8udUANxUxlZahxBBj9L9Lbo+QG1P9fHTvOPl8bujxfnbD0wD7Nlate
NJXSgQmMuncrV6Rd+zJiqbQh7k3J/BZ2vABAYbtVcOOwhOpF18u4UD2SiZExmdXA
WX0itG3tyIleSbUqcieXKgJvXRCAnPkRgrMnuyqYvVHVIDTpShVeyBqh0utTNLcm
b1OWrRMni5P+i/sresE6JIm2uBKtlb3l3L866jMYf+Ppy4kvvSFbXJ1rZxPhA9zq
5YzaYcB0x1VaVn/rjLfu9G6mP5Adb9MYDJBQ8RX9P6wtoWs1048Shai+8wu834dj
rvb/K6PcM4J3wG+J/OKtJIbK94iMt1iPMdiQynLe//Z5214hQ5o7xeYgSinEpFzd
XmLpkewIp+oyRzoT01h93moz1RrA201R7Mjs13n+NyIpJE5C/XoI9S1T/oa5+CQR
ijWiWLCsmWckEH7FLJezgCQjN5/01p318G/KJfmVjeqjljKgQz+DcOEUSL2TcyQz
L9PJRmeysUG+D5WymGxw/jnTi9BSbz0qAllswz7oEVOp1p82nwGFqoCGKd8J4/6o
osrmCSsPh5DXVgXCXpa55TFqiHBbkf0+LpCZr1+nW9L6FMANIpPRXnKHbbHMXTfa
+ZN34CUkmACqB10XLxrYmnnEAAvUBHKnt1qoyWCbEjcyhE0qiTwpb5ZmKsH/F3nJ
/Tht8O2txQjaHXScdwzvZ+92ooKjBpFgpHXnEdF/gsfustTXzNkeHp5qbOjT17ZY
9WQK7vjxEF9GZwJqty6OEbjCDYI1qauH9lUXw/1WxnB1grhP+IPms5QNc4W2afNd
2tlPoLnb9xI1PUGo2HrrbUze6V9D4rGjPYAfPexjHtyJVaUB8QEfAYpS3pAw0x7p
ce88ukv3Tal0WPQrTCokVLdwxg+WFDTM/unzCRmmntwMPPtp+n8QiM9DfJUrPLOU
yVb8RIW06RM5xXnUEgNC4Go+67R0R338dpgueNXb9aoxiz1rmE8XNSSpIGvpz8TJ
5nZ39D/tEsxuf+jofFcOLZ3LzCx4VFnP1dTqA8cK986akfss/WmoyH3610LcMSUO
u4Srlb1cgJf5WSNLthCjeFz5hNaAkaT7ShjmCvzX9D6iNTV89ZDvl8lWjzwdxlDZ
68xwg7Ail6ZLkyOUQQJrjyyg8xYz20PYwnUO4DBlwj7NzD35lV0XnhnitVxy4wVA
d4b2QUUaq+QC9iuVQG6BTpu1CpwCWZ9AMOhGn8mTyVDNopV4s1bhDupcgPBfgVet
gQ4qm82sI+tmQgvN6oGzwZkzawPnSvkDsx4fC9CcWKS0f7SR1TyOPqhiZ2vgjfmD
fBF7Il3RnHZ9hhuFbJLI1NmTTYSedYH7PAfsPdX6aIR5z++TtPe+gUT9II0Db3T1
TB8H4YqicFGeSgW8iJE+Ce2xWrI9QrYl72Z8UMqhCChgjf5YwnND6oaqelaB9wWG
iFQh1zH380dSqhuGrBpdjz6ANZBQGDF5qFvkpls2NohCAUvcO2+DMzi1YZBbdvbw
RRJtgsWm/LOZENBvLZK099KYecX1OMsfHUDydcE7Q4pCHK48u0f7PRGuwezs5t9T
C/AUWMlXVS1LGNFDvFMXW+0SP5fjVPe56zNcqEtCRvui6uzwlOSv7PWG1a4BU3ud
ThLY6f7yNDGCpsYW+aAPx85T8JnRHCxE9vmZuqjjsFQ5CPkpUdOUe0a7uuZ040lm
EwC9ny1SG15tTbnF0xxQt8nFjY00R5wNf0eO01ruAhPGjzDPVAChsM6XuGUdTcdN
/bbN5qNP1Wq3aMmJd9tlcU0WszEe4PQ8SOobUXMde7EpNHVAKyS4SPbd8rCfaC4+
8LFpCNvIYxOE70R/+3DmY65E1KwfJIrnSU4izhm6o0JDcmxvGa1agwnqKNu6PIxo
bkBAJgPG7CJ2YkyuJSVK8vQFVoDDvz7Pvj9glYdcJVrDjUkJhWUlEIhzsz6jaMPC
lKNQOzFgGuvmwtVuy+nq+mVEZ477ohW8+pIPewrFQJvCFO4EPy2SgNoAYecxpHj9
hT8XvWJ/RH7xMUuMzEdweR6hMGBNxw8y3ZJMYgyiJ4tjRVegaAImuZnvCdlnS+iv
gtQGzBRThNarwJtsO2OrV6sxr/QWTOMEN98cGAD+u3g/+hxhvXfEFEVJ+TKh0Zpg
41PP8Wg1YGt5m7eLSyJoyiVgf7MsLfQ2bZnwIXyoY/cdmSy74J8gwtJcpc5nuqw+
jlpQShq1z+3FEogDQekUIODDc8vIYmEeXl6BT4utXceZVGKtOqHsRbCZVybgzPxw
IeTT3fv17GzVktvS9zSiAS0yBbjxnodaKJvacCMNk38tgZTwKvzBi7qZA79YyRlc
+6ZjH3OPqYUTc7XSG8A9mFUaBhwB9lLqKZKgDQ0MpyTAUooEvAIx6xO4YXXyIAnY
ZsbaZJhxDj26Yq8LANlsUQcbhO1mHyS6OkfJugGXtNW9rl1dc6zhxDy+Sp3YaVeV
Gojx18QvkfvYdhEDBn+56/V9azrhSIEI1qFE80/RlCU5bCuAig+pdExQM/Edid3t
e3TCRjCtLeaaYI/kZVHenrqyLgkxO+jt4OCiyQN7cpD/d8+sT508XJWXzCdCtBHO
n/lbeDg22YWjXtC6oN5FZCd9N1gKigiu/LfciWN0QBnObFHt2haaAAJip67jzrQY
DBcdejpspxg70L+qDzI7dRf2pxoMj4JAAGcy+kBxeFp4ANL/qY8AUYTZu3lwqgH0
Ogerxaa/7O5auhS27zmk3XgJkJV1dZbVb40fkzRzgPj9trrjNyUJ4tXnET8LG01t
qncwBh5Rys+zcqvUFmBcZRXuVSyY/Mt5UyLXR1nH+lOWDsa4huNaFQ2MPr/uPJKs
cRF7poPCJTiBM7CZlHyz8Lo2SbD7cgYAYvEvhBHRNdHlZFl6Eek1JcU00tBKtJjF
G0MkRh8+EbHMwdghkh0uVkKKS2wZHSKzc9P7G2dQPK22H8SKFC02GeTjh82cd2W2
W8C/2uoQrKHHyVcmnXFTDlnX7hb2PD5CfSVtEkg6ofiV9Mj90MQW8JrfYdKylRrm
t6d9cX8PhLewJwLHyiZsicjyVKvm3c3mvSoT15/1+itTuG+HmdP4x6mMI5EoOwlO
H5hAhUoI4i5czuLnn7dGcx+TCmKeGO9Ae/Ya+ATHfCviSO3XqQOUDRlXx+US5t1f
oIGwupUJTrOnxDfFw69QqP5Qt0dwnMnytQFEeSeWLPmiUmml+ZouESqGPmzpNESi
kL43lvByhQBFzmIaQJWxGa6TV23udC+jpdjt4Rc0IDzZ1xOqjTmv1ewAae9J+djQ
sSMqwEtdvRF/PxujL5XHhDyUr8v4r8ZNjd62euEPSl79UBZd8ATtEVlPbGXIwz8o
hS7+snW2JJkPWPyXAw2ROrIBMPEVdnwEioDP8CkE00c7IpScnq2JwTIn0aYx5yLA
Savj/qy8GtBif78/RthgfZUfS37Y2CdtfHj+CZbN2vsZ2MGi/lNO58H4DS1soJ8W
/ffr6T8nB7BfuMZtI44omzHmL7n8KSNvIlw9bFghMuuriPMPlolMwmohQbGOKrt0
HLYG80kI4cZ/tUEv8S9I9teP8pNxTZ1uohLToWQttLJz1hl4XD7/p7MhjriQkHWb
qTYzgYzLlAyxc834bJLUnBmm6Q2vgvMwb5DKe350e+ZIyJGhQRsOKHrQFi9y0VDo
SvOrM0hWEPmzS0ePWKEPg1SScinlfTQn5a3l0y+La14B+Jy+q8rfMrr7GgMtSpB4
6bGtFeIDnnqKveXQ2kewV4Hxva/q9fgQZWJEEeu/GBzCJ7Zt1uIjO1dnjSzdyqBx
5i7srQBcebyackCsgcoAbCUirgAqsH3n1kAGbRJTaa6Atq8itw9sZLo/Sfzpm7N3
a1/s6y/v3A7W83ySOn8JzsuuDpy3+cs2MWwNP/1xwYsCZtbXB4k+GljkOLlvvBre
lx5CuISpgLauZ/7AS3IKmn4XZElJYimf2WvEOjvDAAvNk2K0rN/STYZCF/y4VXWR
tpFFm1mBf6OWq/OBUdKqJHlkwC6WZzIl6+oD7C6ZFBOb0epagd8T9wZvHwOvgSPT
vJvglUX1P6SEmUezRyAx1t8GfQ17BGcgaFii1uuUzJZHVywbd1xPS0qNzz1cHNXC
PfUddxyEGF5Yf4Q2kbUADnhL3E7E3shkhHgDjDjOHKAYZby1M21O+nMrXP7YUwSu
n9KlYoJ/xhJEC4X4WXBFYXYZGCEPdF3uiGfLpuSi2DFF5qH8BFbEGC+pMQh7gY/+
mpAfurmLL1GFtFNq+rDoF7iYxlGt3xlj/QZzTE/PshSvtk64j6iCRwfQ7tr0k9x7
DiygIQf5K782WhvarJN7sTsXOsIkxSK2l06JkYWuIMXSBRb/OG3MhKQySCI94iKP
DUnFm7e9GlqHE7sA7ELVjIYiKWpLxM+ewl/LiGEKr/eo+90mkr6i8Ro7OupebIEy
wkv+dU3nr+8RvxcuBMbv+HLrQxQaTLtYcsey2GZMFjiIj29+x7HWFks4dYy4bzfg
0SbvBwK1Sn+wI2eeHpUPyVN6F4ZlXbSBx1kfIo7BW4oArCWoBE6T/snS/Z31DoPz
u/1qQEOtOdO8ijnS4t6HW7Lovmz1HxOegOYUYsVr9uawwNl7HB6B1l5HCibqf5ch
Uf+1r65O3SEOumj8jrTmMJuW7qzYrCdf+8hMsURvfno01gRwoXnUi1MlP+htJOuq
aY8J4sTM41mgcduTA9D2wqKNDx9iQjG4zbDaOCnfM23MHr/3ZvXjVtjPWg9ghjEj
acVs8wj6Pw9PVRSJtg9gLLFaFVAYjlrtGb5Qhr6T4FnQl0EN93X9I55uS2rhCm/m
qT1JhoIs/fexXAlA45P3pCdziSz9sXdZM2jfSBD3xfX+H5A7UQbWpE3Z1CSGpgoV
RCKpn/fKxTm8ZT58a92o633tULdoTh6PRCqL4Enhu0awpY++hEa+4sl4ij6YfZzM
mZwCCvESzzTB9w2XtJekKdYqsAy7EpFO43DkaMJn+N1Zc7Qz0+qIp9T14cREhCMK
H8lLvx2abzFzKeOA7S85+BacDttBVb3WGtwiGR176qOHt1vm6mwdLebaNNTe5uLi
zjhLdEqCS32UNcBr5SCTbFXtvQTrCDTt5dRtHojhn0ERpxTqSfI3kN9eclCyhtnH
c67UJmnUdeDGof6OvLQYOBfGaSD1XIghxYXGwIgVHLyjDdgsQ1pAxxgIPjkdcON8
ILl1Nu0GjnOmG35+ISOSvY/rSRjmEigalcBnoukO3jG+75TvVH+RgQy8qkfeW+GB
pSQCQ08H1cZt+X4O1dD9F4pD9XhbKUn5fBJVRPNxzgCf+5wQ58eMn6k0XzeepcC2
V0KQ7X+hT18HqiDa1MBIcS3b8w+Jf0TjXQgQ3HOl+i0ayCRoypGXqZdFp2QEEiFD
lHjKsWvReYIeS7Uu8yW0zkZSWV+boFKXn7KY/JGuzaEJ+8op+uj6r+5j8nJKNcCB
W442k76s1pSVBjSeU3HDFTFGbGpfb7nncyPCdSMEn4BUypdFZrR0oih6TiwZS4N6
dHYSK7FkKaHm7Sixr7Qw6vSUuGvWBIjx4xWHi7FbShiCQbdmDRAlXXk3FrRyp2Un
i5YJil2BF2cEgN28C1tBDWtcaneiqkVIDpIddqLlYyIeAM2VgfDahwO4DrVcvkfN
LaUn9w5I/mMTNglrEiGG5mJVtJ7KJ9Rgbx+ImF+qbr8dCqpdYaQkMvAPERlnYOmC
GBLXybh6qoUNvjz+6hx6cVKzryI3fA7lDIUMmU9LP5GoBk139TEA2TGxovxX/DNI
+G+IXSsc1mTyLhMfgo0aT/KeWHVqmb7+7TmYH8GAbLYSjI3PRjhDPhYowNOwyiYr
p9zqgz7KE8IRdJumRMNnGIFz6GVedolLvPVy//kOQuCtaEoAu/yPadohueIn16sX
ks4xa2N5jH15lPmu8VgojGp2r8hDQ/Zid70k9B/29aab33o+ZNuq2jOIgMDVKdgL
qlHlxkSL9uUndP6fnYDp7eUPiU50U8RA6ilQdYFqSW7J8TJ+tshgbeWFsmP1rPe0
1VvBjdCU51ZomkrWY2mB/rPN+tf5XBCDMC45MKAvwXJHY+RZKscsaD/gxUDZOsZm
NvC+tCLuUjf6oO5y/9QutCmk/y/R9T+cziLnIyFCdMvX1MV1MYxYq0xcR3QIwOL9
f9orZaPBZO3yQqkusHtDKknP+gGy0wUJWLVapzAjk1NV5ObLsZvBQ9oKkubbI3sk
zF8DJWgzJdPqEeGfYweCPjQTsp8Ow6V3R6OuRQ7c7TORTbOqgruoD5USerwKC2Ln
B3qKPxEXWpQTNLgQNZupZTPN3od2R+Tu8qC3MEbZjnY6X0AaLcn5gWFUE2MU042X
29UgBWBldDKnAytveOX2UBd8ofTIUmjMNQ3/FSquZeXFxQ/sIraKDbap9sWq50pO
NkVT0U98PqfACS+K9tvys+QVMLflLtrGo6klHwSE27MtI3LLTtCxJQHpUROw4h9W
S2MPPTcIVpth+SznPHUz6695d3fHaPt8LR4aewXYBdUUR1pDApOs4lvHvUMXZQ1n
FOsSJ0RWJ6oA9QofW9WOMwd6IU6aZrkr/LCRayTH1ItXgZ8FjLWNc3JuBANpVqhG
QUFKs6qOIrBB0bO2QWShlERdCo07cuA8e8Chgdo/OdNOLj4jXdZjN3UbYii6qsBd
4nRGjU6HVftsq86OwNc/yAz1IJhZh8bwjMTWwlQsx2ze85Y9f8/cn0PbctBpYWKO
svVSgTAMvT/rjqN7Ud/oLDRCL3VZgUWrj0TxqXN5ZZaMML9M7DS+42tg39fRYbS3
eUp3cjhRYAE7KRevbldFBFCABB+b6wAFXY85oAF3piXEAkDDizfJk2wJDczt8mgn
GNYWebd08ngIqS8kJPP10IuvSp25Eq4naemXgjwLiCA8XA+6bX7EogWe+jJzwZZc
E7UzJWp17miMmnEK65nro+VLOdwuXBTLXVvXfsWwMzr2MPEP9ah++Pgq5uoASuBX
Q5RKt7UqhfvjEnr99wN5WqkGzvS3XtF5R5CQm4Ra1f8hEdOe0lzPA/tUSEk6LVbu
Cy2YLvmqRHAtOVLn/y4DS10jZrQrmHzn+YJW6cZSLGm0yXwcNbphKDt0lmzpp7UB
mHBA/RWZ1UxW49k54NIhD6aqe5VuhxS8TkDWqhBKbrL1dAd0DVCtAZMxs2D52oZD
pUtQt/jUo+Jx2j1QTZki49GFi+T7mFjhP+G+W8CsQQ+YjvPTJEeIVGPhwQWaw43H
XZUMAuhbhfHo7O7hXGQoSVOIP3cK20fWy6unDQdDGzJkBPbkSgWnqqWK91vV9V1g
f5x1oQNFjaqT7mTw2RABynzGc+EcVyadgpV60Jt+GpMiTFYBasIcM+BnThRYEko9
QHwqUkCxLZLR7ubbS93U3Oex3LdQ8riZvLcbZCTRe1gBH2SiOR1DvOvKClOdsOuw
8+aBOmPXtoLYnhjzO96HZu3dVpQtr+Wsbhg/9o90kTMuajpn0npc1xA+R6o+Nspq
zZ2X1j0FNJWbLptKodCXOKjkO8KADtCGoLz8dj5aO28yDrkcp+3blm6s1ZQGh/xZ
JHqxwgYsfnBPaR92rjWT9b0MkYQAhJNuGWekVS9apNGXjp1I39yoYKUgjwN9oXP/
j0LTK7zEvKoj1ACptYTaDkMP5dU3NSq+iDFuA852Lp7u4L34o+26WG+viCLkJF1J
GwOmUgY6taQ9Za1QRySOJBhhOQCNNVESfvFg0Jl+XpxcmfMp0EawCcyLM/kDzPmx
nr3V5Doaoh/ij//8oniJiaRWsItPzJ3AlLy3sbO5667pY5USt1aW6jUjPm+6FhQC
LmqUNsu6LWrQOBBvyHrSZdw8HS5OTlyqXwgv7iofflUAR6lslhe6hl4kDYDxlyjt
0X33aoHd+hwr6DYm9o/0f3hRyzQ+mQZtJk6vYIutDVcH9QnZoMbTowxB4TbzPTRM
cu8PfWG2m0/utmDh71Y9YgknRGHtgzH2HpGs0WbxJ8GeBfbBaB9qKI0yJL5RU4Xf
dQcHOOT7PTKTLyEuGP7OMmO6pb57pL19Z1J6NWo3XKnyjpbkMxsDWLwV8B6Rbfq0
xVXfjq6IChuyiJhzz8OfCY7QucCcMcSOBeCsHqyIUtp4h34dpA3TQgwjCg3vLFwJ
PpdCWMNNTjmMDdTmFS8xIimKAprasN0kduu+ivhGyJEocsk7wf8Lz56Xvtj5u/6C
bTArUcqG2GR+0KW2x8K6XGdoto/iIg3nTlEPGxPRIoG34V/oYDhty666ZDO4xDrE
rbcOSKxE/SrAOg5qaO+8nFT5omCj5i6L6xXGsxTx35i6TBXMzrDUZB9hEIFsGDr6
krhXzR0/nvdbfM3GrSAY5mQxTvLwBVmiR3eL/FmjF+LLC25vpf/5BrPg5hCdkvPH
ZoiSHKaxFD6P7a69uMEgvommTf35uFusKqTiHML7m6y0KJSgJKIWZzoKyBk6lKmA
zS2r/9OT7ENuVmXlFHoMGIHVij7Xds54hQO5jMMciT2oZ0dxeL9oM9oH+CWsZ6JG
odJ1MMw+qm0OjzdUhfoO8TlxcTkelYfhobI4AedfN5AWmDpcCZbIpCyXCH7WF4T5
KmzIh3Avkz7BQvCV14yWZ/X2B/5PP4vH/+81Z8s4wZDNFeopAM5/NulPEKAp90WW
rUKz+NHrpeNG1CF6RhEoCE5ZlVvqZofVDLgF271RcUUVmFOg9+8e6lYvtzlR+72E
ORpngHmVgR1VTsUiiFw/L8CAdrZfZWZ1ltlC6vBlaKGpsJ2txxw4Zs9hzwZXOsMB
ueEtAMpQE+PYN7oSSOhhpVA0Si2pI6lsxaRVGxKGzLyekF2Pg6+7WYVHsTfQbimU
YEmF5aKsZBjjWe0sijSLKlyCsuJT0Es5arNYLIl2ULcAC4n2u+X2Ot7K2AheOrNp
IBrRtlO7sdraC99GTVZLyd3UV9yCWeAKRvl92dTmR2nFgQL+BCbdWb8PlL91pj2w
dB7+aDjaE3rF0I6skqYvAxGXoEkU/HmfsIF5K8pDPnU8TwRVpDG26+QuoRNV4PL3
UyfTVkMfXYVbbGoRgf1U+gB/qU9PFM/7rVD4H8NQKGEm9HMSHotVugO6jPSLluXf
ViBVar72hnNsLShz4kN+fiXX/QfzBgsCeGgyMnot1/LS4Kq7rAOXphp3UvfwSu3o
ZvIVvVCGQ/fP8ItQeemY6OqljlmshHC+QYtM4VDIgRJLjN064HQLFeyn0JSQ2K6i
E5vxeYZEbNAPfM6ZMJEXJ4cqoEGA9AeQJ90cXDKyJNU8q2sf+RXef/1OxUGkkkUL
kejs4rqRwe2b8pNenRyI0sUCvhtQ5QLCg8CmDcTUa8iIdUrONSAENjDppbBdeDx7
N7NzFbolYIjo++iddr4fOJsbyyENVW7FrzD7I6e7MsinpfQS0ar1CF9aCwLbcnlW
TsoZnJm2dPdieeHT9bjwCqTlR9ulKBCSxa0kdilzBKyD/K8XJaGFdks4OF1zcEtD
Tp1qp01m4y8bbq3JLE4pR7yTaqszEJn92bLOjLSjYzoGhNFC1nG/scKUYKLM+Lvu
4sf8ghiCrCcpK/VCppHWAi7JQfiPYxYl5xaOq8YqPDKRb1TnoAJj5ew0mhmRx/4Y
lQ/34x0bhClD7c9zEp82QyCtWJViqCQZxQG1CVsP8GFj0zF3pavrEg0wGBY7Kv/+
rv7UBihRl45AbU3dsm3e9zpRzKHTtmvYhRYGwlXElj2dpTI9obtTxAcjUTmjRlPV
/bj3psBSPtOK0aAfFbViLo5DZHbBz6djdN8Rgv/GO9Jo5cZoB2UmjGJUxB3Yvbxw
Ylv1/CN3qSeCCosA25JOIDV3ebFt3V0f54+GgNWNa1w5//QprWQqEygV+BuQFOnV
s/PI8GZZU8mPYAKBqZiw4wxHGkUT258wjLbCimLV8KBOFWweuqadePVkoLczt50/
Mwc4Rs8oNVhv5QjQZiZBgkaKGGZ4NNYYTL0r25Bsbm9vvHZ84zUvY2fPKeSEDL3S
T6XUz6AoSE3vSnENcXW/VCNljqmW+QAqwzwIzjhc159JrfZKqIR6E3jp1b54oanC
MaRk09CAZC4NjZ0PwCATvqL6qD5YS7rKwExVheUL8n23yMQT5hXXyg3AhjuQHnXt
GTO+yrZqT69EztXZUlCEj5j7qAQte5qZVxD6v7SZhpVJHArToM1ZCTE7VK6dcGAO
IFqhN977NgkDySYeoVrAM3hL7iQzyL4rHKzH31Wu32oEWlNGDX6z6NspeqdXFzkT
Wy9OxDdxezTe8gnFxpYSIcESTC+/KYHAKrOSLW1SUa4Alw4gq0W4x/wf48OL2SY6
YcIgg/lEyurVzNM+4qCZmjQzWomcdZ04dkdVUOPJiK0VE/keIzMHkvyoZIz66Xch
st/D9gKLsNE5K4B+htcKUF5d6oHAscpAC6reNEzBYroOMObI01H27TtuR1obNOlJ
yA30fC5gUHQa8NurejMcKlJCtsnWv8kmMw727SPCSBJq14omloI6/KHKMwhkEgdN
n5ks0CXqR7TUhwWXTCfN9tWVktEXMvuMfXkSi/AI/QgJ1dq3UqxyGuIAsiotE8/D
0Y+LkpX8CQKe/Gq3epbqxeqmHgSKSFRV0Qla8Oors9kmLhwHdCsYEhdbVxtOUux0
YjQuAOaJZ+d7zynsrG59pC4PdQHj79nQ8o0xeFRVUXm6sW2G9hisEP1LT+Q+pI4K
gj8maOXq7CHj2YP3+7nYnVbu2/FJ/yfEL3hj12ZiK5d5EPggk5CxybjQncZnbVs6
+daCuy2L/wnD9wx/I4jAiRfAYDWcEM588U9YGBg6BTahDwPpDx1kAd/mU0Xl38g3
nQwQXNzYLuc/b8EPhBqPRNJPRSYRJWp2durqiO9QP7M+m6dRDia0+ml2Lf6J9xjh
rHrDTWeu9zZKj2tpdeiRMJJnMPZBnyWdQUOMEtkY1b7XcojNAq6JiCjqvRe0CIax
Z857u2tmAaUVoPSezjfVcgCI4pPxXwg1oQh7bZa0945EyOp+MAJzDAfQ9gOaxRcY
oUTJe6H0eHL1P6M0zc5sjfwSIhZzsPX+NcB0lJzQSreaYZQ5EiBW1hOjcooNKyWJ
2Jp97ejM1eXsnGCCK4W8zmSAjNY5z2OAlE8+lvyyKodzWDi0PH8cyWEONP08ppGU
iEGlwIVJQZ6mEHYUgNzvTJlx4rReJ78PniLvtNlaPmjjqniZjJQdWN0j65JhfSqo
I5xNmzAhKyb2T5MncD6StudUEdnHMzj3Uv92tJA575PtBnToWOGM4/Z9V9SdJ4Wp
PboES5pYcdIpjQFn3gK1W1mbHJDD/xdYGLYLLlpzd8yxyQjvOcTr5KA+DRv6YjRz
UdKF+LKvnm6nuFoz0fxpup3CCuciaZhj5bw0z9OgBZwPR/MIliMx2VGZ5hSqSHyf
TnTVhfzXTXJBV+5QQxKmK/K3fsWNuwBAk+KotTkawpeYC8+1WZj8ePq9KJbF7ZrQ
8PRtdluTZBm07E30KFLOIDUmxP4zLeQsEhkyitIlE0ZlFWv8dgO2tWUyo9UDJyyI
eU0Gxkvty44hE+jUwNdbmEbEpEz5wpe1I2v98aSvsduaSOggRP90eJxLIJkRk+uO
hIeIVpuHx09Vu7BoKygwOqIWSGYpuNiuNr+mQOR8R8/KFvdbqhm+D8/XNWjuJ2YZ
RVb8PqIakKKyHx7VqcbIjvBHYWSsevv3lNZ0ALxYZZHDpwc1LxBV8cK8v+A3/SIB
DkwaAelkUmADXgIjlN49B5q05RLm/oYy3Hx21ATxjBFcVVq4Mg9WgHePM7m41chC
7dtKs4dS75kXyQ6a6QibOQ/DuRIuUJ4upF0nxeZ5alISjzEGHcC3+Dp/DMwTsGRM
K9QOFhi2eORhx811eB4gnGitEQ7+bxtqYuFpk1QhH4YpuhuwPJY01JTbnYZyZjDX
ex89cCZS+ACfzYOyaujSyqPj7fhRLiP53Il19u/kzvS47JnVfQ59QIiXk/XXLCw3
gngm3KOQA4NDnT+V5ecTeNqL4+0DxReF/0bzu6KawH2PTpDMm3UhvQqZRVvOH5Q+
ZsHUHhf7BxliPhIiowTC9thsZnAGtCMyoGwMcUtH5q/xuHPL/yWmHWN/TpYoigiQ
AmbUNClmlAKk6wbXMhM/5Mpm/ITLYqQcuwkUMPrbJME9bBCdVYa0Em7+wnmfENoB
WoWkBvekgAYDyuQbD5wsAFPB2W+oS5TnAxMu7feFrNpoUpLdeftP7aaByh5/s7uj
8VM5JZii3d4KHoC6W/Zilz1+wa7SflZ+AkVfxQ6NTXKB2vEOOtTcKBslZSXmECo9
vO6rMdNgcBMjngZc1Zw+GiaQr3r2y3hXn5C0w64w9tK2Gs9M6s8SWcPSveUHj8hj
M5JAKhRrY/5jZHoDj3KhNMKaN7a/mszyFocvFdV07i6gwJQdYzU0M1ygURCs9BXC
pji7d7/X/bWXEUL1u3u1UVQYUK44d/Jl8mRhDs4CWc6sosoFb6xXUjRHl2Ym7VCC
584lSGrETDgvaMKnUibgJOBtilpkln7BxsO9I2B1mPqV/kFxojLBU0s0bf3cW3du
0wxKsP7EGryA5w4uQGedJT+Z6QdZYCC5lHpPS9UkjsJ6ZanKusg3usibFEpnmTDS
wImuB1EiC7FZPi41fF4kSTGo6ioj+/8Das16v53Hozj8b5codZiJEa1VcDsrxOHe
ivnKcPx0qYr0RxTy0iCl4H5woVHo4BaY0cXhk10e5Oz3YgNfR+affpR+lQoRxpWq
hzXeSxdjmUjoKnwnOfem+I1WmyFotakDJFILzF/RmPMKVMP6Rh59FOmtkZHAIRyJ
b5XKXc3BBHPrfYAZYWWU6z2bNz87a6GPJl9mKRca/U3mK06z/PaH3AV3C7MXVdKj
+Zc13TAZHpb/9E4PfuyCL6xbawA4I3XbunWe6JA9rTPP1yzG99gADrf0qiS9wpFi
fS8DHa9yisZI1W42OOr9nYVSZ5pak5Use69dVjD9yXgEhFaNpwDvmWUHuWkoR1q5
2TizQOfracGaTzs1DmNPPemh1KUuz1tbWxZVslBPtcpRXJ5U/X29reOF+AgjLEz9
CdqCMCI0MvsIEbaP08ke5BCiT+mAUy2xr9PgSZa/37J42v39El0KbqPiDc6BKBgv
Ls88iFb63P8hfwprRa7czmSNDHcHc8/3ZxGP3bFWk8pJ1vkl1yMzePdlH9S+bhlf
6omTdgKWzl/GKxNhf8I63ehnnS+DLqaa7CXzvkoh/CKxrm5W1yIfdqXHe/9Bmugf
Rj/ug/X4WmyGQ9/cFDt+wlQxU/O81MdGFr2I65kM8E593IOHvrRjCioy3SokraLc
oPlBPgyFd1NiXmY3z8/lPwtlExQEqPdl4oP1AXoGFqkowsOtQjMxRB3Mz80NUa5A
MDuEYbocvHR04b7eOFSWSo4TkYtp8fW8mGEyWzZC7EwBFu+y1aW0+BuF+Y4/LFcK
K+/rA5vW5IJW7ESiQmQRNV+WlkmyXdHM+r2oEN7jr9ZBLyeeDwSPXKZxI9tdrtpF
Ps0T+j5W6BrznGz7BZxilIcTri1ZJz3o5KaSBOWFblBsbGWGkvcQB9D+yYqpbCy5
t1D92yM/BFeZHQCTN2GI9hDhe83GuaBdu0uqUXGihqUSLbucbERjzozfAXfuiwbI
lGMTQGtuGhK4v9aOp1Xj0MvW596a18MJ4VfOdIBEQm0y1/5PLtpG4diHRDk1kAN8
18txUP7GZfvAcfswfin5Rrff+q/pxqASBxEhZIjihG+0TyGZw/CfXt2xzo6/VVmL
Fr2us/wvKBSuPf0MR4jAzb9Pls+H2EXNnE3QdyBW/C3oS53oaBPiIGGtDPWN29cr
qQ2Cs43KISnMZARgqyi7SzKl020+m+VkY1z+nBXeDdgbTgW3Rhi7kaw/OmzO8Wlv
ERk9ou7J8KcLjXnyl3hVq55FB0vgWrDjl3dENhYju01n9jC8/N6aRkeqcxY2mt5U
oVSsq9CD+nosRMZUnyeB353oI1mW3QQfw5DmdKIoaEcXPdLOIqT8TfBdFq20jIZa
Zl5uowkIQNPRZSjcis0WJsK1MZUmCTwx+HwAk3NUiX70ixHZQtv7zCA6TjHVcVpC
3QgMwYawkLmU/3/DNcY3k/WCGlCu1vz3RXlnPo2D/0rkvRTZo/0dlIQ3d+WkrWw7
nVYEhNg3v/kuURYMil2mFdZTILoU8xRRKMIRnDlm15+n3YthbxG0nN6vIbI/gHrg
CkiP64WLyfZW035NTlVBvJg51WkPX5owzikKFG3yR3W68KgFEvpz+ytBXf2aYtme
AmRPAEwmcOYXHCF6ALxCnnMzNef7+9Qa7H8smo4DlzQXNC01ww2aallXRk2YbXsM
mt4UYwgz29aEkN6mhkS/VxJ7ebCpSSpPbo2KD/Qx92ZBIZxe2ETpUXYcneEW5fFR
735MdX6/tMAZdRAcnF/5lB1owvurCDz2e6BQ+KTf04xJqC5uAvUpyztA5YyYS5gD
UR2HK/Ns+1pcsj2drdwRqq3HS6PQ+iJ37Ys3D7+wre8OmJGtLtyUDNzdfPjJ39xf
MGJ04kcEXe6vTjX4fLQSIKl14o0fNIaHVKDNz34rkYU+kkOAA5D0kLHHcV8pMPXJ
kkzlqLPZ+pGebFDYWpZmCiVDK6DaI+6rcqPjA22g4v5pFJjQwk1HF59O65E8pcmF
RN1YKgDpsv8Vkc1L2eIkkkimFg9DTf+B8m7Ek91ho5bQjztgLbNtg+QFxHPE303t
M/NV1oJ9QzzZpmOanrmQp988fYSWZak7AZhWuD+C1Ewn9f2vMv1jHAfoy0c+Snip
XwIx8dgdtiIxYMuDJZR+uFCyMP4KuLJ1+3zIZx1LCwKecZBH14032E2vkfMuP0lQ
mVFfR4PwdJ9NOjreQ9RbW0Dajz2RSfquufzsMsJrTZMpHXltQCGAdXqV40eGP6T/
Lhac3TCyQhO/aim2neeFkXvAtlH/0PQ4PXw0rJ6v/vEyMsCq7K9NwFVg49gte1St
QI7YlQPSbxC+B+FG9/hIw+q8hfATLwTfJJznnJuPja4OWsnTR6ARy+Lx1EMq/xDj
AHZUDi38QedrTnXQM4aqcy82sEOMTuoSYDhqs6e61mtcNuUZHtw/rvzZhWyia7+d
tx0YkSs8x+Z+Zgoh0mjK8F/v4bEe0/bdBHl/5bgdHjgdCc+3uhRHZ7qLqS+YlwbF
x5vCBoEDDmzVQJ1DKi3SPxTzRMQXmqPGcXawLFnZffTaNccmLOqpDeKpPk9LgRV8
7AVYSlkQe4tpEnvtCcRUbRzkt5BzggEyswXIO+602rIu1cKacj0I2D3/y332Z1jC
90YXL6fjscdjg++sMm1cSqIsNy8NMm0iKrE2ONy1lGy28K/RQ9pKMm13VljStTgO
grDHsdxRwfgIhIQzQ6uCcYRNePNv4r+zF5fiY1N16uweqAQs/3NdysBvIEANL/t5
GTLRPAgMIulknYCQ4Hd2kutZ5t04GayqDEaKLjtOKA4DGEMx+6jI6/BeKBTgETm9
a0ba9giDXou4bPwy4YzASW6g2hsWkRdl2IcN1xeCohtIz057THEPugf9iTeM2Rwx
f6kbO0lwoedzhYknHV/icn+R4AlIw0Zm912xUSpS8Q9fxdBvrwW4pdmtPK9lVlO6
esoqd/YYIcYO/XH4akS4bYWd5BFM9WdLI1WTkyEQnfl2VnKIagEqyhRNQVCmhuzD
kl76+iUU6T0v00kfa+meoFCwlwhh4yB0bQjQayZ5LI+NaAS09aStxmM7LPBVaqmx
UwdEj1AzFbHok1ztImdzDwWwq7seg0tTA7gaQs9L4nxf39462NbWoQZad7cw6wDy
mntZ/PgKdgqminlpdPcopPN9e9pJlNSJzC2oGygO/eABu+V8VieGSsX+54C12VgF
ZjHc/Ssue03BiBzknPyoyXWnoitZopMKkycMONIJmHO/73TOIH6xHImvwWa45kv1
yQXwGVoZ3CRisy9k1ki7ic5CV5JvZGTEeJsa/Kynk7SN/kwNNA4veHBEkpkWapBK
k0cZmoMTw5ZBmXFCA2ujvm0ddNbo3Os5ux5O+ZDdfITkzy/zAh7U+zhL9CNjpuha
MY3P9kwRw7VoGUEyg17Jdt5UEdpKvIOtkBtTJn8tGlx0Gul3eQ5fmgHj1S+ZK5Nh
1Q9mpf2CcBt6Gshlv9zYoMo4WDQfJxvON99Bb5Hr9KFq/NJfGSfQwohojgqWO/t3
dnTVXnU6LRK8uHykHfINVWSwmiU6Lnn3exYq93ke1LgxF82Za8zbULgHO0MRzAoT
0H76s5bYo9fCmmBNe4I8MzjBwA8/3JrVffeGsiU5ibu98qTRXOFZfQntrXDAkQWD
/ci0u+dVfp5fJjSisqHtQEMhdvRCALSACizmhfcjONAt8pFqfLm+tPi9lARjHArn
Jyj+8IIe8SXcUbL2E2vngZoWw72BnYIdOQ/WwEWEoK4jUZpDMHBADQCODNFvZFtL
S57R2vWQ2JmOJoMSVY+ObSXJ3Tj/U9mSUWsBKq+J+n0sES5AZpW6bbroI3o+KoED
nVWVtSFnP5tto9DGFwUAfX7Bo0SZAz54flv3UNcy7FKdOnXZvndGj5h50HjxKLWX
Px++retQMfol/ZuuqMI5pYQJaeUo+rof4kxM8pgVJke+r5RDC5ONrrs4HqpX++z1
mD2CUMtApjiEE9MwWd8iq7vjBGLNJMhUBnsFng15OG6dscxb2luOesgeuwhAwY3L
Lnd27wiB072G6RBVyzaZ5oL+/iwnIY5DZDizWdTSaZvrb2zJPHlx9yv2T3KO4qSq
QM4O3XAsrv1qZqTFjGClrruycAMJJiYtDIhAF3Uvql2pFSHdi3bTzic2xf9NWNdC
1lurlom1GoARzJYw03r6W0oVCmqvN3zwCANrCs5uj2Zb5mlwzUEzAQKhHbLuGJhU
zOwuc7a0ng71Xe2MXnijoZvS/WhX60qpw+ve2iTcBtrCu/MsyNZZ6WrMiZE9OPAg
SVtANCuyhWR8Kg3alTwsLAJoRR+mReyzW41oTlXnJJNrxf6JseH993lVd4XhMfGR
N/LBpmYpLwmTwjqWuJ0R9Pwq4i1oz4rMRHh5F6QJYIyjZEuXy4nOBl+4z43St2Yc
6dqi97f8/HYFNDms3vf0toPn56FeAOCIIXeb6R6VG0bj1x4RyLPhdfCCiXqwrH2D
y34n8lAx2aADsuY/zxHYRWMhO91RJQsTtdrVqAf0yg4U3WMYRrF8zG2G/tyw9nFl
o8C6qByBtiCYTOGLAcVvmNdo46yb+4AsL2O7/cmgqMWt72h3ULafZl58A1FiyExb
faxDQFTyht98WgDGGHaRlUhoVXkuIv7dtaEERIZe2Aa6Z7XlmnoinP+XiaPCyItI
bvbdQWFNhkti4ecrz/MkN5lZXTVt43SqayKOFEJHsfgU0lDAK/nqtHPeL96CNbva
+FuqUIudiY7I+bxSW3MUsKS3L49tPQA7zz+3lTdY/gNRcwmWFbBbKn1nfJIJXBmy
IosRs2UwySODHITlJ7xXWR73RszYjQK2M1Yuj1PKmz1H86sv1OqF4ppQZVqeaYI/
C/uLIPkdE9/uUrCgUuK9T5OpZJXXfxYoyUvhXZrfiPZ/ZgEvydmrFwqf7aswG/Xm
Et7qLLaiXjFga8UYuzUmdsOxoe4LSjWWH/rElxdZI+45y6sDuxjDT0wteyzUTfA7
r2yypnqd7wabtVi9GcGHfS0oV00t5Nnron8/nJzfUkihaxOKe4NlKaPBa639Ics7
aYwGr/TxDaUt934Gg37RjJCooGULiCldhxN5rZx8+iMsjpOprhDk5uYmQ8Eny8LD
84nzJSdk42nhjrhXVXw6CZ6Z8vjjpZVtPXaKrv3If2rqvUkfao1j9CCjv/HQ9OrP
xMLly6Tr31AMJkALa8tdw887S642lzOWjMRmpzPOEcmvm5afvxrzD0xjH4Hl3xMu
2qsTiW6CAOn+um0fQDljhRtP8GVKZW2Ki6mvDu18COnGJXko1Y1HZxtUyX7dWxmG
8+JWc6AXhlYxflLd5X2PfIFt7ttmfaIw3OdowpLQ2YmSDajmuPXfl50aDDxinY2P
Gesy/elEqjkRwKCNrwJfkoB4BWx9iVghRvWattpor809N1ybgXLNQ0+GE28bXFS7
2zbj+UK9Da3TnH7licjhk6tCxaB84MA17NxAj7QZPJCAJTmsB/faiE9iBrCelf4x
YGDiFuZQ18yzBtXYfwUbTJtignEyqO7zJuurnjb8zzIxsWUO2r7kTTSneVWtN3cU
QDy1yWVJPp9qLHmIUORJUvu8CMNEdUNdqcyWYODqiVTZbaJEA9AEvG2ZrxXZe7yO
ucnlDOaPnzNZB2Qf8qNkudGW2u4or+RNT2B+HtfIWgvFQw1+WpXNJD30dKMCgpmK
TsYsMmKsbAJ5ngWY0kMIFZXDv+tSjrO7VwUPddA5YN8YBR3XDj/AxT2ziMWDwDk2
kOxAnpplQeyRhv9s8hJDR02ZYAYgupGv8OywhTNyCET4kWXxnAQz11pYAFZLgZTn
3DxBfWbUtp01DAu084s+INc7MQ/IobIAUwT9xnQiGxj9a0irJBzGmuYZELAlyhc6
Gwa70s2WwuVNohOncFytTcTrXcMiirpDYBJxo343aleuFzomA7rVeMKjgWSINnvG
J/3sVmWVptJAhIHzpYT6s/ibdBKsysKXF+tiUmmnfP5y7K/Vx+RHFVMwykz+JZ71
olM/HeqKh6uIjenNeKxrVip7WxXKF17LjmQ2jBAa6GGo4Z4fzXTykbJF3kiZuDx0
QnUyhXoOH7kvsBhFMvjZmW/QEkWaBHOX4Mh/+52Dabt/K+gPRu3vhZaHIAwHGpwB
fXxk7yK78tOpMsf9auZIwUZ37O+OMn5gJRap9AUTObmNzvjN9diqkLhCd93c1QFV
1oQGse2I9qNbmJkoFeuf6maXs0lXsL4SVku4Dn0qkqKhMkkdxrtVAOJFaTYI0yW2
+H0J1OuLqBPiwG38aEk8thcqhXwVCiUrrQ1S26e5shy44ZiVwyBY7FepeYPA1Qim
r5fzhsCPR+BCkIA9smF+FBNJojJT/WFaTKo/xGKuhAYtvl7kdYzchOzFQ1wUBYfu
Fmju1uXmZsAOP2ybcAMdIJq1PIapp901PO11DSnMaSdi8ZH3LfSpqlqV8PVmOAMN
z+LAYlwFffX0MxPiGh/jXn8Z1ChQMUD/Qzzi8t0/mDdmqtKzotk3Gowp1QWxxtSY
TnM39TnO8fiyRLdp/GBGpgGyzKcSdH1gG7u6vMKtlU3QaY32ypTKGZYRug2hnZ+s
dJN1Puk2wAnSjgMmn872OTZ5iKobWthtoXVhHF6KnZtL2zug0FisPhmWttfw+4wU
jdEvJgednniHG+KowCbaw7zrWjqs3S5WMW5y+RBiGvm8HHvtFgRgxfK/lrdKzsc+
Mrf52mDpfvsQ/eptSWpfJ8FKa8ZQeatbZ4KWhtS28RUjGrvJktbls/FzlfGoqx9b
BkdHArOXVvKSrqTHfVo/UdO3R5/XoLMNX4yZ5eOGtMk6uHYt8zzTLewkjslSJxXv
y4/0SWqs/6AsohY76XaY953ei7URGHzd+ZshJYyX0fyVQuM6KEjSnctYtj0pJ6+c
1xkNPepH6wapfpUhBoaiiKZ3CKaUScDtCDC2BKtqxLm3EOgjJML6j8MzSe0AEHXx
2ZzVYctdfJCsbJLxn1S4r5+3V3phhlvRsTwQQx2v/YnHQQ3Z7Qw2IbE6DO0PQY98
BxPmAX+0Q8bWAf+CQz0yhoQa3pi5su3pQEx7yXazAcFj2rpmxFvF7VbL2Ry3AHNE
cSrH7esC7CJqW4L82zVsj2ox2fXZq7Eecsp5wV985eayF6ONDZZSth0N5m4yhm1c
2QQcK5r+ZpibalaVAKqNoNy7t5g+PWqfI6pYJAD60PYPyLilkMq9FsxrBs0OYJHp
Y8cqy8HiPy1KctWjlDUu1Lf3pSNS1GMMPvySLSevKlaDU2XnHncfzOkrfvETf5II
4O2VZwYKyNDhUctrpjZc57YSc9KPVnK3kCxN/bFm85W/Kfxx3bB5Kt1LdG4GsTj0
SzkA+eWB3+/V5bFc90gOx0a6y5cooevnU+KYLAIgrdVOfjqyA6iXLzaNxr8SB4Mv
woZjb9h6TFdN4d2NltSkjfdMcrklZ7umGh4G7O5QYacquTod3Z7vI8wdAFKU2/Wo
QCaWaIjFW7nd6ITOFLZ1PnDnSA7gZiSy5dD84a1cHpibnyjv5n/LLWnlHEKXT1tN
tnMTpY91qFcxFvyxQNNK10K4XhTiCxybzytOWxHmRLXpPiLHHp3eohL7Tul20fcR
4SdxQQ/sdjXfxt1UZ4a40ZJX6igrdmQS5pYx7XObA/R9CwjZ0kA/SkUrPgSRKznW
S9KtmGZgj411wWgojqHk/TW+Pvnnwd83KDjeu9ZgdjNG4Mr648Y0zXnTlmgonDaF
tz2EP9s7/3/hZgj5yzl7EmWRSLGqvaFCZMJ5MS90Uiie2e2U0ZOaUyDjbllKll3T
NysYv8NpNdk+5grecm3s45SUifwVNifuDT5S3QeUa6Uc9PNuhE95O1ZviuAWLD2n
2spjOs4XTAe0G5IpXGbfV0xy42mA7miEv3NzBfzYrF5VcvVCzLQYBLsX3zm4t9Uq
aJbszeIQnaS5bhOHMT7YvPpHfp+d52YeONDbi8AkBXicg6daVaNBUhbxTBUBvpR2
1ZjGZd2fLdbo0eAyLj8nJz/IaQFgEcdgsghKRrjJp48Bn5g/vWgNn8oriVWl89p3
REb5z2md7pBQLa4n1BQ0JZvzPACbqKt94nVPxnAX2SmsewGOYfNUweqbVcTXMqr8
vwVwYFHpT0yhSz500kya6Etyh8t1ZGLV4U3PyklmsXvSGFEryQvmrCA7O2DNea8f
9Oo2D6C8Yh/2m1VriPFyY5H/b9C/8HdSyLTlDPUt9SAyfogI8uA+2XkZmZF0xl83
NkKkTX3AGyTSeELrINaHWo8FeC7P38KWgkDUNbXCcIO1WK9J8QCN+LH1mnuqjISD
F0cdRbWNAKGSurhiS2D9v0i3S33CJ+zcu8sCzT1ldXbgEfup8e0sHY3cEJUue6Wp
MKyMablcL3SPfmsbwU3Af26wtqkXNQVDZwuqTfdgs2ca4FpyXTCMx1vlHr0M8aws
l0S3m1YSakRD5P0J1PDmEQ+mwjDl3vHWW0NMP2syD8PNuU1zAJVfe+algY21hYXH
X56bBLBBKA4F+ZqvhIDmqOuo1RBY/O1zQispH0oGUejLs90wi1D9HZDjhEEG3szN
34D1ctOza1iX81Q7fTdofSzffvuaEbA9Idn7MpCQG0DWs4xs4FKHQuaCoJOSUkzE
yPxp4xIbAHgL7ErL06BBPAiTgIms2Ff7hBWoktKs+LMCnbZhzobqmNV61T740xSM
8HmhCLoJ1PzNOvJqKJG1woPrkKtuBYBctyWKkCyEuYjHDzA/qKis8eFR2ZLlUGmx
FxAejo20zAX9VnkXTK/QREMU6DITRUDM8lB56+kCP3EkM5DrN/NX+fzQLx6+Erue
Tt7xM7BDlEtthGp6CYsKEZOkb/b5hK32my1dL6IgfQ8QZTQfUcFxJqeSomVm8LED
eZo08sfMKIhREJXUwwHV21eGeVUZgbO6jqIVPxNnMK0Q15ZqDUMbP36Ne3ovPilJ
A7PLiENkBO+Lh3/P2fhl70jXwoWzz8Sfmv8+wgiPWK1joHzNqsqO4PaPDuUG6xLX
aepNCovJTEtxqtqfQ/bjihBhztGBxbvyUSYj3iQNINrncR6wfGDOZFdfMrprJgvL
4RzNtjVED98dERQVWwiFY3NH22k9W6tpf/K+kO7qhS+QOKe800Q7xTRaehva6PMl
4OlHXCKyMizDi+A+MFY0Tvt3WlsIddsxLGuWpDCO2wy83kfoq0DpFux21+Ck1YFR
I8tuSuGftVoiKFlErt4ym0jN/YTdF3Ozj5wcNXNhNmzyuWHBjgK8Ujpoef2L7RZn
zVS5DRyfYMHRRY4F2cuEaArqXsT5S4fltP4gIm2Fo9f4RpXpdw/vFmV4NrvhLAa/
HmqpcXXn3O9tqd6K3mHv0Jo9dO9Dgf5DGCAG6L0IBXZfU35zBTU1rL3/NMum20aR
JvhHiFAd3AkkfOpcC+IU85O+50nyK2+mdo3V5/KrCY5mbF1WjEEPxYJQKntDWp9G
4bpv0RZp1TaHu4LmLhbtTYeV+YUDm0v7KXlzMY2ikKjJp+Kh56WzmC1/gPGMX4ul
eTrXj4h/K2VlEOCcmcW64MVMqwv8mX+AKsrm36HQFiUjcrB/5v61XLqzuBKYKe1J
vDpAjA2jS1PLnGScuWQFfwLZx0/GTT61DwNGlnCHmpY0QHCejRLrh9AHuziS4o+n
eoO+Rt76xFdBuIwFIpW01rZQwi1VObQH9JmvUmenDq2458HkZF1JDdEk4lsYRs3e
w291WocuHnpM3X1pLtgPfnvgbFlDFOOutqqw1kvCfCTPrl7DFTLeGm/JuagxuzdZ
VOmeqsKdDpibrUemosZq4NBWLJ9koZhPj1KCIDW+toAvhMtPLYChQi8flO/EtFLT
Ad0QTjuvmEbfDyFrh7Yw4FTCZgXAV4pq4UCSp56beVlEMYFJas+gNS5ck11w6MJH
N6JbMlxxa46JhHh6CqQJcWSUp5AeOksIEh39owjZZHgUrffh4bNG9rnLFF606I3O
EHj7fawhVQmBVt5lM54F2ld2mwM/36UgCMjpCqR25UsRGjnkgjU5GBXH35yMXDms
GxBNdnbiSSMZahewhFCs9qrAOOir7EBs0T/xSpN+BAU5gWEtMjEXg+Igw80UAcHI
BXsQcFf4QmzOLU/Mac7ft7sUMzvBqLKluWwfHm0RCW4SVWFJNKHIcx4yn86GWe/7
NdCXHUqTrfEWav2Cdh7oUAZLKOMozfpZZqJLoiFdL+MORl5XD6hd6z51/QpZgNcT
9ucpPk3qFGSOicujnLPr8zkjjy6vJxrDXcG9JbVPn6BAwQ4/2tMrMNftgt64jecA
BJ9CMABZFctRDBwLw/rxVAWmoWl30th8EBv/7WdVZ18TzPsWqbrpmofsDo+ZNWDk
K13akUaxkKsUSfBj0My3s3y/qqknhzHRLDmeotw+KPaVlRB6qy8ORJL8yXLGW9E/
IjTATucWF/QWCuqEg/2oTK1r0kVu3s8vtz3Z/XoaTZenjq+4uGPB7HA+A7m6BP4t
wlJwIdtw/svZJXIyLvuM1eNHTBkDQqTWKDdJEClP6Sw9LoR8swSiK5eyH2SLQsnd
yw+ThdLvQtpO8e//KD101kYkserEKjEUKP3It3jmu4ivBX6YBo4fxBpdHhGI8Olu
09ci/CjQN6jf9K7JdLSbGEpDt9XDFYFjSLHXcnb71BYznnSU5TnA6OTlKIotf+o7
lWjuhI2tLmTDw4HtGJDrhV4wzDiRX4Pe5K9MGum6ZXB0sZMR7HmUoOJac0OA7wD+
trCDyHhD/3CIhxA4N0E4axGnd9ozp48+rHOpH5j1guhWiyLCjo142IFU75WwFjil
N2gB5r9GtRU+rk96tezXqiFeecOijwAfwQt6EGfre5Cz+EjqFixl+9YSu8dNOmUI
9GRPi3HL5JsC6ATiV/yNOIX5CVDtQVBRxKa4hfkSyPCb+IX+8dJYgyGF46MdsuST
zHiuUe8lMuJkqi+t2iceqAtXVxjzkxb8jHiuFuogbiVkDNpHoJcEq3eSX1iZZiMd
MxRmUhcih9dsPPILgIjNbxUDSHUCqaLMSP/7Xcy71okza+W7k4MqQ9taGmJ/RRRt
PKcoObTu7QwLIvmZD+fGHeR1rsJHKJ3YMVIdxi5DJwnjPRITINbgwXznvFvZBg7C
wrCtLTomdsptR0fW50uTVQfDAQ2sXIWHLq3Kvc8tpv1PO99arWSP/jNDiF+VWQTB
bybC9mvieXQnz7wLoQ2MziPJlKqztrhyTGjMvUBn/30vCoAocya+OLz/54yWp6gx
IcupfKhXrOu7UY4CjwbxDuAqQLSaM+KHaIx8ZFr79YZ3wtELx+JMrsZVwT8k5+d2
SiUvuz2TXSkyXbRdSY+Gr/aZw8DMM6d2T0IXRa4R/PdNl/6upFHoBDeVifQqZ85x
aQtt68nJRZWVU1l1tdfdzoPStqHDMkxFWbIbuBF3b1uUzI4deZrb99aR1hvFTYjz
FJ+K4UxAj42VuGPElUEmkQjmrExpn5jTGRK48BVEdms0IrvLNh8P5qGIzElY1Lz+
kKs90lmGpi+5PAI682evgPf/XUg7IlwAo7dtneL+lMmC89RBfjS2lGpeAZeqUIhR
UOiB87elpYQ16l13JnB1aG9578SqXhCIUazOGym5mqgh3gL6FpFP5j3btFZDq7WL
Y+PY0HDFv8ycjSAxKGWb6Vgv6H4AZ5YaoottvSQhjv55vHNqR6QE7GjW86wS9rEb
qyguUJDAPvJFWV+w59vjjJK2Euaje6iYL8L1eSHCuD7L7jvRbnj4T4RbXuANwuKx
AUf29NcuuVsCTYbLrqv9YTwUYPhLWJxwiXwvDt01DRx8LniUt79oziJZ3KeZhuv4
9owqTIPP9G6zlmP7BwF1/m1k84h207QYUk6On/e7+Li0DoldmE0XQXlKaP9uy75j
xoRBdCMvJDk/7aSDL0jBk1jU/9SFYW44uizvspc9OZ8Z9AcCtlkm4WjVkUPy3zcV
rvBxR4f//7V7MUarUTrWbx4uWoVgsE10f0zZQMkZyRI4xAAUxK6Y5u5WT43+rIGs
wwYdpeVynGWKxL7b9bJAH4VvHd+K/1oUs28q0lzoEEQUZuH/Qmy57EFe4gNPx7Qo
0JxQzaGWPX5U+YxuXj8KVccczklrzwkOKWKd/hkdpNJmlK8rjtAm0f6m8vABjeqH
PB5evH+2jPqi7JBVVTFZt5Hmkei1tj0SKp6TKLY1UmZPnDcskHLDXtkn9HMVd0b5
t6QWoKOg/Qgrw0lAB5s/s1evbv3AfcsSXghksLYAxauRK0ilewfEntCcydAw56xF
u5G5HFInmSpmZt8oI5lT1N7s/r+K1lZYimCq6iTg5OrgCpX2CHhCLqnCa20xvkDL
lkDee0Prafkqz5CSxq6/hOHV2dS+u0xm//K6b6I4TY7sYQU40Q5pFelycUxkKLze
d6QERwldAvOoBlUu/bgfL2ThewajZY0Pxp9uPZ+21NPKV6JticLlAQXLyLEteve5
Z2Ld0/Lg2UHvAFg/z8xMmjLsUlAQM5f5khrHXtKoFZeMmOoCq8u+483N5B+Ahwub
s4syz1DBzGVoTorc0UEHdyt5bgLG2pEO0Wvg4u4wtEpGp+NP7zNXM1Yx9YOrCXmD
3CVKZv0zl3nAtQcVYf6JKyrOOoQtDAgfg4+DwqqKlUOp4tLSqyrwB2Y+WMl+Ba8O
6DfxTPF++u7zC/A41o69FLwcPzQHgYbpdoPIwYXGMVOBca2sJBO8XW0CkD6H24st
PUOMQw7tgOI7SO/R9yk9TZ0NsTTtlJymCLfgtLsZm/w3ZZYDNwn2n1dwRGuWK7JF
gXvjTNRPwz+w7NyondjRKtrvB9xpWySTrSIO0q5m6sIyhgDHtwDv87j+4Ps0oFfS
F2GgOtCZIEJEEPdC9wGr3oTmNFsjsMO7ImYRICnFiVrhoy+KIR/iQUz5RucBVCM4
t+mM8N+ueaBq2Owa+t+3PMcKxFMTwQWQRa5lfniNMVzmZjaAFMAZnl9dys+c/sHr
2nrhED1jfPYpPtGcn5QxFvhftFL8h9RWEJD9vFjZqt5K1E70qfKGigGNWXkK87VE
Q5kKzW3HTi3fzcXr7dhETNyMlM16D7hieLXgk+VOHtW8194dJ+lnipaRmAFC7bYx
O9ZnUBMT/OnFQApp/Cic1Gkp5w/ssR/W7Tf7SUyXJQdHQKQq15THtdhNGKKyJ5oM
DaS5d9OLqG/XmCaGNQnKRFlAyO5mkwQ4p+t3Bz7ejktCB9eJgVdksYvwCSyFwYDl
xEyObdf6RH5SKPGOGe/p+DrWlpSiTJM0O0z47c7MSPFXUjBC2BwZCXub3HUS9uP2
ujolg0ns/o5Jj75yYfkdvrQsyYxVzyvyOBe0xcBfRYLQdebd1v5KAoCnoNYqWkuy
vHjaKJw69wub3djcJEoqomxaOOE+X8e0noGJEMT1xHcALwzcUxpTRYlUoNqPX8wi
vGqsI6ffpvNV6E94qEgfTRlN8oOYVYRBaAtOlFwqeDyr4wTVGATi/tAipENTt724
YgYFruCc7314168NP5jrulksCcYgziUJvAPHbED239SxHXHYb8uNNiQ7FcxgwmTt
XsJOQ2eIm1iMTvVjbo0JxCAI2QOGLoQbQhrGOxkabLN+JqZ/VUjLa6mt2EJ6O7mu
kTk+eTWv71iMMUe50rDIvqHEk5myQOtIrDwlEGeELbMhy4nj0o58hmOdHYmG1FZF
RKsV3fLd6xmLnGYuTZx9o/AWrPWyDv64yjJsMX5jx3ipVVaO2Fjpmf8knDOnNxAc
UZOryKF5cdTJp8KWGORn+NeVz2xHKVB0CygYGCkYh7APtqe4FmxBGJtBvCjVu+UU
igZ3p1bkWREk+56f7QreJEQ4+/dy6ljEojBOx3szGCFHfA8iAgTLAHBn8CpqQbvV
s8FgSEmfc9Kylh+0ZelQrO17/4grJFjEuuJ5es/9hkEyNeEsNMPsIMK0PcSe5Ndr
cbW3ihWw0CbQIfg2ZdFzUt6LSuD5+Bw5AkV5+U9H+c3QG1n8K3SaTHR9/K9k/L//
qyi3+lij5eazSUYvbkWMRvW5bvJJ0jJ0Bv0a2ary9hOBXNgypcYMUz4A7ApLO2A7
GCC2CEHzEz4muIBn+7DtqIaga4otN2a4OJjRXHFvB3gyjszewt4fe7Hd6yCxuZ0N
EK8Nytf//4MgjDPVrukmS7TKxbJYslKjDtMkHFCEhJQcS0+lonRjcgSq7AyUQLK2
UocdMNISlwFs41z10L74azgA7OlR8st09MNeCQLqvIpQpN5GYMzHzk7ilNH2cP/x
RulbpQJDje81cr52aist6KzeCG+Rcfxx6VzFddnV2JBF5L/6X3Euh8SifdpdOLda
IlxHJVwu0WNBSPG4pkNKAOgqFXBa6+RyW/XkcmQJtX2XMWvkwJG5qMvCRuj/Ut9X
3IFuLiK/wXEBLFhPrN6O4GADwT2YZ1OqU1Uw4JbfRth8qqSgb7rH2cHwgui65jCU
+92azNeei4WIu3yx8zaHb00O5okNuwKKQPjyfciSF/shMGqPcKOhNQ6yt3hAd3Ne
otFAAt6v1LYtmtWHhoJ8/GSK6WJz3DZsA/Bo9NSTAINE4SYFcB1MWqK1S4Krdghr
lxfwJ28Nw3RiLTxQqVUlWLVSLFYleVkwgA4A4YPhL++iH4Ea/c+f3h+WLMG3ifat
zm1ocjPWZaEFWscAA5vgC1aLPbmC7WSUbyXby1crzVKakQX3WlMnx13SK6AfQOEw
V81OCcBMSxkBcorT4Yap33mah+FEGd4LtJ6i+egWYVhDbPaT1Ia6Wbr4qaqx3r8/
KxW+cDrPhu/55ZN/lMLF/7mGcFTJo4HJ/GRxgUeNPFolrUnAfYDHNiB8D3/9q/lU
bRuasDbrhm7OL9pcp8TvuK7kDl+p5lXVdRIx2vf0voMqAQBMQYaTXIsXOiZxeUXD
Wmb92/53fZrio00Na1LIy6ZoSaV0fTciZAlw2mGOIVgDZhhGFwiVhfO6oTN6Ta1U
SpCtczIlAEvBhxP9YbAxj3wHaDfHEgskfrT3qvJ1qfwcKbMmlK+Sg2y0wW9nPc2n
YKl7qT7f9kX7cSh6ta7a/PgsRxjNvZDXdlxqapVo1MGoCiGGYf4BaqnLmSqTw+V/
zzBwlyQxOHUY/pjkQ/F+e2r5rtdYa18zpY72mUYpfLH5LUDyeZkt23UA/Bnk/5fO
UTjq1eFCRhXny2T33uZQYPOiJR29VIWgV9/J0SNxZPOWlhAjwKfQcHf+6gZsw/+k
mutn21OrOVswhmP+4V74CCWejoD3mno21yrgQ+NSmdfXY/i4pnWb/StSlUiGL92b
sgZAbl9Uk9bwh5nLWPxMM5NwdLqTrX+WZQTe1ennAi8tyDNPd5FJifBN7QFF9nTM
0qxCmEXVFoWqyMP5+YTovVrZEo0jBmlQATNE8amSDTvpBjvD7RvtUYYslj4it0uW
30/UdqjlgLxCy9XWjX1quC3aG5naje00+awrq3t9pqa6MSi9ctaK1h4ypwrJUXau
Be7DiTPlOXlVrSWR5Ynj+kWGP+gk1uxUMP1eAhB/8Sdhciedt2C3RxIkYq+mSzAm
XujOBKA6MC9GBb6bGZN+ttuxCVkJoSZz24b2MoO9yI9FL3EckPV/OG0Kp3rtAMTg
3yTM+unhEA3frI+UUDj7+Apbnb6LRmVfd6FtaxwV7tLkBkuhSWlUeg2C73k/hIw2
GkJnd7s8ls+1whaLlnNcHDwBD/gAkhQ7kJilNHKV6UnXmvE970hkrAhS1detIKnC
VkMhCVd+XHmC38UbB/Yh5o9IjsOZ2ORHL9rmV4rr/gti8bHlsiaADhuy2g6eMIYA
+qUt1KWNK2UAwZAigkikrXLAd4V0qvdLmXwQvc4Tb4ETf/HY1ryIjDm7y7Sr5W+x
Anm42bFxdQgIttPGKwsrCYu787+5PZG/CuVo599GZGRJAYCrcH3mqzHIPPuirOaW
I+jJr6GcqfVRjYdjVa3bFqByO0zySSB/VkswPFXCvQiWHNinw90za+BrCXNkqATb
W5YnxPomWpM1Jaq1H7G4yDiyT0RgeMfkXab/VpjFleOMFgXKBzblpw/79vOzLzf0
URMzbSQyIf1dWBSdJKeWL8KudV6PZlOf6ET8yx5uOJs+F1ud1cbQdM4XIQdKxxkr
3G4txbRmRWYsiUYknBt4UJQ3x/zGJXhltRBEWN+kPvEqeuFdGx64+dXc2TAZsOzv
lsjfkm5DdfkMi3/leq8HsBXYdmN/6c83YHY4COmUKCYh9/Qa4UupgkeKwf0lVggM
UPRxGWBtSkflonW6KF8QxdetBbM3HBSVXzhq++wDqhuSJhv8YDRBYPWiak22fmb1
fpVMV1Cs4Ywi1yqFlR+xnklW12K9je9bK9Nt3oi77b60bgiDjhXDd4IczQt1J7Ol
vX3vVcvbxiNaEfCWwf5YLjlYfU7LipCek+GCXnERbShQDyUOlGzqJAG/HPhjYc4D
qCEs19PCQwqs3qFMTjcZ+lgM2D61jBTyFYhxRTj45dSMMLkTPHS+Au/iAISfozhn
OgdH6mfg8BlPFlfQDrqoIKFIiVZ3kCKr6e+m8XzywIyVppUekqhvvdh7YZ4grL5a
NIwgAN1XIDnH+zOhJ03fq2OnwXDCMU/OBTojBeh8TD75kMSPIyv5nOIjLJu1CrYe
Msn6QgJFLEz9XP3cD+Fx9sp1aYMuoES5eP5SPs7/vjSMrfye05xO0S5G1Qs8SIZE
K+k2TMhVgALheQ9eAG1G7/KCJmgwkj4NRsWLslbEAHQ4RG8l3HwfwM7MMbKEanl/
JNdYnzpUvD0Lo0bWG/334Td3hz5Su9iCKk1NFbPeWXHPQR3DqRiEQVTeepOUJZcd
H9/nApn/t7diLor7WqDXKd/fKNmUPXZfHtigIvYmuv77c4vkdQ9jcK7+PrUaJDSL
XaLXdA8F2PTsO++2bGOYNCZRBTLHSyVkP7Y2WhzS9LUwibslV/vxBBbbPLxIzwKa
stS+nNlXiOzzKG9tp3PO1C5JzEXjuRNvRbSVBsDKsQpGPGNFdwBZj3vyT+Rs5Y47
Ol5G2CLDHzmsLapZqpEYeor3I/UNW/i75AaxVYWxCN06dzvRE47zNhayXhWZ5R1B
zKlx+nrWY+B9EeSACQnbdD/oM8R0nisZfEHsucT2zfR0QwVdb7J/HslUiLHezK2i
b9uyUyTu8Z3TJ/jzWBrtB+44TAnJHa4rD5ICC7I8ISMY2LDoA4tJR7Aa28pObcrj
DZoYTVWPJE2+j5j+7wnswHHEl8e0JxoKLSra/paxDvyAK+Uoqj8msGBAp7LhzfaJ
hCboVbJKO6nS8G4jZ6/Jpwz7/JHHrYCeyVSSTmICVMJGLyUKToYkQZbnlHoh3KiI
V0uPVLoSvl4FD6Ebp3/S6SdTLbqYwxQgoRraD3tO/JeNR0LC6TSGeERiWDkFcg+v
LKTmrNWRP2ugG16FQwabjXavlA6BLM3pKO1luuUICz5HJj4ZIhnRohFTglVbAmEZ
esbN22FN36OZSxhhalCIpMMf6xHYu3h5r7OMUeZvd55iwA7kibVGkUmqh5aSGwGb
DBB4H0l+TQvwl+FfzBv6sVkjyibSqCWkOk8Vi+/VLERXAdGiKSArNbiPxlaXXSIc
Fux9aFUdBe2pCPD73MeQPfb10y6oci9Rl5IDVR1eC/0guQaYIO8OvKZyXt5eQOhR
F6FNUhkVudpravQwW1l8GVDFj9JFyGD/7bJYWXDaqKjnSoYmtSIDIcBJfZk89bwy
6mDjUI8kU/aA1l853Wi8DBuApPkzx1PQmZer2ywE7iV1ZMIxQLk8esjQL5wO144A
hgvb08/GjGXyicGw+cTAfhZ/lX1arh/Kv+5JHOHyZiPERSR84ZuM4aIBA5miwWIs
f4bqobXeDEA4EfmcMkWasPO8vXu0h1i26bi9ZJyICb9vAWmuAy0T5o9jq1t4B/vm
bW4saIa7u0zdXPHyc22Gj5gX3rj7+6FTQHUuMQO3i1VHgB+A9EXmD6LP6oEU7r7o
JLWX3nYIlXueESzSV+Kao0aO6K6G92Qvuy0MQaw3RMDUT4fkXzy9wuwriyhkIHxx
o2JjMH4wSEf65BLsxTNt0acQBihiZ+jQK2HXnIAEUkX3DBa8SxatamnIbbAYfPvT
oSDryAxlZGJEexU3uoe17RgQFbGd8iCfbdsaYauD65ETJGNQH6WLtuUEsEq9Z26v
VDxpnzDW/DU65uETFbrhv4RdZ8+7tahE9Bw5X99ctU+mNOrCeLa7QiGADcDqOHP7
YQCn9MVlvVh2CxnmgGhgiO04eUgIIQbHKsx5ge4m+LZhNYIAGAFRJgIm4jBZyn5B
xP1TsJ4LBVec6XF/UslASg6XJDPm3DjeXS8aAW/OIS1iz2qIsdZHSRC4kU+LaDUx
O45eFdKenBi7q77Q/q8lUMF0mt0GFhkts0RTWj1OiYGs7ihN8xGlr8bWV7llViNN
3JcEQTDwph+HnildBZ4ZTDnlm4McYmgZbH2ay7DXogagi8cTYLPZUhfUuGtBwARl
dVbEQjkB5d2WN9Z5kLlOihLSiQAPE63nOWyWft9LZe5QPClXJiQEdDGYUxUol3++
DcU3BHBBSemwoiAcx4tPDbtSVFWfPTVtVfAJknKFvn4nTuz6hxe1QptuCjbNTFsI
KnfKgPT6ZeNs5xtDZIzeajTeUUUlMuR2Gr5KjIUz/Enf/8T0xcjM0mpma1EiLpnf
LyPXqsJp2vRH1iV1uzuX7xZbafB42y8Mn+T/ZM99sjKkiIQtc2Epdlx0I5E//JVo
Gb7WUWw3XZ4futGVJ/Bd20cqjT2Qj1sZX109YOFSay7gR83q7IMKV7kXOzaNwelP
Phzu3ZP9mCTEgttojVZ9Y9n4EltQyucVxiqtwHoZxxMi7OewW1JfCOzCOfY7EIpb
aZZCQpY6qEGVaUEvuZ4IRMHYKUNX92yLOjJVM9zzqAC8cJCcFpsHjRi1m6mSCfBW
rOLH2FSdpxy+1zwvmiwqP1ivdJJJ0HevVrxHCi3AE4xZsLG3p6BbxLr2/3AkJPiC
XIcUZV7UWDCWqMN+R6uUWNiGL8ZrQtXaBqVFkEL1tvH5DGFn0j0u3ugCFzQNrQTl
d+OfQ84x4DKJVpM0PPFhJRnlX08kMTpCOpsP0smAV31EEK67BixmV7IzdS7bMPJt
SiEA0/+TKM0fBveg6fmPIHa9DGNP+59dohQX7HCBIWFb6mHRdoOJxT2Ht38dtoIK
VrvlR342RJEgpz2gj4gt6Knk0yjjtr40u+yBz8N9A2pICnkep0KoBohPHaKs5qcv
tb5TOw2NQrRBjDB4bCe+jkFFR3TEa+eVbv6kItHDfSNu7yCedxE5DnZ5VGqB6kBb
M+KQCHtGnSXTQPOncIuv2Sb51JLq2ud9K0A+flELYBoCHjXaDaYiPmu50FCRWa4h
03xTuF5ZtQkDlLoOISWeCbCnOkAcX3svfwuADxROmvyYhJ0uEdTCjvBv/HxnpbbZ
MhVm8kIbSlbccDmjZ0MhBYF0VsY9P4sE66ARakW52DA2mSrvJ4iWveX9wfQ1Ulz2
Yaj9DUngwhcnFmGiz4CyhxNKyE/0Smtk36I+It0rwciuY+q4wzv52K0PZRg5+KDR
Gl2sacx4XYNAtI57mdQdRkCc/y9DgyF2L+YU4OuGKKDZHQOxUNhrl0W/B/bnvnlo
VXFb1ySMbNIdMRCmmH0Zegpudbm8WUkuJWHmlBEWvvNhLnD6jfDcaOnYheFY7Jjo
ivf/4j8wjypSMQbMd/yKf0/EEz/mNhTu2h52VD35v2sqx/etZy+aoBjGMF1v/qoS
96oPzm4e3exnX16mLj3yUJ7LdO15sHYXoO+HgvQRqMj3wS7hsNbzMprnEc4H1P1w
yiopu7dwJM7bL6mqLBqPK6RmuYYd4yYk00rILLF46l8YvqXA3o68x2+sjHVz64pI
ibxFD+Eed64710HV7tF0DTnAEhjA8zQOmUGpJRzpuSBu5G0jgzVTIoc9pRCtdJUL
oAD6TKrFmn3vmfX90OhRg/12X4o9MURVhKxNElVrZiJ7RhXQSeeQj3EvzfKH3ktw
MSz3aCMmvZVwFW0H62LycDBXMVvyXBbeMnM6nW5FGofgyW6tAxxNttjPYgyAhwiK
Y36hW0R8CN8ZXjkJvE5vihqYRWMjhs3QBic5tFBhuXtutIz0P1QMDqSjfZjxO8lP
4AT9q070PMnJ9ygOeI7vCf5Bv+AH+BNL5FK/I3W0re/9D2w5txWnDB0ka6r5CdGs
cYF++7pVyM1xc+0rN5NfmDOfdsmjWKYnZETNuf57xLQViSTtGQ/ziP4iui3Po96a
dDoxMYNeNU66F9+N4Gg554PV9dxZwxHBuLg7DFXksmA4sSuEo/G9p+g6llrIdSML
G7gT639kzZNJ7NzS322wetzQzVPK8/srDJ/KTVstVEXq7OUOaNUQp+Rvp3gvlahr
71Pq655yyPJoW6Kjg43oBb03Lsr5K6Ty9bQcZz/YcKpiRdsLIme7OBC4UriwOFzW
RRUtYf4sfmewedGiJebxZRy4mEb9pEOUAmlsnbfTbHlCSIVYcrtgJ62sqQmw/n2z
UvI58jB6cbe3xLGVDOR35EbyUK7cDzs29+KtENQ4fjMsA6XLk+sjV2YKwZPPp+cp
7c7Ti//NOa2Pgr3sLh3IdlwjDQLBqj1Srd8DYXspjQGPwM8g2iEbw/QOHIng0pf/
jsoLnpoL5GtziMth7q2fe7w7kvM5sarAcFXKHKlM0VISngggzhWq/tB0p7CsJhEE
RaFzac/PlOsGxVvI5xIdU5pcY3LbfXAtH0Tkw2sC7asjmpA7xBePFUps9GsxLasw
cyw4U3GOiizmiVHpsaalwHAR73Mnai9v+nWs1lYKiwlD5sDVTEdvns0RghIH9mnz
QbPG1a6PfKOGXfuEsrDeTPoUfAGZHxG+UeXQVu704BQEIJ6A5+6SxYEjJ3TNT+Q+
igI/JUEeUQDTDVQJHCmVROVl+0X/WoWqt4Gc6MKZW0AyjZrNheGRKiDCws3cRcjz
2eRH9egqfYhUHFgasVs8vmJ5DnYTxKzfIOKASYyw5V8Us5fE9E0fQms0iNlqgm1N
dgHS+UqGu6WeUA5ndzlkjTQ6cwS0QIAxnzRl0j0Ew9bcqaGOE2G+Nf0ssVfbUj24
gPVzKsqn8GYfBOmgLUUUWgooNrm7eLs7KvzDEKr+Qte90IYJK3eDmH4WtllCB+Ew
ShNoI/yIlNFEfJjiMStwzx9pWT+dyMxN3M4Jriy7CLG/O5QzP8SNwVGKsco8aHNk
1pg2790aj5kR/lo02coB7PLFjCJxGbuCYtHGdJxK/IeP4EQDSFBTyTxuORIs7wUs
1/2o9qvpmu2hdVE5ovtlNjmiNSdwbSqFEgcVN5pNrsUzLfYSeRoJUu158pgMz9F2
BVoEBJpnvyefJy++n8g0VOkVtqStAzr2V5eFA4peSD0B2CAIfPWkM5mWE+akAU1X
b5wrvI3ZbTg4zc29ag+CPNZMC7Z/cSfcDSHIUkykWI27KsfkaJ8kX7VgwvoS2Ho6
DEVf9P9XnrBIgImLSKl/Z39m/i+s8HmPSYAAnmg73chhW9n9z6R1Ua/aogGbmdBx
o0pku13ZqqAfn5qBa9o2zKJgLaVrDJkUhXxiV8tXm4ltrO/bXny/PzIvfJcKM0Cq
IB9W7+XE5LZegycSXK1RX51zHm0oGvGWNUTFnMAtDGkAA4a7ZEdjf5+JBKDLVU96
62aU2RXZs4TxdhxPpqQEUAFeNHXikvRfkUYjyJ2E+JwnYugRp3XLMur9YH68bH7X
Gjv5SwLyQumVKdB96gus5AYUVEX6HZAM+9r/XHmCw5BhjQIWuR/ZHUVMUzJKNfMJ
he+dnosT0ZPtznBg6WvM2gMbENV1eK+1cKuWaraZ5RWTQ6tQWzmQ/HnwF8ePXO5t
48gFNDlc8dGX7bKL/fl1hfipPTdc/4nqVquYwGd/YJT97bMDLJd3oT0aScY/WRzr
j3tj8/20iCjTia68MtFqA0NLXa8Je+By7Fuw5emR27zUjdNzcm5meuztY74YN4RY
FX0BQedoTqNNAaJ5jQsDRPeR8qzheXhssKoj/ttAWukveseS4nNPhyvruu2/ND4u
ZtqA1uQ9HH+bmp4pCMCsBPucnmZkB0WXrAJjvOPj4GugavCCELnyjrxfGG3hGhyf
6BpFY6Z9Qq2/aqBcFZ6jlKcaLSwuIwunaXhlGk9inDnNC3Le0tNNveGpDhYS2AZX
NcdZCW55ScxLv2of7BE2iGIZu00x9U4LjqZlHOKlNQroiXm8KsDFy8GFI+QmXJUr
e020+QhcAZC72RLCJa+uV4ZCY1pcwqQogwFgW4eeU/4iJo1IuQ0msPTtIyJayWTv
Pejh6oBdtbejVSOsLiCId2dJuNFjVh5jLdjZ1MgdzNBkUF+l+y8Sy9IFzOd/wxng
Jq+0tGj/G4hygCwJ2l8Vd0g3honouQlb3oXfZhFOReEfLFtlg6wSPgDr6d7+vTBj
pFuMmXdr67KTtPNQZ6LB4QcBoH5J9LkXLrfejKaq6ex9bKPaL/pOblVFevGobO08
Ujo4eAy9zrevLlEKovOO+qSmeVs6sIAgritlRiPBbnRRHxoD1VbkEZwktCSTuGm0
tuEfnGEr6TzXZsr62p0r3xuuATVZX9WbDb9pRevJ7zPlIAeouXrOBxQlY0dZ+YAL
amjvz6tAmBDmvEXFY4cPV4dSW548xucAS6JF/u+vbu2RV6iJ25Zr6R/dZBHMtzij
EBHHkLjBMvAyfOXVoZASsPhaL4mRjuQihpMTEnDaLHkIj9ULt8zoNuVKw258pfew
zjMAsGE1bQDxjS6u67mHR3HtKKp2zfVOrtGx7atG9XPqje5xDuM58UqNwKS/8HfN
jNTmIDQLZqcue6pIxOmhR60rtmoRDJfSnpdQWZ/AGHxXBOOtdLJIaHDJHYi8oPQh
NTI7MvEZ462FhOTb2YtIYb0qiG7QreWTGIvIM9rK6vhAmQo3o9i31P5hUcXwpRQ7
CKXkqaipEUhmEDnKqEG1k6NreLnq+YD0JlVsdQVyVbaaxhMt9tec0hBxGjLoKlhc
P6R8SD8ph2EqS1gzgYaVgwOdFhmEj5tfFwBRxmvTn4j/xlGvCgnArC/PV8/cEQCq
CXU6wElHzQb0J0bft0dEv6+iBoRmd5jb4d0YnDejhHr9f6fp+fW03yPImKzS8L3T
BRB8sEsu8Ew6mC/i6KAbR7hHt3HM7/O4IlAV2DDicfXsk4rVjTgNHIFDeRRi7Oqu
wweUUF6JEKZ28fO0GrGIclo9N+RIMATfNolvp8v8IoY2Nwdxb+sIz4GZsg2j2bQH
hZPjD+OXX9KetpAau2rgBIvie98H2k3BmvwMjBPbTqQsTdgh1H2u7WledrP+KLC8
bYrDS5DBfHLd8dKtOUmJBdsvgV6jSAYczL1ZXivaqQOi1Ipu5S2vjk3FXpT8nvC2
4cWU8EHjRsrwQ5OQgyabFqBKoFRBGUFAoxX5zOOfzm/JQ93kTslSS6QRCjyf5NJq
BMq4fA+ZezivwTKorHa5pxsr2XB/kGBa7EEc25f03LNO727OAZLSnA41FHKPqQkP
Tqdooqw+Vv8peyDcAf+OCYlv0fRAd2jDakfm96c7lURCBz4TpIBoKf8TDoY5zEO4
sQxUdZNo81Te8wVWr+UYj8OodMXgxFu5YKLd/Zqz4iDPW0IEOnfJYeDHAGkszQEF
pg/hMbGpCnCdZToI2i3ri4Vb1W3FsThT/XWk56PyuKypsNcjF1gyRitq026D+Xdy
myGFae+Qxturg9eYOF2rTUHVR+swZJUNAr3nw6EY9wJra16nDQFtyNJFz/ziyvfh
86GXLW5ex9UyLv1fZ8f7rYa41//3CgOie1LlwPepqh43tAZINrSOkTducVGqoysG
Q423OGGyiF7k7156meLRVFhtAUDsf7+YcIqbWAMuIA/uGUI66oI6VzpLR5QDgO1D
jeYrFk53AviHtflADGygmnFFEUqClUTLFwN0yNdmxjORaupizF2g4twSHgigkAPh
eAnhygAcy++uwHWILD99eqZlVJwMB4H3nBe1AXfEFffskVNQjki0HjTdn/fW5MU5
U0xGd4GGkoNFs9ynvPWdoitZZXnaRMnb6MbQM77NLsf3jXe73SozekcecAhCafHL
NHwnvy5OrBUuFzKuBSY7rFsKw9eB4aN0CibGV2Jj9XAv0m//4FmO0fOuoLkB9wle
7kkYnOl9bKEMte3W+gN/pwymWRant+qEe/Fr/J0dkUkXJkO5EQsAeoR1KDt+cOZ7
uvQRlciEF+xNxa+R05Nlg/IKek5FQL/6n91bgTTxscyXfJTC0JyTFwJyg7X9UDQ7
tXy/UQSMYIfqOPlnauhuV1BizxXdY8O5Xj9ywzrCNjs6f6G6LyfnKTSjwiB4bD6M
h95iIs/PRk8/FORoqE3Gmm0Muto/41SzQxtEreoRwNx7CESPYA2s4vvsqeC51z2W
cT9iaxIhxlDSrdZ8TY1I/LqxKBXX9LSMx5w6Z1qt4aAA1ME+i9ZReWpPzAxQPPVY
/lTEx7g2yXKV/3BV/qlxw+FjpixMwPfDyc3xpu6fj/BiQ8+jN29PnpTupet1PKKb
bSQafQbNrymvBqHBvSv62y0+cYWl38m38EVcYwOSgN0or7tW7S9G1N55dOO2RDng
PpTcg9e2odSuGYGi1OBTy/VRirz5KL130NMkeQcI4XjEg88nx1t9VRR39al25JIO
Q8svP2Lvwek4VgN6B+A3JfJ57a5MjA8NxVrwbQALOsu6+FTu8TZVyrNLyUDRnKaI
0q+IrmkUKdePR65cQy0yYUYY9dtaamNZarZwbPsfpcJtL14PZeZ/EGk6yk3YeMEr
kff4bfaDiUd873qSCWMqJViqJAwPgI4HcStopAWDMplr/RxFqKZu0icZ/a5p/8cG
F61BwQoBRGW8YQ4iew/lc90Are5iFaGz+tkLo3h2IFI7xjJfMkfyZKSajE1UsGZC
4qAdHAonh4eQ10em5Lq09AAHj4Jk6ODIfXGxJmsHwjxeP0sh1/CX60HviL0K4Uoh
JcKWm52w+SV1nshLWfCE2ZjV3NoP0gCzj6gCdKD1ODyAMsyakEyO6z3UL4jUzW4Z
fjcN3d84Yd7vKbIpFQt0KJunMCRU2nesmAkLkLyhGs0EghMtTST8XQtT/6gcUrev
5if8nP57L1zk8oGJzKAr5hIRHzgr1y7jBtH+w9RwO/TiB3rcrTDL6YsnrtLZ44iq
Mqria/sXrR1lwvRNZJvwiqmN0c3Nm5OlLVneme3H+jAKkP03QdfGCzBqZyGMauRY
C8qziFOihJoALORm28GlVeur9pOswrw3JKYl6ogQL4nO6bm6cIUo0pvf0Z1esa65
tEdBBL8HdeYjc/Y7NUHmFPzOHtsLek9eabogUhkZ/BrhgumnLAmICgYBtq52i3wm
8XVpXp4qgqFR0ck23IU+Py7EYltkChw8WPDwInCopM8BLATm7KomyF8QEeKcNKdL
6zjVCk1MuR1TYf90uKUCLAU1WNAv8RfZ0UhUx88h4Lhkf+P5Z8ffw3ESh/7wn/kW
4U1RuHSyCRgTpgiwWYzDwGXbshTXJNR2iCMqVDh5icPpHcIJaqTDVdJmU/q2MNw4
2SlVN1U5s38u7E552GZxvjqqDOPzUoom9U4BFKRiyMBjhNXn5xwYE/3PdVhpSOCd
7iZe/0xay3VRbyXGGK3a8XuF5pxGA3NYSOpLSm7QOoVUaavt8Cd1nI+8V1O22/if
Y6dIe22QTj6Dfm/wAtYWSKLeqBdlQbQqb+KnD7nEWNsalEKMdFMH93lRoPuwdWr8
4JLVOkq1zcNSoHNmpCxYtiw7oaFPpKDxqrbydFK6GRDsQJZ/coX8Ep0dWmtipekd
BVuWvrhHI6nm4xJYz02Nu8bOKIw7nbadb24N3rLPCA2eWAbU/iklwiEX6JUu7jhw
Bsy1/GLEFvgqlWDUP746EjdSKarHmclvQALqmVmZ8uKVuXmovs5kvCCxkQ1K7Qap
gtSyyQo5+hpdQUbVwWKN5/OSdcf8iY2B9IEkJ5sYMWQDz/ftqKgUlPlf6YvIqhiB
YEoMGywPC5VflbNqMeoxbFv5dmC0CYrXKTAkHPz3zHTaKpDNroKWhrdhBcfLq2m/
Gd9b0uWXjCh20yeh59Xm3QEKCd2bSOvTCylfsgYqintVXYy+VKDd5rs9cA6KtG4X
3IivTU2PV9XjF+/EaNcPk+/hn3Qfs+hOHbwxLI51HaG4i0cyIG0aLnpWq+lFwjGG
Nbf1jCAYQVHK/FJA2jqI/I5JsIYJ5W3l++TG1M/QoKKp32BChOJ8oPPkFGVZdhDg
LBm5mWlKjX+G1iTF0WGwi/hhvremF81sUTfj5tUBNqLagRbgiP0CIeboNQz+UiTt
S41gEOUv3SWYeuvn+6u8NRCRQoqJ4OJglGz08rs6VInNO0KBrizprSebPtdWPEyp
dJQrFFAiTkpeyuPYGYWzJdoTon7LyG4+RBhDgmof5/U3gBhQojS5liXBT1NecEly
8amJYxzmmOWWkHr0gAGL9+B5KV/rYzt6VK0Di23VAOLRyRzv2MFdi92CwWSDCS4l
G/DJGf5npV7pFxBCLHG/TD5Ch/FUZ7a2pyj0zlXIBj1kzSCuDW5jw+pzuN+tu/yq
au3xhK7B5KQRHgDj9SSbPdTaz9L/KTwF1UgxVlJVHzeBKlTvZFFSTJ8JlexTFOUG
drGO4RVJQH488B4AZSc8rRDir0xRMUEOIQ4g2mDtmxy6pKMl2AXoXfh3xgrCGR1O
nr7K8jR2PjWaEEd6h/9O5bYm8Tg3R385FF3RDAgJlxXfZJy+45pMwHxNqi/R8pkU
9+PxXyytdajcXbdbWwOCA0F0EbKRBZp5Lm+8UphhRIL3IYZxYDpKjvDlXeVsfP0J
H0GbBW6DDgkDtb0kGhvrxLHGfBDw/FmVb80b3tYvyUZDJUpcyE/tFTrxdqdYSEw7
d8Yos4bzNbsht0Ih7ksfFCe0jpO2USDGEkrsDhlX5MEHlUvYDOqTIJVIAz3HqJYJ
3qDfHqlRONweQYsjfWhe8SEAYOOIp7zi6sAHoz7HLHRrJEWzTkXnemvoUcyCeIau
YfCsNVramA2KuJ9uoryf3BvaflbJ/AWPASO6kGafw57byQUcrlVy0DpMKhNakIhl
lQKHgT5ilvPuzaUw4l+d9Vcr1gaZA9rDq37unryCf6mniIPHLyY6rUeof6yE3yRO
T+/wiQYd+8cSqOEbJrixrzVmEnIGPrCphJptNBfifhCqg3tHgkCjesOdY4n7g6wU
wq4e0ueD2wc2aIZvZW0UjcVXQvdKsLTxyR36yUvMvuerIGYfbqVcSHKfXJMNuqOz
Q4mi9lAO6uWD0K0UPD3aKudh8QrixCf6TlLMxiztENP8ce3eWNUpWHWftcBeXu0F
D20gZh5l5iZ5Ifkbqcm44udBoXBm3sSr0oGasIcspl51Ie7d27HoPUUGhmocE4sG
OZpG3OJ0DCjfcYQA7Q9diiFbVA5PpgciFlICgqBXB7KscOsi58Wkyl5Slv092dPi
6KVHP2p0Q1N+BHZcuYVZdaDUQVpb/aGIqxgE8xTo0/U+PF6Qgs+xx6gromk6kzas
0QkCzfdhcdbWox2jaab7iml85Cmfq1c6+hn4YjnmN3ZaFWSjKB2STndM9E7i05YY
c+sTJWfj0+SmvKrWF5hXPIjN0daCEo7T8zyA7AQa5aIMKr/4z2bIIJhyPupFFW/y
fI9YlDjXen1t6RTZlcRKpUnolf/Rm/J+WZOwi+i8h0sEZh97GZyN+7bEYdJdgeks
9pRfBmEmYmkezgg8txcFN6i2zt6ErIxmSi6NFfxkMqcHKBRy0FLUDSL4N4owy0DN
zdth9Aqi+whcAcrbkk6eV2FboFXEuuDE6VIc9ltyhoid37J71nUpZ4//9XMjIIKU
7+X948O9lg2uTtxTA62PoZtqFNFdLnsdjsg8JfrMSLsgEKZkd+dGulUtKQhRDdA1
hKb6f4TUWRYj6UhUGHZ+5vEZub66ZX962WC1srwaOVph+CGwM5Ln8jXfvUg9Fikq
xcgS3ndDuWJSB6hceSwp4Ct/MtPu/4jPdi9VXfL0HG/bQgsqkfkvK2h4ggmr1YWz
UB6HqGePpO21wivW/FS3F1y7hAESxwR3Ei+aTF1j97QxnvK/IZ/xdjayxQUn2lUG
9YfWNYZvXoOBMETE+jPYnjmZ6eIjzwjW5eFr6PrPF+j/Y2bGfTi12UVwq2eTp3lt
3/4PblAOOhgdzuXWq/SuluiuOSuNNcYbgShLkZ2qrbctBedcyt8ZADMQuea0JjdI
p02j7BQ3kUmvBsa3yNhoNchw35vbcZB9zcGK4d5oQrx7xJ5oKokOnN2hQoG7yEWG
ziEbaiEpE0cuQQIz/Xzk2Hhdnfqqt8g+Ul5F6MNrduYvQzhCRfCdGMCPj5KnZnk7
ILQbcc63kVj2V2L5mpqtQ3LgruI+ZNlnZK7+ryQbrOl7+OPncrJ3A4y9l1vry9bm
UNvMEtAfje2bSE4U3B37l1RwXc0VR59ItMH41uEIOmeOnPdvQ8EanN0biw3TLKxL
G2P4dBBaZQWP99MF785gcr13k/TN8tO04jkQSSvQeHJX3YFeHiUIrWu0ziFcaTC4
dD1wyoLcT0TWH6daf0dDWCGa55PZSn9pBP+JAMxkWEUuDgZcCOPdGjL/borjDYBI
Jhh9AANsMYS4wFyEq0rXKkC7jJMp3i+bgshzWwhk+h1kP9z1yPv5apRFYn1BOn7h
xdrNM3+KX/1fj/CpX/cxz2MYNMOFVhL5qe6qp0subtZKHbdBJLnB7egcg6+3LosI
/l7hWGkKclHcAKPJ4aqUj3JXoXImVDfPMZFmcE9s4i2iRY188YKLJNmhMKokHmTI
3xDfjkwqazK6j/4xIj+cBTmLC8QTflQbMg9Gz6vCPtCijyqchB2orIMBea9ZDbH0
VXE1KzvQoM+vxHRSZcS9fZPXKn3bMhYsB0w1XG+WDEkXZFUrZxCckqtCjnA28v4m
9/M+j6NKR2ARuUbbjmepVPxxrIbvmT4+cr6nOrFrJX4k2NGisQ7X4Z9xVr/Sk13o
F/a5+FyzXh0XQuKh4S5PCHphynbnP2nX8WLMKhySLsVbMhMC9aaaDmxD3zcUdRv1
9935bjhsqW4QVxK++BORKArkE9zH6CGQbXkDeD5fRPV+3SPeC7rVEllYX5NHnX2o
thTyY0R7q8i6qrSz+tlJWNR+wzNNWXB1zUMn+6cf2mmzmNQsoJhWHJaJzn3MkwQL
L2qnrgBC2+oAykOf2gZjtqKH4i7v/xII4Z/L49UvaQIcYcBLGLArcdQIiJWkqngF
McARcqIDofzsiQnbNgnzfApt1hgkcwBcMeLu9cieF4EPMp+DfgYwcjpX7guBNA/5
DplkdsIqnoahw29fBMERZQSnVVNAtVIqtMqntUl4jTyvBJ8v3Q+CgIIB0aatpPgz
W8SVfpJkWmorgSa/RY+yRyOjXdOU3UZVfn4lWE6lwjgsH7J25ew+u/1nMA1syTDK
s1SZ0QdbMezfOk+gZaaLR4jnFkFpfICEJCsHu+4Xf05utIJFHv+9wb9AtljEy5sc
tK6LagDE7gFA/MkSurvTIENkaGY9FP/JaogrjGmY7p38nN48T+jednkJhlXHGUq+
VrN3oeeEA6hu0QVyVBkQU3MhLVAlt6Isn7PdyXcrLk/LPviL+Q5lwarPICIwJesl
4fMSrWhRJyfrg2W0PXtPux6+Ho26rWJNKzFQGYtXPdV33yvlUKZI/jeh/7RRsvjY
FiwjjPYh+iRcGMlLn8lipBebrWK0k0wv3AN1jgsdBEKpRU2Avy85mt8TQ7GWATk2
cT0jRteZRVY0JiJ0chcy6FX6gBHEoEkNVYwr1OGlUhBnuyDQQHkiXEkqv3892v1y
ULADoUd8JGWJNkaX3c8XOMVC7/cSArWMoBZk53YjZntBF3UeQCIo/hrvf3hfA0No
f7Ylj5ZSW6JroCI1OHdg9s4jG6z/lSUpvStaTVwQCyXMnV0p93Mjyzovz/myQTO0
B8zKyQgDfWSSHEZ9Yq2fRVn/ZyVBusGzPXeYrd3whpq2ERRATRHsP3+Ti3OaIjAZ
5HrzlxKxYSPFloWUdxc41ExlFntS+BSQhCx6psq/Sb32OR1EIHhvSUSqsVKnjySS
MsW6u4sAoElJBgP7aE5yqLzOjsldSai8999RUB5AeISlSYeoPMds+n0DgcqfBlNV
Bz896r3h/IedsGfB5UtyuYmDq1NvvuNSKJ4fuBd5eyfASZtGZrzMW700wiVE/UQi
zESs9c7Q0QnCOdbqrjJIM4DmnEf6icK2iXfw/jTIZbnrwGVtQ1D3+Gk/d1zA+Rnl
fzG+ZvJqdrPt9zEx9uQyuk1kXQrRbxZb5AFh7FpgeFWnwnZQGDRi/wGlCqGxMuTU
jTVUS7UH7DppmeEghZ5D2jKt2oNThZ1xSAGCUn2A9STAk8tLTtP6miGcRtek/DAt
n8sjaUDs9YFSCWk2JQnJRCH5Zn7WaEs/LnriE2kiNkfaVofE0CzowbltVeqjXzPm
MSBkkT15w0e7LOv6rneJw1NVZMlq5yxe/ZueW30tn4xPyogB5Krhza6fZXkbAFhi
mkKkgLnHM98dUoBEvS0aYf1/ZmfEBMiFM9UKC7isbroBzzepcXWuH08FHROJZ1fh
OItwD/JBXo1OLHzR+v5KGqhaLpG8aXOpXNWOIaqprsdZYjrk1hJa5M+CGhok5BMK
Ka5oUAKcr4skyia+FBeHPzrR4jq4+ayg1USOOckqM6CVq8Bn5NEYJTruUIxk8PBw
dr9JUlqR+PyecUG31B3uxpOFd+EnBNyaEWtKUOdPRpjUYUnfe2SGJHuk2SIypK1Z
REMPcUMYdijRL7M9s4GEfoNigOAPEk9353CBHXB95Pzdd0VRjpQJ7yajQyvfjgqD
wzsccYrqJyOELs+vrMfKFaq8gCXd57VezWJJOfvqd5IQtsrarH1Cg/eFn6LBc1Zg
CF+0RDyd4kDAl1bB+Afvj4BPLcYherGXI1no/cF/u7uRS1wJvc57s/PKaHo89cm1
vBOYhNAI1ADrlCZL0RWH9tlUPZiozg2+2VwC4JmmxlvE595pTFqWufMOSn/9TmPn
+yLb4zowz+lWlPAz3iLeVy+4wooJGkPudFDYltzD/xsRVrUqreh8D2RS9IXQKyDB
tM1kZdod32pypkDLDd3lZc+n7DRhqmS5SkDTpxHB0t2pkUSg03zTGKWtkZ3FsYJ2
qrkoRVjAe9iWbAHefm0tNHJEMw6CHSmTx3Sou52Kc3uDEg9Io/Eul5KcHLqXEuU1
vW7DPHmbQlkxnxnufjRJeShz4nmY6R4pdKtwyxzsoPABasZZ1a2VWs8zAyqKGvq3
MnqO4VIhEFplmJiTrGjx0O4V+vPd7e4L83Qbi8dVrvP+yXEV95JwIkQGFqsg35tC
sLwutnUnM1VLVfkE0THL5Y+aSoeOKULkR39MhPbYB8tjX/PKNvhaQHJsuTYeE2p1
6SXKV+YZ5hFos+6YPltjycR9SXnX4XpBuGhKl6OhDvOw+unuuEmt5HTdtM3DRY5A
fy7+nc8UdW9OmEcSYFWOM0I4NVU7msW9gVLwlnN+v/wZNHMY1qVyZtZ/hxtOijPy
OtMXPpbUDBMCYSUS39OY1JQImb3u/RLBiufS648Zq1Zghx6N/pIvQ/bAVdhJAcTo
SpLAbhlLZXMGb8hyc8VNgj1LiAEMqSP611P90g4B/XkRnzGLXU/U8/eqklZaIviX
qiQyke9RnUmn/2bpKhBjrNBrCKoaLS+STzEswf9YLPZurAFVY0h74Pfe3r+Dzhcw
rLS5Tl0OVhTTXheUoSBXSuL1JuN6evugrauZ0pA/5sU7dmZJHfi9RZkeN/2srwLl
hH5aNeT2wmi9mb2kQPooIO3CU1amiWAuoV2PGLYL5xnQp7J7mh/nq31m+0GdmEhf
POkOD9N5HQYCE8UEI0BnuKy3RhewZeDISXXS/Ht44NRYocLDFhfyIGZfl25xUQtA
z0UiZcjUTEOWbm84q2R12IfptddZUQ5ifrOzrQ84d8UoVSzgnR/B6SIRIfXgrRgs
mVDsTeu4GqHWnnvC4V3etcff+30queDgjDqY6Afda3hZJSRqzIGByS5MPBXOtOKM
wU/+VkE//twDRGyg6Gh4EAC0AQftTbIdLPjlVQdnj4yaxUeyCHMwu/Og8L0n/msa
RM/BMooajdbGTjbAerlrvjNtJSrQbiW/JKLQbGxZrr6lWrQOZxcnosZ5q98/VpQu
Cd1dphIcDROXXbGoW+pO4yycGptnCweyHCikdzI0KoBuqW3UIbqWCPs7wTTSse54
NIL51jMTWFHMHhh97y1mXzFf1fziJcC7/30zdmV5pvrI7pmaPHM/JAntHHAZKOlk
gsDeKrdp/BOMGidEsN480o0vX3StH/WY7KpVoLiQeWRzikxsf+i+YGSGL1qf2mH/
xNDaxfQ71+zCbb93jYK37tAypj0F+DSnbu0V5Qu8a+S283tTzEmRJJEpRViAAQk8
6XustzYjq8uF8YJt+wEGcx/T7YQBivRNrVokuuciBVDfkPMl/6IMFwqtmEznKp5Y
zz698UBSSpBVQaE/FfFWngeV9g0kJiMLVy65YbzQWPL0pICnDwqckz38hpimPGDa
hkS3AF8B8XckT2OLqGA4J5dvUpUEkXgY0IMAZ3vEg1wQT/n0CQmC1lX6awOLA6M3
Ga8ASVNfatHS9D/nBdjKeesVFsEoHTw8ADH4vEb2z01wLzllcl3lUVDLh7ifYRV/
oeH/4b1rj6zadZ5Fwf66j517dAZkEUISB9nIWqRMYWv3FTPSGje8HlNt3nA7uAjT
j7RgKOiPRT2y8nkOtF5O9jpsK1Zqk+4EYu5xZRaHkhbiZMdmboA8k4JJZJa51zbR
HdctGkYp12Drf6LcvamnVxY5+CV960n4xUM17hf2PBR/dw9UZAE4zXYgVOFY6O2L
I9yU4bKNZCP8Fey8on+3hdiEnUrDHeRIWPQy90EuxK4+7HC9aVX6vup0OC8X6SqW
kt4L6TJBNIR6lWN+5azOS8xtwy1L2WwIGI1CRzDYzpnN2HeYlO2u6+tj8m0rptoZ
0Cz/gjMemB8jujvuO+Bvu3oJzsY818eYt+tLKbahfNpaEPVcjq9Vg7NI7Ca9eZh5
7WfnNAgXqlA5mjEkNNs/dqLy5LvBClmRdhDS0z8xE58S+h8dpLnmeu5sn/q6CpDg
IHlJLB74s0N2FC9vFLJCpV9hteT7XiIwM5ntAtDKOJ6ppcS4me3TRXnDW7/DL5+R
CbZngcfedfsIMwZyajCd31hulMTs+w2OuyVvC8noZNv3mCmGxVVoOk/nSCVefn2A
WyTmZLDEnPGuLOOnmfLVEPh1Qu8ZlqUPFCKABsClivi1dJDyMXcljXdjPlsAkj/N
B74FsTKREJnaBOWaRhjRwnK+H1f76QbrVZsXmKja8do2YEy8ldO7kYEy6CE1yqjW
4N1u0otEs1cmPyXBnpQ7uxrFeGAHDroBlabRoE7tVzJm0YVREgri/ci+K6LAG/Z3
/hiYQgvy/NFGqK6Z60zMYCiO6WN32/Xdm2mQoY7pwzCJYVY0puIZ0JXdQHQJa50m
8RZfPqau8/9hBfnBSH0ocqjjgHgoGYdQFx8ALNw8hGitYVQl1G9sP/7xnm2YM1uL
23Swu+x2U+PSFx+baTt6e+fbwe3djZn3vjf1kD5KgWml6bTd5iL+SRg9CV8s/VP2
AHDEDmGviUQTfKxLeVtIZiE4GT+uBnhsZ1ldC/lHxjSiQ5f7TGuaZZuSl8K83JE1
C2TRy14grqyd7o1GsuhXoHOkYHJ5mDAGK0D3MfRV28U3uiloQ4caTz4dkozRTVAu
C+r7uv4mSygnyTcA5VxWd5EIyoGjslw3Op+5/pp/9aXeedW3Zdz998Ara9TIGEE4
lYm6vPgXUMgdXcOuBOfZULrUj15GOkeQ3rXqjYkaVMsco1lF8oSgt6PWuh+RT+VT
kXpWjbd1ZWwVamYfbTkFPJeF3MQqWMatYXLIjFmuBkSoKEf0pBaLe6R3p/shQhpg
wQOw2CyrC+KbXaXogECd1MgvsrSgARmFypABzraBR2Hxqmq/sQTxoKtMhOxK36IW
ITzjt9ZPhCDqwA69HP9PuSdLPse8kLaV6ish3SQguHrgRYIQPiy7nw7L/vZ4bq1R
VU8kkI+m6j6KMUysqzDzUiH1EkwlMZcoQEKXKtFQoZ+dT/4Fhf+DA04ehefX9MWB
KErUP5NZ3VpaccnklFQeAOeammQlwj375VJV/c0lCpSimBaTGrDz9S5Mg9fH4yyY
J728BOXGJh+741Ln8IU8vwogktkGQeCAZw+8jG3Gdfyi1neGcLytjDm5DXPBtVik
MQHtdzAIpfDpPMq3qi3g+TPbX3XmOTLVcEeGggAJvH2irxtkXziHxGKi4zV+KVRO
V1j7qGeQu2OfhsamK+LwDnMWnTGgoWOEN4avyO4MPj58j11Xn42QG6opZ8sk2y0W
1LkW34RheoIkLd8JdyWdyY85GItFZ5aSy805wISowbJQP0GfS8oWE3SyrK8+0/Wo
XZQET4UP2Fw264IqCeohWAF2e/Wijhgb+2BuS6/7+g3nvJYLzDkIvD3RoSFyqUs1
4rwOKxcLYIkO/CaiILqKicPNFghW6QLnNgff1jZR9XAbBqFjh1vZ9fJYCyZeCO9V
V2o//u2yTc0vzUhjBhxzFEAbBRkuWayD3DqQJ45hlG8jYBknp4c80WNhfEhg8XKc
WFEg/KhftGZBMvRaMnAmEgI76BsZ7eOMeKDWzLStKSHbXonGMXel1Qh6Aimh8TIr
lH+aOOve8rLmxf9c1Ez3PvlAs2bXvWs/nn7g6+Ea0l0Xn4/bM0SXxyqZgpkXY8N8
yid62SA806WL0YTOSdy+lY09feHrNuyH6tvOvgkF+2xOxqkLbtVfET9OPNsrr8WO
zt7niHY3gcZ6EQsbL3cZlLijs6n3MzEgk4gYmku7ZlSVut6afJN7UB4wT5KBRgb+
7I+CHxGB75xM3bptD33z3mwL8tjphBBKewEHAwMUNT1JQCFLOtPq3cavPDyGTaCz
+3H5bmIiL3cwVmL9SFB+lsjvpnFF9JCyt6rM5JLIlcm4ufViAi7VaYM0eBsJCBBg
k4L6UaR6yixq5OSbalwgsAoG2k7ho/QDpyWRduwWmZjocRovmXRrwY+V2OGM4IAf
LwPsSqNx5npgVIBuRCPHYc3twYTEZxN+k76f1azRFeKJ25bHKnqEmfBLEl32lvKJ
9Wbfm9BdXgclFlzIFjc0fTPro55Uegy2/gIvxJedI2NKRtsNpZMlBhA1mNJRzcu3
6FalZsPVZ4/ntiP1nxlHvX2//lYLbcdgunOT3/L3OojOd4jHaZuhepZCdSET749V
k1m/j2vtxG7C511iA4XgXvnKYV6K65e0lQryzU1ZCcZD6bab65L3SQs6WCGuPDf/
VE80j9DzcUQRUcczzt53pPSjs/6tkRIk+Cl256cJ0mdyBAHEjvXl6sbkKyFPpvJp
utlWOzTuJequVRmM7eDePVy45HWB3kX+weYobZ6qAzwkssCiTodAgtVKSXUnXJ2w
JrVfnO7gaE5az5dHqag2tRC8CpPC26ylzS+DbrUBST4HT6r1xy8zMKcS/qXGlfkm
WCCzndrQ37cNMtQkjb/vlVnfPYxakvb429KsHv000qrn/e5kZUGlioyC6amAzQ41
qg+bN6FyeWEiPAbvb139NbpMvpH+zFP/V+nmOl6PtnZ4Nwq/tA7EMYT+GfVXNK1x
nGWuVCmuANR83l3WbyjAdY+XsHsgAomIqeSmigurxsdOD3tbIYcTGIfC99UVWhps
Hx1yKmHMTPhpyUSkY6AbAgAGSYOKa41ZEPkQv1aT9+f86mhSkES844cjas+izlRN
qGu1e6WIb4trBpBQNn7VjN/RFN+PGuHQPWLqsf2HRpJtjbBz7s79wF4wvygtlVMy
FTSlEwnJTuVhwvCUYEw4XIZHk38+vq+s2KK5sC+8zlmg3UqdWYFavqTscKodx5To
XOTHdcd5QhXVaET8cgt4KGDRqBOpx7cxdbYkuECW3FOl7bGMLcbEh0ThF31nFtPX
Uyg2HDeuXxyl588hybLJrZxs3Jm47on0OugA3z5GRA0rXbmnIhXpJQqcr89XhyH1
m3lT+PxZO/LlBWUsf227nQ+Jeyw3Fd9HeGYOPkepUo/5ILsGP9fhDs3kRLl7jj3d
mlOfQT82eTVf1RcpxK+Z4SwiEZjTdIn+DzD3jlAjYCPcoI+cvmoXHmuWxCVqQpdX
exmQhzC9rw4RNyVvP7XdLEZ4Zyyry16RRwANfOQdRaUC6fBM2SoOfzEjBcK5vrxR
0E8nIk9iIKkiLvcT3x2NsRMlRmD549LattOEUOQpsRTN7vXU7MgSA5v/NrpUPaCJ
uNE6thKvrC9N3d8JCCy6BSmmpbTn8DkhJvdOtJZGtiE0/zqQnXLCzfKHiShSs54G
OWGFt+KSHsbVrM6ewpCu0+QKFIavRkJLEvG1uoH5gS5m0mK2RTn7Cu2pgZ7TV//V
g3Mufnkr431fEKx6w5C6/nqgn/UQoGE6NDgd0gUZZ5c4jL4l3VsyTqqOpfOQmIUn
bUuGUBh3cxYFiMC+CT9+Vy0vZSdyXtAqp0mOiVHQh4S+ttLQZyvmnMb0kuN9nxHO
Xwd4kfq49wQYa8jcfXfyuwVeOZB7w3trULpbsY+RJobu+7s5reaaQFx9GWAUwNgJ
PwyBAzwyH59Jopoq7NRURcdbRz9f/GHHKFCgXAqAqgX4TNvCmLvsNIbN0fTBKce2
YqG4KP4UKDnrWtcCk/w40x0VvrIRxPXaeBRsPDBNDwO+xrSa/J+Yy4m5IEtWVHOl
xn/Y2pUuxgkj0SDJ70YQDRgrAeDcj0BGW+Us2HyDAwRasbVV94jAgWoNUf1aOkNr
RZTs0CgM3VanZChkA7jfl2c1BLDhX7JkBF6z57L7WVkx0NCQZnKwdwzltgMZBXRY
QCtrugGIYlJgtDrYvV4aHBZdbdFC8hHhCA0BVH1w7UnEra2oW/7LGt1dvpcpsOkM
igemJc27CgZ2w+mKYgD25z9Yzqp4fABkBF3zDsKWh6u4kXkxUG6ewVc0cUSORL/A
eiK3Ccuew40F33xWONNiiInNdd+XMXjG61pqxrbBKwlSv7PNS4u/sjmc7GFWWKC8
ISo5sbOqMiMswsFbB6LmvmUvEvSzhq0bSEhFJbVibwoxZL6Ky989cobxsnw2YKLK
jq3A4MM7vB91LL5NtGC7FX/LSBjocFQQE7kQz4ZqfTvClRCersV+rm8S4htLglfs
y5pXb8gbKgj0kbjpTX8i+vEBhnXEQkoJV+0wIYloONJAZZ6rEALqHMef8yeZlTTP
nK0SFH6NZregG3xiFJDrIHwgrVYzIyg4pPwZCqxN82UGJAapKq+A2nevmiMcu5QF
inO68emEprRWXmw5G+sTxJKT8Z4iKh/JqbgZlfttYAF+hfWGDfPzyvJkkFqrezW9
6EPTa0HsNcKjGnFNhUC/L583RwRY3hpQqcivMT78ifHhhrrsLAhDgYoZu9ypdf/c
26R/Zmn3xn+Dq2GNjIjs882jFGgvI3tKprSwmXfuBYSczqmlcDpc8GHqb1kiRiK8
bNg9igo7ChUzqg1nawMR9eUx8Dhgu/fbDt7f/ufkdFu8BwncajCSCz9ED4NwEk6/
O+1NiLvRn1Zo4/SV+AbLlMmWS+HlSSbiwCHwbDOCaWXC8QE7B2zm29XcYLeqm1Ot
PK7ZBFv/r37Zfmk9aW1QTMOqZBwAKoD+1wNJ1221R/5tNbYN3HGfPQjm2EKfxVV7
QDBJL0DlE7AKcw9N84swr2Lvy/3vf3kae/Dp55ppisUBgydrbR28sRrgb94nOpLc
e3+JV4MJ1hA2R7Z5qWsB4rmb221VYh0Hz6G1Gxos4XsCRwMbS6EcVXSqXkwZ5MuC
W2qKUPkagj/FwpvYJu8lHetcZ5SJjZ9RO2VexbOPhWUOoNzrhrFONvocyUaqbCCE
+kZu7EMrtIFNJUIjPAu5mSKxxGODrniMu3CZBgZM8AmIcJ3TkNh42xuyKJa6gnc2
B4TwfMDsT5LOR3Im03cjYbirLtFyoK0kFUvjkqsHGDb5qXDWq/a5FkeXX0X0Qm3H
cXUyOTCxCAc4wHeBGN9QgPCMND/IS93toKc+IyKR83jRdzZBab3lPLofJITWXb+U
QzQrgvVtz3TuhflWB6UWqx3FJeNuhYvRkzC4lNLpiraXEQ66pSCP/1PJ3J/DYAWu
zPWkac4UXijPMw6DygIoTq9G34O/AGfPwXF+dFFoV1zkHT0EX8dCojzt8Lvtsiu7
UNkjc5HfbfcJyIqWaKx3PZe/D19rWY/5aU4lSr7Kg89xVKyI86QaELTARpcLAc08
S3gJJY6ZCmi1di+YFnsEAU23K8alfOpuMsL2QTutNv0XWWqzIF+5Y1DzHKit/oUr
y0OUgzjnPSkWN8ZP6IGrmwvKm/Z0N/Lt3LcfaPQQjYlH7LGbqwXp3ycYsGfHAFDj
UXT0FqBiV7rgM9z8YdIrtRwu6ibgnoSeI+np2VjzYfHY+1j3zaUx0g+3i94yJPIL
OUT2uPmjKm6K+XfO53pzQPNaH2Ln0ab6YFEmBqqte8xhbectkuKRMHvJsIcbsUJ8
JCBEw5/oCiYH3aYFNQdn8n9KP1JYsme2ZdM3ym9Rn1mzYKsQiE7BGhv4gghtBkat
jV6h12IarDCJnMDNs9YTCfmIpxwKq1f+R4FBFI1mFs/+Xd0xZr2bfWm3Ur2Jyeow
435glNZefMmyskxdTag3lEtiH/iGz+Z1/i3+kAul3NZpVR71ySLvuTRPWblbxVch
Ix2pepPioYi87CSlam1/FpJpa6m3QMUOQbN3dePcxpKYtVVMaiOJNzOvC2xtYlvs
+PyrHl8Qw1RtBOSLi2Ch0ih4HB4TdKoMfWZVcKrj5K1E7p6HTwyuV5yZQb1d5Iqy
s54r2PKlMXC2ovnemiqRJK3zKP05rYLYYBxgCG0v7DX+Ftjq7mJXlAuKhofaDcrf
Jvfs1evpMde2IYxqgiBa7h/Z0yyrJEmH2P2gFy7JQRw97bL+Y3Oh0tQWPVXffWQv
MPDrGi3Fi2DJ5IiSjCrmtbGjdSqmGuTvWcD51ax0WdbWlBTz8yDJnoT3zxbSWxYM
IxYNaSJRpfyoDYRtR15DCleQAjnAMF0/sNtxHq1gQYh+Wl7jClhIEO0LTXLKSYeq
w2LyvR/o7eSKcr8L0KC/+M3QPVFM9iEYJuO7BMcSeHd2h2kqb2Z4fqtAGXBdZ8Ne
IE/vnVsk5LhVDzEO1Q3BeauxPH5oOgnV6JMWP3iZtwixaIOLg/qv2vu6K4UvzIeW
q1O9XKSqqcr6vvxGOnIJ8svumH+kvSo1IljN8JicoyxRSnJDu7x/GxzI9iC/U7f2
MbVTUg6BxPfH35NOMvQFHNBQx9QKN5SttJLkNcqVUoxIgojoAkxV79ZyP9j7YD1E
4yIXu8jJL0lIV45hnf/0dMRW1z5U/zvxfHi91m9GjokYgsM1jn4iH3OSHz4u5nbd
/VnmP5Ps6DFx7IkFSpKYaviiNn0h6HXM72tB00H+fYWyQRBz6HB6El4VBHdIYz6c
rPP9WqB5JL7lccGhwtfUwxDdTlEumDPd4LHttUx3WL8i9Ehz5MkzU0A9z0jlwmFG
EU0FhHvmYj8jbuEp+meh/3zCarMwo57ycY2+r1nyFecB6XdBsXk0tm1aP5bM7JQP
A/r8dJPmjUkJVH2JxEPvz1bZxjk+F3S2qGTOnT6GDZjiyuiA52Zxe0FBvT3lrbb6
olq3Rztb7dZ7HIturo0taMePaNevlcXz+sFLEj5R2mJTB2FSY+qTYcsBlDR4ou5k
dMioTnoClAdWQEHoxGHyw8MtzFC5IZ/naXqQZvEYE6bML5lJpzIeGm+wTSQP484n
MMdnrCP4v3ugC5J0Usgq1J0jLUYbadt14S2A2r5KqA9gzr6E2bzUoeTF6Xrvqt2w
qP5eSKc8uj8V0YQ3PDvioVA40l4vRiUaL6Ob3ZLE380AK+knRNJuO/E3jmgETPVg
w2umNKcVwuD99D76Ou0coAPHPVwsz1w3QKWc8yipcJyb+aLZETKvZo30nezlZq+H
2QIVNV4cdqWscK7tPpH4aAh7RGgJyKeGiB3AF9EpdFcfxSiu82tt8kjlI/wzVmMO
dW2syjqE0yJ4zpin6HBrNdlDj8sYbY4bZD2O0ZbY8p9PIwZ74OlkVPNmx9R+LEoO
om/dV2QnTpWDo/yOxnBVfNufBphZs2DFM+tpeIorX0GHo9giNGea9E/TDGgdpVjt
akW8+HS7brS663YARlY0tmRlKIsjWkczCZfPDVR0iPfv1g/FZL9SVNr5dOhzeUzi
Lsx8bIo0krdVCLEmA4z79BKrhTYrwpNepW6TO+doC3RC9p1LVEE42rZ2+hPD2mfT
oYH5fIpx9PMvVUPzuf3t6UQYsmutPIbp780/kmSjm4ho4CZe9696tUBjJ4KX6sOA
UIHOeq4hDVd7du9KxRfO2jaaPAybOYmvpbk9d35MXJvIZiJ0mAG0xTH2funJNm0Y
jjOqKdbWVQsLALLgdlNKDZ5t/4r0XoZcfuAp8frsQNheP5jbIfcRlAOHREZosnKj
DqM7R5oXY9B+ADDktYqhOKTs6+5Rl+Rh1YQN32jKEI3bEK6tPN+jg7redCizj3G5
9OBIhymctU/lYgAaGLCl4RABtIiJkCOFtHPCJ6rD8Z897pPqSJwPeekH9NsE748B
/fJwbKG1RBzRIZBJ6qv9BHnCMP3+6vKxOr5WcBCSd+q5rTU5+U1iTK7Y2Sw3WD2X
i3V1rZhsHWX149M8/JNEFOzpkfDNKdBW8E+C6yv2lkmTLXYAelxbR1s8HaxVbB9r
yeHXktagos+pDpPwO/dexSXw8DVMHf0rbPIpWCLJWeQvK9GkE0baVioRnklY8IOx
lkSySKdaawigKYekmrB6RqvExM4eBlY6fw2Al+tCLT9P2TvFFycnkRVCv4v67MrN
Ywf/0EU3oBH3A7m+zDUvG2/PQV1Wz0FtoMb4PN9+6mbz/z7WUuA18HryqwINbtQw
xMvOTHmwzaUmr3Mo9VF0uIr8e3651fCllo+g7g8ogtJqUHm/fpD0rwJPsrgHmf6D
FrdVvGjktUCxE2dUcasPVNwwvULU2CpSj6TM1PUrUYuswD8F7kXeuyLpp3Deb0Ng
0QZPm0M/ePV3vhKGrFESOat8aq+whoaA1c7J+mWC9QIfRU9v1I4oi4M28fa3kib3
yjdLMiCC6+YTBdZJL8TngvvesJMS/c3f+Yq9pKpYO0X2mJePAfdOOpU20GrEHgEG
89P3FtmEwSof+3OE/b3c1yphZmb62DLKf2iIki8WpWEPiL0+sIjgzZcnH2mQ+IZE
AI47g0YLm15UqJKqxRIkETD16bYt/3VaHb2VrYbeeqte7ozUzhN4Y01X5EKobyyM
WCmBF4v5MmyVJ8ikWkCSBi3EwwBNCa/Y0JsaKatHJOsYblIMtJQ+CWFV6Mf0uc9t
jyel1qJgaNlcAHk4JDD8KLzCaeq1L65j61qRXy3VS6E3kV7YtcTe31fCu3gXRvJD
FuBGYi1ukgtt9bJrHEAVVEE9eI7LC17kxikJAWHVO0EcMWgcSwLPheUP1W6dsWVP
WSDKGHpRcTcYgd+YiP7wBWMiJDeiDU7sz62/feqkWeltxlkh8WVAuAb4kp/AsMdj
zcADiECVSUbLmCcICQHD9uO6ug8H3XhEKWrRL89NBPtNOK8X7S4yQIxRzgBpYNAg
ci+WcCIOGO366wUghCX6SYutDv/Gk7RTuzQEC4+v3y/0htyWs3H62gErADq4a6+r
pC6tM4wLtwNFMDXr0y4I9EWz7YnJk25DgnvANduOg8s7Ypst1N4FLTQwTOJU8fDX
IMdv+IawUEL/jSFb2EM0ssw5rL03gEsjwLDbSiumkegHspe7gOhqvmac1Dso+y2R
B3eCnbWnSiVreG4FJr9dqF72efVzB1XjBd2ZCO6IP038XHdQMAilWBpLKNJd0IXP
g2y0YlEk+xcs1/lZjkiMQXldC4LQAjwWCo2zVH3GFaYzS4vuMqgujhVni4yMy7P8
yi4GM7ud8WHWLEp8VUxXK/qAiJOuASzBk12r8x44FsSdcx3QRxMSq+Czwcop4+Ie
LcmqLSPrB6Pf5xpD3L/g3/tZBVagUb6u9V/YRTMcGs+F85WORCwyskMF6TqNcaix
Jg7O7yJxu2KvrnyY5q10aqLLCUznpbnffbC1DmWO6ASOb7EF/x3+/ipsEMxRSooH
kIXXnMJmuZE1pt4A3ToNz0LV4JOVTSzh0Rn2b4zOahtQ8PH66yanaUE5ZK4J0WJx
J/Ba+LBro0OkobFTcLCIaBPEYXYUnqab058DsbUZAWR1usxJUd5JpFaxxHzEjdsb
iL/Kfp64Sb/JuSwmbg/BYP9KcM6EVlsVx1YqIvJ8CErpVQ+mgRWhck8NkTceC7op
4kqls5q+JD7C6b24gom2uXtLUmc/W7sAbY+pKDDNPTEs/WQoZHK49EnUE/zKR6Ws
TODjDf8zfhDCJ+wns4rhjpXVCf4D4n2dpU1BJdkM0DzQx3TeKbxM0rqo6scSWmoT
BY+w3/ojTFv78lH559UDOOZyO15Z7D8XMbGIOaFyODPaLN2koo1mftx7ZOG3WC4W
9Quu9v5bUsRMsEVAkr4W9dS5IO8aX+ArMc6qTLpEy9FO2oZb2en2zmf4Rc7EDuy8
wpdqE9JapgKbr7uISGQGKInKW0wHPdwwoepcUPV/cScj2/8WyNBfgCCNiP3l2CSW
sQy0/TeFqPECE0DDGLKyBkY/Py9WCOG+xEIW5GVlwq4iFmXBzJCXlADZlJyKmkHK
UukKIioFM/7B6ic0nYgT1+e0o2AxiXmvnYhDafmYEbVsoYFAYXo8VpCM+32VQhWv
NL7QE6NCu3flZFsTIXmE+R/4RrHIpVMKKH3vADKt3zKH9JDE9i9p0pYNm+h866Jd
UtQSuzyejib/Y2mx9uB+asaHkp/xWk0m+SY2PBQ0qAA5rR0/lVC2Tqs/wxvEhLhC
JRo2ALQwSwwqpsuyjkMfm9R8HIDSETukjevAG08GZtol9q2QeitR/iyL0fJct8VU
dPWXm9YKEOmStI6B1JSkMVowcOi0hqC8i26xD9zML/eizwPoW4PnX/MmSAYk8f6k
P8sJr2KWdutpJ4mogilYIHMHutgyP3TFtDxmNS8BfSk7mszk0goztcIWKxxI+M/L
XHaJyhYpXggpBj6tP2gpuoHHIdCTJTvcCBFwEB0pOMI8FMY7M40qQFuIpOFpSZ70
wo9n6yMw4u4rcrAY9F3NHSKI8KdN81oo/8PWbR1PvvsLn1xXQcISxJHUPFTvxZ+G
iuZ8cKq32gXQnOP84mWcxScRduR8fP8dI9l6g88I/PMGy96Qg9OMfxderqZ/jutv
CetzPTAAfxT7wZhXJWBsER37xoN03dDwPkAMnQ7QCDtLYTXlhtO6mqi1li+H4N/H
8wQ+ni/UxZqPvxcrdVzVOn/GDfIwEKTyGNBew7z52m1ITPN+725VkZeoU11CWBg4
Z6tPiZU17v7yiR6CrMM8vtiqINQyrkD62MP2gRpoLak12Uc8K4h/upUJPhaiCEsC
ttecrD9rWD+JmW8f0uxB6n5zSabCE4GmQxhR208+mjQFvHM1KKdWP8dNDfhgaOGi
EXaxZ6b8SWw1s3kQPNIlZLUWXNRNGywLomQC590/dqmTRUa623ft/PrTPOdBRllR
TKhafMpxbvRFFWxYTxNJx+OESyex67inl2u8SO9MoYQ63ymI7JprfyNXeL0RLalL
WjPcXmwZ5BN5c+oB/KPhBL4+wC/X8mDuXA4xGbddBCl+NDBMPaYLh8DN0qUKNbkX
/2S0kd/CL7BjiGEZhfsw8fTH2/jrYkYfJIGblV3P8I8O1E1fVumsPp1Rd311VRgV
UVxtUIyiROmnEZfB/gyDhxF7s1rj9kU0PwhllER7/8PRnHUJUQnISghrz3+4akpX
6TKWlVOlbAPVamwX6QEFqopfBY3Hbltyh8h999bvIqBsXAkptfyiv3aFP3uyF9AQ
JGKMV8tNsppGRWhEHuUBGnJ0/qLRrMuJ4ePdaUOrasqZjBslD3aZhNXEilS5WDny
HDJyNYAyuDrv0MUy8Xr28m7wefr04fXiE4oIQSBpciQDceHDg+k8fUwDsNDrmNPT
h6N9aUDF90elEPmCmhylLuDuY298cPo+1y54aq6Co2gnaVRlXMerH3TCZhFN5Ak/
izkjTkciHVxI3NztkJVLN/SuXm+57Nt4UTOZunSrvW5h9WR+ikxZlAwmxkZxEzMp
ocZLBdSlDaveUiRSXQsemzC8RypsFn587NYq85EdXythOuAEdAguYokxXo1kqzfl
BHBPf5B0XW1xnlbOHsLoXx1NCqxna0aIjslychDe21xdI75BspFkacHUKLDDQHeL
VKQucwOysXNPccC8CpEHFa9t/ok8XfZWPHs/4d4yrRolcobDqWUiRwi02JQo460r
yxd/PmUYxOPSqdHWZHCa4PRjlyiiLqT85UZ2SEbzBFQ8gFrbJWrYnrmHBibo+oUX
DlcW1pbqIhnoQAMfXMtctfP+XgKZpoWYeim5KzSj16hJu2c37pgSS3ccV/HLsTSy
ilG0gIM75U6zjWgWQJ9ot70idDmOR1LPmoR1uKGhPnjB0+Grt42qwbLVLmoZl+Q/
jVubWodzrrp6ZffqVDAGW27hphQOqE6/gtj2YCxwOozvmgZnj8KQQ1n3wcwpKcvr
Pew8CG0RF7ywqP1pRUmtYV4JeQs2tbVmEZtsvKBliYU7UsA2ydD7JHI9mwtFku0C
NCaFYu3xPFBixzptJqrWEEQs+cbYDwEAaGKL9g/82oTxw8PCM8qsa1B55DJ0FsEB
tFfRnKbvL+EtT0MjlbtIu6QWNdPWxdCyP/sPARM+IiE4RwiAhTIuTSmy41mfxh8r
0CD037MMAi0liINR+skpRht3xtB3QJPHJ+bXj/6Bv8+XTdTuNsfLgbcVoRT+h7Hy
HvhDA5OKDBlAVKqPz/3iLLJ7zGUkmpo8qWyrlNUg+6PDmbP4Z2YnPRpDbrlCKQrD
FLVLPcbQlbD590lR/k4lccGAQtIEKlCdp+i0aWTO2u7weERNqkpZpof1BEdGqg4G
evdp5bkEMELLQSVXF5aTl91HFShXEJyT0myn+NxF56yCCH1EFFghzrlU2ai44w8S
PF0VCEMAnxAPfC4IYeaZjmIJnKi6743iOKUfM6SWQ/w8RW/M54Ia0JqrfeeTkYsE
ug8Q7/noJzLBE4ZF08sMPFyBed7L/5dZG9GpLhufnMU7TAX1tlqe//Ll2AzAWP9K
wK29dVarnJKC+jRhDyhgXJvOf9tKrPAFkboASSxtEdDsk13ycC8C+6xO0jEWlmJ+
u9vsJ39q8iDfVwM/Wnqhg06gxgu1J5vIabtWRJ9P+5faaJJxR48nAnzAF5rEwG9K
anCeRkiG1CZrhJTHns/omhHLQMc94w1bfLKBAGtQpmuUyxdkxtVssuwJIKWcDdhQ
W+R/zdFgSaEWAc9zaJOy4BnSRWUoeVAQOapGtUMha4ftL5q3fleIgrJ6DjiRWMBm
vV8mw496FevUGLrnygqf/oAfJ+4AM0KvqvWCdKYBF2DNzPf/ikUiMoR0IIIevv1c
3HBALX0H/2jv3zqahsDZz3yw/d2OOxe9jUQB3LeDXgcSL2AVmJMbSSV3RIxRLSEV
5j1iIXWorzgxApLBZr6UBn1eXZ9b3lYzJ0obWdJnPUBi+iVbUz2ak2Uc3vgN1YGu
A4WaZpfDbviYNKA6/lSMQmi1hTThnKk6W/IWqHNh1yt5MSNoKmlUjlxGlhsp+yGI
6X1Z+0y3sSe7EihS43mrPGd7wWK5MJ111z3JGVO8qWJ4UkTcwrP1VQssqZdmvA5S
2U49Jg+u2TxaJM8mAj0NRNOShz0vDr+pT5WShXt4CCVu/9ZeqEj6Pnq/QPq7m99x
A2uNtcyXbiiy0VZ9fpzu1nZ/0J0rCLAx3hqouvQN/Fq6DQZ2S+yY6EwvDQksAqfU
TOmGtRHgQEbcTTHltK96dy5X07XX/Y8I6oemURcZn+Ok84c/vNiwEJuNGhw2a+gD
OvJrBfsGdsPYzTby8HqA2KkvO6pPra8NiW2bBv3mQ9irA0MRaSeNYNnzlC1TwkRA
aFtgGxuYi0eVX2AOK8PtHxXErZ9WW1j+RbXKUOQTclhPPl6B/YEsFTLJ4WuAtiXY
fYRyHTOMTIuQx/FsCJt3xrcUcolxwc2x4pRVPhfpPSuYIjp0qFzisLW7RbbuUv74
drh1qnep7S/xoicTBha1Ljpk+P4xUor7LjXLG3IbnZ5ZmDso1FucJrUZcT95/dJ1
B1Ugzks5BlnPGe30/maW9RTEsJuM2sJnRJLAfbQvydPKU7Ym1RoVhjp13PmBOy+I
+pcNSQ1u4HvBrR11eNFxB5EBFLnGpKtIDNXkP+xrq73gvIk3+tnKqworAO/mF0AA
S6S2VyDf6DgWal8A5aGYRTfz+prJ4pKEAOLuFu3di04vdM/fYdovi5kO1tz/ZA8+
iI0Dqi8MfZE+Gn1AO0WrQXZmDekFOggATcNXROg+P39sD9pd+ZODjPMX9F/9Whk5
+8Z2/BXM/CIfg9ZInrntySjk3pC+c1T6u8vHz1jBmoNv7R1VQ64Df9MUsp2oOUBB
smMF1Z15GxhBnWqVBmMwSM0CbI4oaDGqr3u/GkQ8M2/NsL4Xf8The64rxpNgP2TP
MG0ezYQIQHMLOPX8k7K3+Q7/qLLBblCOMe+3MfixCeWhd7baxbeU2UOI1KnJW0lz
b8kr2eoxF5J17WO4DGC6tqDjOury6fTrs2ZSL0S1JzaI7pTo30s9HTtCwkYEu0cY
icyc8YrsF5NbJVSvfqnmQQgtFKXFcDd8i0TsMbmppoxheXFilP7SisnrsmeE5fj2
r4RDrdwkTujUh71CTu6QdjUFGJhtlV8ABMenytGIP3W3uHWiLgcbekAPJ2xYpT6l
k75V4QmRtb7I+TjOt0BnaSzFnCXU9HLA3TyutTjv0aUbsDoTia14iCeXQkh0iptT
b/W7j2YOyEXxPU+++eylJaHqN40PERc2pR32urvxT35QOqHRdaWKg1lDvZXF60DJ
0ADaWdC3cJYl6OnOu6KcrtnOBHbnZo/cZDNx9eN1ccha84dQkNRpMtPth4OOx2ph
fCfAAi/D3IHbivv9WFiWxrT9Ftw+BeY6lMFSE2Gp9cIphUlLGpyLMIk4eiLDzwHJ
EIop95odXD0vMO0FsAldcSSMUQSfWB3Jx1dO7ApsMH8vgR4H0s4lfPNLfEHhT484
r5N4IpVewSr4ViHj3iob8wWXDxlIgoD1h7cvR8zMBBfhqSs2EA+It8+A0H22Iv/9
pVwxHth3UjzEbiDbnuotm3K3ZSVGX2TeSCiKFbnnmxpI9OebLHODNumfneVqmkGE
E1yrfV0OGugcuNLbacIqakEmVyOI0std0NmBH8Ztzrq+23iAQOj09pF8nIUA0w69
HtE/EI5262TonCzP9prhi1KpQAXLpje/716D0LgFKA02N4SdSnp5nWFdTlse2Wrn
lOxlRyDM63nJBTC+eBGG5uWbaM+Ye9U9UdT64cdDqMhqTVdG7phPVpcMBzcBldCH
W64+2GMfrgtsEOdoNkUXABHcZavdoC5DIo+q1+UCd/9lxGsarVVL35UFhKjTrCmG
qHQOUIu6PGPl+GsHWAU77+9besY4qep4Jc5HyOExG9/dx7xxwLRUFllsvUEEeTHI
sRB5FcaB5WDn7mwu4/743Y4L9OlOMqxvlGQWYleBeApPOGYrmub4syCBP24nHNHv
oE+LROateMhmMPRhk8OnD0c6Lhs4x0/2smxPGb0Dw1z1eJUiPL1FrB3QMDZjUnKq
J4OkkJwTcFUuHfdqJWj+++HW0MVE1T97nEkx+cMuKfW7/dZvKqOAAsVuawMDRXIP
2ONeKsPm3MOtlStAyHfMDoEhYhgbmnDKrWWrR/pcX7MRsDbR3xZuusUpbDxJPvzr
w1/9HUEGbloTfxQKSBAD6NEeyLKv9n/C37YZ5E6GwIXOEoULKz5o94LYb2+eMO6R
UxZESqpnkjWgqmr0bB1SSOota/Fh04Nr26Sm5vL2PozN5BTo0vbqnYJJjtD0wlMh
vxdEoFw358zteL9z6efF0bwv9i+00sq0MoqgpKdAV9lmDybJVcfQcAkUCbaaOZHF
dp2YJQM6U+hw2II1OwnuaMygv4aBobjEyX1thXx7HoPt6eBcI/GPGIGuhg8RhFPo
BwFW8GR6CoMNLPzCcTQoA4Cs0yO4y2SqYqctqIr3qk5eCf4m/+/EzWG1MwsIPH5q
nqR8vuHddP4UWQQ4C3C9RfBY+r/Z5LBrxiiKQ0CQaBkEXfEeKENfJGCWeyrUUU9C
QIaSdTvveyXnfYizrJWI0ep6+1S5BRQfXsslQT3cYOrNTbrCg2gWEj51gOFrJ2UH
mIzBQYEhAGN3e0799t9AMzCBhnqnUhI/biH+Q+l6Djc/tGv/57uPK5yP2Nyfj8Si
z48HKQmIA4DcrNTcXjeoH33x+ieKJ9zSI01o4KQqjZuWajMtn6AXoRWM3tc8Vk3s
Y8NGz2uAMoKTB3kXduviK7ACEqIrvG04UGfvOg/x6den0xUB17yCyuAiASSDK9SW
FUCC07htd6ySdA64dSJqJzRP/VwhytozPF1X7hKhlfDLHOn1xlJsqmp2LLgYQVVu
PcOapxS4Hw1Jy1yBeR0JuPz3huN5F/eTezeaSZFiTLuQor10/0++qddtAIqsbwny
ujVjKud4W4q69+t1xJiHkuHdDq12tlNcvEdmGpjTCvmLWCt3olB9Y4mK6Io2VGAT
qHeaE+DTWTcsnIbZLfPYcCIShTQ0VaAyH4C1114Tcy9guSOw1e9h93iIuoJ5vniT
hiX2DTIBCUsjz0upk0uzitpO7vIkl0LlhsdPq28o10hzEhLrT8lRr5kNU9QAm/Cc
aYXqy6fDYzRbau+nRA8LhHk51cdnG+2gxujwBA7UAr+uwfL/T8+Z1dDFAd3R4LBp
FnDOEzuMnjZ3vPRpw8Jw1OYH/1/lf0wCc1ftmssZHSYPoU+htSxqJhO8R4y1Z9ls
o579wOuKlCUEMqbYeoSeoEZrVx5STnRvL4jGjGovQMBU+yJXEB2mqZousiTiOudJ
BD4fYJHdIPEnBnmZ9/lrWeOnTB3BopHPh19fsmpXA+bM/KxYAoLbtmyia17UU7SX
/C7tI67lopSMvVfMvMdA/MJee0OLCZlGOdnjAPkjaut2UTugZ47D0me1Bnjx/OVA
gTiuP+B5Vml1j8gXoWevszQ7MfnukQFx3pSCRn290TZHVtZxAOmR+8X2XQOzspwV
85NqQieG69uIvQVfyKqpSMXb04VDc80NDGC+7BYv9Jm56FXuy4OcKgAhHGTlzdK3
tP6hnEuRQwTVQpdQ99ftiQhHgf0gIG/64yRPM7u1CYJAnGTsMDQNG1YnPfaSuzgL
cS1hRfAMaYEGlCJWTyin0b7BsfKWn6BrboqmbUEYGGzfYNQs8FkfKBquDZmUfzpN
LN+FmAFKndtzwIHETPorL5a/oNi/8652ReQlRneVBbqjGZZoKav475zqZHzbTX+a
10m7BjwF4ynQ5PatwfDXI14xxbVJUefxdFJAQB8XzXSB03HXJlATdiX19X8f25TQ
g/bx/q+6dgZg/Pl/CL31nwBdZYHc/Dj2ghyen1AxNpJIFtQa48r85N7aaEH5FlQ9
6SPkfCQuzu4oRo8dZzWnqzl+DB6U1HHQYPgaev95tRoWtIlhVfMMhEDVJmjvMnd7
NnhE3poQQlB/o00860cFgGQ9jsApWmkkg1fBXPJ5+qAvu6yCdrV9CeQzDR7C0Yrv
i2tJcXgYADM0Q25zsWrYmXTrztAfsDUehRNJ2sUYiDN8q0s51+qmoDVijw+B8GBV
vC/0BzaWr8Ll9RNmh1L9Y3In1FEU7Qo4raZpz8+HWN4aGd2vHyUEdsX5ce9kYUP5
Ghx/UNYpxpAyrv0EwkbQe/rOVnN4KkgftlCdBLttxFhYnxaWaprQXzKzPeRSO/Rr
1C5J5V1ojSIG8h+RkGeObe/xmWPqUG7w9zR8umKAy6wXksWoqok3kHMhMNXzKbKx
zMHpLWEqyGwFHak6cZvrejIP2R1Rd6OXXfjrXhZ3YdUNnWFDEUbdJyGVEBeFuayE
a8yeMzJbt0zDay4M2jKzJ1JJYtNEKq9lgiccYuDmwMC6N9VbvkKTqznezfGQMzcB
7NYcageyPXxFgHnD0z89XW5PiCEAU94F6KxXfappgIJhfzm/cuTJg/nZYTXt6IbL
Ks6CYtR+gBuqFsPBB31bW3OL4CcJOsQsd4BBzZr6MF4B0zvPrialIkgH9x1bVlPq
tgG7VH05/cjWMrTWm2+GQVQceQhXi9nfIXqaBJZwifh5g0F/mL5CKjgj5rbX51XI
SsgA1hsQthidBNR3hHAo5MD3m5tTceuSgi/MjIZN7VAVMhepDx5DI1xtqJZ6PRPA
Z4R3MkKa2olktou7b3nC26LfSD4spoz0NI3QFOhONrtdM+ML90y1aCVpCIdG5G4w
da3E/db+NvKeuBoqeDt84/VmujdnEseRqdjtVuhMERI89j3x3vp+BMXsmwjs9rRM
HTPbot1drhffL1jkqr+hBSCoiQzm0BvCOzfYJ590HvzoKRS7AEDLWJPKYpZW40ty
qwMsLcYZNxFGff+fS/SicpoIZoJSk/V00GH7clmfedPazKrSq8AycQMTYCm4ijlv
Kd3OOtxSRlGFgjKNUk690VIn8cja4KSdNl4bV8eScf8+wm6paHnzEoA88kzQAjox
wQnpI30zcsxwr5SAYwvdmG3OktvfxNu+vpUAM7R499QZwN5mDvqGGwiewccXWFnT
4QuiVRSNvBwTICvyn7TQdHhERT1aTztd9tO0KR+uXgqkBpSxxkNiNHvjb10LUo+e
ri7w7e/8FRppwZDxsbO2MSSK5Tm6KneIsDWuC20CO/e9yx/gPAvLZJ7KalRNkulc
897ZM34oQOTl2ayfha16+ah9DsEMOFUGuc1P5v8u+D9i81rhn2CnOFXaDz5eoDtv
D7khspir/e3WBxaLy3Ebd7TZVi25uHuZ5APZveMdXSgpvX8wvtdw5GrKi1/Gh18P
3zr59mAvwNp9cFMlZZUfewn0WTzqBZvIiGL+Q7YbIFzuij06Q0jaAQ5nYcOriY/g
mBJkRLXWmn8XgcqvDRyyLxaDRIHoVFPP+jteLz4+joGnQ+n2s4C5iXVfyYzfcb7J
xYhd0HcuNSZRtN+fwGC7uoJXIm/IcvtQaPcVbOHf/6WEDbX0Ls2LQUOoMC2wqwrC
wnt1AaE0E7Di+3PVoMMZ2lZuMedp+I/vWkPYsC5s+Id9t662UV1dT4ziqDffYX26
6jaH6XpqGUHV8oizJBbvNyVQfW6VZhbOGYcF2bgMknf6IBwo19BTdu2kCqqnHOVL
1h4hub4b134iaT8iadv7GBKsljfI2kX7WKi+oYpHinVwPJFR4YKU+OWepsz9OBt3
kLJbB6fZ1NniqP9m4VBoTD2ouxH4K6ActcMTN8xAZtG30gAV1ufYE+CeyyEubw/M
8lJsO2+emv7NZflT/k+d6JRrzM3YvLRHLomlGZdVlaNwL56px6s9amvW47Jql4Tq
CQSIaCAhjFdRieAAC4H9+nR5duXWuVPsCnbzLHQGttQS6jqqH3rPzrCRdz52ajvn
QUXxmkl31Z/Mz9f3TpEaOVR/j92UI/t0DhSkm/fslBoAIIdq0VKO2CnEp0qMSq6V
aAVolLADKt39rgqxStuDDSdhu3a5eHgP36lJ5XtEGvx3wXIixp36kOsH6NzCmDHe
cNop0ILyNr8tcTNmrw3EdMMR+imGVJuUqP0zDKUe8wspk4ONvKQkMlzLVZYUFhYm
3fTpA4fzq1D+Vt3w08cYKKrwj4gM5JhtohRv23kdvI23F2Hv4m2iF/Xx+E1z8v/2
EbBBVLupSupXrS4tlNJ162nIzyKqj+nckbuS7Va6Mfre7OPnUMJL0FIsCtivrG5v
T7Hwxqbxdd/894+oZMgaIS2azJhO87XiercvjwO7z1LaoCS2VpJoicr+6vPxzwvH
8ud+hfaZkukUDtEt2q6PFDc2AFBc/Bp1ewFrI3zghDUBrl3+CDEdvLeoG+CdQnfU
3ZLAqgOCbL0RnLYuXxhHpj5Hg880OSPPF34fVSah24RUMDTVauksvqUodL/EwZMc
Pe4IhSzrXTl497A87E/N06X6bbOhnQY9csZpSCEKvAqlwOrVNEq/zVt+7V2aY+Go
RRTQC//ks5/k8RIlmLVO9K0LQhR8eCsn6Zqll2unYGrHj9Xg+w9a/e0Iz5AeBRpZ
mxLqFJkQkPey6kgYv9rx+1SBQtt0uefTQ771kq5YUpME1qJK1URETfrA2YeycWwZ
178OWpLci7cKXRGUH/85/takDSafZL16kKyNqrzGjAgfxLzokKpk/iAmfWPjvx6W
HtIiyJqjan8SHohHoRrmpi4PdgBH081GM2evbx+IVHgAB4nGrAvOhG7NyX2tOyPb
xJ6vCUxsXE+m+weYqMBm8WzncbRw5OGhLCsSnuRqZfimk8O1fkGs+OKIMkEJIpvJ
pxNiDJ0LulwNWnN4CeSNt8B0l450rzvYfxLSkKHWt76Qv5zMu788qGDDWV/OE8k4
DZOxw66E4PkfTpERAzOW2x4C/W0+VixB4CpvKNuEBUCgErgNYEOpUj3GxLuEZbxr
S2NUWRYhC5qf+FevDUbwltBGMchbiUQMiEJv2EvYl0U9zOkvzwgOSZyOQooh+olv
xnoCEA5T2frLYhcOmxuIXVexyEQbStuFVLZ8RpD60GvKse6HwoMPCficdQSscPxL
v8C0zypA5pSu4tjw2vlHY7FIy+iYAqwA0h5cIP0PGzPLA7lo40lbUFu5Afcf2KIo
Ishq4TN/jpD9pRPsCtryX3cetx80WMPVEVXFZgFiL2cX/eCLfRvdCsSlG2zWd/HB
fS/09XDFeKiRiP0hGS6GHpbajYVdf6Maz6es2p15Lob53699e6mO0XBZNNPZ8p/5
31TH8BJCVLdJk456tcI1/M1a5sZAJhEKIeucAnR3ItAGipCSMSPy3Ae3X0Em6ntT
QAaeIAqmreCaUFOLkjOojIRwn2eDV/HXuRyFBzv8v/PNxAawSUffxthqjmNT7EfY
9vPz6nUgXdNOUMor4xakmYHNeKdaLaI8a1IYF+DNAVqiu/TI2zWDPnIofYsg3j3U
GO+IPe0UAJBPilC9okacHbUed0Pnqz9vUCW+LnRfcGlhZ28a31aC9gvYxfLSABi2
BR8u9QZQQUgraZb65uppqDgKZ6YrRRHCYF7luoNygdTpkXGkSEt0JM8QuyomnWuy
yVdHLjZipZ9yvruUBDxY6GjC4BV6EOoJU87liFdXCTKF5tqwibzJX6SmHmoBwo2m
e84fpTm8FcaXkabgxZsAFI0YfLvp9BCYUUPQg+NixVb1fQKdjGFfNrSY022cOqiC
uFFenwNNnUVEloX0BTBSSbY99ze3xWGljoj9hQru/HLBEg51B25kxsLO4+Re84NF
LVp57nr9y7bfJou4FkEJ3G7uUqg0pf2COJxP8i3ErT0ZW+egqCR95jDyp7DEmay6
ufCYJxVMijPFIL8AFayROS+GxNxOqny8BpBz7jDEuVcbfDmURVe6gHLDit+sPDmX
6SbCCU5DbItPlES/YKuMJOFVCVbRAOlfJacqRCzS3PI9nDy92P5Fs/P1kcuF6SM2
9NGIHyAT1eWEO8Ix5WXKjijIETm2MWpTwJPV+d7I80VuynTp6fe2Ju7YtRSYfuhg
wsukWjJUIAbnkeBYg3pZNLvnyxjYNCxS/3cKsxjz35/uf5C2wF3SiKEiw+vCp1O+
tbhWDH9IVHSGJv7N2aFKtDbsjOAdFqTz0jO64j6wWqeDc/ybRJLkunpgZHGa4iCa
EQ+aL5aQUuPpzrYjL+IFCvZJI+PKc/DItFJ9l586sXD3YHlejLe7I0alpc5ycctG
S+8LsejJrEmSji1YgrQOM7SGUH95FUQ/gLHshcRUZULX1m23YcUFu6tlvgzOWqeL
Trqc+6G3N5ID5789Ds9FLC/dwNsWoNRajwDecXxq6s+6HsVUGFXtVSZrZ7xJKtJt
1dEZvREFXoqUPXglAi2dgSus2LUf4iVyE64l6v/E/Y9VaLd6/PhA8e3wAVlRZP10
Xdivr7gvJIovcuj1GRwT6nHNuEsQetjksRrdWRkuU6T/TpMGf/MpJT8XamcdyylG
8ZPMY0ahj+dEMJ/oppSDwSV4zwDHkF4bNUf8KZLXcmD4B3w3aWWdyP0SoZJ3/OLm
f+YhONI8L0/volIsMghgXjwCR9AmeolqK14nYFLD16Kh4o0WpCjZtQGyDIIdzysc
FIOL0IwCyDwdKqNGYTYdefgZGnUGMhgCBObdA8bzFGrQkQUFL+CYf9B17dg3cuQC
vN11EwfCYBVEBT5p9HSKNUxyJXMgUqDYKZbTkfTGZXbqaJT4N2NIs7SbA5lh4cU4
I7NsIKwU/FiQV0p4JD0bpI8mvVXXg5YyMS99WFoskjP0+Iph+CNlAq+yn5f+j789
DVaKzQJQdf/qrH53P7bA6kCbx9Mm1bfv/btjuO3D9Ha0++rmhbE7h8WjiUxkcfOK
6jd6TiHp0WEaezEdsa/th9s9DMBlR2uHEw0hnAFZ4s3G1JzVkANwJFHCc3hZUGnI
APeyl71GCSfUjJYflu2Q7s/LQ/BXggnXQNzj+wnf3TtZK5pZh/he0zxaOoYexNMc
pMek/GQ1JTqL/TnsmsU1RLmQbhZod8B7UwXrYIJsk4UHTj+vwM9oqdOAHRUP8MT9
kKs5WwYwUhupxeH2JC3rqVrgFSnzZfD8rpCA1Qw7e6mVEAd8gGANTY5QV8uO/LfM
XGcdZDFplF31b7K3Ue8h5mZ/dLz0T3ajg7WmW6i/lkkT13301hxP81V43or7yGfp
3zTUAKa7vORRWRC+Ye2fO0nao2a8LkRUCJuXaGFurj9gVy/S45O5MCaBvq3LZHsf
UzObv1oN/zv1wd+g4EsLFqni4KWhyPCBgNScsAQvU6JIq+mYLgni2hW/kSJpoxaf
EU8HAUV29r3bmrmgYdV750K59VLwZVJ+UrokZQE+rtJetljWGOdWp34+NmF5kmCA
oKwYZsJjXkKeYDWK4R+lNeMhG8VjzU2H8oA5cUsqcXxsrXVGPP5IrC1QKJpHW9Bk
1NZUjWyFJJAxvtk0oIC5zAUa1LdAUTorlbqBqz1eHGkZ6tfg8kqbHaEWSLS183py
EohycWfvnMrCWHWDAZKpPsRJzMQzUdX9UImM8JHlkHcHweFLXIsmjBT60HNO/ras
bMYO1g5fXqUnjKCW1cRYYhORaZlXkb0uewMx6n9IJvtQtZf+cvHtAeXYTlzrWgqR
SwStAA/v82OGQE4HfcP+1K/emLJTCo+uPgtVrmpJAEhfHfqWYdIogK3dSUgFzNAN
EhDOH4wBMWdSJkoWMXFaNH3aPVQ+nQyHc2I3429jfaFQTvhvC6GIiJ9ISCjGGXQc
QU0H1mMAlv5KKa+1mkK9rCEbdtd2UL8Sp4p8ADLePAdjMKiEtCQq5gz0LtsZC/A7
X4v3sBGDBI9gBp+psgZzIGc4M8u8WrTWl/xm+uD7DQViq/EtiB0Epu+oD/2CSjmn
KV2oA1XVRA9/ZWZPUFDIPOvr1HtaZ3MpvlwqnmAw1amEKDJa0I1NzlvD+0uT9utv
s3G78fBoUV6ampL8uJXe8qdWid94jTFkdfockpGRIRbUZXTPmI47mU2dNG+NdJ3E
WkvH3HoQmOHQAux/3UPROVbT4iymInfijvkhlsqUXsE3eDxQF2VLGQPmvgHIUoYL
O0cAUw3K8Owuh/C5iBAaVgg1aBqQXch4qPvgYDtJrZYOwnZVCu0cVmiTSd1u06gj
Ew+5eLxkRd5ECS/fN+RWZtp5qVdFU0nYZVYjEgu/WlzWM/Y/4j5nrri1GpI4TP+a
MZJVDFMixXjfyhrFyLBDNdPCnS1xBq3ih07+cadfid85r7cP8DISNrTaOH41ui7v
e5UvP4i34N6noYqiByEKpGo9W1tojBeF6SdRlitdt05OthpDBkG+eml01yiWvqgZ
bndjlhPwaAcpTnmsvFrkovm44l/dXzsMtD9xAgMCOdOPzpIkNluJpOhNuSoF8QCl
vOqrRH9jCA7LM2ACpcSDmDNyhb6wJvD/NsdL99hwJIazjjPTNdL0BHFUPSpY8shy
NG/t1hXuAjFML34u3UQY7dHVQ8qhtIXgGlNGgGdHsfqYxg/J6cZdCx2kuSaf9liD
rkJNKUQ+R5IKvs0Ep8+aIPd1BsjyXB+W+T+VRYlqZxqwSMPaxWRjJbrFPArvs5Qj
oCg7kxfgEqK+CT7TNxdjcwONVjyDmosN2fsIAxqTl0KEnrKQfdp/p76xKNEfKJ6N
RWlL/C3qEFcwNYFlglzVHczpCCcSCn8548UlN7hNyFQGmF6aWQ3QpoPTahVmvEMv
wDQ3ZaYkTuCIKHtwlpFkdAO9pdv0Ukjqo+2I7JfTA5QkNqdITj00Eoa/gMciq5Qv
UEQi3/0sn9fM2GypfoHVEmH9dRM8RQspo1GylE+m/Cua/G4LNla/bvZt+xiuHg/2
gQ068SWMFnf2/Ivj8IPZFAWgzcWNnUlvNfNkfcYljus23+T0MFBxw9jQ1aFFQfg3
NYHs31jPS4Mg4+3kUVIy4xoQmDBtMzhV4SwhVLLfOjUeJhLYy76rVK99JbAuCM0P
LzTDr9qmmYQ2h55e2y7fsJpsjcNsF2daZAANptPbNny1RqRdXwAhN01T0YcV013Y
nzlMUiAi/lUCaQzK5KSFz4AvW7h0Ljxdzmd68Y6tiR9LgcBNJdOcFD9/RJsLwgCV
4cDCVH2eQJnqWoX1T4XSHb0mhaLACX8mAGifvPkgu+j7qo/z7Gd2XryGNPLJ6Tm3
G1AuSvpErsMJdLx2IdQVSw9Q8/15xnlb9pWmiHBfABYt7sXc0izW+zKdZBf4PqFQ
VuyaC7NvCAUGkMp/esNiUQ4m4Y6tCVq0dTOI5VI0NEgUDVTtlIMGCgeIgI5RkMyz
fpsnifYY4hWg6hTz/AVu6DylcmCBG5qYHSJCGbHx4n/8B8dyzCmTbkwllJwbVRpD
EETcpkYy6jFdLNyfNaNtwWyImgJ9bbIwi6WwHdIS6T03siRa/OkChTmK0i+PJ257
QNpIuDlnwL3oVNAsyzzL8lhnngAbjkWiGQaqtkMSDlBRm37Z7PZkEY7MQo3Jho5O
3KrGoSYGeqKted3la7P7lXr6+E8k5LDABfU1Q9JHgU+zIim/FBBn/CHtOGGu65P2
jqTm7saaNd1DiCgV1kXifuwxiZF5E7Ftn5lhqqaTA/xmZ412UHdFHzN4nUDeGzIp
QKMMiPdEAMGUuilfldKIDoJcWpFHyTyvR1Q0imHHw5QpiiHI1LYomXrqFJBHADMW
tAFy8ygDt7oIlMCAoomUA180o25vADsT+qfMg0aZRGAwq1QGFDt5WKzXf1BZlcq4
3ybyKiZzVSPlGYyO4jgv86MZbsQ4jwmLDbhnW5ZI63qM0BTc5m0Pzc9+vynRTwp9
H9Atimx3J9E9FL32mO47RX42GXCuUyUgfq7HVLvV5EQjKE7j/N3oI2PSfBGGC0dZ
IXyztMmGeQuMO6EgFk7UX5NicCFn0yGKUoziE44m8IiODFmRc3v/I+CdpaLJWNCV
AOeRG+Y8RSRSBe2ilm/Ls4b90NFN5k6Ly446RY97hGrCzHOfPLVG9n8ZumfZnurw
652vurVDXD6LM6Tprvmh7P8P+NQR4SSan270z/c0zjEaa3B6dM7qhbEKGBNA8JxO
gpFubXPAzFx3bBUEBVwhL+CduF2VECbqda/JBh/TV3uzDwIfiZ38+Ir4cH/8DkON
cYyIEfdHvTj4c5i7qjr4TqdVxU+DPXFQovT3JboO1trZ9B8YCwTXGYEcdnH96V/G
Of3wK6AiAaggjUHINJq8KqwoE8WDoglV8FKJPLgCyf1Ug2p3M13pjea9fF8Z9DWE
Yk7lPH9+wB6ugVdXicmDvMAJ8yeLJlI3lpj7pDiQMfqrhZuN+iz0J2t8AWeoO+7f
H2U8j4PsUa/HA0ahPFc3z/umOwMl3ubOAVFfuWVgOPgh+3bk7VzWedPWZznCT0h/
09QOBj9vtgnfAMVF3+lxKqSkRGAeoDdagBIWMOJmJ34tAzFVfqiH8/os1V9m1+UG
WpuN9W4JyxXoxVgWjduJHLkP/T3x5sKdtCSQ76AMiKozuhPyHwlUTII2uz5hHT1f
AsRY/chU7UpgCJxFiA96t8B0K8o1JwzJkAOu7Wqrddg0SCEk482YO8sCXCJx1z9Y
ZJ3hFYozh8xCFrz3we2nwygogu1Dv/pV/LsettrpG4oqG0m7geZa8MXABioBRhAH
1HGfdB/NQvZr6nTT85P5zM9s3N9wQWXmVwUjJLzI5VdCVPHLRzllRvWUfEmx1QV2
aHlmYoTNd5HFPOBiWBkbeu2LXNHamq74SHhC3r9xuOjfWS/isp/QujAJ/i7X37Tr
QPph/pRjewx6jxKsLoDnvYe4bWDeUSsiGdcBaIedAabcOWuiDInPqDyrrE0i38Nx
8Cp9euESZYHB8fScSF7X54iFGyyEHhpKnIv2MjYQFTngzzjjYusJtuLWLCebgb4c
X7PU6n3J2WOpgW40tXevX/jANQmXPqhLA4Dhw8VXka9Efu4sNFeTDGMlH/ApmjJT
tssElyhEBeGNDki43XbVJrSlw9t+gtLcllJ0OcvPcKVi60o69NEjs1wrv/ZH3FPu
A6EV5N5vmj75NYVh6Jf5Ds5PoDGGcdpkdO2nd7Als5rSDB5saAlf842s53M1kNZk
Q8kVqvwxvbQvzzrbt3wRRaBf7+q+uXHP1BXc83csiqWQ7LGXfcJxkedjwgjnBFTw
k/NRjKsB6QDmnlL6eR9Tsw9mpQIln1VeGqb/Fc1NdwwK8jhaSP52AVnXn4CXfLZ4
6rEVNOzH8mwn2XE2/fPoQh1PxDeUP/nPUOEoE5u54Di18hZSO2kubEB5pxkOwvA5
/i7f8fxSEATkdrDqQGPuKPHrMdfAZYl2zOxjldqscWz4+VWgSqXrsRBTLruGb3el
eZM3a84aNAxHYvxJzEbe7hHQUCa3aJpw8qCsaIov4hpyDyBa95sF1iQ69OJIHMGI
oHDzff8u7r55OOoCpR+3WiuiN9yf7XH0Q6TetLFYbOasF0eyj4ZBAKhNosv4X179
mlnz7tVQc3KFL8t/hnn8T/E82NQ/xNMK1w+uiAEAzR3asmN2mLeST9vcWlK4vFqv
24kgtQ49nHBCm+LZJGIKYh1/u2IBAxunpAhO/VhLShxmPgwLnS2Dp7W9yOpTnDE0
2e51YLXKPnWu1gRUI4TLMmiNw1xdkdpolZGeuFtgGpsKTau6BqW+8KXsv4RRT2yo
NHh5T6r8zDBM8vBRVMn6HY3z4iHtaKtvVYR6jL8rpjQrnWtTmiX14tiKsCvIVv9Z
oTvtBXGCRCGx/cQl3DfooP/K5O9CYupw6mibEcG28HeUf/wQ5oihEJ5WWXCq1ll2
2/2be0KjrihRCkltx+CvF66k2iU9P0WtxiCIvm7ch8EhMQMDoeQnPFkK+eZwapsB
WYE17S5WXGkJtGx9GC5SZSAhVeA6glfuY2Zzs957WBeeP3zpFG1A3/UaVffB84wY
LiZxSaErQgfS7V3rXdw7HBIl4csZcy0t/6GIJPPkm4HQJDOGHbFB82O0UWW5xnYa
8Cm/l9OOf+ZdpEuzqW8vz+SjoJC7QGQ5q1wpSCbu4rkE7PvYVAVB2xzPpgR+lctv
aew8Wv0IBz0mtN388f8miyH7/VP5NymKOp2ndPPRNU4BUUx/ZNkmb7Ae5eE2tILW
Y+24nCLTFQNPPgaE9Toinh/In7Ubj5X1wZ+5m6D2ipyX2hJ0o+DvggRDIDuYpq3s
1OqvSAW3VjR8Iu0GqUeXHCcK+29/JJFpVycmo54DfxcwP3z+hdjRgkUwXuudSL9O
Vgg5/Ui22oZpHcEy3Xxzh/KcE0sv+PK0A7Qb4GMuJe3Q19nafUK/YClDIKk+VDaO
UcdhfsPY4dJ80rrwTt+PycN6he5E0IqExTtNe1FqjCb/InvEmKqvbKnFF81fVwXH
JFk/WAVdH+OOeLNH8B0ugqmIa6G7XhYH1WStKmyRp/0GxjYhtGVK3Ok4yl8BtFqq
EAyLlb3E1MoWEOeTI+inldTA6a2OhtmDCODJQM+ZsM5139mCE3zkGawetg5wD3iP
mcOuggq+/4AZrVPelcchqjVweu+tv9w7m1gGJn2GtqslF6MAD1YspTgQmbTOT6c8
xWLRynSHFfFHz5XC41TNAfl+nBMT6xRk1cKY24k43RBWbkAj12lumwTIslnn1qNU
hhDn4U/9dADvTG05RRD4TY7DQNBOiJfVQJCQH5kl/asgcA20VGkxpBzyoz4yMNoB
efxtCjTbnVSV8Ib8uYeQiCXob3qPjFAPPoP9rWExzq2Z6Fl48R2P1z5IMOa1U2E4
ZBzs00JSQeDpSRlhMV4qVl8mvSPxo6gmkbUCTu/4/76x+USg6CGzErWb/Vg4rB+x
Qfg5cjqrxhjElzW5dL/QWVQ/Nq6eB5F1s47CuGioCRxH+gSsy8lyp7+8ljqDEeCC
tAYsQusopMY3H9pRmSkDbqtbKBxkbrU6YzTXIo+K+GK9h5gXwLA/6yv8Pl/y+YRY
yutXoVA19vO0Y+HHtQdG4LFCRRzfRFTpU5s7vnFhcVABstJFEvbeDXUCrWRzqIg0
73U6FVIn8gD8sM2IJrhGzhFn81PP1ffcB/kBAKdLeLG0Wf5gnjwYuntqP8D1pLhR
74HIFCqhJSFDAuN/b47hVKEsOo/iF7zv2iGFQTUMhZt/2bEKIYCWQGt2UPXDEhnc
YJ9lXp+dntmWFHSmFGlHClL0qi7m4iiwtFVhLP6IjtBzILL+k7lSDBPNkXWymoBu
fHu1yF2CkwJzm6gEtziccWv6WmifEH5UMqDNXkEckS5He5uiwnpKrUX0hum7jPxU
OqfPZA0Fl6e37id0z12KZSqpmvtaUC4wVhWJFU0pbjkCAOjlzqcScm3AJ3BkIKVC
BNlDGdqofiB5GD8eZSWVGrIlRg3hkUMN/xjm1le/UzftXXeD1ET0SPmw8R42Is9O
MY72Yi8FslT2XVKCX06CvQ79XqwiI921OeBcywTJvSplNGfAFvyszYh5lUXCMcOJ
muyO+HwnXgAElq64MZ38nr6cszEkPR+IYW5N+oa3mtjWULcY73wCSE/MNuWdN2SI
p1w55YgSA4qUM/L61Thqewt4mmlJ1m4dYUd0ANwKtYsdhk4d14I12oUpHO0TLVgo
J1kRpcZWhhmZXdkMQ2UnArkTycqwtkwOzwgWAEk3Q3nnc7NFGOhRifajzg8T19Uw
k378akYRW7GFF9qn2eOuXl8IVfuGOY5XnXGM3K3TiW/0oae/SIJfZfL7+bjP8zf3
5Rwkl1kxgimE+rYhGPRP0BlEBhsVRSJL2d/eRcauo4I3Ommyom8fmrmEeuNFDEF0
UHsQFGkI3Tv7b/vMhU6meSZwF8LX30p1LngCgZ6pGbvRAgiIosPa7rbGB2muBVrs
KywLDH/PjCdwBCx8T+1JiIM9wSCNTrs0szHsLMzpkT9KWDKE4hISHyZZOGgbqFXC
e2dRhAN3iRTKNP2QS0KS7ELmx3RAZg4jMTsQ9RX9/wJzgMFG6xK1H6rD0no/ylsD
aQqbcBU24VyQelKl+z5xkfv9ej5GCt7BvYyZqG5WGC1x4vLYu4Ibq9eHE1yv5mvp
9N4cYhxEHHRYOb76OW9lzXLHo1qICzWs8gFtlpzRyFIqK4ImIs3Ys5BeM23ep6ZS
6mx8Vhda62HUlN75nmOGxZEQA+ShH77KdEnpieRcqH3jQQYeq7WM9xyE905JdOF1
6jQ7ceetBNa/hNrKyAMV3DO/khyaSH22PI69vKEsx4/9i2pKivSiHLkRZKb+krCk
U3HhOUZ6W0QUmdUIZpSZ4v04jvAfWKii13+mo4Q7fZescsHCsgVSmqxjpeV3ytrR
EykJp1kiGgBWeI3LrGhc/LBwakSxCaVS159iea/CLwCmu30tvbv8dgDQRzmGi3t2
2q0NQ9z22DairMQvJ/bUggRWE+HqYKJuswk8WztY+XgnpajFYTPv8IfEdmRj+W0F
Dg+Vp3R2LoNkpfldvBJSaE0jx//URL13doe3ucoGFzJHEbGxQ1apjYsuOxaC4O/8
CrIr9Ut2MSF30kQVNmuNfix1F+V25qnWZA6nSPUA/kk/ih4sdG1sBZFIcj1GduAy
rkQE5QqNw+MB7OgLyNqwWrRakz4opY4VDEZ9TxhZWP++8jAjnk1NwApruHbpgvcd
3BxuiWyz/n9Opbv1QROOAjQsdiseAluQOJczK5ZEQefttYVXbyOihVZXgPyOF6PI
NtDYgTPKsp6mgJEY1paV5fITuF9fjssPzUFBntU2yG5cUNFcA4US7wEtSNyvMiyO
cbFaUy4FPcadcvUWXaglfqdRLAdZ/D6S6D0eqCYIaNjT2H754Tusjo2cW7vZXE6G
7e6NPiPhQ+KORRn3++JLjN1xwJRcrJUAjn1D+9+yaOjmDpNy/mEA9upAd1QsxUBH
djrTDA/Ll/h/ET4V9d9CR104j9xFVwbiteInqj7vwo5ZJnUdWtBFPgcumjNFIpiX
iTnGqmTmuvdA9kJB7HB+m/8g3uVCSldzeF4aqYpkSLGVmT+nNssEnnmWrVQR0Bdf
j07HReoQeuMDn+rhA6dgc5J++ZdYi+AFDBQ8ARCkj++cv9t9YhKgeCs9k65RwfnB
yfBSG8mUR48+H7sTrZdqFX+qSI2QDsy2EAj5vhsedq3k5chiC3mi7sFU5F+HzV9x
wWg7IkJnOOCXFEiKssoASIt5CkUODaItSPQB9O5i2bWzgVv/8UQaQLYmwEevPtsL
goAqI/tMHQGg0xY6wMtBHfVW1dw04+9zjGMXRMzEdAR0COrlpo8j3JfucItkrk+7
jRLmJMUAfNNW6wSCxhz6MXX/mazYeoUQKtmg9qLkCe+hYpp/HCYHj9hSGM6sNMTJ
nVLfYhJC9rc4ir7a+NDqaSwWFDejck65FRx6sR875d5OLBhOZsn3K08shJ7BO+qt
xd9XvQcSsW6uENmnP8ZnSokL3etR2wHk9d+E5r2kPPgkMq57XAc5t1HTKFtsS7dH
kEwJL1Q+IAJh0sgkrYj1satimYZIzx0XQnBP0a8r5xJSCIMu+eCh5NIvHd/1JJz0
esktSIldN+NJHs92umgDELYfuT6ExuCWM0FYrtckh0Swfi4WbyUCIqitCjdS2qrY
fvhd1Cu4G9zCTuXA13cWJgoaOuKhUQDDf4JD8S8d6bg29fjFsfEdaywqf+G+DdDu
bqnx5cVOzHpaOcXASHw1M/3WKcOAuD66vvU9hZWqvah30qRoJ/GH41CyrPQh+OEJ
uZPKLM9PHXWBIKo7BGMYY7qbewguY9EaIN/AEMc0kVWVSE1eiyCd/BDmLIUU9bbq
Sf2xvIaeVyO9OM5r+Gkw9iIaHQt6sGCiNhAmlbbTx/4Mlee/oE2TSdmuvjNkyusq
Sxp7k/+kvir/W2XdJO33pWlUedS+H1ljCF3MOwWygM7JjTgkVTAiNGWstZXZ91fl
9FazJvvQxNzHfG6la+uIp5mnlRiJMjofhm+MK+5kNjLjav8v+VfDJKHSfoBG56Yv
Yg8P91h7zooQXQYbNXjnteIsN8W8gHtvaVTWhZGTPIUuiMnxDr7bu2dikKHumXa5
VnwW01NPBcnynRxskkq/4gQ/DTIH5clPlCveVxF78A7Hd4fm/ITicTDImjNSVY92
se7FegEJ+CENecFK6tvdHRnwXy/YJSSSesZwike3e7k1T8SLZYqV3I3aVQSBke2T
SjSk540jpDswNehjWNh2TW67cy7zVQ57Ab/yyUHzUqEnXc6YmTga5MunntXNVa2Q
e6rYHqX3aTAleu/LuMbkW52YYDkkx2mcuQpG6AwrYVwq/+DJh8cL9uxA39leQoAT
zWcPvrp0gdyFKbdDMC9bwYJgvT5f+0IIa/bFPwoSLKV5KDgccDT/Vrf9nsKxK/5l
svWeu/aRA7GsULyVjxvYwr3i1oCogRhD2mkXu3e3ezK/s9PinbgLY54uKRTStXP4
B2UYXE1jI6CvmOZ3KalrtYi9BgmEUphMgcEec4ecV6DqQsavbAfErDZ0AqpH+3XW
SDhHiCuQ7ImGQltC4Hp6zJg0XRtrhXPgl1UIhdUKbftbrL4lS0hoNG17irG7neDr
tgMPt9/HzTrEWCDEA90orkAwt2Ix/ky/Py46W8n05P06XZOI72DiGazpoK5HDhrg
qEVddb/Nuxuje4IbKLkT4ted9JXU8aIk+DX/wWyrXCKGOs05nPSaH5/GqO89noxZ
UTGParN7rh1qieozWoVk5rYmG4ylbedC8qTnTO42MMlAxziotfzAqLYPXb5XjtYx
Yhv/HRMc2IO+H7ij6LaTE9XpOwpZuyhZSSMPLeyO6Z5f88uxVJdV0fj9WMk7fXA6
37qS0FVMxoUDKUvXhl5WV1j5IR55/CvUJUoC1ET8ksYZh3gLuMXTepZS/ki6J3M6
Zh/Ede7YhJ18Heb96ncHUZV6A9D9EFJikJOSp3fgrQsJb9vP64jVrLjTaCpev1H9
7+JMMiHiJer3thOang/vhqz+Bj4eklMzwBAbGZo9X/wkGKKUvQsQLHgKktBUskoU
ZxsnlrjY36qlTj364xhjpcnq/zgOSPGVCZfFpwuu1fJ+1SqHhagJ9JZCXSbX2i5a
Tp9TjrIzsv5Nsc3iskHqIXpLfbjQ8rvfofFvw6uFk0/nTtpDq628aq8DXi+2bDCS
Htym1/9j10kBhqYCTxbN7YNfg+/iyM3D6nj/H3g5mztZTOP7XTcgsfBrfmFGIjlt
cHIaggW5Vwwb6Fknu2mI1tZKTl6qp5Vl82nbQvSN2jKCYoTumWwIe6d4klxm78Pm
WrxuD7KhI6b2qbYyXPqApfQRQJBos/FH02mSwkh8I6Tre4jPK+fCkaeCR9Mau2Dm
uuYTY/WliD4U0icWDPRG2fhWdOOtSUwSCoeGQ1pdm+PuK7l6mMuhzvQe8/3Tt/nn
YhRjV1uH/OIFiYZfBpOLaoIhVC9NcjHQECktc6+PdRLnWIRPR9S7jLpBuWe3ArmA
M6Y3Ch3mhzL5hzHxrwT84E6ZPukWthTDcoRZ++2nTtvy9VmRNRZAQ8xJ5ow3eB7+
OB1QpIWfXheOw2BjWhV6Vo89qGpEaP0oeAfF6t1tjvexChEj4zdFNkl96xaLo79p
4WNjtdXv7g6IlrKCr6zIfEhms6j2AbXjkkUdfZTeqZP7kAyheFKACWlAZX+vh5Zd
2MBcDsE+6CQ9Y735UxrXNULmaSdgNQNsmc7bV8A5fSEhngqKXEXN6bHYQpLn8O6o
KBb4wv7kmxEXF3gcPq2nC3hR8pDRIl1QXdMYLl//GbB280B3QosapnaldiC/opjB
dcx42QDEJUHmhQ/j8klSej/9ORR8AXt9LDqz/7RRF+06UmlF+iYQipPnbyfpcJJp
EVFj7+HMctS+IZUGZm2CmjehbWN7DseMoI+pnP+TleqK7Stzawxan8oIQnqiXJqg
ofdErt73KZPV/Q+SmdPFnGpKHzS/ruAsd/vEIWAZp0lgC33D+DhU8HzyZxWqV51N
B8U7ofaB0ResF+apwLU8/Atk83X7+0VyDz/I9u7BjUxrSytLgRK6G8hTC2/aA9Z3
83766eEMj1HEfbZ2aEHWBFJ4IHLs9HfS/J7OWevS2tCupuEqoYMg18qkuRoMa7sK
nQi2YJn/8SZpLvGfF8hf7vmjXFt1+e0YBtfYPP8f51sI0BKH8e2KyFfocbm9WILz
PdjnabMLEdXQPRuZm9Hu18xpBKkgKVVEHD5CUQwSj9CcyeOl2Sx6zcpvYR3wUwin
nufP7oOY29FwymWItHLBH+2KvV1B04WhmzoP5ZNwxDOO0WoMAaCydE4wgeYzZoaE
42dY9DNNyDuZHDO/xEYAao2o4Qc3K3qPDOHBOEG8pDs0+Rcls6V4iu/def9jERjo
m934SoM/qaHtrzIrD1xNuTrO0u2iR+CzUq9RiCu6YoiGf7ZuB9GVggExt1jCdx1L
jfwAMmth1xgJeqjGu3VRuDORGOnpUbkRWSnrpV+FoGGzP4vD1vdSMJoh7HE114GI
k9rW8UvvawuJ97DIU0tw+B+PcfKyXn/a046dxUrXicLNR8/IQsD234yRro6/GYgz
p+iDBlRgfz81KltnghAw7fojAd2TETF+tBCoygBGmM4KU9r3B2Uo0ayqSRRxQo46
I/0+uKC9bdKdCTca5dObzpzKEalWrHANI6/ANbcN+GK0kwm8TlqIrET4UhzJTIs7
8AYL9v9bCLZ204KADOvkzLS+xqaFrS/gwpouy1CQu7lBKzggsqBa+YxVqwdffJzz
yVm1iJPq9PeACGhh0yqFunbseuzJIO4amQ8HvroRxeh0L10Q3rvhOf7ixhBtz8Rc
CO05VUBIx+zKn98I0/YwCc2RGQznSlQCzgmUzsKDF0iMh/9SO4fQOQv2mxcnx9yx
5R0QO1RrAmUlpR0rKU+jMg5+vu1ZGW5JxkeVtdnJv0OV4dC/ZcEOMrRw90ymxF/4
J4M4bKVch370mj0sdQoWlYreudZwS3kpR+2UgDNQMV/yQklChjfsJ0t2d1eWda8Q
ie5l3gZzVO1JzTqwLJIa+Q/SO2nxXHl+tVKgMDbNrl01z1lY7UsoCAdVmoEJEwnZ
nbsta+fbplG/H95dBbv4Wr/uQL+6JMQSvyBV0YT9Zsh7bpiSyBzED8g9/7LMM3tN
6MpUirR+uJB7kd+WF/oyOrkFujgq/ZGHN3yG9znqJmXzPKicQ7jyGUm1fmQC98xB
IbaQAEVSpSVAB4AwoYgQt9ykk4M7LuObq2FZL91HUc1yUNRgTT0ZarUFvGq9cDHG
+aUbGBXBInTmW/K+aV1PBB5a2/C4iPlS5wu1/Yru5abAdAIFkWSQyoLZw9bkOW2k
dxTNoGY/0C8ECCTVRGil7Lmlv2jJV6UJyaInGz5FVdEOF0TojrtMknMKde6QYavK
ra89D/ICuOhH29tDFhIVTYhkWOHIVmQjE7fdoiDmC8ji7HqZfruycryeC2VvZyfH
C7nCHiWO+hZe6aFV21PP7ySKdnEJ7EXx+YkJ/tbuLjiLfi4/D0QTk1ngKTXiHrwf
7PCVk6wEzLV7piNY4rv+zfjCwfcoBwiSsIG8AIJ7fRMWE3kbmyvZWPl7R9wXmR35
pfjglrV7xkgfua6sFMglP51T8aDvy/96kWBeU1DbYIdIrLvj5a6FL4bIPp1Lst4O
lHO0ICKxbMWF6sYGH3gNRvmwR+QEl9aTAmVicuwlpdnKiUeYDt8VewYehvQ1+a8A
mke7pOUhCvLNmOlpLdqygYeTCiJQhcQ1WVUCCK6InyxqQ2ICUJZ6Ex3IuMtKFXgz
riJ2WbetoERjrPOIS4ldzniLxw4Vix/FIkkx6lqZ8dAjE424jSvJj7shrM0lguLx
WX57ygMYoU3TTD7H3D6gjgypgVRddc6X6lxuJffR8LHfr1lQPa3SXH3RE1w93QZG
h/qxc1tmTDzFzlSYp7VuKwjrDHrUguvUJHSZt+oYDAVS/Urw57EziscuHDCAr8KN
ecKY3TQZMgLZ/k4ywTPx/Hb32Ir/JuzKSO40UkFZXae4kF7k4u0ImwIiLlKCvlxl
TfqlHkrXKbSHB00t/Z5LrTwEU3pFNcAmFq35BogEi8BuR9dLtp6zqVGOTOo3me/e
9fB/KHtyF614i+KQyxCDSqyldpuCR4k3xjbUVFChJKFgiXy6g4qL1b+BEqTSRpH8
A/taZOEUJIAHFqwyjkp/vCG0QtLaNFvSHTeNw5O3Z/Va/vQpUJ2VySoT2jLco0X2
7tPn9V/DornrMRuEdQEENgot9JvGgQQ2/FhiODEx3wo9fENhpSokIPYf50ju+zFS
c+gQglWNxMxGWWefWVT98BA/HRN4sMqJ/IieaggsHVdHupxZCFBseYfYXyml2w17
5i1P2i2p2yOUsKKEs417f2d+YNAozSkhVaIrPBq5IauG9uo9/46iuN58tK/UstC5
aXO2sU4VqAqNQ7tSmKCoY9yIOrUktlJ05OymMKzsf9Rwk+qzEo9dOtwrCk/MVWHG
GNF88qk+WqEsFYpsGwnJmWmoxdEEmOFtfMmoEov96HSWMzQZz5stQxc4BQ8hkMSd
pW7hp8cHuLpUkhLiAsAMzL2oID6gpKvVADfVJZL/QVyu2fPxkmxh83fD3Rza361D
s6gsRnpQvl2WhhL5ykwV/Ia1awbDcyMv6Kozdnm0AWdtWTvluToh7WXDFjZp260e
r58KT61eS6/8N+QqG5BCcW+GPixuQYx65g0fq7wZ/xp1y5ttUPj1H0qTuSwE9o3n
nEh5//lnia3CfE7JenNkF9qQK9owuVf5sE/pF4K2qVj4QSi63QsD5rVp8pxIW2U0
d0kzCNcId8vfRAtfPpv0Eo9ll9CyIi6aCK9E/j9kosV2QLdD01yCneK1uhnUe5Af
ujSatfgTECKVepVbba56JkSBIq5BAziqC8hBvNHMjVNsEvAfNyzmuAEsKXuWR+aH
P2EStR1iWXzqxGy8Jdj3eGTbPZweS34Zw7WSKXfxzEcMvmbByBMVzZ8k5OWVBDBD
f5U95XWWtjcL7wQOk8rgZ+5KP76tTO8QEA7Paz9BZYrA5nBGcPzpaieYvLrtMbbt
ExCpQoAUnfluGGKnVfB/qHH+KFfI0ji5JejBJXsNYpAgmxZt6Pwoztlvp/bh7BFz
uHDmdOyjcvGhrRtwZv1gqzfe9Pxcdc3MINuHnhWWNahspYPflFMN/0Merh8v6LG2
uU5hgypRHprWnGqvDqOjkp9AaK4fuGg9UPBjR90r5SC0lNiXOSWgIJRci3QmTk+X
CDLABM5mLv8pXzGkWe6muje/6UY4Wj2wv4UxzEYfdn8hxn0wQR3Cdgpu1Xw5OMbf
ILZIZPffbY/Jbz/erCtd4WBW8j2ek0VRlw3zILy8azOVCcRS3vxVqRlyeuSxeZC/
C8G1lVLoypaGgp5nA7KLCVsw+Ob4xS52F8yw0taklIRRo3/KJNFysIvszuw+AM69
/PvIl2FPI7R0NhPwXiMdHJ+1HUNbxqLzFKiPLkruMzpxiW3T4TVyg4Gb4gxaQD5A
AhRi3n+h/wAXRyzKn0TvnZ8GuwxbsA3HEWxu9hbpVKvsiAGMpya0rXcuEcA5BncW
+tC7hxToWTE8Hq2WlCQHIMFhvYd+C6qu0i+w3eBrWLPI1vsRlBq3YPVnkR4jcrq0
Q7utKB5BCy4DAPKrPLQNjmrAUr/lNxgw5WOiGvrQz5TdOWW4oK9lUcHUvqofAqz2
+HY+yfKS13h2UPn13bQGGcEU1nePPCXG4+Gl3VJBuulSMd7HVR1Q/7RvNaHeNZOy
AtR6Z82KDxVV0nqtfM1SwQHwnm0YjKtj85KibMtPsTWr23ZRqHZM8gkBcm1W/fxl
VpOq/bse9AUPZKXOTVeLgG53ZwA0xhNOtYOaECU/erWpqdIauANCyRMC5W8Et0an
Axmxp9mh+1kvd7b6wNEHok4R6cQ1I8yB4t0R2yIvK0OrelrdBa/gDTjwFuBgXtFV
LbTWMxEguNpnNx6I2kni0A1L8n6vo3J+ShA1rGzrA5JENynnD4qLH5Naji7cXE+k
zA0ncxS5p4uPKv+9h1fqEbJkmeOsYvQh0p7IZMBz9qt1M+bKE5nKdKbrerbCSv5c
CEJa1wMcqiIaYkPJb1sC2K5hhiqOUlyU3ykCMVmAgSQQzmD+SpbB6JAeck3GbJWq
w7a53VMT35bhJV/VxJMO0JYQI+tiYQW9YOujqWRNoAlK4WSPv1xQCuKvSJiPedhu
yZWZGmJDn1sDIxjG0THZSXU/yJ2V1pUpHLsZTbfBzMYhpdPHAFGGe/U636jGvV7p
5PeyjyxNyurqwRoho3TZPcWIO349vYXC/gUeoG4aXtNQSGpef9SXXgXqNqwVeFrN
40vvNCc+dT0KrsK62bYUqlz1n+18S/Cgd1qBrEd4OJ3w+7Hufy50bgDRSp2rFufh
cz5bsa1hQ+DnTfi2XJenILEnu7YpmSqQ+ZS6U4HivPF6DKW3RPfJ5OegErDkZtmK
kzjwyASYVUffR6fZN9EOodF6aLmaa3yf2jg1eYnEZviLGMB4bM5TUI29CclfJzbf
pEuCnNpa0FdAddPF3OR46tMuwk51pe+x/WqmHzBpstgT1sXocVDn+iN3o5EhPSju
D85Xz7PupBKwBDieIIVrY5Wjc1NY3pYhR/v9La2XOtNZ/2jq8QqsHKbmo16HNuDW
wx8920ycqOzscJntUbNqQB4cK+GO+PD0uc0i92n7iFfF7/+FAB3jU9ZqQQLmtirY
3thdqotuL8m1lGoTfydw1QuyYt94VgQ9h8YMd4h3bh1hOTKHb6x0nscGxCZK7CqS
uHB4O41LWxyq+iqAvy8DW5j4eG8OFZZoUimVlH11ECBD5U3dTXWWn+Iti2zozyxR
rAAx7nFS5IhUZHaf30ODH0HSe6LwrOu5Ti90M4SVjdSDDg27P/1KRUWGhkaWf7zF
nQCSMuF+7ToRdp8FEDoN54B+jb6VuCsL2sjGPbNFqSTPSGKBctFWmAqYDfTfk8sI
Z5CZR58T+01ivaMzU4Sk9SDvClXTlQf0dJU2yZlNbrkXV0i38I2pcbem6sMcps64
5odP021cvmPfMfX/J3SuaniZhNoWasvWktZJOsdqJRxm/RGEV32IwE1CV+9ARxOA
QirXbWbsKuorKO+GRwavWGYe9Ih9nRpbys5MDLdncJqWSI8RTGqhkJ8N2SNWCfiE
YK5Ox7Xm73/nmrlZh73572Ksuoj/tuBMg3kTyyqZIKmw2unhrt0OXZbmi9Zi/ewd
APqKX7ktH71kwJNV3WDkuthfhMVrVbumc254FxI02+bIN1xO/p9+26jfT1PdNz8P
XtnAQm7n5RDnAy+leQcZZJzzXtytFmrH6xO99dW1jj8uhKcDvpQe8ELm/iugjhq3
fUzPL5nU9EywO2IcnJ6ktuFnbebNSW7W4IIwqCW2lg55/dlEKiMF6rj6FirW2qc/
uiQ2S3EdqA8YAI/YR4g++FBpaI9jK3U+RezUdne4PLmy9FHoeFUbQed8T/jA+kDh
VDE7OTuzlbAFpI1UY1rPw4BhoU1SLqZeuKljB/Gq7Sk2DwvCQFU0Itjb7Zf2TqMF
oJs7SOhOt8MGAEV4FaKUfwuNu23NMY84yunIZq33+1BAO/uDGRYAIKIUBb2qOOp2
N0ssnlxsOOSw3Hjf4AhySxFw4a/WLTa0r1ZCeTqgAZ85mNJU7Dv2AsTC7FLzAalv
lmdB8MUOkUcsSVheU3zhqH3izyHjMCb+M5xGGNUmCdF06LjxQmulSszCV2qEk8e3
qCDmCI5nsX40kly5T1jvE3UHfrwc2gYYkdgTz/LEIYJFv9lqpBD4CDmqXpiVTYm7
UErxmbNvd9yX3MjK8vz0SyttxpcaOxK69haCK1ASJXe6fTdhMg+H8FaSo+KSNMwq
jQDMcK+h/RKofrvmcW10Y82EnAji/hTLmCvEE/zCAXCLbaujY4WOQKLCrDI2+wuH
n5LEQrHedv8IT/jE6npICc/zH8ZEZxP9RrXL9gaQftxrSGGksRfJ/oZYL5nbNOqv
lZKRxSKKXEBqJggPCcShqHRxjX9n/ZEOvkEJsdeHPo1+5GpF4XEvzYOWzUZl2ONq
EqQGlxrmDKkgZ2s+SzS4zZIwqsAwTiYcMuVy+Y7Tir6V/sBDDGqzyXgCSX9qP+ZN
jH2d1Yk80b3sRXbBHN/felqYSYFTqWJpiG5rbEy+wA4lkVgm39pd/TX7hcudqZaY
kZ+GutQc4RqD40+XpUhfuQe2Hdy9LSH74C9Dag7sim2y+eZGs9KLqcYbQVqhvMpQ
fmX4aPCOIW7RH6QzLhRYldixtcolyxkV63xeBgYhrycmPuD54KPgSJGQ3PgUmXeY
q9pu6JpRcwB+Fi0nnTANzTw8jWOthVJPcoBeFQckRrZ8Fap5mBO08qqnlUA970/v
yuR5aV4Z6pPU88YEXFLfChyGTnitYhze+/E6ZoRgPh1/ov7o5j/Z+m2ha//hTe0q
P9SX2+r1bKZSPlJkrpgS7X1e7dcTtXTuYSMh3jkJ6StsKs9cXCHEc/ACsNsUMkkd
uB/bNTDWB2f0JPn/JcxxxdGDcUCdDCypJAJaN1uckDiWpB7Msun4+W3JyeKe+EMc
S/vobPjTvyLarHja2sZA0WI70WmTBLSqjAvRD8pI40GdDy1WW+ikja1Icep0Aki4
28gb2T0aHGBueJxbEp3ONzICTNbWnk4Yac8TfbnJRiVLaVtXVROp9Yg8i22gLHgl
pAy8NdfYri1/kv56XNv4G+dqXpKaH5WTGP+7D1CjixXABzyY+2YrTZ2pf0fsIbPf
WNVxcxJoNHaFb2wLW126mQeBI0flOJVefxj9BEH9dmKQOet6lEbi7/j+msc+tk7f
tv0lcji0aD6OItaLiGVmzEh0bsmpCCDruNy0lgnkdPzINSgawDOg5kHmyvmY21zV
HqT+4gCONKUy9BbJI1rqVjhrVcRAnDbkuyATX3gouEO4mcKl5PGIWV25FNXuLiy4
DDyhmN6UHDszbS9oMpFLVxHzB5lKU9q6MCwkmpz6o/2MI0bVnu5dViT/I4p58Phg
GreErrkYqD6EmsTIjXTXay9zObChzCrlv4ZUgVHuzZH6GAXnCv4F7DWmldK9dSSM
67pN4BeVAQZxH1fkAfC6gRAdWF5R0BbejXUVdYRHZLV06hLJiZLZEXrSwfqdqaP7
+3MXbUUao48LqXOJE0uxzezU6BeWYQlKOmjXKpyBf7bwdf0AGX7EVgmS9yij/8Eh
eUEKSxo/TU7e2h/hnTsRNkFrYwIXivaPla0smMbLIeZ1Z2RXs8aMNWPIa6dbZiKB
0981kULoms36nCXcs2Q29ad7jpFp8W8wrNuOGYKx1dlbssKdNeIU8OxZSMcj6a9x
B1AVcxIVdhq7MVMiid/j9XlRcIp1MdALiRPuBQBC17yhEyb1AQmTCZPtJiekoHK7
+zF2sm1pH6ajOgzfMS85Kmy2ffYZXmgCulsoJLIniqwrmoWum86ucpSOOLd1axnV
pNfEzyTOX1+xVvH0iVDLMOv7O5Ikw62HYbBqKe/dHGzR8izDM7gDZ1O6eUHJvbZz
4lEPDWc13b3J05Jk3CTwgtf0X5nSKmxWC7vKumdxgZCWUNAdn4gJvzJsjLPA+QuI
cAbfReVNjPhHOjdffrViTpFYVeYDzk+4hZxPK3RGtZzBTO0uO3ixutLdsniqyRf9
eAfv7toTQy8M2sXpJz5yAqshoszs8OAoOOoIzbYZWyif2lifzusaVIRq/tajzaBH
alrZVs5W45OJkBhCkNzGwuBDdod74IU4fmcSlJTJHT9h6PbboL3Bqm/0BvZGTXJ/
M1lXJ+sOXL/LZbmrP/Eg3faTxnaE9z+WVlsL2ePURU0x7MXkyQW4pSu8YlfJaaS2
qXigalv2BjOstfuJSQJ4APxByDuaH+6Nv797RqbdwC9BdW/JratBA6VfV+IKJk58
wxCyJ89SQB6PgvbIdoFPhI3yQQdwvIwYahneq+0qmhl42eSofLTLaBXFnxs69Idr
rbj3VzcNhdSa47RfGvRenE0zIUnIMNWOEUmL4qV0vQfLHBWoWfEvlnSQmV2tPQfA
Fs3KlYUUNcz4LLYIc/Ph65zf36aXvopZk6en9TaQcLiyFrqHZljgN+LKMD/nXvee
BEHvFjWQYKbEaTNBYFl3GYP/aJYe6dC+Py55d9B5W+JQwnkzhtGe2UeBFanBWYn4
ZAbJugk3UoF9vGIKCeMpN9O880EkejYTlrTjxijjosxMw0dQMmY2wWco4OCV8SuT
Rsj7h7Y1ATbZ1eHM/jZQsPtIn2JLUblDaSbALcRBuaBTCEu6rUqOwwREGwf2PlmG
BH6JnNW0zETLm6eX1S7rxj8rpd8Pt2a1sixXbB/a+/2q2KOE4WVlj99ifulZ1exd
XdOKeddeeq6hy1+cZj4o7hl9NgA2wCQH5T786/rOD2P9NvBDSoG/rOxZzhq6kzcO
HTnfj4MJlyLCfS7wxT083bmz2E5b+xTfeydcsWhiWROjspdl8iPe/xVDuLjeanh/
d43l3C/oO3gQxr5JPSFsckXH1sL3MV5hWZf/n2Mt/BweYav6MyrObg6G88fPceTw
ZjNBe74tVTb3qPLNEBbV/4jYWqrs6pOdGbUxkC5LNJqrTealkVEzbIyfHecJDVIj
Q0ZItLLKsLHzHyujAV9VjIl3pCfKtUik4mWjDaalgOYRXDiRYAesf4NBFwuE1T5W
sK6xg6saBhSFWD7UZifumYObZL8sVAznyhZCs2Vsfpuesq/7ydCPOpU/i/tdHETV
p/EEAdkMZ2tdwYgqp224p0JRBRwzI/or1oTExY/6KcOCxlQ5OewppYhCEJzfs6YO
nabIDJ0n2rKEPbNNLa6SgFBEpDfyt4xkTjfkwk3R9y5sLBRvunZES6BRkA9k0MZ3
9EVG+eFQZx8u/33U4W9dp7CTMrdroqVj+gYKTtcGqZxxY9XuCP/k+iq8iCOdCHOi
GVuPAABmzSjkiTIMNaZZQP73cuZ6U5Aoy7GezQdChyICg3Ga4ZIeNlPLqUX5zMKb
FX/BHieEReuMW9wokHI35UcX67KpWUx9tE1BjVpJ/11YOZQVW056gP6YHpkkyO2R
qujvGbnlBNeqxBpRafwj8R7eAcn71x3SOs+rWK5t8w4i9+17QtkF8OBxPYPVkCPk
zQyJVRoyyeliCr7n7p2CwJY/dNuG3x1/5Xu78Ur5mCDGfq/seJL/IOzOoI+KklEb
U1DpEi+ygp1Rdg0urNBp5gXtXEAzdjA5LyBU1eBQaBXmWHL9zP1R7awQfQWj/l56
n9tch7de6O6AqCypTi0dV/SM7APc64qjGg8HBP5sN0HDzNCJYCXxRdGpwNzk4jR4
yteXlPmkXzlptfDwYKDlEf2kVOf6W0NADY2tz6CbbtYukpHXWK1DWvWBlmKaNGEI
IvEeqdBs33JGobXomcFLJ2vQYxHZUDPgA+MOji8aHrNc06W35XQG9H/sQq/QaZ8h
VMVtmKH03FQKzGX0X3yNy5lD0FnITIQt+ecQxtZ7Zc6VnbSrKID37m4DW/WlQNav
M011owWinFsjDNYIndDv+gPfFQgVddc4Zsmuz0k4iAK9U776pYCSSAdOuUhnkTws
B9oFULUOWV2Y0seqVXDHl1J2bans9MNed2Tem4JNg83c6fAw36Ii1vVbghN2eRAc
wufEovYS82cmHWMdMgH9AnAFDCWH8G0ad+DL64S3hdMimAAGn4zBlgPkQRhWeU2A
qBPdx7DDzHNFlNIca8WUgPq09D1VzkP2h5gb5DpcYry1A1ynRr1tEWvuQkcVV/Ba
a/FvZhddRwS/nNuiSqjRVf+R4ZvpefMVBCICXOp+NQBvNAcUGraJ+kyEW5hiD5K5
kUb97UKabNHWBRTRZ40XHJfXL9PKXDUAnnYI+aBVmkGFHBR6o2ySzWlSRU92eOrS
1vno3bcHPMN7vGpVPoT6ytfhifdRQ+78is6rhnUr+3hjG7i6lKaAenN7uS6Uw6XF
owyciupUObMDBE5HoOXmk/lSsoH2h1S7wiY5OO3LnCUmk4BLCL3Anc9hSzCW09nB
cvCZ5OlwUpL/6IC+AYCasjqMe/dXBjwWSLUAd/bomrgsJXddiETXs5WKWPM2iqjp
J1ykRFLfiW3MEHidHu/nWJuFIal3F/m4hAx4TmG1bpzdDwU95ObrPbEpFZgMNFxR
TVl/LiMgb8oYDt7uP+dk5LM3IFmHB9nhWKdp3S3w6GrlGIUIheHVQFLns7o11XSc
ttDTRvC42MR58OxX6yRMCJNhKL+/1db13MOCs1FCqhUhp3mnDryuUFOGXn3TeXPK
zoX3v0vBAH/Qkndmf2yFzScISl2T2388yeg4ynlwbGCyCCO0Sbq8dwrhryLjRmGL
SwizJ1M0nml6VPZiDQM8dnAf+qRSJJoYFPzAMmD11VlHBzj9YxGEtroDC+glo6kP
1Q8tfpTWLRhj+P6VSvP1CvLbBAzQwF0eI/xgPs24LNWJWIZ51mXVsWPeZxWgGPQq
JAK3go+a/KvvNLkS7mDIYfXjrzkwDwQ7A/AQfqXHR4rQRxrJ5oY9OCgeIPZjVThY
9QNwu+9llSOuOkD5gWCFPahwzZqJy7TcNhEzSGUD+cSl1D3fVijXfclBvXGzo+ED
VO8WJLPxKCGot58xf0S+wo079shy9j5BpUuh1tmuAfcyGXyqrnIU7EkjkbGvxmXJ
33ovdRqcg9QQ78H2H9PdSgiCxWF3zoD0KlPDi9JQ8/qbZQW6PM7bPm0rwD4vxx7K
9yQXko5P34nlOvKPNrtO/pMCP2pQAMaf5D1kt5WaO/cbLjSZPq37prkhyWcW3/BW
nMyX1ilRi1SevDPl8jGGmb8Eh8uHowJz5azMT1Ud1Gj0i9ps+KRVo1fC91VZV2tO
j8iGv35DzcLbVviERC52Ii/OzACMnA4Pxj4SIY/eCqYP5BOU0e/MLlCm2/lOY17/
z5u/+WovbUHSH8ZpnUpzeTxDQHon6qVISq8YXqhCvG53A6agcdag4ZkjGagGpA0Z
L5sQypMVJqNPFxC2HvJGwjSjmT5YWW31Iqk3loOIDL3XK/ocRN7m3idiAVCgySOv
fGJJNpso0rYe2tXMoAI3AuHS6vz5jmOkVZHh4MbwINxaJOT10XPQu2BaWO73XWqb
e3pMuMe/FMdwueJ1VQ3YZPbLlyBuVznOSPFrUJ8tjzzSlHEiVWsPWAK5rqZLwMnF
JvQ1QMJmXRkh2ynqqF75LxF3IEEyRxEbE8PGy9bjvuZjFwdq58Hl3OfnY86aUaOS
KFEC25U2klYYZAQpdgNcl1Q5q87u0hvOdrUNe7QLKqjNz2ENs8fIJcxt5sVAVfvb
pMQyqOsDdUwuaNuzL9aSHgGXJz9fEK+uBYGeKrrxkfjtiHDcQ9ZkC5wiHQJUrXvm
AnHDHDJVSU2tv3oHaL85tXp740/+qL4s2P5mZw2tZZ86jTTeusgeapfUPRGhjnS3
EuKW0nRpV7YNAtx6f129+Q3S5gN12hM69ijZ2o3hKc35fD2CT3TY91xnS7KbwzAd
XgneF5PAdXhNhjy2vk0ivesS6uqLAz+wUpNWR1jS+bRmYxJCb7n2tK0i8erDXE9g
amLWS092aEQZXuB7bPzeTtPhF5GESPFMvx+OnhC33/hcg+x3fJ9KcO0LtS7A6x8h
7IL/bV3moMYKai4EiX3oI4+Pl1DEkFJulW+xI4jx0ypjM8BBcbXmtQx1f58ywY44
WYQ2QRWIdrucSl9QOCYrVdp07VrvZQpzpcy63JsOQJuHxKBmfXeCD1c3rTyZmMSn
PdNeN5ZH9j9RxuWJLXjHBhnJ8hlckzLMMEcXa1pmfropuWeBQNoTdGsPLV2/xjqC
dxKdglwc2hUrmNPp1gsaGqWtVwU4YCUXuJm9THriNhTRrEbT99q6IB21ntyEcbQV
i7S8VgWT/9sZApjHmfVbU3f/TVAF5gLlvIi4Qxt2kwE8+mABh2f34jwiIHXNmlIM
fFluVtdfsYNq1sN1rBlgJYXaoWIiFA8obuJwlHnE+FdIPuiDZrcca16Q104JbrlF
g1LtUoawUcfWIe/rpHFChpsxLSyG8hawtd46RhynMJ6EnFFuq/p2oqZuffErT14+
CXx1+IQSxyWpt63rtm8phuZO5eYaeEW/oW3hlyWPJGHsNZJf4X9Jh4hdHVimzv4i
zQQj1kKbihF5Sp/PTPxJ0n80fE0MnfgBfnlBPrK4UGa9inBLEL1AAHjthtGEHF2w
6JLeBg7OesmvC/uZC2Oeqjn0l1xsspEwfW7hgppUcZyRIyrGJ5XNrqQmtr0+hLal
YvmPmrlVbmcX2aqNY2ty5b31+HsAAUUU6VPcujlJsSTqt8rems5g+h60mKDZoEfJ
HhlEbLxTZ6+cPnaCWRmojpfzCWv16F7fp7TQBmlDeIYi68bq4QTW1XGKO1SsXwWx
sZwk/tnqMrafXInQZ6jlr9yz3fR8FYA8thFvqbsA8DBuI2OH7vn0laPvq/OTYpQ3
RTTQsk5K6lYmAUzjy02pvroT3zrm71DTy68mlyroK+3AwqUAeJhsHVe1WrXG+CFx
VNT3DFVXxWe+9aFrHrvKmlbPXADooA4DXN85Pp8qiE52iOg94o0wt9zvhykZnc06
auhFpc772+eRRJrt/xNeru/TWf0KoDKhMIHCKjcjLSyAj1id9L7fW8LSHCRfrbLr
CTpiwPkr5JkaKxGuuov2pFmGHGHcIhTvuHA4zj/m04o1JgeCmgIFX2gA3LMtf0Ys
/idIkYlTCRdnHl8yuUSGZQIwdP4U4ulctpgdAEaQdEMoL6lOUoiyzb46+aEp2tAB
yGAS+F+L0RDsPcNZXDI7GpDkOdybFB7yW7PjbGFk22v0wdcTrA3RN8txseq+9Ldr
UT25NC/wJrlzwIWPB3DiNut9vQPvySX8cc0ZkWIyQwivn5BzVtjExLly2IypZLPT
yxX5P2aL6MNnBZVMEAkoTht0nfowTqGpyoBZknXvk4cIYc0UcpjNIKS7iFQrFlZF
rjdqcD4wxeZMu10yrcS+5CliiiD8OaZMlyEXb2vPHNC9W6r4N7forVsQ5GP9Cf8Y
xudhZKq0dnRHKuLF+bLxA915ZZU2wmibGuXQrTCaZJknF1EV7eEjFl8M6I31rxnm
JizL5XvnuVS/hDxEJ3gVMKH/cIdsMladD7YR126Z8M4pmRe/hukWJAkcbUAVNBN/
pmkEg164gYCJX3+6r+5LPos/7K977fQ+8KJ9/V+DzZSxhVOBduTNXAhnjxIwhRZ0
BJy+WOtLPy28z336EvJH+ixglJCdKua72J/lYtFkCE/LyhGz0d4XGP/0IF091zAL
+K33yKu37f8URLa1+BPjGLlk9SMdp3ICxmJXq4Yo0FOiz0UwnmkLXFxtmWnZsIfd
qsHUEh19UOfeBE2PtV41XcYtFuWwT/i4hrTRrPw4S7iKDkRbes1iGreKikp0+2Tu
Uii3DlvFCW5e1putpY9CFXeAJskz68lLeIVmvaBLLEKgNWuBjN0hCp8t8Bbw/Bpr
qgVeOiyRSOBMnz8SJzoSkdtBHj0ofDF8LClvtR3IJZGUcI7NOS8HCFWwEvfx8QtU
hKYG+I8nvZFLULjFB7Kuq+ONnpAJl7cFLGwBeMGQk2XleopA3o/2m6NhO3nHk91F
scIR1ROJtoX2kLFqkIK/HG8t0CRIigqGBrwxm+Vb7brRhbthGDkbGyCTl6chkVMY
aQCgKcURe4ikQScl3EqQF9HikaJmolAMnQoemacg5YtVXO57Dd9GOafVIFrc6D46
LJVv9mLFdCRSewV2pC4bgIfZfuiYxhgHvW5A7VLJD9t2FufL57FVYXyJa5Vpk0+C
bHMeoWQREFXab//+3OFekLtpL2A9fNl1HIPqBxpuDGgMC8aqXcjGqIju16mz4Ka9
IdyTsTkWmSFmmYT0DsGPuqrsyyuARE4JpqvAU3ryDWXNv3qcJSSS4drARbfaYFEP
zjc8N/a7R4yiODkk7wnxImGPIMvIG0gmR3/iJu6iJoDa+6aE01JeCwrMHlVZ8H1W
qh1uamp+1cIFK02WYhmgOiO7xvpuVBNWCuQNJS6PRB32ZnNkNRCY/RC8cpDxIPbj
0rtrpYDgCkuUFnffRdyBIrbKFcL8nIoaH5jH+ADvzXWEIJJjFqAxnsfjK1Z4PCU9
3GOxm18pimsZY4bQ1vOYTxyMZc6/jDy+cLQzBxRlcWqHetQawIVD+AblKRdzvGuv
+tRa93419gShoim4DEOD+3F0TZZXBHmyePaE5LyHVs5AZcyI4qt8M0RxvOqtC756
AI1qznCy3HPbjsMk4g2nkCdUdnHZ6jcFouEmqeGnUQp6y/wPFQUfUDgPQpbLPufA
mhaszH1pPTx30SvsgFlqUb3gs5A0EeYBO8CeV2G5MEBbvIi+equFbDhU+5sWK8JC
Ex1soQIfAIH8Nydl7i28I975XDU/pqx6Hmj8dYDz9q9l+J1zgfYAjZuXY5J/qRO0
oj7T5dP4ughPDtgtGKxXeGgsAHNg+JmqaEorwvnymey7Pmi1+RClpSdrsjUAFDI5
ys75KfwhU5QDiQipLpnnj+AicvH/E3VqFYKi760PWt2Gdg0JfZduM4Hoidcw3Np2
OClmcXk1Wl4Hf1WgGo6QisVn5l7YykLGO97e/rXOOLOUVSpw0oEBIqomKuRSX1WC
LkpTACa4xMnDQfhNcj9J5xrOT435l9bVnN8ae7f+1uzC3QLW1WdoPAJkZ1eNkfRT
UQXY89rZwcVEDGKnQ8KSds7nztWHnO7rgcPnDDXH8dAVasbKDN3uzadL2JUExQlb
SGcY7FWZxL6H7WAv5G8x8ZzRTXgKmPJoCqPkbRkrjoDr7cEK9ZzD5WLTF4KlcdU7
9Tpj4whxkUYLk6mObIhOAAE6f5t0SMxCl8Fz3FpK01BczoN+I0anmGwzVsFaFtaf
U43jnI1MYwiaqtiqRCHB71HgtUJQFziyuCNGjR7Ot9u5a3g9NChTr4rCCI/Vww7+
81COX0pkqMeN/4vaRwd+T/ECgP2sdJ81zJA7rHVqmgaGXXW146duGzqgHWSiD0UZ
VV2SvNp/L/1y39Qlx2m8iIhfTpIH3uIKNIcUM7tpBGiiWWJ5T+F96iXT4j7BJceW
0KOlGJMxrNssE4De158wL6AO4ogq0HJliwVYjCqANir9gRweQcTAavW5Mq41d19A
XCfkUadY0TrC4TNlw+9RbvX3y7mgA4q7lCAiOUVFYYwGf7NjstcG3ttgtGX3EYvq
g5jaGMk3ep1QyObgNI6axTT/SYqcB+gt513EL8rnnAShL0Ww4+ChW4oe1oHxuD+H
nxiapu5gCExo64XMQ8+Nv2PlKXI/TYfM9c0i+u6w173WYHvADjFk6oAjNFe7mDyS
QwwQfhM0lxbDhebliAcwWNFJTEh0MY3On8SPIKRrs+eaFgJmlsFf0fR8kJ3nVVGh
eiMfM5ieZNXqNv7fDDGr03L1W3QOTOm66Q4XqIRnZN+BI9O29XnmdCq3eN2pHYdn
Xgufk6soq6zuzgnLfP3ihBoh6r0GY2kl1BEhVG7A1XYVPbRmREf2iqdCSz+fuLn/
BhAG4xkpKQIFh5/aOsTT5XJdjl1XGBem3eLWVAijpgd5CxnC3nGvaSzAbM0IRTcs
jGbZsvNqq65LQYAEbdT/1pS1Gh8tX+ImMtEezNLNHwQEc1uo8v7ircKiyf0PyjUM
GIUkSB4IVmxjENSr9t0gFwAzlwixjd2l35u6pcuqrvsgDuOFv+KsZDJ3gfFYG4xs
hMFz+7wTTVlv1xrAquOcKXI08nq2tLFc4o/cInmbALnKpSEw1rAv1XlPfrjZm8Fk
+i6OSkf83Tk8Jl5wBY/5WYowMnOUyV+/RROordp4noei9WBte2wqGE/37urB3vTg
ioCeQBtKgRwoep0E7Vd5wGc5xIRZlGHMo6vnRDfLj3rhAykg9YZNZ/Sy1C1dBr0+
PjwLi/AW0ToQszwfkd2mRfYoLZS4gZHTHfhnRH7gfIe6in4wkYB4FjY414U5sPwy
emGhr39uTPfMY3W+wxqsCQrq8GHMSFcTHcyScA3sp9iywtJf10jLvDnpcQN7oIYe
bSAgS4kykDmwRqC00+8RAOY4BJjFqG+EMOP76P8bDlwZRKh0+lCJRhD4kHRF59w8
9YTzmYGF25AKLPHCR9rf2DYYSV0MNY38pvMV8AyZpV0HaP9LxP2Z2NCLX/Wyp34A
dt5y1bKaTk3Zzqx8JbLOex0VYTtKMEdnc3BdQP0eENpZDnlvFbWIxfOvoPpI08pp
2KACQejMQwdpry3+m17r6fmx+v2Jy2+oRpVQnbyfEZS2UPyeHjuJgxlLAxlgoBbZ
fxbE+f5UXDpuZthcPMWrDqALjNmcI7b/qJ9aEpnDafRglsvOgGasmtNm60SSLWK6
PKN7ytjfSFURC0SNDxuGKmmG5/kECYrmRHfmN3xs/zra4hsr8IKApYKwmePirXHh
V0IDCGcscUnxZobbLefgeTV2MLVZJdc2RawCFCvpxlCqSQZk+Q8t4Ireem9Oqmjl
u710OV3mtBJqlepNgpzuzAnirWsWH12vNzztIg1KVOVncpXKTsISvLob21lyEld2
lLY5VX8GjhRjusN0uMaNpE7OqW7dpy9x4c8U3fhxODHqDF0XNR0tbuHJKwI5NHsG
ijhVpfCRlrKb+irEAdh29IrdW7ccdCvU5zWfyQl+bm1Meia3rHPnddbpGaKOw53X
rPIiPhuXxVDERteCWrpNbfShbpgif1sFTUkUru9HDFjJ6+ykixHtGp0Zy9R4Akdw
E5njHXdAFwUZNO8+tM+5RqpUf+EgG+TP5UX+k+As2R0Zz+bD1LPUV96Q3CTdU+EV
pexbt/yNbf30M5Wgkq75qQbr8FtYCdRcWgRWwbiLPX6aJ1Rd98YVakIhTxJkfNSB
2auk6ZLAiqWQC4r7hXlT78XbM3Io1r5qouGlHJnI/CNMziWZuVjUipND30s9vDA9
05lHkNNAMqr7Ct2R9J+9yK2SpUOkqJQswmtZyGjA3TgCloDsAeVUhkW7UhrTAMtU
hf3QeVbP8uhknG23WvhPIxRkavXGcyG4x/hASKuqpQQUHdBTtrrPS7W+W1DWS0hO
9TrpATDdi7F8mgR25HBzH9LQXvN6N2k6R8AVf239bGNBUkh8ZrukLsfuGCztaezh
7RL6MpPaaN4P8vNA3IoKjr7mRiPp5AA9dA1I+4qYBg6SUrizbg8FWbbHtHG+sPB/
dcLK44lSo/Vdexzc8HbaazSd/slMUs7+VIHrghzxPKJleMQ49RyW6yhGoepXZf/t
WSA2bBWFf95UPTK2Uxo0eOcZyZtRcFnXfo8HDdOv5MMMFf7+Pg0dRXrtvsRZejnk
yyhvlrGuQ7o/Hz26XvejQsygQfEtpCHeKGYD+hvlZiBBoyNGQMSs787kv8xprLch
AXNLDOdMX2e14a2hR+lbai+61muRqI5xDqnObdPQqOABM7AVBJ3oYWZecCglwtOT
mMkCkTAtWbNpxkTA1W6khLzocOoACxU80gi5Tf1JAZBjRkAxuMUIX26UA1v9kDfn
19cNDTlhwH5QEDGTLrHPbfGfj8YUd+dxxZhETcWZicjzBn7qWsavEWme7ALKk3L1
hrA3wz/JAvvAlv6St0/viHYQJsvRP46k0PDTMp3iMkRn9rfInBqgZIld0z2GchKt
AEUDFYQIjscWSIwEFFRbMbBlNF9OlyGOpPjcAJN34I4LUmkAFieT1ZL4NLsq9xcN
LeCs7cVZ1oKN3htLxSG7Me6lvLzZjy5AzSkwXLamTUS6+asTtxkLaTB70dyD+KH/
hEIaqxCh5vAL3nDkLXtri3Ti/VleOtfVkb64SoCJt5Q7Lnr8HxGM1IBlO48BQMIe
pd07UQqMSHKBGtODFWEh5G4dO7BeSDmiw6uioU9aM6FKchqqtcWRmmic/vqKkvL2
s4/m1PxBeiOB2dufy/oJ3mxIEZBpZm1l8TINBlfvLZRaMFpMVn9KPqJYbGqzXYb9
qaS2YdZMCvmk3xeWnHIKFAp+tUApw5e1PjBooiOuKhVVedAtQHPgZYGiJfVoRK/T
SgeWctLGhAsFmi6Knqc33Bwl4edgxhyni/rBcuCkNUyRNn6MqY2YSf+vuS2xvIuw
iFtT6Lng2l5qYRGC+gMdG286IsiNXkarSe88oFySZJmyx2eRKx+3jtPs3Kt58rtN
bYkM5ZT88KrZSXRwSs/T6KgTA29Fwv6laUdTkN/39UUBBlatIy2a4xddzs997ZMj
LQgCIr3YVDUJQ1JpfkAatZmnHE0U+IBwg/C95qsdlBklqLvsffxVudnnrllZX30Z
fDxv3apnXvIIWpHmatJCtmR1DrGMT2vUc3vvEwA/+d/JzZarral3o8Yjjni3g4Au
iHcbyjJAHttijCp+o/BEpfHndtlMWV15KRS7pdKMFxnWOKKDFKP0ylXJEHfw9zW0
KHIrS+tza6807GnHODLrUVBkKWvA/R3XjRxAPYJJLu9JSIaoJPqm+8bKoFnlTA4r
yb8Q1wPb8+PFpmhk7uw11oQH0ed7PLyzMrQJDYQwvwiLPkHFYua0h5IU1Krr1zHQ
jBHot8oaqdwS6QYYrMCKG845qymSw8w+X/J2VD/gSrePzlFTA+ZP/TsfcRrjn798
NjmGyc/H8bLJ/acat6B5NYOLG4t021pF3r0EmjWuu6jM6e4Rsxy1DgIDJ/wIn1f4
9pVyeoHtRcwVR38pX0oEjpkxg8RUSe3HnIIh+xrVPMdL114jwyMKYup641FQzVCs
36S2JvJGJxUFykhg3nc5oJjQMh46PI9rcHaERlvCY6+6D44g0IZ8Y5aslBov0r6V
w8VX3n/4acJn5rjZrqxjxOx5XW+vAki7d0UGHziWaW9R9PrmVyAeHtYrwbQvNYji
nd2gTn+JK7jMmcepJDhl4rW1tKE3HXv+qvJDMVjJIDHL56fNxPfGTOBdEXLBdjAR
zlro7Te0x+yhbvawTdPmKZYCciRIBVOwNtV4Ue1nh1tT37aEBLIlOPdCASHpw4/F
eyRioVmsSvDvhKAuUU3FcEw5m3H4xhuHs3WrE2ZiOL+BNIc/COF8cdGrCiMVNP9h
dOuLB5sLNdqDfCtPb//BjuX/0ClDt9GKhjXgsrWfeusVxdOEEUEspscE4nNKMJUd
chFlMD2K0hQsU96+XdeJDsbda3JYp8xurn3WxK8lFPz+02DujfQYRsZNVHLpSO0W
p10Oz0YuOdW5Bp0GtBsWAgLnEoF1yBFhdytu7RW+UZy+M1uiVdgytH/C+bxy/QBw
PsJSaWswaEwR+scvPRrI0nBybgABfVDXG5xWj0ox9BlfTZV3kmHOy4gly3cJscGJ
XWgqmUSX5PY+jzfSGyVfErtyOjjoGKe2weBfRPgZV8xcLKgzeoJNVgMkgqKf4OEI
PfFO/ymCp1c/o9OmxvfFtaSQZzNX50fxZZr6oFy1ZNF7hizIokNa3n2vKVxLtRGU
tmnESIipxlXfNoEIbzKzp+G//qdkB2dpMVCkIITz7qWZmBQdhAKO5s7pwMLvFiuQ
n8CFGJ5GEykLZWzOD+TFHqY42xCvUNhjfYmX6hUkuoElmpqtY2Ou2UlFysar2GXg
BG9RJAW2e7nuqsHmIYb1mJ0caXxZvkNRmjy1nlokKH7eyLEvOrzoCR5fOhO5g1cn
3dHsmeIktAvpRDHKXMafnjuA4NPen2tsPwOJ5Rajdhgss3dEanfps/bHFWYWVEgd
ucJQowSoppVF+GzdKqwf7+xJh04cL+gThKZe36J0OrHkQBflqxrGE775bSMvI2oT
MLx1FgZYhCqEHDe2tIa9VHRikcEc8IYVhtRFeESAHcnNh0IkapZ+1KPsP618VuLq
cV+1x8acQrKDfAB/P735lJL+5/gH5hZpiRq9y8jIcUgFdhlM8WQ4L7vzgy8p3GZ1
v53EmRfimaqgJ5P8ICqjHaJ6+biv3wL7m25kXjsusDtVP4NdEzh3FFdGNAVMnbEe
C7iK1VXDpisQLa75GNVx/j0HyF6NUxzo8I6NlFONdHRqguShKnWkvXPz2OTJaTJ6
GxOPakTDrKBa0wmzyIDSe620M6vItf/pJTmt32Gm3ZrPpxEG9vOWexazWNFxA1f4
az8OcAQk9iRN6beVS4SGYs0xH26FREyM+hMulge9Hj36C2xshNkwvXAh5tZJlpfB
4JFDLpPoBa20F6DmXGBUBDJBjnXzm9vToI3GuucLJF874vCRA4Klw8h5Gz9y353d
ze33wj/JvRPsw9fZCL9QIWjyyLOciVPSuI7ArH/5w+bZlGuFQlN4snFB1aRBJqJO
6o+3Sz+8zLQ7xh8/GJyV4VaHqHXpDOf9yj6PBxuXZvTCfkakr49dT50Afhw0ua9z
kLtOOQp3+55BuPuIccLxYVFKJjCFnInN6PML4m+7guJS6RPV6SpDg3f3seiZL4iq
aUyy4z1pVVXGVLzuusDqsv/yjNKSaFO14kM0JXntRxiqov9RHwDUjekp5W+xdHzt
ZKNl2ii6EvI/BmAPX63udyFrYTckbCC8oy5zKxX8l+onufYcRNdF1/xsaoOWcWBz
lcypZsMu/6lO24wQj1iGPT0AvfFndQp265S9f1bO9GH2AsxHgNKjl6J9ESX6xHvA
DPzq8iLSmkrUsiKLl9GPuoWzCeXnYM9+Kd8ShMNqaYMLhI/yRjxjdeXqJE6EjKG1
JZMMJxtQjoN7UtT5KpRgXbLPgyQ36mFOYVb/3JP4gMjkxDeA4/QRgq1v1OsQuLyl
y7cNpjIzmUUty+J8yoZ83MhOoLLu0s2CS2CYAYp7LLdt2oyxNKju5CvE6DZ3PR0F
M9a0TguWDi+a8dYuWqVUe5dk2CGfg+kvV/4Au9RpZ0l7bqaHxtVa0Mp4yFcaorc4
e1Rma6sAvaAgWDbU61+0cCj4gAFt1B2gkkosw5vKM4E5T/MbW1pDW2YCUlvc/p9s
nX7smM/eOwkgUokSMoFLjIZaLkCPXjhRo9AN//YFEyvP+DHo+k/gMbX+65ysqftt
2o5ZE31kX5Afs9eIXpRrdLAnVGyY9JHQXlH/yLT7MyXyTpEJqgaNd0CilNJaa9ke
bJ4KawH17nbfAlnsvXhGuCTuJxtDfkfO5lhapuxgGr6coyjF+QjAVbN9r9SmuJm6
rkgPpFqXlO2mWHOYhQSX4lYQgwOqYKBSvbsLJDKHIfYlD7L/QrLYM71Tn0E8eLr3
nxTAH/9+eh3DCrqzzKFJTVn9JI6CZU/1hxkNXhGo1ovP1uIHLBORj8J4iQH4Z8RW
d7l7h3W/y2WEY0K21wzFBEGhFddIUr5gnZOKZlHNksHogVYmfltxGXs7LV3zRcpK
JilgIgctltjhMVgnOCupUTUqkQ88PEXOVrCsdlqOapHHrJaiZOzL5bpmMdnUt79k
DcgL3GoSJwUhapFLbUBuQ+l17JYqI9IiZTYDZGucZA+Y9mIN9y6re313htq0Om/K
1I+p3qjVUihZI6sLEFjEgXeyM4/IYY94Du3y6zaI4+moapcqPV79NBdNrf3R6YeP
X1GtVq3taTYQuoebGzqgBRO6sXAHIRmarqSNo3jxLxTdTivPyT+/zcQoVuyy4NQs
CeFAz+g1wdqV5cZ+8g3EW8ZgU/xeUS6z0fuh2R8HMK236ce8M2jAPjtpzV3qr7lT
yG9taynVXKz6T7Ic/+LukVX8ByJM6zDQIOPuP2H2KHjqVE+EmqSJJ1TMJsCQI2UA
OpqaZTXSREnYSRLYusm4IkthEv9CJsomffD5unpYOlRXfnjob+tZdhq9nbn2nL1K
lSN20uEnouDoNrI+WwnJrH77VAfetqA5XSLafIBIkTkYZiO9SBiF28/YOmNzwd+r
8li1X8V/MktVcADWqGZE7MQmXSx2W/gepQT6AchD0VZyYbsgguHE5qQnrdqXKoJ7
6MgYRCOSux/ZX4AzrIWGw167B7Dvtp+yKQYZiSOORrL7eTKq5F4ubMuCKuu8y+bI
14N7V2r6GqevjC6DbLJZHVD1ZYsJ2T2wGZzxWXR8UzjdN53IEHgU752qFuZFKi3/
ygOGJa8Ds9c4cQBPebOg+VYHl8XwGFKtp2N01GY0xWHndBoEvKGaHq2X+E0MAMx0
8LTRQAtEy+WYRpj6y4db6+V/8KyB3Huqq2QfvnGd8fy13nzhbgr2HQjpXA0NVbnp
V+uW2hcyeBtGrgQZqfNxx6q22uG1M2PSHYd5PC8Qt7lIXdl1NfLPPrG4sEj3BKhq
Zob3nEKnoFsXnRySOU62H6eiSVQRQ0y6DYmFdohzW6R3Cu785doXP5RMvYxfBohP
bEWJUAGognsi4Z/yxgLKYqd7tozrfwO+JamzZbN/QCQGR1E37NSKmj4aJMzeoG8M
PvccKl5azXGmV2JbEc/fk2vPqXQz+SVxLxib8vRWD8xFDZMJe0WwCpij/ZO33hlp
nDwv/ef2w7cI4vziuz7gL55u8fdAPJ2Cu/GD4Sci1bjYLMo4WWVt26XC1DVkYv8a
SQmAo7x69K4BtxW8jFUmQQGsRUWZ8ahWKTc4XxWvAR7SBn6GuhnklgUAZ+ak3/iJ
BViDZuBDLAMYPXZRXzZyBS/FZQGdDK7fiCOBOqubz8nUmX4yrtwpM4n37JnsD3lA
OHw70Caadj0oCmUui/mXCGkSPmeTBhZYVZRlw6de7gyjohQ2wTmpDPpNEl9sV+Bi
/tNxFFgwImCp0S6n6/BUK45QvliyJH0slBEWWUlFrmVcP6GEWsp+mTepAUhisYto
WX8oEPoedbaZ3SN/DW8siQxpcqEf9tMuYM4EjnvrxZqQb6pS/UOUjARFp8CMYmw/
Gz2200U02ubXUr5YwUustWBVbV4mZrdjjYTSUtxsV6bTUkQkE97gf8q+MEeUFU+q
nPpdzv+YpMUK5DXdFS1zXW6DNkerZg1ELAHCe4d9+ykr5Bn5zzN0Lui2iVVm3Rp3
ZZ+kG4rlbGS7p2IA+8UIqHPye920TrodtyQBsxfsbr1pGmmPaoPLt5mnAT6NlmVP
YZz2rh+0DGOk0bKscOCLR41QpJz3Swz3xfRvdF+DVKXep6LfKpEmcyoxlpeDN527
ed1YYx64HqjQdKo+8x1DPTv/XDn+yDV49p8US+AuaBw50K/utlk4/frnhUJqukP8
6zLHFyigjw5BWbeczioPHms9/oQfgPH/KQe2oFhgsjwdkCDRrcokKItxuYJ+UVbU
uOAgFcjcAiM0q1IcwgW7sGJ3lowC83cugoV9gj0S5fASiSSeji4r9UFwVw0dqL2R
esuJzf2DGA1BUSaxjPb72mOCWJMoZyB0pSSmx4ANTA30F8+DeRUKXOU6d+471YR3
F2GChRrayfO0C0/sGCA7Rb1wu2FjbJvAqf9Z2MRDDxzmxYlwvOaGbJeWMhJPYotG
bvRuJw/xpVfhVFqtWlz7ReGQQ4S6x/ZdDl92tC6Ow/70Mib4t+lIwgtY9SPDijos
JqmpMOyhVWhUgNkqwna2IqcacHlsGwuivtLuZWWUoGSh7WUMTTIEIh2KUFchPZcv
L8MDsguN6MiAU2fpqdd+7VhZzAM6+Nb92V4dYMypldLhTkBe3SpNn/WnCwSZvVFI
mY0i91AMs4ghaIKwlmJLjyBMZ54mH0zDZ4nXwqZduTx3wU6VdYWkt8PdN1KDE4AM
nU3QY7zpqnVcVqg0veUMcHxOUPkRX88MY1/iQTXnIP0bZDm3y7ra7xTdqtmcK+GX
+G5NcCrT7MfR8hWAlH5Qs5sZWNVPBmbIKfI44eusnTRjt2cuHmyjkvg31Vx42JD+
KNiIK9lRL0BJT0/1faPT+zH3QGMs//92z56fobMfO7CWeNofLexSTjPf0SEMp+qU
BW8krUtY0QISPwthvsrWA1UbdKJF9LWjLnk8TPiAz7dYZJZhN0nNavxoOybXzPQd
vtQpyk6QJqgKpxv5lfBNAOukpv6Y+FM2iEjqU4dU7KLPGxk6qaoYR6ilb/QDMEIX
uziEfhZp6pdmawqxhCgDHdZ2OS17iinJ7LVeSFMgQVDCoQawVTI3w1T05SD36JFU
QSren0qrk8YSJ9AQn5g3xuFofIZvuhB5yKT3sccKFF9FsjWttyWTBSc/YL24Q7PY
RjpJbvIEWmpJkdwPCqsDOJRebtwoUNWZplJzteAdMVDT8ehGPpsykncNgRb1W7K9
RjQOejg74WX0tzN5R722U4KzXKSBvyO7xXlamcXGMruNEQIhQgrSM/14i/MnFrb1
jH+FO/xrjzQkt2CWlquU00Xs8sSKtiqxL4CkBtALZ8qGyX9oWxYcI6BrYGgkYifV
8l+6xLFteAGhU7fQ9c/ggoaShkkrd8EEM4C1i7g2Z61cCTcXl8PI+6xyEVHf50Hr
u0PdRnCvFbArlZTvwUYSoZk7O6fO0pD+aTsjA63+wPnh395pICEa0cUskBX1T6ZU
KHiiC6DAOcGLP8hn4lAIfK92Bc4S1PLZGmktB0tr/WM8jmaLbKhpGOWdxvzfCpgU
SaBY/+/8yMLRZo2vWO7VvMjZYN38L9QAZzhQ9aJ202KQPsKrtf/29hOZX9v2YyPj
MtbZA9vKxXvX1Y5UuyAIWQeeVEyQewp07thOTJE6xmhfdR+UPjd36nuolZLbUheY
KzpdTQFIZK5zkj+R6lutnLqgq91+vDbd1PpnaXL9M69U50O4gVHC2qdD76npmhXv
yUeKVGanxShfqg0bQCH7+WRcQl0eRQmPKQjL5+QlxWDwhAp0zQHIIVSg5g1xzATI
qsXRgB66WhgCScCYC/VCB8Rm2mz1JskHn2I8myu0268DzokY4zeqThGJO7BrcG74
INsR+uVStqCBa5H4auRRYdd/U03cUFdZDklJiHmqv4KbnNPc1XxGDBCUXUpDGuHv
a4RejIyyNNZ4+xWzNy6JgwU/dI08CRMISFCv/sXlTN/DlMNyQ41gT6R0EywcZlEc
moZkz921Gpbz5+Xdni62gBo3/ljtoyzl2/4JG+lNQP5QbK+U6yUFjksoje1gYjx+
4GA8QBXnje8N4oiO4rAStTH/JDcEbvKzuJLoaOMb1mwnl8z2eza4NCOo0/lPm4AZ
DsTVt2sTzLhpA/NbpSAEpaFKwER+LDGWno0lBeWwT7RbdQvjc4S98J7dtm95Puqx
T6zVPjl02Kqdf63THRYhXjUF/v0xOdHXGUPhvbFvjnP/DoksD2yLP8TZxIN6Xfht
KDMziGuUBJBIBd3f2+5sgWEzrMwOmO06wy8QATNlPzKiMat1xTL44yHUqBEL1yNF
QPLZK0PZ0v/Zk+Lzo6woh66JQdeReZqR83HNCKCyLDG9KN9wfUKmYOLFjj5Lp0Il
5b89RDmZOWMqyV+NbhFcNYsBOMdScEQclvaSAgWKyWKPl4Lqzj1vD9EVZLwQ35T+
dn0yuUyuSFALvAzzt8Qk/O6nvbBnYOMe2bLeLD+Sv+oUzdIqRpNBLqaekwsfBWcv
pb8SecNS+FnBPSljnOSwDKQ2kBecTdA8dnscMjf38e2emtvTzyhq+p3zWkePtumS
JcgxS9/kvmwK0Y2T90uDlR3knYuJTLiu0A7tXqTUbgv9Ud1p4WT7SaHsVlNz7UvU
QSbDLmaKWrLmXIkdeMkH+A/RDbBskb+gPlkl43KaWUWXtQohHSJolchHqTbK44wc
Ddpjvf4vl6/jNi4d/EBBlULGtzOcBZbl/t3o0i0nTBHohi7sHZBdymJYJTN6pH47
Lc4F0M2u9VZTlWVSLGZSyNrxb3tErtYXaAKRmLNCIYZo1Ftlrnxlmu2MvQX3zttb
VJ5SOiQR29GhDTljbpK40wRBZ62CU/iZZzjXZ08vm3Q/POIhLOhBh0pdGGOZk76S
2w7VrxNiucuxWpvyBR6v1eN2QFUg4+6AiAYAi48zz/4R2/hVwiIUDHcpH07luMXV
FHYbya1wHutdJe7UzS/MeZZRygmPYFu40rHOKQQL5mqPysIuX/O3OxuFAsTsJ83C
xDfZu8d7uimmos67DMKjrFS8729LV9xqAFLibAL9hsjnJ2uSaDBsEnOxuU9T7Sy5
UEb8ZHqsPqwJw9pCeJltyRvOHawQGFNeheXvgFPurR3NNHTwdVLGnuhmGh9DLjM6
4PA8FLmDKN0Aa9LFAieZVeSkuZvVuqRgCch6l0qoujvsdqjHoGislKWu/NCumEe3
P2WFi0fKS77JWNqUVpUPGHOmGDfE3l16dnsivNR/as8DlMah5C0l0H+YMlM2P/cu
i8eh7/dHgiLzROWr9Kt3IVf2DaxetKNdnkVbqk88mGpR5N3btgAkzr4pFXUlKTCv
dasxxRIAescz/Bz/cUyTxZwrkKy1InySU0k9DXHFkTlKHIC0GwEiNF2yzc1JQZa9
0rfizu/KkN4CSa0Fv9PQrd6QGNR5kzoHZaIAzWyhmsetiOo5UonodfBffurlC17E
SkkbpcX7ci6ATkZvmM9Np13h/LPO8Rc4xg9727HPtQl1VMepAOLZvoHM61jcZnx/
fsz1sR86wo/sRgPIVbC7yCDuthMIeFRwhuHOUsyntOXUjEV1oPufW9OPhC56PH5S
P3/MxZxHbaHFHvsbIRowa3Pe+eO6DD4Q47YgAukImDrlM3A2+3PIxkNBVl4Dzr50
TUtfL0iPgtlg4jgqZ8woa5mgNIm3hgfz0G/XaChoLoidCtvfjeQXiYuoGbPgN25U
p7VEpnnuyr3l3yS5HQsU3XwpDcp528CXU0R++40WTKSZ+gdWMsmWQS56SN3M+/ND
/GRxvEua0kfD6pVqaCn0ajPw6zy5Gvivseor3zoascAqblH24ubdA2nLc3R97T80
9g43PrdZvWcSUMfI4BP/WVxqyzWTY7e7X93T9L1z+kLz5fPHoXvaPv/ACqjsWneo
dy0BuSVc/gmPd1pW0BaSzroAr2zdEGkZ08KvnopRTWfjGe+5huDWY37DIRlpxrSE
K+WluonNo86QNifj7wVfUvYWKkPcfv+4ekd+gl5nheYZC1yQ83IT1SyjtXBwTBM6
sX/WOseNkg3DNlbdggLpU2gFSeYLnbp3GGq2WCF1bh3tiZLWgslZGMUN5gA9LxR/
5YUV7Symvl84TulocE+jhOruMA9WMxspO9dq93bCjhakDZu8BZJhm6DVdEQASFa3
dSKts/waYdPHqqSCclrTUpKrgkHHq5cyqkHcQQHHEEg/o3DcqbgWzw4C1Z1s6TDK
lo5Yu029s9wtJFFttGiEM1EMcQyrH3UPZPPkDn0UOUCvgO8JH7/c8juIAI2swnbn
n9hS4UF7lFOBwAAWyHwGRNi6fFy7aQyq41Bx+nmH/tn2VCCSHiIeOSGGUxtvBAsU
H+32Xxgni2qilbatVDaNJ8qxxsGoBAmsrG3ZTUX5Geq1FNeBmpHkgQaF1t6rGmD1
sWHOiYlax+edJKlXTG/4pcqIzYRVT6DJk0+7Yrs7Zi2sHw7iG7D8cD1YheVwnxOY
3SghmF4UMIsWYz5i+ncKFrdYER19xufR5Ah1ZUsrxk1rJTbzB1Znz1eKh9pfBGMW
8Kil2XBtI9pwdymUIsrYoFt9X91FwPNAzj9l3S2esfa3X8E+MsteFJFuv4wYj0Zq
NbXrT9byWxt/nsqt0IC3PGZB6hoWtEqcs8lkkPwfzL4UpjJbphARps7yQgDoJDH6
XM85nvHw4tV7vgSRxEiwAvCho25xn4CFU/tULG+lolCL31bS+M80Wd61/g/xcljp
c69Z0PZ5o13scK1Wp1J8SJFqsKAJrIMsiqV8oGwFcBE3zkIObckEkPrQxJjcxtsk
fyEdI+UJiU0j98DaVMhe//WxcNYyIxmjPlZI4vItNuWR7tPWoSta1U/tw1fJZyYM
T8r6XbnGnMNqT2DEoHR1Idc3tgydOkXr31CWXX/6d7d48S2UmAc3/Y16AjT/jo5J
q8sNbwAg66PR7ZplAu0hhp3wUvnc/9QBBo2RGH2hkfsuBi2dRVGa9h6iSgl9l6Gl
PMuJK9sDhDCkRb1CuJ76WHJaB+3468YrWEGkCHBDitO+rqB2yN8N548qqqhkY+XP
XMrg7JA+rsW3OLGR7Gi8dhkT/CyLuzYkNjao0lSg+LTtK+fDSwDOq4RIZrwdPfzv
5H1Kica11ekYTkx6LSeHLE/CcUllFaIKuxfa3baqODR9y185nKDSK1wWncVy60CH
45+aat50kLmRqnvCOYjKJcriX1gUP/xYaMYbiP8SyvX+8JEWgqOlmQDfv/io+T92
UsseRm/V0I1HD2p0hP/QrgmgSdonyT+CX3Y/2zNIbP2reDyYBvJUFGrsRwL+BL1B
gBm+9LDcyakkApFsCaTyFhQgC2GbvyGGjGrccc4XlBH+JIxT5gwntqBNdhJE/Lyj
PDXZ9BP8tXaa3iLPvGovAfKbs2EP5mPEuD8VPYMJbYwburYymOzWnjzCjZkl/IiJ
cWSg0fipGLat3t9l8f6zPTYxl/GvESyRGnEkVwH4xKxLUgseIcDz8p6+hc9mSMLP
80/Yngg7tP/sEvePpM/q+uWt5pWgrXYuzJbEHZAzEh96fxuH7JW1q0fb8OVcomnS
3b32KhuJ4H6IndIgc5pD3tqrBhv9Crov1lKVeqO7g1KY0tctTtAT1jUOaIY4L4cd
LgFNxyDrQcGDRqX/jOGJO7sBzZHRJxTE+96UmHG5sN0St4jZgauxLk+zH7e5dw8C
UvVEp6JE9uUwLcThYvNa8hdwcbDXxgYAgX3qIbbPYxKQjgCPCml89PSEd6Nu+yFr
k3oyAHWsNz/umLoXVSg41i1zXSFRVjiDf63GrIOHe7X5MTSKm37BJ6rh2qtkSeXw
3OFaogqA27uuv7vcki4zAfkooxEE46r9xZRtxIlCW/Lq0wrMOW+U6yEt1x/2J2KQ
zc0kcV36gMehVYnsRQGkfHIhbPvrDHmW8r1cMZf7SzhwBCfmURNvCDdlnCGivvOM
Xqkwp6Grx4NFNHPGUApuIAP+ouF+OP+QOUHCBaLGq3lolABlPECVG1kOFq+aLTfr
vhtvyKXhHRm7pEUO22IxBmEENzNWHRvaHcK6oJHBTXVkONOGXY0DoxRu85DZCRpN
xLXk9YcRkJWUhmP1ih+XuMDhQdiDe/IcyT4kQ0ARdAOxmWgTHJ2WQnGjhPJ4R8Pa
bO2SeIJkuNrZ5SuyIAWrIFnEN6LE4PCKam3WYdeoemEriuaBLNb4k7iZ+F2jsHPo
RgkDDsP3psgjNVY0XPDGi2Uv7EHNGA0iotibFSwOUUTsrE2Z+dxy0DMClz4s5PSF
9H+HBHsCBQWtMuyNfRw6LolaAkaRqmbuveMTXb3GtF9+h3LO8AhwrcUjH/eTA0Wh
vVd49nIun8XQyUvUNxSPan2cSWaqdlQBFK2UyNHXqWSlXh/oP7Zqpo6663Gdwuey
/DXOSkMqqX9F+Bh9LlRTtI5EX4allh9LIBtMeBTaSIorA5NpK1jR7q8kkM/fGSDZ
i7BUVug9327J0zMYT6kuORIMNADP/iZh0gtNriEw7LdOmPmpqGYcHmERoeZ5jR2W
LKgD0rbrvFqiNYqX9xxZCD414M6/KmKsFf6F4FACGoUaOfpCcV49iTW5ZdgcHvGG
IxPV7FyzahyFBrUNQrr/u+mu3gGgGJ4ZOCrv5yR6NDtjMVlfpWDVls3fQgma0UQd
DA0JlwMhtMIZw0Qk2BvXHY5U9I/2PtDRHCH829PkMIZcmsY6cYPqOmKFfRl2Gkry
TKj9XvuUEGmJSRYDweIW6Ytv5kpVB4JY8Z3MP8R8S1Yut9ISUlv4HonAzhnvXrSa
k64lgq5VppGe+9YneXqHSOW55kW6e9E6Cw8kDt4HyB04h2/sroi9cXXCEEbc5NDR
GMawRi0o6x98BsGJerr7aO+/ifd3wn5nhde7CU0T0PVpPIppQmJa7MWc2BYiDACT
FoRLemmevPHlLhw2c0WuPUa1Bd31HjAzKCMBgzADTHuba4nWc7j+NN0qj3TAHbU5
/MB5+6gkgOKlgKYLVHvTuqgdfkcsSi/EHbQx4SZgm+Jj+nW+KaaqcJcEE0YTBjJb
EVPlnt4DT/9MWJ8mvizKxnGJaLjOWNABmgUHcysrYt0hBFSOq83djsRH6Q9ivx6x
ZrzncHfbNv4ysdojn7qNRY+hc17E1L8Pfz4ngKcEhK9QeG4JrNITULd4Dn8U5lhp
OAeg7IF/UQkK+c/wa09mjjyp9/yq9xcf3EuC1y8795rYbrqs6R1YVPilqqx2DqxW
pE8OmYRaksXmHgETGNm8pGTkwZ/uG+p3wXgWWNad25FQrSx5nPwBdsk4TZPp7+kU
wx87swDMPywijOwcVA+Y18QSJQUC4+QxW8rojN6/DHP5nBnhGhUHEJPAKfKdQ71I
r9vzwf0DVMBLBwl8qIJ1dqPxDfLbqMu+Dkt42oCnRU8zlbUNLv8HP6uJLN402NDK
r1SZOZ3du4M3BcQH4EdVE1SxzUtaQpyP+lWRIJygpc1NZ633wwW1YHRKeVu3k8B9
2GqXsvNZA94S2uhAUTHYCcpQBJXeo39ZubpI2Bz/Is42sUP79uSN72nc0ijDRxEM
7S4RxGpZZpI6oSEOtJ6/tsc7Q4Jqru5UQD2YsWsBviBPEyFWkmieggMZaRwSSSuQ
PE/tzqLCtc3v03hw1pfxFIJ0hMmiuHnOY3dCPyfg8Ny/+h6RuI6eQk6OJaB0h0xt
7AAccwLq1/u7m1gpwSa6MzMPsPvwOWeYFJhPd2ONIQ53E90jJqNzt1ciH09u1k7z
tOrR4+OfTLHIjtAvNmESAKZc1aCxZG2Z9kuzBNVeHX2emaKeGr0o45f9+ltTXNg0
k8lJyTj9VvY5tKDTFmfLM9z/oUcrIXpsE+fCnzUdihm1H9cwtJuGU8s/r7W26ifZ
1mEcGmFSiy+iz8Ord+xZ1fLbGzb7YcDqRQA8vecYBiCqUek0SyG5D8cFsY38ydHI
/mFSbPbywj7z2GpvVRGpTvljIO3yvF0zpojAZtOOD9J4HG87GyPtjQ1LFwZ9z7nb
SLrgMTDKY8lETf4hilqg/h5BVNvzKG9HJ2b0H7MO8CJHAOo20xuAs1cpl8Ap/fdK
2nmARxfjizqCdQF8nkNOg9x735qeCup/hTcHCUAFkQJvG17D0hLRXqjqjJowgh3w
g82zu5nzYjTigxnNUkEMCapygInKcIdvoQK6hMq1KPCEvwPNCCA9Rwi6PrAddZY3
qrqvDSA0Yj5CJvyguqZcfkxOByvr638LMl11jhzeixGxXT5YAdJUoceIDYzisVfQ
crV5874PwGenxxR0sBLSnDykXYgP4KORmLvmAHjkGBIQ547wuQ8l3hFJy2o5fFi8
6P40Wuq7hHLYeA3pj/aLYZfWkuA9D/2nKE9YLUDRO0mQq8JWEqLQyrotx6YPwwjJ
jDDoDqEPCZ00GFHPAzt9oueDrT0kIKHzd5HFXay8uVmpNUNH2MpYh4jaGlwWf8HN
IotsWi/4s7nVkvMlKMidb5grpSWEWqLEivhyel+3w8rU8k3hC7hdVnPspRJA0Ys3
AR+yqGfaSYTZKqYp7oxVygHsjZy2gUyuMvC6aYs/h4RUpfeGtFMLT0hrulEC95qC
VeN5lxsg8ZTLS+EhAb3UJhOVxyx8rXJkOqmhTo4xMAB5MLU9tjRZsd1ryyWq4Nhf
qb/02IWzWRgwdph2GmpqZ1QV8x1WHFv5nGmvg/iYYlyu6xDvbcsZ923aL6kOiEgC
nq0x2nh2G0P6bsiPP31h5trYjcPbBup6xyNUR0WrFJZ2FNC2N0t2dBlwb5Fj/0k5
9CZesT8pfAoimzMO0zkjRzLiQPmPR/ibOwvT1n8wvnT9jwGCS9aYZLs2mxERTC7R
uUOBan1kc1LeDZGEOvFS9yYZpmWngI/fWkcMTx7zFbCY2EZj23pGAqllGLn7ufAs
j2z4Zw2hOlXLP5X1V5zbLFkHo921SRsOjyTC32KVMzGdTOtObY8Yw6ZeDhbClDfY
cpyL+77G8YJuQXR1iNuJS0kM5Qsmh3qCz4zIa5Ca5YNs5zDWC/LqIgyDCH84He84
+4Mn3SLndxwfdu6NVEPkYx7sMEjURvjfxKrZVqf0/ywDyc7gP+S5hc6hipAb6q1v
aSZ5MUbP7IXpB7ScT+/YAR5JMOTg3iKj3aX4TSBCUbmOeAtrW8h65c463j+UeLxL
jehlu/JXvYVc6AH2Gtt4jB2SsxM/8AiwBPjl+4x58glLboQhdJ5bSVCaCEhdR9sn
dZVWHSp2wEFcY22STv8CgtDCfqHs4GV1Mua5dHbqaRj4l+qln63AsISX+/b8IzB/
lM6uEM0a7/BpL+Oy0rKhLGUE8uRU2HEj/ag4TTKyLd+Lnp9qsGdezU1CFR3qCrLr
ROmQYdDEd23zNx4xAR+HH4xu8fp2kAGxxG+BMe84r6F8aa2I8ZH6pyg/sJbC1RRb
cJ4Uj0i3AFZP0J4lDjTb7i2C2YwKBr5LSKhG5kHNP+4W8PQdpQuf99jUAWPNYy9N
sY7SOnrKrsWzOnXoe+I57P8cTTMLczTjuqw7aUPV90dvP67EpIMdLCaFfRdC2AC0
SwwiVbmkKFKmf+cqskKzYM/FRWaL624hB+0UGfJPjSjpzzPAL5HhoMrGUs77SfC4
piuaElO5OVLlz1bHUbWtjP27sxTY6OEqaORb/6qUtXFgGB7zhOb7my9eF1g5RtCT
rDHGEiUw4wZxrU2iUC49ixs9F7LNw3wpgOC/D+LLc03ZeEkVs450gmHGXom8W5wW
V33AG0b0+a6ygOpd/pGv9ue2m9hRSLPZdL6nsIpW4epKurrP2F9WMTUQ/g1a3Oly
VzEozEGHIz2wjkN0dPhe8D7DcDjxeqBpRQdXHpi7vzZ+zf3HB9ey73g+a9gGdwoB
FqbFIUxwrqtz2xnIpVUwjcACwAA8N+6FkKNG549ivWwNUHURON520bKd3gNf/nsr
ozGum4mSDD0h2NcsD45HQjDGapZbi2P5SdBaYSP+/LsFf90Uhsv5ShMGxgnPGrA9
4060iWsTGviJuZis4rdXIzM0FG78Xw8CyivobGDsxcdz7kYgxzdGHKrOHOF3qheE
WIa+ka9G99OPNRCdF8SGcAw8ZoZmXtnGztsYjS4XV3RkKGUMwwKJaL0yp2jloCKg
xhMtUE5HcKwgigTlTYtMmMb70Xm9LFKEhU1yL3f1jixQerZqJk7rhWOfb+J0LiVc
qM/R8KpE1+y7zXZBZbbnfwX1w/14d32oo9x94DEAI5QfVIKQ1OiW6PMafle9o5Eh
B+OCaMAgGyPdDlPpuU5Cq+sWrQuxF9j0l31WnnTijpr++lErDap4WPwRUjYGa6JG
7kAI8cUfgl9J/qrD070ulJyQJzciTRl+TVtZ1cyhhySYkg+nDWXt4z2PRRjCfzh2
oXL0Zyt26j07ClcCzS519Z+jnL0UwqDOBMN9ezxSSUnN7BCkNoMtn6jgMtwcMyDl
jeqn4Kwp7W01XCMu9DYzbeDBfat8hmHmlVOUH0KdHMqDZQJktrCtiK+pwkcdg1MR
pQtEY9z8dQKXeCp3p0S1VdYaOoAayrX8XYHUIM0arEAhuFeFtN7HbYsgNL9ulnGU
pkEXwMGfBmA8+LxkLMt2SmHRBJTrh2g0IjM7QlXLF04y63jLdw77OJSgR4H8zeCr
8fYGuRftnkTvE3A5vLv73MIzoxSRlMrkSAEZp2PidEqR+mpt4960c32hQxpyTdTZ
xyyCNc17//ehWpFBiKsVUGX0LQod2CEtT5fYam3Vtg95sq2A5/i7PvNQl1ASttwr
po3ONbHBmbuNtfcZNZWparWQuk+y0Yz71KpuFJER4VsgEMPQMJM8So/ve1kEws0d
N/xK5hCRZ7AO1LtyrCJs0SO30RIO1uhDRzyRE7SnFnrKhSJIa4P2e3jJQ3J8BTMk
aC2GmITFFj1+Gdv6GsxywSVlZdvbfVBItdMocFdF80HUnbyBpH7TYRzpvppElo67
17yRDJNBNIYMjdfj6WfmA/orswm7lKw50V9RqplOw9Qca8Ti4urJmgWIkYzihRc3
59fxaHODL+LcYFQs6es6w+5IVRVlyebS2JbRnccrdCFOWGorZYFMnV3dcvnSgDEO
dZ016euSOcpMV3Uom1L26BWZqeRK0dz518qhwHaQKwCruNfcCYvFOBl0yh+YRb5V
QOBo4A3RmKwqQ4ALOWYal1t8RGPw9JYgsx/UZsnYQtuReV8nkZlgRaiIMrjbeV1h
AG4/k1Urp39ktY94Pk6u0fix72fD3xwtw+k+YVde6GQMzWM3KEQt5MG0qonimefq
yXljTgQqtPtlolhkHDUX93lseyDSOoMpdH0sU6LPZ63YjS7tC1ixSIueOofpq+hS
GgrHeWfyJobbarx/+6AgPXMM/6OAN/H/PzT4lqh78CsLBy+PixIRqoHKGw78/mkH
H+vzPzJ2pRHhNUCE9qe4hQ2f7P+AnVAzM5CI/+/7dxTIcfEH06X9bhMCTBRVXRdY
xxyCa/zYUbRiw7L9yEfcnCZuhTQd1VKJ9da1XKCVmTfL7ymWPA+Ccc62dGoSnho5
bdjLKfDWEIIUA6Q7Rh4QzLf3BWX3FXA+iRD1dFqy/AkNRlGtncCa1UC8e7quW5c0
Gxg7GXxrqYdebcUgMoAs77rT7vFUQuF7juGd2fQZzM4kRAWFKsMp+ZCai09INjpY
FbIxUubSzeCFLN7nsC4KdbJbWDnICHuADxvKEZ0xw0Yigq4dY4YTxIEwdF3w4Ev1
/xBhIVO8Ezj0ZDTgLGhV1qRy30CR29iWQf++SiPgCp6Tc3je8YnoAl6qJRohMGt6
52EWfzxRl69WHMQGs3tZqFCn8c0FhNgXk5O9nGxzddKaZ4jUF4zl4YxVE7orXzz/
S5SQBAlQSZ2CxHXClg0EF21n6p5Y4JXwT0cNrHNq1NFM+RFxZwBvzk8K1vhugPWk
CFEHbejel7vtEchixCvXfXJdv6EeftaItOTmMWT2MfkKJHx7aDu3glO6HhzeCOQ2
uCZsmtt5x6tBCyiTzEG7BZGa3c8Bu3zQErjj9x6TOButXGp8OOvI28GmpaLnRrHw
IbGmxFLRsDDFGhyZ5HoJml73vejbrDWg4VvnraESWRSlV3hyQbhXjOJRZfdmri04
mpHTQmfB/EUMSNp3m66rHgXbaMHX+crhJJRzm12XWDWrjQg9uyf8XxRg5okb5vXs
02ayJiPE5BydnGhyDwa5Qof9vQGpPneTKp5wBaYJMnIAN/KxYU5b1lmOicHXzM4B
RV8jVPvu08Qon5zLndMtkZRQF6bBrovWSn7LBjJUeOdrFicBgs5M7i1Y+waOso44
UM825Y/UzzwEvPro+qMZE24Ew7o617iYEffbPfaIpxiaQk2Cj94MlvbQo2S7sq/2
G48dcg0cgcrnAuowwQMLvATCjjRTuSK29ofoHfmOYIH31Ms9l3VFmaVQVmq571Nk
oksazcY//6msQQaM9BdUXlERdn1xzDHF+MqyyY65D+k724hP2r2DYcqxRu7Jfd8U
F8GwIa6+ElGojsxa8YRYx3esdEn0LJRovik2ypifs2oeC0XRh5S/Xsq9HKQWwIel
aN2f6i3tNTH76AhQIcIyGVoVh/KWT3mjLz9lKiTrmLAjVFt/G7WVXt60lW4xOlUb
kuO6Ol3li28o8G0l8ANsEUrUbPHiNS2tZsY/JeGVFd8YllFUvHHIRkwpH5qp7lzQ
5kEXCydF9UnPxJEgUsQP2mZxiKfa0TMw80eRyJIKTr5lWgQlcHnDu67KZy9HnsjQ
Vg8lxgDqexfGNJADlYsxO1sGOb7uocFCjDVA67IVdRKHiT0Wlh+KxOAJ0sRRDz35
0cOALfDIgHYhnAVengFLjt+FcGZXtK6l5CZ1U1pt9gh1dsG00Iq923Z357ijDvgD
GqYIrl3ARr4HAYAsi6I3X72dHfc2J4HBYPs5krN8vo7hKum1MYVmSPtoZ75czV2K
7dXuE8FwuUlM6apPGYXK+mJx5bEzsdrNGlTpN5sVllvfD2TO2zwQL0CvP1K9qDnS
1kynTwqlZocB8EwnrYXH2new3XSdzqXbunzWmuG0dSS7+u6k/sW8HDkzSLopFXnJ
blCnSWiBxDVPoFg41bga5WtBGcEnqQe3WuejT4hq6EmabBYEG//7nMFeDT6mr0Uk
9MPwMUZccg5uYhPOW0HEtgHK1n6Ez6JD1Z4B09uMPLBzxKN6tAZThW4BnEObadCe
JqIPWUEfCo5r4YQD5t/ZVz+ZPF8kXQoW0P8k2WXgIU5S2e0fY+OXlWeBzM1bcedM
hnDOywBDtzIBocnnVTLnUtfZPUBbcZHzK9WrdZhg2A1z0lj5gy8/kawCbm85SkJQ
Lcn9S0vA/4RNRXUZAA3/rVOVgezAf1fejdyLWHUufD5q02/g1Eey/HWQ1SLkQRjW
+1MozGHE7p2eI1dZdfPcBdFhD6fLYdwXPI5Pxvosqg5oXE4qpZNhigsBSRnoKGbl
h3tWXqMVcJ4sloPodTvRpGiZUfm7379RFfE1a2RUdCfXNnDfuoOXZpffU5isSNQY
UfDAhEvLGy7Zr1z25IqV/b6ElIkF1dzDyFZPveL2OmEb3mKI3DqAnHk8g/gbsGQk
ZHlb9LplM14UsMja+smknQHsWXqzu7NrctrnvSabfFHHFmPBDW+2sl5nNgYGddwU
dXQK2FMM+EbtoHcWmo8alFNqZu5j+SoU52wSZ9w6YEfdHgtgFwb4oOPfC0vmnP23
vTmIyxfvFJRHHEpHYuLg92El+EcC/OAbqwjJCxE7O8lZqEmOd8zvRge1Dj+GjWMu
AyDssLm+lvJfxxxvodhwuClin5vgNcfM//it3ui6nUDw7vjgiGLetT0hrkf1xrcF
tLPTLqPASesgZg2y2mLmV5GnWyRQEH4Y/f/PY4uQfQNvXp8+qkFAUorpeL9TMZlN
b6FbcDmuxf2BlI8tOhkuDwt0JPHN/b0LN8DxW0gI4CmOr4QJjrOxT5rW9DXHkZmo
AWcCT+4yboYetZBk2EdQR9al1VSx62snVv3Txk8EK/jgw42iRQMjvhkokZU82TJr
Yuh7cBrsJYl4YwNUJ/wX+X/ozO7ckHf9hjxaNOfdojk0E4hDxelj+YORq+oQpuAH
S/5IjiLAds/7BHQsPGhorYweNsgpuA5yo01crVj9I3YMAjO8/NtncaBedHImDuyk
AaFuYHJAS3S4HELPLfNhRfg5tWQXxNouTf88nXryCQo+6Yr9o9C8TvmOD/CKfzKy
zxe1YpwNXbB1Dp8mrzNzcv/gzxluPKSmYheZMH3bLBGQmDioK2tIuHNtyhof/kI8
kRzwsylWDf9RbmAYVP4UQoUClNAeyabnLzc77QWaC7bgnnKuTwz/0ymyKLtP8r7H
a0MUuQHPML0rBB3iuyToD+vnUNEULox8pXZ+HqP+fIRqNGVAgFpYX7JnhFLILl1z
/nWvnaYn//KkkNEk/Re9nEDwlKRzAeUj7YuMH2b2e7/614wHAyi/KzLV/3bWZ6vC
Ir8/Yls8BOSxcrhr/admCGgfQq/3cmCM+iUrvzW5AOyK5R+ZrzAa40MZez0+Zo9+
iSBFwfHcMTtZpPhfOnNkqGPK3/Qhh1PJn4NEuNxKyDWiIf2i141/Tt/1fdupU9aS
Epw2BemlYCw2O/6r/fJlBoHcdUrK0Wr4EcIOJfMHaBNMZ0GiW/yoQLM50XI1UAjB
pyuZTsT13rPM+ULdEdR3rTQ6Y3LtBtSQhmNxEjGBzwaW4YKWc5YT+KO5hscEqdbU
034RhKicwuPOWLshRmg7o+0H7r2ruYy0UuRS1FQD4uQXu1AM/2Pzpv74P8RTqiIX
44qujUxqOst5uiPgX3feqt4tr7mV1u3xKF/cyZoV9jUabks4S3cThBOsvX1fscXK
LpnWWNmUtxYKLqXxe9KfdUVq8/ypoAT4W+5sMfCuD9JXJobxSqWKdB2CVWoZ4zcm
xMv5EAjkNHE/l6mPOCYrg+LKnU6H0v3TkdHQCHTxMqr2y3MTrUNb68Cgo1pUZfew
kCFW3iebdVCpcrxPQZNO3QzRy2JnQffoHT5fHUk3itVFPojm/yowf2zAjcQHoGSW
pxeEXAEpz1CRDVVpEQyWgmu4+/zYwIAirXdWx5HkHyJdIV0SyHHxkzwNOnQryLjY
WAL+WxP73UNGvNwwLjNsa3zzyBPFU+O4vo0qb04Zp7+cuLdB5IX8r+F/rO3hbz/R
0XpUtnoizRNJ+rPm6zuv9CRKEbhlc5O03F2pKPYR2wZhJ5LpPs8SgzD/CCYUJdDY
R/muZUH5jYQvesbODXdeiGWi/TEeoazYva/pYyTF9+mpy3yv2R8lb6Tc2rGnxsuh
e4y3Poai0Bqy/+8uSFUqL/JMf+2Cxxz3h7iahG1qHHwRDMN1lctj+XUUFLkr7VJU
g6VGXstTtzuCfd65r1q+u4s9xGkeOV11q7mbRaSLeSyQKWDgSStbTWDkMCebddN4
mdTqg5rGUnKMTq0jUxMGYumekVzsvd8PwafJ77L99f9CHgsPBWHUvYh2fpcD5CKr
vS4Px8rFXeeik2D6AdE3HQ/rYYFuM8Xz3Uq/kHkdJEzrr5+bMvt0HzFjR5QBkAS8
2hAzPCzjvzZxSf6zkQRfR8vNomQm+NqLdc/+u5qE5j9f4P8n3X6LjSKFBYAGvdna
6zl+DOKGzvWwIqkNUPFgKRfEeqNffWyPZWSJ7a7YXYbz4yLe+TLJH2O6T4fr1OIE
un+9z1XaX3n8a8sudnVuZ07oFiWvbunFEpHGXq2iLvOXtHVliCoMItV9+wxSe0qH
96oqiEkcJs+t2qzPxtz+VcWKXuO8Q+toSqbt8Z0vR8btL3BIpTF1HqixASU+RTs5
YZgntcbBnQDd/JSOiWmktGzEBlGwPlEGoBpJQS6jUmN0pl5X4GI4M/5tJOaXxQt+
pkRUUPn8VBuxMZKVWP5Iz9dgGT1Q++cgchq6R20u90sva7ysz/0Z/e1hCAJq7xG/
Hvttur4KrJAx5QR16kml1wF1BrzgeI8c78IkcHNYGibSxZwhfAApI7dynvPxl4Ef
Kqii3H4gmXSi8ALkIAnNnsUrZY/kstsk2UGbill3rzIaZbyFScWix1QQ1UUYSE4v
RyRoKYQMyfVTn3tSh/sTTUJE/P1/nfpjgWBjPJp2pzdNnq1V+RrQBBgrOzP312hE
lwlnpNRnXkjnjoVsx8AgBX+T++oc2AWEga2vyYm/C62yh1/VekRDeW2PPYnSxS3W
N8qoFusr3IYjRUSteykaPFFr9KPeNwsYIzzcyF2ErEVMbpTNCVLYSMNQikNDWRG8
7MM2X20+Q6lNXeoa8GwQpp928URfzUzW/ljyY2omBafPkOHKZ2zoli4GqRP06tDr
Q0mXPcmVPOSxxpAeFzXS06LoCQDMisrwsBgw0EHn3fKDfhq2IrX0G33oXFxZK+Ct
QjEV49UFXC5WSKOSaUxvb/SZ5kT+BLQnnuRTcBsA0XVVPkvPAwEZKfqYMXGjnkJv
R/6+udhb/eGm1PlUEV377YoMgILR7xsXp7CGW+G5w0FfGo1Tx09z69wymJpTXdi2
DfSOSVBz51kQwn2oBxB0A/+Ui1lxMxKW8+ImTe9L3TDuNa8Sy3GUBRaxetsJMmZn
szkola+q87+lGdnmalm6ylvgHbtqgG8iWfBY2FfnAKyMPektWthcbKUP7Hz8fkLt
hnUedwDlvzi8vbjTUQpCB6I/ETjhe1SoCtOPYaNAQUVgrNN0L7CntxszxXTl2Y0s
zGUEIRIHz3o+2hK5f2uVQKsz4Lhc6KzyXrDJSxM1n1Rnst11ZbPnvOXpKCCNMydF
gLu1nhP8bE67czikeNb/JzipsZT/VHPe6D3U2c5eL2XyydeouOhhSGB1PhCyFOa/
zIx9JMpdOlIlhfxhFx5vPekuLVG6WpgEKbfRMHEbHqabMZz0q6bNtHNCBN6qN9re
gNlcpRNcq8KD78NaDuEsCit9mL52LPEqitJbibi6j2w5/DP6Cla38Pgas1ThUJ8h
dmT5vNRiDW/0Nu+xiWfdDm6LFUDItG1dtrmTl8EoNVrD9kSke+Kg0haVb/EI2H8h
BjZY7kqfEiCoz7Puo4DQP3NHabK7+di7oBEvjBUnY9MKxOutwmE+PXDh+TATXfE6
qm6UvbOCFCIHwMSIvvh9Wex0FroH13eAQGXXcyeRJE1FvXzXlGuY835yfq1qKQ6I
qBRsSqO4MHP9l1Q8f0N8an+rV0rTumC4hVS4ismcphT0VF9RjPKzYPk5rwkAs5GR
4sXrB0oJYjyQrc7buAzR+1Bqb+nZ3mfuomk6AhWqXacR3HuFYD+mkadMHPcGy+Si
me/XACPJcQ4IK5pW3cdvdAleSFs9LEeQ59T7N0p0M8S2CHvjeIcrGEtPsMWYIuzi
Tb0BTULLhHOXJ9hYxtYYqYr8VTvvxsgaXgOjEpsP72kufDNsr++48wN5jh9pR0bt
NfNGchnodFA6ZPEokL5p5dkkENDabDk0rVDstgd1dTgjBiIt58eirbNAs3CFOe6C
sL/x3Eu8S1wBK0RIan7oa5d9LOg6UxZhDjazuz8/xJfDhpQ5fCINCpCwrne7gsmk
MZzmLQsijph0dDe7mZGvKyYtvQre8we8Ydp405dE3rGnSTLETCX8eD2HJKPLHaWM
Px+Y64ZzMwxX+WBNujbKank0nGzTGU8bTd3fnjqCvA0SQDexWjx3JrKPeIb4X7B+
wKk6Z8uq4NVow06xLrmELu9AMIIXgLHswNdSYyGAxxqfU03EsdKc0b7BkdkcfWx4
124BjnX/Znmg5Taq/A5eDFYXjzsJTbG8tPrTZNREgDlFikGk//sBCSD8tyQ7DErA
c7oveZzODFnAqL5tIHsYPOTWwhefvju3k2KMj5mw0YHqEvG4NauVYWBy4joPBPq3
FA1t5+PaTbJqt7OaZz8V/L7DeWSUXtwyv+u+O2tUgvoIoRhB3GHL9F2XPT6GOQQd
zxL6f/5rQPVN4y5Z2mAICdrxdUvIweOeXxsvxdRPJk+IIjqp/36dLwnKevWUGjvK
gMHu5lqozrtHHeXFoS2DilY+kcN2e7mxQG2TQebaSiYfzht02ZaxEYERAaNZgYr2
9cW3LxcYHF5SMGuhInFPqcR2CRfbOTZaX67RZxeN8VqLPgO1tkd2DJtr1QBed9HB
dkMFYBGCAXoFHBaOzO2Zr3y8MKBZrWN+jOVrMDGkwngW5myWCnf7myQNkCegTeYz
J6t85e78SaqHpWTC2opyrlTMXKsmDlWCvR/NkuAyXtfNAwTruYgaND4IUltl1vU3
PGlbhvuCVqYE0waJMZfsfp8uSOJdcaQqON3pSHqCUFYFNhNUrdm65bQRfIaqM3UW
SBFPysEY1meVeSfSDMEZWr7zYCkBpUucIt9uJ5uPa4SeE5oEkBTqnGuqj1cnw6EV
dJNa6hOtabUov9/kA1vYnaIABl4+uUXQJ0OnW88FEebi/b+g1a33tmsquKGO3ffz
jkK0gBndyo+isLMPO+I9x9RgNN8SPN8QmKn1L1mX5bOFwVEluwFIrkYu7aGlXPjl
P5g+BjJ5GDIqbfk7nQ/qejLi1utseZsVn19EARVmZPbwfC+sfy80YU0GxIwpxk6e
ME8lJfnhdyl0dXbezi9RyLrACd76uaYQFdGg6AwcV/MgnbiTFmyaI6TiJkvoEQDw
b9cg67kbi7XJquHC1jcHMN6mwfUmEKx2Roaxcgdpt7Z8DznuTXvp7OqjLkqf8AsW
5z3Z5Fr3vyRlNsD+1bdv6vGq8Pk3pxTLFjyAOiLctyW0DcG6MAGgmQgjCE3fZCI2
KoEFSvefiyG2Q9weIzEAlsXVeO665DNSg/LdYYWVfaMrInuTokHVnUqFp1J3fLwY
G05eIi/4h9GcxScy9B07VGiAhkWV3YApIZcJ1XUSdejf3r18mLHo15UjCsM5GhTk
FMOw2tD3ZZ/4hgWTFb+pGqzpEKoDR7ndYNKDtZ1Z5+AvndCAmlGoQ9PxwBJ+q4Uu
GBCB1kF4+HYzrD1zZZ0Wag7Xw0+paz3gJxXBVbUQDicYT3UIrjWGUq1taU0j8mhT
XY09n+ma34LODvCa/s4oWYtfofvLa3jm5Jp8U9gXvAS1zvQBk7UPGkpOh/sE/PtR
fWkt+Fm3aeaBIu4GuN8QNGRGN6DWrWG0mVuWffTYANoaDycJAIbAx1XO9qBAAZWh
LnjI6EAjrPYKrw/8hQbkncXbGRSsYgEyibSiTc8CtJ6epFAdU0mF28PaWWpS05UV
caenEHCH5f4Z541u86wjUd9DUMTu7vXTmkJLddazoWLX9o/3UkTwCpSadBRiYW8F
NbZLCA7uMfP63Zb7ECfCUcmEVb6lyZHh8821G2Xh1bgzjk1HY3EbPv/JVMg9vrxo
cdyMVTGzMd5EBZth03jsYYE/JKrpaJse9RdjNguhS4SJI+oRcg0FlSpz9OGoW0CM
BZOsLLFg05BmfnPzHSlRhIZVZL59R+UOyduGA4S3doPRIUfTbaZTDfpMqn2Fi7xR
Y59FuLPASllsyGKPNLBvMB8fxFi9w/mGIstX997cQ4RZj/aY+QkfCco/Rma86XtX
J/bI4ajitm56Bx+q+68Yk/iTapqfAbbIIsI2aAtlkPT8CgtIwGjqw54jfPz+drz1
+EEqQA9M6xuSr08p6S0MFTNuL2ccmhWKReK+HWUliPlNxsrd7/3cT7xQMSyHlefG
NUn17L6TEna2g4B+PajuML9Pif4cGfFtdHjjX5Nc21+rghM1iFKSE2aY3myEC44d
sx2+xf4CEYbLCQaBHSlGxfSELqpjCNBqwFwrbVA8NtLCA/IqqNRRTMA81foStlIJ
ApbS5XitEcI2uFCM1b1T4fmZ6d8t4hd6zBMD4Zp47ASESvaFzA0/qRH/ybDFD5R2
xBhNLWIPrxwu4dv+Q0GDfX6tQBFk/0a9oBZNuduktZjJL9HriI6suT5YS7+5QpXE
CLxb/YcL9ecHUrayLhs030nsGSgbxk5faNMhptJO752YdRBi3I8NlpiSa9tpWaWc
NkPsqvZmohalvl7+PqFycbA9ARkyEW8VeYuhu7jX4ys2AMK3UjTCnPooZLC/pqYV
OE9/y+T4DkKERU2uZoS0c7wTk3/bsiCb6ZiIHtCzhfCRmVcCPs9dIOds8dXczRMX
eH8FJ8hkz8Fad8VFvmhX9nwAL2jvRcMfAxooCO5DAhjwve+pGfq6Zab8MyK8cDbo
Al0WufBVzcD74P8SFA2y8PwGPQLPRMcMKYSx+S1f/FuaEBam8q/RAFPItocQV7Qt
BWPW8WEvV+lZG4AxOKW39XnhWfVsod5Z61Kq8B9uHaJoRznXU6rdfdr15ocVHEqh
VwYUSB+zfLC0GK7c1VIl/hgPsD8QX2smCAPWeatbxIDAMLeJwFQ1joG8u8SRpNp6
2QwU95VzzhUX/72WoBLhdpmqbPdTJv+ZdCGWTL6kbTw2TClVAC5oaGFd4eOE945X
AHah2zwfXWrso5zVHAGy6pimHcO5MDlxBXtIkAy7r+X13EfbGuoAwTZGvFnKXbx3
CgC7Rmosu4Jk+F2Og5ur6FLPSpj/FF5/ZZ0DI2j+xAHGVTUk5b+djhM8Too3XDP5
1VEd+Dxf/kxy2QjEo8YETQdIlKP6PVR4LNos9u+zXNSdsFBUvMEmB4FcwmCXp/lS
p1f+m2vF+XuOwBhMLjtuTVBq3feuruYlsIWYdd7mAW8RkJJtTm15aoGhtWvpwqI+
4THkK/WGeYZZRbTVFFK6oPC1bhRxvij9avQdsc+zn3+5hRbeH27mzhMREym79cv0
04d/QKg8OGLQL1cXN1pYnAjZp7OB6yy8LKmCBPcq/EBDsGmnmVOf8kLXEEvfq9p2
QM8idQY6Db2MBC+rA2JX8CDbnfZzkvk8zijWwQlh9AYYIidn0a44B7U/PFe9pA1n
bJJH/p/HPRdWLU89enf+f44yX+kcZfD94mQAjsBRqES44rzaBvmIeg7LPpev7OiZ
yALfNAMzV4JGJT+ZalD6RxPDyIVXX4HlJzcARQPF/MhW8tIzovO3WdruedVAqJ/f
o0bolTAtBP8qPfLH4P8aMe/cwRO0iYyJUYGvN8cP8whxoZwZvCxLnGqLtUzvtm/U
IrwMkzyU8jrG9LB4NHUIXR7VGfaErPRMlUGDstenvLT4oYEPGY8KhFtYglAZyYLf
iFefHYaXA+Y/h05pw01xokQrC4oPc2C+SCtM2XAECRekmvaklrvz738mTZ09I0Xr
xveW6ODCKz1kDFNWhkNvPSTTxw/rIpthmuzOrqdZUxHcUE0eRiNEEIVM/HmkY2VU
BCl0C7GV3QL1qh3dTZAC8Y2D0rH/A1f7p1QwAi+WULgc97svEDq5YoZ8EhckoJsK
5tUYRwU+tFpNyGMA+IckJudOGoQ/QMy1WFdDxHHq8O2WRtW3+jz0sGISyg0kZy1D
V1Vt2yfy7VHmHyDO6lpyLTn9CyFLRHH/kiyRWiOZ4LTn4RmHLVG8GfrOkx0ALF6+
/PS/SrPL1MtbzEMluaJJHKq4lJzbK7368Y8usH9gRq2DgqVfMfj1/V8J1Qhz4xup
e5g4GEVIaZb6LwidVYyE9Ll1pWGYj9xDv9+i9hU+XZuLKgLUD2k4AkWdVSzYKmIL
6q4jRTy1QdnOjgEHILA/msEQhfdaKRJGUYJmg1/I9gyYzc8tj4kcl8ah2H+Iim/r
vhOPeke4j0i2Ll4AVgLOcm9bzQ37X3omcCaeYiugMBBxKbUzJzuiz+iQNaomXg28
Fj45LmdoFndCvR8zU7+NY5wsBknZ5haJWiZhTKaBeyNvgRJiWl1or94mkFZ7KAXt
afkxv23ceD9Dx7AvYWsL+VUyLip4uH8kf03JpYxuUHkEQm8BS8zQAu12iIh6iZaq
Bh+iwUv9O7oWb4KHOk0LASI4vGTjPv/EA2n1YA+QpJ8RX/+79JsE3MQ0l+OWH07B
TqnaxPrLi5i+EgmywGDgjE7dUe5eoM5+gwNLsN7UpEeKLU4rNFQ8eTKuJIhsOuMr
ePznzFt0U+OvzT7DK8wSaK2aJeQgTV4FZxyUQnpBnR5UsRbhfi9NcASP6nZZvcas
ArVdLIfeYU3hcNUhKwYA3jrHrdKk9P9oXLdFKcC0wGG1wKyXMqdX6hDayQaOIETH
HFdvaERwYMzIvmbcZM7WAe+lFr+nzeNkXD23HFQ5DsXImyrb+TteKYgBbgce4AuV
kcq0u8kTir4fcHFh4S69O8vhR1oxvVDt9JCXjGtlGfUpnHy8PhauRmzYS5jW44nL
pmOPoAqNEwNISBC83X+1THz5Dqn48JUcw6XKZZpbuBVhzIaCykkUKkiVeop7cZj+
jLdkxWpmd2xZfyrSAT4O3RumDByVpkCz1lgy5NoXDx8L96Bn34z57j9zQHRXjXUO
SnhwFVAOVyWA00w/TenJx/toZYocQVgYalfdxmGOwsGtLsA4lR9XLbSLXK0vCQMu
wNLZ1vBsQKx9cQCIYuO5CL+rN2oGYvuA+kRwYw/4ZtJv1x4O0vc1fvA8NvjvoIRH
2+78dbO6lc4wSKqW/XwNnUIQLDvaaNcPo9Mj3Zm8nuI5TJbcwtcIsVz8nchJl8Yj
RZRo6byv8ozWCbfPbaqbLKz2JJtWl7JvXikLSJASgGKoW0VHvSVMB0s6tIggsjET
SJqPokHDHi9o3360mQDZO0/evr4oekPAzkt7Ap2P2zuD17dQ06Lh8TYb7waLgPOH
f736vvGV4RxP7/Pn4tl1axextyXn2v6uYfeeLWHLAqbUaKqpAF2Ay5O2rMJ1kfK4
GgZLrJbFHiC/Kn4GmR7GevHJGpf+z0DhoD5fQ9SoReCBtWfe2p9f5wh0qv+iHB4X
uDtdMfk+9H+BTdqboBMzf/Una+m9hGGo9H2XwIU4ZvOKiULV1xfuIqSFW1WVRWPs
0SVL8L8bhTg9bmSw1Fvq61Xcb4z6D8SRhWW6+mxxUUUz57xlWsuVhfYdVu08fqvO
W3jVf8Inv6l+Kr8N+91sPFM2KhhOo4NU6FHVN6jsBUeHE5N1hpwhPRRF+SpGDXbi
sub+W8ysuruQ2hPkH+2dAjyfu0NUtAvqB8VBru0owNNjfC+3WRnBveocl/8PVjiR
2ErCr4XHy7s7vIClZ57oqTd9uzfl5ATPkLnk7y7P4VkCtRf03+ZeOqwLraqb0li+
5NleGZgGIe84rM7P8vuonajlaqhI4u6oeKG8dZBsmz0tx4lsQoVk+HLp2zRLnCpL
qi3cx5YWAx31InigOwK510ASSmO6gS5LuRsei+4C/BJE4AUmu2J+m8sJ4+xWqbWV
cV4r6KJeAnBSaf7KC63WhkFLVUgq4mDmbnypNAR7WHQq0QmqiDSfGaY9cIYsQN+2
DkzhZX1UqC7M4kgd4s2dw8Ect8HhY9+L0eMHbbgEKQ9ZeblNhW5MPwpwowLgHRvv
AT7Iyaj4u5S/+jHKetsUAAf8yLvRuc1hLUKPrJ4dqbB8VaBjLykJ4efwbyadLhIK
Kn5oulogch1rK07uB1EfeyhSFxySycpx5+QA56t2Xit2aknoZnD8DfgzzLqZLH4a
3Ud/hH7gKAy49MiWV97/tHydbaFN8mLSFFEHQ8hrwxig/yPC89ka2GhGZ5YKA1gL
bau3+ttK4KIsUVPzs6Q7/ibcECxLUc18pznhkkrPc85oLyVEkcwYc954duVNLjHk
7rhd/71V7Pw7NvgSUoxa/2Za9oSfPCJKGp8V7bQFLbKWZcHQa3uAzpRn63BDcDcX
kfkpVHazHaPNHUYs76hWDsSX3nQyjDB7gf2tBh5PiSczMHDLzhh6L5xO5GU1azlH
S2g+WDA0Ls46MTiXk+eOSQvTzKmqcpFvxTBbSUdVaUIPDbX+Bdo2BE3UTl3ImN1u
8UqN070G80qsDpqF21DnMeivHRowwjNLsXXhAmMciVNZKkmGu/HI1sliVtyurp4H
ioYgItnkqnL7YR/SMjCSl/2CXXW3ydNDWWwnXH7P4Qqc2Dl6mtTTQphSqxQ60OKa
l/CvyzAlHJL+DpRBAl+YJ5Bu7A646CaKnlwliJ4TNqQ4qEdxBDfJaGfle6JW4cku
B/4kGAwRD9mUBhpmIiN9e0jsixxaVz1hjbz7MndAQi4Hg1gA8uhBf8L7EXK3UlKE
PlQvR/fJaXrcmjVEe1VhRjkC+IuVSHpTIQylGJBuq+gQbqCF3XtHkmKyOy47vhLw
rBfBwMbbv7Td7LVuWuD5mPtgY6nEeLjkykC2gyB8rFNdcM7nnCRlt2Q1kmOJkPoi
rX9uPEl7iSDIxXQt8fb/BdNY+JKk0wzw30aCKaMJna5jDOgcB0CLB/zQeiixzbK6
wZwhJIjYMbZ6YdIHEyVf0mc8ytiUIXRRCkw1DtNdRCwYuQ2+qgLMdGZZStD7fC0p
ZumHk2IIciRK5aJ6gYe441SWFTfdEtu3hjyPbasdL5eRpeeRUKaDcOlzNC0dj3I9
gM0kBNiw5yo4JiRS3gv1U4Ojg1HlIHrAq0DYPMpTthcS9v5FJoLt/DuVsOGF7CyZ
c4Zuf1NyCSxJ7+nz1HLG4krpCwNR1q0tr+dcEZhzIAxbzFSsimD6UkbuMdGF8BNG
caxCkHdkUVZOUxtrgSNtLxVVL6wtt80aGFZ0VjC0BD2bjRRCEzk4tSbSD25U8+hS
x28h8pu/OIOpuaFr4C/SwizeVBxDEgDz7dayUKD5B5KG83YaUMyAfQUM4p0obGTK
zJhpBLuFJwqeGcHr2qK6X2/yQyZHDGzO87oQ74PU0CttiJTIAy17pArGGj9n86oX
rZ+CjFhUUxvoiGIKu3nW4i9KoYMnQnzaIgeRaM6LTGIaakynJC12xIMxv7WICubD
xvQDi61QhXmUaM1aJyhD1kzPUiuDDDLN8IeiapOWo6zTQ3lVAp2EQJmX72QloSw7
KoibYxIQgDFQBgcZoPQFoM7AKt242yfwY/B8aCS2bRAZlKcNbbsqSsuwu9UzA2yD
6HDnTqJhxZN4avYXC75VjyoC5CczMouRsxVm0tdaGbnxd4ncCFYGesCcd5WdY/3e
wGsJHkp7HRmHvIQgbqoNCqcBVfy913weo68E+jJkuSR5jrsxyGkE7xX7hEH/M5oK
m/IxP5xP1DqThTr+XZPWK0f9k0vaBTeiYJuSZ7OMjvmFLZs89wYStN8J+Jfp/+9y
XM5apCherkNLvHvQ31eFOla7diwJ8TJukQM+DuncmWlAhuZAYMQ52RDKMStD5Ahl
zI2fFBwhGKP5+t4eHEWEDminrlGnbA6Um/RtpxndQkimRThgY0ia/6yYI/TnkWyG
43LyvFclU2i7LJqXBje2XpDtj/tCWfkC8VZQ6k9bQ7ueMDMJ5+0MjDNXvVqAgLff
CK3++pL9MUw6MbpO1MwaCZGle8MycYUryXSGScsLQsnxUlOHpjiECP93hI8LBxq3
Xk0QM3Hr74V6/ia2fmMWB8jxpsG2GIWaexiupmXU9MdBR31x6YNST976kP2998Xp
cPkReHErguxMbZ5DWWG+liuD/cvGGYXLmASIBgotdTx1XiPsT4wdYwcuBeYkrXBc
DIJEV89K7A72cSal6MVnuupEFReElLwj8QKgQjNisn3C3QbG3GXdg7Fa6vJl6uLd
rj/SyC2V82TKhBg3VQxm4jjITL/AQOuEc7ef50maKbKbXveCIu2PfD72HZk7qqzL
ybyCDYieErNPgrvp2N+CCKj7QWCrOORHL499WIu/YJyw1yNukuQsl7BXvOtBUffz
JfuonEcsPuADEbD1pe3atJzVOvKE3eBFWFnGlZerwjiW+aIG+fAIX828k9pYDboN
oe+Yr1difZul+uhJbijT/y+gBxn/4z+gZp+6DRYOG9CFZvCAruumno8/NMv7FIth
QSKM04wABlkgTktcbTUb5uXHcXMhFGk+sQBpiare+UKzpfMPR+DktkYhyepPxk/2
BfzWIpLDNv5RZsJogh47CbopFdMIgGI4cPm8zbz53rAZMNIvO4txAem329CMYPC3
TwQEpQcAelPJn2tSNih2YPIcNGfDH2ocLku72oIiG4xR+i3rRmXSkw5L0ECm2FMg
Eqnz3xmIDNW1M8YVb2W59oFF4VJ1Ptct6FU/oB3ycohyUKkKC7ViGuOpijptsSXO
326irDRZ1SYSSOQzoEapqbsPlKih5cyUZk6UVZWPSXnblaLjtkQUKSqO6tGAeafT
bIFqgvcGUm37/yQ0gBSXq8HX+AxC31fEzb7N2uHSnMdXYO0IWxpy0eldbvk2rjnF
Xw9Jba+HTFbbrQ10N1CHPxZjXrfOdWlfpcZTKM+uH4eWWtj/6R+qj1Uqc594zjWp
1B4xXgMzZUQb4YIWCcToTpAVKimKZ1AzeLvfYKcB9WgAw0ytTCs2zVSEp+dtwddx
C0E6kt5uTpSNVTkopolHVKkh/KYwzbzkQ6Pf75to6AEhzf/G07gzTVYcfO6yNuyL
h3KNaT+oZJGVPARXHkEKzHHVUFqJvB5wsepFEwGuAHg6fsZOP5vLSxB02sc9mVig
fCNsXCVzW8u3XBvnJHvLEoN7cY7w6F+rnTFN9RgfJl0lAqG4DhTZf9UInXzy98LX
dX9GnDIOFk2Zm7uBg7D9lxjQsslPOqjVLKHsUUHCtknvZBjAQLk6LcqZf9rYmB0S
EvVVSaR/06ein//FOSb4Q192sHzlFkaSbgYE8DDmNMcr0BL2zeaTpqwoTBs5pFIH
Q4iZj4A1HKxfVwKTfB7ETw6LqabeaYYe97Gi3J6Y4uiMDoAK1eA01BCC0vV/ugl2
pkSHate5qwVBNtLMCW1XzX7e+ZyhbWZgSxrnxHL8Yn4CO+P9Dc92+ll+ntIyTjnB
GSRiNl+58yfpVyetjA0ct2OU6gRPCPZjXuWlfSwBsk8nsl609lQsbbg6x1/NHMWb
pVx9BXVPc6MD433b7rw8vlgo5Ftt7cgohjA+GNgsfAIr480unwMDYrkAyO0U7KL5
a8bJT1aUZdzDJDvy9xIb/ohipG5aUbrOoMVl38STN/qwHbIFxtXE9QrpRwaPetKW
k52BNt0TcfgWKq5U+t4eP4x1QpS4ZlSlwKPV8IJqhBUrOyfP8z+9hKv011m/Ctal
3czC3qmD25iWiTf4kWQJ37viMy98h3MpXUOci8cZ/n4F4Ylr6P8DTpdiThjWa7Fy
ioGVTAwJid4XgyJmb1lagIB0KJmzG73uL/undNcdNnhA5cFx5pOmF1XErteWmM9a
mFLInsvpjnh8aikPRgJOc+QHOttWCSw+Rgbo2+XczEmckeGCJsXKPH1ttjmqElbx
pQ/J2uaW7TwESVKjPnhXRyYRGBaEjCbo4elYZMOeIlt54BGMbIZnY+DKFGM6Qsvz
8EM/FOTDKt9q/dheu50FJunUroGBC9TokFM21npoWjhT6WzBtnFS17EI8ttcqst7
MaXuAMlXY8LBf5Cq1tpCUollRzzXqrEHuKpGv79TUCmNtBVaETnBS+y2jGMh5R1q
l/vHwcVbesoss5xblkj5xYsIOyEYuVOFoMxG6hZAL2xu01T1APQfi4zFk2m2uwUC
aBz5+LspaTCbQP9Lrbx0yxB63WCC+gbSvmbx4Q6hm9pHiTktl7U78cOfzrEGo7U4
A7ArgAhePhZpXPDu2/oUptG2GIvq6a6nHrBgcWtkd5hZwBdvCoy5Fs5irvGaV/dF
AcUso0gMm9/M3Szyatbav/URUmh34FKltBmYmI3eCAkZtgY0Zu01zTq4GQKsUrvv
59ukigqNOCxrD6xmryEkqCz1UXk6KgtiNUDspMBlZM5G03eRFG2lZbPBnMxcBPLE
BGTygyHLJQkjKRmkGYSvPLLbzyBbBeZC23o9iGQ6gSy43Mnysjnltedd1Qqj2PqK
rcx20PWATC5j07RoC1MK99jKmGw15xdQqS1emoqJe4MgXvDq+Lpbbckh+vMvazjc
uIqWpAC+bppfyjM0lrmb0H8Q/mHnJ/Ni7cnHLHzlL0iAjuveKyJFxqVuQz/M1jjH
9IzytWu+Hc4ipDGCPZPfXdr/7FK6TVcMiisw35XzYCML1ZlIhKh7bjL9B12z70gg
JEFFWiX05F3uMocn4bPsiP11+XxPK/OSvSSBtQ+Rb3NmZjfYnV0LwPdvVJmprKAg
5buL2yS2c9R53454jPAoTxGlYeLX3jkzwc+N++E0kPBncwh3iauYBAnmvIWX2Ka5
sGlz5d8Q4rVymWfH9FQxv+XXpt3Z5Fz+GxukEiXcWgHptjuc8GEqeX3zHOUDthg6
fcu2RbhI098X9g0eCE7q4bg26/Drfi0imS71FvWIuGkxxngTydUZH7e5J2EM+J2m
I+z0GBfYTneuR5EISL+yhJ2KoFXC5nk6ZwglMj0VMzOFKIHZdykeUYMjaQgHujeJ
z7k0AFKSRg9knucKvFDJspf2/jKUy++uNB4sl+UlAleuuzMs7NtLAPoGRteXEFTl
/rjwTFy60BmHvsUrVRHduFC18Wxz7mGR9iXMigPas2jM7Xm05wrcpCA0QhdzNARR
VOgiLDmey/FH/VStbkY9bhKSmj6DhJa5lZxG8M5VlkRgg5wqt1hFec++f/VpZL5f
claB1fcFeiu0z+0H9zrw+kKxBTokS3oVGEhDaH5uku6/hcuVW68/GqP0jzmygFE6
9XGH0wEVylNZlZFRWr39B6BbBCWbfrSo5QVmmHUlclQ0BDx1MdDn/i6KCP16otYN
+tsZoUClqcRLeIDK0MwP6ewjGYSHZXMHHSj0KCYu7xWizD14PiqkZn2OT2K39B2f
IPeeexUhSMnS1UKbkE6J6etP/YHTsz/ps4niXvMAoe+3MLxvR7ms6bjT6QDpgi3h
d42y7QUYWUCZCSSI7fkNsUkhqamBs0ZwuWyJbxSG2tGVZ10bgszDkM+Rze2QY2Z+
58C5LrrthxN86Z1KLNYLaqd7Yc1lwfrNEF+eaGQS50tsqaEEXRMSwhZ05adLVA9T
bD271zD/YP4SldhCJ0uKQe2jn0Ks/7/k9J7MOuYflHPUsMZaxZzzRnaYnsOO4qzZ
X+0na3Q8+mVlqSbac4AbMGOM4Fg57+0Km7qGsLS96moVFZVAMPRxxl52lLd7UX0Y
hhgAoSNIa0gwcnpzOomVmJ+t6S6V6SYG9pdrWkSQw7JRe4EZ13gGqrExXhVGegma
KjdoxPm2P8LKxJ0aeNccRsJ9ZpSPSfvTuZDPjM9OG+5sSUnfOn9RyYJLtf74PzNn
u/rNBwP4W3SEgOIkKd/wvpnm7k4tEi4+Ka/kvweTCK2prAFj35lGosn918xWWoOw
6Ai9irGai6pJmXtp9w9LBvBGY9twdrS87rPT/WqiTz0PwiJdE631mq/UuQuuCfGa
0cX5VLXaXZ5JTpO84pz5zS0eImbPMKVy010qIfkT6kCVAJ3cWgM57P8sPqjDLSOI
3Hu3ougcdahBI61QHcFCGLEFN9HkePRtU58XryEnzBHDAJy3CwdUpkv2ZNSVD409
xCanI1ovgPpGGcK31jwhrlEoMZ1mW3uxhCVYBvicWFBPSSclQ4eLzl7Mwq3RvuR2
+ISoNlZUgY2lavhW4Lb1ATyViDVcyZH+sFymAoP62LnbqxMq123/UsUaIYkW1gez
dRhISiITNngVhTt4cLBt+eVpZCMdqUxeZh/w9hfjg1KF+YO4k0my8k7borSc8n3i
RFAc1BZ8irrFKEGe0CHy4UOeqDMC0490p5e74QuVcsahmTqb3Dbfvjb4KAzLbKPc
Ym5cTrPhhiKwTqcRjRzBE9BgG6CR/hPlDfQkfNIsz6L+95+JT565kNfYvxptj+19
+hPYYS6HkJGvbVQtfDu8yDjlMm8NWDwgK+ty/Skj3DJvSk0DUxnwJ4//G/zeMvsb
eAMO1oRT82hZKB2gVMV9e9p8hZj4WWf2ZYcVgz540wCuK8fbFyS2o4w7nsiLZTey
A3564M+/oSCBNiZgH1DeaZh3bzFZ+3AuE4GZQsF7b3qIfg47sMJ/M93oy4Sy7J8U
7zrXxxfyjpYy6T/3WzQAfCY3Rwcf7+yclp5isJGlFWEGZrskxhzINxoT3tNIHzDo
TSyLedB+nyQJQSjFlGLxUNNzMMsJw23L9Jhbn3e1DqAQIPSSAcpzvkiiK/grhQME
dUBbVaFYsioGr9wdg1MVm3EKxjjarQfcp6cYJgNU5dVT0jAqICZzkWNtm5AIOzaw
Puoe0qwGP13GngZOLipWJLHcFx/mnmWXppv08pyZo9+ARVhfbG6niBvqylAh7YFc
8xWa6yjVzzoBf5Y8HcjomQ+wTAMrwGVnlTVmtBkMMSzv6eeW3ouoaET+rvUfrPjf
eqd8JbFL2q6jwPv2NfJJAv0QQ3YFJyqj6kLEDk7g75uDgHli/iIGiH1tpc4tANEm
6fGLduTft4AB4a9pA95WtMiXOM2VcLi1U2tN/Q8P89F0voZQ67gSBkbmexTyKWGF
wf1bHGmGiYwEH0OR12FBfF97o/wtq7Gr8GGX9yQAJcShhoTH1nCxgN4GBnjxbEq5
EBBlnFz4g6y9lhHaWJk0nLgl2XMSHswMsnW7gadqu0/dkZAc4baQK82DaxljLjtM
0s/sIsptmC/aK2ZaiTGsh5joc8L8Bw5CeZinrQWsHM/xYz7M39wVQVPb8b6Wg3R4
0dWdscB3GOFXpjLxH03peLFeWEDtgQhO56G9xhW+60hmXjZReYHkoyIOmABFlBOI
a5l5Jr5Fvuy54y867fWDtvh4nAm8PRT8fqddQKMgUxuskmU9Hu2Xhm1kZ9XgGR2v
A4lRhxuSCrstJeHBraVITnBQ1WJftdvIn46GmSAeMgRWT5AmXIROylYOP5jrjad5
zlywrG+rgpdmXzr4weoh6pjXY9YxGKl1lEKOwuWjqEaaJgD0WgrSSA1ubWEwuGie
HFRjTemQPDZDmAUqj0e0dXJnMjOmvMJobcLCAZfHSffJ1rJ4ZG1RQvkVsZTI0QRU
y7DclYLPD9XPaIL+D9gby+XPMIUaX/qRF9szxplRCdPT2a4kehKLDNafuEEfvhCv
T+EZh5ZEtqFKrKl0JANLmWMH9yNHOwy1DZcuLd68P9yBnCLZO6uJsnncrcTfGEpK
IaqcGNj0IdJnzQbWag0c0+FAyZQMA/mBfPgcA5RErX+K5FJhM7qf64e9SXnn6uHP
ke+ITwYZq+gxiRRgQLferDtkbpFimFAW6j8W5MSS5foFt0mrryDQjndyOQfyirrc
QTnW91FDMr1ycLxuaoQXn/jpIszEa9ug0yRjWdyz26fvyj6reb7SgQOmRpkLm6H9
rnugqP7vj0sdY2EL5Q2VnSBtG0wDeSTzCn+HshF3XZE03ZA3DeMRAAOGLmrXsfxO
FkUouYsFjhWW06I9rsw53txN/VEEk0PfH9f2qmZBubqxk83yDU1t68kGUWPPqIFD
hi1GrW8jq3MkW/0cNlhzjste+2+srHY8S0vXSEeulqZtcTGRTwpXjDbBrte57xXC
UeUMBu7zDRvX369phw2K4TgKjcNdEcS9DJYeguPt0IcsMAHD6nlbzLoekI+QHMEB
MD30jJCNwBl+X3qsPy5pP9a+nM92WVBjOT8HZBOTmLyFDpLruFRZ4Cnr6v4UC+CA
IKbsWtQH/JimoNZerBv8OViN+ERPrk90zYY4vb1cp2ykz7rdjhyt+EgPznO7sD0t
uS2msmWtohisZ6mqrWOem6jWTIaa/Cj9/zf3l5NQV0Hn9GiQZLBIKA5Q/HZE/8bl
t1lfxEvf8FBQAqGEn+Q9OZ7v7H2hLyQmL/H6d6mDoyUP7rv+L0GFtBw49jebrPVw
YaJQZ4/NSWsGiPm0AVHNbDPhqk4JuMpbtaB4PAa6HlyqXXa48yniP1dQadRrQGti
G2/q+kL4sdkloKDGjfbt8H3T3VfdEEIlkE7kcA07FnXDgrJfXQO96hkrUL27tebA
63GXn3baeuj4tBVvtSW6jWa6qGEcYlUozKd0qqOKn5nRiAWuu0f/KIYDWSF9gDPq
o1OS9iPvwFrdNosnuhDXyqzBNRnqKbEp8jPh71E1U/6LP//Ok2OowM39F5dDxpMb
7FAqHPuubRe8WD5I4Cbj4LHD8xj7dn9WxS/Agjv19ehfjtHSdhvPHS1LMxn/0tIt
q8wQuh7wpBCpNXMW+hM4Xm55AUOT0e6UhU27Xy/zEBwbroST9wX/EPDNfupIei6H
oiz8ZDz4/xz9YNYucgVZiVX/iWljzn6dizDwIv2S8M+L9vaq5D2f9KPN46VjQ3jz
upCV8IPAXiYUYwj1QYnVknPdIcpyTOXg4P1FStRiVKTBlGYAj7Yhmmlqk4WK1Ehw
4K4F6Kafh+aj29iEIG8PHgj0meMMbBcv5tXvL1iw8Xr3QS27vmgDVDV943cxranI
9x3DcKV7WKk/5160ThxFdiYuAcCdFfC++6jhjV06iMR4WajJu98S3Hr9crvP5FUJ
nlce/MJkhU5fId/Y0n8L2DgWBrAc0s5+iKDlmBdY6cNWMdbxIp7e3RxITKMbomtT
18zGBTJsvMm+e7t8MsFKeEnJ0xCQTKQqAFJu2KN4jGN3TRSszRLACu0BT5Az0iUj
tvk8Z20MfOK3df7mlhk3zWhHrvxzH6Dhx4lZNPx8GlNgNih7JLzHY8f4IQtuHcDq
9I9TMXOawajhXZzPzK2lWWOswdPPBPNWlLHMCkMobEt3fmPwwYQcCPkzkr+Ug0sz
C3YTaMRaF7CshKsQwUzX3VGj1X/zQJbu+j13SOG8eDDUfhM2sIBfd+n75AwPxYgM
Va0Znctxx3+HVPGIWLcgiDm5EJfczFjzGows/8LfUU7PvICl55H9XLxOy/ziXdzf
/V7QsYQykNilBtf6VSmMmmovqGEiQrlntHJHCyEwz+PEGlqrWzTfNZNKvJBK1Q3y
X56DbBpGwgRPSbD/xFgv1J3mFUIxAhqEJTB2BDmBpub0kEmBgrUR2g/HK0M1ir7O
QQyorznJhntC7sPpJH2XiH9O0sRRdsNnfCOoV3vkyMy17DX+tzuUrdPzFlNQfq9m
zduuUVpYo+MVEYyfQCJITBxD8KoplZ7bofj9vrQSQocKFMSL/1qKPGPDDgfZ5ufr
Va1Mgc9md802wWAp669GLAUOZ+bB2r+JUusXTgV8n4QAkx6BY3ICqMWLXNrsO5g+
vQqed2QvEWy46n5+xXa5ecrGWICBJNuG87uIHOOhdJJnmzz1TJjUvWhqZRshqQxA
X1C2NlOWigY4rOP/Z9wMQ/MBDT2teRrVoU0+Wkq+ZoQiRXtbTWecnYG6AP75VswR
g5FKIkaEYvPpUxjrDdnJuB4rEqrhKBtZkDLCK2UrDq97o8LJwadrKo7/JkgKBZdU
/LLHa3GqjIiHE8jFScYi9ZqYdQJgnd0SuU1wIkUOSwWrvCbQEIeMCKX8DKLtf7YK
esRRzhxeyJ6xOy0VFGeyJ3oOZcwHRgk9edBEKRdXiSot0V2bK42bc6v/qfcOt38k
Z19rLRJlglaePXxSGRIhSRXNKJ6x7vRiflsCHfyCDs7yTqmnpBEqn1g7aJ7lQqr/
iq/rorWL8VUWYODe93Qi35ctNBrz1ueXY+lZMXm45wFHtKbWAV1Kql9l6QKy02nD
S728xMLmADIEY4Cl9ooZRDwMvd3pa5pYCux2XLXX9dBbFW9GtD+QrvCOZAbDRtkM
+SguguaKlh8kO5ioSd5ID16fSItYxrYkuomcjG525ZBXWKDle+7kM0/FalLopUNV
P5HL+zS+QDLLBdelp0QuRBEOumiMIRsaBsuV8+IXTsZt5e4VZ63zOROiBXbk5Hw2
hwxBX/oRbgm68H1QHJZXq4w230AysNQhv80tRbvbPahRlROjFURWxJZNZ4F4YpZv
++830BLQ/XQxSzkTxoyYtVpIdwlQhcN0+f/eiCVpm0Ku1yJVuWF85wsOuQm6hbgQ
rXXhZR1CIBOt9b18ZdZ0x5f30eIgxrdolIdf/5FlHdAqWy72sS761P1uIh4E5RAR
Cz5GtF+Cd9Y/tXcRPeL8HE972slIdLU1GoW6JbVgMFbvto5WAoWqRz4WD0zuOLJ+
Mfir/a4WeX1bwT16JJtcPiNyDicQhijnOtpvS9SAcrARhaOWoOclmdzhYsgboH/O
SPE1P0aO8kVotC2XPWiekHcJuh46jiSSdKjerVkUwLg9kTBTt6W0f9KRLrZecu5i
SQpLWWuLI++iYENbN0rhexIriNBINcFJLdpQDudeBK/Sf3ijyofKID+Xmb9eeBaG
kC8YlDGCyueyuovhtBZDzJTK9elKLSdL/UlyPWCdJnR/gu1D53ggvZla3YYJlSD9
DVNtp31Yd6hIfrYFtEFUdAwXNCSkNcuSVumZmrAeeh97fUdUFoAkBgevtpsF6x/m
Kj7ltbydv/zlPQzCTagjnhnasPncQRQ505ffVOwvUYofwPTHp+6zbBQnHChZ2tPS
rHEzDsiQkgV8THjjSBSwQCHdiN3WPm05XBu1x/vvVd805SBqinicMAd03Ar/2Bfi
0fo7CM2LqdZyELJ4gDcpJGHS0xF12vKXFaB+Yj6kSwKTwJD3zhP8iB3ZK008gX8O
YrP2O9KlrinIPEbTKwrGLqpHlMVnLqrL1U+q6ZNS3LJ1pNmU6Pc6MlB+aW1ALVhA
8klP8Gqlms5968BPIrBEywXst/AeA3zlNAwXUrIov74+aHxG6NLa5Q9895m1US2z
4CIg8CzGmIRZ+TRrrXDARPL4oieby73EpuC1tVJJBxnxpejRynbKqBX/wMwTd8sd
/CQ1z3TaY3QQiCim54rI71S5lvQHy/a6Hf+uat5IeE9Ev1N9AZ1uoag/3oOErWoI
N1Ed0b7R+D/KO1jPu3CzczfkGAIr6s5cn3BoAyzLWrVat5yk8PvVpA5q3iThuX71
dfF6+rBtk7OrdQ1iPLjygMpX6VlcyKWXbfqVWHt6Q6CtQh7VjCAKcvo/OOLX7rGE
C6a7e4TVQvR/w1wICNko10sQToL8Ao7su+1kLUwX990BDg35UNEyVYdyF0ZgVshK
z/OMPJzg46mkooN50n7idn/l4lhLW7ieZBdo/SIQRb3cxMCjSgT08YscvN5rmARc
diRszpZwKEFpaHQ8GQF5Zjr8g47bOrape5RbYBUBIM1D4J9Q6LBCbPM8hivA61SC
9wrcuiqoFEO2mkN1WFAHgk6fBtPpa++XWkJmzABQU7HkSSMuOubuQwcB2ocWv69l
0/bUEZp3dfqIN2htYPVyF2qIVHPSbAA4DutmgkIMmcSXquc2fy05CggsM1W3L0T2
wQWzUnCzvGw2pGWnsKSbjHsd9Kt0VcslL848tA1UFYs7vALi45sG8d1af/VD2fvw
lZ6CeUzNqvsA/uze22igjf21h6q19Jr8V0GvSPIVfBGUPbwPsA62Jz1ePLeH4C0F
3gsjvcu5b7yASQ/ykaJfqX4BuJP+i2Mdeo79bJvHs2yQ89ZMlwXSzRBVCg376Drp
i+x21OQM2A+jly+akP4k0S7bBE+W8+rZTbGQX7Kd46lapeGYNYCCnZPQ1/FCRJ4i
FFnl+IaY67x4rwDlFxd21gQAaqGIiEWe8tAc7H8d67x/CN1GpZgMWEz75liaF/cd
YPQo1nDPhTIr8yHbbpzWbKaaB4za6JvKm8qITjuvfS7cOI3Of48MMeSGzquzEWp2
BMlltuPVQ3iu1sgnBNnqGT+1yPU/Nl5buGF2UuADwyCNhMqlFazBKjb74VHIPsS4
bTEXTT0qkjEAAhh1BDP9b9MeO7lrQYOKJyMt7uQVl0Vf2jbxQEZYw/YhkzAp0pXL
7R3HoVXwoZlZUE3xKzM3DyV+dTI2YUTswLrzkiYimbdPJ0+8+U2sv/gOUgEc9EZ2
HrDjclrlRv++4JT96IUawNvJL1iOrnbbFOj7h3vdBTECvmjgXbVcueQGvCKRlQ9J
UAgxXcR0PWzAkO/KULPSZNdlZS4YRtSCZDR6aVk6PNnjeNcroz/8loP/K21GO9DI
qjpM2H7YJpXM/VlepB+xYBc/TUlrRVin9Jai2+TdeCLazbzq3f+3Jd49Lre/q3iX
yVXCeT3OpAoDDmIRQTsM7DXf9M7wlPfo/k9y/SRrq2HUamaJKtl/3jIDqZwJTVHc
550P2iP9dlqVdFr/2qjpUyDOONTI3AJ8UalXLfsUsyc5a1cHucvypJtv4AiUx5pa
1nR2w88QpyrJdY+Vsfjrb6LnKY6L0MOwIVGcDSYabdi5P7e5Qzoro8HEfJAIN522
cVAxCYssgJyFdaSYdMR18LZS9JvxQtprNLy/rFf7QTwYtDByQzvq6vaLKcX/piui
RozoFosmXXeRaIaNnL/8uhF6qfX52cBWNxXL6QsdUkRO6oH8+XL5xRj2Q3+aSJHX
R2ntyPmPHpiryzTV5WW89zU4YutvB6W3snkRTDznfw3EyC1IPmtgESI25ydfd+Nd
xrU+Az7s8oNMr7d2ReBcHWxEwBHsYcblcwWemv5D2Jo7/IEP/XFzhA8aRO1CrAzZ
UOGpM6ElBd1YGmixl5+QjhMcHZdcLxBqqYonqDITAaDBgwgGY/rsDjpLUmr5TnLL
i6M8qRIksHY72buzsaFO70LRHFxocql53T8RlRodKB6BpVsTtOJdk+tKmNXcKsbz
aazmJoBx0toKbiC6WtXDd8tW/Agv1NuIJc1BVLANjUMeC73TPLldYwmwXeVZdGGJ
zLuKoGxJ51666cAqRCv2M1ZsnjVaQqgQwvQ9Bcb/aOSmiajtkI8ru6p7yR5FdfI/
lDQzwEMtb5XDHcMCi9fXvjOSc3VQSdU/XpWmJan3y+Xe3m99vtugwKYNOIqlLAUG
eqZKA1kOgEoOSdjBdyVCVgXwvpFOnd888XwfEA3Q79vjZuFlwz+ItxZceHzC0nr8
O7mS/5pD7y6O7x5NbQTYjgQKCNHLrB2yZ3vuZ8mdRCNRd4402/qCg5rxIpHcGJs7
0Dj4O3uQlfQT1PvllHnmCnrb+lVFX2w7nocddB6+x1WQ64NgXuoNnuQXEIRGvpsM
eRB6eupkKrc3dPQ2d562MBQrcuhwrn+0g9xK7TAi/9/+SyJwW8YVJkLs9am1+j95
an3S3vlgZ+9K9cu6JwVptg1NxX84US6sgy2bz3bdRElbd/iDRT3FlU9JGqlGCPrG
P7a7GNGYrmSx4WIsHXCKgzY1c67fL6jacyrJa0xX3ho+W/XF7VsIbCVWNvBII3nf
JdIfjJxJxKxe1c9GyYQpeoX4ZOocWJ8gvQjRZVIXHEvqi38GKitJSb71cbSfS26w
1SfaRO3i4WwVbtUXmD1qwGSbIo+2VNj1qA3zM4zDaeAARoBcvjWgb+Fz4H4K5s2v
AOl9e6h8lsRFfgMcaCYc3stGRUsoH9XEuJhxf9d86snjgnuMuGBYdX6YoueFQLrB
iM5ayuKQc2zhxQ6AhIYpjUld9JC6H/kxw7tGjUfxWufjQDZMso4Bpm1tvDLPznlo
/hzHyCYB9S/q3/R9adKmqmc/09JPO3FK3uwgFQ/RdV/FFC3JAx8vycchiUTP9DUe
o1BbddwO9ahgXNmbFrTes1KN5rW6GlTwC6T5hZcwu7UGHgPrC1sjqrVakzIUFzZj
SsBeHHNoKPEykbC9DPj/wJxIn048OTgrpBgp9OXqAJqiSApyGoQMwJhhT5pugDk0
hKjui56ajvTFvRrA4wA/iVFanACmqtjj/wBZZBaNK7GN1FS2YfxrorJvP7WTfMhT
TRITezCaaJP6DQ5ciBjeM4qTBuYs2RXYgWxnfYF7g1yX5/FOh9FeHwNLkypn1wyx
QAVvEGWIccFoQVw0NZEDDhbw+3pK6tfJSAIPWtc1Qss2oT3S6t6ryPjYgheC+GyU
2ZWVbg55TUnQ+sf9YGd8Q7LD4jk/Eu+BiGCmJjxvbKox1PMGpKXfi0UK8MyfhbiR
snzluojHVP2wDapjJG58BGjvbbM3B3e+Qp1BMs2y8HTCHzqAb001t3L/TD5HY6oi
3MWufgn3TfR+9WXQQOFCGpSy7y3GlVzq5r1kVe296WMQ/9tpJi2XonvLPSr6MQHh
f04+CLQSIPyb1c38xel3/odu7HRH2JYQQXFZDGJ19QepMRk2AUfj7vMdCunaC51A
m3Rs6bvKdoplY7YQxyzIa4rfqrqZnkrHvmK+yw6mMElPWBk7Ba9qbUkIpNE9Agxy
iqvOnvRgfkp8CQXD9XOF8OMvVkb5zaBNsQY/M+gv/bbr9wBFZZsjR4uXhBqQXZdr
SU5Y5xyPDU4+VzlfIqlAw2XaPgUkeVN+Yajt5MYZAoIGSztVdOgGw6OQKfmqxjiS
CXL9HSmMSQIGJ13f4tRn/k0JrBTQ5OQguV9+tbyzE0fA12INF8y3E9V+UuEGRk5h
fyuUpjJp7vCVBktD7zpUFCm/NKiaBf9rlwNe2JGGXe53tYiJX/1gCH0dO2W35TDZ
V2KgexUlVgu9u7lIRlrZQeAx6/wP1bB+oWD7vcjz5zve9vgGYF6Npz6p9ntBg8nW
LKTcCgILQfCcbtc3Zps7/PttoUyobv2rS7ORM2XPk/LAnhA8ghAVBzcikzTP8v0Q
frC4LrVzerjZd7MGvAbp+AYEL7+/cjFx3JIGYW8v+WTI/gTOMRNJT/BeqR+uZPAs
1/j5WglI6sVXzGKachqwb4ryOob48J0PNzZMBg+0mVqaDYKNsrElEubrOufzcTJ3
3UQo7q3ZYdIpwYu2pFcrVyTUMqQSyN74NH1/gaXB/dyxw/PNAWvPn/4QN1ueP+HT
Z68UWFWyBtgegO/aJ8MA6e2h7sHgvEuC59jaiZmTTKVphRAzid3RUJwNMDk9eQSu
wNzAEarycfozx9zQNnTgNIzT2p4CgIEJ6Pwdll+/qx1dVYSc44bkKDYjq6oE1G10
nt224D98rZv1UoOFdWF2yBgUQl8QakT3Eaf5El6AF7gCKO1mO9wzHPzdVmqUtbS+
B41ll7P9HI4n7Eq6nHL7eaCRR5XEW6nnQSMH2jeKUcK3nFnQKNKReFEz0LLjC5+c
lbXHLT9vI3/XOjCWoHIhMkYPf/rGq2byvfu5JEK9bCGbXZztIq6mFLP0cIOBPsPC
f+KYdh8gX00cUgmlh/fs1hBdLCKk2g10HbBpKUcayEAdfpiowVoQE2tvTjiNderv
AjRuZungEEl0nxYVkvKTOsxOjn3OyG77TVrZDIuaHOFmwzENPQZvuix1HEKF5VI5
Jr37yDfgcE0MCP+zh+rAibUA+68oEa4hvoAhkSL5oRjWYJ/XUipkXrdGArO4lrIO
J6+6MsFCro56oq90gCnka4FcReTba2m1+IjBO3AKfZ491EI5q40EdPYH1s5YDr6A
ouSPgswq+PMUDX8K2xw65OgbKZ/IxBdAjs6zlHWnBU1lIBeCJKkU3eWdyrEA3+1T
B6b3ZPYO2sMDcel6j2YSEukvxUihlDakBLlKWxX9XxOK/3T8TOERScNcXVhrCQ0q
DkZTa2Do9nSLzPefXMfRgU6MK3/Cc02RC19zg85S6PWIEYP3VRilHcNPB5ANlUZj
9AsU3IVg3Z1eZN9AfcE+4LfPDTwrRK9Vws0WuTswXKMTF3EHPe9a7Sb/jztC85pJ
jZpatQhXhE5NUUQ/mXTzhXwDuHllgsj4ldE6sTR16qiwc7I12eXPjxu8JHKWHQyP
7D03guHc/EAX6QWryOvjdCb7USeDx2fF7+pbCVTiaLLlsEMC8dJXcO5RTglFiFwY
QpxZZOmgvXqBHALzOy4vdGj5vhGAwkoYDDm2K0UW7EjnOZiFc7OuypW/j0sZoxOM
C05NK0V+5TJvHHI2xoyyUNjmCHhC6R1brLfTKyjDDN69ecLNMpZc3jhDSlw4oggu
DTT/tnWJVMrhKczcwRLbkJHxbHf79ZRSzalnLig7RQBpAkgQfwHJwA3DE7jl4YvV
XAtGmjHakJieHC9wduQvGW5M4em032G05UghwsRnksf2g/fbXugYkyUPo1zHv8Ws
CIIQQpw6uNEgBQMDf2ktthWhptd23edTLzevbJ72htR/3yknXM6P2st7ZQ3Kqes0
6oHTTkRgdyy6hf8vbhjnstP7EjoJxe8o3cRD7JEUtaz+CjKE6pfwWtibz+/A7dKk
IqFQbVOo1rmYimhHX58cx+E3VIvDRUUpI9xqWf8LFTqI4yy17DWFggYxGgyPMfuP
v5ixXG/aT9YrU43J6QGHbGFmElnSOs6xYx2TiCX9EeRKsfol/220jqidTkKR+yHP
WellEoePyzk4Qe62zo9UmxCuvAApQvF5cjaEQYKRdc7j3ABW6GjXPQCSdO4ojI90
ElPhM2qHhAM+9Dtcqs7/osUP2y0iQikAceG/FkzIwJeLzVYpj9LmWmzehXXwDj3q
Q3Rz/oJrBPQ/33OA3Jc793zWyr15dHSGrNPnbtnXbcAi8eogNBwulUuuTuQDHojn
YxzJ5dM89VB/ruaDDvR5lq6EP6isthZgPUU+RTv3ofIPTIsQf4rZ78mKqj0WyfWT
rCWm+z0ysQEJNEtlK2BHFV/aH0XeExyX8jpkaPbwD8C29bPiIxFftR251wzNc5Zs
CUdJsu+3ou/G4rMBS3ydL6WgUqeInEesjcwC3F+FDiBlfbvbDViWMch8FJcvgUhi
fJp+dIDirzWuSVKMWvElBxQF3Wi9BrpUkGI6uwjDzyX0EiTJMEG4ILu7F9diuMSh
Og3ezXvS5TK7CcPpnbQ4lDPIBFtVbwZqT6HLOmLVF3a4ilM2K10QlA3N71nu9u9k
lr56LIl2WAD5CW3oTgCTp+wrdGr9UKxZc+a9nfkcLQ0Blpb1n358UZc5V7IM3qgA
Hsgu7sYsNiMuEBuLt6xXvGBRX2oNKoeH+aDMnebM4hqO0Fcsc3yANeCb9FZASjix
CkVAiwwgkVj3UM1P8JBADQhAEhUBoRSkmI1Y7V+gvNp4URb4uCbwJJC/0OAJbeon
IJeNlX61Xrxp2esIt9+VlmYZlhVblqhUIN+8F/SWwV0fGDAzkauMxb68Nkf5CxGs
4ymDGsHnz/FLfAd4nbk26teMbKGQpLAhEzYo3pzYdVn/NM2aYxZe8mKqHZdRKgo0
jiEz6OW1KRcsEQSjncKkFwMIuRnkxLiSdHcTAuF49kRaqOaELy76hxn9UMpkeJX5
F9/SIznrSzYShP5DdFtD128yMk9fI84MPIt35mz8zn8LKcT3GGWCzusHykpTV40x
D9qu7Y2y8Z7mATYQBZVTkGX4NbbXRyaPI6znQPEK3G0mJsCznOuB0lttzmKGv1wy
VEfbT25ln+kiGX+xilZrJOcLS4fyYw0Xx07PDERwojuoeqf9uFGWfCLhqQ6Q/d0e
KdhGPxauZh/gpuBMKiJSl9seetaol+BpvnraMFbQEYiVgSuqSjrJu6bnORfwCcgB
YQrVfsSABPBFaa5VJs1KZp5L22D6+mR9ixFwfbR2QhUrU7okWNc7PdlQGeOzsgot
ckYUeV8KF6MY4npakJCeZ9npCQ59/0aII1D9DbgfsvJEw4KwVoQ/EbRRckx2+2rH
Cqn+yITG802QLszagH4SdaZhvrU7j9mSGKuX4eXH3i9F9ChMtnRW27P1Z5QPifkS
C9Pl16yjfIY3nAm4PfrY5/FOviPATSUJVl0jXd/AjBWP9hKdGymo8LLo4ZU/tLaA
qnwZHXfDgpPuu2Bhy9m8adILQIOteRnwSWX6pyb3MiNCNf6ZImneDQW0Y5+wXsKU
INrKzMUotc7F8S+eo0y6Eu4kdqPnVb8Q/+XtYdJmufTTdzodEIR1i2X79UEv8RRk
fMawYCtptsBFPj+94SQEyx/PYpCrOaLF3+g+64kEN9PyNlAmwMitNf04t2I8rtjx
0/51d9Ph7JPEXPX2xN8hZQTkEhk++5PBiDgD6Lf+QOqqImNGoIrT0O3L652xlsgI
Nh8681TC4aI8ZAq2rgKz2W5ZeGecP3EmhjRtg4rfjsdVcr6+7uLBXEb4EdABSpNa
FrfxfRzox/jc5sSmVbzoTB+vF7P1KyKdRDl6b179JnM8bsn0rz0H2HejWHcrrb+n
NYHiu2rkoWAzYwtS8ihOUHvCGVKsgJ/81lb5kwmYHz2dcPwrI+RVP488NXacGbZj
6EHBvvln+bfbsrlHojipAbXK39VwJ83COUtipLaP4WDhj4J6NuV/zI7qwmSGsfhz
IAk5DevNcqPojxQA+Z/Bs1BHByPWGEf+CyCpXaW6MVeMpsq6kMqFp8TpB3DVZNL2
0olTwllYPV1IjRTB40IidW7/laQVbs2wZYGWFxefZWnyTZfw1k0STe4+N+7H4xJx
JzKSbEF63z/ScJLcl6DpqOkZycJXn6vLzFuwl+bvPhMgTjxOj6jWW3SQkEHuXPN/
zas0C+S5AltqjvCgBR2YFCCozY19HXZFnE9VMeult5UVOeK3hUBxKzDrr+wNl5CL
KLsyWpt+n256hiGBLiHtX1b8u70PMNEL1O4UjlVWXoLUs+eiB5QrfgIe7L0T4Uc7
NpiraiPTz3C1PcYjM1K/rvq6mdzhh2t68QeFuERNh3obKNDO+3EikFjvCpWAUKDK
6t7xgRb+ocO6ZI7wOdso8ohDZVEjKedJgIt7ulv8Uppc9wyMALgSW/8Jt5W/Hli6
H17R0gFl+vEmYWc3DF0xd+HAP/urRqEb1bLSAdBQTyphQ9jnW8gYSW75EenUGUB5
yvBzy/2hx4vb2AM93D/S9r0ezNjnTORcJcNfoIsyo01sW6Wuwzyiv34DetU0KteW
SIQBE2Ufkp4g1OYF0XOSttHj4JWg2OnniLdtcIxlMFbghk48b7iz0TnHhn+qwT3T
EI945Vs6T2BayfxxY/21O102nzU4rXqqY1TPk1uwlKwRP9wWqJjYD7eSqKteoHRy
v31Bpy2NAmlza6oRKDO9Ehru17Pb1wy8dbbvbpSHRFi/Nxm1Z7hkyH7aVpr1Ash2
XEn7I+GXHptX6Y8QSEW45TweC3bWjYNwutuehZ8Os/7XR09X6Vnr+I0iXwtp8OY7
ydpi24dlxEnXklu2YEGN1Qi10zHzohNvMO5BsoYVBKDZs2WtIkdqgBKhCKs/Xtlj
0rgx3z/g3gV7+5ybXEU2ToXFtmk6OgnFgTZU5w/HovTifDD/Ur8usCvlXGkx/XIl
J1TfhykIElyH9tY24D8LA86uRJzo8N7BaN4yt8vyPASbtFmzvs7qI5eYcpdu8feX
Q05VXCIFw/qZUtPGo24SqsdCMrgJ5QiaSIsmnxdq+tECU1R03wLHTQ2tNCX/5Qv6
AuXiE5lB1J/Eh4+7ZM23Ja2t5pZThkZn81tOJ1ON/EtXrSkiaYwpl7xbXyAr3UJS
ZMKWLL+WYYoqWSW2FcVMRhJXc425ky+q7rznD0Us1voWjwWFVF7m7izeJEEAwqn/
GhPHiURrGCQ90/CJ08wToWrRJ2NrPCETOK04XrmCgSrIBB8Nh9SGQEYn7l8iiQQr
Brv0zXbzih2fs1ovhjpJvQEqk7Gi7OwS/FGkgYP6aHSno8c4ny4FWRUvVuqgUrZJ
1MMmOqdJxzRE0psKPmk275tS10Qfi44nhrRPVXR6G8aXYTYwWJR3KxVY6FyRDrOK
fCsucyx2McdfIVZxeU/rtou8tpHg1hpHyk99bdAzDaR3LbDUJTmXYkqTPQtiVGqV
/7xaeCdTvw9mr2aBm8Yp83s87n0DIkYVkESeasnnQy6DWjIlEJA0ZsGO6XEvlYQJ
fvX9fH9s4e2vqhvoQPavh/mXyY5HRedcBodh/YqrHIFh/gF8/eyUZpJHKOPHxUD4
KnlNhnj03AvX9XpJWBOOeRqdT7pgnbI432AZ+iX2OUbnyLoDYZGJ8epzH3uRqIZq
dYVWP01yhlEvAaKAuLAwYllV2ZUqpXvlO+/hDA+ksJcaEYN7guuWqZRajK6c7dSW
tC7GTDtqRhJ2x52O7d7gyLUOplXZzZVnC2iwwrznq/I/j91jscGyCd/tvAQzWcmb
nYVs4z/FII1wNVDYkCKyV34Giucv/rRAdwsmY2Ph42kkeZWY7AMzGMw8kelR2uF3
QgcJX4EUyHnKdS27wi/azhrNyCGA5mbGf7f/LlzF252EhUr7FCLHr+1fiSjjhPRN
85wANTb+fhIr9Txg/O710l2XPnxLXwzjfogfZNEQPFkfp6elKrAipM4nmMip2DeX
jTL/qyatHd1KG8XWCfcKkFbs+oMcIM4wBXj5AjiBpzb9irG0qdzyLRaQ77Nyp1G0
SCRcMPUJyvEGGwGUaBCToh7+LAgrjqePmUeFAT3nkCCOeBCoEi6U3Z9QfGvaZ7xv
pGAIFN5aNDZTCZ6ECpYmpB+Z/m9I5tG9STTwaUYWFQI+beRZb96Kz+Xwr2e1JuLx
CWiQ/o8j5UxzjRB9GZGCJe2oGe8Zx/EFM+lOAi758vyv/pnyqKaR0Kq+9KLsnxLM
IFlGVi303ORFyVzsR6BGdaw7WPy+0o7D0AH2sZKhexUIqYrW1FuneLZ8PVCVJr/i
E+gqp2dqx+2WUTK3R05wEEy2mMtVDw7APAGvSR4ncK03mffisHQ6s8QcpYRv+/q6
9Zzt+ZfiHkEeX9IITUZQ3XvuL0+KQ009EsXeyyM5sCx1S+cGyob7ym5sKIH4WQFp
mj+8tTsmNvsinB6a8Jw+XJnTRhbSrhAnZBc9VCyO88ptYZy5lq+KkpiL3++6Nb47
wBB2NvGUeCoGIjXqyL2sXunVVZ1F/J73JyzQTkiDkdItDY0k+YxOmrZM6TzgpNKz
46HbIQpWitr8ZwBRwMzmCGVHfI05RsFr4f5TJ5q4YGtKOvV7ojtI3I5rp1w/UrM2
/bzZ6h6y/4ZIo9+HQwEbgV6T5VIP7bcZUM4NHLhAWEI6jOmY1Xu/DTjXmlaNVwdw
5u0jHiAtljTaf751HvQFzMLqOSKqBQ8w+TNnf+XDDNC86n3MCpc97xLjFbtO8weX
Br87wKLczKEqokjzRh4lT+kcoW2GPO8rxygNc2ACR7qiCPM/1KJiIiEZLYBEj7Zl
i8hQZcjvAw4TdDAH9iHBFcQwY/hgnNb+SG23A29GhgnsqHkB10nqTlkKsfJK149E
/u9Q8Sh7OAgdeTSnbYJtPNiBm91zf6CJbqf/hhcokoPYZ4iniT2nNeBRHybOalyN
iduia/GzcLfqmXWJIxKe5y1x1IdJ62UzGalCPyy5SECMkqMFTV6+nalKjNhbqNSz
r/JCQVknOXdbpIQ0OBjcDRikuyEGg1YkpQpJjOEBkbGA1XtT385QwlP7utSMiO3N
eBeyVvJYiBpg6npQIAJV8fLDQQyv2nByaknVoobbJ0dPN/XinIXMzd0LVwuRKquf
o5ZYn2pbnpEYSfl6S28UvhywFoAtDuGaA/H3K+KQ6o75nW0Rx6E+TlJvmH1mEMHG
J1wjgDO+RxCCXZaKlteeKvnYq8vP4RhS8zMEGhIzTsHlVqKDK8nY7ENGUTLEuR9h
NbjDV95dGyniS2yH/qeAy+S6aHq6UzkAw5XxfYykKiw9BUufutj+177DU/KKLKyj
kae2pzEsFreRoRxeAwjPxiUSKUoadsmSndjpj+2OqfKj3nz/6An4lvbs9g4Pg4+R
SOk7sZjEvN7G4Rzw77yV8/66cqBAFLphlUPwV3H/yQWRU+4u/uOVdX3LwGVbBuZn
NxgPI1Y3uXPCRtph4wbwq/nyjI1LWGBm536UZDggVB7WGPtTCo1GMheCo23ZTFqX
BnMeKJBuEG7TDLutDw5H+vk1l4+qmXxuO45u2+fTg+kGfz2m6kGV7Pyx0v3Fb+/O
a/qCN5W2WbZb65bSN9uF6SeTHCd+C8/ZAR2B5GKNadjXv37xtwTP26Cyf2CphzWc
Hnn0bco19kA8KGtIlopWjKIlj1Aoi98SIN5t8I9OmoDXlgEz5sk8p2QW3uglewKj
7RHhPu4oQDkeCqjfKKud4wZ1fd4d0EmdaLdqZgvf6druoqTIzOBPR25hci7woPK2
57ewGrH+VC3M/bov9Sq/FAQsU9/uZT4gbpTYgkq3CMOiG2yXuHQYPLMt7dQ+0Lrt
HYpG4Z8yEdT0Muz07nxaBL3RiszckeWj/sNwQ/gzQrXSx0rhP2L6F2PC0MiUNvse
BaX0BgSmri/J38bajo8hfE4+955QCebJPx1sbX5J/lfhx0d0rDugBqZergIjDoub
dPyi+JBz1PpS/kaZWiUj9MJbmbivg9BFp00hAEbdMB8b5hRdWZ1dFHxs7J+su8QV
ndQyKt3qjYSn6NnNtBg/oyP4jLaFK9ddWy+F1TH9WhOVea5sI9U/iin8empAElpV
wVlS2gqNmiTdFE36XrSpw8PiDMHnegVNHQ1xfuxXceW0LoXTaDBFLpXF6f3+TMB+
ZYa5s45V32YMXNyLEwN9yy72RgFZgWv8Fi/Yb2TSgp2UJqzCDVPNJvheNQzRKCBL
XhR3iVV28ryiEDK+gyV/9+QI2Dyy//w2varBsh86paAwTX2x0m8mIgvw+O94gsDa
anwSErHa6Ej4M8KvhKUjZkSulehgiesHM5VTBM/QNUYfMtdW/ey0lUgv2uifyLxQ
nfG2ufH59TmvFlrSkO3XIQXi3lmxY2t93oF0Emcny6oF/UZmuDb1Z1M1tFPy4+tA
onkRIM/Xc3AKc7p0UK5HupOBOqPFuA15TVY9ifzJeBzcVDRGWr6v8UqR6Rlf6/gm
U5iez7m3aLw5F8/1IfFbyhuns9C8hUN/yAoa6IqkRzf9fM7oQru074VXX0x/pMD2
RYDfJgEBcz7NKBzjWbyKKm2Nm8HyCzImvcOsyRcZRi0nxbmDU2Ern9M5mDJPR6iD
Il1cWYuFeiOXpCvbcDu+HJ20aftchc0KL7azLirEc2odjmdflF48jR3ZbxOvsrG2
FdMcPBix0Eifo8so1i+SBzb865/tBQh/VzGpqR1OCstJZRsFDi6Ey5KbgoY2mbMf
x8+XFr61L99fPN/CUatrDBUlg1+N6iCBIKAcBt493hakUCrvfzThfeLl68CdODBi
sl3UmsDp+zS6uZiXZlX+OozlN0GfaYFUVTKMXFy3CF41xScEVDQnM21C3PoR5cTx
uB5vdPg3Mv03NLrsvVp8iAW0TH0/Q+8GUcWfU3TsxllwPWl+w0ob7UlFWUP59uL1
sjldbshTelC0TeRHjfZWzAuO3l89Bb5OTh8yVFKO3OpXN5WO/bdIjqqw6kfjy5ts
DT3rHrU7h7yvZG39ONXP7RL41Yotf41kZo/t7Gr6U9vm75zvXLF/9ABNrW8zt84q
h8e9SJyWtnH4B8ICpyTm5tIDstdpX8dBd8IdF8yHuBb5UF0Oye7c0M7D9lhLdnoJ
p2O2SuqCjk4bFh1Oi2vKrn3DPhnk9qa+IGUSA/+16YbJjWh8cj6z3umwZVzW7ao1
Cb5Y1v9r20EQNAjXBwDdugk7VRoPZRNt5gB2mauz1Ho80CV649w6Ebt55gHgmpjr
R62BvD/AtIhxGBjinX02jQ8iHIYwpRKdhsPQc79GO2hzhYVqpHoboLlwRLsfL7tj
KOFkARFtJeYRjq5Z8GCIrzaiIpEw6gAbmfpJBKS1+zPrasfnMNO2KifcYd0zqYGl
4RDiKpGRzPDZllnVcUkRfkilbXJ9Nwq7dm0HjFNirdqX2QjhcRnAENpSHYY3JNjf
DMHdGMdkzHFZWeuFzYj1dI8fG8gxqAo7+BiXPsg8b6Y5TOh+elm58UVF0DMQVEcu
8CIFoTHqiuBBcvBw1arJZD2vPmOQzmaGXSqxGuA4IAZdW0rTmU8n6+QEo+XhIoNh
kPf0bjS2dcv0Ch+VuadOQofZRA7v3FSrdI1P/+mJ1ii1mpedu0lo8mz3h8S1HEZF
3+G0tXQYCLIb9VQ0RCEWSSJOczsWkBBCZRglgYsiqUKifY4b7+F1aqfPRAIpvgsZ
EWha2nH/eF3abP0vf/d6Yxww5OKkWfTjaaF2mthYATrzInrWUMzzKat6YI3wYW1t
uRdbtY5LUfhZhURGErJZUA+Eo2K3jinVhJW4OebBdwKj3PeqRaFUWu5zo3KGaT0O
ndK/p0hx9gTS4F0QmReYisEiKH1iiVUWDOJi/cKOeDy06DMnMwTjhhyTzBeyP1bd
fAKRlz26jGzUZNKT6xS/jJ6D58Fw+Rl4B2jwDZG8zQHN+6X1iPFOaV57+L5ftMGS
mQ3dTkaW8uYK4xbP4rESNUFcxrmA6bfnalPWO/tZ2Yd6EMN0Y55QzjaupKw0BX/f
nUTuExxZQuTgVK9not4IpqjBfiJeVQQrlHnbvNlvvEFjAhr4gf8PrJ6HLruaI7mf
8zKd6R4TxDaM1AvyI29xT54PHaOFJRGGj7mvDaMsv4xQvvC4d+V8lxcWCBcKHUgr
gzHXNubCQX9/3toK62X3ga4VSoTQTN2XH8Iq/tGtZ8x6QKVXvgCmwftrf3Pnvql0
WXKRBYA22MY8CQK1zajDgL8t/kAevlmYi//H6QhAymX/OV04R4OJZUzqObdtfw/n
Qwjx8JoGPEC2Rp8wcQGygjq9zC6VORaZRI9yJJH3SdIF58ub5bd9hUSG2G17FsUB
vEOT9/8etXxnC1bNx5lnzh4D1PQU98ekSoga0VwhaHf8S79hAm4UkKO5GEDjtR4I
51+1e2s1ddiNKlp+Q3xrudguKoazG8tTaToa2AqNGYrPVTsOqGocOT+BK1Vv062A
636lsIXB28pEAlVXMrtjzBn1GelZ7lf6fbukzADP9v3qyfcIn2HiseOG666BQVUf
PUVXVK4yReMxVvomjpmn888YCNzYBIqwuhvvAy/Eq675XTEmXCl/5B0OyJpf78pd
I+2fqKpCIzqF8XrxKFthsVC4lNJj8mBRtJ6tGI5EcNr2zMBMG7hB3kXAeBxiPoFf
aP8L2O3Mk6bv4nYf0idHBi/8bsDwD+xrV7vi/hU3VzxcanPI8elc/c4I7BYCvcve
eBNoL6vnsisI61Iyl5+H+B4yGhPXFm6jXhFixZtRMSInj+msQGYjr8+PcMDBEwYs
fHqPsLLG2dZ8zNDYA+U+4idCgQY9ycMoLE8N63pHVTkTfzR9eBG+yA+H8iAT4j4p
oeNyqsMU0w8wzIwuJI+7L751lnqjnoQ1BZ79dv357hnE49VQTt5oQaEEEXhe11sN
t9zHvQZvS2eKVN9SpFpw++qQNyW0zuNO2TyXIujIf/mE1k6co5sbJz2k9vpWezYy
VEEQoIYE/HlxYQbflao8du4kHC6nOD+8Mfk2EMAG272eKLe9olKBYQseLnYJfiof
zsSqtXYPlXZGsyqDrjrDL/vbmg/lMZcZB3UJ369mWAkNMPiEaRezdZ4+d2pyNREo
rGLB1iq+Xh7+PLwFv//YZbzqNHGwb0ZAbWVaMWOd0Vlq0u1DKM/lD2xap2wQMyGx
WV9kpOvaLkuZeVU9VGrqC4zzlRogTEIEywMTA16vAPmfIZlHjJIQ+mb3xIoo0hVw
QX4g3dr7ByciwViO/upoYZOy+VaVwRKBzqqbvkAC0B0vUI0+tF5RW2QhW1NFy4K8
BD8rwAlp68Ef2AShshQzHPlZZbQPpJgfxCIfZ6CEb1CKpI/DYWw+0HOG2mhmCn1N
o7wSRuWiFUVVzknjL29U2v/itlJVm01CwQC97jjUlks/s6hvwAz4NpBL6ftoJg3U
3A1DPGN7kr4yCJvMmLDQTJkdWRdKeLSc/BA320Uskq4cHYIDUg88zIxj15Syp45d
Dvth0svGpFS07LKWGShJX0KQuKsRpg9GMR2bgny/cbZ491sizWzBzenifzeALo2m
5bJDqgFBbrIR8WYDAPDTBdX8VLx4uRa/sZs3SJ6MeCqXHqglvC6djP9kU80sRYX0
N5XoDjV1sWQw9F44pJOgsRRqfXbQoeBE+x2lFQ7ubiZtRhHHK2t2PwGsiA+TmeRs
B9+25s2bGeNFBXQ27gN5B/AECk/70X7bY3yVLCjc2zbF0q7oNTmPQrEHdW1S29hR
MlNolTkPR5i9DYmEoqUVdtk2QNy26N63ySA6cORH8axVrjEkt88TccvneKbW/jgn
AHlL/8gtN5a30FJAozJkukkg6HqobnhS/QV6zvicKbfalvssbQqEB8ZkcltAG7eO
ryIkOEQ+JvxwwiZ9DWcH3hQ8ndcs3fpQaJiSjLIRNoR7H/mh9cTpieIvzOnkB+PK
FNtD8MIaBX9ksIkPPlM9qUnysA2orlfPujrtoMCbBDg0ln8AblJveRtRJK3BVWsO
K/tkv5r1/O3MY6GfFklPKdHXbvDrJK/CfyWB897kNCSjjr6D0xtCqDOHpD8tzpB0
MdAUVsztVbm1wr5jZdxjg/z66kGmwNqjiyvJ1PidpQs1SfJO7k2q8GC5hKGHRtu7
3cP+Us4P9bONkw7T5oWi8di0hWcPrVLLQJimsoiAKz8RckXZQABhgMZcUa0QzvFA
bY7++f0H2WtRlGlMiZ0P3+3k4lvbOliCxLX7Tgu0k3EYQjKUdw8ep+fJZ7Zu2SkV
8vB5MB6ncA28NH40DAGJbVKeH6BGiTd0YywLJDitWDO41yGZ85tr7o1uZcm6WR3a
y7/IN4Q7JOjR0OkTWMg4g5wNjsOQl7SkDjxsygwBJuj/sew4MRNfnuGSxNTgEgK/
/Pt1AhU8gvTpAsEYEUxlC3axVUc5gOWK9RFpcgk8dPAJPjJh9ut7avfb/agm2dXC
RdiF0n2JnB8A1SsEHjWuBh3uOZt2BMtHiKHIwLqikizBOtNFDjcx+NnuU7x69+0M
M+T6900P0DfNivAb+ytwOMTNl2ZHBsjAHMjcN4qbZ9XRdbQrrJKvRHqUcT84MAV1
pJoVdygQFLvZXe+/GD4fkk3sv+AbRWnBeXndE4gynkzPXdyAuGBTr7u0W3TykVHO
ENRUcj8tnEk/A6V40MZwY7YFPBTcMYB9xUIkShlCy4BTwBJPqVMoAFalAMw3SEcJ
qmd3MhvMS4BgYYnX2yHOyQZVCQx54sE6Z3uKaiN/I72b8B6G/oJ2DEOc2+4+Kcvx
X6wol3w52CKz0Ml4e7C0wMJbN6YlNmNT0qnEdswqA0O3egNG7166U1LBBeaMM6M2
IQWaxjIpmcx1PtkFBOZPuQYAtIZO4QydyLLnpUiqvw54grxh4VX2o4lbDxTlrdSE
3UiGhd8aA988pi0sI4+zUBH8MfsWK9N3OqMpRfq9Va0x5GKdKpuZHITVFcKasxNX
DVY0bd7KG72pghNqXaxeTNmNNXzYTm+ytDDREGxWiXsQZuaSNZui7tjCYSrVTTQr
nMqPrpbbNGJ77Uwk3iFcTBxzpkxzdeC+sOsLg1daRcfwl339DUZD/BZq9PsMOBwv
NHdar0w1umxNtjQWt/cjkiyZhypwmvoVnF72SURxKlw106D86uUjG3jdwVrr5ikp
iEO99DFzywoMj81lg44wGYCg+/ixJoVW2mrFk1nDtDEoNg0pjw1Ur7j3umD/TGu5
7lJiFe78LTNwkA11isd3SO3ZwJBoekOMeWyXv+jGMH/hSZNOJQ2lb+fcqL75gIXB
ycu4MPc2Kl5lT/gvenyVb8erRyMZKEWijPHrwyKMlJ212XewKsxkOIBvsm0B/9vN
4o3oKrJly7SdWxm3Oi+RL8izt9QdKWXcK1wK2W67I6tkgphzOuB0ma99TFNAI0Cg
sSORTs15uTIcfZySYr8JoLPRA/SonM5A6aRfCmLv7bwisMrL1QlC+IUof4YPL/UF
GzoKOPVp+pEJVyHiw16O7F9aTQiGBuh6SUN++4NijhmX15HEHI0MmTzJiZ02EHvJ
0uRuZqb6K+YMMLUe3epJOFNOkD/vfFxLVySDAOBiItKeNuPh727I2Qq3/DHL7a6I
Aw3cSts7faWrUQEZORJMnGTEHPa8pyuKyTo4O7fPaNk+ATYUAt7hG99Y59DaZfLD
SmftGxPXEcOc9/fxyw8f2dhM/aq472T8gzvBV7Taf9BMpXVDSTjf4gCkeV1LE1zZ
vt1qXLt3YcVhGspU5+jEvbM49bGMiASO23DrNTMuKzvGnuXk2QK3DWhwgOqc1KDN
C2u+v42Sco9Kc4k8MTusamA4Hel6s8Q8M48cCB3Q8ZnlXP2yF1ePzssd/SeY4QBr
IUGFwMmEblbgbWnggfS4ooL4siHLWNG7TMG6R95lNhdvesd/4uE0IzMHBOa+klKJ
q+ULiuG71qewWPgmLCb3hVX+29mpar7pVzOe1kCZjfRncogDBghkXtWjvQkMef2X
pWlMbu99tKp9rzdj4KG52oCRDn8blbei9GTEuU9f0/sbd9NV8Sln3UnD0rhPVzKH
8E+vjYB6yszL8wcSLqlceE8/XzZbhAwhsykhPur2p1xNgqsv82PnY0okczNv93Gu
a5m3hxqlTUHP8XPNAxSiYfBEpsLBmB1rTKU7mkSV9yPs/sWUPrRb0V4zQfcoDM2I
Z8QJjn/cpi0zapr45CkNVqi//QtDdvE0t3ESlLlha4EatolYLaMNnjst+us9tI1U
kiGzNk3x/+KdfeRcT7blU8Gki55l8K8wBkGEYOg3RxDfd9EDosVzX9CGVHOQYVg8
R4cv98LVBuL96MXBzAkYKpGvi6bUpsTgPrgF9nEjJilzaQSarLlH1KAGUK11h1C9
bqeY9bOLFsoN0HMFvVz8va6KBBcQuqL4hR2BSR1dV/qCF05VMKGnZLiZUfk5JsYP
7ZA7zrZPuU9ph/lCPxHg92gf2z7zaLvvNod/cGGf6VRQ1KN+3DW9VwAUIG7Y1h7p
ZIrYDUF9hgMaCsxumVEYANppelODLq2I77oiZEAoMGvbKhPQqoOXo+VSGSfSuH/C
jw6bGxwSET+IPjpPYL2mdLDE0xyllfHdVD0RYdGSTS2Ou0d0I+Z16vpO141XEjvx
e0KRirZjOaCrFdEdpGF7zuGcB5v667myeiQXoPr9rmDheOgSiHI+7wras+bAeRaB
aVjuoIRGCB1ZwMnyQv9sbQXuoEeUJ+SNdlQ6zuWoeezxqbxlyw250eJ1yAML2+z1
cJ9el4jpxRUzWPSe8xdVR9OfSCZsrv8SBBPs0oh+xc/YfGNiX63MQns06gNMHmbA
9EeInbLzJ0cOAI5jlIm+oN3KxpZTrGqdGwyZpKvra1jS+tzFpqD9DFlqTnb72GFE
Gs03NjfG6G+4EUCPoSSXS7JkXUJesnkeIwL7HQeadhN2l5FUDRCu/Q6AkwYFHfXi
O3NiJ+WRAWEioGCCujiYuxDD0mOtDZ8voB9qkkODqrgUivblY+PKilxNmGd/Dazk
MxLq1dpSdhA4GxcJig4Gw0iUuTdBOsrWIbI1Dqf1lo+LHnl/B/3qSUNLl1SKuqdf
5+qu1W6iVcSkNcykeq0X4dNBkE/ET+HHhXxyrKj4XjebiMRlPykjUnKlJTl9iZbc
k5nr6OeHgiQGTSVRW2gil6rFSJX6orQk7PtDV0Z49cPINy5jGQ8ec279jLtCWs6/
nHMoSQUfXn2fVCQ2ohPlE/93ZAr7sfgYSDDdPdu+Uq+/83ZGI4vWFg2wibSzW4ro
i5xuGwncQqG7IHjm7xEOc5PSh0fLxkiypXU4FzVSgUNQq2H40+h8q0VSXvgjS+ru
7kKqPlKwgJ2FoSulU8u5h+zcbyOTGa+IiGZl76HZddkTGKZnZ6eb5+GQ2NHExG2N
0ojwiP0scJ3HdXBgw6VSHasPJtsGhd/ywDxodVju8MoVaWmmXlFa6YseQoxUNYFb
GnBb+jyWAW07vu/rEbTNRzwVH8DtEtzQOEBwnhfZ+LJHflBxzLHA7p4iDY/7lTew
htRNNl/aNuTFM6UUEC863PsUUld7Jn3aOO68YD5QPfPb4qxEn0fcY2JYd7PD7Hnm
NJ/7MJFlfVgiS08mJKCU5TdgeErJ2BIPZJwtUl7nqldcOcgLWF0CE3ySAaQKQqCD
IbXfWYohRxQrjRSjllJkjmr3HgsqP9MvSbl9TqYe5NPc7A7j2sKULSVJhQY76JNA
it0o6EacvWO6eTgyOc5uyMB2Fg3bCRcYguhAXrZbrvgnp69CgEpxKdJGwjVNHPlD
aMSp6pJ+x1gBW4X4hRqhRkYqux4hfm7tkMP0UCJkdPsZt3Awbi8X0r34/VqX0Lt3
qjY5pNo0KFuqcL7JhGQ06OloGpIatVie3+e5/ox5undXhglU8sCVwcakSJ4u7Bsp
kKO0liYWlbQ7Zm0O1sFTsrDiRTRLeEs4vsDNJE0nt8yu09d/7UfghcRNuCRZoSrz
LSC02UCFEDsVTjJJlCu9hnxaQKp7KWvVl00vfFacIoZB1gjvh/ZH4cg+8u6jA3WD
U11kqcSaqXMKu6kqjkzVu2nIrc6tYTTGG5uU2oV2j0j+X/h1i14IaGqeP+ouZBzs
lCfNGbW2FdI66Y5OYqlbi5RBFGfyVOI3RbycrJMKtAQR3b86Bc5/cwoxLwjqFXSL
iOIwouAjd68NMkd2gcljlesPXgZKe3ew8o7kZSanZa/U53apPohazuG+A7OsYDmW
1zbI1LmBogEVUqzpuIiZVUBUXIYq+MSQATwDWp56ALsL1MaBX15l51N3/R8sJyLi
HpOxxdi9lHstxDCdo1WfKGML8FGa57ubIxGE/zlnYJsnyL/FEOr9zK1FmzZexTjp
n4TvzPuhZP04qbNDwuTJWyjK6HtuPO8w1IOhdJh4QERFeUL6TygniUPkqLKfrDRD
DsiL3rbD9t5PVBbTcK8Ht0nR8V3KeICqYfMxecUeo30eDF2UVCksXHGTf5c1Ep+J
bUG1DZqdjzkqhmrKQevSMZmnS9wmmjk5m3iuTUkl2jlhkNyK7prhjZTQSLqK0H1J
IAkNtHaDg2qCbPvZE/27I4I4+NSHa+sy7xnXRpB3CJhFKd5XFrCJr8R6BWzMouWg
q7spD1e2YL9cI+NNwgJVVhSGBZVFU/foQGMrZw+TKvRheFljlmGewFO5L4wYO5Yg
kEHrME1//S5VNahsiq0ni9XBtwxLxmFQ3mOuYOBQW0SA0rtcWBPlFGwjMlRPL7aF
9ParGizIycWe6ZJjUIFYO6Hx2dSwLyd4G7MXjaCC1+berFvcldN747yncw2Etkqg
ozLbQZOmXorK4tGhLqgCscMTfWM95RKfIJiH6OgRr2QEcrkhqT1E4ezIUKftPbFz
P9PdJsmM7vG4wQpLyElZ2eOx1Z5EiZILQk3/Im939ojS9XknKfZBJMLeARfeOxPj
LaRuvpjDhTuAcTa6yDP776Ivi7/2PUNs1EKLQQ70bur9qXHvUxi9D4KPQGkRrAIP
JRK0QjgqGaZCrtMbfva0yU9dds/v+lAcD2kaJXIMxgFouIu6Ob+I4hCHHEpQ6JP3
9/XgIngZP80MvM49mTa45PrKVuoj4vPqcMLmCcqJ9rOWiUBB3evUuJx1FpQjm9oM
A1XYIlDPa4PinneZYfoJ92ZCeCwQa2fXcbVwmvLc0+8OyHAybVfAj9AIIpZdDzlF
Y2ezB+P6xBOWWTCJfiR2eCdnih+PVES3D9ZkPRsZoKqnYjeBV58lsnF+XfwxIqD8
gbn2HO9rSrPM0FOf6t1T8AWZOVn9R83YAKZQJF6j52I1a+Vu4Rt/HyHUwFBWgLWl
4bSJwt1jmbcuFJ2383l0AJ1wt1tcAwwfOrIQUrg6VNkDqfIHKGws90HKPb29hbkN
i6lzyjkJ02JGHkTIcH7XURnehS5tBhg4zcAskdmgVksDfyIaFrEijBvRorBjWoqa
U6Y1ckdFFaAhNrMb1o0vZOtkvryWK+ceE4czaIzcVeNAw3/jdOdiKLIhPh/Ub17R
5r45IBjo041VK11O4NCWUpq/2DM7rBXzQm0ddu8ecmS8WCIn+EXZoHoIFsAVYYRO
TGZafXqSEhsz/NFqDd8hdAjghA5DYKRRdQPWjNvOqiF63DRMgLrmiF12+e4yibw7
1GKUFy3DdwYtZQIblF/M82KKvkKnUJrV1gau6NiB3fKQVLOZXBJhT/280Gp+aolo
+Puyi8Ht/PjsA9+czN4Sfl3pftOZjv/jDhUFntM1Wi5NqPYgkwSyjiUt7GQCPu8x
yN2SXe15i44Ajy6yW0lBYyiTP3svn5tGLY8Z/mm8iIbaRoIQtIL2N+2p2LZEvpr3
mdRP2IeV6s2WKFfmDfyMoqLLjjg8s4UMnFcpZOp8c7mvxfN0jGqAS/YTbmYTyTwE
+prxwinRYxxk1g+h6D1q0fN7vXors6bbyzoVS9vczIy3HsXLGxO0JjX23wQ291fv
E9Nu2g2DETMRlK5aJbp1qQ93J9eGqgx2ljd1jWoxwNc+BooNR6YCGXE0RvkwQuwp
ed6c11xxIGIBZHBjwPiAC6lFMk5LGLyZPlqwqiNpHouxooNPv2iUI7Cby2LDSho/
Wa5qn8pkrCg5iy451YuvbFKJmzop5sppBhiI+iRRn6p92/QaVO41/EbDpDFptTx9
jhiSlBtYfwHCzyaZDVhooCapIRzUpsz7qjpkchuD5mDgAeGJmGT6WJzMeKqqkxu1
ZfHWFJj8Y9ANwK5HiopsIUGxgkyI4hGPylObFWgrWKDuyDvFnZrWD/Y2Xin/lIq8
+pU+i4ftI1TbhnoJuJDGz97q/kveR3GTKRg/oW8aNh/fDnyFQWl+xoZbg/TC6MS4
+hX0ocYg7OX7AZRfQGVJNAGmdM0zAds1W6zztw50Ijva+t6XDzDOwsg2i1pjoxe+
EMEB2S/fO4qKk9yNijSCcB3kXp1Y/l8a6Qg8wyCRZp1LLvtxuvRLI5e1+ReIEeX0
YQviVk+805LGPSXhUsFGw9sTv4j+Yb23cZSDNc4Iw0lFVqchsL39Xua18xJLzl94
mlMyhnUL/Ul/OHNMkbvcYm9AzSbHT+UK0Xto5FR4PUA2RC9hg/m6h7A9NFI0cilb
ZExKXy++J1lh3KNLGAuR0AC/3eW3t6DlZyEgs+e+/OihAZLSlYW7WrBXmLoVtx2r
4AYrrRZTnMMdV1ODO6A9Q5EmBRWpl/N3yHKg9cstMD6nsiS/+EzY/ZKYXqBDZDpA
NjENguXRhyfmeJJUega7nVsbmLijqvcJWXR5nh8xKFEAjHMHSbwIIJTVchXL/YYD
o8xSp6DnG2EDWKN9sMnmrXpRuzjyZtuk6vxrxg+5T+BVRPVbHvORP5Ykge8GeLTG
1v6jfzpmAO98XM5/Ij6FDfvdeLlPFPY/XS2v49NRngJPzouEgwIzahqLJfAjrFr2
g8/KOXjNhYXE8Wx+ncqkLObpqjEvVH/f28rGT9nhhUfS6PdxmTkzAeR//AmdzAal
ga72V+ilLzFvb3Dp9C/OPOZjK/c5zYCaR/TlhaMwCoiy2AanZh7oAKZG+TVCnY4w
mo/Kp2Zrkf+u23690he1RuaFVbOMS+dJLquzvyBxRH2cJOZx7WjTW1mA6UxTflqC
RSNuArdAwzSzd6YeWJNCWF0hENKd+ROce3FBu9nk5qWp6uiIKefywe+AY9I7g79R
bRh/IZkQ9owWdgJhl9ql73zePW0F0mcb0RL1f+O0PZHBSTXpBssPt8KWCtySBEpn
bpvXoB2HhKzkQQKBSx9dwiRrUN84Rf8YLVGP5ljJxSAP2yH1UFY5fedv2kJedSkZ
Ic4ww3E8M2/QtjVtDrnpnQgwHsw0O9foe4flh63B4Bi9nudYZaKw8ZssR6HrBRf3
e7i1fMIAHVabcrOg3IWLBLTvpY7Ji/LSSYoP8iedHZ3HvHYqHJ6c1rz3nUEhpDAK
wYY9jLCBMx53frOqMzBPnxumsp0q5NNgaw9zdfRq4snG6yFpAg0PElvRQ5v1q8by
8dQL8GJYYK/CVmnjiz8mEteitP3IzNtC4rdUdkoGSiRQHN8QfRPb+TDVgjBoS9Op
PFdpCXi8Lk5koPUUG1wCTYLcCzSdy9R7CiyMiaJvwXeCPFddMvZjftLnIrcOyjl6
Wllwd4sQSuDkZojRN0n0m/6tS4zfWJV3FUW0cyCe9kyLs98p2MVbl/K3P4i3gp+4
E54MNF+XwEb9QnQaeB5XPABxblWdlVbiWR+FSEz/AmtzZFceTko8D9sH6nSV/GwZ
msQoRSAzRbIGiYBsd1X6O+7hP6up1PXOx7GPo0FQ2jirSkZTy3/s6BAP0zBJg06Y
PAJODI5LP9ise6+jnlh4Kp2v9D+6w7hYWQ7Ilfj7o1mV7ib7no/gE9wL+xeQyffa
L9dsXRTEQe5KC2SKkG8zmmtCUHk4wg/Kjre4OpbBw0eb2aJiOR5IcZd3oCEum5h1
PVSpK+JXgKd1BcHp1b180OvqT3nQV+MgqV6PpdKglFlBoMGXDoZFYccTWUHN4rTt
c/OFUK/swhl2XBjVzJZb7P4YVvCILFFHyIsED/nnHwKLv/FNc2iK9lmmlWufOi0n
eRvtMnX+DWzNzFM1erAvO5WEgt7ObHDmoethTg8jiolZcPZmP14cUCscI2gJpjNW
ReqYSLpJhxnVq1mrlJwtUWeuZ0cgBHhzqYb7fDTJLz1ZRcJqrr0qQID/1bL1RHq6
Bhg8aUfzMoHGyXJiDAR0sz1qRv1P7IudON5IIBoAw5Sg+FGoueCD+/S6Ru14pS/G
/g7ISIENgfExomdyabafQALfsy9ZCr+EJWB6LIU0Gm3PuaTvDUnkwnqHSYwMTyTv
hYH1rHWyogzm8RSiCMc5DuOdpMzkh0TlhqFvnqZTHBvkGJSqGYqnyrib7MtwKwRD
RsJy/jZ32racXaNry6WTiJo+C4NDqbvhm3xfUPImBcV/nnUBLqNeGOwxT+B4+G4O
B03BJRv8NJNC3EGFObae0V4Wko4ehTYgsQ+J+nuTkpCYe5Y8rS70QBl8xZLkiZl4
7Ia4r8Uh4UQa1BLmnH3q313yJm/ak2E1Ovv3IiecGVZC6peq2s1tWb4IL+cNYPaP
U3uDuQJTI9bCLc+X/INRS9HS0gXqmHKsAVAPCHvR6aFBGYS2yZCwnP2zkybVelmR
MeEPF4lXQycQHgZNj8fP8JGn7hvAXRTRGoRjzBBShWNOzVuKogxCtf9YxZpfsCuB
bgRwih8TSs3/XeuzrjZ3TrNo42wijEZgieMywydKpKXQxvUp4uSlEkjMcflN6H/K
HdG+Wwz91e5UuvyTWJEAb1mE1EtlXdTU9Enp7rSVzFOQGjlTlDcD9/Bv4IoU8Ga6
F4dGxn916rHRLVn9/ZoVcDNIplcwvo0Mo7poHLX161tNAzrH9waAzw31962yAT0c
9zjcOIPSAKJp4suIVBSn1XQ2EBmNyTq4msprKdURcMzZL4R3R04cdYzrdpLcigO3
g9YIvz49YcRwl/PXs7b9kpX4f3n4RByPg2rOIWiwl5qnnDx1L8eNqmPVaXeoHOLB
xCkUCk4Pdool2zoUxsxcIXTjzkDPF591PDTKII/5R2tLg6OpoAE3H3C01RSnoUFc
b7Rf1Af4AmIrQCZL5q4n35TsuBHRiBCeeqOPDsxQ548IEx/9XiI9Y9U4kCCpJFMN
XuDjZ8vrluvs+6+z61AMAMfllbMNAbYHA2lhxzYE2rqukLCpDo36O3VeHuPjRqju
08GOxtgFb6r2qvx/fr9oHxEhMgR+Mic3pRkihOihoTMUeGthJwcoRoVaK8Xo6Xzv
q/7Ofjg+7BLEbr9mrL0m21hdJQipVaJmHmIldPHwCxx26urE0vsOI3Y7II/T4hph
GlH5se4acIvf+RSMNFWHe8u6n+jVMp26Bp4QVNIStBi1TaXLSffHKA5UTBirfAuW
6XlOEKO1ILu95Z5b/kolV4XxJGiYx/NcR/CWX9p4dqG3rBxFdbuUNHmX0nguAT18
pZIfF2DzepKVeQAJpRvpC57e//StqoPASQzqtHqWvr+NVMCJtBl92Exv6uihRFBd
Zc3YN9TPY5aFMQ1Fa6hBHCnAA63ZbzI9VWGv3JoDPHIpUtVewF1tVRMkp0ccAL+1
wePz/MRSViMccHQlBd/wsHorDNfza29y0vgl7YXiDT0ORcu2twmAdQGktukopVHK
F0z6EyO0ByeAJhUGQdGQIc+FprDkytA80RrCBozLvDfuUVWwGTfu6JEV8qAtFgQd
Hu3/n8CI96bkG2Uqhk5AKnQS0aeIps11xL2dwrfSvedsF5Gw1alug8eAnm8qjOXr
i6Xc3GTPAaexu4fkXh8JDJ6klRU4OSue1glPuPapgHJY1MkcMgeDBND5Q6mW3nuh
1HBimuQBPi5tLVnRFEdpiOcsNIv0XuCk44FMyLXYyLKAjzn/V0WrUJAH+cMSrAPz
5FxBLs2eizTi8QRwDuKw/TsB0jJ1pADtjyppxBqnxmLc/dqejtBZve2SWv+RegE8
fTrBGajtgP7tez7i8Ldf9SI+RA3J+cO5+1JgA77uJ17/UFV4dF+I+A9jBsyACDJh
3Yk/uZIUReW/lLjHwUoMUo340ZVJqH/CjlR04NWEJoH+7p7HTdsllVBKcz0xFVg1
lO3NUmuUJygSAbk9xxOKtZpaJajWLQ/k3mKt6ZJy4+3vYRkcpkANGdtwIS/cTLlj
HOKE5rOl8JVCbFWbGwITyGWxe8QLkU5/MtWNvMZ3aqmNssItAp8RMKFP5HeV/Bre
zFJMZrrTBBOpTUIMf+HNs72CBJ2WEiCFLRmjq8TZp2skQ+VPZ9utYSGkvc71cPox
JaNl6QHE1sQ5bfpzmluuijrtOLKLNC4spB9QKyMbz6/A8YT6ReOGixXFuPPQ+w1y
sLIXWV+1Xd5k/nf0eaDr/WUEc0EPrIfWa63RYZqqsKztc9YOQT30GzUMrv6txBNX
jknckDW+SRTYcR+yxAl5hRZ9idACQ0U7uW4ljABk/WzK+1zJqOtd5FCmcjEdd/fD
tZ/DL4bVQDHW5H3ug9mIiOwrFPO3egQnj8i9Ew1AEnAItwJMDOu+rxTnbZeyCnf4
/gdpEm6uMU4TnNTlYkb6k2ausDP3whY4dQI0x0UrGNEZy6IuJWEHCWc4VEDnps4t
UJGMZeHtdOCQUBHQ/Leb7JH3Rgpl73C+c0ljXl3z/wbuykfVHEaRQ8QTC8HP3g0E
Prly00KgZ7LmwcyU6I3wU+mNjZCKuWujH+ckeLaBSpqDp6aDPLjwop+Glzh1UpUd
YIijJEYmF+Zk9Gp97DutspcLUP+KbM0orxQRHdDu3kOQJ1LbU+/eD1acqaytXPDo
oDtA5Zi0yfPvTVhlICwYmcAC/mLFnn03GPGIYqizg22zgHU/N1Z1erdc5If6IXfe
aJaMYaY4DamNe1p35uPtuIt0l65C19YHCz5vQUAEfSu6TSeCowLxGqsyAvQzXx4C
ysjN4geZF4dHVFjJ910kfqb5IuISRN6Gw1QBHyqtxvA0fjOUGGoY51x5Jor+9JDB
T784Vt7/eAEZb1ilXK7T+U2gvzIsE62Jx0FFrPuDe4TdJZGKVoFvWtM1gX+XIKtk
d+TnP6guV4cBaum4WjJ0wbt860tWqOMxnkUQ8SATNQDNpeQEBRlRes0qcXQCndhH
5hTyzi8eidpNweKRox3PMhdw4mJqkzwtj2O4glowI74b+einukBBIFL0i28ApFlt
yBc91A40L4cZKcL2yyi+QO6Q27e1nreoSJD3/7XFG9S9/uB/AE+BZ0ruOmgF9QtR
8xxw9onijBXTcxWMhd6kEA4Qp2u4ARJHGRQBvlAXeWPq0R3yP+G8g1OGUoNbDdXE
nZTaGC1WfjwCigpT/IQFmuT1IjptUgBO3sqjpn/7mMl5T22dT7LtPn2tpstxEWfD
NMzPcID6QdjR/n/CX2Wr3qgCuwct/a9HbCb22uYG18ihv7qEDcTEpwUTepmuypJB
Z3/L4gi8kiluuZb5LAcwrioBL02IpWlKxA//A8ZEnc63JnVcxqU10rBBGHgga1YS
19OaSouj9HDADQ27PaiCHSrgZE+P1yjdnpqKtxZjqJ9mip8EMJd/u3j9BKePOpz+
dcYqGOoY0eNisTrIfkA3V3ARTEjhBB1f3B11BnRaIS8S8C3NnaqHOQbEVYJXqZlh
RAAZnTAtvRSUh/K0pjvvfyHXHPdVEQTMnZ2g0XZfC6flRhXTPE5xfXMMbfz6zpxl
BJBLvV4z+BlcfC4ahb4n6dG5LccIg9rKn7q6Q+J4aJtlcFk7+qBY3i20rfB8R8Zm
da4pQmK2HhNcet17N7mJfyPZ4L9A0gtN0ZA8arf1OXY4+3CHEjKakhf8klomMBZe
ke1F9TdbOvYTaixt3/nvL7FFlfHoUxysjEYzpGvY2P4KuJZBH7taLyROFtDrZged
bcCwL2KNbXss18HaCwzZm7ZAHlrmbDtLyLWxczWvSNYlxZ9S8PtRmkTqAszjN8bu
78JglZJc4nKpzXYaJrn1yBTD7C43nVs8L2w0X7fyoUAXEYhgAVxMCsQarWr8bQ3f
shFv/YD+CXqCUImdE0wTqRrb5LUwNy2Z5pcYtF5Ly3atMG3bhzo6AlztszlJOQ2R
y2W2/Hi5pxXQMFuggORwUvcFYnldg37C3mWCnNsA6RBfWDdtpye/03+yGd3uiIiS
SUH1vPimt/Fbdtr1zf2Aswhk5uS8zD9VxRjsucBbIfXp23lH0LE2/KIVHKIGpb26
Ym0Jpf8H/wHLCvQXcpcFJ+P7cRWYZw97ng39FljZiXVJapRZwTHs0H4rTYpL2pxE
BaCs5si9BOHThkxsJrvsrr3l5BkOtvVbOfG0J0UwEjpni20alVnwM2m9QUznxCYE
0yHzDi8N65mQCFnAJzJfQiOBdFafIRAhf7uJnI4niY0JLYm8wsgVrC4HQee6KiRx
N3hLFZUFHYL3+hksSoFJsY4vExwrZoQIJxi8UUaS5lWc1SGk6QSxMTuMrC3sl6YM
EEYtLcRDGnuU9K35GaHJXHxVLZWTpqRQCaUbL4loiywdUXOHjiQJWiCL71+Lq5P5
PSi8etLtwasvYMB6wt2yVw3/SNfFELM1QNm6NkljD+rB66p3zyFTdSuV48nZINLm
Ne6pH8itU1TTqzVx4uLjkVB1MmmTuWo+cGF2JKBR+Sfr+489i4WKivRHIFcVjG6U
7SQVBg1/S7g68GPPqD2rVJuLnM36wwkHNyHcor4UWW0w1PFsdF6gJyXI2v8o17+h
W0DHh3YHJnR0yTxB1pk4T9qpd3em3+Zra6y65MSNog0VofwRWhy71p6DLx0Q4uQS
P/XnXm+aTM+Ob2mwU827JXaTKNjjFqPaRlLEojRLAWUvbobBO3iOT6EAF246n4wI
pcTKyqQi9iJyo2U2qyIpOXIIaedJy622GqUJ6YMT4n593zsndM6r7YS6yewi4C9p
Iq+RJ9312grMGHscMcM0laaTbC/w+rUZiDpmTSmuRTYXqJBI7zvgkfRVfPsx0TXn
E0yw6MdEohLeyx2xr3Z73YYhA2SFEUHzNpVRS8bon8ge3bxcJ+IJeV3v5gQD78JV
rprVhYLd40TS69sSJIR5dWZ39K0IqdxPjkxFZQPeKrpFP8WyRDQDLP0860hR74v2
9kkIvY+ICwQMQe+X6l8gYC2DylKzPVZ1JnTz7aCrvK/c+EFAv9BsX8tLEGpzslhW
f6uvlZkKlx+LeEG6tTzFeRba1M5Uj/PhzsfaQwxiVlS4bYCSv7cKW8wy1NktexlG
7/oDmPaj1Kk1fb9cjB9jiNNVKFrIEqw57hO8RvxGRz3JWVGJi2/AkU9O/C76xf1m
2yk+epo7HKx2heqwWVBsLa4u0tX9xHvImT8IX7L4h+K3Z0a3n8Tw+4zmKJq9vPfp
SVHWsxVTrecHNPYs6ZbUyhJa9EofMCvobkf9wMuaY4j9mi1uWBnZ6fRGsMfUjaYw
CwpQTbCJv+kox9JrWUmbzYAJqGxCgft1AHKWiiofhdSsGuvNHq8NtifWFZH2qnQU
CG5y5k8ekOHHabQtdok2Q8G8ZWaK7Xni/XYwmygnj/jYy9xbcAiu7BEMQn/Ursme
5hR+7LQ8qcWQIDTLEWsJ3eVm/5Q18gJeVVhWy+mTo6b95ycoQyC/67IrSSPOlwRp
PeU/YjG3c11ArKk6fIln80t7JR/QDH1/eltSAJiG0JVTPB9CpHERC+2S50ZBL4RW
+c96d6Bx4XmXzYuJEWp93cth50vxUV8UzahwgSAhkZRCnNXQTycvv9bHAgXKlqyP
oJg8tlZSPuDuis6/5QfBITkj7sDtQWJX6PZlldds8g7Uc7TrIR7MR6Owg7rkTs7t
mJ3/ofjbzaqIwy5PWxOZaB79BjrLxCvfgBIz0nXLMomFCRk8cnTplgfenMEtiF7L
MiwgIvBsSZ2Sjl46BCJNXkWfYG4Y8F9n87qLRF+9jcYx16HxtD87BSuctDsqjGWW
EMxKUTNhF2VF+KpyDB7U8+4N6FRXT+AvnZsrgcafZpuJE3txTqKrzIY+JAW+kA5l
+UQ/cMWplBjLj3EdbmnWtIx/u2IeOWfhVOXvUvzUiDH+oTanreikE8HHWEyTGSoN
YQYT60YwfYGA6owJUtA69UZlkRzSm8uiffdsB6/n0ID+bRIIIVhi0hJAKfJ8otqW
HJfpTiu8NRboYOh7es3fF3AZlv0bsfZ0zTcZyfOqUleOIgc9IaxJCYopcoTdyRQp
N6RekFvyirql+oCpcrveVRyTlavqPDyIAY//KvTUs4b8zuRustsIc1zxR8bOTZFP
IrneffOfzgeJXOvaKQ392pVaq4xwW+Wa395ODd9QpZ2hh2O3U5xvYzoxmxf4/gou
UuWs8VpoOciJlQoZ8tlNwQs85wXL57LwvZGt0mz5/O+e6EC6HkfUjNVFVyY2RMWf
RtK8xVK+njP/ZAB7lAFdQGU18AP0oSTIbFXeLN7hLSosT8DxZJ8yUBmnUq3hUQy2
95qVq28q672AOxFUHlM1p+mSkX4dnyC9T1jDvqdCAUJ6yq8uF7eNtwipo6EkTu/Q
kb9CgG2iXnxPlS6Y9/kCyDjn9y1gPapNQ+ojETlr2sdgkE79Xf7ntiS7jf81DbJg
xlC5anm/hxugDzP7aICIyP2UKxOMJ1NXJRdP5xWZnKjMyGSh6pQzwzV2HjHgmJRt
JiqWFnbz1qw8D5zNIns4P9EHqvUg1RNROjFxsFRbanMbiv5afJYPQafyz7dGsppX
0I5oPLmCieAfqAJUgSovNHrB/hw+B7AobxIIYcpsWtuKjNgc167rPCA8EXt9zp5R
ISdTkgw76kE/bFauH0S+ipFyFnkjBZo9Gix42o/uUuAaelsLy9mlY6VIw7FDbwhj
WxYlg3XE7hTDZdcK/7c4rq4ycEtJTb0i2GwXcHmJkD6GNRU2tT3jycqCU3oRJum1
Pg9EL6gUdx/NoMWSLmyUIYu6AJkoGFsODbj6Exlliv4npJWsTzYlFl8/GM8IyTw3
hopqzuBwlLzfVWsq1KpmhT5wWM3x3gkWxYKcd5R0DgLWvpsBkPSKVe02n+Hhxhrv
kHYfiFs+fXTttMvVxg/rqUoUyOsLhR7dNEaPHluQogfXn4LxkynqmrCSi52pdiXA
PehiLa6vhj7cyh2yJsXPkWf6BxQbhxgTjCYi1QtXgamHooJSAexVFPsKEX9O8nv0
0LKfbwQnpPfSzFeY6yJ9BoqFxOoU+7HTQN3zyf+gGcoJL7bzX0eVlK+feRT5SAjs
kpxjCMppXUFaEQMM4lEdIwROOlvuyH++8MdthexMD7l8VzNFfv6PoKBfelTt58lu
/db8pjAfnPUoFTdVfLNoJd4NUDDVs9TQoFn6/1ndH+VcIPH2fOHWIF7IQbX4lxNX
JIzsuNeuFYaXlduCew/Od06IdL1Ic3XX2DaWD3wH7QsR4qe8CJdiCfCzz+8zXH2a
3hFEt7/iY5TUztxGA2Qhjbr0eQYIdcIXKQGKdixLWBN1qmVv5fByTAXlFLzYyU2C
+nzUyZls1tjo9ZTE/BKKQ7cwInsyHo++bVZWhmGFQQhMpevYGd+rKEvzrZsSC7tC
2Mt3Gp7KCJYIP4MIjNiodHKdKmE/jHLoubADPn1sQp8q1cA1f7MEUo4rSkPjt9KI
/AmXk0RQ8GvPNxyNbxNZKuxUY3levMpbN9iuItz77az6VUVyZB10Mv1iGzRDTXjw
eP7ykKXnoUzQQblwOXaiKKNQoWvD3GWFu5l03hxSpOT+KW5H4QdkP+CHbEEFOAeX
oCBWKBgEZdvNq8nL5fb2kXEInery+Z3qlBpGXS5DZGZ8GW82G4vJPPpmPIgSdWfb
i+NcNz/rODLShUqUd0FQMYoxJLDKH32HWflh+y7ZtMixB6KXg0SgGN78Oi0kLXMy
bq8hmAnB0iz2v+VYlFG+z7nCAOww8PhQBzf1aZl2/y4pG3S/pAg9dGRkxhMRsRjb
LCX7SMJFAiBTrucGvlkeh5enJX/Lz9fYuEQMRaem6bOKgCzAu66ah+9GNM9vbwS+
nOtwHqOAMlJykaf7vXSowdL2X37JyDK7nWXnlecSEjL0Wkg47KsKqiKU0QjEa4HC
AheBFKaml43tJ2yZI0AuGfTPah/vMgczBmC4+3dxYQ2ySOjmke4WpYB6OWcqUMji
xVlcquCUlo9SMmdNKJ/7TKVZMjx0gIAf18zJJpvQ9kQofpsdZf0ZjwkNCdY5W3iY
LDh3+X/MIRQoIWWDopbb5+nE8VqrUiHHXRhrspDgbm92pWHZxvI/ZvRBCnw1iywK
EEW9crjt5F3eTNASP6WPBfS3pOQYD/8Z83fs7xrcfmhDLh5MiLSSxEaHWQkgN4A7
ZbI6uaDweJ6+HZ1SUQ1tlXjh5FN0zderCCjONDnc7Bkdg3JqMx6j8Gm7D5oGSsLC
poiIa7R2p9JW7myV+5be3I43I49QDEqMiRgir7fnNKDuIOnMkOhq3wWNgcV5slHa
B1PqjoZ6h6yqn4xGJa2jRfYItmGYo2SAQpIxfr4NfYAjbOfV3OjlXkKmzKGfKpG/
USNO8n+xyoCJ9INqCss9VjnCt/O/gaoIrvNCSLfkRxcohML261eW1tqCaGoasg4t
vZIb2oJEegIZUIrWNCNqXsD3IbGpfpm+6S3aTXhSw6/SNgurbmvCzq6+iSzbaIuT
KtCRBYH/8pDuWE/9j3cyEtuMmZGndh3id+BU84v3HPQeoq9moDJd4qF2FU3TY60U
rS8ehoCTr5/UrJ2bJPVkhZtZp98BLYfybaNM9YwupFeh2difRMq3Xw1061qfn46v
zn5Q39fpfPAV9kl94/SmB4Yw3sH2NRvAYCqB28kN/18cqRzy8GpX+xWw8W7d8YlU
jHLfZ9fh9A18GPU8y385B8dPZ3CnAt2i+h+0nd3ODF4xefhsY8d4euGVKA/uHRT5
ohcB14rb6b5xjbO8YCwMWxCXuMXzAV/wRMnIlOJ9jPg45ytLFEDyKNwRaEaXAOLO
JW2BR5T0qFVE8ltU1XSIdcKBBU30DkVshrbEkPw3RyO6/LMqEbFEIlE+kveQBc/w
JuTkVbUdqsWOvuApdtP+egKnuVY4TSUPL1AMTPLa9omlGILYhp1HFHFwmtkR6qi/
Qn7Xtb7b+mrIdSZq48JMn65a71j+xO72N0b1JBxDGerrOOtb5UsZgtRCK/Hp8Hc5
saW327Y+nR0kTanXSqWvx75Yuhdh23pLoxGX3MnRD9WwSwfWvb+UNiNMC16F29r/
vl+CakYV6688ElfsiPKh+8q+23+b92xNBiqHU6Po1AYjnLHk/80E0o3xn08KovJR
LUUr8nxZ0wff6jUH+aikcsvqKg/pkPyqyq5aXRSTPXv4IQRPl11hJfg90SBM/EG4
DPPiae4lwDHrkLJTDo19v9cJF2d8chNW/NH0XDYPOKv5iEYFzgpsjG48QOSxLu6M
SyI25vGyzlrgTfMzpkUg3Osl5p0gncVdTWc60WA/UlBOZCz9IZSqBSxAQ+yh3jai
ZWwvbTlAuQyd6m3k5GNEp1A0xf+SvVmhl9o7BFmWmHoC1RFPf8WxH74enSbZEH6O
Iz/SjqaNbZH3dEr0KQmT/CACRdFAbBLTyStRwcIKh/UlTC7zukZMpmDDorNIMevZ
VxP2X23bbRJ5nw1WxWtOuRRRaiYRzBfEtzJ68Sh85FSa+3mp1VmnIpQ+H4diVkR7
L/hUKcRTRYCbAqiymtp9z1OvyVQ6ys4XP/i/NiCcEk1ILTfoYS0kiLLhGm0PoAI3
E69dwyLbpSaQoJ5Mqt4YLfUkRAncwu47JsAP50IC3xvUU/xm+IOWWKoLi0ByJyEZ
kqZWo0Ai4PWQc/wmrG3u0ugqO0HvJJSMmzyoUJqAngQPJBQ0BvZuSZrHlogmdd+f
XUOkhlhvWfZ5Y+WsWXcWIH9zhksiMLgGdGj536h8uoPmhYgbk/j1NyU+NmlD/th/
0yru3MjG254lCodQRozi6vRWXjuVwXW8InnwMKieeokVyMOLn7Tov37PPNs39eFo
eXl0J+W5jYD3Q2rVT92RPVfyV7yR9u38TX6PTYPeX3H+XQlx6V0b0Ctye713pjPu
/nXJLf+i7zAVWdPDQH7/sf1GOgn+mNGGoecE6kVoKOnH4aLHy1doqOM4gE3JKCpE
xLUJm1PdTbo4ry8xATn0X66ghuRNNOnn2Pr6jMlP0YYBeMtYrcHdKXoR9Q8dHPtP
nn5L7h2u7k6Ykixnd/jF4O1IIxa4tGGfKiyqEijrazLcZlDm8/3mb5Ef9gBoapSJ
2EIVmF5Lm1iQkqRG5DDWomxB6R+MhPkElCUI79shW93l798DYrpIYHgR0rhdedGI
cohUBmGcoU2vJOOwANKSaWSd1n4I4BAxPFEGHtApyMxBPpJqMPPqQxCoLQRjN2jy
2lAfMlRN9dMSmVWA05PK6/HS0NAxGLznrjK5NnqNOMvfixMVD8dEHVhHoOXWQR5N
7LcBrAuxGNg/2sOlk71k4EUBK9M/donFWQs/1LOiyxpn4oeYMxfNYSSETfKlxINd
kCzGuxGWPbjvCrSyWwVMofN2xwDXR4zi+N4/zOCeURdiWCPFC7d7s7rU9BSquVqd
xPWLeRbQ1Ll0UsDZbYMsLDVRMTByvZPg8+LgOpRbbM7kgM4aLuEJQd7NPhzxqv0l
q+wb6nBrWZ3LBblXOCps7wFVpK1iF13ova9oStf2S6pnKxRhWrGpav92QCYi0DxY
NDoaCScmrENX7z4dcpTOfmZ5L2AZ5UubdUDkpj8VaPPqI28WM9CsQYvN01NQZrNO
9Znmmo5OXYAm6JkriTTr4NBe7FYYsqEzzOIFkOZZF8kMmt04UAI3Kpw4+4Ss2WQA
EwjgEwFRlCwutBRRK3ARW5AxjNbfTZW1AfhJzFxI8axaKKRpOuAGVYHam9qhu1PM
2ytcOgAbCPxlFVn3BumfPDACH1bjCdWhHK7oVf6px9/hGLQt+gQxQWkaSRl2Ljgr
eE10LtDkvysI7BmcuIXJBPJsi8wgOu1saZdRXMmD8fBFFz+g+py2RaetnZvNsHAI
uQuchkhGdeFcN8mtjm2xp7b+LkxFhejQBIDQ4nR01z80nfPKj7I+OQ69b8+LpEJx
6cqD3hsQkPc/tdclgpDP5SaGeT+YFTXOZAjYRfnYTk5KJHlfgH7CCz10nQA4ELRv
FNiFQHgfxPccQoZGhVjjEgTcpBTQ0dA3c3VOGGNOSa/LxKn1ac2QKgvX1thju++u
OwFYc3IjWIdnHwqPVnI4aJoV5xDSq4Wg4faZEmrCiXkYQ3l6aB52yCtDilql2ygV
J24CDAFPQoBBzghHlH3oYfPAS9v10sMeA2HVJISI8OBxPtd/HrG1EnebfPhgiwgi
FNGBMIL+OGacSMvLOtnOz1JFtyUm9ZGrcdQUKzzfEDrhpMw27lwhAnBtSEoELPxO
XyPMmWnF5cPWDtWibGHEmZ46WDh7avmgO1SKurz9H+Ro1d9v4L1ERYhf6893qtTg
6scbmSa1BbWfXs45A5KRtuj5eJZaPedz3tIggQFS+bzYO2UF4o25qtBG2NJvzhsK
YOK1uldtcXs2sKJgxnFbezqB6ZzindatcAnR3p9n64AgxmIzEv7hNhiFhjojBH1V
5orBH5Ywu6V9CWmx9waXr2VEU2STvxHZJjq+I4JLJpvw7i6kbdrKzPq8te4EnHd7
OJQrrYQ5QMgSrpix2//aFdcQubBlShyoHvSyRfGUSK8K/yisbiZm0xP/YpWPFzm0
nnOHlQfkgJIE5Yct6Lu5RZe5cUj2oyAjVXelQtbQcX/KXSbDfFU/k/9z7q4UfE2a
PG3WLrITNkgubhiP818KxekYITFt5nmisac4rmSehs9DVh8eT6WcMfb9js9ZEEeG
QDqRfDJ8VJGxcTYI7av2yaUvRxmrV6yrY/sS9gqVzqcbQ4d7OXyYmoxXA1KtaC7b
tERkRS7WhHZOMOywzqZ0YOUcjPHV21+qJ64zn7C8r2aAZFae6YnNM7ieIzqsEVTy
wpRmi3YinCjxPYTTeVcKkDRe0w6sRmg4YRIoCLWeB94hwDVOEQFMeFRDqL1ORRcU
HmP+TSj/lx2SI3ytT/4EBxurMpW8SbSXbJmziC9eZzb0/AA3DFAbI0Pp0UqQpf0o
CJogu4Co3jHFWZmbL1gU7xUJAXUsLMpux0RzvEVmOZ8tf5lOSTmLyiVoHKZyABaH
JF6uoAM7GZtN7mxT5DtEJfUGNNp0k+Z50CKl5dIjz/BGREpdsoYfK0bG4M5fQuzO
xMV0SZt4m9ChDg7kGCSyMH0v8bIXgxOsRTB4MI8u3dpjBPHIYbvz7m6CO3hszfm+
VYFD+IX6sA6GFYDc62jckyjSkSq7LIYxBYyItC/8NALEeJ6U6qhf3jFDrec0oX8j
Ql8PsX6BKfPf8V9vd73KN60B2So+m7QlN74FVqE8eUGE3mho4kNdZj7DjjScFxfh
UTiaYPtCNr7OhW7ElJsDxfKAyUoDP1v3yTd9StDefFcXcK2rCGNSjjnxfGJjKjOG
GGKJc4XOlBVlVTFsX6xNM39E6biwmuAeYIt990khwR+mU34bQMzadu3Gz4OZ63x9
VrQv+aqNjcvhhjaaK/jGJETtFjgSIgpckWHhmEjreykq3u1kLdK8180arJZBwmIt
qNMBihimsjli38fGxF1HDujZ5eas8HQrppXm0w73e3VCqzidE8I4AzWvLB9+wuDc
84wngDHeCY5yMsU40ez3bM8MVroR677OZHdX1Whrvxi87IcwAhkVpfn+FZphYa4Y
7nvMqNEhPyvvW7j6LIpWaZntxMSmvynMLBqMMjPgeqHLg/6G1efeMKRyzcsWeJ3N
+uNqd6d1jLxmivfSjJ8xvDYGOqds8xM0binPDby5OFETtt3/xHRRICcqRgrJJDnf
OVmnG3FKTLXtvwGd/DSQnsLWUMQ9ts/qZpEJQWfetTlh5BED50Xq+58PCW/PYBUG
CjMcOQCUDHmuwrOhNfLVCmEThjWGEEnbqdGwez1jnh3o0p1Qlgpk7QUcHBhUAHWD
IEaXNaI1hTWJTkKUQBPyNU/jA+0M9H9POaT63sIBuEhXFADGkgBUf6VpxKLtsbxG
ybqu7GtTxcRvS18YETk0eg8+Hc9EtfSS2o1YiCiPLZ4xOb+AVnBG/ZMB3CTgkvNo
j1adKJUUf8AYD6UD217JYTd+w24bw038gOZl5qgXUIR+veM72anGHzxjuU6L/5qT
ncpk3ZvhW6m/W23TU2t1baUcUs+z2ES7pJnrjWI14P2Y+bKnovLTCaVzeVCnaHO4
blQESqLu4g1fH3PomCFBLTf8hImVB3vvMfiEOGzbDFEADrrm81hsAz5fxFNGoFu1
8Pdeyt43fd0GVy4B1A1AyJgF3uCjH5/o8Ts2ea1E/gH1Y77E7Al23yqs//Dey4JM
L3DBOcYamBV5mo8oDPurObsxomPrOLcuHJ1vWlY2XpAVrA53up53bH2jU+O7zAYw
6ZU1WEG97QPSckZpfrrAQ3FWhQfbf3n+irsfbHmNWFsud6UbeWlXgDuyYc7zR7EC
WYqBTA2npeKxnzeZV9ctsaIjQq4mJvwjAexj9Dkm3WPfn931glnIEuS73SwunhZ9
sSaSSc5ACpjRKXpcN/0WSu7FX2itJB/+/z+vnOpJaOrWmsl4z3mImf7P/vJigyz2
qi5In999k8zSezm7ANwMR5RRACe0ttprqoGxN90ZNB/HqOP/GauqyQ0a8jQa4T2X
adn4OsSHK4l4ppkrqxzZTShz59A02Lhm5QjcWgYEKr/8BxZ1p9+IoYWuWBTVA/r3
4QtJ1Dg7zZm674uW19KM1CIRefsvWV0A6pXcSv0uGEqsn5ypgT4a7lSgtO4HzFa8
0sgitPPoZg2LdQi9sAiNXm2hDlme4vLnxdFXu91uZmAiJaTxI5C3FFmxtcNiNpjc
pYjDBGrDlIClkvsNneL4sCGRI2iiY2tdxPyPcg0oas0nenq9CJ2KcK4GCXKX/3e1
2z3pzw0nDI6JvcOWxtC1tp6dzWLUwCYZMU1WHiZ0Ht0JY1iF2PJbKdh9MLAHsSGZ
5bkdc5IlqvaoLOLbT4ASBJ0OAi+buJGARtQBPnaM/RFOjYHjfprHnOjTMutioSQh
wmZ1SwuQDloekNwBeaNOShtNWhHhdrmwCxTA09jJfPMtmAbNlJFBPe5jXKAlqZXS
qG+Ap1AkzX4ls9W3cGiVlYGNDIhTx6cSiox5413zD+weUelvLH3GOp/jyk1Z6Fy1
z81ZwY2NjDm2bkMLNoX5wicucul5p0BYHcKBoeg5QKlef99n1RLQJlbzeKsKGqC+
Di7Df0nsb691hza+Tcq3mruQYAl2JI2oXWZRGnSEbJFQwzN7w0yNxCNT5c/LpSjo
iV6k6n7yAW+FhQIPceXfYtNdmWftInRfzbCrfDW8/6pzQeLDg2qDVwaKxDq/FPPw
K+8ZrHUz78NwtE/F7+PlkV0Hxy6EJioVwrcu+8gT6yv2h2DNq7vZDlGWQgrVxld/
2JzUNmjenEiO3ukzEal0SBTxtEvHh68hG3EqGOsuQHG/AyU0AffLjXi+DXgaw9gy
nzYCtRK/nGLaNai+FdMTwKpQdi+rxzB4csps/KPhuk7K0+c+rjbNYiwMf1MXTFUZ
XqbnVzo9p7jXoFNjthD7Pn+vyitg9F5z4WrOm5PSYENXmR1G1Ih3cYFaaLEdF8fB
j4Pg3KW/z9yYnKRcMj+9mgJhLkJ8EBzQX+oZuvLV1xM7jmvpCfJAmM53V/kM6UbD
w9v/BZLVkzu86Fy0dcCi8Bper7oYLCxj+xeamfUnio+VKjTQB9wYNncFERoH0U8f
XmR9Hh5gR7dfaQZ3IerX7D4d4rrR6j8ySzuzoX0yzZd+aWk3HFqjyXPMq1GPUEVy
+gqgBDURuGGjJ6l0uNzbHf9N5gPnDAZ0qSD2Azv+cnchPPQXSQai6B4HlMm6qSMu
i4JZIaKvDnVyQqIylivkzO45GWQ03BHXT7/9XGhaEk+t1IihE8SKe24F1a9IlepB
QbYCKaBJaENJgvTi3KDtxPw6m2qPzhkAnqJhKSmNKCwv/cdd2KXtFz6pcRs964wc
05OF3VS2R9jhjCx7L1bC6N/nVu/kkxeJXCVjnyOfZgaK/ct8sS/MUbZwI4az70wq
rvoTGBUDTTM3DdHqKBPMqP+9JrhUdQOjVcevxzxd7h4NW9VZjn4I/ylbhzk8q3BK
Y07kyX2pOEAT4wYpQp94huDNYB3IRecmNjj3CX+VxLupwNgWaeMfNDEgK2EMrQwN
vXgoP7osfmzUWHAtKuNA5icFocVwqvnHZDHVWqN29e+lvPjeuTiDNhMfrIoPsbVJ
zFKxiUIc0pv3z2exyQNeuc6lQPiafF45HsTShEfdOTkhxxeRmXDhrGruhE/cJz82
i0ydz9GNbbODe0J1XDNsZMRiOKtOAx6vWL8l9qFMR/IkcMXehAYnE443v+ik9sJf
mn5qQ61zLZH5pknSRvwBpbMV4mWZFP8dXF6LRHXAO00oak9+gIow4HCXc5WJPppB
7FE0wroEpl/BR1XK0OTl07QN9R5zsjmLIza6mv2ZsHcI0Nekc2xuwARiNSVBaU/W
6eoDJB8PrJRGDGaBJqDu2eKpQqAF1gcMLTG1mE15HiZNNwl3dZiH7Cp4vqeqm49Z
6xOblyuufYaYFF0M+7LX3XhXjTPu56vT2gJIqtEjwyWtZxKP8MvO+CiT+rMGsq7v
Dbya7waB8wK9/iz2ToNUqV+2zj329fmTDsdpOKk/8MbpAaafvcTNdXuNQWQsVv6r
uIB0iFjldYcigK1LTbQ+0J5hapbrhFpv+GkHW32pTquH9Bnv6kg1kKsQp+F4WtDs
0AK/AGTXPGIRMoGFKdYHDjyeGWtujtf1ONLMAl8qo8yvOVaAf0ww1Tyi/paRA5bq
U4ZcqCXVQnw4QjV8poEUSFfWmAwb3A1yw3dwTx24jF//H7IR1V6iXI1IVDyVppkm
5+gb8FInDY0FrZU2uwuvGUNuCuLx+LQYHI2tYLpZyQSOhMzkxS+1Ea8tdyV+TeAK
2fqtnD5C5N9ZFLvuNrUsZk+96HJUXyBIj+VrtGcpo0kK6WMkDXWrh2oJSKC8AII6
P6PX5ij6MDQ30FBn9aXNMEXHmzyQGWew4wnCTfaS8KlAu6vyudTpnRXhAmEubgQa
0rMDMZSCX64WCIXAxmmpfx10LWqyCiq/ZvnWkzm+QQzSGOEq0FwUQoKr3V/2/MaG
lWUQLIe3UR9I67CslqredPhqhIH3rpJeXfDHVLmMzmjaWtGZXQXHLy6riYgrPYfe
PfbkeeMyjL91xjtjPiID4831dnO2T319EO04eptMYUL+AjxRLe/22C+JmFBMXn+r
fBy7d4i/9kPe+vzago1XR+Qhy8fBpsU2KjNxbU3S4Uf3Qy5Ct6dB13rL25It664K
6ZHRCODQ5rFC0hqAB9MttgifcXuhlVQUQYgviLBOUktwmeNOrR6r9BnlX3d125mA
7PqkKzBvVxdcYoErDFAHxQErbeUT3Aq6Z8ZQj16eguh21N88GF6+WpaMsnebuV0d
Y5/C2plMaGtar9ELSVCF6ghVKw0EsapceL0vCc+nw58xOdN8D6LVPRR+5SKkk5AT
iX71uY+A6HfoAFMTIjRolJb5FLpgN1y2/wBkPFJzeknYy6p/u6pjjvuM8mjRjwID
kvwUhe1kswc5Xxt91LLTBn+TuWJ9/xCLg5QrLK3vaZk5IF/pIejvMIBzftv0QnXH
En6FA/C3xgTUjfVnpDq4Q8oO0hmM4iihpHRC09vFASQu6zn2jxoCRFigIMi5I+xt
hHdsOIyIKtKw2zz/GXXXrxAemgaBtEhn0gT9JNO+mImkSTjJ1vC8z3uPKyn3nIjH
fXKxRV1kGxdGcnjD5xuED+gkj01cF1W+eHqxtPwRqlNCo0kRaFZp/cpCDtd7pj1i
/rAP3jvPOJGfmZ4VDNLn6OGfZfdnvjgHH71bEicGULl7qV3qOG7O8ONKhnW9t/6L
Gklc+4HICRe2Bz09mToFYpOU5DEShPwa3bwlGxIIr2DrfD7tC3ECxxdt9oe6wNDz
Dk6nJnRQSI4NcTE7AcJlYna4L/dpzzjWOwwHO6oernbSTWlIZhaACRVCoCBs0GQQ
4mOx8YLXtB/EqU1JZWVV9lh396gERU78/k411VFKUDbEgqA/5a6nGMVyncgu22pW
tUE+75X0c3i8elDucuoyXPrnDB+w/YIzmXKjnLDnKcckv4wFv33VfMNzQpbS5Is2
LOLd7toD5khaCTwfvmpdHfq0MOzAHSeT/00LMwPIVs0xsB1v2SeK0CbZmRsNoogE
2qHBySarzVAJFHuUIVkxqn3WgIW5cYPbWn4/5kKcOHDdEmht0R+Cz2JtHDUdse25
VOp+AEBH9XXQDMXnXi/2BvJvIH/AQst+11if3HiFT9x6EdId7uQm+lrwCmDMquKM
+72LCvcfm/ba6KWLaSLy7V2guY5y3IOfTkzwExJlowSPhcbxlYH24zjLJdAkyU0n
hPMu5FWkRqFXd39TcH4SBOVpu1vBj8Hnh5FUKizPn7J99ZGjFGEUTfRkxjYFb2W1
nPCDTvNXnUhxN6VU+an4IQY4Axzk5RSw1ko1F81vm8P5fpAT/iRQvi4PngqDpLGn
q3gRVElCvC6yN6wJQp9VSxIhH6LrTFJVECcyRE1C67QnilLRJHFGlWUlIyjSeoee
7BlfYsTo9Gec/vZbkP0gclEVHA+EZFiL4T78JX4MudQQZQGdg3DVXS1e2VON+2cy
hCCwrKQnRJV0YZvwygXhDxxKGNx5He4m9c0KkvQ2BPpzTSBBShtobRQz+ogkRDM8
sX7lgbT8RSwAqYIh66O9HRBQEhlQk3rbEAP0wOBpgshp2EKIseUZSUkyCZuXXgh4
ykkc/e52M6U4MJs7tHcvD0/sdHhhRfLEBoeKT1ehxHloa7T0Lnp+70hohq8ijFxh
eaHYU+tH4wij/0VvZh2Ek8gXpjViwNBOeoKxldsN2AofJmRXuW9VPj5td9aJuG22
jzuS53jufS9mU7NzRaKf7/pUy+bXyNw91tbhHf8xlzix8WOxF2FbDPoBmSATWiYq
/OmQ252FuzN9B2qHsP1lBaMbj1EkooTe8EfGlyaw5HmPOP/FKBymg4YJSTeSRddo
pnuToauwjhpsbxWf4pUbUSlMkgU2/wzqqNW9gp5b3h3FV7R2pxmiLOKhd6aNrZF/
c83gO03pZY1opvcLXt1pILh5xwgkWn4WMGsj+ETm/sJVTDiWqVjF0yYTkvo/L1A7
I5Jt4ddDWseOuJ95IJ/bPKEPo5gmavS/dhoFw02Y++WpBBfCcldp5q37XzkJQZhS
cimgLMmYo3ALhjsCa/Mi2XTW7zj3wN/KUF9j+yDIOVb53na4gBrB/5LIys+SwTjD
noov4pEFgPNi6ucOskHESnkGn0Q2QHJraeF70TZ876ALqKuv7yjmPz6olPXVLBIM
EY2NPSd3Frpnv5/4Xrfu7abXpUjHxRYVu7ZgMDqnsL0n7mkMN3mZhMVwxEai8tkp
fQ8xa4ug7EiKtEaawOpbWIG3kAA1deVx/YXgFkpQcAMdAmu8bozIMf/smUbogxjF
9nnNYfVXw4a7/wkr9DuW8RzKpZN0Txo1ZXWVxJseQJrH6I+lu5Hoewsv9cei1xgU
kU2QMrHydxoY/ODuZQyVMakXzVXkdE1lBPQVznFvq4VGySHlg5g8TxBwy1oFIZc7
7hMtzBvqc43peAG4wJ9Sd5LZ21zh3eXKo7ginUuaG7Q2b3jPL+M6ZVpKk9bBv1oy
NuZgJj/NdVgVxsTr1idp++zxCqd6GL9nn8skFih66AqJIc0aX/YTrGm6SsMNI1fj
RQYwuRaiRsW4x1ZNeujH5AXbiXVwBK5rqZktIyjIOUdkIbpdz5w57N6Bx0j4WQ9Y
fspf6MkN9zbJXTiEi/0tuB28KQh3h96h7VKFym5uAaLBSPiQpYvJ1HBHgTXhGY5k
8tLQ0UDKSNqctr32wnII1GL5uV2tWr0Ah54BOmoPPwwICWDE9HZFY4naQ8+mJuzD
mKQU1nUmJkOI4CFv6rQHM/yJubyeGMC9b/CYA0s7uLskiOiE8DEUfG/pz049AwS3
yp8pWQ02hfTBy+5JsTFTJMAgKlst8GC6XGcSQkIjITiTGX4H5EBS/L5BkPsyMkH3
Nt6uELKCDs2Zot7ISCZBVlI1Y6YbN2q9FJbRzgfkXT0aoYprMn1W+LBH0HUclPG+
HU6Ag62oKX7u8n7opScaH+KmNp0N9qZI9k3+IOyUJLwNrn1FKqRRwCxbuiW9bjlx
5jRaTgqZ8gvUdf1iTJMM8Cz4rVmT+SuoIEULpd9qD978TYHU3b4n5WAext1OYIkC
LFZPaaflZsa/lf0INi4oZdqGRLd9+61STD1G89teViNg3tyFrFL2iKEboXXN1R9a
0IwScXjjInPc0t8XQ/i7CudxorW8gICxknaw1FZXhYoCfmUdgvXCCOL55SKpsmYN
MrTS7lvzkLmPZlWNDKtzzzj816/0RkCJ9dE+XDg5pY2uwV9VZLwKwGjS7c9ukJ1A
KSljC78fl4gd0yKmCnVJWlu2DeP8y6swMWUJWC21uc4dV2f5RjvlTkKKtR8GIJD/
qoQHm4Az27azQtjwhEbmbeni7nIH+7eKO6fKHsJsU/ccgKdD7GMnXEHPm53IW3LR
Orp0YVY0gzqTi48TEabUgSIY9fn0fQlWR0KYEnWFzxiHFLe0uXEjKMzaxxgNcX9+
QY6Av9uH8VC9R4nVQ7kxFx4Bg1rUWRoZYMfJonqIxBspxbYzZKYdaMRCD3pexbot
y4c8Cst7YPT87i+IoRKKl9Alp6XqmeX75s/MjP6uZvXDxG+ocVKKDNA6SZGekr1U
EEAD3LEYJc9PC5QlwR6uaO3PejMu6k8iasouc7Q2n5hrvxx1TU1nF03PELKx8yUX
6ongsQaXOz+zM3sNfKGj1Q3KaRbGhA1WkKHP3Rx8W1LgSI3kxcScCs5nDZxeAvLj
zlrXx7RDvG35G0fjuZ8gGVxSCn9eFdF8MT1+19tWnalGbxuRaA8crSdzE8A/P/lA
nKS95mhq/V/tVcCCxjShmYZRVdjt0nYH1gv3Vm5K9DuxGflgLybyELE25bZ8l3fF
lWkVneruQYzJhuU051zw0tlWaBg1qvE5OOeFBSO7l2kXMEbF7781jM7dyjWuzWx6
grodNLw9mZ64o2x6udPxZ7nSBk7Ltw8DGqFL9IHtzJWOKKnkYhcHgBr2JBqUubXn
BdLDVx9bQBbRQ598CZBZ5osp3ODcx6TliAdHbb8camjAsNW1NpGNkXtNyUBBCnNP
2gB/5s1KX/QaHKZgahnLJpx4h3DKDpzwE9VW82U8Ckn5ovV6zzduXmQR0Sbgx4IA
JqP/A+bex5QZ7crQ7zaEWWhjZYSw2W3Kvt4IW9I3F+Td9iTw2fdyW2QYzd27TGMr
ypgqIRDNXlbsWP71E44HdT1YgU0xxs30X5NeTN1Y/ofY63Bgci91a1hcuiEjrnwA
5gM2BrgTL4KzUngg+weurZyDtUqQIXfTaYrxHYGGE+nD91xBmJ2xuRZKvkrElLEq
axpktGVWCJNEMJysnAO6UAXOJn/h4JE+FrZxaSqlPlFeZF4zlvSBa3f2uLh44/eD
gQb7VToy9qxsTBD4HBbInH/6A0UVjoO6V3lATFXvFw3oez2bDCQjMO/xBLPKCsf/
IonfdpKm5470RZ/Y0ahWuHzv1uwzbTqZXTykgvuSUbN4orliV4LntoeOClVuG7eX
ZGCOk+gFVK/NTU1529Ghwbr9xV/aCWWAb29Pvs97O7ItrqCQxBwwaAr1Bu6VoAKY
cSUEr27BJuA4kd8QgC/6WKCNia62FTruE9ncEfSdxXZr1rigZMHhXOaun+goMM84
0a6anR7yoEvb8w30JyxIpMcFLELPKkowg8yhUE75QpfqRVCLJvqipTMpzct62CoY
A7dNdhGP5TbmAaA6qKGCDy1H87OpUHQGw+aoosL1jnXp/iFj2dPa3G1lD+1tvq1v
A0VwDrpzo4JFkylcuNLvOwcxxj1qMRKx3HekT8/JDbCIeYdOKS4aX8OTZD9fD12/
mW2jcO5bG0Cvj29SyhHjYrVl8Rmte4AdGUs7u4ZYe5rB99jyYZoz/rCrFMEcKOK7
kJY4L6He/NliptWOoKQ7/elWRh9A9qYcX21dex/lL1v4bTbXmqzkT7Jtcflu7w+t
y9nAOhCZ8sktED/X4mRgSLFcdnCg9Yfpap2W0Ou1gjf8eNB6ycJmpuPD8F42SPhT
kODOm6bg0y0Ot9qiZDjTSUZBjY2GyduaEYCKP57dVVwKozXAUy9p833WiZ85bw9b
WCdT/JBM6mPPxS7/Z4+4/ZJZ7lKz1rjkofC7MtH+Enc+pfx0W2OKQdkCEb06810X
L6W/86+w96LKCcwVt/tjT2GAIuMeDAezhviHWMur7rfeEUnlTS/52oCGFx//v2mV
yeC9/LbIvzky9WVkhDcRX67GANGHrBZ4aeJw6bUxLdhKUHF53M5U0hAl4WD7JWGR
F01Uljpv4Ki+iEQ4MEshxuMk+ugqAcWNyBqb7JwJ+9a4ouquW2YzmzuDb1sAawfS
MZpy63I4uiKFmTogWCiou4palaCqlJG8pkL/YAPcmwbY5WDltI69JcRqOvp2NFUI
OJnwdETuv8MyBYcpm89tdJXH9TMpr8s3YN/Ca3Yf4xWEyE7xdt0dk0ZsxLp8Hnzo
GslxU8fzAFduu6b+6gP1EHRt7Jfa4PXSl+3KNSHJoK9oHcHFz3MI7xNRh8uoGJJC
M8eZXPhkWTdh7gAES7nADTmfwm/XtXIQ8KDTYjeKjz/dP0PEQKqX7oM1yqFbLmPA
AYnjYgSJh7Agg7D/o39jvoyuH+z7i4qp2uGss65/NH5cKdG24+roa01Zr/Rusq8w
CMNyluaC0osf0TPkxmejSTFzCfVIIihxG8rhy4ARaahNFKgP9O6pP8XXoOj2vYuO
SG7k9Yq7IKPLuQrd/tBLp+EJYPsGyKrFnOCgEj1uMzXIjSt3xFx76DE3GTpdtxp2
eYuMMxWMFUZtPlHVNuUI9RGltVnzKB6DF66MadJaqtymSimiPGHDC4VwYoeXuU0v
P/VROE3fweuFF3zcVvwD8a5MbmX4q/Zj8o1oUumsAKxPtYIyjAHSYk9cnBU+G5qo
9z8g18X7GXnG5S5wWSXhpy8D/w5KZSTTm8m8dVkQRrQDLJ4om+KkGLky/sT/coIm
btxnnD99hp6eILvUTZ45ho9Vuoi2ApfRF2E9Vjh6vNxNHlrBMN8Ri2RHiHUvLrfs
+2Zr6YhyNsmyvrzfPcX3PeGdIeUmqI0q0BUQHCS/WZlyWM8O+rNBOK24rRdDMqWa
+bU5F0gJpJgnIYFkGxM9ZUokcYCpss/hmSWkIzfjx32f6j1r8JVXyXjLUAAPUzrW
dW/wyRIU0oKJvAx0vONKu8kyXTPcxX4R4WZRdZlzI5QzY95qh0mIIswmxMA0ko7s
pbv8C7iXuBeBlo4yMn8ZGw2Ehkdk9kqaMDyL/dWR8/3ec2vdZcTjRlConRRJ35NG
K+xq0+sJty6IMP0odUKOiztHsqcXybjJEcaGFbhxLHkxOKl7W99+PIcVzr+Dl+/2
DL7ywnSHebr0DosHBnjVCk1aQiHLJkfEi4WJAZOIp2Ywvd4VKNjVjbW+4wUs/N7v
GO/6wfqRh2BHSs2CuOsIOWQy3hjqakyXKHrSdGRKyUTjqZkzZChoEt946KBPwziB
gAXF+4uTpubJZ8ngwbvKHc9B9CmBjCrFrvntZzNknx9L1MxW+1ieYWWViN/n2WBn
P10aRULpboBFHO/sOlPrJkl+a7wrpJLqRtyC0Fa7RJDYVmqTaXwPygUglibNQSHL
FZ6JvLQDAUhcYFGQR9rbghcjEAIy8+LUk26qjvOlRvlYo17LzOEorNyE33+pwDXV
cMZ0wyneKCbzLmDO/pzlUwJFQwGT0nLvZZOzHNheQR2A+SlyI/W0JyUL82hM+TJR
9+7aFz6qz3872T19OAxs9WewwNE8YNhzsCMmLFlUpRs8zHDwwdb15MD7NPAhMPyr
EHRjnn+H8SitVgK2GiTSjmDB0zsBt7GcLY+OiUCMqjJ766gMeKCHvl6zMuazshD5
ormXabH2/ZNL1aEAm5swieqG+HgGDyekFuBffkDYGkkVIt8qBlz6qRQferuHljBf
IkjTzADJs+jS0JXjD2hnNfh7gHoJ7Fr+I41OrvUJGbMERkeCeIGEzAJT0Ncmu/Gi
54R0eC72yF7zuJ8+IN7iJlbRBrsonKq/ML54vc5i8dOtMxzwHy3zyU1E9DQNg99v
c9ARWE0Miu4NNkuSqA7Dccj9gfETu5monEBhtazK3wBmhX7oXadxZ3aMnoXU+UU8
VfTgUH7FujoGVjp9GJt/0SGadYUllxN3UagtIQTatnCeaC2sjHfHHWQT40DYi8yT
Vtajh1nDJGOt5pensJXHbrSNnH9a71t45jV50aQ/NWC7bjH3aSlb5f1JfbAoZVuV
IMhgjfsTUlv4mFiKKTq6LE8/NOYgtDINwQSktrI1mg0oY7ztEubMdm+SU475yawG
cYawkrHiilPzQN1Ayoabq7x5BnZY0ueuFXk2ad5iZnHFLCVVykOLkGo14h5qSEH1
ummNolwYnd/yI9guKbvVyr3EY1gRPscAp1cskiIzNyzm0OM3M0zdSBSeM3bwaDZx
IfmgdbyLY6IzMZMNAx7YtoDnNByF5hP0YJsGmWiiqD2k6SMSdy2D3FvqRRhMLIGF
EHhePmicEl4pN+wBf+uUdoSJGLydS3DQWG8niesZVsNA0pWiZqK3KRUYwau+u/iS
2KU8x63GCk9FiBkmQPyxKwdoJR/93NM0SfqBkyIc8PzZsvoCfJOf4Y9PcHJM6nZS
TsqvIJuHkQuA5tvJtTBll6PC7uP85RIXhwasPecyUrCag67EfMobcAjMN8T4VPTy
5/YH6CZ/qvosWhogB1apA2+fmYyjZNGbM4JywErP8UTrY7WEYU+s9M0lbRnE90mp
1dcGXhGQlnu1w8STfJRCV2wazC+18FKI65MUOQtKF3tBkffpueI32qb11g20jYm1
MOImtnK9dwKMzbGmsRA9oJAmrgH7zudifyy6hQh5jAv4MO3Vo2InDW44/niqXiIS
9mpS1atllS5ie/APhp91Uq+Btyu+ycfUIRvJVEKxuRKT4CWAgna2x23hTXLXp+EQ
W6ZnqpuOR2BDNEuW3yI5GKooPKo+QCjVLQWuVeGTo6AltUVZi7K5J4qnZgVSsZI3
ABlmPW6NtQj9O1Htykni0MH09Ge8x8XyelDd1ioTpv4wTrPX6dXTtOQ+h4vGJmNn
MKCwearBS3esWFIfpBLKOzbLQxE7+XO249wat60+8unip7TtaQPueKhoeL7VQh54
p9L0dKBtyYBw05BFvuVRgrxRC9PNOub7yRjwU6KIYeYDQQlpr4e3A3ZvWGJ90sz2
HnayIhFgL/MqjPaTNdgXu9OgqhO/OUOdwLqLpJUF/qa6C/tyRNssLsf3l8kNk+vT
IUS0K9zVJHB6r44qqI3k8ViuZslO+M/IYf86pJoDH3E0tUdif0whs9k9F8JZzmin
pZCcJcHRbowIzoJkbYrlJkLISbqHfBVzLLMZGxuZOyrnDQYnkqAXX/OduQOF8iYx
EMAzIHIcMafW4SoPX1KDnCWciiYI6tQj0Dn8zeUb93cMS4PfOrvL+XKPgn0kg7IM
Up3xO1iagAXSOpJv94uTJOAsJuF3gF5WKwyWS83l27GtlUnfqHTETQlcbj+5WckK
HuZt6U+3QojQ5EbBvS0wYbXKcETywpqmMllidj5UfFnbuK4S9r4NufkYfkQVWSkA
DT81CFtYc0cZgkMPHRp/wlnNscOMPHBmJSmKSvdl1I5A5NDsFhPWDkWx5Jxd14+o
bBcXIw9m0DgAEdapvy60qO6BrxpeAb7cFf3njPhsjUkul7XiD9RlEAT1IBH1Hpgq
QAq1yom+fAjDzCeOunhJKScHPIdhFe/G+2gDL6LJ+EY1dbL7Zo1zlG1us8m35sg7
0tvXc0rbYVWbtrrAF0nvpegX5b5FAljpDRPugjRglc19SC/JJGGWLlqfUe9o7eT2
Drn5NPcwfYaENuAjFpJ1l9yc2qOA5nj/6jOTjKHs10B9TABBCR54nGGW9E2JEoht
2YdS4fVs9W8d0z6rs7Nhv7l9b0tAr939ngZNSA0s7QV6iDSEVX/2yk/TgAjqtDw+
+p9ZdYChqs382NvWhkVnXePKoojP7yqxDYEDbTNzY+Gr/RvgKWWZvQ3+l8fF4Tav
7FnywULbZLcniljom1qbVYzaGGy6+PfkE5riA8JToyKPbSaYw+jgZgI1hLN6CSYS
/BgNb4TpDVBe1HHyiUOozKSVxWv79fmq8XM7fOewAVoydaXKDWaJq9zzoRurdFnm
ytbNETUK2zSLquEWAKtpTmVTaIY7Os1CP7NWKFZ3sNN1WTIQvK9ehsJkiomameUy
nRx09fQVcRWBBTD4TuIYbbJbYA0f3mGj4Kd694rPpN0Gnp8VkSquEZX1jqd2kA+A
OEZL1yVvAdLEsz8MciCaDNxYxSpp8UU6XOwimL3crdPu385AlGrwa8X/JSKZiq5F
d/UODvZvxtncU8REgqzAKMBzT/Xr6SxOtll5VfXMrWYwtNlv8cbdzo5OpXrKPYVZ
eLFcQ1qs+oemmnljr78xb2po0q0wwcc5ccawkQ9pZg4IL/789PUeIMM0DNWsIKWi
/qpQYo5WS0lQKz0XptkaaDwPBRMq72r+eDRiWZ8RiKXrRauWZJLWRuDLy5zJlmbe
aKIw3075iFk3TZB2N+Hg7LzuzEo6u8+DEDUBxRtAeI+ch+ox5xX+PZ62GpUmmUgN
wEuIMfCRoKeIuHZLMwbWltKBNDRyQ9WEcnpEOzbAvlvAx2SHRDUEe/9UC/1G5Yd5
NCI5LfPzkm7DIaoGzKGcJ/AjclzhNPYRbn3Hm7C+xqsXmY3+9txkxCXieKszg/3Y
sI16HKDPvApG09VyMDV8Zo1iXpCzkOKTBLtK326Vhb5TCdtngAVdj4xlRcE3+7eX
C0kUe/QO3dsZqh8g7uaTVg6oJvSdBnOX4YGH/KL54Xn97BywpjpDfvJmd0BrAxoP
GGmSWrDzzMdC4nRhMySBIPDFRdJghdRB4vW1AYLcvcDcmNcjNXaPlAXAmdNIH7uh
P9mnDFjrXbVUXt5eKcfhvbIoAH3Jj2NNAcZXJMpn4CgzCMD4ve+RDDcvyoLuJmRh
NYBIGDOvEo9n4I0fPY71kgVloAntNnQa0U4TaRmJfOD0yvZcwaG1U674kZHWdryJ
XOKXE6/3cY4D9TulrNjxyW7NXBeR03TMilhoe6n6BnDd5vN1YzmW5Gob9lykqbdL
rtsr2Ouf0k9JFQiuTEFx6UhUI4IbR26nOziAjGkymdcXo1qnDH6OYnUDJZVd8lMO
N9FX35evQ61fVG+jIOBuMVUTIsS9ykJ+XesGPxQED70nkQvb/TmEAYDLM+ic8gTh
ou0nTX6TL3bcxeqgkyl9uqTRg0VG3kU4sot+RHtgm5WPNaed8lOYs90P3Ya/gX/8
MStzTJehKegpNMtRaDzMg1GV/K0NEwE6fjZ0tXZcMJ5k6qhJEVwHWc7mZ1PhnkJf
dC/qVmWhCSj0VgHcI8ek/zAs8EHcqfOXWvZRs/LftwozxHD5aC9O63F0nb3qg6Ge
7lA5QM74ReGfAhf3M4RkZ8Uc10u3YT/25g0oIFBdsfwzJPJYq5HClgRXRPl2Qezi
rKIpvhKPE8KYr8GJcxCGGiSGXH4Y3Rg9/spncPsyXb+qsveCiWVTMSHcyOjOzdPo
VG9M4MAAaOLGleQU9yjbcPU00X3mX0VofYOU4FCHiRoI1QA6gkN9mK/kvtv3jKKx
IWbMHGUtRUrAJixPs4Ieu3NvSygUc93QqzXdc9B1WKbX0jOkSV09BTLQOjP+pFFp
8A9VCgmek5/2D282kNNeXV77a6vflLPL926EfwTLyXrhNZS5ujgjeyGtL0emXG/q
yUSPcyg3HAv+BZK8iRsfLaYfx08wVUVdQA8QO52/yqLeh6Kg6xAAmEgPtv2uFAP8
CCyh0Ont3uVWdTn+iIiA8ixJp2ZqEbJHKOl9n1LG9dYkzvVTWqkmFljoJVBKn1dV
onhE1hyTfWUmuLAm3t8heZwMqMZcuaZlBoarVmLv1rrBvDMJrShFKkaiGUdpAbj3
Xo1w2tcfU1n1WSqoxLuKrxsHMSafHrGLZhz69j6PCT8T7Pbo+k67ZawaswS5zLGo
ANkyTBS9ZVXfcAtJoO972XzkUbhtBuRL1cMhdRDV8zOMA7/NuicG4Nda9RGKaI5a
a7Dr4ZWbTdyZISQrOMHCbN55vwBN8VZWii9uEJYQcPAC5wW11oddqDTwMKZgm/Ds
sWjkAu2r8fBmWsTzlztSqFxhk7JiBxmRmQKdh3rvYfS3grqi/nFNsJFyJih3GwAM
ejDtDG7vBT/bn/PAlTh32PphkPBNGnA7W+nI94groiMzYZy1um1tc44BJ95ofk9Z
x/YUzpKH95cCYsu8a3R7UMUyCgZo+YA3Mk30hFeIoCSib4Gtep8/wrwOErdg0T5Z
yJbx/Tl4LG9bX/g/LR3lBbxFVZR0n2al8kOVrwT2Z/XXgT/rshBkZo4Ebd3CWWfM
cGh89njA4V1TzZxZ1H6n7Y59RierU4wgRWzgZkecH/hpm8JHUxk3Tr1Yi8W53Qnd
9219MRCRfEDQ3gL8PmuD8zlIwzXCfMrpmi1uPnhKNQOJ2s07umknhGCaoiydv6PH
HSM8Xm2lSAfmtDewQTlIPZDnZPiN/eOzMKxPXtICbxT8gmsOJb3vEooxyhOqJFi+
xnZTZfMPoh5YtWqOr5KjXtBIbUbWPJ1p4Dj+Hm0rIpTMDnpAMZsR62PZpFIgxKPH
QP3OYtnw2u0PrChKIb0YX6YFS8cxPH2G+l8wKjDLl9ugcdAyZBKo61rZEti6veWz
WGxd7LVmh/3V5fiUGKIQDaNHjZHJgMI17t99qV6U8xGJ916MEEI6dS+vH3/mqWkL
oryz6eQKe+3zKL5d+MindblPYRM8coHX1HSSdUfWPxWwpDnuIWmNoHx3oXA/N8xK
xjiXeb0S3Pf+jhTzxwnoni57rryBu+kpU67JcZWq0MSOy4vacRATrkPZpl2COeTD
PeCQ1d6sO+Lkqw+SSlq22VpM6f9AWphVM0uSVjSjKqT5eGXF4TfEfMfNVIQeOxh+
xqdflwkW7dG1oUtc6XIG2Jnf3pwhSGTzMvwrcaQF5e3t2NtLX61mNaIppFRJzUNh
sfkgzi+DZ3VjmaHaFXDvSEAauIC917b17xwaU+ZN2LsQxpeOk9cjMlVKuCgti7Mz
tOD+kZdzpi64Yr5yfCtzT3tYiLjZpPrqhwcsp7hbw54rd772DHtnemFc6YpI4pHY
CFbQJLCNTDNlwMsmGNtLLFh2fUfNeyWsFFpE8cBBQz4gy/aFGwj4mjeCVp911x2c
oi1jcbsn6bABV8GVAign8dVb1kzUJVRieQQ+u+K+N4bMashHNGLyYGVgFiWBnVWa
KHJkmcMAr2VWCyFvRX/zgbanjO9uvNKLgiOqGT2SbJ7z+/eSse5w90wuEOzO7qUT
/ICfdje/iMCkbKDgxZrVHBpiZBnV1T65s99ppz+W5FEpiZKbxznuGmxU3syntJbC
ChwZUTMu9zO60Hj/tHsD8BRuJ2J50hMP8YmcqKxRq/D5xvZyHyv8EYK1JIVc7AFM
p4tYOcJpxvOgGklkAUXDynI0EOPiuE1w3P58dg2bvbykubxZ/TpZr0JS9PG4ikBA
RDt0duFNDMpEjzlJDlYMb2kfjCle7Za4nFZREvzsNOcK4vGxPnXprrQM5nbb9b7b
YsWrot75VpSCHTocmcVeOmZXxuP8CA6Gsxv8cYscSnhBJEtYY8AQq+NuqLt8gcNI
ivLTlRbH+MMVkr0qvi3TkG1+WdqLaBwa/7s2MtibJke5fheOpUsz5dB6id32y22i
EEtGsc+LyNO7SxS3mgup8r9saTi1+TwuN0+UTZW65t5+b2hlSTgNfZuIkf6fb4B7
eh4DIKK3qr+51Al51qEoqh39tW7XBeJ7iONS40rmCuowGXe2dHU/TqNIgaB15E/O
ecWom8bOzPTqH8QIVvDP3Uiww1GT4DjW8UndNa45ztkao2J0/qHLvh/PglQT5Uo1
o0uxj35AjwhS73IpykAakMTO8o3+EeGQTSAFb4MxFDitGgshc6h9dNQ9Yj0uP/KM
mnI4Amg+PUFSbKn3qkup3RXuFhFkVapb0i7D3OS6MjQG0f1vlkf33syeh0islRaV
oepgkranEaDfims/AGqmMw4cTg3QMvsBzID3nnbjgHolpjgTaA8uQaGf9NEmbaTv
zTnWyGG3Apt0azVbhcdk2UPlYN9QrmtkeXcJm1ibAdtjNHVLOGznAtGtZYzQ1spH
m+qJCTCaIyJY0daBcUgqhiJsW+SPxFdJidt3xgZFhW9O3E9X0igmjaDP2UGnvitx
3/dXh9osTqpwAxbKP15fgk58XaoZQiCJMBi0i2uYARMY4pQC9RwZDQfcRJoIvrxN
+0V1UokD2TSUmipGbboZV/QJ1cos92OM45j/2QIuNMh3ZYjCZkVAXz0wT0eaBQV4
BXiNutEVMJ2b7EBeVQ0tasy3dKg7j2I/gH7stYUUv8W9/ZY82M+HRUW7tDIDF0/G
pIrDtsPqnQN3AqmO/EP8fZPZQBDdBDphLjzsSgsmmanZC+ZHaI6O+jjjwZy1cK4k
KQ6Zi+g/kQp4bQg1YzjbKZMEVOe5jgep2PjslbWHbtsnmbm9rwl/yivdDR7mRAFc
rCdWcxj0Jr0iRLgojK89zVVAiEtYNwvILL2bPGSDjydSAe+ZenuAyoUKDxJDl8Wv
vWyyrR28AAAfb2QQX34ECI+4aF8dybq5xfRZ/CcJF/QoS5OC7g0fR4um0dajgQdF
zNgKj4j3JYs2mEGfmXKkJ+tFzl3Q32N/Rvw3zrdIcPfctMoVHg8D1MYalqRh47KX
P2pFDeJp7xC+j6AzxiKGWsDqoC28ZsgS0WWecAjcBkPbsgRIGiEkskvmYbdrA1qM
h58JclzMyr8hjVezwmCbDlIIKITQ1mvkg3oUdtMzWa5i08nJxehzBdFHO8pi93D0
3aJFq27Ynopw3WU9W3Lh28jTUNuYlfH7nK7/6Nj6ueflpuZLSjaE3/xpM9XIDJl0
BrqW5CFOlY6Efa6OqET1B7XoQP1VnWC0/TZhDF0FwUtguabw9hisNtbVfJhiKnC5
y6UEi5ae3Se6LRmnjwnkMOOVmbnlTkIETA9w030uMdwx/4Nv6qmYGsA18SBv56vq
zZ2NBG1Zj4FS71mB9Qv+m49s3+nyDMEsBwCIHRJIh8luzx7FIkL3Kk+hjIGIBXR7
ALgvRdXXTyLt+9e1BpQ+AQzu26Xqz1ge5Ec6L6Dh21vUHxBjsQkhxm7MSlEyQBA+
2dow8W1NT8yqoD8dl5ZqBKxBxkiL8M/hNG2WzLE36eHbsCjMfHwGCFL3YVyluVkz
b9O0JKQoUK9uX4UJLQAJQ+3OxFSUnA0JYdfD0BeRxoO4kqvE33G7/yJkMak84L/S
fvpvCP0URrEtsNZZuqgDmdU2DtrO4MEr5jo/eACTWMTMGowy0U9ZwROUzQH3fNzk
L29Zqwdcmz9ecR70ahyw8gzRZcLMzE0r7qlvf+pjquR+aZis7SILDSlpoIt+wK9O
63Zm4+pARL+O34YfRh6dElrjEFCCFG2xyo3QCrLtwWXRQ6AxK+H0MOg3v9Mjr4lS
LQBTsPNvJX4C4X4ob+J3t1/dkeRT1KxCT+Ijupy+k1DNnUxKngOfZvj0QG4QIlZU
iNj5OQJF5m7QfkNNACsfmw4sQyCYtm9G+RudC79W7m33LSRW8Imqym3EyzuzoqUt
asUNdWbCO5SLkH+JmpvhSbGgIZ0Rw06VREUaVeryWyggFNG7zmKnSzOZ/Pq8DpOb
YobjtPStyaCESNK8oErxKEMGwnPW3DNHGkXqh5zVFSQvTcl+GyGyrXIS0awXKDYp
u/7UBCrEtQD/DthnPqcE0OLE3uz9MSDUi8ZcCrloBI8AKk1XIG+RXZnIsSitfiB0
oQs9cdwcobs4fZr7xxIR+oSnT8Li8EOJNPSDPpnb+mml8cA8QqcLh0hilVtqpi1V
cAChLgyowz1oIw4xYGGn21nYg+pTwFI9VYRt/fX/ev9CVhfaYwzPyCtxIm/jK3+n
UyHJpITs8o81Zqj+qAq2rQvjLa7lEd0/GdOE/ataNEGMKVNu7OehVLFTVPmuQ132
eRgNwVQPq9BMzDpV8cME3bqZJwxAT3tn610gYfarjlHx6GSQh8rLx8z2EX5p/nvW
l8fr5ra84b5yrPjp5g5eAn06Wrr7tUQgxNEqn6Bl3H0Uv3DBXBgcf1avP1EPn3M4
4uvu4i1FSkKUMazMEkBX+fgTnZ63nd/U0o/t0RBF/gXnnwt35chq5fiERqvDMgIU
ysN8IcUbUIKoIUQ1RrgTAmdWDTF96HAh3LZp6hGtwOLfK5beYrhASNOIQAnw55Un
LE/olIbpu+bBk2sktJ931VvhjKpTJ43eCdVbc0HWgXA6TcTpExc2WwIaGXJAElUM
L/WM3XB8K2gVufrCBzl60O4suIkCu82qaCzUo0xqfoSdtY3lQOrQRDPq4XVlQNY2
6BZuhy41Kl/VQ5qhqZfpd+020Afz+qgRDD+hXtD/EZ3YdHu0eDN6rQoaHZTMwGUf
p8qB7TLGkajxsZ3cHeBV8Lr+l6VtrnGTPy5Qgg61dNVQDo7x9H7e2mCYn/PMNz/P
NstN9YWqYkp83M6hlN7bMqxGivrve2a8z0QNr9d8DSYwhLFlsv1T7skSfNtqpMji
POe+PIwubmhJNwOl2zQIyBWYdZsC8iaLck4ZlNM5mkv9J6L7UvBSC/oozBLfj7ZC
ngTl1ximVqIySv0BegAkYNKNBxw5TxSu2fu8dQs4F1mRZg5ORFa66LAmco9/C4ER
atMAc0XG5PP+ow0Ce4KTsDx/HHQ0iUoeY9wez7+nBHBAoZ79wT8aOF1iTPKoWAMI
F1uQ50HkyP/IcL03ACEVDTDVn66ycaMySQ9aMTUjqTSZ3sjrhlDyfdfg5ZiFUMgf
LauE8n+cvfCKQOCPGPG4VIy9co8oum5XsgHWDI9cfcRSs8cMVeq6W0aWjiD9JIQt
6tqAbyB57APPRk9cfbE0YMOFQ/Jm91xXE7gd+BmfhzAcqhz1fN3l5oSMkbIx10XZ
yeFOFlx4NMj7UUwQn37CD2Rla9wIKpWwwlw1gGHFssx/vFtl7H+j3vazR/Qpfkb8
pAdWdzK5F2b+HVctgr3ESM9IOObXb2/HzAfrNxZSu5eL5QsCpzo8IJQtV74snmoS
oZ1hlkja8da+3FXkBRi0ohPhINunfxZ5UScgn4YMcyDozQtSNUJGO176jN7e2IzU
FfSB/TCqcgF6I+czRLhEIh0itA/d92DGnPdDsZOBPB3B9SG4NADUw6D2jPvhsVNG
kIaOblx7AK0QYEC0CJrHnYD+pQkxPDtH9jmkNLmUF1jwcDAGXscMcVj9NJDWf0w0
NMguqG+XcrYaPMLEbm/vXSLmsfF+mwbnl27hTZti6GTpSsaZInrI1j/Uqjz1ys8l
JwDxVh+8bgRCHSB46Lbl15ZTJ+j8/CmG5MDlBXI0Olq7Sux/x0GYFdFAcqNGU5kM
kxH4POqZpWNdiOCaaQD+1kM5bHi+eUmgQN7dIKv96PQPi9eaUB9nqKNvv+mfgInj
7lG3RQhZ8hDuxItdv+Xw058kZcxqweizjWxxgsZo13BHBqf9j2OQmlkek4HIAY3l
zPEgYD2d0d2Ubv37PCh2t5vTkz1Cy3mrxCdSjQd4JVe6c/4OkoNJnlvH+s1hF9lk
MqxrFj+naUZn7JsQHukRYuhBPrDqWAdcrqYqFlP/WtjGES58FS1p+OqL8r8bu9+f
9eKa1wEzdZKsfTsKiX47oc6+i5tdvLaTb640DuR37Sm68lpb30pIZi5q1ZrhFBY+
MOyQHJiOVeeIIyydn2ukExeAG42JSIsRBim6w+Lhmr9NMz44zvAJKxI3FDkbE2Sx
NYlC6vkGPLLgHz/LBn+BTiT0x7sbk+LQd0oVn70ZPgHd1HhTcrF9gU4TPhK0R+Lg
GnspSsO5nkoUs74OYqn8/4LaPsLSZd9/hhAoVIz/JA3NpAmDZx0BDkJNSQOGYFYb
4uWQ8yq7/7k93VNd5ip4Aacbq+X4BRa1D71QHFq5GXParGj5Ju4woynt8F9CMFJs
NnRvup1vuuOF548HdznvI8dzJypjWkrjZGGlk3nIwRJDj087wog5CpY14FPO9OTC
C2gpYbTO9Z/10RutZSsyc+OmT4C2MrW5dlR1ws67JEQsBw9ReruCwmZhIhAHBkbS
wkfes8Ea9aW3rdUh1z6DKBB/ke7Nz6JlK9+HyS1buf6whu5p4xUUGSwNSP/Te6ee
INNeNOw0Tw/Rng7yevoXtBMdR0svx8hpBa0bSpwxIZgieNBCXDaLhUy35N2CACCY
YY4L7SDQWC87kKI/ejTTqzXNMIyI2zPcgBZuhZu2hQPqi3ghIKUVixOaYavPWAFb
4CpDvTt6Y8CUQ4/lRc7fYHVz0U2NM7a0UIE84qUPB/QxsxG2mUqc1ZxMdySMYQrD
Yjavy8KJx4g1HfM6XRuAz9R9pJT2R2EocykMeaFLi0dxfy+M3Uc6APxKPwxyEpTN
6bbasab9qYQeUjggbPt4p6vwVWSXOJmu6DEFGSbFAj5ftRxi0zLBoZamqA8BuA2G
XfLAsqlMUUxjKNlQvfrh3kMi68XdJov3d2gTCabTL8gwX+xqKYvxs32AtWLzEnFF
mBCIdvaxzXcbNueiHWhT6WJdT3D3/b6Ggnp3Nw0qPXQ85E/knFk+Y1DEA5asNA5Q
5QIqxknWif14+oWbHv8ScoFQXXTOWYynoYkt+GjO78vRndurvCLuLq6zHZJuo616
l5//c3AnbLSYlG1Ajz5CXvaNbBE+wX5GUgpP579L1urhcT25xRVI21+mkKrQBja/
m7dXt6xnj2DAqAosa0qRMcYUntSHggydNc8gpjbVEQxQquEgg7EyBeLH0+dpQPr7
wHEQvo9ZMj5yo5Tl01fLtOHgOe3eseADaImSsFmm3ArrxoqSonxQSijgSgSSuhbd
aRqNBw6PNnorZ2IBsvTLIkf3LamJtzDZeACsUZxA4ds4Lz7b6c7aWJ5jzlPEfHkQ
epXXLCDNATkg4fbvg40a0aFuTAwsBp1xNNX28wzN7G2aJ5ipHWA0d/g8MuM7dht1
CyNG3klX7MoPlUmwMdtFnEwxCqkJL9H3DxhDwctq2OhqbAphV8Aaenn0T1+ITQfU
euaoDgX1ZuSL/+vuJEhWFkFuOPj/+PlTw0XKjEqo7whxdJVH8oKa2w4oxPy1eo24
0qP2pvYZlfeZIBnrHcNu37AB7w5L8vkSxfqXGm5tFXKQtt0+oYZk37jt0DM557mB
2lymFzFcw6kp9cAh4FIvfKE2l3RYC2tcn5chJkskUKwWzmySnq1BIq5DyTsihadE
Bvy4KA+arLnw/RK27lnkhfec8ZEtIac34lN/YJnK0dHBIBG1rleyE2NAvnw1qN43
PhzcdvL2q0W0a7Jd0JNQG/TppzSB5AD6GUpz9Y7PgTGJZy6NXQZn2n63DmGZiMOh
e8wyliblwPiprMaka0vdNssMv0PfMrb+TXBxoeg1DCGNkzk10ukWEi00U0M9i7aQ
2T3v8fnup5XrOAq7EFQ/pjKB0uredRRbLMZhUMNr5HXf5LDfvw2S/viCJQGPP2l5
pZ2l/SqSE9WDKFbx1Qrl8pMocLxl3LdFKM/SM0+2EQ6uCE0AFp/kGLiwxSW0RbAk
/n6CviGISHuiWOnH/y1QMpikiNO1L+mD6Hgm64rpnVgjLYHNFXQKfeMa0rWSqr7m
AhrD6aiUWdyQJUbYsPWXRTMnMm+TXjjxzU7sUHsHw5raoWAY370K8Q8unuFKml21
iqbIiVEEM9SKER+bZrehtj5Stl4ba1YKY6vkMdI/C9KnQ55ln5J/SJ5PD/dhUxy6
GLG/zBZ2q1i6rAs5ZCCZBqkUIpCfn78ZfSYOORss1kRXZp1yI1xYjlC4u5bpbeCp
Rs1m8MGbese/mA3w6LEWrvMORfo2ARGCsvbm6ETUMiePjC9lQixxPf7/z1/Re2fG
W1hq5BRDH4J+svanuOO4oIjLajPz4TQt6t5roTpjASxDcXHPYbi3ccETyxxbXZAh
IDZ6e6NM8Fn/B0yLUWwsxCQNK41BSKPnq18rFzS4CL3EpjfYeAN1JCljW8buOuRd
Q5WQxZBz4RIJFqeP1SCuDlFY5OrgFu4NSU9BTnA/7vD/FiLHVeSJ18f7aVOjDVvz
b0W7q5oQfEqYaBlqwh1OqVXcOHIw5ho1UD2Q+ozCWweWqkEsCOHGv1K9xE5uMkzu
kd1oKRb6B43yLbZhex2SWjH+Ptn9hMGqmVp0kO+LvyjRevbXfcuSED9uRAY44mRu
BACZyEKdC2DklM1TwDsjo8H7NM6faDDro+/UCZESII32EzFoeL8uh1WjaaoCx/9I
+luo5GiAzQwjuqNblwEwXg2I5WKYmbPr2TjtACnGJB7fleqN6z4eqEAqzVU96Ipk
zU+cqn6FudY41bW+xC9akgY1hF62EzbWXmtrjI6jHXIKEMIxXFWFa5+K8xaQ0CZu
OMulDKcd0X2lDfjjMoIw/lSOkTh+Iffc/lK1l3EWBmW7g7YoMQ37Wx20i96DwoiD
isphdOMRmChPtqAY60di/ADtVBO9NDqp3BlkbCJ/USFzDnOVQahEjlOT5SImVsel
2VOUEKRNcfTZGZt/oUShrhVOhoDn8yIKY0J0tZHxSDcowCfCCz8Td2NdEBrNyyH8
5tLSwwQ0t+HW7XK/dDuzpqxIpDQGvHMoCyE77Q4bLBidEJbZ4HiKRiG8tQ/Yaa29
/WanNYk7ClUqpLt1jSWWw9wX6NbmNFD/Fdgb5+OjZ3MhfY7SRqfbI6l9jfAZqSlb
RCzIw+achz/4F2UstMCMKI75Qq8SX9/5sVXMoNYHAGVA61jvMBIjC91mYTwGS03P
fLniFckC4S5dllW1kuDoJZ9NaMTOOAM8w8EhQlmd5H2AWAhRmzK2OE9tdTObWvsY
K3UUOqEqQipAftXCAcuTyDzH1f6Orzfu0VDs4DxWkfS5WGfL5TT0VhyR6s6LXagg
XtgnvRGOSvuCoQFk9m4MdXf1P0w5eZMGfpXpUncMjl1w5YZioqNtShoY5d1+KGUk
JFhu27xXTNcKHjEKF6H4ltqGWx7TQtSM35josCiV3uGHSN17yfT3wroyPZjbZLCP
xDVG+UHH9Wle7Vuu8s1UF46mU2748QEa/NovtQgBM75OUqeldenLfp1qwVOJ2sVN
eOeA03ZS6v1qkunfuCzbNJHOP1+PS+UP1a5Pw/JuJc2ItisCCXcnxEdgWQpVefWI
VqcTm/xoCij1fSIgAJCCtqk0MEIz6iC5bXQUwYPaAOfW7jWlaadm/xA3BCv/le+F
mqDjNib5unCjc7tJmonMNJ30ksMsDXL7Y5sYnJ7dGIwafV3BrQCiERFl/doNGJsA
tvp0Myrr0M6hBSPSleaS0GtMYhPIMnnBfqWvg6pbfrXlOws7YMrew0WhNZVDYp12
LCgQAT/kJmIiuDkO6NbIz63o7xyly1PNiJ+QAi0giROE/kZroyyNqBkmMh70CJu2
jN/3VFph85P8KjqetkZTPuwdygd17tqCIhk4DRVLmLjmXZLX5DaRiyGoRqLlkb/7
rEE/f2Ygy75BrUD/YLJS7FkJBs+kZhuxoj/hMl74DbaUTic/8OD2tVDf5g6/LHjU
TRlKQTUDU6z+luVbVf3TIpgWXKSiKJFAZ0gOBxEfk6dL5Tf3y5hEnuGJeUPmgzQp
0o7uxIiQIBlVtN3gckerfxV5mXzPpH8J6O/KjfJuvN3bFHoWdmEgqZUZeNthQ9Gj
r2bidJx1d1rgZXfILygIlL1iXxl3QICfXDBMo43RGb+FeGyVnMXujAXvFUm53Udu
wEvfcxjUAMXUyD9GfnDXgbBxIy1nRyz3AhgY2zgXu3YHpJ82S8SycRYeKowkV4uZ
2r8ne5nQIjLFAKaRUG9n1AOAmsmAi0pN84VeyyMBF2o54SP71QFDwcZQUAG4kUpX
kj/Xwgclxo58lc9V6t8cNkhuUZrI3dtcwVOhTiI2Sl5UL28pe7QaKj/ONdE45Y5I
cR4cxDBMpAZdpy3e6TLHYIn3mu7joIQ5v7dPVT3+SAhd9V0L8vzAI4GVZkErfM5D
phbFbA4uHCjW7F7IrZFtqupCzuaB5+rZG2jy7AsvaJTS4HudmBdpfMPi0Pq5agjM
zC8vbWy7ld1XHoM2Vp37fKeXjXn1pVtfRjQZyp0Yb8frpCJzx4ysZaeDJtO7yZDe
KwwmnxWPuOvgbc0qoqESMyzNa6bCotwzi0gcHMb5WBM+ddo86VZ8b3qHrJnxAWeO
oqmgdFdK5te1YV7aVblaCBGE65FmaqphcnrlayStNUSSrmMS2tbt25K1xrViDwrK
NdYSvwSCO9pU7PqD+jgfurBTxV7dQBZahf79mukbeuI4PXpqABheI9JOQ4r3t9qO
FvY33b8zCf3GrFnbJAywqAhnZGIMTGpijhPjGuJYCVW7ytQOTqpC2dHdS19FZg5b
8DgFGUwbWtWpqntro+oKS9MspJef5FVCwrUrkrDpPsa3POgy6oPSlKAdJ3Pq3dQV
M7m1rBinIBrv8Lv6eNKDrjWUCQGOoKXrxR6fzOJJVpSx0sESItkIVPX5nrqJioUT
uTgYHSChM/cu6js7rquUHuXBAa5oDPivueKJIPZJYqMLr4AP2jSFTdn0Bcngq5aZ
Fjc1xNRw62ZmfLeqs9Y8l0O4WksibHdYsLqQB4t281pBfTiDwcdXziAolhzIVHUI
xaSuZyv7arv5WceOFq8x6yzdTYUZdZD7YXs+DJZxe6nzh52+u42Dl1cB/7lwF2Im
UirFSHSzVxatw+zI9OTnNUcC9f6a8VkQ0hfKMMa0Nx2dEVOP3bgZJWjgy/wRiEoT
qqlEfqrY6lsRewlbA/fNDxkB3y98bSx6qd+w7SdHrZ71OW91Lb98poJAkhFK7lS9
/17BpvIQ0ZZD9GB01MjzX1mToT0LnUpuLCSX+25RvHmqER7GGYUcE8pIAqqqaIdW
boFyEqnxDXIFjfYmPHVpRwQ1/yApICIGjEHp7IOBrOQook1BHmECIADxqaCDFzNK
Qu/PM7oWlOsgfX8nY8fr+XZ8C0WC79VSS6G5Mb75MtLx88oNtEcE2fyyKQ2rZdyK
GNipvqffs75soD4nxXl1F4vDXlgPM0ZVOX3kk4TS4NKC+GiMgBppl0FR/T10awc4
Mr35YgIHw8hdgArhH1qoxyfnf+DDJUdEOufRR4bVbEgbzaEQNsnbXxfOOT6WT14f
ezCY5DvwMaDO+ZNxAIC1nKIZWMj5+KbZyM/q4c04Cc8GTGMcXRrXiDsS53RIG3Ij
wIKIYh2oIijil6JPqm5S8wryacCL7NkZzaLatPCppLB+f8vi8heu7eFyzv625uhs
zbVPXtcAJCwl0MlCRaNJwHEPR9etY7vrXpd91MqopYaGH+I398KuG0e7U+KwH0L7
PrxXaDfosplJ5mEJxt3ZlXxn1fFmURUy27ghVZAw1I/DtywdZzTrsPvbwhRyBAbm
eH8OvorQubyoIgGX4hfGyv4I5nFKEFaN1ihyFqQ0aMbKcM53bwnFvFfj62SLynqP
ZWYmywBiSOkpNDNOTHvlAOQODfoxvS/WhXVDJkAwdykEzwOO6bUqWTxyVMLpkSqg
qlG56Sdv9IepGIoFtmYGoFm2qdaDzTKo1/dY8jQl1GrDgKiQy36NSwSr2n0Qasa1
okAg3G1C11T/EEKP3MMsyyiLRBD8cw0TvBjivqKn7vDi48cy6xHwg0IqbYrmRWS0
Iho/A4NPpsoUySHg/ZJE46l3C32Ks1+6MARw/tbyHP7zRarHBaXLtB7Zdwr7DsE3
hPI+ZzqA6UIHnQlCut9llj7SKzsljIVRgiEtOEjbyH6BArOBgq/HdaErh/i30u6+
Xl8sTUvaDGflEvdpxpYZPGajuYJ6UArvDUNrqfix+BWOfsyXbRusmbHHW1AnSqvN
gm/Iw5AiInD2Day8yDmftNuT7tityCBb2xVP8iprHUQfraR27tezJZJ/y6JhAi8x
trPgos557p0aeKIivJ+Ebv9F01jrrudxloAhYAXBynLPG3iYq9yxQX4t5M6+MllP
eyPvOMea151eKpAN9EBzZPIVFOc/p0cwRYZEypTWsGzsHg3pv3xnlhUM6YtkWjCp
06CtDxdnAE3hSnUTw75gfzFtv3CFZv7WQnzWbYPWeBMe/udIeeFYQEo18xNsPT4d
QNuJlGR2lytE7wMeONic4/ADsVcR4Ao8DmAFl4xmwAaAGMc1AIVCRZELzOSQCgRZ
KRQOV/dhk64/6O2WsfwP9t/MttLIQ2xXzjrDGxwzhMIeyG4RzXjCA8z1iaWU6aLN
+jrFubCxYrsQGZKLOF1NJrxlR4Bb2/D7dTHFiMVjMG/7Yl9omF07pFJMXUX1rgxM
aU+5Fi8cql7WM6D80thzaFIioRnQWcBeIhHN5R6uBNDKBKGXPv1hqRoF+JS8pm+E
fQ6DgYho587M1ZVwbmRjOhwOxlwIuS/UqQqtN8filMbf8Zv6i9c/kvwRp+r/wJ7P
d9wlQqsSeucN6QdC1Bv2PLtq4MLtquWMV+e0hiMxtKfLIF5Hn0Ug+ANY/mx02wdf
X6z2eNWWR0B9L0vQutJZu6IDHOK8yzCKt1RCJsiCfjcuZKt718xHjQm4FetTB/Px
a1KxdKxA2Ii6/X8AsLFkxMharNzcQeH0E+hOMPgzaKqTvHIRxzqxi6mt+SfZ35+6
dzmcPuOfQ+aLCk+BEAmqsQQ2ZVQkzxhCxZU0k2M0yuMlVA0/6XUIWM4TVVm1StbJ
IaEDphNGLIbqbGZBetsfAwZg01Lg47foU073Gmsl7vLdmGo7g4bo7PYE5KS/8FwD
2783dZAODvU7bvC+yphZpCUQ+U1+o1997t7vY5+sYBYB2gbdDQZ6ziVET/AenntW
Lb1jP+UDbAkXf8H5bdDAMe0tHh6jntWvo/sYwYLByPYnLYDDXDgwBPy4bykPgEeu
T5FQcAjGV5/loN2NurvuSni9E3bosnMSzAG+f0uvoUzKNtno1HLSXUnUHI9Jt5TG
J9Ass2Fd/rLbkAYytO7ZlNSri10eFGAML3xsaU7FO6Ch5I3Hbg831DX1/q6Lc5XR
OniSDwzQDgnIbuptR67Mloue+JqXhln+30QMyTd2hFjHWHFECBnCZF/U2X7hHW31
0kYxHXMqxXAppLyjj5oARQQk4mjZUyudEUorNjmvWJuPDQ3MgVvzf2BA+st3fi+x
VSwoXhF4SbsYOFiO2wrba29sQgXwMX2j2zRcqqIBqYdCFbvpYww+Wk+JVuGp1lMe
gTbfRnUTBVhZxnGGmdZTbXSOzy2MhHVB+sD21mS4Uns9tkXi+u19KQxVVeFKXRGV
L1TA++kEeISCOO3SJc4ckOPfUqo2Urx9bYdyxKkBYX7CXGkm9U9FKjCzFBrAf9hN
X/OtxfIFGIPjHyIueNv/HCaRU0ZeL+vVLX0YxNImGtiz/DLJPMZ98OMzyZqhZMA7
pVXX6IL5kCgIehdot6JpK94KJo7zyMOkFhWnXFYE3UHEdv/xBk+8MIPginpr2v7I
6QPp6QgPAkSWjbCZ8g30qApl2T3dBpsxBuzDOp7sAddQwnFSyDE8dUu3E7/pPKvl
T0H78oI3n9s9NhTz+0FQCpAHj6T/IRnCy28F077ci5dILMuWyHpEK2e8quZ2VDyP
s2S9e56ffilaX2WV24mo+nvAh4xZf9TWC+8E6xBFTIubJk3zm+E4C6ah8kodjPw8
9nAZ7MLdar5lNZDF6uEdsdvhTwz1JuC3wSnblEBMVwGlpl2ImJO2SCzYENwkA2gl
PcAG2+pra1+ZyS9Caos9NFKLSzDty25eTXJp6BYObZ/wNTBDNaoRf7KexeeakxDz
D+hcNEakZieywOGdZSzvb6JiPWynu9phRWqt66Xb+4r1CsAN5oZahx4PJ0xPf+ui
vgc8pCVMlJXF82wzKq+3A7WsfAtWxV+a97jsDNexp7OG+WRzOg9MsGat0NlOHn9A
h8J9ZLZwZ1IjvCvkocdwJq+wOUBHoJkuf93JtGY9zTAaqSHi5SlsH8g4JbrMSuuZ
WQw1c52+lHRwADF66u6DZYrbJD6DSn07dSWBEM7uUQhwreGdpNl83ENhpM5muUb7
bbI+lQpI7uB32jNQuCqXGyGFh5JJ5YlPGxdpm78gczx98F6E1QW0Pj5wfcTAEfNh
DZa8Z/v0FeWXSAAivIxs3DHODVNsLJVVtKOKwWvk0PIm74CHYsvlhEt/O83GuiOz
y5A2DvhFbkTMVQnmV3HVGX0RFv/NbumnAnf8fAY7eLidbupia11TRWU3YM0kuFpo
s8Um/aD7Iksd/i2rV5lSLMyAgitIOlVr2W0iro2YyWP0TXaKHY3QSkSf9aRySGPw
02Ujm25zpvv68kJVC6ALvk41URMM6YYLShtFX52CvNNHT69xZ7OqTPXzM6I0Oj6W
1/JXN87TLm1aXYTIkx/mjP6Pc3rriaQLgRfSf7bNsRSlJcGrl9vA4IK/Lv1bTwz8
wL+w11t/kuEagqGYfJHUsaA/1WGiiM0EUTq1gpqisYFD2z6rfqC7v303Zdey/ODE
Z+tyU0Rd02YLkNZ4xjHbDD9TctqWbE9M8uJHARJde5VrHheSqXtGjAMRf/SwTqEm
YmNCMZjjCjk+PADOnIpZzKYmbI3okl2qwUHtemm83U0NVuubFDhGdDy95FM2JRST
CZ44GfB309t1pToucxG02DXE7FqVXfk6XxwI1X7Mx/40jT0JL7QjXGvG7SDJYZYa
FDZQMoNIHXlSM/sxhW+bXNb+FECEy9VbZwfn2BvsG72i0y0h3SL5ywiTVCTLCBNk
MkD9J7VqQLHXDQQAs/Ab/mW/BnWi2F/LVQa3gkc63gpqaYg9+pubh13k/Kc0Lt60
+r9dQiT8whElhykUwqekiMybbdmR9edNHwEz8ixmawC9PYTUIdWVTZ/acjmzonPa
wGEGH82iesfl9CvpgDl0mjwdekCFIAvnEXe7avoAj0HoOGMGREdsprYoYzsjGJAp
9gp6PNH/FuFHgLaXCNPeOjY63iXa8ZXfH1pP6lHjYXIMqbK0DKdtm8wQ+pOy415E
dVK1O4mwuURJUkNgNCbjVtbCDKHWFnFiLfcjqhuY3gd7eCy3+z9TCD4kt4N2+NFc
P8/KRraxBB4ItwfMCdcyRkDXUkOQJXthOiFCBbwiioSrF62/2Vjl9st8oM/k5wCe
/cQkloSnCdUjtAfevtHYNk84qU8d0e5uvTfqoo3QKm54YhNI7lSmfoqdE3aExJmN
iDy1lfIssqmpNhNF4NfDf1BdC5szaLnARZOfRupGaNeLLV1mPDq1Gf+9EpMKtIBA
jZeNCKX6klyvip97G3LbwpsH3d4SG/x4amK7TlNz5Ap1EaC5ZbVC5FPjEK7MKdit
hyohhGdAl6RED2YGc+pvRYs6/2JdPxMlWts2BX3ol1r5m0XAe0SQgm/HEHH1c3ZE
UD1pmXIfpLX90YyVtJ6/iaaIVqRELl7UUgLGNtTLfrz1qD1+sJNWy7biwwQJO3HF
Cb9h0oQI2oQhxC0g7aQGTfrCn5ahFHvwLgjyIBhXln5odfu05hlBmv0KS9dIqBwp
MdyC/a4c2MJU+DIMbncgXIf0/H9co8MOtFuIchz30jbwtKLclNPNBP699+TYXnrF
j7oOihOEuOWdHBRVK/EfU7A2+Ow2l17pYR6R/3qHzT7J/X4s6y2ZhBOUMIBHA1kp
tnPAUZ+SgmpI5hkoRmXgLVpJSM7YZ37xAaKAJfkJpgKaAdLDxWGDRfZeCmprq37a
QPrzvqfwdUyIU2dy7m81bj/QsrF70jcmL8F1BpizKc73iMagPaRkHMk6YRwJJL/e
vPq1S6pj/wDfjXdvHuEdhx/zUQBlufGUwQFzHFLKjdDKsPVfyU4GAak4UjIE1X7u
+3cK5IYHrDye4qua1F+lqHmtAAFEusQ8GBXPH6ex4in9oHLDuHvpsVWvLP0owCEL
eA8Gwk58Cqoke25ESfjR/jLaGfZGNa0fD6Kv8rnQAc5rZqnHH0tvnuU0U/Jm01e7
KIbGqmPnwODzgmoTuujohgBYLFk/D3ZFe8g9xOGldOYilbnzDD7L97zZuNsT2bLu
gkopESRJEYcK4XNrBH4GRST5FKQ7lW4EbpP6zbKNfC7cSUSwyBDvRCtMUKIZUVv0
sqDWzfItChhJOzh8/r0YBj41clM6xY5b7J9e4SXc3mLQuYnB1LjvWsILqMg3PhCR
kske2XHptBReXlER63DqPTn+w09br2TLFQE8exlVJicOPpW2Mrx7JlTFixPYrShU
7hZ0/HOyx1fGTa06ookW6a1ktT1YtpqLS5zDRLVuv5nMwUz9C9FUGz45zlC5Y61+
VwoYVuGz0VPIrM9j46K2AmhEK1R77LokZ81lOwFWpciTE5Jl35zuzs2x/8d42vTL
43zZp5SoMxePrwAqeWJhehKNfeoPrJpys6sMff8yoiarWF3txUSmqQ0XgOyYoNL0
8R0YWw6SKKFIOtQ/+mhZ55OYUAqeBjpzdNtz1oc6VBltolTuIrARyyn8WP54XQli
uJ3SewaeiQxpPI8ZMfozeBRCFR67wYcxtePi2LDjCtBa90homWJR+zl7YPWznlhw
eV0spWNwm7iAHtDzhcj5dicnrJ+AABksnW/Jn9F7x9RYT9c0lhiw9wM7KFDvWcv+
J0jjG/8oPSl+2E+HCUQDL0/BlnmtwFv0KyGSGwSe8LLb4ors5sHNvwlmaPrP2Uc1
P+0051s3fEkzuiyOkxW/Z2/nzpqjiVtKNY8dFDW/l41d/cVv/pxdPwWz4flFq0z4
S3FgnZwnAbQjxFhE7BAL3u1juFBJNjSeLuoTymt6LV5Urtzhw5zidYIOILVrwxTg
jwYdqDVM0zOiq442Lb7hkiG33Zwf4AlWpbzN7ukdRubfncCYW/J0gPzis8olJGZZ
6/WJdRqIqeHkWMEFHoYfb3+r0TTeCDJcW9ywskXXldW85S8UGP8NZ55/1b5xDXcD
+kF1p89nGa5sh5vCRfnrlqFwhkwhcTLYDDxPAJovuS5a4MWQKK1bpJT/MdpMjaoh
F3cDXsiXsrYpw9/yzq/Pyoc9j7lr9hhJ0mw9CXQmRehu3j152tx+hfJc7EmIKJcv
3F7qWjKJCO34Y7b2YZo1v9BKMJth9Z2c8iMzbZ3QDNHkUGGswnlGPVHOlKhPEakP
nV5EWrBEmXYk7DEUitukfrb7Vet54crUVdlqDRyuV5CgzzyoB5+QWhZ9g7oaNqOw
ZbFB4bqjtqMHOPScTMpl+vf2BBcMyqbULhcl37mM/4p30LyrInHCuYLHkjpQYcUt
s7VYe45wIZYoj5SDW/FpVkyuBGQpoXRguUF0kdmK3IhwfgZLh717aG5miFcGe+mv
5RU/RlIw5Tv3ORuK0TsaZ1k2GXOMo6Vypk9afn8LWQvRtztmt+bm8X+DqPQUhob5
kgoO1irhjXXp5U4rasSSgSjUdxT9MwY0QU5SsArgW5oo+nwyeKAPQ+ts7nuDzniE
rNgnJTLPbivRzNbOZtD84t1Hg10whYRAK3n1ya0LrlGAfqqBaBcMUwD3S6fVdLHn
OgKxgp1OXcgMBAd1SqqKo+p6ZidqiLpP1paXtTPLYyIUSe7UdF9hFRo5hmjD13QL
/N9SSJbMrEpC7F3STbi+C6sC7gkeTC2O5GAr1TtIpGMV5tcD9t/fTVs5lmlQJWEE
Ov6aWTtSy2bNUlk/rH1Bw/QueXfzeMuchi1wcdo2CjJTpv/+J2sDk7JtzLrhIcNo
h/3w8/sQueYmbRVsVrZUfqAkkzg/9u6+cA9/SMYBj6aySbecCXIICc5k7DVulEqw
mbRKYQ8eEQ63yWXCgso5yygOXY82DDPk2qaPR2B+FZvn8ZEPGzZ9WNXiOBTvN2k+
WnvDr12pTFJtmIbxhXh5xTs135zlOnLzHJl9XC3a5Yt7RVZoYzFfMhOd1TB0Gbbn
WCvn9x3MxWKbsF9TOTzagp6qr4JgKPB5vqYxTHX9jNpbIIL0+1zukTabtAsy+9kw
uT92r9mogMFgcqFoBKEM8lialsniM8d6sxeLaHedrI57iXVwzugpNps723Ylcpnj
ISnY+RI3dqY/pqiNbeQN/rYBxL7gcaYIx615tKHF0MkngtYm+OJke2kte1cxgEf2
spDCMH9xJfYh+KMOTYk33tYWAJloTKssZdMFMONUFjGqyItSK2T6YketUN4Bjf2n
jtk5Zow4DK/QbTZSsntvZu8pBvoLIlaZW6BlPYbJX+zKHgHM7ZNpyyjk5kEc/CjM
rVh1HFI6aP+phcQUkdO8w3dfuB7k+Gq651t7Tpv8xIHNZdYQSoQtswKm1PMgqnub
4XsqRX++T4H4zvPvbL3ZUwwMynong9E725Lcw5JNfC1HlznxzyvCaMCSl5v1nqbj
5ZHTzbSaJzWwn0nQov+Rah+BRY5HVkZslukjeTz63/rIWcsIw5ir10VFGFm/2PVs
EpRtzcLKUm3AGbUKouS5E3V5X0Xn0nfBBVwFmhJw4H1iemCaWuiZEUVs0jAsLpt8
NjPIT/HAgb9Nji2MTyNQXIZ/qJhTkoti4dSRkSOHjxFpHu+ksyKMZygcVbXprB3x
iF8Hp/Zl7pjL08VAQA+vZXG7v6BnYSt0nYSwfOl9pFLYL9Bg40eABFVDApTiuXQd
sJfvVpI0rmDdbE/NMvbYLs8dbuhBQy7MB1RX017jfkX5W3xvK3VTwg443vdCZTO6
a15c+4wRvFEIQzDxLqqVId3o2pRUe/Y/nhlj8vppkMcQO2QEpwFmPVLlbshuKlyI
sKTxDOUiOLiMpx0jBp+Ufhk3xOpzRYPFZhC3dsDP2E2bjK6BQJluKGWZTkM+n++r
qhYeOg9cyIi1yJcoJKeAgt4RwKPVnQdcCH7O/34GoK/itqZrPE9Lvk2IhYpftuYJ
XSK9Ely70o+YuUVarRch25LaDbZGyjwy4YSKqnNnpJKjb82zpoF2+F5lUhMd8++f
ud6ccgFZZ4RKv4/gzX7P03reJKFyTd6vDvcSH1Q5BmhwPStx6Vwsm2jiSEeyfO8f
ka9rZOu4qWHkKxKO4+nF++plMj8/YxW5xV3eLwBUGHPm3MSthaNgeqI5Av+P+ruT
l602v9KTmA9RC6FZVTMEFHoT/4yoDSxrMcx3kWnchlxJz4cU6tA5FMu6ee6WTI5/
JcM4usJLrhPAdDcvoNm+DJhfgztmrmvVeM3QUAhnLHbPK1FXo++Y5D7SksBBCTRq
ARqXq5reGwizW2VFIVGXnR73cHC2HKvQ83baXwQw1MKJ75n82E6O0nVyiL5emMgH
5oU3y4XHHRkYxrt+rjjGdFK1fTPSuD68rkRMXJKbpRswFvQwGBN0ijAR+UzRvvCk
0yzc5JztaF7l3ipsK1vqXmGhAUmz+7bYOQadp/CjlyJMNhkHPRb+pY9ay0CwAM9Y
n77DcIe3iURh8CajfbnKvA0hyc5OEfWsfSN4DJEkUDYcXl6dUdyMeUmN1BebBpzj
D6LajKzgAOJb5qI1hk/eTRM04qGMyztPkKGJEpJnyBqxLSjxe7+dAshNm5bLp/KM
/7XnDo1IQKzehG+dhdHYOugzYofOuZ/tVakn7cfBoDwVMCgHBT8f8UkmZf6Vy+6k
Ir5MrGYpmL3NJXeckQCNvlyI1FZCdkL5R9OlYpv+1L0yLursOA41gQy5lLA3q7Mx
L3Pk7hLWTcnrF/A2rn89rN5Ae6d/6k8Jp8ivVCk3MLhKMDovPayzO04Rl3bV8rck
1G28QQqgFW7K3GowqlP7LJ3+jGyTbToUpl1CAT7h6+OhgKgj83CJYR+6BV8Zqf9K
8kgztHoj31Ybhh33vkppx10D0WJbpcH2UGlMx52K9KCT4zTYPxCK/fGYeXAC7QWt
wlbT9cUFAPJG+pVnvZNmQH8K0BODjYdiIrNQW9jAbN4xcm02iPgVNOsxbjvNwhth
PPmKtvPrS98/2avieh/9A51fKdUyi4imJxf1vodWRQuauUT/Ao79El8aWRPwo4Zf
sxIuTeVRe+IJKW3Y+DaEgxeIxF6TXlobQ9rBrnksx0Yd/SfzZvvDLJuZwUoL4TV5
AINVaZw9cvwsfUmsUY15SgrYHOKTq8N1A1REmgwF9mLIywF+oHO9aT4d+g7Ej2h2
lZYn2Fwu2yJmkcQ+30GCz28B5DW/HcuBw5tyz0LQgH5HxsEKPUwwpeL6J6y3SaeT
gN2vmjcc5wYfu9nUgsbHvo4CpVSZbc+kb9HuDffbBlPrKaLiwsevwSI0+h21bZq/
beYOci3AtJ8SwSdd9o0tlzxUcPdVb9z4h5KqFnChhYcQE5/nBu2Jzre1EVUPqtWW
dHvoLKLycCMC0hKYd1k1toAsu+bt0rH5Li6rRkvWt7RKVUN3k6pzj/P+ugy53vSM
8p6fxeFepg3SCWgeI8ETKETTJn71TRtZctdDeIwX42unPspM7ukgVDqs5dnfgalA
XyDNHo7gZeCxrf1/jcbujOND3fcwbtpVP9rnIvVKVmyN9GcISDhb79fPd5eThmV9
fayTXKjWsVj1pKQ+tOmuy2KnPMZhLRg9dHJhuacVgRTuzFcRg+QE+N7fP5WZs6Gj
748fqcp3FZg9f8St0+BlWERy7sIbsPX7of03u36fNjaa6KkpRGQ1CMRjE8IphfIr
6cxT658tKiXMnTflLes/7WIYcnrjktn/BieeVqiopFZgs5i3aOsVeUHw+z8yTats
4xon5pDaeU/X35ZGBxa6z3/U8+WCRuITFRdCH65upEjPg7BFkqSXvqjvrwnpTb+A
VmbF81S1weIH4jloMwX9XEO0DEwlh9veNufnND5D7La88uGBBmptFDGtxzWtMCov
KC06b/VDLri1So/5OmVrntA3MReNPv+qkEDevmeEl0JFdZWmFbBaxMsgPLgu02r2
W8jR/lJXwpwTbobGJSXeYFY6ZL6FZzuv7aRQkm9E2Nwel2fNI9DUdVcBTh5I8XMo
+LLoH6siNRHynvFFgNi87hufsYsUzsx/sL5bpRe3vhCAzffrA7WnJRqp/418T0pI
RK4B1dq7oQou15pmU5MVwcg1c5ONACLuRMPhB4RiPcBb2ZVhMWDBIdkfpaa97NNK
r0CVE5oZPWriAzAK1w1fVXeuajQcCg9U34gtN9P4U6Ayeh3A9f1+IXsPLVk6ipi1
YL7MtoRRfPjt348LnVIIXzjWMHqOkcGh7clFV5KAOqFaS8UqfKWeZP4R7Cl80+2q
JydcbKJOX89i5t8VNVt9Q9XmpyJVIVg0BER38Cnz51OVg6bDJYlNco72rV+uBptq
f0YEJmbHHrzDf/j+8VeyL/c4j6WHEzmjFVojdGnH3OrDjS4PjJcqw7cAQyMlDxNI
oU+bcVmcFdVeVPIy1rVor0Ufu2YmXfvNcjLfT1snxPZ2KoSxlp8nrce5nYBXSnaX
jN5EQF7yVYWIRrWyZ3IYxzMRTWYEgbAc0cnlCsmV5uUR03fS3RBmSHX7lz2UUKwd
jxSADfgG7Cuzgcqu+DjWlM4Z1h+CGqB8JddQGcjsWz12WNVP/xUd4yWNAUn62CVa
VhGjw0SMBGQqV84zEls6jWwSkZlcw4Q3NcPMha/vkVyWaRqGIQCfKXXudQWzvF8I
deRqxrYhkS4vkudLU9iGlqacEdNA5RSp4o/HPJWldGSyLJvsoCa2rBuggyegRq6J
0ASs7Uce03hyPwl2MPFFb8nVD5z5DXrVxpZDy8+KAU/pTHQbNaNJGIBu/BZXGqpA
2Xo4V9TfuaRNu+xqDJ11QRwk9TSnPXwcAiurxi4vPzaqB0F53h5+Vpwb0Q1OnUM1
AoePnhfZLquNJeemGnOAQv2KOStqWTHhHMxdTIT1afPiAFcgSdf7MFmXoIwxtQrn
B8Ui2WWgI+rQ7yXq7v9Ke1nY0Wzcw+y6kcKLXoQNIL10v2Vc21k9hm2WQW0I3P0p
ncqG38MVhhtsVukPaoc08cT917vQnX9llcSLgUU/2Ew/1zCZluijCH98lSrz42Sq
DXcRcYcclkQig9B2ZOMmgeD/OdIJQwzVnMleqrWOM8XhdCnyfQ91oVR1IQs+MWbh
moQkRSxfFOlKSENt26hwe0+x3e5khDtXLPsKvyU2HHaJ7t7XVa/PPS34rRUQ5559
K0c/OrQ4g1HwDA0IE9ocsjBM1RKauLSpfmoYvyhYMtHo9rRxFF0fEGevy26MMCk8
ImlPOUHb/5uHVvOlA+a3e8AH4zvOf1gfQWkAVQ9Yrn547YE92E3TPPgf706X2qQd
QxS8Z6/Xz73o0u16gI0r1ACapK5sVnpI+Jtxvru/NJXk+APiQC4KIV79cEYbNfAH
acH7ZPuMB/3jJDf0QWIWSChN8I+MSz6Tlfq+BG+/ON22oiX+teU9oQQcPQoASkqO
pE8xTSVibQ/vIsODUvtv6Mq0vnvIVLeynJ86hby1LuaQJar5DqejQqyGY1td3NHV
eoSlO9hjZbP43dIINQRobGf7WrdVo/JXmw19ioQgSCQ5Fo/N3bRdOPf/dXf0RApN
kqT7Bs+2iwc3gqGSx1UcvkzE0/XvratU+3c/ga3Lu7k5gH9q3BQUboJEcGUiljaw
o8lvNDdGM7sKEBmBMy3vwBk5Mf9mTNPUvCUer7c/tF1I9H+q+/nhheH/dAEiPWOy
UZQcLSFM2rTvLpr1KCAlm9ubGROTe0V1xWN4L5njxAU4tidSQuesBHc0ufhDp9yQ
s+55+wSoJcJG5vC02c7yoHZuZyWkrVBnW8GEd5RFiAT06paQ6iSVscf4bKkA4hpc
Va9xyLDkbLnP5a1VsG3bOuxb0WS60OEdrHW/1PlV5bVe7cZj91cGXm+I155I2Pmv
Zfng6tdiFosooNQHMP/HIQJu8vEpqhFnw5FygjnW49bqJTZ9KXzwqlQBJ0mhB9jK
WZXpGsSyvZkArZBfw+8vdO+ZAyfgffVkm4dzaL7oT/BaUeIPnt4cBp5FJ1525ki5
r/KauwNkVcp5fqRPK6YEOPBZvKfrTT+BUHKFJX0dKtKMTpChmrIYmzOILCruIV7N
g+7GAiFOpKVsy5RUPweRfRLPd5BykTo/7+Xg9lEm+KqweY0iT6hesJ2Ad6+tCsg0
2JUlROVM0WHfSFTcDz8ol3sN1ZSufJOQ1PSFzEelplt3oKOcmWzoLuh/9GOjMNWF
e6JQ/Df8E8Zj5ST3TjelnLqZJeRmW+KiwkYrSmIWsqsPn7p8J7MNNzNqQRHyQFTZ
XE3Po1klj1387uE4rdpZx20puOt8PTrTbYWCTIQf0HzN/2PDJzIu6TxpXaKpg0h5
JQG7F56ciefZr6b1HP8S9rtcdTVes3pcqs3P7mCA46N1wDYSC+T1KdkLV3uMD9gP
l/9uEVchM2zn+qWmSt7aqm43pfQ7UyILQr0XnojobCY5GbOM4nBOPVuzaOjEWWP4
UnNgCc6Ago21uKt/gKxvUGkQgeEIgZeXacaAFM3y+88QakQ8Vd3B/ZcunUFmQ3HV
mf+h8C4Q/4sETKG7/CBhpaLMxyHrv1y+eAjMLn/T4dopRVwCZG8HGb4lZwU5DBJ3
0VexzupDz+wlR61Kj8PoTvT4Xj3bwBMS28GoSUO7H0JctFhxYu0Om5NJhTm6fVyD
QmCNGXm7TShNuEqOqPlSpiZYw508ahIfrcdPwMo3Utd2KoI4FqlyQcYnd2BqfNft
yocs3x2tqywy4gzp7W4B+Mx2r9H3XDqJXAnlZhWXeI0R7ozlFF1LayL+mWqoYJnD
sZllTIbHvxQImIpoaUqiXCJmnSQMkmBvE1WYIbD6n7pJxWWf0OZj0/jb36Ttgp6R
VC9hJCbJQnCR7vmgoaG1SmneSsGXDFegZZFGJ6nw5EoopgfXv/jdgf9euUn/PeOb
4RwzgFiFR4MOUJsA2haNmO8t8qqa+i5LwXs7nIA9KDwCB/3++f0cusx3Rdemfe9z
CFshfbQalhBI1JhGKMKa3iEZKGCB3Mp5ZbTx5GoTm/13OyZnNmZqmTcy5VXRacdC
Se4vh9Mano9eGWE1+WndEgSd6YCIobi2VGfmkc/9XsXNAdDXudu3f0gm+9XwLUAK
4dwNFRp4LjHjH+lGQiwEhWD5yxdiiPJhkLQBXIcaop/330N5jjSREBzaLbYCNxDl
UaIglm39M7XNGdO6YjZt9bNSCWkte8XlDJ2KVh2iP7ov3mSaP5uR/JieweS7PYE/
ERk6RU4ZQ80BZ9Lh1/MZPLHNi3L2I9TMtuFfE+ro/TvKYDLwbjFw8MZwiylLR/Hz
IpZXWBtiajeQ8rC1aydgBUzx/apYXTRs1RfN1QoiLZGJaWSGTkSXNkgcKHpVdo4N
6mjGslxssn/ZDWEFbfn6Vbb66uu2HTZK8N4pqbk0O/uRpRNDHsLunJZ2vmv/eDte
+4UX3A/SyXi31zeEmQqAygY/+1yBUY9iHZmm5GG4DEwSvgcNWcyAiUH7/nGsPpPb
Cs/EXJrxTF1+TWoEATZH/vFotzr+2lciUdLS8JsDg4KoBbvbgngCIhXAOdUElPEl
mJydIOHWXU7ns2PFPgSrsrYGqiU8yEme8t63VQ6FXWqsxFvCjV+GpU8+c3fDN2iM
8YX1pqcAl4CF1OTv+EbFz7h5//NClJ2OzRHX4pCSVCGvIveO3dOVgqsSKHEmRhri
act89Sas1iSlJU+TSX+Gljgy4Gak1iF9gs6OfAtKGcNVorgC71WDrHK+XsuUSqvh
dE7Lr3LY1nwY/hLQXsEbJiv5wUOdtO5XvwlvzsgoP1qtYixsGUKzPynNmzaeGmZf
HxrSuwk5nKigKfmuSj0Jp81KIBW1ROdR6VeY82WleU2NbIVc0oalehjZD5l5ncxG
O2D6QryYv19STKE67iDKPsus8IcCeFTNhhGHp9H3TN1beB40PXs7+nEFUfkUdgX6
KsmSWBz6is3JKx07onBUJUSQS7XPiBF9vKB346B/U+t+34vbZ8zzrdxrRrJSHxvY
WqTxLQg62SL1Brhfz2rJgo8joZBd5WX/blv40WpgivuQXoMUyB+wKFsh5MUhdArQ
haTSCPdT/BOZGZBviUTAZS0ITzIShpAl8DlzGZtOWAtc+Zp5ZrkQwkHB7h2EvoOF
jOLcLBwlsJaTI4AGB0Y7dTuEP4rPUvCpBV5G9Fl8EW4idkqmcKst8kqYDK5yVshD
KgiieGlHADbhnZsnGVAyI5wV7fhAE/P/f0BbuLpAVB2rCA6hey2gnWeygoBfRDX1
deZ1effDZvYpFWmGmcTxvD+Gc5jDX3O+rRMDonvmastCEQQzYtEdr8s6iU13U1V/
dKXdMtPP4r7M2tZdVkXvBAt2l1y4O5idxIDIkSvoTnJfJgadc7H6gmtwUZz91DMu
4eqL+E0CN/gu267Yf5QXuQ1CxRzj6Bdqa3jzywdUlNY13wU01Y7n0hL6egCozZMT
NsyD2CkV3Mv443XCf7cVVAUmz/aLzMTYzGhWqej6Qx3C3mr3Zv/BLQ2d7npri1fj
OxxRBwvmSQcb+H7wSlJrXAe1c7sBc1YOWUAMkpIIC0Nl7w3TJVoSHVXFEDwoNlWs
7OktqrrNmQActz/L01mnJOVyOuUgKS2kFBGwjnFqCWpj1IGXPD+hgEIitemE5YcA
XhjuZMkyEQRgvMAGE1GwmV949YS7X6sqAIVgThXmJJfdh4FwuT3xRzK3C0Gprbzp
LCzF482t54qUqa9m9v5+sly99H3/xEhx/QOqpnRvShrftG3YyH9+gQV/KqzquuTo
JEKe9lqQ/DGrz8y7Yc+Zbti6gsfN1FgoTqx9ocX0+0gykC4av9Uk9SubiOv0O096
CdM5Zq9zk7SuhPu+ikSwFLFbmAJPsMnmXzUks/LqZ2PkRC2f0vIVtR7eks5RHsOT
d7QW5lXWxXZYqCszuup8Za8bMqCLq770fV9jTjWCT5G00Ofj6BDGhNz1sYUAidTX
CYSRPBSPJgXX9Oy2utRpNoyRCXExZHOar6XgAN19rnwKByEwL/KzD45IwaJM3OjE
5jFZAfCl6heMxhtEbsNwEvmAL7AWbhBdtwJUq8bpUzza86j5xMXa8deGmu8PWPoK
S33B8aUxUYcRa5zf3S69Yxjb+y5WklthZnZVgEuwplJ+Z5/NvF4uFQLze8sjbXDc
NrrEYSys8Q3K1utYEPqFLnbwHadMxEciBKmqdy+JK1wUkmTHI/ipftGntO342/gR
yPXyQgmd07Hs3IeHOr8PWzW46j91uM+LzKi1d45sU/4lpbWQRDt8I6UfOZcoT6Nr
tOCX+sFZ68ZEDaMDOJARuub0sfNkwmpoDF39qTiu1g8azsylaJF70RkoIs30DTBZ
uI7m+nItpImQNq4udfZj1jWbfXHSZ86IPNfpmTmy2sw0X8fkOVoX0/dmZxtOau8p
VW9FlVrltbahNTTnNNJMk0Ojdd5DSju4JYCTTZSDp660iUlpG2jGGz1XTCMggsxh
gkYeAgQeVqe1SRYaJsfBxyXCcoz2WbkVrONFb1k4ceHtlaW3uxcoOVVOtEYSh6rr
foJyYMe5o21PoInCNfh39ICkC1cZ4OLFRfEeM6wLH0bG1YRrpGaEEwLN/+vnT7Yd
SbhV/3PIeUM+zpZ/bMFmsxiEMKvIeCImfd+c1MyLaf+c2ex3XAv1lbNr767d8cke
RFErhYlTB/Ah4EWhnaJv5coVRcwRLY3dYkoE2jFUbY4Bc58JSKitq/KjIlek4z4s
qlfFrZ5USabSUnFFV5iX/K84Mu+YNH/I/cGrtPstNN06GwqLWoUeqKZDC/Ig+iqA
9vU5WeI2TAPJj0h+TUk1XouNo56eh7CNlsvCJsj4fl9bcIA35vmQxenckqHSVXRO
6YKoywiIZSnw8cPRnOcY+E6SGqzLUMq3x0pa7H/Ts5EGxutOJikcBFoiQ1gMpDwj
rMORSh2+1oeIBa4Z72kWND3BAYVMvOEvjguJZreD5GAWDmAocdqRr1evW1ye19Mb
bDIqqjO6XxaxAHiBGAPWKbxPlVKFT2L6Ong5G9JUkJVJu00W9IA2ateJPg6x196l
Uc9/N1TSGtkcckllm859GLWXaFSXrBREMtBxyfmigi9PQ9GeRwFMANyVy4ktxtXG
hzl+ocYXD0H5eLZAPrh2yYY4UijywktWqBPew9qEbubmjFGwiaibdvvp0zSteqIh
QsCHynQWptyGfShtqSg06WViW/Dhw174HMKoS0zYG6wDZFOkNBQ/jZ0vUPmly8Zw
sTUGJxEncnkigJG9fWo4tc0bXP2EGdHBFYVflTP+HEuwJ+6hVg9trmumXAXCpo8U
1+KJCCtcFd4wjOoaAtqMNpZvpIFsA7LdWYVGFua1PscxHdgNCRofYZ5m31g7FxL3
Hb2yezxz4ZhEMGtnRRJ8f+JFOCRFOiykL3haioP5evARTOkm0wUYB9jt4cdjduZ4
MGOUVyWhqY/nRdLTO3Md8BG9aRXVwNnHe97LmFAGvrRO0UWnh2kWPIPXMBLysnp9
K+HXxNotL93MkRjuT7UyJofe3eBLrU5IetfxiZMB3Z1glBQuv1Iz0FDUr/5O4VoN
u7I/pf4SaepGy6KrqbMt/UxdHy03o4xU8jlCs06XZ4vPdOnqU/Nq/zlcJD7EAd+9
rpXrHs4hvfBx51Tlgu86KCbyHx32kACIqbV6qtlZhw2qGfU5JYpN/9LHnJ2Squ5z
Vc1vhivtQIcbbfkbsGbSvPId/AaPsS/bX5l3+VWhyf2HsXJ+qihgSaG6qTXfXoLz
CGcbljnoSziZ5K3nJDmKSBfbNtpWYqBswbj5XB58sa3qcrihZAoMhUlTZgSxSNZE
LnwDpQqvpVkQcbBOM1umI4Gzh4lcTMgyaGnT7+oSqN3LMFn5kmhWenBTc4ra+IL6
shuF5NrO8zyGGzCNkdXFP+gdY2stnhs3ow5QEkHDYuwjwM5GJwZdZUoRdglC+Bu3
HO5W/kuu/HYvWZYVjuWelGbVvGOHfGH6t2p8X+IBcwphsgxeF73EbbvbHy+yzpth
kbpYr6Cylvr33SRdkmCQgzWrsZR/omjTxyoh3z7cDcIU7gCWxDQKdZXspO69uNLp
81nICyYc1HK9e27wsQQEyuYFhpLbCR+Vld3SIW9TsPt6KN6eR+OgAgTPSMzBpC2q
sLg6hwJ92dKAgbgXNvpka4e5jxmVOaixqMWlzq3kT4lTYPcWrBt8W4xQ0IA6roK2
wwnOU+zdMnkGB2EFH2bXHzpmwmOTn0LguHiNGDkvXDkDarLUP3IPlXQ7AlocjEC+
3GLUAKaeuyIEK3bJE4Zyu6AnN8Dv2RBK7p4sAkjLhXiz/OdVYqfJouYSJ1LRTo/6
phswyVLrUOObKVwZpHx2gflf2PjrWHADOmzjJjVwfzYWoMcQ41vSml2hYIb5oVHM
n4xG8ZeaAsGM7fesepZIKpTtjQ9C5pA5uwSl2yseDOqSuzzItXAu5DU1kOpjLSai
DkfsvXGKFvwd5ngQ0eyZFDcXEMgi6NTG+WnLlbpvNij7wvp/LBm1nh2cTeAISu8M
FHvy8cL7mZTBdA5XFqd0nADyuM+o/gbKbBrpsuSCyBFQpAz5wLuc9oyBdQaji9qv
BA3fl/3Q4EabOLcgM+YO5OkQaWA+lc7BfaLfWy1odb9jEUf8IAXkjg8QYcmsQPn1
d2wpVlQEWherzDp6hNwN/8i+RhcgsBgLYq91STTrLd9xdOFcJqrxvAfGurxZH9U7
RWcCfesQdoKt2BRwDKSyObFwaVwXO3hAtAlctTYK+qF4kasV7ocf7F3ganmK/kLP
V+LncF9kzr84jSGDjJsn1Lvt1bUshcEcl5vPeA5kl+gtJtjAb07hrOsZ2qrJjtzl
OlGRVl2vo26WxZYuwgD19CAVCrHkTObq6wrEcyzVA2mO+L2020icLmRwURYoPPG2
LhFcRPSpo+Rzsoq58Mq8FBAzVYwG3136C70/BpFggw4lcvFuhU+Cl2kMoBvas1KQ
GFTtlHlCdt7GszH+/G3c6Pn4QYQF+m5RZ8yrhLKg4M9ANy5q142OrK2SgvaQt+74
AKiTuNurPahiSu5TyCU8J+7/JaO+ISTUdGu9CvpR55wN6kQk0qqevMOebMOtsMIy
hPYSEpbf6jHnWeMqCMYhJHKWyqYsDPRAewKpYZW9VU2ycBuZaQgbvj7s7HBwIk1+
5t3yvYbHNejJcDOazvqhIppFKm9hK0gUN6Sv0PR2y/4rDiMrlTZ4ESVSwh52NeTH
j/TStroJ3Keh0aam2nwnDypDwtyIBfdC6QUrxEKNbxKxCkpJW8M/xdArY2WWy4Xo
rETfBsIndaHRVaNfcmNEPziN31wQZujGfUfh4lnN6ywgKNAHnRbo8AKiUnX0EiH3
j4/bC6A1PTbug47AW0r7orcT1sU4zhifUFKHGRo4S+6P2CBJsROcJDmJ0UDBpAOc
+g58sBZNCAWddZdJEr9mXNGgJPKIckdo/ACEzX8WpLeUMG4LbGs8cCc8793u2KvC
fiJ9pNWnLxP0hfsHD3ZsCDqOnXZWukS0kDUEnq2zKFAyhWMq6Pf647XrV/imGcsE
TjZbPbtW4vRzEYJxgx9cbPETeUJ7TbcldR074O9ZVykuM2xTe4olMnGQfbYg2qmN
yOebuoBhRTw1B9exmSmykUDcwc3YZzS9UX8nisTDn70O61HNIeHgtUlWFOlAjrmu
DidGGQBAZLOuQsX7eZenxpTcZRUwyEiLAWzWAAC9zXIXnN8jTnBRtX1BB9Qid2vE
zS2M/D+O0jvuWpDvz6M+cLq4RK/Dc7fQCtdD7BRksKi4t3KMgxt1I59514l5D5HI
hUXAZ5J++DjiJKPrsND8S0rkfhtXZ38WpnKPKRJaU9mu7g854VYHKaBeLhy5aza1
dxdc4mdR31p7RDP1DLXa04jGfmUJbDsuRC40yPSIJCbHacqkJ70IkePfZF1xzx5V
ck80/AeYgYUJLh9OOamjt6xzhQ1wsY8BnMQ2hI0ihyujWmd8SVxuc3MLr8cwEDRk
jxaTeB5Zm/n5b6dAf+P122cZ9IMAVfQ3+8ja8ZJLxTNRfwq8iI+p6NTvKXq3UPiW
5Lbqq1meb2VEvApRPt1QoEnKmiJ9nw+Xx9aDNvsnueMUoC6gmmVbuzrIYROrT99W
VCCCNLM5SDyxqEv0GJZdiGyCZfrm7Hw96eK3mRntDa9edt0HN07k5Y83shS3DhXL
wjW0ta8nPbOLZ2GlWNI8UcqxlQhH5KnKUi9QxSGllbgUGo+fBE6wYBRjlbfi6fGV
jnciAJr2DLMmeN3YEGAWi6DMNYyTooi55Jr7JRJhPRsmCytEUX/pRnp3f8jdIOX6
f+FMXTekshyJ3U4VTpbwAtMj/9Q6IIOwh9cLXx0mHzqGd4cz4ext30FXlyTpaspK
k9RBH28OgSNoT/lmjnydFrULt0W5h49LnxxT9jPBrPkgV/Oj0ZsWwMovPJC+RbiH
/tnOIb/UrmTIWU5MOmsE1n7lNzeGKpR1FFQRhb6oQ+EKvgqj79hEFYlb7SbEv/67
RwmZNAomq/HTjaEZHhwPZeq3UfB4lY+bEo2xvla8/VjsdBt6PqGxD3GHSqhgDYHl
2L8kiWMW19ow+RRUO3YR44JoQRrJqNpgnofvNM1ks7jHlF+AGT41R/mVOUtoz4wD
CEuX03LmLJp+f9E5yR3EfUfkHTfAK4QR1OF9sLsVfrU3pRTX2J6Hn++6WInG2C+v
UWYNJGxVmsRPNJalKBGn4bJ35pSBJ24vXHbRKEAGpSJDLTbT8IGXYAbdMz7CZCAy
KsGDE+M0nvY4Zb3GKfDWI//Xbg/4IquLxDwooaxOIMSFDGiMUp6rs0Hv5tRowlAS
x6oisg1mVgM3SPLcZdL+Ft2qoS4otBFKGz4/avI5iUlJQs8Q7D8a0wGHsnwVCuZC
vkG1hTL+5q+FQL1Pqmlf4Pjyn/R969AuG/AZ5jWls3rEWY4jORc3RRDI1/VAoQ5i
J4RCxweFVMNyQeq57oStHTIB7OupREp/hxzsRUO4XEXPLkOCBN4uDzamQDeZUbjX
Uc8RVtTFSQQshLAIEP8LaFtaY3bJqhvnqVXL8FRxuMOBzPoEdSEJHIaybzP0Esls
c/8WHXtaSzhEOOz2DedMvUxVTK9wxDw9OYdfk/QKh0heYqHlEXHoyQ8ORaTLLTKo
gKr5WJCL0CtI8QzQUBwWj2H6CHib0jTZ2DAovIS29cGHUwT3NdUasB7FK3mG16Kd
thdNwzLwmPivUiLcQ3M7siTm9AW+5bSL/tBBohiTNMBE/TaBv+FYjpM3CtYuv7/+
lydUgoHaBFuZU1M2psDepYToTLgXh9uX5lBQinLZyApF9Rkg7cVkYOpzbbTPUaAk
v1JMZmuHl9rcVx5r2Kv6mAPgTu8PHUDutdeDYraf3SFmcszMK+5JD+KGQvKRGVS/
xvPkGCuptVO9xYpPHATxygezd8dJPeVpFuGfyD9QncegdpLmadcGRfo66Ti9nzcE
Jwd3MqS24C5HhoIOr7rWkWWg6yB3s/8pC5NLLMaO0iR9wKLYZNfX2Wd+nQHuiZ2j
PLdd2ET79bs+vdp/hiWs7mbPN0pEfb3TYOtvtzausEw2hxt5ShfwpjPKyWk+6HMS
5bfpa7TwQ3p15sNsc9vl83sQYKxYzPxhsrisNYQeoOt0ANp99HlaaECRC87aZBkK
i9ZdIUvaTDlfg7avQA8qKJmqF2vspPxyNjSMFg8hzKVEJu9W6KtWhKVSmMjWQ+3s
aVKgghcrl24NM1sGJ1asPqL9z4RSQogz2sx3qMNAntHxrhc574uSkWi5ZujqonkE
uuWloUVqP4FQmug4BqWsUSiYM9Z7sExCM7DRI+1xU+fNLIoD5FnigAOSJKpgdDaR
GTtX/j0fa9iXJcOyXS6AlTBILl43qjcjIXaI6rDJjW5uUIJMIVXDvWPujU99VN05
gq/kkobSHuToxtXKJPz+Jcio8dZh5+fbph2eoAFJH9iwObOG1B/e6qQKW4UGfq7k
cb4oypbuUDoqhujVPp+C0pwFsNSXSiUNjAe6HIwjIPhy/BYlLUEvmmkZVbxsLe18
dBf9aPo4ojiHT8VDx44v7Gzm+we33JHz3Cyang3FVi+K5acTsN3+9dvoBj05oOoX
brfWGMT4pIpiePXBuXt2Ky+lz0G/YnyezAua44Y+r094sscGTrmMPiQcgvbGP31N
03IT+5b/hIfZc7zYuT7OvdGYIOh35lKSGDEqonQj1LJuc9NjtVTJ1KGQUJA4cnDD
ZtUa22qsLa1ugHNMEFSpMNILn4o9ImB7eV/75RiK1v1LFzEiB7pYumnVr8/d+3Of
8AHVl/qAJho2kmgtVev40zgMfnLo+rl83k4k+XZfE/Rxfy+M+Ey+JEz0rXr091vc
tmDcfpcYCwlPY0ulbcAUnGSMM+NdMa8zj6oLj1T39dILpYDHO0UPaZbsHQ2sV/nF
nxWDSWtwhfqMsApH7O3hD7d3MzLzRS3b8Tv7BR4bVfv+xWPNcWe/qKuqwLsue2Te
U5wy+1w8IqCzwj5HFc7TmVkFWbfvm2125nzSM/EHD6iyth7seiZJuOtafSVP1bZh
gFOVgWKX514KZjxjfDW42df5fVSX5xWBroIP4I9i1rFvwy+LfJgmcJ6cyXF4QcMw
ydOprsXNKGiQ8soaU1TY5EKhjFmuptHvYA1ZfmddyBcS6gBltQYrFuAWUBHPXml5
T8OcAtYgyqMPHtt60wFDcw3M5OswLbadDPlXfo14qp+bh/oG/HLClOM+CoZyDRiK
kuqDk4i2Z1NC5kzXIGIqHB+NB3e9cpALTHXLxaRtnoXqZcS1eg4dyIP1eyIS7XI+
77Xsc3pzeAIJeg42UCLFjnqJO6Jw+NHz6FT2L4+5NXMuj55k1gcTic0TNMC3gMo2
9CAV4GxLSPvDFXJx10WrhcZSvGk+j606Wx0N6l2QLgrdrW7Q3uvygOliTZtgJwHs
C6M6LuclI5Fzs1FQknlnQQ4ureMEd/oayaWkrynaj6AA9ZwM9AB9TY1vRJgWUv/+
mbGEXRZvhP8hCBp97YDJWDfw3Ojj9N7X5EaxuhUbyW/FujSDs2BCTL+0Fh5bizSh
6SmgbWzZxy6P2PS+sKb8kcnCazSre7Yc5ESblFbwgWBMoQJXDtIKI8Ur4tHCE+3j
T2QFMD3U/uYg7F93b627gYxob0iZ3yMfC486mEDmurDz2CWRubCeGQ9MWXJOoAtP
1+bxGaax40ebrwiWYD2sGFa+9WYxPk7ScZk6P4nNY4mPI34TlmLhp4uOd3kah87B
In/gCIGn7+P0Bn5jamFrETzKnYPZgJYd7P3Fmn72U/IHyFe1pQgo518iDSxPiGEb
J1DxK6AzuNfGKB0hg9AXzkHfVd9jkUYUW7ow60RNCPoYN2gNoG1NoaF3ubG/eJGm
7cxUibsvvoOaf35lYcCSeAEXanjWc9s68sLb6RbOpA6KwEY4meAe4kFxpXWTRHKf
BU88bNLfqglYna58J7KdiT0cZSDloOP+w1wfNOdKF//mow2GQM938GIbHwAhwoB5
PmJ6mRH6akMpYXr4UTcF7hGdWLCAUb1dzE2ntZSqwYLDbP0ZfSJEFkpSYuiheNJh
NNHNMpi+uhprriZr/p19jrDqPHXBfkz6Drsx9x1lPNX1xd7G6oCyGMUkpn7P2UKL
wB7SAjUEooWw4l0VrBf+AtqBq54EcVFWTbC1Pwa4AW2Xo8/ZCaLGZg4w6XbHL6V/
ECBBMX/mdk/6sWyCYGBCAzJW6FIhgP6DMVWtXNHUHeXSAfSJ3yg9lW1T+mCCeJ67
kO2xckW/qQf0qqV5RcJ6nfdRs+ReDl5bhy3fC+jzz0yrjwEXQzVlKm+nQYB8eH53
LqLoItG3dM1/KG9NzasMP3/JKRB2PTWnIMbE78ID4qbIjL37C7gHA5wxuiZ1YIc8
z7Ay5+qpQ/7J4TpJNwKzLH3y6z+O0gQIPHnp6OPEY3QxHYLy91zO0QF1I8zFUXWf
r3AruvhUhV/bEKbFQbs1LA726tp8mxF6YEkuYxymqCyxorulmJRYf7sxm21DfG5w
LoaWSoOBODnxruv+7yQdIPWy3yHR24CFuxbvunhXX46v/D7kk7qJkJYCohjTGOx6
rcNHWeBA7gf9OozeO79A/7u+Xm3VVQupSP897JtSHNYtDkBxYXBcjnwroqdFDHoq
Vb9GzilCVDNaNawNWgicqdia8k+Qi3G1gzSI5GyG0fbSgF4UCnxibotbr2cWgB2F
okBGdMRC56cD/DL0Z5fZZhVLXNKKNJzae0MNXTaCet1d5uVhuAcWszjn0T5gpCwZ
V3YnHhWYi8kFlUdgC4UOrHxzGdAEwcvdD1amU3GYiRzUsQ8D+CNDw+zo38Cv4C7V
ZxQu5t5HiuYUwFpG2Z7gZP3OEggRTuX6NjFVZ96WkS2eS1RiUOxnMphSEWzL2jpX
jWqyePFPvZXHpSxXV841bMEVh68f3UzogJQ3zOVgAPYrPb1sU4PuOSImFzP+ZmbU
tJfWoVOsnl651XJzHhDl8tttQY0gOyTQbIXqAg2Bayzrc9goiFpm0wtlA3Ftc7iq
aVugn9qu0XuhsDNHf53tZmwgEnrOxg6Hi7FJcgVlB1NCP5mSXyzfOigN17gc1LU5
zuGUEMBp/G0FczuUr8xdd2MmgQ54+5ec21jBTr/VJ8jxrHMx+EaQVP0tMyYKfyo+
IxrgjW8XDxoUq/W0aWFBLPY07SzoT9WZbJ7reEQzKhINBjgibXiNlnFXPTWZEzxX
ON0SueTjdKqR6+iYwEMpDrQk0bB3w9fpkFFBa7BG2PGTQnDDPI62OC32qSr22bBs
zoPorLQ96F/8vWjrdihNWjztAEBU0cjdQBmo2f82WOGyiGOoZzS6l4d0LSYspy+R
Xd8kihkS4xJsnmi1ThQhIzW68RkSP6lLiRbsVjvJLM2z4ujJn5vUUO09dyleVh0w
gv7MpRsyS6eMiU3oDEtnEd6AYp4KLtfIrPMtf7+HjiGcTPRSvAh49PUgbhN/ytj2
uPbWlPERwcXFhRP7eD9BadV8O/DGSwo8jBwHRm0rhYRvn8cO1if6gHSz/K19ONnM
JBOdfVtQ9lTusL2VColAh/VA+hLnWkpqlPibqtHJbOw2zt464P5JqGZM1/JVEcz9
bcjudXZCjHzc0HVjyCZqz1NqwI9Qt3O+YWWKek6Df5Cwdi7RSeQMmnWWVezDMtq8
/qjL2f7FOaOI4lzMOYbD4UoTYGpZ1WyJTRUeZlyZAsVITLeXri0T7baO8iRieTK/
NE6ovh1jkxuj5mirXCjYy2ZO5uZc6Lgk2ehsGdgiiZRM3zcrTXTgNmS0qPACh/52
oWUVV5D69W//i75cst/jgU/yDSxNedxqaPJUyf+CUCKDbSKRfPuHVMGfp2lvV2Jc
SoQv0GK/bZNcGwdHeN6eMMc8rV5JAxYmHYdjGiido07lOdIN1xMVSLSeoq8GtBAI
asbxkDB9fA1909o8hHes66g0lrZqQswNGZ+Tal6bAZKEO4NRFuze/uZ+vsMR55b7
JzrbMIplPGhRdppyUu7V/fbMe4OD+nEaIzRbuXm8M0AUh35r6HljUbNJ1ei2Qw3M
NS6+5QfbSRmJ0zHrIhzgJYJ+9zCryoaUuq+/q1Ep2/eUP0VoZ/lIGNAAFT65g7hO
GXyxVeQGVXeBqKvvBluZEE19HF5mTHzskcELajEHF81dFuF/U1gnHvlh2MqHuPKg
G0a+0MGzbsg5DsrBFtEgq6Bg4VFm/JmGLzxiWBsgdHYFYVBwtZKsVMyG6jl5T3oU
mdSjinIONJUt4meq8fj2pgqQQEG+mjJXBfvHm5un7sQGokUEfnJVOy1FARWOAY4/
ovbbeiRk9ZwWZf7DadFYronKZ3V+/LNu8qXRDKboeS75pgaEfzu9tKrUgErNC9KD
F7YLtLdUA+EdjkodBF1mYtghkzs20Jbzr77c2GCnGKDwmKJ+JjQdlO0cm1YO5965
F9f9iQnXzcXJPMafEkP9PkH4okuFM20mVlS+/mCiZCSedF826KD9EMIGPz4SylOX
fJ8RNz1RTsnNEPPyEzU+1m6UnDzfQsW7W8lVWgavh0I0Bli+TQfo56xr9qNRpPOr
idPEgy13a2aiOKBxbKwWRwlCXKzvHoHETDau4dkjl/nQd6+R9TiLCzQ+8b9rUSek
W5wsJbcGlpiKnekZSUqvxpY7dRDXMRZb+2FHKH9/MDYTeb829A+CBz+E9SPQYKkr
1GiqOz14FOGlnpA/YlFbz9bUnhxanecpkEAsDjTLyFphdaVIAeIHLiiCsGwiwkoK
9zI7S3MdQ15DiLg6cESAXWAJ9/ae34wgFbVsjPJOT0D/qWvZDNCxpzqBjU/Q449P
0LvwYt8xH4nYCh6B32kIrNIHn/7dvsbAmY8pGmpv6XUdQPw/MVbf7bo61+fVS3y+
9Ty9p0DNgy2QdEoiCAcFT8/NiJ3GutRsccd6S/l+ghFxIuIHzSbCxe177tmE9AJ8
FWub3jz3ch7u9o4dHUUjHMBv4nd1RqO11p9QUAzKRphu3Bh+DUJgmeSWWM1iYx/c
O1Jf+Ontny2c3+wN0hGIa+ip8zc4u8QVpr1hkYjdn14buqu1f7YS93/FT5/JHnsN
gjMgHXP3tSXwrqJs/H30d3NKStX5s1mqXkyLiIrDrccGvNk3woCti/wLpSH0V3Ek
r3A9N1VvYXunwt8wjRuiq+qAEPM9e/5KwQZAhZsX4bVVRJk0tpTubEJjsMfZ/8FB
m4wpovDCyLBdeU7a+aDX4aZsLcMpuvuyt8EDls3tcCwUzcc2/0Ql8cVZeP7v5ooj
KXq2bx9ve7Ev0RS+e2ouRIf4M7h35WLkZ7HPc0RlYwfFJguhNvUcz3nBfd29AmvQ
ulFmZQocRVfpppU8Q8jgwxT+Jz3mtofhLzRyrm/5dvmpBSyvbQYnPMfKYoNHKuv0
GiEWcbZ0QJfRcz8J41f/2/Wlr0NwP6TWFHKPg1rgH2oUjhBbbPQeYw+zIBzw+Y0+
vbkitQtp5JSzJrSVJ4ydbGVUwfEx5EDvRfArPYDBCQ2xcETVScwk/tzrKl+A8GWn
XZ6l0ckrj/0ZOdntvvpjt/fnSGibArCz9KZFLk+JwaCK4Lb37BnETtCVdoKgXLe1
qtZ78M19Jp1Seln/1E1obtUiZBNNuYAOEZP9XPTIoDqeOqMugoaw1fVk0jwV/F7m
CqBIRo4ysyKNOQZ35HlDkqVkEQik3yptCNd4U/vJtNS+AJOW6KUrWwuiGPie11in
63ThuppRIJqX90+kC+MBn4wPyO4op9pwW7d0ek7HL2ssfZWqIy26I7JxjfW2Iy3a
A4DYce1/lKh8hKYsASU7hHPzw1iD4scVbMbcH+q871etzeTzOI2uy0CFtV7fgM+n
Sf+7vTuRZWEKT9LrR4t8czZz1zzDnQlRJLTwsJJYDspuDPbzhBSuNBxbW4nt6naC
DEz9pt6D9IGmSIiyrjppyjEfWFKZtg5S6kHBF8hTV2WBjrcsxAl51w/JEGp+Bd+v
PSoR7VDdclyUjvCp3J2cKjvjsSR3dHhJPRBI1bF7wq0sJuStaWjefH6kK3UpOJUy
7kil6OqvxuplEKd/XXii1Tm4TE4nztHcaVcslKn0NNELsAZn2iCp0B+X/J0vOvbN
F2hPDe+nom3v9CNuSesmBfi64/Jjf5/Sb4sf8WyIll451BOPibDXxExJOy6JDjtW
2RHRQT03BwO8Ug9l5KbE0WRQpkGYpkpsrz0OwmiTE8sUyfOER8UxLX1fRQHOfoJu
4zirRgowDM9LgFgjwqCBupVROW9pEIaeHtvsKpZ6WOvPkcF71KwtcwPz7S8cspK7
EDPCXUTmrsOF1QgMKtztJwK5yAC6YniABABJxkEQrWH0Rbv9cwipxR2h5Xp1wTeI
Eq/ZriizzcWsIPUxdOoHHv3PDyj13mOmoOkDJaw9QkLUF13P4JY+CsrOvSlh+LI6
Dpny953PzLlv3/xsXRt2nQiqf+H0vM9xp+blZQQjuTsxJu40nGY12AGFqguwlfNl
WQChS5LRNeY8rsmmQ9L0Tj7yblC7aKK0kT8ybuxD2BWdIoFWpZOjAiGbngAzQK2Y
VpxJ9nsG9FkgJdRUdaWE1w03BlYrmmRmOFyif3pPMMwl6djELk0gj7uSFfjWdlxg
jvtHq0RGXeXVDF9vAT1omTpcwcbsfBh6glqZnACHovE1YZHll/vVOs6Y8s9Gn/FO
k+dlDTq6AnyW6GquswvPaVaR90gKeaxfuqYTSu6RPiGJv6Opi7no+OhQhmNCS5he
Ysu8L7dL/vfKDLAbAvEX/LRJcRGD0avaX5c0dtJ4CZuBl5CkOsuqgXK8zgnhZkaG
0oJuHG804VokPbg1H46w+ntivnoQ7cMI4jP9PHhiTIAsv8KX4TtrGkNwjTfWXFOr
PqVpf1U7h4ZZ6l5zqVIBQ/ENOqzUWdTvfT4ccSgV60qB5L67JzzLEnxTFcpeMLPO
45R/4OwRJcdw3pp47JjznJC6OIk7wcGThErttID8dvaM6/K7wLDOHZ7KY9gRCfWO
P55oDhOWwUfpEIJkdWss95HEKiUixiVjflngj2cxDQ5fxFzEwUqTc1E6kBKSqIjq
5ctsDNmiJkKd10pZfxaeVJHZiJSEoGppdmvae3f068At0NE1WtVa4C4ouqx/Dgzj
6u43oyszoRZ37pCHaT8xwVwMGdHpUqGj9Az6r9po+GGbJcDxR+jtyoTGFJgjkLfX
93DiVs/q1z/hKxzhl4ybC/3J9h2pENvMi6whdrMh1bwOxVuleiGs1Tvs0VjsAicD
UzkR9lR+NXFqLXgM0SskJK4uoLbgUPJDDo2r4Ib4Dare9hQ/wETWZqKOaowLa76J
iuaOqSnosGszg7Sh45DphgEGOZ3GjL6274tCD+AcR6mDAvWd7C39kcD6BUc+Ziiq
jKXovUH607jsiKoBYBCqOOFq9gC2Hr0nDUMXEP686W5CyelalSuInHiR8zLBpQAc
ak1Dy++rXBrkw6ZfFksKPGJaDoZatsW98QBN14JpnPZQ+Jw4fvH4Cu5/59pUkoTY
7DlrBTK5NNTV/kYnLgIM016VnCSf8Mx38qbdFVbdiiKeAzCAQXpHlg/mUSlq63a1
AwG3Dk8l1iU7DevT7jqpjd7X4bnllJg73HCcNcYAgin4aFXIv3v28aCZdKTB7jBR
DUs0xgZN/xFHcfX3QhXlsxqOaw4qGyANWVqx9IpF3TQobm64yt1GqvpwCZAj4/4T
x92YonsGR8QzY3Pw8HAEQChm5UoHE3Z9E8uefy1/AI7WhsKkArdD2rJ58XM5UwAr
BEM4lhiSz+N42K0VDRNeWRCSZwkvdXuOTpEuuqaHCCuJyq60qrUMpxNb14eBvHFA
5QicgCrjLbClmfeDTciaEFTqWRwfe6uHl2gK0Awsg7krrHzUlNls6UX5oSOuSZMW
7lVM34poukq1g1S3AEgdCfer401ySsL2l5SmwWmX/PHbj7+Dl3gNGEgDxwozhdic
LtlXy7QE4jkrOUWPrvXGln8YY7Ow8kh9ib3uqjzfUe7YqOuXUPf/anr4txwSaw2O
/x21TNBj7JVSGCONvEHACFaP6eS0bvRFlLwdIyhXyjjk3sGAcEKXhhzrFtrnwvZp
qdt8AmIVcrIshyqINenye5WOlkgrNAU+IBejF9BcDNnV46LHFhTNoaqQvQawInx4
RVFrw6mM6YU4zyAgClO4kkhzxfU1yOSlFeFTGJT785UeKeKJ5BhCBjZSlkXhRpY4
qynOWdqbi4p3aYn9tTKl65IMAY2DuI5Yuomg1pw4Z+KYCJmjTQ6HH3+mgg8+EeCO
E4VwWhJyzMuzAfBOFNLLG5BLnu1QzthxjUErGs9tvIFJ6ulW1FgJF2thMZL59j7H
1fO/SBtmIytBhxFJdztCoUIKtHxwpl+/n0DEkdOBGXBCt1zev3w6n4HQ4gZyimXx
pxCTAKbCT47+yptlXoO0THmipFNqW2mHwACoqi/PPPuOuD/aTfwSRhN71u39djE7
df6YXKFTJBs6IKU70s6mIumj/Yqqt9Rlar2M4bs+emlPL9+8NdfaBtZlap8zfwMY
j9BdNuyE9Mq4Xp8MQrrYQbsIvr4/so9+ynUnARDqkKya6idaknwjT4s7y5t0s9KD
5yS8RddaX1cWwQScE4aLl6jPLxqrrmTSdYXaexDC+D236w25KSnHGygtex+pqjJo
SVn0IC7wrYpHdDJF2TLQgFzlNdOiWs7uXSVCFnGLKDdgN7McvSxWgQwsWxKFCfCh
LbIxzg1DTB5S3jn4CzUxtayLszLhBkb8cIx1ZkzASdpeija7xfChMgo9T09Hf1dY
vGOIshxEbkBHJtNFtmVoieGnEMWyGN7cj8a/q51H9GvHA7LMuNAqv2XkDEN2OkDi
l47149oowNnHFUZ5dvbigRN6ReE67dRMke1z7gI9ITl7GX01m3f9Zv45HoWRRopc
MZI+6+FwOu9HZ/jgMtuet5AcRZxYKzXC1QONdwna5iKIBUBK8XvXqiGzVGUcqPs+
7bfhDCfBEsm1TGL0spO+bm8u9yRt7kwfpSKe21GhCsBAp49Dda9e0BNpXdHrLWzM
4Ne8ZsABNIJeYNztIeTsxuwN5W+lmidRrorQlOykCHcqkFhb9WsEdaQrYCqb33U3
3nA0wDTdUqnfz24F0yO6mGPn9YA2OeYPlANyIjRR3tY8eiL4MHP22XJRARL/cmK5
RNgjiofyhapBnV57QP9aBPyGRhgxQyvGkG7DrWxEt6aqhY3lfDA7XngArlM4molc
C7y/hrcm9CFb9tNwdTzT+m9oJFXhvCFxGly412uUXwh5ZRghx4eUc4pA6uAELXW6
nLNAr3Wluznx3w+wW4LB8RF3DAfFJS2lCM7eNNH6vdtj/belfHK26HfmHoLCmKHA
RHNBdUiB2CTCfth0LaLJAnJtKKhSHD2LakdCdzp87GhLMbFCLCYspI3QoYCtpLx6
ryqvWQOHxQvy1qRCRBTz3wnJJpi1USt+CaLKbRdHyhrr29gcW+cjwCbqvSZHeofr
g0H9VPYKgHWpsPsk1qGjpNHjwWRspiH7ZliziyMMWiYIndSRmKwn2LPHUm2Xx4ch
mAewnF1UHhHMjN4vryMWVdiTnztKNOJ/kClwacNprClQfgi2be34Q/uDN8n48YG2
MGbzW+LutSr9YE4vzaNXASNX7ZLTa+3AWhn0LZgJCrqwgH5Yf10cmxxI26oKmZDw
neKcMXkC8lQsh1gdqzQqFRCmNqJ5oQlaR+F5MIy/DBS7u4u1W/6bpYh7yRvUWKqK
41Ty7uHyzHQw3b5s4cHYUo+3h9hDeHue7h810ySyf5ansehJftC+ou5Rj6mUBjCZ
LT3o5MlNM6mR5UcRd7GghBuZQC1kKualETJHS9zI5cb1LRWBKO0pJ/ZQgTMbug8S
qhzwO/QEewuAUYQ6XBHusUxsvG0i6EajJ9fW5qzV5T+qQu/zLB5wZWQJXh4qZmO3
cL7zj0dMZvHnQbnO1E+U7Qqo9qo3t4rJxkIfTy8Ut1uiUg7GVDapDAgx+6upFGr4
bkjurpTj20seT8ooIr/I1Gz1TrqIaw+V+1sAjAg3MXEvKWNneZoDLeQYE0nSnOGj
fULrxZU866jOjb370QrVL/+dLY4HdnmduhqTK1/igyaYhY86b4TwaP0xwgHnsI2+
N3kBd1mviPrBYLwFIPAHWFvXarGAZs/U/ZOUInh1cu1jGYNBq6nJDrS4v6konCKh
ozsviGBSbcOSddzSMtRIH+MI59sRkbYIVovW0ZBXgoMhJ0lACNZ+pMC/4wdwrSyI
Y5JJZPdV543Z3OTth2Rcj48/uqT2CRSAs/X+5hhdWUkDkIgvjWWGuFCqy6ngo7l4
yzwRKXVxbUXZHnmkSA8Y+t2CekgqKMzTnPRYzy7PGr82dlAz9a9OAvbOWKTf50gY
5CcYTspTo1aB2tmtW1sUmYv4uFGllRjHMbYhFErfXKptQ6Ol/39W5Fm0bZog0Vmj
oWe/RXAhzNECe5QAFRVkn9vfofl9FJ4uEMxYRee2wwxzQ9eIJHRpotBZdFtreY6D
qOzwN+QF6wNBnfasqWAbQoUg29J/DQxQxm8OkFjR9x84n+eCl9MDpfwoiXh4XsS9
+VlJxLJOQ8S5pcpos2pmSBDZbsPA7KQNC8BcdwUS2IGQNZ5ax9LUC8OysurgGxrV
fDHem/WYbGall8sYwtCkgubpRhXiCbbOvHG9zpq9+tf59kwY3rbZAP0x4eEG1Ahg
F6W1Q16oUKfCoG9/TJ7PVa+x6Wang+U8xEAe1wObTV/w29ytu4LJH0gpP/t1Qpm6
7xR4TN1aT1K1FUKkG+6jWOcTjwmqHXYA/079eAYk5aosTwnn4QEeA7Acqr9Xrdy+
cWbblf7euH1nOwFhqILl6JAjqqqC2UzytMVoUJQ/ILHwj1HJgA3sGj2uN9cXbgA3
/MdPPml1Hr08lvGCtrUgwzSNQf5vzWBjE58vCYKO+2RURgCW85pclEGvdLw1dT58
hztJDzoyEnyhRBsoMMn2VKj2zKsMv4OpKl16PoQv3w7bkzjfEzM1h6rBDkRm3cg6
8V6I1aHTI6PMZhq6/yQo+p6mnhv+A2sGpEdz6WNhj24+s67XF0tsVwesj8XJjYrV
jkrLACYVQAUeZrnwO7JxZlBEaVdflCjCRD8gJzzJ6IocqIhIqF9gPl5s4cVMlwQm
jekXBHPpgLRA4m2bsIDcKK8oljZ7QDmUfRKIVwE21adJsrvvJBTHam23MI4LaRT3
Xxc8YxtD63Gj3FGgPwSIrXQJ0svUn+TrWpx23oa7pdIPEzJXOhzetX6qALR0Dgxp
tu4WI0H5uaRkWDTs43SQr8AAkAew9/CfFeyfT/cHqRQ6z2V2ca+K2EnNF+Vwdqk6
SKbpWYQJlp2aTP9hyyMLiGOFKqKmpBHWrbSwPfRGUar+0yyUs4TKM75lOq3UDpL7
4rPdavofrkmwixg+RZ/5hxs5iwrulbjSq4u8eSFMSYvUnCYkDfm++2jfHOydfnKG
7Q2tO5gL1ZdOuS58aJMfr61lG3Rkk0gyvnEw5T+q7fo9ra0zcO/CRSYeCD//guxO
HAkELR4ButFLdZbi1ZoT5zOW6evePOfcDcsvMPunUC6LCy4TDXazJN0HT3/ho7Gr
u4LWTssLdE52LJ5G6n4GTgUYhN6BKlNAYLhttyuDGh0u29cBlhgVBDKrOj69Yogy
Qvs7N3ui9OIZn3UT2w0wTgv2a8SNN30oGX3v4y/et0QNWYqLCcANrccIPT3CixnZ
P3/8Cf8FJEFHsn97gFebEB3vnxLJ2W2fLG09Xa84Ffl8MUavX3tI4kHkdxfhDmZ6
ymwVX2IzYIu32nNqqWN22ooPqzsJQw2QiLeVdTU4YNZZtTO4t4/ZMHDGBNaLbaRl
W2+KPyUnz5rF5cp7LeFsfdLO7rMzsH33HFqYBgl2vWOmjxSzzd7IbYv2cr5a35f4
H94q41RDqKIMOnXMZIkwA6/cGxXlJ/83F31QBHOdZCGJi7NEJz9o0WINc+aOQZfH
ttJoJF6xuiIiVy77B5l/Y6c0hhoAJi9q6BpRF6KJGpTPX4odxWuDphRPlkF06Cpa
C3UQO7K/gsxtEjwM0KukFr6VIr6FMJ+DoetO7PO+2A0naylxtKOwPg5cTDwSpc+4
hYFnZI20sqhS6FGYvohZu/aVaw7JuGDG/AIlQPST9/3dNWrVBqunLbTkZqUw3LFn
6gvFXzhZKPKTs818T01eP2Je56+gmdiPamJDu8KOtX+mqaUxoXKqfsY0bVZh+8zd
7rFtvJiqyIbU3GlGg8Brj5tXJZSF65uyrhkKcgfzfokMdZmInTaqFMjL5dvzO4rm
Ss0SMC60Bq1QVIL2ogPr6XFKiIvvfvluWdQokwUcNfBqWn8dw62jXjNv0B+5/QfB
0+ilX7ed7eBMSl1brNnlf1ovNGU/wvzaoJ/fwBXKohz+Y+ieh0ArDMavw7Fjg+t/
CgzYFW7suKv523NM/OyqcR1Ej+vsGIHNTEE4BqK6Qisk+hXw/P5Rk4t7DQvTIy1q
LdKh713Man7NVS93sSSb65+4euFItR4nJA4SrGDY07EQbc9VBRko+nV8jFG93Fcn
am0h8Xfq0FYUSQzCmErQyas88t+HuYnMV+Xhdq4G71VcEeSR2n3qBgRlJRUibHe1
J+4yK30Mvs4hfrDl0fw9PB/sZ18tsEUneXSNG+Hf1oTidR3+LUmga0qG71U0u+vC
syk0Wr4Axu6Lw64eVzI0qD/CFH1cdGWda/5fhntMWnuMpPdom/tDQbMxwPWwIoFL
hzSKIB/Wfyoh98gcFXXkZwDQuEI5onwTZ+y5Uefriw62wWPho+tbb3LwLaP44S48
LakZUq0nAHc/F/y8Vax5xYAs7IZgZC/rz+QCJfQiA2ISbrjNjWq3PnUOiOspCl/r
Acds7px3jnx9KAM5OznI4eiAO5yQKXVKxv0/UZCOIBtA5YGy0xeAAHIBGsuFKcci
BZ5+ufawCd3FAU3F3NIMKbpnT8FQ6tXBvoRFGKUrGZM9JsXy+vrmGBGF86VdRgO4
bMg44dhyizrpDx25cmU8cyf5YlO4nP+g9Tn7+rvifEn2lTn4Vx3MYDkGXpv9xvJJ
QmzlWrs0LR5jpGObtw8yS8AVHiNk/hsrSJb1/EOreoGBV+pcCcpjL65qqnP6Ymdi
E5s1Qv3WVMhTG31bHvVPAeBO1Lbpz0OoxU+33FHnRnj3RC88njDNR5VOawegBuLi
XK0SzTS4X22BJEVQGnFyfan+PvzgkDN3lVGiDSLwJivXACeMuCs+Xw1se2s06AZE
ffOWr/dc0W91qoadK5f6g5UClvl+eslV5aZ3+HX7Jy0t3c8LC5k27k7AiqSbV4P9
nxp/o8i0dAFzIXLfDUhTKd3eY1ojZUr3fsAxKqQDMHxRfhwb+rnNvjUfF2wJ/CZc
fWsGrBwMFdUiOpj0w61+0vY7u4zCgTXM6ex7C3r1oixPvxRDzCBGeWjqHV2QgNS0
kzvjAdvF5OshDdjos9kswlBXDtebmwxntcyUs+H7xWJFFL0LL9PZiFGlPUBiCgFb
fX5KgoruDlTKktwK5i3p24cMfgqbMC5GFG6W9UY8WOcVfCv6iadx7mTvG4IvgTqB
JjINlIURPJWRKlbHquHEshCaxxkkz4GmvpJd6PWyd4KWIFN9ouxaqVgINhRrdG4e
fu5HKU+vS1WzvEf3VkDA1jT3tjOSc8LEY6k6IV1HfBlzd+jqSr3AM81W0WBjImPc
8fwsTJpC/8SQhGYpLRxUxY6u/X0AL8AmgFJyAyp9nb6zikuETl3c0R/3TapICFVm
dcWmy/GnBfpQrVgkfccEjNBawvSkLOiY1a+AYYPvls376sVjN3FpVhdis5PfmwQ8
o35pmS73k4DWsP3j1+5Mb4vIkPrBqINvy4hrxOp6SWknc1Uhdry7+OnhYX6z7uhi
7wC8Q4/DX2nCMBDofgc3gFQDoczMc0fo77rGzUykd7uCRa7/cTpNFT4iAfy5gbas
v1vdVaZaeVtFAI8blP9uMNeulVhNwD13MSkOnhviupTelOThqm7uUvYfxy64NOeA
5wZFn5dCiVLskcF1JPWLeTQRjVKZoEWMn87E1f4vz9LXbQHjxV+wQ0GeTtWQ6PcF
ar5vigxdSxxzWeoL/5Svi4h0CT0qxVocwhJ6UJDjeGruurawp4OiVGg5PntSd5jM
/ZHODNSa3jtTz2daiE/HsjTQLDUiUrx41zwQ6qaqy2/8MCyu6JW3W5yzmE6fF2Fp
3wqgK76U+eES6To7GgheniT6FCYZOG71wy3LzC1XgEkWYzYcigp2fykFRzxB5ar4
1qG3a6V4JvI26eqTlps8U/e6j9yWhxdPaamBu3K585tTm4D6R9xL2qRNZVepnWgf
Rii5bEWwdGmOWMnNc2c5DeJwnYGuBr+Yt4h/pXdnhifthnCjgjuz8abuLLsEGVJ2
QMPyeHiWiS7edNOy8psA4XrmtjrDhxqM70DqUL8ekOIRmaPAuHjAKpAh5p0JJZom
tHJOzDtnCivdcPmVYhuHqRuW65iFKssgccr4yU8pxc+Lf9OwE5EwR8wWmJRb49j2
5WC1ebuVGXiQmeffMVqK59fO7spuiP8OJnKrEuYUgdxCjQ3428uLSrbr3cnjl63Z
+cGpoQpBcplJaCIVZPeOJaoqccSejSo7eaQvVtoigTx0nHP2Uf3wQrLx6slsKeK1
i/1q+yVP51YvimyH93Th/u2p5ZTALWw0QK04lVTvIh5PfgJjNYSq5fCnPK/lcOU5
HHmpL9TavcBofUe7jZei6CicTKRR/UFnNL5rOUZ9iT/CoqpV5nuT4YpTf5tiEJNz
ahIColzqSDwz9v66YhgG3jX0dMO2vMJy/Pi58iHJ43GDYwMhRjelOvByLYQwk7Wk
aXpOjyJgPC5z+KfuzTs9vF1FT4Df1lcp/uwN3oqwAb3NROYzGyrH+QFiywBQYyTv
vAERCnXIsoSE/Ek9L5hFk4zD0LD+nNFOxFgrzNdQAVMla34yf7V/5Xkw6RMmx7tn
/r6wmimv9tDG0PCX3U6UPFBpfWma7dUSdo3AHApaqeGh01wkUF/Hct080ouyqhYx
ZaiQQPxPWKiph0P1a++LUIUm1ELqHMIwerwHuk7wW9eAu9o6oIpnzcekCLaH4DPk
ZqzaBdrB6818K9Pj5FeBrItG/DyWeFPJBl+UODvgv1DbWofehHfuuo6biGCDmPVu
+SjeRbP0c7PzI2P3U0hHsErRE3RIvZbT8OtBKkgcMbcSgDfmQbDTX8dSK4pxJwfp
Buu27yTb3GhD0Ibv4Q2/4rRN7nj+YUCs3quRyB1I38R3W6ljEacx4Wd794KxV3KI
Ejx0ZTBHq4Jf73uczE3UbGlo8JzoSgeRp/Ffo+Xbu3W0/JiEwq3Ihhen01bc2wB7
/F0eHvyl4THTh23wuSEpUCLA9DP528IBVFf80Cp2fmlvaBRjs6b8zA0WqQfUrGJH
ePY0ytjjT/kK8aEteGweSTMK6vFAgIJdO1dsz10b6LxoaiiHAMK9K47YzGs8WPW+
3jfyvptwjhfdfNEab+dbN9YQDHIFP1RCH7+MNbNPRH4HQKZTUsNazW7J6EjLf/so
NWx0KapMyz3k3FtcVi7Ici8XC05oGIWrI7lLapjl3WtbtWJQ28g2WQGUCsJO/BB7
DyRrrTFJ0LTpvZB8ACY5MijjglgPuqAGtriuUI4ENhy5hf3212KJ5RmargbepxAT
FHMb9w+1lOhxHDN3Ykjndu9rOokWgK/S4qE5VBkOo/N+QWZr8y4bVsqziJWmHmQ3
smkbVmZQCFM4gisjPgQgPdsWKRq4DSPjoVOrZHmc7ssPv+RIXNJQIIGCrUta1MDZ
NornuozznhJOPO7fbWPIbn4E02ilOqhcJKTJ+mvHIy0NtsWIYOaXZReDhWxwRLUl
o2IKQyxGkRNCrriOl6VgL+1m/gE43FdemcOy/vQgZ+UoydvQg+Av+cayDBNDYNF5
rYJ6AjdQQObnMxNCgBvWGSLI27lN6Sh7vYsiLXk0rMVLh7u/NWJzfFBx04dV1158
CeH0dE4zD7r/c7d+X5k5jskmTnUGNtvmhnLtQ+Hefr+fLRORnMvnE9tOEzrVS7xy
QLYg9rBevz9P6qQZcQwfGhym08rE4rJ/wz0MtynLChZYKDgqBF3b2EyPbmKkbKe0
5oSyNelwvyddrHEx3qHHyng5QZFx2X0ffRkomQy4dU4zkh/C8tuQYD8CoWSYtz+u
R5ozeABwgaA3WwK/6hnQbN6n68xoldiSn1WCHH7anQHd43hOobioMLdnqsbNeKrN
Ry7sOfgdWTu23Dd5se6CRr+SgZrR6HNHN9CZ3LI1H33ONAxjY8eC/VwCsjy2EIza
t98tnC94YkEvO0UMKe4MuxsPs+BPDRK+ikdr5WLW2x0ef/fmKhYaLuo0vmQ0qf3X
081lFw1bDyLvcSyV/aM7GvI88UPV0eN7tbFoWEVr4wRXdBlggaPPom9iOYh5qG1O
kqyqrDbA+zQqGml9LIKxsWCQbvXyHjNiZdXKlqNvCg3vEBa5ldhm9/YjhBbWxSWm
8LSQfjQhc6j1wS4jWIm1vobAdVIyOqPamCvtEqxWtQ0a3vw63fHvFIpCda85uxsX
LtQtatAz2n6ji6mRge2sSz1IbDGEgVvXlN2mawXrzlzxfIb1z/6j4MvuuFauiU9w
e6xAGgSAbetp83UJnH0DKaxrYXvR/MR8npmvrAnBuTtvvzWa1mhTo5KCfBGBQou2
Guy7bFWizGm+LHO/hswK/PZS+es4P2qXeLknTH7afi2pUQfjUDReTF5F2pweyzII
dq+LjSktL/srxheNVBMzLLPZEa/hyAO6Ycrvot1r+fpw+MHtv57+eiNWemkkJVjw
BhSES8xFTJrsARDn7Bvr7axn8jbZzaiFpFpIaOA9RXlWqJinrIiwsvGYnc71P8wr
u7J0GIzPDPphoFvqts3b57MYnBs9e/CDPaCsDAT9jnEIHkmlCpeGzlm+GMUoWr+j
bf5fNKAcWoS8nc2N0vVK0LHz+IGZnQkiEKXiq2QOPGzearMNbcW2Pje8Zd0/d5I0
It/oWeJaWcWxFisbmiraxOJS6lUAB2uUyay1+SarUCqkosHgkG42SW5If9kSU3KQ
+cOKAeFJWbWpuovjB8hqKMd03BZV+xPmU3f10etTfPgYtoxC8LeCFw5/NETls7m8
N3t+4i0xf9amzAEl1zoV4lPdDDP+2oA7piyrs37lHQFRtSBaGemGCBmS2az7njdU
6R7IeRGQ4WHJ1+Gkpyz2Wy/A+qPlq8yVi0HrJNwoeeRj0KKCPus5yIc1e1NZxoX9
KlMSASrk/BCR45ssxecjqGUwYLqjw7zoe+Wh5JW2c6PnAoJCItzHBRAJX+CVnEvt
MyaiWY9hNz+jUPAdwcpnrm3wmnsON1MtMjIcgHsHqOVas+VRC6hbBiyKcyCHHu7l
MKQWiWtCcuH22GFRHj468y8z3bviCqBLOmoYacLcXMM8N0sfTnByZPaTwW7a8Dk1
c7UzSCuO8gkEoumqZ1VcueFXrZzhoBWHiwTRVXNDeUpU/zzK6f5+rgExXn5RLTRx
uBCGoscfA4V6dznPgmvdIiONpM2menSCS7G1VgfWi4Kv/jumj9PJHj/jd5TmpO4d
SKc1PydF+adOvhrEVc/ZxAnkDPZ+05l1gajdQ9AVTwliVPF6XopEj1gkjanO8JYd
FV0rvX+Qa1se5h+WyaLX/EMl7sRBUwRqPwX/DZAIbb+r02nQKiUcazgRp8koxUlo
etTAh7J8c5+V0kxlmg3byc7AsN85Jpbbv+xDEkohX2/QC79nsnlb8x0D8phc5sMs
CdGeEXbPrHOiMCiTrG7Adpw/aUf6gDy3G2WYM4188D+57ubaRvj8qy7nXy2rDMno
/m8eiLgt1w9C9PTama0a2Ao8Zwp9kTzz0Ly/enGqAJzrD3TRfme5OSg2sb3T/L/G
IQTKXzNdlntUFp/1bWuFvjJVUAvTpjBnSEr8DsPvhh7ooIwr7FqtuHXCXFvROhRh
UDxk6o3Arc8tbgelSe9AjxEsi2OlZBdNWgcARXpy+AZRMX7eSFCjrZXP2nzqepu/
v0cVCCmgxsSJuSvOsX4Pt00750Vu4jnj4uyv8wYQcXpSbtHwEqq2efwRTbPn/HNB
3BFIk8++id2IFsZN45+SqvNJC1MJ1DuZMxfcmDVhbe1Vlcr1sGsAyRJXdoza9TWI
b01csb8MFr2PlOmdnQUNkL0MEdA1OemTaK7RCNKT3UXqjVRFOB0B6HWV2sC3NRll
Npjnrch6FfuK+4r5vrGfsE7fos7aEgcqzUK4Md8+dh53Dw5ZG5IErN5K4ok4mBo0
xFF+UmP5XCjbu3XfO08WFjVBkuVMx68BUpYApEjQw78tR+wBs35SZDCbwT/j+kT/
aD1R44nzmng8osZw302nE2oJGk0bQ2g3qO9f0+LJsh0qq7fVICyi0BugTzJvJyTB
ivdMMCHzhnxT11RxE81Wekanj5iKILutf6uhPPX0W+LfNGoeI9aj7ucp7ionNTiS
jMjcA5X0n3Hy11xy3L6aRjhi0HfD71Gru4zroda4KA0qwMMxRSpo06zCFtLeR5Ll
pYU3G7Q9rW891IeEUITqactN9ZZGflSwX9MGpOTqB0KXKdCn4SQCfXWzg2RAwQpa
8nyzn7DzAQVsogfitPyK7Y0tbgW5/+9Wwhi4t3wxrkzoeypT0e/BUZ3a95r3ljOj
WdWsw8lXwuz7J9GpZenAK/LORHUftZaNF0kmLlphglLenYODJqpSHvXy40Pbn7St
3K6kqiOuIOgVvdqMitwmZutI8Q75Ob+vzuB8kkVBBYuDhLbwQVQd0ZhauH91h6ZI
1c0qSJyXpvFTYzk7/dYNnvsxliTYzBxJpxBFhpU3SNn1ab/CVcKOAhKzDm3yXziw
4OyqYe9/XWx025Y6RxyBd8cKMSXaIy8r1BvbdHarPAXL5ZzFlT6d0CvGrkUjnDe6
bOtqcX2gMMJWqCpMpwpwlY/YoOTxExzkt4H1LW3jlANtQUnK8zhmpQXYD/a/Qr/t
gN0aCnFlCeyzKmCAC/5SS0PcGpYaNhpOfRXsC4TiJiE8aKiKEyg16oEMnygzIx8o
wc2J6OibVkzaugG2yypYpRLTn0dEMpPcNiHnFoUG8estbGkqDvQJEzZbLnPNzm5I
85Rg8Jy9HLkIMGMfjgpEPDInMPbFm/49RlPix+sDjQzqFc0eC87q2fhYRTSQCEPJ
mLzxAcCGkPB2j6GaJwCRUUia1fDWwX2QxmU3RsClcCgJtU5ltrKq8UAYA02rgQXj
nqn6JdfXTCtxk5fRYXdy9TXUD1bs/9CrO4f7Up2FmMTR+r1TxS1DYWfLjB1joJcy
XrGn/c14C8RSH57rL33ntO6cAFb5snLpi+37NyMRvpac1sbN5yMQhNx60s7Vie15
9dkIPzBBs5en8qhUI5do4yzfS7RWR4fG7RpRnIojAy67ZhKRVE/73eTI0zJQalnO
qWXCbfYVwIoBuhqFhxttbeUxHHD/qZFbVvL3eaTnT2iAxggxpcx6rcoviX0l6gDa
o5jQZW+9VYDAnFGJZi+nQ9obhgpndb7k+evEEHCmqqQCj9O8C8gTK4BNSRUZ9a6I
C2WUeWJGzh4R5ZR+lgeRK3EXh6x674MTpS3PckYzhRNkafDwodd/opt19Vd9QueN
ijKOaX4sU9MNuNcOEzTSRPnY4q0QmU9hph+RvZe2bE4Apm9uOMAp6aYUvNWASvwM
4f8mmpElQf346neBb7twYsJiwr2R0HLj+FqDedThJWOhj1Ovp8irpLaB5lT5YYD+
5x1gVcuqaF5VSa4PMtkv8dKvnEz1IE8mnG9sfibmM3D33E76VwOuQmZ9igJaQfD3
EAxmxWCJDVY4XY+hC+oE9aoKnMVbZCjqzxE0UTNn9FboAT2MIwvVfLha0YOp8YUW
s2UfQ6eH0xq1dgWvJmv6ZfXHKGzyF9EjWF87342c0MvQIOi5Pj3Gizuvj25e2eBU
YSBb4DpHhrwhZ2sSK9ONLhgU4sOR9Vb7dpa7VhMQ7wtvfCDDJotfzcnSCdl+DvFR
zJ2TvAWJINjIU/25qUW4P7Tm0knFWCde6cNpiZ4MStqTR1bIFO/5gbeMInCWl2vw
b7Q6x8H+uakoTq/TQqwkjPc+foz6A7NRcczDzCQo9fw36zATdgdCO1e921tRK/mC
KIbavyrqKB4UbPga5HlL7zH8ghSBjCsF8/tCjFrSqRFWapz0OEl6b94yLwwburlz
JK5Y/KesY6LYqaMaV11uclzCnn5nszVlfkMtxDmUd3N2KKgskYO48cA8PybEIf5P
gmZWeJbG4hmcNFmhsy5CkcR7XrJ5YLonENZpiTSs66BAlD+jK8edhcsdLnce5g6N
U0JO7MA299duOto9IlQE12CEt2XYejS541QzjzjojMfB9SQbzPt8jQROItZJYLq0
n9z8Ktf5zWDLNCen3ipa2W0MtHVWrynfPZVuaWrUkvwaHj/hv14OoTdS5XBRAMIx
gmUcKvGTtp5uuWnwAWbwOflXzqwcjuIwDBfgOCErVi9dyeRHjWjDRtnbviZZbNEK
4y94no8ewcTAZYgu+vRuAQOr48mBswNMuGxZ+FmK/aKcLSQZjYoPv7SGcPR2FmTr
EbYQ4c3YbXierekgl2OvLDrqJdX5uTMOlpvSmvm5GrqcZ1QTE5BHrabZjCjHvJHU
WND6jcE0bTz3DjwUHpSOldJplDIwS54TYe7FiF50l0el3QlR0pdeMKlG3VoiwhpX
P5Q9zOjRk/FSUG71IWZlgt7XVoARIEY4r28qi+FWWc6sit0hHNkD4/6VETP1vjsJ
jGfwHqz2+Ber5XvgrT3ElAfVjJmnyIy8I0RMS0BLPyxx/WDXSYeZ5MExDo13aNbw
n9P/ACeKkIqL1C/UG1ezXQVmiJKe6CbCl9DhEv2HUlpLge5Sr+FpQr/osKEWFKI5
XJkNqiIeVP3BKxmawQ/pXCrV3ISDfTPuvOZmrYeegRcVIjIQHdYKOvSeDZv9iA8W
P/bwvjhIdHe/4F03x7O7MJGMLoZ1zqs+hDp2L9USH+6cGYHTsNoZHegTj3fKHhm2
CWeXGDP1v4x2iD7G+18uLZySbpKwhSdM3GNlCHKUg07KAxez5iy3EqFZOoW+m0jX
5mcS62OjMDAaKuSbxKmU8n8WN/XI2stDQ99lvLOJ+n7OB+XOnln23fhGTTLAI442
o7bgigqdetxpThI8nua6wDGI+7gQhM7eLSyKN+O08uCzfc2Bkq6Zl4yq2yJUv8Xa
HWoICTZqh1PFZvOhxW5H2UaxALAao2lHh4aMneZt9dv2vmon8Pw6xSHaSE+wab5N
G+RwxMZ9tKVtofK3EUHs1Yrh0/cWApDAvwfC0DKwgOtdeKShXcjKqv5syM8H64st
T+teB6aQPKaJDP6ix05fmmxvdTIW6+q3VXLcbdIzDvPkNIVqGNQ7106/hBHARCfU
Du5qpRT/KBq96y9lRv400F23yXI0v+twPfDnx050yStXI9zIXudsY/MmBPVGdm3q
A1V3kHUX7IEAIYl78Od14sbWm6tt9ELWYHmZZYIjDS7+zQJxAA5oYeoCiWqIj2/q
9kajSz6ezMuFhLHntKy1GuQW5wSYHGdZhu1tZa7DXUp9McY1Ugmw2r5aGWRaP2oG
iGj0rDa0vsW+/Sh+UMceJyPOHKmmGkbk/aqHcwLZ2S5TUAImjjK0AK2ISYYE2bGM
clAmrDxn1uY3ZX1SbLARtrqMl8i6qNEVhFtTSDzvxzHKKHGB0V8IOroP6opmCYbW
Caz+VNoXZUprmXmXHucAknPaqpeixeAcujFNR3sUKt8FL9dW8aOkPnAXT+4qJgBy
0FHE7ormEmFy1EzXQiF8m1VNqA/Xf4FZEgnv1LW6YwZX9k0vrlE4J09xvX6yiO8z
oCUf2itWrmoYmoA5Ykbl67Hayfb7iuAjvvoc0rHkSd8Y05qIUgE2/gM6ash5tR77
D/woiMjNZytnIKv/BqKycQpmYtSnxPqE/bHiZHETdOur1s6bDjbfQ8gngk4mh/WQ
9RK9vokXWJFf9MkHhsgi1F7iie7XV7sP7ptLNRVmlYIbifE34/CO/qNXDzYssvuR
mdClJIU0pYS5lgsDgx1Ak57YEsLu9hEcgiXYwR0+hoZ9PQZSARWNBVoYu0rtG6Eo
a525ooSpIPnhjVtpGIDCQEfbxTFNidWNmq3/wPwwQr6rMJvmbRdWVg1wHnHarFxr
3ITMdnakAUEonLAc3u3662CO8ntCrsAJfN/L4SbD8cHZTDgHMh1fmfHoJQuHBCIy
HA8kMad+BeCaqgJjTbdPwiyu01dHaQLtePqQbRJOD9nkfxV4dV+HtF20X5b8vu3f
rGZpMxPYVNC9QUCiZASqn9apP1n6G3KTPiL5s4+NYLuI/PluZEhtE8hp3SbP+Gsp
9zyPA+L7ofbE8JqytpONvtGC0v1u3hPrv0w/1R/XQrmsVy7ZBwBOcGgcsmio0cHu
s1crplnDUiNuQcifBNGPs2TWy0nF+SG4bDrO7VGyi9EtFGFqPVUtq+qitk8Pi0xY
mZIvE28kiY1k0icV7KPYWCIdZCyd4/mweysENqdYWA9OxYpoLzwRYzeZ46VDGZVR
r0NP6Z3+v5DlAjD6X7cX2eZ8avY5eaPbf47toMessiw7zvFY95nE7sedGmjOGej4
N+9b26Oz6Ftkq6SdE1J4Ceff0h455YJSG62/wptSJPj0yZYiRBAHIqy9idX7shDc
/bG263Mdr2NzmY0y4qZMnjGdkR8h7F9taSGqIbV2//O+It0AqTIwJbXD/FtVO3Nn
hVfA0AtC3Dd8aTWgroijeJtkKpU9sfkPK/4A+GPixqT8+x9Q/yuDyr5dbW0WtzPi
9zJ9w/umDCz2eoejCNPEmOtyqspi4MSR2SJlki0oEI8/CqkLdKBYOKrf+b3YXKP3
jF96OzuEM/QGZ7fhq9YJl1zRf23TiioIuTZlvDfxP3Pg3ISZw2R6oAAcXTz/Dc6Q
9WhjqtujaWT7F5Qi9EWrfURLh3sJDff25jr+ZNlTqroRVpASVXtnSu6pIR6qnW6e
ATr0LlkU4Ns3uh4wRlSNh3DA0eN3+q8nc9x/t3nsDAC+YAJkrG3Zlz4XNwsX1Cu8
Xffs9GbAmAJaHhTo6UcPlogFRRityUeuMX3ArtECOidjYx5GOzBQIZtiYczy3gDm
JESyOCWfC87tYwjaufmXOB16yV6SdAvFjz2p34mE+U8pM2mmea21kTnY3YZGjmVp
Zq8wZHUFxhVb26Qyk2JGfTLkpaDw8zXbbRwMUcyQ4VrdvidWbMcS74e/358KhBx3
r43kJO7Uf7mUJaq+GCj+sYU+XiZMCR/xGurIBCLardUiSqoap/BbECy1saIerMY4
ZCBu76MFkxFmYy5forq8p8eWTDZBEizzYFIn1LEYDlvBjYK3ktBbdNph/uohsb9n
Wv5P2+5A1ot0IJwXqsljBoqyjvh0HsW1EixUKoTS7fvTNe0rzcyrHsLNQvpTrRe1
jl+xe9KY7dYGkYtHqwNcGDSTjCrRAF2biRKl6+OtdBczIhXJo4oU20uOelluWD/b
7pMkeoXnH9Vz5CmXnbKTE/+i/HS9w75c7PPOVhf0mk9FNfVuWWSkXfGyKqETB1KZ
qq1rcc0CaotKigoukqIOco8Zv9XcorhDignRw7msM1zZfEbYrkqAcZA4HO2N4QIZ
NHxBO1xd0gaXxugFql2TUg8SpBQwBOIxrwqVm1cxT0H7YePZGLqmNj9eG++SJSaL
RAHHYwZIRxnRPMvmP/eMOHacgnZEATgoCgPCtgMZf5p4xW6939n/+PLWtJCelIlj
k3EI2XuZDCkAygzc0yXPRXv+kjBTkz9ufM4k4p9rg9r5/5yKO00SJCED8BJFLvqi
2II5OyATJamSlTc5ZBKlO7Es3FBvoo8J0oiNoJE7kHxPBT/8Zw47tGpXjVa5THiC
NeZotp77TSh9g3k6YPa3/3dh0MF93LFaPhuQcBL/G4un6idClpOGsg2ENRNFmS0W
AV5NJG7llLXYPnc8yiu5UV71X9LFHYmBD6o2eITbzcfUjzFN8tBeyqbNITz2Ynol
lbg+O8I/A6EZ/oMSLpN3S8hXC548lQUlX6SarGXlajKpfrT3PaOT2Rm24tqPmdDL
kjce5J1GAT9Qgc/FotA28I3Y/auWjoNDRuai96jjx31kuyyQuhpJoxxHH6IdieoP
Wh1Y7ksRDyOjmTbKLAI0nQc00HPsA2q79i7Et7cS2it4tc8jAXdkCaLPmwQna1dG
rU7tu9H3BgeQDnQTDECHXg9jzG988kfY0HAFpmEaU+zPUDGUHbXv+QN4ixWemTXM
jmsF8+/ZYrS0QN1Jh1axb3JBa2paIzZmtMmoWR3/Bzkbz0jUkcI5iPqZhvI0zElT
xFG+dPQq/FAx93jgMhOXg7mTYduqGV/iEE+SnOuTFNkLY7VXFyZgQp2LyKDZ+hQu
46fRGbUc7dTVZNQUDConxvgfOWggNOat+YH+Fr/yE3oDfG3MENPzikvcvw+mhLpH
K/oC2plHvb46iYmTFjPzgpP8VqozrWAf2C6me9bfOyYDxHiL918CnlSB6eHXSMk/
sbWl+SyBXoZWsqbVKENisGYVqi/XWRO4iDpqOQtKswc+jw39NSAUfVDGwmGe+kZ0
HfqqcE3tuffoxi7frxMKEOTEwpZZRAZNp2BYTqkcw4yPFNQsY3q5jNoqhOgDRFEL
9ujIq5F2UNT0Njj0cTMfhqahs4IWQdgFdwG1KWDdpE+lgjYqQM1i4cj7VhPMMtuq
4ALhiD+/U4dpijMGHe6x0oE8AjSusjUmL9Pe7i4laHIM48v/4D0DJQgcjA4rAV2M
jtj/620SLcoFSDMt4xOsvc1aIjGP90aKSr4uoqycgGFzXo9tDVkcQ0/o16O/Xpgq
xC7JtbT6aK0qpaDcwhN3y69r8lDGxzb71AvqBOxEGZb4SXj8BuQfbShD+CtrkLXt
s3U9OfkaVT5vucLFeeg1PMfRZa5som4JJ/XNx8A4V+WqVCIhNVsoq0Wj8ZN9aAzq
8n6i650fkjxN/z4wUTiaI19i4TtH0hIdv1IEsNUrE7CYoId1jLz0G56M20DfR2p7
MTcXhHacLTOSDpLPRpphT3w4u6aMQsmXEh6Sx+Fon0ROifx13Z/1IMOhjQDeS+Qq
GFEuNyXCuvRccnydLA5KMn2gAxrREhsaVtCPjE77T9zygKBrKyX+n0xSBCxyEgiq
y0aNFsshFMRg0b4joICd/0BbzJkdFbyUhAdY5lFEtlrdgUolYjwSsUg3HCNC/r7I
NDX0nIIKLvb57M+YpRk2gB4vKifgAwO/w6dYEeLYcZS0IQXiMYIoAo91kMAyj/Z2
U/OX0je+vTLUV//eVFfqOUDIt/Crfq9WheX08FFnD2NL1nivVgVcCuNYhHpTkW5A
TsNFI+pv0aUFer2M1bP5lHjSNSmAycVw2Dak2S/UsaOxg7IGmLrymYzV/veKscWJ
NE/C/4Yiy1LTHrAf++PmrtJhNHr39JifIWohD8vXS/zGzemYel3IJ2I/i+66Sgv/
d6DJTmoeXQb5esUAZiQpZQtJZVKxhM6BEjBZr6Yk/gx+ffwjta9W/shfWua4WB+9
dHc1dvUuoB6g+dybrpUsZr5jh6BQig8IWzvdhnpRrcKWur4YGxw5Q8G4AnZdZAkh
Id2PyNN0iAEz0ddCTWk03Oh6IwhsE2VMdeHyIjBtzeNbi3C4XAGXI4Ed8bVhuAHE
Z9Kf2Sp+BdhPsLAheEX5J5hs5LswfmVQceNWlvu3bBwQygLbFn0z99sdVFmyXpMy
9WLOC3LOEBoLLF2VTudM7iCuD0SqGA0dUPrvdt7F/d7uNhztvfRjaZFJLehEe8/d
QBEe9QrF0gtMYZVnV7rZZC+gSBn7/BBbej+UjoBkuA0/JGC53p9rudquNoodQdRZ
Nb5Bt1LrsjrKB+wIDvA3JeJTiqAfTdPRs+D6QardOTgoHHFx9tBKRDWd8DkvjJN6
Go0gUSX37yv55unEZTTOX8mNn8rho/r+F4SWO+Gzi2ha/YbjKOC91U2paxsftz8w
zwP4vqNeFrxS212PvxYMZZnDoaInSG+73Kk56EaKiDC1OxZOfDNaKqNNMncoZEH6
B/Nbv5TQ5XvJ2bKGKBcgG13gqCYvymfgEVKlPPSMaUBKuibX0GX0CSmyQ76CxBC8
UoO/Y/w6r0S/ctVwhn2uhnsaUjnpekx9KMnui6y2/bTQdNZe3SeTLfBM5WK61HBx
2G4wGNxspUtwc3Ow0E/diqeYA/9mFPQdY0rHux+D4rGLEcyrFnWwM15egL42HgRR
jn538hhiXp8xoLmPWCd5wHk3OSY4wsLsym7RAFVUrHIivsf4wKt1XogvU5BkoX0V
V0refdhyJqAu4Nhfkv/J34coPbwmZpYbEMUiq7sKM9G8aRbQ5fWiVLa8UJ0Kd2Oc
7mqvctf1HHVD6OYaBmiLNcHDQdDP9Clujd4FyeUD7hO/8q9oaA9lEeBiPyePn5DN
HUfPvF5dxBy+EOR4abAktauHKLFuKFJSyupiN8AQxkPS90DRKQlmiT8NS6cIslG4
E4uQNrL6UoAGLQy/mDdH6p9awnhkqxGSTNZUfCdJntXJHND9J/KCdOolhzR3MlrL
Gn6WKhDzDy6Eg91N2PtETQSJk5+kASQ3zGLi6Jy36Z0v/XuWwvm4wG3MfyZ+j0xb
JbN2UzfZmvwbanQvykr8RxvfLGS7ts72TmYAmrEzvwq8ffEVjP/mbcSxSIiOgWui
IAI5Odd8R/tnuE5E8XAzw+XxjPOMmUHsvqa8Eejz7tO3JIRKJfITXpH/GSf4/Q30
DGE77Jl0D6oPJDqBlnD8oMMx//KS7MwWtq4CWXbOFKP4nfw9Wy3AAl3uOiwilmbf
UwBDvp6FY/GUK2UFxdKJdE7mv+HK9tM8YPQFRX+QzeUR6FSAGR2pFd8+bX/U+BOU
NG7BRdVkiGat9qkDj7Os24u9DE5voZ+EgfofHy23GGVyKRQKkftP5+GTX9U9j9Aq
Cw+/hurdV0xyvRyjTPfaXbfyuR+RN2e6Q057TvQXAKx7Y22xTFDc6iECgnhGvCig
ZyFaDZ+i7HuUIzZfIV11E94zD193LEaEKYszTEj6mxtEPfyj4JwPp6i7Y5ahhrDy
jeMsjvrh1gnJ6ZdqtUq/XMlTdogiOwDGppjLOM1AM/ue+gXPYXAVlVP6+hzNmUbr
EQaYywfuCxdJSjTw8WzdpsHrFTAV7B0F/zV0FmbgK10cceGns4H+Q2VylewRYSUN
pskJePdwKjAHg2NreNaGSBh4MF1ttwlBNBUVoUlVZW7c2tC904tyi520ZayfbZhb
a7CjYEEurdXI5TowV9ga/8r5WWIBCOgZdrjeMPhbBO589MYfWQPfQdiuRIPuus0w
lTnWL+Hqzn6XnRu7zTGfgt7CNgASlHEraP2JfX/PjuExjbaBKZ2P2ixgKLqJo93k
xInIt4/RY5ujlHWZD4xMYXQZH/SA3H5wKDXSot3NCHvm0xcv5xQkUPQW/P9YsP4x
PcMTDq0uf6cSEMS9EthhnilWfOJ6F3OyVWYoksiW9wk4Bb8XFuqjrV+95oabgefm
eW/CPH1rtOTeOMTv17+xjwLuA17EjrTSF2dWTA+/b2D5A3OoUH1BGnsFHhYeS2aG
YzzCL2yqElQ7ZN2K9AefmwZMUPqRzJZ+RTuDh/RyAiMi06WMlFdsZpM4SeyZINqA
7W+ndbSTnvN+/MQ7CYjnmbSIg8QMYxpvf2BpFcKmuR3k7a87DAQhD9fUQbkMDZNQ
b841E2AaokrtPF/1Q4cz4Yw6oLNe+LAh/ngTl3mQSvYmbEpHWjJvbtLVpJpkjXqF
PRnuLHqWCLiz7D3EWQfHbHQkUFXuRa3VxSTiBxSY7VsLIvIRHfl9iOzLvaACRKe9
KhvdlKGDtvLelzES+FQ2Vtrx8H9HZ8vVQGTE2Vv4cw+AeI1z4TGa2CxJQYnajWr9
qD5Rg26SzbJsVy3MVm2YFMV+ufvQlDhbVV/j1fWsCXw9Otg2DBJcpizQWJ48jWpV
wtP46pjOnSp6X6IWcy/fhTVC7ExP/l7tXC8c39oGJXHrd4Rtu7wiPRiYziLkcCb0
oK1EK3arm4VWvwZVAe3S8kPaDrV/FD6FqyOdnSUU6DApBxo7b1N+59Tfk73H+IrA
8LPer7cozC/eSEkTdCcmflI1Uarv4aBfmRsc4i1XWTH5K9HvMzErWPRzmN2wMdSM
Rwn/bsNhYwTboNe1Se8wNCessfnp1wj5WeWVTB1z5Rmr5yJSsLFrkg2SJ9NeH1Te
q2hU5Doq6jDrGPjzG/I3nedo9Kjs754XiUnp3zakD0D0HkLoXcSy0MzgrIi15dTq
S4xfGGUlieiehD3XKN9kCatMOkm+wjAsmg/qWrcNUZ8CegFTG4S9TGGLdzhD9H23
H0l3ayWZlKZhedeck7quIbWwE0B+i4hAM8oV/FwAeE/2oT2JE/RX3xyxEAJf3+yE
zqNXH8fMcVoeg9GbvphhnXDq78Cyo1MvxhLtIdBPdsH/cAuwInMX/yRt+s4EQUh2
eqLILwa3tUG/JPEd1glmtK/wimztC/cwKhGRhIRy5OP9TjyMJUy+dGgbNBUAEKZQ
ilrJviudmb0xhrUMAeQ+BpW7z5s+2qOKgQrcxSLWoSftY6T7T2A5IwcJ9O7bonTY
COtB/SgGY333KNAjcfUKoIgF+svHEknjj2yikuLNH0xZtz9L5mQunlGmBDQ7OGUy
lUvE8D19FUBQxEhJNvP1hFpAWk8jDVw/qFgU1/VfBBSzyY/ruhBMp71aNLAy8Am9
S2VrEOT1WkswBtD1UDQdgxQ/ZaSvqGWaJQqFR3PepBbNThknHyBUiDW+U3m9bB4E
UNFRu0kXAtUUVMnAfu08Ks+r4BQ5WUMZX8yuWWM9Dj+qaeSDbxrigp7rb7pbYYN9
xvVyetVmn+j9kyb1kaQX4D5cAg+LAQ1QUBgwB6O4NycraoZ7kfdg3LLXvO20BtlK
7mWXwkB2CssgcQt+m/Z1z+0s3lvCTnb2xcXQzg4hmevHiza/ABnPz/HZdqQPKNDr
u6VWvNyZ2jtLmebgtjs391aP3YvPuQZbhS9msuZ+HfKLha5aEeCAPNdbUSs7Zrb1
A7r6B8GBwwlSDWaEe91WMy39vIZG5HRmk3oy5S8tFK4Uyg31T1lwAgGwgDpOrhGD
QgYJruO6mjHAgVzN+U+IQ8PNMYDrHh8Kn9l/QpyYsoPliRh6tMcIKdttItHicIRf
CaAg9DwZgRRBABN8NgqUHMZRp269XabhF4MYd/xQbzMRc+CDw20tZNKAx0Zjmgo3
nYzyRba2b5I8e6lO1bdhznGGsoH5YZrpPEwMElMgY4csASpu2bLupV2Lu5imrHZs
/KUPAPlBBv650lnYfpVox+9Eg3qIAJCiPFE8KRB7v2CSKhjA8YhwS3pfDXo1Jccu
UJIbgyCcOWacrBCFW87o6nYqPh/fQF5L8I/4r2vEdMgazQhwkvB6ByCUTpnlXqxz
nA+n2yC8JbZknCPgY4r2ktIT3idyEIUDgp4v9NX2dLvmQfOOvWfzF9LmFdYqfNYf
ihh9A7AXc5oFQWlTHWuF+ryJ1vLY/EeKGx6kieIVx1Srx/sfUNiBDiE/N8iSMa6u
qsPMjBlWAAG/F0j8i92SmjxYybn7lpRHNLt8izUwnolSIkMr2o1Jp++4IoMOZrt2
ivIRm7rHJlaxpp7FZ2k20La+09eFGj4ZrG8KxOmflYHOIMFgdMrJk/nm3MoknLAu
Yk9ugPb7xAL9gNSHBm2XV4mk9B1uoz8hnK0/sPNm31OsZpFaA1vaUa3YBtibiKXV
RmEztFgHt+6nVHQSDi4neIKZIXlZkNe83WmrRnGRL9Xhcs8nm4sYEzyiDjuNUrbn
NBdKOpyly6C2v7D51J+2MbcQYtpwJayAVWTD73fcaOfmLhu8lsprrhiTQRrwdJQc
qFqVv+h2bszLEJJAvksZlo/NM54GxbPTyiQB/Yw2HjA+h+HHXAYkGTv0dEzVIJRy
PRRXXkb2aU/oYo3LJu+MIFsRXtPsqjKcB7pwMX7INJRlHojx4YDdEcc8PvfPT3xA
TEhHdB/7CMYBUaWDMaY5SJfKrkoZaTA7zYmwB16UDOCt6jfmMOgqVqnaKyf2OTsC
VVd0Wydw0WrvcDwBumt/xKTt1VuK9te1b6IGMjS/blevqyHaTl2bcSuVs9wvCSRS
Of7JnJr9+zy/oND7PAXRAV7GLlc/eL82T0X+gqLmMKRZWVdl8yijH7UBJFIe7KGi
tNr18m7JZgEnNZaC8J3NbaGJ3DKW4O4Au6JU8bbym+pMEStNPHh9LIjuko6hqL3S
GmpcBR/I2XeS17noftBGKKiEeqx80SSXC/piccMo7dqDpo4ktQdE3hararaqx97n
h/xAZbgnXyzBby6lZuajbMFmSWfqr2DNx6DUouoL33ej9ijup0QjVtLQHsLQ0Xmr
bQOwJc4wlEyASxFkPwgw5TQFqOfKjv+4yV9MeiudhiXqKyn9m8YkQ8dqfNiDRILn
Qbp0hykB6yxNAMD2oSf8YSzDR+Z/vZycvrs9WX516Y3ThR/iLYtRdArXGSoJcScU
6zvwRGFe4r+uMB1bk8/37lLkSnm24hMzL1KE3ddz9t2M2++zY5ZAul7APLu4+Jh/
TbCFmofBtHDh6WdOgeOuXV1qI8H00rjr+bkTKo65CBQG2j9/kU9V64Vgfk4Imzxs
qWSLknkNHfH5sTupy+V6umcxPIbcCnR2MNKj01jKrlYVdlDFGeAWYHk2T2OD11ts
bCIq5C1gDrwF9MGFcYNIYEjjGlXZgnvAybxEcnrrvfNFcw0lQQrqs0F3JY85FMUA
Qyn5bVGWAO08Dfou1XH8n0y9+zsujjBWkI2loioRQJ430r/z4JOFmWGzgLsgPaF5
TJv6qqShXS4lcfISGcxJ2xNUH54oZ45yE6f1QMBPHuwuFZuKV23v3g8fg1kj41iq
YG9/WsAZCC9ndCsB5FQmDeOD0vJNX7vAa49rN5VPLfYeAMSBARmNS0K9kmwfK7C4
QRdDSnJ+t2G2leY/ZcF4u0M0VqBk+5/QxFa/gctr1jM0R8oPiw+DWxFCT41MkBh+
qpHF6k/bKiazzvXt9hFrr6/GOCO12sag3ndKjXxP6pwz9myHaGScypNLh0CDWNWw
m5sHH+BfbylF29rhGQwDu1ic45q/+DH0kDqGjkFnFqPvvYTLyq3guv+tAnX5maFc
z9vuoZsLvenYcW5Zf9/zmRCXTjXmdvxD1Own5WZ8bO0JM+GCmKb1cq5EWbbCoNKn
x/3HU7cqFbe0DOLhaifzdSdKg2htBLgZosO8POEJ+/vAgrUsTe3Si28WXMMMv/v8
fYi5OCC6al5ChlTikX5lDGzvd9HEqA9uo0nANpCccHFbnJJ8wt6sI3NfllaqfFqS
dYByB3+ZIT4GrBraMXA+CGHLCH01sHMBdGOE2u1isNHaTNCOkpfNcvP+S9DUNrLd
quW53KIy58gS+n9Phu5x0wOnX/RB/oSXO0f3nVigL+Gpv5ncauNVqok9OAU9/P4a
vHJwldDJtYfHOAGhyKc+Fo3p80C/ZuUBQYtuKRd3hLmLWwTvv1CyuoR6pGg2Oiuu
9385t2fKiyGG/7bp2hMd3rXAV2L0TJ5rrNZnJKha1vvUedzZvgtdYzWrxZxaVwhD
KSDm4Zb6SQOJAuFD4MfwB8Ll0iq0VxBgI+y3KUAFVVOfUnBZo/xojvVCwn//VLz4
ohp/r5gnMaAYKttnbH9W63Ha4z+nST18bazNZabTzCVeEw4pk4jyFC2dB5S+TYSq
pXvdUsOgUH8VpvfMhZ9amxTFEBJ8nPyFtxxxmxobyoEKYIjnGK0b87Up7h0NejdF
mEJ+u2RizaCD6kEzd51+ACU+l3NSInh5BByex1IKkvX/rPR9NAT8n9lBbz5JOA1M
S5qNr+4fLoFHNOzIFsozhZQgdZbj3TaQXPnYTYHHUARmQ0ScfnFVUuFHJnMHl2Jc
GLFBhitwRGfYvanep0uACu07MRkCTua01Fomln8jHLHOIvd6EInvOd47Vl0iLtFy
IN5sO3Gr4qI8F0saklTrXYlIdG6NjCkXKnXKSIqfcAHYXWH/MVdBP5qQGiwUnvXR
0AI38cWR7zVpqhByKsnpXyec+X5mPPfDxDS5X9cwcCBGPCCWm+2glSxAiaHwXoV2
CcGD0ewVZx9pC2GQO3I/4aXauNBsW4m4uBbf90vtOCSr9c0s22ggNtfDjN2/N+Xv
MYLOtx1IA6X3vV0z1x31RhdY6vY/OH8Kdj8uteJNm0ZghpsPTwUxXgJpfRy4LkK0
Vk5AqOysFd/q27eotGTFbGS7jY/LqiQF/QjWbhZCY2eVCGn5c2cad5sm1Xej6y2r
kCCRplvtDdQ8E/e/r1XyEDYVp4Zzs7S1l6jZVqXNmRRip4i+BAssLEQPLICSGlnV
9sk2Vz1LEI1MvHqGf6bq36mIenLnL5PoO+fIZGjh+I9g6hUIKir1u7DDA4tsuS7v
zeOYjo1RgKHj+tBJf0wtAvKJp3v/fDRjIeXWuWzvsE7iR1qmSnEP21prhTxxylMN
Wv3g/oV2TrRcqWQ0ezUZkF40+XqI//cFWMxy4hOB7yNH1QRlheR3XkX7/ZCFDUJM
Pt76rCLSJIFHNeXSpJbN9r/PDi/3l60cNQvNvs4uqEzQnQ+6aP91ha4eCCVCAzV3
Nwjf3y6HieN50xEEe2cy24pLuj0MCeHLg05NTHH1jOIM87vIpUrkdy88ytIA6pRJ
tWRqtme9iv2r6t0EBLVw7se4pt0ZidYXoEFhPAsDMWd+1hySHxbOy6SwxKK2fdZf
h6Px1JHhw/NKc1Mp5D1jC2Bu3h+Gkf2XFYccxVZIqGI5dpS4DFJ5hHisOM1Z8fSF
7ULLKuwefHiEDhT5fa8DjvVsDXdp1OGxLyXV8HptAGFk9MZ3eyNZBLnAtX83OL6u
Rdn8/gx7KC5LOg489s6msMEQMgn9RqVRBUkF3nfaELZ2+tacXtQz5PxxY9Pe+t3M
KCOcuea8Vlpa75MFdfjYn0O2pXJ+Lrq4H4YJs+rwbQYpOtEpacyu9ziJGUasLno/
LTClkymlTf+Zy0paDXRUCU6ZEBdObwPYrHZOj/a5UNXcZUBnLQ3Zmgv77icbIU1P
evpM7SqwhoX0iK3wM1TKI5NvmGmCYT0aNQqffRPbjI1oTdRHGgx8YB8cfPNzZqPa
8YEszDCgoXAYsowPcQj3SZfox48Mn36M7vcTcWp+iDAYt+RyW7GNISD49l3IsT6n
fOcZIChVDLj2aI2SwpwuV3kAvtnu5pjyIqFVsk0PqhmhM1nXiwWl7XVCMejoK5z2
9ijBHeSz3GPTdcNerjO+iwZubDB28l1Smvp5Z/Rf4CqU142yB9kBOAMqodUL7W+v
paHQbtpsufWe6HRgXAPR7FWnr8/GpmwyFu5LcEJ9+3OLuCwUVy2DYFl1GC4umeTU
PJX6kDJ8m52E3hsPE7VHOhfLaSyRp8MHWkubEcFggsgc0dXE+cpknVLjOvYsr3t3
+1wQ1jrZBGShPIgdgq9GmxeOX2hnLbbq4F0/V9ZLCWkEAGuiZAgx42PZG880Aq2D
orxFDCwoPrQ5oo9sQJMcGdlBAW7O19YujXbOgYaij74UM2FyCqlRPhC4sssYUj53
qzfWZWNpvJpxIBwZ5bKR88W4UEzKRp0jxd3pVm+eBvHesL2mF+dgvwAQRLK4Gr7d
UCZKl+KcqVF5RQEJqxY26onvCYssp4xCvJrqv8iKGjODUPmBB9QTZeFFwUqq0KDp
YcPFz6POOMV+W3AFOZb+vqnjb/n31KZCzM5LKuvy7ZCJGQq/8apl7P+MxhjEFPKB
qcShv4gMv5nLX4WLvJD0q4VBO3TrgObWdD+k5Jw7gaW4xJXpeOtQng/kmkw4p8r8
tSLlb07fHLNXCI/IZf69Ot0R3jw/Fk98S/UeBtAl5H6hvncoPMqZRX0dWwyHKUUr
cI4z/1sP9BROkdlCZa0bKHRuAdkAYlYKoM058PkeSmDagOlOMTl3EqLdf8n8VugU
UsZXDpWf4MvHxe5b6IdyD/S1ZWpCzlJkFP1uPVQi2n50UlLUOB/k9bZv0ek6+dFk
pwRWPeXK4jvewqXkRdrorXdAvTHsje+IiK+Z6MiDqm1UAFIDZlNN9lZi1YDxPfZw
nLmjywT1PTtiOCyJL7DVvRTv5nsb9NzIHXhiGqN01FV/9wVDgvzC6hPSwI1Z26b7
5mtagW5nOwafHs87Z8B9Ls+vsm2Ob78AsnlLOWITXlNahEBwuoIsdoPTr3MwPYXO
8Zobn8Px2RTVJWLw9PQLv/5qJE9N0HNCNp+famelm8C4AaB8bD32h0IOERSwIAkV
xmmOxXnOkiheNU8NW9VTkT19ktuplGAw7S9O7VV7i+BhiGHtnw8fcfYG8K0CvosZ
Ua3l7q7JTk0IO6AHPxlKtths50ZRnjNZBa+150KmkblR5kfJEKLaf5unUrYVLo1T
zXw83Llj3suZs6z7gvh+qWn3u57SLnlzTWyXCuXUaQGsLg6JuS/XCEvEzg6GCNPj
l7o7Vhs8AK12NbBEmFR0vjkZE/zS4LD2dHYlyrheOToLl9ga+BL0iYRr+qGpm6Ky
GoCdZFgcUN0qhUqEQXMnmIKjL5EEHeJLH/dQqMuVuR9NWR6RtPvuy8BEwAEhZX27
A19Gvh5IpHJKuHYiGz5O3tRp6yweKeN+yTLBSMnosxyb8CqhZNOwLgLzMRCS3mDA
P7Ju6NRYoYvX1uoQLQvPSF2omL3BYo1lk8UZtmP+u6WJ8wI+OQC/305AspDj/JXh
a1EEba0LzojWrNJ4dwUMfPVbx8EcDxC+q+hw+I+PdMGYRd7ViM0fJ3Jczgk4aF7V
NreeFthUrv+qemM9HCccgylleU8sMm8hcWWDblqgIQ0wo+xY2IRueo6nNZpiHnac
I6NRIzB86nWrXhVTOisY2QMKJ8stXYAa3cgZb7kAP6Njy2Ve6ryzBDMp+Lq8S5LL
eSECIW6qBcX7dgH/Qdv2cI5wjo5atHEYkzneNDrUtEHp1HNsLUzwgUAx64Ka2J29
/6AW+RQFS3hc6fwh7DqcPnZr4qVjg2EN7MqM9z5UPYzDvyqV9fTNhA1iVCUidKmN
uTsfzmI8rEX3/RnGu3OuaA0RhqtNrSGIsz2gswexDkQF6p98SQNqe1c6gvjJ+J9z
eDm97ebCfIMNqJZYNLyoiOGtqTNif4pbf6GyZQ/C6kj44n1LNUYWiyVKM0UgVzqG
O3Dh5VArNPd+WquhJdGCcDn+u4lDsCBErh7ys1l9LJwssoHBlgF6b0FYAAWsYJ/B
sJP1osSQ2aGtn0K4ZK65xEBJh3XG3bw1EGbDCg6tYsfD2HJgTIasSv2lUiSFPNyP
EbzmleJKy+DaVA57KKEmwjO/0WC/8qtKry9OeCXZMraOjaMvU2fDGc5S9PoNvFWs
X0SJbop0fmuKukQAZcf847OCiQ7WuPHXt3B9+6LvVDC6FeRqScuPvA21TwRvG0U8
mCR1ffEYF3qo6XjK//FT7HcU+zorzVG+XYrAfLlU6pV5/DPECijws8uYGuDo67ix
sF3ju08VqIcaWTgv3Mhpd3VkqdYI/SzvnohzHjdNhmLg7BtQ2Rqr9mUDBDxNT6v7
jNOyHN/hNzqcCCzakrm7yBbrBYyvX7/oTqcFg0uhSSNeUY1NGAVK/L7yGsdAiZvx
Z6I1IXhGy8SifThbvRz3VYLWnAp8Nxv7FCx5YIELxDAd+8zY8iHBQxpzRNAh85Ke
NAIn2sXg2PoBymjMqY8mhFy6i5SMxxrY0rkKrXkSsH0m3reRCDhmF/wVnwTD+hgT
aYUm70de3I9kGcAfdpgf2iPT8cwwO4K67FTthc9eD7IeKIlceImhti5dcFKMjdSW
0bh6GoMgHprbUw/31B9U9wXJs+6dFQyp3+1JvA48NhyfulEcYBrq6Hth+72a7QWd
xvr1w71PNY885tVu58YISkFUBX3jYV0BPirluT18/plp8gWBlDD0R9/2IEc0k3T+
GvZ/FXaKukDDyjwL709XhI7a5pQy37SwOPU00yZE6pJpoqQ6gdx2uH8XyCRlfZaw
l8I3LmaSkiI4gv+h7k37rXeWY3QtzftmvjTPv5bDYd7NZ8Q8s2uH+U3MJ131LsOx
yrwKP3xPnbMWEnArOf088LND03Ike0tappzz6rD9khefKtYRvkBvNVBWnVuN5R2A
wzw3G9+DMaFXsB9fdqhPcoITUrVH1l9hFX+VOtQZdSD2Y+fTNVED5mfmFebvdePu
bz5WVnkNg1UUDEQUj4Egf4s+GReDAVe5tFi6OYrX0OZw3+MVQFeGjFGchoqBJ/v6
J2x9yDCfaboT13kVb5k10gmhp1mOBNP8NhQMWZpHRYMoH2REtA1vUINrqIzvz1iM
kAWmmg4kh4nykMdfPpc0QRo3Gk7kvq1r9SMTEdOEtvE7andwcctAWaptDUv87Ydm
nvpcz7/bANNV4G0WWefekFAuInBtn9XL0RvcVTYoDNFwgDnSwI9T7N/N8iWIp1yL
o5AFhfQge7N7p6TPfwlG8Kr0cbKX9s+SC7X/YLNx1V+xSIvN8y6/2B8VZPT/KCBf
zsAkT2VSl/YGXQFjsjQcNBc6YwM+ClxFNPKWqV8MAkJdSi/1f/8NGgkZTEGqVrml
cz/qVW3OkfzBwE5SauSoNIIbt6wPQW9vLyHbNEKjVhAnFWar4DSaB02iFz79BrXC
6ouomtcIQ8dqNg9llnXd2UBEdM0AYoEVUhnZf+CCDhCz0WUj6M7qXVvVAN6G9VWK
fooBjNw1xsp/l8x/r/6NPrHJWvLlbu25HxX8bBi1RzHReH1983RBu2cPG5xYDLwV
ZQY5Ip4PCtyC1tTV4hedw4R11nSI63tAsEKvddawiup6bv6D0Bdj0vv0IW3HoPJl
5C3FUnu4Ra2cAfuX6iTQTLXX53BZSOviXDRyGIvCQ9YqNbxix8UE+9NsfB6w3dcU
qXTq/FZy+HhxlG/qtRLIoZY+H4zCk59wMqtBXDjKT2NgT/OUMyNdmdeTx4g5JtYI
3A6MG+wWbAZnhINVChtFXag+ewN/ts13gjjWjaGB9c4wmIC06YpFungXhrXnZ8SG
s4LR3rJKrakFoyc4rXXB/wtUAfhp5vOo8nMRrCXO9QapJ+w/5V6Sf+a0M0pvoxfT
BRevfsLa6oCHNjBK8TcPSL3j4U2EC0iF4lltjFCH1jZwWOJ/PQO6i4fIoUsa/7XY
j7eqMsqQj+HlpmETgkFoLdN7wZqAAFE5y6mB9nD8Fpnn4JYocJT97lCo7h50abdG
lpu7pVdFC6q4/G99lwV3cY6+M/GAR1U4karCqAmXMysZJLElO85uJhhx22kkXcva
kpsWFTOYLxOfFUx9PsSAadI94lR8uXSGjQ0RljmIVmyX4s3T1gAJRDRbU5dacpaa
gmCNODQTBBZIDJxqU5rxrRMQMWc+wBqug5N6YrAiZT/w+8zjPPVuyZW3cyi4/LdX
TJrPBbvjpeFly6/bl7GMCd0j7KVf0kk35B5Ca3tcL1BjlMdAwf45bVOl7gRYr/ia
c8QEKGG5dfSA6tCZsQdifOXiC79LDO09JIUcvzD5SdbEpFcbKUz7EKdXjATYo46C
aE8lEecZ5HSx+NFpxtKQkVqJRYArkcn6ZDUELA0R7MxIGPBaTzYeI2LH+M4KBzvk
i2aO7XgcAq/tHiOqMPVDJJIaoCbHM7Lxc0Gk5X6ZqhspRKA/ZxfIgoEZ5oFyTnvn
IzCRjy1jv4xa4LtvIHAHA5oMxF9SbU9JX/huMuQ7bgF4ei0GWvyDHSfds2e7QAP5
YtfP6k3ovv5c+GGxt89B8s4xE9vXlrqDh0bPbHtVrTGQYGEzd+RILLTge74W6CYp
xaFZooAvUEcmZ/CBUtva0fcRS3oddoM7WI6FwINPB3CJ+iR+1Y8oqCeJz3IboiEZ
DfYpOIlxU70ymdVpee7dDg7TMwJZWFch4HR8asvKR71S8E7ixFHrTZjJcOlSl/qY
UFMwC7aGSASN+vgryOlvbRbE9FKPIqk5INgsTzx+irVbg1MRVGEJqbvrt+/Ud7fK
HkWWDnq510yGfCBFpUSnpnjXpqiza/886DF5t1D+IjRR+kLyJ+aPHUWu0QAsBeMd
EDDGR41JZVFqXvF8CeFv2KDOG2LUFMsZo1EMxY0qpdMdSe8hSFnsvWjYOxhHMiqT
B2ooIW24258hyPxwH9g6f18dcpFyh0tWPE6QF7AsuH7SKQ/AY4qGIHHogXfBXwrK
qSyHlr4/OlfhuVDUYf7XZXWujT90Nf3iZHUZ7Ji2HLAnjpq3GFNUAsVtjbje6x5P
G9QNKVFPfxoXQKZnGjdVCqlISUk31vY1bC35ZScxKWHEGmquQEhl/E+1Ww33CLJQ
Tuqdrx71URldA34mM7ut/nKdAcXWEUV7S2JJhJDAyGNyz5/ZCGuzJ0V/BnqDmyuE
beNyAtD03VBQAFHCUVLVYULei3+jcZOUhQrO0uvNtWPY8b4xoeKOq6wzKCaCZYdk
DiJvjL3m3SJTCjeoGr9PYsQVN4sPwP/pVj7cwHJakN2x1H87T6C6/xZn5xtGeiKk
sowg5aWhh+HiYmDMAyNNKz762tRI8HcETKzkwCAAq7ZKE589RyReZTvMqrclVrN9
uptKJiUQZSq7mEkCFiOPd7BZmcA1E1o5+mVyU2+lN1Uwm+DjRdp6A8gcSPWCj45J
g8/VCjCefqXHHJOl9AdvYwPp94dHFEzK26JY41JMYcr2h48SAGygP/lcD9TmaaWA
BgJuFFGApFzYtyohGLXbzmbQRW9cP7bxQAvV/9rjyFQuGL5MfwIaLrDMA7lZia8t
a3P+peoz1Z/0zbXNQ5xGCPWFBJAtdOMjaKMgEictR1GREjZZyv0ZAYDqBlvwxzb+
g0W7Bi/Hi5TfoUHlCgAmbjedTP/xHXiP9QCu987z+WGEmh1PpD+9NtProM3cqA1L
QMZyUjNmnswm3MyjcgyceS61b1e1FgJ3WvCEN17fqhhxrU6xH8zy3+jJOw7BkJqU
Ofsxt8VP9moQmf4rSQ281Xeu4KWOeOuHFz14VUZLu1tPTCzdTingaYOLYNA0o4ku
kaiVUtlM+PHuJpdzzY2rKQ1YcKxh8NLbIQg7Ii4xuwmi56YdKX6DMo9mAARJgLNJ
S4YFietqD6WkmiaGAU8gLZBoXuxZ0X0N9DE7dg/60lB0wwt1tDCc1ieJ79w+/Aok
MRSJESoDyiEP/1AS66amuhlsbbFmfekE1kAUha3m7zJJ78rNQesZnxJRvJ6X4FPP
4vUTmu0bWsu9YXfN+gzTu6/RBtWKB42NaWG/sUYRdSEXdeaqtnSlVrk8k7bzrRVR
vrFCutDyAvz0+WN7yzmzvdgouPYjIXRiGrepp1dM2UTvUabE6HOlbylLo6Z17JKQ
tKBhlxNp/6SCP2J6cYiXfv1vWm8WqoJBsrRR6ocQdGlCzwJy69pU/WPnJuqD05NW
VPJpwyb14267rI//nkGyZKMMUTKkYZG1gesrZ7/17So2/yGJN6W/EWyHdCaqaCKw
8PPaM2ajpAXkNtBhF1yvxKB5KUQjnjBTd2XOQn+3VdNqiLCZN7Za0+lOEIaHt/5M
zwHuBbqbEsLbR00k0Pt58X3hKp1tdUv2Ol1f0FZp8aw5ykGrUNRug3N896FeGNg6
ktdwoil8TZYwr+cWs6z0HwO0bEXBaj6OHW4bD30m/EJZ7aHdTv2QQXKummCLBr+6
03ZTAVZ96at130g1XouhCpNyv7UOfXrm/SETmbPb65fqa/N/QyVSjjI5zSWidhlC
v80Nqb6asazfsEuQaY4UbHOKMbOjp0rUDTs4V38LSVp3DbjbD0wpYd9oNR9tja6S
omxyvYTJbgJ5+Pnc3ACgYY+1iZ/OXSzIRkEjpKVG1dEJ49HNLZbXIfOkniR7OxEU
x8+PRRk6f92JCJ+O4Qfk6NZmnx/mktOMVAveiBLdhaQ70id/q59gRypDTikbtgNq
KivUnEzpdXdElnqGMd10pe6TzBwco+XDrDl/eT86WEH0EhBKlbMLrJD1inG+fX88
dbxyFvJeqSsohOg8dOC/GwLKbNQFPo0tufaLlpjDIvg4Bv4kwbM6KUWDxfTNqyXo
hkhDxWB2+GKFz3Koo1lkZIcCvG0vjc4TL0B0BPr3GcDB0Rf12d/gtSAwNXOudktV
syhWgPHTdXS2+XI8y1Dlfu8JaKoEcOIfyG/JRmyU79hMQ+BJ9NezRBWziFXMtCMn
gP+8qL+5OxsmLiuUTZqluARqj9CL6UOV2cUykC1Bq8wKyQPi+KxK+gzEy4ffYoNV
RcpxQeOV+iAzHOT7O0nQvmVWcg+hKsIr/TsaGI4oEtc3y+abatuN6Lo2KtDCbyZZ
cM+GLgrlDopxZsCE1T36TBQMwHDJFjrcR30yAhLeTervabn/h1Z1ahAC2kOFrt3Q
9Qe3dq3xRs3AnLmE3k8C0mmHsyW/8YfztlK5/wMqQ8rfUDg+NumeNFar+/ph+zso
EuByd1Y1F4pZ8t7mEdFOvOR4faIzgpiS69PijX9ZlDtW9xuGqba8SbXc/XvbINFA
w1d9I52pBxeahf4CrdKhCGLvT1VTEQi+Jb87SxJ/gyNg7PTtc4YAX43bYotqLJm5
biLD3mWBeoy+j++4CkOew56tU1xRxD+rwWYR9WrniDFx6GszqdUpE1EA+c0EjQk6
6G4lIq1AgvzLF9o0UGBsRaoZEG1IuM8h//tXU24yWrh+3w1KITgwDqEV5FnXljVG
gDkyMc3Zj7Y9L9M7b2dLPjB6rJ4v/rE0w7xjzVtOVDcwcvKG+tEIlyfHqdkA0MpE
hqFGhJP2h3Qj/AYSyzfvstGk2fNs7lrPI2oj1AU4J+a1/IOdXtab0kdjzK0ZVMxA
xEbVWvxbXnLZirMoAQs1okE/0RRuxD4A6LNdRrmAjehhbRMmle3d1gxegDRpYzGq
J0tBXhoMVR97fi78O0u6fnpgEOyytzQ/lSpL6nQRkwr2v5hbf/FSRx+lp2OFuWQz
Hxqx54F2rolTMZqah3vT5qILfTIFyYuPkW0lVpj5MhoigkaW8a1/9crQjgHHPoiW
ueDceNC72LfUitqeQCIps/KeuhvWUJcTuSnL5YStReOq3ECQhL+LctY7X4Gak779
QW0yahaEFNAYEDz8b2cAE2PZIr2dFItlAVTa4PsH1ukXXBSIu0Mm+H5OS+bABPPY
ap6WDdq8gcF2M7YOwUnLU+Ykfa4OyO6Xeqa7eu1rsZx7MEyAKNMakkn9ZB5jl4HZ
RgTk9GeWlMnX4LJsokCVw3WGt3lzUfp5UkZW+iiweRrkndH+4WirCZjagfobNU9a
cxQn9ypUAe2a5MIt2ZsjYh3uZzjCQyQhyTmuWz6dE/4vhaVcZJiLIH4Fo2OirstZ
ibAE5hY8c5vZSP4+vyk6m44d4DLzn0tc448fRa4FFI9vMNyfV704GHhTn3/Hj8vN
8CeUtLtxZYbi+PU9dsP53Vm6htmVOicdfmF4X5ldt3SJguud05lnJMAHF74vmcMi
g9ckJJ0PXHbQuC+sF+qH9P+5bN7r5T+zJuEN95G90u8KxMkAQk0Ia+IC4X5U2XYN
hIzGhe58mWKrzyjz+VeU4oRxtw6uHKjCBL7dzpjwBtoyKGcGIATT4Iezaf1NQXXr
0926doxI4jyZMvmQwodkM2JxNmI1RdVmCozSI8Ul4sJZg6PSH117e5X9Kl4YQbNv
0YuQwiPvoOuqwhMhjuqQ1rEGQfUMiAVml+lYbFul6YNiNP14z1PlQ8Q9Ws7/GH0T
vrYn3gNveEcC6n9DqEXnTUzf5nZCclaoI8KVg6pMdYD7kCXcrf5KS9C92n8yMysi
X1tDNQ4Fy6TeyMqTBc+yRp62ZnyDJfUG+MdQmXOU8env+0XZuQsPrryJ/qgKaJU8
2d+o0SKG9JT8MIIJJA3b0hr0j5TMqrxBEW7aj9iQ2XFvHCjLDCSa/XK6cQ+DzBis
8KLPvs5Uy+NeIFiXqeaRnHD+HOQUvGQ0fhqbrnbTTgsHh77ukNwMf6DbYs1SGX5l
k04YZh2J16GDH7+/oRc9Oto7iOMzrx5gZGzjCEUWxHTbfmeg3qELI7aMQ+1d5lK1
7RH3P3fxFTnVg/vBfgeCVylhAoiez3Z0TiX57n7NWIzZrrBLStW9g/3lIKvie7EO
eRibMkOW1eJlDsJ2T+Go4KJnJ8Q+EminHZFY1XY//Qnv5M3jZP3sNF19JKymM+hW
DRaH7AouDp+o5mVkibRpUwXBdZeIiZwRqXhgBdj82TgDc43v8d3+kjTroiwZW/Hf
jzl1e7rTARxWz1UAAKHO1MirPuj+TVUfEbUBVx4Gs7qqADxeBEQVyaai0HfHMQNo
2pJU0Sw/x2L0w35C4CfXYvyxTVZ/f4hHVrCpRhhcK4y1C/1/QKtSsiTvPhrkOhJ2
R6qbKPW7LWViFG7R4jIq1V9NDvmmhP1/Wher0XwsWhbFxsrJnFfiDUtSqmtmKVlA
JJvJVcy7mIWe7RjSMsLOTvj0nGDrufIJUx78JQcVc0nZ1KiGPv97z+lIEwi195WS
rCQlEsejL3MdFbvrZUj12uhTk6D6X/Qtbp26zNcpKSYe3+YtzA3vgkS+YB0zS/0i
oRxmaWmiyjaNRahjf+g8VSkkJRUFTCPmgnGcYlAyOPL4NYL69cD7ao5r1RAqhen5
geiHqCWxEcB+VI55vAI8fR5qFsQW+IhaEH5GhLmY55kgn0HF9xzfTG9E0Kr0ZfVL
QNXENrKbVgCsKmnQzfP7vxY9iRpgNvyWS/eFV9ZZTL+cOhcK5OyDSfb80hx1smNG
oV4tTvVLRPd2PDmyfGPzPwFTlcuknIkOM50asx6BbbAaxnmnV8YESFQL3gJ5bqXf
gaojEpIl1qpNZOJtnVpdH18qESHO+xdp4aggEci4sEV7yCTb9iIrbMxrTCuwmVBJ
8hZOG95viS0keAxVZZ1jFYYmjq1DVOb9ufuW6+r98CvOjNZanpWvHD/hKYQ9bchG
gFHn70h5i7Vw7tCj1OjwNqSjNfYX11XL8p9r/AqlEyo6HEGno4VveoRBjdUks41x
bXqBBaRzzJASIOFNijAKNvpjr+oKLAqKzyWqeXSxjOmTfkZ0gQ8pK0WCVb47n/6E
oAdEqlQMWDfxEQAYMKL7iMDwMOet9V5QgxBD/sbThkTM5bzKZeUVSlQSkgSqeU6X
Tqq8dTnZlEbC/PPdcFCp0CTTUX11Kz00di4sFqplhiirktIT5RQNOkMYxOB04/KF
KocZbvn6jbwobp/xGGaftfyr6k+PSuAF0MSLnzDH2N/gmpYL6EVcnQw+7hjrNeru
iZGmISv5hyMya4AgpwqqrsKs+4ehXZtxCrZkYeTrWJm18KxbeB1S7TYfZaZBqtvp
0KOMz1QFT/9s2XSN+860haFRWO3aI4kc1qPI6YEy/Pevk8RroUpkJBQzGufNHC5l
un9yMtd8sEekOaWZuYBEeVYv1/JZ4vF3VzvzxRMY+WDRUwc9olELKq72GOVscHo3
JsLVgvgJdML1pKjBxWRxQxDFkI1BywzXEa/5O9q6c5P5cmO5ghHvVEOmjlmHFfsh
gJRXvWUhDG10RSNUk8+lUtERajm/cu3lvce6SXASRDrHs4Twb67l6z5M+QHs+0zD
irvE+tTp8xR9JVS3jmXCl1xbzvbX1UiGzRmiHjT51JYFAhE5sTAQk2Knxdg02/I2
WftZO7K/+iNvFpekd1Gr7LljE15fFViPUJafhRUVqvCk6H0iam8/aZKUXDRjj/wd
SjV1HrP8lPtBnYrp9nMkY6mjgjlJJUfZt5QtjsWhKnZMjk9Tzsp/cRO7L/E914xB
1GNea2Vvn/7mZ0Wxyo/fr1wW+Oo4XLpfjzqR6R9U6qBBFQcdWkCXbtN1RPR4yoG/
zSvK8IMYHD/mPoQPhn/DZxOS8eqmEOTPTjMucqclG+APbLZg9F8H4Eh6w//V3ets
DuR/QzxT3dHrLk591ta7dppEMyDZ0v8vCUXeBaLG2VxxZl4sO+KOfUDHtwj8RqRv
v9oNB3mELAOy/tgpbqJq1QoTYzkmelq2Q2HPJ9eVZ58AIMt9sFJ5lXAh+SHHcssH
Dml4ddzUe8gk2UOmfOJEdx+4gfnTvlDDwQ5SJXdGRmejSxnEARFrB8L9ms/noM1+
ukKIEyz01QxZPZoVaQhUnRmvD2Nr+4TN0VB086+GlfCK+To/pMHwkWIaVOWtAc+X
figLWMdY8JvUOmBC4YOZk4iP9LkNY3YFZoySdEVCXowgAQD/KDaReMqjd49yV/ph
Jc2oqYd7anPE9y0lotrjrvBlKdB3Oj3SQhT78RRp1ldEoiZFZclOjW1mYItH5Jaz
CiFlYJYVO9BAllW93aDrMVDxhxV8QmoSFLuwAgUl8fmYGkrIGK7vA1lCY9yoeZcy
KVJTcJ9gi2KKOGZttQbDMDSniO16re61Di+ykOHts5DNWUIAAJ83Y9J2oeFRcg2z
EuKuygEkEzO7gwxOvCmv6aBLbPm41brhAWmlgy0A7XpwDSwf4PuuHoS3S8EneMTK
wgsHBwHZFCd0OuB/1zFbciwayTMgrTbvvPSh//UHlBUc1n4ln5CiNyf6Yeiyug27
K5vLLLRPazlHZKZJqYw6GsYHbhY4Mrf3lxY3Ax7eeTK7y5+oJtP8KP3ZvvfVeOaI
G8zogglt+4wF3X0Ht2vsmI5gAl8JvKWnfPUzGd6VbJ5yJMiIjlTNf9WgVE1xN31J
uouYKxxCnKFJBZxEXap9Tsn5KXSbJeaYe/F2QfB45UvaGUi3Wv3aH3TjckmxJc48
raoH+X07/E2g5aeEN8n5P+BHQxj8mR5xPdtn1fwUo/QRauR+Td+TkMOT9/sPkinL
WfuOpGRvVBT+Ct78ZuPzanxL2vq04Ln8KawiqGv++AY0Tq0HfXJ7eFcyF3hEvbNe
gk60ZPTQST61q9d8QaPdiz90VMifATHPG7nJ/MDQQ7T0ZD9MduettvlqIjYbzaae
VEKirXL9K5UyBlLmWlN1ritxjXw6bSTnodbCnaW/g/ijvmbUbW2vWGaR7T/5Mdil
mHSG4NTa7AXkOSojkEXpzp5l8E1fr+QF3FR3LyXGiYjIkSTD9nCC3pBt5mzghviq
CMG2untAvtPa0Xfkj6nWEJ8LZHUxGT/B9Kxbmg+9diSHVcgd7CvtO13CPJ/sPkpI
pdxttRo5jO0XmuStC+k95hPHMx9iqjbWfDIIKiiT0LSa8hj8s+x9Yz5Xg/MKjxZi
xavBoT0xOJ845bgjGYsAshz7Wi4OPTgjcwX3aB5ymV5zo9PFNybTa/Ouv/4opiBh
/xBYzAgbjLTez46hyMm1Viy/N+Q4o4dWXNhK0O93kHswMfa1r93G+B3avgrD4P6y
WapMOCxjIHU15nY9RVl+4BKQsw+37PR0FKPyWy7GS71AZdCWfOAK2N5m0Z+W5jIq
sfHdk/Strg6qLfQ3gPtFIoiBXSLSOnB1itamCkHC4HTvlob0lO7TzBYxJTv64Bwb
wdVCqx+tfxom3ri95p8JOqY0agkjmaaNPVygJt6uwgFqTMV09pgOKh8epCu/c3UP
BhXe7Kha4DBWXL72DFKKSEYc9OZQI1nGdNQuYuFgq/MDPJm7owRqGY55+gYmDmzw
rlUIETktq8xIWSifPDnBYKlCVwr+INzYTldA3uzfc38U3cUy45cYZV/QTB+Gw9uR
3hZeBaRhSRKQLL3BD62jfnAeNhCwExHvetANm9VoZbLRAzg8SQBbfy8gjejNTIgt
o5yr9SY0eL7iwdLlXPAiAF9KzlwyhEKQ5HZXcPt9R4rg5bpQ56NQD+R3JO2MBfGE
DzZYNZ2tO3Xibra7d4/RF+FyNHV7E0wY0A+lBKhKXrcf9bdmCzWjzget0IVb+Yqm
PeaDme/bmnsE0F2QgQGv5OR8edDls0gu8mRIS+nUpTpFJfw1VQ2YtO+6Zm6xjcyv
ta/Cj3noIXiNpcy7A1MKWB96rmIydWI+SYnW12sycNYfXkvktHq5EwYNiRW/DupM
FhyHKZ7bsy/MLglUwCZhN7RpESZYOfCH4NPFW30LXazeeqbShMI/tOoa1rkJVI9X
DAby8hgmU2PZLlHoJ62TCKy/PJaYLQe4iavPvRGvYL8lQdMGzH8uAnHjPkXBPhjO
SqCmmCn1AcqITAfnEMltnHlkp6HHApXQEjLEfvgaGrB9eWN78/ZIvfvA8I0cy6ai
pfYnZpFjjnwk427MlOVjBElAwwm3YjXcCzjkOGBj2bP+sFq0ED1kFwRGHm0ciTzB
d2qMMYKVA9b3BBO4XhZ37CN2LM0Qq6OczK63kwxaWRa+X34zJiPsTDLbaXQzkK4w
k4KUQ0Mm817x0lvLwfuPenT3HnfIXU5oVog+xW0Xxcm/y6/O5Jb6EwOjrqDL+hR0
HnsiaWowDllY0orkAHWIepeiWNUThRSMyEFTtpHu7IN5KrNTUNGGX1ipY9IMgoF7
XXP+v7yM5e9SbnoXk1TVF6iteKZ8gRRupRTYE9EGCqvVZmMjFsuhtMKTYi5N8RAW
sFkjBLcYUTve0oleaFEEnTjREqR+9Nk/M70nMKKJqjw5U0UQnLXAfJAFSiBN6J2x
yoeE0uJgOFQ3ZA+26IWhe+WpMiH5tPWN5mIVoA6ncatOWrXgFxbca4EKMIpFZVQW
32qtYbzeMLEwxKA5m89ZSu4Cz0/Ag6DY3bJIgdpXCHxdYMKEB0LKhoDYMcIjUqJi
82GDk8M0imWNbCRiVe3MQMEfdubK7TalMVyuj/fzAZvqqQu9v8mnrM2UZMTpSZ+a
13FwBvdfgMQLAN1kFZ+4BEVUY6Dy6kWwAQBz6LkINcpRdoPMsE1VFikfD4+tc2t2
PCjjvW7MU5r2F1x4YS2IC7depj2/ZhmD2aqEb6yLHHJT6a/sxakYPMLOGJEZMOdq
ERnx8kjuDP4kFkLdZxqTE9N/WIAbMtaG+cJYStXTeaPv9Wl7pJ3IMPCI+K2A7qoA
l9uj/krtWSHPyH0dlGT79grzWkwBqC2+45VQz21tVXXioAyrSiOTefjD4F7pmIQv
2ouHGekx0M+8A+RolBsDKPIbnPFy429/DSppBDrME/IvVhEGh7vhxa3aPr8Qs03W
AIwTti7m4d9GOZJrBy9GSZ0iePemo0i2NkI4Tavf4xqh7lW/2S0LvJYcXcFbulSa
4O50hD3daxqgK3Vf4HYMUhm8jGQi8wwEG80P/6RzpU85IurhsKSAuCftorIjRhpP
ijK5FTOOwCCEalZKH/C7nboSLEMNJukAuHDkdFs71L4m64Y7cWaykqrweDfYzhn4
R09iKB7jn5bUWTBueNAxOSp24A4Fgm/tFPGZZVF5Qfi/KrxwB9U+N/vX1vQr8V5S
DpPpAovEAbolaQY2QOxCWl4S7kg7UQMD0Y8XKtGbwrYRHCuo7cNJ1UbiXSSwBDsr
sU24t+GC+42LSLKLHkZ/Ro8w2spmzmKkW5am2LlanCeVPjgKlq1BEdYbi19/WRVH
BF0Sa2x3PopxTU4/dcx0xV/uRBtrFLnXOaAwxUOxRmHSb0hr+HVhpm/iMYii5Ai4
+NTggNQOV+beeivIOWqGPeIZIhtiDj2zmVy+/qWdoqCwWNzV1Yz+dwTafecdZvnh
i0ooNsJlI4vNjfb3tpbggr71YPqcrdAD3Jsrq+hC7yUzbGo0kBl8BnzO8S6lMuv5
dAGGAazO/D/jsZDdSlT5ZtG2eI/U5Aw8+zPS6A7zl41XqLdycq7bKk3Ldyoj7fve
qkUluuXs/Su73eGeYJoxbE9hHEagelSJqGqP04Svd2LqJNzyI5ADKR12IqfQ997U
MtHnP7wIy2Bc6lMyy33OkmHzsJKiQKAl80eUElLsnkGFeD4UUqUIX4BQBFCvD67m
2u2famD/kyF3GmvJx1JKS5A6IVoSXiiJyTn0//+giGcMwp4PtxcnvMt6aSmDYx60
/OyRQBkbyvMTUTXrrBuZVD94ABO8lZNrhLIkBSWl+EDIH7iHw4hI5zVTanbupbBt
MA8GIKsDyDrrXZ2dU6SE8Y1O1VMKdR7N6XgRWzgD4kZ38Bd9/hnw2HPedXPzVwLd
wKSdEfweuifkQeEi4XN83MCvJ2Jig7nAsdQGAgWD6JjLSs6lFNfjXHvi3AzRKl00
M39u/rku8PBPX5bmyoxLnufysZfY94jqe76eZIBEjxsnPcg2pD+UyW87EkDTczYe
hkw+UdfAi8/XAhaxom12vvnSF/qw+k+gzY4Jn6znKgZSzoK3Z1rg/DyKp0b56YXP
+56wk7RzdI8B80kxwjowIw9eqBI48RHwfXGBDJJfeQQBBnaqO6Zh6fBdvs0HOlY7
CAmDY0+7Ae22MDtpB6zT+Of6BiA3Ldgl7W/Bs8kQJ9LTRYKFsI0Kp3BGbC2L9fi9
Bis4yDo8rTtz1TD//87mVZowBksnqQEPJTV5/TbyhU29GmwQx3J0YgknPirSZ9ry
EcVnBx/qqV5mKLt83vHb/HEnMD2qhb/r27gMEyN3fM6eh781xZPaxzenECw2uxf+
RWXNxWWCqomz3uJ8S2p+92ekUK6amAJaP6DFH9dz3SFN3kYytal2CQp56IXLC25V
K0d/lpvR9p0CatnAEq5EIHuAQcSUK9sQd9hMv7rGigG7uQzP/aTy2Hg1vdYTpuvk
39Aw1zIRNLtSQG1MXFjdNFsogu0byQtXI7ww7tl9qM5Oo+rDU0yDkbu4gqhcjaSZ
LZJqmnB+ruJNvO0oA8lHKExgWBt9/5oiQOn489TXa9QhsV7diq7YyeB+k95wb8hc
y6ykyEeyxBXBG8y9vNr4pKmVWIdk9YzFeQc+jEuZpZ0HF+sJ3gQDCyBpnNoa6X70
PQFd+7uKFNYOug1l+pqRqMH9I9M10TdRi8sPEYtqpZogJrcLqP1Lly8+IK58ndgC
9lhANlzqV0Ojz7bZroL8DEwYV0edfBBYtVWZh/fq1Vdk9T2kW+h1uSH/mBmfZX8v
3VlOGHAZI2D/ev7HjnhnaT3pobmnimCCYIHpvdzuzVbQC4z4ISBQJ1vqD1VbKZWR
831hWxFli4W42n+RcU5leloA4X9Eu5cLf3LgH2hMpipOjRWbofrEf4TXz+xvttdn
YPgX+7O/k1Q8epXvEcoac3nWZnYDNn/jFlb6tKT4hu1xPAweqEJ8/yfuDOayqNYH
ASorThb/5onrogQ2ZiTDTb7OOSA13OJeezF4OAhftNA2L5hqJ5HqLEfxlNnTv6jg
l3zhYkd+I+z1A0yQIfmBCHZLSeIE6aSG/kTf354LrEAM+IFmC+EwiAGOESvKHzp4
ehPs4I2LA48QB7BmFmm4QMq/kRH2Q59j91l14jEJScHQI8jMZ9uYSW4GobRAsIwW
eq4PP9ZurEwecxlnru+k7CZghp8bSm3lyZk5S2ql/aVYdmOXieGxFGgy9RFnC0zk
7atMV5r5XWKlKInoxBvjNdQRDcf4q316GmYuxsdLnUTs+CnlzPzgDrx+B4JKPOB/
jefhhZhFZ7DhI5bTpaLAglM1/THRUrW6apS5vN6G4B430Ax4XJcEQqBZg6SiFREb
ldDc49rgBsudxDetZlsG+EzFQvXMvIFrTsd64CmzTldDBAHvvebUxQGN72pJxk+G
HEuSkyRQgfnuE6B8cMpaKgzPw67j0vAUAmx4niaEcQMQv0975X02RvundTSsNvYk
RD0EFmYKcjWT/Eleg9MQJRgWXjNH0s2p+lefx5TYu8C+2iYE7XsNooqEoGVCb5MC
1KocrfSJhhe/85kQDgU1ztQAbnma93zw7NEZ7eq8tjm7inGE9a+6NKIVejy/pBae
j1/S27fNliBOEJFWtOMcSmMUxopG/nKfR2pf0G131f6cAcz4qlDBmJ7uCUBwSHl+
CRogDCivjaj83gqTBTYFrpSylHH7raBlvy1o07VtfxxCMf93vhzVylNDLLRKGaoA
2SMFVJ64886GB3DhataNDlEDTgwb9S16+F3LD8L/CLSzAd16s9SX1xph0mZcj0/r
HBx4vxOBBwqcaaYk24pO/wuOByXUQNUSigbK4vAOa2l+8KE11+i2c7EPs937xh3t
4qHw0gU17UUhtVW9bLEHaab5Ms7yIH7sxBnzgSX/x1J9TO2dcorPki1IZk7eFcsv
dBZDRDIHjoe47StpgjfvoOuhGIchHNH9Cdotx5rqy7rKEA6slsUeB6K4/QyYcsEP
nRVj4DMZBItyL3X/jD0usRv4lBMBew5SzckvmzYje+VMiE7mr58PJ2Ed92g5eChi
oi8rQPR1bIaOThVVBWHAR8wjAUNHhYF4JhGXliINyNGuh7Prdf7jF4yqnUL9nwkS
LxDwWWkUVRubtVJgpMg70FazwS4EE+CQLfHjMPvpIFp6uZhakmTJpzjY17GSqT67
QwjFbHx9axEtAXUj9JtqrjUv1SBeQXr6+Jtb3wAbeMNjeJWLKtFOxz9CgQiPybeh
MRRxXJGEXFVyDdpkeToY388ygYWGpprAzq7+faoIJjDgXOlpn38WGDdX162+/r+x
U6dS1Tu1hWx5bUE9pEZu9evSw7US8NMkmn/NXFGO0Jy0L4qLVwAN2XIfdC7Hl5wB
tQFmyYh1C5no3t2ciehuOHrhx3zbzlwCYADURmD24ox4aGCTmTp5c0DwpHQeN71M
NQozE3UZrZfM18dSP/KoZjn0zT9KqQyoDQolOAbwHXH/2kwIC4U/ltqx0sSPCnRF
y+1YvgIt/2LgGeUV4ajhPS7NdUBt+guTYQTayUwd13g3ymBvX5Ke7MhMfYhrB19A
z6sN2gxV/sMJ34qosZOWUxMfuV19DHxh5grjcQuHRzK2+izAe64CJiVOfROX97TZ
BnaL0M2DirbhZL93iTs71OwpRvz1QseVRBuRadbk46UQrOdiss5P9pceFaOad/X5
2h7kHAqmfK0jB7wu6PXl3ZHUSvUZ/rQWzid7KyTu3NE7BftbxKD8SyRlZY7ZZIVR
hFMU/yJ4mgEeq57Tq+tt2bAbRTw9BObgYMtbjNrIwp6Z4mqYBcCf4LT5Vey4bPPQ
z58cXM1HQjpA7feGQrFu+ArXdxlTvffrJ+mx0iqr3CLiTMiLLasbmEaM5wpnbsuJ
JuEXdQU3Yruri1EM5I5gLITM6JPdRMEfCDbpj3ftmOzVvFn6IcOXmgzw1e+puzNO
xK8HN/3fxESzIBMm/WXPlDAjtCJyb3IWLMIWDqxV5tmJfMy2zYqnWHQmc8+/3/Zt
TvnvJmKBx5qfooA2z5JwkfhcY94/RvWm5nYIssgAnIEaalfQrYa1Gh7jOMpN4ou5
DP7jloGylfgVX2+xreU+NWIXq0/Tpt9eogLWIYhcZTtAuGIm6KY/QYJoRD1ydFpA
UdvNnmjPNGiM5gqCYiAHCmiafKikZ3dFpGNEgXC/Rw5ua3Q7lAimqtgAKHDYR1ZF
Yc0O229g9gRMnDN5iVPJ5+OcleFg125A3IVp9GUhJnbfKJ5fRmbu4EOIv0PTnmGr
Qvi9jy/MDFow9Xhk4Bq54dzXXZ3axH8eCkomxXQEHHmiGeeoeCwiFpIvWF6H0zCg
vlzQshahAL0rAOFIs0/4BH96zv95giBNhdSl8lnP7iwkRNzp2/QkotBYVItazLlL
135J8MkiCMBQdDARS+sDAMFRhtIPvqHHFg0VHsknQ3LLgTzeS+7OFnscw4xLlHHT
cvmeE7tp3MZsQ17kAepKwNdU1i9dDv/l6EyKR3wAbqSWdQoYaE9IwwGY2S4Eqx3b
OuKNfNYVHgTQG1q3TkIHRDyuRcvFTBcfUZ6474u0MawQ1GhCEcRnlX8Dw+OxgCwu
lSW13QB4HTK5gu1TQ4K2MmJIrK5i7I+eRmGg2x/IVQnIrKMI7jRi+f6CtYBV4GWN
I9coro80aMNADbfANr/8IztYbVZ4c3D+6DWi9ZO2VXd5oVny2FoqXaKNmNuiXRvd
TZzJY9WhG1l2n1jbWxrpJxqUHjeurWXVlJLNYl2nvRO9hqoCJzUoCMwWGVP3i77E
w6QkitfOLBSlmJ0eNtjOpdNpgSuHKK7wBVmkUHYwxXus3nZEi4XODRXPcJnDKo6C
0Pprc/0T+WVAKKUwNM8WynMssngllqk5YPwFJFrrAnr7ROMgX24itYC4vuTvnB/L
HC+oSCrbvQYt6bQgdCasS87BxYTLA9bWB+5dFeW3N1NY+M0GgwSr1FzQ4T2j7Aic
8NXp402Mwa7F723d6l1xkBL2D2bxXCTP0IOl4VrqiBraKdxr+8cto6Pu1A0yCSnP
RIepn5lng4/qeVlJr0WPAJqGtb6B2tC5agBcYZUK07OkLYfxY5wKEP8OVtIIrxMP
5MFME61gdM2bmzn89abHvctq1Z7afZSAcS8/CoXB9/lbWm6Kr0YzBJyqo8eoUK1f
2M0tyRIgbfcLepmvRl5uP9nWE/XtbmhWxAJLdUaS9hNa+R/aMo1Tph63C414IPqk
S0x/zDKoM8Q1aZSTFr3pM4WCKS1PrUmComk27fSLYrQcpcDsVAplY1x49jc24jyW
uk3ROMftSHileogrPdjE4osq3Ukvjom5ORjmwz/EHma4zne7AXTdoeUt7z+1kbDB
eLn4/7uunK7qxylctWrDCXsdUXeIP8c4ncTjD1XVNxi2WzNH6P59njXlKB5KCqPb
BZTf74PCecVwXMs0ZV1j0EGKGd3MR71yzo7LGiDZLF/fQ3LHaNS2SmPQ83WmaJme
LPOGxdBWujStWC1T0psMml4x70W6j3oNdIHz+QdedfC7hl7RyYA1np4vF67z+nY0
+rRW0C9Y40IqObDofwolNBEhIz5vJeaKMvgZSGKcHuBHWZNxpCYXAAQshD1tHMV9
Y3U0xPcoWVjYJ0nytusWW/rlyFSQQpn+/Koq1PAQzpuRrGoCNAu4ndUMfkotckBm
0Xb9K5ciwHgdWtFHNPlZQprp/bDYw0fQrKDGvzeFi3NBnD/rQSKdoo8ZN3pzL/Kn
hQd3vLaIBBA1TMO/FZEuTLqulz7+z+p+KSDrMlwTXA5zLUUy9yEI0+JKUHoJ4lfg
tMLKai11vcM5u4lHyS+DPYvS0gOo3p1bGmrEGJH41HNNCBpGg5Hi+v6el847CfsZ
ENlxBi21sY+8zUzmv9SN+zh4/HEetWIto7xOy7YUVhJa+XbBGcdFxGP+CuCDYKCD
2IJYz213UA/GkQsRMSwdjtRwxRSuQgHUc5rx5gxkAAuXtUMQPzscKw//R1kZ1cmW
bDE/1w0S+MyHh67f3njGkGgKM7V/+4Y0xdyjDGzkEjDvKSQhBWv1i8vqcpotzVhi
3iGJnUFGV2DcOG8sbemyZWTcrYz/JOQ7kml+jfZFNLWe3Pf4zAkDpGA5mnYRwDiW
EJRL8DJ2TLU00wISCMn1utDHAi0K8h3T/t0sPmQIXfJICLc6k5cS8D+tLZ1Hj9ko
8nGLWMXHvKql3IlbzMWSy3iranM76gv1qSfLs7gAooyL5bbROdc5NkKDIUPkisht
3fT0zLoao5TnnuS0lDbtLl/LE8Kd8bvrFqbpep4NFnh9j2sj3fJ9Q/0AZ2wtTpKb
v9fNrxrJOg3k7pi4Csh6BSJkmEZ4CKL/FNLkSb25SrOv3IAGQjA/bIDx5Kfofcg7
hPl6rnizU1r46HpjG7qRqSrAp2aEDTT5zQo59m4AkQ+2Xtl5yFCSyihXL/h3+FRk
zPNc38oMqiqRD5YNtv4P1Hn10cCvWvdlASAdcUa/bxXA5BFSlACAPp02d6WQ91et
4lKkeJu+LEflrBBTiszjHReLpYz7iRYrh+iiChDpYr38/RxXnegOCHdq2Nn4/2Wz
BjVcngPq8aTQI9DkzT3JcpW/vJex1WbJutfoxjPQRiSgkagxyucCPtL2IcZwJT+T
SXupuz8hofh61+6dEHN1xF2HOSTvrNl/KlWJMU0my4658mLW+BaqwzF52SFSwohQ
Oe4qf2tFWxVrTFC9UN/gswiGCrYdRVvczNvAmc1QWmx2qhY3vg6paLu18mqjmWfM
eqkjJ06dd8GJ+FckPHgfVu4yRJFWZ1e4XkWqb2Go/u+pSrJ/pKnqu6GmkkoBkZ7A
5wYPxqmHwf0t8CU0XuAs8gW3jYdfJ7uSzqVEVUC57WFwVvbotIyesZqg44lGfrzh
xmN4mAWDf6PgRICrTVHZt78HVQSseTKAaXEWEIlHyHWokPBdkinVUFiD5EX/9LKl
InzFSuVvMEu+4V9wbQuzaW4D752JiuUVAyjzUTDZ++mdewrhjudQaAJVA6KD9Yeh
tvVll8eF15fqHMoZ0W7XqsKpQwe6YWFwpGLk+cJ0ao4Pyq0B1cKJCcKCHop6/Cph
HeH4heXadCIJOV9ADzhHGtrkw7gWT1wc8Yk8AUDV4ayUbfi9rphhnTempGpL006E
RtkzJKO+6JI21SLgPSJ6W6YQWquJJTTaqF3WHvxlw9tvEMph2FpuZhpV9dWc19bu
1hPhPTkw4KxdkXZqQq+4THuqasJV8tp7ZzXw9Z8hd31pZToCuj21H/aJG95ZwfE5
6G8RDhwhEVN0KX377aW+BjmsqzXrOAhEB789axVT+YETTqIsHEGtmeCFob2Ki8l4
Je2H15jWi+UCb0Wru4sSeAUFc9w3pfO7KJCqXom6K3t6bErzmSz9wwSrdlfT4bWu
brdcYT078mhICeHWkQWGuVZfaMmO2VcGRqdKYnnqFsRTo4+v2/Aamw4U5QfvrHSy
901KZZATi1ZmzOJr/t3iRC52PNCqqp2a56jfxJQ9OjZJ0uUueSwxhonGZ5hC5tne
6gFIV2UfL6A922rViDRAchJnavUYs33dUjekqhNOc1Pfgyq7bBxzbwHFnwhIhXUX
EemJ53UWR38PbOtmI0sjQrSZkEJy9B0DnTN75lnpDhPYPlqFGuY9SeqtHkdQiCU6
oqJAwoJt0jtWBPRIW8uIs4OXmmpn3s1iS0GKSiFB/n4O/bvBME5dwLG2McO4Gg30
GQ1TOA/3A1QSFtt9SByux1tuJCBC8GfsABWe9FZvSb77HY6ktv0w7jBUlipNiwia
LPlIZXgwjlLfZiCwjQBSM+PDWl01f+KuANgTMxgTW5xkVjOCNkD1QHqYh4jiHSfQ
LlRXCBAtuwjIWMTTmDQ1Rg7p9KzLX4lxuz+1/4aZulkOmC1Q5uKCUVbczIfT2Aor
muGJHQ1F6Zrmix95JqedLe4zqpIZ0L4jOEfOF4Jz0M2b35X1WLXPPC2vzNe9njlG
ClvSsG0u5XbohNrGzB4u9j/xqXki9ZxXyy8RI+AOWeRHeTTzU5/51YuI/EE/wTvF
Q6Ij8AQ2gVieVVKYiLtFtGR6ONJJIqqg3YKaWAvZCh8iFIHjJvzVyHUAbQfT1qfq
27G0Y5/A/b4w0w/IWnRUuWXsj5Mrw2pRLtV7qnW79+Cq8e/0OwKiVtuW4oIR1eFh
rD/MODsa3k6UHcDP6CayHgJiairjV891ls0zkZl8nYDOnI68aGpsrw4It/wm56Ve
ve4SDET13Q7pzIi5APISFNXl3ksrq0zFUT4Ske+wCJcpkrhaDwYe9wqKsU30/Te5
Lmdpt9h28GdEAbeWXnnUjKFiW+rwyQhSKZPP+pLy0SfUFcPxuqejjdmhX/aVEzDX
kqqGZrD36pzCL5g1Ng8Yh1ViCC04dGB0leMVscLxGy9qwCSSx6DteZuQsNTV4hLd
omF4rMdbg6XHmtLXgwwzFIYVJlCUz5W346V2YChlUEiai3yj/4KGr50p8AgA0mlm
5LqkXmfoj9HplL71aIBU8YcnQtElS8Pn0SSccVHVIreYYWgPSVeqCAwe66NcFunM
x5jr/nCgm73viM/ouqvYF934XzV5vWsmhpQmTLIJLkdmctPigwy3yOMKXt1xjxfP
0UhXsk0s6IW8VkGCxsnZCT4hx5LVDeVGcH2FkH6ZpurxRgVqs2I3Q7KJOhn28zli
4KFcLSZN8J6lqrt80aLx+d8WgKg0HZp9BSbrplrDX3032MyTUYN3vieWKFBjTUYX
Zns/i+ZJKbSD3WKr2OEqiUNs0FHs/2zDDUN4xTXrX1AE7fR2H0Td1NeU9eX0mch+
X3wdc6etbkMklScPvXYZ2AsAURJYcJJkjDucAHiwn/wRF2RBrSDiLI3Kzr076LzW
r4HNkPLftCLjoR6I9l782rxCLbYCzi04eEECZ6ecTPZ1yXM4g3aS05NdLDcOhc6t
HQcTqXjoX/EGpy0OLWIqkwwq2MFpL+PBTZIxsYSkv++nit6OyRHpPkmlq8HO0bRk
ajpDfxWcVW5ZMoIpT1J023ypEGTXzYzIefQoSOzmjKEZebT4R6343Y2thPmKVx1J
FPmX41NIoPaoFT2Zm2epXATo1wnWufXiDmYKSBmtEygOIp8Kp2jgK9Ujokz4Vwcr
mROIKkdL6QVl1leRLVaOtxLxhbGcMXV91L9Fl8G5MlObuu9EzDxVfsO7yhul0eo/
0vRfjxTN/a35MITGQoOGLGDC+mWi85/gazGmooMznJ0k6VP/U9EBgqJmSCSsATlR
0XdkKaeu5V4sJ0ZHfdJ9FW9YlEJ8os4TxVFKvSB6QuXygKd0Zcp2/e3IkBXTUwko
dUlqMx3P7ZsorJNCLGQWyUtc+xsgaLmGJZruJsqJwng404AEDNweDt98pQkDNEk6
963Mt5T5EGYxqquWnY9rcOp0bk5E6HAnGjmrARTnxvVt4SBZ3Tyz519AarpAARDR
9nOTn8cP624M8gi2Fi39ZLQk4u4x5daM2OzVC1Fku0xdyZAEi778MPa5iQsc5iTm
+a3GepFKdqcMtMNbmcxKFtpZ4uhDvFChWJPxStGZpjjipEquxkUtztNqSBnl9Fz9
sFIfhzsqgQLExyrbXMXPeARMTxd/cVmRU1PYWZ/LxbTKth3oHPL4aA2HrenTmoav
U+ihGF47dyz98qYICnZhstBGvXT4RMFD4/fqRcGgGCirTD4ThN6Di9hs2AzV/14W
CuOOskOwQL0kLyMX3JCiJsxoxQ/ORqgl0+kmqbrppI2Ik5CZFntCcEbf7sdhdnas
Q56MltfA+o0ormWoigtiJX50u5/97npa5VFOQ76ZEVD0Mi3fWxdhISVXHBv/AAhf
qO3OcLYBP8MltUifVUpmXnQlhQSM9lmX3YMPxaZivR3EPciSCBRwCmrKmlcwxT5i
jHc5JiG0A6H0UJPygIYb42v7JChSnsdefqZjnVnUeVwv0OoxQAtIcdnoGS+7i1VO
NUOCbwn5lv/Jh3sCnJMXAAG8u1GUo2q0UA+PIIY5VGFhaKrCgtE/hjBxf8ClUvAb
XurMAvueIasUz4ZfOeDXLSKD4CsnQga4qMqQNZPiM14AdkbL7ldb5mUPHKgt2JSC
HICWmOAjSf9tB5Ab0iA1ChNJTJzZd/U9ne3ZXZ8HMROu+3N4hwW6Ib98O1unbjx9
uTxXo280aRkbJfg/k/TrnBIvd6E5p0gh8syUjP7UxEWJhFZd0bzYJNlHt+y0Zitm
GLeM3PVeOO6Gpa/GKe7bZGDvkXRi90GAExoJ03WZ0KmCqfHddeGsZaC/zIbmQZGF
5i+XAdyjzVKEPS8Qlf96fNIy30TFBJIkbBLtMHakTrUKE6tdyZdom1qnLysyaVEB
cIHXmxJZyFM1Yo7W0GCFOe9DNDYXXa6Ox5DS9HWejenGlt3qmOpCYTDSycZ9mMBK
n3gCyaDPBt6G41npoSHnvSYLH/Asp4Yt7cax/Er3XAphzUZuHJsv67S71OmykNkj
ksG5UMdl2i14S0Pu5B/Zp2NGHoEwuwzatCVn3WimB1+BmLL89IT4ELOoBeqMRRW3
b1Mu4PG0J9MxOdwQ6Il7WWRzEHZWBKwHFsuYoFLG5PLH8OTZKQfnZpYsh/XSIcK9
jo7/aG/7L3Qcqp/vcWIQY8YwKP3iI/oFx8YTzMaOkjRiVxxFGD+wLW9gnjv8b2Bs
M0rFwwEYRPsky99IT3WLm4m5K8neoVHeqRStGQr4QhLS03JS8uBNEnSXNPyNz2Zb
05Or54q6MN5AU902ksG3gDCPPG9clvSgoh1OjRgLJ75J+OB5MtBtLMjiHzvzzZZD
ZoWioYLveN10uVyh7I8leUVwOJfVPpOR63B99PNegttIl2gXtY7w9Q6lIx7mwPvZ
T01i509feC87k2lb9dHpiI/7ivjgCYA+NnRi1fIGyz/5C+TBtyUtrnE+j4OPSJ6b
hGoJ8/2qTRUFJ29NHen4Ia0dfNil/9aGhrvNBg+vprpAzdDv9p7lpKk6h7rHExpz
cx7XYrDhP+r78frb0cyzH1Oru7NiWadT5mbLuxuHul0ARjGhykrI6nEHje/LvxAz
jgFi/Bxu7WBFN67GQOaSk2L0IbGm3bkhZTWac/u/u8qGET1Paz5R/jTt7mhG8rmq
fbq/GnXKNzX1bZynbkq+5fE/GBVzyj0KrHUrmOCI5Uxx9/gLQj8sPpuSU90rYuAX
cWJbCj3Fzd5ZFSMnPVlawVGC9yoTezcer6RaUJZjpbNq/udjyx+PcP9hZKw+jNCX
geuv4lwtl4DmmFl04ufYbEfJujTYO+zA10yT2Dm1kO2HJCATqZ903LUjLxo/DHvb
vBeBP2uRZSz0AkHpK8P9xtElALi7GO5qnlonv1SxNkF2OLv6vC3veVLxLyhZPNqA
WqnEwFBPL3nINTOrHSQkV85VjaWliEiIkq7+Q5hVGXulKSYe0/QpG9Smg1dAPQ3J
VyoZXdQJ7OO/oAg5szaZJyjVcViDPZ3CvnCQ4X3aC67x0C2SWRMmGRf98Us+DEPE
C3CNgDYxqMgPhIAlTcKwVfPMDgX3/5SfHJzhYzoiocCcAH3iGprPzhHI+Kh5TQJF
N8ulunCbumRE1QLpCuq6DC8Gx/9ngOV71QoL9uJ9G2b1V/X0Uqt/C+02OXoRRxTD
CTQLl6MW7xvyHJZDiWan1MITJzDGV9CFnJW0qeqney8t87V3fC31wZF3+RZ7LOOV
bsQjrvfrYwaLrnHHFceTIziPmzBeBE7HxYjIR9PL0A5hWPhWQm3JL+SWLfsUxv/f
cJ+LWWVRuBgprZjE94rRhE1/L832M7eRDz0+aeaZC7Zh8NGum7k7dhpG4uHjnCEW
VqWIKwrAXTs3GarlQvmT84FKuiPp2X67bE8ZFEJc0+oLhRQQCs2G4SZJxj/XofWt
hKjZEWu2TIpvvG236Flnqk43MH60igpA6Ep9FiU+YhrgEId1Ty4r0EHcsj72ua5l
qw+kwXa3dGmsJMG72ueJ97BYpgUyU74cq5FTRGXELGIDmUOdicvB2ePviUDR4BwJ
Txx9Ce+WwqGhjxAc8zCNuJdI8kN7ERThYuOrMSa7vftOYXYbFrg57bBJBOcWjAzQ
GMcsK03er4EEBa2xwreHYAI8zzhkTjEON5Twww5WIIYknV7NalctdJ4MaukozkXq
P8UDc/rBGh4nvBsmSOR5FLrFa0b2w5pl74MIVrKsDr2cPcLAnK8kLRSzIldWp38K
SPlHdzxIH/4xHhJulpex0eVse6ZowaImuliMUWoRbDvlrqhc4YDAUyaCgIcOcFGI
EHP9iJkVep4R0StwKEUamGS4wDbJbSeDectLT8kTBNyxx76PdCVft64+qzRQzdWH
98/FnF9CCNLTxfsEoA0nKuaNpPCiDNw30UPMaR199oqTUPEjtHsfniWK6uFTCzkn
aMeDP1q10SabmdYEXRZpsdSx84mwPzjh6kxEs6POb3Zp+JGyxIuu945sQrMc+3TO
70yT2g/z13UMXO/JpxUKwFEwXqOEFvn8yrp+m+jkZB60e2TzYIo0EJnNFrsd9Sii
hc5I3arlZS36/YdQ6n/LXRYLHpE5+MM+DJvPJuJx4fSZ9NWB8wJP0eg3rl9KN72l
LdeLHhN2rocILVn8Ue8biLzfpv7CMkNM2baNZi7dB/a7r6Z1ugtPKvUySTTQ2tKZ
E22xFwPlxRHBCD9x5NT6NTdREDgJXJFbppm5wZXjeYMsjQi5LDBL+/8VZix8V0Nt
GZP+0JPgpIJTbrccuri7Sxa/DmvUJLQ5Zw/UjmK7vci0NLwNQIcpKMKK+Fm+8WAZ
rqs5pjRZJUbIwHQ149C90MNSNx3LWerGCsm64UyrR1ADg6NzhhCTHLSwqE+5mfG2
ZgcORbagLc0lU8yCwfxvCIy1y4QNA5583m5EStR2RYkHCLZpEFxXc93eFLCWHHT4
lr74qLcJ8lnBNif0P1COloz/0XBVK8qNmuouKjBdYMzL55RIfy6A93eg1mLV5yMc
Wwq+wvoFcYjsJa2PtNjtUx8ERrlXbxQdbN+UmfitBhiXdXfJ69lVJovUtgD5CvwR
Cj0+rK5Xpcmtpa0XBhfAAT2M8J7KEQtdZqPoxoDQaDRHIsB+jHa9TgH+mIKO3hGB
JFXzhbsq/vrrO6OQRKPDw14xg9axl14fzE5dBM6ZUeUxtKHSb9FRKiRE3yUhgJdP
Km2I2FT26evz5/mjmh8GpbZJyiVxv8U8++/SEXuQA6PvD7YKdZDSVmVMyHEo53qY
k8TjRIfMW5rYXKassspDMO3sJtVcRzbAJZ+OLxfPBhqwKM5Lz+oTfBQCuGtgSCUd
vz3bjiyhc5flE4YSZ8psHn5BdCrgwxDJzmcMNIJxaeUPjo6/rPnm3CWPe2zH+4J/
J2XKrhgRPIZigd6zKQ2Ku6W/jMshpbeVlyhg5m6D/pq0YySEqpykh5uiwn4HrwhK
x9GHJCEXY4DThhPrFetXzbHWWeavVTiR17l3VyU1ucyuNYyyi++Sha8wBI5Zdrfi
7M3ioSVVZIRgbX06NgIx63BIRmV6FQzGdNWOKp8XNRyT/ldkhMP1HjAq1lUCKAd5
7LdL/fL3ZRN60Wrw6ddsSa5tPEEqrMAsqpx90wBPwMYXY8wZJfPMTU4E1GHCwm6Y
NX/ZFQ2SfMnqDlydgL4GVJTJmX/NA3HZAoDg6slCZacb5RFpD60bfxQ0t/fj+/mG
a8LkEoQrA1DgRQrneO/CGQPZl0/TWhyuPlLczoIZFGl5J+nVo/wi/IiC3LQmUJdT
Bq+9MbJPnyUfrIiKAqyL4EBCtKNTZlcrI0Pj6GydGCb1w2QrQc9iUGqChgXLtudB
ZV9D9hoaf9JPp/RmWCb72VVZnfoFyJUqzIHRCspt3xHiJjy5ktditFtETUTu9W7+
HbCLDeq4e4NUQkDZy/GHqlPU47v0mmYjc3SMBbO17Xqdo/qrWQ35x6TC2SfvZRdw
rvT8fHLatj3DZYWhOKnlqKHwNUNqoLseKzO2Wle3qURryCPQLFebycoH7wxcMHjL
lIs0pmNKmN5M8ACNbLXj7xJDrLtU7MwIHsM0TplnEpe46JIicRadLufxINyuKC/0
7X6xYg6OvH5XCb7D9pG0QbETHE4tOOdhtfU+5dkQvoCAftYV9otdc9hrNvrpPJFX
ecdZJUNDTKGEA+DEXk+e09z/x2agLiK+W+6ckv4oaN3gAWEdFwGm6zvgWfNj0daH
ruVnnEydzBCqooogKC4oOsL/uOrNouMpbEG9DeV3F/QiUkOpfllqV4qjZMOnXYBP
qqkf3EnpUEr1xFnCuqu3pl1kGsXMxA4KgaspzG9fmtoH7rDEmclh966iKXXg2yax
mfy9KsGwhw5MKAeV9/F5dxbVGXfKbf8Rf6Evwp4t/wXVp26iO4BsD1aAXgC4tsh5
InYWm8guvy++nhvm2E5t50SODsz1MrUncOtXZ2uEUkIdCKCMkRk5BZPYUVyc/LeQ
5NgcfVStTU0GVxg/NNoQfUurkthspQngzHoww3xC3oeRkmE92oDAvU3OZzivMg/M
OlCmiRiMQGx78KWwuAe3P+16Hu+y/iwO3q232o1cRMTPXI9LnoxgE3GQNlVOJf0E
8EpKVaP5PFdxkYam75u4npxhHXud2J7VJ+UfvMPFy3toViQ6abpSyeDnLocuT56t
Js+6CaFwqlmAJSNKc77WI5jsf23seta0NvdYtBzbXA0qhsDqz2VIxdTmvAa0C8s1
IoDV9KOepFIHQUJAtndetOf7GD0rBMjyp9iQ7VUyvsuJs8IJakFR/eTgd4e4GHxy
+A1caRcZ6yI+lUo+DFGN1AgWdLpY8BFwWdel0sD0GYki7KN0ZHi4G7o0n6rKwZZs
c0gq599YzYX4EpBbpUpsOQMjd8YmlRv2PGTCiznw1wQDEh9FJrwbEoPiSGYYuEFA
UcjwkDvj8M19UbslqWDDzZnB/Xa5PGsGmWnNpNT0L6OCcNqYpteW+T8/mYGIXukb
+I6nPOh3+gAtNvBURAke0XRaI1IPQyFQ4KvTD4kQKFmMq9iCpIY3Vkm9DoVUnEGj
6k1jW4wJf9LBtg377SGDMRGl0O0y43MR2mHK589p4Vxv/iBnfSRF9idibjGq/+wM
nyRRHR4Y1nn93SM/6B10S49kyTU8WvttKtR3Ctf28MOwSVRp3larsc+5Rqm+eTF4
MDTUnFKy3uA75vUx6CI+KzVz5FwfS4XZqCgoaIVi7J7xOY6e9b1K6GJhGAuRNJCh
pwylfULSzERFk9b2drRxhAGOdIdw+1QxfYk2Lnl/pfJ79gYvMsMBi2J9ivKk0h6S
ki+p94xK92ZMpGahyhvQZOwDbJcpWTg648HoO85ILnh2fQvnUy19Xf6l7FH2A3z0
bcYnVYIS+at2kFCXnhP8jHlrfIPAAwFC+ELzQV+AdvgMPeWDytQ+tbNhseDtI5RI
75gck18TwBGOB/T/VOxxni4wexlNUt5YCAZsJoSLHi3j7cIxyPNTRyMFD/Dp5UWD
H2w+YU4b8e7GnJsQ4fQJsnzsW+Ep2iPgm69QKqPzYNagz8NZzNNXtySWR3/SFuH6
UYrRqGKwDKb48wnV1BxYIAi6XjLPAd82cv7362oW5JMh4VZcxdFYTU5f0n7/0d28
zN9TCKC5ltMHFcug6LaQOd2UAvE20pWUN/bkzrvsXDKhR8DRuhlGFMPVmQFXyoV3
Z4XjyCtevhaCLd7dQlxnUcTfx4ATCueosUguR6ZS4mAfF7DWXed768WRHh9cFLBR
u0RndCg7EEtnDkorZj0fhDlsqB0dtnpksMZwVGT5YFAyveK6uQGzljPJCkyD7h3N
J+cY98XQVXVN4Cf8i78TrvFrqDXPPLkARXXjUOtbVLv9L9UrlE22igpmaaEm2N87
EmsIWnCG40TSy+kIW+ah15rOX7t22nhOzY88G8qasK5BgdcuU3Jb6101hqtjDm6n
B9aZoL+oN7bsFpP8gYLQhjE+wrP//FdBvmCn8VsQ1DxvKQe9DQGTULI2G15VQnzw
c04hryvC4fOIiA6WBSbVlVk28DMwVFgN3vCDYQ+OJIIoMzbFcvXqDtSQw9F7Uedr
98RQ9YhhyXKHA7VjAbPlG3WnClZacK8N7hqdJ+BthK8+xFgkEiSWdLHi1FhwSpxT
Amdg6CT6nQRlKJ7w7U2a/DtcGFJADj0qXUeVNZu/GwTpvXEjXKLadnhGwccq3qnc
HfhUSHmFA6ohyX0pvmM6CzllSbz/ZPOLc2MIyQiC2unRHH9AUrG/0kRRcYWW+d5k
6+T6POX19/8StWdlP0U5+4W7DdvOc5Nb7zZE2Ahm4/Tpea1FSx1cCbfAWM+vtkAa
3LRW/vLbhYy6C5ggV5Ftw4ZNVX2HJDSzblkfq52yGNaz/XWAX//jS1zhNL57X84C
3BCD/ucQMkqkz4hP6e7yFJ80AZlyhlqNBxLQVv7kFXDzLJi5CEDMBOLeqYfFN2u2
x05v4qRnd2mKj9q7/ARRo7xxpo+wPfCSGS8n6MCylNo/DjWtTn7kswIFlWvWqFp5
cs+e+BDoikLJgSeCLhIQHuqHjpfH0GRLPDd8y1o1LMig3LD93HL9mSyoJhxoS6G1
UghnQ/103KzbFmj7C1JxyYkHTf7tXrLR739k5eFftcr6Fqlqd9LaPDCkXA1OaduH
fLDUvMOr6cpQLCUlg8zItXGnMHTSPvWXHBqOczFAoUbrCBQRvFvuMOTpbrluT1Kv
1nIgJ0VVKUAmoJGl+BcN5BtemtC6L9bTwNv8KZSnuHK9QUtkM6gcFLAI7MDyG35E
GkrxOIOnJ/tocelGpsymu6wm3wJvc2sM2no/g2wLnVHMyK6US6LKi4PO/4Jnpvz0
6flO58ntRoUjOWEflY6OegI0khF2V8GlVdXEA6mno58upzeFsDsasE2xl73pTR0E
d9nn9FZ8gfPnwZLSChIUvZ3C+1qMzn066XgLVZ6jBaFlJ9TDrnJBbOY+1g2uI3nM
lciiQlEhlhTahGrBl1I46qa1jHzt+d3hyVAKU/gp57rTd7ty8/GQojBQN5OIlIfa
hjITaYIrmP3d2SlXggWgAFUzTKFkSmo8+kxuQPl3nmc5Mic6IImTN6Om8FJQUam4
L16m/y1MKoq6IMB6Y43WI4X0XaAH+AuEf5BInS5v9lR+lgOPTbMSxPEOvfL5zrl1
Thh9MkcVGQWoF2sloQBLiRZObXgkviaoV6M09Xwq6gAq58PywgUsFcHoB7WVtjya
TZLpPp9IqpBmSKBEuYAOpPIl7M2A7ixvxcojXA+g9u0FlbHKlns/SyGeHaQCa1kn
I7AWOfmqE8L2gyqRXKP5zb4x0H0C4CKXRmOKx1LC11XLn1nJhYO976MIlhuy+PCf
wk3sO/EPl50XDJxhMt3S/ZdgqSGrKE9VDoA9RqvRXGj/jgQCTPkzP/MW/w/5DEJl
67YYkgHvLXpKqj2HqBrrJacNq4Ua7gt/p9qbyP9VTMU3HCqKAUkOWuM2i6mqN5qY
cfos7AVisSGJxaUoWnLP2v89luTeLdtM01MaQi/CDxB4WHBSNUa3TRGCQJteK3wt
XdT+P4LHYcy+wQKBnTD//3/fTP03m/LfKZklDwc2tHvNXsPXkfCXM74QR5ZIw4z1
/glPQBW164dIpvCcYSHEqJeBHRvAtaRzKxe3MpfCJpRmrt955UhjM0wvSzvN/MCg
TkzL1rTOoHLUMJnipi6vCATEXGcjuxJ1u9DeYmJdvNvBADrWVnhKBg9O/l1FDPsA
9L35V3JoM75H2mlwRSPjiSSUTIlQR/DoCwGEUdiaseBC83652QGBoLLmtslIldGv
3DYhvz2ZA5L4zSn/Q+PZ38yYxrpQqYf+yRMgQNc5EbnRkV7JuxKBuGXQlMWbM0pv
P1cbVmIAQ/0S64EWUn9fvBf5DVMmfXFUdrvx85K6t8H90PFkwLXtO8abVw7lGczF
zligk0ouCtjJCsM/RvP+sM6QnEgr2cEYVLW/oWifFOhcVpxhtD9g/H/FXaMZtonm
Nmz8Pn5kJzbwmVBNYUu722F1EyBmstP2pU47Kf+jtA43XIG2LKh2DwUL0TfqwQkd
JBmNzgByD/7aW7MaD47tyC9VwnmVkXh31r5mbFFJbkDvhXVkF+1PgAV3E/ywenPl
3EN/O7JHutg2ebNsFYS+ER9w/pkGAmZJbrkpUf67DbVZenFTArKJdhh3Td9sj6m9
oZLm8BTsHYAfkPb09rytgkXJbyMz7WnxYVJ85CpSzaEc6LFo9XehVFOfHPWEy+e7
V/TEDKdoKtHzdX03P9xcIqiwqrGcDMPNGfXjzlwIHJBQoABArUdIPdKU16iQO/Xw
jrRf4qiSVeKWBEkqK6PH5EJQHxVnK06/3elTQZIoEs5n9cGM36S2qCK97gs7CCVu
cxuhbxme1yY3bOz9sYJlisNgSKQPG4SPeB9BNLUYS6/UM+ciFqhQ+QJVIEldnA+L
AqbhkB3CvOIZcHv+nE8RJXD9KamDUO/wtkDpkaa+/b7BnCVRJ26Sy8oozKgS3HS7
gZgN/N5FJE4uqbtQbM3My/EnE3QclFA6CDPbrfQaiFGxPhZiWywKQX7Ics9z0A0x
pvVsza0cApgv14GoDnSPQv5l+ar0jJ+2RY7dCjMd+eq+QfmeNG1qR5RUcVyx5pSM
yAD2Ov7CQkd3JsDoqV7H4XUAlH/oyMqgImHYvFn2lDObyVX3Nf1cogZ6WTnxRHSw
CWR1aIv4SqvkdbcyMz/0St6V/XzDcXEGdIlE8z1WZqfSV0JJp1hhK3VM6TUaCKzA
KwHO4/xDUTJ9FWcrA2WNEsHddhMkmXxHHmmLum1+o2+K9o442GcOYgQ6Vmaps+AR
VD7DtNRBuOSKWhrSRvIVlQREy0ObLQNdM4MZZeUDSHvpIHz5pvfiNZDME0z8T27a
4jUZWc20Xa+6PieMJ4HfK0FxNIkXwq1dVI4/E9tuxgLP9GT0r6XoCdv8dKHsbOgq
7kat29apocBlPNCSYGczvmMmQgLnVWUMjhr1NoENAdMwfEURnd8naC+bPxvKUgn1
mRBJEiMNStYLkBBGzwCvd44JkwAHVHfCS3iEuNSYVKr5b+FJkyQbkwzyfdEEsA9W
ul+/paraBPhZVBqiINPBNTjtsZNTawdIgI7bcQodlVRfsyh6A5VOS3aDqZRBD34e
q0Hq3bqY15cTkgc7I61wsACfec9ijZAUo1qmg69IrpJF/mcpy3Ev0fNikfEPjhWx
w4a4vtxT2bF1dqb0QOAjO9+OmyafPr6Fstp30eX553Yhmzv2vwI42Z1nhcEt/LBf
lyqQiTrHp4jjqJ7sGF0WCdNn941CAdm/CZ1nQQJ/bGU84GIgSAMA2wiZPkIBZK24
ZnQX9W9kVKLDE6+9wDhmNfahfewb4VGDWTfEt0qL88IzdGw6j99ZHT5b5yUTZ6pb
WCScuEuQnfQUpY+mshNB9Tmm2kGjp7XxJ8XxjjohAGIjo1US0hQQ2db7jsq8c2kW
ivvcyMCMdvnaEbEsMEesEyUoE3rdPSCQCtGJnnL0a3qW5Ljb23B7j62aSF5anOQl
1xRP8sRxtr160++RcxZ8WsY6JrjrRZPXqOIZ7K0CFa052pUoyoMtC6uOSOUYzxN0
o34SnLdbXtHezexOwGtpkTyiGNWMm0ZZpsDM1pmuz+nFexYHhxN3zXOghSjnykYh
PcKwAzzynY0tCx/ui4U3+rmQ1gTflVWHPWL2/zQl1L8wV6Hrd12jI11zzhjid1Qs
PlRuUXMi/H+BFPMYr5fIO0l/rROpBMAQQAFAmzjIux8iJYtpdtb+EVJ6Eb1dQF/s
s/HmgdmtwcwfbPdsYVZzdOSCJfzIFgnIYNLs5NrOEUQyxhH7mONaPA+hlPD9YbAW
ZicOVgw+yT2u/jYjFQMNbh/AbIb7OXRYosrvR0n6Sy/t5IQ692CrnJTi2mwtpRpS
QkrlGpoiwn4ji7vfTC7VcLe4cX6Q0L2L9vm2V95N1yJ5moRTKvk81wAlWjgPDRtH
LTjnsWzsWirjkvgzLzXZtXpIARsVKR0/6PED9eh5f1f3R/IN3m1WiEFnZc0lz5bP
n9/1rJ7O9g8LWLROYwYuhUXdGhFnnkkW/kC2lP8y8ijeFz32d2BJCcLB3HIZRXAp
dkmBYscXVEuYNBWLf0CZ2DNuq3gEVEdZYAn4IzFG3ax0GSUgQwbquxo/m1mvblo7
GFn6xlHOoCGpm+PjEWBbXHOrAs9ZqcbLTWpsER3U1Rb9n5BPToafCjR+v126YZIu
/WMmBqHpdUxxb/ablq6whmLKSZKWUc8p4l/H8Y4ST74dVWK/XWBT7OBE+mnKbCj2
OPhlEBPVhAG4OPsPJLXn+Az/x4rhjdxiC9lipkA10UjJCyPr/dRtqGHg7q/SYHEV
pW9O9jUPDzhri9PAHYqyiF2R8MuHhBEipY83i99bUPiqXEelNdD03nsooSBfxyDZ
8kDRpS+Dq9/SyVxf0TV1iWZfdosRMQUaUvEOYBFguIx8lg34Du7Kk/RiWFNSZkt3
de58A+KzZXQswcgiCMc4cumh827J9j+rj2yVqCKBNLsKuoCWkfEiyMx56YhB+j7O
q34CBMxsOTxK0L+drhHauWT//qLa/5zDlXuwNzEuwgXjGp7vHs9EoXXU9BFXBNg5
OBnZU86v4N3sVQ20YQ+77TVDnvfVcaKbd8Ar4A2bV9ZYgp0iSZV1ehE4spQTnVXh
CSCtBACZMqB/4cb9IKGzeavI7YptzlKRWQU+z8SMLtKyIrLqo3I6a6ITClGZBnUY
g4/irK3SaLHnWrE3zdCx5BPzBP5xsurDt5JksgW6WVkRiqVwamhwOFOfMe9EYlzA
57ZZ4U5db0b7lJSxyKOPUMPFmdV/JV3eTHwJSYIr9y3HX1rbP4K5KoGGyIwm/PfZ
4ecAahHjxVYtSnHWyQ49GkC3o6TSydZ9sdhzS5U+N7Dlz6I7GPVj44a/97tc1YtR
YqlJOePUGKrDgpV05bi4XGKYk170rZgIbVrPkgKn7hcotxR0Ul5dgHl4Fn2uk9KZ
CZhrL3Drgn1J+C9xBBIQ2wThpiVZIU92Jj8baiuCoNI717hZzo9hRddtP+M96GWv
NEZvzuICu24oJ81fPWtT2TXJ3MHDJenq8oaaw97BoJEgY1OWmDg1aKvSu6Tgo8IF
GNFmsgminVJcDpX06li5ZTiViaPb6qutnad8Gu1+2wkly/EUz7IxW8tYxcGk1o58
i/NY7HKcuaT0YaDaI+OXOv7yP0J1OTRL1JTTEE9eSk7Wn+o+lNNV32bORRSLqBig
xNYzhimxV2mpKIqO2FiRXI/qudqky8ebCuFLbcGoI+p1nhtDFFKbiEFqbWeqmuq4
BKjyp8ZogpBmOH1c9N6aXNXtd4ISzwcdeUtK0dnpzVLlLCHTs9+vUzTomD2vBl1p
HYd6qopGq49MabWVdh7TqAg0piGIsWltFEhLO44u3TqwknKJp22OQoWv65UefUNS
7WzjMczY9jsg0lAkgLqfnS8K7vZDgqfFXP+Xov/mFvWQ8+OgQu0aaP7wVlRs2jCJ
q2Y+My4GWW3fZzzBCK0J1i8KNY5VjLPjzs/37jFWoIqTtZKLulHKgCULDOpj8bE8
ECbdtWedCzr3X4uIWqG+K3JF15pZlbHRHYXf/9FdIHvClzc8q6IoMAFu7XgpnR9L
V0FpAQ6g5OsU2Q4kLMGgF+XUZ80V6X2rYiq5Z6ubn6CrWmb413Rm91CBygnSny6g
pBW6NvAVueV+v3WlIPour+UXN6raX/iQ8XqtkK6yz1KG/Fmyo/a7JyO2fehuzty0
Bf1qlP4CQ/OIQfEr5VOmQ4imdTg7Hp5cxUsb5JZ+eEuNM2Js5yhlTHPFJ6VZ0ARZ
knyCZSfggoNjX/+l6pOEWNIHstYm5mphELHHSLignW/XP0mcYZZxff9PptKgK8bu
dvqRmmIDuIvxoTdijTDJYrOapnySGnDogOpXqgunU9+W9xFMduIW9dz1eTULJuOW
KwFqj87Ti17ASR5vJBPokOZb06OCIwbFw6vbjXb2YpWaVbLAAkEAoxxusP6vzYHS
j0/KBKVEKEEPmxXXdPaKHVUtpC7BpeTgC5oHsx+OP4bNmRHMLEfJvo3b4+R5O/Gw
/giRdMk/cUvytATWlyfmOahhVUu3VoYnTwXSlIWigJ92O7Hl1LuqFWwyVFWKxHLN
yneRXo5PSUv5bjWmFgVEyAhOUPlQPioSVmD9scokw9oTKck1+KXAiiSLgsgRpol+
hoUNjutymD+lrVt19q5OBd0ALu8/PL8Mdi+aT+ZDK8ba9br5P34y2ZrJnWmI0Z1T
AcJuIOSHgUKuEAaymQlxZK/ZghIAad3OaY6kANzxP3Kh01rqiKK6FZxAMvwJMqEJ
Y7apT2fTB39OYG4AMR43M+eurZa3aXktNmYHCd22b1DY0vWFNDEYQEezdhX0vkuD
tSn13m7tuMlFE54YG/tJWrpq49GOR9fVo71durGlEYoI9gWNAVjsirA1gzlX8vFM
6ExAXfmB23UXhUbT7yCQ+3sikvJYihFeHB3ttgvNKhlaWD/QpowGX0aRbwrC+5DL
imcG5WE9nb9NLcxik9NxDubECatojle4DavxjFbOyyAojH9sq94DckfWEIkn8yjk
EVO/ETWsOU4yEkbcvhyhiCei9PgriaT/VIOAItJE/xZzSAz22ghWlQVnYDOedIpZ
U1rjpyZUgdc/6sY3NPj/nv3PeA4mC+RdUVawt3A9eFZUqK5TRiG72hNOO6HD9eCP
IYVC4XmDerYeMSQIMI/OZN7b7NfbCpbSYUOBsLJHH27HXkTgaIlbkeBnG+TIalMn
vdQy0olSTXLsDxH62lvsqnOGsZ54ZH+M3v+HnElMdT7bohTV/1MGlCDj8Z2fQ4s1
eq9bHQSP2MJMh4KafLSppLzTLX7qM/5tDecjU8oyZHYpJuSL0Y9TcQOxnju852NR
xSCpGaezNGegogQ3abN82XPJRllEhqK7RfbWpsjJ/tEGHBmZPWLIruzLdDDxOjGE
mjqLbMy0J58p5yqMhXfL86SFCbVyfZB60IgM0qP9AeYkzetUCeS6mzim/yLPV4+k
a1ppIMZ0Mhct1KW3UP2CmEBY4tUL/Z/dWvDbfDKxlmEGx/ii7KcN5i2Fj/4VY1A1
yJArI67VnxEgEGPSk4jQQ2FozT8hgro3vD1xYpFNRrwuf4EZ/flAcFlWUTu+0lm7
o54LXd+WZs3ewaENAO8r4JlviIpMPVT4SAXl040crXYZrZY8DuRahbadiDH/UbPF
qkY/P22GNh/D6emjHHeG9+C7kc4BjTKULt8pOlTs1sti5DkAE+HQjEKZds0BS4sb
Pg0tDNo6/wNxVrtNhy835iILSGPVhH3K6ASQEsJuq6jhx3zDBGhROEqWveZYBvxs
duSHghcFJt+U9tsLOtw3L8qcmnsl3uiQ7WOEwcywKbYQnrESk79xKnrym21A66Qb
Eq6S2NIGSa4jQOrItvJWn4+B7ztR4EV1DLAoyJCmGb0Ld8MNw0hgQOxrA66CsM+B
FbohcEP6GPRZWoQjDxkQtI8/oFxqzHq495GNw+4ZasB8ZihbMOOF48ukZpoDOqnt
i9tb/ompnU/vRrnf4sasHMrOPEeMP8bM05eCCZ9HXRHFlubKv77YRhmFHGvrskM0
/s+FBxjfJWvQjBKmDf4d6wxgGe1vw9Dt2f2XJiwd5bQeOEViDT+lyrdj+hikbzd1
aJG7XtloK9zt9QXfZ32Cav8vXagtS1Fawk66DcywTTHoxQg66wUw1GWfgKohfjjB
h52zMjLp8U2A7ymyv+4Y5jI7wrlD6DRmzsPb5tkjWPS/V5xSq2Es5TlumflhNR++
fnAnktUo0MJlRm40nkMPiSIkdSUtQJCvZaygpwR1Z26WIYd7X7P/TIAZ6YTtqxNr
eGge1s4mpoFXstGySQg/tNlRPTPLpZt5y1O7qNgA9I7Bh38gyInQWFNzQ8XWdmDK
qXfNQnD4RbNXquMVsteHmsMrRd5V96TUQo+JWlZ5ZtwXaot0zLWTaneJFp2/VMFu
FRk5s14ibRaNwOjyKOeZzopOWxOQ9IKSk/e27I5oehX6naiC/3tRR4M8SvGLIoGL
MyAK7u2W/qlnQDuYCoeiMq8kXBgJYoemhItB+pXQiRgebBKZd1KYHMsXiVVPmX/Y
It8yyJ0r528UTswEH007332DXTKlKL50ti3r0+vs5NiCe07RM51f9IGu+Ij7Wlp3
ljoSdWTDbON4Wi2yX8lhfWPXUeDu3KdHMBTqR26hsB3ZkioDdusOLdAY8au4cnOd
JNsF0BcZOWj7ywI4UAQBEI6cjpqbFxWfn26HfWdwg+csgwlTgzdAEDcjSQ/HBXtL
X6rVu2bquGnke7fDxLW7QhOFoJBbZpaG/tBmHvrs/VSUHprfBZLDHufu9esRIUHq
49J0cAD5EYINDfIayGzlHu9Dh77m0ZPJVRlPipLYYSrn4oKZdRQgGhg1fDhOoHjC
1fsF81sQjSwnbWjw0fpERVA8tIXvFn094QzgmF3RIneyOQkVPTMJuMGFMWMWGkRS
X7s8kZI2MuOjRkQr+r6HmJ6TWyvizI18tNmu2Lx3RbWjxH5ZRL9t3AdDcS3+cUFo
HnRPe+O1sUxlXVe1jKkzaFybjvvxs3XI9oiz7yyGMlA+FVAi0kbiMGAiFLzpuNfI
gWHoGD6lKXlxIL25oLT4tdhHcMAp9gRdxmcRbVJi6k1qpCmADlB4SPaHj8B6/smd
WLan+a80qB6+SzwjN3zbm2m/yvQCdLYjGRA1HVFx8M2++s4ca+YqGBKBe9erbVBV
F1QiTfTaZfoP0EzsZGxMeNLenOeE5BUTBpreyyM4X4io8ChqKZQXlgKntfM8utBD
kt41W3tOJHyB/1212e114AmPqDb1V3kd1dKHcui75ftQYNYmH2/LnL46oUwIpFNe
q5twZ3sAGePBX01byvvqcNKCGsDfV80wwB9b/MCzJ6QAg36B4fIfjeQI7N7ci7UB
Xag2wSblOb5qgO8THBfgYn4nomhLyNdCg3AuTKuIrpkrHl0VOq9mMTqwbdLPLcMp
8m7y9JSEWU6hhS2q/0JGpXibp4NrcfX+Qh/3nU45DoloWg00ca+66NvFS7snbeFW
otGZH/TKRKChKRPwetHbPidAnSixRR+vpUqHYdrKS0nyYccm+BuArrlvbgGbm+gl
YulO5OgUHLmxNURp9oykdpXozRxKkPj5oiYAnDxAdVKR/g9PfB58N14AaNtE99YZ
LRmDYBICSdcPaPnhxduPxtf6wOeWWhkEf4k1dBurPnOZcOHbVKqj++pHPwiMz4ZT
825SFx4OQeP03DK47Bvpace4bxUeDYczInG78gsFTrKXbIQHEd18UQ1gU1crNGFB
ZuCh+C3wPYWamr8Le5DTWx5EVz/aX010r5GLBdow5xqeqO2l4ldgbPnm0alXCeCL
9VnsrQtN7Hlqg8vUWWsuuFy33lnA1q+jvwqgbcgKnmXXZx3HjZn896xwdjW8v0lG
TOqyUOwlf2lpmatJkkBMI+IyGdwJ92zfVNdfOJ6KZoH+ESK2ajAtucI2M0EuE6xh
P0JQEJxIEnao31kqRWFfGbNTXDrO02K62cNnsiaalFrOpaidRwt5EQ1uDUlvrDSO
wAzixFwQ+8fyXs7C76PZOpGaOTrVZ85NBBnbGmE4o99q6WWOZkLTRsYKZ5zazUrG
zZ3FC6kL/FqnKQwfEleNNv3wokzLZCEUa8jhloFJ1UU1vGAcuywFeGk2KOfIvKSd
8aeVMc93ZLWFSMx+kx4iEbaoL64x/HKjwVKo/K0rYWafMhO9HxvVDVfwChjnPjt/
XlOWVVQWPen0tzrS1HTXxHT51MRPUjKvMLCvFHcQ8l5FyaPhMnwvc16ljc9IPhbn
5grxhEuf76wheOSn9aQIvilh80aIgL3F8CpgbAhySXvdmggK42A4PRIej8KOl+ZB
a8sp9FnoLpVO7l+esgYlTROn7xHwC6B1D/onS/Y2zuOcv61s9DUCe6DAyVtFQJrT
jvXrWl00w4EeO+7uy6qDrTDLWL18cO0EfWDsQZcf52VH0DC7PCtBOqgLwk2Rs6d8
pGNEkJd8BkiVX3JETGX5HTexyd3nJb4dHpGsu2DduNP46oBNbgCdcjeUiKZe8WwR
9uY8g4WOXy1nAiLKko7QAY+2JQLqb3tafHcVHtUTAhOzivM/ZAFfNqBDPf4MJmKz
Vz0iPFUl+aac7N6GM1MVfPjRLWTZO/7wuY3BT9FJI+BPMtObJpO9MKKtZY8GZO8o
5JU+o3xK1NDErWwO9j0Kre/XHxHxJEICBSctMhVa5QW58a82spqTsqJUKiNApKGR
1SpQu8BIbRjrk3abl3F4wSbRDmQe2b1ka6is5TN3UIYsvXi5CSIl8oIEgvgvKwL2
5bjmknkXRPhb7S7SIYFKVRmXtsz29F0S4aqofr+z/npScAAf8xm7f3dtLl7TgbxO
7mWKLmkHHaeoLd7PeHQywW3JjU2sOfK+MmTOOrP08p3yPw9ts8wp0WWveQ21Wk7C
aEu6wMlCQ1yz8DNE0IuTFqE/z1cySogMWBBu7W3JEmWnqGcEOchmqX+tQdAFOI21
18TvvLToHtUJGOnVFxCFSQ7dxBwryOA/HcbHfRrY5gnwuTKyrvdq6OdxtiTEiBVJ
A0pubnPWcAKesRCwao70E2Nb/39IgP0KXKsCDUpj+LOIthh9tkICm50vAyXto2Mn
9obIsYn4W+r8y+wR2so8+FXMRy/Eh/0lZhURcoIqnDJNy9a8WwoSR4Q9QmkUsGp8
orpHEH1sULOqt9c2rH/ZM9WBEw8jKZk/xE96xqTCHLLCJYUQk+zNYBPWhBJ+VICq
z5AolNl8FWLKx76iWJVShaT1iJFM15thBELa6Ay+ivJZtymYW9jalee2fU5pK6N1
NXxSdTIiN/0i+Rj+U6uzhvvSJZpKZQuyixen/C82B1iwiJSTlhiTChosMMPewZZT
Z4TMhnRPzBarwrS1qKGkIBdCbxQTCDw3cUGH8zOCkuksN0M8cfQVnS7RoTm5z7T0
Sh3pBm8RHsdHPd5ePuYnBWqlrGJ30i5iKa/uLwFPM/g1I299/a2fovAVyqFQxfrE
dcAwquRbBS4OhBvdlXuWcvdg0wvtJom4L9e9UiZTpn4xJj4Hrhjs1KM/CRaHhF6u
dM4mhTl7L2ZeMOVW5Mnoxy7A2C+LVUVVUUMplYuj50pJk7vtoKlSnHWzmQt+kNNu
/fsCi/PBlKkgGt6ZGJJTcl3k12aeM0Xj88Rdo+as1JFXJwrec6l58SjJmlxbqMuw
LgPhtQsJO+UIp/vYe4dzbQ0rMLCGC+KnwshC0jCQ2PtwEvX/9cbPcRvN00q8z5zn
y0DBPV9MFf/vjA6k/n/xrLL0ofId58Z3qSfKswzwAtpe7RDQlKyGh5xxMD4jT/FQ
HEdEzM/A3/VsDxCzXR0frUVNF0WHfTaA2bgG6SD4B2DOtc/vxJ80F1xUj/QnvTxt
1LREI9NUruu4GbmCYYmv/vBfBSbF8UCR5muKjOLVF80pxVHoSUfsCiXsmunTHJ65
fHY1i1YqHeTd+E1bW+egUcQpPOkMwKuJhpwJ8yQ4vXGAcqijx7OG99TjDVLD2jBY
e6G3f91M6oTqbolNWsLSOMMD56QhXInhnN54cXIp//CDXMSqTRuWRHcshFGgYJgr
257RpGnNhsST11a29m4xaOM4UOQNREOiogyKnja1Q+6xDCpWrPN90tQoes0tBrmq
jY3fICfDVWAJ1ZESb5TMzl+A10DZK/VrkcUfSLaJPKV/gOU7xry2oN6T3RQGfPvt
oWjKZujA/lNBhk8/nXvophPBUjp+KRQMAWxCxydituuWvRsDGHv0BcsvscdKoua1
xuV7pJNQiHeJKQ0ggkwT2+QjnW3Q40QBxnfdC7u8gMcQwxf88mvQEqoMNkbyhUkN
EnLZrN8xkWRxELA30xIYnVTOFf/K5771QY/eYWXVn9C10mmMZr6Xbj8hIVEeZq6C
x+uP0+bWJdtdKiYrhcCDdJqqo0wIVHqfEptHDuYu4KvkE5YCxWVKFolYSSw3jomr
REMZ7jc9RbTDlzrBslNQWcndtD0ocz7z1x4PsA/hmleH0OtRRp/YfPtvirm7a3y6
n22nysK2nGO3yxxI3OchYWAGbCS5uzUsxsdCLLk+76KgNobM8p3jJ6E5lEQHMglB
WAk4Fb8LdfZTDxv6mU1UpjTVkuk69LWiGX+rngvUm/AMUqvEWu1TycYoS1agd1h8
hB4WMZDjzeKKq82cz+E9SugXEMZvSnJ898RIAlKJxC7/u6ONygGjEvPzEXoiBv3F
1lW3+O7HZsjLDvUy+JRRf3eIUADsruqCIoiBZh0BcRXSxJKV0oZg5FBql7rBdDTq
uOLZxwoYutJNaY8oDHPUjW4ERdOWv95Pi/j4GYkHfMaNeQhP/Ev1AGfxfYsBMXkd
5ygKlyvzzjLymuLx6jjw4Eh462wHhxXPVtBJDyS80UhvzRDNu+UJlI5q2qI4ZLNi
r7dtw1Df8AVdw7Uv7ABX9OJTcA8Nabv/MQvVIl6x/whnkOb+80gvq94vl6unhYEl
p5udVfiHCSjAHZuBq3RwQo9Jtf355Sc7qXrvY8aMTr4s5NxXtLzjy98j1slBuJAm
78db0Fb44VGsQo3Bigt4ktD0tebCj8g6sCDK4rsXgUJuPwfVftGlblGWBXciMzky
OFmy4CqfTTb3MiWnCFmaonqkMSrUHbNiUNLKL5sjlG8MnVY+DBoxSByiFaPDDWA6
TG6vYJZGwgtTfgSFcwlBVc9xXvqMxuoHVN+OpJJG4jtCU3A5+3dL26uWKBt3xmif
hfQD0rqNEB40Is+RgaJLuRMwO0atptlYRWpSbfcyUzjpV4TS1UHD4307g34xphnn
uCdkf25pCP/vRP6Owyyp0TTvSV1Bapu5rjZJyavWq4eXnh/H1t2BB6rxuas5IT0v
SlEofi+gWxX2nmbx6HZlU2erhBONT/pQ0A1tJcSN81rOry8RRj9I/17VW3//4Kz1
ZDZxA7EAV88na1+1l7VZycSfg7Auu8nBBy8fClxg4Maj9YKon34S911lytLMppvI
iXZIKgnRaJa0PUQm5qO3TVjAzlKftyUd88R2MLxBTdQ3ThqZFGmBX8djAhXdD251
hUT+S8pUg/ZL7XiYLD0+prGA+wvIuEuHkRlxd/DruRZs8kts4/XH44FBjE29rBTj
WxVLzxLPIy3rIGVwHFe5bMRS43pxdw/Z5jhW4n8T8h7dbARDhzx92YYZD2hUXxwz
igSXBteiKD49jPibsnxVAvbJ/4Nx611Z8FbYkktO7TbmnTz/IiHwaDhCmUEtiwNe
NWBAEJlfJWAVT7l3PiAdAFfoGwYM25M2pY5XRVYQ2gk69Vsyl22N1YFpEoYEGAPn
E/DiogfIcC4kRwJ+5xrG+bg0MMGTOalQDR78ZJoX/ErgdCAputPP/wh+FrXRy+7F
/bdfw3GExgYaTlScqJtZtPpMf0MR9PZ9o/Uec8RKGNN0EpE4iNH8nEx3w/02XSpW
qZgPEJjGDVRkAh34dCNhCZfFUQhm4A5jOIgSLXwu4+UC1wL59qJAaF6ZzTnrChyv
ovnP0y1+kT+laJ+xQo3HjD2dYHXQeG1Hk5wzARhKfzdqyxIYjLka+9c0j5bxOvM+
/HIpydpyOq7p2rgg9/XNrKnF0X0Th5j9JX9sXuX521ofPJHskN7pwAHynewpJQIo
zX6BsX/3YXMCdEVj/lePnNWgmWCWM9VdXrV9PbKHQGDJGi+vUOtmwn7ev9GGSpUI
yMUFJIhKJco1P0eHjVvzYVTwDRPK99sbNgUHbrWaELuZSC4fNbjZUO0jb8Z0NxT9
4gbDdnOMTtieu0SCSsUJ9FfRWldN3Jm5zfXJqdzwFAY/B7sL9T9LT7r5EWN7WS6s
vBbaAgasVdhWQSD8fMLKt7XOhqEkiEh9ChTT/+B3ierpvVYTrHqUWX6U3ksOabBZ
amiwvNGOmuQOqDGXzMBAzWd5vvKzUdlYXXMRC51+sNMMObYbOvVbW6aIB9+OVEcv
tjH1sfM+ta77dXhx817TdDwXh5O0TuCbOsSUwha3KhcSbEuVGGdjfLg4TAw5aM0e
6ygsfHRC+m5YaFt1rOvByrb7+gu7sJn7GHWdZ+AFVZWpULHy4N9gRNe5K5qkNnyp
/DJP7BSGtKIjjl6Mi2A0hHjfQsvonF7tbIh59qHmvCibK+GzE4PjU6+/Giiwq+Kd
4YiyIWWbccaPA817vrwrQJT7vf86XNpyG8Ewxc2cVsK8TC4R1gf5gI0Q8Z0Vv5FL
xQEl9uEkZkGJbEyX9EQYZklyKYYmv+W+MKM86drLX3KoW/bXYFXuPdQ12fGHElEQ
3DOPac0xzcS1K1Zo55OK5zVUb6+sCaJyeutWqE7VBipt9Q5A0VnVUUZJ+HypT6FQ
inapkFk3Tr5V8a9nXUkhXcbVxLWqZODwRoEbIoCuza5w/7pD4lorDmVqjk0z+gjq
GpUfzV4odIjHtRfP4cYzx72Iz1MNEGo3xTpWwSXzjJVajKJzeaMFWEd6l7U3enek
TyxvPkkTZalBdDuXhbnircaqSKMG1CrezLSBD1/U7JlTP1/rwfVAJznYKWB6ko7E
jsOecUOZIxN+SaJuBw8mpKDeCEVtAgGrFnpQltRLoJKFF8Zq5mhz1fcIEwPTeR24
DxWcwVi5dOvOFGL8Wv14hqyXe59Ltrkwmqj9HQSIGXNkLe6YlIs/0YSw9ciLu8f+
00q3hF14+icM3+A7Qzqv0X7BaUuqmbUCMhVdiC0E+5jScnzof34nyuHWFUjzB9O5
kZPN+K6XU7889jgbCqih/rRlW0km7VVn6YMdpyJpf+u5JfreCBRbowWAKqEpybUV
70CMCrAYi/EzIFZW4EUMIBZM3y6FndNSVJgwfKSr3vW+FGxV8ojkUef33AC+nwRZ
A8ik8NpjbMHO2wTMwtk8BM8JAvP8IsMRsEImiNvD7zaTvlwL6cd/68H+TWk9gEx1
p2a7L14/foXPGVpOCUtMcXdET0W2aJQkFbQXyCfiZPA7ijmISdubHoQxith3Uamg
2E2kIxf+fWvaWsxl0jYcHVMMpz8d1H/i+vZUr03l24lv5mI9H5ZN+wwlQhfwvhsC
u6N1xnIWiXyQe8EpnRROhiYPiWpbb55pmlh7JzHMnwF22YP0Jd1w/MJFYxa9ikeu
w2i6N5Cplpebw318/u8X7uo6Bxkg3Tw10NHg5b4AJEQHLnHV6qZNnWg7VYT9RF9K
eKP+UPsjPMidl5wy0bOyyhWmD/Q5EMlNPnl/fGOLaBAb+tODARFOsUd1SBPWW3pI
r+YdQH36qYN4GVO/culFfJxrWrkMhbGWa/55VD7wyw3IfvzqwmXPiPPdR8ax1MO6
nPggs8/7V2bGs6QSnAKMb9kbODawqfRELlmvAWRgPtRR6eKUDJ3o6MdzKtcbw9/Q
vqcH4NDuR+lAvBi1dQhnJw8wKsvqfxzdMPk2Wrf+FD2qunSkGVcA7AaVJMHA+syx
Isd+N5wL229ptQ5dSXOw2JScDaR4iPgvKOkMMMskdu1zJdaJaCObiTD5LsenyBQA
JfhOF/CrbY2d+ctludmgyDcDHQfdUp5X8Yq1AhX/CbIKwnLIYKrb0amaBoGdgKF5
td1fmPd7WlflXzxa+t3DcJDcyGA9xDU5q7w9r4Kwu56+5jvfuCFJjakPYMI9TWm1
I5oI5Je9M/h8oisRgY16CAnxn25D3/BJ3Xb6uL9biYsAJo3FJQpqKfbx1cu3cQLv
qyQhBSpdsUV0S60t2phcGdA8TRH/qZzK4SuQ2jiEco0h6Hvw2iV/bUGDww5RsrkI
AaW4IfeKaG3s5wjdVOjcBCdEffOYIVPuxmittUyTo1t3q5jrKqM3lsn6CpydEPMp
F4/b5Smd4+D7D4jnFHNVGZQNfRGlJZOtlVsEGi82a45ThSJVOqiJRtHGcLwn8AIX
nOmd/izzRRGaGZdTrM3B0yF0Xhr5zzqI6WzjetG3eNPWGaFsxdOYMpIQBgzdsl3V
NUz7DZbwbuYzCrZxkH14RJQXVDHRlA2HaHXAQ/B1XMvtt1Vu42uXdgOSkh0Z4SY3
6RqtUScXFHofTZiwddypgyIRQVYZ8TznIxMW7OxJ8hQQFnZMW+QNX7HK4+1sq7oS
L1SjqYiX8L2qI14FbFv2OrTnYCLmh4IRhcc+ZUBAxRI8g46+bCZrg+GUo+lnwqRI
m8M8nmVUGHzwULBAfE16oEhs9ZTmNTZPs7Oy7CxWGqGnKAsdfGOAeEIW+Ub7SI6m
KDkXViu9rdfb9/jF3okmX3C5nHYvTRf7nzzwcTpp6ytQdmlpwBt3fpdbLhCxgsjt
4xr1quRUtzU/sXoOwjazFe8Zti0rBzf8DGQfUGcYXYCcq1zRaW8O7jPQJhrj7lV0
FDN/0jIsw8iBKePEJ4fMn2Gdrkts8EBdteqkrLOF1L9h9l1wSguLsbpGNloYhH46
g8/+h+EYYGzqSyIvjdFe5Ghd6crWQvC9+yhtYsEvWdcX/Wfw5xhueCpdNpPXdH1A
FEozaXpx5yXdceyw1dMM7jNqHIwNsSGbmNyMSDUOuYToY9/LMbulhlW7P8dXv9ia
j+jzva3V/KGaZUzvV377gl+HAA3RTAgL7dKg5vYg0GDwSvUTSNk7/znC9ZqJZhFl
bp+btpSqNnPRyy2W5N8CbFkNkd2R2u2cqJM2Z6xtdCgZnIWrE4+Lu6mLuqfLdT0/
OnQO0wGX+LjSKHQZa+EjERJZNzuLkOSEBASmuROeC6F2q5LhUycwSQQ4wgJ1/xfM
MJHCd2lhWqlhx32LafXPCzO9Ho6k8735C0iq7rq718QOogHlMuXRbpA5MO0C/ijI
jchKzI/L0KzEj4XA/ABIJUWq7cPuUhY28TSpxwK9qF0PGURF1vnloFXVUpBiikxY
X2vWt85AEJxweDGYIn6AH0vtPI9w8L52G+3lUY1/PXYXxyI5SCvca49BlT5cOhBs
KJqC2h8jJ/4StGFfblszK/6wtwvvGWyc7TKJkVfnrxqZgmB2nXxvxxBr8RFTiSi+
GMN7CbxerEFP4a1ql9xhMGZsj5lhJjus/oFFoTl/CXSkM1gf3IPgzvaZtSvkJhSj
k9y7xR4KLbhViVzXHl8NsaJ1W35o6Sh0OS/hK8C6AfFkxa6TCvHbN7GV0WIAQjBY
7bEij1navMOpnvj52DJdtJcNBYh7k01IlPl4nVa7h2BqKJFnTEd7I/UMN1yCGU+R
De3pUENff/9k++6n4jV2/SLzDVmLvfr7/WJGJyxAgys5sj2sZnw9gI/KBChVC16G
YKq8uaecmygZlFl7v93d6kLAB94L6LPQbr57ys80336GgsSsleMaNo3tRjxgilZx
oBNm10RrTn8WTA84W+UzU+ouNtu36A0SBHntwIjTMGwazy5DlJXC5Zow0l+UW9GW
X26kj18CCNUwdOO9570xcCl683h5Z34Q5dXcC3M/8y497wvLwOEajJWDmzFqnkg+
H0DVLnQBwXe/84nPMfF093FBaMCA88BYJGG+LnTwqHRBUfMiMyO90IOuHmJg0NHA
HQpqr56n0IFRsEPhXH1nKE0BawffSVOds5B5CnU9i8D6JCKq4ciWdcKe1xk3mvL6
wTRITsmldQzIIJIdOAFIWzHZ7nExr316NL5kYWxw1lxc/y4wjmk6fvSzhiZ29Cx4
pCTd7IFTeZCPLyygds+L/+pZcQWOc7+G+U0GcekgzbXcEg7D/dtiuUrLPX3Lg73v
E5NgnZCNJLVUciHQcuLoZxYcOU/ZI4qbqcoRN0YmccS6xkeyGymVbbQN3tv0cfSR
s3RB7+XpqgjI3tpOtCoRAvol2GFGRE/XNj1kF7ipv2KWAvYd/OJC5Xn2zRZOOHUg
5XVjOHw4id2efdXvfZUUhPzg4Bc5xBgH0mxZ0dWoKzWyHn3MPOUkR1WKTapCy7Pa
S+ZLsBoc5f3FQkb1y8FaU0hnuLyRYvANMwaq7OWeqSYvdB7WNyY72Hbm11aJiAZV
78cRWTnV2pJ0K4Vr7CZKv7ZPfHFwNxCnCb1RNRL/L9vVaBfu+HfXK5rcPTnEG5Ub
8KzM7n63/Pgs+CTS8mP7qWiMhJ5IbVjarrlmtqh7tDbSYdNWmDYov2+dso8s4VrD
bd21sLPe3cJkCzOhVieXGOjuXyRRhaATglOk9Tbh8DXlY7y3dI4fx76tlqst3ecf
5xS3dORUICxoscFsjcSIUXNFe17lLtXRO5go03C/8W2pM0joime0yZDayLR8xstT
/2HnGoOLPCzDGdeVvRNlIUTEIVJMDnBowK6yftjEFp0UdCnEsR57olvJQW1pfv72
a+8frfKBRDLEoWHLfBWhCg3rjlFtdMgYd55KOEjHtiVYP28aPpw9nhVTORDPRY8Q
FNdKINi71uCmXMPhnMgF/qXeuuXQ3l5OCJR7zl7K0ABmdJ+4nQWmy/0zjHHqhvlV
9wEfsKCm3HMTWE7C9OlyX0eee+FZbXTTzE3SclQ8ElpnB2s+uJasdJL+LKwkDFy8
Odh3FZyduSWg4RA1aZffhSd27+6K+z4tKLuX2AqaqvKC1GHWHTUVtJnssVhigUQX
73opr2QgAiIkDpyqmdPuN4La+2qg4d5EczlNpqM8KRE9cdumHHCMZ5yluJOCEK0p
xw1yHA5H5hIsLyI+DxrR3Ud/U9rzV/DHWr5zDi2C2APc+oD7WsPBDtKLKYH3GfuJ
TshqNFbha36b/tK1BubMDiKUxVVnD4uIhJPzre7n9Nw9yIA44tM/gNdKeYMuWMc9
T+xIWP1C7g5bg0C5ZG1iF8ZiRiOlTpMKkDbOiZN4k7ssI02WfCDx2C+0ZIwTAT6d
CloQ3NEp3qENFp0wLULnx9ushYvEuS7bgdUde8XCmP5zvQ7VsHVMNseq5Sk8H/MV
cUH1DG8KjzDXOwL0Uj/f9cI7vDuPPavoemvcc9bk7Pdl/pE3Futc6N2BlL9B2uup
gVCgETkZjol5M4CYyYH1WKfKaOv0pzfYy2M7ff+IBUxCMoH4b10iQdVbF8JQnkc2
1HeIMQKBncJYXJeX59935IicMfxWuAyAqqpEboWSp4uYLilwieNJ+xpvk42FV+7T
AKXqgz9djj4qJEXMQA40ZOjTl2a5WoHPkyVGI/UcpBmtsZXrn9qGLAXx9dkCSdmS
NRkk5aYp4tGFc7YbLvU2Eb4iVvMgnN7KEhe0lOrnppUeKSe+cmLyJip7DK/+r2/L
8kJxaj3YQsJfoJmxMLhvt6JIfROoMopvZi+qUt57/urVnMZOI5c7d8Z9PoB/tYiE
/Zzf86If0Ja7VKmnCI1eSHVc3vfFVu8IPGyddy7mwHxf2gpnRw48YWPrw2V2N1CJ
aiAZwpRj8O8vqzXzwxW+YuC8OyQV9hJa02kimabLzl5soV3uzZL3vzqSpmEEio0f
PNfi6CB+4q8eyfJpZWT7iL0ZSfb8GJkZFvJoUXltwByZPU4puJYxY2T/mZUFEyNY
l2N2JwC8CVRTQCMQDChRRXszCKRgvFSjuPpfHH3rd+o4+/eSIVPWCC1l3FZmLl7O
TMm8062AWXgHzU89VPlXTpHLuiySrTRe2IHIK7P+fV812ZkdxrnrbzPGOI5bq3wY
moeAz5k5RwuGz2Z3UPTcPzf4CVrSzh3H/QmXHFfFeb27VfQzAcb223IwHC2mrJTJ
TWdaPHu3NFj5DUFgUTGUgeVoWOhY6nplCfqqU9D9u0bUM1cREvN/uDU6NXUpSzGH
tiiS366UvXdmLJtbwMYdesT5JMUUO04Z/iya/ukRGycrL1zumscU/RmogdQnxM35
USh50+j42g2mOoCYLW+cgZ7MeYXt9Vd68sz1uFGjKetTPqhnnJPHTWzUfjmnGQbq
dsyWaVNM9i/lyR56EZxCYHS7nHIZ8oBVrkdICv3Sx80cTijYer3Isbo8/rdOGszR
3c64Cbt+kWAKl4+yqFIJfKuKC1l7GrrOkug8GmRswNOvfmzWiJX/sRcoFgXbpnLA
mlW18rCb5pYVBn1P5MDW6QSUVjZw8Zk53zhcFf30URZfLU3hIOg33NyaEJ8v2KD2
FhQNmurk/fZPuaXeMgoLmcZlvUSHKAkw0m1RAZMPePOssSSQHltYaNJx5V5uvyS9
ZEXdKEiw6QPARe2mkks8SyJ2IeVwMFtsZ1m518RLT4aqQ6H28T+o//2i4eimLila
iUKtO0ksBPnT747DwHir3WThmbvZoODGI873gZLc+v4G9XlRDViBD+aBddaG6voi
d/pYbM0u31Fq5EewdHxNQHXSwgzUPlj1/W4YmTiQiTUSZXWaKqh/sIN5VwEm3pyi
e1TnDxiXgq278X23ounJUmoioHKmV/t5Js5sq/TXjQlpls1pODrwubrgz3WpLuNy
sjistVaTkUhvy02/FsxNo3NSMvp83Rdg7yGEfe3vGEaTKkwgHrD5GGgs71jaagp1
GIByOeR1eUIuB/Fe6yvQxsJM16CoxQAcdZxIFKlyBVN+f5P4LauAsRh+CSTr3lIK
evhY3AU38RoYdEpU675GlfWo5D/OIR3QhIpvVVnaZk+6oNskSe/SfjOmzCseOzs3
B1ee9Ce1yKv2RojXRfiFC1r601ZYjPuhWnsgXTpnos7SbI6rP0/d4FHNM93BWaq3
8HCCEc5sSrqHdMbogSCxGkElkXKEdcoRP4gvqOVWV0fr6RUMGVXPFvsCjV63c40Y
I4HanHanHQ37pu0TfmGz7h7hpTgaQImNkBTYRIJo4x7SYRhtIvtE1ZWIH3+sZeHw
rRrHFZdYnKNfhgA99ZqBM4CUjgH9i80D7SSQ1bjhdSJiXweLnfRI1L0r+W1yCvYI
kE0zdSAPtDZlphQuojE9HM0dAljfpWbrgy+tKQ6kCjsP1DiPbFI/1rsmligGrkCV
PjLsfG+KFJ1T2YCRJjpnbg7ZqV7xqat3qu6qw2um/hYot2Ga4REwHnLeFgO6KfCG
OSBWksyHqATjMB7u/TsG/dB4wWDSCRqdSwYdhC/V/gKx1LQ86DY9q0suBgYVqTLV
Lc6RYjhS8H+holBrB1mkQPgKsuxvRH6CXlfQTwYE7HbJbhP3QXjpowQLMW/xVaJa
1T/szVbkuRUQnikTZuREWeO9G70He17RCJ1IHKBQuaLxBrUgJg/Jxyc6HbH7y+6y
BB0JVBrG06+w4gZx4lUDLZXCexityK+vdEzvY+HpFUiq/Pb2YyESnxHAi1fCuMD1
VzWlhcH0A994noY8ACYoDp61x2ZQQSWWrsaYVHCWI3NHrnxE4U7XHFPvxRSR47Z4
h4wqI4G4g5Kpbp4KqdU1glmuJwCy8bnBkSPMuRdgxR44WoYfQxmxf6yHCxVAZZlC
M6rP+gihbifNDIePlIFpWOqHFHDSbaWJzyJZO8xit+J1v/VNZ6EGz4eGcMeAf4k7
pzu8Cw8mLIfnr/qqN+YA67X0m1gQ0WcWaXOCGUT180zt82+ENyt/OPjfkqispPuN
uxere9ErjDAnrBkMYVcYZA7MX+TEC/PgseELoCSuxP/hcG4BzuvL8HE+u/FtIB2h
3nI29oEM4HhDCri6dC27lG1Vas3nvPxb0ZbGRjkm41f/HlrRga2cw7IiWkmhAzoo
HbGQoHbozaNHf3JJm/E7aGPnQFoVLtI14+ADeSDUXLHziNck+Ge5XDkninCMOZ7Q
lmOT4K05vS1F3ZImRjwV95bAZiPnEcdZRE0bRao2h4oULLa+ihuQW90n3bWaTMDM
NMdpZmjsmlut3tQlHqlsDlihBc+AMWlWr+KgCBqvKdRclqP66xyqBevamRqjNyKo
Tz1J/Jv0k/46JWu1+wjQUJyLtORPc5HHdDbK/c8J6KDIHom6rYqNjh1YrArh77h7
oMhuc24L4LIydcw9nqftPiFrl2FurlLnOVIt/5PA6eSjc0FjnGJ4A6Bm2u6BGIOi
8TzzTWLZ6t40QKwu4cndRBZtwhcyFEbDF8sOWcbtr1XaqCgR/P1CveY4UGPVYfOb
32IOEU72RlkfyEr5SpDPnD3g0Uj3aKAsg1Vp0+aLX60wQ9SvGk6p/hl4BBCEJyvy
LXW4MVi8DqHiMEqBs8rviSxsTotZSg5qg2nxu/onvnTV76OZm26yYxncAZbTUNWY
+Ym8NxdewW/+H6y8Iej8vXknKdHnhJwFrc2os+NBb8+acdWfhtB3cVotBCxpMCpf
vizCP7+ZfoRvcrSzOtNA8oFFAaluxEpgOTKLxKoNjUwMrH0XvvJHMw/lJcCR8epm
JXo7OJ1Xc86DmAyIrvdeJcw+W97ttxaMfjc9UQIz96wE/YJf03voZqwZrMiQKAFy
r5K9F3WzoiK9/49PHIXKtt5T6/RsEICmS3Suo5VsfoCkoaT5RbcR+HbxO9eilNKJ
G6aO9f7P/AInmEk1VYHfM3mxPQ4gKVJ+Mgjl8jSkGUrDeQfRl2tZW9XH0rBBU8ua
PTWtASahWXaCI++jmvKE7IU3s9DCvtuouoQ8GxkZEkFRZxPekgn07QaFL66DWFVe
MEX81nHPTCZN1bFzuvuU39G0xAX16e5IJ/IUREmD/ImNtGj6j++X9yY1aYFr0xCG
yknBSPnt7eOpBOWbNNNTTuaH1jVWvI+3CS+gKJDMfQ74JUR8HpPCwZ/pcxGENYpR
nuM1T/SuUezu3LsnRNBJi5KEgyH/5x4jGi/GfR/iybK8fQIO/a0mp6TPe2tsncTI
kGTK2ccPFhoD1ihV4tDtsU+3x5DU70wdpZkivJdBR8TPYPjO2P6TlxqUqJaeUS2/
iha0ffqEjsZUI6AiyVpkHcMr6xJF5KVjx9dN03n60d2UiyTytb9aG5+rFwpKGoU8
wy0WmCWfPAYgE2HwW9i4VeonO5+e91VJHgclXQQfdXDAGzQUjDcv6Mr7mBdoBtlT
xP1dmNvXFDSwP548LI1KD+GbAB9klihsVlYtsFaL7I5SbGhWvttO/UdRUvw6bPQ5
b3Q4NOTFLVDzcF/TW2NbUY8Z1L9azK4dB9BI7Iv14QZFjYVMV+vfi1SaZ2mO2YA3
RYlyfXADGCRCZAc8bFRrRjJ2FcOlUuM4EBcfqUSNs5z8R61ED0FvPEDWMHGPz60E
KSNavTKGN2tBg3H1KxktZKy4L5b0lrGD69uVs1gL5neQB5yK5xCuCkdePe7fVdJo
kJ3d7HQ0Mw94aL4NKECeV8fZuBQog4rd+aD/N1062IGILwRHUxx+xnRTWjrC0oH9
PlLl9KIgDbn8Qp/ET03I8SHWS853bGNQuS5qN6Xy/v5yUwsBAN5XaiRgKN5TsbsJ
ry7fnXfp98Y1lU+Za8QAoInrooYCXjIwdc0nbF1LEZ/tZjPF66JXeRZg4YiOoQn4
gf4iHt3nc2e/Hwzcps1tQkmiJ/y1tl57Q1mCBBh9Z/g6CBOjqph5fwPibiiw/7Cg
DYyxnNbKHqi/ZJg1Wh1RQK7B8F8oYrdzhiYdKIt8teGrK6k2donuNewJuYYBi7tX
+0bL46mxRFNmmnd7XDKIbi/T+d9fTNMtKCPb3WqbXIEIOZeUO5P36i2I9KRUWGsT
G5jXj+ysQMbC1EgHkNulS1tV0kORmAhMBduAaP7OalDDYryG96tNSuIVWcPCl2eH
WJPT0SYlPVcoA8wYNHoWVH+TEugbtSG2HDR6fMY9WW/SUGPNRHfiJ9PWT+8qksMW
srfQtAfKCzO5yO+u+3RUJ1isYvfxbykmF3B5k1/Na70sIHwm6MDx5DG7MYmfd/n8
OZI1cLpltPiMslY3hVkIKaPHXXQeI9dJ0rMV3h8C+NtJ0zsDz8azh79F6Z9im+DY
eevvvI1recKTOwm7ZSRAcQw88XGjbeoI8mDZIM1dM30BtgE/fthXXfoIl0tZCgm+
n8REMjOBgs2PM29JMmb3fqjOcnbqDc8oehZhse/rKkCZjcymM0jbP+5VMx5KOFuU
hbX1ixmm2Bago0DMW6lKPHc6ZRXF87gWHLo5MBC88rkxcZaWhELlYbvyJGm1S+o3
/wNGVEGUfjL5/CNzfUj9FEvPQGRBubSZ+LCEQACtBv86fQDl6O/nFFxkfra9W6rr
plbNKd+XCdC5tnE7L+Gc8lsVLmgR172/xGn8k6KX68JzLvLZBtE4ZjE817ukp/3R
w0OSxgVAn64BExGe4RgR7u+y0eJ2tgM8WHHspLUaS8xt5pMDPTwl7oGobOWTVa5T
/nXEp6P+cYYqwQi3FY8qs2/3nQzcrMPcwvlGMr0ZRYhvog7N/JgGaYu+DetghMr4
i2ICZO1znQUsDT0sB8zQGIbhQHMmMrerclMhcEqkK4YgrPxMkHaSDEtsdjrQutIS
NLHg4KrZcFzmFpZ+LSS2Y01zZ40IoNmCZ4XpnZD4J323029MbeKIBD4DhrqQUnzP
qSxioAWFDRJRb6jUDkzUH9n+SgIBPYYkKmkRId85TM3t8SnrmyCpfc/OK9YUd81f
Q1OtsZfOeL742dXw4CCA9GTmLB3TcFuYEzouS+fAnknFZ2qKEw2YhMutK9/0MTTC
4kP7opkqcjZQxdj7n9mzAus8dufjl28cglimMOtGCaDbmcOhEidGoZgItZNzCpCK
gjFdMenj85UVT0nOJr8ml+UFyCIApyAR+ObapnU4EeWnu2Sl8n5w8W45S/bK0HaH
qkeERrzkwexNKWm7rcWcqMqk3g4WduqaBDeRJd6Qb+vuyZlhjxsKRp8Emes/hlce
CQ5ooFWCnixkgjv+73IJHSZrD1wbprPtpsUJ/KOfIN43GtE6AUvJ9rrLjfAEfczc
SrFZB6zMDXbNeM0UFpRyeEnJNnLBazbBpxEcEY08lpHAJ9nM/p0R1Fmrsn/aWYC/
xgO/MnIz9CkcKH1bAdf1uACreMcaOHGcx8kzJK1+5GwDVatxu8qw37qE7owe0Lwe
0u83dZNJolZdWKkSZDJ8prQ0Un/vu4FztfkjQJNHY6ux9GrJ1R76ELqt3y59BlQv
RY4AGqh61trPzWbmF1CyNTulgnJiYsYCh9f4zSucE/8OHZXdaZaGubGht+wXMmL0
wNTNMrt4QIdFXYNnnJxoZxE5xnx2JtIpvYdsYSVZ6V/RzL2fQBwXTNHFl2T2RTbI
2W12eRC26eleGOZ2kb8y/CH3Ga2GRBbNpBBa82UdqyF6I6k25JVzc9g8BQh0I/5O
RIiXbuQXxwhCMvDGJvJPtWcwI1M1ePhdyx72DpbL1SRm+vD37UyZEPJqFUN1hM6f
iaFl4yArJEC/9nLP6JXu7vX25AK7dNdqSNF5BRD1ixNMAervMmHD3uXcnaETWLNp
hILrA9U4GuQaf9Zq9OIOkCE9xVnlklcVVPLyptr7CGShbBGyTWG2/y4pSyZzNBup
35LcHAvRGud0Ku2aUHXjDhJC7GFdy/FZNUVMUy+G7Ig5A0Brx8H1wwt1vdOTH45x
409BFUUNiZIP1iAv2vKoC8d7p81UCgKKaHNBKbY7gCob7b//5KdPv++T1LzO4SIf
sTDr7HmY165zQWq4uDKwUgINoMC0xJzVQLYi5F8XT0IvhIGAkwGPpBVBj2jAb+FT
5RIG7EW3+aGUhIsY1J8NCHz6XFlwY/povN+PRfo21W4/EU3nwR9mM7H5nU+YQ2v8
PO89kv0oyTAgd6QG4z6pCT2gYBypbfY3f0URWGpvXjLoZ38G3IZCOYFQ1Sk1OnCl
gBBbnLJqf9Hrxhfl8FW/FrXUEBzTJf81vVlSz+D6mrUQDjNs4guXbg2KgVnm3Ry6
tg3s+OgTITPUUALAn2OYZDOTSnd4oc7oUW9tGHGoC1pURkErmkVsS79d2XueRZqI
Jj3rpqrvXgVsfG7CT5JF5IJGQJyKdpkG/YGdro/U+OF5wAMJG3rckK0hKhbL0WS7
b+JAKXFkSPBFNrxqMp7Wuvgm6f61qwuIJJK/nmGn+yVGVSTQMs/pMCWPyqOgnZcB
377i55n099hJYamZnqTNlFho5ntjZrOZXJVNVBJKkQVqu1nm9o8YsQHykGNjGrkc
CryQPhbIUILrah6/ijjtUjkBQf22S62KxpJUgJ6BuxXo+fgdjLwvAdUwvH6aVrsy
+mNC/1RpJKDjoBrrk1g/fgZ7RhtXQUj3xBHsYUlr0bf4ed1GYwo9Fkv85fxvIZ3F
F67kwUFXS3Jw5U8pNNOsFi0JV/vGSvwtvepbHcO8xtD+6uCD5VXft1v31/ZwPHrc
qy35kdCnkBmUq6wwU0nYLmY9u3itKkLn5ZesAFjk1k/5xJzfh5gpgBNV7fblTjrP
D/gwvzZMPlTYuxZanJiZEqwYc9E07YrCe0/PaOEJYZqaqncjZW22T1mgvrJF6pFZ
L9YVKsxVDjUE+RL+P3CjAFgoCaSE0JVdXS0xp8GHG00NAc+XqFN9YAjSfMQcHt0D
vGgzvXjVin8lhQ++zvVHsW2yeBvNKUyXDtc7FAaRJzmOS66ruDaKo/u/KRO3FB0b
VZdlchO7wF/XjuMXxjlVVe49Zzu7EOjAv53n6ZU5nn4iO/mk3a3iBSCJ0VxCYAxq
kNAF5zab/RKGApgFMoJxWbvt+aasapIdkFyAvUJixjvrd5CEkRIOnQzqKNIEEw98
cJe9GLMGRIKfYpjJOGe7p2Y6blpx5WGZFgqr7ubluK7xPGWm4xb5cKLaLZ0lCyin
FaPUqY66JhCdMoaAkVF1gvyQaXnMVfI6d0PAeFOhfj2rUzof2RhjAsOW8JaU38IN
xZpyelS5nVTmocaAwzzGtxdmSc8IEc2DWJHeu7tQnRHaHfUoUX9Jp9OkFueho6zG
4WQSbJZFZpjYOmQVjqSfsuv6pzqIJBfe9atWxsbWuAaac/9e+3LXhWij0lt/WN3y
TEF2sySCw9/thWc/9vr+hXAG/8pXdQUW7ViO0jJpE44R7bIBaiCr1VDuOaW/+U6d
NzlYecuERjc0lRN3b+9Lly5pxq6IQUZAYb8yiy4iN45ppAKsd9L/mG2Xm1KZ5rAl
335RJVBvkaRkEygIxetkI2DSdcrveFQU1Q78smA49PCvJ8buZC4x4VIdyiCO4Tcs
m7HK8tIuSOrHtf1Qb6xw3Vz+1Q9SItfHF9Vv/An+7DW4jYhXD3Im0dxvzYlOKUkj
vmNZobQ89aVc746NlkjQlsyVO8A7EO0ih4harsWKWBdyrBScLUesV3iRs+dmcqvo
qjct3f3ochIyl9Zc+1giwdWTcgMrtbEy4PN4anqk6B/y0fN3iHLZynfOWQAv3XR/
nDWKxKJAqfSEVWhF26wyk9edW38CPS0AM5fWj3oPi0Mq3DroMoIeoRQWyrR8dqmL
azZayIXyoih4pVa/cjzRg4KpNjjTaljawHo2cL5/OqdxB25O4crNNRG54l4/r7Ma
vK1bFAj3Fukrrc10xH21zTVQgO+lMqU3ARaHWk4vVfo+9T0Unl5SswrgRXs1/2H6
owcA4oL/Dvk+fVZ4WKRIVbng4vi40vfm+FUszflo+tIPdh6Ip3Tf8hKIadRfdbu+
cZgKuaKHpcVebjTOCZbfXBlGvYPrH5P84KneNKb8zQUWLO38LnMSw3QbuCn3Muix
LiGEhOzDxpb6livewoP/BdkvU3BYe4a3u2MXMGF0G4KbxFxPxdi2vS/DXBR735PO
XqAQbxMZ5dnlZw4bGrbaPTdC0f55jinvg9pf3PaO7teMhigMZnvY53NI+EAE4Xla
0pQFlkr1IoE/04yystnHkqn5xW7WeQbEXVXkVEmfGNMLwhx/Wf6F/T6RqnmGEEtM
CYMxZFhRuPqtNNzwAYZsBxcSttN+D98s7SDxkaQeCyzp+eF29pAtvz4+sivOBmrb
DphCHTQ6bvGMT5Cd/o1Ke8YRWhdiL3hLfdYabSWEXQCWr53XuuSCuFMjvYEEzoPj
mYjMqzT27GK9PH9lcsiKCUibwrqdzxaciglPQMMQ3GC0Fm/UjK5beLxs10kZPXO2
sliUbQVv5lintk12rFn3YjDTmGsRybp+2RWGQELVa3uFV41wGjQycxrEwDwdYzoW
BacGAAY2ZMdLcSNe7S2Mk69jqCkfg3rkfUCnz1bJQoPjiWnJf1hEUCAFlmJSD30Q
5LQaMCnAUsc8y9L6OeDmEiNnM7v4Ov4dlDGs5XRGKfquyEKPJgx2WnmzlqiSf5FS
l2+lgD5oRxVxRPwk8Zr94WN9tci4D3cjqJrKSYaAnqT/hlDFHWAkqSFQ30kD0Xah
ortlS4d0Cp5zR/8y+A16a9NW9TfCQOjlEd+djH5UpOO+/sYEh2QEUJIIlG2guz1K
L8cGs4+YUBrBNDEyK+aLkI31879KMXZX/HlpTEJBjDacPojM8YQU5foy3TabmeD1
HfJpD4Wyq5EE3Dzgog8uxpLGHZfmlWgmcO3gAn/5mRuvZeECydfRVOtwhVcFYjMu
GHn0hqfhHvo042ADstPAPEgcVbCQar7iXaPL6X0NGx/SbJk4Hr3eVoAeZCpzQoZw
ol0x992Bskcwy96B4DRlpHFrydwefDZPkcDRByAUiiQmYjXlzbeTFcUxbN4sbSJt
zX34TGcrFj2qB/vsmnl2LrNXyHvMncjeDFjLn6H5cMmm4M1dssp7pAagFOx6zyMw
QRGQMTHU6JeRglh+4UzXkObDzusWSylHBl4FdUEHLqhAVXoTen/ednq/Q07ByTk7
32mk5QFQtOeSb2xMryB7veVMPsLiPIjPVD4k5R/725MXijX61d7uxKg2Br06IfNb
odkHMJhpBEl1ACyCe5BYpLwHHeLPDxaEeiyBjJ3wCY5h8+P2eaKUQ4IKKJlG91X4
bvYn+XeB70X8khBJr7RIMjLuRPT8rA3aFnkF4EAyqFUMluO9QAFb2vos0ONdpbjq
ZbXEpABgVDNM1tT+A4iegvmlqI+YNeglJBR0pC0HeSX2MYrPLHjZqpCXeDZPkoKo
Thlb3Yok8I2LpmKbJGcR06SiQYp/tey6REzh/GDzCskJJSRrBruQSudMkeGshSJG
ZhvxcXvny6fT9oJSp80eBcaLDMLjPHjR978FzUY1372KCL4pw+HiCpOKGmNza2Fk
gCIXMosuEdezG5FeRwbPIyJ5XyqaMf6fimSbPAW6s0ud84gV0nUkVI/iPcrARnj4
fvIlfiNen4zq1P7OoAbb4NgyOrOsTBEsVmFAfceTdOuOadYSp7ACp14P4JVcYt9S
s40ejtrFbbWzrxtD88IuSE3hMWEf5HqVk3RW84T+zw4D0f0eRRKwbX6X95Gop3az
1EnXv1fUyP/8FaN70XaeFtFacF496WpN8HVtLYUGpQa3388SM9FXMQj1SPhqyUUE
V6A00wXljkPrDGUICgwKdC+QTvK7XH/KyFB6KDUe4ibo6TY2zabo2/edBxXT8jwt
2BMAKGH6k2ouRrZ4Y8R9veZcRY6cZP7+bFSoC6Dcz7Fzga7RYTOXUk+ZSLnxOnwl
+rxIlOOTXBRdc+ydb08XtMGuzyd9sAqV3UcyyEK0cQPkzwNuKtrr4D2ylQM2BvBJ
MlM338jGpCQHgMC+i2OwpNdY0CFW/bd5CmA8v8F9bibr1jGBUemm0I5D81JAjIPi
W70HKUTdxXMAZG1faFdOf70E6Ju+/gKBJreRtEhspRZioFQxKVU2tlCgsYyzxN3D
ClXzn9uBXzQrz6r8kUlHS2wmY3iJgoUnSG6HilQutl3kroP0Svi1WGsQ1VnKumD1
zPYY5OZA9cpz+bj1GhkmC5kN7C37TEvGCbKyV01iLpg8PJtcLNU3ZQIF89TJ6vrA
DQTQS1zOtYi/DfKZkZhSWLq48VoONS68xZ1byBM0DOEoucRmRUp7thV19sOqCffX
xS/CRbHSPUiPFcvONz7+5V7Lik96F5kOHogbWdKA3bh2Xb91oa2lgEMyvfFjCwJb
jHSC9Pxnjos4jCQBQrNRhtPxTXiyCshFeywqoqOtBKwWY90cEBg+hRbA7tkas4f/
xTcBvPbhPRASkq1TlB4/RNawUOU7az4gdMFFmF2AjwpL5LNbp6FxNhmjoWdJpvsq
0mKfWHLa77rrTOeyLZcnnBjbBfa6POVrTFBryfN9GRhHpheafH/bWpsW2I/GW79D
IItJpvqFLv6jyBlMaxqsT9i6To7wXKlm0S5mmBPH6rbYfZSXEg1ZYiXOewkgPMfW
yn+gci/oCgEJULcvVvbQ0zqAassSRgSiPDOVmBwh6eSmBOArOK0TwCpk5UlzfFgp
6ZrpU4qOi8UETtjPXzhARTcYZ1tI0rJDIer3LrSlYE1F0Y4k1aJyDe093wZ/noIE
HGPQuMH8OizWv1tHM6K03MrSaRvAq5svFIq+CS4xutdaEORsZRexo3krfujuPKoQ
XsizRJ+elRh1pF6CV6QddXcLPDoA54xfVmatT+bZTQLbVTjrJXBrRwbL463Rfd1c
gLjwl2BsaTqzUZaI1PyN1Ord+DQ9HiuuyvbgjCRu8r4HjKN7c1Q93Q+wHZNMEZwf
/1oPF/ECblmrNN52tUnh3UopeRSFo9Ey7N2rseO3bAOo7AxarSb/yYbmVdPFqliA
RNEjLxBP/dXnh6NGX43JluHYlVvO044QFMLMb1RQ2iHzzylnYPrw0E9lwl+OkdW/
3Z57QhVqQGRHzqa2cT35IGL2DvXJ6VPcvaZBj93Jo3shtIEJvkIBK9hnN5KkGvBd
SA2FNw+MBKtPKAbWf3+5O8dd0Dr0C3EGvidK4ydxK/1Jcf7uD/4iSSS4mmAks9S9
X/SV3qX2ixoZ+z+mrC+LGLL6xLV0fTau+iCyHsLILBI7onETk+ZvQJ6YE1KAhmyk
fVet3At7A/PT56wab2HWCnIWCQDexGRouQoOuS87FduLGPf7L7IBzT0wd9+cAUa8
uSUYaXupdYesJHvje3GoZdw6OHrsgpyfKf82i9gpxTZkKI3QC2+mEPwLCXF5q9pp
pQJefFzsmH0tmwnBmFMvvbv3RJI2k4OFLUo/SjC7+JSUeRttEtpUcn0CSTMoKXK9
VGHQiJgMZVXveZ7BPKRj7ReNg+kIdym2Lpv9hpsxeDw8v/0K/+V2awKzehJChD4O
2H6iElM5xi0soY83zRGCd71JkGp0fYFoMncTrXsIdwuUcSNwNa4p6PvQ/vXFg5NY
GWUIv/69qEKTDh7AkXBTPPl3ucxZcQqxVoQq2YsnGouECE/GXRx4O+SNIlcWFqVp
zvHXWQM9QSin0fsIc7+Lysz+dKVvGs4RAOLw4jCtvgxZO63vQjVg6ZlT3LadwrhL
/JzrnpnoXlHbmNijBPhhArrEAKL+PP2q9COI+zD4c/ltc2xDmQVKjHH7V5UmBHWG
21XEJ7i5947K6bowrmXGRZN5ERRhGOVbKronvXCYCIlmTHqf1v9mHiqGLKUeAtDf
O41R7XIpehrFQydFOaQ2VLAcqjAdlkLLQd6l7P74bZVxcAG1a1NgkpusSF4vcd5O
HuMoh8SbRNxGS2+ibVye5Wr20XwrqeScCSIQ1Zj7LuUHvJn5BXny9tll6lHivAyT
EQuY2zhBlRCISxWvGZgCr+lzTvD5NS9oX8XFT9meUK2nitUZWyyYrzikW0Ajiwdd
6ybGEBtzojkmnWG6ui0Zy49JKYcnWvlpNYDtkTd0WfGTdKy1N9z9LEyUgd+t8Al0
ZMgQ1YBZ3vP+Fp7B3kzOY34ry4tdYC8a9IklNTRc/huihT/P6wyqN/o5xp6TP4tP
84xf25BcNDbALuHnaXVlBBn9vckts7q1LDN+SKCrzQC0IcRMNmNziUofsAc+Zkwm
DHMuiJ8HCvTiSd7hiqTvcl0rumTVIBFlCWBHadjSflX63PRwrKzV3qccl/MNmq+v
tshrCh9sz1TjUJIIaTZYhazvDO5eWS9sezroUbMJNq6oNbx1AaASwkAjD35H8ZV8
z5cPRalNNqH3dYFXaeSUDfBYVxjACvGI8SBvthtl0t5txnZlBYWEMvfRr8zG9Kac
pytVjs98GEYvIrvEGJ8RY0NmRgpn00l2BefgxCGsP6w0HAtmWfeMQkt65NacTdye
FnGrTZhxIpkvRYY4lcG9pJh3ZW1fpLMNg5YyRFhzRWtcBw2sNDifEz5VNZB31Ohh
/lg7q4zElguPpZwcXgiNDS5hTesPY/iNElm6UMQAgFx05DozlYlG9Tu2DoANVVuL
Kp2s2nDN9XMVB87pX5ilzyiFQLBZfh1eRkj1qEEjFp8W/bO9qAGi1cOeTcJ485wd
D95rZ3xGgTeJLK5abgrDoMHo6Q2o00zv2RS1sAqWOkZXJiLGpyZqOAUOWTANguoo
PjCN+C+0aFx4ZjmmeeTupXzbSdHkzZoJmACSHnm93OEurZxAaER64ZORfQKCpcW0
d71lV7/jMX5pBIe1yubwYNsJxUFywJRnfWtmVXdn5Wfa3s19Mq838i8bXuWs8xeY
ScwPAt742D2+oI7l4gchND8SbvykJelEdowPs2Gy+AnImHeuwLY8Ek34LQClN36A
doVnFSEBhVIVMaKMElR7UX59m8UjNr01N5q5Alb7MLaz329ISxTNGFVHZvuRUkvP
mjOJ8+4d6Ps9c+wGpDqfYZxXnR2rfBkfcf33NsKtqm8/FM/YSq0T6LnYEMMx4Pf/
Nq4MSTP+blGnHdiawBjaNXKJQhT6fGN2ZClei68zpNI97JD0ypbQxnv4QlxnbEHX
RzOU5R76dEoolgjfVEO2IS8MhemFlkc7TplX6vnmnWXN0+We3toWDkDDwE5F/Gib
s28GIeVtOpzX9BPD6vRww0hacWBpyIuRiJv4cINuAkpnjsq7U86aiZE18VrAafH2
0Sg3wWeXt7euz/CqCOugeoGXXFwWdBb7quDJQl2kzRBxQ81OD2qOP7djVmlGxlWu
3oflDbskz2oFSlGCsCxWBPILD6WnSE5BPvV01SvT6FZ32xA4syRXlUauvh4Hakho
bR4ztkrea2g6KgxQT7MWLjbyxt7GCnNxSSqcfyQhHJCroOb3wfCvKC6/keecipvc
3FxeGJt8DTAQNmszC5FlwIFAefYYaKaAcM3XIAUMcRfZMTE/RcPnl0634Qbp0/eg
bZ/TJLYUaJiGnDcVFmPCOIPweinqdE+2etcm4wI6grgnzOvb2vYDqQdOvLE67GPx
7A5TpMPKNVNDxThrwX47dAsYS3BgLN3qd5xIboCZLawkmKh7XiEcBHH2biOMyana
1H9ybfZkmaS8KyqtvxUD0CC2RlJkKR/8HiSCN4AGECXxrdwB3Tl9rNpCa0fjoPQ6
K7eqTbGTh7hoICisrbnuavqPzUqcJL38YsGO/c0i0iMF4gEOOqpEwDzhtJrFU0MM
+DLiG9vlK8fYMl70i4pWBeT/8dSVlz5J0odVd6GmpA7uwRMmCq4wSjV2uJaSlqog
qhC33mPl2VG4I4hwc4vlVD7L7SuOTnJnlUHj7kzIQUVpcTX7vTQK7Qgs3ajp+QfC
V54qsAPknFJkUxk1uX9CE/vYn2WPD3NR+F2i/y1Ap4vOr+3lgjE84PR7gvKA6rXe
as+qJhwWngTKz2vXOVnqZ7lIOTqDF31n/tjSZAkCx0UdlWhtCBCOE/661qRlJUuN
83bhxXHgnofmPcxBJS3LFXRX2MF6sEgzNfFvSL8aTKmEghSz63YvQrX1rqN66bqr
wdx3A8WSUJkqvfo2XYMqNA190Vo8Ry3H6U/L86jPahk8r7U8LqoT97tft06sSrkO
ka8IdF4LrSu6Ddu6OajJgYjbnYRiLJ65V2GhBZ8Lmml1QC3+FFIvTeIwJQG7XQuo
j0pRdDD+dAfoGzpAPKTJ3cU3Jvm+OwUbbrVIEZpGoz6MHBTJpz7QY6iCxHnSeRIR
QG5Eyals4clrgBCv0oRWbNZ/7d6fcTqTgp+2gPkFt5hx9QfCuiomY5QIHCxTreKT
YI5yZEhKoo1sGg0dETurWKfR+uy1hllfaMBWUAgMmIDDnaeiDxmHCqPPFT6760PS
3T3OdMh8rkMBfhSByWVOdFQtdumbQq7mpqgPF8j0wH6YBpjjMAIiSjrN1lKLrz5A
6NNubPsnUzO0kNJJHAYHhcEVkl28kIe+61QQ2s3N1eVeMDsA2h63Q9UFro5VAx66
Pt4VgGyUjLzRE/ZFkg/8iXL0wofSRkBXFBUI0aKYHrVKu2reSHwi+8xQBLrCTwjp
z/cxwr4e1GS1dNtEQnlkN+ybUJseumPZpBsqRvT6oxTyzJ+4VaaPTp1X+c4sTrbx
OvY7DaN/8MdXwcs/pPpR6jdlRxpkDTzwuznFuattmAHLDnleKqlrLc6daaJAljJX
dY78WxtmGKGImHZVQ6bWVvc1v9QFo2mvSQqHseNrgDApgOs0CMR68g+IDFgXkx6c
FY3LEnVRjKXLwR9+rV7yvTZwPnkR5J+dR6XNfsKy9qIOBf76dsRxcneEMpuxVm13
Ff6ApnglnkYKCoM8iColTl6JrEm1qKRf+7Z8QGtJuweJfOsBhH/FOkzxxfLBjegT
/EdJLofnvXbbNRKrTFzO6WJkuhq80iA7HJdBiR1tURSe1fFt91s9wFI6i0jUzwWD
079tkeej7jZbYFbEYW65eUOrCu5zzLzZZJAj2DMyW2r/KFQ+AAFYCYqHa/Gtqqu7
7PtQoMmeBKcewLiw/wNAhQ3UyDpoFM9vyWx8XbA7w1znCLVMhhjnhO8nDsKq7w/3
P8h++zqE+9bdNqFID4IAa9P5CNt2Hqmgjomn5NX+ar30+0q0XAZObrI8+0idAUVp
1rDilT8Yl/z6xEIFPRWqLTxz7jiaSf9CawA6fHWgt3bGr8IBJjULIi8rLkZ6ByMq
OJ2xr6+7wQt1R2+XT0J0u4A4wXPa77ZXskZtqqz8yQo3ls3iHyXtLoupqlQCr8MU
acgx5OOrY6dLAY7TLMsrvxcT9Ey5vXxhGH5rHnNh7cv8Jp+fTJJcs+5BElKI30RF
5HeOgNFg1bIbfZeaA7Ebbz6Yx1tYe3YjACdiqnx+eeHUBC5SubhWyJGn88X0lSpj
kST0eW+cPv1+vHsYxo/VAUUOj1Rn26iesvpObIJhxsSPqOVGv3GUXUmRSJNZZ8nV
LiJuMSq8mUk9C/904TNQwsXh5VGDhRs5IEYkgMnIf3F1YhfRMkQnV0LASFtbUZy0
8giceYg3Rq230UIX2LGTpEECW0ZMID1dgGxTWKhIyMZ2VL44A+VygJpjrWARMj75
SZ5KA9t6gO77IylbvoqxgCVm4n46EOW0Y97SXNDPFHz9OAh7ljvwaH8SYAuP90rF
iwnj1CM8Fjs1kAbs0pNwi+3bvmm2H2+fLFJkVFMBtmvQ6UN2HBu4ZR9twRmpjolf
Bpf6a2jPfsT1HKFUfCSG8cQOKREgn6jZz6p9y2D/BgJwjE+DxYxf9vV46xBxjWMm
0I12cFA9NvNXZDl7ovKHDzkTSAOvy4t/1GJ8XA/EQcBkB7HN+HE5YINeQqOSAYnO
B5eNA/hP5IyTRzI7ZF95ovR6K1CWidmNuJPCw5s+TcJVTWvA2uXAPzxeEtmnhkzd
Fn/J5uSee9o54zVmjUwij6XUVodYcgRZPr/id8S6vRTzuk+cro3uf+KU6l8UWPXZ
mvqLU1F8/xqMZHf9206gauAm+jTwFl88XpHYa7FCSjyWCT1crUXy7inHHQkOswxL
GCf3u89BGZ/0gjK5IvJk32HEeVcx82gz1o3tv8SmyDyuDEbamvLldfrTFska93Se
+CgfnrV/WE/Cx+pqXmQDZveYtAtx8vImLCIuk03jPnXDxRHBZw8el7tHsS915llg
SFOEIOrlaDGx5udFBHdDfxsg87YRGP0032axRcxWqXz14jC6FL7hXWs32GTAygR6
ZCGQdfjwhGQMexVL78guE2eZ4igadKdwiYHPsVcSyglftw192YxI2EsodCv1DxK+
oWlI/NX6ru2PLC/Kn1TGBCcD48xTGUwy69Jeu8gkWi6YplMe0oMHV4mgYQnbTA2f
81U+wpBE2yNcFs+Esa7YplZfnJf5tl3+zQgwL1jku35j1Ti8/Luu7E2kUpOmIDHW
PSK3MijfW5o5HPO+XXiQVJUgR7iia8durKfyiCJakiA2eyuFjcuLHYUI/cYI2WTl
Fn7mMQyAojgbaEBR+MtxK9N8iV6nWFn0aa5481my+QeXAgO5HXH4l0c4XTLTnITj
YinO4g8WV4PVHWAOtIRsuHAQOcolPx4Vk7EFgljqmhCzpzAz/MT5WkkKt3xjj3/6
SQ6D1z49WspL4elVJE190O/kc7rQ2Vwd6g5Qgz4DbjkVnqGVSA0D35oo2O419KoZ
FxUWGXD/5E/2DDPzmtG3wURZRYKSyDS9/ke8QGhBxU2nmG0XXv1mkb3VnmGe2pxC
8M0Xr9gOHy0MtLp94YLsfUaYpKdRRXFkZQkJAT9s7DLcGGloP60lr0R00QGHBsM+
JjA93najrkZ8OhKeroYmebiobTGhBMbcDxdjoZQb88WAqDwVFDmgmatjSP71ffXC
UuzEHvc1AHVEc66eVGqYArjHbci0QwbSsl9Jj2LDT/ywCojVHjxsazql5STGdZeT
5SMeqhdSB1LBktfoz3YTGmpnl7K9wby3CKe7yTzAcgpgrIJWM0JWChSwLzNa8A2k
mqA/vqEt8e0yrl7nq98hCqU+qRkzVPBgvh0LDiamyiZGuUblL/z41gGBXxU2r3zr
lxHPxIWI6n2IFNmh5Si83sTalNZP38qI/20Hax/J0w3+xh25DqDDPVcpsF2efn1n
ssWVtuZoXG4CjcXL+hoojLYcbPWhCP9evVyRrySXZbpt7i7xqB+Jy9D1bgncTyKw
95mn0kpMa2i651X++q2PzhCtRlZ+h0lU4nEBQCz7v/akhxnY/3jy8k3FOEZ6Rdrm
4hktfZt8SIe+oNaNVa5KcAHObf5Vnyno+lGfvGbOaCmrLwCbJKV0/m8ooQS/MKdP
PM8RctSQvoeMwLhBrWhr2yxiikrLl87zRVI2aBI/ivDVrW1rq6Y7CbQCijktUQH3
tLGreab3PHiV3AAY/kgGtM87hqPGH5bat+MpsIVHK+kDb70661jk8Q1364W5fRuA
UBX9ITmeJK0JLy1izKAOReWfAt0ibP1xMN3MEQ5hyuKod0m3nqsb/LNkCfp4ADd4
KDhe/DNk4z5eb3RolA068DsTtZ6xtRgyjTCZuu4M57KK0EHDy6j/XCGslThPKo3+
HNXoKq447ytOfGh0G/JILtkq+1SBE8bw5LwMdldd15vZ8T/kHp4FhM9y/5BZdbfl
vBygDyocg68rxiufh/4bP13jrXQyYl5/O2lOMNP9Ga4Hs26lN/o4eXkOsyqljf9G
OsqNTcrMq5xvT9ntjqDI/22U4lx/gByduApOOi3AJT3uSE9bAOCh7LHpyGJOOjVY
Ykd9vxVCMWFE4KiXuvE3x4QXg1ZK296gSH53Gg7AnJIxGf8GJoh+NFBqoTkCO8OD
8Ssxj9XAV9Bln/aboQPUk8NMyBMLVKR5+fuvpPFmXoSQdupbiUJ6l1TBshb1d1T9
e6uVr+97DwIOTU7uaYGaHnvJ8EU1WMTfa4NHzYT7kl6AJcjtxKT+MiRlkRdgGbdo
AgudLWirM/Y+gIm6xrzyD3rXwO7xC/gqIBC6YiuOGd93q1O5wu6QI3YbITGq1QHG
msoVc0rRLDUM6xXcGKLSm0hvH0/hDHaJHjMMzJJBJ4opeisZOv9h+WK7A3VdCWTT
6qn3chAOJsIIosI9zATcW4tcd+SEqVIRtw46VELrhgGHIT/zoXMaDn6Bkk4BlX3J
CP+oQdYxGm9QRp5iyEgqefnz1ydqsGIu880SSu2SpDxoqxLieiSf9Dc6xbRb/njc
bvBUPw1CvdfncB55umG20FTQNjAElGRrt3LwbDYsMAWV/Jv7RDzcSZPOvMUKogBQ
QRD+jprdLD/ABh8W+HIUxCEz5NSjzsvyCpx3DwGkq3z2qtI+OPazTOqPA1ROlnV0
h+8bYnttJDPj94ZvOHKeDd7l3FtgSosrHKJwWAxtXTYUSXxRvOHMcrb5xdXpvSm5
AXJnSwpIV92h3Ve95+unchz7mBGjZx116foU2lApfbeUHp/zZMC6Nzgis9vmyUSX
HDrdUbiBkEDE3ZUyci1TYGiScklPmPRgcelH5ZmffcHLlnz8NzI+77E1HY0nGyxX
oHf8oKIlamMaAWmlAD0T0JpRxsh2X9rOOf0frOpxq60BAy+GHke3wqaKmsKqPk93
fBUDpTgjKrlVgoOR/9ezEMMOnzqS7rID2Uqu/8sHCjcFkA4aNDmDZ9YJarZkMfya
/zFe8F/vVq8zkuP6QaxOxV7UxZvwScWCIUGGI1u1Ndpa9s4Kve9z3qXprTtK3KLg
+XTWuIAMC+rn8RXJZ3KSCBFvApcpi4Hyssg1I1sqsvfcwaPcAMUXdcNN5Wt55HzX
dpEyFUy1jtkGVid6I/a0xaUa2J7YYtWfWdPTz7cNCRtnMyfxmMK8AOfI8W50YaiS
P9i2D38BnaK86u6zfR2uNRqWZEXvm63g0uGrfNTi67fNMOusK2dDwq1qKioR6H8Y
ZuXt21vCTDNUWFdXnAkJOpmEj14yAD+T/SIJqW6VCtgd/EpJubPfTsER+BmE/Din
6UWi3aK4h8coyQkFJFAwFuLbUqG3hdikhaGL7Y2FJLKDXiTZVIaNoi2Lx4fJ6dEr
vJ7VDXKDmXQOzDfQGbPtdXBpjd4NZEgR02PymQn6bsZLnw4MbwOF1fWucqCWzsGi
rEhGFj2PgfcISlVtjb2fb1eym3fPif+zYMCPrYgkYPQqJsRDNFynWwXqVP2ahEVz
K2lIVYzDOXppaQPAPRwIeBAsVTwfiUoyIv8zQiM0L7DRHKLt7mRWmDH48JHWGT7p
L8om0z5u/XkSIgt7ti0A6D/WXkk2zHQyyOwlwZrYdYTQqTFG6Ft05J7fATHP3V+q
fz1jj2EK+Tgrm605q/AQbbWtAc4bVnK9ZOoLejhZyGi1NB/FqEaNzaPgt0tl+ffm
KWIniYIhcNLoIAHCKGnIkIFvXZwdv3rAUQ5M+CAV2VMV3w/S3Wdjcwcz0EwY0pRy
ALpbBw3V4IH+3IVs0rabKXGZO8FPfhtnZGYrUcv6j2qB5aQtCklFB5bBTuq+vwS3
E48Vc3oFoS+vDZ6n8iZ92/aFqoTKUYaYZsof09shH1eehg49eTg2OufAckp8KGWg
cF81ShDzOh06fCyV8nxkL00YcGFJ8br7GWdKcncuJMRwqilvwHVpzstKKZ2oo/3T
+jtba5DuY1P9OSvEa4KzlLzXrM/e1hWgdjcbh4ORi+PRkSYVKOCQfl+AH1ZJdBHN
u+9+rzlrzjebPH+ckTofKyZe4/JfYZ1RRDityyjBRVA77HpnbmSSPdqi6hWHbtoh
CE6Cm5/fvNJs0x6a7dVhoIrcUdqu9v8br/DF/8TsMRf4/OYyKgzqfVLKfIBlfDXs
hD/sDFaV6JwWUIrfFMrvA0pOJq3J9tck5vEmW46XVvK1s3fwmAo5Nkyz3ByyaZTM
XhcwDERa7mUyY2DTLHsUG16Z4EIKwPgE7F36hgSMy8egZdusirmIkOpg6Fyhjhuh
e/STj4i2kOSpL11czielVPnCs9awa4PJQiGonJOfggzvV0RedRm7Tm4xQXzkNqRn
OZL+cZMfkDW7Vd14FR3UbkGw0NCsR24ORz2ACua6SJWwNl6r5Pt1Ivx1hSy5BdOj
5yzU/y6k1YirI+tkYlon8DbvXAFzOHZTYIry0wnnSuHnNj6YE5E63s9LNaycMfOs
PaAwjc2VIxyYItHGOf5VVNi30LFolHaH0LAt0bi7M+ppwnWjYk2ljcVaNwLdWz0l
6sTX/TSGSw37Z0estAeheAiGyWBjs3lCFWDnVNN1PjfOvVCZvChz4Zy7T3OSdxlT
8Qy+ZlGiaH+SWHKBSv3oFm3qZDB8IpQbd+jDbGobNEmWn/ugb4V2iwYG5DJSqScJ
6LVrIGRsnEB2HEqcSdBFbesapcxRg0Be7IZCy7y/ZhJwYSUWqT9rufrsh9FqgK/g
f6NPwxWWPVqjBYLt5uSvieydH2boWmBDSuIuX7izKdYLRtEoA+qQxzQmdmWDbqeo
fDTJCu7S46Ou3Vq+GbNhvioQTVMcTRqVbC3v7yD+TE/1zosUpXimIqMWRqQTMIPJ
+hkUtp3GvQ4e6DOOnllls/oonLeZkio3+Nyjt5AfFxf1kf1u4mCcSU/1qkeKIFrK
qPYNesX+pVw5s+4EzQkv7W6HbZf+9n2CeM7q08O0JtZrmqaSrxTYyo9U842amoF1
TNH9lJihHF/aa3kra9VbDcYOUueaZqs6UExCyLKH0ZSav7wGuIuccD195i8AwbBr
+3cxRwQKLWbupwd2AlAzkwbxzHdfkGef+Pg96eL+kTbyNa2VfSEREjUztlTlkgIc
68umRns9qP7wFcADSOgnrx4yPBjPbcsPFbVAWs32m0Iyi+cQuxxAv/5eTBz1qcYn
r4wFkhrNbauFCLOubbDDtaFQeGuRBGIAWuycCM8lLbcUW+jk6S36e9+BYevubn1G
wqE4T/Crk709BeK1yEz9kLY3t7YBTF1CFoXexLOgGpx8bnYSL/544SjV9TJUMDWo
K/vrkEscVlxTen8qPQbRBoMX5vQLD/ewUqK3U9k5HSAAuq6VgUy+Hjjd5rUDZzZJ
h+cgYgSc6ItQwhZkX41pD41yvxkeos+Ul1IsJmNFtz6Tf+sOqyMJhRMtc+AOnl0b
n47JuCdq6JCKnAf74N9riRXoVBwWOCixblteGdAJXyKKX1ZYtSVxTBHmiM8Hcvba
s8frsjz/Thv9Br4YXKRoXKIMjdZsgNubtLnFg9JaeQYRnEWfEhO62Qvgq5LR/Lwb
MEr+Bp/5sy2+7br00CCPScB6MdAm8Ty7SPgmvaF3DoZo2SnQDuUWCAbhuuDct+9s
LfYYKsfh4qBeLPHEua2qsseNJvEgaNo5I0ZfeIjG9ANcrHMYntfklbDCTfQnaV4o
YBtv2T2n7WzIvGwkb2H1dnM5X6JES9yejuBE1qfZ77fAjmAE8Yvbo+W82F4bihDN
/Xnl5H2vGtLpT8f1BIQ+GYRS8XYnzh3RHalO8juVNHhxV4I8ofp1UoN/0G1DePH5
Vq2kDDc/fJ7BfimQKYdWbFxlZPnWqljupUNn7e/Cl/lnNguyjVHBvB7Rkw/tljXP
K/UY16sTTOAVp47evHDrcwXx8oOFU1DnuDsZPWGnv4Gbp3osk+c+PYm/hQIqkJmx
gp1RJuGqalV4il7Fdgb09zt+BLtMTBm1LbNfcSZjCL4fTue6vguWBqYMFzydft3y
bT8fghHLH8e45askTKV0JtEizaF5FVFHeoYqgHgbWgZiyV4R/4xCSCpjdoElL22h
YKUiM6sykjlm5dVZ9fnxB7Tcsmp+Ch7z1gQprKcQ5QTTzWgcwCTQjplrZUNy3HIa
Z4bysieGNXntVbRmtvJGICG7ZeWUGZ84C103LXdYwrD0LGik1M7wbmFdoMDmauZd
zMsz+/nECDf30HRvNJPUdWZwhBNnxxvGNl41bhDXhmhakmA5ChrImTPj2jH4EA0b
s0DI4HIajXXE3lws+oecyIrkhjNtvPMOoxL9yK2KbFiA49vRbvq9BkpZej4INP7e
0tUOOJNODU6XRJjQJJOKX6TOfkKfE1yT+gY4gm47DethxlmRDUTKTWwV6gKPiuyc
FyNbcDA4HcTMKoPGAavpdRFeIv1J8T+RZZrKyFeWHtQbZa8/uqh0+U9M2AC4MqFu
8efp4siVcjDQC8w7hPAyBtc+if/Bo1u54HfNpdtJiw0h6pgMy1BcJQzcB1T1JOhy
iEOTRklwLkzzGPv2C1aGhX+DfoB4M3c0b88ZDtyPALJMCMG/pV1EGS8Ihm95F0tT
L/soAEHt6T3q9wIDopOhOj+7OrLJxZKMnyLMdmF9QHjx0UEIFINq7bktunJf77lU
NyHN62lJ5RDg9vgx0bgue2nBuLnxaL+7mYVxTi1lZSwpuTFFZoCPmtAhQPmLnLjc
cNAJXSmFx8bdsSasHpkbqooUa6fJba2h7F1wJZmmiYqs4wfruUj98PvPqqUfLWxQ
1ruvg0CZHKUYkV9LeReFbFYzi7QaBNESl2UMIifNB5d8FMQ3aOUO8CYLRcJZwInV
zugSgxFyJJ0w2oOU2BAoOIe836QUsxafyqR7bfp7Q6VwkeZqQ4ujtNQe41StkPlk
hwFS0FXMIy7u3jqfe9Pfi4Xv71tY9SV533/O8BzqA+bW2sD8s5y9r5J0B0Y5v0fH
zQ0pttirqUfbVcdANJ1kHlPE8jiKMzB4JZYuKFRi4IomkEnuecAAgvOR/Aix7u7Z
WprAiBe+CNQ7ku1nUoDkNJfvJTF4EI/cd1B9bU3dOYEdkYD3Tvz29fygOE2TZuO/
sA6mEK6apzcaB6RVBj9iCqLXcCEKXfEc3zwY1hhwkKeux66dGovo78FD4XzK5/n0
knTKubP6owoEPD+wdQ1OY8qmYlVhlpkZFF3e1Pe/SCSQshZC1OKBSzZPEVMnupER
rjQc/+NHVPdlaaveu5vgDOPXsRaEyF0osIKjGeGrB9LpJn+U+UMqok+oh1E/OrK9
crstDi1B+Fn0SkxPLZC3leKnVN9g5HCUnoT+GbLLYFSl8D3sARyFHtaoSY/GseHM
6SwxDjVIbwcfGlu9+06dSKQCQWNaBPejvzXz45EJjxM3HXUHNAwrNA1oGk68tsoR
ZqsY84TWR4Tecmeogs/oRezin6ITT/j0zS+NbPE6ALwAD7sY+AWFPf+t3fX6pHI1
igj+xTrX3K0OSk9PReQnRwjOdRLG8Q3kcDP0YSTsP6qwX21zXTnDEyTogWEm85Qd
kXV5OfmwoppCoLCw0g30uluqFMwROeSBsMpVOVA2RXsZT9v2XyBeFk3Qx8AXjVf2
2g4iD5WaXskd7U1ZYosHv84ceKTGYpQZg0+Xxio+Cwk/YqlZ/pRLJzl43jhOgp1w
1X5L5tAu+AFhBgfzqjYN+SuvJAvW725jnQYa6im3XG9j6i9aML68C9lF6mYltrlJ
34uYqTgqbtpa5Eh7CgXvl9PVU2nPQyfLnajXE4bWw/D8+JOArxUIb/fEeFIFAVqI
tCP4oGa5DSK2vJJrLpu+c3gMwNdzLJxIRfBaBnpQmvV05l9DfF0lekiUcw5C/ouE
+2i2wticeY0gVBgchVIzUdecc6ggd9K7QABS37/Ln/VW/b21VQHSdjXaBQNBj0fA
+Hy+ExU52NQa8ONIJV63kLD6Sjl4x5KlOE8PBI2D76GCMPk3rPZgVXhhy8d4pbgQ
kHpeRCuF40idOt1fOHnxRg6rP9QiLrAyF8tD/2m8qYmxRSi0L26kAtl0IYmML68c
biZILsekLEaABlhEN7FUzQN7KdIO22XiPNCXIASXF5oRf7KxxhsGxbLkMnDXrZYr
3r3WyoMU0JcmoP65F2/Z9e6mWrMpvnvXICoGrjFsAH7aXMsJJNRV98G/cfl664JC
ABg1XZruMSYKjYlMDO/bBYqFSY4n+Ix+mQHgYKc5cd+IKqJyiqkvKRvJmqAzIC/q
0jHhLjl5t3/lN3QNdeBwkQ8wq7AzAmOFILX09ln1xTJeSk+gQHiyKWIcXWYnmEOb
1RH9Clb2n2slR6+Tq7LQ9phIHgu2HuajNCO/iWkV3ospPTXW4lydnAl+TxECNlOF
gwvjoSjrOgAqAMogjhIPVrqRpAadyuL6WPuRRBtWSspohZWGkpvH5529JG3IY7nP
rbjQEmTxjDEn2IK6+po5GUlm4s+U+lbXBiLpQXOTafIo0VOexhlEUqeGGVHt1ZHZ
JXh6opGDJqv5e1cRtFChuGW49rjvo5ON3aW9MKAqN0NH+PsN1nfMqHe2++Pt50/M
kLkq3jrxaZTaSD6kquIzve3RN1+Nf5SUCZI2VJ6w7yzpdITN5T43r4WwT2EESX1r
d+aoSgfsjXZXqCx/6PwoU9lE0ZTU5T565pB7IV9EgF5bBiudDJx6QIvD2T2ZI+wd
zxxk3si0LLZ1wWwZmysg9YiyBMNGUxWzRi0JOrkSI0QzJhvjoNpUK6DJQD9yeCM+
LJvIbErMndC7UEgtV3YoYL7xOjgpi4OS5RdkDe3/7s/6F/aX7TfhORfMGUm3tn99
dKNqfCETKJNkem5eb8xfSsDZ1eBY9RgbfPhXdCwDv6uYcKPeTHUVRDf3pVB3/1dP
8nMzec8CUB44jfv8DmuuQ0SDUFyZhzodLpMyVkW2cV0wcv2F95ZENbcE6RXskhNk
2lYhIHfb3opgJLBJ2P1X9CpR/57SlmNvb8+3uaZ0INuaGqlAPC7iIJD2u+2/4Vb1
Z3mQpqJf+vn9zlDX1BXicmnLrBBO6GkC4oD0JLt2Yy3ozJU8KARdUZ4p/HcXJ96K
u5VuJaEfxIzNh/VORr751dfbyUjFEObhFzjCX6TOecs/EXtMVkBxLV3ybyt82Wlc
zg3+0Tm0OVGiFsJhWLeloY0YE0nRh5ITLJ048faNjdgU6G1ljAa/iVR5iYmclaDQ
gEQczPrQHeUYArZMbybQ/AuPrCnox1o24iffi4SDPy0EsiwF61AAozWcwUYSDWvS
/6CXXFaYudFMlaQb+JU7jjGe+kayhW7KDppMl3VJkRvw7B4bYptAkRy/7WZSgWkD
i9nZGieJJZ177ACh4t6jMlaJOX74ae6BrBT1vNb+ylplObEfRGLUZGYWtjSc8cyK
08znYd0srk8krJ7z2kXVeZ300ZNOWlqMBVSRLWFRGyJ0L1ilBubdev4rbM5lO0h7
fRIgWG+KfNZH9N3y91B9HQHuc8w0iF1bLwd9DtC+GFp1ufHESCfy7SvoL+vZ1iIM
pX9eP7vlCEYHGw9ctYhc23STrz1ICXhIbFW3rCRHdSiCsRTyAm9KIYHUAAj8+3wd
z43anDx3qTUfV4/6g24UKrprsfS8/HZ6Cx+f+3mNyIglcBFKeDZZgwy7T55eXgCr
VQFm/R6hzFiCPaWccxRMUA+HPV0GP32LfW6HuOdd/f6GqccmL+8bssm7ZJejon8K
2UaKgj5EtnUMnyO2Cpsc9c2guY3xZjbMziIVTNP+kSDBTSY49AXD6AoO1Ogz8yMb
8QPA4z00Z0kIGHS7zDUo6b0a+myow/MtbCXjqwJKNJao5/gjV6fpqiPYyXbaEeEY
kpmnOArFAW0n7pBXGJWeJokLY4BaMjZi5ReTE9vlaM06mVo2F6QdO7ZJWQTNd/rX
rbOD/DUNNF50ywre7s837WYdJAxRYAxdoJDqXzYNfL9WLpTgbCVwRpZClri0xmoG
y1dAzwIZvfyPi92P9SK9WDIr9F58/I4+AnyfMLJ7WLn3kbyAF5W58ZjcWV4A1IAd
mYLJdOuh8/oJgmI2G5TMEvfTsSAk2frp5os2j+qwYcGZgSyn1vLc5bHtMMFWKQ9o
zClOv0FCquoQVik0pCRsSEbZiBlKY0DptdKRuFFGNf2IhQAzpZKyIS+5TCboslSq
B1P110U3rK+Ls67iuSljO2iP/WGn5+5dZODjTvGFTyme3E84aFApFnez6JzLLxaR
dEhpgUkk5Yy+5gLSWjcy/h6rCoXr9lFtVS9cO91nXO5w10u80kltT9DKeyVj3VGE
1V8hkakioTkesuc82DVseRV/XfB3ZA/1zxDR/r2sl5Cmc85dDU1ynrLzl9Kqk+m+
S+DUP11CREQc0HttQ5oUYRwa3W1gWYcapR+Y/KAEvV5Tm3GPy9O19Ok+zVk06jOL
8TZvC7c4hL33IkFEh3XUdVIoFZOwOAWj6YtwsAYi7l1uFotLUjZXEb1MCAbviMxe
nkX4961sPCKShk5pbFoVXdHX+oJuxiS1Kj7akkBvorCIaaSSkRLLHctB4K1RAmki
eorLQoea1QnITsP268wAJfcMt/hunY5sLZZT6gy5OIGQtMj58LNPaCqmdY5d3rJG
0hejjz6u3sn7tqG5NQLo9n2pA0IaYIP8ATkiSFV7pF3TqUTweLRI3gOZGGBCEVP2
9E2Rsp72DyBPqvmcPEkONMrhZs2Gx1yqxyXuP8Hb0Zg0vvj83ry8/0pLZZGQnQBD
YnUsy/fsc/2WidxqdK6TOpJZm3bYxbdcZzuVhpQQQUIMD89JGTWl/OyHLbQ0O5BE
HqJRU2+BPeNPxqx6VrLwTkfiZo06s1cainwg+Yc4UyHuqy8vV30t6DohBJcx8/+R
06xVd+BN139pVHowl/G1l4QLPv5KQa1DyC5BjecaDLBRNM0bkTHyEo0aWZQdwZ/N
GZcu7tOkxN09bPZJTE0VqtoKNjMSAnapNmKd98y7fVcaxtO3UovQYxMx7/jVAnZf
BbROU2Vs8JgVtcnl7cnBn/gZHnT4FYZSQxIFT52+XtIfGVSFKj2AblFjjLzOzDeF
ynYCzKhB674kvojt8IsYbWRm+a/obyiJAh9Zod0kmMnSn2ji1Hh4e+O8o609qV4J
RFubyCAvHIKc2oZSPnQ3/hssiWQWpuYRDZ447oCAS+eikn0E8h4sZG4w1fRlAW0A
bAHkz6kMXqBSVQo5Haqy2PgyOmZSizd/6f/GnUQNtQKSVhLx37jwcmO2KbAJKiJo
fZ0DVzpmzFK49HO45xG68EJ6UIH2RPKUIIsTvcfeidzj+XDD6618dLMzTuDgxJ6D
4KCfSHYPJtYwYKrEzDZPjq3Rd6Bn6X9UyauaqnZG2IRVqXLyuHxR9XvEoleO1koQ
FGoDZLec7gFf27qfuEZkpNC4Mvre1ViAHL3TGZiKmTLsBF2qX10mY0t4E3vmDS8w
waLLHu0GfFNX68JPa6nWIAemtDot2Y2pcp3LDGWatijxOCcCMeiBMxhltZMjAfBd
CVQYlTpI3AHI1lsdD6INV4DyDvUdXtYDE5bG341RHgnSjPeIYTbE5aOV0iInDOVF
32aKaF8bKDDArcknLXD4/l3mDxcQctLcOazRqkhjfX0zsIGbLoKjrf2AbT8rqChp
bRF8QEEY9Cc9OytUJ02rqQuY66dkqliSjENMSSZSUQ3vYzB7IQ2ajV8HYMDy4n5f
KrZZk2DHe782et1j/5EQz7tk1tDbHLXL1PeWP32Ai+cpEc63Crei+Drm9c4srw3d
MDm8F7f0c1FEV96XZPqGMXw2WXfgbmt97osVDGwZ5xefmonuKv4L29+GQLtNN8k5
aHjbF/TlD9+xM9OlQjqqfyd8HIBrmacDS8pcxnJzTk9bTpZc1IK219IkTxPsu/JA
ywuZBE41fcUvXpUyI9se9a/R/fgrVdHSi5T3iPAGyIbjOgPAxlAw+FLcOKW+HKzb
dKhbFNta0cZHhbsVsKjvWGEQoBBXqXjT6L6vOz46Q+sGvKaT5vSzedbDdt5FNMxR
KAb8RVCqbdJPNw6zmp5y9TcIwMdgf2XP7X3lNsYf6aFXiWFXs+9vsJmacBrB5u3I
AiImqgz0GmoL1HaHN8ZVBpOOVnc6dEjxcc3oUo5n7S9bs167NJvo4qFksTdOIcI5
TGcg4U3pH8q6MiWVqQfzwTXXO/lJ3PupOR5OcpoXFP2lvZEI2Wqe7Q3hsAVCMWN1
yUxLSZFn/3fPUlLh8e0zPqqKi/eQ/IGCuNizy8fgqekpwO/QO/vWeJ7/Is/rItFn
uQMEhmu+rWttxcTTi/4v5BA9p1LH3fu2P/VJ/V8vvDvJikmyp88w4aLrfifWQsSB
hHzIMDwaFHYEIz2rozmBijxraHouBOc+3RQEqkS7zDVw5uNQx0auyZAyjEWzpgym
rYBqYDAE7w1YFn2QPxSkzx3xhXzVZHhCp2tG8H/661MdZ9yFota8u0IOjTBMvODl
eLojjnVdSKhfkmSAE6FCkEj93UGHni5QL9PeZO2qJoafJjNEVNRF1eIKS7SxfirD
64U8koEOZu8JH6h3KtmSR8gkdiYsTJxncYKo1+7CTsEsXyAcguUaEMLOqE4HTTsU
p0jUWbwxRvs5PcM5wvYhgTaXSENgrk2Sn4MP9Vgwv5bx2iA5oNpIjKMUwOIPdxMO
XFVxkco8bwqdsLJcCw6wtN7rrTO5x4FelPAw1Ln2uMbB7bqvc52BBp98+T5Y7vzD
h7nDzJIqK9ew8L1KG+tig24PqXrXCSjRKL99pl/uv3od4PfMVvM69UNdL29JE4t1
/7aSCntDNUFwNO1nHFT1SgTZaHpSZ7TlnNElpVDsc3n84vCckPL/jiOJ93TnYHKY
+AhvVIpDY8kcsObYGQu9UNKuEH4P5vSsY0/8ltv5vXZh0+SBsOkvAdLXnlXJxXpg
jZFVoSSzRpZeO23+PnlII6VucXITTCKAdqmcjOdp7CXEDrIe1mf8DBvy1M+bhrn4
TnG6s9QDV28FiHn24GB7ZIpOADV3+hsqg8ffVl1nq4sgy5R4qXN/yDsoL1L5Uf4q
bIxqMVJXpyQMlXCiUdTV0QWCzkYqSkpVuvuf/2uza6bGVymrnXsjTjjxjVzilXwI
5mnoTIMu+E+HifKQk8eX62i7U9o8MRslQs32sdjDJivKPgsFFK6Yu7Erd3sUjwhv
95WRJNIp0Rg833sy2/GtBkBjkHHqlI7MrCZnp4zLUp9c/bZec8MnsGKF/pZW6rZQ
S1tkL6KL1rPTAbKGNd993N251hPyzlIQfGu0oG/IJDZ7m39D/Z2BLtrD+VM2KXEm
R6vYKcstZC+VVFfiZ2ZrTxG2QN0y2mtGKv5UOA9rh9BQkVhMV3dfr6ya5lF+9N5P
iQw3Y6RQHdJTtPoxs8j+9EABoceaGnLVq3CUj97Hfhk6H496J3xB88TYyuhvWIYd
GrWB6mjqzsLNXyb7E0PbyHMCqZeEaF3LHVqvDgJy/ccq1HHbE26cHl7W6Jl7sfp0
NXPIFm7MIyRkzbMqRkNhW48f2ajMrvw15wuPa/F9y3VcEHMNq1GLrLOgyyTd/i73
f3d59RhTSyjed0+oXAsajxHu+TLMt3m2YF+J0i1uoRMYVDOeuQyjpDPp/Kmvsyg/
W/D7MW81QkL0xty6/ytBtzeyj8hwMhDZEx9O0YMZbDVkglhJ5VsGTAxwMyXgvGjH
T2HS6G8H8yHnpMaWUMIcB2QuzLupyijhwgC0hW5HzdVUUC1OGYstJIWn3eiP+T/2
3uSyTCzNrnC3+Q7ZBjiILAtzJ71lsqiYt3KJybP6b9miY/375f6b7eLgWC+3qPlV
Jzz/Sm8ABkE+dOuzSosGMB6n9Cr4FVkOPx4qGHfQpsPHQ6TJfQ/eH86PeF1Ux6BK
njSXbXgsCkUUvreWqP5w/WmRCqYhjXX4+wJ0BdVslEjhDInURziGsPgQ7I4g5LVP
f2ng1VNJMHb+B1Li40kXqxUXcgzbe1zhhHSqElDqBtaOAbSXz9rN0afx99YPbqke
AW2iVykvRfGZNV5/xPZeU9Hy6w5ihn0+JYC9ZYvHVLxhQufzW+Fo4ug1mxc0m2O8
Ez/nj3AOhvt2Rzq5/xLrlS5qeUSHAbr1BOfHyN1FNc5Bxr1tiNJ2uvrvJuYaqzRm
P60JJAIc2N/UHsu67KEot987MdbiO7YK8aIo8dSlYnCPYwmI3Ad3kn0DrlN98SEU
duoJyCBVPeJ6UESFQgrQxUVGh7YhOKMZaHy2Gw/Jk4ClBhexa+Y9oJOh5g0POZiQ
GYqkMoLA+ubGtSDAdvm5BIVlJh33BNqNCfiV6naiywXlm6uCP0wVWYGRgCh2gilf
Ak+wuBmsKKSGuHX71KXqM8Md6qXPROZ2cBqlKjLmc0JBKnFYet9R2nxsUe6iy0L2
ju8QhdWN/wpvTbRZcNJa0XCFggRdSFtxLf1kwyWiIDTp/hcfkx7kcLbs0aZU7rEX
YKGN4oM8TmuddZ9NV80JL+RNpYsYVxwf7xhF2aU+vsSKOrozSSz2K2NzvK3shTnG
K5l1xDH7ykPQFJZsXRrnCx7QiJwWW6WTFzNuai3J2JDaTlFJsUpQ/CdhoMxw8SYJ
sUrGzdykSjvlr4zsUEHRIfBQcwNptLpZnROBCcvCchvn5wOP0FwFMCrdaWpz+zrg
KXqV66xn7DulTSv8oQOu0sczY4Pu9sDi8W0ckjcKIYhJe3VGw7/YpSLgl3iySSrk
TJEM2+tyHalCU3688B0TJ6VhTuWx7RxDW7YXih2CkPdWb4erNae6SSJR621HCY46
F44WKYKfmYdEuFIth+RC+mJ/I6Ed8uGpQsfZd+Nso3CcguJStIc3opijlyVFHmrx
ax+X7iGiK39xlr03bqkMOm3hQCFj3ph3+fjgrOg84oanVBhjhlB7R04VViFcdGFO
qqPLQZMsZKdruzKVsvQ//igrKDN43vPLzGEsA33eiLPNpIUZudpvLgmPlXktAvhA
91JZzltZg2IQDSOWo1eVsNpQHAooJyIwWw9rf3hPt3USUucDHIgEAoLk9mko39J+
yJfaD7hw2ehfNq5dZbPHysr4ndAFP+gPwsBk03c9Ws5dIQey3E1CeSFPD/pOvXpE
wTKQV+iu+hDR914q2nj0vKapKUqn1As8WAVniDBkhH70JwGCRnoKOzNLPh9+tK/m
RIVpF1F0NA4mtpvI51iIOyL0ikCAPua7UsnKW3AToGr7CdCmiuTizJXRfoxnTGy9
ThkptK5LHlTLMY0V2QSb9CJlk35zoUzyeRdV9GT1K0V6z4asRl5dpxyek44sGl7S
26FUM+Zx2UwX05n1V3NYAHwFbPrSvmVGzHyinE/dtnnsMEQFLxoOjrBINdjCEu0R
xLkjN4B2f3aWEL/pZg7QK81jxzPqskDj6TjyoBW62bCzAfxQ/AenV712zGrs7wuR
6jjweqpoU7AhAgyoeaavbL/cx3dexFk46o8evVqoxH1tuzUpPTMdlopA6zCNpqDG
pNbF/mJ8LOcZ5bRintf374Bql3ciHR5BwIXD3l7CDZqFnJagCJPzA86Lnis1GyvG
JEV64BdC3ltnJ6hfU7eIQ0TIiY4Jik+I9J93cWAaS+KJW+Geoc1VJDAKtWq5DqUy
hdoVVQPoMcKPodfbqXv2P4521YGosNSguUmF/97981pxGwSv2ZimL59O35poRKkQ
FBMDYKbycBoSdz+p34rcP75EJwADmFyfBbw1FceEMVmpRN0mn7GgVkpj5XuXLmrt
5BHQttmu6QfWW0RJa2VsJ6C3SeK5WnfkpaX+gs7BGrhynj4V5O5OizafQOU3MVJ8
dfL5oCrFYBpY/KWXJb2aqKWJcsR1WBjKDzE2T+kPnm5IIPeAzWP5PQdyEdKqVqe/
EUVKl9D05SJ5BsCxC6mvy73ZHoq/oitI2E6I9C2sBjgBCA9xvgY5tAlWrwA18iUE
mAc/4B9wGM2Z2Jm+AIVRk/3JMAHPMXV3RzDd/uV9IaaOZtcoKg0MHxSmPI6iiPhw
SGsS6OIryTW783uw1/lmU4u+jiPUOrDXxptoUNYLbeFpZWHu5cBo2d9wsDcedKub
C4WDbYrHKW5Cye3rQI/yDFuEBS4nxyrvQtI3/bd0JbKkfWDyu6gvXve9QSk4thvr
v0bgNYQw14jJnQq7U31eWmu+8WrLmbX7eVTA6CU2yYwrOG+m5WELmd0OjqFfpAt6
65xlD5icSnv++2VPIIvlC8pVHskfDAW0X3hPCT1VNNgkv/JmCOJ4G9NHbVo97vzE
/1DXZFjaRHPNDIl01MvKWeGAMIwR1fmVeUmOo+xY94NBKn7Wg3PZmMnKAAUaNDay
eB/TjwH17oA1h4XhnvXPAW9YS9Av2kgDNnMRljlsCBxGujaRvKbi0bRW4lsGBrgB
Dqepc8eUl+PluiSqk7a8zqyubXT1kNosIgP9XM4zWtUOyf6XB55Zj3zlr/Zq9oP+
gHCRW0CaYaEse8NHvCDhw94Fl8ZwO2yD4C9rjj2o1xswQDxK6PSY3iCEzAPqaNTq
VPcxXJoSvRl+tJcebUbp0pegSEt+51LuJOhncWPAFUGwLXwX0PpqIipAhJ6dVd1D
Q/4XL9KhtpIcXFaYL7FvP8MZMUk7tv6JEoelRHzANeujNbQgs1VJPq5x+fOpD6ts
M+IubkjAL6yotbfYyfEsP1LUJ86fnXV5SgfHq9dEVTLJWWcn3D4jYp8CowrQBPw7
P9gK/UeWpp2hoh7vFxwP/12aallOEI7odt9I+Nd8IXP9dEUrF/yEANF+dR50SVT9
jaiAfSE2qwxGnOj4oPec9Njb782QM8asYY9pq7VPzmkiio4KcGpkGXDnR5U064Xd
6b94LjOTio8bQ1P6xytEXX75TFeAHtEz3hT2obM756xm57NPL8Q9b3sTq2YQDudl
NqqbsCQCZ0zqNu8M8Dvp2qrfsaIiCkSHx0hthWtlcc2tjisYKtnbnfuTW+fIhzbn
KyO98hyBzLCq7q8SnFmJb9Bc8Ihnj8eiWtJRelT6p8Eyl7T+ZzKXJzbkvujsgHwA
P7dboKdnXYgr9FjTjIvZK4VvHGSI9FGz9afRYQVRy+SBydhcP9Idpc1lNsDIZtex
Z/OAaIh1HHOemHV1D6rciScGze5lSX3lXg915ELOoMGd+JKkBJyBASW4anU7ZC5h
xhiJXlkXMPQNem+suyIJ0z2A9wknpNVgBTLzPbHPuUlAcHRp/bIPw92m2odPZs1U
b8qpDnOIK7oYiXMzDk3ECbn33xy2Iwg19tuCv6+u4mxVVeth29W58Aoum+nIgLzE
YNWHUndxiE+1+MoDFsJxUEuIcIfFjNh0DHc9sKwlVJfdlt4sBlITEpV+KEsIsyhk
Flgl6KN05dqbcHNLYf/3hHWSY6hBxBr9dwY84cdpC3F9qZF2Dg6J8w/+WaWEeOAA
3K62zB+sk2fsFB0YDgSRJccl11VBuSQQCumZ94p0Li3sgFMuTzAihJkDJLTc4TVx
rHSDkcswcApb52PYfsvBTDPSo/oyATjr19R9ObHC8FYEe9ZCehqWlfhjrGkxTNIe
hL560SQM3Y+16lfAMDyGVh77PGdhUgV+UT3DStPR2MT9vq18Sfxjb42tJMEegV8i
FNIki6eyTFJtT6gmj++dL+7ktHA1fpDUvcMx11UJZtuaR9By+nczdVD/luKDVXhy
/x19iBs+6rhAKTaRPSE2N5uPM5iGQWJhnkt+kG4YCMPsBZMlXZ6T5I2DPHet4VRJ
2tqNuUfC+3Ie2BvPB+gSimqVAu7fHOxwAYTE9EJHKKNJ9cCTQV/MAWtGG1VGIIfz
6H8cpqwIss66gDEy9Ppi0Brg83M1KUdSB9yt15idgzhDeX1FxDtnEy1SqFxNPlDA
dBJQ/0P5RSATgG2dEGIvjoFO1OiQ/O1s0M9ewjmC2AgXUDDcc68HMGOKxTKIDzl3
3b2X+JbvYQUxH8ASiAe0F1hggJLcw7XngTR3RSzmRkORGpthZ9gZU/QzHTEOqZop
C4nDr/A45ytDsuGMQDFGqT4VNRsawbrYzXfNALiA9mTRTTsB1wYjt+m4wbrGN2sz
2Y4eV3ss9dQA8nkH+k/NHxSFRGs/m8l03lh9nqzMDOwNUa6aSNBRtfDUWD8IESYi
foqzcei0FlzLRcZcHWE/BF88GWX/AN8Nk7xTZRhP0l7a59HM88V33Cp+j3c1Gd85
6tRg6oriTUMCNvzjuFv25EQ6CkuLOHUMWN3EJlu8t+7tdsh9uLrV6WX7L8gsAXRC
ubGOGK5kd9R9vea+QbZf99lCA6eMzyPQ6iQypYCAU8+03j1q3vwa3leL7RcMIjC7
sHbGspaJxNRD5Mny/zii12CQ/mgEQheYHiVMZC5HETw0CKNwtAny07y+5rfxpica
nXGMUI4T0INRk5D8zPbxkEUVFUlBrDlXMpghosOcLDibZXjr4AZ6x2SgTO56osSq
vbe1pQyq3XoubZ6ESn1q3UtbxCec8iLDVN1JLzGHGgrUH8xCi42Ob7yD19BNkfCx
r+e7QuhjBxd8tfpR5bDoMW5wpg8CcQvBdtBhXZKvKS+z9jVYipNRkn0el/Dd0DJy
AHg0PVXb/0BRBJXEixINv5tTFDn+7sul2BaYIQCkk2P3u1X7xwwm7icF2pUtHb8J
+f5sK8sevToE6UFkfBzwpxrIQzlXN7wZtaEDtksQ4YLsF9wS87i+Ys4EK3OfGsmC
r2iH94mfKRq+hDJCV9Z9/WHMKWCk6blh9/hhTsuUQijOBzSpnsXWmMP+KnaKRMHw
vNqOn0aOguoexiRNwkcWhDe4oO7dCAZm9+e9W5skOeTLoY+j+WZYlEZ7WqpyiJb+
Z1sQgVkxL369r+1oErZcccPe6AHOjUjnx1M3le+jhIGyEghNM8xbaKv0SpBrF3+n
tWkd18cqQjhTxMqjDklO4MutGpK8/HWa0ZhfvvnQxGk0sAPuXCw3/XMpMfGqkQ08
6QnIXAMXB3tx9CwIGtUIzDxgkrZYl9GwpEoQQbGJGOLH2hrIOg3X7mdpSE1M7Pnj
D1W0rN75CRZXarh6ps1/JzNa6M0G9FkydROoqLDAqCEuMmr+kdSm9NjjF3KMu0JN
5ef551jQm4pcjswqQyK0DIkE2VMtm8Wl/K5P67raaNJBfhzUtvRuKVgJ9Ab6QWl2
hfl2DpW1LLJSGSdJc2LBOlQzVzqTnUnhxgqUuNELuUAjTSK/C1zjBI3jZg7mD9k7
eDHDFuRdLB4csDzndlsQzHSKiw710fb0jlcERwyDNzL1W+Y4PqwUnBUN4PmF0G3Z
FIGA401p1YgD41OUG+7cMaoNh70ybldt/XHCFLW2gaY1sR2tT9VpUFHCu7Qz7bt6
+IpnT1N0f+0Jbs1jFCWrwC4uKl03yV4X6PoZwwcSm5K8SWDJTfRGezDU9FL3CU1M
AGhJFKlr4QzPi1dXkCiaRKBsX0Y87e4SLe5rETYcenQXY3Q1sRd8Ls+G3jSgLumw
aKYioM9xJmNm2fcGvQRai1xbh3bQfrwEGNqV4sDX68LIcIOBodiHBnBwtwI+/CVN
4w26lw0tYah9k9FKzTpq+i2Y84O9zjiW3NRFTxng2bs4vaqtwei1ZIgGelna3NfM
0HFj76urQWhvnnkhIpWbFCpB9KvReP9D9/gkh4dU1SB0BYwCHnrUnfNEnD8R/ifF
RLI04wvqAMB/EGGoW4AXN4iCddQ++3L/uKfJaLwsvHZoux6c5Xlv4IMKPRVmmhEX
IFGtFa6vKEaTsNi4OrkEZKg0gA1VVzXEAKMytIXVNkURsZ0Xv/4D2JQB8uiDufia
XZnAXNt2iWmyHsWsezZvUx8dn3Gg0XOPixytU/fl/J5itWSq6u6Kej1KooeARWxH
a5i/aHCuiCygVMReHIM2pQfF8pegeXfxNMXczDW/DcKjCL8/XN12ePItYa+0gwFD
9VABnzldR9fXUjK+KamNDG3UKUN/9IpoNP/D+75zJF1BROag+HdbdkmcNZqKjToC
dZCpu3wtzSZwS7QDyYYGiKkHdS9IhYixUT2w7rJl+ZQY3oVCpwMHnzR5J+SwuMe7
6tcGMO3Ccd9ByqXAhE2i/x4JT6bCjC1gqqUstoo4+PAtAvNnfJ+Nd389I9CQMLAG
PS3YuMznH+1DgOTzhca1ypTheKcvZh6nSb1ooqfIHS9zcuLL4DdRLs6gMI4B6Kmh
nKYEPAGO2L9gQwKeKE+GQFRQtqxAlvzZEV18huLh5o5Vv8qVc7Bmg0JEGaslDHis
LlYIHBG8PEUwDzNCBeUli02RyeK+xg3+rgsj6tGlF/B6fbWEhOujcltXJICEa8zN
eRWKD6hu2iqRrbLIK4f2yCX0R1xAiYmq9djqlaVUzeRZIzfDfcDAqSJZ3cuEYoZy
QradHGxE8GWasbcj58ak4nofqZZWsrhglVc2Vr/lMj0fmB9UgpgB/L8748NDJBE9
CMIm54pF8b7cMG5sZ6D7lNUoCRe2xFukLPeNkFKjGW9nUgb+kSNUns8Kd17wAw3q
ZTTkxE8MPMy/YqdeQNWwlOag6YduzWPtUd0z7vjo08Ij8W1r4X1g49lZjpajwA1z
LL+5wkFeBjA4+pJ4/4oobca2X4++4xTTZUM/7azCzk5nBRcLdUil2Qi5MFFqb0bf
lGxwDnBk+HlVGTa2jHxzfsTn8uBnhL35WatUUZvS629RGQvNtal20ZVBDlsUM42i
sCpRaHuQCR+rzlkFLDPksSdPthqj26/iaG2UX2HNdUdaC5bqK+w4B2OufDKhyeC1
zvu5FDTq6yT0tMe87cgaBi56UKEbS/k8UNMcixCe1v1zc8pSoD0FVI716+s4P175
CxoETZYZILD1rqnOnS1dII9S3i1hLVbkJCba9BZocCVexErZJ1rfzRWTCkonDr85
OLQPtm2oGMnfn1fT92ZfALclonxkAejV/OEDZ4XfUlThAqfRaqUqNJmOVStNhqJD
hg1UTt2wykaqjTx/dR1e1CgC4GeSiZGPoFUClcgI3ayq3ynt2MiR/gu2vmU7YGnm
iD5OXYn7BTiEjF1l+byONbwTKrzJVUI/oW0dFl/WI+jMrlMkdQMwdk+ZFh+9xuV6
BdzGSTmgyQSMwzvjsCLYJ6a68xWGggJ1zGPwmfSa8YE8qqcyJfa392IFL1OM40+/
6X8tbxq4Ocv4x3g/VxXRdNy1jPaj2Pb1e8vGHIMhjSC85p12LsU/i8AgB/37IlO7
6Jlzidjia0biaQ1gk3f/IJvh935Jf6XUWgu+tM60eyx5rx01DM2D/T4BcfkGgS3s
y+VtrylT5e0Yyfq7fAUuo87lR6kkaa2L4EcNS2htF8be0AU/rZRHv6dyfBc0XIxj
N2HPhWUWpRCqTHvPoK3MM5WoKBAMEbz1JHyKLOOiEtKyz70oHjQiEonBnJQrKB2C
VKSOtx+Cn++ZNQYQIyOsFBG95zKkwrhkWhpD+b3lE4VhQCvlsaz+4H68AiCzDUl5
x1lKueeduPPZHhmH5eoqW2FNuv8CNVyYd7Tyr0xMcAtOYTOm5KCtzLj6JFIcoy1y
b7ttKRJRPS9Qgy5KuZPwIusk9od06LtmgME7JdtO0xbaqaDpVcmVHiDGj2b54dbG
XkSF5Lz/HWHGe/jj81GR8BoPE+EdKuogB9J0lpdm0cCZ//LhNiRbeT2n8XPRR21f
qW0wL+KDwR+cIFVFZ/6WxVNPVkPjnCbn5Y5hwNyTzSwcYtvdLE2H+SOlQ58UL0UH
x2O8qsetUnny7NekZhTuBgdR3vBCGtbG8tNTqB6naIlucTxXBbJhumdGcTypYT64
2eeMcUNmVXqJEUzmIFih+U30mv3eQFVoC/7RkT/5g3vsTXKr0OnU/vW94eG7hvAc
T6Vtp+9LO9+gx1gObqrzbIrgTNtaTpGni9SydLJVBpy0CZjaYkxHcHWEt8Fg7afS
KpWFtFHlxCsXYLD4Av7zzs3j1FAmXJ3GSsV97Tp2J5ceWsofll4ygJWkangHKBSe
nWm+peQjPgqTTF+SA9dMCFT19bV1MKPTkPK0HDtRoyu3U+CSXyz+Ia2tbxzwkPJn
5tcLRBafE99snK4YIlKrSdLyIATosgTWt1uWM3MuVZaWGbIh1q4qyDt6Q1foIAHW
Gbi4mA5dBG5uU/GI4O00Pk30mnRIbqVcccmI6hwgHo0iOQXVyB78DwyVJTQzVzDM
TdS/mKHZBSG7ksge4Fm+D2SJeiOi5y/gO4wNZpL5yyimrJhCt2IFf+IkieoUUMTy
nNoGQbgYFBl4Q67vn4ZE/3p630IKtqExQfSn/ebdU0vww4TzkR2D/HoOQHXX+n6Q
X90pfFg+sjlyf7etLElDctK53BjV9fwUelywavBDCfduR4Jufky8iWqB0Hhc9GlP
/zjPDt+Trr7EEWBJUOMiqFhBGdvmu3WNDNLaAblCRezNIBMBqaNTG+GRK07j3eHI
ZKxtm323tpiEv8Lx1WgJNQ/RcQ6l/QO7ry8keiL3JFoTEHp0Es+irFoQDgqA3GZ4
x2Mh8teM+4hJLeVeu5dnay7IOxi4uiX9tE05T7RKL4ERODb9pXkd6pg9WYenSFFp
GpAjJ0vI5bOjKlOlnhaXxwd3HLWZJkgHbhswTnEqzJExVfRXhVK0Ihqr76xscIo3
uv0CPl3Xmb9jmFsVheBmTbeF+LyMZqCWeF826+DhpTJcNEDfNoReCMuJto6oYwcn
4juGpdvMwm8Sxturtd2UB09qvO64EqI97ZyefJU/BhK1ItiERMksbRuSMBX9wDii
Y2SZBJjrq6WhC7kbNfmIuHyKxoLtG2LBWZmcUd1lU95vp3eCtq1mkhInC5xMC7Hm
eBcsqV2Be9xnG4BJKv0LCs4iqv+flOFyuqTCfDsFJjeAMQT+yGt0sYeTOMJhFUPJ
Z2iNqkRZ60gTfPjEbJrBDa8BvLW3VIoFD3nztK1NzJyd0pYlPOF72hqsswNBB3HM
UPErMdWlrlqjKolCQ8PuD3CY54SnfJSWuLS7Wj15mRu8ZeCI+EmJsO1MWitCn1+C
raZW3e2caIMVL5FtcnltYr3d2dAfy+KPMGmKBABl5zOjAsO1rI2jlHGyL2miMjCU
M4NZ1VU9Z8J0Old9LL2/J5yt5ClZ+O2Y6aLtyT8hWcTncSFlye1f8yL3YqYt9PIz
NQYJ+mW8yfJnYp2/Dxu+eclNYiijsK0nCeGVU++lfG3N2wT7NXQNFRH6yNvGRL2m
hb/qN4x/cPRkBEICGeEvSs/AF0WUyOy4y3DyC0pOyZ8ylgqE31Cb9YpnVru9ixVK
PS/N5Sx24UV6Rwi8sOfmXcgo6jm0JmO9iFoNMH0x5KR/Wwf1GU69op9m2t8nDFA7
dh3keN/1nnDkCfhGhWjdFSz+O3KlDFWk9i59FPNQSuBnWusHJ22RENnldN8sqajC
MBPfX3bWVPaGysuc3YkS/Z/oMMtCYWnn1uKvHQ2uHCTZAdRgaRIGhaewhW0qPRU6
9LdRwi1Tq4KXA+Y3GHBU5+iM6Q91ZcbkgQYF3CNDtiZfPigOQz+efowrGk/AFkac
KilHdE5/rFj5tPeXFKU+kIc7/drVmuT0jh4gMCgV6WBmRaBZ92/Z1OVnxEWSYlWQ
gfsVPXrqy5mwSJm8EBGaG1fWPhyHYD073hlRxIuGKE2UdlgUtjSggcIWVR/2vI4M
23PStuD9qt6W387mQLjG93O6v6Hq8ZVA4X1PVZig/Nepi6sXkOmAKeCBsoq0pLQg
07qmkQiqRRNQjQx8gXlKyxERbXB6db5nLXGtZKsmqjUjwdCNjO6ppduKojK9LuWF
HkzVIkDOqkxLL6PmNXZo2rP9jcwAn3wciczY2128QeMUf1Vtd+VJTq/KUIZCUbER
5zmqpMQfU+xm23ooQQQqtq9yvRi2XVtPjDMb0soKgfJRvYPiPSzLU0jE13NSmJd3
zdB5wOW02lpGv1wQicTeaOINHVgIrMi0TJfHoC6XFHLdI24hnuqC8//y6fNvGeGy
UcKXjcuoZA8KPWS3Izv61xv3XSVcWa5kcBxjVAZ8eQvou4s+TQDyhtyOvcKkT4Zb
n0dNVvFf5cB3hVdqqOJsptzfKRPMllGucS2EqxWlPNvxm4ttLpWD7myfnMoHZ7IW
uA+lhkDEHpZktYNxQ/qdA/34i8vqLKnMSWbNE5Izykxp3+TRFCOa+l5UE+yDIXDl
Em4zYlLe2igcKb3H27IpR1fRYvoCTQalyEP6mUoSWAZvZY01KthkD3i0hDPHByvX
dTGbyb4BYOCY70JeBAkitsM2v1tLjvKAasrPfjrfckkzqu8DiGUA3MsEIjQ3hvUm
2080dBuZ7k7dJP9P3RefDS/xYQIXrdi1Nqu9ET19YyXOiwy6Q93Go7Zw2/LGAWor
xTlHbp7bIk5XM1+FESy74aMmdcpEE8swSTmkNLw9Z5MQfNxiIxWB23H3hX/wSqK3
/YX7JGfKHUCoxCu4LBMxR35z9/6Q4z6ij//rR37k2dBCKIn2G94SqqNyZu32ZNM4
Mrei0OVCVlNPYDU3gtAB2G/j2mJeSydBl+fL8lXefU9syJsM1xSFlVPO223ANv4W
b70O5PuKi7KzzTnOogNI7uBrujmZyxRCY8DzmevuVRdwyxlogilV0P2IQN3ziGuP
0By8otxOSqf1rpnrMVC1F0vC1Y+mYdNteYE3BHEAeHhmTHx+R1MyRtPgYZGheXb7
zy2cSRVqev7bafZpH0KItKhLEN14QdrtLLzfOjTnu6BTYBEWHSzomoc+m+tUkL4d
tkCtV0YXoXO53Fz8nMacEhvpEZQdcAu6YjDegU2baNi0LChNgsRceQhY9BeCg2yk
K1KgLxkE5A88X2/XjpPtG3AtU/L5Zwka0Nty4xEKtMKkNloyDWmUHkMOCmzXOXF1
Hxp4YdpY/afnFwetkwpRXhqfA9DHSdp0t2yyxmzdvFt+cqIv9GXKsvEp9m0Wxf0l
ZlJaO9hTd2S4V+673qIgJA5GF9X2jvn5oEutGhGyUnzzqwrfjQSF+7slLClcd9Eg
irdTBnx/onXZtZ3Op9nKgm3AsMeEWc/A8Xbe/F4h6lhRHa4uth3h4dyrWP5zYy5s
FisyVa/4AJ2H/Gv/69a4hvYfyjVglE+rr1kY1v7ykbw1DnjRJXcXA02QqL2DNPAG
jO0Ep8UY0CYjRUixbccUxk7NjLGLd9sM7RmR/Y3FEWtfxNjNZIbYs4mjI/v3uCkZ
RIKm9eBGmEU8ZvvYsVkV5c0vAuCGEHsq56iwsnOZD5Ak2V35dhQuCoc32U1d7gUu
TPNx8LCa8eQAUpItYbJdF2xmD+CEs1C86n2CNDAPJKzxgOBMN5KMmGrWRyNu+1dJ
V3TICONavVPGv8HA46a/68R1/ezISXAsQM8KGzm8JeRjmj7+DDG5Q12Ktcq6zRiC
PTofV4EVbCQH2u3LN4q6mi4njUVsLIZMByKWhGhiC2EoIh9FoKBKoaoCyCKZrcq6
3orpEwHEk/lmgODAy3G9zUHnkf8nGxbCVkM06zu9+SOGBADiIL27q1KYuvZVXENs
J27iyz1kp3PiM77xMkcKn5R/Ml7oAF1fJEbWDIducsl0UNgQUqO4dsNW4QYBirtw
fX96pbkiLEJk5udZRuKY+QxglGD170fqXdMSI0dzqxrHNFejDpTz/3wOy8BxDyFY
ZgpZyzikayf8VewU1bi676AHTFR3HGbTd8GIn2/K9uUQU1o+YGKzZI5XznyKbs8g
duylxNF2tQ2Qyq4NU90Y7yNPw0hzZpLrQlmmfF2AVx8p/DZKFzgofp+nAzyN82sy
aY62Bz1pAxyYJVfnRr07V5/UeCCgJunB/gSM75Rdm8BJ96WCRNWibBSVJL7JNrvw
Us3boVQ1MaMOE3rCuCVmp6L4KmYl/jAsfFUvibwqVuw83ajBB0OV1si1O9k1hlEK
R/sO4FWNPFH+xfG4AW4HQB/QuAuEjhj3vN6RIIzY06VWK7nSVRy5X/AZcJMMMCb9
p0gUwQNAUC7R29byu/7kyoi8Wn27zIygwz6Dzxnsc7UTECp0LWAE82TPP3f/MC+L
xxTFNf6rswQ5QFrjJdTKNk5S4u9IhJJzcv0gDwqpQOGpmMdFlRD23wOv1kd1nDN6
4zHRr2aAXtBUW1LYcxN3dnav02jbKjrULE+uJt0ArIuuEj7GEc6uuCqANOOfwWFb
36IIY3+qrtORRiwXukpQWC23a33jc8yk6uR4mll7D/AtUsnWGgELEPv0vtWIWEer
hVtZLHDJACi5nOwwvR9WjHhLNVEfQwJOvF1kFBljZo2qvljPp7faS6dz+niXhSnl
vm8DnvAjX7u63ZEvEpO8PSHcwtxByuA1y/ls1Xu982IOu4BphRJafPL+l5UMcS/o
45fmfjA3B9tOalojcSF+r8nGYrDgBDL0lmQdd+By2EL2Rudnho5B3SmHligZO+KN
iagG00E/b8nEgrn6GOpuvyog7F9uTNDt5Bmq013N6up4tNwNiczrJ/99REdR9wfD
6HvzMl2NCLp8FcvEiQkzTEuahByBNZ/wSOTggnUwr9J+zHELaVA0Tk3e6cJ87AJp
PhyxMdgE5cYKKJjquXUEL90Td4Fhd2cYudd0CBGV3RpB9C+hblFZmjZ6KsZUoyWI
m9HcuVbTyrEhTrlohKOALR0t4BvigWbxS6mkY658OY3PXHT/HUXd554cf9De6r95
hMg5D8kq3gX3qt35X6C2G/b2ZkT8KrlOaxqCxWrkb30IaPADsTZWuz8fZaTdJdRX
8brVj/VDAEJcVM4Nf+o9886gaJoMpHl0AXHECwVU2vw/6ZtmfyCfSmBaAJMcX8Ig
KlHPH+ybC9TmfL/n7SEVmSrMFUqt4Smkwfn1ckOwJJQnMBzimnEKIGb5MKss+B0W
5Kpe2oLql6lP1yhhcuayvE3ZDYLQ9M7j0+3Lhh48C96PLExCZbpEoekX1Ug45Qih
Undn8jlk+OUZCT/mnIZhK6Hley1h5AfKRTG4nYVcHHTGAenzZ/jOXM8V9vhENroP
G+gbinIYUHddtoj3IW1fUQ+jYYSjduYm5zwzULxsf5UsznupNACCz0PRTw2t3JC8
OT5VOvfHemEGYPbdtATO8hvp8Q+i82ve/5TDkCifAv4vOOzig8bjkgYAVOCJ0BBz
cKnhkZZq1H7XyVjcXWLR1exCRRF74yMl7csWg3jAA2iPhBN5BdvIDP9lX/s/lVqS
5GmaV2VdJ268mnGsRO0atiSEIWJYPtH3/G++jpp/ZdW6Rv6nmHex5TuE/LPfTYEl
e74PjI9iQ/lOf4oS6Pxl/sek2/ZtndNz2TILW94E32S94+16POcLgTus4iZkj9pR
xyp10ypdgqUZ/0CFoGZap2W+po5K4I6J9MB4TUh9ubHVgDRvi3zv3r7bHykOsOLN
LM0mPbFbzYdSdl1nXUOTCMuCJM2Kmi/qR1FqTMjSDvJDXcOzRVItRrpPeZH+GyX0
pu9WaZ0yw8TSxfotNliaFRV+cYXr3D+Y5HSMU5Wo7L+Ot1uPO65FfIjKucWtNsh9
tZiJVcbvb2p+RTh0Iez5ReaFkU8hqd+/kDWuhuKVXmlmXr6M7658Cx+jG+EZAXEc
O7wgqm9f7eAHnKEELOmYwnxyeJEXvgOf0cM8PacmojoPX/2PcR56CNKfGbxJumnN
qhxd2IcIJ1rXSwdRsVGavf/5iFiYyYnWcPRVifyR2EIaLrEJBpJAIoQCTEQsq5MR
+lOd6MH3fh/FFqQoIF1oTJygS0WG+UXnivAcE7vIzmEw7a16W/NYetDmHEUn4jtP
dEzMVfCmp0o75/erzp3qegqmfoOwlPBgBCoGKNK7o0Kf9xAymXR6qMcBFReutOu5
/Oo9Newo323ZME59XPrBr1Y3eTuhDavRgOr3ukwkYwijGSXw6YmONJuCB4uKLJQ8
f+TELxTFVzevvbZmiOt33/LCiZsCkJMwI/NRlJeVffzi8CCQyetdtgCD8IaOfI0W
dkDud61nsXEuLTJgxVU39rMrTIQMf2o5vftCF3+H0AQ1llb8DZGUhft7nbrEuv80
O2MHqWo2RSEgzKeHGTCct8p8fEe0FVz+7rB67c5dVtcmbRfu/BHt4Mxs7MJR18ja
8QBUr3ceAJrkajOuKK2zeUQNXakw6dX/SCfVHaTi6azFnQcbU1Qp2fdzsFKFkybq
4cJsEcjN4MBtpSe6Xq1B8xtLb47Yo553wkkjI718OKBVowd6/u4gyf/1gO4zhEAy
1hRGEWFY+f46ECuprUwp97JzdAeHXRmw/oXgSDTzuElbqWrROSLSP141O8NAOo1x
7eYiiCrmYo1rsYyStrKYZpY9bOe54MN0mGCjG6ns4adCEHyJgjsh6rdmsnvMclbA
+LfjOR0XiazitbjFZmg6YJTGqjwklGWpYMVnRHAsfNCsL1byNLUjmlMdKOc8546Y
YisN3dht8MCsiprT8IzRZH1mG43ctwHmNTkIKOzEVHKRXK1Ty+tFa+tFjUzcn9DI
ZOOqdZqLe5HrM8LtA1D8+74M8YpVeaqMER7ThFcvxsdSjyyI8f0uY5oF8VZPUnq0
1S5cc+2HfHkloP6oOa94RyDrKCxeDCSDw6FpLBs1IxVNPjKibmVZE8ou+EfEB/A4
nZxehVcl28XmenVCoxUsRbovtkTjA+PKIEwCGrivJvkRGir399BTcBiZNWvK6T67
UsEWduc9XbWUw/BQL3moxqLIWVIGdusOCZRPwjzQJAK0WbHE4q0b3kQTFkLiBhKk
Mu6txz9FNvotyuagYKRVPkyHEEg/+9Cly3PFdtVDXsP9AHzMbIa/ncDJbovs+RAT
uR6TgU9eG5NYIeMn2Dka9QpafHTug5riiSgnbbXLcI79sbcoJk/AK7cuGnkL+Y/Z
5+UA5vsyBD4I7fKrBwBQzc0hwVCc0Nof4Z7FDHSquHvaQI4ya1p6wuN44V5S5HPy
Qa7aehLTcpELr/m1iEcS1apaGpE/K/uFG8m9nOCfRTqtHoOBpCmuYbfXA9SXsQlK
2mxXep/0ycCoIUOOeTxS+gIVWoc8fswXX41Y1PXTFYDGyfvaHs55WDC+4VwDbH1Z
2mRdC/B2EKy13laAc++of697o74UtUoJLKaml+AY96E626SE1jxLaB9R3M0OB+bc
O/hKfe44tWjM+BtfpPdTby7wfwU4rANspJpe8mTXjLWtvfZotauj8ed1KrN8xN1/
NVIX+IpLAZqtDkgAEd2k8IUSSEd92H+Liqz6Ok30cLepSSEjikPnrEr+LK/oUDDN
3SZbMrLhl8Aed9dtTIlX1qYSr68z2wVeCAznTGW4GKCksKmhJ520GwE50dxULhLC
bmMyEbgnJHnz5DzcCBG6+aMbzfi/wQitOTJ0igUTHm92WDgMAmhPKuZjhP0HMmPk
3iKpx68JDkxaewO78KT3NXElukESi8goK2e+SlkdnukgM3wlpqbQNY/JtxTwevCf
baVznyRUjI2dpCOe3+PYl8LQkG4aAIWHjaPGseo5Wgez66GgDiQyLnr1gxLd01YX
Bj3ChhnaKB/5LY8MaZ5UVQ27EBH/C6lWxAMf+nslUrd52Vd4kwE2H/J1eaHCOi+T
usVWiqjmG3l9SBwq/xYCUF/Xm3Ol+oQGvqTHuQ3I5ZljeXwje5HqjMC9MQ1c+iM+
vUp26frRtDkD+eJzFbF7reZL5cek0ikAhYCobsjV/bHjW6enWvNkszoqRezG+kpo
Rmw9NvkostzrSUswa9DdplWUYvKp8JxiukbEmrBj0sKxb4TTfKGG+Mhukr85mLMB
MLhcl8pd5+rfNkLI4JbSHFb5ItZFXs6ryweyQvhCVza8k7OcsPjuHPQnx7TsK3/n
379P0TmC9EyDbhDcC+0aqtPFVZL8YYwvl480JTvqw/DUoeMKUbg5HvUc4GhA8wCG
EHrT8FzEM/AR95Ka1cf+n5vEl22KMTB3RH0bLn8H1e5UH0WxDFZLBRbiyIRSG4Pg
to08D5fK51fZpmTZclpkksWVhfpxN8oEmlzT1rBfF40kzCK+35JaHh5NP0DlGrdN
qtGfulrKHY1ikN/UnPtfKx5IwVW/VFf3JDUnydp43EDnc8cEpZ1VInUWlfcQzaU7
01f5T4NA85g0kNVyv9AzztfOAritI+KhE2/d0W7BGRynbgwJo+rXUJE6atT4mFMz
c3kDVn3lo/ptrYtYFroLppe91Bjc0E7TgsBocLFgkUhd0N05mF7leLVU0PpLxj20
CIH1RIA0DrYhq0VMdOMKsdZr6s9TR0LH/+vMGosD9wBAP58/LeklGFX76ZHF6yTk
5WzxKIBYagHf6Wnxgh/XovWQQ8RCuKoCs2FskkqJCV70Wnz0WO7hRLWgQIzkJgyj
YIJBQDAJ86v32A2hZ9IbiSaltU1J544RanYLPpy4sF4S+ZrYJ7Umn6PTxP+EHUJR
KIiNI4Oio4am6klY1dLESQkucL4mWqDdj9E05U+6OfNEuR70E45eGnA5qZ3yU/d4
w3Fyg0twI5PNFpn4DQY6WtVGlk/UgUfAoVmNurVUrVvk1Cro2BfioPc7wnKL0Xvj
J6QUrHhja2Xs7PYkTGHZBjpwHK4A3UydIsgaqA2FAWfginbh5CjBClkw/k+KR4bK
uxs2gi1T8nfprLGbWnFgFKwuIRqabY8n2UTYUvdnvcLmXTm+0t3PlfMysEUdNceQ
GpA4re13Ef6XcqpS8N1QiriMkjcm6uoMjTwqqO3pZaXwHgs8zJANCVmANJ/Isz0W
3jVSZXCz1A0suVY2UqZOx1mFSAFRPfW1f1gWjxRsZMR3LE8CbNO5DcX6BeyZm41W
OIkDmSrBMd0cFNilLBs0asKZ0a4KsxOmqQv4T8I/aa6ql2w0sTqL5fAOg1icLFhG
FRjIK8e/aOAqfOrxjKpcePBRhO9AGqTQINOtqSMrZWH7yeNX3sEO4jgPHKOxLIud
gFjZR9NOOQ+sQ5M/8+BJ66CL54jJqSPB7xQCRO3TxL5joN+hCNAthOJw+g2yXCWg
gQ92ZVrpLX8vpJFMd9hK0E4A3o8HNfkW9dSpdin08dfgdp9zI/smdegYrMbVT0vE
mE8hreXV/CtQ++K+L6K9Ph1Cn+hH3xTd25jHdp2BG5BPgPvE9j8TgJc9vZJ31gen
hrywNyjbvCT+sBUQBYr4BamGTtcOlAQFJW4SbCjAsQHkMHUK7F/f0b4klWNm860W
Ppo5X3WdCeUDMUNvaVpT7lg54crMkUWQca2FBeznNgHIzeZoa43DVa3e6KDCmcc0
NkNXj2zTBDdizsY5lIfNLWJEHWWeeaqYm8jncESH/fV1oUYAhZ5GNHOrENXv+EJz
qTksdTcsasGUcCfKoXqH+cZ6Sc8xhlKj3XqXlN7T0ULQVDGxbh+AzKCONJpKJtl5
2N3AOc0iQltgJhIoAo5sdTiaKBZJ6PV8k+Rc9OJgpCL1hg9iW2nsMWw71LTJOQiZ
8Iw6vVaDwUcWUAZUzk12ZxlWWccb1MTFTEms5mowOZZ/Qz8/2DulnI7gu9qQ6QAt
iuzvzCR6N/NMupgQKK2bJcOzH6AF55FSEMzC2P8yqtF6+H+UXMfXrRUOswDioQtp
VOvc21j8mw0cq52PAjiGXPQa4oQY0wfEfAlrzuJSCViUElotrKMC/Yl0unMC37TG
HOZeUtZ54r5WqE+7pJsP76Zxf+yutsWHcDqKLBeKc/qdSSaOVf0BqosyK7DYSdjD
q702H6vtkOvjaat/AZddBLBpnDDXPQx2BrEjQeenBm2dw+U59tEvuvQcWHW4WWYS
rL/1yFL/P1GPxyH6Dm7NKCqO74m+HWocI7s2e1CVoRfgzB964VgG6VV8xKHh97sL
yXnXnnc/I+mJBCkJoT6xqfq5vbFfVtwZwwTRSDQX5ri4A7EslBr3UgZTRZGE4FiU
E+Nn6xXO9cAf69v/ZjMqZkQ4WPiJG6KCmHVIEWGf7YmDhjQPkQHnj1xyguCsSo4g
7ofK6ZZq6MFzivjnS3TAcK4sI73rPrlYF/r9xtfQSJXrxClr1mEpoZ8r2V9K1A7G
2GWxDKcJopdXyut/S3zQ3KPCw/+a/EDD2kvsiQz8o7bO+l/MryRgxOonU3Et31c5
BWewEIIaVRBdVoA2a7kQouLSRJhAmhW9rIMXvdsfJXSN1ESHpQZo88UT1uGFofnE
OBg+m6Gp8tSHIOiyuXOkBzogu1gg1CGC1dHN241gltDz0jSXTtYkgvdH8VMTo8xA
qAteojXOzkF/Luym6MorFiWqkp7vUEMzy7OjcNgiK6ekvYzRr2/MCOy5AFiHshMD
qJJ/D4AiNBuKjNSkNdI945EM/iHyiuZjBgfpMLXtTB2/bgP/mYzUGQovI9goLaIi
WUeMDLnObN5oFs34TpyuUcoPmlkjalemzJsU8iBasojuVg/8BdN6USWZbOYxzFpe
yGsbpvvmEmahr9jolzgbyNGamL0AedwkfFmE9oYAEb1Dg4TiJP6RoXqdFSpLWjqc
5YS+UvPTegSTea4o07RY7waX4LAEZh0kHVIdsd+1gvqN+9i6hN5ATg8C1WnkPlGq
XrW9Nd7yYtMXHyp9l1aJ+xCdyyhjrd0Z/GK3xDx0g0+oooTx8DDaiA/pnxh7nGYy
P0UIUNh6YFH9TlPg8whQFIIGR8cNDn/k61wBbA+frFzrTzDkKYhCYC2AeyA836aP
APRTww0l0wsPA3OVZQojDzzg1XFBKZ6qwkqKLWzlBGfAQjSLVBnLYpilAyA/SKcL
JPSW0SqZGY7J2HekU5n6eJWTTqsJ20m4WIFOczf9nfQDW1lCRcCr1Fs+oKjgTZ3K
KVGeQCKEDVrtfMWjlO74/I7s23c1k7ZtNiOZev5emfpkMB7oGDME+uduYjmQeKIp
OFKQVXrrmrYyu0PaOQG2UbVFKvfEgsFNWSeKIr16chbN+UjnkOK3CLPlmnWKQMJU
FGJH2rsEXXU8KovIyKhH2NZOxUGZp2QUo8VRtb2Qo3S3yuwshpKQ9WICO5XBzLaQ
CeQkSvkZ+tiyPjBKfqxEvM4Pdjf8BTJETlpZA3e+Qu9kh/SsnWjTpxZYOX9j86gi
9I3IrBBLqzQbz7Hfm7VoBwvgLoKMx3s7h1lhLaXbNjO0Em4Nfk+np1yT+2+ax3Ec
PU4KNWTo1U1XLyOr3PHDVi43E50cus1Z8oPdDqRvhVq+cuVg/xCht1qlnemjJTsN
O9geMVBare+Dsk0aNAzO/5XUC2/KZIbV9N8Bc3cnjK8o/lstvIA+PfKhBPuNKOqM
ff0uAvmowS78azGb67+V3gpXpu1njQVRLkIL5KQ94Q7zjaSwmG1B1ETUACoNB/ea
zRqjQvz5LBbnJTr+BK6jgZX1p3aJp63DKMeqSN+1kVCUrxobM+DAma4Ky2xAnk8k
hC7psvsevIkpyanUB9DvdQLT5y+kaPJdX2hSKen8EGD6velOkcpWDOma5ywhRS9z
Q5NQT2xUa/j81SK4FBRi6FAOFM70d5n9Gf+v/tbnnYkPNznIwTRnuAtBPcKvwVO3
w1oxhEZGOlUb1+z/YaWiR+7RWLCN+jtRsn2WXpp/mUXnKeBvnQH9yGARllJY7Dn0
1AmALithr32oaMuJgya29HuVXlPkB7y7zPjkf8OPC06OTBEghKN/GKztqMUPikD/
d4sl+rLWowpNrVUClclwXt7GKXaO4d6gPRIncnmbcpGHcuLJSTau1UBtkpE0zQwm
bSHsw6gcLLdLtPtTbPy0dKWX5ty+Qar2lqvUNuUpbAhdW64cLpD/NK963RQsJgjk
dttsjZBzTUpYvx1gCaeB5w2WWyhXZL5OTyG3WkZrhDhSbEKkj4CT3XCAqRNgyiRN
pLSENoxxau28EdxMEE0oRYJXeiD0U5L2flURL0+xoP8OtN5Ble3g/BNUbV45ShbC
x+oiDvgH/T2p/2SdW7CB7tNRY/uS2AUdmjrjONFMFlFaRxQ7kEdLngG/FLAAMxTM
wECrEaPu5FUiRvzqhP4ys/hx1pihn5cfvsznmplptIKdmapxqr5+S1DmiHwWGzjc
atJvL6rxq7LGyFhNL2rDOoIAeUEGldYBa5EPg1xfvFZwhWUoehHA7HolWcpBRkw5
kpHsJuSVvkxkaqO4o+85sFklMWl3dIoLO9hrdRGxOtQkLNswKHIf/6pXWOEai/dn
eyP2JRj4wljyXli8kOo+asQAZdSaDOAii5F/uBth17h6QAtcthTpnYi7bgyiPMFC
+gl+ZAGgyB9xSiU4s9aFCUqdS2Tw/0WTdIjsV+KvUWg9E8Qt7Abs9AUHB2zS9Qm/
DlW1c21yP25wPQZT+Zgl0oLIhxr/lOV9/sCu/2OObNdrSioCV9AOkwwEwUq6In9N
vAKI+hmc55hln7DEVQgmVQayIGvt1O3rRLJkNyzFndVZ+9HiIl37IQsn/eWfi2dT
dfPMQekboNASBm0V/iGFoi8v0TQmj0Sc16QqT1kneSM68uErB4RT78Sit40fOq8o
fT7/+im70mp+jK8KVXsrYfph48YrkP4dA9Plz/RdTLc2oXvbOZIcT916qrTSG+Mx
fn27PMJiKh8+H7tEEHcC4CJyZnCNGR5ec91ZXk8tMXvEol+uqArGMWXiXU2Nvpjo
0i3aYnFXVMMpP/2c6buGHuRhAPQBPki5lc+HxXwZo7sxQjzEtIakaEpA5SkinOEP
myS7S6ETKCgxn2txPn+lEbvle0mW0jtUHsavhjKlyKl2e0Gg6ry0bc2CIHQj88fL
Y0YXYml1mst0WSRf83ngDgPUS0Nv+3ExB5VYOIFpvaFUpme+tpec2KoM9li+koLV
xibN933cLc4utgrmz0jFRZpRJrZ8z1lYm8oi/tnchJaIefO5dRLE72xTL6DYsjbh
sOfAWtTdaI3CTU0wcuH5rRjHUE/h6mnR6eKyI1jqLau4g6SqXLVdkrozRDLKxCkL
DxJ1BMwfGCtLZLkw0Xfoc2XBhEEOZzoFEn1wBPuNyk1VNrXfHFiISFlEVWBDKBO0
KqWWo5IkVZbOxWV1BUSBLZvX6T/INJxjH/XSVBqlRAIaWNtjpL3a0z//1ct7v3TL
gthQqb3dXMsbRd2scyGT5ILG8rwdWgYhobeNJugRa2lowU4hMvELroS5Jc8ROq3O
REO077eSrK3woAsz3xjI5OJ2VxEAkj8FQ2+F8FCAi99n7whl0XwHsXS2zCiFGz0M
Z/HKa7l9nIoHgNwXZTp/INKXOMpjAJFzp4uwQVMmYPa9HN/jiD8Xu6BRcx0mi6aw
R997ou/VxU94B+D0dzHlykZJhHBOKrN6TvmWN0Rrx/SX0N65jSlgJomG5+6ngMiT
4oI6P/dXZjanAfTIyOtYT4/QQ/MiJjyvWAM/yNhU0fqXYrhs+JW1Uzt1Zda828m4
IEX8+8OWcew5O/bjpvNkYQsdXzP3riGsVhUpyL/wx13eqGHFJdxVcaTAsDeOIH+V
U4t6j2k47qsx845SyGyZHTWPkoaKOKumEiLFbfAW5QtB8z16WNZK+AlG8rVzuqD2
F/qG/bc3+N3OHd3GEq4L+83ClKvREuxvP61aMMdWe+NDsdz+DcqHKtwZDzvcLGiy
HBiO42CM6Cc0ZtnosusbKWaB955hOAkerJ+JhoRwU6DCnQrZ6dDu1L6J2sv2alRc
tSzP0CFWJ0vTWm5znf1OIrmG+N9ERV9tGzA0Y5Ghz8MzYz2RUtE7R0qq84YALkXx
4doTsIuPXCD8xh/Sk+dwe8e7QOJborB+OHbv+r0s3ozmNYZaJ5jpA9mT0Evy8sN6
hyugAzXiJwtUQ/zdw0/uutGWs0q1UALuv9Y2MPg3FnR7Aw06SCozUz7JX120ENvp
DOkkMPQSYOhdRPVoxIam2UPRGSvzlO69G7CyPEhDWcncAKW4eDA4Wu8nMoSVj/SM
3NvUzl6T3AtMY8tYx446T6jcopgetfa6sJFYBK1nP3kHqNcoau6rE8/nhwKJ/rWc
umaepznBou9+anvv6g9WTCIkyy08IrFAR+Q9ZEJqyHP2qPRyMAoLAqHjBvfCLK9+
3I2+/o088E7NzSfCXP77jkkFZ74b0geiK3AkXwSgBoZTTiI6KOth2udbJM9yeqCB
++g0OA0vJXYH5HffvkLhT5PNheWcsyzAHy9o5DddUjckbIKob8DFh1vijwwp91sr
gOeb+DDB1ky5PE3HiU4CHxFwUkbRa/OgGAJjfQXIOpxqhxsT8WfH9M9KjIw/iEAG
wMWL2a3KaxuhUqVCL3NPnTaoxPSOx0oqNCuc329wWBFTvvqRUV2FOszA2AJcenUU
OmSJVjevsSZAw5oUHchfLGMG/FHFLVu6xciJWXV/pelvvRlRS73KOvDJCqbhT1pC
X3gTjyqR0iV0ci7NSyUeyYiiKQoqgoB6+EtfXF9R97+CdhyRi/dB+nGn/Qi+u6fw
fYildKjOucSgbajz4+P/ftS5nLLXJf3JNOdUDnDVtzcm/KKbXbKLDA1wCfZttPVx
oJTkMGJaJrkNDrhPzX2+/xCKIGM/aULmMNK9M/K0feJ70huhRDMotAc8C2c5RhUO
7AS+sKvX/4yMk+faAYcA0+4fg1yXh83pKshW2VE2ul2cJXUpQRLu0RJ0ejb2I2M0
ogv4DqczVggtVJFLhu0j2wHfdGm70yLhuRqjxTCyoTwXloUcE45VfLVIUPyQyI3E
rXsJDljG3weFMTu/6SxKDaHi8P/S9qck0qBtj2lxL9FYZZtnzhzXklqb0PhNzAxM
jhyUc8f5glquoPdHLZtMbAM80pa7gDyzpLFNHGD44/CzQ4ypnSdSOmS/KUkWnKMq
5P0tMDDA19Z6pS/uEFD7G16Q80GXpTiCZlAAljBDb+f9HIsoacyPBzJnDDDaVj+i
423gTU16S6zF++9cWtB5Xp3vHKtacgOyjHGXX4SNETFN42sboLbYuqIgfTZbo1tB
YucqkCw8jQuw41KaedExxyd/2h/hsIFXyuET5BtVtp4YocxvyA2hWqexQN0TshEf
7zi+q/x5fOwJ7ce+RU0+HsnYFP0taLq4MdQPeGCFEGcak0bLs4xbLmCE+QD2lKT3
ktEF/VKwh+Z9ewvASCnK8J4vCxPK1QGkDNBEzY7ozLwwEznoKTyR0+Umb5Og77R0
X5Ks+vVx0L0g2tlP/3lmbZDlJR6rTxm4/47Oh2jZF9A3EjvshEsqolAVN3q2xRPi
qBlV0yTdSMaKAMkC0yuflgWz2Dhua15zpmPTh7TS3OqjuR/J/+Zcpm/TV69OyAdC
5WVkX2VjhDhs1dEj2uKVK3KUTQ72ADKamYftuZAbdjxzfVZ2OZcOkxQACII53GAS
S6vF0vMeCld93qbDfUxlxEzdhYhv8Fqa9xdTbzLtZti2kOGP5qdFElP0OMhHJfqF
2ZZ2kb0YTGG9JY8KO+pQ92wPXpv5Y6CV8z06ubaZ/N1CWPm4/x+O+Vnwijah7EIM
/vio28llaXwlHLI1lRXsCX7l12es9mbKTQMaQexYwvGWhiq+1GBSAwDThibgQLI9
jxmab3f0BnTtgjyP6v126UOpX21Lf8vnuRABK4BCedpqdnHGERspCkz8FO1Ok97U
NICZX9+QLX/GORhKmGebF4AJJpvN/M75MMkP6vVNj9R8vxrLPSSKnFg64VHuwX0P
BjsvwJ31RhxCj8Yyt0GU5bURkKF3MXGmCb7ro8jRbOlM+BzU39iyfAofGYudgOqB
ZPIeqwAlkm1uPEOjfq4wguiEys63iCUrZ5U4fdzXkiG+C162UGvoy/iL8pY/BbmN
4S9Q7fnHFb5Cc9L2qagPdpcEQYNRHztQe7YoZokjpHs3Bpu4a6Xvcu7qDddv1ryG
rYuYFuV/NhMvCcm75HCUzvWD2qLLS1lOcozFLyXJmwt1sPGziOtPvUgM75Hufrxx
Nzc7Scx16d7VAc+10WuTZa+hGMX3Lk9+CSzWA9H4CNgsVW25P9aCu5VoCj8tfYzR
2Lk7o3lRxr2AKu1MK9og9Ar9LZdo3LO4tFw2hLDbFRgQ1D5WoKJarCTWLMSEkvmv
bvvu7cmDgPvRRCUgoJl93neCiC+9yL5HVfwtqSHbigNZEIRtLK2/vxBNWZnkYjAA
wUH28MqCAEWC9IzN5pVd0nQgzzUR/Xf2zdjBOYmwQzwAtIzdTTAGzDrXyaqcrmp6
czHNP5853whKJqxv4d008tt4LY6j06xYHgm6C3TYxyXPSJI6OkRTTvi3eeOIS0/3
mXm0EDniGEXz5CGbAPSPLaGOYwULrui7gCqFxyRox2NdM6EbqLaTOmBeUSvdqzM7
Syg6QIIvY3hqZUNSbQ8dzbScEqYWFKInSeAUBX6QyCTC9EiFV5PCzbcFYWMue4Op
OxXx3xvoVB4ms6dS5h5EVD39XGM7jC4Z94R3H+colhOG9JGAaGyV4sjgCNyXF4mC
puDD65Tbth2R3yrorAAcg+u/bTKFzDDc9qvZmNPFyfw7BYpKMTFTMsSxTpSybxrw
T6WIui8XwPWJQPEGA3NG9/lD3QyUUkQ+sH8O3Uh/NCcLHMReHdyom6Mxi868DLZr
5N+J5d3sSLnkrSTgDZqM2A98HjarLihIINvv8j0Vk3Aa/Aq/4/1AVbdtKy8htV+f
27pldyug3kwCzGyaBc7+oRs5ScT3CE0LlJ3Jegt8mAxTOh7+UhBy608C5HBXP9w+
rTwmADf+MI2fwOu9Kej/NQnlNVv8073h2IodHT+KUVVC6k8XuE1ef3uYuxQfJane
oqBpZrNekxJBHY56au9mAPNr6kcTGuxOt4F4NWLjVdLwk+skRrc+04LU1/0QGu+F
/1SIIa43Y/MtqjrUmMEzFIVDaIPb5Zf3F4y/LpqWXxOxeYklkEcdRXzkFolV1NnR
UktRi4bRp2A+o7OHxvmSjxX9M2eavdL9QxMAVuJh744T+235juAQrS3t6oWnzX9h
FSOEtmnqPj961YrXTeUEzrX8soZrAsZxKwV0s+5fkYcFNhi1pKVNvGn8bqARgBNO
j09lftq5pWv0Qaq8Y7wT2NaHtV6IfS6RJmxA7O6CfgaBox03wpw14zhyGxHHDW6o
RxGH/LLDutdg+J9kMg1571n50OQ4K3+dRlBnS0PAfKvG3+jQCBgJSWPWDr5dQuk0
kYaK4fl0m7cBJwvkmLmLQBjXxWAf1uKYIozWsnz61g1lkkHYnDl+9NjDul6T8Hqw
gK6G8uip+FDCgKfOd26HkuRHp7kdpiojtoZogSEtVkCUOMetiuTa01SRtkHiQAh8
sp4X/CH9sM46c7vDKBVQ3pwemTQPQg2yuc2ZU7PY/URhk1/hMIVY2RT83BITv1uT
/fyzJRu6PpkRI9KcRYCVdF+c4FSwLe+EzLu8LaFdCrDTFdaTBOqS3J+ZRXXseREJ
b7kO6UYTUkRMWvdUsu7/k5EoThmK4xohTX6vGwZjfaY6QBKCh3nQZm2LNUI+ar6z
eYwPyud52nqQUDI0+9hkLi6vxaVwPxCGcGWBxN2NDDUy5FFnZH/OBJ8dbuZdUxFw
/XMkvHVOBilf32csozVTNLknBGTa7M45t4V5PjddiQng670zdi+4JwJzI++GIR5m
wtGNezhUuFhyQ/4uknaTMe4nPWgo+gXlhiO9Q7rfC/RqNPrMH1p/yuSn6bDwyBhM
ByrE0ndZR0UC15eoslOpSF7O/gi7b/yljecFw4x2aWYiOiDXMy5Dn4QMK9OMtTnr
iu+3b0ntwh1TAKZg94se8Asou8kAa392DtmnzPXMb/89fesyCsuYDMm8n6B3rcFl
7TtKBs6tFJFxitxzH8h8EN0x+XAmhqAdBad6r2G1O7jLRZyb0fTqbrlZkyDPYZUH
RoUmwX9u8+576Lhrd/GyW4ZLoTceZPrpC13hD+041Z7QXZ0PbOCP7Tem3mYaIw4+
uUeb6cu6LaGu/wL9xlIRtdMFCIBVlcublq3kYtuqDDh1Lff62/0DTYxfKVdPy299
Fl/OOymElFebYFD9kwqwnf/Et9wACaMbhlKjfebYoXj1vWysjgjCGod7Ndo4424N
L1+YcbA5GhiteeKVkQWkArO3DTXdgND0zobMdru/grPjs0Anb8kSkVDtrBbWMRUY
t6J+QUfK4PMpMzH24dVb69G+x0o7j+jyc3a0kJJs7UQ3FDkUwBMKEtE6xJv3eLqn
tAvOLAGwhXrI/XdnxKaZnqiCwHK52Hx6XUDaBQg66Ajf0O8/kLo53hDWhWk5z9NH
doZLeH1G1WXLpyUcvPC0dT1TXwnKQtA5FjnGc3KRL6YmFOZc14BCmS6iUtFH4iQV
qoaZgZOoZ+pxKvZBKqXbuJ5D3opZWyJA2Zjmea/ZUMZv93N0rGmQKrmgGJmlOgFx
aA+33FuNaCIAkw9uqT0EYyuFHF0zx5YLlMGkYHux5qlkpQRDrSnzkr27MyYfgQOW
1YNWZ5xYr9e8pnE8Lk4wMHhqUWNfHkF93FxFJo2SqUnpLBbVvaIFenzL6gdIOkaB
hfBZLwSYLMJMYFJxCAXddIyjNzuwY8d+CpQHHcZvIojtfHpIpJ1OrQEgze875YkJ
tysS2HlQ4NgaQSb9CtN9BuHzjsprwHFBqBQPZIjx808ZRiofmOjb/oByPI1b/Ji4
mR7T8sJBsxh9DaV3QpBdRJSLDa0dhn612NhX25Rbvs6ygjh5lOJ08qJRlKVL5kI2
Xu0H4W4BOnV08QAuPRbtBEOeCx1a6E2CJ1pGVnDr3ybcVx+B5STHD5YR7oT2ihyh
YcOB8tRnsy0u4ew7mTB+hq17U54s35MOXOGMKurpLge4J/tyxhND8/iI/fNwd6Rl
Z11Jv9E7z7NfDm8AVh8bJPyle/aUaYcZ+Af8RVHVluIKaDxtHqcuVTu2e7SpRWDH
+5NbQcBB5wi1VQtKJzePeLogkBi5AjiNNmh6cpgXA4d3gXFrBsLgayIK6f3lWhDV
8CHQUOslCjLnZnv0EjBb/q3dKpm9C+vzyyZJ2fzRwbxfFSRPWB2iXC0gWAVPnlcF
O1VVUhZKVRUdgwqvy/wQb2//SAeWTt1i4PZrIWEZv6PeHHd3iIzxHJG0N5sgVmNm
/jXFJvYo12YLfKH680lMD3cQ6jlMlQ1gmReXZMnydxylZDXgXhaN8L3HUBIk6Ctd
pFMcTDeia++nd7CX0cj0Pe9v8RDrmSQV/Pmj1l0o9HccbBEPFdkAGnMSa4Fuo+v3
qzt9Q5IPxGF/lGQRrAr37A+8ewzD0xbnnwDYC/lVnzB376XXD86sgCZPErG5+XcO
ELjeHRMbuoVxdkga6JotqI0MLHbtFY3JCNHBcW3oeL9QjdbWXS8dqQN3K02/kzmn
iR0kwxWjlgkXA7Suej4RrUojV4WJb/ihvZCkdrHSyIP17TUJ41ylmbNkjeptloZE
VshGG1MqhZ1DHmwGCSfdOpmi/9LiJYZe7cwE+vjkhGVObYEJTYINPvisQBT1XQ/K
4/EFUnQ+hbauNracQNco1PkwcaXpgjINEraNz5T7fDf42wkmZPm4Jr7P94KKeidN
n1Dl0d6PigkW4bHd84hyHc7uY5MFmg+wihOXe/2ahqHFVN2y6dr7DpCHegrLNXfg
n+g480edvfb7PPmIsOzvj037v8CbCbRUWqEntQr8uF6To+zUTGVoceDLh/BA3oEz
97aYS+CsFWp9TXs9P2v5ty1+5Gu1/yM7M/izVBV7mKXNBUFs2Bw8W15P/H+mJ24/
nqlPxS0DjUMiaZGuuFARv669KMYyrtLsDXhXRobZol0+INlzKJWcsNt7LQEfJy8D
rGaY4/Z+nImeAZ7ggIuKFIJdjHR1VbbOj1gYMFZonKQm1WXLjiXiHY4Fv8h8RczK
jfBtvZb7BFCPLWUqfzZlyBGEJL8UumSeoYxHSskcz3om6Et+VurjuvyXf+2jNtfv
w7w9j1WwTlppBM5O41dgzGBr57B+WzNc2m3g507WTx+ZkPnaO82vZ9FbW+39lcgD
qVxFdezkd3uxWrgJNJqRV+IzxPl+2iPTelNB1YRsPhnx7+rgDhBTdaOQUQJmnEal
q+7sgj6Y1TKWD/imY/vVAum8G2L/ipBpLFhwB0SawvrGm3CK/okPANC44QkrSjdA
s+5zM/CoT/G4A4ajUyQuEJt2L7dx3JRYLEUtYpVutDh8UVcIOF4KvrckvEi8IO6J
MnBOABIwvjFbv7HslsvlwLsk/Fr98DTb78Y/8Q0G05ANEsSYzFj7ksZdiHiv9LDf
VZuTjF3AYADP8KjFP/o3qLqQp5mo7Pz57lGg89jOiK3GOGrMsSikEgcPz3ZpIBTb
wEO7cf2wuDoaCPYjFZqLY8MtpOiLQliv74z5cnQZRxiBkOL5tFbkHTiXcgrLgd5p
GJ1MhRO9mcgZ+P4o/JzkMR68zKsWDMmYcOpK/muQElace2m9gshzmmKQ1bX9OrJd
L4Gj0Mtfh7IhPZ+Ptr2QNKep7eY4Yj5vbsrjxdmkrTmfEDzOqA4cqjPQkZEvtbBv
US7rhRcyyJAOQiKMkHpCf5EMZr8B9h7NkpIyoZF01yL3UyeUoDO9Yd7rGznxW2h/
3vGgP5p3+CpF4YH4fGOhjCGor/jmRZhQEeqTSCYxXpURWo7DhuEglgLELQmemxVM
OK0Fyzixi1WTkU3FaJPDIuqxm+2hEtg6+87jGeqxv1MOkLBRy0gT+0JCQSFWvcZ5
ZRkg8kDaTHEg/ljbWdJEm6vrudZ6yC4DPwAUhZhbtv+CKQR7KKIsgG8DT0UlKIow
fHyyl1bKrIklkDxxClD4Z52HI379KhO002CF8pWoZReaZNYWZkmed2E3ErunsOHR
s+a5FOJ3ukyUIQe9RI5F7Z7JVlf23wDKCwghJoawpro+IteG+e4htIcFZ55uG2ZN
WABuKcUJoU1HZIo57kUbD60sqnPsKxIW6x4AG5Waqikl4wGkLUvhHTrUdVl5Kvv/
yxSC8yhizBJL9p49o4YJAzJUDL+MXroHQFI5gWUYS380LBvxXEh13G9hbM2WeWa/
SJfWfWqblVFu5dzhGvJAwFUd24DeXy699SvjAAb5iWxiCvfyZV3j3trXtpCVxdZe
mwcz5YvOQa9sfhu4ZI/eosdzowL0Zro+6cJAMinxpXM/VYLrGEpFW/5M/jhBMo+9
3svntJCbIGAtsKb8f8aXqEje8KkrnYTeVXLf2DeXIcUXGMfbKx0zc+PZjlNK+qBj
/GZmcFwQneH23Tk+l4dQn4plZttjv7LDese98zTZgYrCYRahLA+K48dfr8XyD61E
P7HeC3/JzbEt08SzcEnkWmTPehoDglJ1CrfbCcKIzsvFTkxR0Gwjg7bWiA+e9GIX
7zy91KQd4oJqJth63fhanpKXGj86IevmwNF4o5/g9CBg5wQVbM60W5jnMjWadAhF
LksQ6yP/SqC3jiUMx1Y3zofjS04lA0ZFhp3pYwdN7F9vKGsAJTp+Aczxum7DlhTJ
71TTFQts8whW6YQvIluLWZVKcCFLYC73MWCyL+r1GjF4FBwgeteHoxGUTHRSdMht
TlX6ovHPAUMWce3/8deASomOzg7fJkOCP6Zd0Bmp31eP8zxMTUqxuozgGBVKYNOE
nTjFfSuyaorKM5pgShC8j3gaXzXwm8wOKgErsctVPa0UffH2weFyy33Yj+jA45DS
9Hs9p70EbhHDaPwjWyVv/61DAFqluFxUKJhC8wZQyzbZsn1ZC/5P2nE74qQ0zE1S
XEROkLEeHFciijyqTiOO5d01BHYmgg8yh/e+EgoJZI4ptH818BW4NUtNkcSM5d3N
hYOhOQ4uzJIMNQILtNMXJTrR7yLilLfguy7KEgDzOnVxtFB3/+5icR4N0VFVBZMo
E8fy76cRL4nwg4U8gNYLFdDhVkvSPB3b4vBdr+QEGGncPhpxuc4uq60EXhDLiOB2
iCYtXpMd5lvmDEeSsxYCQqyBp//htrTdAfN9rPUoKFHG48cTvAEtdlh6uKKk/A8z
brz/6pw57w4WfcVz81GVwZ/XRuouzzOHXodmV1sEH2iW7vKnrq36n46p0gwlLoIt
zmq2Rbwa2HuBtOBLavDQt5DBm9mUrFRB2QGc7mWuPw7suPZMUFVvOuG7337dRM9O
CTpFoScp3O1bvGGE1a2sKZZomb8XnA9e1MM49dsY+jwnSThwAaqN+wpMc75BOZRG
bMPko5a0XK9Ir/mNaBVq5Wdwco75VBEllocKMh3rN6r5trA28yC+S2lGZpPtm67Y
ZiGfkzhA4rr6enudCLLvX8CSBUhRF7A2k/1F43gF1rY5yJwodHyWkewtCfYpF3/k
mG+d0g8Ni1wbI/1f1ZuPjqQWmejKIqUH7Hf3z0ikvdwzOiJJK9GMBzvCLZf5EcPe
8gDbw6fY8RiD26CGLTOe4nBgZ09e57Ob69WwAEewJljfPB/za/jb5MkRATPv/u7U
R11u9Ptoc9Vah0QRSerWv48UpD8dlXuTQXU94TttOdeNIK5Djm3q3aEbHP9czu3e
ezRy3psKLLkT8hznszbL+9txL3WEmFHUIYlV4CxGYeg+wyzFxFIBVI3IQnG1hFKR
faflM55mMHXcWF3Vw4aNMxGhfkZOeOwLcyaPdobcRJE6m8AlFlnbUC3NsAKHHX/8
cnqN52mYjOgteMSkBbWqBygBNIo8o8JJUO5w8EfR2KMGsUHbCxhYP0FaHju+e3XG
1iSP/4j+REAyV67p6I431AWKxgumIEpLe7W0ingUyAK7CZMQf0l1F6bUNL9a1HyX
F9r6mSxNN7V66eXUH7Gpai8QnW+WYKcNt1vnRtZVrRWyoPRhae/HT7fbXY7wJ4PH
elcL99O5+B8pUdPyS85wRhrsBa0SVt1bQJ6J+cqYVIYJZ1urizTv0uKHTb9mOo9F
obUn/hVt5YgZzzFfBdSD4HvYNNOrpJtH6/RQ8RgRjNY2XBqskThJpQoD4Phnz0X7
j0zYX+GEICxuB+VHkpK8Oo9hmdyQ7bh4rVOsO/CkmgN4geuC/bmxFCmCgb66nYQx
yS+QQCDBvu1/ALWXVcHawAk+RRAGBhoXAzjFQc/Qf5dVGKnnyyacF2TUR2oqyj49
iFR55Y9w8jganl2v8e0kGt8zSC6fEVfueGbTp5lbT1qIRQThePZiqFYbm55Hmj96
m+JkQiIgBrBtlHiJAWC3rDRciKIwJ2qYS9NhWMBhFBSdzaz97detTbsW19l83oNY
42Ayvec6JDvB4vdI5h8cLyEfFhKt5CssWz/V9vMrkox0Aw6PIDz+JMQa/oaNMFcM
7wDTBgQ2LgRUUTI8iMYH7UcqxLm1qjHZgoWOUft7r0wlQPJi6Z8jFzvP6MqjWdJN
iAqHgkD8HDIbXoOF349NiTOcdZpHVMgTK9AKILMstFHQKJGJF6reZsqmFicjN8cT
UwWNYWGbYQywIP2AfkadVqD99uWm4dTCz3elDfGVxp7KFmu+AVpIsXqorcW5okwU
t9OF0pAj2uplaaBy2NKbqvDceBdxcd3wtuh9zIu4xZcZi/Mle12Iim95ay19SYgl
+HHyuTU28vnVczQbidi6GKRU7BYvp39dSABNaHW6JWX+VPfbhhYeUieHiEei48Ah
m0i9DSToHTfIrj5bk4MUJKPheSTQoNEYVkvSMQ5TwfzznIXXvesJ7JtRanwN7p1C
+cBbTc4cbiHKPaU2OkxIEmKxsCTkWgSOeYkfzQOLWCrSB/J2ySAZ4OUxC5Cluq32
B8Ex8yOEMxMDt7k35s4uy68C78VeDrDdNWs2sPYV8x6bVVshBHZ0CiAPEKaO5dcr
quum7aHamvUo+2DrNyqjYWoaUCkzhI33FNL9tdh3ro5Ie9VGFA/q2JqjykFUzhE/
ShhrryBMi8Gib4MXYnU4CI6C7/3CFhHLltdLL4uJEXAAQetrySsbrxKe3YPW1ozi
2nwqRLG/DKMZIIWJV+XsC7fZ/IQ/Nzo4PdSJ4Xw6sShv67/Hg0V1POKQD0cWCvUz
y5+QWy6hFKe87Gv4Rnc5NTTtptco1eDY82EM6mdmjoBIMggT+3SviYYtgcpGqlHI
h6rxydEBeSVpsfhqQn2g5TQ7DqWjNBorKwE/Ny3hzkvpZli+Da9RVNj4VWXOic46
580SffcjXasbwRxSp6guRE6xkvqQ/wcx6zNAL+dX7R4tLDMoeoZt2/hh7m7vdEgy
NMQf3RevCh4WOxeXsE1ZdDgOELQjDN9Buh4dHz8wPyr9RuXmEkm6r30JWmZeO9lZ
kbEXlohWyyJu93V8+3QobV6YJrUEhNteD1l5rxBTh2kFz6QWQXB33GOHJagxM/8c
Nz4+OfHY9YAxRnfSA1Xi5YCLy8+/D9cKOkfemumsO3H74o7vhxKdNa5iA0wbIG0L
IRwoql/pLN9d3FPDkKbJQlLwtgjqfufJGmzWnRhs8ByV1YAubU+v2qoUOeSCjyf0
cIwgzLnyUh0bbSqWmDLDncBW8da9U/sb4s9CwzCOwQLCumxqvtPpTPcZLjGfHlX3
hOEC3CPAIPMX+ayoQaecPwAhILJqLbgttPvp9ooB2a2YL+A38Hvs5TlUqM2308jb
WMmT2J5iNqkfvjpi7DwdGcHsLdpLhZQJ1o7UlBfGdy7FfFXlW3HV9xu23c7aPTz6
cjscVQSq/BLS/22uYAoApdpKAKkpRQtlaRXDHmLOVJMAVTAOOO6teWLN0c8kuGPN
LBZZVJr4jHHg47FYOz6JcN5ETZsdtQh/pxJD1/Z7NdFbmwcW7zf+nCHYO39uMC5G
V95IdPtb4/W+qC4iN5vSGc/dvGf1aA3JiC3sEA2/uBqOlzg7e40NwdQoZJvtFVuZ
Ra5KKHfqfSvOcN3B+8rvUsbZRmpYy19HkxiVcGIL8ROEoUJIr9OrZBEvYd3RDDDe
TXV9Vluzm2X5j96rJ9k0+ev5w+vWuSLW5Jn8Ndgx53we9ZPspFNnDHIEEVMaDLCw
7GlGk/Rs5AT1N9HRODzUTos2UlSitJy8NAIyQdVoIJhOCApXzfG7y6ljRLN3xY3/
HysCpMEOoxkVE6h3fWurdceXjc9QTxllmLR/c++aXG8zP1e0c9qfKIW+sCSfA0id
Hw4C26U/q/BCS6sxCN5MNFuHnRoz0oNvUAdGkhCqmDaOEcxACj9QMGUKV0jY8olG
j+9ZpVoma36e6H/HF7w8uN5e/oVZDio6LhDGe9EgW00HCFpl4krydc5jk3v6CJos
TRWYkbWw9cwttLHzNTlVw5ez31IISEmqcM4N/sni+HY5OFTOx8y9Ava5oGaXrzkW
9klhUG22maRc4PTbkmY35xvKLNiPHsjLKwaUrrn+1H0Zs9pGK6pkqZaRXKqUxnaP
tM9FSBTRmPlRic2W+jdT11kSNHKH/JIpeuD1MhFLPJwOg/TFFKbDfyga8julwamf
+QcaOwnTrjgYJ7vGY156nZjdHEuQI4T614l1rQe6RrsCs3PrJeulGvts6y0EvbC5
9wDugfwmqp6OAncWdAXekWQXu6MUoNJ76Y7hiLoSQAwy3OEahubixjlVe+lIOEmr
zf3EO94eYl9oPSkzU9YfSxrlVnA8pKDVvwkAmZuguOt7amMWb+L7R/sCAcbKT5GR
hOjXtRuSRjRAmgJEYzEj82E4gt+nIrJjPw0e6IFGD1sMiWEGqUY7WjWmcK8+C9lc
OxD4qz79fmHF5Z57N6DRN+TVg6kXn+aF5wjhBsXJOhQDz/qykbpIRjh9zl6m19pn
qf9ntDwLfrVKbl7SWOj2dHRBwrLUep2tvnnp5lYzmlpoHquueZoaRKvYCApCohgb
DzX5b745vchQvkJrhbe8PwA38Ju+el5tU4SteJd+0fFHq0lCVM4Dq0aYdm+TJdsN
mX1B/CdRG/jitZZpvwl9P0NE51NVE6eDzKTvYT7hFebLu5aMdN98NTZM1ACNB27Y
x29jO34KlhxDJwdtwheOvEx2MFr7Q5MXeMBxxdcvK4TOsU4RoeZuVfHx9qKyLFSc
+MPlKEzSscXto7FMGti44oaslaybb/r4p0NYl3O+YHS4tjsCvNTdaFNd12AxW7aZ
wQxK1fS59Uy5rloZGr3cu6RGb7rYZHawkBsxG+fdKP3UHOg6xtenzei+KclEo8qw
9sQesMZ0eJFmdS+eQ9Camed6kqfxUbeq+ifsic8AzXfoPqx8H8OGzXjSn6wPbvW4
vqB5iQhKSQ+fHHsw4/jdDxsD/7TfDtcJhaZ77GlQJF34ZfX2EH1joj21wfTNt0n6
ZeQ/E0v6m+xDzt9JovrEZRJTY8vSVpYrp7RIIhmof1z8hNhHfHd0C6yK525IM41D
P3DhE8ORXZafqgF4zFh7yNrekLM2H3f7i12vBRW2HrzL20mm5QFOgVDXVOT5HLSp
+nw/H8YBPrZpjHXh+FJ3maP1ga5hodb02tEvAAJG2yduyrjW3IV+nCix3FfUlxaq
Whta/oOh6CaEzsou6Tz/mIqEDvy8xWWwd91JpT931HTi+s9BSnUfCNwDs497uLix
ePPTB0S9sax7n8vmQ3xuYdulG8hVxzcCxMxTLWFYAxOUR75e3h/KH7wPEoZMvlNz
AUuWb5j27UmXHQJan5sAQQFfeyE12xY1SUbiCK5r+N7M44ML4EZ/M2pkn6mZqBaz
hafyOw6TSdAi3SH6n1bM3GlNW67eEATUXrNl7BHPvC98yvtWpQEVev0le+Y463vr
/ZS9hKfuLpJ1sV98GGCoxZJdyiwNqjGbOi1nZ5fOyh7xntaa1GZ4nUYMglc+UeP0
WoPcm+qTbkYTehPLDp+VR4adj1gSUmp8FIaLkfHu3snUuZsKw6N3x6G24AnEshIu
9sKB8R0Mm22dMr3obyAU7BfrOxc5V5x+Fqsu1vITv7vTs7dTCn0pgw7C9nIDPxH0
JIXDqhHqk33GcKg9PbdlyVn+77Nj/e2NBdFKRuiQhfnjqNLexXMxlWT4SRWWc+4R
IS2iPeErv2udY4TvfnI318lCEw4Rm36KQ8oYVGN1hKbOz7IOhRteXN3hukUeCl5q
MZ+biVJgpCz2Av0Nnby1e4vL2SboB+OU+wozSiKmTh6niWwgE17xk5vIgLvZG5SH
drjOEAPVbxUEyvMqwtwLdG6dToNT36SocaQOEtalRZxPq5HhWn059VxOHC5jAQz/
7h/8CIsow62ybeCdRzlZzPX2SwP/Lnspb1hUdrpHCeJ3c1Br4yqInV9hY8XIOuwI
mkiJavb26TYxtn0VKf5M99TEBwJVhP/CM1vWiRxQot9FuS48T384iJmY4B7iFpWP
/nduClUK2Calmany2+c5Jy0SO0rR3/VJfVVRJS5P80+DI7nJv+Z3YCuGzF/ie42g
Uj/41HQsrA4r9fk0Tkt3DxHCK5roaKgz4emP91hfsTYGM067QQwIDBzBqM8V/9ko
vSXxOZI3unk/ZALnWmZ/wnD+tM1IriO9nvwCZHWakqPlRAaONuRSG8oqiFJIfB4T
iC2KJDP+HO52Hn7LfXhdG+jNCWfxZT3vIbKGfvIxV88InT2J+wjeJ8zFNYUQbda5
gycAUc2t/mmD4a6JLzmN5bH9uhkHMxcGZUgNCaGnj22jvqp/iAWGb9n3l/P/g/3r
WEzx8IaVgyz/G0Rx18M5ZbQ0iTMUu6oIpxYaCtkrfPw5LmUd6VatYXkklVKZ5gz6
akZV1Jqf1ArcekW1r93l5C1RjUYZ0mdNFNaRCGzdJhjQ4z0MInejGFODDqLk7De0
1aNnISPrY7nVJ4jfFb/3TaWsMHE0dPYJn+F9ps/ACrli6WKphkzYxvexV23F4Thp
+JPOY9p864sjnR15ppU/LNLNRX2yzbqoy36uwcf/gbjyOeNfjuTYJ2KyZDHGxhTz
AjABxptjmK5DOQErFYlFWby9GEGP+zV1VFc0KNbwdYGTDLtSdKF6iygXqvNSi8go
TQpbQEErYBuvP+oagd+LVCeSarVMiag6JVD7GudLoxpAhPE9gpmrHbLxi8QwU1Ux
tCuCf7KmT3GAQoUKfBpBFOtxsPLIOd38gRtK8xoVDpoFnB+2GrWQ01lQ1oQu7JgR
KtXzcrpjrrZ3l05NioXJj/Eo/9DTz45YhF6q8Ms+QzPnaPmGEa67pJ0Af0frpOfX
91PES8OAh1iza7ohHpQu1M/tcjWSTDChHffvb5+zLG6fmBvPbt+H0Ldgk8y7nSrg
5de9ot/5PzYKr+keJL9Pk9NSQwL3CaZPIZ5bkJPJ0/T5OIzR4Q0vinZ7J/aeXFIW
ms+L9K0RwiP5GQQxyvpmZDxz8iD0zLGRuNMgZR2Ss/OZWzkNGKvCY3GJeLWBxhnc
hF9ldcaolDZfY7adhZAD0ehn+XJkcCXKYCCgCd5/LU6UGO5zUCNRu+/viEkfsnbo
xOVzApHfv/9g9LfM/LfEDWvVl+lTbvQzoBsgUAQhhEqdvO27T4J3RTLSokAPQuhB
UXvG4bSYIq/alUfJeMU72ZIX1WOsUidwb24MOm4OCulX4F8jYOGATk0DFidNXshe
DaHHoJ78x/lwTpSOqbXofjj5lfYDN6if6R5pc9CUgs+qgvLzHv+Bi6u8QoAd7fQr
S5b34J0e1E3poWEkpgxi0EDloKrLxzU0pBoe+5rwMvH0ibCsEaJpdQU0klldKsVq
C426fdc8qR6FrJAHVz23XJIach/uumHOXwfkkawF5oSXnIVDBGCAwP3jJpHNRLUJ
Ywjl2FBM8X4y0SO45buLPqyHHP+DYdpgFxe8LQC6Uu55cLILRPQhFcecuchbqXRI
X6Cj5HjSXc44WI1SFj6fyge4Rk0C04D3hhnqyjJwwzSCaxiybqOJhibVa/eRKyK9
LRg5WjvSqeoUoUfSMC6w079mjWMw5Zm0I/bwbjHUW211frLT+BU2fwcKztSG0vdn
mCKtMZRbTz+HFjngqowJD5m0hCRz//E6VmesEaEH73oQRREsJiySXFm583gX7UBM
UYfoxdCE5ukERnoMQtQNyptozLJjXXA36bqmb0khlFKBmWpugtTnZTy021a1sMkF
OTa9KPuZiL+WSNDcuIfkNBXamDlGtI1Uswx0nnE39f/8smbgvYh7xi5QqaCGnBcX
IDatYC33ZZ4SoCn4s80timzYiD2H7KuGEljPgkYuYBj3wz6CpxsYFglv1vn85e7d
Fq/uKiwCufb1pj+WopJUCtTeysxvSP62lVGLTXWzVygoi4hkpKDvHY5EoKwL4bfL
G1F++de6R0s4Y0sxaMSi25NlZCLu6doacTpDdtJBf57diop47blwmp1KGOnG3G9a
lGToi6NIJCP+evwtyiVi0wWhfHS23av3xWONnSqFPX79QG8GZhZ8vMdBtFdYogNV
iskPXh6ry31QCfxLT1Ku9mlFX0UjNmgzOY3C5ni5wlrU4eon4JP7DOXReO7ErguX
wt+WK7ONbU68dweuGOG0hRP9sCQwMyFHQqEB6roh9exDxHWHLq+enH3tE1YbJ1Ke
fOWpH455i+kQWRf8SBLgSMJwAMNcQafrhFTfhWhUWWzTtbA+rO7JTs3GJITbSZyQ
YaXlIMuSL2o81dZMmt+ql7kKFuSk0lt1v6Ogga5wJVhiDYxHNbGubXW3voa0Kwy7
6tOH2xDKBDGJS+/IBZF4H6GUexjthnLJCVu/UHnc3KVxZVTdQ1tOVFuCoRdYT6KW
oU5zMnQLDrYNsQ/MgyCQ0oMryIPk6nPr4JKzCRMNDSJ04uVO7oFLK/Ef2WZMZfoP
brMHsEcnbU5pm3EKNkW2zRL8l9spjHBYpmKTOr92ATek+LiqcKiV1nav+olJkjNB
tOigky4MDyTQUj6nH6klOezzYvgxDdszQfb8bGSh8FOtjM4RQ0HNnasg85E3R2Ui
XqX4tagSUC2+6Dwi8mT+A3FZtuanJOOFj4B0vZRxcZVJQ1FDAXj2NFEJTuxwCrvA
zM4bfNwuFikML4q2kCA9cNmLI0FoKIRrnfSeMuw/KusZufyKt5jo6EU0NQW4TjbO
oW/+84vkgXmV4yr5osQA5FnOefnW2z3sIp5Q1hGnHpL5iXSVLEfT5VcjUzutr3XF
neTyGkRhkBpzjqc4UaPANijRbI1omWQxfQwX1JygRGWl4IZVrEFIbdqMIuokQ3LF
8htXovK2uSHEoEL9/NrcRO/oYHKQqx1OIXiAWFBSXq4LOM3TlGr7mt/kJ3+n0+fg
/8aeicvR/cwvygXXLh8QytQLHDbjk1dU4ePabZPrLly+kA2l2AOYyaaCFEXz4EKs
ed58XiLDxCOWKhduRfIo0n6DGmLuwJU1t3ziXa3/lBAhC16vng7aDF3xmfdIG0hq
I9k/sOdKwZVfbTWaDvQRg7/04O0VHELoxr0AxJZxoionIJGa4e7WCwsVXLYes92b
NFO6u9vOCCViZeVkKXfgDt2SGYlr+VzGqPSYUI3EdRHhLTEbYbyoh1VNWhLQeIH/
OaXMBimQIeWIv14kHbuBw2HhDeekCloe/2CwiAe193u/WgDyyevmI478eC7QjJiR
cKZTwIkQUe0KEOVXYhS8RqBNwK46751Hdueaup5IDAR08IHS8xmoezbLKvLmAfuM
bNf+DUSlTfVA3e3B3cSU60Vra0KC7045ze16wOeRkdetW5W4OGWi2L+XEjo5B9Ez
jwm5WD5927yl1xLXR4amQ9ODZskjkzy/sqkd4N4IK4MNGhv4ihxLvT8OzESwJZfp
cmR4nEm7Mo1v92mJnHcI1H998c76cj1HrmMJu+RjX6AzuZnHxoeoRVvnqML9CSAH
YlV9qQTruK9HOF0IdJVkI6rTukSDwI/YmxKUOLcwGXf+W3ix6T6oWzi6JrAJU/f4
Sf8yefo9aO3omhNDyW8kU3gfwuD8GCcnT9U3YCqbdGgv+wiCdpVKh6SLVv4f04by
9wCb/64byx1+4YFIVeGfQNZx27wk+Zqp77XU7JSRaRW7aBsA+bALNef7Pv1LyRU6
JTMm59stZTUkwBXKItlSgbeFOvPwOMOlCKJeuDHvt5XsueCrFDTzxZssnyn1szJH
zNpjv/CHVci72PDK6fMKmAIPn9L2QekFuMwIGeMXCNjVValRJNvOAtMwk7C7Mav6
ayGE9MBBoovPSgZku6bEsN4vZawOu0ONs5znrf42jDPFivXooUYr7uBwfyGEIRRs
TjQmH99FWV/KSqy8iTPCiCK2fQt07nAtclc3aVFBfFLeppjHUSIGvTxSWLwfSTcy
13jpJV1nDE1IGldhO43HTWQnFH4q3cu0A9MjTqF9qdsXb6SU2o4bItkmMSa5sWM4
uVcSvz5yXZUY86sbGsJTbA+Rg56bf3CCGhmbc0+s9MiKNyqDz9YMgxDdlGQy0U3P
9H5XNEPENn1APAeW/eqio5BjgYIZmy0HqdK+bwrBRA0iNquNWUXolQUFefVG1cuY
2pk0+kGGAnMiqOTLdUNPmwREO3IJUE1wmwBSuZpjYauaiy2vfjqBgmAX/qkLIJCC
8rd4EsuNc+/rewWp3ebzEd9BOw92DmXvoKr5rp993ofw27GXWmw6lTE4cUn+nKwY
z+hRA6ZG83RqLMyv+S66Nag23n+1MtPIr2joYMQzAi7QxHYDCCo6HB7ymhWFelLk
p3UNrC680FKz58hrCxhC1AtOJfV0Ww6DUkgdvRDsMSfoduQmk8PyFuzh690ZcIHn
EiqRFQyIyCvaaLqN7Ge6zQPvjnVL2PHJTtF3AkEhnopgcZVVyPVVtCNP5TpFOw6y
YGLgZOUSj94NvKUe0XtUimc+6feTfiNbTPhc1KcMAMqj+cq3QaLLWwZiu/8NZwso
LKk8k/OynBsZIFyu0Kv822yetziOFyZHHMg0kEUus54mkAkOt+Ey5B+OkmH4ONAN
2Dr2qcdgCLuf4SjK9NgGQVnFbBgsetgvvvemc4z5mjO0imjwQ0qeTfuQnRLhSZYJ
Sbw8fNt19j/a2uyVv35WBdzR4FmdJQPqRkwW7NdCf7eYppf8J/89RTVpsQWzQGQ9
6qkLQl2yl9zUv4ScuAu8/BB7OsRKAwgelNcXSovkYQ0jWZ1MoD6iyR1sVD/JAxSJ
kka1FfnAEc+f9MAP1t3//wBGykxracwn2QsQGOPEKjCVejFULXN76RtT4eluSVM0
gl21k3IpnfCXmJ8fSt2Yj8mqj9mIXnnKhpA+xDCB071zxxrB7owYj45dtkuU195w
VRpKxW7uJixpNzYTX7ohxffpHWL+wG/X6ht+sAiUUYgeiGW9zvoo8y/EV0hy9o+Y
GbbEzxDS5tJohlEORDkG6Z8kAuxYHZjIQPHozvF5fOAnsqSK1T1v7+NU8MMOfc2e
ewHuDEgyrWcGhJ8Upwd8/wbe6ZAvRRj39qwdmngtU3LWGTGNPYe6M13eQHO0Qk1N
0ToN8FDBOI7Uta47RvyIpB3C0uoyTR8F1KAoPfITX36zF0fMGiuOGu5jK3kiIrx7
KrAiStr2Ul4oWHD5CTfDFsQpCJAzgAtwXFngkCiZ4UnWzvp7v3dw5coH6XzqOBYy
sLn1KvK89Nvp1qy//cTE+ixPvG0UyvounA4Fd54jhCErDAiH9PxHDd7Y0cWoyaPH
7Dv9nehmzjjGJOmLBhrIiSm+wfxNPbsjxY3KPVuGQ5LgrGOLXW1ExPawOruLIjLM
9C/5hd3cm4zqESTK7FbQDLk9Lbz0WAQfHdMvXR5Vu8ne+gNNFX3HKg3vbLVgtc5v
B/Emo2Qz6XHfkU2O8dBgC6u5kWCerhdxun2aoif1jVuBoierO08SJ5Fh0OaQFNim
MQ9pkga/yWZGksoTRcqxM5ONd04i4521b/pnhzs75eetuNDA23fYcvI+XgqaPCS8
TKzk8k5IQT4IV/+gsPjIFTsYjLAPEjfcocodhhfHRkAoLG9JCPswFknXEKSOXKRc
Wgn6r9GxnxEfiWpU809MhsiwMXZ5ak/bBHt5NAS4axeuT1L3pEGgfs+rJgtnLg0p
tdFZUr/ct3XvEYDYs1sf47SvaC0uKYTpaGnIEwifdbrlzd3VIk2uVqgQpUTp81c6
EEZnru9kso8w4qPSq/z2u2xnHcT4Z8VP7f4PYuKUmVqbBF1KAZmMKqe32dlXHO0S
udkBEEjuTsSJDkzh5cUIqk8fmoI9ySdKx2ANfGGCFabq5u9lUPS0dmETUeHz4/ke
bz9OPckmJiia+AQK0LBRxlyDmZKAGzjnO7HVARAr1FGl4oaT35I2CqTTcxm5Zmyl
7IwHQiADODuqZhs3M3X9apUWWBbhe+VTDEck2uYVWmbv4P6jvY1AoDPP0/9v48PV
Fdi5hKkIxa5/k0x9rIoWS7G6+ZKq5nBp7+nedNHsUHq/yfNpkPebXeFfZSrpmg8f
2AQ0v238xSv9+E4xdqBxEwXPDqeEt21qRMvtKWF0/+DXl+YjHX+klb4IyepqbFd6
lX1gc8oeYOlI8qXnKbs3bx1HS8hPs53XqEA5tBFgQeEeXoY+oq+xEnskYGYBAN/U
gw5lZS2yzLukP9kMs4l2BB5pmNy+EPJgUqA2M85zMaI37YIe2QCb3+m/Q0ZUMzj6
ORtp/de8FehRiegdzyz6jO+IZkNYoRZe+0uZBGQ5+NC+ZCZhLmkZkk9kCKRJHN7n
4bG5fuozuzJg76QGKa39/xH6NOpjCbEnGgQJcQmdBKlPbwYLAGMFknGL+o9Y311F
G+hslj1Ay7fCKm4JSn+mrtDMs4cfEdBs5amSMeHI3MA4pDsPISJlkT6oCTwY88OE
YGKQsA2QqgquBg53+oKyLO8GHa4jYIdwBI1Rqo1o5bFFJj+71yN93wR8Tq+ZDd65
01ngmmuraai6C/GtAmx9PuTZvdoE2KfpGdRvdW1FLPBPA+9sTapyc9VzC2F1YSrR
r/y3kyvAhyyBFnBttL42sYf/sSc11n8OT6CADrbPKgkw1GKON4qumzJTXNbtNRWn
xhwSUtZjWAMLKxvpHiYPnp0x4oaar4Br5ip50ERcq94Ptmi3qjTLmmruvzubqSPf
jHi+ECeRe3+vcoilra2G/sQEI/O43L1PGBHTdR6mPM3MX76xcVnJgEwVddUYL4dQ
BiDkEfMV6Z+yvRj3DD8AxVzXlDL3I/rJQsFF2nwy4/1cGPPFwfMZB3psCP/7HxdW
bPGJy3PD2qB+0Rs625rg2mnQ1vL+4+euzsTofXG77qR7+dDEcumFOk2CxoC4YTzr
iOY/83TN31t1Ey+xyBn1zkrqA7EILAe2QHUZuuyb5SbUOxp/NSP5UBIh7AhRJ64w
DFsSeySQ1dqNbxrp0N23QYOf5XLQrGSh4c7N8WOdBUzlRnVCNJbD/OJs9MnB2omN
Wpjb1b7sHTbvIatzJo6gVq9+CWScEKtI8e6OdorjuJABc/tTwuhlITonDt3dvcUH
HQYQNrcN8Rgv+n7Zt3AMy5iKs8q48juNJs+2xE+Y0oIbQ1gguD8JwY2//51r0mKp
p+iBvv2aaeIcaM6/z0a3QOKLwKEYiTXWMj6xOvr3ldNbFUUhe72Egab1PjZbQBLH
oI7UCj13wQtgx0SP3H5dII73uQjkQVpewFwaBMEsw4slfseutGTGJWbcU99ZZF6T
580ydmK8Wgr+VQvguwPjANLhRPI5HYDxKG1FALST28RLMOidm2IyyYOUkXNfBe7D
LToGaIotYPsfZYzy1nTLuS9sCmcmK9CJcdOgclCpYUQqUqMT1Q8diX7jb+uZIJFU
0cw7KghRYlU8nUmIi3lSVkgxtKW25y87cd8Ia3xLlYIRrtL1YewCisGwxdT68rFO
y+9YFwx/utSlzEKy+d94FBqrk/xRMjQ62ZrA8LCRH0xDkIymdPNLE2n5nkEaX1/s
xp+0VS0DR3Yj1YUkpYiz82n26o9T2CRlmyOKB3yb+xo5ux+uWu4aFMKcrAGS9nrL
06BE157tz9z2Mj5cRVWcTxRk8sCl/yIe/BEwDKpS7Kc0bCxlaqcBuinq55u5+1nr
YGZURk7i2vWkTYWSYij/4NCpXG+cxQtqay8dlMmbi6xfsAToE7ADUIzHrOE1QMNZ
Jsx5ugvega63N/QByrepyiN8mEphOS1hWnmiwmaJJRMjO2lyID72n7bTxjx8TC7+
wbIdKU2mUkWmrlQlALZ5eRfj3bND+qMCohTRmIlPIWH9HfFWOs7xA7BgZsnbpqIu
6+7wXDjWXPI424SDziKAJzKmnY+uuEh1Z/6PhsWhKXWCEexXcwNtlGiI48WSqn3u
cKxg8PRqGJDqlesLK4VEEIbPA/2SWkEf2Nw6k3zc+piHRcjkbgeGmRte7Bk6ZLSd
WiHKoijMtwiP1om6Bor39KyGciHyQaQcLaEVE5+c5kKdE2i+AhCULnS+w02jlhiD
npPzZFw52UTmNFGfL6XJ2c6W5uooctY7SenqQM39hEEvcH5EQ10ddSPuDRv0Vkgc
jOjZwRbWZHHMTvuwwqzDKJ540E91RaZviS/+gk0CKINzmGcODdXk3BFTBB+C0yal
4YKLUn/JTBJOe33/MhXvBl2Hw/jp6MUg+5rlnJEdjCZWcQGkcolp9tPR8sdBSlPg
lH/NhRy3xbVRWnmLgOJcd/Woh3Vfxljlqc+FOkw46dFCj9IyeMSyS73wMy4UWIQn
t453bH+PNiLrxbOakQjlIEdg4fZiJ8NJ3WQi/XBdeIM0KV1Nc7bIOBALMXzdmIp7
EP7R323eO3MLGwcyrId+rOHx01l4Fa1ZhGFH34+JdEoZjiBu8yffsu1uCbNjqcSw
8hZNZ/Br8wQJtX1Kf6SlXeUD2pKo8HHSpT/3JW8y3l3AwHGVBd5U08xftPv8PVzC
GXrqESbDF6GP+y5CFbANLqde3r3vBYN5qGSDhzFqEOFRkrKzdxyZNMfuZ0vIUMLr
b7unEfKQruIhvSQ50xP79ZustVMTi6R4kPQRfH5BzFvcCKGF55RN8irxD7o2Vpbr
eTkuuBY2D4iGvngxOvBkDQDECq7JA+iHP8c8ZhQGpBnhKY6PelESqQuN8biJt4/B
hmqFzu6F7nC0dB2trjdi+8qze54Nt5ijZlw7ZdyHRJU45JBDpDuUJ+v9HFCaRwCD
d4LYQm7R+oB0lbj0njgE49/mWFL8eV+AaR4FyizYTvk2GQJkNbrK0jq9XOezKpLX
ShWebE9rqk9uPZ2p3k57pqoY4CnnYR4xTlCBjvntwDwLfpMextEmTyBl+h7G8L4r
U3UPIPkyu3t4DoPExuw0j5+fZ3nmsjkTjqDQvyTjhVO/ePhQNXVaMps+YCCoBQtD
4ORbQz3mKRWPI6sZSwOfDyiIbVgI1LSQPjCPbcCqLYqSFHTsRzpXjDDa+XWExt2s
ogidEwKHHK+4GlQ+QUoSw0GnLYoMUaSRzw2dO6MpIltmuiHVGHjfMIHG8cUtSnwJ
KNeABummdRsduW2WM/nqtThVVrCr5AM/cQSSwAPVFyTgT0GZLitISN8ekKEEv6mU
rxtT8T33gcUenLezXbjl5C8hNLofdrrEMLqkzxQW/0s7GP8vUgzhbgCJ1rcgl5fE
Aj5uPBDvH0GkhWPqq+xQYw9sXQO3l0vhM1drlsYbLZElbbYAumDHXXR9knwK1GVo
wFBWBubw7xnWydkgbijXuKdScAS9FfZIQ9aWZwrWsBjP5R9ivziviaE1hRtQJiRb
lU7bWtlLNrcb6/864Td/kj6dBWAl53n+nNFmPVYJtGFe7+A4iVd049gVwkSiVqTN
RRBGon8ZtBmszeXR/l2ZI5wLIEKuWJTD+m1lqcitqjQces9sUsJoZWvGC2QYi49R
x7uUvZjv2ovWTBq45P69yNB/Ok0P2Kini5ICvydD8ntGU3C/KxaIdfMH4bd8J3Dq
z3VQR2rRGYBAe1GPWCCOVouWRq34y0B5wOh2scxumAA07fMq9I4XHySDx1hiZM5+
K8dLbRvV2B4gU1KCmEoSXAKQ6D1CqS36Xdm2C9gFvjqYcULvthNOJkmlPwDfCnSM
PY2sqLWHXnu13WUhRaIVcleIF2QhHrkz4bzg0tcgqiepXqGyi60W+jOoR1hiGOZo
84PVizwK7BI+bp+99csUu95DT6SVN8YsUglySJMxOX1H4oKKIXG4D7qUj2TnFcyu
MM7B61KJmkjPOilKBpyCZzwCayU8MIuEfD+MKvpiE5pveFB02YJ+72iAYZ06/yOu
IXccZdJd5eY3s1cRMgtc0I48YrQPpnqikUCFJJIyUlSoJy2iP7clDqsZRokeFgeV
FeoF6h/1PP4pZl2SC5HzNQkcGqMtJRs6TR5Xo47XXm55Qs1611rClRTgKcQuwhyB
9w/zySY4KSRs1SvOt4affMq7nmKaYsneHHqhd4aEKnTHmTIlYNsk1FaCPpKEcuJu
kaxFFmSNPwwqIrWMh3IRmeoNEUFY4Ifh/d5dgEKRwZTU0sQPe8/f2P7eK8k2Y/gZ
prNDCzdwl2oXdSsqFo5L1lterYweR92juNcxuQZgb9P3lS3hLXCvXyH1FGbeNWvS
9eWOXgBkD339LkeUscRK8Hi8X4QGp+r/WHaMja0zsaxQIQr+YDaPWIFxDZ+Bt3E3
A/NGmFyvW4pmajcsJtEg0sqWKFlGwH2/Twlzj/JHqOmbkLkKScaX/vOqTdQcCKQE
ApDtGhqlAJ8QqoO4NXgQZIXTAZBQbRbYz/53jNsZFyScwy9uXTBxblgTELMP7gGH
bWFk9erJCSjbz24q5ANjIgsRhoF/oq0Co+dM5RMX0HJ1ePSpyUqZuuJarpayKaxb
pE0NyKshFL9E0Xe1KkBSR8p1zP7ClpOGNYiUUFloSBa1pqoYKaVfL0oeBc+CCWGE
iNrzXIBSVrwtTl4FJdrQzRHqd8m42O0qjF2FAtCjkq6Wxmdcf946bjx/++GVkOpx
NFZRVOj7YsmWLl/fhYn07ATLhxJYbd4by/BbGviVFaf9c1SdBUdWPsnbKdYf8n5c
tTb+qrOJH8vIxTTT8w5PcDkFr6lrmvYmag/HC2NacZ4Cl0yfT28fVqMuNV0Quq+Q
sO3M0L2VHOrMVUudFXCUfFBSti6WTiAZBr0hCGq45GAKXJNYA4r7SDTyX3OHM7Vp
fK+HFTGgnq6lLDwNYXI+rSK6fRKaFetmoNaIiR5RJSPBk8nnX0cL4FUY+VgVtdjj
TgC15vFJQxFgUo/IkYu6ZGY3Bp0EyHJ9hPsXfMvvNMBdCQeZQ5gyMaLIrMmg0nmt
Alof2qMX93thMb6aryBu0CeL0uf+10V4ARtGkRP7m9X3dgd8vG00oX3S43R0Fcmx
+1zRMUfmiFqNJXlV96l5DkonYPQ5m5iR/jt29zo03Rlv5TuEVGd2W6esSKwCHvcj
vveBbhwsMt2C/YMnrd1/LK5Sv6eFnUGNSLHN/6yizYZb9/0CJ4ZeFp2hBzOmgHt9
eN8A3lQG7+RSU8CuMh2Btx6Jrq8sui+596hOekq9pyfVD9/11DveWXvd50Z/Jq0k
MLKBwjbiz/HTET/tdzhwyhVFzSsWlFnXxTXAQ769rhZeZjz3Be1Loe1lqoAjQxnW
6Gt7Pau0NVj03iKyl8jVWYv6rKMGbzD00NOdvHX9lXGWEHQmTxAyuQx8oPO/QiD9
LnpJxZaaP/LGnxdY0xaGkpe/osY0rcoNY0NwFNyPM9fKJQvCO9jRUZVKk/QkRX8a
zjOrcSq0kysSQemORHyY8XOcrovSHqidCyOFHOkESSMHMXYCmMEvJ7XiQYWYuwzO
B1tqtEi7G1/ZT3owCGeGUjunstaFZzKKo4+NS417B8nw9s8MK8FY+0FyNhrogTzb
lG89bMV/sBb88w+XLl/BXbSVx17jVHz+4CBxmMNXT4Gp5aw+pfcXEaVY7lqCBZtI
NshbJwYFx9lEBl7UcDsi0AfJyBmgrVH9h82fFXbVJhjTKgONvE4FRKd+IgTJx39O
PNztKo7/8ijI0jxwvKmyDVHytPBZYPMVS/YwPhnkm66JB9MEcd5PddZD3YdYd3hF
GpeFdZ9uxVv1UjZxbs+EZ7vdg+mTVreIZ3HRG+CuY9CM0u2aza2LlghRp845JJUN
pvJUOX8pJFS9roe8xa09e609UkbLq8xuyNVxZL3tGOua/wwc/fOhdpq3JtnEJ1in
+fTBRtHJMKjmV84IIKRNbeyse4PsVgyp5v4QZbrPk/9YrojPEYXEHGG2h6kAVooM
ezul4Qtd4ZeiePfsBp0KHBH7smpWSadRopY0v8aZb93qIYW8dr+NXcQOGieG6QUa
OXxZx2Knf/nhMTxUhM17H89Alhc7UQVtndRQLgfTocEwCF9cPdTo4+oNmzM+S70q
0Un2tzS4xN+h3NjehrMzPAWyPqWLa9LzIoJ747GbiXfMO+XF/1wV5pHu4WzO3eQy
XwWtmP4ycKViqm8d0bp3DiFUsWT7yGRJ5Ajsxlg7/0Fszq7yns0ZhtFunKN1EBns
xPa3BwlReTHo4ETie//+t1cPuhv8Qephv1MZKdNeLpI9Dk4Q3NPRvmEphXbBRmyL
uY1/75FYoj9zeScsOCDndMpBcr7tDDJIlWDgaOTiNgSGZ3Xt2FG5niyyWdcWi6mL
RR6cflmr+9br2xjzaQeKQf2520ZnjwSkysrmquLorwxUIA5ZyBdFNdIOJvlYJ/io
1xq4YKUqt8NXS9j9kmWOORfY0iZoe6itfUU4Eq8Howv/HM+C7js7T6Iy8qTmzWfz
JGkZTLpHWBoJze0XPGyIiO8d9rCBDHVTDK52Hu5ajTayEjQigZxz/pjTGC90jAlA
DuU1S4yLcm1+p3SbgZQIDWHjzKY2N7O4BX+1BSFlRcbvzR3auFPWCQoSC9+7A8L/
FmMSuT0w4EmlDHT4t5WX+EXGlABzt9uyjVtR7qxbohOSHpIhjl3D5YmsQS38sAvS
/Ub2iFj2MjhLoMYnWNu7uwctGLGbU67gavskacgWiUyDXyc2SD6E1ALqueVmfkI0
1ZGDy3tavUZIZAO2vNRcCiYPjX0F4M6spAb33gl0kXkVT/H10Qnl+RHjWHl85fE+
mkJRdEMkXf2ewDutuLTzbjJtWznMxbFv/r3u+Md/HyXUgVfUXk0oW7pO93QtyNAj
6Spufk7kflRm2SYic4ushqlD5hprz3NHhwirVESAqzg4EroDqvmcGWYidh4OUguk
xmL9OfB28lM5isEvphmKp7b5Is5pnl3SMG7bbBW8E4pyY59MKqd9/h6GtnPpF7Ne
cOF8vb1SSbBOzhBz2B2o7upOYT/kUTMjXL7qqRAotN+jrib1jYvForj0579zV4nQ
kJCS7un4IiKzNhU3Jo8w5dtVQJkIvV7S0FAZ5FViKP5VoCW6QmsGsad+nnczuXBU
n5YTyRMnEfpJk5B/LOdPnQoay6Voe6G8VOWhbY7r0SM4l3Fx+nS6dyEBhChFWgUD
fVi7eUpqlm3xevnmSn0l1dD/vgfo8swJoSDpNAwvOnZcyUk3IMWwJfPjONE9Sfzb
bYiV+MpE3k8TC25Gps7lUgBqxniyAK6tKq/am6zZj9gkghaCd7WPZdHDvD80zy4s
jJ8ii09PROrQShNxDfPE8IfR5Au7eSDyb4RyJ8MGiL+bXp0W2trbetvg5pRitGMZ
0JyO6b+6vw1LI1V+7Waf38HrzJIdRlyzW785QG/oF3Yd4eZwjI5NRvMJtbkAbJM+
5bWw4yw6w6ZA2PZzcEX8ClJheiNf8vfEtS0bz3WqmUF28Kmz9VYbZ4jRQcYj28yd
Gn9HqypdjuilyXduyNoZZ2fttVYb/rFUdqM8vRVn5d3QHrleQnEXTqRS8LCUtkvn
yxqjMN1nAKp4nkaAVbfwmmC7EuiZ1qzQEMnrVQmlESXoMbGbjPSIqrOj5beUrC09
lbVNkO8KmmioH2I6mKJ28puo5j4F3ZFzoMMRSEaUkjE14Wu4XtcOTM8OtDmmq5UX
jm6LB4lQhxRlzhTS/0dgMh9IyHh5TNxGnbUIQ4K/mXsxMUv7tFif+SUrf4VD7blX
y/mQQ9qz55hcRvVku/Quy5PUQRM9n9S5kPCrdQrlRLwqiO3h7fjKBQ9wXPDnN403
AWrXirjA4ZVEHyVD9na84Z6TigUsuAIlxyUxpQ/5okDPGfotH2RfEKj73uTK49sz
Wb2I3jSnvlFe6GWvt3dVHlVOMxikwyo8kAnOcxASviIOq5glXbSI336sGl1D+Sh6
5avJy2AukOZdJyqttpfwrmwcamuxkmtysCKsJt7K9aQa/JC1Paiw01tLnZSSaITe
qoIxfmAZ5BZI+FjcdflVCDrS5UG9SYfpZas6hfVC7KuD3ZJGB6zBBwZ7w2ogjjg9
brpsOrLSJHHYxnSzetKr4bjNhg1g66uG6fOD5+vmegeFUr9SLYAu1gSlvpK0j1Wy
Y+I3hQ090qUiWx5op/9GP6qdRP6M9/QhiGWKDByge2ARAHCDzE9d/sz4A+5ozjd1
MU0FwrYutyAswLp0KLvsAlDkTbpm6ijJi6fYWx4SwEphgehcbXp/J05LiIqYJqMu
DHxU3xL4tq653S6IF8/5sNxYYyIl1HjeKO2AFtA/9ROYV8xCQWljv/SAbJ7hjs9s
1NsqJqD4it3T1OR7hQrzs/klWqsVwNuWch9TiGNgcXM1FPRXO3azEQ0y6A4rUPsS
LpRIKS9xv2vMwcYROF6118Gumrhnj3XyPJQWOSnFhwkhtvUE4fooUKHnmPVifnYs
hEXbqS1URs0bfzVUQ6S0ieD2ZrxXv5Gn4duSBdFGSBBQ0t6WV3RtpLP9f7Sk6UNw
ORW26LMu8LffAcSWy/ZJf2YzyI6JoHb8JZMKohSSiEw/vpvYuKgdhTJnVKbJwTVK
VlJgJ5bzqQDS4d3IhSX+I6/YzCC+EhvmM/Jj1KJXf4CphqMrP8A8V1ZMQprHdMHo
i9QX8UOOnp0HVMPYJ+VyXEQAmQWj4NmZUWO/89gL7pkbg7VHKrxT2q5JM6o/WG8T
pw6dqt2oOliHuFYAuY/CIkTNG3cyQgnq1Yev0+0tWOpYKhfdvMkOhLTiOW3EFyUS
0MJpEiBH1cmDufYJziAw2PtlKAun7vIS3mbb2eRkt6EDMafBM/3xbgCyHPaBOYEl
Zf0Jt2FR1w6028or7GjLeS35aYo4lIt6WX4YOoIcYq+FCuD/2LyF89V0s4bTK6Dt
cx/6rGkWEqqSIUy4OUHUndJ7ZtL02u0CfLdZnJB6i88E7PIroBvPzTqNABHa4xix
AAsjqdjCrJQ5pNy/vQjP3vFCb9yDTtvGjtNvtxj2CrB0y1jknyFhQRMX6BX8x9fQ
7mLb1LqJs+OT5d3Xhnjx28B52RXf7mulSJNrL/6PVWnDDrXLbx39HOeWqO4l808g
EYKiLntKAsNQ9GD7ZbJWsoxkCTqgNJZpEyLbcKRwGIBwXShhgAKecm6ihSuCij+S
EcWhX7U2VCqECbbQriU3UBOKWayIymgVgCbAHPxuer0nX01vWmFngNGHWgt/wsEf
A6wowq7qFdjIfPDpwW+grT7yf20ohLFTKcYOMtDhqL3OWJpehwk4foRZ3sQJUfMQ
hqlPZQczoIZZgQF96xX0lc/JR+wbtyOT1OKVS26oMHnT7BZuC7HXknM2kbIZhDQc
lcysYXfpm5y1hhQS6jlt4HQEUMun6mciFKe6/aVm8OeARZe990HPE2YLfE8Ekr1O
xIfgxZeAF/Xyv0HRshtePECuco+LiaERXUn19aqaWHKaOtBTYRw/2OPkj8WwiVcA
1CtL45YQp/FYfZy5aUC2m5eXt/iSops3VJHcD9xr4rlUNxLxMKWRyKow8/O3F2DO
tv5KAcwY/Lrekk1UbLYxIGlTkmhOZytUmlaiUaDy/zzViyzag43of8mnmhaum7pg
OFHdIakhCM8BQlDeEaBN2PJ2t0jhT05c5V4oWB8+0dHxE2DuwbduQ34FuAGG06JL
e2pGGLu+Y3pvONPI1Vsse4I4UlAzuJ6rcA60iTYbBDykFV01ZccAeUMxIz//qcqe
J5ZUMGRFibqRBw7dTNN2EIkA9gv3XYdKqdSnYRplZ0uF1SW7+miN2N+WNnSeim4n
aS+OI7U3CCu4sCKrk+yBi9f3tY6QjZcA1REugsmled8BhmhZEct7LYDoCopvlnQ4
AbtLP0kKw4ON2OMPj2YhnAZrK+8680zxZL3ANbMkCcR2VE2J340CMAQu8WD0PhoD
gIqk0kNNEv6DyBQB76BCo9IvWtqSW8SdGo7nPlltATxhpssUjBiy8tYlOxFyZsp2
yvjcFzFKfr6k3JDY2Gu3jaeIfemzexFqKhm+Qh1pYatniQfum86L1JC+EqGxCS/O
QfoIM1h90+Rx+VemHddMsAklnC+2cfRDTbIVgP3QGyzqVKM67V4MEVBEqXmFFbkD
4kbmOt0UIRShMSIIMWeayPv6W6WvJYTAlKwNj1jtDWgySuLgAnRlDwxZYKVYyOBZ
SgIAb2NvTkwiY7cynplhlawqMwQDn4ucJS1KJJfsliqF/Rnly5xtoTPRglAhakH3
KR4R5GtZ9q+4fSjhtU83HJ0ihAntmHQ7BTRTUps0DzU01dVYSnv/hEhJO4w82TQA
x4V3gcB8rAm3tvulATAPiF6VAwEY5EiVFNraEzq6QklE9WbklNrTD29zsie5cokf
VsLztfuJo5VEgiOnLqgAPOKN9y2csEXRUfNrTwSJ7kn38MY/a15kcg16K7KccBmo
kM3KS9Qp4Lo8u7xx9N7fxT5ixvZprmiDdNnMTkqPIdLZFqyJCLj3NWWbdiSY7q9d
EUEsZ2NI0vh7m+1EG90neCfF1ew0Y1UcvuSomrtzpon6iWacZcMw6LrT2gDMcqbo
nqaNgjN+qoU8n2N0PTlw0vC10GDxhcmRTgJX4H71IUcVq5tAxmBrcBxtgpd/OmWK
PAEZv8nQyzYkPeiuZRSetGPVBGglbudWZsophll8caWL1XAo9W4gLp4PfPdrsPrR
C/dGcPVi3hsxRasVx1kBlHaoDOCdvfNZ1a5wbk2pE0xZuKbolRRaEE48C7EwF8Js
9Ge0o8XOYkQY3C6Y1GW66jmS90Eny7vLKFqGokYI4y+ZBUNo+xESFyQUxW0j4Nir
PHhx4xJCyuI6ZgeE8Q3aPh2Glk7DojQLv6ZMVdJim6FldqsoHk+eXs12Q5IR0/38
CvcbRhvXyVvwF1DnPWQVNi/vsj4d/0pJQx5ydwKP2hWiylwZc/NCJz8G3ZrO5Ea8
fHZGz25uOqIyqkY87lMXEq/phER/WvM09yHgmz3GiobVMSTEVQHiLm+Cxe/EPsyR
vKb0WcPp38Jgd6Z5EkgRrbKZLtjj8gyWSlHNT1TzaBrmQUXaz9TbSZFi/MOC2s5B
rSKvToy8hbSVXU5T+dsI2FVIRe+YSYkC0lAmR+kL4sTc7FEy5IhGHsOguWLIPbM0
wMy3584MSMUjDvjD4glW+M1HhGDHETubStCYoxp4N1E1mRjJRryIFfxPVYhl8EIC
4dtvtQCp8kJUr2LIy8GmOg7I0YG7DA85qg22BaevsgUded4OsQStV63vW4gWSlj6
bnmzq8EZPY0ImIJIrbuQVcsqAVHFVV/2hPDVavfRXtoZEPMxth5RyO6mjOOlwk4k
DJyimXXCxwU30pQfeTjsF8o9bZtVLnLGursWf1WFvYc2TVvusbbX7qMR9byXEi4L
CTrLLcIhoag3rUrSYHxHH7YRsTw+z/YrN6YnqNrweg40JQsCfgWPWkFxDXLfrdxi
QM2DUEnZrCoubjSek/5sOMW8ZTXbb0kkrO1Bv8BV4XwzJOSSe818k9rmFJuXXS19
ak3FpaRMDL5b2d6IxASqUh3f2qidqNyBBfBz+wWGCSfD85jLvUfcE+0uqHXVzLyc
p5AM1Mm+J5sfNA/QCP7/dvumUjOloXpApGaS++n0UnHuZgS4rfTuc+Hskdy1wYXm
XSKui+h2lqINYWXjRW5bbVmaYaB+J0MQkp41SGlmAduuHTi04xs0gZvfuM0Hs4xh
OXHKKW12pCirhpiJ9nECGrMw4FpsweIG0pMVmJ8PI2bJKobuPMJ4c+gdPh7TtDkH
mSCu17cMZ7JtSJfeWdPHpcGGd2VatpwAgmWgDRDj2R3BVis2gggQzCiYaevwoxyg
WflA1wVzQxVISScGaF5evbQCjToAhJgpya1qInYWYVzZL8X7JNK8dvbaqOGrzYCF
ujTReqfWoihltGUDxB+HQOLB9l9/7f/WtNN9lZzqm7mfAozomSaXnn9Cuqm/GNwl
ovipI2HCeW99qz2BwB7UvhP5sn7eG4NOcDnSZMCoHMQOYmGmGuld3Ir2gIDKKbGo
GTQkFW27Wl7/t6XnpqHC9jP7rbuzx+wlFkwD6qBztAS8E4l1TULEa1uCdqREeR9R
j8o+fb6eKwXk097z+P/uUFPkrzVRxltmlumhgunLGiDi5A6HcRU2qBBZVMMSiGjq
K9W4zgC4XOnf5hfPAMk5fvXfARPsJ49+vDRXUovmcJuX5wfWrFY7ExOswxjEY4Ry
06n1SsfUhHnEZ2oOq8dqMcAwFcMWdYty9NJBUrNVfxwus7HiEwlXp/owq/XJGegz
yFCbidrm1SrAEJx2TMEoUY/7JI3RotqxuSfQwwRr+Cn+P3EG7llfw3VqaXE74lPL
UXbLv2o2YkUkhkC1P61jBxCTC1mWKHMo5SC07FHJn9Xan58lOuzaoI9kCOBxD+jW
a5a2n9GevE35eoM0uMWgxxk8+tGAL8NnSd78836VINLWr3OMLyuNgwG7PA/DhqPD
FNaGYH2OOgSwzVJ6f3eun5JCAakEQzy9sw6V74laSiwDVkK03ymjY2dgS7OQADoY
pcJKZGAxGS9REh7NOkhd36QcsTD/27kxyJ7RIDWDwhaCVn/FLvzf3fKBY1P4qYYh
2I8L+aslPidTBYaSL0uutpIfa74TPVa9zSMQPCdJo+J6H3DfEPsM+itZyWANJ75N
zn865S9NEcbzPinIHDshDhWY4+NanNWorXK1vx2giSf3WDmxxhrV0zjR0rLcqu/6
g5JqvlhqdaJB0nFwudvnTnU4qiGdbG1JSBtvz0Bmdz7loAytlV40IR9MMRfPUfur
XrTUEukiLYLNAmSw5ETv6RywjaZeBYAn0JUYkFAmwh+vBFxR9iUvVyvXj46RtjuI
VkgiuED1wGQn5LSSNQXQjDDo6AiOBuIGx63LV8ePdc2nwCl+BvWrjMQl3MuOp1bY
J6MZYqGePo7saoTT25KqRZk8VY8csIHHp3dR3pqlbPAbJ4MTHVeEPr6+Qp0dHyja
V0DYg8127zRl/HsZDza5jr9r/jarc/tLKmqw0P1KD+J80XpX9UkbF7uys0y0eHuN
UP/bTSOSZ80ljKuJ+VliY25Ah0yqa1Rl2Tz1NiFarv/3N1kYM0Cvlz0GmV/8Y2iA
UJktMKjFOQKvydhRnjsYO4ZYhpdO4zs6hRysQ+cjA3+cZTOBPOduaWCZQsCOVVui
h8AeJbWcf4LdP6C9+GcGYHxKpK7c6F3r4QK9tiSwJNhNzj+KGY6D1qP2YDWMMzXB
NLz+5iuLJjNoQjR6iOLhfjs6gMpkv/hMP1797bKd6pE4QYNhm0Z1CCLTvJFIZf7t
zoMoiLUPMt63Y4pcE/HsUzjQ9ahrfQtkHK3GaY/2hch6lupAIQNmb9bkF3TJKAIa
b3WTW0H/5hnR6Ry8chMvIt2fdTl3NNFZDTrS9fi1ml2dcQOtGzg2ELPbwpRKYqUs
cu3fYRQAThpT7NymZaQygxoQAw0nC9Jk24k1wFGzQcfGQ6Q9KCmW2mysIkHwYr9j
1bJGFCerGJA42xhNkL/RzeeEkeF+B+Hrp8dujMqRnJRG+jaxEKWSvHBKlj5/pDvx
l212aG3bNd0WSWXERs5VMbgx6Ut76gvaxUZHfGugt5OPkSbwYQQ+uPNLFjSQzJvG
9rijwz73DnrutQtb4n/jLOYFNdGebmn2XQLujIYJyG7e/QsrgiPze1iUNE/XQ1ir
zC0pedOfFVJGqUM/7T5dyqZkqnRWFcm4+wkfrERrsb87BEHKbDy/VwM1JGX0E7za
UeLcNhcnnFN+qYOhs8vaQxZsHjNWj3o214hOfnwJVPxbXhl7ERjHcSO2b6LtIrX7
k+ZVtgxJQgHHGy/aQeKmM6EGrGcNDuKCWt2cW4O+3oqf5ZyVu+L1rJgTFBgakHPD
emuri7zEVWGJSun65SZZ/ZY9jiKXIKlmYEXad32GaXCos7AgLK2ni/YBMHDES9Dw
2b1Q4R/xSfslg6LBHEqht+X3hfC5vFNKbSTD/QAyRgtS95dm5vt9PlwOlHKAppkW
k17LyvcxP+3vrd6l3P6Vccj7lSYpI5UFZHj/bOsFP4S8zbfKC2kqLXFRrAWvMpXD
GOObnweZdR7fC/ZB47+BXyG/Kjb3O5iAAiP+1p2gZmXUgxFZMBCANxmbx9uTm/9j
o+zhRPDznw1tP6tDPoGznfhWCDmpH0RYwLGuYBkfDMX9s3qkoCbHL0II+AGy7kIV
TRWwbXZ0voOoZigQl3IBlLE3tRpx2AccvazakK4PAiga1Kj9EH58a2XayZa9o6wn
CdUHfF2OTv1WAQIW1b5ffW5krkFQeW92dPGX/tu2rmIh2piUSfrxlAXhcRwpECAX
RbKlWdTme9Z+FeVeIv/jcQZ6/WYG5YeMjmWZcPCnnxcbwGoKw4Y2sYB6wSmwmT9O
2eELBUXtT1NsiYI9kPzNdiC+Bv9pydpKqvLLi5iGRcYiHQTrkrNWs+7Pxa8RFYoW
0yd6KM504BOqJHdepwkcHrVz0+T/Vuvwa5uVRd3eUJ4I/M+UL8Q1xBql9632ibZD
L1TPRaNpP6dMafLCnqS9Q2ZilA0yeScBV0hZuU8WITsowFRma3oAyQxj/jRd+Pgp
ERZNVqlLt4xmU0bL+md3/KF6/ugyJ9fSt6kZY91PJcUF2Ff8mVdIMvH16rwUAdi/
zWq9fwiEIozHdvVqLunQC18xB9T1XzoMvKvPT+xjJviDBOKmg25GoTI3vPa0mChp
VAH/5B293uYYsa1CkXPFpw7kgCKoie7hi7Uhex4RT8yuj1LwN1gaC9n6zfa80rbO
He1ygaAyK3ReSeTs/UO7KOf69bMDXgkxRK2E9Ljvkaghm6APj28nowWMsS/m/rtL
KMCYId3+l3hgdJi/D+uq9aIclBZ8Q91WmAI3HscK299F5GiZxCDUJdMmJPI5KPOe
dpR9ImjczBAseZz1XnN3k24PMU9tSeqI4XYC3J1RH6u0hGzlEhbTq1y5N49/lUOq
LFkjOfD1hDSiqhgQClTPOVM1Xzyce0bsnJn55VXQz9LCLrW/BuC++BTOhXGyXKaT
xpvPE11r13LrcGS8onNGy1se7ucQRY2b1SaG2ktJj9isvXGucOS+OvJrAtE29inp
OgcDhid517NNZW9SIGO1H8DHA8xnJ16Viy1OYqwFWEpTrKgDQ3soWqS8mBamoxuA
ZQj8aV3eEmMmLFAGBYiFGyj1sm+2IUXuE8bM9h8hn4BR+LFzK4dc/2pGL70Suoom
+PjVvBuwecnjO0Oj9thGl5um0iR5gyj6SOqJwc7Zge10KiO3D7TCylwgE59ambbM
4ar2Qvz6y/kaLbVo14CRbCgenY9qS88U20cn5cXLHnaKPE3CJgbxxtraz7qlK7gG
1/s2cNZD3k3g2uVuIHlF60ynHJS33qMxMzmKTs0WA/ALJshOLCOqGL2aWk13TySv
bGIraqcu3Y//yMMHXD+n7y1dUKuRRYIacy32h3mkQoQsqFrzqbHJ830bW+MmqU7t
zb3MV7DQGgRKIqWE0JonFMfp0wFpKkNKyjAJYJ8IINDhGRan6RACgDxfOV7+ERfS
Vsa5NgjmG10+kUlkNkH3IVLBjarJM0Xn+FRyNiVFyYEfD10Bw3PdGt0cq+cteO1f
loq9rahUvBw/1jgrJ4C9TGQUiOF4g2WCYiZKkcg9nW8ZieLkBjlvsYwSz8v/PoIc
Xkv2WKUHWtyEzm9zfePvTKVzRwDFCC9FPASTe1UDYuMpROvC9l/SsZp//e1kzAgZ
vc8zU1R/bN4N5RkM3w3b8gh//zf4lqEtyi8KSiFD0O4jOM8gWL6xhFz3mxQyCXjx
lMQfKrtZrD13bYYyJbbk8134OR918P9lfo4m48imKNvLdNetjBPEBuBbRmzDQx/f
B5Xw4pEkie6M3J+bo2eDMwaZujn1EGwFZfb4EIlzFNKh/rdJrUnkioNtD7uSFZoe
0AFBdKHHwM6igut+AZyb3YvvkVZQKLyAgjjdEykruLA09mVBaW6OJ8Hve2mAZasQ
NcZ+gWwN28CTn8qCGZ+7BFQuli85yy+puJXwe382yqFstFYbixfpD4eT0xWoEjoM
hn4abN0/3Anaa4TzNd7dWb4ZabFYTTMtTCd65Y0/DEsxUck2uvO4db3x+z2zs4RB
OeoQ1mRKs1oINOCZdwJDqUt3UBQ1GYUZ7jnYxekfP+Vvw76Icy4ihT52h26LMAuV
YU+HqER0PAU5CcWl+w6cL6afgfJHmin+VGw/D7tgERODwms0NufRC/foF3ebUmFd
acl1tMqhD6vq6GTSfOaFCF67hka2sV50s3z8i9OMkYm5IE7+MZIOHR8qA5QfRfbl
aVswEXEdTR+HdWZ1QSMF5TgR2+UtQ2EEjOb6fXHjPqiBk1T+uSPoHj8VwCVWvV5j
9HyVDJDb+9pYA8EuaGywgB1M8EbaHHnIGd+YIVXpw1mA7xILgq+cW9kmy3IIqiMB
yq0jW1T8YvQlWHoG7xuiOl9cjhmsvK/iUh0IrH8xI5/AVuzuwlu/4WnY+IzK8Dxa
sP/TdgRdVGI9qoytvdSGJuMECSORQ7bIjDtlh0zL5rwui40385Cs0O8c4dUQTkwm
MB0+asScbbkEdq2M4C9me/9UlBK9WfgohyI8C//CtC8p4oGIMayMuRSCsG+7jfld
EwdMGt4wwpsFdbIHxXWkLMWrU413eLV8o1D5TyF93c/WLz8/A+bR3Gasuq8nTiUb
pWmtJJu289prKUDbXYxKMtVrAhqXR7nnmaafIPAnZvYNn6Sd5gqocpNqDS6P/rpx
33vvYYiogIHtJjT/4CL+pvCbwF6J107fn96/3i30YFYmtQD2IRyEUT8gOAzU/maE
eJ24HmR9dEdlI+yDrHyZNBnFTH9YN6Ev07v5Ofrgxsfkj+c/N3GSxiW4CW7ArHLQ
BDCMiG6KtAwfAcsOQyA4n59syMRJ1E4KF2o4RN5D3X+yEqME/juBk6Hs5txKsuuk
hMOZ8i9iTMezShQujRQvpEXahcwKv3bHiLUFHt920md4u3bZOJqY2lBspVG2bs87
huchw+0PbH/u8118lc1vK8F+3jW0keoNSWLlhYRLC7cOy4WjkWS7sfoPuaFuAriV
W0F9ElvCGraNPDQTydEBQdjDWdUYJGzclQSsQMFvkL5MWNpIzHByqluQQT5FOwMu
qemyAoRPfrhSqdlA2N8Au/TCOIdOQhJ03awWlcwo6F0R9t6KSwRl5jBqyz9msXkk
9ULpOxpInoFRUZ1qgJ4ji9oyYI4Uy6xzQDZhwnIYCfw48/lMy2mWAFkxGsLkv6cF
0VA0IAPvSCH6hHYOrp61zPi7JXuIx7bZ4EXpY9khpGU8EItj7k1DewYIoIjuVye5
yAdz8xbrRdo9zFGJ40T7p4qjTr7MVbjzPKeL7P7y9C2Mxa4H1PI2WnpLor2DEA/o
QrfJ2kZnScwMhWqUFQop3FO8jxIUCc9dYrLyJV17iy3/LO3kr4aO23dftXzRnV4M
coo2pHzLTN1HouWpvlIKZCBiDuE/O9ruuMqzYlt7x0VFm0zUVPsd82vqjOLWDeAF
iPy/zYgrsNKCF4Siy3W4EK64idUUKQy0dy6TzWVPbEI/yflZZcOpey1c6TMlSbci
GqARcHyjApafJ68aqsIJHeLY1gi3z1E8w8s1K0tc3oSCMAFXtwWwWYxM9b8WHa++
kYtAX5MWy3gYMyUe6GVllGFejFMsIodIUi8wNp6L6qY+rn9MYuJVkQPSvgoqvt4O
VerLP3e/KAsNtYOopD3ntOSHLiVff/vLGC4bNCl8YyaFG/oC6tzsS4eB3n+L1jUm
xPmXpBxJVPXmbfJm9Amz0rw+6+tW6/qROb43XoiA29wQdLIw6yuBaOxCkmTUhAa3
XtZYxlYCzU4jgh/UckqrKlkB4XW5ncjPubA9dSG1+Gf0NUSB6/+nfxbATEpp8fqR
3ImY7iGKsefNVCrvdPBij1GZlamjQj44s0VmQdy0UF88t2MbiaZAhevsI6u34Rb5
MPz62EDxEXQJPx/QHvivqF/KK2wrxOP6axV7timy+hEBqaf3G2suGw5xvCxt5aCv
xQ/dFKJVxGZxOf4JNvii1kyXDkQ/UKIhAkzcPik0a2bNNDxBPJcxn9YirPAOdPcw
R4Sr8EIhN5wQE4UEg2VZOx7duMH9eCq0RZi9x5upI51B4IV+jPYecYdVRW0URXWo
1w/6hxFmLtvUlrW3yPItyiHRwMKA6p1zayaJEsa17wVh1Fnd2ipd/gcfKN2WJr0+
zfD2P66vXTC05j3Dhvy0WIq0piYc3h3f6lKSlqVXc0caLk5X2a4+zLRlVQ8VcUEG
ELkLcifN3sM0TWg1Rfmecw4mymr3l429lwCrTDRqSl4Evz285rxp2/7UdXmuTauV
EoDMGbFUMcs0XmQ/HskywnfL1LOED2+vcOyovPP9qhranQZoSvvps3DXj5e6tyv3
4OsetnRX27OHvWC183xIoE6kJmvdUkdvFPJlpJdLr+TENqd6gBxPAuh6wzLR9OVl
5gORLneiChXZZeIbrDAMQPE1Wt3If8iUrAi+faIHhyKco/o2Tp0nOmu2i586R7fq
EuBLPWbsz83K33r19d0of02+cAa3hYjvXpz00ZWXdGRfcfGqpA2sH2JIxNCKJuLR
ECduRvza4kxRb9xj7rYCNmL4ALo+NqUxpisIjUoCUurEl0QwDPRgcxLd9mJ/EHbf
ohPvHK9RAHD2NySwioD/W4mRpvdxcT/nyfTdoOwvIyO8nyOIqx5DcbMuHhVhXpmm
Zc+VzJ6UulH2fBiI8ALsfvS2Hkht5tDQuZWqeEcsF6tbPUffkO8URcSw0ihooCOf
/bm/PzQ+wSt44rNLaQCLYjE4ekbho0z6fdRMUUCM9BfIuPr8gzTw8wwfUuOs1B/j
OGotXhOGjfrIRD871OTAhfLpFcNfdXCHxpSp7o3xG5FfJcBe3xhoiH2t24HnEDIv
gDvdvs2YksyCe6R5O+7LQtatixR8+QTMS7YBP28z/Ug+apKadAuLlkiyogPDdQQQ
+PfDmnau2Y1O84j2zYj9eh0O+BFxMZH0VM7wOIpGa9Y/XCkxDYm6IMND9eza83Mh
YZbSIREGyGtxWcpq5gRGHoAtGgxuXq9jxT5ZU8zr3fpk0Ny2RWLosWpw6IGcyL2w
UFiURmJ4I88uu4FonHT0qPa75p9wxP7bRO3/Ot6qKn87DPgzYxGkxb5vU+vG/lSV
d5ZoJhxQ0XRMEn5IcNOcQcOY/L5cwhXFCEWHEr5D1zVdNBnYY0Y1HRYUU2/VfVvM
eoHhWd61NYYpI+F47lne6Y5eZFxdlXSYq4mK7m9bV1yvRariXGn1QDH79ZpWGYgd
Ielij4J9oZlMteG86Q6RCkdkO7ERgB2XSAae67liKOVz/Iow95fnY8Z5Y9KYUQ9a
ncYnHTja8tVuIu12GiucKpQykZf9SttgzdpOY1GJi/KBqAz8dP/fEysRwrR1idnD
EiMcfDHWuIgjWwtz+tub8+uKC2t6MP0rmQRIcjXrsItKIf43yKQCJaQy7Hx+DWKv
c6/AgDwQAMs4GEkbwiDT2QBHjKX/cl4peuR41LxzZpE44iNHrdQ77bvRj63eBuLT
m/vC+MrSHRTlzRtI69Fieo4NjvtFUsDHyXM0oI+Kpl31tCIag7kcwVCd3AWn0Haw
GLjma21RfyGdKlnbZdKKGF4dWx2lQuiEA/xsVxGhpZJUSCodJLtxg1tMNtik0L96
0E0ILv0tXQy5xiwir4qfh4pXTDn5qQkOFKgWfmM0jknOqBg04FK4nLxu+OpDnFNi
PxC5r+hbPapgxVTLotl6CW8TJf8gBRhqSM7CXIfAJ+2jf8zDFBLWm6JtFY8wuDeB
XzMCo8CNvm/KdWnJZj6bmeP3uo3gIQUxx4B0YtcBkScetiHxFxDFzo+ufaTamna/
VpWybrxEJ4AockhYSJpX0kwdltF5+K0HPd8HBbLGXZidElZSM1yj378Ddr81Nwu1
BkwVYxWF3qJl+/mWJ/zIv0fXL7ajFmOsDg5CrfSq8nUExH4Ee/un0XmCqTJLfQ+j
X21W1xhVZBDGb11XeThiuI6UHbmD7DnoCsXjhiJqcPtpHdQv4XQy6WflgyY2BRb0
9vTzy7fHytrUzYBgrcHdFTRmqhjAkKgfwrLMdvgQnJTWVAKpGsWh+W0NPtD0q9MB
Ee5uc7f3Airu5KcnpmXC7ozjF9zjsKEAyzJUJ3jF89F8qpztaYYEfcJ4RQFhebos
gC8AErlrbEc17/c1+NI1SnP4jcOqz/A+f5bqNjHcwsoGZ80IP3EuGjgDx9h8l/h8
J609nsbWaYYYDFbL1CFpPaSQnJw58qUGM772/oHcL2Fg+iRdTcTXobB1xvkDz7EF
gUYb2aFQYE5YOWDJDXbyokoU3ON+UnXkFlgsOEieeYjilBF/GEKiypTgOkS6WxWJ
ZmXV7Hh0TNoFb5+cwBeE8PImhKPZJZsDWTjOxF35ZR/QW9e+mN72088iMw983m5R
3Z/x4ww7ep98XYZjanqkvrquwmwwSmd1AluGzc8ho5XiJA1WpI4mQwW6ByD6Sj8W
l9GTnWST06wBgUHSDrOMz++ba0rjSEj+169QkkdKjdnnpgwCmuNhs4awi9JSAlWI
rq7gjXi7d249m5z1DYd8Vk5hFlBMyza2Zios9EIfA2dtW0+17yNxpF6aMTPKK2Z5
Jcz5Y2zaZsF/ujN8GllzvH8DZIxkDyotYmx0EegWkui2khyh66z2zqSErCWdodg6
nR5X63AGrd1lfz3oPySZc6TBiM/qFeHNXCqaPT78UPOSlIO2D+B8r8c2q6W15cV8
q/XO2tVUIUWt7jVgid4Ikxxgn6db1KLOaO426boWruJsjc9jvAPM3DmV9UbqfCDm
YT2X7xhHFqIbafJWFXdTWVibz9HpKcxsYr9GX3+fL3P8G6kgoFG1vGuR1SBvtu3H
pKWlswsiztDSYvkufxbbXb5jIPxkt+YuwEAK/IpJnWmlPPi+JV0FGXTsdZ4o5zZn
D7ke9zCMtD0u8EtfB2lgUZLNUCmPuU2wqoHDCORI3yBlSlGPlmuFTpZV8zsAmR69
7J3AfmhvmNRk3nMZBsHLLKHVhwo84jMVeZUALPNph1+96ZEecUn0pm4H+aOXDs7K
RNJ9RmrSeL7CuwDWyCmUR5i2V7u4xIk0OiGA1VFDgTyMezX+J0s05m+Yfd2EYy8D
mI47wezc3aFsqxqntm7/ZZddcJ3kDCiqtuzXdNRxWN0sCi/vOJ7aiNYlm9EoyKBK
3AHcmMKuIwaMVNuy6oCPtHnDPLU+aViu0PB1WgcAH0J/ElekS6iiA0iG0Nr/h0mO
yQb7BTc2nAcvcfu7YJPsf1Up6duJs99kkR6e4MAMMN41ZmtlVDXGcly7N16zRxZu
ieGjVi5zcnlVltVoXvpVx6iozprFCtdNhBiBG6IKNSRfdFyTtsH/2TX85lZpO+Dv
gojvnAW7aFgISRi1DPUDZ3ZgwRluv/taI3c+Hcu43SQ8+0DuWtz4hxDcGjDXeJS/
Tc9zcTCkDu7RAyu057LeCQ3anidk1wVqageQcM6Mxy2U6rOF4KK3yxBHsw0SDoFU
3j+yTTsqMQe0DcG1ge5O2yF8yLWBouHY+w8zNRXqHSc1l7HxMt9+TIe8EeX+jhGb
imIChDTUqcEYRasNZxRzXrYjaQBKfCIw6TfeANpjiAmZmjlFjKZtZPoxDF6FzUd0
pdl62tuFS5SMMJrhGI3M8B8YKfM1MUFKw7Gw3N3jp2O0vVbCIiR0dEwfCEGMKvjJ
hSqGzEnuohJk1Sn46gbxNzjjnM3McSaB7mV6/Geh08FGLUtNdkK9TkGnMEqk8AkY
5Dbq26XbKbxQ0oFq2F+dkGFYdNZUCJi1MZ7mYEI4Isx2UT+9ADclqgjM0Omn7gPu
RoYwIowyBr42ovslxzScG+2Y1/bC2KmBIlJb23RIOdnasmi6sv0m6E4SL+0oXuqw
PrT2fsTli6fLmBc65sT8IGSwP+1G4uT6lW/G4brlsRyIEFpXuGiSyqCtGUuDbCom
YIOyILUeB3oKimfqtlySBiaNQcisZURALpj+D3LPr9uhHeinCmFzzQON5og/HzJX
IlbJiO9wnik9oHKd5+zegNvmuIaZiYRqYT2jMefu5Qej8HnbCh0Dom1X4mWnFWvX
CQepV6dwm4TAExy202tSd65HihMdviQodE9oL9imvc93V/LtjwHzAyeKnLOi36iR
e5XRhZ+5hUpUBWUFJQzJelNo6GRLHo6+IAM5nl2vIT53vuvwUmNnIS40SkzaRsfu
jvZoo7JU618bqhBYDtSvsZqTIyeGbyCr3SuaM3rRtNYAc7vE0HqQcoB2vEg5moV2
Iz0xy2Eddl3w7T+hsfNi4e2jc4nhOG3nqKeVLZou/rJwJCizGfmNCEb3YVdc+/59
wx8zsyvSn2mX0hxObcbGSRvyjlcRnLmHPkwDa0ptiMta1t93NRAInqmibxx2ka12
gY+Gqvcbjlbxq4THGe4CHYK6wWCrtIcP6c0g3BgkIHcKU6TXLqKFalCTM7tpKAIk
8kH62YsO5cZ+suEk87mZ9Kfg3ZcaGygRtEnfwvTJ71B8Axk6VJ3U5pUJYYsliyA/
NM1Bft/Z4YoYHMjL8qGviWBpILYP6yvPkv+ZwODo5TLl07hEY7Ac/0j8cyu68enH
NvW0/UaGd9hNZwMMxQ9Vdbul4F3cXM6sUSdFSC5N5qhqLSyf/XZdcxyhcNXTmmwD
EQpmgg20yJdD3QQPBINHh+lGo3yJctSBCKEakPLXP87gmkhIukSWP+i+F2aAmR+L
dpMYAcsdqB7Ie5x/i41ikmWeGlAzXHMmdTYvNWA1NHCjpKRlv9iI7lde6+sjLNz9
qapINd4COwOtEhDRgaTo4THSrHmEqbsQDYy/BHYgMNXUwsWmOE/kY6V85mN99t9t
d0pug22k/G+ACMAe5HO3xNYk6Y8mivdYmcVBvsNjQtWnNekLkdZLV8nvfwjZo+hj
DBIWvEeQPD8EjFQ0IngFb+9i5i2mW6NANNwO5wIZOOy6nQPWPmMzgv8BVVsH8Z7q
2Fp0Gt3tb3LvkdNGTPNvQ/HSIQf3hKLmOeGRUoLf5FbfKYN2V7HBsOJ9y5r/01vu
fN2VVH/QHYidKlV6IKaqBL/AQjW0f2mPNwzOBtyyUrOeAOGTmBRBriNCC58vICRh
GtvZVLT7283WDsom00PvoLURytn97jdo8KA8nuWkMV/DiRC3q+yGoPdpCSN7tCW8
RLmjb2T5pWZ23iMciaFubjf3fDDWWN//5i6fjqBRkE8WNzNRPBVfacmzSUK5hOiL
v1w7+nhyLx9v0CLIF1YGwjEspcr+a5JJjyIIrdUtaVB5Wp6UYYkTru8lvs51S6xm
9E/Y57md6B/xJwMswF3fpnWOxN+IIItyvq1ePVAfT0aByTNHoEaCnT4PpmFChrHX
KK6KX+zlNEC1XlB+iRtY+iVW9pc1BzTwtzhOC9A9FnOcehDyj0PTDr39aImjEOIQ
ebVIaOAEEHQk919RTZwNTuMwaoOd2mBnahAenJ7bgD95nm698bhKHuQVSPnEO84f
oBKhlgOs4KCzUXQHliggrB1Hc2SkCBMglWbe8E7pthGYU+MBsyokM4Ttbt/hMb2/
ckwMdnZ4NRpYu5RbOBQ8CYUOGluN2lmWVqJu2JmO5W8PaDsRHNRCrFA6EHJ3S9pH
hYd5/OPXOBzx52HEGEg7tyzQF7c4M8wEhI7XxzQYLF359cAgSUaJgM5YR86OVPJ4
s7Mb8nZ54RhahULEyYyL322+jpU9q5R6QvCqMnB02i36rsymGZnGa0bANNl/YoN4
G0NLA77eQhtXNcANaU5Xaa8114MXli6NlqgbLmnBML75zfJHV0Drg+TDWFkBrpO5
HkXW9Qj7PoUxgAzkg1JduYS5Id3MzWRrWr06tpUoyL8VywR+SvPjKSpO8yRF2yFG
GSHBoGXLB0QxBWmpazNHU/OGeqTcldU3J6ui67uJT6SdXnFDP6nrx8lGgHMP7N8G
cijmyrrH0wPkB4aiqYe4H2rcGYwPLx8Y9aWCZ8QG570aunMdsvXKG/29eQ9tCqFL
Dvf31hmjfpx1XltwikVZTturb1xYkUq2v1nPg3w86tBBHqX0c+WHzekmqY9cjYum
W3DNQP65OJLTCcJh0cQmEpoz6Bs1MuRQtt/d2j+/5g5l1J7j4FJN4xk04HlE3ejX
TZ4tOdioauZiMR/x6njhKY6Mobxwr8H22P6olgq2oU7jnNUEmsOaoUcJ83G6K43a
HXSuc/BJ75bZ8cWEsarV1qsw5wKtWazFaqlzf5u5KSzCmxXg60KZADvdeStKkY7c
0FD7T06e107xkjGKV/Jmq+tZ9OiCX7p2djJSPe6tHSbcS3N6t/PBNj5uHxRcOBAN
B0tJf7WorawN4WrfNVRSl4wZiUYBxI+ciunRQyHBYD9WsyG6TLSFVKV4bdosfK2C
X0LOMCX/y6Pu1Tus/nAnh3WybABYHPf7ngXH7QRdjLsTh1iGHPk10MS9iGTKZamP
3NRpiVrrzYvY7IMx0M2J2G3NxdkDsiJv5N09eHHcSZSsjpUOWWaf2/0/MmXy3TTd
FSM3HzWx5QsKMFLL/PpCvvNdIKfFk+qMB+JG8EgxsqtlCVyunPhaXOBuQ+fKsqUa
J8c5m7WmZUBaQP3pcw/6ozLkBbACNMylNAEJR3dr4mz3PpJJoVTudbWm43eBkW/q
Jj9rXk56mazQ2y9bmU9nyjuQlL9Hyc60ShrblrdCZYRVAUzbw4e8JUe3mOwNRYNp
KQbJg4ylY0LC9TDVILkvkfkLNuOAyrYjkppgLTDci3y35mOKZ/IK1Wc7w9CHRFHY
+8sRVs4w/pNi33EXwg68poOpo1Zl5tviz2pOkqfXQzP8rBV8lHBFEaVh3JVT85jM
ktmiprgzjy92vTZB721YJ26tURCshCbKWWr6C1L4wkxK2/qptSI+UCtcXIdxMrTi
1Q88wSDh0T2JzKWr2YN7cBRf9qmDqaWrj3KefkH5LAV4MXfcSe7raxX9T+979q3O
4+xqsg5QdPKj8RGtDD5NQ/jw2w/A3JyH7rcLeCJpKcUqyyTXLEji1XgKZ8tjGoT+
W6Y0eH+qp876mEjlxwmBh0dXSqhQrmrtRVs69h/E3spaM78vPIvhb925wtI/WhWU
yv2lEOgv4BK5qnl2aL4zyMT7QciDMcPxswY7mMJHBVt3TZSXJpph23HsGaEhhHem
a6iwlrzCKiNYywvv6jzYmqQluMCa/q0tkc1iFgixUyq5aVZS8KwdPHixCQed5Ssn
0mtg8WG6SxzatK1ZWRReyDoowOSaOlnTEqtPoPcJL6kz9GGYI6c4RAPiddhXI4gP
v4QlwWKudCKn4sGTzBEN9LTNxnRnNlrf1ZuIj9Ht1Ye3lOtM+70XJkPUJ40rDYzD
16Z+kDpQ8RpOnA55BrUtdIIpceLjAGKWRmJBw3hdZ59Lar2uY5DxqN3SQy3+xlK6
q1aLPQ83gyrc6O+5j28FyuERyxrCYah+EDYpojs+741+75/+AAt11Aes5+Aufp+h
ecyLgg64J9extCxbWm4261vIbF9w0hkvCkmkfUYmaRvMWCvU3WVSIgdmKZL5Xajb
JF6IB8XRP/pRkuQq2VLoNRcjcbFB2PtORNnghPp+IoKuBbcC2HJOW1egRxTDnV+c
VV5n3b8VnkljFGU5ZUU3Nz09VYKQfDOcBHQ8A5hXg+enXuBqWn4EYH1swiYe6Sv/
Gy6lWGvwW+QqOiugxqeWwDp2bRAxaEDft1cCMW7h++hR37G9rF0Tjt48xTzMCBe/
IgMJSDsnxKXu6gO5pfz4xRIpxRoZ8Qsw6v+cxCTzcp5KVmtuVtjQecdvh3D6FhJy
zlQQjWujG4q0LKczc3oU/igGX5zHQGUNu41UQub4cJD3vtvN5kRd4gh0F81kTohI
hH+yJpN0YV7Q2+RyPrszMgrEsTfPzbkKog5Ow7lhvaCoQS6z8n+GHB/EJ7SsJrhe
sqcKDlq65mJtO1w0hWBlKIy8zK0U3bMKt0MqhtvYmQfw270w1pn/qXGQdIXewzDh
qDP+NrFpURgSZA7EmwaO/Ifb5+7eUrQxHAHlS5VogiAP4mEMMlSlhIaavccMnaZe
319zHDnoqrzSylQYAAE405jBhmz41oNh2IFBA/ZdlMwZyHCGcn9h+pyK/2ZXkmmQ
eHKwjMMKr1FJnkWnA5uQSBrMzebJroszhj1QxRdvYfWaBMFyY2qGotz87q8C/qQ2
BSxmjm3LqySVJZFKa+Gasez46d5tGLelmhtuUXB9+Ee3QFMgK0dyXpkgoAob0xh/
cfiSzzs34U+8aaUpWJHmurgrjivTHjpjzjYismZRUpDx2wgUd/gVDJdxAiSHeaTr
9H0eGpdPs12U45O11l8v+oz45GRD4qX0oIQ7tokcHHb1q1tw18YC8haIaP4pdZI2
d6XyECx5WGh4UyJe+9SaIau6oWUV1bn8nZTm7nqbY+0mfUUauMJ3aMiytqLX7+0l
h0yPEguwsmfWDPa+c4o3JwxyMmWBbDOTXuj4OXlaNpGh/7Gx8/cUBSU7eUrrBZlc
Nph7/ImpVuVlf3VXdn+/RWzAXdF7JOmHucVgXJdTaxvbXEFxa/L+qDwSZdnsp8D8
G+nkgLtZpw5lDc54Fh4XeW8wExpxatwA20V5/BbE/CEPg/Y4sMgQibdCEj+To52C
spxyyqKCBlfevaxsVJYYRXIe+5xGO5JH7cdw8T7Ytzw8CG8/rXRlyAu3pH2GJy+o
SSPC7pXiydprtYkml0Hz0M5lKLGctkWpArc0ilVj0VxUqzYeB4/GOXTSuZaPqVry
9ewXWGjLW/iYjHLJjUi1ghXz/0+1T25mGObHHkEslfipmdQcA4CyBOhKIiGsm6ed
L32qt6o3jFrbURTFSHdLBkjbWmp8BF60RQl4xyzwwKLmlA7kjBU+2JDaJWTKzKVi
xZzRBXc+hgwC350dL9hEFVCWqfgzfNT2RWqfsRxaTGIRDL9iojS32bDx69fozuyy
53d4rTw9XpEMIpSXZHboK5LZOEekfZoi11RMD5mHcdtYnLWlAD2fQxX9UqT4+IDt
Vud5FEArWSqmQy4u/GZJsWB6tQ1JqaUDX4ZYYv9Pvuwf6YbDutc+tqKKhygt2jDb
NiMVX3x0wpYBkKjaJglc+FTQx1pPLKcWTM4LVM3IxPYqT1/Sr+2duvRPzeICmALa
4nFPeW4HD8dcaXPB9GEB5qHZrM8114i3sV5/O4lTw0FlrQGDOVj905IpsYaZBcCm
8dvNHNq5HyKKRxm8hiuqQQRhZ7DSu0O7342PetmgHUynZ8f9t/4Z9TWDUqc9AszA
Ujqwq7g389L30OOs/fwNQAP/r57Gh4mcYuslAcQEWAm5LTxb19lgVbT0Z8SKllLn
DT5/A1S7cOqyiDq/7dctfomQ/zT5Cuf++P29KTrUQ1Vu+bXUjXj/5I6hmUcL0Nt1
unQQSaGrLhS0dljte9+RONlLiF6Mowo+bbKwDVPzTJD6OCWb0wHcvxVJMy/FqXWv
0yzdjJ8VChRgcFODFyQ2YXytC/O6/a46T4kU+xNm/ubHpmPGkZo++7lC+36Iq+Q4
QcgZXha1myf4jzwgEQlBj4g86axs6Xh5qP365SOgFIFPr1yfqCh++drK+d/gUox7
YRB5K1yZvGOlJptzYLtgU17Mpac86bdIYCuiBht7Oawe8NhEJHRHylAkD91A/9aG
xnFdoAcYX9BcuGnuqAaQXgJUB6AqRawqDCvFAMAXbPHUn6rJrXT/RLMHb7qS4iN7
rKa1PPZF8LEE7f86Byb7TDGlahwrjBtWDYHv0axQXw+jVC4t+pCUhrpPXPXgkv8k
DzoFvTPqLIYkyUShGsZBYCjm1u5SCMP76LgWO65TpYEBQK9NrvxMJUdYk2j6KuFg
q4Q5ESt6hjQo0d1FobNOu/lXtVyyrEc1T7Q3bawnmCl4GtP89oSFoAy01wGn95h6
8/+wpvOPSxfdERCsTtLfmur7JTz7DQuFedeEUGaHbB8onog2nzJT/mHBpw/27Otx
XbDmljY2nfSjYBeoOZGU2jQNBDHdMD5iDPTNGgpAHn6KpZ64gwg4I/Onzmq+XCvC
ajinmTAloCEfxkAjlBEfLm5iuMGgdasBTgSbeCzXQRT2/Se3qhzVLsM99IgEdyVN
yUY9PfOhQt7DIUy4mF05SDKniZWmdRHSKvhcH1OctSOmhg0nyL2Qpmz4IQoip3Bg
8sVzgizx5rVn7xuxp/0mmk5s5X7xsPznX34n72y5RfSpa1OsLsSB0HdZq9KeGKdC
fgLGi9GR9MU3NDNl0lfn2mpAA7QkXh1JZeqM6IYkvtui3jT2AzqarIKFs7SDJdnC
4Wq27Cipv0yJ0cJ1iP9S0e3M26LChm6Y2gk1seQA/5G5bvLEjIDo5UlGGeEX8PI9
N1758ZgPdxih79ZbSVDm5+OPgkqveoV2FlGK1Ymqsm3WLRw9VA0vWFra46ZzSciv
ez3Vw/AMSplO2IgFIGIwV5+HoB6gQn96ysZWZjeWazS/J9Ei3h95Eh1Wjw22dfNF
/AmE4dUcXe+SfwTSIm4UC2tmmv1SsNesW7PbwvQ5OycazBYZo46e9YvlvIgjpceb
rxhrKif9ARxIziUbiqdn5Vxgumntw83sD3LTJEjxb8zXIlv0hifhsCxEpX/VJoVP
hJm5VmKJn7bhYJOTa4KFc3Q1IzggDCC0asTM3kOKoq3/2okDRfYW7Ewc3LBMefGm
kU+VSa5zw9geXvm86lIICGDlWB3hDVGND9GUZN28MBg3R2tZmpZwFf7TrjjO4Up9
PoDfI+KXOQ+gqYeyJecn0rA/UOcVv7OSro6o3uyiAJae47ChU7zk5MBvvOcfFIEB
C+/NKIriptEP4+SQWpNIPeQ6TBM1A9r9Oi2WJVYYTObA7jlcc/0T+jKwIBe0WpDc
qwtAQK4OmLIJJas5uuhkN02pS6zIzWHop7k+FVLNq7gfBU0YIWH8tF1sGoSwOL7U
hqYFHzshDH3TI84Repw1CqMMIiZ1s7nlH9wLtDplTaDUigQGFOGa8fVXkEnZYadI
jWfBxh6poNvu43EHi9s1+ne+1Nm9gJmG6k+gJe8R59x/vTFfT9g4mJhBDRLfD5N9
vgurd0OCnmypiAoj9tqRfT5lcMKNOPLVfeMeTIjf42cfQbYkT94eC4ZewpgywgHm
u5Z0+d30ntg+7Hco5AviUp48R5Y8esU/f80Dy/B0lzSSlwEAoMSsBzv5jPjp5xsk
/JFNOzkMPLmYaLCD9nreMtzUG1ErbZgt5R0SIhMXsTTUS9PT0Jdkwzom8CjEVmST
NBI9qz+3c0Fu32xpxvkA2fvzUsrUmBHWuvReu3gZsCsR5sxlHaT/Qt/Fy34j8kHH
qcN9lEHdpL2NzcI2Wx8Y+YI/grfKTw4wEpnxab05CID0N7BmCI+zdA42436X2iUL
PL1QHx8tUscn5obqgbf7x+l5ZzjBLTYDuP4wCfD7mYx8h7NQolb0Ws8puQSVzqmU
BBTqvVDmOsY29KVpjt7tpfpztt4FPuncys9RrYrA6h5jwlHY+CsrUkOF1QRSxt/B
gym0PX72PAH7pKaGI8PpoIsHHRTLXoj46GGIvc5XKMG8WG6LF8MY037G9ZopXCgQ
+40h7mKH7h3TDiekm6Q+TpJbpKGCueLlHx1toDqE6/urNzEgnSIzN7pfCKXRSDwO
Ti0gi/iBbYDQjCeTp6vCux4RZG7vwK21Rtf2MFY56Hcrz7UU+SpcfS07siyeAGTf
20pLLaISSoATzknANSp1FhNEwr24HO+aqS8YAABldIDvi+MWen2Sp0wPQGVN2MIi
pj1ZKhn6evDqxwqtPyojPRWRi4OMZrMsK8QxZDr18RBFAQ2MVO00SNJqB7dFxpOz
fMBDseFubDNw+a022ZejonKrmlFuTH2OQ/GWl8vi1Xi5Sq61UeQMclYFXIxbqrXk
CgOehnJo//pybWpiquHGVQZBPbPkdXwk6vi1Xh1MoxugooWIzJjuxPa/caMq3jET
Pdhd1gsAmxNon+bGSxnz3lNCvlcqya8/jxxPbO4KxOrLOnie79aw8O8HzSu8qBel
Wes6Lnar3V7hTjAy5dL6h0rvuFm0E89kkxepm7vDozLapHtiRVvQcwHc0tFoUZxG
3GEDI0Sv2PXJYvjzhIsEG21KWZZL2McBb44tpk8GOIUqmiwz0wZDbOaQUAMrhcNL
cdjxSL5LYtd9tdBCZ6YFWBYOK4NgilJHe2ffZETL5Xghfwe2Mkk/NlFe3+8ONrzu
uwoEvqQ3ZmdV2g/XdJE6ET2c+cwhpsH+2m66wj9cOMBNhavS55sbHwTJSlv0qW5Y
KcTsNpz/r2pLfPZv8qYYSjrn9OO2s021+xFpglp2T+GM57EAY1qm8co2/QMXgWv+
d1JfmODF0WgsbIZTTxvKjO0F9vKqn6j13Wo7Fyt8xJVpK3zQ8jfudrj3HhBv8vI2
XL3GNVN9VfLde3Gq6W/GtgQMrAs6UdXJW0huc/sNDoDsyuG6p5qbEcMucLi3/OMD
mWQ89rnwkuWTWTAREntqBjbNT7Zzm5IFBNCwuR29I7cDcjHCphzhWVn5a3dtSUGl
dpH7o0IVbhZj7Xr6rTR+VDH9SoL8FwQoJuT9LBrCoz5mGAK9PjroypoFeRDuSs3O
yfO9P+oIUMtIQJtI/LQ/ljxaGb5MKFHFsYV3ijuKs5qfAAkgUQFlKuCN6llvcQS8
FsqTL1Z957CbHMsX29LmQ8OuVRs8UXe4cPHUqTFVIogPMr9jQCwAzo1fViqhncN3
TXp5ww0aHmgDAwYHFzSplaZbzZaJ5Mt+hr0dD3t5gsCfndLn69jho9zPeTROVN4Z
EC2Rw3ltcLOtnxQbv0eXq+QlCmdQHK3+AwRXljjUrlwoU7Jj+cGYtW5o1vvi0Q70
34BW6My9Y91NsADJ+tsxSmCE6fpryp5UkX8iveqOU5BW4b7/TUsbtP5XPovi2HT7
bRCAg7PX7WFNu797YtvT9ka7ALAbyxcAUlf+7A+FZ64B1I7G/80o49dYhT5LuE25
qDX6L4hdVRNI29yStQueML3An4sAu3Zb2jYad71mGzvAEZE6B0aBC4D3/GGXS/w3
7veyaAk781ynZLBlB9F2m+VmAlmHQPZt86zw4qHzNf1/VTXpgDfivE/xqITrxwSx
s8tO+bxd7vLgCOLgqWB+9ShnKwvDMUGu1JCWcEBCN/ACJ/MkATxDWn0SZwr2XqvF
ro36e+hXHpkenehjO/zzwnF67X9Hyvk7W0hsQ/J4JN/wahhBXywbH4IV5nXHe8Fx
oDrNRWncvqltOKUhxr10CXfr95RAdVoS8yrjLj3lyUmQ79qIodfu0HeTavM6Dp5b
fu4/vJbFHFImXcrhIHj1xu7UPJuW6VvOKZ53tKWauZbjidRg1GFu2yvqjrgqyNrl
RCTDMy/i14Owr+IKqfD98E/WVtkYqY1veCY9TseTYoAhpAhwbXyMqcDJ179S9zxn
omEUqzoqQ2FoBJDRsoJyhKlru67ZDENns2ONMioIZU3D4ruWLkUY+/qMjaSJsLev
eIvKkbFeu0hzSG6i4bRFgJeQRXKL1ed9PTZfuEtNPYxEAdglXkVqnKPnjKs9DeOY
MP1YeoHbSM+wfg8dvWgPvFAJN70gXObiqsvnU5+vezG9qEYr1LrkQrIozpt8hE16
wQgVBYbnZvFSZ5ANosUfkFIypjr/k3ZPbGWc3hJf5fQg74IQPVyQVaonn+615kOo
z4edBGC9HFgiPo/Tg0xzwAtD37cXFzu8Y7zNZcP6kJEnHpqr3c5tPZummRjJ6rq6
TZzJwDEfWAs6tzvyDLBdO+rwJS0wraRoascZH//R96+d23UNIJqwpJfyEfU1SGWt
riAoCA6xLU6bb2C6NkoDRoXr5hpaqRqHhNi+lEZ99+fOfZr8krbc6Wp0SP7V7XJ+
YavB0R/YNtpd5iDJL5B5d9a/adwwM5DS5NbPibHdf5CfLZAA6ZbwI/mG9bNnYWnT
lzxeyb3E9naRiIdRLboV8M1yWSYo8kyiVDgnfqqOXmu+HCKtNcerBAW3ttKB4JJd
LgZXTy7VDwGsjUqaKpuEYOdK9+ACQmhVdMj0+qyJ/cDnvz3wfUrMgxnEPTOWmywR
3M8bgNTXFitd55G7XI9npb8bBr8sDqEK7Ou915EVLERRP3sZ4sXVjufE1doG9C4P
TGhmiOeBSOGNr3HIF9vXcem659dUM03zdME9UuaT5gL/XF5VGTnTi3P14CgvbrRV
9cY8ciWhr6a26+h604WULUaMBK+u3Y4ykq5dzeneyQ2aZx4tAz1qU/33BUolrvIl
7ivJIIlRjkRmKQBm5HAOM8Fgx/EyZvUzfCYCwvaN5snf2TAT4uTaacjJcYgo0vwS
WkQzD3+ZGx98F/uN12sNZNZ7W4zI+TQULfsq8lZHsWcct8WypAVqA9Q+zOh7jJUZ
GyEsvLQCm5gVBmLr/SO/UfOzhGFZjBoyO4WUCN0Q5cT/bD9S3+zl6ddQ51uNKZao
Y4a9NLPE0H0iY3RmxmZKtye2qGWtDkv43oVwiCQX9Fpmqanna0D8Mr51HETjcUb5
6kAAPmRZyXuK8EN/aJAeoiYOk/mgsaHmzzvN4T+GwYFOioEBCFsVB6aVNMq2Bhdq
Kk1SPKov3+B0ed55vP5r0z9b0VQMktj7BNSMk3U6snFieU4vgC3Z5gIrcqLXF8te
Lev4ZfZ4cxFQdqI+R5PDaEPFM6oVWYkvzLnlusDSMjihVTUwX+QuyYi7herLPYhj
nzy5SXTQgtOYCZISYq5xaXrzIX8MCjNBLEjBeMRvaG4pT49QkZSAl+TtAqfZ2dst
CFsjWawspa01xYwN7+9JTMWCYF3McaTL7IA5aykqh6ZgljoFRfL2dgn0hd18/Udn
WbEsfnSkpNj5/RRYl0+xohmbk3Jl2NwzYaupbLVwJsT/Lxt0akuv3lDK1QeFLvAr
Lur5I3tD7mN6cTCq5uKqp0ulFkOF1sb2jk78Z5pTI21gBu9sFjOr8bV5ELoV/xwB
SEGNvSoF3rfLNiK5pyJaAnAlKT4eUKe212KIgU1+O41e1ruNH/xjZTt+/p9VkS97
fMZ352bdB6cYGF9oBNsUNHYId0phY7b1cKw9nQ334JNEhdqyjFA5ZBBvN0Tn1CJi
V2xSAHG2NDm/3kuEDVVUUnYUdK+wJaAuOvugk0NvHVSSe/VByTAPGxFA0d7gK1gt
0+/cDshq6ZtZ+kCp+e05MfV9HSJ4Mrrap/O4u130jSy0TBHP2Nla7BmNQqiIl82X
HgiFcoPv5vZ+IO3j9HyeT2jvIlni/gydynNsX2jqMogPJ8I+doYuOUxmzicehxYU
2eBhjwyqloG/pqAXeu3l26qCbkAv5nh1Z1xJFbH7LBpBFCTiyyztCKYdyhCTgdM8
CeVE+EwEeFWK5j5g4GYADiNN1YCmDB0XNxCYD3Vpfa0mgSDlthFojlwk61UBX9bf
xKBiO8O3SMWrASHyEfydUZhNFqtoSk+hNa1vZnAaVE0n7Tl9VX5rP5TKAzMfInNp
boU4EKMnX1jSUshjiRjqL1fp2DwU3usAHBZ7OMnBq+zRtYFNET2c4E8ZuMZXMrh6
+bJStbgulSuFdAo+Hw9Xx8wHLB3xnUIcLI+8uKcgf69PdEA2t81gnmt554CLMwgi
IqLnuhHVtP3N0JMwSvvNe0iJRmMVS6l6wfFippKeIhY9GXv/MKZiIPw13QSM/5NC
ZZnr2XAvwPYevbnPozzfnW5tXNgX59iIGMazNI9CqCM7u4FwpsA1EiLaKyjzM1y/
+2U4dMIynMFx/hfeytZLAufjmNqu+ps1Kc/qrVXonS/7ZzBg+eqoDqFzhIaSAt+Z
qY1e1vgGUtPuspuKEkGy+BYBV3N5yybwtmeMNeanQVUkuU4rW4MWQ5C3dUKzJiUQ
+LBxTrZZV0h5lwoQugzmuhdHi9SeGR7+HgcaRID1+Qgc/zFwKi52YNlM8CrvDCJ5
cCrHxs7BbrgyiE5C9fLiiRZ9Wl59R/OfI1+YlIvhQEafyUfzhZlwWJB/eKFFTSVC
sRHgnll6D2DSJvUS0TIJA9DiU91354SHDycU2Q5xGRZtkbecbUDjMSLbUNguSB+Z
4dzPNNdq1WgKe1TwjxR9pJqgBwaKhWidXxJuCXOadExK9p5EW89daNsZwlhu6DYZ
cY41eYmrDWkkTK8xVxy7kFqWG44e+szomsiu6h4xahL4yA/b2w93UtBzH01dyegV
EfNg74YANALLRLnWY/AgKAz1XK/1so/yNn+s9CnKM6C+X6VtRZXxG48OvqnBBTWY
pvzUBPGDyLulyN4coePP36A4mZwYv5VlQYAf7hOgVx2WyQPqNDSoVLcT1yoS2FnU
AB6Kxj1wW+i6qbqbEzFgw0voxwauEskaDg2fqpSqX50GUSF6t+rPzVeTyml27sBy
OnTcShOoq+RvcoEIqfC2E6oiF6mXuX1rtNULtcX/FT1vjQ7ZdcSk9Fsuv1Y+2VSL
tI5sUAMdCmJA+VBZleFZPb+UO5zz8udpUEAyaeLnodSwlOnB2RNcvBQXi9KtgWcM
9WvMcrNkp4GwsrgElhy6d1LP18/x4gpiGjzZ1yyLTkjnpon9NufEpy36c4+YtsU2
TESJgtpPDyG2AvL5f1nnxHXLq3ZpzwWW84pTDKxvCOvM01bo4n0y++bn7jzvjeDA
IA8/teVuB1gqvssVUcVJAzwC+3OVb5JYZgeW8gsKZIjDm/EHNEDbelLxbtg83Rar
OgYThcbXUMEeQydiatNtIv0aAyJxbkEhEvKo5U1/r/wW2gXdGa952z+I3Hv4orid
dQA3aEEsI27ZwAe5jeBnP63sYWqGCYkpQ9QRb242BjsnE+W7x8brYB5Yanultqs8
6BPUBzUiDtZfjhawC+MHefRgqgM52ObDKfjGAEZ/Vbo8AAxhkySU5J3U5GPavIXZ
blgD0UKfKYS5OfBDa89C6XSsknDmayHb04LZUzcvgQ/JCQ2odPIYK7TVeg6hWi0O
SvoDkEN9MlHP1VlSj2oJrpnZzo8s9/l3yNRz4tcA7XMTrRrERSUrT+ojbChYwy22
2qDQzI2jUVO++zio7/W1fdUbqD3PmatAFL941jLNUrA8W5OXrS37kN56+/dMFVAK
gMaN18WSOoC6gfUuGf7nFnw3tGb2fhMezPf69SfzSy+29Tuym9jtIbezYdp0O5de
0Nm6sWmM1lCtfoOptarhxx9EnhxvfjTWCEgcldc3JaXRGg0BgZycGiyUU3hMV40Q
I+/oqjZMWWL5kxRmgUT+jZTwa44PmLGoCJ4pjBWbCCnTncz73O3/P/7aizYAPOgt
DTDdZ4AQTBdLABSW/eISR78u3s4xGHRLF8QCT9TEEDrfzyszBk/F49+kB7hMab3K
bCitESLzxAH5kYylg/caYJ6zCx2n2+6yIr+hyZR+En9npmNMigy8t+pDn+iRKfte
wZwbxoZvKn4cVS/2p7VpFRPUT45krv7fGasSudlJmE3sGXlz+x6/UgMU1149VzZB
zBpBjfbJK5oYP9zKu1JSQbckqYPiAiIRCEKaFR+mSWjtQRhsMagl7qi8LBU+Kr94
m7T6eJ1Cf+5+z/EjOp+Z37ahShdp3U+9R8gt5DtOJvJuiO6rWP9dQe285cOUwGzE
w5C2INlGjvUf/cJLPZViXSPapycpckq5Go3Dz+GGztS86bNHHaUp1T8EVAZWId7V
KxLuNVG8VcI939q3lT9ogF6P7Mqr+QNtPXlS5vFCEYrE9heP3hVx47I38y8coF0o
b2RlB4BjmNGhHU7ciJaYn11oQORJB5b1uwYGuALgaDA5onP1KSCI61S6xsHlDfd6
MDnX1q4xcsUQ0XMSv05l6aVMKbyee6fJVfdmvKL6ptJxa1vBJ4OrM/zlFAQt+A3I
QQusiis44WHxlbe+ttD6r2hjGH1OW2YLBgZwhiL0jtJIM+Fne3JmuYE3it/wIy0g
TuAIj/laySNQxEcp5jsXMrp7DM7iKEHdBNWWtBmlv1u/uyBSVsf2nJxmUSW4UNO1
1yGM+eYW5e4BKHFiDnH4w5TqFlLg9HhkTlSFKUIZPQGE6NGnvFxZ+kBANJieikfn
SPgNXX1zd3ZE6nsjLpkZMiX/XxYH/NmBvqSb0ji8bRT7zFtDH4Twk4BtVl1C6g8x
WSjO+UB0XdI4cST2kXOilZ2oe6+vlTZnBwtkfPNVvR1qEy2D69CcnMbLVCUa+Ieh
PUY9HdQOYrEEGrTKfO5+rz0YZN3Vsj9yWOuqihSG5qYkTXLBvo/pKnO1rK64GofF
P0GfhGZXhe07DB4PBD4xEvRgzts6Qfc5icSSodeS62UIlxip+nhxcXKGk5x21RTx
y5h7n0ZD7XitUGXDen9c8QtAON6C6cmDDy7qYjIQybWT+hL4LrUvpeAwR9MhbHsa
sF1nlphkDgT6espelsTcQfziTPgYPbHAB0+Ivq1KjSxahXCi+6B9RGCxVSBzAd8D
SmS8idhtZ+pbobxiQw0wLNdMvbJYj1DBMbFUI/vZW5gH0ssXkl50te76B1VjtU2p
9xhiut1v35c0MHeEaQREXERiGW2qGNjVLOHZE9CbBh4tl+uxEH23IxkbfeGdMrKT
ZH5FQqm4mmOrgEN+f3VzqoaMImHlTbtpRDPNo6emYTTuPp8rH3eQpeC9Y/Z3sAAg
BFdCezme22aPEmt3uWpGnogchv+UzSKwdiYs0bM5Js617Xc9L7czOfFgUhKW8iwG
xXFK5GM+ygnYcPMJ+UBCLrYz7ntDY2eNy28Lq1g9EqTRG/uxl5XtBybakUdNdZIA
+X2AwvZKXw+zL5Fb3zXNAARi+IIv21+AQWr/kSOZ74nXjs/4Zp9uAALJGvbGQaXW
VHqLN9gUiq5FT6CCt9Cl08HxzBJzJAgkAx/KnsIhNKv28MOrFSbGbJ5cw330blcZ
NOW3RjlhmVxlSqecOhSvF0YHv9YAdxIt/y9Opw5dNfTBVG52pmbtTfAxW1AiKRvY
4RIxA6igLBZFjAr3kQJxaOMnom3JjFekBISSWEE61PzRtW2xD3SeKWeV/jsmkYE8
dfkfUu1qWUuqsa0jXEvRnjvbMKX+kNQ0PVLbInPTDwWvCVTigiXdEjyvI8Wu4bKW
Ovrntzf7riHhwz2s40Wm+RXpaZsoSTl2lrEdMVcSdvKDOYdMV+TFpY7m8AOsrsCe
FulUYRK+N7pczBykPziZk/E/ZNY9tNml3cc6lM2kwNTweykGbAvCo9R3XAzUs1yU
WiusYK3/wxnTux1vE2ulJl3pgoNjG0bWRj6qN3sYnn0+NsOXoG3rKEM+13VRblIJ
D035bghZsurHrgJ/fNDnQ8tum/TsqvAZIrPVXuXNQtlsvD4PDfHB5KVKt8UcdCZV
CGPWgoNTsQfE1Y6g1VGRvxbqTa9zekv2vLNH9f2MEJKB2Uzs7jCarqYcZIMTOEQd
sVyd8nowTqoeDlqfMzllaXcPMgHEu//ygUp8oyhLP+MHrGyEaoO+EHhP6serz22D
xj+utZRzNWy8HOA19rfTR8fwf9HSU1qrqkboN1sqbzlWmZRnFNRTuGwS6hZStRKy
XIjhDukkVzob0sEbwODabpYcmfgxUbmXTVizPA4kqR5yqi4ksCvTA9qct+RX1sTp
xpAdUvZnQhNPwdzMQ3ksMjtJlQr5Yz2JN81JJgZ9vw4RC26vKlebmE2H9u4a/Ul5
GTt4ALFNdhy9J0Jqd4/H7GjBuyjRUTJiBvbEY5euHrfoc3Y2PK/DcWNvnW/P4Bd8
ntGsktz2I+dFurmmhRzTq8bhpXOAEJwSmpbztyNeSWodQE6EZEGj7i3eE9icTWmO
B/pU+9ffoTuF78L75DWhT5vu1iaMNm/RkKgOTjpxlRyZADVG9yRPt/Wj36+5nju7
qo1pJUA10FmtZNe+AKQfpvhOd/gfTFFG4HapVYcScRxtuPRuAhkWEIUB/fHcvZ8W
uaCA5hPlRh+Ct+4Tu1NiVYNIKK/yZL4GGfzv3gyvI5/zsBfpdXVLAnw4ZiW74kdO
eKoqmXFkfMXWnRSeyLHDfAVQF7fZcdqihjSQuYQCB3PMfHFRnq1vUinuAObOKqqE
k6wytVuIzYqkwQnzH0kDPnf45v31HYGe5ddxpcjxx6Tt8CYMmJttczBpL5mI6ZFi
+DpVXrpqK0iOKRe+O8js15fu0L+HjVHZS2a4gfgRJknAfffA2w23L9oZ0vFGzZyQ
H/umlKF15Job5Nbr6uhi6hXQjAdTpuVJLjkMmJ5q4c25025j8APNzeDMCjLF+AwH
VawSY341+FXYZ/qHwCjPKE2u6kcD+zvRiFrkAT4Wg3Z3Nd/GZTlDQW7b++EM3SHs
6gCCyKWO9tPcQtVTDfp4rCOdkeYYQRTvjSCBZNe2JKfo+6YR7J9fw0UPMGuiK0oz
adzstiIsnQ3ejnrWQYe9VXWrnAYySKDVXvZnIDUQ8XGr8ywx71ZTgIMetRPHqs/W
F5RhAhTN+vUdtME9pl1zHHMZw1V/j5hH4OBiJpgn3w7dGYB0sH1q1VMSQhtURmgD
15+mNq0y6vjwNApVen73az+BCG9Q3cJnKe+y2HiU6w9QTYHU0fEV/CVcz8TefQBR
j8ViRZBBdsISqnytUMDUwnA6eNrxFKSz6Ns9L5o58GpX0LGXtK2Umcd1ZEEEaQjO
87arIHCAL3rRVvP8ncTbAJRk/CELqpgKZ+uqAIb1zJdugKJ80qWWH16xozpq9XNF
IL2Kaajxsc12qdM1LhZ6CflJ5wr4VdOfJ7Y6kjmrnnu8jRNFTxdRFayxZDELPumo
IlHbreH0OIRwxt8G4lz+okTnFd9z+9u1nLnBwIDvJqrMmme6CH4kqxBF9VGa0z0J
JQRwOo2qSft9Er07p4iF0TG1NQvo4cjhoUY3d/n6UenRS3hW7tzKQAs1pAvmMhyD
T/Y+MtVk0br6UjFAoccugxysQMkXx/EKenrHad0umyL3L/wQxmBxNCLs1NUux9Wf
Mk0/3CGWkTRwdFvUzdBmmvl3UYk5rq8sPWDaXl/1n2tGWimyKv3qqGEfSm9owKpN
A8/LxUTvGCdZmPRbs07aUaGOXZziIwA2sfJEOw4fs4LMdx4+eJcxDM/EfvX0Nndj
Z783BpuEhmLFabUUSHg18PeD+TeRiIf9T6gz1tKfQfNG2k1m5mD6rC5KdXVBU01V
ifCsUMXKbliX+SngPBxB2cBFN7xK1iuYi/ykn3VKALXpegzrlZKBINANkm5/7rj3
3OHUE2WooY796IOpD+8DaYAithGG6DVz6vAl692Uba6kKaReNzCb41q6IV8azFnn
GYfKYmfmMyW/fT5pYkAcV18wubISBCeundWCIY9x/WJGlh1epmUPSSsE2JXixCC8
TlHDhQmdacXz3GLfD1cD3gdnmS1oltl6GkaLJRPPZf17BMtcZI7X0KGwBFAH2SYG
p0c1fEpVG2qq7YuxhR9gHOEKRn2ZT+uk7qXl/ReMB+UQRoHiKjsg5XBfBTOL0s1V
w+nKu6/SNbwfy4dNNAVapCyOVpPlTAHotAY6YFuMHNUS30GO5Z06dkNnelGksJRp
xzathyFpOgtklLVHS973tfottfr4dDMwKti/IHmWC7ZD1OMPtIhUvMpYtw3X3GdT
vO8dEzkxq/1/qzDVOjAEiuiNCKOTxMRxgBzk2KnF+OMhYYACOzrSkcngkA6lscCW
SKzIE8/O8L+BmU+VZKf9xYvOx1mDCmVQPQVGKIUy9mH7t1oVRAg+jkf88v/y8UKN
0QnR5rKdFkcI9ouowXedUS95DeWz+cpw+I26Nvt/AovxLe9sHSfv17yvk2P77KVq
gOW37/4fhtrQNtpf2ePukl45E1MnUtC2KmNA0cQCuzvvk3/A0+v9uq5frQCiPrYP
iYlx0uvxwFcSwtPJO2OI3NXCPJbQXiN1wEPBEcM5+Vges/W8oYS1p9+rVI2dIbBz
Azs3wtkAq6n7sna6e0o/XGoiST76ZDfwXc6bMjrLqS50DAtHErB3OMTCEpT5+U4J
6smMUjlPDO3aDoOVQf3p1lCGhI+opsPrEsAhjtq2JedwyDC4DLphRse0N/Ws+BHW
tsHK/OlctJYivlEfu8u0qRkewoPAk+xgTPJulr0ga/JoXR6nWAKUSbciS8hPaspD
9WUUbhH5U9RXunajBVo7f5SjjyFx2XrWU+ujCVx1dBlGI1fnxiDZFZ+T16EFfSSH
lOb701QSuSET1+CV8eHBo2c4viNI1CuwHP5k75adecvkObL+uNEgQ31kwRH0m7nZ
j9EkKhckpTif6MKp+Q3lugofWAZcdT8AqkOmrIfvnSHFiMbm4USiM9qf7l9YGl23
LpmoVkW8NNPJykq11HqEacjgmqEubhNxrexfIV7dlBtsUKQC368C1hojMits9+1Y
+jPtLx3B+DjnZgqr9OWsXGDYslUl6U6llh5DFFz25ubzY2PBh+RPEmzdslvZ/fZm
fSi88nXzTU/8TXxsC3j5iv3mXeVZD1f7n4WcHtf65cOwSVZFmtt6KKRVdjMQpWN3
l8SlhDcmxAx+3HNmDcywxbXrVvj2SHyQ9h/SLaIdEAjEFBdbh2/GcxDNEEQ5oYsQ
xEsnJBqV0A6+LAcWKzoy54mewIa7KQBs0UdNWuCXhgs5ygp5ERrC+v7ChouoVvKm
2Ga0caC3Z+yWuzvQw21lPOX3bpnFAsBJzx5NTh+Ug2UPwj6i5ZmzuBHbbzH/qMNc
p4lBpJOcQ3Z9Qc4jMu08g59ZWaR7fXJqZYHvYtz2c7LI0uRuGFqBm81uiKXNcN8p
nOO+X74EShLlskOij58MF213hp6xgfuX+X48HkSH3BpqCasbdfD1w9+AuUvDbnhJ
w3pE5p6eWl7wfw8vEH07VJqSGYqHg3/KvW1GX/NqjpSW7W+KBzTNpedAtZI3Ondh
pPSs41QYJMyfFwF0RmSYVsbIggkQjIYidvLpi14H7FwsywRgAtlANvOk4hrhVES9
J4PREIIWX6qb/RfQfwd4hZvgGKZCb4YmKBQDUkynXr/kw3h2r5aQAmrDhW/oRISw
YR5ZMO4JmMQIOVGBAugmwXpYv418P8+7D/jimE3YKCaWnX0SCY9iy6ZkAhIGRcRx
Br905c+USPHJtZflBC4JYep3fvI4ag/u9d1JBo54p0Kx7wAmOggfY6FA5Pg2GpMF
bRNerIHEoLKAbXBdjp1Ihb/PDB31elpOUQVpvE5Y/rqxOe4NsSYuXzjE7LKqBxAT
aQ7guAW/Up/Ei+3+iE7r6QNnThQ63MhqrR6BjDagR4kdKdvjkqN3A4BJ5J/QjEgJ
Pi8fWHvNcn12rERj2KdeGn1eQus9bX31T+4+GUtyEMtBWa8K2nfr7n/7EsHWZvTj
RyAPrHIorSscy8wfo3VvoAU0e8YsWj4lvGqE5cqqQMpW79b7sntPqrOkY1wthR4w
SApiF3trHGKF7lRA6I3uEiU30kkKCb/bm36x+cK0WyD36TqlDfud9XBD2SZuKzt6
e8oZD8z9U++n4BRilJKim4TSoOTi3mvIhEC28lpvMW5Fkox3pFSHW2EvGYBD5bq6
MK6BHsRurz+HTefwqy9TbNxr0u8bmgR2Hz/Hheb1RoHNn5a6hwQkYm0JHpXStaQh
X4m0DO5Ws+KEZh/tiEOA7jrxIO3Xy6C7lPnX2Y1s6jEvAJEZ07NPM2y+BPIPlwa7
gZcVXlzWQMnb9d6q0pYXs+RnCO/I1v4wt7oZTDHJIlLxibPluAiVdpVQqdf00YyR
BiyvpFJlbiAyDDrr8iyhgjTBAnXXgbxksj6YAXrJKP4pOpKoEMEPda9WrCaQv+B2
cmCXsqTJmQmiHKFtcVOSVBkeQMo6ben5q523CbMJxHA0aoFaBpsHsyFKb6sSwMXv
73nHKI2YrzP85WDZxX6ydUAZ5auLgsn6j+QNbcwS1O/253tjz0gqzoFkCC20ymmh
kaNOmfT1T6gipSNR4e2/I/JEuvKpDSu7lRzeq8hyogbcPRSJVe5Z6UNdBRFNCuTK
PtGtEbjGq/lW6LjgVvMJvwdghkJG/s45SLSg06oqN4l/G73KyRNs+sS5x8iW5EHC
hp1NgFswfcoT017dWzwghuCe3NXpZYe+CI6gGuCQoTz3vpiL5jRdinBivO+MKM9U
41EvOwhlu6PfRTcpm8HgD2D/LvgyZZbvoaQnfC3psI8qOXALKE2OMmD61Sy3LH7s
Wu+vCsynZn2R/NasZ9Huof0grcVROBzz7U5FDIL6URgT70E1f856bQu6jO8NZmOD
joCA7vEwmoVvOMx50SFkHt8Ea25bKVb7gPK0TI8Jvf300sWYm8iKQjAHWyxykSHo
4/0+wu9fsED2CIA0HVq2lDIuRH7rO084dvNkjyIqy66uuwNdFn3ZVXa4O0sxtrHQ
FYvP31btBmmcVI/UGYeK9ZrW99VnFgorpSB/dsAqZfGb4k4JIYSYnRvS9A3NQNLR
Jeg30EFBBZKWI15SbN9VSslPgE+7ZQvyk+xfZECC2OjIJyhdQ5880SQ9v1Cz0xBv
LM7c/izbMAZevjV6xT8hJKuKtjUapDt+oQh3aEC9g6UcaHuMgw4/Fs1CB0l/4xBp
YhCQfinEALThK280gpvJ+HyO55cDA2MEaG0t9+rvT4ipxVfLjONNLApUtQX0QG0S
dGeJmbSrfNpHoBTyWmwiXMptI6gxBl26/tYYBtTkqm3hYhxeYSf2BaJxEp7Xlyd0
9Ek4xQ+K7gRgX8/ioUfpzYg3ySsOKdBfbLe+XHYh+yMpTqbr05iHL4WBnPl8Ofno
CHEdl63I/KUfC/yKJ97zGQBqW/uSmmnWL/I9qKEJwpTixFTBg/vwMzQrRHJFErhK
3HCq/Wx91WrIxnCYo/a7mfdbJRJUak+oZIh12YjNAUVMhjBMFin5wRvPT2rLbpky
NEUtCNzhCIECo4MmlaBPBdArImmd3sglKtmAtBErVEOsIdJw/YqgFMBVL5fgnR7b
a9oiPKHUd1ys64nQDI7F8kVOLlfKap7YKw9PYjihoIpJVd3kh3lxaJF3JMW4vYOM
etKu3Bmc1211xe8U31E5AeDbr/qwcZwe1UdA0llyLbOJez8zq3s/cafTzQnDbpSA
4LsOBjIF7ljZ7pMJjtFSp/Uelh2/1vRWidPhZTu2CPFVA14xOaSdDGX3POGimHgM
Pl2qRUxydTJmm0eiO9VipBDhORuJIQzuYNxec9aOLpgCZashbSQLEh3FAC59uRXR
eFauz8jvxPOjAQkRLH04F3SVfaGq22YzqkmEe+WH7VDnkzF5cDDS8Anqpq+iNGRP
E7PF8TsuOPLJzVrw5+l7/BPEQSv5JRFUPv4Pob2TIdhQ0Dd8sXwIyw6RijYFe7XG
3YdVkdyO+nnHfCQXS9wFKM+fCk7UI2izXi73W4qw7o4Gl25dBy79TBSTSY7kYkLM
iJVVQgYT1bQZp2m0ssAaA4h2qFMZlDG3tZNHJmb6XXkDUWeeKXGOhOHBaqBOkytz
JwjE/J0y55z37iRwRCIwy2+/KZwHYsZyLHcljkLhHcD6FK3Xu7aLDF1uzr8J3SFu
rtRvGk7kDPW0uaanU9PgNq4lMrP+6p+3GDLvTfcplQI6LbAB1vO3WTVDQk5RLUmc
Eoi763jlarI4SNu1MLM/WsPH8Q42245AKNxTaYxh4LvCMlfNET6D4KHYmtLv8Aah
+B+aRyvuiYJdj5xb8ujyVTi1df4cIa4DhrYb+PZVw+oQE3yHF+dRgcWaApiPsu/j
8GN/+lRjmFgzY+mcD9qpD4CIKIkWatLe4SuBk3gOODXIlKzDC/v731NLnNkQZ+6V
Ga4zSddfyVLbjmvjXrD9426jIk64yv5oz9yQNE8e/UBoD8dTKM1HRKVxbEqOgv1H
jXrNz/22lgYQf6RrBfbITzQs8WGIvz8RTL4XTbzcWs/vFbgQHgi0dX7q1WJq93ss
r9gwTCWvgaTowt79wEC3UdG4NmY1uqBwVTLqEtn65hzr9MZPJO/5F30dymAUZFfb
aVpQnfmyoVFyk0N7t0Lh7jaxFha9DJIx2n/fQYk/JOhoY87Abw5oBoQB9os94z+1
SFoJ0zhKKDJ9gPNdrUzuXgPFHgJ34JoMVQsJxGiBdqrAJdfpkXB5eCM+IETg+RKO
oDJE2wwuORhxf2hHJBRgp6sfZ1NaTs7Aesi6eenssBmuI/75WfQNaU3h+Wk+vu3e
9FDks1zP4hmvDln7/wT8HgkBAIx2tnCFAqm/dSv/dphp/tfDxn2K9vyNFRMgL/e+
P/7aXioWp4+2BK5/+DWvhZ/PTpTVym/CeAFIQfoTTXqxGYT6UyLGz1tgpcyZyShq
senT6BaYsp1n7HdS4ZymwYBUYZyJH48g9zWcWgf5DCqY+zKwR/jWGIWd9Sf3dmya
gYeyrIVzNnaYVGhCHaWEjjLIcJF3z8aGF7FyKNkbnDwf12WrGrwrt1wCNozupkC4
+kykuqmQSJ0jwDcv9HgsVhlSCDeTyOo9DKUz5a8QS8+L21ABEGTs0gJ5443CvFfH
y0edV2Q3WYs7VlJPpaxpSABVRKb3Cn1gLv2MWswiUT2JG0JW6C8281wki5hJfo5J
+Wckz18JEmZwrPb/b8jwIh7QU9bxZ37YA1StRJw1gqpFMUksYCs1fCyb4A9l8RqO
sdhCrkJTGghuqpryRFuO/8RPv0pDBDeOYB1kYGlE+yOnh77F4zEiVAb84d6JNrML
vBjL+sLNy/YkE5kK3ENO8Uulm6Q9ULHbxVN9F7kKdPOEQUVzhyImSr+DEc09AkSc
/iuzMwdgpK7sKUoEUT/dL9o+2JV2yvEpOcL0pB0df8+IU7TBS1nQbFn7dpX0X6lM
6NpRrreMJ/pX6dHomBMrVIU987+vg2Rj0Fr1iLDtj9Jo3FuOqNsz6a4SGFm/sElR
0Ju+PZ0Sy1dlLloyDKAK6w0acblVLhheZ5gF+kJGq8wnRJIzx3KI7CAY/pt7qSVJ
xi/rPKQ7aT5k7fNGZAY92QtwriiVarj7uF5xDGsy24MC5Kj3Z6jWsdWllwKqdYyN
YffIDnLbyo+ZNvM2htG+6UJBjRdBiUZ42dLu1AEz4PM0LvmrOnR+mWpnJmNbuSyc
3Plo3WhmEYjL1BBmk+qDce976V7IKhIpCrHIuvdKj56Pc23+1pp2/j2SrMZQixJV
jqyd7fn5+e0Z1HPacYhamXO1hPpAG3NM1Z8PAYD63O94/4yAwA4mdj5OWYi9rUlr
kMgUs2HJIsnZZDr/YMqMERKCpR/mvRjrh2np6lEZiMaFCN1X90SMd25ELr/myZyR
M+Zk4E+i8PXHuPGvLUv2wkiIpFNYA7s+04X2V3N7BzkAbo9UEpT0WAwrTd+VQxab
q5xT4N08bRf/KpUXkdebBIhh5Cf903mzmndlWS/kiCw0SGww5B8eBQ1+Ic+INgwT
S7iRGAObZGw66/wH0IRJOcTd8xyiAO+RzDtRGj4y4HxSYM/MxWnVBUb2tePukuUz
gIXouHrLg5flSWoPTGGHuX4G21BVENW3XC0o/+5s60J2Qym6Xfyj7gGQKImkQ3Dq
7+sz0Mbq5IgCZ/MUe1c/k9ofFuEKzpqvENF0nmpUx6yDXNMWxrp2VAD0pUut3GGU
cAnG8/KB0k5GzMSPpmv/4dJAZjEYPqvCPz7SwCaj2+qFc3ibP5IkJNma2jgZiIyS
S0OEeA7aLZcH4kg4CX6FCJm4yij0Og5kUepxYTCj9LoxdbFdPKQRC2tasngDNX76
A7seHRzHVzvcqrmhW6r9Fuye0N5DH6pzWeoDRtA4zorvt2h3p2pkrvF/dH2FIfOc
rTmhXn7TEekqR38Sj81B+7kQYo1WOas4WDCBSHFolyFiXHHdhPjJRL6Z72jbRNVd
bi+28jJHmC9W/kGmuqjDYcb/F5BLsHIYsTKGNkIYuYo9GQnKCWZE4zDSdyS9adjW
aARpr2RmYKeAGS9cDxWCxKpqtlWX9DDMwIfqFFP1Mk+xp9/0M4YoqqDZOS0uuqxP
ek4cqO13TAULf2dUoYUOwaG1uYIcwF3/utWDMH1hhFxJWOLqo5tqjqLpxV5eVD1H
Oo9elMSNWlsXhEQuhYTiL7RBCBkUcqGA6R22BaMEZMG3bLJlJgXAz06rLrTEESW+
VwrCOgN9IzR6sSitxspd3RDQT1xBDdEFNpzTkKQmzObWiEfV3M7BLYACS0otU9JE
ZakKJGCXypZCuMvlCIck8nNhYfsqesV2Kyka0OBOzENqylBrBB6cU5cGxkve14VB
3FyWUmzGGzaWAJ2wlggdJgi93Z2VBoAJ6mAzToSwD6NSs1Y4NEeMsQPS/DZKFNCv
rAX/wRXgS/Ukpz/QLSa1ASPb6pCgQSvPenhMnLCO/CreDh1pR6igiaA5AtrSoD+u
OZ3CrYsFLWEuKVPWqXm+70LdTRWBmAqV7RjtN80vgAonNDDmPHfIFbIr8OlT6CY8
X78VbgFXzIFUI1TnKbhnb6aiL8upvtLGvvzynlHDXm8FKsDNhvXNaHmAMGTwNfXg
i5d5fB9BiyaLVwD++7l2dHutStLVYzBVowZ0WVBMUU/yZVL/136aXa94y/LnjQEA
sjf6vwtNcE+LwSMwgKgbEMtV9kHGrZL9T1w77i10Lt8TFlrAvQkYA6CpyMtxQ6HE
eDc45p0+WBFmPDdcztNYD2ybf26uCFHKQBhB1lTZQ3lOIKK3WEAka/j2xU9j9zqG
ANnyAnk+gyIBPoV5xBkqAwbmTGyQ9Ubj8l6dR9XIn004JqZFJy2NToF2x4/dXLAK
6dsEf6oxFJBTN4ClGZvrICiT9/LIGKtZPvsXbn+9qIi0QhPJYmq2Lq5fUruYnWbK
pbTGS7MHoq0vjvdt+VB7dNxT5St53oWJ/lP3fB2HTdQ772g7ZxoI7clZ/2FQ7Sn8
zYRyXz+LLWfo5ys3swssJmYafPdInG285Dy5A12OQtZobyzGJZK4wIoHKexxzxTf
P0jZqrvRSr2IYXWcadEPJmV5Eg5qx7mKFh84pWIP2+udY1sOMnlAWGClJID7EyYD
SN6DgSIqmN9J7dSszbNDUy9X90JVFtsqDWyTzyTLNAzFiI+EvyLjxis4AVQQyR41
OBubp79ixRRIBtv4Ie7du/GTkmKPvwuTo9qkZwS8EvisN6flQjKR2vxbQtiGyYpx
5Omgn0yrWT55dGsI4GWtcjIik98iZHD7xURWG+Z3rbSQOVpbJT6Aq51dNoKN9sr6
jY6fkf+LGxtzoi02yUnF7k5MVxm3/pW3F5fSbI5h6Z3PwzYP1KVrOV2ASzHVR0LH
be0sA7rKJvWOVECEWvzL1+txy7XWydbS+m2/npsani0vabiOsJlI15I4uw7EfF6F
q1DyRWcJ/B6qqOHdKyWOVQtw+zg/S/oTRxnzHopV+QCFsQkeh1doXPe7M9aUlWJ1
/vZAaITWMeXZ/qCztWEezO7WK2I+tUaqRrqOSz/Rv1+Jy24KS0ieIKx7qwbwduIF
+vYZhmsy4HGO6KDuAmQdb25mheCn+ZzTmGd9G96bXFh+/AFUHXb7EeRQLgUFeMa0
lD5agolsdQVlpvsxAT/pPYrSgmzEMgovVYMkm/FjAfUJ5ktDsB84YkXxZYAaCxdr
SrOSpSVGlA8TP7rltLKKaYHIJokXb1xEl+0NoR8Jt3k9kyGYMa5zR6jqAqOlGlOb
3BNa7Zu0GixaW6N1yb9GG9gw36T6woAX7a575Wrmgnd1WkWBb++lQcM2T7iv7DPb
JqH9FIwsieg8T3yhk2CiK/fRBuZmgGEpOg/4yf5+nm+fg4FczXIDUfNMbNyaD46e
dxAOutZ+uJGV1DHoiMrKmdLGGk7MlYG148sAK/raPAwk2UFPtLYTdykJfWhou8Cy
NnEezIjWGST1GDqhNLJfxrgE0r1vH6CJ4ug4Oght8dMd0mmRqnE90bER7MZcbfpa
JhK+eDS+XgTI4qZAc+4Mh6t5mZco2udDLSgYh8ZhoDyGexjLQeendIHaAMalVHmf
5B38ufCqlYZuBvuk+/Pp+7K2zsg22OF6liMkWA0nvz8DDNdWh++SVabo/YHSuNRK
+RUW9xfjY7dWcH83rPSccLPqpjwhiA8R1o/gj2V+uvCQlCOLXMUeYp/wPR23BOw+
hRE3cOJUXCoJxjwFu6/ytkBWP0Ia1TB1PVqm4k+0bHkhKEVajvNZ9Pdhw/IfiW4Q
WyOTq/MGbXeTvC7QZ1EKHHca2ekfGbtJSJkhEVnok5KSWCrAwzaXbd42aTzd7BOn
+aSNg7Bo0wS9ss4SyBhAegcrsB+l/bxCgWTz8aK4wDqirtAhxT20C/NOc+2+TYcQ
U7cYfVdALL2tgBRRN2Qke00nEQsOt0A/wOWjSIwf05InsxX8r/kY+fiiuAWW1aQa
aPcGd0RlQdwCX4hDkyS6+ZxU1IpB2KQrCtdQ5CHbgxQsddJgX6MFpPzARgAKcAoa
oRpXTIB+h1fkc5YMJMMCvOu9sD+MMbUK+5KDTXBid+pSFnA2EPx5kiBQKLbBf9bb
Ci2SyuTt/z8qsv/2w2o0gFGFDoAj7qlpwuM8onjMwNpBwGh9LTaeSldJEN+Lu28w
5quN5FvJ85zFVSXUysQDyFMbmMVCPDoDzDF8CNAxqPXT9ewtzdl8fMzmqu2EB67f
t/c0c3yn0MAZ9DigK78vTqFVw+xs5ef5LyHQdtSOZPDSklqX20BoYTbNgPnIB+5H
m8czOUe9thXm3VBrCaW7eJmNy9uYkxZKx3X3IgKib2EkSSoLRnFcF/2EEOxmBnNd
pFS3M+8zkaCl/86S85ezrP7XzRZCXnjf209KzvXwL0Y967HuuKZn+bU5kM940bUP
S10F63+bac437uGBVtR/ULEKBzrt+PZgVUHsxokKAR7sYJ/FVBNKH2xDZHDHIItF
h9px65RTdGhN6Dp7S+1lD7tBU64Ucuxp2x7tN98PWJe/mrzN/SedHLy2LO/SD+kU
DcSUWWWnT/Bv+hAYKXBiAT82QF6Y7rD1/HcnH31OXsk6ZnERgUAYhKDinPHQojnm
ZFnKPUCzrhBGOLGwhRulW4q32Gdxg+P+mVseiCYTrrtbNphLFWpvuH+VkXfQdwty
GwFpOdrXm6s/dokjBU2mw/Z5bejgUHsXXfQ9LTb2X6zBEm2TcH0n5idNyGlJ58GW
VSV0FB0zp4ZcMz8aoEhCP3tnlxDkVfAzeB0Wa6oc0gaKDm9h7rSzOmvjwAXvtB2n
pEvqtrUQavy/DS6FDfeWkNY3/sp6msidTr8rkoJTPT0r2Rg2FXF50noJ65Y+XDss
37krzntHu9OfUfx/AadTtZywwSwgkBcOG3etW8hg7BSiQrXQ8ZCFgU7drkwrksy0
wmN0JikLIsTEW81splFl0f1wARCUYJMw9n1VY94IFtvgzGjEys0dV2DIJykvVbzN
zwqN/hR6QYNXRpnb8I4BRQAXFGSpn6MGJdLGDqJirNMTjpwJ0ilwBcMOCDZbmMq7
j4VCuNH2LciIYcpP7JfyhxfLoee0UYwt3zM4q1EKV0YwwVc40OAOF3KaogevI/RM
+QqZ4rGM5i4gdvx/TfhBFfC5Q5Gw1GC3P7ISlowBqGT9fwicKvVUV/vQVxVXnzFU
W8RTZ1Dhs7d+4tjt/IyGiMYiUXiAys7qMjrMtyk4kmYkWKafsfX/3BYT8P518w+V
MXyjdARYKTcISotg2PIY4QEOuvPmuk/iXH9/NT3JcN9gZWaFc7lTg5Z9EWXvc8Yn
AQrAHNJOcxNWk52Y3B3Sunxlx3tqM9zM2yUdHxocyYmpe75+Es1gHyHnB3qZ/crc
udaB2NQkL5LvwojQyly3yviGtmud1KcPT1Vhfdxh1bVc11SjNXlUl6BWKsCSguYF
PPAR3Vqj2HDWIukofRTlBhsN2oGxpm9WWrg+stM2LsEDL0GmwPyZKWwkTtbyUtc8
oTDmMnQAeM+ikOPQprTDLK9r1rCaG/UNM0zJOXBVcyNx384sAO/thp8Zqu9t/2g4
IRGOe4G+WMDV6AxIoGNBUot31Y17QbAq9grOCaVivRcANUbRMdDoFuCnP5Vzt29r
pvsZ/bsjlEUfs3DMklX8dTbbm8OB3dfPNqQU1hDDA7ECXrbwWvgJPmuaDyM6kmgQ
aAwAfBTBAO9uPGSix4W3pMDrx6o5RtsffBA/B32KsCAv2FwhYaJziAI3YqNH8Cqx
z5r71ggvsDmuS700Ky8Sz8iGh6nopchPYwt/rUFyfcqFoqV5x3IR721D4Qf0oWRa
XsTOEw/yJWWZ/B8BRJfFqamvNl/TVOid8O2r8VZ9kBlxXJaHC1FhoaME+1LDaQNH
VnHwZu1329nY9ZRoekglyyqvgg401eG7HeZz9sM/VelQTTfkvK39tcI6fvLArGvy
JakYPP7lAm04Jlf+Roj8rf0pJf0foOxeQi2NwXZeKHNpgQqyf6KyV9/6Zi/vqRCg
EyMnAqfUvMYRX3wBQ6/DX30UJb0P+XbpAwKkWUQXxZoBL+2tPRDWTgpadbL3++fS
NE4lGx6EUDUx2Dq50wpfHsk1JJp5rQWA/lIfId4S88EwFaXmhDPIIDibmvZLpI6V
+a7okavKYfCCzgVvp2142kBUI7xPSU8RVtneUSfz9Nu0KfNB+Jl+TZLiPmgYSv09
D7JQiF8s07MLtGYlR5Txznko7b8e/etm0OFvNf3C9m4/xA0caxaS8IhFgAC7uOr2
SPNsMqKiqRkO5cz8yV4lMujqMy7M9I+WKLcySpDVatkbjxADM135Yf3bpg5YAp8e
1ikcZvzC9XKCKiRb8Ofl2W8C34zCfd9hZ12GCGS365IB9EPC7AkH4i6wTpPJ9+oV
Byn0N8/fdyuHr8evFH2UtsT5qTJzLQrR6MgzhK9nM1WoqrOWbPb9ezqSDG7JS31F
Q7IdYNEKdWgmmUpB9KHPQtypRPo6pQFjdbz59UeKE6H6eQ3aKUwgqXIRI22yNzgR
XQnaYD1yz6IbvEn7dbWorV3hKcfn9xJ6s7H/j1pnOev9k+jmwQy9zzf8/wE1WFni
P9eeaOEJPpVvaarzRXvSfIl8vFZw40+MnQPVsHGPM1pu/n+9hZ9H0gUyS1HinXCA
2KEnC9e6pMzjsejJOrtVcKFp38DbMGO4Zau+sqfy/f+KvIx3A4Mf8Ha8iyGBLBqC
SyReLwlitJs6nj2Dpc++IRTvYHwaDqvPK9K1/Zzd0f00Aa0WnRRi7TeCnSJhrolc
HIUwJtY04ycKKeXH5B4UYWUazLU/6LY2FMbkzoSmhpaQP8R1f8ZRVFePGmP9VcCh
QPC9qoyTkjs8JaDF6+VxO68izXirdWQUK+dlRL1e9bVCo6HJx/34ZVx+19q7fca+
E02QvoLKRDAm3o4UPGeu9G97Mb1GQmhrM9NhWNe5wv/LSORoeGVQ/exT4DzcnEUb
Qnn6PcQl3GUCTkolIRgaBrnL2xkPwnnis+wyCUobEFQE2pwI6J0SFw0i3tDqQO73
yXQF6OcnmJl9qTM/f1wouCcGHXO3OweIZoijp69cCK5agU01IgMpDCiflZiwje+Z
GYGIqZBRqDcp1/3bHhs/JyAjw7Qju3vkFWBh0ZsMoDUPj9pS0xLQwjOjpQI3OgFM
/3Y3toMQy2LurFHV6zjCnVC4q7R66ZP+GVgA+aWLvymxKOXY/uMdWE3wPrznlvLa
ddi9ki/vTBgEWppGXj3dTiVV26k/Knqs/USAEomGKqS6vasLpPYRo9aithSiRDax
38/lfZVljSSy6DnXv/1s+MJquyeoNydUnagvBCX9znBNi5VOPM8usyKCysdD6nOr
j5OJUMlyZPL2mjToUMzWKFZoLJiw5ZIHl2CNQqdy6Tc502qJWsbqlmzjLv1dXcdA
tU/N1j7nu/nVC3y9VeksM9zwzJkvkL6dkMUlimyDEZ1CYFYywcdQVJi4ycA97LQr
RVyrf9soi+2PDNKKEuVpmAHB9QqOXKbIjOyXQpM9w6Zb2UQSoSSY5Vt7BHiK+gYW
OutTiBnsYyMhC+JGZDtqOuDrhMgMFBrxTAGAcJdYS+XJ3XW3edxB0ibY9wb1ot0d
giB5WQZH66+ZBQXBgdm3ZaO33GRvIgdROqaEF69/VnHtBB5mtRFSizCgMS+YrgKL
GCEHJH13c/YNTOF3VwLD/8XgPUMXz0nt9CPr2WjaE0JcPqvhM+qEOBq21h7SMBAk
84jZ4Mob55+hcw6KGHfku1OxQ+uO68TbdojhP7OkJbfrLkfMtukwHtp/6GVcSJ6C
m//osDT+tTlG8Molc1wY4x0bZStTtWqq3UbkQpJlXswWS3LBvNdjUWHqaVgLYwdU
SldHYXzEPAsCu3Oz24BaGVKU9JgKMxR9/1NpmW+GCjjWo3sK55n4N9hIvhyh2RTU
+O0crmts1WHT9yEdmJzl3h4Sb2cfCPALlluoSSbL3wYqQ2nW2PRwaZKysF9YH3Ab
h+PFUXETVK9ZQDyRWks3NWXM9dAVPdesomSedOU2OVOTZCUl3YtzzUde43qe1jk3
l73u++oA3WTJ5UTpUBaOwZKdP6ThtVW9lcldeAS/WEmQ8qqRJ/SN5NHsh9AObCIh
GgQ7KevD+35QqTJsKKtbprTcVcxnpX3DBO1rPUpYVHrFEuxBqb/+tUQR2wa5pmLu
gzYTjjC+D4+ZVUve/jWuQsDNniunZ4UByl4dM6CmeMS6lcVKi7UVwtU0fJ/m91Cf
sw0MLAz+MabjUKfyVkcWY9OgHaA6gFxjErbZNLPara/oq8LxaKc6G+/3H+hmQe0z
R8Kj0qM4J6c7OP+pFS2eyv7ZqaH4qE5Mc+Uz1okubJ/Meif0H02s6V8nulwsEcYO
GSA1o0fuUvdeoogpA2rZ1ZlgN5cjMyii/NiiqIp+7Im57LoDiOVaeZBNbrkYTzpD
2MrsJq1smGevMdxjZjEuGnubOhm+RSKSwpo5oGc6qSG2F1p0I2z+aUrmqLubLf6p
rTHEra3kGW9Twt0h39ZGhmPe5KT/kqakj7Qq7eGTB1ykdBbA2bu8OD8qQjtWpfkY
LVUEQyvLROV+TiKAKLTmRUIrliEHxiFzoccYCJj9xsV3DAPIx4GKAPYFg7hd9kC/
i44n6/o8o7gJT2fyzhAnnNJtMRw+qpfw/xqQ1BD+w2W3Udo3eELRzIuHL0H2NRF7
wfVWtSjrU+hoNCI90P/7Zkj3vhywWgi1mzAhWA42fqffiSWMIAnAovyhLQKz6K8f
LMawRugJIzkmKwux1yt1nhTJh3fpP1/v7aGOwQPIU1TYRV02diEhL8M24RkoroWq
KGTURqef5j4XnnPWYiOQQ4TlNtVFvWE9FcY7JrnFUR/A+CD2tJot5Z4JYpfEM9sm
Fp1yECyzNBeMOkfWqda8iw8lCQ+Dd5iCii53+3uXuxqpbGS1NkrX5Y0Cx8Y4jI/B
aVVu8z4+NE3OCLz3nwQrvKcQVV9eaWcCqmGfDRAwXkRSHW7EMbFSN2HwymCLsqd/
ldaoGGGCoh+UhAp99KEmC9ZZh7JR4PvEq6HC1RvJLff9PP1tfRVIt9KDAMeuH/v3
4JGvjpxqfnDKULo1kMfzSY0DLtm7hvCYuSXxg0IsnI+KEgOLagIc1y5RwlyLH6Wx
vBiOKXBf5xqGNk0KndOPqXJI+v5ULbYLl3da0zTgRS/hBF1x55WvT8vrHRHpeHgT
n2r0N9hSE3DE9/jJayjbAHmgnniudqjkhP/PqUvA4VtmefrqEGSkuoVKc32FOUMc
/vtjy4UO3zz01tAQpr2ceh+u6G+0Sj4v3rNUadVNcTd0BTmoG5UlAt7YAFZ3Ft52
tDgShqJyRb03HN2X9Zwa7ZQ28xYoJai781vGjkLdinS90umSfN60d3jG97cDA25C
cKl2bdh3vn7XLvx99iUoW5cpJj4ccMntNBpI/Uev2Q4lGeEcroJfbdmiurf09ngu
hNQYchcSxV0jqhi5q3xlH3UPRgXkBR42hwe2f+uZFtwae7h18V+ZbTN2l9Hlj7Cl
J6PkSCevwkLHss6qH2FZ7E1JnXmwrNlsJ7xPLBwdmU2Dwfo23toLClKoYH0c6wSG
p+Bl6FQBAAVr7Kx/KqwWMpHRbVIF76pXGHtUwwPoE3p+auEdk/dt1wSync5pTlT2
oI/Yc6heGp+Bt1mx8P8lI2URNwEwPC/F4dsc6qRrRLYAoKMcaWtk3OeCqUuFHWGY
44mjUNvbE5f4U7saYIrNXt0SmbnOqAEf7uFcA9zp5A2ExFmunb4l6zTzPsJWFWZq
12q7RNz51QZr4RtoY/7f/hRkDRLeNnFMt2Q1CzgfP6UeTIi5bAturY7v6j3zzwJh
//aOgeCnJUp91qQs6b9NY8X059nQd9Sk4asHGs8y32yxbr4d42Hfyf4P7g+J3kBZ
EKDI9SlSOln6gfp7HjM+FaiDPBwigxXyKWfGIBxAzfYCNT8o/smG/tAwMj0VKUUn
QLdpSJqzEwdnWhqBgHExT9A2m57vnxEFpvEdMJK4uyLp7G7W6uetk2KGq9C4H+/d
FsPtlBnAiz8BqGS9Pn+uoO5l2ZTWqoZeOnTnPs1zWaFlPe3zZMaSa9/+/EmgW+Jn
midFwBtlBJXLeRTRSa0PhNO9pKxN94RRseFJE1JP3frw62rLYbsGylCRlMzRaKib
wm9yHLVQpFVQj316qSm6wp4FJpxrnNNQwxjhS/HdswzsQFxqJ/mueL7EOSJ8aZzw
RuHg+c/x33OsnFgRo7zeDlGQZgX9XJJfBC9tw8GsIDZR6+JQ9Ni3MFXzfuAND6+M
0Xe5LMTADIuItHSy8HhZoKA3q3K4ICjlUBrnfvMwAjD3tVFq2cKSZe+20MvE4qAv
pOw7IAM9LDcb4F2/Kt0+/zDnUjsprtJhIjXRk4XkwBdvptsCZwphW/Rqt0JRiytG
mCnAlX5iFeLjOK6UIv9peuce1oJ2aHA2cmNStycM06ZRng/vDth9CQPg43LJM0t8
2D5AHt9/CvfWEsTlEE8vuRnnmpKw0RyyG62VTxZzeItQKglBDZyHya79NRbT0Sz/
eVYu+Z8i60IzSmUsha+Y/Wtyyj1giZ2Y4smqasFmxsIfzcIVZEl3Wx4UHYzz42xo
e3H5+Ra0GAf+bdc5g3rnB01mc6/7CevvfBwhIzwC64cPAFEsK6fPZy5ncTfrWqYb
YnQKapQSbV0/WcoV3BzwFGyHn/7Dx/+EdzmZDL7VFJYjlwXl9pqLqnDFPQzAQhSb
NdfP4jB80LsEBox/feOSWNaiVGWWRLIhBQ8DTZFK2gLGa+8nKQE6D6i6BoUyM1V6
1fsByAwKGgptapiedWI1DZwEjTnKlCoJN0PIkQJDMHFDG/iYWrIHI190bHcG5WAx
1tglpuAnM2c0EL3t/tB4ov4ldlQOMTRlA6EfxRPmpxPvzoIdqqAm5d/xBPrQYK0q
o4Z4POBbkag1GMZ6R3IYG/8LH7uMC9EAlld/yuQNSMIVlKfD61DGLRBXVf2VaFTh
YxGWUt3wOk/SbSkpNn/+xH2cOXYOOcjHEpgUEv/o6DTUZ1U3oFMwB8K3t20YGnbM
kYBNTR/bk2tLnf5zULu5epvnAhkAbieMDWe7feMUAOJ/+6nwrhKO8+Ki5ZrlTEbA
GleBkj+W0SheoB7Qrjrk9RbDJ/rTB/lxhJ9wDc44dKnzR2lDfhFYfq/7PDzbenPt
DxcRsbeH4CMXqxEVQmlBqTlnVb/yy8qf028eGxFkMS42iCm5k3UosyHCpaVrCgRT
K8cGcRjcOwgI2VrRAnfPXe6qHKaHngxOvbGnsQt+Fg00Ukcv7rRH+Gq4lpcyAmye
jH68XIfYQErgD9jsqXj4K2n5ig1qMtdFDc4bfUsbe+sYKO/CdvmIXZhF96rxr541
gRPWxkrOBlzHnLJHPSilf/6AvcHiH6UzjPXowbAF8vrKLTFFgDRdkwhIEa5nOyjg
aeW8JQzlHeBcKzBKrZk0l2ITNHVisEdeTYPqO7BWI0wVHb+t0xPrMao4vtHPhviG
JeURgRsELXnHlmTUj7Ch3XMbUbVi8JOxypnoMwGcujoJvEyNkJ6iVwlBolfJuqpK
X4TKDM9Aytv2OTBAt1BB75lg5c+dYsZHrtEBOZD7mCpTl2TB8nWIi6NUl6iPagSn
YuctXyQUbjzp/NeiPsYAeCdDpjoAf0bGzqwOI1TG6eLpuV8TXMP6gfC1BF1GqcY1
T6jiMmkKr1Rb6tW1PUA5OqA27P6Kdnj0U1es/qy2GGA/ZdAEg0MBBfkjXvj2Irus
UCwkHpjIvQkbDZlqX+1Q739yQjpBuQGgH14zX9+5p01uIaING0jlGxI0VKRj0/KA
5SWCspoQUJ8HNNSpLY6PIiote61slFc1AoMp19RY3cqT1Txdd+fHCMZ85UXxf/IM
C1UHgkpPoPfT16sug1lngMOjCP53Rd8ist5KzwLNh6f3UXSr9NSYV1ljX/gqxSBp
xC4HsnLvi4zTLyRaA4zia3+FlvtrVpUxXNY1xZeemu0dTZwQzvgkdOMcvTAb9LrW
/INY3XM19k7+n2HBeyxNYzRtqQMJhUDEoyiLa631VZPw98IWirP+w5lTrynlFlsa
PrxvZHL0ml9WK83KsVYJIdy8pOHrPUZR1NGERFl6BHSDzIzQBQkHfOStpF/mZy2c
8nDRD2QkIrc86VE43pohbh/vTWRGpfZMRXq5ASBBTTXiLCUJVDOsXKZYFe3myQoV
WFvb2hQhP4K/j8hCUaImMvtwfb7EKPLiGbOQn0k/tNm3PzIFCCZcPqlCWRyhKHxz
F0aDJLgnzuvMU79IaVTaDlqUC8lwXOf07W0CVA27DWxlNynWpSh0i+t8T894med0
m1pUH59Lvc0ba9HaMm0SqaxfEpNw4JAnaBy4AIc+cW5h60GrhdH64IQOUXOF//GJ
Ht/9ASH+nFbDCZb75shN6G+QkfYwxyIPFwvfofpHMACvuztMJJ/h+wA/w19LQBJi
PuSiYGxjKmbKinOdPFYFm4P6hsF0fK89OpO2qn2LPu0N/IhyIGl2x1Ooj+J9KwPt
kFdWaNjnS/lUngl43GfnJh6jzA52WBBZYEXA68q23Ofg0jCOpcgHonrJiENBytOl
7W6ytYsU4/tZRIFviE6S6qlOvKVt0qXDKMrAdzk2CvqFYjbswyzN//ks0CgmZXbj
nl+GFjo4hxBj//sXt5qNgLtQLtG/a2N5VKmNx/HbNvvd00rB02VAXj4c7LI1kF29
POzeJss0kmsel+Pj2Z2jSemTVFL89Ndhi/IRYHDoBRKW62xO+md8586FWhDEGiq5
ZF9y29BY5PJYCutTrGdRhYS+5zBUxPTq/MNeZcTGpKDewKYNqPyOIUVak3YlVNhb
2TsEtTaRLFFVqAVrG31iloJ0XYNYNhFh7D3V1cTuod0nm+dIqFAmR9kDDzqjFs9c
73TvgkPRJSZnB5g9FODscu8r0QHoIWL18nwyeyW0yLxEzlSbWnAoY3/RWcDcKrHR
5N4vPWiN4q5eJB2nom+eKY+O+8Py+yicymb8+etwKNxBFX69TuDyOYEMCEqhtXa/
uO/LRGhpvXbfyeSvu2CiRcjVLMuDLmoPNNhpGVOQcjdXSo6emze9EgIpw4nPge43
0ppaMVaOHZueIOET1t0axZvYjCtstHdwHii3s8JXGsth738QKTFu50xPhDy38hBf
mQ/YOnBDAdmu4sIpZmGTmHZmN7tVaGhpGHn6vypaowadh0+x1VCVTSfhzKjWJrMg
C6vMEHOH8eflBCGacVZw6oNt3hVvKN7ia6p5VN9heytCXNgCRyUsK493KhYVbAve
3a/jp+uKlt/6fvjgTkxpJTx+DANyL50pIeu+aQOAjxX51zQNHbd4w/S9mya3ytLl
eBSYpJonCkiUxpfurM19AqSmZ+pADM0hnx79FCnAPe14zlcGxAfwfEXR6OW+x/Xd
BvjGmKVh2IynZMLzzjMpYdNceyhMHCIhJsEKgleQMOS3dAiXYUn+QRpwGMnpy4iz
SS8o6ZLGqZoboXRnqsRuST4cumCeTP3OBcRwFDZYNE4XZpEAPaFrQ5MrSmzRHAZ4
WkaTAAI9Oa8cKweG7FM+8WeU10LF4wORoQ9vjtSHPWrSNrfpKzFS8d3Wtvy6IB/W
q5yKGxFDgzydgeUX/e8ESw6WrqYK4ZGWsk94w4r2sgE426KWvFV5mrcT2eullBZa
zL38bb2C7SIgFBN5rBRLy9LpZPIrzsv9SM5Ullia3Mk04eJ06IboGfCCiIBPbywM
5I1Nx1206lLUWUdtBCDiAYCovw3v2lDAG95YP4vxGklRTnF6EF1SUObOzKZYamGr
4sHTRjaxmGhkv+tmXFE7LgKLKIt2/h5stDO3Qs0yDMObrbreBSzPFDYjVFI2pQsu
mRmx+bgdFSfbuCXh9CHByZqNVuWPW7LeJvOZAVq31ZweIIkp57ye66wg8hFY9p6H
zFp0y+sl6tMnygkwiL6SEJ4yQlVupHRj9BMtxM3OjVLmjAOWivOc3+4j/BgiykUI
6sS6P9cjV9Tpz0RFbiDUl75VNqMD84BHxo1IAuB2WsoOvjJtDsFCIQTr9M0SSO4C
jeY4Hjq/wIoABOkq4SzVWQ7om9G7/WdXMxWqPhWtFSfMDG31GeeWWOATHswLtsCY
8zv0MCAiaFy4+nufu34x/Be6b3UK9h/rAd2o2M3T/CwAzJMa/+lL9H8JGMoHdLL9
NQd78c3thzQrMOP/oJF7o7P5gXcMaN96hcRAxrwa7jCrCaUwP2ZEo7Svs3O+ZOR0
k89TL9lLykPSJ1xwBjCkf0HtmWx5A66vPazk1Cvquqh3bkn6vN4tJX7TU9HeZKlT
Op3pfnU3GejmmH0K3UpZAVW5DPCbyGEMs2py5CCBPs2V/Nmcf1Y4fJmHtBMr0sXE
YkltYFIYv1VO/iuJefug4iBQyDnA1dETOJursIeHKmxPH7KgOOZNwdS7BhkI8XjA
ctRreLGLsbnbkVqSON4IxVz0gH38mhBQW0b+67tYo4Wn9GPSopBHuXDnQJnnpCGP
OAwBSz8MCC5xUWX6Fxs7a0y8Mo+WhxudLjrFnD5ANY6tAf943XFdsRUl85os2N4j
XxsXIZzU4HaDrEFB2NRGgpfL6X9qWg/ipkpBEwR/h0EF6PhmA/VRfCfFg1veSUff
w7BeguWIEQBR4Yn4fO9P1qOzfBu/e52CvmllnnJ+CJiw1WbML5yFTVOUclHk2I06
c4BwWax+XrmVrBf1936jW2U5rEP+Tan8pIUCAnwtks3OnNlabj7HQq71Vp/adZ+9
lifcIbP3LjIe6o+SU3OB1TVZsVJxavOQJTM4wqsAUztC1RuVdbys3r4vbfxJO67+
bDJ0oOSTsq2R4d9UKRoly3yHQLpWoPW7PP0U2oN3hDhTSzAlEzAMCxxsbC0mE/HP
hJHyIfAHLFOHQQH1QmQZu8wo0ihGsmFqd5OirtBJur3xMIlgqZponqQ1XaPoJFop
GAL4foDvwQ7tTZH3+CehcVdNyRtJT+/oAnFNPKfVaiLXyNuEIs0Q197Kbev/6zXG
kjTG9bdfWz7r3QzrxaoQygu+MdWY3DkACpN4kOQklPf8IMmg8xahi4kFSFgKKIvt
6W314ZSYKi63NGEBCogW99E/9v8MaX4g/ImTd6uW1Qsku1ZcD1BffUydRn2fIrFc
/GTFaMWwU6E960yomUmjxStGyFmz6u2MPUQ/7rKxQ4kRJgY63RKv45tcJxyBSAs7
tVLVG8bYsiOIswr0spKKSPv32WQ7Ic5Z2SmfGtdswioBUYj6TMN/UedRJFiOWAsl
G/vX+L6G4/TQxIaWPrVsy+V90/Dw/O+6R+TxwOqb4+jT4R9liMfdsg4hR1YgSqDi
mQ5X/w8bX/qqfDC/hXaihwsTBoEE541NaEwL+rvjQIE9/uBaKetSVkJhKqbdW3N7
Gqgf0kep070hkTtDwXA6cvz5kzMGetTVUP8t/wQgvGYpXFRxJ/CeATIf04DkbXEp
0b+evd5eu3ZcR9qrHz1dx5ie+QZF2ZGfysTjN6/A8HUZ6G9MXEnoVLlaHFnaszDZ
Y/xBSL54xye2/2oPlHyQxqFiW12L40QQnySXhW5M+K2D9OEK45QOezUqSHQvRgwY
UKGyX16/a4+bQRHU4lFxJbjaTtFuc9cvN+PxAojFfgkx7Oxp43mKiFmEVEKDhU+F
vCNbdSDwmhgx+1NAcGwyftbagmAR40N6hggOMMr/Uun4UL/xppQr1I5UHJNtICF0
nmDgciKi2KIKazTA4fWtd9nKsnAb69k4YXJE0ABpkmsT6a7YLjMVNsP8fNGEZFYR
woPRJScr3NdyPkjA+ljsqDlwLxVLIud3I90sHWz1WeS1t3Gh2yl9eYv4MPfHvKIr
iKu/fB2Wvr+KreOYirEaV/PeHwc85AIEyWxwZkLQxGO4Kvnbc5GsYf0caYsuuh+F
/DyrgQqaBYUpoXilckEA29tG3oJSX/qb2q3cHtF9+r6toNpnPJOFfbeR+cCmv2HT
bMAFtwXUcGUADpAH93R+Y8GC2DwBmVNFzp8kmr67iunqiu/YyNH/Vdb+BNAZ2OkL
VnzwPiIcQjH8K4Q8gi8MsGp2us6uUL3MEXf9pnE12LL3up9rsUZT/9HShWIzwDKJ
WiILUxsRJnrhYRbMs6OkvT5XYHSSYQUu6qwdPZJaVeI16ULXuyTsmvNo/MG9mDSh
fFAd31JFn4WY/hii2C8G0dTf85NMVG40vkZ0lhcydTmagBomTkvFssH9lklBG7Y/
99bjX68B4HD82VhFSUPuBZmUILr5QHOQ59Yh7Jsq4Y6HLt6QDiAEs1Ox8J/57Mwa
2i86Bi5OUuB6DuQtOFV7jTqltDEsYCA8Z84sapA5SGhqIHgit1+V8ZaIpKmn8odV
mJiFixLf2eF79DVqGAXJQPjDv39afyeSSB8mRiMSEHSo74zlXhnAlKHNVGfI5RLH
eIFbTy67cYpNapRR03p6xLWLEhsnJTy83VeDQh+iXzvcjjW9l6Rc9s0TcwJ9kaK2
aKI8pWJMlwlDFMNzLE7kXumMI0GkMFtzTV7vkMenpmJDPydPlhSn3BL5Bi/JHJ+B
lfy/ilg04a8oX1JjmF7IMSlRmQdYxa5mRMzGE/B0gaPpPRjaidAyfsTIDfqp49R7
7nk0Tp9wlUYYdBIXuCaUyRO5NGug9GPt9S5WKG8LioS0oHqXWZee3UZ0JLd1rJIK
5cE1uxrgoSyrWcjaMAz0aKDGeEeO2UhWttqhlNLuXfrgNzWVOsZVaEBKDPMjVbNA
IQWOmpCguyi7U478sIZgeZE749u+WKo1XNAoty1NEeipsugX+LK39oN7vDkFiD61
Z0XE/XNqtTRZThveYucOQTcuyRDLdl/JJ7yxAFdLxemdv3lU6q4t6+TSGqkozdVJ
EbRBKcHwy9qpk2XjBYF+5rLsDn8+Fu/smJ6hzbCfdcBYxsJgL3aJSa9RkabK74cU
ii0W2DCdPBoyiY/cWSse3qyKuOgvjXP0j7Y5UqPcvHyet+fOhzh53AzBNReq1i0/
Xpwioh3WQCIzbjcytzzcakEEQ6Gjpj3cHV7XR8KRxQj4iap0TTl7w38MorIPRgNg
6JAxntRF+xjDrXKaHalxjBT37TI6E3VdnWUoGEAbNVzyvfssqnI0alJNlM2pyEqr
4A/uEg48SuQKl+5++IQ40ocknCiGUjLmiCRNACUr10wxS6mm5zhI2Wsq6+JJbTWX
n+jbgYFlKv7D5TQl6pgKtajPIEku39RGdL87pOJGzAziRfcazYOQ3+wM8rTNRLb3
NA8qtJMY6b+UY7LEHZ47rufWq8HD3aChxWMV3fNY/Ezvc6O7PMyrBgDUnoA8sYUW
m+vUfqSU9YRzBOuT9j7W1pkqoCZBM2kRFIUgS2NEWltiNLD24YinY2R0+GkX0DR1
E/qppgYHB38vAxeCSVq0/2uuTijDYsfhJa7kcMI+JLNfJ6xrNEoQ8XL8z25YTKZf
7CqB73d1I2sMjjDlq+sgKyGg8+choXW0WlHbpigW73+QdzmweDYdUC2IzhtmYlzH
dDyAICguwflir8ox3B0MTVLJeWvPy6Fs2BWrxSTdjOpF4+tBEo50Co0NBb8dbssa
FMdbcUWzqNl/iVM8ZdLsxnuN+ETXUO1STRybz3hbtDJhlqcCfSfMmP0x2MLMEAr7
yoXa9Y0dwicVDETsedqRrPfgdtqlRBfRJlE2G1urKOMHQGz5qlHGrUjK3PnBL9qg
YRexWGm+8y1XyMQ0u8pkF72etFMWMt/L7gujZiUcNl3+V8Lb/6EyhQ2YWc7z+HNS
1cY2qU9Si2T+pDfVmOQNadTuLjhpWVCSVXMYFRNIs3i96xkdMpYzImVP83sDn6YK
nLjcaRNbQi4jBAGha3sjW3ifJ3FDnzLz5bS+RO8+0yunueNQJALxO1Po6MfDsFao
GlUbTYg+I3km7o57uo0ToAaKL31nyfOWt4JBPdO32suxON1Ak802B6igEyKNmNQN
J/JbnWsMWqgCuvT0iONw7v7g57IFJH+IsZkvYimBHMuudkuh0Ro7s24nd/9nYVM9
UxaYub0uLPN2NjFJsDlp8E933ySNZLWovD8+Ja+E7XFKQuhZKIa2zODUulQedZYT
P5OFKwVc4yZH6XVGYuErrEyyEuMOUSTsuTX7ygShuqJJPFT7i85z5IarkyLwUhtB
MMd0iU38wUTgOq8/JAcYKZjw1W0UQgAJ203Gt6VtRjdn1C/VTibQi+/pnB1fyx3q
flQOKifbnXRF+h7FY+GMrlWDjASa8ibFpX/mRGzW/4I7umksHYA3H8Bxy7plUAIc
iM6tX4D9/oOht1GiqV5J+/0kIgZXMI/nponOBL3D1E3FUn69dQyKVSvhIMj+qsVy
0RTQckkfqaNQKCBc6jBziLgvsP5SQsq2FdaaovIrAm7l4vWBluuPYfHQT88ZymtF
zkqxcxs0KKys5M9Pmlt5JMD27dMQNlX3ml/dtX8+2eZbyNGZOmS039QHrV6YJttv
ktdnzDH0kVHM8UnYxtlIE7G20ogwkFi2VjrZ/Fq4FTd9bYKlKJsNaGlOzP5PZRpW
xrWiAWEM6N/HLxUSbMYeDAaNhwUz0tCF0EPmiat+RCnYAFumGa5ab1LJXGlqgGQ6
h6Fg9iLfxMaqKSOEjXth9rE+M2u8JdrqUXajN9V25gS75IHWWt1r7OSUE9mkYFxJ
31EM+XfjnYCmRkhr/PLbFATJSnp1ruCHlvL1bMqJkB51ExecnEOg+uk1mG8DiN+G
hGjuEjCNej3bsU5RkCRd/PLfWpf2Jj3CCNOFDkuia3fG7iARfJL6jPqtCRKKYxov
SJWypNgjv5Oyu3dN6rm+9EGKVrMAuqH5LO4WhgTT2GwNC3GRAVfSSIHNIk/WhSzS
3bspdHwywTLqkAUiKrbTuYV6lnPh5fcSUlDCcbwPcQzRHlWhawK6URiRiPY8SBHD
vwg8crZB90s91GQAoNskmGXRP+mf5XrDbCPZVtEv6/os/WLLrxAGEh3K1x6Y1mkf
R8bhLv08jOSTWiWCpcmuAy2v6HGW/OdMYBZ1ce/zAN7BOKYuikHJGYXW+hWCdVNv
yifEsZD2hywVEE1y1kvRK773qdAWRebAcrvVN+bgqdYWtHDEfEwR+4fSrH/1UT51
TMbaKAWaoQXVCoKPhOcNk41Bgu9LtbzYe98zYiXktky6jmITsh+W722qdHnsUrc6
eoohzlAFxj9BVnQI9yOekW08kNEiipmqE4f6wkDbDwKRMUDK400IdML1Eo3DpUfh
lrJ8Gv3Ntx0TJQv2YGpWqpWHpbqv7+1Qsw70A+BBft2anww51JxBgoMs14cLpVLl
TAdiMv5gSwtasht1GqLBl2tYyYV2kRI42cjKI93tRMfF/TXZVo5rl4u7/KEdnkVC
IRcSiFbGkCvG2nD5EcW94PJL4cSNW261KeZuvIia8I8HBjhdDnBPZ56yF+JXhZyp
mHEypKUHe2YbFMIyP9aOl0LIFUCyGiV7fMOYM5CoR+j2qL/84S77xB3o38BnuwKo
LjnHUijvwvzVH+Sya0mbrKQfqFF6GfgXwSGSt7HVHMnetSEk5DuXxXxR+bQfheRi
64ZyhtcWa9BYGGbxg14h9LBItP1Kvbada2IDN7HzI/TRSfpB76oaV/onVWqYOWZJ
4a52OpGNdzPaXSuoACFhJhayVxTwEN0YWGCFRviY1VuOb5SuTSTGmlngcmDNsUQJ
AN5c3kVxUyUue7M1WBH2JGLeCOSxxoJ56BIoRMT6jtul12Cl3v+y9gtlEN9KvNRL
h5zjhksUmtNdR3slC2hN2fqgXeIPE/R8PB5XLRUjf13zaUh4DYyKPxzZJDuKVvqH
frXr6/8jAKc4Piq5XibiLkFqfEybaC0VHCf+RcuZDiUmknFQwSzRUD4jdsIWXJyz
iKpHB2G85m7ke8zw7o3oGz0Xc5UB8c7wMyHXgyEMNZv7Nwtw1MUJoN3Jp5bkRDNS
KEtprK3TrIYtTqjsDq4AcjDCUsfc0IvMUN6wKxUqckOVL7V9aUsfOuZh6/aaSA2J
6E+96YqHdi3Lx/j4JT8m08wWOwiu6818MfWdLmD3Cd31LEeEhhwX8YQmbwKA9NTL
rbZTk+u85lawffHzO1KsH0CksIcYYiOmd50N8OCj3Z9LEePWmM6TFm69uSle/7GO
meqPxCRY1XoY/g0xFaL+RQGwVpInk5PEpEs2QvikZxOYJVUQ1Tzb4NOvCHf5Yu6t
gGINXZULpBoYGciMj0MqBgnPm1hDGcrC71fd9Z0mVIgYciiabl9vBVb8jUoHgTrU
ccorEoBLdbZps6HEAoEpVEJsEyN2xVHlhi2ljVSIMnchIvSHWzmQ3F+4nJ0I16I1
rff8bPzUPbrYRckcIYfqbGFeoapby0EP8ZPAjOBAR6sBOtG4rrr5OippIAByN6i3
DOm9UDdmtnG/rmE1AGCGj4+rT/OPClg1CbLsdemSHPUMCEYjLd8Ldx9eD7Zpm9IB
fwdu2t9zJuST+3mMVy44NfzhCmUX9l4hYH0WfhzssrUnN3EJI5MOXw0DSmwETYtz
VWh4fagwMOYFe9NF3IckyDwWnveDYe2MojjRAkPZs5R8uwsUqBu2I2DHODZu8BII
bPE0chtxC1TaY5pPvboBfc/NOXlhaV4indEe9nlM81GpkYstdswsTbtiquzjIt55
EzyDI2YRXO2nQ3U5YMqLqBBKvSAdeIoZIue1ma47oycFCpOeJobk3TFid8+opWF1
qzu+P3Ozjjtj3cgVGC3yyybOd7qctbvo9lELJu4cpF3QA6jmi/lefIyHWQitLpqt
KAjiyRB3Ojt834eH33uFJkz0NBhzL1APAJdzo/QTha++8Q7zKPWfEYseG6a2TCRK
ovhLDlizWoBYP31mtM7OR0eDgl8toOgWQrvfvV20KOpLDl1WSons86NFBUbz1EG6
N5Jumc78XqQOzsc0fCGsDuB7b9kaXdrYMTFtamdK/BGsyCHhHr73j3YpEwScPjkH
QtQFbLyQS4ns7wqs8HCEEHiaeWPQI/nlBMj0uayPLVM3lZ8hNe9aXaPeDZL1Ano4
bv7E1KmNnrZWpQ8EyBhlk99pSHoYH6V5hNwCm6TEfdt+/TtHfZIcFBu3zmAl5P5x
w/lVKbS1G14gf5o5P9onOJb7XXQJQAtafHrwhk2r8YOWpbZBg2sq5gJNcqjFU08J
gyOoatVBcbnSJc7e1UuuBZ7ec/YWYREjADoZLVI66SskqDjZV/fItcWPtZK4MjYU
GP6UNp2tt2lkLR+Bh2Q5F+uKRIFhaW1YAH4U1zOOczUfGh5Ggs6Sr2nH80EedM4L
4M8eW7We/LzUd8/cGa/POtusoZxCMKwRtHeHLb/mogqPgF8W41lcMLlbWBfF/EgX
ZGveaiEefqUxr3Thf5Mwyz7fMmuMe5EGiEvq2Q8AM8iLjFSpgsb0Rm05Dg1Afn5A
kzdxB55/2ysL1mgNBvrPLJ25wHtfr9CQqHeVHPIv39JnsHUP8TKWubwlQ37ACoOM
nhd3yV+8fV7WKMXesBeixqFr3v0+05/BQ9cnW7HMrwDe3uqvnqQzd92mhHEQflCR
FG3jK++85WjbFZc574XTA8s8T6wjqqYbG3zlYYYiUbWsRc4Z+fnCtnA9MT5zg1kx
TB1BPROBMPRgfauAMwPJfMwVllsDoKdhOjadxoZWJJmPPUaiPB09G9sjpY8XcyZC
t1YSBlEMsOON160WNjqcWw1HlWQ88tWXmYOsUGoE7100UzOafuJXM8jyiezk0V7R
1YUV6SQNqncnq4yXOyMjlAq0n/fyH5S0R6mSwVYyXfxczdSyJbrHArFi0uK9Xw9g
bIxihR3lQZUXwQ0igy7oM77ElpkhcT/ezWQvZy6NZlnhTCLjoNqXz81g8WRc52gQ
pjjjmiCgBYil06BLzjUydZMDQk/eT5FibRwM4PLw9JWYZqShS6t0iTd0EA9An6uy
8r8Q7svwrFlDQNOG3GLGrVVYaqwjydawIOqTibARK2rsSOQKblTK/xWKTqWhjszL
MIoalIvzUCHmMNMZSyI6M6r3tFhFfhnw8ZgGUieNsVt5/5LPHWtStkJeh5DIGL4d
itEG5/1xKsv+qXkdxKii+ue/c6Lgypzl0CKe9iU1BkOD6/MmwanZb1MqSV71CnXF
ai3aMSh4U0lT7A0spUzd1w3yeQSLAwCdfoSJfyCXcKHxMtwtH77SwDPy7if9gLcJ
KGS8zja1ToZQq633Ejeoq4WtJE24yhq3yAbQjCFhvBAtJuBGplIdnfBeUChHW57R
TiyVMTPoDHdEfGgVUcw+apgHDjpcNR1cLa8fHsNJrBGanLfAo2EMWfAIvgSATDlq
pKWrf397hHFsrvF6YxqrFXRuFmTu6rVVNu/Gq4ERocztZLP8HcrF3rsIVsK+buh3
0gMHhicWw3VNB535PlV+Oy55iKGJwq8gUSXT7CbDsnylN0d6bLJw9FeVTbmB/Sck
qOjxDlNusN6MqhaSTJqbqaPSruwvmNM5cXAIBf9KGP9z5NORCfeer8zdcG4XxqRS
vJrq74Eok5Z/0kKqWuyu3NCCCtnA9g31jqeqwQ0IjLc8vdQir/Ka6bkirUE4u8Wm
hK90XTlCX8q45lrLOvUHEnzMJWlGpvR9Bo5GDmRaUD2s37Wa4BU2CGwExQFJuEEX
a8jS9DPXJwAmvyXOQiZLKcnBs0RaCD+8ORJLgmGnuOXIYr++IwGxNcU7Q2J7rygC
2qO4faXekme72RYSyXJunW9TY1JNUC98PZjNXtcOgiNRgY0813DJyYcV5boqTBZU
mToSuERjZPPnU94cov5F7Bn4AflHeB5Q3oXbXOkzYIu+YpaDjR+j/GxqW1fHkII4
PSyeoPvWsiU/AGtXA03Vow9ovwQnZ+EVW25Yc5LSlMpRRizV2CW0TrqIsdWQPs31
t+LIwhd3cdG4oahPS+jO24+2cTUpLsARejAGdRCHrv8kR2YJko6JiqxWOPd/PWru
ayclRKEDwNyUjlFip+FVI7UX1scWDouYMcEbORwb6dj54rRyT1W8GW4rw9sTAN+O
fM3ynBk6o5PLcXuVF2rVLsPVbDYjnyxsZzJ6toOPySZIVU+VZaOSC5TRzeh3VRAC
DA9pGCJz2sRh8HDy3r1t93E2mK+DMkW82mbSqGDqkHSiXJuVNju/3IE/VPyPx/vY
WXWkfhtqrS0QFQ04KYcC2UyqMSmhVboDycrcQ2IA9HCZHIDagUsOKxYN2y71akWJ
ETgb7p3UD9v0aqiCQIqwdteiIF3d/cnDY+vMIADi3eT3GleMuw9Bk3Nw4pLzBJLu
+IZyY8DMdVBdqVaQdwuwDaGN5NbImn6bUX5Hg/EPVFDLWaZAGFbBVfgTKtFp6S+U
xsR8TLJObP+JY3yrPav530ZvDphdGMiXv9/x/54bxWApCu0hjXS0GfBqkbeifX/E
XjPfDt4J1xOqrUZO14np5Z7WQUbQoe5vEvhK5IVzAVw/n7IkgoDgH3WmZZ2TkfRP
YH8+rV2jEVPZcRHej/VZsCCMyGJ0wgnsm6yL2ltnTuwQ7w2q38QXPEz2OSFgOxnt
GPksCDQLjbf7nTh5xht3H9MdQ/SxuG6GJpH+yr6WnnumdaW+59IOXbURDYJ81wPk
AMkyowm76jheRgtfBfFfEH2XIjf53RbrMpTTPJgvjmXLABRqiAl6cWOHqhLiBcV9
RPTCXiUVDlWSVOVMbEE47JI71qkM7HqVOMAfynstFsBi52mZ1io9CoDrkcvv5CT5
9xJ+pgz/6/tSR+RJ8e85Kg5vhsHSErZ+8f1qJaD7RN0YyDsdmSuvo5qsCvXZhQJ0
L5lMJBat+MUV/oDEDIyXCEYfkaF8sKoF8ldoqU+fusNApfRwsBsfwcWQ5AzbFAxU
togwjC1t9OsY5FT3yl8Iv2l/RqMrqd0ZixI9+y2CO5oNctKHhHRl0z9I8XISIxck
6tjUDCQdX9UlTek5C7qJv2WD7uBWh3jmjO7uMFftcFmvSSq4d0SrugsiIR9pzkpr
EvTgJZRv+qNzQYTkLRzHt22N3IyRWWo//YCnbkkkUhjXOaS4HJHnDfwWgXgI3BVm
6pPVw8dtVfrV5t0Eo7wcuiQRW7Ngj06DAztn+c8KC0gehlPJimCFRFR5NQxMNT7S
ER5+wFA5L5IDIDcGuoL1te7hmdxiFCqmK88JigAsgEuKRpBmnt+rDWHzK0QBQobu
KlPsQOxttMBGKjg4kV+P5UWERyY3EHTmT6QVCzb0tbREZOdJSRxCnPILg9aJPlOB
YVMCE3TuoU1YVbSiKrp4/LPQwb4C7rIrnCrkGg2e9VU2YM7B8CennqAe/KU2j6pW
iKH+AsZML+Jgx7G+aLE85bewR3AbeFeI7ZDeihV7MWuJYnCZrSmfACdLprWPJuLt
i12GtjbP6M1qMUYeLJ6UM43jbRz46PVZ4r87Ua19A0VuZB3Mb5p5PcvbEMdC62k/
YibB1m1erw+ametD350NPN5CV1Acn5m8YqHYM7zKnvg6rOEe/R1NFyx+K1/pOYB1
K8BymtmbXt2tHsiD+IojyVgLPqMw0DIz8Ah/58rpeRBvDWLayOy/zrk7K6/3y/7A
4z/hNodWwlhJyxHtAxlPupuOhIl3WuDvgCC9E0vEdAMFo4XDa9BJ3pfGFZ8L3fhK
Ra/nhIvjcHyAJ9+FRRmRTRBkz+I2vkXeVYJFZaHkHGLGoUbXcTTVtItRQBASoMH7
JIg/nU9tfg8qXCqbk3CEMdJ9Kvwu6pNjFfgAAjyL+rkgNQQUED74PQFsigGZFD2/
nrDxprS/fQvTy7gz1hypCGVXHUThlXMI8y25Zn4JGxKJhwAPZKa7GXGjj9iEB2Cj
WJe3UhFcwW36rsALJOKNg5iY4DJMxj79ErVuIQoo5BtHZNYaGJcLoSsyuT7YtMaT
/cqYyD/jtjvuNzcjKQAGExQ8xPfgPxGt8++Xyo98TdObS2/mSBFhDnckQUy+YxCQ
fblirb2JK5fDOeWy+91s3sbXScJ6sdsMvEk88JG4XSpAUBD0lw64Eg3VbzluiVH5
FzV39oHj7ZvDOfbFbLsIJ3iY1HPdJFpLJgjt//Rlx80N8qw7+h47n6eh9Ae6TXTm
RadhC0jDw+Kja75psIl9kda1hCPeOsryWDjoSkBiKuoSJQTVYNQKLFt/Mh2jF214
cWA83plSma13ktHV1igYISeUX8BLvxYetgV3TiS5SzdtYGYpk/xrmPme/kkRn1G5
xxJ1w3EHfzRA4/revT0wusurbcfF285avz/UfHRtxr8yapr8BwCTnniYQK2VZpuj
bGsX7MCqaKPHn1WSdHJ9Cx2hoUJtdwntI/PMmQCPldmRyk9QU2c8+AiQsPbAfumE
ZDvsvaKsEJ2jJMQzV9WdmWp+pnOpIKdYqJ9ZxgQFn1MiiR0CKpovrWv4BnMST9od
RFFIOCj1UnWh14an9JluETtqEpuCbvsRd4d9ybdiCOvgpMbh00pwLPNkLlFxmNEY
eKZ/LTT7rVhhJSej3kMzhRw2WI/M6OA2i2vrV0gyjVV/WeBlkWGyCYCEg6YwmiH0
20dTw2RvoQplyjC63wsrsZZ9jehZtdeaj2a6C44oIHoxodXkfQC1DC4+EjUqhJDP
UV6reKIaepdbjsTOzeWaohaZKLRnJ28woo/P3UGHCzycvly3rCTbIWbwb58YPzOn
j1dA3AkS4lOORHrQYe0Vl5A4jGHwHMtulB12H9kWvonipKxoTfXnhrEj/2BoXtzv
tVI09+s5AfOcf320WHX4hnH45EQ2JHzmna6jWSCWPxgS7nMFeGnF0adAXyE+f/S3
aU5vfSA0fDTwTYgXzMUYS6GcFSr6vvzHUGYtfms0vF4rnIwio+19Unbz9kIpyfBm
Qaa4jxQ3UJIv2vhMGacLiX6f0KMQQzpG/yYWLKSWIoADhh9ijuy7aKT2iuL7H9yU
yGc1MxQtkj4O5R0pqdvNDWx0ExOU183eWjHeOm+BAMIPx5Cqt/uGId/mGo1Ny+ct
lHDoNo/rJfs96lW0oqwmKuGPOPLXBrApHVBcOrgga7F/3/t9p2lODTfS880geFaI
TXzt0e8HxxxMOSSqkOMWJkccjTQEHig5RkozoIChsEmoJO77t9M1OFAK+Q2Ubssm
vkiYrtn2rJqyjm54T1m1OUwcgoWbsyUaO5QJKTLvGxn6Sn36IsSP/J/VqgfCuHlT
XgS6ubudr5VmPegSwYxzZ1560UKJwsxiXI0+O+1kj+pG6fGTSQoo4u2CVqjVVfxv
FgYMVVVX41nhj/HhLpjnleL/6cL0va0FvqmTS2bM8xsnliW7c+WCw0wv61D/1r1B
AQJcBWa011OJ7jv8IzQIl8gCe9u1hh72DM60c0O9JJ/89uSNVNaTNZWWyzte5Yov
/3oW8vZRZkSBQEFeYOVDqjtcglqkd3ZwLKupmP15D5s2r/5B6rUdLz8FkTh4+nO2
jWXhZd3k50iErf+XqSIH3PsYh5592bGhm6FJEiU9mH5ok9bA/EvepDsJN+rSyFKo
V7MBbFIwX3FPvw4v5m4orDvkpIWrSfgXwV9sL9rQQ02KnaWHc/JmZ30XT6U7h9d8
gKjBPaFPf+iIpV8BJoSiW+a4ei6V3T25e4v+D5feowBX4r80uhB9UAB69zMiPAfq
6V+gqHPFgx2bY16NQ11XhrM4XwSFdU4M7I+PVd7IXUndYY9GiBLMIqRYaDoSLxTi
PzkkCJ1ipIVZkOJJoS2XBK4lT0pwnM33iuISN+g4q1yn6UO21WSI1J/HxiiZNb3r
aCSaxjbOvNeH7SalVqKSmnKHK555kdp3f3a5Ax0htp3pZgdCg796skD5yHpC80qa
kIwWuwRz9IZSvGRcifDMnszBETIK4Mko2Q4lWHmPqZaNPBTBDTlgauiTqXJngKSf
CgcdjgA1f9SN/jbgZ2iWU+kbqhI2rGfZnPsA89qGyOC30WEt9ULVx03I7PoXLBSC
gIEa/vSMlItECdi4/WqFU22Ep/e9qZfOrPgIs2BpE/xFGNLyTRXrmXzV/dWonipp
q+sC82adazBx8/JsY43a6gHqpxDaA0mHLS0hBHApzn3M7Qp9LXqpVG8J6x6oAYei
yaz+8wnqQi3/ajStO/q1QZ88vRTDTPL+o8AAybsotM0PNMR8S4gNGJloKYL7Him0
0cemw88KnH6Rm3kzFHZKFmt+450T44wgq18tQ6fY8z3X+0hWwWqCxnujRQU1aUk3
1J/0eV92yd/e+CnIabJLAVSeaPAhczZNJezKrJLxaLr8+8S5IrdVn5D4OOfK/Ft6
+WkKNippqJ7jHjq2N34pTuZH6Tx1310BvmUgXp2fnCrpK3fDBy2w7OvYfAMJtRA7
GU4Lzhj8XNFLdb4UtLeYxoMl7DifWMcsXfKNNQDAFiI80u1MxqTu5cQEce+SqnWR
NAh5+bYZN1XWhtcUQHaSpVemSE9aE43Ldld1A764p5/7AwO94Z7hz+ZqKkL/54zE
k3hazb5naj2g2XORxUpV+GlKjvr70ah5F2oPhUNTeEQHk4oc16NC627EWbbKPEQ+
bogshnDyAH6lUD3TcnD4YPqCa2fm93PwFq/xLqVWPaLEUOG3NJMuQvSGTcNbuoTC
skOzQMNV4CeOJTPoXt4qHpoZ1jhdgU6IbYOz8PRN4Tql35+H99ygZH6Rt/XDjY7J
bgLTggFshsP9qcAWwWd8r0JeMkmfbik1cLzZghaMiPVj1MydVAaw3EbUNildwWKw
HDS8zy4MIBobm7uSti7YUUP8XFuOpm+ssJJeLg6AVm+b8/7bvNNNYCnSAybRLLA/
VQPY/pqAyC94QvpyzIpPh5fCfI2IMGKn9mvyMOLth0UvZ/w7iWY6DBIpQNflh7jY
RkizeHuS52yjAhXjtQVWT0vKGAaJJE6hBNBK/GLZV7dR2goI0RguCGrdkUAxVxVP
C1Xqbz7DWqBuG9ECgEQhnQReXBvMnL04oGD46cVw5dOBI4Ir0kD0J8RoioM8EwUx
t7266w+QAdoRSRzU3ObfxuDCdfnKidtfuGqcE24Z6FMUMN0CUjckfHnlraqN/bw8
JiAbUB20ONKT5CIuQs7krlGVZy5MwAkYWLbyx52NDx5RBUjEZOOGOEb/Q4drIeJL
DnIjmjFgAarZ5x3T1DBvgfG6xb8NduXGVdvTLEdvEa/NfQBWPhpp12yUm0sFR9vT
wnQOdzC81mbSqG329hQ96wGmrIDygfJN6R/EU5QDnmq4ptOlhuLpWTUGZJyUsMTk
Tg2Tkvkde9qBw1sv4MXxHZSeGb4tqR4WKEz/JIz6xtR3OhAWK0SAVnTCA1Ir4daq
bfbF3nYyc8ZWW0/O63AxZ0KX4tBi3l8RZmHd5zZ4mvm3yhR1krBfEast2rtHfBKc
2695bgkF7eKyXHxvlC8nJ4j2zdoqUqctuXnuMHNiKhS6XMOSeZRRhxhWZEaU8snF
Nx/94PYe0bEdnYqPbCxcSUMwqwb23Lv+0vpF07TqhTUclNTjlM6jq0SwH3JNYs9Z
5d+pJjs8j6j2MzRGt1xU7Iuh2mpg5LDBmiycdoRBCtkl+ENVix/W0BDYAxcxnZIR
/cQ0sEXsDKVLUaxdj20pqKlS4Lv4anEd++uaiIW48apRFAIfat/WIe9ZLcYG4IvQ
j62gX79fsw4UE5wmnIzTBdBWnBfVORvcu0l6ipbz6npEIzy0cY0SJnG/bxpXWiE4
hs8nt+I/9QK33nZU6GbLd/xCLudVg8XBIkK14lHtCig+cYES71Fr1pxNwigmG+nk
PhE7Kk/kvDhm15JvU256bxSZjf2cxK7BXuFTDM1D8f1LbZ1OumUnnx5PqJDjuG3t
p4kP35a3Yne03AtG/KT+aoljVNVXb2KNvIuF3nMiNL6ROIMOfVn92HUPDbkCR1ZH
eYIvKZNBACNzRxwBWCESk2PaD7kx3jEo2fwoiYRakeIZhDARZM0T6V9cf4eaOxxl
Z2NwF1Czb9Mhn+Xd1x3wlsxHU+bGwvvD0POInEGs9JlSqomYJcRcxv5nUWAE0vp3
JvPIHdH3fc6E/7ChQwEJdRFnlb2ktYTSIcHNQ+Y1JSJ711sxydMCpZkckfv3SKiR
iT+1mk99J9/tqhxbfQDJYVcl0bHEZ386FR4AiZwS54bg60k2KnRZ2a+w8BPIm1Rd
8sXN46MI/mh3aJjO53Hvfbqw8A4CbLHjy5x61vmiXOk3XY9zA2bSS1aE9oma9CA7
YSFkVzYqkbEZZsgHK1Ma4LETX9lvMwCPOx+dZvCiGPb9lalif8lBNqlGZsDaAoRp
wcQ8Q0vEZnofqTWTB+JNbYYAj9QD1DJ8yLmjlQXvGh4lT+VkQ/ZkB8dxtSCtt5i1
cZW8tC4Z9ny1eHu7knkncnhM3bXt2EFX1DnOPd6iQqr/DFGuhEFln+wjhzzCUPUe
NEJJqdWTZsGNlXaLVjWca/FfQyWxuECi4SY2FdKJj4+yGA9d3ArVZYa9RBI5VNCp
oUwQQ8H7V9CadxKMduC18jFifwWQdBBYk5QtT648YOl5Cz849o/bB8xUCjlhE8D3
MyvEgUzLj+nqZQ7OFC/Bt9kR2Aosj8okLPIxwPIuM1ZBTpfA5JdOU+FmhdK+MKlh
UFweGQDO/WHYBcBd0cwioBtIxd/yDpeWV/PELmiP2lQ/cj939WctmGOzK9zC5mlm
ni8Dg+Nd5jhB7jLobh/TgyaadPKsiskgK10s3dh0nZdvHgbZuq0xkf1Y03Q1KFvL
8Wk4vTHQm5LYqHy7jvEezxjPWmUI+mb+uyH7L/a5i1EOcWW3QrerWQoMmct80Lqp
utXZmEpCFZQ/+w4BiTM0tjuEvI5JJSWMzKmbsWIClgpxDCr8zc68KpqAQ/f3VtGT
Vxps8qXs0AJWusWA5ESXI4auovqQKkzzEU3DFpGnLNd9TNWEixe4zv73JCfE3hpZ
OHMxXi/AFrf6iDUkfj2GNhVWhmjl9YsJse3SCDuKjY5roB+IkvHVavcfLRS5Jsi1
vjYH/+lvWdCYsFOHobe3sBoYzTburUaW8tq+KU0G5E8rZNXKDMj77Roab+guHVPN
HCKoKNjSuQJtQBCUXJ9RzSlv4nm62wSGVtDoJlaIG1OpGmZ+TvK/R+YqxnFgGLnn
btVjJMtkuQwpuYJB0Y21P32uqXUX1H4X9kK4lurVV3ghrzmTkQDm4bH6fZzgC7+A
Z3Mcv2AQZUQmPXX/HX3hTfxr2JCIhdR1XiIxF1aKEF2mH6Nfn4aKeOYqgXvAVC/i
94vStv6eAuk7Fk0UdnmBrn7N6vOfmwH+jQ4WZAnnAjjADdXTiYULbGdvRY2AZkhe
TRkve0KHvPy1UKBa+FBm/OjZsyD1LJzE0wStkgJmIMhNTg29GlZq1geNeL2zO4pp
FjK3rxxacaAs+ERoyt5PzplzAm3sUX1QHOhokoEnH0tfFYT/q7BgcHOfsEHh1xSS
4cCbdeTjSC+HoHLhAZTIHMU0Zr72GOc44PQXbc67YBQdyb97c2lXSqSEppcP72XX
KdSRZcoTbMJYf6877tpqolcizZ/e6xQWe9fQoy7ckBG/fVspwxv8W/ZXquj1XK0u
xgWKbcWTMGIMj9uNo5WMWnUvscf2Ih1HSWBTfJtPkcsWZR91iUde2GpbusiDM2g4
dqQW4PBZ9Z09G3+jjV0ZABs3npW1l+yC6SoMWtj8PG8/ruceNLyv2Nt4HnEm+C40
lxxVQvNlsbuSJ2y58+xguJZ5tvz9tywDQAxaEHTj5G2AipDYH3/uzTAKwQ3vzvKk
yCUV8NxmMTSkf5jBAlNZqFIAAmjObfQp+kA2IJ5eQg0fJlSRpO+Gqg9wpN2upFwd
0Wy/sIZ5U7ZpVilWDNjep2bDUibVeaTysBX28sJg76FPtDaw+hn/JlguW4ppK8OF
AxsOdOLqNtRU3oul7q09D5rNLz3eN48JiXv670UMdrWjwz98YXW+y5yCQpBZ3OQU
jtBHd8aVKzkyWRpVXpLs4DNqTiGmtzMHyBIFKsj7NsbzcCB2zYCqKGD4EBcc+p/W
FuKTqrqYGF83fh5a0JrW/TTzTfXbUeRNdJHlEvVG+Bw2HQmNUwBL2h+9rg8c+JB3
uwa8cplh+D6I+prQSvKmYDtmm0dfMLbCTdHWxU5QDMGjYXEptIR9oVgbah2IuFjb
fKKoe0MwbQtX8ZpGd8/4U0u66RmUmCRg703ENxQbmxgKXFRQSdAxS5mYxufac+AE
TwCBUy9ivq45HVcHHuhH/Bynic7kyEZCkDhh+wXOCw8+4Nq//fMAQF5x4kwA5XKH
mw6+EaQy0CjKhVZUmdfaA6/XXfOrBCZhmRqSMLz4d+MXCCDIahf0ClyZR+hMvJEd
p3meBmrpGj2fKYU63QCfnZP3Zhn0afjbiK74yEQBfR5pAiMwmKpnniFj5/3EO3QL
HKdUSEnQZRluZR+cXg9ro9QP4TfIprYgkjqWzTVdj0IWKedQQLgWTmyT9HOUTp8F
lctD0jGw5M/6ovOlu7NYVnWxVq5BmTKP494v3PGBy4+Fzq0IEsI3uap8rC3hY0jC
YLxjLxS+kO2IHJaMSfQ9KSI/jIiXxx44wKZ3pEfrNM3SsLt1eWgDkgXXhQqL/ILn
FqKQIB9DnGbnbcMlPx/4dXyk+NMY9IvRbN2qW+B1kqJTMMwBloo9vGWMVll5+rCV
B1dIOnqClw/k7v8bLBol8Viqv6hH6BvKrBUdTEKK3yXfQ4hN4BdQnzjR1hpFzOtx
X8JC+0B2cSTmx3BH2Aa31GbCXRM6IDf4seui0wAqbCySEJvZKQmjV1YiI22tbS2y
vF6aS1p4+294taGvhRChCgNTOWoqiNlQ65/tyObg3RHZ7xoIkU40fi1XeXiwyVkU
QdY36ml+zLtLIgAtl+gb3gyuxCKZ9CLCBpqNacUneFtH0tMTa0nIY7hkszWwe65b
GK/iXGUDuYbR9gJFuWLNY/zCUnrI+7BIriAomZA86jTkWx0HB3HXiLfsj9IGGbo5
tEety8QGrO9eB8UluvwXOvET5VD2aWUSoCCSz0NNfPRZ5qZPTJmh0STQjfIUFfqW
MTcPNaSapBOBjAnfjt5Hjmg2WzD1CWLaKP3wLOXU7a7TzJHLNVZNU/moePniDl4/
khXgSViJ32atjnNS6vTRmVT/20PnQwOIZMuV1W2/Sdsjorig6UDwoL8hSQ9ThI7G
aJhEFpAkGSjqRn+yHhXWpzSP3bZjA1OSLPkyqIBBNafdYwR70ypS2faT6AUwJ8uG
Md+qYqFabr/hX57qhtr4m5QHtbvgwuuOiY7hr9JtH9E3QqXNqohc9RQLJKk76LEh
cJfUL52H1HJVJN01u2EDYqQsFfLWgf2WA6w+L9xBAAE55SuRHDBxpkrbDWz0Jom8
+WtXHFkGSlQQd9iyvkJexUHW5G3ybzg6BliBK00bDzyLXTMHeiKFNiYQybUlxCTm
FYMH2JL6yl3OSGLXdXlm0dYfMY2Zv6SXfTwZ5zA/x9xwwvwBTpfH8oNFkqA9rAOY
hk6E4LpZZV5EmA7prXDQpoIEdbvtQjB0plZ5kNEabFSmMaqOGyAP2furcEtGW8/2
tEK8b0RAyQMrrSnkPSCgL7aEJq6fo/Grmne9tiThwqvVaoSYTcig/1mck5pmgGOq
AakrJfbZfub/J4drCjyUHrTUM3knmlOHWTW9AS/4a1VVzB2Htf3/jy70z6imPvDo
up6mWzwxwl3620DZFU/vi6vDy3mvMJAtpkadYhjlb6NXv85QwPb4i19Qsbu3Fybr
Hyt/yXGjsWGTFCsE/CcCrxSZYMF5IjYdt7WW4wMM1XVWh9jQZZlQ4fk/Y2u1cQQs
9nwsNhUH2IIIb+bKdBFw43BBSxUZSAsGnyeS1sH6TJGrETIuogHHpFzzfXaOsKDJ
iw9qaDg53WNU6GmYcbwFVx6B8OyxcrkWrK/Swl6P1B4bIQpfcFMKUKhMvg6l5PoV
ul75mxKxmCsmlXZVAfHzQ9ggheI1kUrS3MWbMzB04lu+Ife5qh0LS1M3Cw6Nf5Zf
UzbQg6V27VYLNh+eACaDH8G4m2eyw5RPAs9dy8NUnVuoU3fazz67irUZbqLiuWAv
2r+NSKcRigl4s/PmZSuDiClh0eCgSg7NFYBRO4fW5ArT8Bxfg8+wht9t/aR67T1B
lm2cUTcS2OZnlhZ5rSgBNemJbjbY77o1oSLB9pjAzr/A1msaj2CjwjTZKaLq9H/A
EA8+4iLO80yEjRfdSgRW7TcfOdHL9+QGn8Wx5mDPauJe/bgMAljiQGDfTniB+75W
9FSn5sg+IPoVq9CpaM9NUIP8xiVgCVtnztnSUtkLHURNi9Itp7+6D0o77wpdnjEf
H/GjmFkmeMfV5FKEneSXLYQrSsIZsZGbZIp1d+LXX6jbvKUdBYypComhLM8lW+5/
pj99gNvpHSAsCQtGeXwYJK/M97Aifu7bwHc7BJ5qi8BL2H/WHIsbR4GZPdMUJ7WK
vsue8gJks3mWu2kLxK82jBU38k3lujEl44SlOHnT1klBhZpItfQhW2KbZUIRCauA
+Vp0g6SASXUbVSpMC+vXBX9NRADsFf1lkdOWBOC5O4zoHBUwQ7avBQsm+lNo2bu/
tnYAjrYRmPBnfsaLQn+wXzKD3FwD68PW38MoSqL2+cnWO0tv/brJSFGnU4YrQzY2
93EqQehYMY4SM3j5gqeU80mCdlsAd1iS2x+6bpbTcJ/6rB4rH4N30b1O471lqC4D
yqCFfguFOC6VsI68lbH3/tjdAIWHDnnj92N3L2ac+C54WpMgoJen4fALoVySETiT
+rIb4ec9UXW4+kH2Eb837EW3WPru33Lg704f/qZA9kHUL3bEFqYtk67Ba5XrBxJa
SAO7xp+B0Mjegjd2plUwzn7lDdpq374kuRtVQztbovMbNgNka53VSSmJoyvudwoS
ayGaTrFpwkO2GK3Hk+JT2iNAUQpsOFh/09cc71KuBSEH9uinSUlohbVOgKc5KYwM
UhAAGHOy9tuZJoTWcAsjJj08sguq9xadPH3nqe2muP0g5dP3vuzHUgQdb8KYHm/U
+5pJ267GnfJfkMBThzU99sIP3D33l4ytk8y7307hZkCU2l9N5Bh92Z+XyeIX+K9l
qLk7VylfvCQGl3++3V75phy3LNVrbMyl3Q1SBaAeXiCcw5H5dJtgiF7sw1EiDQvH
ykdnFzn+nZ9lGfjaVq/W3LU/csm+prndTmbAlUs3fYpiBaK5/dcJ1Th85ITINIFJ
ICca8IyHwB6h4c5Yjcc7O5Wt+8G3FruPB2w+jM7LrQPKx7C69Kp5Kn97myLcTDG8
GNu+YB6vSAipTOmjZjzBKEyNn5+gbTl2bsHb4IlPT62qcfa6lgLqTIB523arnE4+
s9QAEYW862FPGt+PgjPBdAITDkShhJK9FYihwOJMhEGWo389irPyHTu7Byj5pDPe
f5Amr+sr6xnWp6LRbAxDhXh+vSaHlOXvxJGmkTovkRLmAzWuOTMGszTT0vElNVPR
n+cTUfusjkqwRb3Dxan+PHZ0Q+Im8Y9tD8Fi1iBQxy+EsUY5ONWONZl71c1Mx8d+
pUAoahMYRVsIVDU1EfwobqmwQ+Te7WDkRYQMH0g/wbUpZ9V4uXu24y+2ww6Hgz78
cYmlroxA5FcHCVNpwe5pOQVDBTeem/sNX4OwC88/3VsX9CLflHZ03BDbc0DGp3Rv
uIFloBxcttBDUuJh5PcKweb1+iekTUJKvVdvph6TsXMXV0OILROaI54DjrBapAZF
7Il9XOreVw7c0voW2ug+FGNDLvOCdu7UsIfQ9ZCEY45b+ULB+hCbupqnR1bD3dha
Wxn6ndvtJY5WQREUbUPXhfWXeei2Jx+wS/LF0s7+eoiNn3E3l9FzGbH5U5gdpswP
fAvtViueqemgxKWIf7p1BDMyzRkYSW7yjAbnXylZQq4F9HasgLon2ucBku7WFIoq
rB76dVBa0nkkQsNB/Sfq7/BohJ2eUJN9xkOZKR/jZeQb9t2WHILjXBPVojYwNR90
RGAhuf94hsmNhqKYFhL6m6NPShlC7BsmVhMT+VmZ0XG8SRbP3zD3hDHH1ZTtDVam
3TO46M5hhjtfdatNeARUoQxcLYH9mpCPGyfkC7Rac+Bjto7SSuDAo/iPb/PeVW7x
UuWxEYKnMljmCUPtoNVvjqrxy+SRwer8T12RebqaHMkrVUrryIEose+BY7XIrGQd
CdaZJqB4bHmfLZYVxYQO9DFeq2K2FzFqiHgaf4baMJ698byRVPUbtQp7mP5p3gum
4xZ18optWeDjXRM2Ij2WEATfpWpXtR9G7Sn/KRrG1gb+YiVhTpf2kpcpNhKpgGc1
9LzzJGW8kFvA8zyWffwe0L0BZ3nq+VG6CrJOuBD6tuJ5YUxaVlcuKSw45Jmn+2KA
7mGLq7BevvgmKQ6V/T7NPx0aEKBAlzyN6XfUgOJNDB1pxNkn370dpjVfEHFjQRg2
k8glw7RAV2dSnZlJtEr329PAIthDw0BD5vFGvkxMiQpMV+yvCl1bjEhkzWwJ/q1+
65gHM0NM35FNREY/VWM0RucN3eklCIK+Vi+9Wx9kRiM1595/IyigueLz2N75dIhB
LZywjfThusx3hiTErlyUTopqjAf4FjKJ2o5Ff1kzxSqtmjyS0z5WG1fashhCoU1D
62VR24e8ws75o+msZj22qg+YehF1N47oVprdIA/JZFchn5F9ggnTwHAubRrPTlmh
86lBz68EwfQB3rXlQIF6RH1PGap87oYBYAnpmxY7acQ+/fYCm9K1tOEE+cRFji6A
BKfRl9fam+u9rdCoKmiMDcFQdtahlcAXr551yzD5n09UQJSO0sKqwXZcC9cE5JaG
8Y3UG9mov6qRlgP5geOkK1/ECCvJ01Ga1s1vcghMecv3ktXbtY4FlBC5or+6u4R3
/4Ru7L9/5Ogx0nLTHwXZojk4LQRhR9dAe3GkBQIbnMt7UpU1v+I9DEzIE1Cb28xg
6Pwrvc1hUQBrJnZ0/uWCjbLAWwdjh7OSBxCaD6ZlPzASyT/efwmMQ82dWhoxnhG+
XyqXGm89nb31mXiIuKaeQIsvxIuMf5AD374wBJ0xI5KJSOW97pZnVUrG0TiaEO9l
CDbgYUQ8pvEbh+YNFI1OloKmnLuy+rD4rejW2khFMGX5VWnufPAu8FbpzKJfIl0c
JcsWDqyCSzsWMOsHCKcnLE96hrX7rfb5JoNZYPBzmhM5ZMRltx7X+KPz7U2IAtod
y52XHjLpHHtuLYAVh1RsLRmnI+2dy4vMxDxdJR5bbmCEtq7PgcRiR0mj0l3WHY17
hZ+sEukK2hddL1XCxjbtJA+DI1S/R0EtRfkqpj02knBlaF42I8wYbSzLrTRGL+cM
3+HdWu6KD12F9i5jO0dXLBrD7awsco6tRfA3J6U/JF2nsAz6Fm/LdZcvHUYYuN+J
ZBBkSkm529uFqNEKPZlYA7eelDCnSltT/erQ8CtwKYTbVlFE58CJJPUJqwybiyrv
rkJ5DEG3TD+9Ioz0EJv1chRv1L7+c+iRslHz+UzYeEi40JKQZ5zTDhgxdmgllrA2
dKfffsM4cKzLx9kEdhL86OvgX58+BP6gYR5YAb7WGCR+7OsIm50bPIrKSrVs2bgl
9UC8R/COwHM/3IyX2IUCG8TBmT2cA3CNPsloUuMPISebun4PBy3rca/H6JJ89s2q
SHyonpvLovP1+9Zp/HwYK1EynebxxZbXy4+Z6fuiKmnK6tE1HCaZY3yjO10wXo68
/5OIQo7EbNr80ZTnkdNUMSuC1dExCUFOfTO2ibt0+oobFDYHyuPhsCjF7lBg9TrH
B1C+7bsyLKkwQG704C5lpQawYz2oWYn2S8Ln94bI9/fGMik+G5BqNMdogORSTnuf
ZGJX0WPVuCClmU1MDJxSm8RQkwcJhnr/FY1g++BN/8ZRg+8YpXg5xsTGf3178Na8
amqpOEzTnarwwTN1q3YbXiJyXgRU10R0Rcm4+4Ek67a7blUy+hMDnX8KT2UGQITl
mIpacCAEaOLY2w8rkh9eSG/eLV3+QN+ueeo+s+s9n5KGg3UIPuD0Xy/uqc57XgMW
9SSP8p4jCOrT9ABlyLKy33gkM+AVdvAvMj4FeVmJbNJkmxsrtsuZZyYw/kXb8ybW
AU607DYNijKLO7KqgzpMnUzxalyAOYXxohTHFfAtyqJVGxhoFLJCL/fAREtqniHX
WQkS1RR20IbdIjZzA+kjgk2kwZEJ5z7lylJKPELnUN0SibhiFohMEDup3iQIHr5+
SXpMvEL/J3fwPgKr4Ojku6lOMKB10vD9ghI/TxGBWSt15Jsn1jF9fLpkVVusb5JX
TPLuJ4B8Db9kmjSjZF3ln1NHgoK6ZxgtpcEfslZvl51fywzf04owfYLSd6XQLJoW
QVC3sTkBOv61I2zIrGDJgeFk2hbvz/cq3F6TOj6L5Dl9/m8cc+G8eu1ty7JY1ZG9
BPiCmnJagSXQsjYaZ4EV+dc0B9ogT/fkBcMu+Y01tTE7PCj1ANIC0Oai6PZKmX+h
VzNqZVCtyrbc32RvSRxbyslfSv1mqf012QZUNqHZPXofWvu5PUO7u/liSVRbpw4q
t6JipcyL6GQBdQ2wLEBiR3XNQYboYVlBXO7GLNj0yHQNmjCV1u6lwVNw2R8HdztG
U4GwC+EcSoRtBt1omqjwTRxTJpaJIeUOSTnigd3LrGpeIMw+ocxXD6ZRhYnyuX2K
wezacbA0S+qKtU/sCogtcmYpjo4RG6KhV4VIEjFr6zFFVirz6D6auhy7h/YNMNTz
ImmGE7JjNp0hgarihBbcy3HyEUqUE840N9xY80EACDqFr44MUhW+EWCNP3DH5/oJ
JLr8ZuxhG4c7dE9wUcB3MttfLUne1oBLl2IStr57Wl5zM1A/h4qTotXpyy4SHKgE
nV58M0eTGQSfqixbz9spEJaJGe16mC03mS22jPIfnIh70rBjdjpE04QYKL19ktYY
T7Tl52jgiVAPo5NJNQYHtXW/L0vIjF9YRv1eKoagvDe53Zs0ZMCROBoDkVQVgf4N
cPmo9HA6dUnRBdKZfsp5BA8KjFz47uI8CyK0WGJWCZKrP4iFqaxUQISzg6sEqzSd
rTqj5mB1DXOGCrtHJMiykcf0ryw+0KW0xvy2h+c6IdRjP7xKRFnL1899g1xokfMb
P9wR93czBX7zt4LYK8XvnWsyUg0m1qKEQteg0G4sBo0jvwLWWnJ3AeOTyTVvmxv/
1LmHk3PV8Da/IBe1A4x6ew0vWOW3knHNbtJYMKFiG+zqYq+hwAGk5uu7Wb8WlCOg
dpyjeY+OCLhC/+z4qLusupcTrle/0M4AxZ4ru5TnVS3CfJ4hQ1+XS5HqcAmROFTT
gXZqTMCkXKyyd4z4L4YG4y5vJjbk0J+WpaV1X23YbXee+QSMbjOCbTHxGe/oQTmU
m1BkYBidkeRrsgsodJ/fCeNKmTzv1XCigVpl0N6SgVrbL6VBm+Q5s+vqpeJ9uUeO
s4/fFIKq77aXcgtiqJ0HuSGpUcQZ5aQou1dl+XsgRsv1KeGiD2Qlnp5wGGElTxNn
qDBmVjidUzfectkGxUr01Yg1bgf/pHQayTCdiP9+5BEYlyBW76s8B0cVhyhKFsYe
NNXoYkz16ruCHY2pTX8tBExOYb7RuyZBJFDMyZiZjG8boFX0fNBrzXoVJPZV8neT
swj+T2JYuptD8/cFegpT2dCgxbaH4d1/IXA9gkCr54aE3LbTIbaxN8k6Nbt3cJpH
7QAXh38kBh1O38fLbwVI7AyruDYEOZB3QCUI/3PmEKDYTp8HGdnyFFCSRuOs4ErJ
8itkEjXmD08PH+xzP3G6+Ghs+jm9BeURqa1NNocMt6tJRwnfw2yJoMpPs8Jwd5Gv
mV9THiWDTgwMRnU0I1N6U6uYv26LJQEWzImD5At0bgyS73y7BTZ80h4aye3Dq6Xl
+Zh3401MQQsl4tBOHxQ5l7ZKzcQAfM2aWiXWn0M2QeOjI2BikquE1a7Ht3/l0IvF
/YhdWTNw+7jgjQT8Z4La7jkkioND546/D2ssbSh7LllnIMwIp8l3U6kFbfBKHP8q
OGKmcT9eiVaKij3SHnjjSlMXriZhgVwFMOhSTzfvHsYw3lqfFYYjDukG/vFmPJCR
lVe2vWqabqDTKEThOiAf20CXBqEEJ6a0NkR2yVKP5vY3e9LNcpuGPpHlTT/kw4Hr
Uf1N435sGZ1aOya1Z8Knv//TMsGcerENeNhE/gaokFUV/CekehpFZGN3YCpieMYM
l8pUHeEK+cRySfmMSD6sQAod0GL/of6ZuPtVSD4mf0WOJavqMleRL0LlupqNOOf4
XpJpkr2xWAQE1gdNA18HhjEOexgCDtCGsldnoA9mpfuKr65N7w4zT/qp7kXiTcjS
MiEi/B0EFCWiXTDK63FBPPNMbsoIOmfNBiE74IuSkcCftYefcrOuRGHrCVEuhv/6
6VWGyPQxc83CTYcSqnjr1X6e1KX3tDURSqIGhWjyy3+axi0gdYrQaUYdYmybbiKD
2SMUft80ECByZJZNQTPNAufrWM9uT2hXZXPhCr8ynmh5/caBTF0ZgQtFsnlWwcQw
3tdSRHFdhYQKDYAm7Fd0/ld2k5EvaURatdo2hCelFZNFcHPJngyPJnnKDLpw+8RX
INs1zYcgsXzziXO9ohjRAuRvY1HYVCBy1yuDifQpFaMHQPVYwMrYa5CoyCUQJZUg
oartsioASH3nBafuhVxX1G1ncEGX7igCOa9vCbCtPu6FHhPTXixIeR9L6+SB+foM
dbk4K5WfUxOdFopdFIEl87BTOBiw/ltCsVdAYkTkarp0x3GKh4M3CJBw1acyz04k
HWLgV0g7uGqteoNXZvoa4iUklmwwguC3+EMz7v6A35/QmSvFgf3Ui6B5s6VgJtZu
JsDotJFBrNfPgG+1fHSABz6i1u4nAuMIhMVVDCZ7c10olHAbC60F0betQu+uEtHF
1t61gyVKuJ/l06gQir+hzIbtLTrOzGVMn4kBNDT1QAFdj3Tp11jNbuts6QP4dcoL
Mdlyqz3u8YuZcf0dI1FuQBAr01P4Ppl3OsHYrjubb1xoA2hBffBRGYdPEKsplhfP
jGGSnMmpRJr4Wl1Va1U306L4NT1OsEYam+9BIw8LJj5H0/ddE2PBsmfj7QsSzmEK
Md95S3mDLKB4nxmMJoFOJlUxbmyF8UtEpv1Hl8OD/8YtGH9h7XnhFtJB4mYGDRWo
3ciKLe2BaAp9LXKg1pPETgy9Qemle3UBQZbqHj5i8Tj7a+qsVzVjGNvwNvApTMX0
piG4DuAom64vr2I0PRHOgVxlAYP7Njbd4QL4gZl+RSDuQzSWyEBImB7AHNaGKys9
moW4PzOggGV3+VJWRj4n/ql8H5WptWM09QnsmhqXK0C3EhReR1L1H6VHJasKDs+T
rX2wgi04TCeMWFHKmnSK/DwaM12lcrImh+GNdD1IRv+1fiJkaE4zZAsfFo5LtdVd
tq6/w6oWyJG78NIcuFuIBgfh5Vwl6XRDKT6PTK+gwhAaum48L+tuIvcwCAO6M/aC
rQHrU3NgSNog5RQHJ2useQ0o4NwhzR6VPQodZnnuzmaNQAc/IqJy8MEE2UOmI9FF
65KMaeqhdWDMczYp11bkSY7g1BFKDi2J+OHFIiyzGqOJZVIIV3emEZsorEUK9U3G
OwtdP542Cj98lodQz3dVoA7wn1bT4dq8WE7fOz0j3ALkoecTTwgrujakdKiluSaF
z1hR81I4RubCHB4W4BV9AgjvNsGfH+W2q2R9qfhMaGx6SoeObhSWCzpO8A9HrTsX
vcE2+CnUbhmGrYW70D6bc87GYY+WtU2d1ZCXLmPMy310aUsALQqsVyyfSGobBAWo
PIBht6ZX0qbh+c3YJ0NbBLrIMFMt8HuyssGhwig6++YUWVyM7KnAwSX0WbmN4cpr
7mdCxUEKvJvs9CzPJgX0kGMb+Q45hO01duxCdtyJMRb63BjWGnjHGQJvwN0byEkg
0/VidTI7ZD6sQlSLGoL0iBN9RV1PJgO+0jJO+5wG5Yj3isC8td/Wvy+HQrUo86dv
RlWyozp93bj96G1jkWu4SJC93SsORWuDk42W2o7iwrYP8AFz+LuAlm/6iBVMbQT6
Tk8OA33fGnqo8w4a6oiE1WbgD5ciE04uchj9mnMrDLwKiBi8BlPHleFHXW16MAaX
zU2PjbSPbDE+GaDCXyOjacDAFQBX8NeFYzUUowhHMsNAGrUCZQV8M7iaYVBlv/nt
mb+57QFijPYdkkHqSyutWu/YoSlKC9d+oJhpa7izrfc2jtf+9KYT8W1+pdB+wtJB
AGwKrofqTtnack70FudaWncUaB6TU81JzXzmFaiQQTNvn8lxbMOccmhKNXrcxETd
JWti/HCTOMa0yvgArYHajZGEj+kb1jIYQt+tqDM59coD/tfdqkn8z7pkPLIskEoi
QcKMVTrxUUff2Er3DDds1Zx6j07cg5TVoSxOd6orQ8pR9ivrU0SQReDA7r2OFaIN
FJ67ogZKJ716s38ZgZqCZmgOon7h+V5teBmgMQrCIsJ+TfnlH+DuVF5CWrGmqTms
S65vOtQKfWdrZps5BaCRLhDU4RMcitcFEAfJlgo8m96WYBbXU+k7dkMfbrmHyJ7G
NIB/TG/plABWrUYSK5xp3rI2rF1JGRYnptBDDL2te+OtBB+hoHoHBBQSRxxMFgzK
VFsbG9M/qSb04sx7o+Ph/uuZXERPAaemGXv7vJiNFbhf/np5/BfGDuAo4lO4Iu1b
oVUGtkUlsyb9A1DKsRRaXEc2eEoicWr4HP+m+TSuMqDNnpv2QDYZOCXtbLvLC/oA
CIZHERoCwBKavSL8iLjZsGLJExsW+dymPYVG5XQ15tvCJmxfqDPzqILf8oDysbUN
zOaoqSpLqe0888448hs2EozYVrjn4oZ0vQ0kvM4NM9cL1FldsPlgdWk+tD19WDqP
dmP1mwXynRffxVypOxuAVI48e73kqY1utyHyx9Gmof8XsR09Go3/6r1UXhi3kS0j
ZRL9fQjbhbHsqXxqWcXv7nue6tLVgxngZrECwuPMgKAUCi3QSvyafpMFd48GBDg7
opISrSWHSp0CtRkXY6uMPFTBWfq/5sqU6Oc/bUQ/ONTYjHO7b+VyPu/VAh/oTB5p
x/hDcZddYwmrwq63fTPVCdTXExZcKxj3Eh+J2qTwFMh68+bNUKjMsdpNp/wAPrJC
HRY+yvhyvPSOB9Ok+1KSN9UQqPb1v7F7VFChM+8Od+Lv5QKD79nDAqhx63IXW16u
U+ARE0tIaHtuZiJnjmo7w/zXZBYJQQ7g4qi51nEDB8eBTiy2BLWAawNFqJ+vjl9w
JtzkVWX0GoShnZuM8bRVb+LPw8XuLkbsSopzu4B/MAGoY06Ork9cuwj43P0wWdma
EYOnzvKI8B/+9JJPaq0wuEXOw1K+ndu/Wv2pQAh4ZycnC8j0C26mzmXEd8ldrYqj
OA2nJwRdL5mTrwijMlqmPOqrtYH0fHmWSm35utcpNssLPPbwP32Cn2Fq7sxcHZQW
k1eobMrKvULlkGgCcaeu7RMSr+Au37kWVCDIVNU8xjRdgBdXoexO37NvARFlA5ZO
VgoHfooa8vCCX1s0E+T0EnQf1hkM0EvaUTaxujRY0Q2JSTVq7zIsrRvjnVwskh+K
wvv7dXKkLXUr2uporxt17/ViXxbHnquNyLchb7TXJF+ncux+Rrrm48jtt69Y4cSe
XamLU2hUzsd5KXc+KnzUPVamjRwBZn822NE1WhMkd3V2kYs6YxZXK5hG4++eOqO8
c0Km2DhedQ9ZsKICUON2xrzLzpYLUwoTy3B94zbJR0W8KfMkQHnXefuS7BHZYMy1
Ri/3d1qWQB3XF2pT3aDDnxd1mIDfk/DsX7DWrWNghD3pBdYWYiFNvTPndwiWEPbO
cWUzWAIvpHr/G3W69pPfn1SMWWy01vANN4+2d03/hmdFeP1feseM9e6L+hAjYqc2
rEkmFHw1ivSgM/N+4kbghrr7PJoYYcCT2MxHI5QvlJpeEHAsm37KTdyJ7GCl/LB2
imWklKiG7lpLyGM84R8Jp6WVzob8BRgws0slku6CxluSDFAXKJ6d2f6Q3GErM+1p
sBGVkcPJJRTjcdDRMeyTJNi3K3fDCBJqGw3e1IThbk4O38pU7qmqYjF1rne6koqF
iUU5Zh1kTCveT20rIOI+OAHkh6MTUQXXD8w4vd9VnsghIeH62ii+0S85OS5Rmb/F
zJTaD6EkOrJBuF9Vgm6zW9EdKBJcjIhX2LAku3RmFHX4uR/AUbt5wijo4D55B4qX
pprNFTJaHHERkyV2Jze5Y/nsKhSacVTS/Oz2qMDElPcZy7j15TT+XEfF6OpfsgEH
vhdlOMQPuZ4+AobqfjoasEa9TAcUpTGnv4FMnEPX6f8t2r0b7LHib3IXDusfKjVJ
NCn7Yos9ClKPe8ZTG08f5mZubJr5XKfuX/JoCx62Pfx/NKIqV0ATarhcZ40D/07m
E7QlGDP7hV5TqEvryTDt0tccQ5LZBAI6zg6bW//1pfLHwxvQK84FJAlOjyi6CJYX
qwGcdTS77fIjFOEY8NBT+mm078Akg/N6LzZrbGjIzvs4vIK5lr90Ek+Gme7LG3Zy
5yrvQS3mnW9L31uFUhKmKQGMz7AxYPAY/Apppqb/YAtK62VO1PZE1SocWgSfQiaz
wwllHciqthyEBW73YEgC7qNp6wKlRfticGPtUA7RGffS+IgvYYiFSnufO8JGnoPK
9LhWHT3RRf1kVazkD57v5bBkpHzHAuSNoTgs2eqZRu28JFxhwEiNOfURNDv6UqnC
gP2YOa1jtWrO7a/8kwmzPn0vJIa/ib+s5fEgEH4Mo9OwK/pW90IAU3CVG8HRDA50
aAOfR9j1CADqYYoDj33jaciS4e+pVtUweNhK1HBu2yVrMKZvSyTUf0VlbcwcMUHh
FOVMjG8vx8tcKr04GGR5j7tTQ5/xbxrmEIswae2uby+jN2fcZfBCpGrW6l2rAGkD
G9zHSEF57HyIx3ExQxXze/pj7HKQREqNSCEoz2jkX6eFLEBjmZyss+pzJ/xai5Oy
1tDjp6CgnBfhpClQfXNxL84NH6Y6ela5Cx94rY1hCYH2DeURZsP/sdHYR4dhctVS
AYkTbrxv2ZNRN305iC77U/DFvaHKL26K2MFVqoC14AS0D+q8GW2NZyjgN+xqPhKC
+NsWx0ZiOYxP9D+X146sKV7ukS60HhdVDLyVu/7CBjugQ5GjaFaS80Qvxx5eSrNV
ODakub6J6ftjrSUKwfGTL9nmJ2SINCKgWbtos9lYF/fXg9kxjtJYMTgH9pipr4KR
Kycrt9tmEmDtkVikzLDG9dVj7vGk7ofJZKb446n/qiBm0sYqRr6BorqIHsJUsTGr
uVa6Zq1W1VdhD/C2bYL96eRFchNYg+7SvO/deEMIY3kqeIGE5UhaoMT4cvKucktR
WMEc3b9uUr+cGGRkXQyLr0oFhZdtjO/+aSKT22rZroPxpoRu9kidECtQYg6YVXnH
p3hTklFlReoAkqYpawZbM8jAXf/Nvf0KMmMwuSHk8m4t+TAKThrmDMlTNKu1Vrui
KIshafVMsFL6kMkDObX2db2CBTNaGbfR2lstbb+ealuqDwIeUZVW8c5FdVD9aFqq
m/Eg1gYgQVx0H0x5DAlxK/rTEKcpYp870n/zzF82o8J/hkVnd+SWdB3Xcqbknr68
TxsWJ+D5g/sGn0lmtjRDQKwjv9Wm95n0WzdUsrcFCWM7NrFISqdCNRCRNT5pGqZG
9p/6vNEHmpIMh8UIGFyS/GGSj22yBDNpDH4x0eZnpqJhzgKfI4kZ4PPNMGNU5qXF
7mWJIgnisN8mI9kcb4kKIC8iTfcMgSvHKDyevFPytuC7tb49NmEkiqMezu+BBWdb
W9i9LHgyr9/A+7RJFIOapQKLgcQ3a5j8T9mDPYYCMnfP3y9LjqBxpgIS4v1y9Zja
mbbP0vFSlfz7w9OjOZ2xp2n1P8y23lwwcMU/UfLb5lLv78R7NdxZVP2GJSrJEW0Z
v+N5kgpnKNZN12+3/kfTePiF0jAzRPcQ6NjVf5KiGKyKBeZ7HNPd/t+V6WMq61WX
xahsXMQDjvTxVVlFhV2osLv02nwqQCkIrOayVTk5gzqTdGigFtfyLXHXr39Zx6co
76ZBj7LUHXHcMS+DQ1HaE3ugLxeEMNpRxsUPkHI9Gb2o2eUSyxWdwyC+Rm/U46EY
QmDNccQEjmDFtq1rUoLwSna8XSNKD00hLJARYHZeKBQqZh1lj6fQzAKtvN2c8Ien
uLfq4Oj782qmzx5GQD1C+ttoxc83v3gmSUUsPRywtV+s0iokQMvDmixuKxNQycPw
EVgWwdwnaBDNM4Mvms6WIgj7/6zxKsiLDdp8kSx/Q7GcuP23yjKUOzKnQXhlSWC/
uGzaioZGDneSg3xMhnHXgs9ORDnv1K24zWGsCMp9320WcYQLw0tAvF1RImZamJ9Q
mwioh0Eu2E7ViJ4SLZbr2IbNDLp9sHo+YepntgDvzrf0weTS/CMPcQUsmkNgp5QG
yuU71Ok9IDkXNRAFVzvutDugWKl0A2mE2sSn9359BeFxjGc8bBw1AnCJbpkFRxRm
bSlJo8nOoZUS4Hy6x6wy7M6kPX1AclTAXWxe8cSQaWn9VGktjkLGzppFjSI27aoC
yn9sQXdXp9nq2pBi7YUCCfyu7VoDN5PCVJrPt9IeGqTqcuFChO8zQJm7+/84cuzf
YvYYeDzcjLq3KoJFPFuoKW/8ETKcHQchxidUosg4TnXAfUaa9Ovo8hy9ileYUvbS
Sz86vLtZgJvnvgPtniLH/KfeuUSVFqf207rFWrVsjzr+x308qnGpnlQ3exFEIEFu
TzAHew2cpkxQcSkLiF1dQf8LSdcn7MHO0H/diUQuaVoWU9Nv//PPtrZqc4cGjR7H
YgjbRCzLqCcqzlsp4peDC7kihxOrPW2m4+Ydn9Yvk5gfGo3L3gDgtpP7ico3gy/0
qBNyA0yJS1W3tsVh2Bf1ka4pUh/D2uMhqcn083ZhAboe6MBlPjrdXgSnqEP7D9eq
wpdk7RFdEYBcQKrm8ct/6BaOCc4ZFU007zGBJYM9q/BkMZXtkhDkBhdIpLriySjZ
fD9y55ggggOhqyaWVPQ20wv6AL6YTBNM6gYov30DLoWqwuDKdV/4u7bzNa/ygcQK
+S3z1dVE1SWFAW/y8lTJVL45uTk853cM0MTdmkCG+JOKrFzV69up7nG3/3gMfsEP
rQbknVLh5yjaFNSWgbbBzJsNFcDZYt3nNtGmW6R9I7za1EHXvhM41e6liWsgHsG8
0cItUa77RZ4EDuwe6TVT89mVg5q9KQbs7aUKHIsVjtUsBv3AM89QhJ6ojamc8zW3
ZoRMnUPEOf/5hMHBT8Ot2C+4Ba9NOMNFvDtUfGc8qYfxabqFZ9u4s35n8e6mHB+s
Le9g+BQ95NlRqvGF81ulvQTqQDHIrGIDzDTUTyu0Xf1rks+TM5LD47b6ULYD0utx
uqWmXGvP8TWO6tNc33zyp37z3rZBBxlTJ/ZED5inRqY8vXk97wifuLhoyBdyRBP/
dWXvxjb5zEICsXgzRRza8c4XHxL7ARE7m1S8TekZN+3UiJxDni824P8vNwBItVQY
tB1XBWVwwfgSr8+RX3a/nNFAttRPWgIA5boWwz0aLddO+i/r7nHrWmLURK40HhCM
tuJsfT/weF0po4VVYXDSLDMMR4V7aX305XiikzqP6eRxy+hOl3Y9Nqmqof8ZcI6u
J8qvViJVzPTiBNtht/JktYjOQN4PCC0v+yRMfkL8lGq3eDZrB+HRKntwgiXP4kqr
A9kW73qNdwHh2M/8nyX1bAAWUBDQHJN5Zk1KMKe9UR+bQzr0/xDS38q4XS0Q0aYC
bAM5f7efGnLh5kAP09rhCyWCDKeyjBAsUgA/RJBWLejRSujbBBjL9XhktABlsWb+
CZNeSEqBEl46t6Nqho6ibcO22Kii/eAVVh2EkNJ+lQkGQMb1bYzu9K0MXf114P7H
AHqfhAh7rjNzmbXypxOQ9QbC8GepwVxOCYxOWJvoLDvqkmW6RDI0DFfn+yqBM5J9
OBinjOxwba+E6azgx92JA6ywyzOSc2sK2Xb2QTvaW+qS8P0ksPLOsJaJ3mPAbKg8
IJj5yt3f9JJMrtRJvfJeAzFJDOd7hoFHv1ZTknS2WrKr8EZVNRhX+wICJMPHmTnP
o/smiTLo6QwPCRr2RAFWarfroB1bkAcIMAszMZqMKCSh1rAg+SkX0p34bBZw/ObA
Va/Is1m9EstzhoUqlTxQm7DF8LzIrC53/42OUMrYuPNYHdRI5um6u1Ri2I4p3vYt
oeH5pBtj+D9rUEJ5JsduUw1zQRpPMu2fTVEVaVI5tHB9RUX9jrG7VX+YlKcf/cyB
tOELy7zsyTzPycEzxeYsHwkHTYOx4PaK99VmP/PWtm4qrO4os74D59Y+5CkAJyy6
tMxg5UUr97sJzaJCSwcO/RvFBqiTIuHqfFRshe24ln7pUxTJ1+/V9knLgQefIDF1
ohPR9uRBLhTi2xnnLNQaogQN6nT8Y9lUfuUlx+vxG4WktLoipJk+wZWydfi6EswC
vdax9Gys5wcDunp8H9n/A2WCtR14t21sV53LYKGWMcSev8JpcU6lKht6MZlRtr5B
bSVS+FW2feI/2CLbBbmB4RA4fr6KoRGpGyYFCuSfIqa3yhzy1os0UrIttFd8jX4Y
74xyl8DsejmwuHS2ngGRNo+5WC/W+j9UxfFBz/r6pvu4IHDwmhfTjdqrXv79Vh0R
3iWDgzXRu1rSpjIZUasocJfTX1j3wpdACTl4oE1pFNDiGnhXB57rlLd9iY+JQO5T
/+CEwJxxfDVTAJNqdMkwFHoGQtjy+iNiu6j0e83l22qFfby8NwMHuLw3mQRWYLHN
FVgGLrP9WLDWjF+eLUMsgy1xWHjIcAzgo10Ocq3Fz99vcHfnw/AGnfwSOO1Vy8UT
FJ9Icbva07TMftYZg97lkHszUYkXu2YMVIfL6f1TXs5Sd8yzGOjPwtTshXb+SxLc
nVatFxewzwutsp78IOc9ngonyLIhMQzYaw8rEO9nb/6+Y1qBn9g6uBWw0XtfVUsj
xA7KHoo2CXc9cmR81osMz0db/zvMiPMxAS5z01WWQ7UrR6QD/rZZXbR4tHOR5S5F
lHOD+wWHv1/F71Lh2We3Zx72RYA20D2OO/UQenZYs0Xl8KAiwejOJh4ZhiNC7BYF
1V1Qff0yBBKYQNXGTw6tVkt8Sji0VGczzQwed0lwKLiS+w1Ei+qbKckoMYRz78vo
ThgasUbHxdN/d8E9CU8PE3yYGN1GSbH93JqWb4a5/gm7RGDxNnutzAGuUVbHZjCI
RN11IL4506wNA7DQW+oTMlaoHLmgwSpJtPyhXMqnFo3NO780wGYD8sikO6ChZIFi
bNMGwPxC0Esv/t6Q8RTu4yvD/bYCUG0rNxTIlY6p1o2OPy3yh7H/LkcznZ6GvUNj
tnVBOOjYF0kTwT8weM3rv7A5iJzKSrUrkg53eLB1gJ4vJIHUbHChtiIC5cm4l7n6
LFoGDWKocTk5DoCSNgT48iFcptxWO/1fl90A+JMilDqTyDtdQ1GpVN29fbHgQSrv
xMOiTem/JZtD82WMZi1UtnCP9G/5UJbsPrcNothKNJQeJZyt2EhJpD4ucSYB7LrC
FdqwfpbHUg/mskG0gBoO1uh4OXN4aMFbf+v1f9/rbr7nuVlWfV5EgQoGsFa6xjJq
HFc7tcD5trS8DGRnhb55j4ZnwZJwU+IFmJqpngRPWFqUMWxPzdxu19HQgzJvyed5
1Wkd8S9POzJifcTVH0r+rcA3MNpHxEwGmGRVi/FFk1BufFejfzcc0F826kK9pNrj
vAEjE1q7/5x8bIgyvlEeGiKODOeOvd8Q+0MPtTf+zgZkDQ5oAt5PW1ZLfvI2U5hY
IqzWr5nTAtA6bqqZ8TYGdbhXUZi5H2lkNnz3U2PjmzubpJayJekrQ+TYMk2QK7yb
m9cqox/fivLxshkiQP3CsoeZdwodvhfvZ7QMe8mNQo320m0dnitSp7H2LacDXg9/
ukxdpt5fDlF+YQd9v3oYWBo/ipJJzcWbnJpIkqQiJcl8gLgkiAztM4C96OfNGNTq
tcHTro3zx4gBOgYNdAua3mmsb9BP+EmVrQK8yuqa7kFY24zB0RAEMiBwH/4FNc5G
hVfD9y1ffi0JFzzyNsSGyZTB6D6V3PQ0F55/bekTfIJFGmwnFwcAJIHBaC/JbUxa
IQ8t0N4ILBIcCPvJaB9MmUEOswmZjJW7kmdAMlu3sdVSPAZtytx8fIYpkv9GmCcb
zws6WSKqG/UCwhq7enKGx6909TqFG4QI5opPsyh8+lhZfPaVC0p80BWuxmrwa+mG
mTUT/5MQ0niLwepcZQ5Rdz3v5M01vKrtAZFRCj6iy8Qh7k12vkBMWDmc4Zcb3uPb
BFSIj53Qrpx40uFfRY5B7ajZM/bY/DjHnFStoxdDtFg1wFizfwx3UW6RkqquRdOC
Yow3LJqnQv11nf71+NH0EoI4AUahg5RNPi6YMsdpLBwAPBzqUoWquHhJPZKK2U8o
iyZs9Xd3JtYEDgdSkaApWjSbFvTtoOuBHqPnoC4kDClJyB3aeStyodUfU7171GsJ
JprDbBb/SgrkB2lcT8PM/YHdnNGGpbh9Www+VLV1gldcIrJGSgVHxta1hPgHmpGm
sjxK6AE45oiT7YDQuBFmTsarzco8lavMG7rQU0dPB8O4f+fFstlU+aK+QkGTCs/W
M5CGlCqr0qx1ixVpZgw6OyZCdw9+LX7Ukq7ImL7WmAv5GTw0OgH8Ejoecwg4jYyv
tzJGGkgFM5vQ07GO30mVGrR6GLzcvzC+Rez8X0gQe5CYolBvWyl+soLH1YHSBcgQ
HrXr9l+06vBzMaqmthR6OjjWLDyZ8Vt/JdXrp5Pq4OSEDXcSpPjkHt2jKUW4KkU7
pMLMJQtz93ryPirOJJ3i5BgbaEVj3BWeEF7wwW2Oxbw+Fc5bv/luc0j6HuK8UOhd
/vsddadNvYNkhYopqApk70H9vSOiB+VoPcVTwWmY1NBM1/Y0XUZeRjadIEhf46dE
gMzLyGYg6ttdcjtZUj7LmRYqw5rPTK0RiXh1iKDUHXLeG/+k5C06HgFjNAN8J69A
7Qc4VlG4VGZw42kaJS7gmr9reU6T5+OvAZRipdDprrBH5F3tageV7hzWZ4yX5XNO
ANVh/dOHV2aSZ12VgN2bmab4eJ60FuXBvZCy3widjbK9TtiUXMET7Ws+6i3YDASM
H7Itvwc5sdWQS1bELHW3KM5jRt8oiUQqOADREProcEdqZ4sPlDV1hr3cWA5YyTuq
kCvwYHmc1VqGsodNYLpro4qQ26igtErhsFzzuVOiz5RCi8aFIwCMhg9xDAZHp2L6
3DZ2TnS3JNscnY1SXI1gZ1z2belaZQcgWW4xyXcR+yXJkamzoe09YobpYAvoXnG7
1CLdlVeJ9z3L7Ru6urKRopf5iH/XYuyKmU9vXpmlyRXQPbMKSjt5iBghS9XBUf2S
i+fxvjeqWJIOMA8rN+aXs4YghlmY4ZOFoyn50l+IvZqr+GwGZ1Dg6s3pouMKt0G/
WjKnQXmakvfgHFx3lbQfQcqnzyzj+uWjymR3GQ6OW1TWpGzxRC/btwSx8390nIdh
QQLQmFUz+a8bkx7wv5BVVy+ZidecEXAhsWLuspIUnLVVuXg4ScspOfP/ONt18aGl
T8u1HplMJDwgXElp5m4inckxQ5JsbyACcNM57V8tV5O7Lb5PDeFGiNymVujQU68V
mXFZj5LoHFzob+Z/VhUYu6ZjgN7HK4SMcG3PQF0SNpqiIRSY+N4sUdcHE0FewniB
18SRKjvyKz/ph5gWL9JTjPTndFeRtrplcr0pqdFbVSBFYtlSUp3BJpLiWgsMaHBi
1yfvCbpJ/TY69Y66hUYZJQpblrHCsVSZUlV+O8pxNTMer3hBjA++aiqlw35OqHiY
u+8K1FFHdUA9kZVm9IFdOi5gMRaQMlx2Ud8CQmQ9im/+fLh8doCxeba9fVOBnixk
R5GGl+pkLBeFQGUO4zznv7LxzfL7lxKTmE/n4FO7bfbDpJoalHnXeStoVtDlCCwi
PTp7vhO52sXHJeqgGaNLOOEVt1QX3n4glqxSEzSH1WLtQtg7qsPQPUzze4VCf/tM
nmbxxrDXvK6UPTp/jSUbYxTGyy1cykmMuVU1cWn2cRlA55BGSPSFt6Vc8p1AUfGr
IfJkLsSZ377hckdI0ruBgGC7uEtXKk6tMMaSL2jjAoRH68fRTayOm26G7oyjvAOp
UyfWzMoZ2RZrB/oLm0HmGJNtFalWKq5oyueeYRDNTdijt0gTEwTJAMPIgcfDOQAN
POp33BMXpMzthIJxDAzKcNglHO1SNx5cmbTsNB6HosIxrhPU8uQA6lAtrKj6nZAX
hq1zY8Ia3adNI1PEHyhME6QYHJme5OrbZKYiWn5JYPSp89Em/N4nA7S1OupIXPId
+a1sqM2gnNQrJzqJ7FUWnTg892Xf2xrBRA5YS3YVIdsvX0jVNjYJ9X/Vi3BC0hdj
7FQgY9UuHND2AgJWQV4CrFhYMRcqqFyFMtB5rUafWJKwO1+t1BfVLQKQOcKdkYYl
JzzlDTUyE+3mPNll9lMB0lAJpK9bu9EkBUKs7Vv/Y3wNCIiWHs1vc8rMGPXGpDxw
xtB6DBBsXfPTCKkeL0Q+CSaG1v2vRZaNX+fzFKLUS3aThxfVFhLTTDIw26RXdNTH
uXFYyI3TO7jh54Jx1eropfgu9v0xgQc4QXjtTxfGBV1C7+EeDiFEhFd9ABS7xT1/
FjSZ79Mdc/5EBVwrOz5X2zaI4460VmUHhCgwNgCs7MJflW8gePzYpATMqxsXU4e8
4fxhbmf8jyDL5xJXRdFdEVMK4cB/OPAUfKPDB4ISTWCigi8XVdtknaFCA8UBy4XB
uiOBjOj5etcnJLwmGkMEGnDnWT0H32MEZyLvqqCuxOEZQvMAI1AUVZW6ZF+xczRl
bZ6Rh0UkanHcHoFogA9/mkrrnzto1CPpfPAYwL7KImidevYXes9GiTl6/Rxr5vMQ
gnQD+P8hmLZ9oISV0CDq0+KZ7Ge9HIbrsltc7pamz++TuA1O1PjJbQxSrcnlLPLt
M+RhfPYrIPRDCGSY1okxiqLRae0GtS3NY5KAKB+m0w5IyUnu6EF8/UsnT+i8qIdI
rWeXMOYAwgwXm3Ebw/VYfFDSCvx/7jp0ZgxUdc6TQWTz7gcCA7vaOOUtPwPX474d
37hi5SWf6ZWtFANWb9gz/8+Uv+G9A9YhjxqQehHWBZsoCIOmJPgoRUCkzdUZX2B2
lCnVKYtl9I9YltjYhgFJ4pQ/glIyGGagbJDMz2cRakP9dtpgIhvbHPKa+O5MoQhz
71vi7D+bpFENR9cGTjp7cKNvH5/E5mRGeEMMgi8Puxg71HqnxwOngK00B1jZxTk6
qAjV2rgzdmC54uAa+2qAMddEeBBmjZJDz6H+8UJnOUBEBPwXDhg4+U0NqFuU472K
b18qOtYFNEnc5wr3ZWvbdyrNHxTiM3nwaywHNqhHyZO//F5u1U760AtyFycIj2Lh
wId44I93r5oO4Iu09bWvDmxGvRCM1ZgAxjr8Mgx9C6t014WitvLekzxXaLXGkvrW
S3ZvbjCStT7n39YPap27Mv9Ubk3xVIChFr7uUGOnE7OvSzFl52YZlEYhtJaxOet/
RtLFH5kW62y3VHdkUVRD+ESkCDLGfhT//HdaZ6rceT/g58SAaWtDtKbync9ttnqR
ypoMpUHDPB9IOASp8+08YAH/ZqBw4jAqAUlDp2S4asfKl8RDbjr6E1MKlg4Q+PxQ
gyPSBHxaJDiyPIWHLAsGqCaZDTr/iP08Cel9iWvgWH4DImDmN4QbNDVTB6NDokue
H7KYV5ROHouUgXuw2/ITDS2TWKd4jvJD0sBVOZEug57A5+GslZPffKRkqkCA/XYA
XtK4+SaBf1+BbWpUK0dvEYQCX12e0BqZVDCkaMTcvfMYFSsThPBQYxs4oOvRviUA
o87x46vIZ/YPgeF52bMWBrGgJhqWTAmPkHR/HUwJZvLTCSQ27h3FkvPitSe6KGxm
GneJGBOpmVOYTVc8h/f11t4+pMe9FBQulTtcuLZRdRM/P3ckfibi5GYIi/DD+5NN
XMQO4sUsk8mtaT1qra9DBkhg0baZKtu4hTF5gmyN212gLFYyO3K4fTnXY73ZMiHd
a4uBZ7YoycIychxbPdIgtsBHNQuQaMRkODiXzBLku85grUQcjVSYLXlVdq/gWXIa
oPdkorFcNNY6nsv7ms4UBY7VWzf7GRvaBhZogg2NcfEU4S7CxXQUOMTU1iSM4Cbu
NDnPBNTlUVRDyOy/b7Z0XG8WFdD/rDDvkqfGxYWZ9HsCIHRmIV+A/S9qoc/TRQrs
N2qWJizkUceXzlP5daMi2MMc/Wnf+O1N58l8QyhOshLkbj+Qt6f2PxdyBCM3zOYm
hoSWhR13lD7JQ7mgd/ii7ZVICeBKia7OhYu5K8KiNd+CPGV+RKAiuzdhygHE4pR8
2dqvM4A3zvubLyAiY4I3YSTaY9evRHT7yt8aBVERJznszB+L7rudMiz2lzU98mVL
XptgIzGiKIyRpoYz523byVbBeJakSgirNSjMox82/qjCx9wbKDnGAWp6K5bgU2eJ
nOa4h/Sm99hA7aOjscjo8qmUYBGVbVolqhQUWqlWIV/ePzeTSm8xQQD2hbVzgj/6
Hjc4bemlTuaNbHj/qjTQrzI8AU6PV1R04AXNrfk7eKUjEWrTa/AYEdG6W9OuNOD2
cu4Qnv0E2UMVaZJEEeQklXRYcfD9zJX44qVjvFC0Q7i1pOkLGHmnf2AZjk3h/HrY
mN05RKUGfoxwWq9LfD1e1APiBLxqlgwdgRxmqBULItDvm7i3BQSZw3nt9CwGZSFX
g4XhloS4k4PuHbY71+ChiV6DsSnIlkYC56ajftOo4zVBZXqycrOLI1FdzTPqcoPm
QuKeGDG/S68tP1DDfixad/rt2g+G/LA4ElsPWmXtCO+tM2PNToctrGe2L5k8LS2i
Eu5cpho0YaKA5H8AH6OkGILdzahsr6YLWgyIwE3UNKFD+yaLSGdth0hhUc38nftu
OmtoNkKCfv5PTZNuhilp1mfGXHsPAYbfwN8tx+QRa9PqNvAxRDDv/JEtAtkvzwv8
W1bEkazm1tLcfe2a1jEuGZmtlTceh80bOt5A70+/GCOJlMfh81Y8yL3McE2V73g4
LWrZR7KDP2rbTgbeXDmnm00CmsKnlyDWrTGa+zBP9sImOyeYMDgavbKJgelM7Hc1
O/R9oodpf6UpTPu+v1C+FVme35znvzp/T0oG9AlHdCenpyeWgSp37EawoC6mUJVL
zlweq6G/3ANl5KMEKzkhMnTMkrhEZlNS/epnhRh/m51gkYc+H4ZwXK/QiLHfTiux
UJvw5QIFzwOnqyKmOWVPzaaC3Rg8+k6GSPlZjKogucCo+shArgM45472S681rNXM
b63ULKcRdPntr/R8otPDV8AHCaPF31fmjCWwk/UZbq9O0Pu51kJ8RtEH5l2ftpFs
Crh47QOkvVxoPHxrWJVeaJphlrKTx4RO6Mk7UYAyWa7nvf6vrk/yKwjc0Xwo1/Fd
lP+X0Lv5eCGvIdYIysiotsKR+DVBoi/HE4onfvdcIALeM621o4BSNf2S1ahSxSEW
JJXNS+BmTIdSLEZaELqsb9GyH3ezTfHarQ7Q0lk1rAdpBM1hxvN7ntyhUCjDjckD
hIM3ubNafiGPSriHMvTk1mAqdkoKYHSRZIvzPAmkI9Zr4s3rhDc7ip8p5CdAxEbx
f7jpcUcTEmbhuTajE38ehkE6/9w8q22e2+PGwFv37jRXfQvLlXisHVdaYa+lzVwE
iSbVWx9WC1d4LZ+n/bRcnx0rr/c76FC7WhvWdldoUrxCfE6FxJwLpH09Kz5o1kwE
rrXRdCHaga9Ecr98f0ez+JQiRbN0+CVB6AJTeQWjEgT9MfkAgMQH+V+3/kPkBqeA
Z/ckmzYXKzLVf1f69YTFkBUau3RAR3l4jzAKFH8IzQs6Ynxn7QG8GJ1g5R9MqhM7
2LcwzL4QdcN3lxLzvwx387IlBNj//cG9FjDGFsaHR//YZqx06y/j056uN8BWvjzZ
yHOhwD3fs/A4+b9CpPIfCJYJMBscYH4k3vKcsAc0Vh+s2qHUDkgF2luxjYTRjbyd
V8o3i/OjGDJd8u/00xw5O/eMFK9TcZ88pcedDW7ddD97jqA45oQo4JjBlSUNa5JB
2/tBuhnvDpKRUvGuGiD3bR5y8PahcjiRal/THEdDzTN3KDxzd79qPIArxLSFgaqe
OLgsiO7SnEVTxy6fegepWZxmFGZdyZO+V2PS/Vmmt+kxhdoohNXKXmfD4m7dnoHd
GpecYiIO403CReWuggUP4Vn1+VFGkfJ+vboZgAdbFUg69JlvnrsK9Nb1K6nUm2fr
IeplZ6lg2j1ThUQ4ES1zjpKQZmHT7dAR95iMDI2d2Fa+BbYanMORnK+IAbBTSI0T
54tE/e1cFzD/ShTEQIPOavnie2ZoGuGbcUFo2O97I8fITumYZNS6yCh0m3yjtk6T
sSyxPkRaW4xSb1yAX2EllirxgvJO9KjFpwW4e/wsWM6F1vUQySk3dcZiKn3Ac8dR
b9aJ1gQ52LO7Sc0UfzCTEzCKGc3+DsZ6RKdNXEqPsewFbtGeuyujDrngABc7InUg
QhFfKdajOu5aXbxbA9Uq1esA4VRcHoWY/U3QfRODT47sU1Rhphg7EL3l40AysX7K
VnUJvYthsDBkvzL44n9n3/QNnE0NDOv2nHtkZY4JMKAIRTk9RdU+3Z4zZfXlMidu
MTNT+1xzHYJLsDmKAxTzm80NSvhI15OyUFgEL3l97PZvv5NYx64k/JV2N2BTwBBY
smN9hyz5grssdMe2x+K/5QllUQrvRLRyVCHtvm85/5bDPbv9WKxwR2BTOx3QAgbq
Qft2+GPCByp5MfBeT/DDbd0LcRO0kQbtksD/gB+CpaSH69TyglqB0MMcuX3p8ySz
Xx7TpyCo+IJtoEFzDYsFQpnNZ6TrNdU/oxjhRbuW7se/so3FY8jxxD2EtUwfn5Ad
WmsYSyamPCEdNvKbP8x7tzqr5w3ZBmUlRwad5FkELr1HREYot+xLaxO7mzJfEhf4
lLKxrKMpsOY7wL8dSmch7imF9fiAvBFz7Jsa3igaQqUYk0j2ynzO7XytgS2kLNeZ
ki9O0Bm14cCy98PH2GEdSuPYtLI5oD7T2eImjCIN2hhyDaVyKicIUUFAhUPZJocY
eFzN0YV7p1Y36CHhcnr87Wart/hX6YASfM9W/4lBi/36HHH8V8OT8SepD4MkFZVM
lh+MWBF446Xwjf82rc0qYNmqGaTytjY+6PByFc0iRoMnap3u+vgqH+nhqXv+2BAQ
uzltILVtyX0YaIg1eAZW9hvO4j4XF5ejIysSq0qnRBLuVmCBiTENrr73KRI3RwKq
T58iHvS3IDguvPDV5L8KUs6Lu1S24vMQjuVLk3sUN0YW+jQnOFuv4IRQe/mrtdpy
brsuENr7iVJ9jTyjY9AmLWwpKFHTQdaL6voNQvvb5fQIY2/qKJ4x3VhGpbLs5DPx
u8zsQDpVumPRGoFZ5ivVkMOxuL9/r0ISZtkn/ZXT6nEaoFgL8koKAC1tQEmb5Wdx
WRAyFauozTwzNeNhzQRWNbdV5YlzOcMzRYlF/WWAmfDFM/b7TxOeiclkfriFUUnX
7RQHfSdbmxHDI4Nmcfc+ITGBvHmzN7CSr/D86c2s7/rQ4+Fl9wymRM/P18jkHigK
IByoYVbfiZcNXY3OTx2URraceUX+1icrKeBzEFhV9Eq0HteAvZvLo+86OkY6Gj6q
ElWDvqKnV8s6LBC6zRn/4GJtsV+GZw6H2mESSQJgtfbW4Ciy1LrsBSotHgy6XI5S
zlzIkKDVYflYhYb47FVIxerp4ynjhDvAFMzJhVpxOMqEo21vZnrkYfO6451S0mFh
xb1/oh16Pm2VSKoT+/u9jmGuPBtX/u3gNfgTioJFRU/HSyV/Y84XYoT2swrDB0JI
GN3rqPl8hzod91YkWM3U00h3M9UYUC6bLz9CcmfEO9YoQzbUCgskwMS/DZ0xyLfc
e+0BcApIQ+tEshhHPnMwzWxuQv6C4vs+MSSd/8f4AM/AhukRljGr6J1EguSD6ZSo
HjMOg4sJuoIzNEh5PfcJ8GDpKLd6womUQWPVfmXSe0EU6osJQ3lKALTgMmp/JGs4
TxBe+olX7ljeRDaKETOqHrzmYfk86T/9hkMqqCodh5Nd2fb1z/UqaM+blnDuORRM
jU82pDGv/tp44E956Hjoav7TVfSXt74/mqYE/vxpW3KWTalwXRtTKXhVHh2DrMJW
HzccB7kIkZeq0kWNvwStSigBUP1VFFEUz4k0yKxX77TSc1dp0YESy2r4TqJAS/yS
R0irLPyENA9T/Jov6tKtnJCPyQbzsOK0jWuiYcxt4mXRGSiidL+SAFJ36XXv+Kbi
fMmfJXN8b1/CNOllFiWuGuSZW6ctOy8PS09JHFKWUhQQGwebzUDTqNrG1Po81x5E
NRj64TIwzsAma7uiwXbdadzPOO0kO8m0fgn0RuDdPPGh3IBMJBn5p1q1hGrwNth5
Z8LGOzyessCl7rP26taFjJ5eh3/dgvP0FdgY4IOV7iRyC8ekzWfrQ0Yb+AWP9UVr
SGus1r0HKLvYmQzBXaBy05ktGkLjQ62v956kc2YG2HxUTAKoyNscIlQdUt+d6A2i
Ooho/7uDvb37xuSJstbit/wtADThiXDY2wmzKJfa26l6F3nuFHUrcFEvoKkNRSci
wd+Ga9I/4y/zSHCzS4/OjCI+PqoXNdbnuZj+A+Gmda0HORooy6GBc8hirsF+dmKb
TbhHrNjQyx2Qit3pJvIsKvy6KZh/b/9uytuYqZpbsDlrJGPZ9Z6rS54UtK+VYLej
Ep7h5yeWr320c1xX0fS71QL46Go/AkIsz5b6UXFDG4GneeEvesj+U/TN1cp6EPG8
QcGOg2wtGBPd7TNbIo60Gmpk6koiTBAghulge9mhN8Ex/SHZad50gmoPMuAhqYAm
E94a+kHs4KEy3Gxj+G4QP7s+z4dBnUQww+sUE/HMhWNnGCc7bKQ/Dy5MS1Y4QZ23
2WK71E4PAm4eWu6C+Vmw7W3eBWeoGqtbcTVVb19HVHmRCCxSY1stMC6EKfsesiiV
GZqTv0g3IIlgs5HpXvkMxXk57EKOnYjiG69ZmplFcXaDZqqv3OfpWCQFuXMPxrHg
UJecKF+rshof4lnvTV+TujKythvM7j/BNU5pFhdbJTi1EDI4lZ74L8W8hYXNE/Ev
MEqS7FMcWfOMF94JrU9LvOepwLzXP2HjybpYVqzsZkCSlN5l4mfuSB9znuiCPzLV
jCwFvmw9xjkGmWx5pP5fS6pvx+SGMqSNN4V3iKPbj3b6ER+JkSl4zEAF4Nu+GJsb
IhRgFSBxBbiLmwP2q5pd62iF6i4junyoIdvmKIVDbktojSySZvkOKISW/ZopMhIo
LLtOta1ERX3VjfTFtmRGFnYpdgjWEriubLlD6Uf0ESqYOu6SSqQJIMC/p8w5wMbD
WBiJVjBiRQAkig1CeAdX6IcCu9WnkJ7WM+Di12nh0QwWb2BCRX8CY8VNUd086qqu
mGyaehKLFLGKieAYOAP1lW5Ok0ZkHZ2RZjSiNSQ0kQqSipucrlM+Vtt3MXiZBDy9
tl/1Cu19zn4PjjPrtTGwNqKxzJJXJuyqjCU8UbCy+DRSkuUOsZQg/zzMAEvzPHlN
TrEATN+W4N1gsUDawT4iyn5tZ9+wnz/lMozfvKAJ5tIDFymQBTPHxuyEuV16QfaI
KKmckwQ7ivUAbLJ7lEG0F7UApQc0QwSpBsADZ/L0NMalGVuVvo3H6cchmtAhmtCL
nxIArxgzYx8Y+/brlFmhjlqqjY2x7fSY2744DkzlODukH5QFVliC9h6E0ujGk2Io
1pEPH6Yh+sVhuDTcjSwlbGU/tslRW2RXA5ut75JQWkA1SeSNTMB2JUWOBzU2/baZ
1y+Aie+kH0CX5xxj9ixAPUKM2YtSUg95FUa01t5yvGzhg4ImRj9aisidvVtB45be
6FhoqgBfsGp0k0ueBeeMMiE5m+cQkIM8CE8ox8lV1dFi3IbkoJmlQEykn1RRuk1c
yBN3XhFHSa7VDoNCd9oJzBZTA/3vnrb2HmMUsoUyn3KIq+qix3zbh6xK5jnvKjSg
Uzw3skVrWWOy/sMHnwDuzB3fvsFd09gr3KdmXmwcVIwQ9WVSmv4u19tGKy+w7CGi
DFoYDY5zfXXSE20auV4WxUjgZHmdiHZhx2oDldVo6m6QyDOoJYtOX1NML1ALHQPb
rXTwhT6mOFvsWXRyAL6NweISC6c7oRhTfeJEUOF3mzypj9iqoQqc0gp8Mc4ezKvX
aWQwg1Vl451ko6X1RYJRcV38Pv3XZZvuxbksm9xMQgIekH4m6+uWbhKwYOwbUEwt
PfmQwYeCxHi4iihSToXYBAnojvC6vUaGHn3gTa5xQmcPlxAthAgxv1Sp40c6gXZu
ROecDTlvdNyD1eNm+vC3lWxbM6FvBo4wQ7hczimV0yal6d/xWUBdlrOWfSd8qRbJ
IgcFTNCnwqpar6KniiG/zoAbUm+tc5oZH+4mCt7VAfcCreb4xTGqIZDslZygJsoT
VxhOAy2XsUCTp83/G69j23vlpkEpmSo8jRCvDyQIt9XlpbyIaadAvGLuAxhubgEM
iGLin4y7W5tOH1y2x/5nep8xgBX+cL+sW5n+9tksoih/nZBqGQStGlE6dG7KrBFw
nGlzL6Ni+wKo9YdwudiCyNjjv2GDRY6blcljen21aai37PxLyU0sNHtxDzrYiyiJ
DdAhcuCOXmdTOrsXZNLdWPPojSVYAoxSzWHFUmV4q8qIr5LFYb7godBR+nhVbqLv
lniccK/tZ2fY4kIT17aM0rEXan+uJiPWaJjlN21t6gXi1Gwnoyo8mg7JNiCCWwBG
rBqyjWaivTEC93EabsaMwSkWQMQ9p+0Ktb8uX03y3C9lOJKEU6155SXwtWgdJBph
J5lqHe/VXT+rlRntQ7KGuz9QJu4qTkUOR8bI8Zj+Y7xnGBDx2fRBmPb9rgTMuTnv
AL9iL64eBjHabIqT6GLbIfvKUFqJQY/GfJHC36SlzRR60QEXpzfrLcfjZ149a4DF
rbEbDVbAG11RdV6evGM0NJbbUPQtGdwKoomxZDeDj0jkbSv85iHA5haDuUShGpT3
5/cjZiOq4NT0+SV9ycnzqWme7KTAYi3T2A3lnpc9h5EYuc6LsRqfXfdJivrwWOmf
Ihe/3lXspvxiCISzeDBSElpmg0ijbId42IYOM5Joi2f5PgtTHj75lsfh76bOdSaY
IEA3iXTTqIhrb9Swe3bO19RkOdF9B15FA2pVCte8bw16tAwMFvyHTDnTaJhOxElG
yRiAUp9bzY++NhFVeVRMN+KzrxGmkbKffyWp7ErCeeXWWpKMICx6PmoqPYsA+NP4
xag5nFZAxoDPcCeBQdbJednem7KKBaxVlyJhk0eQ7KtXgL+4zECas1YcCzSgIY06
jHG7R5HXLqfjIk8DX+RhUmYbxwLCp238IobOb/HICTVXe2AI9d7E2G7lh8iskaO+
ThaSIakf95wGIb+ct/YvYRDjlwl9l2/XzyagcXKSicfUAAxERHW6J1EjUVyZdhg5
s9ZstmGNHZqVEaVTTuRuXSgD6nd6NGH0HRs+8nat1+pCDGJtDV5p57FkwdsBvCcO
SzrlrpWDsXcpvqZ9PP8og+ndtoAyPJT1b1it8Zdw2KD8qgKzRzu31bn+6FD2c1EG
2bGE5CpDwbnaO6DeAmzKHyxQhM/qF3bi0WwMaJCoPZZ+fdo+rntlxapJhP8rJ5A3
7bWwZSOTf7uhC9gE+4lP1mJ9Ewg4rSwQtYchmkNK7LL9cKec1qPqTxKGP2y/CmqC
jIwjP5oEHKqCNSpzCNNCZGz+cXGDp4+pGsufdDTrYih9lCSJEmEW6AKLP/d4pp/J
mThIMGvzESp1d77ON/Yn0aZT4IUN/Of6yzS8+AhzBYXPb+NM8nnoEyXNGQU6tX1w
WP+2BTJpBjEMlYO4rrZnJR+LGJYEtpr/DELQsPEfF4NhcTINcAKjeVm6/i+lHRxt
5yBSLAtFVUblk+ff9YIbjCuK8g91B1smVyC/Nh+RcL1helk5Oz9NnSPA+56f4EYl
Bu8LHtJmL2/X8tAecB4AV0Xpty/Tv7OMIKSQMq5MfrIpSdyBOB42EpJux0VYTieG
MjYKdvEPVU4sHUD1kRAsSF9RwshjqBuJc+5pYp6zdCLzgl9DKhy86U7sgTFM37L8
7Pe0cBf0xtqisrK0eJo13JPnHHcvRhEwdEL77kg/PDD7ImsApmOr9eLj/Bzeh+M7
QPcSMpRVoCJ3KNRKwCFUPCYy1RSccWYzX72RBk4z3J473Ioe3oy8kgyoJVdjYxc+
/D5EIOjH52ef/wf3f7mIXgVcgjrr8b0bnBzW2Uk8zXiHZ9npJ1cQokAFNa1cz1CH
tLkPqndxYAx2QQOIbm5IJClntxg13coD/rXZHGFLHzcsi+uCiHBn6q5fmOaeVfFw
nTyVlWWPhwTypSBZoYYTne5R1Ze83YAGDFLQU2NgaZm9ylk9z+kFmgvQmZRNp0Gb
djq95VlPR61OahjqLZriepv+X0T30NUdDb4I2eg61PfuScwTp+iHO0mHtLFFrEm9
sB6TWcU7u4igMD9yujU7raApnZxUbr01XKSYDyNxN67Wmy/qUBIEqHAx41CykuoQ
Ja6nTuU8111RI/nBH8Phxu6QGkwa7PwXdRxjdPVGeQLz4gycSHRRw7loNkY1nZR8
3zB5BYE/pF0zlTXVdPDHrkFOGkCt8fkbGyY6Jq7h0U+rS5cHCjHLNXBBeqhaorY1
qpUqaixbVN1OaPOoiQJE+IE+h6EM5zXwOuoHzGvNCSHl5Go1gksU9jM8jeaPYmyx
VgrjmQmeJy+Ls3n9Qy0GdqKHGHIb8CPhEUnJ89fRahf3byt6xQWXcw600sJaCaMX
rvkiRgblp9CfwPs8b5Pm+r0mEFbgTiuC29xDsqTjrz+Q3j6KgHtY7BL0/2s4LU4c
KZjZtFuWokYdo6qK6nShVRHng6xgj4WdG3L5O3281Y/+mbb1kI+V0yPufHN4rCi5
gdB3SH1mzYYnAs77j95rUT7V4mIKB+Aby5sQWcA9GbDk59ys9ywEWHxo3jmfeMLR
6LO4jx9ubGjC1AhoKg5pywSnQwUoGP3I7uZSM2sM73ZAq7l6MPYUzq5BI1LC+7QI
fks3wW2BtL5RWW5Pkjpyr2MtqX8/HySrAJU62I6sZs8DCQyahFnPaHu1IGWSIwkK
DiSQDDu8XMyD1O9DgYEeGgTq0yz8POyt52YBGFPtSdv/s+8y/KR6sjvYkvjITU7p
lknQrAEmVT5HLI1P2vcE+yQ1vVULFKSBnrn/ECX9Iyx5t0ifcGf4FrcJVWGhoQOD
+obZx67yvVO6CERqfLLYkWkgt0lqvyeKAZqDrTa/adPTspdZOSv4GHqiSNPs26nh
/v0GFnO8tgqkKPP5V4Pfx1cNGZwOj604h6mLL8yQd3El8z8ElD3QrGVcg+PlfzNy
rN6Xen6CWs7SJeudOswa2rEavkkve6hbwii10hO0w3r3YfAuMY+mf3uwMrFNwRqB
mSYLGR4SOP7cQ78WDAq2E6BF4e8fgSY8Ci9ssMNnGOJsmEBQ9YOK4gmeXhaCHJXz
dh/tPbpTxmmeRdfx2zuq+GVvfBETQ7NJjuLibd0OFs0RBsEtSH9oGUIWDOTMTPJg
mCeUEsYc/89V4QeDK6ZjxuEf7/mFIJKptlvhwieYt9SN19lvhula7d5HPpDmQizc
+PfD2+3zpWLMA2y0qdc3gGR0OMchkcx1CIoyAIilXP5/abrG1THyTNQ3ZDrHgYAY
ipfyxLudnHHQ3II17y4EWmK0s6jnNZR0jGrffKQ0jS3hwi7t9E9Tx2Hq4J2ThLLu
TU2W527Quykjv56Ftm8XJT/aH79aG5epycYbgui4bO0BYDJO+8i6/BcboJbn09No
PyRe/BrBMNPRACmpQaYhE8zblTQWMYhrOqMY6Bz0rcpczsJzJeApvmavvRZgsdNM
lxbGD/4KgTAcU9Us+OMfL8yy58mOdxUGMgGMa9nq9A1CqKLAb6Cxnt7d8TEBdicC
LHqyYa0ViwRRZKKB8DYQYPKYHFqoNMYiyKEg3csGfdnJLzw5+ZgPb3/YqqPgd8Eo
wqyc2GqOyLt3MshUoARMJwwDwH0XCvHaSYs2y6qUZo+4HAeGtEQdesp67iyqkt39
WZ3t9ZDiY1BI/JJp3VMt2/yuEsFwtnRxuB0wWquKuwytLe6guUXbxTzce1u/uYSD
5OnSrMeRykYnmSK+QhE5day2udw0S7264WQYqGEGqJ9geuSKNOc3MZ54VTaKi9JA
+WwQfOX2R1DLp8ELA4Iqgo4UY9IxfC7HQNLDUb4RAu//q9QJ4GPmlHepcMMR+Ovk
TNHtXhYcuYIxSEOUdBpRKW7OPdSquTCB7BoEf3ulXD95FI14X9VyPqtYQIukfoTs
e8+s+X9WakReeJ1Dro4JlFPlm+dn6HzbRKke+gXRdH9I9Awh+Bj82M7N1m/Dpro1
6/lcr/WHlp+YtCOQYL1xvSvHYc2gI7JuoAfXBJ8yG6zUj11AvN7cKh0W7nOE+6xs
f/tfSyNx8G98F3ZPWFHFbipcKJZqeDURcMrWAl6oFtONsDMuhVAirq18xei0Rusx
kwT3OiNhDOPIKW/pHdL0OTr1n3NlF5ie8viloBw1EYB6oY8t+bX6V5Qnb3J5lodG
cJHpYQ1w0chmGC3N+mLe/If3bM8yMYhjlm90wjG88gj94dR3DkyICTPcvtKicaC6
6ko0/IpRawlMZa8Z/O+d5fV7bcKWwSEKZar4AMRQkejhHn5mvB9zuDXI9pvKbRJ7
0qyqfD3ctsYCkMopuK8DvkhvXjwE+mZDS66695cAf31AczCdSGkDGYIc4FfEjy6W
qzRmaqqkZqxzVRwiTF9Ds+WSqgUoLntIGx4Vg2EYqqE16zNw1vJf2EbeiyGGmDNX
GaI6bztaXs0tH69FwIEhG++dyL11pIuu3VIYgEO2ftojGD7SXdhjyzhwE7tQtQGw
nk+QfBkbYo6QDjoAPUNFnz6C0t3YkIsEHT+D7vvqzzb8dpQEufBwBqB4au/mZcR7
JlQjkyHzw+jGlarmyVZW34EQ+oYwZgyKZ3Aj2pSPpl9W3XMZwiZ1ZyETaPISjCkT
dIns6yTdb0QDtnAiLqDvMDdyeg9P4dY939638dpwPk4BszTT2QDFCGVgmdGFthOe
s57LKAkLqDefzVNf1d/73vjxc5EhOGb5Nfqx7dMctJHjoUAj83d+ekEy6cbNA5AX
F33gsJ3fU6U2e0LOzatr6T9zDVdGWEOnuoVBmwA5Ci23f8q6LrNPI5JSXNsYPQWP
1V93YPk5FDZ0E3ayMWZCVkHk1ATtnTNzAEJn8403IgAlt4+ArrY4Irgn+5+7JmUY
WLd3AJPWeTtb6MlFPV3CTWYfRtCySpmNDJ9p9wwQTiwMJrAoqDeSR2PmkUNxemct
AR9dPtE7TVoGAY0qEvFFRlkRFysE3rujyIxH3F7sq8zX0Wy672chxIk7qoQgHOhh
xNFYTbe4p9WxT04Zs77hoeXhK2dlM0rsNKGSiytfBtkkHnP11NDy+79wlGrd2Bp2
KdbWfg/GfS3IKFfeoMMgOLeMh3D42/SATLfeoZQRvHvDSgj4v76vIFHei+e+TAK8
1Ll1jWno71WivOU2xPvFBErlIfAYifEiK2+ZBU2TYfzIL7mC1Xf1V9o8maRwTRA3
l93m2xivffFY4SohoTHLOJuinqcfQzOuz6/jpFK/8mILds/ANwwn8IxboHcCQwnr
dAsBrknMjv/fpLd1uLRQMfHp0gaVI2IGgw9tTTw1qVyzZOmy5kpARc8bglHasw0r
xGrGfG/IUYl1iQiAxSC8Kja8PXJRQe7ljSHcS2ttQV9n/GTmjDiWtR7P6disouhz
YNb3jtUoIZTXE0znejsoBCNQsMqGjz6GD9t8AhJJjx7ZKBiUhfNEVyXptthKOCso
9i5WO89mTutMShWp7gmt0gQCwuqFYagWwGtkerYwPAA+Fy/EPvMJm9R4amOOhJpk
/fwVe4YIkVIgCYXXjgiLB/VZ6uuG4ASUMOOhjSY+NnEW9F+uVkjw+mnXHv71kRYY
TauIZaSiWoyeSaFFeOM5OLxBnHfqoY+14lZgv5Vb9LdWZvTjfhR4ml6EJvY85XSg
cwo1z/Et4HmX0z8HXaYradLaeNxluM8jvXksZ/BqFhD2nT1WFrnbDvzU0blbE5s2
kXvddzT6kxaK3V5YKbKtYHkDOq8E5VxyxD1gGIN9yZlWBksQbxHfesP9f6ZwaNhe
XUQDJcn3eLqxqeYoAApUkNQQ92EqfmUUJFkxSVtGaWtIt3SDMH5YqZwAzbjPJt1/
TyS+M4D+btyIUj4oLyikEOl/m1H8oNFv1Tl6EJEtl4P1tZPqTn9FI7W7FwtJlGST
pNL9gVcujMXozO0bpzQhmciNQcLT7B4peME07JFtDSxjZrUlvQSJ1dVr9mLvI5Hb
AGUJKkWft2ECP9psW0ddYFjGQdQPPAmBA+rup/6q4YUt5m3O5v0+Y7g7S//kvZJo
ejr2d5o67hIqA/S1ahypfsNahPWJ3RRGpKEsYIqoNhY9x/LB80Et1lWfiwpBCE1Z
PpXBaXo6j+hzlimrS6XwnOZw5Ujl7LyhBLkOfgc8vYrvm8gyAcmdMefs46v+c4f2
RuKwiEL8g5v54qZiujayvAHR8TXWuHroJ9+QEsOk+GGkupkR6Q7rVO9n2IRi59+C
hZu8Kxsuu2PkDv3xW19g1NsxCoYdv22j7WhXJDseA9DTINsz0d8lkOY4GyKWJ80g
ih3/nHy0CgyVah6VIoxfH6i+QVyNLg3qDxZp16mPRe06kG+XdjeNqpUjvd+7RXUO
EKVpolSAqrZLRi3zKoT+02ydQLQ9aY7wYx0+pPAD+QVmgDc8CKs+8p7BFhppkNFJ
Bcxvb2xwXVeiwW1J2EWNgX98u17Ifl/fVzW+MKbMUGGr23Tsi3PF6NJlKk3MwF3P
Vy0s0IvKMDDNgXTPLognFD9iCJkC4ceTrL8D64Qsl+70HbY8I8svF2MR34P6FdFs
giZ9Wa35SomDZFEc72dyHA6yZjSQeoS/cgWNMgfBP6fFsI26W2hVP1iktyWuMtF5
zfzbvgK+ykilG6S306hWxkRh8ztzNotBEXLVw3Fme4KAHW92sxWo31k2P1FgjX9l
EMs17+/dskDaV8cpXGn3xDMLyqrK4fYoxfr2E0RQWaPHX6tB0cKJdj1f5gPIgmWT
QrawWEkdjJbIkEdRcPGYBsf0iaHIpKtwFDNtwadwLgTkGEjdtU9ikmN3K0KtKii1
rgvAYNFopJpDXpjxBACWSFWNb0DqTlIXk6AirU2CRw8fjtr/xvqvbpdNhSv+46Nb
06/hWIvCzkfkoe2f2FctOtkb6pxop2gCobiQ+G7o3JVBsg7zDpDct11H67imEB+0
MbBv4VVcQ9evY0izrMcoTlUuM04O3wcMQchq015OMiLMPY0DKXr5luwKz8RGFV5j
7pOGHdue+5/6+p0nkbDGO3mNHcjpitnAXaty/pltDNzDPLLKB8F6C1WLs7J4t/uz
9s02ZoVEQjD7nS86cIQgvpsRfkkBagoJj+xRCfnkpUyPCAwbu3sAOiAzNBFWeAVK
cxe1RUM8+7hZo9KKl12u7wmvcTVXb0mRhcsNM4jco1AiFQm49jtYbCtCU5Xmnzcx
djvznpV7VxtcLzGNVzr1FKDsFbybTZGCwNSquTDF8Q0WSVNm3UJwOabbM9R0hbAi
fQtpy0GTENE570DSI96+MHp04X7qGIAwvVyURA9ahBgkXQuDXW5x20JIVVtiHgl0
6MQ+OMExVxYaLydrl/o08ywZnhj5WaesM4DRgY6f1WrU1yKqOCEWuw6xIFpywLYn
6O7rT34s6XxIWQNW1IG1Lt9KGTNFTSpXqHxFH2osOrJR49IqGF4MxhvcHZiIZj/b
2BH9k09Sbq5sfbIb2hNzvmdL6q7TAHb9Ikfazde6PfKwZlG5SsoSekhggabWYMgm
lSsNLDlWJpYO5WfUVYKIaWQ8uy0AZlbX+9ohBddWFdQpquGvjPfPUGNoerh0waVz
53TDU2FusD9XayYWD4A0TDpx+JmVvMZOzTfxumcbX6eWyC1HUCIrbuUq/CoWM+8b
Y8vNGO2+61d/kxd723AJt1xFqvmo3g05mPIR1cOQFVcbqbaB/uN6hzD+MwnSz592
Ws0C379+wmCUU1IRecoFC3xqdUZy2sCnj2V2MwZGIaY7Ta9WWJnncwtIz9J5jaiQ
3afmDxPxDwLZTriZt7n0ei7aztv0BjFkbd2BCr/N9bzX/qKVznQKHi/qknTYKZlS
BpvJmVIU/CeMfOkZoHlOLaO8eIlj0fH/GNsFGNfpHqainWUOFBBL7GmTwx/LbLPE
tBs2alLhP9k5CZe9mNs8eVEFGEIBxFTmhjWBXA/onDSMBAjZ+cXfFGW1gFPxyRIo
qyZjIPn+hVnSLIbGxkmhNyA9UvALz+LX938rTRUvWwS8Px/aPDFDxquIeWdutnMO
MfWXJE4Nk2D2jhkfgDDc/uwPcqnF6mhoNeu93MFlayLOybVGhY9uXWUyHXC0MQrs
k3QCYftv6Os6g92lMKWee0fIMuaMeqf7/e2c6yvvbrgTQrUyXHttfgHCDXQP1bwj
45FbvFrtRREafiW1BfqJirIpXLbjFZ+Fx+8Ky17zQUQEeaEgCgSWsLln/I3eK84X
sRcpc5fHxfKSfgrvDTq9sxHsTTBwqRZ1X/pqbY+LWwUtYS1xdWgUITZPCFM/lAka
7mo2PZuwIsQ94y2TFooiIJ1pNDPKJrFWFobxWHiPYpWPhBinpX1d2xxOC6n8sL/J
OmXyb8UPdAyE9LN6GD64DHMWS+XNFGrwhsMbICFFaDjz4+MtfJzBiyhPZsa9Ci/P
abTOgveG3yyfnObqr/u/m8faBHixb2YO1pJdRAyr0uyBYo6Npn8rU+XTkSDOpbBg
kmzxT3puuG8suqV+eZGAdj5bpZqeyFgXyBMEo42HCtXI3e4W4v4yHK2vlquCUEno
WvpBMwgPBEsnC5DbmsAKt31061ZfxWnXUC9G4J9ZW5C8LbJjHFQoopl1TSyOm6vD
nwikYB0vkdPJvBaeMiIAGXxi3K9WjbzCoHe/ftKjPa3cxcDLMWPDeKvaDWI3J6MF
x6IjXEUrDds94qAGISrY6SNnypONJCJ9Jr3W6kSp+WPeTKugXRHLcSt5JCT70z9Z
+8SYhrv2GNSnEZXqLLQKfROCNqhLa8i7mNGG1QgyjgAsCGpi+uUgQ9GAaxUFTrlW
oGstzk1VbwT0AfeiI4AYOj3FyPQf3AJW0WzjDuAmEKrF/uKUuDxy70RuyfoobwMW
mfCQt11ov1+297W6A1zJJIcjOm1F2uyyFZT7PtSlWB5oJ0njpnzXrzfV3Y5SpD+R
d+t7rVgrr7RPpW6ZZS8EsUrzxXfXlgRgJMKD7YDwo+6/0zwFJtPcb1vIgbfSrqV+
uohEHDaGJe6n+lwd8OxJVw/o16Sm2XXmVgldKXNKy0ItlcKaWhW95F9GScuJQMGw
0Vwpsk0L838XskoOVtTNJFQsH7r0kJoEdHMwJVORMc10s/y5BZrX6fvp3yRaxV5W
7Nr4jA8kGwN5TPKSv/rYEg27ONbp07IwqUa6pt4+hV8pfj0V4Sf2b9edJbwbGB+K
jiDEVB33ZUwp22VBO39PahY/S4U0lkqEYi5wVh17aSbvCpLscAONGLD4pSL8OchZ
HWRknfbnLZ/ymITWq4qq4aHszY36V28J7BchlFD6dUJB2O/BUha69PRBz7cthhQm
Cwdq2hDo924fuqpoJXgf2SXRbO0SLEJIScmCtz5rpFMYlEal12Q8BZGfihw6rUT/
kSIpGoJiY0MVP0Pekdz2GAC1uTnNH4NF09fmu+flwOQAR4Pz0O31NDRqR+5zzS9F
CGB3lmY7rG3GSOoqkDx9rpaZ8cdlDQAlXiTj3JOrLz1TZ53shEQJCIqmwDAn+Wmi
pENB5xrZZq+XUmBw98exBREKEWNZH45YX58aCT2hecZG3kFl/ikcpjJ26RQNvGkw
HxGERSZjzJrnSiSqkVDA0Dkuqx2EGQKLnTU1QNKxuYv9U/DzPPNpOpW4uEIIG0DK
srJ2erP3gdpCXysn1Fc+lBwtLyOdfOpe+It0SlQKYpIWkpKuZ+2z9B1jxgP9nCiw
M6aT7wZL3pztkaf7XKhsMrHkJ1TZycOrB4En6ndvVc+Wr+R+1Mzec3/93mAC9kyc
Vk0LCOMGO2ypo4qg8FC+Ofo1BlqyuKDBM3QI7bR9PS7Of2OV07HBHp5vEaiJeAgh
3AFqO0mEqNuqNF+6BHKVkhKsatdmMKv8kVU/RKPdvQHVdVX0XW2n62DUsmO+BwVt
/QhL3DodDTVvlOo4nAiHxp+PmOKhCl8ZbhahJP6tIqz3fZHDtcV7ki27PbBJM5mE
DJLsEzNzl6X5f8/84pyS86bsKuuhMb1iJJIlMemDSikRYW7sFW5tVbjexTNk1wBm
i6O5Kr7erk7zzQ7AVPcF+/oSyv2CJCIt8rGwpN4/NJePQZFWxY9WGRkGWJLV4OKp
PnklqEheZFaKrWYqFPL3wmtadcfXT7uXuVmkHz3w2oNYo3grcRdHMBKw4wgaSeR5
iTHkAByp5yJKTnXQZz14+fNUUopHM8ZUgaiikb8ojdcGy7QUFKUYIPIFdZY+OlO5
3g0FBSCERoTfks81P/IMQwieKgz0BHTXPxHzLSUGoNRX5qMq5SxKHQtqFfpbv+VO
Vbv7oTzjxB37VlYtnXTBsnv6VwK9d53FjDm8twC4DqpIJV8uCqfcfXB4b6dGHnSw
0h/G4UQx0s3z1ir4JmbSRElHP/6689HN6xu7et9Bf3UblreyigLGNRqeK4igDGck
8AACBnSlmTs30TZxvYHdnP3S1YxRgA9fa9FuJ1abL/tpafdwWErD52vX6+PafssJ
z3YbSaXCX+B9CY09ra2HAk/uSAYt7KZpueujSCmp2ngdCNGj7zddYve8yezkeYTz
228CEk/q3UyDbc+XftiEi79iVsYmpCOjxbI8r1Jt41f7MJHTx/19PitUJrIsM3gy
NZxEVXcrN2fbTAkCsVQkYqCsMd4ECWgFPbn8ZrcPEjP+YHDefG1BlB/2ECTYA/kD
MFwI8GpVgWWQsLToKLT9mInTSGirK3ggxY8MsAt3v1kIk/+3lHsA2Z+ZnTz85K+j
AOXHsva36t++b8mdW5f0g5FYvNzJV7/jMIzrgjQLhlu0VCQM6WH3n9MkRvqgYIQq
OBVXOM1EAtV6YWpHS0EI7gjqG38JGxH9wBB4I1Qqc9dm1/sx2F2sW2wpAI6qFrNP
TbMRg9MM+1avr1iD2Rzykv65Knbdlpu6msoFKq2QBsFXyD+czbcjnbGVyPcbwUFz
mHOtOf6DzTQTjg3POhg/GWDJkWyqHaUB9KcoodPYEjAVpZ0h2HK4quQthEq2QTO5
mP2qepxtPRbUiIztLaqkHE10CNVzbQwr9uPSCtWHhcVgLBOqRpAzvnMYwpcQRE3n
Yqy2Z51PmX8tMVlFJWRfFLFuHn/evX4InPacMNm3YDk8WM0aMHb70tN768t4ZIb7
ltmmacXdEAw0f56V2o9AUr63VZ1A1Utoq6C2jKAbidLaexgx9fXoOTneEfQyFmDH
FB6eIRv6aRoS+QkJnqwfNyeWawQfIW4COTWBMTORMv3edhywkQYB3P12gTJLK/k8
R1yetOKynC49nd85g5lnS/wzn2zyIh36Lv0AXWyNie0FsNUPWrnUSc9gz0fuJNFu
byGRZdSBNJAMEkq80aFYKpYdSqaiNDCpgce5OSRpYqJdauqcRTUtnti9nEJRYeA5
OwYQKwRYlrGCf07ig10Abc4b2NZ18srOqFOcNJX14VHLTm4qcdeVe2Wstm6iy2Uz
IijGz3b9KsuTyxI9PYSHcDTBVzQJMq9XqND5pA8dp0miCOZ77XWfnKyk/X+9Uf8K
b37euXLZpeS+yzViKPpWOIbhpkoZRkzvMwV63vrTfLPlmpfhwb5kf8Rhg+ODOLtP
UAM1kUtURDBC3/zbPf1cN4NDlPgfyjrbqjNldE+rQsMFJneZbkr9b1q70oQBxmH4
P+UtJug5n1jqioVD1KyU//PRVj1X/ZuHLXIcHoD1AX+Gs0sR8SSqgqpespfDd9C9
sYxb74DVWAti5xElva2LnL6AX000QDasVK8oxh7S1y30s3TNV6vhzMO0MgvGxhMl
CKY0eMVuRQi1HZS+w1Eu1lTJKvBL87j0pJyedLh97DMOqXY+b210pRorR301PBK5
FuLcbR28RY+xeHPtw3yaHb1lzpFwj2lET/9EHRKhpv3VOKIvGg+WjmQ8BWfmJqEw
YjiEQjhPmZV0qncAIvz8uSbNhZAniWLwEJqe/ie4jOLO9PQ2oZdfNgxEap4BT8Ox
VQvKyrDmjJIM2zcyZot7xS5td1HZnzd5Pq7t3dmXpC2beeytq+bIJthP7INiAaCK
0oG1vsZC3rS+X7RQbw/3t06GASkUWhq0kOYfXBN0F7FkkPPROPUgJNCC31ZZoBkw
QNCPlaflS6Rc9cUzyP6BMcUtCNi1oJs7Lxvj/kfuQRyalzmzM+YjwTLDfG1SCRbo
ZqCK6qdit55o/EgNoMIC3yrEPq9pcQHqCCDkdJobMPOmYUYngc58jrjOqdBkbaA+
IXwgJMDlDAKJstt7TUtB+TOiNbHMu9PWgZOlzpNtMwolgZM8h+GAs8Gt/PSIJVdu
Vym28IYdOsIwh4haZS+Jma5UegwHweYqf9JAgmOByUm9vRB4mez6A/n5wlLzLCdS
9hHMp7vPQaSpMvLwH3r0sdBvQRwKIo+4ShqciWvh5Ey25Rk0swbrPa0u6th+7NJm
TOMZBIwSo8CFBpx6rx99oXggUM0Tu+QwNU8bEfADDmBWDKmhNqsQOG3WQVr86Va5
VOaww+t7AEloPlpKotJySuG0BNPaxW1ovm2W79y7AX+77woLuoq7bswI0ri/RDos
Mych1bwazzrXl4wmaYtOarGamFkLAKRAgSyy70AE43Xnxyhxv12wPFCERa5w8/Hk
XgQYuMeLLODykudaVWqEJ1AhUokZRLJf9JxcDypJnQzCpYZDpw++6HxRkkVchcsq
6xA6CK8dgKg234dIL7AEQt1M122s3MF0t934j+2JUd7lKM2eaLEjwTdSMeWp+1n1
mhewwDQuyW4lvPSM69028bIeJD0SiepzU7JpbQHnNZpxoknouvX6z5ZD8NvbrhGk
dIuEzbZO18b40pp7RqCdT/Rn5sHOrkfgPQOOkJE7cYsU1iFCjSCCOd/OsWzTfTVV
Zgcf2jQ4deJhy3ekDVU+ZH/aN1s6pfYMZ1gjXp5n5BJLTNt31li0X+KTI25vngSk
8kh+ZRzh73eE3ms8QRLCaQSU8zJh1D6iJuck8JEEQBtzdCG8SVl1gvovj/T/WTux
bKboxMYuOPj60GHobpfP22XwHDgV+G5Gm+YuYqVs9v3tIYcWUAtjQNXUJAKnMTYJ
7ImO0WNbvowRB/zxXSmVxqICepRysiFsE9bx4aOdLbtrQ70SDI5Z1X+TUwLI5yYX
JXL62slhN3ClB+eWtklaswd4TksLYwM/sLDKzYrBEeRNJa1TPFSC77n3UMi1Eb7d
KtqdMd5EEfXahat6kTcLscoU6pPaipPoLhMx0Ksv8I/jeW77rGTOJVtJwRx4UgYo
BOCq+2fgvw8qjdVJOUKTsrDZzR9m9CvC5QQp7zJ65xNRztaT///I7u8SNU6CrF50
CMnz1q8Gq+2jRRL7vq9KbAR30QzCZ9+0hybomMcaqG6WTEG1i4p4502TNgB6hY6K
Z0flAErUKeESiVK58HMU6kTn1uf4Ua54UtyK4J25wewya1gYEEOZxt6U4Gl88MgJ
YVZWaRejaxb0RU6X+zX8w6K7o/dgMxNFJOCDlCRn9qS++r3dz1xlVbRVsAeT+AIE
FKgd9bi7xawll5d46vwcJLke1+kL0oMzG5DNmmyPus/ReFuYI0IX40K6pE05QT/T
VyLio1Q+OVBdz3nTU0tgo0ftOKlCrcLWjkNuk1bTGGkEF7YbhSrlg0TATxbRb+Uc
evg8Q1KEG5TlnzK8brxeng7ywOGbYjYCqaHmpTu5Bwkr+ZNAunQpjMVXwJCVeFkv
0syi3wB5XEw7NAnyC80n5oVXKmfKUt8EcnRSEGpwf1+zoU04v9R4ujNMOxulDJ0s
/2xhQ5rEAqxdh8nz3llQVffa8PxloH1gKsQiImCe+RYj0ECX2s/KyFoCTnyGaBx/
CRLGExNQyaQjG6IA7lmiAZHeNPUAC5XpgZd6ru3xMacD4wKzUeSUU304Qkr3zdUS
V1/dtEn1yuK3rdsdYrVRPNzwb7CJDgQE+W8We+rVdCeGcUaAicxLBhlJWqsiVxzV
rWZ8UFqXYxHazbQO/p40lYZII8jcM5I4ocGilxXayTdethf6WlLeorJWkgaacAlN
vxLbiv6YKLczUkBVKy50WRehHXv5k8NXaMMZPrPTRiT65PfXa7unGpROpsQGH6yE
vrlVHGY4YkfDAXuHr6vv/RA85lm+8tkqZF8LUhanSzWvi1TKLznqwS9RDLp0V4mB
Df7ECkP3VdByDDv5DbUiVu/lrReYb7zfW4ff2QY3rCz8mUxs46t/afnWW2PxkFNo
vWIb6hqtUb1vD6Og1xKmGXdJf82u2Zu3sQonSrzYXP3i5+EhrnXo7OaUpHXiYxW7
scxteqtcevNrhSXFZ9yNt220rrAO+PBAC5GVBxshgbDHZN0tIbUmj0vZQnqj3gjp
YLEk7EWlSikccXy9NnBvuMFwHVRX5hWcALcxa8d+/xfB03kauE91TJuBCf4r89Rc
lliak5Dk2zmk9+z+CIhJr97ZxQVo9WTjRBqNemrjbRKuU3Z3BAPi/6CkmGOXOKza
JBPEjekLXaYA7kfMsv1e8152jk3k82yG7rjgoXvaYnDIRpmFl+czCbghUKu+SnNa
Sp/Z+6h7VlueonLVDyoWCLmr0caK/2s4Mz30jrV1qnjcbS8MElolMFfWanFZ6/Nu
BwXZBJ6SGZB/f1lOtTR/beQBPnLdjJ6BAxzLYCkUUveOA1klddr7iX2DZsCjKwec
kfzZUCNXh118Ztwvw/DUILkhOVtc4CGTrqSqmTI7ti4jpp8X0rXXKC8+aJw0hjmP
VKPKRyF7YAlMaDjnhRap60ZwUWyu0Vd0vqDKt6kJIfZQgiN9lPATDQ3vMrVR949F
j2K0PKrbM0Xo9o3xYNh12H27Q3JR7wBlvhA2Bp/OGq+W5kxgVTOR1jXmHakDBqRD
23zWFOTObPGRtSs8BX/X0Oz43cznOrFn/I16lLGwkwY1JKBpzpO/EEJA+9Xseh2n
vkoyFZ9Qj9/gXjoYfmUGuPw/RPaayy/ghqcK87qE//BsaSEuOFyliND9Pl7dTDB8
piYQoHwa7nNz0t7wWAR3nVmK8T1qZbPbEMpo0AYpeSq8ojhNV5oh+3ILfSiLqZRu
yGirSiUlFGDMGn9Z+TFusiKZa8XNVchuyl56bmQRy5pP9p/QT2UlSMCE02urTN53
JL0GuBLrdCmubASYwaYSfsahRT09DumRpdskk/nleXf9axZ/QbkIVWb8TSawr4cs
R1z+UTMJew8N4eDPL49DZOesR3R0UIck+zZqy5z1DheDbrnaIg5xIHx6uKZOmiAG
aPCbaR9+UoxSqA4LFViNddKQV2clO9DhvPVNNd0OXCuo/Z5zxkN67qPv4RrMFq6e
p5/DYTz/NZ+ihXmzQqP+WAUmMTlnBh56x3yMOLU8WQDhJccmZRSwHCa/2FIvsWjk
FlS3IJlbQsCxTkWHfIrQ9psIFvuOqyXUY6XXRZwDURqdQJNL1933cqFt612B7c9H
+LHzLzKC8gvMYpIS9hSAtdAGmBaNHhaErvLJhJUML/qTKMm06/aTnINotJ0YN4BL
kjLHGt322Zzh25flHW5IqPd4j6Zh5hMSDmBFygT7/zl5KCyP4HNmV5Z2CqwW8jxr
nv9B7GGN+aFeydG/dCmwcB086TUjyZvJ8mq0gJqmNgTGys0BCFScpHhk6bOOlzs0
Dk+yMCo0Rrp94XX0KPjyjArkHSrj1f4rC5Yb85L3xAdqNuIDjOP15fqfD8p9ixMh
FkbGByyg5T3Y1wbaLnfzZ9gATgMyAayv6HnefIWbpU0waNJUygEZ8acBTFBElgUh
z2iGXU+tg+j7W2lAqH6nFhrcq5rY2SjRzTc9a2SD0uUniJBtcgZDr5ikuSTPvrW6
YfCIOe5McUrk+FXN0Gd68NeIKzIoh0lFT6D4PHwLDdneYbAaQopj0YaCp6JHa0l+
m0igfmyeCwgdGy1Gyk8pSodvzJw3swZna2Sp280LEhs1Ak7VvgUGX5qg97B6Gwi8
jWI0ZMrmi2xxMffQIylhfwF8JW5vMLUzrNruksX/6JEIB7Wet9YjofICpYTiXFBE
iIgV0VZOcJSav4Dho5GSs6GcRl3Y+mtmk41bIa+qz3QZZ37DgpoMLK7nuLGnodoM
iyRjUtlpBPO95g3Mzvsx9R28Z2u0z/NyX9h6gTUsi/4toRYou3C8upmFu1MdNvDa
0Xm/D/kAdNWUMRhU1x/QHw9smI5nu1OCl/DB+wStbTPs/qoV7HsTJvMLuqZB1xx0
BftY4PqFuEAf67iL5vu/UJIevWkvZ/bCN8LL2sUWH+UDM7K6ZQiy2bRbFIPxH63U
EViR9JYTDhg7R9ewN451FgGFxBMidte2pb1P8yXHe/2he/iYQKKI7WkEhTnsWdwK
LJEZSPzDu6G++JSQ9Wqg5EFRejxPuk4FlxQXjrGQlzTdHoBwIlhq1UGbytfgOT20
ZDYZNCLCJ9qYS1/S5gGCrGFHSIKcDtDh9N2vgjri1ncSkcx4skfLfy7SL0VYft3Z
OPmPkt6oQYjKRmIcHtvcF9NDh+PWPQZYy3vajzXM+NoarbvT4Kc68ksrc4sRJsXS
WsYcMsf6KDQEI8dG8zCil5CsOmaW0T6B1ouvLX6w4O9VT6kJZ8UU0XBp2TTBp4YA
sei/PUG0pQVAYINqtEa2ukm/w8SfKQ93krmdsNWR+18HxJVrC2Guu9pI9AOxtvqE
QCax44TxmMFie4rqrkWPcVw+IDWDMZQWqEn8EK7MLR+vbZeYOs6J5dKCR/fMh9lG
t7n2LlapOUaITPebLvSiFwfqJ/Nrk+XjU3Kb1rD3FVTcv5Z2Rhop0GZy59ddnmC9
69Vfks3ridc07y2AcCiFW5HK3Yp+giKMQKAsD/6HtrZmPaMv7znfq6zEZ6ED0aM7
Bk6xq7Kru+r+c3C/89Qp2ixydH1Nrb0Lw4pyjlsrMNP8VxdAQtkGlKvJ87J6hcHI
1+A643HJCMGgiCsajUh7DuopLyQwltw9deBMKJzniHhkJd9Zy0fGAiZmnZ2YEhKQ
e/uXxv0g9aLlVumMy3mOAc4nse0BTdNp/yEI41HTtK5WvQI4eKpEFGjKz7w/iCaE
9iShPddwmxfYnXXP8/oI3jXoRIAlVyfMtE/lzUnOrVmCf8GPtvTiRXS0U4kVTy47
7/4Iz3eFsRaZdYHF0o/7GV3pM5SJ2xdwP3tsITYciEG/dPD8fKNQeldapkmNLCXz
pXn5MkRrJBmU8MWzJopSwogXcA4cZ5/A2KscseO9hyP+4I5Vy6kYWQ+jWPSDUm51
EVbjJ5H26EZiX6uUwYtjGIBkAU+srDV7K1djjYJVMzsKrJDGPB88M4fOllliXxQP
M7J8rzuIp/0c+vaYEjY2haainZobg1ZAjAe/zTYEnQ1cApq5/HAeKfy8jL7/iR0G
0AzTn51vPfKGFGLGC9xYDxhqycw+SgNcZzos5HZpHONXahCv9KjnIcWhOHVqFjgU
Cj1cz3E/6gCeQ9UcNqGMoeeUq51emhNpACzPplr2912qVPJw+FKzpX840UjIdbJg
4GZFD3A+sCiHHNaQpDsRyZXOyUPZTnbZxQoq/tBP+CkQTVBoHXvHZN5RH9/dv2bK
+qycw04W9FX8dAmRnNWzeku0apOGoxNOLKVe3ye25uSRbjyPm4UGjl0zN0kgIIiU
ER2kvfLfsT/mN8V5DcbzSubVnz6UQualW1irOFSFqNcNmEHYk8bZQRv8Q4blYLNO
0sPxvB7BNN3vRUf9gjhhaiUGYe6Fa8Kl36k8qEyK03ylQUv0MWBJHJH9wWzNNJPs
FCxsh8OiolH3qjPNA8f8OfXQAUmKlQ+lAoxI19v/KzbAST7S5Lqs00yB8ZMD4drM
3gnmqq8uYtKowRCHmLsu/DdIZfIvlTNf/lDxeYF9GAV21bzBwrbgpbQ64cdv+XMM
j1RqYtLhoTlrfE4uu/UnoMNqZ51c3scg6A0dEWPkxoB2F8bs0S1cNQ+9ojj/HkKJ
d1GgL6vs6W3uLf2U42oXmSgNr3mJ+iP9ImbNwZE3O8FQHXhnXMblpi3b03NokX21
HhlYyfQvpoWaLnv2PiPRD+vmThdZPISHppfIoQCpCSgDZFGeXQPOxieRA+fJfNxm
SRUEts2k7FyXQzejH3YOe8WpPKSVOGiXfWYymKdJF1IPUaF0r67dvXXVBUCPbEbw
5usC9lQ98NVanaiPo0QIHrRvJcWpiWO1XEfuVM1IQ8mYymeLV5H6oCrp6jxBetfs
LEsDF9ucB2NCBzR6YYgawyzaMUtGAvf0HmGZU2EJB+7Vped6VeewFVay03IaHY7k
ilSA1+s3Kdy7jNCOlSK5OCY59rP3hkt3pv8SC2Gb7UyC+3NhLaUlFFMqzNLLy5IS
BdudDJBH0izhtnYo5gWwHLRKtpSCYgQdHWsuXm+mrHLkbQWXsU9PFhR1+Ae+wdu6
K9tI7JQ5cgCiqBESHbSkxphEmzed/6v/Xr7Rjwcx5YmDuH6e4Xpn8vOuNN4WBHyj
FJMflF3IPlZ7FcVWu7cXG4EP3HIc/6yS9hXzcYP5skYgD27JhYnfyKHwyAhO8n3O
70no9HhiMpdmg9B0NuHdWaZpZ6iZFF/EWsFFg43UA1puVb+NUq2ZqpTk5LbGVGNE
e21iwG08zCDvCjrWlvMM0fJfreYHp0qC8B/21oLrBRNwg2a6UDO2CDIL/wz9XmyL
36/7n2Bl26Dxca9FOmsnRqNkJi/df3cZNoDWdbn506GPcrgDg/ZJiAkUg3bjf/ct
tO2P/V6gsOeAFFEeywl/hw2OC2VoMM8AcyqlCp7vjhpHJTTjn3EKYukkgzWanU3U
3+strfqD8X1wFIxNmgIUjnNC5L8LWyBC2EAzOTXNVsQNIP63lNkNlx1v20vj2Knv
1IV81CyycxOXE1zGN7ghVBesaoNRcSWxnZLvM+ZzFLySZntg2ng9dX3YWwb7H4+3
KATjRAGvd87t9OejEOcVLrGC5JcsMKmPcgFbyBNafq2cWfN8KANa1cHl64bjhkUA
kqAIuZolaKQcx5S+xjCx6GY8M1vIPTsgchZxpRt3gDCQrReNTCsxCELhdt4n+Uc+
w3hckK/gkCPazH6P3H++ZZE8FOpZuMXWxTAXoaLfJl4GJRhvh0cR2oXwq/pvaJJ9
ENMW3SBX7n+/9mP060DW3nd0g5LayeN7rDvxHNiSc8UiHSc62dGRchzHq15mIUDK
zfjpQPukSI9gW/pyeBCPeumAMOTBXDqhwYot8+8OfFuDjJ3wI55T3HAZHMGOhC/l
EWuADdG+jZHEmuxDK1qbJ7gkk6BjxepOqqvh8kAmO235gheON0N6uuuXQz9IepxG
z7MJlr4OlDXS+RoFOAodjfpYZUmu1CAgsCv0zVgd7WXggxLGm6LzMB6YPNKm0c6H
SHpNSqcvRykbZ2H3LHop1sLyY5S2JI+3u3FR6pfVFMyws8RF2X+tWIIqM1pwmnGP
fIXJOi2KHXL/aehyrV14avSQpew8+sa/pbjkRBiuL6VkgqSHuFk1qblBbvrTHd6X
I0DCKGp1OJmbNcwtt2cLnoJBMkOxbR7AYaCNzaSZGsePZdz72GqzHfNw53CVXOe7
sQ19swFQz501+ifJ+s4SNL273VmwoHWBHG8joB4yAl4fkUV6yvLif5g5YNl81TB6
18H4FFX7KRBtnqA5Hai14HmRV8uYI4AsB5F/gQjK0LhCw7d0KJKFE1IFt84whbbm
/xAlo5ePuyDJmSfE02ehyKOpM+EyX4N2eBjwOkre1yetCg2cYlotZMN9i9UdnoiK
HMtwqDVJocxOB57drqkvuaYpsApsAAlkztxTZ2HMIoQV9lggjyW0RgUyF34RnfQC
sCh+JsJCnw4Om2skKNsL5wTnga23qn4W+dPvvS7kpCEXFxbwQtt9AKnm9IT5h+zG
zQfpNZhdfPeSiSUBOCtTs+3DvJckcQCyWL+xije04cr1/dO6LtfRN1NYrS0UdbY/
OOpxOymlTyWU15t3+iFHqJWQnroZfKGTTaWEV8fHCvMQqw7vnOYIJyOgmxuuDLat
pHClG4mbGpJtoAnKsvwvIfYt1E6VAsg3gl2N9Lm/SXYAwo0p4TiGtWJ/hEvC6XmI
gPi04vt+hf2OjMO/S9FeBncW01gj6MuBt2+MReYWmgopVznjEStnhHkqBPuSztyd
b09FNhfzYitXO6gvknriT18p0GUuvor8fdEg253mj177TVWsuKnTyVznCRHAddQq
nrJlP3tXsEotPiLUSXN0PEt1BwWVJ1e+0cwJqh0x4HzqQWiijPPoCHBdaqMNyAlj
x2kqIASiw+3/WKbwrLN1WPby8Q8XIZ7R+M6wiOlj7YHN8filn0svGBYHzQTClQdZ
cp0zx5Xxpx88EfeFbAchfJxZEeqZ8RN7yWFJ8bPvE5TkoB/wO5AV5f0le+NkYWhc
Q32dPTzJRjzGrxrEUBKlRAJ2yElnMtOrjyfKf0PQJY25I8N0/tSiQ308vTYaCui4
lOeYet3UBiOpSfbDWNYtFkIetvZqDXZzPAWq8fqvTn/NrAolRm5EwTSL7dCrQF5w
5EFVQZJIOA0e1NfprBQO523RHrD2x52OjvxcnKWrLYq5vyulF/IY1riNaasUSy1k
n201He3XP2juGbZL98xD739yCt25D56nI0zQ0gaOTVcoRPedrfX3KgBeq79kTwq8
p6POh15jRFrnjYntA4tuvxM8Zem0cPPDdoE7aPdd/w6SkHFSoPW8hfgNfKQHo74o
LkVKERLn4uCvwMF3HZXn1WSFczEnH45jjqn2AdhqpxDcrEqHjXsbvzIhpzNJlSai
gvGptRpM+ff34pgtGn1puQWD2urlWAD+dyrDaZVKkfGHHwwNP8ACFdfhveuPUYcy
prlRZ5cNYRazT+d6g4/4JDTUhxjq22yno7zy3XuD3H+Tsl6ldhyU5fSE/pX3TzOx
O5czi39Htrx9n96DltNsb+ysjHN1Kr6HuHY8s6h9bH8m0pYi2TSMvcuEe/qDNR5G
OekQsGhefVwfueQBGE96dc/Nh8aMd31ja1XFkIpx5aBNuQCnp1u23tkKv06z8xLL
3HDOB9dF3aKrt5q9QLh7pYWxXNOY976Zg+YKSuPRKLeJ6M+vIX5Mcpn4xIHj/05o
vziuvlBok0A1jVwUZaX01u7tvIqzb6bhIgk+kBby1NpCEA+tEQHEL7oEUbX57a51
kNFVNZJ8JijBJU2JmCJIodyNwZBtD5/KGLurKtZEuANzpQIYoL18JM5U32OlN+w/
8CDgxVW2rnhBXxLUA8rzyWZ9Ho7Ju0oIgedvlbDLbi+54RiVmzPLeYhlVT/UimF6
KhWoeRIatIk4xB0DBS2uU7/x8u8+ZRy28j6ldIDg1Sv84TzFP9rJp29LDZiQp7j0
ayhMAIFGLKW4UrrS0STyIj+pwKT7Mf2d6WXQsfK3ZTDZFNnyRK+Xr1NqyrSqhDBr
OcG5BjB0l2igZNZnSRwwmEA+nBEFMq2Kz1sjBZZZaJfsWg5qCGL3J97Rj1t/goxc
fnAQ2Ra83CKbQiCofAit7REutW8CCJWOifFuD+azTJ51ykK/FK4ncqfqvJRYbAUs
dHn/zMatfW+cGU6Qy/Z2pSMAnV9HdvvV7ZDVkjdoX4HEKRrnepg/MOkQthlntFfv
nJdLK3btmE2Oe8N8KuSBUkVoDLuIFXU4QXPDeqvvng2uieyQygdrR80q8RJHzAPO
HQ0AI+79nwbO7H8YSPcEsjjM/qWqt4q/4elYu6ZcNsvIoEZt9up3EkEIpYddxyD6
P2QQjbP81L5KSyPxCbM3zcDG9eZQ14Wc8Ub0Oj6NGkIBJWdOsQiUaYWD3sjPpzhY
uURl6YXRVLjV3X7jXGT9GlFf+h9HgqZVOx1lZRd3cgDbRttjWzMMwKmVcIq4AagI
qnrVmnmIRpabtWp39z2Vkr1pGeXTLH2SgssUOwTjVLp+cO+wPB9XjQbWkVjZYPsg
ULvwe/iaGrUDuTRHKttny6iYHVo0SqCFyxf0kKRAxKetveI5VmTIgK9Dg/AsSA1W
4Z0ZzhMlpnendChomWBlf5aEFiUz44fslt+2JEDGR+l4dQzDaHuV7bh1+LQvQYnl
LIvP8a/3BuvAo5cnhlhDH2IhXcMBnQqmvXhOm5a7Cud5is2R4bZOBY1oKZhdslvk
Ha9h3IeLumWEc9T8ujn4Z5GeRTdgvGKDKnmOI0lf5SmR43+R2VBYY+Nvn29+dotJ
zhi4z3bfvkzYTKts3fSibzeAcKLihfKanKwwGvgoERDkZjWCAgVft7IF/z6QzXgo
4s3Sia6mUBWQYZMrIGqHKpT48m6PKexP72ah2KUkIR25asWYN0itOBG9cH03wupt
MrlchPy4/d9v1cUzp1smbGPY/luionk3fiNb40fnK2VuCRdnc/adDIO0+lRswI2b
D6CyqB03qbSM4WMl1Swe9VWq/eZaaSVdtQKvU5+bt5w4vphyyWKyavzZEJuXHYs9
qH2P1QPJVxXZng5q0EFe2RAFWFPO7mhhPxY+y6OLewlEBI05JMFtkX7yHPBPCJbQ
MyIM9MK5d33EFDuoCHPVJiw+JtvMXQWAInEnIsBEz2sS7Nyy+yGGdZee1/ojv8K/
+Qm3+aMTYE3PZN5Ah6Ug8ZqzhmOfk6tM3hP+AqS6/ogxfjGyA6UoZB+F4OSLpqAX
tPnuE6pvHWMCyzXHmbnr9BQBPmfa3ZztWnVklmysVHpcczp6hTlv/yeb7vONS8U/
X6J6hSJuXAFthlUehe7zfwv/F7dNgBuTtMf/N+Pg44iwZJj+VLinqgdIH6gkBTrJ
Nmw6fe+nzUxi3NfT587fS8OYzoDzzMqe9a/mL5aMNvPTV4fPiG9qtZlJiGuitiul
4vSAAIRkmLP/wyFO9QBGit4O9akMfkA4OIQRUmYvau7V0qb7c+iwrUvbHaSZPA7K
6aplfy7U75REMfrWvFEe6UCp7olIlWk8kMS4Jva/k5BC6EVIj8yHoi+F/wP1nhDU
MKr6nO6CPoOw7M2tcuC12+AwPU6EjuuqyMTi69wCCarR89xOLUoVmZhTli19ocnk
Y+hmqq2nui1hnORwmk4/BS401vi4YgPsQPhHwoD66LN5okZYviouttNrkFyAFWT8
5JI3fb0jYsyu1MGDNUUH/GuNZO2pM2duD0Sp1yrwwA90qT3nsAB91EeIXTLcRO5P
yxhwhnpgTQFL0MhmQ14tDpEYCYllK3M/KJlu6UKYzwMwSk7lCob7rlJseYdAJQcS
zRRrQ59KvxCKe4bYSa+PSn4iSi56Rf4/ITHg1DEl1Sg3oSM/V1QcsdRxOr96NHbq
le5yLAz0SUs75oqMhc2bfQaRBf9oS/mgl1UJBcLg9HUOPc5XIM8T5cC9t9Mm9yVa
l8F8b7ZA7mVRGSd+Dckov2UWo/3AhkeBbEyDBxHL9JnFS+3rKYQ8uWjihSx7vDLU
za6kOuLYUiibOrUfv1goq89OsVLuKWDZnRkudgEmg95bOLzdlnexnIsquRP3mCxc
ugMcwdfFZjETYnwru/kKvokt/AGnhFJU9hVhPPQX5ZaaEsAMq/Y/Xpx/gpWHGDxT
IP7Lsjyurnq8lcm1wpyZZTtP9s6erL4brSTcemdZK8ztJbhjLCzd4wuZkx4oI8hS
bsWfjp+qZoLzoLwcn+Jce7n4URHY//2/iz77P4HRexMMjkuAb5xfnTjJ0dDWNnme
am4lqUEdV7QS/dV1T1hCWq52vFdDTxBG6nZfSjuwY/55hwjRZZ02LYa7nRlYixeP
SdAzgK5NUWexAZ4RPz+Oo/VbCic0KWZ0b/qZSW3aU63c0qXP3V5stVfBI1IFMrOg
qMbaJKCEJBfL5aofRlhC3xkFJYX+s5lxBlgRwJVm44jHujSBRwpgQHq9UDw0f2MY
Aan+HgL7dhWRegHcx/j9cw7v/shEY9d/MsiNKWv5MVXYtX3JivoBJo6/3Mv5yzdg
s7NHbCKT5LxZY6sW2kTIy6sH9Quus+02E00oNIdSy671Da4RfYK5WzOxurcqTJGe
3KJOAgaPHrjOzVdocq9X+UTlJldknH5D4aJ9TbyqF1le+idtiJ58v7lZXnStlcjU
RvqyD6pdSANqj5pvYfGkAspazHmFAUPg9qm4T8RlRSI0sDTWDTEQymbz78ZQ32/h
DW9LHgcfz9c7v7noVjYQIq7ETTZ2leHiEV58g9/XEbVntp9jRwuBz2WwRoH6AAxr
+3+LgvWXNEmOez/u9vVgYkgw9a94mprvu/9s7iHHg+uXtc6TEdb6RNZRhhcsAruc
o0vQPFIVM9BS+1votEN0X4Ydpxb5trNG1rcTA/1AUhlPDhP96JBzajDwqSeTXl4O
AkZQEir1pKMUBLKrqWimx/D5+Ia1VD9yzZX2L8ifRubJha7H6aVQCvkHGQL8K1ar
EYb+7OQRnAXhmfTHia7mr7FY1qy7Iw1j5kgIpkIL66NG9+2fVRBPYL2gkX79pcqH
RhP9dn407rBzRNTTI6S7Y7ZtLILWqhRygg9caywWN5Zsvdp/nkZdXiO51j8Nkcwd
9TjmOWMp5xnXhj8X3rHNIm8W8YZnonDeihxdhyIcbSHYKSoIYBNGvVvc+usBoIzs
L9VlgujXtTjj/toHn8nUE8afHEjBMfxL4ulCpJJ+kpN34Haa1usSjvFzQ9tYuepJ
nz2o7Ej+MrvKnsKnGVRAaObbntE7KeHFrEBRjscM4sQpGa5mw23bV6ITE+XAa9OU
9Nd+XMs0VDkJDYn0PUg/4VrmlCFMWO3Q6ygol6XSBebp9ZA0AwWjJ3QX8mtJV1TG
5E/vd7w6Q5AmLSNDKPQNrQ4cANhYnvyJG8scE9P8c/BIRJZ4HLRu/g5SIqFY+XCf
SIDslbWcOzmsZwPZcA/RKq3FGrhJOpho/phFNBIzY8IYSZds1s6oHS8CR08ryb8P
Nt2qJbJOS1YAwUg3yLKlyPqKDfaAWkv3fe7NtwrLY/ZDGQquaQ3sLoeE7MFet/lb
izXkNcPHfE9jhdJKVbVqWcG7ATKDmKMBuIKA1YZ5FwzZC3ceXHvUEj3CZbQxBX5t
T7y/hvsXOznzy96EkTGZB9sOx5r/VqDeyForwiabsW7ejSSE8mZVenCXoPtIANp3
qGEY28BZGWQNdzozs0GyhZweYzm2VnvYWDsrQieLz1Ls0VdmwUoEVCqmaP3fKPSR
g2umM63Vpc3Cdu6ccuYEQauEbg4LmctHytCc/1CU4jyiExYUc+/OYIw2Iao0L/9N
1dWawMiHT7XX2l5MRbHzSA71A7iO3tpnHSXgOn62QVV6oa6vnFhDRBkKOU6dV/Kh
eeWMA4eGoHhG5hPAgpeSGQJjdaoeeMh4YffOWoxTk7yMMc0H6LNko+bEaKBNh/kE
gekWhomxBdxCmVTaNkBgycMRMANacI1ybH2hcgnywDU6p593wzPKiVJfSN9VoPZw
O/EA6hCnXOlXe4j3tmmSPuktLkbOfq5J5Zb350/VPkklEpTDNnckRhBBxoxX+rq8
X1iDKXSN4j/ViAWkOodN1tbYE5aERVdHPU/jt8HU+z60/f3CCCOxiiKsH4CFD4pe
bmLSey56ce6pyLNzfif+mwU5rH93Da3ecWRt/rUGuHvARNYLu5iQx57TcexHdNnw
YXM5ABz3mDdE83RLr47FJk9/hUeMQMgDOnU51YlScwaHMAdAYSMTZrmGsyj3mS8v
U3lhwVu+1vf70eQALgQTguEpB6j7hxA+oS744c9r6hux4OQ+SvjvfDDKZjvPY/38
dFaDs6KgYIfZgvTFowE0FprnHVTxOMQXTA7p9eemBU8pLC8FTtSSGSlp53MkG8Ur
jo8XsZqY+hcbK2IxtDH7Uie4B1UZbdJuh2M/JaLufSAWzfDMd04ORWEcCVzXhgh4
9CIWtBJfy3YRwncjxjFjVPlSNG85R77ipKpjAcNCxx2+j61WwTNwV9xhdAPYfPzc
aXWtD2jy/k5JywOECYLnM2pJfuqazpaJGZ/JtdBHjiZPSXOSt17kODPXOFOGd18t
OLmgurnelZng+Apd1seqk5LUFlJyg8notzbeCugDlyG9d90xQPgPncbBKu5cnNgu
LceY8o13/ajuaPffa7AvDXQhUElLGStxuipHqOFbAjEU3WLluhgpjBFha0U91y7X
6USvyphDjJe6wRjVgazZfn8roEoA4Jyt3tco5yG5gh89y13Gye/wf4t8cY/lPbfA
NfEV1knd6eEF7NXvNO9S0Kbzf+majK9pqsdd/4I4mtquu18gq0PkLnpp8xZM2Ull
y70MQUInJw0Ar23H8o9thdvKI0axU+JKoq7ZRn/LU1BzhpmGO5EEi7Oj2WMdcpkV
gWSwSG45BaOJkHdFkD6PHM5fIyytXulenJTvuxumX16aJlmoKqCwvF0cSCKLphYu
6YxqweOY93yWNblXcTKYUEmDvLe1huTPqdXVL5I+5GP0cLMlBS9blo5TBcvaxPMT
wdQmeasG6llWcOxXp+CoKoMqSWN1nnSLOfT4iTC69u0PNUKmH44Cdidmkqi2gszx
T1rP8I8Gr1E1vzXj8M3F64vEUUdzTe9jxxN/yUz3WbAVmjYWxCstY6mVXA5PrNlZ
HlYXeLcprP537QtMPUpHnv/Go/DICxRjUTc9XcEwQWIU7ascoKT1gYunPA/k8Bhr
Vr+KtNp6cez4VcVjNDk0tg4gBcDG1DhSX1VphqqbUQiHYYUDKB49IYE8W2LKmYgO
En0908CBjaadRX6GlXUjdY5eji94Mre6i/ZbV4iD9YXOxXJ3Z5ZMAllGbNREsbJy
8A/HftQ0/p5D4nNwMPvONjEBWTyYO55uzQ0MzZfWXKFdGvgfEMcCyUT7cwyyiihn
BkQ9e0JEwhiST0lTvswHz2T+3BVxb1NQ48XGMtEs5uguSOQqdMBSTvveGvscnbR3
7cndWQO2I51acvN3tIJBWxVYW9q84E1n8UAO1FelpGioNMMpnWX4ghVWl5a/pf3Y
lShXvwnO4oMRwaZ+OK7f/sBhzSs1hcn2acQTWnCc2C9lqlt2Y+DJ389oLL/yO6PW
EBQFsIyIOBk4kM5gzGnOGWUmih21BSLYvwmknJXryROfmL8sHP6TMS6HzyEZ8ZfI
35xQxKBRPzU5COKmChY/nAZpnh/iG65vFkNoVRf5hOWEwXUuAiMn2disHvjfyBp0
fgE0TNV6mPqFKJalzUJMAtU2XUJpC4i+2lLIO1hKL3ysPqvPY3vzJFjQeVj/EWzy
9Qend34MkwBoplIYMP+CPiEy/vuj6n5ouzYd9/i54EvZCg0KlX+8GUCRLNK11le1
kvxAkc7POPiBrgIKjYAuwnpC+ArQSYxbxREobAVrqGrt/FVlrHvy8fZl+JXa15gy
0+V+kJWmqJ6CupGb645O13YSJtHLvNQmWHwx3cFVCgzoIPRvXa3wpllUg3Zj2fhL
K2A/YO5aZQN3f3FTMNZxdm5muZVEkpa+eBJSdKeCX2KITjvzXVumXw7otnOoSDoU
Ak+xkwx6PvsyKVGFBFX6HP4omIVh00AL9GfGhM3OIqImrtNlF8H2YxOqE0sXXjBd
S8f9ltBi/VyKtbJAKl9pYHBDv0AfnGs++PpVJiEfHOX43A5TazwJHpRiwMY7QJ9G
u7HQFQ4AlGZxfWkrkMPyNqri/TeAZHkWzTlrQHprVSyGK/vr1WWn0ySDTKIBZnKp
NeGzhwZXmenIHqb++gw2RedAVL4fpKtQbj6TQ9DuKnEs5gHDUNkVm7x17Zos+G42
TBzBWbecPYbeSPR6+9cv9Fi5Y2NNW9BJOmhCWz3eTb05qo16LmrfOVjrY/nSoAFg
CHyQDU+p2RuoloxSUZ3HMbCw3V2ZeR0f6ZxnBvOo5jKeeqJpUe2Bgt2u8RttODwQ
IXSu0pXy3tSnEOSmaurnCpJ/w1dhENCvBMlufG8zkD9x0luBkTE0lh+iBnEtHYQ6
NE5A7mjJs5aZ7kKo8oqqUum8WtZ0Euy43xNA4ciJhFL010jrHPX2M1AkwlCpSz2J
6d8ldmX3tViK9/3gDhiwLLLfmV4MSejaUFaNSqCgaR8yH4GSi136FEn4nhq3rOKo
T38G3JOda3Cw9SqawVIDw43rFdmQwCGs5kJDTc4Lo7WSUS+n9lEXSaVAUepMpcgJ
Yl4vLjmMLFQA5HQ0qFIOjMSzhM4rsk4f4z9nUux1aRWWw/QnGikgmUuf607hneEh
siTzLVjYfh/iMhSYqE4yn4E6zGCmIs4BEV9E4QdWxY8WmwIjTnvOoVz5VP+J9bqp
09th45o40IJGZbbler1mIKhGtNAwEAo9WzHAvv7i9IxnrMT50GS2mCilWrCr4tVy
WdyCe3I+EcdB0xMC4q4ZrIWniTY5qPqSvkdQnKlueAxj2MU7K8Tgp7+ybsxZlHuB
uz2fZvNxBSGC9Aju6kFeaDfvJlAIu52ZPgTDxpj4l0AxFeSTdEWZVo9QajkyrnOK
VIHwqzfs6iOaVKbwbn9cFXbSDx/rqOVhOskH2PMSAr2HGZnVTiHaWhMx8EIaq3oi
RZ8HSOut9aGpYJgEShDPlir7vPOVbmCdRPzy05jKMMyIhF1UD/xmQchYt9Pq6OIo
lpvE7jRtozsYfoQXcs/ExObUj+32KWHxVvxiLlVwuM/N8dKmHIuWXJCnNwI0LbNh
heqbMbvlEck5cWaxHubyMWF8Bii5s0rQhcfVjNJrryY6Zzrh6olN8bySLXUQRVin
GbMfe/kqFHVdfeM3rrA6V6sLRxwu/Rf170v5es0XDVCUTSrqUCNaSAzPs4l+59yO
YcU2mu7oWBezZPEqLA6AClB41om/IouiRvXapVqLf0tOj1j5XI+vdef60LrpqV3r
ROOXQ50HwqXbfLmLXuzf8+5SBFZ2ODdPnDFOXzTjwswfq4CeDNqqGTWLcani96BJ
btxIE4lLmLMQEeDrlRIvFhBRgPU5VDISNV+JtWEdvAt5/jPz7Mpk439X92DBD/6d
YjjxEoQzct2hIWiK6HHWQUATaiZhocmVR5noqeSqj0nm0rXHBaJPjq7MzcezHs0F
pQE9WX2KprhtZlIu35OUHwPxeqTBM3Q9OLZtJv3KEBQJjoTF8XdoUBIgHKfkAsAj
a+SKvV/DkUQh8hMKbSrNq+d4AlpPLmUs9JmOgkPgVNiRRZlR73S0vhodfoeDrvmt
oNz78i53uIrGFCDptAWshn9iaJnAeawSgjflo6q6A8Y4DT76J4jh+NrXSKkDgVXz
1Rry7AEJvEeJgU8CmWqxoUMr+f30+kJnigTjYJCQeHeOzjBohqXqKhy6w315C3D5
wW+C+V2CK5VfNIRazqwauJ+PYXOgixfaVMbIJVY3WwBT4eKCSRRdreJMMsnmXoq5
qEzvH2KB0ceuvd78pBPz+6E6KkVCuin/P9BD7gRcIZ1+CJfSIoNoMEHgavEr7tnc
1y5IptLqM/koHW7yUk5rZ7Ia7vp0KBi13hSbaxpwbGLyQ2tjTVFJ2NrYaqT0BgV3
4aQkq1poW9sTRFVXRqgua3n2Uz0orCTqXF6YrcLJZAcjgwA7ANiPRvjlO7C4X+Eu
8MOPX+Nwm9mwxMCUww+oJG1rG/+rQX3UQZuP5PslpFnlIqpW4nwWsW69QY95xrBE
UB3qwHZ4QCXrDgi7zK72D9iR8ivKjLU7V1Xr8vEMSwb8sZObTwj/242w6xOm0ePq
8Sc4DkYlhOzY4OcsjYVV8fXZ/lIJ5CLNcZLWVMSgbDgudMfRO7wnvT5ls5smrYlC
liHsG0ToJMAWvPwTWQgnRmOdv57tQt/MO/yY9KMdb5rBVH5IbflDCD8Jpcnv0Tsx
1qS1uBrHlHOW7gtfBEzGNa94rPwiLMcP1AFjPU32xZId1pd0L1CW8u0v24401syl
Y+evE3uwvRGm/WtcbgjKHOq5JALbtEemg0CVCPpLzbzD1JyNUl3owhVSc52BYd07
Sb7PKRBOeHToEWhk1yh9ye6IRN6YnNyziyLizLAhlyfv6DwKJSszHdL3bxDHYJve
T5pR9Qcairv/Jm4kNsy+zi6kJs6iKdVUjzXZfD7lPKmr1EMw5qLzeaQTFoslV3Gq
gYCzrH9eN23M5/6SH3OShA+0F+o96pxxwmiKvTbR7FnPuA0Q3czRtkipNGMCnTQN
DPq0WzLS5VUbRNeOyFXvXqlqOcE4F3NHHI7D1N+vR4PsCTCvWuUv7eiTKVv3F0hT
J7VUY9Z8O5DuayPntoRGXsFIQ8bUvOtJsbukX+gaP07TpdUt7TR3kstXvZYQpj89
NZoIV+GRcuo1/meC/j/81sNO/lfEOUbyMar9oOlFD1GaYUHF4+XnbCPo0TMF3XJq
Xkjyw5imrBSmzan0paSAqf1bfroe2cbFWlJ1bM8EijepVVT4uY535LocIL5iqQ4w
QmojJ33ApsC95lh/umAONhu9+IxDaUszSQPqTkDqVgkwsljYREwvWkp9ccRLciF7
KVmkTN6sPkULzN5t5Ewvv7yWV7HNdgW9XgpQ5Z+opnUjoC6D3p67+CpVEYmkcKYr
XuwrkLueQfC6Zp4Oj+57ZwZ68OJN+EFk6ymycIoqK5sNSRDURy/z4YLHFg69Fkvd
3Zikobcu0YvUW7xuqHGLgqWKlyibHcvOVMR8vel5kIRi4gH7KutGafVgr7ur91KM
Pi8FVx+SzLHk1thgRgBKZG/7UJwObVK2I83Ge93Wtdh6TXHvNI02Y/PkQOGYsKQb
2+vCKos9DcGA4uoX4RGOshpSkObsoyQdP2E6cptanzF8i2UVPmDCuvZRhi7w8onD
td2fAefPYzGM2Op6ieMfd7pk9p+S685TwI+MBW0i/Q7oe0MWur41hhlhLAy7ZAPn
pBry135g2KGovEcmOtCScOIjvYCzfCwMAKFQ/yDNLfqrZxWqiUsoHy40vYZqX05w
0trIMmP5v4Y+4Mb6qK/Ox6HDPE13svPRXW/wVq+LsMsXNphHGSi6PfwwdZQed/ev
YsnF3YphAG+07rc2FxB4eSAzMhFnGvNzIxT/A9ahHNzwscYxGlTuAxCSJSeHw+Dz
X7ej6FpkpFX1CjXNv9NUh25S99gWxW0R4Y7AnxksVMAUByN8xdd0r4huJrGCy7rk
UKY0lj56CTPxjmSyPxJWgoM2Ne83LneyEoDNhEVlbBB65miVJnVxsKTrse0Jw1OP
c+pSYBgMwtb+K4MUH+/6EnJSrK3LInPti/hUJ2MMbEqtN3Z5vwPWxdv/oLxbdpCr
x3eGjioM+KbOBoBJ9/fNG93CyThjho7XNkB4sBTz+Dof+Q1AmO4G04cTZHr57FRE
ttNcfvhlqKSxh3sylGediHUfTXMChQJu5v5ezAGCqgS+E9uRbSVPI6uOGjkfD7oG
PgdeMHC5E+XX4buHxAdV9KV3e5h9nCEvp6SlAh4HB9UcsJxbnU8A/EvOtqtA/DDn
jrnyW2PnEX9IpTGRImrmL3ds0G4yViVObeLAO0y8UldtqVqWGjUl5P2aN/PwtqH0
jWyKoNLVK7KomG0fbM8om0tKltJrEL4WbFAEot7dNsmLpDFYJtzRQC3dL2AGUkrE
DEix5NswjOpBI/8hvaLQN7VyZvEQpW1/AmUGexbBcaB9LuN9XcA8d8Jy2YLzEw87
UOKTRRlGQ5NQpNlgCaQsVEsZAOE/VugZ2Dhyd9kAJ+acG7FYBl4Ltv3BMspMtwHd
Wkq4mX2atorV9qYQHFC1kNHptQu6p+T3TrW7DGcA0yXBIMDgwAfgrHf+JCBQBwKW
vsRgwIgONuXjQNiBKx+9F5ZO5p+rsU3cGhbOb80761ZIPNrUUKN83tEZCkX5UBpA
B/Sl85x6ox1az5sY86xwqiwPZIQ5crP8wlbkJ74tq+DzsZo4V00v33PlZURB88eC
Ar5j1CZcqbiFKuD5wcFDPY0KNdvTs38za0n/xGBFoJlqhPkURbN6PtFCs3A54NWC
uGaR1CTrMWyGqpokM41AImsHX07BVCbCw+ag4Z4Pa6MjFX3FJ2boKhnlHnx1RncF
S3xNk3j6bd05cPvHwaFj4Ic5ogJvVWoUYBEBA5M0jJaCcnlFaln8RGd9D9TyLdCV
5AFnVyi/ga73Pk38voRxqaI2IZ3216r3zpaeCsVVO55jBbthIU8+goZdrNYY94Fi
NpRIayuela0Q5KKswci+5MVnyOgi0pYhvcnSpxq/KsUrlJf5j4Ybiw//r0ia/G4X
+YUan0K2OAsNff+G4MnCPbTj5Pfwc3bbWIp8gyevvG1Ait8HxrOOi9HKfXgA9YNm
PBWUlmOh/AWsvhmFhdl6p59DFdGTOsMmLQRDZbMQyNpak+TV0VORsZRZ/ozKnrQE
jBFOonIe6lQM81ZCbaFDOcd+Sug/4m5qBMndNITIzlN7XOeuDsgHCW/xT4IWVSNW
ixX+9Pqxpw3HNz6i1F/4K3eU90oYO8PN5CUDKtyeB1bkvqdbXQg33oXoQEClHxQG
eTMI5tw2hG7ep7EvXD2Jg1JlhtEdALsQ15SA7Rt4LR3UgHzpVbN43xVKzh/3g2pj
4HJbHmUQsotO+eMo6a/rfykdsNjZcP4R1zz77G7g1iBJd85QZasYXxcyWxLyR+V3
PNWKRNe83FIq6Mi+KGz53h8lO3/lltqmcdxXGbiW4zREec2s9KXwlPyIQc+48ATv
3J8V0mx4mKKR/lvqzOlSRhWLTYT7EP2YlpREUVNfjlwgvFcwv1TsxFiYwpGZhXGu
HhN/4wbwbl5Wukfx2IAEg4BopsaIYZgjlNRfKJ++POe53PIJRpLigvZNvF8uDygf
baSOONd4Gi46ME8RyeU3OdJxOmeIhl7m+xirhYtssK4c0uWpDnFr7XI3pVpeka1u
FQ2xcLLvbvKcom6Nw3TBPDJe4ocv0UJPG+B2IVIz71ObG+AqvWT14EYHcSaxUM4j
QzhH6QMa/W/duJgkVNax6AllMUx/ABhh9LYxs+idJfvDADZNzEyap78HTUvz1ZVI
cD4TV8TSZYU3Fc84k/IiunoxmwJ6DC5Qr2lKkx/rbkMX0yDwyjFVPdU8HS3hgx3v
kmxhuMnRPstiWmZkDeUieXPTFWq1Pg1k05En9g5euoFDfN6VcU6RNcjuWpmNGObe
B+WDf6Wc4zMHjGmHRkZeS0f1sy7LePs0dKVspVuSGS6Q3wrJypZMe70gTXOKA4Xj
VjIy+xMc8VKeKlrDwClpQh1SBnVl5Q3hb2pRWSU3fU8rcRVsJny5b2TGVC+/SavI
fdjxAh4LDNv/ebgAtZ1H5LzjdDeOZPjjYYGAR5bYgbcawAMOGCiB2Rv6ZjW9nV5O
PswR2nwuxEuqnmtysvlk2AGEGpYC4NrSOU5awM4druyYgl6G/SYv+a/IkMPIvakU
4tgJIfkZsWeOxgFQqX36ykqE5jXi0bPhwfvJOJi4s777ocUiFDoY1qloYJfipI5F
phycNqFtqip1Tax8uHIP1mtGzfVV/4lgkmauY7+4Vw+Zl1fCRJ5Oxsu/pubFBtcO
79CFdG5QUfcGQBFHxxNhu5G245ylltpGDuSkrAxZs0ghRbxLFEa6Surl4hnRB9NR
9TBIR8aTc3SJCfdZ9w6iL20/+LxOAGg0woga885UlfcjfSvFX+cQaaKirS4i6Wkw
dyseIP9QvB9rH0ZQweWLyAbHM7QH02LpGjHgQVnEQFJDi7ZkVaD0nQwf+SWuUOZG
8RnpItn35EH9Uh59KcDaX1bXzn/70IwEVG3aX1w33DLY4oCKWCfJOP71BmXFYhiO
gs3HFyiuoiVAs/oIiV95TVnzVb45no5bGbF1zBBqnztuT/43WPBbRhT97bQ0OILt
0hHRZotHnPln/BDt2sBj42EO/cONI1Jq3HpM3xkXJNtoH5oLBo0TWA4cOs2lqnzn
JXLlitZy3KXOq9iff/zTcSF9dYGTG7K0ZA8HaxT2bstHhsDnnMq4N/a23Gl1Z5iN
g1unY+H18ovozFuM2TkrFvHrt/hAP48beRUM8Ls0rPGhxqwG7YPDB319wHVmegzU
iRWvL2mn7gSZDkP9gAoCZ+vKzbdxeds/1ZcXS0+oS8JwRr6poKA910OuJDxtvqDy
yh3Gb/IgR35SN/bKjovaDQlKw7zS3xDFobhg4UpvJnau4dP+HpRBNpcx2RRLK7Kx
h9GLRS6wWT4ZEzOHaa43Ngp2TBNmL2gXCqV/7xdhiw+svGPFGu6g74wtSG8TCH8j
0Ozj30MK02RW1uRYfAf/Bs3jfTMVHHDRRkB6uvFuYIM1hXo0sH9BwtX8MXTFR23F
GL3YHFTFy2kQwBCtOJGy/bjB4jg3e5RTv2hJqHkItu85r/BD1q0Uu8BvvDZ8/yMd
4cqGfmCl2ZI27xR1z6sDnZUAOMNR04genrExuo5I2WYuFUDeJU/IAGpac2ntSY7t
HruktInECPSDEM7o991JfZt+d1g9H7q8RVKdYI9X6Lpv+s377MDmKjjdUaWC/tr3
rLNSXx3hRo+DC6ODLf/ftRJvp1bE1Bb0raYQrS4Ovc1UmUmd2hlEqxceuVvokp6l
g7UGsp5cDBjY3hcU6dVaQQ49txhaAlFqTCL/Q12PaVeZQ+m7naj93Is12JVmGYf8
FHvX6kEqXpQYtQUEV89SNT+Lx4oDcLLngvBqmpKKR0GxCZzCoWv2GHRSVnH/JLJA
f7LfV4IIh8hfyUlhrLk1G+V75bcWviw4yvXfRpcHKBTkwmhWaB71208k7BOcosZb
QVLLj24WnhNkcvOUVeNtsl7ei+F7Z5FaXVpDy4dtu99ChtGAcABWlW9j1VnuAo1N
1AJpcxw/vikExhY0yqy43IEmnmq7RUZUJHs5hwggInikK7IGIBTYxERtFonRzXe2
16SKNDj+7FxdFgh0vpSE4QQ6gjGvX655Ik/VKA9tC1MG8Qgb/iP2qKE9Cj9YVU4b
ih9fe37uuKAP+JAzsITpyrkWKHnUsigysseaX4+buy/Q5MaaOmevMhmImeVfdni9
tNYkZ5WrQHnYV3jWxMWjA4GspvdARlUCcotwxH3f5YNUbTjPXMNJVctVrD5qp3Is
dabdza+qWrwktrd3ki4sCTg3TzNcQR6QwnDWuCX9SNIr+hyw/RvBgDqpvOXSLAP8
WS2/C/Sqehsxc1p5LPnjExgJi3Zzthkkj3JZKT4zYkENZXlfP9hF8aKqM7ZTfOr9
kg7blPBLDaDnrflMGSyfDSPcWGywguRdW9nj/0/n1XP5AF49wOLiaRCyPpF9/GC9
SO3GKpHEYQN24PGRyYaJAH/EXLZWuNITKRlB6SNWvRTPkxOsd9xiZV4BabDN948y
NpV5xaCx4uLz/v1C3D/+2VdbTgMV0ZXfDwxWAs28lgNwWj1t4Yp9kVH+S9OsAfME
SW6L6EApASFj2X8j4fHNVA4VonQ4TPfldD+z0a/F9idUqnpnRfP0cvM3gTdimVSa
CioBCInx7dlNN2PrpE0HJcLAg59p0YrdtA5QqQTPYOSAQZxsTLPaUxAO9EcIUcDJ
5Km4fpzfQSNfUd5TbigJ0KP+AYPMl+4AbCr7zN1IjbgHdhym+gSfEEfyJP5tbvDA
WZwqeb0mIr5GwSTE3b6JzEc52ALeRbvw0hMvD+/AQvlkE1F887DrheoYkPOQnRCg
M8mSxB+CQlf08ZVQvyKBEAl+t/8q7sliCdgrFFA40pE5sLYwv+agYR6yA5iLb6KU
V/XXDYTbJ/FKucx6DZP0QRvMQtwprgQfiswvVa+0FH6pc5d8UDwPWa22cXin71u/
m4nP8tG4fnkbhwFoL7COeMKOntKPTy0act6B9JZl0cGU1VcWd45iT40wpPsxCwxD
qHAnez0zyx+2IDN20Kq1WkuiRWPnBdAuq6QWAwsumRtWdHfxbGQ4jKThgUyQdwSy
ScXrVFfjyqykkzFYd6MqcQ1UocRFfm/Mj4z616teDDZx61iFSsl8ZYK5EZZcVSRR
CNBfWqTgV3uoLzv1ibOtXPbYNzIEDOFPj0aQ9csecXbSjUOHam7lKNxR/Jykzepw
WKdWaO4fWkKsretafJWycLhHA0QYpvgnZymXcnBt8fGfyjccnlZK0l7esvzAHOTn
FNLq07Gs3kFUGiqxHbp/4FAqg0Es5zws5p+WYT0NizU8u4BA9D953B093ky/3lKa
j/GbQxyiYRJdy24IdGWiDkcI44CmKu/ZTu6XgcK9pSVDobM/lg9KL49X/GYsXZsr
rZfTxYVTuSjh757S/E2AUrPuQwQewWy6E4vpQA54thPwNT2VG1aPbB+1RjNia5uR
O0AGOLUTaHfXkJ9d9yrMQ+cWIBPXCUi69GtXQLl4InI+TYKhYJO9qsG0RWYda1d3
HoRGcPYj3gd0YbsuLYU5YLpCGaAbI10NIAC5MqADRPQr8u//biyYQZ0z8sykryKi
mOwC6o1OlMenNjMZr1DLJ+aBvRko/2wOFt8qfCSB2K8conFy83N0dKh4Si2kWt0n
EaJIttRnBewHx7uVH93GSCAQ68cavKg4iu/Ivq8KvQHmZbuWktIR0WIg2XIOXgmL
7fY6mEtHuwXmxdlKwlKWJOQGq7w1nWXzqDMzBZZuV1Av5gQDtuNRdCON/XL0nX1X
GH7cgMyUDS0x53vAkm9FXZH4rdT8aT9TM8jw80YAzoxDrriUdo8k/I/vJjLZ4LFu
y96o2AY/ejOEgPm9WSV57scqzay6OO+wvv42RVFy3XUHAyt7AOQk9dzab4vNrRVn
CL0Gnatr8K48ReK2CNQINK1k67ye9DwkOL2tuC+z39G4B+DaWnt6nO0jFaSAiZCk
r7/JUjH4uuqvGaGnqowYDSBWAQFz6/drpw+Oc+BJIsuq+aXZN/L9VhYSREBFmV1o
QqDK0HoHYtrYU89Ko+Nu2HB4u4bf58WYE8d/cWbB/iDYsk8onIWIM2DAooh2K6F0
3Y7MxrFAqGbJ9GUefTn30fWwxUaY8T1pcbh3Q6kpROApF4Xol94hQPFB0COyAp7y
XayKvQnq9xCNotVTN7QKcv/tP78JwEfXtZRSfsMq78SqbDXxc6SxjDT0UQLWJoqt
Q9XVVmppWR65hu4qXSJvkiAHMERXT49F6AvwwGAkb4PPUoeFaswN8+cyTNGluIpG
8HaonCjQfXsefjUvTSB0gfuS2IPQwfgekQ251FDfGQDazNeOF/Cwh/g9/UhWzXlt
9W7W+/V132dRTyeJ9Wu9WwXkn4yCkhaO6bzAd6gOzzPqEAVGgcNmToKFoHrhR5Is
EYF1KYwuUyCbsdZGng2ApIZtNj1fz2XXmqEGY/CsBkVg9XWV4QBckQHJNjmtRyqO
R50WXkqJlEo83HJ4ry0O0wO0yFTDWSEK8+QNRUTAmAdv+I48H5GZ5VXvhblM9E90
r+u48xX9XkalIovRNQyYayiEK4MHGPU4Y8ZClLcBSMTSjDE5BuUE805opM3IiOJK
9D0xiluxRUnGq1+vCrtyrKOxpCbZCpUUci7MYTUct7Qg1ZJfWmRS9vGXXqiMtlC9
a6OKTCSUGb1dMmv9M4r4MDU00SPOuQ6pmWhKyErhMPzLcJlF0O3QWugNWtluBVxt
MF16BQkA9kCL9quHjdpL9nqDBoswTjGxhpyX3wRgO5HxlXqA7veIQwfkWeVq2VZP
FLIMAG1AYUYTI3WTHU7zTya8Vqatagbj0MWzDYC8oq1OMcUIYUa/bemmajOfwQL4
TqcbKKSz88dq7dPqziV1C/qFf6p4turPbxQrzuB6QOpwQN8Dg5Oq+LvvR+ua6cbF
/JZNVK9KMUQx3W+TTQZaEu9YEDUfd4A7njv7kLkwfTEoub/X07XkhkKb3PL8YAq0
r7G4DxPZObcsQHMeHg99fhSXH148ABOxJWd/wQPAjoq/zZIM74Ojpe225wXltbHz
hSrlioTcele/AMDYzVdwUbqQHdL9yQ2dvTBlGDyhu3lTStBQsmCZztRuEip6uOZv
pAJIv8BQ7JxMllScmm46foD+ghqSNCOlbKIW40mMGFX2g23LEbJo4DuMgYZhewd4
lopxfx1wTJeMpmLNcmvzrOdTTO88MnCU7+CApdwkMZF8TK2F9DGJyIs6l6XG8oc4
SuyFVyeXBdyl4m4d4+4H4rM8QskT48xMVwawdrNYw2ENs7TFDxxHJgbbfk5j6rFI
vbLkorRXCyP5k85XNrSSYaYbLbS0gvU7J5dpKC1+BQLM0R12bnThiwfpvFPzJ1jX
cF6f/1t76wR9Bnr1aU5RowN1AEimxZpqJlTVNcCbPMOj88SN8pYnQqvZiVc/tc0d
ow9ey6tgiDAfuqVRE3Jq1/UxNQxDnCxTLVBvVpXRk/hpxAuYuQM1quzeAAZrLce/
ikJY1qOtRkZNpbMqueW9qbAoBmuHiiW+GTM7IJM/JySQBzkTJBegRyWgoTQQgHdV
4CETca0W8Y8CXre+AYSDm1aHy+8e4Yr1BiaRSHLMSGoyvJ76QVl8pFbqd7bnjCJS
D0l0zLmf3UipyUuzuFsQUM2KdEJAh3f+Ttaf9HJoBWVnCZPSCnC+QSEguG9lYREb
dygLgCyonRAzFq45pxTy77NlYK9xz4b4cynON667DbFwRfdryAz73tdRwZsWNwq8
ntqBxPsQU8IhkRIEvzR3smGThOzstnPPrItbCXClW5LVSfs2JGYkR1TPfakSjbKV
vP73/SamIFs0Vx7l0s37zKkUizD3OR+2kmKM3nhezkZnqwXQakGXQignne7cZuyW
6dX2i3KzNeKYJqeYu8w8BkE05dbhDehYuIIyrw/xjex/3XNujApRCfqllcg379ay
zMK+DEw1D5HPpwQX4vkkTxNVI4UZrE6jKwPwcp3ubtt4LGJNL0OW6qbPWEbJP15E
R3KWAIs+79lOjoJBt/plBGwWfDaYY8DY/7A3zmK9ct4t2gX5ouxlxXReMqxSFF32
ApC6guMRvahtSk2Ig9yGBrspyjxscZsIERYn2SSBSBrTzY+BqhddjFryrOLebBu3
xjl3oqHsGY1M08LIkfgEL8iE80wmw11pa+KP0JRF8cYiwvfGIfdqC9uHwnvIWhOU
Y2F52QYSlAjc04hM09onbmlAYe/7LwKJqpABe7y9jS/dHjXw0M61cJSJMWvA9J0k
fDWeGUnqXfbrx+gwUHPQ5PhNsdUWZvDwI2J64qvBqMtXSCQDwmPSnKUFY+M0izWp
kkOD57GxqCfcfBgSmGVxD28Y98YZ4Q4ere2Y6Aj5TWukEw/8ceJE43oS6nPNFR5r
KQ9AEzRMB2lsYwUFZyidqRlQ4bZ6p6L+5bC8Pr/UN9E1EVf7dmktGNvJMiiwq33V
QB/ElAU2yXrNfQPKZ/HbX1oa82qPKRA1KtVUvFVpLLiyQCQb4D0xArSP/7s27qvj
KtGQfyZfk4eVz/Ywn9BIAZFKdctwCHHHW8iwcykoo4PMPhzGt9cBsX2LrC5O/uL3
UHSrdbj9jN+IThb2r//a7Y08w83HbUoGKv5FaeU3oEXGzgu/9D8yTDTfJutBI1YL
A/eoQyk3fYIyvlWWjiCk9QlyjPsr9KwLWhIREjKeg6oU+9sNVsvRRSxh9T5K+H8V
V7Bhb4E74iAOAfCMvCZaM0YlDzLvz6MMdylKpVmHW8wvxa1+Fmc56l9rUnTBUsiX
xYNtaC/Q37rlUccZVy6qLMSMz7kEmMmmvIgqccLTVU/z+Eje0vfepWdBiiGgmZxh
5JklqleyXqb0aiy5IUq5aEjlu61qJA495NhSdK3eZlYrI+7m0WO8tu/UPvq5EQ1x
xGvUVmGi8YDCASn+ItGFl/Apl01NGj3wceDkWvDSCpUGtnY7kr2XFroSvu8WWgU2
KVSVmf2sqMOOaSbxLyVrS8F3M+KYcvzvUbvgI0bUbPqP+Ajzy99vBdOqw0utpiSs
QsEzHjdZL/20GMZr0XkhNBdXWc0ocIYpsrsKF3nglPsWdtVwpFRogSzTCx8bPciB
lXaajy86WWktN/tQuDwzVYpIMsbKF33Ul8mkZ9wgZdHLFR4pv5bJ3SjaC6BLXM5G
MyWchNCr52/YkB/4uGzWJC4YxrTHxKW0Ah0sAF7aO1ZqplOem0A8HqirN9zWgHRO
3aVnRBOBQnGR3oGs/Md3hrTbPJsuEadhwJVuMVuT6MI13wGQ/TZ3nqA+UCadXW8v
jsNem70vD1PKm6MzvAhU9Ay84FkZ6h3vFIYqs1mT4XRgyi2t+UBC4lE8PusRZMiQ
sKc0b0h7cSL6fmjJL1AnAyCBnSMWwQRvPKNbRD45nhyAiqN4RJBVj26lqGA6uOaY
0zGhMI+sgM3xZYD7SUKvYVMGnZeBUQusEVsrE/OR6LJwndp/fjMYxNbhrrUuFf7Y
OxozJEu5q6yUbnyOhw4rkANs/wLt5gcG2FJHoCE1bG7RQJL4Wm8OSeF5X7siXNpX
8uj5HLRg4ovk9k+Z7vS5JooxoupeuJ+kosrhchE71shNYPpPf4cc8G19ITAQS+4/
0Ae9tKwBQ/1lClYatd19jKrqdMcNzZJ/XA9j38/GTuQyLHij4R0kB0f0cJLQ9iFW
7Ele3ERl8jAlB6b5KtE1Bl3CRYDyd39H6j4KUe+NjQtNSf9M6tVtavxK8pQKlE3g
x3/CHToUO74hCXJRabyqO4hw7RIE7bSf7ZJFPVkCGGKavF7UX1Bw521/kSFB58g9
r4jfD6qLT0r6g5eyL8Bho57OYA+zCJsjIxD5xlvCTTDvE9MPvWkO+zpYJ/FssNhH
svIAnvPHqS8j87neUIvKIZgce1QKjcMAlA5prz3/OGAbBJCu5VF0hpJUVy1bbAL3
Y9tReVqsebzMjNS+ypd0jhih168PRx2KIqH852Rk77wOJw4YyEuGvkh3tlCVXLO7
e7I3O8KKXGF1SXAZoXLwHrrFKtzkEto6WCI9pmyYChxYIa85NvzvylU1osgrWIS1
pEJw4rnLvFDfF4IPZE0Kx2CE+bV8I6LksyCc9WXuetuuuGoDVf1mcMmMynfeQViH
3mVM+NBRX4jedygDYkpybzSFBINAawsYRaC6uLoG4p0PAR+EStcC9qlof2N0Ln5t
dKMA06VZnX/QAB/7sPRGZCQB5yC49O9sVxMjLegoRK/vRvhfoImDl2GCLAAWRQac
ek0x/oOD19v66JMyuD0A0UIDfTHlRoz3peU8dsOawxbOu4ntHvSlIIeroJwlLtdD
4TCGgYSUIWQ968WqDjEWcBrCrlqxLi4G3Bg3jy9WJnS6ZOQeovsm+TJRDcNoMBqK
7SdUCKxO1exSinFyKjvy3nwdsjX4VDwLjm4+a26XSVAej2y7q6yqaVzFN8m0PUZF
Ib6POTE7Dk/xhJQj/waPZastjsAqRBmB4iSKwzwZ2g5hM1LUj222ws1GTXemxqiQ
srrGW4kpsoccGXH9E4tbrLkUDvvEk8q4fY1UhlVhvRiG3FGpLRD4PWXezwxZgorA
WSGEJhpnXdlQn8WCNzpltz6m/KbTArKqLCSTl95aBP5yRD7zmK+4CBxuPUou6zgs
VatOkIvythWjCWINSLZtCUqJrCSeb3aODZkUevoRaLWmX7AKMHyIipr5/dqDcl3J
tpUr+PQoinMRskEvNVy1+lQq3eXqlnK1YBshvh7l3qBmbmPm8r/t3aRu57FCmOez
mvKDLdQNiIVK1/OSCzyYEDlvSB+UlrJlmrEAHpnn8Aw4IxI/mAoHDJoqlZydrz/G
ICJ+WdRrmlw9NgEr+fJuM5eYCTE84VmdEkv+soS32dsmgyliYqmBrD3BXeT8p54y
xFqyUcCyLJ8fX8WDQ3VlU65B0D7SwDb76TWO8G2Vep8KZl+D/FggehM/rKgFRr1E
TkM+Pyfh4SKJ0LJeO6p696ZyoiNiXf+1QwxeGqqkuXlLzAeTkkdN5b73W9PEtxgM
xVpcoNOCNMg6d4zyCK0em9KTdqDIK2FloPU0nGp6HfaAtT8brP6ymdPcdnF/bkES
aI83UuuOgNJzO0tXECjK0l26iDhxeMArp16fx3v01c4MEXF2YzB9P/f0dtfJ2lQv
Aq1XYXt8P2t4Y5j1UDVfESoNqEb00ef0uDtCODj8I91tJvbW6qKa4C/yax++KZzn
ehrMNH5PjO9f3tlSmhKxqoZR6PDhsx1bCw6xX5m3pUSNBK+90ZIy2CADF5YmFp42
7SPEmwoXdPXaol4xQ8f7LvFWMNZF3kGIbshTXD0DgBvuuWoC4oYq0F9A2XZbd9X5
2z6Fw8vackv0N+YqTWUjM2AMDl+r0grEk5iLxb53/lk4nLU452eTzeYYXeHs4E4Q
8Qj68KD3Jt/um31YcPnrAI/5UtjfLlZm7IqG0wD0VqkmlBQ+ot2vEKg00rIvVy+P
XUKz7BhxbrZ2A/mndLdvWwFxd7De2sOaLcP2c0HWAnxcTfLfYh1Ty079u8EXl3R5
Xp2A5fhl5iT8M9shif5JwKrqyrboNb+VEaQw94n6AKuNls4URB4BKYdHiZaI//Og
hrUa6BN6usNDZNOtKFGs4V/qsbIttj5HYH0xcLzjHGaUL7cHdxMW6UNTXq+b6Dv2
/uGfAz+r5YMCJfYk9ifIUkRp45p7HFzbNuwRKKESl3tcyacw96NOkB5lhvIx2vyN
Jimevh1oD8aHSPzML45t0N6yKxmiG8PA12WWscEZga0SY8yhjPjYPmetcn9ZXjvJ
dLaTEJr6/at3KWAspTPrsaPPukGY6vG/jZkYq+cshJW8dVa01YUj9txMvmKubpwI
chr5CE/LLN8OPXlWhRyV5jbHsldCaER1e8EjdV6EmhghUNF293tJ0tS8CC22V/jb
Fw14Uc0HbnxDXABIgkSu1AiI6lVN9xH3I/IIInnUvHVwWiwW48B2C4HjVQXkXRD/
UjRBaai3kB0c8icdKz9Z8pxKHdXeGTsbfOPfKOUIn29hmEggdtANCgVhb+9DMv6Q
QRLx7e1h8liJEXbq6046syClEXbVJOKu5jnzxFohJM0pegw1wAcR0DhsgRTgf4Pk
XYlkiPZWtHfj39sI70SINgs0TSfk/zslCCwNUWr6SrjeIxsSzTR8gOdU+m8sw7Uj
JWoz4+6X4kyBi5vpPxtKg/yJXDcdmleK1OlDSbN/KXemuUT9CU2QKmblIVRsrNR0
E4n/VeRtbllZ3bt2IdTDqfZGgdyts1lVARu9yJ9YSM7lA7MS9atLYK1u1t3xK8Vn
r3rCsLzORPELx+2Sj26oOzC/3HBFIu3124s/PiWW2apKqshxaMHwiv+lRLcXhjaC
HOBZhz9joYpcm+h8i89yq1lG7s8/0OG+3AF7U2p1gSIu5FcVxLEZ+xDHP81eQAr7
CyIRrkBH/Y/LiuXpbqT6uZ4sK6LB9qAe0OL4LB6rA84a3EcXQW80/HdIGwBKEQaO
NzjGFxwwx2WL5uwg1bW1sFaitlwTDkuYaGxAXxo/8z+L7fFFWnKWYCOfVtaMEGMM
xWX7Lw/5CwaXaTU5f6XtGCaLezdpD2Y/1Ohm4Khr3MjKH4ipfwLNkZJwcZrpKwnY
wliEIKeWSMKWn97zv+kXY4BR0FN39sTpXPWgb3F22Pshtfhza6W8zqm/RKsXOtlC
Gw/f4kQHBu1/ICQk2Y3x/BP0vb7dPjnA3xULlFDIfsQ7mDqu1Ke/PS29NZgKHIKJ
eihgB3oDkWrhozryzAGxIdxVNqNI2QuBAYZh3vkPWcvxZl2IhAQPJHod9RbouMoh
HKd0/PaHpw009FI4JYq/8MDqqrRRwBmRiKyOZspf6LyUFLILwwocS43CP5W6em12
5UrCNl7r8LH7yoJu0nCQtgd7ajVKPMn6qloogPSzaQPZ3PWmf7bgDBwsoMMU24Hz
LS8TjBkUDH0jm6T2z48qEYfpTTW4yKG050vOQyNT+rRENvtZPzux2UbPvNyXMA8Q
WWbJZIEMb6Q0x/SJIoIwSY0h5TLE/c5aAy8x5cjmFqugDQZlK6Wvauqr12NLqnTG
hfiHm48ODvIi7ftX4qxNeeGNdi3gyyJcWkWnpHdO5YvjUDMQrZv/CjW08G6C2fUW
UdAXcA6PECL8esqOQU5cpE8ksR339tDwFvbkwNAtHzDUhzhutFcS9PS4P/DUXptq
PSQLdYZ7QKKJB0+1uSk9LZJFqe7xsWJli4+uRHALQVO/ni2PXLPDzz1BcesB0rao
uIptWHTIKwTmrsQeupxctIKO2NEoB3GfWCLjniswW2F3wBK6sTJGFYwyACcDd0hh
fl3hdMh33FYGd3IDYPbHW7GPd03IXnMXq37JrGmCw6iAjbUouL/vbhfxmrmdBC5C
u40lHQ6oll/rKuZOf7fIza5uwZ01/7AIx3MyGGfUEDq0sI8oR6b7s+HW8BzyjwHE
GwgzCO/2UbQlWqTjVNPf2NM2gjq1humm1A9gOPDGCRwDnREJjh0gEukuLqpl2Nzc
HAwny97wqHdlhaMImhXbxNqXINu905X91A/ftfAZPqqHkw8rodvbZn3avI1+6S0f
1izcJKQOhBXMpTccLhem6wq+WAOSURddT8Lo2EfT0wOb96iY4dqH72fR5XQnNQ94
MWXrZweK9MrrCmSYBn9FYS7/D1OU81lmu4Ci7N7ptPlPMGcQF1Rvp4O/keNehlMo
vgWpawevachFJkw7KuCAHmm0zxvij7iV5tVgTtRU+u1kVrtmlXDSYN8HNhiPTsHo
A5vsmC2rLLt2XlDtMLMuSQY2C+UX9R8s32jFgOVDEvAoX8rY6QDUopz0BHa4NJ5c
y8DFBMozl8t2B2Bep4hf0SSyN+iaaIr3KdHBXq6JIUu41nQ24Xb6JVlMSp39zyaG
K4Lyf9Qiky9rQugeRKF/2J0Mv35n+dCPMU5x6ZTIzER8se0vkdLtCEIUP2B+LkU8
7qlIxjPgqDewcTrpfy1dXTWnJjS4EtzEfDToGn8pbDO17sNDlulioG+J7XX8kVWK
Zfcs2Yom6xDOu8JL3MBbD/hCxjx24jmj5Q+Rl/R2330dT+7Kxk6o/uSxCMK82G+J
ECAKX2ei+3tmE7ktNRbjrdL1OpdKCTwGOnwQa8ClIVU6IecztVMZey8Wdt5jfZ/P
jAkMihd8+edV1jX8gcw8khOgEGWXm7OiPuOucEKFzR4NGEpmYMlBC0LHTUPbX5d3
ohHvnGQJzb3rLvabI6rM7kmUPibenWz9Dgkg+o7F5bJdqbYB1N9zOXamcE/oq8gP
W1K0kw5X7jcBYNnx6eKlKOkVwRp7FDGAckio6JQat3qNatoqjFTPkGUev5doFkHK
Ml6uVRJOmqoMciur6+H8qJlSQLMyLHBIfX5uQnstoDgb8AdEuAkGqCrpXMnqRfKd
3H1Gf+Fot6N9SvhiuB3NOT2Ha5oKf8wzW9Z2bU3w3o8G0jzSDODz+0gda37H4Nin
PmJMi83+FQDfaNlqLwtfF/IqNb7XUHzYD6its2xGnvxJ9w2DygzCKZjVQ8X3G1A+
eiK3Nx14xpd5MBSY7zKAs3Z2KgQbNXCXdA3L8KrYqv/qy9HdsQyZNKvtJbTOVCNG
QvEG160/ki/gCHQDIZHPIzCHT6on1nInZH8vx90xx22KfVTQDBt4oHZKZdtE40+z
CFHXoNF2WVrHerIICBb/qxreLVd4BdtGyxqsyZIn9bqe+8Iq6Hq62KqGvKUvb4I2
NeKU0KdRXxT4ro/Ag7drRMQ0/AF5rA7b/R7KWH1X1LPBTy+K2synAGzAatsD8AX1
1QJCYqhhCVu8xe3kKRT8z045lsKN6K3OSI5tUmXkrOkykOZPTCLfkFiP40j9LsnH
dpkzdgonKmoNj2xWXJb+lxZkeLW0X6w1yMPwKPZ9e/DyVGwpxAIIRlGdZAN9W1A/
79UY/dh5/ZY12KW642Y75ru0NxBTvXKnXJ8S03PRMLbOLxZDyi6MsazCN+LLPI/k
uUlc1NHz3b8aSHF3vbcQBALtud9QnaT2LYJT85d4H79reE+qci6cazgEM2FlIMlb
kpAKvUHE5eR+TMRd1eZaw7phRrxoyiXOe6AQbxDmpYfkXVN2FdzhQqIB4+W8RCRZ
dGv8LPzWKvPYPOlyI5ykvAa/On0v41FkI27xofi6tLdNYNaYRL1ulvp9RzsnsbfB
srbmjq6lkxCICt4MvNLkr4oaHzt/abdCq4e5VV1yrJG/eIRpF8DJuNZ9HNHfAglK
jeQw4u3tzGsidIPUPXUl/8A+VplzIFsARjs/6MLgK/9X8+Yuw+s/6RBwuuTlsJGK
cxKOKxQZ2U9y3kkEYLE5oQ0MaBxF0i1czcNQcRsfF8WPHSxj9KrED9iU4+m91/pl
tgNM5KWfvEobf3uvz4/6SQN3Cvw9NZI0koh29jhAGHnrqq7Ak3VtEs0q4GCHCHUK
Bv79cQ0XqwrsURB/FKB7eWT/m84TyAMupa4Rd2zeaFsgZgWbDPZXvCZwz8LLc1bh
IpI3YsU+GnA59OGws94r7mb8lpR47NSomMAVQJMrbrhmxtbHO8SwOTA+alxs6rDV
dypyd/g7RTmbS0G8gRUedrTPjblpO1dVDmZrBQVcYTo2hp+3YsQhxqVKlB1nm0s/
k8gtqqHzw0Pvf0e9To+Z5JNCb/CPp61Sm+vvCf+MnzEGR7FUx4zh8NN1x00gzcyC
VvGo02QvlwFCPCW3I+47IIDmq1ecN/SULhEMAUTzpvVqrsjVcs5rmUj3MdCMkL77
N4Kjf77qqYe07BYeJ4pNeJR8uT0/sRwmR6piu+6tdLqa2S9av170s3HfcyC5Gvu9
/PdTZ7c/MXc6lvTyLSEH4TERfLVBnGj1dHS6uvJQT0lfWQBt+a0fyWrhOpKMc8Za
iNyzaA95Ykb3JdHJAXd/ADcRAJhgs8pHdJptc4csuqGcgNRrHD4BtkfzhpHG1bRO
223m1fiVidbLwLhZv8Vk6dNVLWA4Mp7lLM8GFC4IFvfKpGLODRgZvAakxXeUSzEt
a6BMssBx0noCiQKk5W2I+1+G68Hq3ujoKZb5bbEN4nB/aM1Ws3pDMRJ5Ec4LBr2Q
bamHLOk7t69+ocRGl5FPdL2Zc+k/oUeyV4lx4pJ+lW+L6L21yV8j1nX62LcH9Bgl
CqVcscHpCgmc6gaQlnjChfwYnbVmbuJfxuOdA/rUlzBn3sLx8GeRSP4gEVyZPObq
9YfSmgEPBbRDOGVjYDwqE0lFNPOSCYPj734uLaC0Om3fIoyfuNAoKYpHSiurb8aO
zuKKRzo2TQdgkKwOhB+BK2eKFzjUVC8rtv9ZC8hGAdl9N60PDEMU32mBjK3RVtvd
F8po3o8viPICQvAkYYjT6mD98L0sVMUbyBg8BHdGpLaB2AHskI+wtlPhYpfz4W4F
DghlUvI2lNcWv6gkcGRFsW4D/qYykozv1unyjRZc/REp44Hh70c8uQPHFg4lz2ez
Hy/i4Qrrg/4k7IrXTnYniuW2aP/CKAd4p+61g8Me+Zt689pWt8vRLoScM6hhWpCW
dW12YhpCs6rt1nR3ycfJWWQrnIg4fe6hGJ/Yalo27tHrgomtdl7QmgVxV5E0lfLv
pLH5DIwVBObbxZVgCkML3tO/buUlFmuSIMREI58NYL9hRkiP5Pfq+FKCxtw7d14P
xx/isWcPzpZ4ScQKsQ91uFBpIPDzCeQE2jgjdN1wawjNtHdIMf0SjkVaFh25nCqx
BFb3nBl/GC3cNoQthRqC7YC1H6ohfRFKMne1EmcdBu8RmvSuLNzMU8LToT8IL5fG
Cz8ECiE7nMFncZbsDkoELSpkhb1xWPX/MkS9+X45AtRW6wO91cPuaytqOPEXNe2n
Xj2hjC1cmMCzzf+4L4VDsSpKvy2ieVyDdCi7c6S4K+5+zLk4XeRJDUg8aXGzL3QR
Cgnzp04+WD4Q2xQTyDr0GN6kmBHfZuYNMlpG9DSuXUAh6/52qChNI/cmI48NgGwY
TQcQ/aZdA008IV3KYo6sADM48queMAtT9JVgkdEvP1bFTlDFtur6whTyiKvQ1xYB
pW0zGMCH4CGn9Xlomm0Hqwxn6kYLkL4KU6dYIeMIoWNQWMiXwMBWbRvMW+YVWTlp
TQbANFHduM0dVI1SQp8qaYVFoI4rck0aESIMU2yj5JZ3SR3VYGO/X+jCY13Wi42f
RFhi/wM1WUZj95y0kq+am6U2w9HJwOTxRcuU6NLxJI0AMQ2eNlztBCRk47BJMYuS
0OPNPTrynLGSTejOHZZFUroLrlcVSe83uwfbCxfb3ix6hNt2prSk3ZMsGUTADJBQ
Bh8MdEnDihTH71zaIgjh8gXUwJLXQw6g4Hscl7TofDVK86Nd21HYJvYLuhtLbkUs
bolS1CB9FLv8R+NphIscJkTZH6TRLFvjzkV/UrOzyJ9zVEpioXhWs4icZFCkj/HP
384PehdTg3t7vtZNan4zhtTptwRnLa15/5+xpA1Z2pJgc1jUzthMzs+gQatFpF66
b0nApTxYrWO7h1CTdng2yTS0uijeAYGeYyQ4TcPfYshXo31B/AvxkRvAJ3FYsJNV
/Hg9izQg5YSzH40U0AnFwET2uhXOQ01+hKZ7pjTRxZHO8lgDGMAw+6QcDcbPFCtU
GblggTT0C6DpZUM3db3vXh8fQdlcVYsO6QVxA1h8oPzqcfl+FTzn5oDfebKgeDf7
HdVVY0vuGKxy2j7oSlfRinEctLXPoRI839XLDFKxIb7AiE9Hu/Ub5AHGuXZsygIH
9SFEmXooLj8xPwYWwZ6hGYHE01003gYsH1Hg0QZxfp7nOGY6pLCTCZKBL1UFvf/2
+mvFBTCBLjp1VzqMWhrbDOhmQvuyPrdlQG9+8A7HaQCZhJpM/0KhFe3oDBH5CJFe
vsJ7sBahhdX/Clo6Mf5usuVhlxwQqAyuBDIp7JlrE6fULI/ffvS22inMmiBu+1jp
y1MkcU4uIuXNqm6u385ZSiD39F3c9TXC6ggtagsV+aDNXv2hBgYq3ugXrPJ0GEzD
cbh5vKsdv4y/ul0U5m0TZv2x9UntWnqC4v0bN0C7OgBFBVEbrke4xYeNU93H79y3
CYuFbiY93o8oYw4cq2WaKsoOUNqbP5x//8Gf1kYMQnJWaOeaZjuZNBgzpYIOnGpG
VIWB6DXC9ZIwBMGnNCQIbn7ZKsFoasAKc+fikc0o/Kran11wiGx2Mfp5EpjOtV92
zKnBOGsUUrF90u8UOeeRJ97U9WDTmQQRhm7XnUQRLeaJYfqnjEx9pZHZd6reCkAJ
9OTG2Jf2xtiQkHX9KX4tstl+PvvPcF80yQ/VfiIEIr3nndQCAPMl6APDNTy0bKAZ
lKAfOWpJ1O0R0snFtCiIu84HOb+Rkio35eCrHQVyH7SLxMlNjHbUlr3yoNcLp844
3l6D8f3N1uksgvYRJ233Q2LKwYsj6pJDSDrPQTNFn2+9w9ShwYx4KcYfKahElgd2
gHWMNv+fPmc+5U8lzRG9wVdrgaJquClfJLLafxrjeqH47P5YTjf76v4cp88F1M/a
GL2O6bZ9H+y2/jYujBwDlqdeZPbhhWThClN/kOAGsPjKh0gKGKwLy+VSFarNc+Gm
2v7fl4gIGdLIhHOBawv3HbMezf+hAByGl5KEST10auw1bBrZS6ayQy0Q/HeqGuWO
kqHq6rp9hvIT6iS38zH2kqLZllGsIltoFkK3NV8clxcZ7DC1NR4mYUjrmfw4d5rG
N3qpPpj32Aq9TEvmzDHQ1htctjRW66eVR8Bzf/GfH9N+EzHA58kB1hRJxoqcXOxD
JmSxF32fgP74/oT+w5yGd6itNYQ5pmqG/l5bxqLeJwCq9krAU/eS/Z8PsixyRLmo
W8ert4Oabp1LeW30A2m/PHcdNv6Z3C3jtsNWTqYjL5eCzSEw52No5M1Kq8NHUqc5
NxsmEz3yAjeOCBUqjmrI+tk2y1UZw9z+aOYxCqmsVz2JQJAJ0aew1TNKprU+vR+S
32aoMdqRC6RgYZmV9DTVhKNUyeVT0sDtDqR8E9fC003N15JEXsWemV3jIDanPDZM
40GeiA+7DZPZMM1oWOL3qWoopr8KaaB59Bn5d+3d/HVKLMLCI19H2A8kIao+vVDn
xHLzfZdkozPMwXx/X+e2kBG2PUv9TmdWuYLFHG4M2R0FH66F/6uBH8ll/zgSS0vy
NiPxFMWvum/rWQzmAfuMudcEOzycgC/c0Dscm+AMoCxW3g5KGpMBs9vYG/wAEBDS
4VrNPx5Xd3hxBK/r4h0q7AP84ZSIqoo1CT8d4cL3q3VCSgaRT6eusjOpicyQpVzn
m+aWUmuvRfYGUPtva18l/zv2rd7FaksGIsHCDYkJu8at0fKAviniAWFaVW4h3yRL
RWbbX+4TFg28OudGfh/phN9dMgdVoRhw3WEXUfoYA1aQI0aPeaqoJtO1JTFN5DCq
yVtovcny7oq1/oZANNJLiYZpoNT6iv3Wf8Fz+U7tLJWocEAkMO+oHCsJZ408N3Dh
ga0T9Gz9GGAzD9hqpv3OZlexzpvDwRvYjhoR5sJ80JGF5a4umXN5r/8ZY+yG0d2N
f/Qz2udSZWcM173dJSsTJieXoNu3OouRodWd3ehpBAArhVhA40+9coD7wmZkRPvg
ZhXLPJXL508d8UDewDtn2dgQuTesqLVaHWGnaGuWCUqcKPrUPRnImbGxOpJNVzry
Va9Y/rztsPJJedvsacyEFOiUEK87xfWJNOj2QqTJJOq4USgLtj19/X6vQ+M6oQki
OqO+uhrRN8iHuAGxDcxthU8N7mLdZ2h/db2ymOd7j90u2Lj8EaRQ701JLniW+FzH
5Ji5js2aI9ZwdgOtUtbeWguddMOBtv5yqlCWgvCVF+Vx3Gb5iLIMFCYcQK9eZS+T
fQlgnatnAPwk9gbhRfneY6EyHyaG1UiTz4iGJ1ZroULpuhNERRsIyy2Sqe8bTLJK
ZeGRhUG0PMT2/uh7pAm/8DLRidhrht3LisuX8JIOLOfe6RWBrnmv2LG725+471kI
rkO4zKA4C27Pr33HpzAEw09vEscDrNYAoMtxQRmO/dnVu983UzLm7QVgnPQsXp8p
mZyPIclJmDTI/d+s4VZRhf2rrFhR+6Dxp0AY8iauadlSjIu1va5l0B1yr3nQ7hnT
atFFm0l3JgYT8LqQr9w4cKHhu6kZ7CtjymLG/pu45YWjZ+a1vRc0s4/3M7LbsAIt
nqQF1bB/1/RMrejF4KD+ScNdYp6Wra/gpTds6Vjs1Nwo2Ee3fHa5cAQpSMHdTDZs
P6DE2ezwPA4brE+OceGQhpK85T0nh4ev/NmQpUxN+mffwxlc0dIKiTaRc8UkgWen
SZV80W9Jv+mDOH8DS0Q1kbFA1izektA+vf/SnFYNpo/+8wUMLcxdMEG/g3l3bLH2
g/8T014vEiiGShnjAxEBos+CX//Sr0ctbttT8K5i1RourbkiddK2LqI/y8R9MUxR
HkXrfoh8tH/3AIWHJafjlcKLknLk6Gt3JTRcglBVsdYww3dIAX21u2jhhsqnmh90
GkUrZRbKG7+X1VuEg/azb3ET5wY2nHAj+V5kqvWnHriwrt4QA75XuKS/LevqIUP7
58V2quFG+o7OrgJNNwwfAWk3L2dU5IVNzaFFTYIFkzaqXIg7J2FmVJvPWgt+Dsa+
+O6PEZzhpRSN10S6kxFzxOe+RFP3h36X1/Z3FBDZIcoeg2Sl9zZwmO7MHyRXfCOz
pHK1t4b2Nb3BnB3YJ8QlKuR3o/83BNHzlIz79N1gKffH/azRXsaTzoeBTWeltK5L
nelSHDkaz7IQZMPXA5uVVOTYiNfL3ejbj8sPyo3hbKskpEhrhP0HyhoxqzQogTC7
gXEfg/lsZZEu7LBc1q2mDOSNuSJ6ZUWsadaXnF209PYvI3DaAQqd21FTPNJE6Dfx
yfqQrkYpNpRdeNY0cs3q6Ba0HWLr88pYWCzi6ID2ii+sO5fD5hohHXBSzRE5M7Jg
y0bUudOSX9/pGpYWPCxZPtBRzXDyTdkNRNi/nDOoY+qylL3Cd1htA7oWc9mWVEba
oBrFfp+fWd/3n8PMcTmxA3Qe6bFBH9wKcEHj0aBxSUvgHmELYWMhDYlnaRfJXbE/
CxYmshMo5tavU+DGwHixd5fvDgDTBbME3aIcm4kRMhgBfvYQ4jCB1goEoiz8lIDS
qAeueGpde+PghVFGDFY8hJoSWBzEErVvjUvQ56PYO3vuwiWPVn6W05+ytc0zc/Wi
nzdxgSL+9mcFGPm+MkWgqPDB11HwsCwC+zmFiiwZuxRJhSkV/2NWvwpGFcr4GKDQ
Pc/ubGMsPj/3q+4UNNSCl/YxFhIKzbY639Bi6CxiZ3WLClGpV49pEk26s6Y0P5nP
uzGolqQ+b53v6T9epUmwu+GIkRN1lkum6ZsQ/JdxmAmtz3rMYWozbOnkETC4c4bS
AuhYxFfyVKQCxviquAEr3Zf9SOAWt/U2s9RK2DBhpQdJKIHpGH8lbp+04E+Pc5D2
O8ylr2nbrj+fRcsawHErm3LWa8BXlhG/yUlcsVYdechwy6QEoUksF9cE6peUf6Je
SiDthxJ0zbrHD7u1S1kwBVHz9y+c21PqFboMb8CJqa2cRsGIOQVf5iCdJkRAWrMH
FxO2S/aHKsNMDMpa5BnMGVaUR35eVHnCSWiXXAUxrL84sr2fQs3MTlMRcmFbGe1q
xMtw3fU+v0VkxpFUKzIdV4sPne6HcZFUfoW8Y4Xu4spxAGTS9oa9Eil3raObxwnF
F8yJD8UnXlEarKhWOrn4KruS3iRV1P/HDZrPzdwEWRXXAb7tysQ+VYguc3murDCF
J9fVR/Lv2Gq4OKKFQFsgMpHaM80qyeguDGYdP/zKqxzGUEzZjSfQLcIyvih7yPJm
E1Zo7v68FhBOOQZRhkyOVcy37LJ83aa5lebPyQDIArY+qLeWAKQPB2yAO9wbvwPH
cMTJGKfbiXW+MMvlfFrC4XlOlZW1ol1Ax5Lxv9bVRVdvWCOXfvfktuUPb5BMtxvw
V/pfNmUbIeqBSFK72KarwXb0qm0FG1iO9mZeVYY7LyWjS80FWkM2NyqmJ6R/QJzb
+CBP58KiVQUCr5TitwOrM7CZtBw3a6eAQk7oCHN3pnn2z9epuXiv7lEug7TaRdjh
GFinM1C+iD7DgiXQx8dt88GXrf2JkZrnTE95axU41rYY0cIs0TtZpPTD7IZaskU/
dk7aEMU9Tkqes5avR6ISpMh+YaAdf23cPq40LKqUWHjH/6DbujUQODObLey2JeQN
DVqV7WO4Bu5dvdwhfmMl3TsES1VfRw4IYxJqkhlrcniIoCaZVTsfbD0adjMUh0Gf
pvjf2TfmvV/CSA8UCspCwN+roPcWzFc9eDpwhq4BK3pMAwWc1hHbpG5vDYEPQPR4
XOM+6Zs0n4kJSkQU1+5IUEOCdjaC0nD74i7P3QQfVAIR+Wh7GlB9o/V99Scjnb9l
HExe7HfxnZkAWDqv0OfX54HRbtgDXPx+Z6Xf/8vQeLWXdWWkJcMGXCbJstKOUxDP
1GEYnVae7wBzfZUHVx9Xm1dgZ+okDh0Amt/E4+VlyImeEDW43HOSaReIv7xStGVt
xH71Fd9PsTF4qsi4bavInCToQNYrZMEMIUwWK8G4TJ9Rv6tBYO/OBSV/M1NDthJc
InjhXcsjxa0Hox/P70V9vXcfAmB6l1KgzVq00kOkX+hDvnIJhrjYCF/ehH8zd8dV
EXm2jBXtp9jidK3g40uiREfr6hF8R2hHA+gHow7WQjMjz68si8W/4/uNUyvdONaz
lGtVpvnpze/72rG0Se7RULNV/NHIzWnw7TiADQmYc0/ynZA7ns1/rpHiA+snq3Wh
RmrruN5hgLjY+V4qw5SlBubDzpRg3jFgBPG9bJhn6apY58mvN0tyR2WFaOBClJ/n
p9Nx1MYTH9D0Q7lF3vuT4elh03jI6Dm36zgi7hkYNlHR9HBehomxx0+rU/bbTR1b
LsOsIH2TW9HejuwVBTcCA+qLC7OyKXmqbn2l7ISwIecPapQdsnsi/7IKcjgyi8yd
irs9s3nMsrn/EX4tTCwraI76s68O/WVLedcYRkTsjaFb/mt8C1/xxcNYvM4IDMPU
hB8ugbvTByEgRyJSCbJWuObrbhDaZcEwCSolqEzXszCqZmdufr5j785z7jzBBfsp
cAuwU2w3rzoto0Ba5SOl+Hp1nt4oXRFIoP7WfjXmAGQ/ckhijyWFkTU+jT8gNUJE
8iXNme6QHEz9cwKYIIOy+lKpixcNiFfsGszIvcnrsO5XV10NpfMSLym62Vzkuq5y
Cl9EDvk04r9NDv8dE24WWVm9f+9dMz8GX4zZThOmPFHTUfIz+cDvRYgM9jBAsFDq
5doPx8jDaph6PtHLFCKP8WnojuG9ST/vG/men/KS6JLgSPrB/8ql9ijaVH2WRB+q
meweQxnqd8vDa7y3MypCClLOsub/VSOvUmHKwyEEXodyBPLlZ/68MLyNBsZyUraa
nI2dT7FsA1wqlRNwA1emC5N9j4TvxySCrMqLP2qDV7sX9LT6SOP2+tHOka6HZEB2
t74TLq+4NC2YePVFmoRf2NiQDLpMirUPii45FsAV/+B1kcJ39g189i7SibyUAkJr
l6XDuRRs5VJMe8tKgjTim2NtsNCU0unDbRQWMoPVf1APpZUBeJZYfwHUrtVbq6g5
34rZ75cBipOq8EJeXAke9xre7EQtYoyPETq/52fqZHd5nX++XjZhzOCJOWl4y+sf
0s9vNRIYy+gXunljZtbr76tkrwzHo1VjofnZ64zS66LJO09pmlMMiLDi6Gn2GSer
HI4dcc4OD/4LPHG+D9tgxmSLiAvZnjmcPmjQw5omJwTL5je5glvUC4PfENDm5G8P
o0M72QVEOVAgBYRvyvUJnMOwXy6bPmST7mdo1kKaHc8g5KmWbINNS9xASgx7AAsH
9wWp/GOj1Jy6cjJ7+1FZ+FHL8RAzgTWcWU8N4Vt/Dbh6IH+yN6nLB8FUFl1HDJkm
pitcQyEjiIbhR7ogSL58RfhdOBLFXDv9XtoBunjvJOEPEkwTCevjnJUlCh8YSzQu
f45bE1gZOBULSLZqMh+4nYt76VjJXVvW64+00kvCQnB5VCWyuxM3t3TFOTMKvpcm
3p9GFLz0+h+tM9BfXx7XCoI2vdsHZnmZ3GklSPgct8ojD/q9OE+zDtZwsmOhIsgE
+4EAYf9Bui9Bgi8TJB6kLT6A1gZGhoa3dsqshJee1Z8SHrjjEBC+VjYOp9LeUnxA
R1RL7TweJPAdxGSbcwYIf+k4o2Tc5STf2Vh99Z0moHDo/8zplESIIyy3Ob/pp1/N
ac7S0aZyXsGU/Z0nESgm9gTaOJ4/yBB78i6tvPDMRMKxeh2xYtNU3a0mkmMc+Iev
dxN3bGAhV7ByubwZop9Md/6Gygr2HuE9qbDEi80+vAaih8ZBgsU5fFL590oPxzQJ
XDVKT5lVq/H0OH+rqvjjVi9OpHoF+bwRbMxDaBFlY0dQZc8E5m5p9OooLcEqLRJZ
RM18mC2/WhIiKV33fGbsbRPEomuc0JNZem4x3qoHszQrolwUOTqd8+Fr0Lq4VQVE
IHfYaJefMiDgzSWMH8HHfg6afoG5YgmWfCtbcw5dudrw8whYUgmRQRwpUiP9DOrM
mxeaaAWDsnyrHohStjIa3U5iL54FgQ5X0C+szvHrkCsJdFG8r1nv3YVO3udQmqK2
TeoHNkU2pTgrLtkEDje90w9MAx+VT5UEhHE0DHm65NKC2NuyI65WTPjphAM3dESQ
8SLnufpelWMjS4n5LAtiZ21/bswi8rSY+frVAC5RLqIBvYCsmqkgyRIYu5GIcKjz
gGwAqE1I3lml5DjEqJfEuLaonU0z8uecxMIj3UNVhjq/FSxPrjX7T/Md8wSbqDO/
qfpp29piLQjPIotM2qaEuS43v1kercG5Vrc7SXspBp53JWEdtczeOQzugSexf/E7
MVkil1QD+7djU4w+n8++ajyBsbi7RM2siq804/ucMLxB96uHYynPOnAB4IqZAOgo
BcjyK6uH3syJVcccx9tCXRy8l0j1PwgnRSQQ7s6PZgZ9z5gA86m+Urn8NZ9hVW1N
g3Jkt0fDHhceOMgd08UUeJuBXnJ76ZM/x6uFSIEkaZsCAFAGlf33hnGE3QiZz/cz
eHNSXP03Auk5gmd3zYO5SVWFqiOOO6pKucCKxf3tL6lP3StNW9s5SkPem9yXbFJR
jFzd4Wt7VxstX345wt44wH6lv9CzBBt/aCcEO3EfN+rG+RGFaPFJXgSIVu/M/oX7
s7KHSn9IkVI3g5gdiliRJMQfnigkS/brySiIvKFZ1LukLVjQu0etjBVooGjy9cq6
SDezYvUfNzYIvUzcojFLhJBpPIt70WNyrYiRhoipdxo2Ma6igH8O/5jMWrpajglN
Xwc9KWk4ckPdQOzcNvAZglqduSaQtiXD5cJhzMiSe3kdB7BqnxMX0r5zoAJZ3ww/
KOp5OM3nVLlQ+l8EQ7ti7RZuabkJiPzXpPijhvsRsyQaBaR8qpPlFZfehTnZwxfl
QfdR8xHYVC1DLWHHVGWceL48zpgukYjUlZsQOUdbwbPAUUNxSiNKijOoTda1mMt6
P/l6sYVZylhqhnMfJZlSL6uAEQp4s2KpNaTUpOTWrFHv1I78blzDSTPXfiIED4Ax
28f0mYbhmQZbO+DSEdTEtM/4nrcvtunvHPlHDMkthfHK2ZjuHmtva+6bW+9pYw/A
nE8DXDrfe13iJ2dMtb04nzNAzH2uy+jRoseeJWCZtUNuguoEX8veAnNtnPM2RDT+
021wdjdo5JbaMdpAfK4k7mEuTWUjIbCHN1M9wxrDjfjphg1RL+FQ3+sQ/ddar1G/
Cxx4L8jgAHxrcNM7kfcefhSmURyjKzda9Hfb3fIgOXFbacbcuN/l+igTj5zUXF3c
qUf334V1WqEoYyImMB4aGzoUdzzEXNsQEjTP9NcCooZwxUNPEUrKhFBa8TL/Sm0/
svBwipIjHwYofe+8Y7f6JJ3gIOirZgtXtc0yJ/UA6i+R9L0l5lW26uDzJg7CuMRC
fZtVemMGm7GmAtoY/utRoZEn+oGuSsT+K7Ywtf9ixxY3hYlA34Xwg0hRwuB1E6Z3
niOmejr9AoerJ1il9JmNAg3zxkgO52rfX+ui0QtyxTUbDTG56NCmjTRtSiSTcWne
e7qXQJiQMytellnjUotB3co7O550lr7gY28UpJnMqattsdGS6N5muNC1BgRJ3hK9
qgMoP/TckfuXIij6G17bW1nRThkuA8OdheI18dfbPbxKqo/pdRIAi3jbI/sOj+Bh
GzCis6Gt8pF2EXzdvoMfiU6B/bxMvaMdRG0VZhAB9+e3yFuhdRog+YTJ4qZn7rIa
LeMLRaW2PXGeQgAZbqic/v0jNRme23PQJPSKdOx9PGKkqr6NO4VZkcrqmxzMoO1V
pQAMnTzCyRxkSsF33fndmz+9YCL3dKvTUJyv0gTCLWnM8WQ1U6dc/1MUp0jOtct9
QliV55SwupZlhA8YmA1D7SwvzQa52wpjocJYp4dT3X1whu2HDuipqQ917DHblhAB
lZx+d3hPhymNoE6oRDgG8blG/Zom7yWJAIdbl0sdt/tzQ3GM9eV6UoH5tSmLsRgw
JDVxiMdVOHFEy8q4gbrQRBmUb1ed5rc8i+X+yU8b0h7Hr+5Zv9S6+PWlGi8er3SO
Uw9NaJaBjcDftiBFayljBQtmj0xjl0Sa3ip14Ey6pt8q4sYt9EisdWBZeJoBfkoB
3luKz8N07nKCdFAptIxryzs6biJ9Nq68iYddi9BddflRhzWEL/0xYkzXFvm102V+
FL62NOYuBSezXhI1uUOHBpuYj+MRGNKG/eVal6yiqLz95Ij606uR5EkxCufH5U4V
usGZKU2UzFCQZYbk5FJxOJPeqeil2Qmiv9aQJ7GOIhD6ZcD5V4QlpG77tgI/INLT
5lai19kccjvsOOaaIRFMUcZEy7GNvrgh5Tp6fP+ZyKmij4ZrK1HphwXHoUV3ywC2
PZy8Z4z4TrBIWBrTLrN0aMCo//7unNc84RoCKdUJ1C+7gdPmyRMQPJWMxxYdmBcZ
I5CpSzZA7krhAsFevcAuNckqwEB1/29Sdf9/iZcyoVHjwonLRLDiPKgsn/yhcp8c
F8N5dwWrqiZSCsK/LkVVFyNgfIQNcopB7DboxJ/PA+XoPJM2++2ytfYsC2qlOkVt
6ouKctmfM9zfnGCoBfdbFP77p1uYiXWvdAx3C3MASKteQzl8DKOHZb8vzaNI5W1l
aZbIVeLwgxMWxiMX+eGnXmogtEPg8b1ifMvwCReCh9/hmHhZJ8d9k5yJLLRXuukP
U0JutWtk6g4pucsc2iSynYmB+P08vPi0gqLjhSCMemSHhyFcP4UZ6RQCkmOl9X40
RxnP94IWs3clHgxMj+UEJXszzzbd6pgebSY1wSP8tFQEKkeyzDeJVMdelNcVExmr
B4N/hxbbxQW5ONUkIs0+xDNV5hPIT0xxxj/LzgdefBFRSD/zZpcjLLF7Afr351o+
XSuw5kDeeH0ccU+BcyZw2SnUVSa96IxFbq3rNLF5mLg8Cry4KFp5P+9OAzsywZkH
MUqvDJATqb3JIEM8rCyroAvrMylDC+IAGBavCEbAWjrjLGf9DQ7twlCL7PUSzPZQ
T7RW+J4STwgjlCfk2k7DViQYaU8hI+fTnJNPzi1b9IPtjw3sRoZ/wfDumwLCf+LY
FRlzi/XkJsoJ4cqjSywadpdpYLfraVvD04lcAd05SFB0xpkGgeuIrttssS7zHKXb
lxgbfV+olbKoWS7mfYoN9mbkWADAb5Mhr9jM21LxrELbKXZ4KjhM7lemv2aw2hag
f0kQ/ScCSKtxaPsONajJlZhkO56jb70OoFkRR6iERob4BbKalRUy5Ly1UVNGfPSF
xMQbFgWXci57A57Un47g7rs/zvt+xdLI3LWeUrEUB7hRs3FuL57gV8qhHlrSZl71
r6FSve7V1CZ/SblB704ygjiOWiMnzWjO8ZmBUpweBiQScRExSZYe36EpQ4x00j64
wdQFKxnw3uJoucgbp7w8mNtmDCv6gXBlGTKKgLMgMutDtV5To/uj0iOeqqri79AE
aXKD1rK3ZhTT4B/DbwAtsYUc5qkSmn3eD1uA4pnIC6poNyU/+2R+6eqPy5je+TMw
ixOaOxFOQFMX5lUnG5vZ7DnuJ7XR4KyFJ0CH5BQiwyRj2PJGKJyrSbcsVu1V5NxV
KoUICJJNHuVHvMPy5xtJxKkC512PD0YaWahxNi1ds5qqgccOeUwx+dNFMgXMg10s
7CL3FcRifAYH8T3/fWhBOFyDJKNkG3yJv4DX9Megxj/rII6DZ199p2dtaDHWk3Hw
xKEiGFzjcjwjBbScPCaYPQ18wavLIWX4jr2Nc+GWIqui2VUzVjpbusBMJi3Q4HDo
0ZYU2b3KGeiKkt+LXErlDG89xo2g1XEBPs6RL/2VrHRgS2VqkTa8irA/ZTbebQbA
NwJ8y+BTuVUQl5DR4TbWIG1j5t40+6NfCKydu5cuipfziMsFv3u5sqS+H6JyaV7d
o5oEvQ/PHI+tFKX9DqzZZtRnrPliUOzGy5cI9P1573rditIsfca1HHjIS17wzj/d
5dnwzjAsfKlxX9EgnPykwoY51krxf1mp9L/sKfhthYwrMCdJiN434zJLql5ABHgD
cAQr/3jMmaU+Pt2fcNaGeMJIIKbBb9Oy6qDD9K1joUGLuu2AvwI7F0+I/Vuufuaj
lUYSWx1RA2yGVFShiVg858nRX6WJxsvVk5+dsTCQDyRmkEhQq2dI9FP9d8tMOxif
YiyoaENQuo3lH8GZHsWrg+iEZK4iyKfq6yKx4oPBXSIIXnDqIdallvI1t7QnObsB
oZ0tg25Vxcvj3qJadF8840YEGKXds6OACp4yNY5ffuKiDb+nuP4HfBvZm4FYjESI
pPV5hWpVFrceSmSJsEYl2DZWRn0AOYb6536tLSCw+lN9aRrbTzgTlepv6NEj+/07
/m4k496ZPKJJ4aC60+OH4n+E/TySVm2xj1OjiJnWbjy01nkbHda/Z3IXBriNjBmE
5R9SnKJl0snQOzLLygopk/TzXNnCOmyO3+Xo2LUjZzrg5cT3hOH/WakzJnNucN4u
DaahI46wwU265kKqmlAzrqDL4zj/KRjW/KVJF5hMjRU6UoNPnPPvUAQtgug1mK8b
Nx/SoOoRLSaG/wiCQx9yjHPs71ixDqHt33hNvZbkFjozaFoGTREPm7fWrOuhyOag
84GILDiYCFXhqumFltfLwF2yeE3Ti/eikIaaz8gUCrPfUVxxjgkaS2Sb0RCuZplp
x6pUQvjZQKBsZsxRrlZrKb5Gf/dfaTAIXGefhbI7GDE0fe/LQx5a4/y14JbQOZRr
2dKTzqpHMFk8KNx3I60lcS3jClsTPKlSoZglaiJOJaryY1nagS+6JHXaTorl1nzA
x9axa6oYHE9VVV2HznzC7PTaP4JMmLd4b1TIoDeQ44arElzsLgnHnZ5dfj3col4F
z3TREBYibyBzMxpDHjIHAuN2ZTwAwekHK9Wf0uijRau5X9qqr9bWUGvjo3K4RBkV
wP//gTZqGLAzEM5gbCcvCl8lhOs+LRnMIuWzYyO8e+SmlY2U+jH4Z6lr0kOjJawA
ohAdUKIDUxRkNpSo6aUbiEDAc4Y50ue/y168xBgZ/MVbz7ZMbtIJd5xJIIAmfrz4
zh/foDIXWOZu0s7mYv+63di5OwiBcnurd7hT5IKKQJIzl0bHjS4l9fKhwvpeyw8z
W0T/lPfREB52yujPV48C3PXFMcu0QqRkyCaSo+k3rvE5hbWFCRG9gKcWB5akb0so
JrzIMMfpb4pv5tsLwpb1yncxkit7FVciE3HAs3zARa5RKC5Cjm4c8bvkmAHFHssZ
NeKDt+BGlRTYMMbw9fxNICCKgCkxe8+a28kdOZb3yMZeqFpnTYtNPwWk8cI8tAdi
VkS9lrb2V6mPF3FcgLYTnA+vwkD3anWANP09FiIM+GEtgnOmFrqLgJD9NLh/uqVO
QmfUUirIiTKJsFrCO2aYKbPLSNMqn/FJNJvsKJN02UBoOwxWdWPjagyRqrqVjxPr
icBjKEF67NxLGqL7nzCCvQuRJAzWZdlkf31XSMrKUQ4IH1cnhC/1L6QsoBfrKnOd
y/tJNXjFM2MFuHoNt0InQZoB6So8bUW7YCtDiPf/3wo7V6YtULq8eT/WeueQsGl9
XqPLgNVJUrAIsoj86M8fOqsEhkdD6Q+nu4QXRxlaJVnsk7FgVofI23juQdb9tmnz
6d8WVP5WEOxpGu175qnplZvZh/iAWDmUG9ptY5dcyVptNIM1SRVX65sKETMiyxss
VHzeYVpwXaqxo7738iCi2tjGDCgHTI/I9ZGV/hEqLxFK5rPd/gO9Vtbd1Z40kXpA
66erUAsY/Luo7lbOLAYnir5wrK06qCYVbYv6R3z8Vh6tGYF8ULXM1EVI+snvQOEs
9K84qXcoqxmfLYC1bNTjMEityg+OsbZyh8HBv/h3pkBs+vuL8b7jOI67R2+yYO6/
HYZvWGjFtl3kr9jZ7Q/PnhH7x+jK9xa3cRv60TjYaq3H9Vf8hcL3SS3kS+7FplVR
Kna8T32Coz/ZScN8R8JNBiPPp+8wae0cio4IY2LbHjW+Cw74zLadKt5qGlC9LJbC
lVLJEniT35BbxEfJK3MIHT4cHAj5g/hKArKbuOmTbYW075gfpoVmQbi1bRtE65ef
KihfCKia24pwQUwMIKNJ5aqz00S2bhr1dgUS1+VX1bIfom0MjJLuZU6iBuGybLS0
HxIxHt0GoPSZXHkmKjWG31D/K4on1pSp626xbGxo/PvZo90pI/eZ2L9pNzYlAUj9
TeGh8LOrSsS3fg+ntNN/UkxrYP+iQNpi3Qt4iWsxOte3vTCv43LXT0HMZ+0vr5CA
9KERB80ZTvS4EdLYztGAMs41CJEBwtn2ttN9RmSQ6x9QwJuAYJiRYabD/2Zj0xnE
wcx1W2dOBykzPQpQPhR/QVzfsSjgF8/cUKmxyv8R+nuzuha7fuf3D2eNhIDhUbF6
oQ8Q9vsX1l0ziW4PWLYi9xaT0rAMx746sDpBF5pRqv/6rAdFkNLV9RIiZUCx15Ov
B9wOnvikMZUAGlYqcKzUUfBUeZIvTh6Q8dvtxpASKQct88YPno2q1/wEI31JvRdR
m79oe9Gt++CauxkiC7areTjRmVxCBykRPgp1v48gdsgjE2KPEhxsBPxLyjfbPU/S
nhwF4gRPkZvborET92cSKsfBY9BEB522LqiH0Wq6asVFrOLPkKSnKayVdQleJhU7
PB5XZFteiW5/U1+IX9aXbOS1jREMr1Fz8VukoevXgIxv9nzfAADFlpZt2ZIB2y3c
zB+Cp+2aAAbdMYILZ6AX/RmsYHWVD96tg4X1Hd4g5YJyYLdZjCReD2k1+PzoACYE
2kb1yvKhqvsNSGpcYcb/AKwjAaf69xhs57FqMPgAh/kRb8QLnvbNYnHajThMrbNO
InnxoT8doiVnhs60v0SW9CQYYV/mOz/JQiGr23Ez/t/VoZ7hOzHC91FzYyBOXJav
0/IlBG41zT0PRB3WfFyTHrU1J/yTJRBaoyJGnkdjXmZXRRi/3GxWgUOfZ1/6HfRi
TDy0VcYJkXoPfd9ORoeouF6jvzTd7frWdL9QiC+a8Yw7Kfu/3CTSBKGjmyapiKHU
56vQ83a8JWAcJ5RzAhxNuRpb/koY/7Rkdk2LdTgiZWk/1WCz6roF5JLOQue2bKmv
/faL7BPfdRW0QDHRzBKFjyFEg9sMAen/w7cIVkxCgUF49h+eMACuN7NSVTnJss55
a+vi6dIlFdWMYFZYKaeS/CWNzGnIJDvTD1QmbkakmVCB6H8bHZidzAHFLNTfKEPL
nIs9TGiSXrxflNYZJTlSriiW+vcOs8Gzc3Iak2LwkPkqdWTHejOqmgcs6KU0ebrb
gmZiWgvPvpZf4e/w5Q66cSdGWtaHcjedkUfLguPlrwr7V1tmsWePo2QUuoDdgnEr
F6dIu4Y4z7j5yuXK4qv1A55b02YYAA2JC2W9bZS9e3xfkt5IOOlWlDYDpk44DL4l
hnEdDTYrdQDKUF8lzShAdvhwOP6xfbh0YuFE0v5RVp+vMLlj2TT5x7zQky9lkzjm
jYuWALqG+H3ngkNPdRRGPEWoRas4/IH06sIIs2tzVob5n8UcxCC2pD6K6lH1me4F
TPfX/gRNqtAq1JizlSj/K0jStAyhvQzB7edJvYVMnvCAqe4xVt2BGA2aILG+1+Ip
K6hiWd0ViaxGD3JdDBiVXTEiwtQfALvlVzxd7FGX/kQ5DbJ3xnbPYsXQOkN7yOJy
s3f51BPP8pM9BMSU6dT4IA4PP0BusjJlVuwR1ROPx/K1Ks9NSpnWVUQQjzaQFkVr
IMD0cZb+K7GhaghqE68hZLitCB9asQ1DYsyhcjEw8Iyl8sbYiV/cMjNTUlKOOnbT
3G1d2wwQWXwfCHN7B/nOc6OMNsnjorOeaRWT4Ykpf7llIezX2+SzJdFo8F5c09Jo
Ov6itTuoaZacRxglkGke/ip0KTW4PpVhKnXvUDHlTRQkRMtmLamo5ypR1TGDfteA
OpGSBsXps/uhMUiCfTXZT66TWaqoMQslr4t9omq1NpgedhKuHT/QbsoBBmbdv5fF
v9hzwPjSVVT/DsH0FsRbTVApb4mUwxIayyE20g6tzxZApVvArcwE/fH47L6YFdZn
gVM/HV0OnDbWsyiV/jozrr/VOcfMoVJSjGZFRIQoqpxe0V23UciITpd8QiqIgQy0
WYHikT4E+6HtneDilmg/Ky/2godEx/NIuPL0OXYfTvasEWIHg1+9mRIUuwYK5YPN
keAAR6rmfuN6LErMv3CVpsJ5AjlNxynbXFGU+NJDZoujEQl0kMo4SejTbzZBE1Pd
arQNqm99btfigVw0uicLu49xf6XhkDdIkhoIm2BMJDZtlUvMXTpJ1oG6zeUkHuc+
qtFnFJcDTEOSQaOdHZQIDzf9ATbhGgMRxgKDfck0ELF0iW1atL3sx73dbfCP8Qp/
24OnxQfxl7tZSip5OvaR10iv5oVYOgjC7bsRgIhQKJ6vCwpzvG3OL6gCMhKvcVCY
OcRY2EMIjYwqEesGPbXRgGzr+K0rGFHIz7VysRTfhclgOJw0AtJBJ0ZPye0p1tp0
68r/F2wfpNoZbApyXk8FpD/1kMilwu0xYJ8didoKBixW/Ycouvim2gqFgG1Cuqif
aedYvPL2iqIlEMY/r//V7QdeeUMpJYxsSl1x3INEVIypTfyTXZr1uJYapY1q+nHy
LrF+gf1FRgsuXSl8AJM23ve4qwx32tbwEtWpcH7ja9omENXaGxnVXpJDdQ1TP21J
H3PN0K2DRuzBfBOq5RXbagU8SH0hgoJaXS90Z9Mqw4MK7ZAvGwatSGF3IlLpF/gj
er92SLuwq4jaKCAY1dlmEydyr9ZcLNx7F3dSE7U7n9+Kxn6dgRvlveSSVA6v7H5y
QVr2GC6+8GkBdWaC4UozzB/gCxSNQb2Bifq/MAAHYQ2D3BwIkj0KY3xkPx1qJMfc
Fsn0CLsl1l4UYJMk4dvsCQSpEd10UQP+6FHWl9240aNd67ewHrkXDN1oHVnWLMDj
MzEp2zjn8Nc3C/zpKbqa5/g5BbWTh/DhjDFNK7b2jEzv0x7325PR4Z3NB7/cs/Uj
9m/YXEMLRXV7I4GaV3enMZV6lenOcTMXZswjCs+cTkqUEqSCahqSDpTh1/RRz9F2
yQZ8xPMCCNjg4W9KnDtcS3CbcT7+Y9PrZpNQqc7916VGK9N3fR46HXZe8Jl240lG
PyMhOIrIDzzfM+xk9a4l/AyQ2XOlI70OzAK3awoXM6ausJVUmuKDy7qDGHhoNL6e
SpQV9MjmdK5MArRrVa/2RgyvZtRZ6EUpX/Pn/KK4F0z/takl/qKZZzkYwa5UM4gT
rTNkipxeDXODdBLfaSnuRRJe6JA7hjQ7KLjRxecRDDT7FBdQ0TBdPzUjJNVRua6/
4FmEAfWG+RfCLloivX4x4AU7uCL5eGjoqAwhSZkz//cW7+/ljWlSzKLWbDcxWx41
jexs0Cjwd9xBvVJeLJkhJp1sUyOSuqAwUxOEKX1VFW556xyif0lMpNQ7vSwQ35Da
kFbhdI6yHKQCBdPGvqslDTW+aP8Ers3YzudiE+c/L2jZmoP06EP91cEiP0Xvx0xl
QwSeY/MeqORY7SNtjuBaLWL3id9K3vXMMNFLhCV3GHdtbFxgvKwIf24o9JJMWNzT
bSkL1Dx2W8cIYpMa24Xct1riitAJrdDoQgIDFURjrZAKuWcQRMAiQ3h1Y8+SiM8w
TBgQ+yAq6DHztH1lyjMKiWeSH2gMhZmNDW8lC+mV43kwCcju6X5ovvnajAHK0nk9
8W3RiajG9waxLk5Mo0WhURCuSjGYsJ7CT9Yw0nACcJgfXh8/vNKwT10vll7VH1u+
P/ZAtA0ktQQDfvCdwGvwIz2Arp55Xf6MVlRMxWhao34i7X2nBoCagsM/JvHdb1Y8
pCoJB6BQK47L/nsriLgAMlqUPd8GukH+fVQ4LZPXMQhDtpt8fRik3S4AZNwGNsaj
KYtmJVAucaUNkX6kfVVL3jxA3lOFGseJEF81cM2Gt5eY04E/bp+C3yodR1It5q4m
3bazUCSVALuHWIadIAB5C+m3VpfEWwJDFBb83S8ujePq/L77a5GV55tq864ayU8a
caIVYMjU+kPDQ38dgyM8H0kqqqo58A3kcrcEuLIDcRUTyetaLsfljtpsNZRHu8WZ
Z1X4MQM9lUjF9S0ZBqE6hqGy3UOHR0dLwdiykBdLQyRTDGWyYdPMmT9eC0v9pnq+
TAtsWeapJKfhpCw+/KJltD7xFr85p1LyXi8eJxT1/rU3ivFjKlH+7OTL/WE0F8TC
Bqjlh8Kn6quK66n13eSyZY4yIik/QHywZaPhdr7UlwaSKdjoDOSOtuowuRUU+e5j
jcT9l9Ql8+Xv1g/c3Sv86u/IQd9SWvlaH0moLCwI3esoab5BgFpkP5cLDWhto7AV
77QzZl3/kz1x45JjiDyOGVH/c5VQySpkih44jg3bVDJnVfAb4//BQlTmsSiaZIIy
qwd9/KRZMmV6Iw3MWkgyuUefupaIy+vF4IysSKOuI9IqA5CfQg6Hhm55QUdoMnSf
vK4yhyC5k27X0aarN9iRlunH5UN7yzLC4tpJ0DKQlXQxXPSqUgb2LCEQexNxIS/J
OKcq/zRMB3mZ/45K6WRqF4M2L27Vo6BiW3uChNCcZuKZ3D4IZjZjjTECL8Y6l25y
Vzm8EwA3gnjL2Rtxb4OYqsbh8ZW5DuX2jyB/rc31pIv6Ya71QYVbMt2j5w21x5VM
ZXp7zJ27pTDbIYCGR3WlHTBMhwrtteXadtlk299jUiIFffXz9ItGOJAeF5npL2WL
Pf4J2v9uHw2msu6AnoD/mmv8HkDU40xCyCRBJWU2DtkhqS7OiL6dj70RmwdHWVGe
gsBqQKtWedQVuck+2DtBhBSMamHoEHPUnNK+GIcPdNhBjExW81M6qrK9NEuBAJQe
TX9/X6JKPYaw4S5IwH1kxW0JRfWMP2Q3kEHfeLjsYnrWijLjusnlu2WflEla25lp
wPY0pJx9pI5wmr5PwqE/GOxf7IP030G79/9XMg3Ri1+dPRMVxq8FdfoxbAjo3zLp
YLiQp6SKVoOaFaYhhlH1i1aTTf2W7BVvWoy4aFYdxU8gXSP7HVSFNb+RJb0o5wKK
ktjwIpW1dMDSjfzDCGrP0WryeALprSEzJie4nSSRKUJGadTSC6r5mjIMuC/Kmjr4
jN2MkjRuZVVx9BJvvE8A7uF8+wHeRtPnjVX2/EtUL3zdb9spkmF9eosB9odlRkNJ
Iw9uSDfj2/I+xK3Pmg2ASICHlXna6Yy23neL0/iq8w7tzGbxlDKcmVNZsgcPPKdF
pKM+TqKIQT047NOo6y2nWKk9TpONEgfXQjdUsXiwPjo4Rzj3lAebihJTmydDNAVR
x2nZZcLbYoIBqCFf0c4Pi9ljWQ4MyTWurdU8hKu2CwD7Ea1bdpAm/cQzvDmRziJg
JsMTmiDsJzAWcZ71Nrg8CEaE6CBDO56OQDNhE1NCQZTzgTdu2MK8OdG6bHAUi50j
XW+VQpwTEoZwwJDlPq6mCwcYgLRdqICzDiPI7eJ9X04iiTkSKW+77y0J+IbVMQZ1
HpW8o1jDXxjuNguIgML8PhEaAR+Jnd7DIFMrDSWEC1B5vWXyL+ZfI3dhIQiQENyA
48oeY3Nkpav3Yw+7GMGb3Hkk01n2DaAUDQMHh3iK9t7TJAkFmpon4n4T4OnrK7hJ
OfGMUZ/iPvkXguO4fMbJQpuBT1TAqNdxMYQhrWawWWzPl+v1DYl+O2aCts0HJO23
gdSEmj3tmgiGVPR03HwVaY/Q3sb2F4+m8YcMIeJBAVMIADZ+RtXn0jSe+xSTvx32
8hoRZHw0Vy7xaH4inM+UO8R3UYKffjq1Xzg37gulQUCuzQFkyV5NB1uXjjakJRs6
S4Grmf6QDnMfD7scxMWWA8f0V7P1hENaNvYXgu+Bz+KJPUeQYjXYtC47Of/iKcK3
086GsKkvy6YpK0mQ++MvlIBe+jX3Wz7e3mmNBFUS2N/XkVmuZa1dq4ETVxM7DL11
J9UR2w56DouwFY+S9tDIlxq1Pz2MwT2arNfPn782RncWvVLt6inoY6c9Px+835M8
g5gMW0D9CziuF0ySLNDqhsc00LjeieKBQdVD2AeD2srR5xXNfHC1cAV7U7PqDHrC
G9txv825X20lAp8H1zFNqHfom081wuLPZm5kTQDgBTl+rHZXqiVLTy4dfHCKWn1Y
FTxYx0GSv/pKebaEhsDgyZZrM1r05zJKWKMWDKczgm/5f9SRmvQmg9BiVBDJxpy0
Aea+XSdJccJulQN/anpkuARJSseUdmCqugGlPWw0jP2vhyPTLn7W32b/zu5HBEUO
oPIYo5WvGmWvPny0Jk8OywCXL5Sd/JrFtpsOuI7+tQKaOlNvgqHD3B9FvsAV6nGn
EnUdl4Wbsn9Q/sEsvONkvVwwra++0O4zeQYeZHxsR/o/macC0Jtz4tDor6MBBmpu
/oztdU6gwrf+FVoWqIlvsXXe/x6fZoKQjQIAHjpvjYZSaysJndnKafvB5JOid2wJ
PwxH1eL0TyYpiAvd94G8mfII+ULTQ1UqW4ASknQSj2sqRZeqZtHfLym2lhSsY7Fx
a062I8Lh9o16ix94+IZxvOWWw3bTvmkixFMmtxsNC9EjR15A71gQ7eJiG+/Hh8PG
fxDdkN8zOt+oZKWTj2OYYXCGlBBjboibxmAbnn89vTBKDL9iIHBbhRClz5yka2ST
d1OjoXWGzmvUy7FzdMxhc1kJBfsk6JdSjNZ4T7zx0QS57+UuzVM9ZZAZl3CiFdSF
Snju9kwY7uG4a3G9pCuOrbURUTHrz6OvMVsZRTSK8kPY6fwjHMf0XziL32FXePY3
bI5fOpJNLsOXoo6/RomB2ZXpDqxWDxigJEuJafHpcte7S+Gwvj0lLdCI3Z8+btQd
hovkugb57g+i5qC4ZdIqUcAT7No3t1NZnc2v/MiAtjFmB+sBvREWfrGbINdvLwXV
edMhV9SUwUt1AiHImy3TnJYbSNb46IIDn5vDxXqw6NypqpX0/4J5eqQJ6jCCFE+f
TsHMdN8fWe5BpB+w1aDLtWTswnZcL7jk8ONvcJZbaOK/6bzgNWBm0yHrNVNt747n
wczOt9lzEUBgQVF9+vriYLb5topuQoSVgmptgD8jkrwp3nM7/bYkqDUwNNcXxRce
FaGOJt6x0xMV01wUahpR+OVnq0cNVlgGuuSyBMmp/2SAvNdkhHrfm4HkLw3G9Wxo
9qay8IZhrZDPa/ZKLD2VLsul75xfmvDuA4V37GN1usW33dss3OIyU1HMJ3sxKZII
DF/ywSrEgLtK2rq2h3Po08T38tuiW8+eDA+URrDu6HzwlH2Q/K5eoqRzbPlkvRa1
Zi/3ej4uFgc7dh6CBW5mYw+eLKlae8Z+Xal8Padi9jAQCR16YFVG6eGHhOj39M72
a7yDm4gYRWWW6tzzFnwGNGhhGfLQGCIEBOAKiuGH/a+fBorHgx2BoD/9nAJ5rTXX
o0FXgiCwbUDOGsJdjg129GKUo5+WY1ghAkFotW7SQ8l8DI2hFvV47vf50XQ24j8l
2ilQ6aqOaBJiF5ZJJeyfhp0OqTVkrqIoHH1RaJmPT5cyxRf6KRELrNwOy4AJHexD
tHtHcWNDMUDVVXNdZamMcJkogaPn2eLChxiVHGULSR/vPTDUEm1PTslnmptcYqh8
SODoGX+RGuct810ESdNb9J9qbTIds8ASPqrJxkekHOYZcemrr0xwpSvbf0nSXlGE
5cdtOqvnzKge4/SYVSdjMsUj+eOLdwAEEhLBeCU9jZkZeYh4THEt2S9L728AtIkO
+mSjY34ZyJebrDTg92Ldxeezu3GmrRjSFgMGCQOORdRM229cKHHbk0mUY+G5rjbJ
hOuCO6y/AZUrsJyO7wav+d0bDhEGAYNxnvnFzivnHF/ND/bfon6fsVuTkf1259/1
aehGeHI7rks37zYGgvUpu6O5QtzMe4HSPd6pX1NGgVdecEjWSNRkoObIdG5gdKl6
ViVHrRCDNRK6rVgfcguD4TwqZJiTpwAHQdIU3SbivtxFOO0CtGiecm9vBKlxOs32
vTIROTYPYvnlf7zneitctJoirKLg7hijEsKw5D2pULWLHpuSqLRzQvRmXuj+wkYz
sWS99kH5OQ4omaFheAeSzn5g2fqaZ/EtKxYg52t5HbMzxmVQouMs6vL6Ymi8kWiW
B+svmwWiet9VFU9jnwNKs2ge0ey+p+zXhIEt3i56qXK9OASFRYxsF82zPtU11vc0
s8Piuj+q4ZbNJx1xhzrOb7JQl5zfuWxEE85LWqSBt0V07ecc2eCbRLUUxWGzvP/5
t9SZMyvYV9qPMRAK3pW738g0MqnHw+CHu3Reu5UtT/UMQKjTNj8ynHtjY5fH5wY/
Z0U3nQBUG80n+NvXC/AdLjbYZ6X1V2JRbhmu/6OFifwGKRDP3tcA34fuxEAF3bqR
UoqN2Z0gZ7/i9WBRf/B7xElSMzXofWYEAuVdM7wKQoThPW70pl/5JfQaW97jajbt
59mng6N6SORThGaMnPq3lkhedkDhq1VDM187CEDmksG+v5dJTy0Tb+gmBkhUkVQM
PsMwmf0+SgcA7CEHTPRaKJdscUHn0RJppNdgyRgoA5/gcP5aRZvPVADD2UUIkbkb
N31iLjV3rzy3Ttqq0lKf2fHJtJigRizf5KhF1AlFZh1MaOWkopS6+/nMuY9/x4Og
9YRSKg6GGG+/bVT3qYzkZ1TlJR9dAYICwAOz3wNcOZbn68Dn6zbLAiNjB+t+otRP
ypF/5yWwlpzEE4HKMbEA+pKcFTmIBfJVe8CmOu4Qt0lgSJ0Auq+Wy9luOD9Q39Q/
c4TlwM9mDFHjLXe4EothSwyNe6wsDCB8KiiI4+EFdOMQC/HfuyFC8H1k6N0KHnST
OvSi10LbnpKEsarqbNX896Gg7cx24g/wPP/UnEmyygjhfJxQiNwzCCFDRanOaTLG
BqZCAyZjdL2hEizODPgfE7g6+U4lN29gMto180QksCw47gJVBdGg6Jd7CpiOnu9F
i8oC4teG3sUrhXSVSBpsleSye3VxGd0B2/PtpyM/Go4QbLf57ADhwrcW2mvx195W
Z5RN7jyTyi4sVk93y66TPcMRfeHa9OGokYbxxzbKwxVmBcUwoRx6YCwybyo8u9XW
mcaHzqkjGuaTE6UW76SSJNoXmWyVGdixHj4ax63Ley5d1umu5+vfXKKyyDCl9v8J
VlGfOGbFJEbngkWd1LVT6IS1kR6iAZf8LTNb+KCXgwjswUKbb6eak7iSmH2Z0w8d
j7AtYzxlmv5AYCXpZBtqbycs9mHVO4YKnL2QMTgojj74aUDw7+seES2KIoct+USw
M1YE7suPx4a96JL4JjLY2oI/pq8ik+XenIvy2Q96JZza8uZGN0Rxl9xnHnSbEqG6
FD00AUVat2poR81RoWx1WO0gjcO47X//RLcs/F/lNMB81KFyVjsiLr3HJHELnw83
22TD9diwB+vkxLDK97uf6vKspmqMV9n/gvNzOEclFAaRSZEiYSPvvadoziNuAERt
20XhtV7IUs7rzaUIN9o3axvKEqfprLjysXOmHnzGV3qU3GQGsNp2j91WXnE0v07j
PuGV0zsjRh6bd6qThM89dAQQYh35MI8w50cSnhYn38xhQJu4ttkLzvncgRMKSxK+
AELqMq4w4ao82INycE7iczu1hh1m11bAoB4rOtdcLKnFW5otidLNfymXDtbMK0ei
gaO9SZi1WEqdtY62pdTeb5We+RqSbz65MdPJdzfYt1TRYm2S11a1PHW+oBZ6bgVF
q3aD2fHxD4g+Ww6MJrwlcOwuLQjxrepFnMMVRJDlk48Mh7ozJxEX+F7ow4z7XKuD
4hHj4kdnjZH+7N1HWOZSGHZ82IZpqWZqInHLsnwA1eXTmPKjOc7ockvWmYyKf+Z8
p8W7HLK8xU8pPnenWccc7+nGS18MpGngVnIdPccK+HlEDvTiNkWk7OCEoKqtMCWW
eOPlWqq+2+UBZQ6MAjhzJodpmDPdpDYUOWsnlCHusVyjot7S+dBANsCh+ypmRdeB
WYcPjejBrDwOB66ueDkK4uJyi03r8afeeSIY2TlzaY58gY4wbfygXbztwM2chgmT
XUwtDZnPiXik++X7Vfa5FXZQxUEAamdE0DtnsbySro0m5BpQYs18Q3eIZYFsr5tK
iUTp+8a2k4OOZhdy1/UWAJi6IVZaBoBctu8OXmpFUwT0UhWJlijeSeMUfp+do5a9
fLWkW1KV3KZuCcxDbvDOSlz4W1kZQh1NgT5V3psbUjTGdFG5oBJu5iCzw9/Sukda
cgcAeu0+k2XLwSvsaoAk082Dx3BdZyVT5w9bRbEwrTaf09SVvR9qDDC4K/+IBk5p
aX9yWgjAuA2ut2+SiVeCIgsgUm1XSFrDZMtK3KDwZzSyqY4ssuStYL0GbEERE5Q3
pcLl1QykrbEPelH/mEdetaHsMcQqicFrAwIpWES+uHU6qHOEF8TM7CQQV5ByGX0f
R8lMx4NqB4KbBjk3qKJHQkDxpmmiVMdkUePWhD4tYrQjUAl0LfDA4lL7zm+Cb19u
OeO4SyrU3dADVRdnaSDZ2CYq/ryW6IOgNEnItGgXsaHbdsmCFBoUsMWiCRumXQu3
7UEz8wjNgTSTTXXpm/LEuaUgyjHFAeieTlobuXVA4YvtFK3Ig3aAW0uQeZ4W1plN
daBGLzBLzHLdigpXZ3vSQqWHSivvjBC4vB9B10BIOHEvJiWMLHRG0psgSZfELKBY
4ZGFmpZyipnIHwjej8vqh0DjYQ9OonnUwe6OIs+g/hqs9A0SrL4iyApVUo4l1pW5
yNc+auL74WVRnPL0hLYiaOtxA8D2yh/7JVTWIgxuAOasCcXq8z3wrnJ+8VjW20aU
Q71NSNvZK6X21FrT4wOBsdYtrxD/+A3MW7Mo8B/y/bYMCYNMuFeIetqKSg6lNGfa
NGj6u7Fk0VAin22Mhbcwhp4fPfuDeWEgBbyDuiv2tfmXIc99tmwB3ic2Sk3sW6Sl
bVGlszOcNNm8YZBedzEBilxFdqvo1BwIR3wVtlfXEHg8Rvel2qd5fjlHc7ga/N0r
xFBBHjsX4B8tb+n8HB9EjLVTqtufuvwPATxUuL+2laOk+shiMFgDsNm+ssctLosK
2KNQeuMqDneVMC/VXQW//nIXAk+ADVVUCWf/jlnEc603hAZ4qoUaIU4IKkI/yN1B
X6xHHk1R2z8r3cA5vc/zQjhlrhw9aCyM/sLq5bjauXRuB88JDkZBwa7j4p3TY404
ecrv1divrJIH/RyKIiCHuRf9ZksztjXF+Jtfeo+JiykgdVjNLm2mwszgduXI8OeR
qxEtOrBGJVGdDTDWtaw5EFgPcqlS/QLahhM2Sf6wIo0sCoTFhgXvkXZjxbjubw8h
Cj2kzT+be0CJW/pYqTAL2Vvsp0Hv3qIEXtHNZPxsaxsPbdPv3tulFG51qU396dv3
//JniPyaVAfUJTqdjGpi8P+ac8k7vtdYJTr/rb1Y+0LKgO/0B5Q1j9P7lSmFdW2D
6Mf2C5wzCm4jOK9nLz5UDKugGsxPlscuZHAmtqJZpU88a9QXjJsKpfyguRRHWaaa
q7bS4cJ0HmdPimPMP9Xpdrl8qQtqjHyFt2Ne9TGApfOfOIt0XFlUTJR7guVI+UWl
q06fWk7JzxgNqDskKZwDKzRPYw6q+DkY4FwQY6nP1VlPQNCUbAogdZtXb1Of8Xmo
71huGMuIFPP+yHjmBFcVZNKheL1ViW53Mp5mJmaiOg6NQ5iZgAzk9Nn+t7Ng8o3o
UnwL+IizHOOBDSX0neL9yNOGXYOBQK5DRU6aCxGt41zBHqHpq3qlv2I1QwbqoKVt
MalHAstggxJ5MReRT6BcPlaYAS5UZMe0vSjiU+xQmrydauwWT6unLDvvjZO8I7pX
bJ2eM81J0+zsverjAgM4ubL7rtXR/J7dKSkif7oXPaierA8gsCnTEjb5uTBlWKrn
YE8B/elC7WD5swfB7A5tcCkIcRQPZFC77RrXdJQJahSqWPlSI6ZLBtnedbI2sc9Y
Pe0uoOKa2G9QhTdaujprMQ4ZLsnAPFxBSKbMV53u/V6k4H5nLG8j7CxxJfR9FtKd
cBAvizY70pqXEyyA5UP3MRxjdVQ/v8/lxSYKkkiBb6PmcALLsopxm5l9kRrb27EI
3AS/V1QEkqY8G1AoWmq+WekPMq0d917gnEnqL8qz4oVQtKhswOyBOVnm/bIRbIx+
kI9aFdcrs1i+Uqk83VWduNvQUocGF0uf6qmzGAQyoqOXbg3XErZZjHsoGn1l09jX
Z0TOw2dD76VLZJceskRYTzORlB8J9qJKqCaTf3msXxZZmDHFl84gMsf6LO+7uzPY
HryKM6h1eVfME4zH4lcOnLmuhdSFKYEt73EXUkJ5R2PLO/1tK6h1Khs8lMzQPvaL
I3mDXdIh1rqb+iqh4dimgHPWl12rXaCQS9oT7DBRCn5t79opnd/TfOpVIy+gVi/j
1xBhyL7UDok7qanJsVgxdyF7lHkVpfRiHRc2kqbF9NJtl1exapS8R9fN4ETrcio3
tI67w0LKkASM8YZXDc4MUqfF/5SnPrjbShLiufxjbJt5HrpCu6Zh9yF70n6v52hP
o6XcYSeg6cVpF4UxF/eMvBBiEIrvrX1rNVLgMIF+Ih3hhxQsDkyRycxoi0ZM5Z+B
B9e2tJriYK3/pA69zvSjcsOsqagrhodiqo8SoPnyaKhS0FRx/tQl7jgsP/WPg3MH
oRqZnLT7JyRd0VbqhwjPNU+wcEuAkSUSh9pUu6mgjFZC6WeHuyvUuwH4RJTX6NC1
PEXV9Ls5TMUgOOX3kcUTqCud3Yw+rQQqKcSy43xXeVt3vyjmq3H8iHGJHbGFo7t/
vb4QBHKzAOSDyQH/ms6xA5nRqwEvAzaJFy57qxbRftaA4RGnM3Wu96/v2RE+W5Yx
d0QwKx5lZEGk8vc2qfKa3Xc5Z2KcjI+CKvKhBxbAW0dpomEaxAeIWS7Zk8na1X/B
R6S2zL9158o9eeQ0Rw5IYcG9Tw77c+v0sm2cHV81Rok35T5V6uycK3zoAtembF71
WOnT6k6uF7+75NAVVsG77p6rpIUGpZ33leVRM/lmW6fKXV7Z3+/gss0ko+QotnGR
QLh016fa8ksPP+o5vt6srGgz2sJe+lNmB8aYi0UlGgz9EnYnP2nbWM6SVKLKiSiU
I1IL9xz8c1gdUcxCHJTNQe1f5WPiJNLtrF6LvarB890hK4GO/zYxcsx0DVK4zFYg
lGS3PTcxQ8DZPfT+0KUk3HmKs+ij2SjZxtAPeQdpV5rh5YJCgUiGAaQTRb1FOJjY
83siDECLhvSrjhuTnmPQIOHGpyocRw+dvDHsSZ3q/qv4dBGbAISj0BQ8+nVbzqVp
wcj+nYQ7zSW+uohArNgLU5ReLK4ybEFMZ2hZuDxJ4SymQ2zR3O+nZXHYQXD80tGo
s5OgGuTKG43XeoBf+DOjQZjp4ohORJg/rECmdM6/UCa2N7ds/DaLy/ClUYxuxF6b
unev8Ctb9NkglosTpQ2OyMo1ZbjTxaL+1DI1V8dmEdp47ybvkRc5kF2YdaieZ1iz
mnWGSaFuxnjQIVfhdStPwCe/8otV5CdmcKNjkvp1NgtdjglHD2Gm163CaTP4Dpe7
R7OPQTedQFKrVy4XWyxeIfN5esPUsQZrxJHmBMkCWu5peq3TxzKoNXg27i2jE2j8
UfCYixNNJFGE3ftmuVbyYeYIC3z7D1mYPYCBXdLAJnZL+Z+D/asYbRFHivXYSI27
b00n5BSXU+iJH/ZmcZ2EXPODS1KsEnMlmp6UMtHhS/lCkgqWHPe3U8RPXNqpJMai
5izyU1QoM/XLD0hMU8kCWgiwzCGAyMGXO/lOyted6p6+7d3v5T38tiRDWntG70N8
vDUr2tQ9eZpQggV4Ep8eONPIeDAktYSZjbYnL9S0sAjzA7ewPTrPT7u9t+a6MAP5
idMycKglMhRATDDIU0eCgtj/1yPZjT3j7B4dHaqtQY7RoBud2h1XAJAqlN/FIXkJ
rz8x5v+WhkeL/KDYB2OMjJZ1cyEZFzvYNw7/6yIkrbBzPeQRlG+KOPYZ92CxFetM
RRMKmNC3V1D+xE27yabCNCsC39qkLrofJcLz/9/mkSZ//zsRUk+Nef+vmvKmfH8C
B+3ywR8cxpepZpI+l7BjIbeiDrC6Cb5o70ymhnaHX9thRSIXaM3fVJjgnMZMwiLv
NHzhQN8UUNCfgRd4QRzzl8NxWMECHFY9j4I+UDHZCmde3jt4vnLrK6rW2xlXBZL1
mX+J6+29wQulAZyqw4vK6um8btRk4CGY/wTcwUrZA6MDFflppFVIOiN7AFWOf6Yx
4zMilrOLOFlbCni8E7As17n16nlILxBk3ETkOqkPpBnBXDvjH0F4wooKVbKzKeuq
XJ8e3SgWyL1/eLaCPCc90IXo5Au6tlk2RZQf6qapc9jeyizxnezHqeP3Umz+M8fo
Bs2Ceyd59MA2yroW0tpskiSyIA9OmEWvXV1k0u8fyHg/5KZaBiy+UnrqlDAUL7r1
SFqaRZTcVF/do1XYkq0AA0r6dIh7jp9rMPRTXaI/wohtr9bZgV5w8e0L3WB/G0yp
WykIWGQAeRqOPS11ZRqqk9lQ/BN8b8vvmzYtqjLEcRGlMI2zYV3pGbShQaaF6xzc
BJFt9Y1+GRJy49RlL52NCwUzlEQBWaWxNuCzWD8ddgf/Z+4YxBwm3onMlw4mO+pJ
9rvUeuvHm9fPENyRHinz21NPXA9AxNE0ovTMvpQbeisQNC7CUDwZ8tVoO3F0Js/J
O6POsGGSXhgrZ+eoAYHP8VF+NAg5s1mhQxHSP9W7MIejVWdH/+SRRYx+TRw2lJhq
PyxC9S73GbJ8S6yMkg20nFdYUWr6RV/dUDvKUCeEPb7By+ue92zDZ2APfbCdlVCN
8vHLNSzzaueCLXQH2rfceN0qw1xwfuX5MKMMKwMEOWj08sJHVUK1PxnLxRaj83xW
5Un5dAbyEoW/nh1MjQf6LeTfWwyHXj/6JsyFBOmqgT9Ak6SwS0w0WDirMNs+R/O1
Z/SNKAziEHN3Wxxg3uXF0yuz1GxH7bZc1HafRKoIQpEbEs3oGCGQz2iwsvs02CbY
MfsoewUhj/87FbomS7OuSspPZw90ofPQQp4dQKp4vvnhlJf5HK0wyuCooD9xG4Nw
PYvl7+dV6tMERjOtHBqwvXM7VOBBceZtDnuz7C4lsi8jik95/Cf0vLnwrveQFi4u
VCN7F34zMFPYVGWYYiqqoM3572epKIRNWWTsA54zCP0jrtZvkkIWOutzebne/4Bl
RQ7KdBMviyo8QZlmXJsIIEdyRMM8JPjv3GZMe6bsLZVPEzb6TXqRPcAeMOc8k4Dh
RDLF4+C7ed4KkIWqh3r0kpcs5VleGIru1uTpgTCOIRq/ZQoBvo/5HqZyoE84c+Cf
1FflkGuanivW0YbbyjcEDsCFimq0SOAHlmDF88eTejWvOxFzCN6zhMlWpyM2d96L
BrTxvQEreiDole6bCKM8jbaJXvdb7wTFTW2eFeX8ZFcM3ubsRBVCC8RNAQ03+ACq
+E/1NP/ph/GStecOt2CyAbsSGVSecAyTLjK+dX+AR0GHRqI9KCyBbokN0w0mlXmM
61R/3pfZaDOUpfkUV31ZcwJYtfx2zt+UX5wBZzS68Ekogb0OULruWvJ06KwrIE0P
F87LOSSHGtStESKuVgpUDTcxVYS2C70afdcZ4uMAwxdxgKVed7ylJRVdOMj7Cjcx
hXVesLC50APflhLQkFQ3fb+ftWdHPbuP2bT76Zz6KnR4CTBzOgbdrh1SyhcdcBSw
+koa/fuJh85IcaLIJ5jBPfzz8rxfJ2ibXP70zGsIqteEm6I6JlffHWPToAa5U/sv
5fGYcX+XtuvN1SkSLU6NdIQnkpKIhOh3EZfRWsgwmJohv/RP9d4Q4BE4185vRGRc
x2RPpv/94hZ/4lwWyBaCVn13S3vW7Zu9VvToIPmzG/sCM5tbL/DLlg3gLPfU15b3
k70GdH9CIcIDPIA5q55adBO7eYSh9LhfZm66GPcxUE6E55LnKxI5N4QCWax3TAxT
MHM+i/EOTj3jY/NawRh+ulhKCz89ZBdLMRTr+cmltp/s+ocgllY3xL7bRpd8WRYY
AyBg9GsWGrVy6klLlR4ESgG/7W8tdvsxNKKIERBeUIqygfpJgpe+beAWWxyZFQcL
8eClEeN69/97GRFqxWFwxPy7UJOOCrTkO5nYLNc/WfwqYyGNR+OZ7JquYOZPsqoe
zQdtUg3HYlPRH5Mu2K21Wtsqm+0sjNIa3saUzPKXa1KHIznZ71TVLyubR5lzl5hj
a0J+2lTYroR6ziQ+f171fc3mJw+Cilr1fLl4CFDgK75dKqWl/iLmpzwJ6ZmpQI0q
zUlRgdGyiNZeJRIth1VNhxKdyCHb68aIrBqS1vRKbEw30pRIQZub2CeMbfPg3hEU
ubFtgDAdAGT5p2WyKhotS77G3otBHTkljconlo11uXZ0qjarE+XumRn4E+j9UKIS
7CpJBRCPPgJYY8mXJCL6OIUI0RTNkX2KdWtoiY+KBZnr1dqTdFWwqt0BKSoLhzgh
myU/CHK+nprWZWIhOzG3RTKuXLsq2+/blhwJFaTuqDnc9c5oOXhEP9hoAqSmzGTy
fvpGH5q8OjXujaAuRkbktRzuYOf9tN2Vw3yVcHRH9JOgnpPHhZ3W2SWVIuhX145k
9EaXrFp26fGeyPotbIeZsLBHB94/uN+dZOGCZT8+D6KFtM6X2U2nTONBLISuKPpY
xKsGpAXsRHOyrEZOmutNMdgrZM/TEMVxvIy1sUg5oioJ4CHlreBcC447NOepHDkN
Iz/glqtbLdYDul3QhW/MnLL+ysHFOaEERg6jjhulKBRj8k6ve6QIEWVNZhmuh0cM
gUJgIHJxvfYGVNywrwaqA0ARp0qgfy4gBWbRmMpftYq7+YiXBgcfsooUKfLRScQr
ggWIMZdGWz80nQ4Gya8aGfa6aGpf0Ky8g/qXG6FLHj3xgxBW1jQL4ZqbZqK0Zw07
9T0TjBhmoHXRRBOl4pJUaIuUSN2rsZuLUb3mt1xa4ybrEGkG4ONNxkWzavVZoL1V
8ZG9W7fm8h4rfU3WNe/u9YcPP58yeqU38DCWg+H6oKutIveTd+x7zjGJdEYMz01v
FNIF93eh/NL5cIAftHtR4zs1FJDc9w+6RDh+6oTC5xVFj7BC52QRIGNvHsoYiAMC
hUv23XQR/KvvpPvuAqdr4SwAT+6Gon1HX9TQN8C7jFT19Au5jEH5MIPh6+9O1GGO
JNaUEVmc4x+B+vMhbyMnLOFbqvZpemhV8rNfck0gBKlZAnlg0e2XElsi00EbCzeC
3Hcyx9GP62PtDn+2qEiLIM3SX85srcw57wRjU0gTLGUWs4JAso6Y0YployJKqqxP
X4Ca4wCZweetNTi9gVBno1mgO4OQul5pIvrcX0k9+ofsE2EZwzmScORSSpgE6sv6
yfeqJZCO7x46KqkpfN3pcLuGwNqXiwcNzVBHpjcDoCs8Gf52aMoMlTa1gCnQmIfX
pqyLIBPGaZyo+q8Axx3rgngL/HOBw8QBsa4MMvM/ZGX7hJZFieg94ZChKzFTExpZ
xdPH5qiWUlwqo7UAGP3lR9GN/d1IulzQgwbYutcUODtouhJxyzYsD+QunWKb0JfJ
nlDzOa/RjjuD5H7tu/4wEyZ/G/SpdHI1figFKcqEf5v4FIs8jG9PTxUckSmbLUHt
xBMhWZA6q4VvQrh2nDlkNuLJ2Rqww4QBmJ0iunuGIG9c67LWYYWblOLXd1NIJrOZ
Hmq0F6w5KLMmsAQtTm03bImR9aOkn0+YfetcBtLEhpHMy1ulaJhUQ6LCA7Kv2O4k
D2JT6mkx8YgLK2T65AFB1w2F5yNVp0SH/nWi3yJHOFyPE+dzrZh6jAIkUurzY5uW
xe2668OK6T1szDiZAiBf9CUDDy/ag+ywZJO4GIruiXnzeTBXSiDc52Llb4Z5kvZ3
UrgRfw1oAKBh2uTeT+ClHYWXrko8V5KvIkVQC9LdHwtJxqCbFfs+VZRSbWOipiRq
Cx2uLgEAWtQUtcyyUMoTQotU4jXRqYr8iCSf8PKMqGQz5p0m2Cw91x6q0funX03Z
60XOOa88CI9N4OBsbIVPmmxrCrNT/PTKcNyuY33TZtcJPQoU5k+oW22m1URcOF38
hw2xc1PB4VsGM1inqCWOPo872xLP8EznOugmmoiPbi1qKoFcwnDOZEALU3ZczEl/
IelbKSw1O4XOBLQ/Ge3IjY0ruMkmKwQYstIiQcmN927f8qfU4s8EZRiWGd/gfvR9
6oex/lJwdMnYjUMRy4vzBovqP2GbqM2Gb6I/X5z9hyqUOXU6cEil+25O3ZspSpHQ
zoNtzMfStMTHkuu6LK4Gxm+wOfdIMAln0v8rWpqSqpZquhrOckD2lFhsGSeCdXfx
rH3ZlDZ72VDeHQg4s5CijZGKgPjnHwpI9OiqE4pSGViISjSkdEgz7Y8RFAzb7E/3
LK97WyaoOxyL6qdiPfD3cyG0FY90SzCgwMwppZ6H9cpfwu/BqdZuy9Ttif30fAoW
MTOjjeaY2U/iK+mReXrbnE/FarRgRoDtVsqAC186tEesmmtvrSULR1mMrLnEaTNw
65FKqF16z5hw7mBx3xJVo276YLTQFDEUGHjrqBSAvdPJF4qjl3kqK1GDpZtDzgAt
wluuO/jgsLT0T3bXL/HqYwxYGeN9TSz+SHe0sBUIPyiVWD88I7pWsXDwRTjme1JX
LBl2HXZ5AlRdLRQqvF0v5g250tO5u/D5nN0hglggeVsSIkGaAsKAkke33lO7foST
ue+6OXid97Rjwh+YjFjSaGNfZtQelXZgZBAl43p5TS6t60YTwgBZNc4JV7DDjnld
CkO1sz2WsioCZ2uXxEF5AUmS4gM8A/9rJpcaZIZYvbHGzo5hlJAItMEzbbzb32p0
/0y0i11IW/kHehuVFE9Dr/7wwAXYYeIAurxf2VwHYmnQ6wJ7kZEoOv2Mt058ac7F
IXpkCrrihkbzOV3z0F3Jl7x7RzUSJ3EtGWj1pCqW9gkkIGEU0He9mtJEvEOd/fmU
XiAPixWtXVH8Cu6TbQWoCNgqkx69Ce7eGNROEEd9oLpFsSI+Kz8RZ9YE2VY+euab
lRjJOD4IIiSHCZNVOakeKsfkvHw/xQhQlO1ugYIjkkX3zycZhrTQj8yuvr0UfrWa
Ld4K+GdSL2TFt2Z3hmuFZ38wfGRJSWnIaC2/l6Hoj9miLqVvpQsiHz0EMokbVxbV
tydT59EuD/ca+6Ybg1KSq+wwvaFGd1kpYJBcDfYWRDHpzQRhHLacIfmW2e8P8q2p
YIOqIaovQD43RlNhIpVaUwRMXHiz01YI8i5irBcg/lrPgQf2SmacUAZZqUKho54B
o5d9KwaUiLvvfBcSOluBpwZHkqOp98vUKIsB0y3IaLaiU2DtvDiwykEybztTf2Sv
IcZ9xnHppf5aRALbsk6Fpt4a+T7uu6pIzjBSH2XGeuLF8HzzhlxULtoN9a9aGjyq
i9j8WEVn+s06kFkUoCMOUv3mdtjmqnHyuMEIs3OvzCy+Lm7Ux8zZfXpWWptl6p3B
0NyG+PkDvK50BpoTBX/zrsEwXEr7mzerNqtMHm9bmB7tkl9Qau7dpzRwYpxICtue
6i5Q952BuJV0prG2QhaozpRtqlK0nxg9Q83uGThQwzrVswNubr5T0vowrRXP3OZ+
Ulw2pnB1/ugPdnYT2I684N5DzQgjVJAlnki3n6QuVkojib9gXvHdWJmZ6msuh6u1
1wrKShp7kcJx1JcUZ4okGSWw83o3V8ZIsG7OQDwtFjIjDHAoQPS7/rkPdymcnsIb
i17DFjkz2IetQvcV7X4/O42O4EEGMcxAe9qMZIgvBGyVrQ3RPOTLvaKRfTLIWDF4
MkWkaUoAy4A7moOaKtJw+cL6lsIw7L6AnahwUXJsRPjIFFM0YqnS9C+WAq5bC603
8B27MylKcvq2seJlRdEkJb4GMKdAhAouWNz3bxaV5c2o3VZqxRR7W5UHL5SRNpWy
owXqk6127WtnxEjkAbsA07G+7eJaBYe8KdtGGdH33R5dyEkEAptvzWH2RM7uG9E/
JqMVrSAKASmUL1CU/4jbzwHFpev279Czc+Sya/FO69HiWyhttxaHkj1HccrRZRoU
pkK4Bca3bENh8V2g8M2LjLsA4iaHG1svbOPw7N4WDPWiFrwHlTkhje3vktIy0/kq
YRhmvgm5C7tkOpdi+TGAHQJ1mPfKB+Bg+VvAnj8obwrPKqXEL3xOSTu9JZAIg4Sn
gdDtubfAjq8IpqaltDhEoU4omgwpQpGoMz34ZcufV23nBdKIS2NcTm8S1PrgYdXz
CZZPi1Q74tSIZNt0WHCupnW9gGcjsa9lbyk2JmQuAhiPITRsQD+sQdK7C0O8dM9F
BaDsj6wIcO/RT4eZirVrJfkOZcqUJec9WtKlZ0OD1HJpUEIVm2ouSZHy11GGb0ej
2KTv022pOp8Se9+EaNPrlb5TupKJwHR/zLxIhbsPMe3dZLDfM3HzBb68/zq8iVpo
1Gd2AJVc9ocBvUkyQfLxMtRfkJEVx4XovbeU+5xPdWccaBfpKWxFbMRf+KZGtzWw
e5bY7PtRnVQ2mRcTUFLtr4dXb6/qojiGrLfX2YIAVhy0C+VETlydFCLCjTpRH1E9
AXSBvtIKPU+YSBzWcGhC35XHQ8J/5ul32aY8SBp5O3GB1fhq6kj/WBPHgGM6s9Fo
VFcEd2+W3qwTBBjTg+5CsF37M8yIDO1IZJmEgBnnNANt1Bu6jQLuDmGvlfgFn1ix
afY1kSyKMk5ac8HsYPlKtFj+p+oWEZRFbjz1X6tRH8NMJnJAW6kKwLNacfyAN0Yw
qvxCPJoVVP9tQ3O8H12Eqr5wxSI75RDRG5JRTsI41oac05dVSF6L4Q7Ibh2HRbwY
YCkc4V7htFiyil5rIKhTrJ9e8zriv3lOEZlI0hiGTKf5c0EbvazwcLJBpCswdsxQ
5416VuvgDbQlQm9W15QB3AOSkzHD3hu0+TzT9ZOAEktZfckIdT5D8rsOEGKlNkxP
BV3Pz40LPXWrQLf8aXlMJtNVSafnhufaam85ZTPaZxDedO7BGB04Cei5jIp3IE0H
lvh96zVxS64oDfYvikvN3H344zwx6nBTETua+9yWEtkqv4IwXzU+y1nkN8gN9fqS
R+SKQGtoiROgMHN4JxtazAzN0T7vYbzVypU0jkLFD516ziW6emJ2H5KdLqLcMCi8
GvSHbBam4XTwBdADHMdKoQYrE6uy7QCBVW6HrkJDtywqkUZVUOWJYvObjjI/ieDI
Jo95hZIC/sdKWDIraq5HSlDo9maOTkGFsFfCIC3UiJoOxVaokvOKNgY54ESs6xdc
cBPEcPu3Tz4++0P/bJZsDrbDpO4JqzaqvmhMN1lJoAEGoHiLbUC2S9WYhQWzB5PQ
nT061xpn2eDEMzYdMmUU9l5Br9cBT6K+RrZOMakZHx6DXTrwgbJVCNiqAY2BmzZ1
MvcMREK6lh+ky08y5dlq09bSrpyNODFHi8lCps4NmHIRUhvE3PQAq8IISXZUEb09
C6820pv+3Siz/Da5TR/oCQ/0UEA6hyHKvdu1jc8eIlNrqZ4v5Ha0baFq0Z9lAkSo
ol+2x6s42oL9VVV6oCu1OMKR8KSQoGFyo7nHZslrWu568SA4Rwc3+7MzmuttoiGf
+Vg86UYrizb8o/DVVEs11rn+0LGeFcaDLehPdOdqzQcT5KXDRP0lzJY0WYXgwLe8
iqe3oQcXWjacrXDvFsnnsSqu/3QM2bIOrh9twYR7/wNyiDwA2HfZXvMjk6ownB/d
AlkQ8QkNJzD5nyThITCJqr5fn7ESCQMU1jnjOQKppFhTA3N7oZBDK66FZIdgy0Ko
9GOMoJFx92JLVuL6NkX48sSmYjkLuZw/Qd3/IhnU+2qTnw/D3J7eY9A9XtBU5EY5
sLatY/D7rRzi1rPoRTHwGelWHsf7BSCB4SYiHi27My0J9r3dzITS7p3oJnT/lcxB
ca93V7JuuIJi2CyPDSw289SkDrlfO09XHMuW11Qp7dhvSgJcJ51VAp6V1JlxVTaJ
39jdSPgHOh11M/0RGN6EY0zMrz0VDU1FU37SiDDqgDrxD1l6W/uQE2XjhwgyWywf
QPkIdebXKiqYLzRGv0hDfrHe1sMjIsrWt53lFlWZJBLyW22alDEw8a8sgTdxF1PS
v2FbzeC+uFORGcPUDajAqPeAd8RUpvIIksNf7Kri5YctrfkFgJmZXM4c2VO0rJGl
ONl967m2hJ+0+U/1vkkF362x+DmoC9B14pQ30Z9wUJTsTMZsuMgkBPfMSnjnig+v
4vr8yW1dy9/XRaUZx1nkN2RDI2C/kNiFL54SBuG0mlJeItHG44sI6Ang4KEzEQkV
iDot38edxlTGoHdiwfZIU281ZRpTIiERDrg+8ebZA3uejMJnMpRQi+Jef+R2lpKC
S2eOAjhWclwbf8Qnnb16SDZfwisQ3Lwy8IRRr1TaYcw9nYjxog8HHIHZB2sFedtJ
fY6NONz6ERByI5ey8a1Ju8r1khXOOhRqk/p87n1khYCukqYXVPcsJePLAsIyihkN
xRwArOrBCVlkGHORg3oOmH0/rr4dLD1XHw/XynOeWObWYwfjuKRSgZLwq/MSECOW
VtA6L1EtVjaNp7OeRT8QjWLUslt/yhJIDbftySaKkMqDbMRIYfa5eXYPJrFRtYQT
+dcwCrkK2FSdXs3bJZPPRbsmXslOl43Y7yrVfNpxilgWFYiqYMVuWo9DxPHYNs8A
aldqi/KSX3Vh6uWDcEZJS3w0luGeqJCDdmvgpPKGFeycoHN6y2/sHoFubXuG71SM
oq5V8E2kjEC3HieVKs7nN6JVV4hIwfnfqgLIT90Ab8lndZ2GJpRs8W2hUTKx2TSM
9ynjUh1ycZADd+Yil/roPKmpxKeysTCvY+nKrp6YD4B7kKtqviGtadZA+A9Q3So3
3F67XIcevSOb5k45JDDZEpqGpiAvoyEUGdYjb+cOivMW5zoZpNqsYAym/E4XaHam
TaGMj52ueM+DykVYIcFsoZV7ErJKlprPJyCzHRu6t8/gWx9u9+wvPzhfn9wtk75Q
itlXSjCdqkbYtv2vtPbIYWzUARtvoy6CiqcCAruVfjnAvI2+i0q4c0xAWfFQUfaN
JHnmSccfrR9eUGbhcZo6dHY15qikjM9nje64Tx6cr4RObcAFqPY2eXhp/UEbEQMz
wDJsWKKM+OfcPv2mvweR43+EovfATv61LLbmgehR/EGUC22IrZDJwG4aQ4kdjfuz
UR1+Zzg3SSU7+B0IfTLl4MBVes/IrQHcHcUHjB8fIyaS1lmWhBlwMA7XZbKfx/dB
tlt6T9qzKRTkq5+0q0XjtKUW6t/cP+z9y/Tf7FQC6sNz9lVIPwGMjssb7XvnHDO5
pPdvXhAv3P62EUkAaaG80Ss5/pCl9Jx+yjeKHIbAVRDVDAwi/Xcad6RdPW8yZEQP
akMjKEvPovFCruOk775vOeV1T1x2OBNwGbJnfAJ1+UrVAYtvrBu3t5HylMfRf9o+
loFaREfFAY3Pd4bPFm1Mr/i49hHKGdae97UjzQmDmPTsMxReSeZ9sZzKgKirwUTY
t4DVk5/CMq9LM0qXD7KqWNa3FkliQJl6fR8mfqLumD9EtgJVWAtpzCMc1iSc72vW
+1S3xjWUK+TyUXYv00kzcPbLkyDkAOhAGTKc8juCi3JvLAnkXoIqirVMJ4w1DQbS
N4WN8UsZVFWRwimEUCWmG24YR7+5USXNZcuPxAMHejSFW41KlPdd/wd8JUulqTKd
7xJCT8UENfWVZ5U2T4lOjJVa5LeqXtAaXYDs539iEPB+hmmKM9EEbnBzj0bB4WGA
w2D/ND8Jrbq8L/E7R8In8idi3yEhe6tLY1cO4CujiuZ2HjAnBuZ36kpR0prYh9MF
6vZE5Ux6mCpnWNSwzxIK6q+YgnO9n+2sNYmmThy1UJ99GXB8kg5RX8QrjU396GEz
CgytgTW33BqEcuCRP/rqZ4CrgkVpa86YQiohmlrWF3NHLo/lgKqoIfI1652pmSbx
dSjnEVRXdzEBvS4bIee0tWZXK8E+7F/GEaCC84NYOGDXMXT2vJh9nydbLCdGUF3K
ifIfoHIJCDFVJnGlMmn652XMzuha6iSHO6rlR0BfrFWp22ix+Xy9m8F4Bkwxvl0w
LKTBAbKPujK9A9BDc0B2Y/m+Xm1sRxn6xaW1IH8A1CT4ULu7kjqspZ7ANj8PW6mm
tFp70f3n3JppU5jYzHI16RrZwUTfaKwf1HZJXpchz5wRbaHRGvSM0qIdEWjSv0m1
aRWnJANzU6aM0rscCx5aLrzKA8Xdyak8zTuNOlDuuFDlkodEv93tBRaDD6sxjAqK
4J1X51cgfftSyNDFzdUoIyyYGnsLA7ZsLn+ACWjBcuJ3EwJyggvAIEb1Ta+OFEoD
xOMjjeqv7dmDQ12QWGBfim0W1AJ3vIXd8+olWpR/5VZ03G/tBIecHxzjB/oD+HM6
KA35d1sXlkRNP013ry+xh+8tkxs3HfgRQELSf+0qh5te+uliRrUFuYQEF0hboliC
4SO4a/sudPt3mWVhJY4OaKVbX3xx79P4q0kQWKe1kveY/BQkzToSlJBsnT4aKqcc
uJfnNqY/IIWwhkzYywCAXQL811EhP4n8DKH0WurIedmlZdrMGmcupQnxPAa0N9wN
Et6KWesSy/EJ3HDFKfpG5gf/K15M5ZyeWf3WmXOlxZdntSE4ZHHbt+A1oPTjL9hl
0buIeOEh0t7mmdtaHT+/0EBMOG05pLKKr5I7GvCCe/8b49zD5q0zl09J3i0GJIOA
tibwq7QbMPMe7nZRbfTsu1d9SIWCMec+isDxNb15mP158qhf/HGIal3n81pX8jEB
XM/xL2qMlH/K0QFL6iC7dv+daSrgZZHxFwe0vZmB3RqyVGqCz/PGoZS4+CWk//IK
/09c1uNcgcWhTlxA8cW6OEnTU3J4vb9r3I0AIM/DWtuJAhHrvA+3KFU3fg0hC0mO
TaOggKTlWPK077TDl+O9mWx1yb6g0ydLR7UEnTvSqQmjnxZM7+D8TVArCWoxcg88
LJFWWaYzibA7FlcyX/WHR2c0wt1+Y/WzyZM1EveTJgRGDedpgTdU7gvW5KxS3gee
AlxPhxkj6RdfFw9Wd9WX7knZqphFhSbrW4SzbGIzDy9jm84Vor3omeDjG3Zk9CAh
ktmBscCTkCs2sVXdX3gaRuH8AHWZepcwlz2/l+NB75BH9Y66t0jRoyl0ubEA1LS9
+gD6YvLGG49Ksv4AmpxOQzv1NxQ6EJJ1u9JgbX5OBZKNidMb0bsZih2I3eQ3d8cU
Ljtyye8wJxrxPw530sZGq2HSrJkS2uJOWCMy1tKqL8xerqAR5arHbkRZgZnXPBXt
tnJuiEc07noohzxgKkiuLNrwQCWmmlQUwGKfNGEhJiiIIKFV6I24mfhMJxzy7VLS
8eZneYBb0HObC6rjMIBAQdYUi8mmS68H8ycmqUYtLxfu+3pWTzjlSPayvi2J3vfl
dd97NUd9R6TL6ZObdk56zpzy9sPL6RP+I6t8Tu1ahUZ++C1dr85fE86wlQSdLxo2
mUAq+VsBgPYzuWOHn2gVvyxHTItZMulOEqx5O25JuffmDGB00CEatg7MYqHz8Zaj
j444qUZCBFiNd35AuFkjkGpLKMsf5nqbV3ughXtzDxh8wv+6W2DhKi/iWvFYz5c/
3rDWfpicF+CXxORuJyHLhoyAD4fXXsYA8zER0XUV8zLq0ezCOf+jGLjPye6ZtcbV
k5rRC82DHUUKBPxQOuCoBW9OESzLBQqpMGiWeZ2HYiX/dyKnf9QO8yt7F+mh+/K+
Ubp2+r+2GjUWiFI+i8isV3eAny8lYT4yaCb29y7WMRlXjJGMEtvIngbPxTR3n4fS
T4kRYZvai2UR1VvBL05zQr3psjR6iniTkxDn3opFiAb6YbXka1Jl0Z2aErdTOwWI
z0OpI5yRcGNeC6WWVGj2XfhTdzc0wyT6bjnmKxtRqBkUtqfdpSE2ja9QWJl8e7+e
H+M/kgzEqpMIWzaZk90x5yLDXIJn22SFmc/FhEiVSFcIQb+fhG9dcsGoCUhluGw9
nEUogfjUyzn4feioS9D2rr6GCMDWw4DpaJv9XVMrCDdgb4SfRGNbEit4vXCsdDPR
THO/m5dR4oJ/MKhe9ALvBU0cycCzdsG+CN3OG8pitLdi+J1DsHe6trCuaV8uqNPK
wk1sYJee271lknKeqV6+vcAAJCWEilEIL6+Z+E7HBWsYzB7B1lwkwWdgLFJ91d/l
5vzbXQDJXCYL3EWsNqdcPWguPU7t4fFkinqgFKb7gg3RTgXBSmn7cSyfNW8e988+
FipPskirdSejGjxvbx7c2Y9mme4hTgMagDcmfwEEiL22M/zUHAPpOu3CPVgCOzMO
jiaE0kmiSwJUtn7h8iv3FtIpSkQzgI2gkhV7kvpO2HOWas1vsarJMI6q7aLWYwcv
ZeLnCmRrC+aQWTM+N9JnPkdoNkTewUBAwM4Aw9M/sl0/wmFpblWf1BhInzQTMa0T
dzDUxbjVgEERieQXSFi0Q5E6tmMAdXumCBetlvN3D1zZTYL8VrpEA4/g1SYu9Vko
60qp+sg/9kkqTYYQbfhb0DsX3nQELCxZT78rRAhwdFTSt8MmIrVX2H9HsldF8Zsj
nvkpcqNwXeTa5H2oB3WbHkwCuOJMXfsydQziM1j6rwfsXT1Kre1qu6ZdvMjLZw4K
PlpE2zJEwmiDvXDrWsXYP2JqLsK+brXcGEMAh31EixiCr6k+f7Z9VGXIYNY4lQr/
CB927Uox5edimg8TnXyq6SzpgF2Lwu8P8w6mMuB74RazK6TcsYGu4mOS7rg2i/fE
6QGfl4RdOIkZTyrJY19F2H4w8k66Qr6DbcXfh4LIYhw6PmJ+ArvXnptpqG4PdB4M
afuywPtqL8mxFZDE/qUqrbFEIXysI1ZAofsdXKKP8ItkpMnNcb3pgO2yLDxMT984
JxZUdPW0Azsf6bsGdkTYpHTOL2GkvN8DvKAsPJaqJfMmf6JbHzyPjO597mSgW9Vf
oDCQd3jGDQvxdMDFClNR5OWX1Ae9pM7Obo+XENBpirFU4+bjFtMweHK5Y1KQoSTF
d/9Tr151RATC4WRepfL8H3zRbrHoLmEoVE4U912pPEcWbe2YGVBztHx2QwuImadp
lT4MgxSvxurfMkLYaanvjlcbj7YYEtOebuUOrTF654w1TrZc5dccH4omWYZzrArN
iEwnQDcs38v5ErWEeOWcvcL6HEOv3ZMWnHIupNDtVjkfm38wz2NwmtlNSe/px6qA
T+f0UchoDZiIJ2E14FhPXKnu4OkCFjp6pMlLAjZQBBB9DXfmgrE9Nkn2qhyi9PDZ
16YUD1Fk2ZzuRXoYVx+QvWLXC/g5D4Ymuqq+RrogNEFrIYZ9NypgmsHfLiRiMlMk
ZsxBV33pAb75h7TLNWVTMapj4uD5V4U5lpMDXFydnHDcTostmbdhHCMEW+T46O8h
UpSs+WrgidOjzzyv2LGNgzptgJOX+u9srG6QACY2MqsQoA5OfuV0i/3Nq88/QPp4
hGwPIVtjaJn87/zcfInF0PNLHKMn5Wp5noPHtxOnTS/mZ1Qdjoh9/NhH8jJgw8rp
67oGr1yLWwk/xAB3eRw7dHdLjvnfBfelS/3kDvAk8P0R7lPnQ8kgoho+7nosukTc
Byy4PZcXOZ3LqHnkoU+VkSsqZzL1kOJRLn9w2Ku26ABuaPuLuLW4kLNveb5IHsW2
psDHp9dsDECed7y90u2DY7BYD8z4uXhXer38kHOTfE5o7a+v5EI235AedJ5acAL9
VCScYGJ+Rvs+WxuLKOaiZODVa+JJ+BqEAzF1Yg9x/xKOIH1Xd0UZ5Gz+bzmSS3lG
ZnjYIe1lMPh5CxJ2yO4sEbcF7g4WmJ0xFnPhfKrkiCQymDYGhus0ExymmxPS8ibg
YxuSgsBIlpwch1c5o2U1E2p6BbgWahzRpXKyfpKovVF9lF6UMIXF5JTi28Wp+XT/
zqE4GzPj5sMMbALyU0RloZPxEDGxPmOWgQqCmqjV7UqaxQKNkb13GrspAnI54Al4
vhUTwiwK2hUqE8Mby0fB1t5Gvz07luCCQDrBswl/LJQ5gML/swIA3kA849fGj5iL
N9TPivwbPsbMqxlf4d+TmEJ77mShtNjp3caZHizjBdndIzYhqRnpS9+XFeGyKLLo
b0EnZGbeNy4/rUkS7Ppa0/c6VUbFW5BK9OWxuSUMixONz8fPbLYA2O6e0sjtCzMh
Y+rJ8qy3/HMnobIjPAm1G2kZdp4Umzl34GcEJKiLep9mUb2Mc6aITqSQc5ar25ZX
UTTNHgoU/3QRD4DCVmS7vNtIc+VEBB0GcYLJQZ6gSHdFze/aTh+zLV4DvlmSlGwC
hTXebqABPAAspePhSrZwafuYbB1gzkOcThqlE5kx/IwtbBaZWc7O0G3pTer/uFTC
V7QT5u5sP5rMWUkvPowwT95rR1r/wIZqL0ZYLsCe0mhiNoar45S0wW8rHP0IJTZA
isp1UVyqZEU/htTbuVXaOgeI1ypOZbjJ8vDYXTxMyxTGvsQrxMhtBibfLC3n6HiB
tLWExVAxJowc6kmKZjHKd6RBRBUSmSxtTDcb0o0Gy4dyZZ3n4Tx7LqxzqkmOeAmO
/K2CjaReK674WBYixeySLOQil4qV/GoQUc3ZoW8MGI3Adwpvbpy4xqjy+QFGziLL
cX1SbIJ824A5CdhAj2ME55teSnKsfG5sYvuCvslHkbouH3Ui5cbZEGTuRH6QoWMW
TBM+JIigwOTnXGkX3ncq1s7m2/P6LnGDWSdsgulXR3TiohEoP5oca7xNZIdeA/FK
LGQl9DzkqavwTBia69f9GaVIq12XNQrfYTAz51jLR5tBsItVyx7Vg624T2daGsYa
GSW7r/XIOUWQX95V5ft1eJyRK6FDZAC6U7pVMm2mlveZwAs9hVL9iI2CD0cikVGu
SxtmHicNdXkw+cXnJhzvdZ3JsJGk+QPRG7CDg1n67Cr71s/lbRhTgR4nBzYFmJHJ
ioiuFfcHkzWRt3xPDvAogXVcopGQ/lmRnyY/EbP1bJN9xYMDHYPS0Zo0mme06b7e
WB/ZIIkxTx8PkWut9GEF11yKcgiAouMZLElpdoCeFXF4Aj7YocNTO6/gy7mc1pXQ
cs3AACW4p+LrZjj/dVlqVwY5zwfjk02TVmLWnyP0Zhk7VEsIiCHxrIaSqCH9SoFH
aznrKQTDUEKgj0k06nKHopqOchKgYbQn7GLqemE8912TkyWPwjbvoPw+/q4IP2Eg
GvWRRwbcEOKk4jNUX2TphNCwYjST8EWdoFspUp6LwJwH9UDftQn2ZKzo6KhJY1z2
JxloM0Ojr2wcyJMpYvHmjyz3cDTuEph67dMvnGUStCCNH5vs0tfasVSCodKct5En
eqLP2BisLosuelnk0c0QgFBenBEb67Iv2K7pJnFrQFr4zWoyyrFrkmhxeUOBWfOD
4YCKj02xRDy47EReICtNrTg1y+hYqFSGEs14V7zAUzYfn0fxFQZzS3MJbWFYBXbd
91CDofQv7gOlaWjY/Q8xuzksDe86fCecBz8HveLFXVvbbRdiCR3gGmy8++x3pTPX
AbYeVT/IOhrwbL7Sw7q733DNZt4lpBjxWwzqHjCD2cYsiYQpJU90SKgygePhP/r6
lE+SZH+648zMAJDIVqY2gh0qRr/UHxjHSZb9q1iq1XIxjYkYw8azxdCFojeqomoN
K9m3Qku5BOYvPA8b1sEiHO3+GNZ7lKGx5C+nPDLCbAdOUYEx4JFJoWKkXbR9z3WF
7mvwalbvtCeX+VSFV+s5Qv3doC+qS/wf1Axn5+hfK3fIyl007ecZDhcUhYj9Kk5U
f8pqZDYyOuj3iqX8MQwhwQUV2nQ1hrPwbZiFbiaPTuqhuWBnHU2eV8hKJqc9Az7k
a5USy0pHbxlJyfx07QGKkvyUXLLZdB1fVwT3bCufYGo0/Gsb8AmjkqLqeIcCebya
ZC0l07bIHdfLEx/vqM/upHdetddyYj6t5HQ/xLKDeXfj4LXozf9TFTTBmynBGr9b
4q5w7LizHr00+5NWLs4qTMc3lwsC6p9qDXYf7VWsb0X0g1x5QXeDDf6HPDyGVBeQ
oQ4ZrKgrwSHZE/ErKaYNpOSexskCrQ+de3gq8PNt+VEoP8zZ106w4ZZ7YsbjLJhY
EXOs5eJlxK0k8RUiZnG2Hp9xwIzZxF3+h9rR+9HWbXKhEJVzXy1L8Hszo1g+wi+d
9QYI9nzFiPh33GLeLdZ/ym9d1jSraLakYy3BlM18X4SEwUXFrea8SRvVt7eVg6JE
2vl9kUco4qGwpQ+C6wE6KWbq8PzyXPV7RjXrk/S4cyhfElMB7U+aYdHf7bmhRuze
7wi3O90gJaHPHYYI/G9Jc3BNb/NRqpqIQ30isNVFqo11ZHTGPDfHrvBx8mCNmDig
1/a2U/b0GdEKQvtkWdijmGN1X1CrF0Gpm0ZTb0XBayIBhBH4Wg/63lJD9Vs+2zM/
1zfL2f8YpkZ5+IKXlsWh2gACYV0d5O71NYfisVvZ52qNLxf8rssTxbFXoVQlrwHa
qB+wxajHA55pjSXCYSLPplf1TEELfE68henz1j24pPk8CvoMR+eV0ZbeeYI/R5kB
JSMhF22wkfz0HN2zgYvgszcclJnuZnLQDgUjadnkqjSV/E4Y5PdA8NjqdfvoUzNj
ZfIPqpCpGm9COvmC35c1D8ZmhyIJAx4MjbFzLZYa4amUhMwmnGvNAa0NAH5ocR84
jGiS0fqEcRBteMY1bN9oSgxdPbGMdVC+l6qvtBnQyMhf8MoWOT6OzMoIvpc+oqEa
8UHl3/aMwhLP1ZJ/ONi9NUMuIbqw7obcnwGfFTXyvrE15GfIwI8oHEM7JXv+uPqr
vXHa45s2jqIfe3JJndxeq/JLvUiPn9t1jRJeRGE5mUo/CBKAHA2KDXRQbEuzcRXy
eJrebahwacMgX0IcSPwL07uvR5vgj067P0EQhypglpiE8qEK3aN+D+I7yBbIlrOy
w21aOtqTehvyyfGFSyYf2kFJQXMH1srrFlA8lGED2JxafjJWadYME344sqzcRlFZ
4ii730eZJhnE8OYEC9IMU4dxpqlTEYGX+m7GJ7BTpSxv7nMELBtFGcAiRJo/bzrM
CRWZ5pAQcbeSveaM/oaMWA0/413+V7sEFARpdQcAgmqIfjvRU5XPtd3Kkl0lDdd7
64A01QAjX9FbqWRKukp+aksH0oCK7Sn7GFzj+2+3+Za9WlEmksJ2d4EgbqOXAKfP
j0J+Lk5EVR+9wtYYy36X38D2Z+tcRzf7jjLhTdsS/XCrIwOFMjpdbZ5Kud/h7Xou
OdiEgdr5eMaSQ7VmENVjznecp8wA3j+vfmDYKGYMX/QrSQJHnKyR59m732mhP9qv
flecBA5WXwkTLOuMImdw0OaIJDlGLpGo3fr4QMn7pYXwO1U2Dl10bDLZUgz9wOCF
h6xggGp+zoCkc5Twzq1/wDvp/d4V748ZVS9L76RTJaXOizUrUBrnrY8gscUjDKzH
ipbD5TICAkewX7141miABaJ1jREP/jS52xsJFl/i/Epdgt8rHwgw4o7c2v6A7nD1
gOk0aQR8EV2eDf+XQQfVVIlIq2O54v7NpNTmeZYmPnojY7zrTPD76zD9tBTKftb8
xybTeYVQ1rTGHbyGeIRDS8o1Q/XZTkIFUibcKcSKtyGB77nL90hGGT8Lp3ZXOh28
/hseqsRjYjfoA0+2teNQBJ+jbbyEfwIljwicwpCMrr4gn5MQfE6gbp7JRQadBiKy
4rLH/MP1E04+DdicosEqt3rVBjRDV2s78XNppDOwjHgUvDXlrs6XNPEHuQHDQj6T
V+jX7o7CYx6wDxiIOx4HAamuQO/W0hXIjwkcWm/rZPZBzf6yz4aopXvhAPLAhd8E
0wLG0jqXJgnUHlC8LqXNOTSiOx4QSvOCfuuxYiESdYOfLsBjQhEnRMH7O+8acRWv
vgazSDJGMr6y8nM2f8lpfh3D9x67oZyNaB6B529bp9qPs/i8c/Jq+9o3CcAPkrrk
Oyb7SDiXT+kNRRRl9XsTX1u5bHSn7Qac6OsO3533RP9+9N2NOy6YJVEEw42ucv64
WcH0TPZesBwXTyTLKnYZjx5FuWLLEEQc1N9+SUO1PKhcv+oVicgoiw2uqdn2FbWb
f+AcVkzsaUIiBNKvcU4RhYsRwB5k5mYlaZVF+pEMsneWQd4HQVwuU/BHbT7OBq0x
r5AaCbjLzU4v93O2JPXcgPZ76tzxAge8rZ1pg7GnZwriQxsEeKvNa9xj5MCrCvE8
8IY8Tf66I9y8BSbXL9CniubQYsUwXnf5rUMA3h/+OIfNDZsL8n1JKYonDHkGUruJ
eFmatKWnO0tR4LQ6gCGVeRIYJt4bxd35pSxoymwzHvBTpE5E0kFKH8AReKlAnb6G
6HAWpxfVQv6FccbaOTKOUrucOE+4y4LjKUKY80XUAUhGNiuiEGdVIA5lN1nAuww5
KIvGu0TAxabZhzQEEq6cRwgQt44kdxoLVWOlvXLehkNGbwmcJJHz6Ihkl/82NuDg
JvmkNCHZN+LfgGnH+MchlXDKnf4nlH/uElxEyc3FK/XPpnHlwdZI8oCfdeEtLJ8f
lfbZ9FbWoC4eg1OE5gBFw3VVBE/2cWiJLWRJobhe7NpjsxbRS8M2UqSbSvETBIZ8
cHfQ91+4JyZTAyaYnAQOaGpYz5xHhCXDbzvATym6K0hsfuWQNWCOZNSn8eZhXanz
N9nY8xFz6icWQm6I/XhB7Pgx+e3dytc2LspK/BgDiGDbsiAZHUPm0q5i95JYZbIh
uJDDJ6JDskt3FRN47rBa7Dw1MfGk+mYDl534yO+XzMVJegwic4IJGLk3q3Oh3EO+
x0M/7l8PsZjzYsoFei4i1EY0AStaAipErXSPO3ja9kUPEfwA/aWQDcqIGEbJod2w
o4UGV2MVfTIsAZuUDJMJnt/hQVy8MHluVErukoTFBDvTkJf8Yrv1dMatv+4IbQDc
o8aVCx0PeE5Z+hh/eSMppIxqCIwhVPkp598x3/cEpUe0pJEz+wxFoYxkh/b597dE
hAExUWPdCP7dCpRybOkj4Rg9jSFNK8HK9QDefokis7FMakEyFCnU4j4on9LqE9o0
lOPT3jGhNbDVQ1Y1h/SJS09Nmo7QWJb9Xh0+FRQqKv/OHlaOZjyy8jopkWjFLtRO
H1EJ/QGjFyMiDeX8YsKjQsFfSXhrgc0TGzeLloH09nVMl7fHdR8D6HJqTWgC8ha1
+bkZ77B26J/hLO/8/FpnnNc5bPA/ToVEKyzaKQhlhiCg8EXP4k+lvAvWLrnnSLxe
+/0588rWdr1kOXnMpH7h3gZ5KfISEgXm2cgxr/LpJNtlcOUPbDNtZk+Ci1U9NFMV
T33yqspIjO5h1nkCbauNCgqyfkmfC4xlfY2YkCTQnib3EREB6fz74rBVacToAZrG
mzIQbx6+qEHCECA3Jj2rrkHj7aYJJM1tLTArIi+M4TC+1kJLqpfvn6ymX79gYNYf
Hio/oF5uYqHjTJlbwMMjqjaPF3/ELO5z+UcvsFwaF1hovlAEyWP0XRH3R4uAYKZ9
o6tiWpY3Cj1u3SuxJea6WPcclVHQILF4w4XeEZXS8QltLjOzGyIT52NyJLD7EU9g
ZnGUv3bd2LyKcF8Q5P19GrxG9UZ1Shfx9+GvIEfkEzYtfUo31FhCP8BanIK+EACC
CAbF7eOvCKDX3KQ+xoASgpSFiWF78p1dJK0KW/Micy2/NuanvWYu4/GhxlUJQaNn
SIIBcsB92MF58O+Bs/q5VQPn5zB/8D/yWr0s7RbPCd6OvilfzLRgFecyRGl+Ti7N
5qbqkKuwqDitlXT1GlLQ82p2GHiQtWTk7xn9drpk11kiix0DTEdbXG7Gt39wbwpO
er9/YagXy4x+zAPgMWV67m2Aq69k3UBatel3qh1+3/EM4ak798qFgO7DP/CGUHo5
D2tAJePXarCyj0zATnB/dD8yEIPBn3mnxYZpi28tNKg/wbGqPLPYNN+8/dqM5MkD
4dNEIKnvZs13MZcaHlAwF6F0Po15GWVIBT3swlzJYoQrFxbZQVvYExGXyQjxQQkT
Q2L/M/CYI6DftKunoDf4tUuVf0bFykYA7oxGOMRzShs6TL3q5sl3Ew30TedjZTPy
/Y5UjSzpMi2PYx0FajP5wjKOcjI/cozuCU4p7BYbAHh5LEXrYhmJzurKzbf7ys+A
5cIEJHmDhczXV77J9yvJ/1Dv2Vw6NASPYISeLNxmYJ4DIxrMERO0pg1Dmw8CaGUZ
L3vgsSR9n5J2U+nuPk61rXv6BC3oSob+ev+kkvkrdnHWp0saQhNj0hB5R8MBvded
P2NmgJiOvJSNY2WHNctD+YUsLYwfjCHJPt+pLXvapKP3FgFAhJY4zDZ7IG2rK5CS
cLvlUb6N3EoJya5Q9LJUyWqF84vVwLjuWMIz/lszVKCF2rGFAmDfmsKr1yAcAU8l
QhDSHDr6XDYt5wryFz653zK6dH5cl83IUPc9alMkc49Pneqk6k0ZB2ongn6oKt0S
9n41vMyP9rwsQN5DUksoEvz9UZfzB8Nj/kJwuTBfZuSP/btWVP7aWZlV9DZi4gsP
grzs6GBwGKruNVbWA7mld1laeXeZh+I+tH9+5HV8uFLhj9eZ2Lwi7+q+ZqHx0iTb
ZTzuUoVVfjreG0mIbBsP09b3ChhpAC2WcAktddy8y3EROOk8BEziEXYbX+xFKARo
I8tjceTTOBUm2SQ8ymRnMdSSnhgZArku9xHFOBbZoi3mX2Fx+wfwVXD6k5T8OQ2F
mIWOAA+ub2LVN2TVpcWbmG2TvyKYYn1R+BEVqO/h7HxlzETjEBSeavLVhQhAfnFq
C49pKnoye5Udm20o7Pwv1+H3m2qXwo3RtEgxqEwLfdouB8/YRqHy4Xyyd3IxCP+O
N5ij6t2azX6BDH9T6neK5VeIg/lNVhKURZWek04l2g44eGtUaGW/XW/q9xCXcyMo
5wCHVIIjS6ZBWitXag13WYxFJ8amF6nr2xwW61EFrJL4rLkVrALJFeB0Yi61SDkx
tMVYt+GMmJA1sYZwEySUHZQL4onnDqFumaXeUQXVY/SJIzNX5zQS1oGi8Gx3yTab
N6yA+0NfCdry5jAlv3LdtEi5xVONrkTlFSQPoN+2MyrfjRcOzJh2M2DSL0pKuiJr
NetfgTUomo5vGx7yZHMiZ6m9kDe3bYQbGUNq3Zk/zMcmudTIKM/5Z/3hAXqSzWIg
xyHr+g/z9be4UvUlRTidxqXFk37XKpJ4JDh3vgIMUZUSVVvxoJWfKYcPddMZBd0Z
N1+Bq0kbcxoaP9d3tWh/LTiF/V2rhqmvfJ0TEnXAHBmZC0oM0DnowM6ViNJQarEO
+jwj7A+71OT2L7kFdA1y9gn4cg4qe6qcyyFw0z1BZ1CdCTN8jWQFwu1v/c63wxQY
ZU/NlFspL3ElmJbXs0sIHaAfw/Bmuj38vUzXPYP3BOqQbzEeiiJM0jGJ/sgKavK1
Vs5Pd9d5uSQssUpIphJBFtoogjMih1dNZspxeOc/rv4HT2Bp0/V501c3oYWREoz9
8d94y95A62RxRVHkcr27wpd/hJviy76nKUb+Sl58YXFIMWgURuYzLVPu2xZXFW/3
7Bn5XkYQ6yMLSxA8JMAys0TYyzpesFK8EFyjGP5jsJhNe2tgqlq/NvrFg+kdcpU5
8AeQxCEmeU2F11dCTgssNRBldxyZduujIwePV0HVn/wkkSPTZK8ahJ4XJVdQTTco
wAPku3Xxkrp+TFXdh4F+OeJTfM64nxoDspim6vvSaAOEL8+n71fSH3H7/hB61O2r
+DCKckymzK83qPSHV4M0I+k91u9JHtPH3n9tOzG7LrQ8YoSqKKCznNStNLaOOWim
Y6nSPlnx84tw63D5qmcs2Vcq+EoSQJsuqc55+cm4LoaCp3Ngc2s3sFTTLG+UNkqJ
/htzi8cVJsU6rnJpVV6XNT/GimCBeob0V9gXgAXAaC0fn1U40gcoNrVK77O5jrCU
Pvdu6EOe3vXYoSYXNDdPyLoehKo6AUt1khzVBrtrz0O7UQNtkngPkU0GXfcen6jL
rBBZWdojomgAY7Yt5so/fbkond69vyFTAyInpmiGcvB1LbyHOwanJb8grq2HxXfC
VAWPKzrxjS1BKexV6JeZEzT9aMhJ7A2gVD9tSvrMlMJKUbtMHmppHtS8fO4MIE+K
WBiBBvptrcx+0CdjDfm/+1KNucpSsjjj7NjJmNCw5z74Jl7m9RkFhluyMpm02xV/
eNKHz2ABHH09IEa4h9TexcIW0+oQVVyG+7e6dppwDydhCSVasbiqggX1CC5rb2v/
YtC9eEuiF4A0lG2ZAZbzbuBkASOR7a2eFW4KV9iZijsjZEq/6uYJ5kVzFXWZcYpK
lLY5RWISS6C9fgkc1WB/7agpDyEDbIbYEDsaRQWbr1QovXe/QttzpCl78unMy8ok
wbLHcWvEcaOuJpPxuqqPX1CCQg/kZ3FhsFz66raa4JnC9LOlyYw1espsYelubc40
zjy8ytPo6OI9r+fY0WjLSuVYyo6g+wJbx/GDzd6BSMu3QYBvH1YAOU9KPAKL+nWx
ZHgKpea7h4IV9CvCTYKd9Ne6N8c35MpJaJxrjwLo4fMM+3gphWyWDuan+1o7ht2y
zkdqTHbTE6l9BnU77GUYSSkujtHKRsy2qHQX7Wcqpj93ZZwvTCtYU+7NkudnAxod
5DcePX5JfZA0iSZ46C9Mkb6cDM8slNTNnSUJQpOzN6B+6/LUKgFSYOum3VFzmmv9
ACO5ICpo0eopTvXTaGDgND9owvuEF/wthbCaEphDh36twktRGPbL+joPFxF0KnSJ
WmRQYMHSLN8k1gLE1Da2j4kqZjaycu1mJiLBWzVk7tob00RKHzgQ4GOadBybbnuY
9+ttcpWiKUcta4XwrCTRouAfEk6VAB3BfZDT8wZnoUx4Cai0KfT2xo28To7MMVDp
hnwf0kKQ7X778rlnzik0V9UbbfnBliPZQSWd9cwpXMlHKXx4OgJSrWdtFH2sj93j
R2AxTs6dQzNpjWt/GR0CdfIg7jVW3iViq8ngoAlZncgsSwJuLs/xVZhC2oK7g50c
8H3YVdZQC9vKspror/g341jD/WKFhl4IAHDx4I7bIm5NK3ildYqOEZW02u2Cm1Cy
YjXfXWjHSuoxXJUymSRx6TCqkmDUNIEQO4TWBQhT0p55Sx4gCSbU10AY89/oolda
I7rdMT0zVldfxrugTnEl94EPzlUCbsjOWJlwLBUNiDZ06t6xPTbKoCRPa1QdekXN
Cms+KNO3bMn+84F2k9GqF+Ox1kKKzTwBgQx6MEp6nM5rlTQjhPe1De/fmnNqOibo
codne2kG8niRUmgNoOxJN7brt9PL2eCKiY3LzExBu6rCHBtNOI4iQ42D1++zIcCi
HFSNRZBHm5yYHoGMBuIAsGiZ5JLnz20pqSsy9P4eghLHMFT3tHixzABXdEmfv6E3
m579PgAdcJMxswwU6seAd7mzrGZJiIQERLtiHxOFXS4fhQFOQlV5NF3KdN5BQfdP
aWM2ZMXLp/gO8NRMaGsZIdhSfYqxUPK+qrvQ9mbTWBYIbePxxVH7qEbrISfAIXZP
O7csroWl1uizOOcVd3OosZnvjbjC01h0B35AKcZp9I8iuUW4iwYAFA2Bsd5qDAz0
Z3dZF69hG1TrusNUnxFqSdno5xgYCTVtkzagNopfRfVfIRdVhIpoDnBpcRcFOgyQ
Ty/RIDodCkBlWzr8jEzDXQJHm2KoM925SyCyQ6i1VavI5JWcJwBIQEejItZFuCo1
Og7QZufN+beYYng2tMTiLyalIFSg197TxvUaBARNYJvCJ4b7wzK6vkt59O+ZYtDE
uzWT6l0yY0ZAc3CRDWOiuKYL1qroCM1wS0z3nKYbgnzXxr5+GQDW4H1QDYRRr9jI
QIDbansVXsyadM/IO0kEtFw8lnVHKKMlaTy5UxzD9J5WqyGHu0WwkrUseGesY9yp
sbq9Xa8/ZbZ6CkJMqQe0ajhwGisSe+IYWlSPo9+VGiKUj7e2y6IU7wfQhvt4x3pA
2mB0SR0+eE+Be+PCDUz2F+vBtncW342k1P1DbKRooDC4PqSViTf4y1PXnbgSR/VP
+QH64fpSgdg9QdpOgXYSUQF6nCbaxj9lZT6ryDv2Klo1oTt2tSscpuo33gOKEt0S
54DVMqxV+mHiH2OBpsyaEx0eM1CN5KOPyzQU+r7oP+2VTdsUouo1p+gfYHblreIU
bQJF4KiabwVHvoC/8+yX94EQhOG0DiRbzneEt9P/bsjYkpYACRSPdkbEvOkxYSel
4QITTQg4BNcXKSy/XntNFEOhOk5wLFNnCWhkjkbvllA9HLlKzW6VlpIlPEOaWim6
4xlrOsBn9x/nJrqUt7xpLv4SodLYX2j+RR0oUwaR00jWBsD9s+BkuR0fIgw2XMWg
OHGpFdEWUtqjIYqH3r3wSf9/CTH7Xsw9e0u51F0SWooYJIL+bIVurciU34HOqSd/
m9BS6JyShg0gRteFHYd5VpsDBxqLCq3r6602P3/lmnxPzHhLAXXcfU7Utq18xABy
hlpKEccQ79mPaqRs586zU2KU54ojrkZi4qMHhoa7kJq6bay7N8L+H+/UvLjgINBB
zqaUWqYZC0IGt6wB8+3AoIQ5+G70nubaMbpf6bwukAuszEDUmqxTBqNUxkjvy8Rw
Lvyio96XjD6X80Qdfb3NB3InjPRSogLehJV7NJB/2aJ3wEn7DPfMoF1ys6I3qPim
l4yADEWheipBDqvpLS1pKEEA8TkqscUSQEul4BrHBXef/WKpuGr2n6+iPuks4igQ
IrN+xBd1F0hTTEmmVYbhjnDR1xReee6T3r37fyQSq5EkTTJb5TR6TMR3lYQpb5+1
pHyrB7WBxr/CZZcliOM11PoauAuu7Um3nxWC0aTOM3Vr17AGmF+H0Cp7Q89CnKrj
uEv9xs2IsNVRB7C76uxeTB7cqRg60s8eGZW+Aav18Vg/PG3WB2EAIPnmSc5r4bnE
zqir2eNl12iHoZimiV0kx2Tzw2jJ8tfdNU1KHQENmbaD+FPP8Hhszs1wUYCT+kdd
Z3+hXWbTG7hcVgedzumwVlrRlxAb2u6/Fyv0GYGsNUxTqnnSiNQuCy+a6frNd86T
sf6/ZmAnIuTMHtjVA2X03J1H40uac5p4GFw/r8jU+QF4SLME7HJLNv6BZ51kS8OG
NkVu7EBpAbeNPamSDv0QGn2WlUlz+31nMp6Q3wr09kt8RntyzR+lzPvhsCiGgBdM
yo5ihwoNzDh9hi9ctRJyGHS2jgF4xDxvqZtYciYPKvz4vNr2qVgXz15AJ3GA6gwi
bOZP+DpvDHfSZWky3z5fWha6xR8tu3yRPdMzFyOpL4R7nWFJOuUErFPbGj3xfcJM
Z5+fEmTvzIijvBXsk+UT7XlWzn0eF8UhQ9iPIFUXPQAydHHNuWwYcdIp2RDe1evt
ePZJF9exoeclTlPliGV3XXwR0GHEmT3n+xn8p+80MB05whl20V+UQgOXoUYkAvK0
DG96pZ4W9LAcBP+OPUoL/FAoOHOoHLfC2NmJyo07EvGIYG37HoC4+DcgplFik1lH
19S6j2MgMhb5PYBkABGk8UdDmKv6Au191uenRatRBgbdlD+c7HSgF2L5AZBTsn5q
nE7zksCmyb6bwK+uOgSfRKuQ+RetOwqCwUMUYJaJFZJ0gQJr1cwIsjXfqpMVXp56
EXS08EKj1zy9ls/9lGs/ZabqgjBUNiciSf92U7YsLeBpJrkVv4iywQmk+8I6/m22
cnZSTjPB/EypDBq23sYDpoczfCNqBQ8yzZ0a0qfcsKXVHxIiecUnk3Pa87GWQh0E
x3uIr4r9fjRCtZ221x2dF0x5hCzs7/ft6XzrBj4bmTJpMhPG8GM5U7R8M8pXtfq6
WXFgee3a0dvDs9X/3dHTr6fJHRvIgzgfoXNVFGlfCF8Z8OPOyYu1SruvfJd2rftI
sAg2ijSZOzyoALOLPciDADqZffhpdorgvB1wO/hVCjH/hT8t5m5lvzW84CkmWKMh
jjjE0XQ42648V3VlRSOs3eY3tkr1MlFb8iRF59RY89Mfb1VWFMGSxqSUpHF7ollj
dz/GShbppHptAoYQAckJ1+AnDtoHJDO6MutGMMdO5jhQC6zDxG5zB9hbiwpQIK5Y
woiF5cJcvc9MfD15PMP+8ci0iLjrnYd+XmjeUvFbTQWeRujBLyhDKpacMM0XELwN
K4/FKgwqZPK3N6HjKEJVYl6k4d4cRLoHP/5bvWf69DfZ7BvdvwT/wnLtySUawIjQ
M0lOpzd47sFUUX0I5CQhK+FjGmYBh5OxPAmoRtjcJGvIG7Nh8KTaPRnciUVAH2ze
CjCxfmnd3IP9Ag8AoLIWG2XlKLJgO5ztBDBE3tzM3ECIxVCiWarF3qSeS//QmI6n
uliOh2QxGe8qZOFSSP9pyMxmau2xOmQEwnY3eCz1DnseaFFjzujmO2I+VeACeJU8
NO+WWnwmp/e1JAi7h9aUBle4XFzLuwJ8tfZpX30qXwccx+a6sP6XvieoE/gIfHXU
XLkHx5yBVrsnt/c7pOm1EoRZtD+k9HKVa1BkNlgpekw29sxDSeUoDMaKNrVNegas
FQiNdE8l/BcFFOregtzFoEVT06tB9y/eWYRmCkbRPPpsC99KmFhKebpmgI8ukRVa
VLdyPueQz/GCQKTzi41jxWsrYQ/s3qG2QP6tlgT3twCa40aEpPBpgrb4deRlL2qz
D/mGYcwW4BlVCP23IJ8ytis1DzmCB3vahABQMXLiOvomFom3I99W7cxlw66zbndS
oJvHWj0fYVkalYLFfLZKUpR+pfWks+AMLT88+bbpbpH7TC63iUcQQq+CiMr08cjo
EVH1jdNWjeCUMpMZYLdPjhwnwvHPVEMJdFTutCkWNGaG/ZGC6bBSFA3m2VT75KjG
LoyrNNYTbRuFW7PBYOTvUSxUo2oqL555CwErKEZQqwZQ155wfVw//isktK63HGgl
SPyk/O6gBqknSA0dGKrJ/LgNvTOX0WYdx0+Op9U/oxl3OLyLnHVoI6shcPCzk3gd
d4dqOh+s5oJrTOoSnEX/x7ctJEaJkgEbQyAiiv/7jPtubtHDstZVPP2hs/tK7EPx
IRuJVDyaslWIpC9f7sS6drlgsDXB4AmV749sFnr7A/2nZlLameDt2AVnJFL9NUXT
9pbh2QdaZkWZCoRgWtYdu5DVqwhJE3wpVUvJO+jfx1Edlod949fhgJgHEokCwiMa
DqacENspbGCaozXqliJO5FArBbkKmyzUN7emyrBGVUS8H62UfugU0XwSFTYmvtlH
WVEEv0hKTBYb5ME+XfAo46+bYfvz7YA610vi7Bx6Xzef72P0lYMZy561EN/Nutl7
5VsNC7FNxwspOz3pOyJMbp2YzKem+k+afKElMSziC0cb6ACBTXhQdapFeI8wuaGy
jIUeZAdmMN2zVnqb9rPPBmUyI2JPjki4QGUMQMaOl9GhOy44G+yI/9sHbvSGO0Y5
ohkgi4XQpaXwOUWKtPecX+5ZE8OPkT8++2IJ5DuR4BPPWA+TC2PHw2MXy7AIKv3Y
b8PMDTJ/nrHJzGf2H3GBGwvHcZasBU+/3bFeGmEaDa2djuVEJyCLf3zMfAlkQpIo
Abn62YDFvblaT62SZz8qewe5zafmNt0E1wAsr7K+ymqcfDLE8O2/VyFlvSPtN11C
w2hcVNoxqdthEqBwJRumzqYGq4Va7V68pj9OzJRWCjbNy9YmeYgFOny0I2Lu5wKL
C/DhuBfjN5G9pD++dcQ+NRHFlsy0T1ZoK3kMCCiMLqHHdIXBi2YnmsOry5d+nxjw
WyumQiuhNEH20TcWMPqsSmUsDZkWqZcqak3Dp/CYqrrKIdEvnIOdIxaNaj7+UiGX
ttdJwFHD7zdOiIDMbloa9/eeJAE/3pLjEXbVMnxFqvhc6r9UXK7VfTCqhUPVFm4a
bgbfK8ncZ12h0DTiIi6ioqLU6SOBpKR97lzD/CMRSmxV16Ww9TadnTuQoW8cLqrh
vpuUdW2Ku1qtP/f9zQU7Ux2vJPssmMIJezWj64RP0AqFgjpLXxT3caiuDB43A0+Z
Xtlxh8WtVQXpAVquRmIhX11Pxi5ge7WdHVHfTL6CI2gkkp3lU707ftk0RAu3TEf2
6OYD1TDt3EF1SIDeqKTAaNoYs6JET34hsyb4MrjOQGnKB3i+Z3ThWqzKiNtP0gE3
BwVzqf8zi094NxLM2sKHoq+3Rw+uPG0s6PafY2pJ/HbOnTU5fJSX2TGDYfDk+dmi
nUxTa7yjI/of4VfJMke4epJIBE9XFbw5go6GP+REcGcR2Um04jF8ZYZ9AxPj0v86
W3UWX2B6GE0lRZckiqAzOfhMYuZtigh8w+bLMKQgnrAL9ZgDoU93oRl9FRvLTTg2
8otr7QWsdLwSRD+aoioCvcDZOjxNVFpy1v9KOV/7Rnl21EtRDzAmPoVU1lMarIGC
IVnFpWwZqEpeiJyY7wIIJ/oTSMvwnd3rqnzCga5+wloi+U/Dd6kAAwWbr5sETjfu
M30n523Q6jnZQjitJuAyHTyOsGY9IR9lOExKUX3A5lx8yjL4JWAUOJll2W2vAF+b
ySetUf/w6m7but51xKnmpcXolBqXsG1ipr05kZZhigUc1R5UzQWem9E1KvXTi54W
U5B0jJ9+0fu9pKpEwythPsyMi41u2KQz004oKzpcq9xRJy4etBO5yiZ4evmvlrJV
KYl0OX9sMz5oVr5cisIAdVIEsqRhK7Bf7cUMnUtiRGJ3tOnw1Bxk/bbg2lsIMQtb
CWCuPmJS4LOB3B1fgH48V4v57HgQwzXBEdlIwbxs+2oEg3HSnXJrQvSB1AtlNhn/
g1PkAIUsPXM7MiWXTxljRZIAEp3KNxogW2tLdGMPpqWYevvPwXK+MFXc0MSuzbrR
pI/p+v1uEpezCM17IgzB5Qfd1Bm/xkp623FDGJ7Paa8J6Hf9gAVaWjo+KTcvcXm0
pl4bFAQ/480fVR5TubQSDV4xFCF1n1bjS2UA2fdCCfTa8rT+l6mR0Ms7pL3uRHh8
IRkWQj6PFUSq7OWsgN/dhDYlZKHzPgQco1GnsluCZuv/nHtym9MhVSigUprFwSOd
A3qtMeUL9DZ27oaAUzD3vDg2SIcZT9C0rfYsx6q8ifiUEBYjxXxSzQ1wSCJND6+a
lFzSDHlM6xOFaBDjRvfE3XFPiBsQEOnwZv/0L3SrC1wTIMdxL2tVrEfrhU+Lot0L
0BxcKqdNDrXAEEWo5o4Vg2+zLz/MXDnlsH4SjmQ/D9DXYf9SbNdCdOcYSNCt/5Wz
dY7CJrwWfwf8Y2ZaY7/+Vq/x97OHjfRvkZeSxQ27433dRmAWSYt6vYNUU3CRpvNo
L53sPW74hddiLnqG6PZcpcEhkzkT4phcDiDk5zvcFEvXn12MYneBczjJp6hACC7u
Nf1mP8rw3QyG0tBigLreZkQ/2k0sNXfNCbApBxg44t9O6Nks/KI2fRxPjZM3u3g6
VMfz3po/pH3Ah9mQAOMorg5WkBweOHSRF9LpOYKnocH/7h/Dwp9kXnz7chcQPFo3
yhFDxiy2ShuL37wIa80pSBQ9nDs+e79TM2Cg2EgbQtdSuqmn7OmbCAmKfPPoTSX6
SlbwowylO/zfzvScoWYnMWWRycxU6ojhUwePc3Jc87YFzmTLKrXPrIe88HoGwr7Z
rRpCLFTFtRmt8JlTjwekrnO/sk83zm3/iBVYo6b0A4CYuojPHMrZz99K8a/tGRhH
80uYsauvRGgvcrpXJdScX7CH1GtcBvJpA5xNnlYDpnhE7XQoC9kaTlhAfMwewgMf
NNJBp3kJEySDJBipywLcsRkkwes4Ks8YT07kk9A3auZob1v7TWlQoC0hfcAbdvs1
O5hvW0/iU2pMvcuFku9k38md/xts9cJeuE+CR0XDOEpM9yLU8vfKphD6UrjYdEeR
XUs7l1AVvjFidIDRkE6llWKrSiaWqTL9+1DBXvoYg1YDRcgsULcd8MYikNZZWKSW
4dXgpSIcEKky8JAUldRRJbF8ejZ4DiGDQtrFykE6ZJkubzXe7ooQSlmQmYNzZmhV
bFrsywXph7tyt82SyU5k0UP0wlrrtgEzaKjICIHxkGrCNBscvZA4xkAZ6t2QXpG4
wt1ibT/qFhnVapCcRQfRdzL1pO3cA8w7Vm+jBVOrYT/oUmF1wbPw7uoSPdcqGqNC
WZWUHp45MIWvMM9F1pGUNz+oYkeWXIIrK+IQq0VEvhQYKQzFcP7qS1YSRiVPWX3d
D2FY/OfKozJ4vpnmCL3aRwm7nxt4mKodyLn0MsfbgV3q/uON8YCpkVJ+yJvuT5nV
kxfGeBSlVNpmLrjvfV95csRw0CJ1RJP2EoEJOpTWlh8XVKEB0dKYL/mcxGzkEt7S
U5zHGdUjDfkWpa9EH4BKu+Y0mNOc7Uk5J0OFL3wtyYVz1ZqqtxWV7jFhXkIeUpLQ
kBu1ziMTEBBAzarvGZ/jPx6kPgmqPAddAoB/mSafGPIR2kYL0toShduEx1RnsSkB
EBXcR6hms3qsWG8Y38Yu12Oe2HbOREbJeiDU4oMIqe7UFngs0ixtoB/0FLopMb0Y
7deJRdsoDwx3gSwppNf5ZzaXPXzNADpL7DB/chZWlNE37mo91qJRuF432Aq5xYuW
r+aUkpV925NP/imBFMaqm6oe9jwTH9gLKbxglNYtk5uwZKAdNAW3InEu9Ix9Rykj
BrAjCequTD0XOHS1IJndeXSg5iuWH6zf+UfCI9uq9EcN3uK/APhrk40E0qohEP/8
sL/9nDYsnLb0NEAJd5sSeUtUJ2eM7xgZ2/YC3jMrx040hUVDvp4RYnj58DNNs9Br
9POP6Saw+cYaDae8XYJErKKcOpzEmDiGK61vXepN0DlFKeMS/iTbR4XN+WRr0Erl
G1BOAiSoJATAZ9VYDzzKTpm25Ky7YzRWUSEcieD237kmrgurPeFWjICdA8rOTVoN
0US88d1szoHWNqvEhfz1nqXiAxGR+nREb/YZhhS6zOIyCjXDnbzMDtE9lVFbBERl
ifRmlAT9sjzDJuoq5CvwG1Q/4CVqEsq/5oCfZoq41glCRC2sKrbgd89nT4Rhi+B8
BpcrNLduj9CqTIwbb4u6GEtEsE/XL5rKiGWznYhBKoOc5W7y81dWud8+kYuRkuAM
8dEnd62qC5Qb90YkMA8Oy2yBFakHwLUG58+8ugeUK9JSbtsal7ICvDZihlmRdUVC
res7qKO9FAJ1EgD3QXbIbM/x+r11jQ5QMPq/ZM/TFN9Ax5kmqp0zd+gzKUUJBuPJ
52STXWCLN5aSae1pjh4Ogp1f2L16JZVVuj9QBgzG0JHkhEOOmew3FmeT5jrDNnzt
jwjQIhiY5qFkm6AE+9jfrJR255SIUe1GDDlq46TlgRsaXv0LrXGKMBseTqVr63VS
VegucyaBj4X7s1Jrfz5wv2BBLPfxD64JeduioQrF5fACGC22ldG/4Ais6VYLssy+
8WKaWHftKd/RTboYY80fJ1BOokXjuWh+yaoGF3T4c7dxfbyygZuzlGbd7LHeuDpd
KbJZK2zTx8ub+vrc29+SXEUPvzTwfJDLHxrIE8qcR2fOkOpcM5ur8QbKiF9ADA9s
MBH0v4NibwnuVCpWbV7aPay0VwbLLJRtILfKMTT4bv8NOwju3ISRCwG3AluAod3y
A36qOEe1JVTLXubdgHz5MQHImtkhEQlpE9qpPUR4dU6UJmc7w0SyUSgrTSocCQy/
vzafAJcM72ibNWs6f1LCbJA9Z1Ia/zOlefeeX8JnYe9nzqZLu76UhceEilHRUQ3O
LS8RdQIwx0lphKwINLeJWbEtdRNmkYMoUGwkS9vIkpnzOsE888xU5SQibvuSca9R
gqgo+qWAQpc70zqOpF23CMwtKk+Dxj16IlgSfE0GrU1cFkELixvI8PU50hRpbRYX
k54Y3Kt4ZsDfbj+fnezZu9K2DdfXEGD3mdGQM9PgLbGcwVULv8ipb9SzT2HXRKGY
uZ8o9XP9xBaqKA5KZaybhWeAYcS0NL6KAXXMDq/oKXpLbrYhKafoutMn32cNBv+k
yKvDHel0mBRkRX0FfvpkjDjUMfNr3pItVNZ7jVOTk5gy9Y0/JQZkzpujy3OiLNC/
17szyqHi5N0zazLdfT7vwfScHdnGycn1In2uN+Fhc323kVKxvVlFu3pCKHdH0/TL
2qalexuS0XbD38x8hQT7k4f7WSU0mdrlOa34sK2Z6F/d1GLQqhdYGwX3KKai5/bX
KCkGaJmnbqyab1LejhYxQk9hyFJnQ2g3AYJiqghvQPWKvhDITxOfXwQIThyGVXRr
zSFy8445YpEWe64aLGafoO3FANAaU9jW237V8FMP5w5vDuxEx+agrUw/WRik0zW/
31W5YCuImD0om8rdz9pnGM0pJtFR4aJ777MolQqB8lgBdLoPzKBt55UV7fcqXzXA
L1cbJa3VLCCv9/W4cMXZ+w7W9xK+sKwkuTjePhMDYGvj2wqJ2OTQq7fO5fTXcbyg
Wj/sxSLs382pC9/2yT/SD79PWxttHX4AB7YL03xyVzbWzxCpszZzmo+vNZRVqVWB
4f8Uq316b5aAjl5mpqE8BujzlI44ZAX2tKOze2CjIIaIbRkm40ql96l6tox5vHBG
0xvJ6vbMlFJPmtib1XTAcXDRohJWHoTWRH4iJ81FlNkyLdcxBL0/aCzBPB26Dg15
twQhL6RUWnyHIozJL2soYrm0mLhGE0Ai3jXHN3HqXFMh0Fbp9MJK2wQ9Jorrq92R
lEKj0n7dECWCbDiIyi8n80QEVI4gjCo8c+Ir5UUFn73/wSElx/EDIBwoKVmE1JkL
K91wbR60MbbGxeV53ZgP0jdUDFqbpitk8qQxR89q98Z1vPVAFSS4e9RGCCn+TGhc
NHy1TBzqtSkAmrcrz/47Ibv5eKZx6TdoRPD8KP6OT4onmKxmLX9PZQ28t58+p0Kx
fPGSYjAH40Vs929v7gcf6xSQO/0caHp8vOtD45NS6hYDxukDo0aIscdSQGwgW3OX
Kv860DmTjP/tYT13sGu7kp3qaBjr+LsJGmIndBl1GShvHBHj3zVXVdTiNpU4LtxI
YzsexMZpeBuVM1vrwWRqEDQ3peDjOfH+zLDUwQ2zwqzEjQScv3gwDNPgNmpvd/vs
7jMSHTmj6bhsO5X18D6DWctmGsiHOyTZxCv2SR+6crWq+5qojM3CAHHzsZDsPyF/
PQJ4Bmgb4wwaXhNhj8SGCWq1TdgKYIFOtN0md16fLjpwEv2YvgnoOfjmbmbiOrXQ
lE/VTbEmIhx8G183KOcLaPvvX0eqm7ThDhZyu8Iq79jpxOymb705oWnSoCKU9Y3t
vC2+Sa+KwQr97bUlXbNvkPbc8TM1KiLu6NgQsKEOFHrLJgS9Eq/ckRMffH252JLh
YALdgwH2akrA8U/2FGz5aYOBFKJ1i843jNlXUbzLWkTEULtIKlHEn1R1MPL8C01l
JyAvtnsT3ZfcThc7HfX0wkRoAg9VitwvMAJGDNxQmF8L3G4zUVQrZTMylZ2RlQ0Y
g7Ppdgx4idBkV8kS+49BFAOwYEoweqvVQrCqB9MQLKW7Tcj55PZ9vI4wSgMZEY9i
WT9rpFW5FJrmjfM8voOUwTtqpOnFiHqCHhWUbzCEzqBmLMc3cedjIkgbdn3HkXxg
8/RGFXiu9oIlyKf9NAX7QwKvhaD/pj1+CyXOS69GHHY3AcrKrHkrNohfTwiaI/5u
OU0huOMfhiyJyqXzpqZ7mVGt3U1ZQR6FgvY3yk+fRGQ2pIseUraoNa9jEP2DHl8J
wFJ2Agcu6DmQ+bwPw8j4+74YfBT2xDt/nLFegI13pVHLKaK1t0HNZcB9M32noaeZ
1J7O6ZrKEne2azztAG8Vr6oc7K4mXHWHsKJhAgPjmah3QdjeItnT132nkkeWTKn/
c7yuciMRwmPjsoWZcFAllMmId7xSqZvCdcjitdbISs7tctqboDqMwl04xDw/7kcU
VsqSWrKPOPP5wYk3X2NAmJy7GhcX6bLlY4ObfitpNhkBMSyqW3VYuH5SsQMkBFw9
b1ybj3gLUh1UmoIYG/E9BeCsoqLFypSwAqqfcrPVUdGfwPNRc47YXQ3XDctVrVJX
WI3mpJzt2ouR0irTp/IPrVo+Z9dtkeOMDLt9Jqxxk3ftbO09dhFraWVnhR8B73E0
Vd+wZqxIe2+/RITYVFH9BtwYc7lOrkZta7SMKgc5DtaErUPQi1OA3S3t3OAQBIva
NzZufprJAaDSlYzXcD/Vxr1Uf6lBuMPOK+JxvmIXh05JEAoTftXID2ROop8Pbvhn
wCIHb+1VhhL/fOXM/eoY3iEihqwX4kZUUTcT/ZLNXU/qtNH3t+Cr820UMosQ1uSs
SCUGjD52YVJSe2zo4BTEUU5f61KOdgB3VoRh+7PkmLbKkyOd2ELBP3yILowzlpTD
RmOOA6VxO1DOn2amV+/T6rnSFwednBnaqg1fHEwKOaYZcDxmLbLBokhrv5ec+h3d
xX1+qSaPqvA1AN2MHrYyv6d9pxsw8rTjyvOMPWSbmXQiT2yjyyDpk1J6bhSF4vCq
EOcHDtaW3xxnxaU6ln9eNtwJp4NvD1AsKnBJ2VDT7xGDnXR7dZoTm8RqPSy6soJ9
vhgGM/1/w3avNOVdKVdcdLV3M4iYc9YYcFbx7oFHaxjg40CaPoIYog7lZLh8ja8N
4AAsNH94pecZGT0StZC02vIrGSkt3JVSdMgBU4FC3DaNeyCLF6xgyDI896GQjldb
Vl9DiMxjUfcZiIMpANl9xnwRWF0lK+iVqDA/oJc1GXL0z1nh3r5oIN7RVFVEOQ+5
C3zAjo3eKuVWO64+hFXEKcF+XwUYdw5ssnazZhOQW/iiqX+WLwxpuU5M75GZsRxI
VG8HsWLVqUJ6sAnINPb9+eSkY4AHtcSrKV7J6LJUe6FI2jHm+NxQnHn2CFkTNmof
ayiDxDUOnqfaoWNpwaIdRPgAsb3UXqeEZ8E7Quzvz4sPnTHpZcoZLvX4ZXtADFUl
kG6zviqbfu+OfUscSs1JySEjBa1rIDE0v/u7ybkK3KGkna/XarZvN868x3nSs/2A
TySfoxZ/ArfkZ1dfXEU2Y+5DoLsC/bBl+EP+AeVfD/3IhxHzwhs+/USP9WENhIU3
2tcuzVTGPklYpSDAbWLzqCQadp+dwK7iLdaB+QdeHIGe9EDpzX+R2syg/R3/7uR4
UpnP18LotlYl+B6ZxNO9vv1rq2XnIs9ov1INVSwiN1bhregm2/I4HOfhbhRsn1Kc
96XrjjrNWXmivCxw6ztM66WvFbuEIfdtVXMYstb8pES+SbonZE8mXVLj/qF+DHwy
LcoR2dnBL3Incq8ug1XdXGU6wFhEHgIgrEkLgaB4sw0WhkGnqp5jAONEeKyLQ4AU
47vizZx728zpY9uyIjVqlgo2I7b3pS7XdBRiatqzRm6vFigBeB4rOVS6c0f95Z96
4Ni6L45mlrNAtHkMUvQVIfYn+L3uQWzLnVhNjPgbf6gYr90pJn33fRfHLd0UrEIK
bT42pL5I5bz7BGhnS7ZKyp75Wf/NZd4BVauMs5CjdfZ/LGgUbJ7otO1dilbHOjKk
TwkiiLZOHuzESk5nbM6OzRt6C3eTQsOhrCVY/if5Z0MM2VkCTA/eoe5xOZc5bqnw
a/9xxYQisMnOIdMzJBT6LG6iWSonjVTYw8WiKi4I90e5p1eR/7JhnU7qknO1JGLB
VfhlkRlZpc6BfDCRYIcBth2GBuWI8Fde54Tdzy+n8rEozeYKM3uTvUAN1cYNtBBA
maEIAmtZILt7pe61vJ/gBrQ5ZTpDPmzYDHPoYovUunUdqyIXTsS1onJYMEh/A2RG
N/E9z46C1ivcA7fK8kDcIdbWUnwcAfeJUe+4G+H+wruNiIoYV1XUmB00VREd+qpI
fm4/0IDzU0MkOidpUtgqvX/v3toZdwNzNOmbir1DyRCC/ARcCAiKjAhr2Y4/34jA
O+TdQrXo5kH2QhwVoPL+O6WhOfbF1oYwdKLerkiBTUr47SbA4WxjX7CX4ci49obv
SWgzKFQs0rkhE0k3GLqvgUYVFBU4jbd4s3UkJw500iKgpL5zF4N9DpJjfDVf+wkZ
tfzWfEyRFC43Agm1FLUacV0Aw3Unv8IKdq7FPejpkAtJ5A5reiOKWwK2bBViZB6K
XwPepVCwOPx79uPynjAv2s5hpiPLlScIyxWl7B1HvyZR2GV6t3Lk4YrRWGuYS/4K
Ubd2xywDWAaBDib6xwZNyr3dkFHR2saPMHrVL/xpgkpJtJrKHF1SW/ihquEhWh6i
JmbTpUM1O1faLTyfHeytUckFjiM4dKSETAn3oMbZ9MuJaaViTdjWgUMROsIUwRuJ
Sy3WzUTsW1cp4Zw0fezd3mJvEP8rLHRM+Emna/nvZ6iPMZLfIohP43UEyaJxz5u9
MGpUnnfyCCQzDdW7CjkT5zAG+eOz1Ejf6Zs/dgfnFSWl2HKtHtARBbt3BaexVSSD
12Se6zORUzO62i9c02r34pMNABBER+pF0bZnBKL4yxAJhm0ea21g+pkpThDzJd+1
RwFaR9cFy1SppNaMUY6ONZypVK3wHh4/0jCaikiUeQ1KVVJc8tnbSsfw3kiMSPae
gDDIRaJtGvs/Ch9lvIFQUy7zw4H7zF3qxNPNzFRTX6FKiYrDsiSGIrCNTjPhl5c+
dj7qydNy7TVshsGeNjeZaNfxkSRKR1e4UTz8lbcJB0Ed4THgC4LP9/Jp7/HCGSay
lb+7OO0IsV9DwCdaoNAP9CZYSVRkAvk7iycx2j19KvR0X0by8Nt1ao0t82uabnZt
IKTInzk/sBV5D8zCLmRww2/fitSCfWv3MCSuMQyx7bOg6QKG6V1nLiY/vJYBXX8B
T5gbIZbAO1EPt6126LAya7ezDBO5he0k+QNtjgaLry+3q6nHw1cq2pHUPDodErw+
8LSZyIpSFh1LmaM4N+hYN9LRPOxsx4TyIfnNHwVwe9f9XOSvkis18LOS57jDEmJn
2dZ3sTyJsz11ro8Du13xz2b5sAGEzSODTugqpgyQjGqFSahVuXdjNvOA3TMv6BZS
CWG3fVYSUWJxvNGR+aTj1ymauzX0o380qtRq+DkSrUST++R0EaGWD44jZlglVTFK
2a6jRj+cIvwivGNDOyeEM/j8KbljoMyPgv0mUapsBG/mIsbxFU6uiNVRwd31uZCO
6zKxnSgyOeCPcdn6XdQdCQZCDLowN5vLf82Q5brwSbmmq66B72iIv9xg/98I9PoG
BHoF5YuaQdoThCCygXNh3nQFWlCqn/fssG7WOEqI/H+LPhAIQ2EXLFEkruRnVmCN
XTS29WQfXpI02gdjrArf543XSjQ84lhAfSX6G/XcrQSGJwJCI9HSJCJM2SrghJux
gGpIC1iYwdkuhCLhLnNEJiLqKBfgIKRCAUtOAPf9maQEcrh1DuMIU6P/t71vxs7z
sJBQlbSs3dQEEvg4/ve0jORqv7YvjaHZ1f68lEj2Sb3PGQ+suN7anf1cQAUsr9Az
e6MOjKoR+TcUjbc8m7c0qXZneUS4B6PMKJqScLbTatDKCRo8E1578msq1HLuLGpi
+qvnqLeIZRdQnNORHFr76r14I23hDs8PIK3HoGK1N6a1RvqnLDWzsH7tLEw8kcgr
DbPegbtoFvlbJ5RTs3qZVUgTDVQ6QgosGjg9Uoy1wzfVkw1CPJM/147TYa8ktmip
WUBwbnASHg80FTWsyxeOnEn+jhYYtYPeRJCkEDW/YK+onZ1no0S6jOoUXJJVjoLs
/UKYNzmAWX1A0SIwbMze0wEhwf4+s7QBkVs9CufsQwv1h82fGu9k+NagNwo37pNY
3bIYvWSkhLeukS2CSYlqUEigjZ8t+KEzBm7Gpc+VKOBAYOje9skeVwD+JUyT/HY+
oY8P1tXR0KcFweyDuGN3DinC4+kKvasQ+V6A8d7PaxWM3klre3SVrWQBAIjTkN9R
YH0Dy99Z8i1s77ozQyi8RRgHRxWiQ3pdWvP7PYASu6WIkqaT33EBd1zEp/XfnSYU
H4KI6nHXlfRk51Z+5UGDZJESww2A3e0jJK+xq/H7je8MXTqO6HzkJwM+JGCaDUdQ
0MeInIZ5pFQrDKwrJl1LM5g6lmEsp0OK1PcS1ECMOE/BL5kFvNaMVF5JwVEvjvyJ
ywtTcUF2LcVLQjgZwFcsalMhqjo8+rLAMqc+TmIQqfvjQ5EHjc0MlVSZnyMqzba5
zzp1Wahh92JhccE/2ZG7IsTmxA3L2BElpQF+PSOdEXgj807ZIHUO3fkm4a758KTE
9BuVAGGsWP2Oxqykl8LdzUOjqzYpjPSf1MnOKmzChzp3m4BKFY8TF04WWZTk0qlS
2bqsdN7cvCXtY6z3ZQT2YfGh6GyEORE0H8xro1WlRnwxl0OEBBHqmZsnOoKNzlq0
zAL8xJ1MiR5Yt/PUiFKgpN1a8L8TsNVZ/+5MVQF+p4LebXHFQl5K3CkTlUd8/sxJ
WOFBgV0XLDABjtgentk2Z0hWeDVr69ZMgPlQ1UNRNsJsE8M6Yc26MPAZhfcFUOAX
v/YsgLufdxt3HU9czs6UHP7mljcm0l/G57CW8URXFBEzyS+Cp+Xaa+vi8WT93R5x
2x1V5dCe6hn9eVjtQ48chwbCbmsK9jvp27QJPn2o0B0PW/WkKseIVxp2hmPWF2Vd
nkR//qJeIRgqoKkuO38NRoFi/Bqjvo+BZAIQZInEwvEqR7ZsjxNrB60qpUUuN1mz
XsEvCtVj+oVGi7spGKXmfuHrXlIolisBqYzJ7uUE4BYFXStmZHBEQO1ruXWoOHbN
B7jhgXdIchFGFETTNTFSZ/xLVXlp4MxzjOQBH9xDWCgwRiMMlq4M4K+77+KYgRa3
mOcwZx3lOEmADPurh3kJ5uxtKBM6w06tQ+SLo2t1W+OYDdVpCTvqd/x7qHHTSY9S
zJrG2gFDV1hK0f90dkra1bKfEa8jJnRnU2U+c2k1b11cV1WpDN7nuXu/rWxOKfhG
SdsZ2hFSRy0Oaf0SMiGNz67IRbcQy6QUHpcJaijINC3OUMcAdM5QDZBlJrKqvePd
X/Wyu8Uqk52NG4pdG4bZYFEEXjQ94T2ZqC4jnZN/UMja1fV8XsPFOQKuqQMVwgpi
OFKwXZ1NSWuun1lqs2qryolVWf4tRLj1GxIkbad/6O4W0TyitkBGhRB3USdha+m3
QAHci10uFQiQZni5pNlSE6+oFY3/SP7cqyqsntwoOxHAd8GpHfodbjb/nIa5BBOA
K/0Dnqa83VTI6gzZAjydYr6BthiU35Ohuo20Lx+Wf01QKaIcYF2Be4KhWlV6pGox
5shlywHk/YcW3By/pulmyOpHD7URw+CIsR3/uadOMB65JTUROvbDihx6g5w6U3sx
/GT/JgED9i35C0myi0Nth8yoUdsb0z/V5oYLEjIwUPNbksH7vq5uWADMYickSoMW
7v/KLakvrAtH2o1ldQUURXGR/tHvA8ON0s1alayEkM2wJimhzb+PUducjoVAuEdi
X08TwfjsaJahFltrF2dF2AZqWJwW/8F/nlsqw+CwnoZJe8QEAyAEx6Wkn6jOXh03
Dp5thsje2M3rMY5yS2hdQMDrl1zI3/2sEDrgpqtUZEPTodDCfTgYt7XzHBt91PO2
D7ra6EfvNjxRLfW68N2I9Pys39Vb/g3Po+/t1LvC310ALay8XGQSJBRqJeqCVasB
pp37FQlBaIVw1QJTGAQRCYby8ycIKmcoYST777QQW/B5Z4Zep6wMJ9S2xFDqCt2u
/6wYoSH0chCcCfzeNcgHletuSISg5hnf0BSnpnrToKI9IHNByXRnzsmQlrCyA/ig
XZ+soLLTsQw5duU4SMOw5b7fPX7iCHBK4LznYSI2vwVAb1PyoFlmqTQnovrXTzOS
Mzpk/3WssCEXda808oNV7ZCiliFDIko3jAM0YYlQu8knYZ9bYNEfQMvRSx3Jx5au
ErVYn9dwtz6Pkc4XDXVoOmqkhyqsvOhAWHJ+ZCVMXMmfDkNRDzUbkYuzz58win7N
R5k2G4mRWifoOGVvXcNleBrrO7K6PwXo8bq82RQYy5T6j14fjm9zil3fHCeS44M4
J+ZNNTsN8/ZLbPslkGzMZYUZwF45WwMyYGI5xNJKzc+01jZD2TK1QClRnjLlsn9T
V78MGMlOLkqq0HUlSkrLnl3Rmpi2MO1rgustJL8njwYM3dRLubgG514SwscYGaqO
9VxxGNYb0bGUr8fpOJCTADH/OpuJZ26vPEs0AUKuMDH6hr1cRGU3aJEUUTgIOexw
1BRQAq/3NDYb2scR2yX+U48OZZzcZGXWIExgAf5XhddAc5ng53tKk1BIblLktfN9
mnB9OFLWF37qAvvG5msJPhubtJp+ag3aX7910Z+fyI4PbeAoJWNX/Luico03LViq
mcbM1LTW3ykwwlMyfRFOHyzhTSp9m+URJ6IQzuPUDfatIe8gjBJ5iMfO2Ynq3jeI
aZg/5d35qkD0zDrk5RZs0u0a7BITdLoaILiWaceo+0ZvSaqUhPc4pD6rC4V7bYNY
fqdNsAsRTa8vGN4w19LQ6KYNkwHnFSMbWHpLmM5wOgNpnuNC75Ijyv3QL9iX1z2g
kP/1Kkp1dzBPKSBDAoCQeL63V5GaAYIjOE9nZlD2ecxh7DCCDsFXmf8lbuPB+Bv+
JXnTTz+QTqFnye6gN8aHNXnTNqRxjI+Zk4r7zbVF5+R+7oPxjCMIqs4qDbsb9Aow
4qbIDR0uJ9lomnDo0tBPm80IqogiNtE9PP9vb0XuqZRoD3hq8DpgjOurDnd+zmTo
JV3OaETk1sVI4SI1LwxarsXajROwt1B51w0dmEOn8dYHGNtO0+xwZO7A1Zn023ii
wyGxGjByPjrcbXHbf+11dbaMk1bIHn/xzEzfHmJbuKwpWvbIfOD+Fb24p13aQgkl
otz8/wNprFDHirsZRoTy8Ep+PyDJGrSLicT6XXgBe0cgMLilMSqB4sfkO3EdImo3
B9627cD1crWOr7GkpftXUERpz0gtDyXYzCD1/9poEqP1DaT0AEtBQsMPE9aF7ETY
Jm+NbTJ/NYiAVK773NuLMghfl0XA5OXLCxs2vfBZXr4ajaorXA9veE47aYWcaYVO
MvjcpB8LhG6kStleEhXCIOHIXr3XVQyuWelRJr8N69sMN0o44QaxiIN2t2CUbCnq
DcSlN5GvlZGrnOWCKBfXIBA/a/cpNd7LwC0MzWOkArF6E5N+NcwXr3dCTxDDZN7V
xOCjYw11e4mwEdwOcIFvnoRGzOFrxjrtLjtz7ubDzb3cIkgF71PlWtasHEHnmZ5Q
ld5Hl/krGPQI3LTWP9tgb1BeS9B1wdT/aPDNIVhDHSiN3nIFgKH4jDRJAZU9fESJ
EPEsc9sg366xrYgWEcfqEyR+hAw2PzRLOLrxF+j7WnbOrQvseb7AMwaYRnjVR0DC
1Ww4DQ27Xfmd5aONPu9N8BcPZ2V12VZNPV+pMZf3eW8dfRTUJigx0qFe+8+NR5PC
V3+LnLt94I4OafyiY62Ox2IvINE28gJB1nIZpSVhx1+sS7Wur6S/I1dzQ7dU4GAS
CfGYceXjCJC2q8vJqis6vmmuT1U/mGrfLvF0YIrqDJRCvzoLJpM90XOeXdBu3nHv
3XVl8oHtTIDItj6X2VxCeg2DRMO+e/XH6cXqB1bX/vlVZxS491axuA/KrUSLgTWf
z1eE142oNEpf2+GC/iGAbQoDPzD5TYKjcDMuLID5uucK0pbfe1bSgCjXZpwW5Eti
TaAvnyYOGFO5ORGp8eaNp4R1/I556LXoxQRgsF+7zcsSpWhaV0wGdYr6jUPIdRcL
clf/feC7Vqgl/afjO219pLwky3nsW6VROigZOxGVUuj3NfrO+DpqiZDI82L/rH3K
LMlNoasHi1rYYoNQwHl59swU1jRsFt9zcPviRt+cQvTUaqkJ+nV/Lf0wumVMYx94
On3MW095kvHGqcXbq8NR//M8pd8fdVVe2TPDJxrrpgl9wzVFCRkcKUNRFr44KW+/
UImFfr0kIiRBLySuCx6747pFm35ol4lDUvfSLkEfECo77B9o+/rPmRFAfejoqZLt
iz1qABdky1IA+R6/Q1vhHiv5MdwW0VsS52hQgXZ89ysBlFLlWi9rzpWyZ9qBKdHm
xwRwxwyGe0Xiwxk/5lN8NKLniyBT83CHLTTgMGgouCPyj3KK7R7FkxYTRZ1yiXNZ
FmVbg3rI5ayy2//+e7ycr/F83SBrswrF44jpLzrAUtSbXdHIQaX61EzjIClvc9QT
QPWe8nms+AHoyWYmU0DCs1Xk9iwOdjDc+X1HjHzxs+oCnMaXY/SwyjMi5VPGltht
FRfWuNBG9JiX0l/ZfBDW0syYvWFKtHL9KoWBk0VHj6Ehb0PBgwZPCvnAYjAKOYhZ
UgilCxGK/Yj07oqwmxl/dmefiJk+1vaT/B0GpxMfOg7u8OLJ7ve0OV9j9xGNin6h
A0ZVhjn5yuIxdfwFa/+2JXas434LAoGS9y8MqQbbcT+uhTRr5qhaoKAz9xNniG/+
aIuGAYOeSGqFv5x1UdBW/JWBNBfyfx0Im6gCEICgc6FTMg3aaPQrNjhDcm2iwAz+
oXDi4fV3pk12iNGVnKRs/Qd0+QRC6+bZcnOOPZ/lqmFc8kh9+VmlRgP7N+VAG1Al
SoEMEvupPzvuAI+TOz4ZFv/QovoD7xgY7WNYBJSGZPVu1/OUofmed3vH3YraWS2G
OeaDkOyqATqR/EQbhpGA09yr3sZFBa70gq6Gwu/7Ifegk9BSutaaG8vv1sOl6vrP
lwr2U3WFQr41FCuu9pNCAg6tx4Fj038Ok+9Bo55iEgXsnhmLptQG99FF+BbXzINS
T2JZoYQu/T7ZV0HoGSjopiJX+BPrSoYFLCcPY//xSbKs3I4tPWVB+VSM4/yXplnt
FnGgTLtDW8AeTTx9pvFTTtD6Iv3Peap3y1BORWRjLbtvNOGTBcHoEujB0ljnpU9M
4ix9PxVReSSXhUCqaH7ZoI7BzTXP6AYofmiMJomSrV+W/mIsqpty4ufSlTKrtkFv
1FWXiJ79Kx6ZM2ojW2lmYFVNKxhdQ7uj8E6FWrntHNJk++DqF2sCTXK6gAEv7yqG
hG8Yo4QHmDTVWluvydXzaHDQOKYlDYlB8OpfZczaKAiT5nue0z4e5OhZGTNpDraa
TwIFm5RQg7FWHxUXUkuT24pWweI7scvOo8gHaN9Uv0Qi0kt9wul3pCkP2x3h4rto
K7i0bpeR5TIQxBDkscAuAtR2CE0cRR+2UINrlk7M42/yFj9650z8ArvK/R5R2JZ6
5jqS85ExeWsK+q8vVDE8IvJsr4Hsdpzfk3gJdeNjVo+MzJ/WVmqAEk3TtCxig0vd
WUT0FUIn41fp/4EUZbZzEiUSs2pq8T7G4V0yy2Am2gWfp4rOAvfd53J1djRFHMG5
THMacFczg7vX1C5YTf6oie+iAd2xiIiRL1wNjs9hUC9XDd5Zz990Wop6NX7RwGAw
OQuQQ6zthWMrAnhzO3zpiVm1R60vFFrhRaR50dnwnXjuZi/vnUyo7SM9BVn6CpFL
htgMOWlZ69lLNLH9mQreu0/bIeswUlMtp5r0THRBv1tPSKUN+jOpUCQVtxeCglZ7
KlLfYfx/8O1qbBq4lOw9kUnsRMlZrcsU/VHutviSw4vjVz8ZYipoF0Uyq224In8W
7b3tzMXWg8XqOErncW4zM/ys1e6TM0oWO/ZrMUsDRSdRhHu1+IbPSlMjJE/M7/63
Y3xxFNkgnTS4XUeEYdu4cgz9MVra9UJWJNx2FE6mDnnjt9ROOUa62cUI4WzU97S8
NhH8F+1diACw3t3ufinUzq74X/PqbsjWGSCikzw7syRlLr1JfJxLQp1dj9/QsbOS
Qgp13Q7rixSJVRHfioEQYG/pdQrpcnDcAm4xH2WA3PYGdqddgO4ZWSW2zmd5s+XI
gwgo20+Rh7StsbD4+jq9pRVyFyvnTmFYnY/+4+YIWujAHArB1aZI5WKQSHioVpVz
a5p3dPJRzFVA9ktnOplIPLOjE3jZVOAN9fVuWZ/Pch4hJCjx7OgwuBPLKOrbZtpw
IHZKfVO777LRS+kBAuKfarAaJT4xd37LsIcdcVfkF92/3I7zKHL1AouoPdLKMQZG
CND5QHsN5qpHghfarBLwHkgg6cNYZRRT6OrE0EiyFoFG3Vc/0LIXskP3bFMQba72
3ppkXJcEdMJJ6TObVmSKLfIGA9dwkU5k+0VdLLfJNgYKwLDDm8MNCXTr7PMl59iG
MagWO5hsUK/x/rDAywi/AxelKWY2I+beTmJvC2S5hwozZBN2nHalnDT6tuxWCUfG
2QAq7VYwQgzXYl2tmu47RVQt44dGBGslgt0EAGavLakrnXCDwM1bE8ACXaFREGTX
LjHGavt1DEIBBLt3dP+rysdC4vY77lIY5kd8h9XcP57u+gb+9rLcTwTJ5FSBvlKF
6RH/NGUNFLwrhJQMbaKPeBVQcbSuuLKxCCK6rebzd8nSo9elhpz9Lny+CHh0mFFk
1AdGdr43oc66L/rlN0i/TzkfRNgRvkrmF1/uJJRrC1VHrT3xWrmounZPlP6/lwqu
o0KPefJ+B0jZ4LBJwsE4gvyjvtOm5aiUt2eTbEoSMNpzvVC/PU+5gNkAKluhQ8CU
NtHgmpJF+pOuLszhODhlQi07XuDjE+6MPzPOxcobNsp6EG0dUDrud/n/AGiF9iO9
RAbUmaFIyNvYMN5dU7sg/3S0BaqrXwR3PjH1iGF3EZDmw9iI79SR7c9q9gukrA+h
QDoBv7OnXU2BkJGNnJUp2rU72RsJSwylfyOcv3io/FEd+FL7m+O3Bmi7aI76IU0a
v6nI7i3TvmHY9DNWvIvFUjybZNsBspn4rqVbtVKG9g7/oQ1k8KD31QApGHNY8DLF
+kY0UaG3FSBZIDh2sQouRHUAsyJ8C3V08HLxO3yfa5a5ioEPtApAO3EcV3gYYcSm
A3ot+tznl2QPmhgbqQupjlDD4NPAXhokwMtXGTBgeGDvOFRWVVPkdkw2gCiXKkPu
5iNM//inlf/hfHvlGAzLlHsLqTMisvbiJMFKK++/JaK3qgDfzIbH7j8OQk2s8NLi
2uILYK/iov/byCOQ+u0F8g5W6Iq+vYCMkx2ZlYJhrFPs1nn8324sLc00abV3HlP2
QTGXWGZQIAaxNm+OLSWzHMF1df6M/Qik/1agifeOHC/28VLB8itqsxuQceD0DuLA
yQbvmHyjgcIgVTUYCqLplCWd0Ws47aJepHg3CtVQBNyNmUtdi99/IjTXgRNwr1U5
YVXDXm1IWLNC0wNd9Tkyf2kWvOBwEJXVGbFfTyaiZ8rqP4gf1xylrcuUKomu80QF
irrNTraPKg56zZFnlBBv9xBUT/7ScADLhjDdAKJ1bgN/QjCzulmqZRImORnBDoJf
Y8qn8MNlT+RtaXWljHsySBdtcVyaxfMiBbXWGga4dI87vekp19zclU5O9mpV/m3K
jQLSkNiaBqRkDpKX9D1anusRIxC3IckQJlAcnSL5eH8yOnLY4y3HkGb/IPnF8qj6
MwB1f5mV1mROd0dlLsHJmuZwGCEC0gLCGgAcOvoq2UPEzm7boyjvoYGEpqkV2r7Q
/kGHmYvCHHDrotcIh0HmRNDwI63BGPp3mToHJ/j4wVc1qVtYKJAwfkpp6DA9hRD+
s89X3XsM2kXVZJvc+91C2qDbuZHxXKcZbRloCK/IoyPOj6EO6dVHDo/uHMQwzbrt
/kwoNWixafcz5rBkn4DUx19seYnrLTfenKqOCL5Ue9otHU1bEdfavpbBNnuB/T4D
DFdrLk+/w996HmoV8Nr0ayXVX4HzY9MJo3BgpXRkj3y1rimxnOYyPnAWEuE6+ZHU
FtXvVs+SHo4Byk4tbCgmNcxknPxktt1XK9328+TDIx3RcxKRVJ6g+pkNWaw9D6Gz
ipK7v5Z1SZBFrB2IpAxlQ1wsXWqOirqfsbikQAwv/rjv4CGp8fhGZLbwjFeHEWsa
kHr0ykHXetw1c4Ho/fVfc2xIMMmLJZ27ZhLJ4bSC6W2ZSSPupgCMRP3YBx9/UrxK
nS9rfHtKR0DSjT8F+AKSzmw1wMOmAz73VtWdcHzhxS5UtrptXh6PBc9vji+iqIzL
om8jhzvQ809iGLe+ASZg2tcXq0Uu5s76Oqn0XH48nCwHX1QLV3MLdGgG+uk6cpVH
NsjuDyBXEYv4LVuYCmv0dqA9uNWt6SmyeCK1OFEiN8BzveJEuKnHa/I4J1Cnrw1o
FQdOFa38h9Di9X0oOcnhUzvLNZl9wg2f2wkPdUB86HKGWDdcQBZUbc9corkFYMae
YjiZ0kHZA394czlvrwMGJvYlqMGDei+1Hv54K5f7cb+GloCE+uimbUZaASEMmW6f
qRvYclY7aXCzNoShgX2NmqjNSvoMxwF+hWzuvZCmAjescH+tMbI5bDEQyi2Ks0Mt
t8ujuR538gkW6L+p9S/4tNr8Jr9YcLGHH+sZEAz6kw9KLpbnb8o/JFXc9VEw355u
NebksWLeKydtOED/KQkJagcTAIQDGe2kArkSFg5KobFDhozQzyZ8wenfu+2EgkRb
LFhOaWlS4ygjkCbwm7vOcDnjOristDnvqxN2ytXn5ItR1Yx7V34nNqoTvOUjq7m/
s4zd+QQ9Oqp1tEyU2DhwgDd5iMmjOB/UpTmFiB/ieCA8Ls4HjbqPsxzHK7FDMyuP
/rOmuU/wn69YyEaqPRd1G+8W3CPKybIkzwBs4cDNzNsrTYOBFnNNu+XBRwSbKreI
MfwcHaJZGfN0UW5551HoFd5JeArsT3mF45MIoytjYsci5KISSOme3ZMfBmEiLGlY
SoX+GqmpC653DUR3c1nQf+gd5/3+ShBGv3YVK5XiUNtYPXH5odQUgiqByUtx7iXM
eX1U7QgWH3SNk9hjQuXCmrUH/TLHEyAY47LetBapxVGXuron5/ZlrjlUrHzbTZSu
IEsE6C5j4W0kWOe7u1Nf9JWel+m7lxSaOyzxs2aTIuwj/AnO3O7QDzdnFnvUvKIV
C2y3lboXtJh7W9y4BTiEXU098MEx+Kb0tIPRpwYz2TF5R6jmtbQMetXFBR3YeEOg
3bWOaeSvoCwumBkqI6ZwmX9ff0qKhsyqz44Zt2NWwKATUDF7J/KTKOOL12kvFVWH
NwfUtlkMX2wZZrvbC2iXIPHYSt2WzULzclBQIyFbpRgaBkK+amIDRFu6JjAvEv5A
i3s8fN0glEoL7MLel1FxlfSYGrKFjKcW2RlVkplE2VFfGeVpkYqSycV3XC3I47JA
Rwxxt1RdobjY4jVjteTN8BPfxHs4jVRds+e7RpHHpyc54n1JRUmgf2J9lxyEwnEa
UPg7rNviyPCyueosp6sLLWLI29fSmWxDR8DL+0sSbhl/dXDrCXjOR/DH8kKFhqCR
a9oaZyt2NJql/A3V9ENQNCdLWjMNiqwTPINFqnEQujQE/aq3A4swz+W72l5wjRmt
PGiBkCVQbEp7NlZep6lA4gX9bdxDnp29/5n73g/UnETTZ/GVr16EAmAS44WA1zKJ
05Ndx+jwYJffKjQoHvz5Phj31PhAzOfPU2BjzQorbFAgRNNfvezgMvR10feoEfFB
waz7Lhr5R4s06gigUrPCk4kYlKcV2aFwLPcOHoe35M8ak+Xj7Pa5aipgWxhtxYtn
XoYeZazcPRFHHoCAERrAMW75tsTduf9qUFzCl1rNjHaTqHy9bmKOW+zDIst5gAfn
HCTunr8Dg8919rMtL9Qjxi3wYKfzrBQxNscReWj9vA8ya36ZupwuTSMMKY65Vnss
2DTCwhFb8sn2X4wq2AXo2qLmRZSs2IsaFZdQCgMqxYsD1Cx6MiALUkT81sG8PfPX
gHJKps9timklJpILCIdJwtwqiUNEcPKIQrQrBLGdVDMoK254vtojQ28nhnkcJFxG
H8Dr4ZFz7lA602ufyyrbIwa4+RySGlAkqgkSzWrMdLUHsW7L3Rd+kD9v13hhs65/
mALl42AzlTX8jTVlQ1hGgYxoc98J4bIVBR/4t73EZUpyFrfK6dNpoZidKzxhMaVO
Wf9ySfDVsRDk7C/sFB+C5UNb5pa5m3Yy/PWWDKgv+SydGmzigxB0WKhGT7D3JL0a
Yoiex45BEx7nooStRN6SJHTYccuFAphitKZb2PBagt+JGqptSd+gsySe5zE++l24
hwR8cz7GH2Q01RRFQsWZB4WgfDnY2oaNn8yE6lgw2P285McGV9uCKDB2BT4OJfsq
BMcLvEAASYCKyvA+Xu+0bRUOvBwFh/2CRr5Xps8eHwbXXa3IRX20MwfMjMSoUr4X
pcUiMXpg1DFQuy91BxHddO7CgdpNG+EnC5I4u9ygvTjrQa6cmu8ep0jJKoBZk8do
69erK02LucSvi8tiVsxqp670c/BAr/XYMqqyfSwKzfJe90I6nyI31BaM3BXf2PgV
wfLY0SIsCT2VCNEZkD8q/C7HlyLYI1L6M0vSEG8t3GI0fPSLwo6mBP2GZYnwlRo4
oBILbIZlsw4ILjbikLVcEFJElwnjVAds8wJXnCGoc03gm6e6tJ0UYuCEJdyXbnTg
bvSRVNeo3gMt+IGm+yC9O39a7jCf8ibsWBKzMDW8tKd0h7NBXTP4w0+lKBg33HD2
OV7PFaZRg1cXizIZYW7Qvpy84ug2xOBMQFRHrwBMQstZOzyG9swG0UmA4+P5xxmG
j3VoDQhVrLvQvKsq/UcUTunvKlMEyUDQqTIC3JtWo4DWFYzWMkTEx1SNCF19aEpT
Xebszd/yhxR01JXLyPOfJfyx1TSQuYwU2GsNjBpJ4Xvx9V+solkJ+pq+HrN1f0b3
8IDzRhHaFdceA0a7t3divM47Q1Roqmf8360w2xyENnyxzh1+s+zzpXudfmJHCaqE
7Hk9O9AZ9tGKy/kkHwYn3igtKS6Aq0QQVKfUtgFu9Jx+sQ800xJrwGSyuaaivQhb
ZmH/f0l4OAYez3NhjD/qEYjACNFrDhiKDfMtWxc4RIjmuECaB19CL6LU7TSU+nc/
8Qp0zGTDqL7b6cIGbBvKSHNzzt96E9J3KsbYEHgnFH0FLwKPpesjgw/WduHL2LOl
d/No1eGwrfndwbtz7kYT/H9c+ivUnO/EvgS968MRnOq3bq/1JAQsLHdvQi3Egcw/
sb7B+I0rl05/QSKPzrYKBL4ii0CGP505kco/dcvCZ9GWs5L0QUx2UZSSko2FQdyP
UWjxiCADv7KYq2d9vOaQBzj2lWx2761qTGnB8ewPSnlEm4GSMnQtE1tUjXyag9Kl
7O4W7kiW3MDf36/IWWvh4eC9C7CxsG4E5RQzwrckys4Hl+Vo6cFR4Gq8xkXEUfGe
7cN6zL6yZsxjIrxatzh552wAOXtTa+6RAcVzTmvelD3s4EeHLnj2lZDIpbR+pWrx
4ncVTlsiju5KI1AxX3w0kg3uIeegBW4RUxGLXLdPFsWK1igep957fSYlNf+vdAOH
OTVUyF1M9hOSlgqnnYGT0R1ASV8so//6eqaToJqUL7OSpfIabWfbjmG6bYbh98v1
eUa2lBIeOQEWcBNP9heOsrw7UUZXJs5MGS0T8yzp14ENCv4GfrhBs+hjxpdqOq2q
ww0N9r/ONRrAWV8saOLK9Lpe1kFHuzD05Rlc9AoqhJ+OAH7mjG7GopZZ8n+tHn9L
UQg0hJitEIxqhrXBrlCzzHr3ROPDpKDgSLvyj7oR+om+BsnmFkGTfI0iyaURsoq8
HxHItNRmHZQJ9lZuiJcN0bNi/Rw+em/kWmqtVcsKaWA7Biov9qbPfvlk7MkKx/yM
HLPfJo/z5DDOg2XNDjd8LQif5zeG3rH2PBs5k+HNzQ0VRJDGLH0UAlwA6mU4tZFK
pSXm1t2QTI4zXaDAbYwG0n+s6DlOz6NjwTCrvCTftdZ8YvKaDEc/Bo6v8QF6y730
vSBdJdGMHXiN3Tdq+nK11YrIQvXcF99rxmsAQY2m2HjChu/K0/PoU8ZCVFkx806Y
iAGP6xF97Y6ZMBB57rlRupih8wpEamKu75XdewvfF6TlV6fY+kSKCFOLN9npbOdV
wukXvNbXnRyUe9TqzUAtoBAA84CkMoPcI57CTp/Y6c15SKPUZdAwAiPfk1Y7ycDs
BjQcNuWtep8KR68zLgRh7MdoGMdIgVs8T5FGFWLgHIsLrR4k4Awq7l6gYksGhxUL
2j7ssX5aj7cwOxcb3F4OEJi7qZt2RguKQF5WHN59azWOMX2g7qdVlZUlq98oHLzu
uVpk0oG1PYMLumZxnjWPKnhivIMPvki2b+2oVMOmOb3p4l8IowJMxtjfbDGJtSGb
4ZLVbppTXzq0iKgXSzk+DaPHor/cah/QdDnREy9SVdAb9InJUu9HwtHkpKlMFGAu
9unbY6+5I0terDFMM86MQDkEieaHozaf3ZqsXSmLgO/fyyLRouHUZsT/REQuHsta
S3bST9kzCBa+QCXAtEBl/iTkkreZ9CiyOGESdI/p+FipzU/ZaLUPvP5XWuuaJh6u
VQ9ihnDA20+SitKDcSMO3ise2PPZDRR8m2McbWEtord4cDGvVcKy8nYOEFsp+HkT
xqdW7qDfaig1m8bc7CEgUjoqaC21DEf6hWC3Dz4RhCkx9SFWUcUM0J9Y4rTNiLWq
o+VOzxGgWMx/JQA7eo9fT2gxup+NSeGBKWVcxx40tU2HerrR5QGLDz/3po3mcMyF
vETV+K/IWrS2m40AuYyp90ztfx0WhbNJiRifm0ZlDcBXboLfp9KnrhLWWc2SS55n
+U5IeLcgNUWAAuaIlkg/aeF+kej+DtGxAwkhu/1ULWd/TRTZsn3sHMV1mh1VpaUV
eOKiZgNvlHSdV5fT3RKAIeogciewd75Q/6dz8ktC/auHAHZHehfbIyYoeA14bQ9k
sU5YD8LwuEqdmjRshmcPJYRUotTvz28ftaNarv8Nmkv8sb/QhPSp7u50vNBTh/aW
L1fEB2HVbUaKSzLtjvQMk1QkVkEB7UG737rGAdeP1/DkAXOZuiNTIMkvd2NwEaSV
OYEr+vHfngg6Irel7eKN04yMGqRVaUdqbuhRFdLTTz91a+zDqiw8Ramoe9DuLpBo
/6Q3YbWSeVPAMP7xodd/+xh+OCyIJCAzRNAcmY2BEAIioTo5gOk6m6qNlmwEZVLK
oKBECYM8apv8PF8bKkrsAEHZ+KWhm7s0m1iLqGc3qPVOlokRLIKodY69IFkGWlV3
KS+0EaMOaDW3/aLUofIOR2ir4YzhUQr5csWEePghBjgyDWBxzrRUnRIpeKLc8zk6
FAGPj4Cz8u4jV6qhr7Rk1i+YcYfs+yXURfV2WwY92IsxqUYmOFErfZo7fP8VPGVh
WtdIbFiNsy0OxefU7rwdtQDTIPriZasxd7HeYpgicRMrDaSrFw5ruYV4/iw0YeO6
hMjuqUEBYBURZSvnwVnjVZgNL7OpJ8cIqqfkPYEBJ2+9fa/tSwWhlRwH+mp9ssqu
d1bXoMPyVmj+hx2NEGEIJE91sd74NjbVoFiZ3u5ggJlcPS7BRuwE1ucx1NJdYScw
q28e1Dzuf6bcrntwzyqbl7a7OT/e2Ft89wefpbZ/mys2Q8ySsv7uiIUPEWRU2gsi
A2K94BBj1e7+A+6sbkgURLZiDpbCGeeYDl7J9+LdXhLLcKybfd/hjPXiOQNdRygJ
JTFGPA+AxcMIR4xmIWmxMLGcdpIWrJcoZN0RzgUwM9b1d1Jh3HiWyjkPQSosK0i7
LRvGLInqw1gnUslpc8cCC2Smo/PWCa40Jc8pcg8t/IkhpZycDnXkuzRSUhqx0lEi
Z4lVpLhtahVhY8GmoNF3GRi40I5r0zOHQgGSuTN95tCPbSEcjMLBZgeWSJ4XLOmu
6bhCXVuOcsz67XZc/gJ73ZDNZOpIHKHLkb7vBH+KpVQmcXvd3ayETB2NKfhxcook
VbdsDogen89bQsQiJISXifXGz3/BjN5/dfIzgyOBogyns14sTNKtN5YahwBBx6tR
F8rMpOfpLbvYS9twpz6NF7ZLjgfNA2/gX5WVhwiCJmy3NezZaFhe2TosU13LXxIJ
zT7B0PgoZojCApDETrMgKyyW649s1G8+gJsdc4NArVbNptf9vXnClUWw0yNnqaP6
WbJ423Fg7rgrMe7IcGOef7tdMib641Rre1sVbShPOcWd46AxLNhvsDqxrDEeivuN
ICCauh7NgD+48vlzdRTABOWGqG5JoZXf1EEox4fWwx/PRzvL8BUD3w6V8B/tXvhn
E7II96z4A3qZsg5QnyDpri6fCfETFqU10XagFr0fr1gcSHYQKheqb13wAtMcvxTQ
Vof4JMIL5lvOTEbqNdnImdyghj52qGZV76ZrKtezP1qxrTSLP2JjhO8nw+bQ9Ygz
7KDOfQQ5Wm2jE2dHrtHSo1UiiXqhjRP8nDc4IkOA3B064Mtwf0xr6XDUQ2uWlsI9
n7zGf+q7k/1ggE/DoFwWucR1uQqNL6QYNOrKLIWgHK5lw8hx+dzx0/SHKs05apmo
R+POmzXzMQ/db4ymI9pt3QR4UanFEg+6VghGLJsk82k23X6lFHAivYyoZrM+X2KK
0LNHzhxcPhin9U+81cxRHIMjhoh3knCnXpZy2s2sFa4OFe1vXQFkPuGiAHkGE6eQ
fitAtWwjgReGSL+h2sctcNjNdkMKSAgzIWjvdgm4Ur26rwSIE6tAkBBHzz0yjtpD
oAiBTc+Qul1Rs7WKinrcLAsRjvbYe4JzpJQ7Vjb+oGqsgxLhQzwWG4fEYofXhjDq
dlJDpcnCkWvEAio0yEPiCBWsO8eolbTkV2Mckk4zqACSMwyu0UmLy0d14C1mOUgu
yW6dop4Edf1WJkGqTO8NaQgJ9t7gC1IQawap63ermagU4LQqWP6SydI1kinFnOuM
Q65Ecre9rhX1ovmlGmSpFfx6+4/q33tPTd3WckW27/mpQG2pMiUFJdZHwxT05mwK
GtKFIesPEvyU61O5hevCH0BHu2VyI2/9p7g5GRjYbxriQJjM11/LJBF73c5uwBuY
NH8jdU0C24q5tvDOOrE6g8X7+UQkYHSQeOI/M3mo31Nv2TTuipULz/yo6kT3bYWf
Jw0DTA3SubqRG5tUnxnW3vDIJRwNx9Jml9uZ8IFDgApVyxkYZ6YqX91MPN+uqzHX
jHmU1P+dIAtUiFMn3RGs+Jo+Co9fZW2OxAi8NgsR1aKUomcXHgokFOudJb4bXes3
jrjxu48gs4KfOE4YgLKjM5P/sJuWvJScw1va68zWa/kz16+EBDiiRMLOWlZp9hNH
SrQBKBBXvYiG8G1ijtb5LSjKxrtOkwEjv8CsEpBjKcahppIVYTOINGS9eVGvfiKB
2bmtdF95Dv2ikA1nmzLfinlvqM4np58IQ2cg2vbRTFMTjWhoitR2wiRatwV12Bur
2VvoIhMjfWcTvBxDY/lxTMlybfU5dzT7+vZQDbo0bw/t9XGRXJRsbvePqV4KiEUQ
vn7pbV2MJMZShk8SSDaovh0LR5B9eb0DT4jY0SM+xukKsnp6Kck12BOh0vU6msOV
RiixLUJYjGz3rpy7YV6PGRXnYW4hKjixwv78gm6gO6HedGGX/8+nLlNuq6ND2/fS
a0rFk4pIXusNUMQHYIIYz3nNUFIy2m6o/Nqoz3LQGcDKRPKbk9smTpgaoWUML41Z
ifWPSnasY5SZm8u2wte6CyihKJzudOTxdnYLGKBaXeMz2lxX3bHbft5jsnXbnD/y
YDt6ttBZDzYas7yrFSSZtrTZleLdUPzeaY8VoIwNrhRv7/ijOc2y73coJz9jrk2D
F62vYBCcMhaVt5o6GsPTfApoOA/kPcw1TJgv6tPQU3OclqqOlZKUyhhQ8oVRkWKN
XZMZNhd/a4ssZ00xPTtz1M/1mdXlx84qwqNifeVHgU5katCL5Xwa6FVU122VhF6A
xsuI1CqIsLGViyaFANfHw4VKx09hNK3fYQPB1aHo0pxS5NNCopEkASM8itDIoN59
Q5xRGod+HPJQwDuUh94x/aHLiUZZaQs2DXHVGKgfNSNAd1kPg3oVrHZjCtj+wERh
MvtBJwJk2Woxtat0LleGFZBX92ZWFasjWI3hgT5km1SQEzlaX0uwRVclRrM4gqsD
IoF1H0tZ/JFlMmTXeTLuuKIq5SFqRPfxH5Y6wJp4mt4lAlry5Dx70ohSJQwBxelE
dykAAMIj1uYs74mFCtRQmY9Sgga34UaQhGoJ6kZ25XahM7pyN0vDDnnLVOdJZ5ya
u1ujQ7h5j5vuMpWWiah4KSF6WstzIwzh6Ck1lsjwN9vI3yuiIsiAhL+1rPxWZEBe
OmPIMKjo0xiiLBwiDJTuc5Aab+bGVxoq/xv6ZxeOwhIGmrrZvQD9xOy0i5Ow/uuO
Ni+UYHRe7AQC3QJV0Qs1agX2ElpZQXMksH4BH0lyKz86z2EEkc70Zqr2btC0yQ6S
MI9WBZ9E8vJ+ZmMpfS8HCaCa6ShGFT0bOzF9wSvA8u/u08u4prjwO6wbeLr2npp8
eccvVo5EQ+PnWPdVvnkmGdx/yMRVFSkEn+e+dfDc+p5Lz7AEc76/O9MnxU0OyC6N
Uzxg9TSlQ8oi+g2tC2VjDAf/L93LDueB4B4qbC4FoBCZ9B73B8B0Fj03LPrz+nj4
FQs40lmyzVjaFoHkMS8NspOCK23OdUkI0uzDlbBpshOoAbWtYjcMKVekivnaIIf0
J2xp9dSHex9f80WZyP+02uMYqr/FZ7D/mtjA8r0ea8Yfp1daHW+EwkRXYPDK9otc
W5Jjm1jwtoLr64z+5bGCF1hOXCNufkKBPJmFM7g34mzd7hUykoGxX+KR+4glSRcy
S6Mz1l3AZgOjqVyJ2f+pSmT5STkLubs/FMPJs6NEj7t8xS3GtfEhvSt8bdp8HbQB
GCi1tRnLMUDb3pwluuragXlh5YNZ0VVL7qXZwO5YMvQgE41xcUqt8Hq+O63kf/lV
x0YdzXkHevRnTGFz1EzhHmUwF+pgNxTmktJJwd8IYYn3qz8u3opQgp73Kn/noLZD
JOmX4l5rAgroPvmVrjX/y9lD2ngasLwzeRkZXKJGjb4vZil4VjGk154WWtbyTePE
p/gJ5OLJzu//qWPT6HyKLJBdLJy8bnXMRc8m2aKzWe2eEpkcVPzXotMOkobx1Byb
7D/bSYDi0NKjQKBf7gQj733YoTfRp691bWSwfbzcbBtljepQ/BeSLK7lW1UsiTji
ikLdaMBdFiq6s4G4xAKCSIcrA11CWxH5dfAeESdTmtoNdf6a20j6GbrF6Pe2Kurs
etjZOh3aZNRiQ/7SXBJd6OY4WlmdLiyzo2ceRUXi4LxDm/IQvdfuz0aJjU0TSIJ8
+Ct2TfIuIQ2HVkApl/XWoUep0emJtV7P6GEWrbiQaeXyQS/BXt5xc3DEAYodcTv5
WNcyuzHpwURuqWyrMCGzLHba8xL0MgLuUpIT7poH5c8ajeuSFjMblusNFDCjSsfB
QvPtzQMcG3Bwta3WXQTLsnadct9zNg3t6iKZXU0wT85T4n/07KTSJmMoMpC+guGx
xodGlNdILv8f3HQ2H4GwD+F4Bklqb0ULb+zo68tSU5qHYGWdjN8Txmc5pJ5GuCA6
oAOsu/O8M2+OnNcrWVfR3VOKOK/X5oBdlBPVD8ekM0k0v2xgO5VZds+7cIFUVhRL
FN+kWfEZcV84MSi9A3fXVQsEchJP4EnXQdkWjMRSlbvhSLs/b0oKyzsv7xpIowu8
aFosGDS+aHp+XZJ31LQE4/E25S3dXx8uQXiJ2BTDN7n5x8E73qnGx2HpU5WSjYm6
/zJuCPGRv+8QLalmEKC7Lqv1DQCUB+Z5DMshhDSiSwrL1Zipx2vs7dDsj2X3su4i
vGbdtXA2AoODQf0ok8eBUBE8Itg1Jjw1BoXj3NVAyis9x91AIX/sht5fglRiIQaq
2xCdZjAB/qdtCwILuBfV5hkXZzf2heeFyCSYfH70Qg9jGLG2DDsrABVfJTLLKflx
+YBtZsvYKI3hDeofs27KlBxEAhXh7fTFJvPUNUUQQ2PRIEkFivo/ORghySau1dtv
oxOhnHsbBEm22QCLb5sq3homwTrQsDetVrwl44wx2ht1N4d2ypJXi7mjqaD1Wkwj
tCZl6FYeUb2UjDF1HKEUAoSZIvOeEdezSwJLNdDO1X99iMzJH38OtnZvbnEhervm
BzIChWiEO7+aRBjy43jE1GulY+NYC3hzKikNxgbm9LIBlafqiFKomBlvoKBFwHZb
wtNnR5McUQ8XMlUi7XiqgMFQFuKQM8HoEkW1IEf1/pSp20czw++4EUgcL9GcqDrT
bI4CKhHHVV0wtKetNs48dyJbT6W3mCkpcG/yW3Hgl7ma9mbWJnpLU/GwwaUqrniS
z1UzTBkBbUxzoknr/4Zpac2z15ZAFLCNyMKP+MsX3lvSNaSKgD24SqVInIBKppGE
lQXbCQOeN8Q+uqN1vKgw4UDcLAUxHxHpG5GZ3hgLTBmvEvrPsc7XNL7UCVeM9qIt
gQXVC9efD9jD4tU5GHK6MtPsuNpf/cJ0zP6MTCgkRGKUETxJV95Fe7vS8tUwHzsA
yDLRWCYuuzYLKS5cmvXqkmkPKWTOO8yu2dc2RHxZ1uM5VD8mZ30y2ks/mWJry7GV
58iw4plrtSxbysx1cftYfctcAZoEI2kQW5wFz1dSHwVu2VjP7s3CZ+PlsdRBCMJo
M8h7GvMQ8ALeSM3x/RPcxnG5ELGsrrxAEkG26mtxQuAuGwmLWAd7Dr8uDNRup5oH
kLGhAb/Ygx7kuKlBU1vDWdbZXlDZ2IMKFjGbKeZD7SyjlFlHKQTeEYbPQ9d5g5Zv
638Ve34AVXPB0NuMCCEosUM7sWrukXyTFQ4RcKpXMOtMMPK7VtQWcP4hCz1+nngd
YTvlntu6Gkm7GXM8/FOHEQjT8j75UvXBrjKKd3NePG0rso4D276PwA1IzMnIeUmN
4Z1zdUfPSBPwiuNpSMYEcg0koU7IgedGxQx/1jqYc59dFqz4+2BC4zIamyNevcjs
9cGBgznoJmrvePm8UymlCoxnN4aHtSTYoUK1tuB/MhXURHxXEDvgGymBksZI0+gW
8BUmz0lh19GqgBswA1thnY47ayW0IurmoT+XiAsydKYJzrJy0N+UCtmNshZ8i3oc
VoS78iFogdwNtjTaD8hSsLfZvfWd4+Vfe6YzlRrhViF4yLYId8JAIFFwf0VFDHfw
WuTQ3tfmZWWiJL7KQ1CG+NQ5EHtQR9/6bD2YtCscTZIvTm2PYKW+t1Wd7o3NIIzf
Ar/6evfaWYv8I5/duW7Xgx7yhEFJYpVEF+ZXTggxtDwpTYJggikzqf0jrRJEyg1a
xtG7u1jggHdLMjH0f+5ye3M7ArsF4wYktYkAoiBkEbiJv6DAqp9H8+dPWkxdrNgI
EZ4BM6mbc7BfgD8qjHM3cQC2/lW0G0PcOIpVM3HCYp4KOY2u7OdMipLXEIN45+gY
LZ5xsXxhCH8wEjuSsnO86AaXDjdBZ2Tugd1ZfmrVuUhD3MSAKZwZzkDFyJa2C5XK
kvx/dnbH1ij1aQJGhVkQLfWaoJSt6JACLNaiNo2G0hkqW0M5kU/3iX/lPLPzThaa
8zcBtQn00Ml1jKAoKGnWFj86v7Sq0huelg6og4IA5CFDf4lN13dEjlxg3FuVoznT
dXs82cCc2zpHSLOoKtfOVqc8ljgWGWA0IKB1KH4p16GJTBsiqKfKV49Ol9l4pAPt
/GqZAGcnGSqHfbjfi0tuP676BHRIxOcSshd7jW/YDU54XOMWgCqLCWEkA3f7dTpj
WGpQLp2i3tkSYee0iTRxCjsyHLQVgFPiG7WcFoAdMalUK51IAsG7PlDeM88LkhWy
rmpbd/6rdJLHeE1VrB2/idLlVXfW21PW3KztaJTStdFkNA5sZAWvJL65j8KFs/2B
Ku5NxfgKOEgT0ykaZ1/+HZp/F74TnKf/xcu6//fy8lYw5pYzWP9pjgZe2Yvo9Ecy
a87mZB4ZYdwX6SMCyT8NZMSFAsHYlAwskSSlfE2wEQwKSM/KiLclmkQcQiGTSFUC
wEpt8Ofe/AwN2dI56IQi7fZYLSjvKdjH6YH7E0jSvxK4VyXA10Ti4pLtmMoWUQdh
Z4Kh/epxfZw8tir8UEOLCbOkJVGYkggVkBTAROUt0LsqkrF+V6SKabdtPE5T4ibg
gr3Cp9A5Nld4Opu6SLe8zwRQS/QOzo+9vjd/MPCveNkKNFDM8CKtzbuMwNqKGe+8
8G2TK9XijNa9e9HbgtbrhDoS5trlvojBF0nHOIhYBBhdUiis+/NP2Sh+1xvFt7dM
Bl7nf5nyqYygfXF0f2iAVCawevW3MbzTPhLeF020K90rLTOUk0bVRQuvScXvrTAc
F6DHsitnybyXgikgP2z821c9HW4zPTmPiX4SInqg1VC/bSljzhBa9zNCkKCf1QCq
dnGWyinvHTXfN58+ePPmBSE3zpcNOXSPMARMLcU91XOtpbR4qLPxL1+bdrdmbncW
1CigKCmfEGc0d0HEwwl8We+kmVtIVSUYFUf8+rTaG+KlbrsH3V9KswbNr6gi+KB4
0EHVdZCyq/Ir86MtIt58pKU/cWZfqOuyYplpDjMuPCsEvNNGfojK/YKByCCXEGXo
vhHGmeuxNpZLjIaAMZB6IORAarDPOK0OMn7mQE3WcgdrwiztWbv8E0A6MeMg/DP1
Q+bz1Ew9tzfORk8utoiEsgzq1q3KzAZ4Lj3iZJc13IoXUFQt1mD/Gd9OZ6/Ndy0z
qUzZsA50KX+vqFYbX1NiksqTmsUfW3DB9I4zDYU93LPDP1P6lZf8eM1U/pD5+xtF
fxP9XqxrN25o20K0TyFYLAzc0v3M3iSZ0+agyD1mQZkazO2+TQgKVTTyFC4uqbpD
QmW/jUX78lWgV1OTiW3+ep+yo9D1r0S01esjtgzgxWHTjVhbp5TL9KwqDfXRY5dW
t5rndRNlTUU59rGue2fuMOcXbEWjgrCm1GV8juh6NlQy6Kid0xBbJ95JNF3HjtUG
hjJZNPE6yGMxL8pr0MsUjs5+B7Q3vdLIyzd6Tw4a8zXc7g+YC7BMjzqN8n44NE0k
VhTr+qcpLjICFyeDiDbxr16LgYa1DA+jWkKtVYa/RMHSVVL27lzYPcKKTCqh8ao+
DxLQtLOL1ByqugxV/epKWCqV//LihshlxAEhaI5Ts4O3exRBXeYT9rlU+QlRWipc
7oUJPMLi7N22Eg6OuPHfcOFx6g/u9fUYCHQhLT2IWE8oX4c0rcrEn2mJcolOcqNm
NP+mSXdPbi5qGbWx1A/uDLyMmHWIKptdSZcqBkFv5TXTjzyGRCxFFbZ8TxpkIZXL
J39pPkQwfR8V8cxpFeWltXb7gxNfdV29SijFj57WOpzBBA1SMGqFSGp569pyZ1Je
C9FOj7V6VjbSYHA1UPLtkkdjmnmBUHP0BOJMrGa05dVjrTyrveezl95Ai4idH2bK
VCfmu8LmlOZ5dn1tvGdDnBS28iWOFJQ8SmgFGBrvnZQvJ7/aHGq3uPzOsIkZVnWh
zsKdusP7nXxP1ltMURmMuEE7nF1OVBuRnh05XXanhNObS/9NvjRJZAWVCrVkgvm+
nNMkOXVBSkEienKPa0j2V8TTxE+7TiajVGGT2cjO5K1wn9VehjEbC6Q6q/SKoJ2F
4UuxO2rGqVyA/PZbXF93wZoBu5ZVOgQKY4bhiiZg0TdkuTgYEjstJd1s/jg9PtPA
zJhknzcv5rR1ffuRDAK05Ct1f6KkuRMTrjhQ1HgedZI3TfXzkhkmW+iKRsF5PeHR
YLJSXYNhUfX4+EZo1AIalS60Y2RmlDjV4MkEA9WcyA2t6VbhH3pBWt7o993iu7MD
84NKSbuQQIJynq4paazdQpPofRiG1hL7/Q+zHWHzLOn2s1z9k/aOBqXn5abTGabG
QwbgpcgOmiaIR8kWhyQsgQPZN/GsfgtwEGMc/j32Hm+6zfTWQb+DRi+wKpZWElW3
AL2nyqVbWPh1IUI/t0dRARm21IPibUuEWRxX22KcQWBScw5I4rpnhvq9e6KJuHuk
9mbDI10FJjNkfUUk5uxNzEsm6xQPMqT82aCYqLAyJuvT7OMWEO4oWR0g+uJpurzU
krBVmMiGdp3+hz0H6UW5tj1EypxfAzfJWmUJcDfUPY2fNXFp91a527W2Q2so3rcx
AyEteSRKiriwqgdIreDn2C7eFw1zfVUyRpvEd3J5d1X70UPBNigCrM0bDA1dfELH
6NPxaKpVq1nh57LVyjYNHK4W9klZYPxMEdxM5Q/qvcTYGVASVYqfasyHlSNUrZp/
yE27PN6EtVxWQ3yeSoS/FFJda/Cahd6S8Pqz9uqNmL+7rWPjjiOXggU8AnQQLCJC
8qeHvNlKIEanpmTEWg/JmLG72xgr05AHoWQ8uzbU8pYqe9GjdeOJ0Idph+rNrPyM
rpYtBMM0fzWzUnUN2AAI5l1QexpcqSrm27NeerBxhuK0CnfRxp01FjlEh2iY6I0T
l/fL3PUr4hoU7A+K64rWKKIPN443fb5hdUdLXcxY5Tcrw42TGHE8j8PJoLKw67Uv
vauBvXIo6d2+szt1zurgC5jtzbK6jnv12eiWDGlM773Jauf3tdngJdv8pHngAwg5
9s24IGbcscCzF9cPCVbEU9ZLsabtrtzRdnFlb1e6u2AD1rpF18kO1Zli/IggS+sV
u5nW0t6lrVW4lEek7h6RJWkab3xyiFeN2oyXdRY2H4cblAbdZP4mJAAqloHg5e0c
+C8pnHKHgWeE8850ZvN9qeb9lWtOQ0vqX4skvx9KclAlrUBNu1K8Sky4uMPGl1/9
fFoaxHX0Xct1i5c23mpf3AnFSaBm02sszz23SETt0fCCO/E1aF6KNZK7UvtdK1mS
+tim7cYPXV4m3EqB1+wNjQkW6NuVbhFNTGzEbSiLUPzH1CFUCAsgqw7EjDzxJUO2
NVJm4bpTF57NFoo1p2Z7jQiIpEUP63uQK829oe/OxEoAuQ0mMkTjWfoJMZvteIMa
ZBO/L9D9Biy32s4aLpZyyyq/ji5X3vVXIgPcF/j0fRa9j64GXrD0bltReD4rxlDD
50U7Xi+QEpaP9Fjs5QTyJ3KBjZ98DbeeTu+CWA5P5Uk9/PuGLvKDPb730qR7+eA9
rUFWU2Jlszx3RJcT3wBWa0sWFbEH/S94ZKt17t1Co6wssfh2kkdJVjO84euqMI6J
vOhRksVkMActzmbT5Luvcbx0/qY4+NzjUiCXi+TzHpfZR32HLQVVmyJjrOwebDNz
JPfIWY4c1MN9r2X+nDK0JBKKP9jVNXrhhnCgqnnehMybH4B3c6yLeIjnbOSknYUt
FhzQ/rKSphaPD4D72+/4sqEXB2z9ksO5GIP5qQWeQGCyPp6WhyzP+Rldu0U5zLTn
CcQZeUg3M1A1FEQwls5urHbxRPqXvkPAUlFY/u0mMsoh4YvKvmLX1kHE6EVDWTYz
NSD/o5HLolSNcy5ewAyCZSgq4a+0XdRAfSdepcspGO/Hy5DlmWptY1xOagbbUapS
6gtXzDqTumuTJHJQvJYVQFhhxkq4Ucd1iSAYxmUc+o1mzsNeCsfnUC2SDeon7+Y6
+J7Six/8Yk7R+5Q45dXTz2RwnJ26hViCOfKXNyKG3peaHIAmJd0wmpY1CncBY4Tb
x+BuTUa8AZaKjwDaNXXaZLPuDmtX69OJluSU26/NfGK3H8PXsx2oxI+r13/jvCbL
DSbnqs0MVdBtF8AzqNEoDvwtCRl3c7PTZ5ZHvXKejUqXzYTPY97uW7jCNf9bCVjM
upyndym6TdlVZoTzT5SFgGa6dOpFqHYlJ+gqyXYxioV3up7BnMmP7l2OoKcldkVT
OzXiEv2NoVYJzErcMxbbchngOmwuSoPepgwEefVIp/65FIYr8VL1uJOLO1vsoMWi
laVtLeMAQvyZxMNoOO2r8RR9KM8PZR+2Fu7vkFxRPZFhLDNR0EX/KC8KjyVel8Ig
5P2S+bKNlIMGJ3mNdL/nDrgkNy8P0+PqvyHWqgPMHzEoGzc6OZUtJ3FJi2ZXT52j
0tLQvRTdSA01fCUCliK0AsIpEe/ign4JO8liC2ei/OXzhLoRoMuJvOeZ3cGsTZkg
ULbY1NfN0dK/sViYBrfaerbDURmMMqEGxwTin7duNnSivFZr7XK6iEr047rs4HhK
zuaYoD+mB4xcs32VpqJgSU56W0nu/vw3oEhetNBkXND+LCPH7Rnv9Qn+5xLMPk0s
LkrLueSgLXvvG7qt/Nsq7JPtN9VCVdVzt9tVAlvY5MJbs6KXli3TKZgP/Zc98rjk
CMIKZzv8zq6AZFJYxsRNJEaQzoBtism6Zi7tBSuhr4bR9y3egJmqcGqRKJoevr31
DUX+0Dmw1QCz6/YWSW5/m5BcS9MlVcd2lyFFJ3L3WROaH8j4oYeVABmjk9WGBsM0
OjNJ02Z4oHyaRuA6pLIC7qW0JFEyChQgAToEXPK2uQHcBU0FwUwGmCm0DWNEvBwa
LTn7IOUFFdPTicsWJYLE46yRaMPPppp2xdfbB6dlrpZsnJV4jyd/Hd7biFENhBmG
byG7kNLASdYkjMVQWE5qF6/iFVT8RynsyVq6W5/bmp1dHEVvXr5IveoyMTCVcUTq
Z6+zZ+NpM4v7LwFxbLS9kKBd2kA8E7GHYY1N7FCaJtPeKXj6X7dK/5tOmNSsUfje
GVAPaDv6+kISOvn5eq+nXz2nszenlnciERoj+4SRAkoATkzYrZH6pooS82bjWyvG
t+rrH6YvZkYHqTAxkKKYMm94uxA9NBVnfp0VccpPJDKMt+uQDbAaXf7Nl1qY0TSZ
d4uy+n0PEUlHklii99ObVnxlrUMEQARMgmvpbDV/zPi9koYHbTKLAwkMkVNuFBvv
0rE9HbJ4SCvp07RPcpeM5T5PZU0YzLrfESX0M2g8q+Urn+2rItWa3TXQkDl6aDd+
HgNl5abYSerC9SLO22g9kSjHakZCjhj0ZCUh8RJO9YU69F+X6MDfXtsZbA3a+V4/
mewAIM+oR/Nax7xuZUQ0AvB/kNg/HfN6mQ4QU5m+YnKUPmHO7RIPhE1kbeTMF1n9
sS6sFcKxLJPQKcL4ZZuzYASbgE0UUKncC/pFPQELuTQhiLfNqFV9ElKuAn3H+KZ7
1fmQLJkwJDLca1C9hB6Z3TBtsh+T91HyufqiuOZkcFH+iifB2vi+lqH1eJH0KrmJ
m/0KRt8gaQlhQ+qMgZR8xKTp5iDcR/s8kQLlsEUOS03S/evhJxXW8DG0dwvH3Tx8
1K81/6+zDsU57KbbdNsAQNGwsKqfip38bM8Z0hFDqNdBZ93WOIwrxd0yuDiJMarH
HhFe52KBbRJF1EAEV0V9G+NozEJwVa/jRlUrqCmfHsiLnvP5WGqTkpLIdvr9I2B0
srXzAA820T7GybhOd+a2BaGMZEm/U/53XN+j3Sy9SdDB8eWdyKcNX07XYDL2K+eA
kaXI2T8BGhWyQKAgskChhhytyquEl04KEZGDpM56e8zPMGw/91v0b88Dt0v5NmKG
wqOfb2qNvWgpnHNRcfe7hXUZD/1CnqxvosqTyh1sd+mQpD2gnXYGPCP3ryI+69sY
yaVgXN5+djBeRvu6i8hyRFw9I2JbvxYqI6AQbNA+XtqlNA5/85MVk1qjV5q6qX+p
ycsv7FqNV/nkBrflOwHF1hmkA3tDQ80+PFu9upL0isrGqqo7BBGG4zBthH2gRoXm
SWN2C5G5HVS0NEACen6r67MD6DPQVkD/KNhLsSfXouS1grtiAsTy+jYwT3avs79X
FxdYGxVv88x0CHrZNwdWqFjV6n11hnYmJprrLWbL3cB1gmvvAJ4/nT7b7+Lfe78S
q3uCV0aw7QV/B0sswkB3QkpXH3XlqLuMh0PCV/0fs0icwRdwmeMCxyMFKdXqXNA3
qC9QRC0UFTIs7AXKXPqtZQ9oGKdNjcFPOuursBTRVZrNhq/UfcyoPPCVr+sUfPle
KnE4CB8TaEJu45rxAh6UWA+oYY6FaBHpAZDVZO/a6nYBLbWdRAzw2Yk4xssIAQnq
KgB+3E7n/maK5A1zPGAhCHX15mOIVzzmdzkRVWhf9qZAP8QzsLUxE7caZlYxC025
pSaaaxPnfzpKLhZ6M3i0dDUFtEGpNSXL9I8K1BlVNaNurd2tjR+nU1n9heTf4A3w
mrG7vxlysjPBzo7a70zsJr+Ic7p6ZCfgGqpsLfWHwUp83pi0/Vf8IidSG/SUETIY
ls4vE9fMs7T5aW9eTrPo7u0aUMyrMrXfVLj9oZXkPeVjFY02O82sR6ibgtYcZnh1
YRlKtk27BCL9KZlj3FPr8oYcvH1oR+wXoKaoatB94nG8EXjRk0ub//CqqeaE97Wm
28rYUxd/iWfjfRKe/J/kyRSn/r4sqxy/I7obqiIyAWfu5Ti/IonQrxem5qmU39QY
y3/LSKhGx49Z3Y16z06OYXHjUVI8d3oI3gz0u7o5MPrHXHcR8KUtNgP2QFG7yBf8
wAZ/Y7DO2K0mZFK0mSBNdWjxEuKuNNqKpeVJ+HZkXlmH++dK3fgB+Tpc3NVUX8la
FOd5Qlgm/YGKGPoeEj1/PqcHIOH+0dDiVmOyr3933U0k9kDwPASgaJeb5dM7HkqU
+PSHGwUuh7dXZGqjGCgcj9LWuPKlZ4iN0k0Axcq5/UPfmvdXvO4jWX0QypigPSbS
Q5oSUG7IBlYr2sJRSf3HFcexF7dvsuSoylis37KmlxkmvTuXV0sknkF44XFASvfy
jjEbxxpj8XAQ8r5fzJ7pDcx9zEViqV4gwEQUmsbc7WHbqUM3fLTA7OF+yasjhLGM
0itNCVthplWkNjU9QtwB0BwobzqMZV3UwaoQ4tieRtY2ct/MVsHlO56rKHecd2Y2
H22C1glsvS5f15UuWiMdgcD3K3aAJ5pEADdWHJ0A1ENKADV/VQOUF/cwdOJen7hl
ZzQoSdIUTwYk5wx9zUXVrQA/ToYJ6yo1NdEu6mGT6y0jtGwp3301HY1WoVBK0/al
80ABzVj48VsHUV3uQWMo73bu0W01rR2DPgaWDOrS/nWHIZ3ZhrXsdXhkt8CdTlkr
dhUjzhEgiEW4QMvGEM4szauucBbmdoP89fADx7lt+kBvhO6AS52/7hZakAK4mVqb
3G+rOgxH2QEpnO0TpSKPpyzZHPgasmLBK7n753knqBWcZTyTHFZKdsTkv8EdGwxd
GaMbNLW4lUBmagnWptX954l8r12EBol85s/BOJ2lbmG6hAOB+J/2i/gGIvAYDEo6
ZO/Gj1sOpAPPPPjFPnrbOQqoexk95TMUfBsgh9MI4/cUrFt2rYVWx3m48MmDp/Sg
Fm1cFC3nG83CPp7i5KaIALj2QjLvp41Nq/cjmI/7HQ5ZvoxhDh9zz62GJYamRLuM
CPq/ZCFdPzgqWBpF+ete4QdIrtdpQjPz4FnR/vQNApesIwtiiJEQiB+EWikLojtt
RXC/G7swAbxTD3P8Ed5f7GskpDykI/ea2yiF0mm9giYbaYCJUGw/HF6RtpZgAJTu
ad24nKW/jvfYl8pgj8H1/SVNj0YaAqnKxjqIhHn2aFmHF8TsrTsqF5FA8emxvucS
m2fEfic9c7DGKXnjXVLQMySNlaptr3dusjyd0+IHA8vLt2p7sUviFvLWrpbXAUIV
LWi+Q1UkzCaslWrSKqNJO9WwBLsOO1mrKyafE+zVtc8w3X+9NlfIcyYxoEdkZ97H
AWIB/8MUjQMchURwXCVOYcYx3VvMYyX5x3eadi83OWrLIBttXqNHX6KU47qqv7+p
/JykrNYLL2EKmqCHZCiQ9mOQWJpDHiLrOEv4QkiZ/T2b89FWDUfDvE+/947UmmaN
fawrVeEwBuE/D3JJzYNex6yNup+tnuhq+CtFPQwo/EdVjuna17IgijWGmNNuxP1Z
oC5xRlgmu4G0nrOYymGmCuPn7GmUcvFjoRcwsFiFXmsmTjh/+uEZgA45jtNGC0oV
snGjKjjHSUuEWeGTEkYISHcAZNssrQAZZRqYKrsbGEvRdHY1d80kkyGdg94DDpDH
e9WzTxK2lSQyOvUKcqi5b4PAQ/cSDT0JIFZRKEz80XLQboISsM4AP8mAgiHcwXB7
deIGFo5jgvk8ywCqwaSTOqVAIImetSFmhVQcKQ5vD8xQ61Ped6VOyUSbANAmu5wC
GXcwNADZk4NYz40Od7PIvRHO7AarC7vE8sOrhZp3gMAFwqW7q8Yydls7/VUyqBnK
s0gYv4wq1l9FtajKEPnGILgZ+QMnt1QxA1xGlaKs2KXc7rjlggmMRvy59cPZ6r7p
fbt7StJJiqpWW2PvTJPon9cxt8PgbntKVx5S84Pq0cHYIAA+ZyTrY5yYBG9Cx59y
hIK+4QFt/CMtf5RMLCth6jL9eQHWtBQy9H0a+fVxm2ltcyKjdg4vx2z2wDUNRXls
yrzCa7e0tdu4obg/CssciTrtmPOpTE/vGFsbYK8IQ4yorqWJb8yxWtOmqx9F4Wwm
9bpxMzzsgYXbbg07gSuGZr0gFXvKKSfzKh0DfsSytlcrOevOgmv3L+1nMfXCH/w7
a0koeuZAVIvdK4mCR3XmMM0irdHfRH/laAewAELG7eR0TcIdSLv5Ac4DjLDRbTIF
9llJDcwoXmxMD8CNGqt0NbFmS846+WnYFymMW/U5gv1rrYWE+wqXeU+JOOPTlK8y
dTC/2froX1BYxgivhqlkgjmgOF3wDaBeTBG5f1fr1pkQ6KqFpk02ir92WbIhxjHK
eWP7pKy4CdVdQZ/o7XqTtJqVUgz+Fg1f9nz18gDFA4Qp0ycByGP8nDqIgeCcTZpC
mTYUMELGAMuOOD5TaTI9jZPj/a6Z1+3aEkD0Gkid6AhFV02F7+U1FdXR1VKDUlxE
PgVmrDm4JEpxHCrPS1tISk2E17ZEu6Crh48wMdr5UwCVAXrjKItTPg/8bEyBOnD7
IQInu+9vjYfNgAh7FmM12yigeDYJEoEYM8BykZ2CqsDx5ZgaDEy3VynB69Mr3m0U
bTKkD33Jg/3xLNJmJJbyhXL7pJus12xrIhycL8gnPLk5O7Tb/0snTokSkCMGKotU
g84a6B+3WHbPLufiGdUAVEZbckAAqsgFjP7QrlNJzxympxSQBxwedZchOP1jNQHY
6l1cshvDCVofylHAFyDbQEvuzW6x1r16gY2OmQm2noRrjzqUeoNjovEC7LlNPNH0
10AM2ceq4dQ9HbYjvDbUrKZLqy6Ji84AdiSX3kFwnwS1q+AAKxY7xbtjUVvzFopn
hMyGmM+GMaGrh3iys9kkLX5mdrDL7mHsfzDg6wtHB4MPCMWHqob79HTInJEm3QBp
sO7fvAICjiBoxagEaETzJTve7sy1UA7xD4jtzWCN3jXjroxdDnEmSGr7t3IXx7pV
IsXHPnOaIiXgh+sXRDegGu+n7y7Aiv39FB6ueOfoCljCCP2dBCTYhgc8hFhByYYr
Zbu/EWSuZQSbuG/yhc953quhsIZzchiPiKDaWLyrkDVvcYIwtGcGHGaOV6a7WliR
DmTwobnnUopp05GdNkeygvA/IOqwjKy3ldp9HcYmmV5v8uhLMIfCD9ch9E4qKRWf
N23PJA/NYaQrUuwlDNJFXS0CI6z+u1z1dK4oiYmCGXaIBFc9k/vTqA6fE8Wyu3qG
+vhrLlwsgaem4A1O50yz6+uTUnpYK7qvSg8rFYdwGKFfz7kXxKqFe/quy2L/w2jN
NBo3dQah/BbR4pcJ8QknEyCrXxRpkG5whRt11JkGqseigHF2aaA/GL7uc2eC3/r7
dWg7RamOrPLGl7nxMeRef1h7mLaxMvp1e4oPs+PTRzvjYVKNXZJfw456UsFMlP0Y
qKuUS3HL0f79bPwvU6/ensWpx13beZcH1ILP5/RszkeckwCjYX4OR1aF5sYdXcqc
+9L24noGrLFFnWPr4N32pR473ZG86J6Nn/f3vjFB2tvYbBOhOLg4UvOZIW1nM4kH
FOiP6iwLhdvhFKXB+IBKJ1uAmNekTSEzGzyxDoTcBnKDPCwcbiJ7Q26davHXOMHw
rKMlvjlpeOU1siPdBb4BMHu1yfmuHbfaycGJCT/rBUCxzTsrneRulP80/dLkDlWt
WnLhX4cotpb905Xxb1FcEuyjf6r1z5PBTgk6UhMyjcw1dIypI6Lh/0sYBeQwkYz8
FQd8HfE2rAu6H+FfWoR8WSOrFlIzSY74iu1NGLpq4dHs721Yrd2xBqbCn9/UrRYP
Dhix9zekB5fmJHc73K6TBy5L6dopti5YsZKsnRHviByh1lyZmV1hzXSB36SrZvPx
1oqkIEIk0tCF/o8N+h+cxCsawhVd5rMySTWchbI4Eptg0ir9D693V/KJnpj50SJ1
JPkSv9PuEO4ufsFWbuoDM7McGAfL8vMlT1Nku3BAX/fsAWdlNaxrzbzzJLMelv+C
lgdTXyexjowCgiS6vFSq0j0Yqso2qKkTDrZmDynUJ71zPuYXTF69edesGhNC6eHe
nrEGyYFEc12y3GUFEBuIX56Yh183e3v/tO3RkPWMSigPZ/HKcdVZh6oecqYaT13y
duS2WmNtJMO9Jpg0c6KFh8+d+z/eOXnd/NCb3K/T+9ok7QxC0xLNhA89V4hGnoXM
13RLxeLen06kYF3uaZdf5rTYa2enYEuC3few622i+pwOxP/y6mkSCkqopZZ2Um30
0HMLbgl94GLW2WIUvKnySn6DMq9dG7ZozoBdmz44mhxbxjqRDMNmo6e5QUuMnVgq
Nc2SeRktrkm/5t/UFDCVvdBCqfJbwgjLz5rajBUWfRfBhEc/PumopU2BDY7dMdbb
x9IxXRYu9//0JTMzcmUv0OFqRcVrj8v1zMU0BIP+Q3P2OQCjyGcAOqyFoxmh+r4t
tyy2sWdsStay4l+Ow50rT0j/NSFohps6spJo/QBcJp33l3aQwhjfo9DHr7SoOfyE
L13+iJJkhcEkDjcNNbP1zoKl/xAw7NE58USxy8iAXK3Cs9KkDhKR0EEa9SxgkJVi
IsP8EMNOHxqi5KbKfaRr2+zx6pKsalLwTCixLt7FDtcI0TobHk9+xyRJpN31gb8b
lCosMPmw6pfGoNszz0oYVMCIRTX3/5AorCrZyMLnfl/iexJN/3r+cmPIabDN5Fzp
7yCdaVtLjDa+nZCacVmDH0j2C+lbZmzPvEfPR4c4pYWcbjL16hkad+UgzhtBakCf
CDNoDLSdKuUWonYV0ndOlp926txsWRNQRZqcx9UDllsnFU62xvKLUe9okwsyc/6k
ulw0qPxfNeQClUyiVDEUt0VRuzIikrvjqpsnSuRIx1XxORDZyIXd8XXMfyH3IkCJ
eWOeQP0vT4f9zvr5rIY31wLh+8AuSkCuzNXqghjyTnEdfwCYvVtrZRFUG/fC2ajT
umo2uY55bwlsLjVn/ASD2dZMh/z4sz3UJaebAammRQlyyDeXEaAKRvbIqxBwmwne
aOtyId9L/OXzaeDwRkMrv9LwQBzRuXYQGdVM3EhT5ECqgUTwXHkolSHXfekNazzD
XrB+VHxvZ1uchwUla+TC7tPdHwkEaZYjozUtd9C8luvxOZY56u7Hck70xHMKls6M
7tamBgjJ/hiJrl0gkLtw65G/NOssmSP2nMBbqnpgOWELsiO9cRzhIom1SlCsE0Rr
ZKbUusAe1iUj4a39P8o0cD3/fK8LQM3ZpE/g1NaZME5b19fKa7lqt3uYGr/z9tEO
y4mfHIzWI4Izqk7Pc2Dbt4JRi0BhcxaI7uX9mFu6N9Xhh0nWvbtY67ic/oSie6Zy
FVkDIgi2TDPnlbbkcev1umhgKcfIocRBhuaArJL247hhjbxWB/3CfXLeiAztvNKW
pWSq3NqxUUmEV2375JN5SJDpsISHn4IiqUyz9ztncTK2VPmAIim33iKM644mPwMs
3se9uH7zQUNflyT1MsmZ6xWjL888mKp2pNfrF4L/swYq2ppON0HjN431w/Cb5OKY
tAfxmFLSnRmfESJIykUsIn/DG8QJMq6kvE8FGgqPLKwZkiHGTOveJnmEfYIrxrUU
YAu75GmLT/L37wC7cu9bcn+/QYJbMqkpqpvi/8G6kLjgA3eGCVA0ocfwu3S7WUhx
Sz8nm1cRMuozvbF+9c/VpWB6e5ltGqWYU6cF54dyI0qkKsDlPghtQUKXkl0IevWc
LFedGGDevrnB0I3MUdRjH1Zf6a6hlhq9wqPVLuu3WrA3WWXEwi3a4uIR4e1IVJE2
8Y1L4IQoCyqePEF1qeVsHYxGIb1CCVdb4zh4QXrz/9vlV2HPalS2jb8tjPXnZ4fl
ym82IAw7BanWOFFgW+S7GXnwakJEMp/9l55mKkKHIWW+iZdP/E0o95dlQRC2ufOo
w3A2eyYb+UNnWzInH92wq3gTJS9P9PfXjB0Arsz91VUg+OEN1JeJjHdYbp1KM9wX
24kGM3oiLv/QE3uAsTAFEW2S0Th3pACJTHIMFvNaoIf+1vPoDyvWS7K8q7bOuHTZ
57KFxpsKJ0Y2WcWJGs0hVEoPvd8neppSAOF/89kmH/Q1YR6VvoFhpehH8zwbZIXc
4dQZHTwjvsDYjRhriYLXEeYff9mccb5nqmGCm9SB50wdajsiSdAdf8HhOleo+nd7
SYZyK+gfh8Z4BDJG8aiL9aEz7eo+iAmaWd6Z1hi9mk00hZRMy3h2ugJGG2O3B8wF
erqYdSze7MYpeIEswKmBgvgkizdXxFZkx9WNPhxLps6d8mzAuFPNreb1IA/MVSAh
cBkZUn5Mf+RM2UC5OdSOJaTlYkzgSUPtruylFEcOYgxDjMYA0lEr6Gvaj58k/4oi
bXdK3uO/SdVAE2zkaqceN6nBFg4w1WNDATP35KkTrB4j17zfzG1sQRDEIn7e6TQN
iP3VLYp3WKNrFkVrbZClWqIocDdsbE5TzxHZTRRN/3mrvoOxEEw6/iXxJ1OFao6+
jVfNp5vw6zpjGEKHxYsts7rzYKDEITc2Y1qyVMfFf2zE1L7dlwzlscJr7HueAZ2r
0hjunOo6SkruVJy407TppZYpKcRzaLsirmTXI0qSr5GPDV4KwNhlpU8w1f80NjVj
4GehGOCxUJdwtPCg03nRCZ4mspM7RJPQHHUBR9JQe2nasddU6aYilGt165TvkLbT
D7Y0hsQwz34jWlOrDvZ3GpzoIqLQOMp0duRJ9t7zixjOb7Qk8hbxmFvnCSB3wNFL
DWej1mT1tEksidP0JAptHfhC/BseIYLF2bJNLHrgFHUR6MI8+f30uwgiJjNyL/ZL
LjsPhF/1e3mXHx4pqduiU722MwwUZtLi7XOZ4NWz2K87OlkxAVVCdU73jqCrd6L2
EQGiMnFUbN3AUwHWOi/mu+A9efp1AjHd/MigTEDO+44qSew8S+fHvy/BuW5aBr7h
LaqiDUYRIYQyStrxAUyb88vOKf0n76IvPqSJJeUZS0Q3EcTAgGeCkiWtfiS2KEwH
undhV4c2Lw5B3YDYuIukJLWhdPQlfqp3C9IztOQuksnE0a/8jBaT2ynNxzLgnqkv
054Ng6miHSqAK/c/uL63I0ex08/e8cnZorCKt4Dgm4/F2XW2hj1ugh+tcIS1XUU2
tQJACYSEMMDfrKn+TtW2idR1b8h42oZexTM4IQOrF4KzHBJQg3xZ55MV9IYy+7+/
pfq0uLAh2AN53/SoKzQOVHLtPxRLYBRfhGtLW7lgRH0opV1bwTI5X9MDiEshoc1q
7fWob6ONbl6aNtFMK1lK+n0H4Nv34r194EVKQdW9jHxvdfcLQzu8pEAWGZJ+kO6t
LuvQgDL80CCfbWcewaHnYVqMAF3RW8Sse3lC37uevAsWHb52Ld/YFkO/1zsaj2GZ
nO81D1ScS12b1hJQi4nevXo5dXPPoD+XiXz8BnvuaMrZgJckxUneuEJmPIngnD02
SNo0lk3HG34JjAsbnken2i+74+NjmC/2I2oRVvug/c62LvA8S1yf4WgFz5Sj6JWn
qoiwRmao2u/J7tsYixyt27M9c9D26HPbLaZgRBgWEqQVRsW0X7zljKFIyaYjuCla
JdRwd+i7tW6waWmuUrhpVtzlzEAEGqNN1JwPJlfOEAq2Wzyh2EOMg+low7vzcYpa
fSeDK42TIA5mnl0QCcESYy/Jk6ASgQO3ZS1hw6+LkumZvXeNc2l+x6HfNqyedDhO
TD0C3Xzgz1bZ6Zqotm7EUBTOdggX5C8/hqMvQDyRQvImD8aMD52PoPit1+gZ/ZnR
iUAB77GDIEk7MoNlyoeTn2QbwhoqcKz+q3rWgkYKWBUIW8q8YH71UFhjsOONje5T
l/2wmzAxE/yUqlwCBN+Fwl07yE66z/8wxIM+MWLLsSAPdi094uLzc2mX5F6/1D1k
GNMw7kOoAet1vwwbS5o5z1r1M1juN4Ok2yeeM/YOcN89lOPZzrUynn7+h1gO/Rq4
XOu77fblfc+R/dvl2UZf7mAulVkqV/vQOo+fDLp+zRgiV1YTVUAMH9XxuDMBXN5D
4vgJNP3eFMm6msQnNf9lTirPbziuJyGkACTPr+iBhKGCqvF/tqI77TxiknkfssE5
oLj8ZjCT9XthxqezngSoeOM7D0tf6IPiFJ3wKPhWk1u1qQzW8Y8wPodb73TijOwF
3H9YdIpVYrlsMp49Lq76Z7yI5PZkLC27Un3h8tQO7jATskOwvPCvk322umtfRo2X
JuMM4pTAlLlP9a7l4VEWYdxYJbQqZC/CySu1qKgvKXdU4FDSz8qIuPNvtsISPhAy
nqhlKnRmZIFqjPIu0z5OuX01RoVSOAuCHqeYV5a317LaXyKq/w8pQIA3cyUgLEN/
rYeaqmVssXYhhK86OfcGDbuAD6JSW//BZ9nniwG7QvyQWcmzrHAvsWq7swfETkni
scY69u/hCBZfMTMhmlmUwEeDHkS2gzhry4diZXLK7J4MJwdyTpHktDZ6w6vSpoIn
zW/p5lK8tIgtBkB38QFthacyS4AmwnjZR6QFxihUR9i/10wcgQmWRFbBXyZ6TTdP
zqImBrTy2pBctevx1R0A7YaC+sjVoF+IXuxktcOO3Kl+3x4yatvzp35iMKDEc9GH
PD8+j+dpmut/esAFHYJ8eqYAxq/XsyXaIotaEYnii3JoXetcDL7OsobxnOAryGKG
eZgg3wiJs0hRBWQUomPdwBNIcwCys7cY48gUSN9BqNM+vUI4HcM/ihmBSPBuO5Ux
+A4bs3b+mpqD/0WVgpumkke/+BCjvRVwZLawaX0nG7F3ieZdlYWjAWLHBu2R6vxJ
87Kx/lXdW8VleR8Pi2hpcw+98Eb2Rh9/BEMF4CF3gKmwqdw/jkNkQPS5GaZ2TrrJ
RlgKvfshKj4fs9I0pJUPc4ehws/D/v7I1xLJMm7eyIlJLnkX7ESKxRC84/1SWMMb
iBI42J4MCrxdouRHWAvx47MGJDZSYYQX7PZ5Ks14Hnu3VP7CbbrsRoj/jGa3CSgp
4GZ4UyO/ViD3Znxal65Zj3qTggfqMlIfxSM5l9ISnqyTT570MitcsRfSnPndJ52r
ufwBg0ZGaXqM82nnM1cyJgxm6Z+TQoZlsbjTGgpyXsux3e7uvg29KfI0DYwR9o1h
VX2JkJY11XRpEY74DJ+xxZIsXlMxzpYnr1CVxlpysEQ+cfJWrpLa+EVLA5ZzzfMA
DtvU+32t7Mkq+Xyyfnhw3lMn2wRBJb9uOtQVQ3BOjDNBz1eN0DNHXLy/wVkHV5P+
KFS9rgE/JOHWWTfBxZZgSEUAx4kYO7M/eD64ljMzgTQUyZwuTw+qJ7Ml8DdpWj9i
UNVK5z9VVZW146Uiy0Rvxqh5r7PBOQj/0JtMYaFiX6UAXT5QLh+FBkaukTFkdlEK
JqmrT2VWM177SCmMGqtbHJcZQs0NCUITSTYH0WufXqgazGaqXAX3OsYOUt9sph1B
Z+Lvpy3ZKv+eWsQMuUHskicLTwqts1PqLp5EwNn9VqNxaFnwoADJm6eGZIwvRSOu
dmw+H15eOsuj1t4eSuAp9F2GNQqcQBYOrB8x+AZW5Ym3UsHoQSw2MTQDqhLaBL5c
m2f1SM+K369Gm//GC5zSIA5SH8qDCveIBUXbvB1d4TwR6Wfba+3g59nEbc5fgA+9
nMWlNUbRVCPUGL7lRHMfJxHe+CiZ0L919Cmcua5Ls9n8RNj2YW5xjVKhkCfuQ34I
5NJyp0Ocs8HQVz0pJbptdg0p0G6dWZAFK9NT01aQ8+QOVNI6OPcGTz08Czd819K5
DhlGterrH0HzUa3a7znzo2ulN+5b0agcVjl6XU1lQdbiTYZwcngm69dYo1mJG739
JQFNCwC+QdrkVmYjHonCScoCgHnzTgdIkOcB16+YjmVo63G75Cxgee0Ko9a1ZRbc
9HY7O4gjh4829z6la4SgstFHmfw0ru6AJola6sjJRVV9/Lq64/KFXxEn24n8jqDf
QRLwaczvQStEJvh/8KXIA6qGm5H8gA37KSFDcFrByH9jIwtqz2BR83iADKGoqWOY
oBTk4poQhTK86A7zzYzaUEIICpdTdTsX+yszHHxIEX97r0UHf/BR3tne2IodFfQ0
FyUeYIm/pBj085p4pKIDJ2vm/zxMjSzwX3tu1wr0GbEh4SHeHnf8FbZzSLTFv+yF
bkZZUqSuPvpKHTwXwskjwe+4ft+vFvqzThvXEeIEmj1laNurNX8S91jMcNw1NvHQ
rZRVVC1mZd7HC0JBacSqsYLDpzFHSo5KtGOpSM7qS8xbl0v4UCt1vujN0badzeZh
QhyvRR9r9DGL9dcYbvuU9Cx4iW+VO2DAc4lBOMob+2vJiY6majBS4ZwEpGUDv9x8
ArD0OIRbWCZFzIzyWJj0Y1I0r1kob7umj3dptpIF8yov7AysZTXMiszsLY4fCjQn
eKd+pXY9CNUmPaEoJzhOp2g6C5+IljCmiqd3B6uh33ztdGeHg4DvVBkxHgchMVmB
MitY0PxdVUOKH9tsQsoQ4XdxCeI+el3JP+fORDPibbepZBykr8PuMfg1F6lQpYhw
3UN3egqrmwgb3AGVHP9ibxCGod4CIbCu43c1d0p/qK3/CVrQR8Yxtxri86jS4Mlu
CjvFXxOvOith2V3jhJZcCwm1w35/Le7FrTaF6UUPCbHWecBe5aB5d1cgtWKmiciT
VY974tAXjcRHrevUOY6klny+Dkyk1TNGSKSCpSetlcc4EIUzW8mWbCE8jE0kDDPQ
zov5wH7SjGHejSBhgqwa5H/jMnPNw5KvEmacu8WYrfmoL16M20JBjiL+h7yzEFOz
x+mQNn+EFahPRnY0//0vjlwVZGyfZFrNu9W47nTs1bLCc60Dhci3XnwsBkVULGpK
QCfw8TcZLr5JbXq+BkuraVB2SF+FF4fXWV1s+HqPOoPqNWfQzEA3o7vLA4Lv2qrI
BD3+J5IueGnvboj0remg40BjhrAqJLWguBCkSXAopHxvqeCvGfwaszbdLVZCjyOU
w1XM3TGgf6RF2yKLsyDute+uBS0TnE9rsLJGUE1M7xfwnlGmx1FBjYhFjk/4Mdkr
ysndOUyS2DRDL3ietPGDoqC5EKr3zc5P+CjUQVWbCf45hbhkoKaprcdFKM7PUI9i
YBX7lUFJDmM8BJ8qZACvF/WPopAIXb2z7aqoAwL479/LxAhd52pnnpwEbIOroMHs
wvQG9v8RPnPT31FljY+J3HUVCsweJNTDoswB41UaJiwwMkhA6ATB8yyNuIwYLWw0
CvWtV8nDIwHvfVPQPjzBMXLoZhbAqurcK2rka87OP8vfIXtf3vH1yciKsANw1ybU
/YLMcxKa1gEK9gB2EaYhsPaT7/8EGqDh82kWFLRWLcAnz1TqFM0JIkycGluHRQiW
OxDkTTRzoFB4QEO7SPuKAw4Tf0lXW9MlO5DR7SFFxxhu8UZKQizdGYKJVuz44fRn
KzQutDPWImDYSRg7XH80LfiK8SPoF53hiX1JEcSWEKc46w/O9ujGUDFrkP9dM7lH
7p1c5SLpi3zP6rRVpEbupyAJceGcqsgq0XdDFW3FjXcfedV72V89cDhVf/ElauI7
KWJS0Oto2rzMG8/KiMG2dN2WkZwvqhhEmSO9VHXgzuyBKhniXdxX4yELiOIKDR+o
MXUjw38aUZ+oWyuSJUO66aKJeny0lDYqDKAgr6zA5Z533IR6phdOCR+mD0hruGXy
YpsG4WbASAhlP6vBlMqFcJaGraEqm6eVi1B+BU79zfRA85nYaWG+oA0QJoKhmbUV
kuQZUnxH18KzqTSS0NUtvEA8FDaYOXVDyZbCr+wMQTlY6lOcdLqAbjqz5JCHrGc4
9hE2B1TVRA3iNQISwpoy6BJPLdYm8H5dzOd1038hcqa0jP6dYDeQfV+zmU4cffCV
a8kW0fLzhwN3IDEYcUCSbOPUdDqJGBlMPfgqPI1abDnPE2yPA/vw9R2LuLObQAfd
OkJj7zl3KGH6PQL3Dy7D1RuRIfsA3SA2oliwi08j+s4klUptEKkNfJPcQFTPZe2x
YX3zV93G8l+9MEKBcZBZlIWGgYhvFA3tAwMtq0wH2jsD4BPtjH1Fzi4ywphiO9Vv
uPb0FmOdv7KLy/0kJNd6eq2Ek17XcVFUmbMOBMHiObCCZYN6jflTARrkMqZZeVXC
Fi7wpYqmc0Nf7/VBzOJgTHhmrT86kMgAcTWS0twDRRR3aXjq6MTsZ61SDSwqWZy5
11QS2I3zrqu4JFrnl//HnBE9fAC5fkFCQj0noHoOJxsfib2ttXaGB7Hv+ev+gVCA
WHEqsLFJ387jVp6GdPVC9FClKpynyGTO0o6FGkELTh6s7CsvsK12s+fdrTS/WqJT
CHXrJ8MAZ2tTbZdx5M1NA6FmAAgsRkuaJvuXvlFk8q9QhwtrEZkWeO+95PvofYFz
QOF9+Ra45drk2kl6Z+Wky3hIgeBa2t62xyCU0Kc4OSeV+9rA7JyXOWrdZ8BeEw/G
a76WmBVEseuSQ95n4ImHlQHO6CFGF2LeIOwMGhZ5+rJ+AxpD2rlrsQ5KC5sqenNk
sYLkBpna21Br2aO2BKVVLGcYuDib1eAcmzxa7tR7/M1GWcZ8HQeL+y/0NoJ5w1A7
JKrBj9uEPflsYe0ImlctmeKE7VJpVTK9JsN6L1k7w33CV6YHPuFvWelIOZ/ia4AV
rXKautDreQ7ARMzujxsGTV/M+dqEx63HLSElRvnpA0m45jrr8gDnHANDIwohojNY
cJMVzlJhQOcVlyUDZcS7do7tNsxGfubh/k8ocr3xYaO+SL89XBCsMxVnJdqufbeN
0nWLWRZO3OIPfb8hfhv2tYdTr9BL82v1J5cibYMUgrZlZDF2B8cChMBxdaEFe9MM
vEQ+XXoVv0OJGHwyu7ilBZgt/QzU/ZCsHKbtwhsq7B94GX7kfP3koEjkCji+WZez
xAs2hqOlo2DQ+B3EfYZXiFjjKJNGDUrS4czI0qO/8UM6F7CnEE14T+s8BiqgriMU
cJzBNYXDWvznjtRK+EOQ2eLAa3XuH4KIGDNg0OyklT1Q91midYSYGCVGO/6/TP0I
q8sY/AC7SEAs0CjLWTGxRTG1DpkANsLSDtkwWE+U4ZohsNbh13CKACldS8MyzX/q
E7roUYxpWjsPO6RUw4iExJEahys95hJN8YJCZ3xAmnuWh7H1Oof7kfgHD3+02zlE
rk2PLv5eIUS34N1IATGHBaVF4Og67enA1ekANuZK2ikAV+3hECCqoW17+cy/YNLe
Q2d5wFqwBQD/QqKaIaWrvk1nYDWZwVnVUOe9vO13g6j4l4sDh/NY6Smcd0ifHJV+
e3SHCYlLtiJkf/7riXr5cApL1YRjGMZ72ArmRl6jrhv0jgClOEEQDYfXO8vHuOtt
Lh9PMx9FhCwm6DZKLNUODgAU71p51RuFkwGDfjWDNhwsbcIJ64XlUOPWc7JYVEhy
HmlOrL2WY7GmNuSzQZnGGQ7+j9Csh7AtlCCzYJ3MPaxkWidbyW1Mb1t4wmnBpIgz
NRKlSdE3VBWRQmGN3aXpipsXfMs91mOireLBMEffmXYZvVVTO/aStH+aY9PDXRJD
mduWX+crUhnCuYyrAQVMPo3uoypkCAEoq7AVrYpHfkHkA/0BiE9fQt8UAgde3DIh
q6b1P/RmCu23I0SbAP8IUFUvHHDP8pFavxR393GxRl3FDV4ljK4+MBhQ8i0sSgP1
T1ZmuvtJ4hsaoNxIKlvewOjSFjxrLcLOsdVGwusgA4337q8BIAzV2SuxtUsbKeWH
QvHxeEt8kJovG5ZS/y1V5E+JgXUdRYVy/kJyAJuaiAIxX3Zbt/WInGsttf6SMsb7
PF3VUcL2hcQL5wbIajBmKYxoJ3hvU/3TcexJvazFk93rDoGZ8NKRKjUFeU46YXhU
WspUh4BmUt/mgl53Ch7haqZxHM7NYK7YiqBhebA3EZWsmumDfDqN1rav86mj2/VH
XMPON4SaMMsJRz+Gg1juPPRAJM+aWDK+StKpMiM0Fi5hRjvmRBb3DB6ghlv1eVVL
fg1ead5IORWyx4YQcvGD+hRk4ElMultVVpW3FHGpHPH0NdAxUtYFT6cPZOarBt1x
q1wHuSFGiIQEuaFWVvXEm72jWxPnOVc04/ZmTcGUcKFzWaDOGKxdYqg+hR2m+/Iq
TccSRqpxijsNE5UB1uwzK416wsKZdUMITWA2w2XaQm96ugcg4CcI2DbbyzXLjo0U
gH2cljPp3XFXHy+cNg57PNDjSiawWB5kEsXzsRo7dQroAzrt/IF7/8ETsIqF2vjS
/WWepaHZ0+/sPq9IuyE1f/W7Ib1Ac12wqqbuinyX8ZgBrcYaNgjzXrPWgCz7KpJ0
cgc9lEYl2MosvwlaYy7xdhOH8rypWiZC1ty9+EzMlkuxg75o6loTTJhdsVINbw43
46bxPZpW01ODF0dVCc0dof5kkbC7nt2+Z0JvKUxCTCe/xuJDN+d6I5ar9pjSh6Bj
7TmukybWhJlB0+memdUJ61P8QqSGNomAxxh3FQ8kLlsQPAn7V9FWIszpECQgbkis
ScP00zknXqGNLnZsMUEZB9vMHA/EbXiwCyEaUwNS2F9c1yGSUexi+Eddm+CcmdSm
aZrNpZmAXaV57mR0RwBCw9GVAotIPTHPNFAR4otZOBucJwvpPj0a3L2WJzA2ilXc
3BGb9UtgS1muhwLR/LERSlvwg5P+tw600gPMvl+pldOMP3bAHoYNMugDABNtlXkv
yj+KFEKfaSdsHEuEe84Tvf2i8Vg//K/XIH9f9/ADK4P12HzTa6Rgu446qsu3O50l
mtFvJuor0/m4NahWLKRfOvgR7QA5OmcpxZNRoc/HysJcgtVxP0Auy4IJdpteAQve
m+mmsn6h23QI3PeGd2xYYFJubiBjVJCms0g2YrtfNgZzHBWQSuSqru+3H5+cLiVd
yYoBmFjFdo7mT78Q6HXIn3rhAc33PiMsRqnySLAa5VQTH5zBuBsFNJL81vDlAMBO
ilkLQdIcEfITA+8hStxAC45L09wjYHfA+a65VgPS1mecc0NuWpShnPd0yuSlKOTJ
gQV9cUEIiisvWKEA/MTOV7Foahj27Jrnmi6F0H70FAIx7StsCfnYtwpLIVciAjDc
LwxfiHI/7HtoFTqomDX8oXLJmsKqMF8dvCxpf0+3CQ7q7VSUjIDNuW37lZqZBmnI
5moX12JxWSgs4ioRZM2yfTz1eW+puGrlSMQsO5UQSCqrl13Zz+ZoJh4YuzxJoztR
HXUeevyklP3XnXyRwduhwaaXe9K2+YfbAip/2D0IT4Z4ZLWErL3fX2E5ZInBkRno
jAd4ec9h4ZRUbf/18qsnVTbZNvQgJlBNpJeMs+C49NQG44pJtPwh8vUlGxf9s20U
k2pF0mjTejEHuhXfhViZ6gpREsX3a8qoIqSayqN2dQ/cKClm2YXZewP1/4ChxN+I
n+r0I35zPDsOvcGJzQckXfUSLJuPnlABvHUyl+LTFkbhFJnDGx3T4EMM813uiadT
nvdrOQd9EXScLlGHwnkdYPHeluhoHsLj5QS9ie1OIpZ2q4NaTNmNmcOX8dwTEKp6
MvQYdOeUXNz+tXuZI9jdeE8JE/djAWfs0ZViEywiS3z4vuoUP0BB6I1u8RcohfRR
Fwrhy7houCA+Hbdj0+WFdTN5KMnFpiKmJTFoyQXOIKaNSD0M+8Xj1Lh4yyJvjCwN
PyP8J/z65aR156lcqcoKVsLP01vZL47nQBJi0Xq/s0d0AmvK18/cN9sZcOHhPnEF
dwR3N7x1K2nqMvz4dGWGx8/KbOVUDQH4tmIVzUBSxrHSivjFaRIEFYQZJIyD0lN5
PVpjyIZCLW/b38gQXxFt9Af5+xFAtmjCb8HA3pzTKXjwXYxjUqK00vOVimvKP2hb
TPp1lEjP8XLBfguAxz2PeFMDVGMLrdsZoB8Hdz5JY8IiWp/SxMp+rV41kG+K/m0d
Kl0u1/Gqcy5h3tGz+z+jEzu4QFA7gvCMdkZKybyB4uATvg5Bp84JWXyZOgpMIA3i
rIUivqO/WarK4KhkXROKMB3gcXWZOqvVpTqU9qigJMXtepiaPdy0dWCxGDDqG6yl
oMoEb3muSseFBkoOdZVEiIOViWMpnjRsL2ldIIC26MLT4GKTFsA9XeWBmNXrthJH
HrqYGKgWeCtwTnFK1OGd0QTrOjxcA5cBJljsu2CT5MLs1XVceHWunTzeOg463gT9
IP/Cdd4eybsink5677boBl8Lr2qhXCuBBbS4iEYTP4sevy3T/d1+nO0q9/NxfyTW
pHxGrZlpHvBz2NtQcibgQb3iPqnFEo4tub7ZjGFQbC6Ppe98W/kOy1ezYVsSahWp
3NhhovG5+vfEt6W1FKVeK+fo9WCYxurCc5A3785Q9t2xtLVtu8KN6KFa4jSBYcc2
p6qncTrMMB/Pu6VOgKrhwb/jEskEJGMCID7MTo/TT1qBcvZNvvwwKgRl6jfWiV+C
LMr6eAWZySQ8ia6KNra3V3nbBZMbcsyO9TwM7ik3jCbkMhbDzSpbbKrc1uuFyfkV
KpFI7kmz6Dl1SY87788cskb6holURZJ6srgb2slpn8Fed2q+eiOviWv54H3eFNq3
VLX4sR7NLpo5JYMZd9iRsWpZT/eFTPOnhw7cGr62KZKGX7dqqZe/93mCfPiZq3qW
MGe3dYnKB9xK7wYkB6dFZeKCBMW3Hn6i/AlixJZGVbWRcRtn4/Dxso6PXi3NAQVM
ZFEhnyCHexJkoPzXpkC9MhoW+mShEz6WNBqHA0IjAnjlAZt/sL1LKKg232KNBihz
Kt11Zm+CajVnHSpid9lA1KkwGaq3f4X1H7nUTeCCNtLVMF1HN612LLR2kpJGRD8J
KTwAsk+horNCQrmy6C3mo995DW60/U17scup3i9qHmjUggS8TTF4NCJLMmOWsuGY
g2oQV+X4vv1u/kxPmX3IWYMrIjXram5BfbC4GFXXV1MOPfOKg1NU9m7cjB6pbPS/
TzkInW2Ph1Mrx1O0PmG+hLArTlGkrobFTMWPeKdTlvcc+438U4t1xAAEK+tqjVE9
kXhIAYoq89gQlxR1l0afNzpt0BDPycQyjg34T6hdwmpQyTvWs1G4ZK5IbhSG3fhc
wkDB1z8jBN0rbiqodLKHzakOTGX+jkC9qxP5b1QRxiRqe0lNBBiDcaaP/3MbAreK
zp/ytZPa02/9DO8EWx6PnecGwN8hYeHbI3aB0GpTSAKYZDwrvq353z5mOeHX5Ew7
wt+d9CBHlyR7UbsmnhAOQt/CuuRXIMhbwphTuXDCD7pUP/De1Bh+18YVy7q4FnOk
/mM6xOfb9TQ5MfLzW/Q3WbUJp/+pNDc0XUsIHil2zV9lHo5oYoFgL5OATfcq9izx
g26tT/Uh+L3FyoAJxOLXSfbmBwB/MR66IZ56YF0UB+I7QxgzaOFZEHGDoJeBasSo
LHq/obhVlBRCFINGfQOho7X0h/kjA/6sdpWFyzSWqcCtrZnZHvh/FxVGn8u3y5vA
dyGK5sw+3yy8dQhgSPpvhoz5CV6w7OOhT984fAZLLfN1FBSg7JxJvwZhfzpEbjQa
BXNm7+OAy+kmf3A4eXLVWjqDMaYV562DuH5xmx4vimswDKCwT4n9dCiP9PFn7huE
aK2i29SKbwfRQ19205qskKN09dNDkE5pFB6YRrqdlQ0Et021EL5uwQZ3pnYatCoi
5rm3PhdP2jkXmFk19SUyKiadP4P/P4Kcdy8uJEpdvBNgVMv0dFhPm1/VZUem+gWB
J5F2lfbf58jUUB49y6lhMxt2FXt+MsUeQXLU3GeUIcDt7vwPzpO8lwWIpCzsX0qP
dJrah7lwT5Hce0bkPP8pj3aQwF16CtDsyx/A3+A7/dqCdkb9Yl9t+c/k6KE4ixm3
i3/iInbe4rGr6QN8v72Nhtp9jSYuRx5p0wSl0YR4D1CpyU20FMSBQelb9gUTqcrC
w14yz8vWd2MQtkOxGVZxN1PkHLXS5zH32y125eLwM/HJxIJB9Hkw+05dKYFD7+6Z
zGO8AFmhQEIQh0uUQ05s6QJR42Z7qzrEfZHX7cAqTHW/SImq3tojvwybKEPJ1mya
FzYXxR+gMFBlSehfLgur7oZ2J8j2aSxoMkVqH2DXhQtm+4str4PnUT63pbr1rdO0
PuzRWoq24i6+Gf4AzkxRAFCIoaLjIootdOmsYHo4k9r1uu0ZuWheGtmE9vkDbMv4
6pNlpIip0ZuoGbsP4nPbhqEpwml10IQtAo+/AtlXPkpnmof0ZBod480VTCGYDlSc
zrkmN+5VBQDgG6wT7XQ84UkC2KP+TRy1PtvWr9EmbKJCSbntWevFO9K+D+7w1fHC
g79FBxblBr23k+jxesUDyibFdXV/qgMdy44ogyQKGxhEBK1+N6pgMQlXVEcU8Voe
2U2i1ZBK85Mzou7cGCksOUZy9E+IkZdNvqvqzU/Lw8nRVOE7RtuGUvpqBxlcQzxV
cw16F4Yfi+zdrY3NmICI7VL/n5YF4UUhAKpXYIhgpBudJLneQt9y3gXCrXJmSeMJ
GxXxZXjBz2x8i3oruysAzImsT/Q9IRuR2OIOB7xxykLr26hHbHL8uwk2D4kZJkuW
b01EHd09YqCxwZf7J6XuOnTECkwyV9bdCq4cU1BejC56UJ+QcuhgD12ZzKDL7opk
Gwdh0ndlqjVy2YEEL4nCcIj0WJN1DpRZaUDcJrxHVdWq76oRQmfZCPlkdE5OhSn3
r5xxgrWqta1QA0M/o0XLoIC7hUBRwrH5+zlEtzNwPJsPULz/JStUP6fnbmouXYRa
TaQlvHcIs1fpM6F0RS7vw2Dklf68qtWV/7AN2AIxm/cycs7wrEk9+rIHAKvV6wbP
TIHAGSvNl5F6VbZ9vWmsQ/fFIo3wTg2ngBtIfcCZpowNJAcDMsI0rbI73lHmLny6
pxmgoafC57Ehvlp4b9ULBVqvT0HnCa7PWHvk7jUNHqEkfRfZ8cAkvuckwSo3gXZC
NIfb+IxjDg0Sr5g4DnKTE9MCl87195KoWMktsmcOFbjkl+tgObJKm3X8Q9OtTTBd
gq/Od65LEfoxhudrN37cD/Xcsfs2P6HHcHf15rxC9BbiHwaNkbuylzhEhwN9Nh0X
Mcood+gO17OsitojV329pq4gJD1MbfV0oHzpZc4J5cATn/XXgcpvau07UXnGVyB/
DAiCp/ExpqC6Gx58KrhcchY5oJIsfmi0JQhphe6iRS+Z3G68ZLobqrVNYdCXQBNN
U/FTaYDzIZZvTPAmeWJlfiKQNkV6sXTEfkx+BEcU0aenbJUHq0YlxkpNzE+bDPo6
zjRbhffDdGca0kG6Go6lrEkAjIYnG/EoU82NtO8+IlQZaDQPa0WWl6Cs4M8z7RN2
N8QreMUAzLLhMHDpRcBhTWdMSJocGVXfx0KJgiJaPTNyxe48m2RX5bK6hLDIpXxE
KUYfNQtBYnXIfc4jKPtLYI9T86+Q6UGE3LSP4dGe/KMR3bWJVkcBESvXrnF0ivkj
QpAXcTpVMTPEt+xJkIB4IZSqUA3NkzhLJSl+HYhCMR9ITkqPMy0zDvk0Nj4NM9Kn
9D38wDoHSGjrr51xhP2wS6/F068m+COkCfEkQUIWNr6KbTORFp5n/GfEkH6wzpy2
qVqHvGWsuSoSi+03Yb3ZvtcXNL+wiKi39gHLj4ZBtSwthctL59CR2j0Psc6rgjAh
pwbgljtb4jHtK+0ohjFujZiDhezPR0sxwsvT+1Br2acDnwz2OcSgugqh2vBrT6+o
41M1Mms0hNR8C7I72t80J0mbf6qD78euo/IIUeCqWVRsACUdMYfEv45HFEshb7Pa
KVO7glKNbz4mwi1pa2zlPKkY7oXGWeEB3y7bDoWjSBAD0bJOrxJ2oUbcztJzHQoO
SUUbnt9w+lQYel9SeT+2FeoYLrA523QX5Bk3OdHjMc2K4v+Wnyc31XfNlrrojKNS
7wIR+toKG1rq6Ozx7sSeYbCUZCyABJ3P/rPRrK4BirMEMzF0EJ1C2Qui/+rLcifF
AyQSw9CnhEprJ8csIPMQKOZpoRfdom9A4nI24My6bLTrrhxOUs72rIQ0F26rLmGi
QpoJTI/JI4ssKx5vhbx5Pfu44L48jlQ1rz93cI5yCTCMpRRSq4qK6tgfp1pHCNxw
znISRs5Qx4xQVgF8/vK5B6sKCM/KTWlhWg5IJxgv/pvLsxU16uCDZqw3VAx/SfvF
EGtQ22tvVq7NfNaMRw9+JS6Cc429LRyM3OyaomwNwo3bJR9gbJhRWaHm8lUBvy1f
hrRpKBTNbeL5/+MdCWXP2lcd4g5NtW8DwdtWLYQzm/NoP3zRL7UhfEaA+5aje+f2
j7jXBIZtLxO1Dut1mzOuB6wTImF9EzJL/KD3my4nkMGNlLyVcFlqwnIoaBG3FjLU
3OxhyZ3tnYpD6mvkKg9IAB8TsJ3puw7+W0qNVuLqvW+++BS7GX7JLnx/bVyebjRp
8SZ9T2hm1Aq4pbC44oFOuuekxf7+k/PowxSLwKwPymH1ytyBmHBt1bgT0oDNYDrw
uaKsnieQ55eDh7YNM2yzcDML99V8xQ61h5WQX1uPXjx3QKO6bqC1muGNMVCKR99d
gLerJiY3u6pk6xWqiYOxrX5D7w6X6ok3bCGHB7DvkiWUcdTLNKk8bloQp4b3QA1q
Lxj2zqZJgfmomN3eL+HJaLLbMlXjsFpjdHxxCiiLBm6BYRyKKV4nPQOTbeFZwLTe
qcZjGLGyOEht6JJ77ngDez9iXqj5pGysBDttgqDVLBGWiOVaYobDmWh7aEK2L3F2
q+yHk9Su0McXbfdcJC9a6a702ApGK6HT90lkjA6GJizw0V8cuY3jU6IbY8X5bzj/
YQD5L/BtKQX6AkaWEJt3/QNupYRBinP0F+lS5w18Sjy++ZrGidfUIkPMKputdUrz
QhZSBiOT6BodEnWIunWtQa3rV+VYjoUhED3JFh/0+KIzesXGUX6Kyo4qjmyVf7hc
XeuQvrQIa0aBKDQpu1yLCGSQFK8ZGn8zOLW5uvsOOUOziT15UE/XEspsj3gjBtji
bnrAVXSY4Wg8xxDV0+dxYPsN5M9seqMdrgbtnU09cJ1AGQlTCPU3Zr6HjQryTO5w
ANsDRLH4EQD1sXRvVzVEjVkZoF8lNhlP4cSRYa9V4+qL0Amq/cfZuNcrlYG6Q9eX
OP6/MG6d08KARfsF/KE1HKvR55y4qSTnwQSkPRBxCWsvVEL8z0OO33Gpb0iDvYff
xh/YMWrWVXqVD4cod6Zc7M/SOdZM+Ymv2nSOsxqV1vBYjvIhGKYt8v6/iGtyEudL
2UMu2uYUgiKQMUKsm0q4ThOexvygjPGu8x8gcs++I4Fc2FraXvJUOjx4706pQix6
McnNlRn7EVLW5zOYIteXps067uZO+JRsvv3CNj7eON5HCpE9R9TzLBSDg5Zn9lrj
rA5djKxeSbr7LlS/r2m08vCTYZxzjd1w1sCs4V5fBDcObzu0oPgo+rI50gexM0Gm
qDurp6Tm+Je5WO74Vhwk3Mf/PGU3aETJxZ8MZn9IMq4/rYl5BBr9cCUqNq/cHCL2
nD1PRPzbsuR13nUJf2QDUuBmwxzKgICfsgOTCCJ2mXqcst+gunrmI0x8zzvUyNFG
DSHwXUxqhpsKYUWF/NfmPsxdIjddu+2+zMbdBnR5ev4dMJQHiNJ860k7nSR3mszv
J6FL1tKckZfnziK6OooFJb4jjaM55ZlKgcy5+W9mVivRdwIMnXTDN8x5dVpG0lpq
59nWbF9vLWMjxI+C2dLBdXoXZTExnDHTGBpicNDAkAgktyt24bNFYVbKDA7iZsjF
XRHQtzgeRo8b8dLLsM9BOckQq3udkNbzuAukMVY/uYn7oe/YZgJ3rxIYsepSn6f+
s9zOn4G44WF5eNkhSw9zp2tbpG7KDxlEXqi72pqBZnSH5vUsKUZhpExyeyAieGXJ
zF3WuxdeoX6F/tGc/nJAn0jRUNAu5za+05eQWB2a9Xj89m5fJAprK7Xh/16q86uP
e+K095bZ5bYaudY13h9P4cCi+S/i1lQAyJyConBRNYvABFr1LLNzQH/TxzCa8aHl
cjTYXQO2S5nqf+mOVMPnaH8bfuFged/M2nkAygePVZ1uF/qFZ8w+/ydAJ+9lNUhS
FSXP1UJVmXmIL/l9dkJUJWSELzVnHLFyGmrZJDFFFaH9rSyVOUDl1+j9RLasg14t
nLmj9TZ4U5x+K/PF/nK7ex67C5wBUFpaRD3JgzsTWVVIA4M5vCmYq2wgb3Oz3rjS
Q6PhMf2tMSdjofmS65yhxyczLWhgbJ/PXxSreO+4hLgBy9gcXs0tjQpl7aDRU9Uf
iWrFtXDwJPcwoqQx+q5M9OAbQFcPcd5zH0o73FzYejrCqKhb+rY5+gmkMRUDGRLb
vrIS5lb9KVIkeRsZdC0ynkILC7aFTZUmQ6AkrckJuZTImaRMXlAEYtFqYm/c3KHJ
jIYvj4VBNoogfUMY+r2EvkaLrOoaEHBN2QMKAXtrkYoaQ3BqGq135SbG2OCecmsf
jzcIAlQDW5O3Nlyk4ab0il0SJr9mi2rJW7amxIlydmuMHt/6EuXfL8XG8+s2C/Pq
SbWW7GJeJ3NtuaG1LfbOm2to/T+V1t77sRf+ZeQDFFMzireYDt991r5aWqndVLS5
VXBDAp+Nk9TCHJ+sOBsKq4plXoj9gtRVYWwZiG7Rfr9eepG5efQiYRxXn2JwZZRm
19Xbe5jjFV/REQq6+9S8o0CCmqZkQ3OhdNQ2PVXCZbtZH5X8Xx5AoPm/NNY9OWs1
sOTWQtgYdmUyINejWxEmsESgwvzdHaDWnI4XZh8FZcJt0Gg52ZojG4Tptuihc1kl
22lUw+J7WtTDOEOEqrH+GxjOcelolzSKjdHeKVUJ6Yg6x3ZXo69w5GJiocs2DNqT
sq67ft6aHOIj2KzBs/fcitDNOXTlMdN3czOg3ormvytuPxaBQ7VITPoMJFIeqWxr
uAvZQft0/lsh1XcL4w3la4uPe39kceX+I4nogNv9sljHYvzpwEPJy+GpXfI2Fk+I
70K7Y/M8fSHnoiIK2F4bJlHgkFuev/sALC9/XBjTGa2WcSoinqwefPWGCmg/H6IU
zZLk71nSnePe8z8ZasSsgWXenCzxMCwf7kZDgTOOdui8HBIe6s3e+BR7XCvXdHsc
kKHk42yWirE2o9pj9dPexYShh1k0prfQ8j3RZkeLCuqoqKoAuCEHkbUmrtJxBtTZ
TSfFcYi3QKrwUCR0LxynSg6jWDKTWij5HAwgQsSVXOfHHuEEbF+LJqSqxU7j5M/j
YEjYdJUEB+xKa9hb2LCEHyuNBHatd/cSU9fSjPkCrgvlLDf7xf0qUNF0VnVPX+D5
3Q45DgasELReG2u+ar4Fg1lboy6dtTiCII/bfGnWphR/DG3qJn4CGfporJ7tydxX
rGFjMz9BX3bTlj/VvAhMw9lQdr98IiSmMbfnM3TZwvyyGuPUs57HYif9E7BXTrbr
Itv8nLfg+uCW/5rbEjOyB9ub2FQCMIAek+O5EfIe6stpoqame6TqlL6okXerotVr
sfqXTkPwpW88ANVLyMD5Pkz4/r7uAyXJBrWEqnwZIs11Z0bSUfAEWFyI6eRB5JYG
XhgxnWX7Bh1B3Y3iEmiOLXcQQohp8cfFXyyjhMobqWgaYQIngDPR/pikr4RpC1Ir
3AsSHrp0vz8ZnQ0AdZMQC9qGoxB2BkUoN92readtrmDhpiOHNBdT9NHOxcRDFQOq
9j/PG/c/OMnKPGl64EEHfkSNN/3kXcbAl+TjvZWWFjMkqvlc0fX8W0rfs2D/Dims
k784N6zKOpC0yLDf9e0GuL2p+0wMPihqP5eMbWkM5o46YyRUKCdbltjFjQ25/7zU
AZb5HRFp0Nx0KmD9GU+NQqL8ASLgaXzXM7cNL2IQruLPYEn4ER8rG/7zrxNgEqn/
LiTcVgDEXOKnfhBmOyJ6Tqg59876ZhqoMdfeyVzKq5EtFUuJhl7jw0LL88qVRkXu
BgN5pUvIs6Q6DXozm9qD3Rppl8XVESpIxWhlBSuE+GCOuVALtChMlKhM+veOsMsI
BqsGRrupkfsd8wNAKptMmVQcvL/zQlWQTANZwTuuJFIbDEDM6t5vzJWvkA3cISpm
RApUpvv0C2j1WqyOo3sLPDoOIRCkdGi6S3h+U+jPwOVoAmaQiMBgk04lFep1OLhy
bkaSTUUjnq2vvWyyowWTn50jNTv4V1an8I935IN5QRfrAn5zSb3HXScu05LodJ0r
tL2mzsSJ6lKplP/CEhImUJVMkmXHKqHZSfQhU9A08XT5SjCzBMnbQW9tLU/LRehM
4Y79F/gGJZgYs8wy4a5iWcaGX17eGn9mFlJVUwS5/0ik7F0Q9gsTImfF2+NtXwYn
bm20+Xwf/rbn6CNmNJLv/ncnBdwQSoc7AQEpEwcvucjxlrkvTsZBid5w2RqPApYM
4NUIYbBdf0c8gRD+B6LGiSTs4BcbBtWXXpxlKfzUD5qSXU444HlhNYQZ+Gd2kM2G
MMpXAKyL5u8WahrA+bbViFD/CVtzSnnAolGTQn8E/Z5uFB+dTkCO2fzyB8oXZJG0
6OHF3Sdy/aYDjB10vKR9Ye+sHWIQZcpOLPF5WRng0KLo1q4+ayqkLz92YcRQpKzN
9E+YuPp2vwhKFOefJBc/MCvp24p3Vj8b5Ygj7apZyY2pkPFWnGdREM8FqDM6U+JQ
LZ+eivF1hG9z9AsuTZHobm8F6xbSamWHzNwbj9td48ODtOmaIEPNXGpZ5QyYoALX
GxSiLPsCpH12msYNgRBYuXh+UP4hVftLE4kYVMXMtx4W6Aw48Xj1nI6HCL0MKKOL
0B9asaXKF/lljtmCiPOn/cn15oD0ut1m0dGdKMiCVItps8BatSM1AUQEwwRpSn1v
f4RE3MFAa4zTAscgBb6wxwgZZxvqe7u7ix2Vv1DRmjm/y7y5cnsg8x8u60mmTk4p
wLjEMO6uQkzYUh9oPEdzTdim1dAXyd6Ingja4q+ZDAO51g0InwDwq9YsglsgqQKR
faxo0Pc/+kSInMbaJRkjeXUcwzDT7QyYjprBxOnD9V0yhfp8lbO8fzg0g8AGOnkj
ZK9dyT1OO+OpXxSzKkukXVOalLaaCrxrdIb/3Z4Zb6I6MHy9EZdEHPZlalbuRCfV
PTgdap038IkFcysoIpOo90kHnZaJK2vwg9WpmEZ02jlomLikMCcxbTwQGIeE6e2u
UtUAaj1Wy3NZGvJtUfrynQd3/H7SG9O+bNqGi5eBjtF9hvEQxK6bmhSgDFeIFfKE
Cbt797v9Gj765zxr2uEos4g8Q0NN3hvYibHx1NLv3/Tpiuhm7ENubvAcNME7Xcfw
yEcaZGhCjzJMwYYrijf9heEoi/tN69sBXfbsUtHpBKEaXjGIIzAm2y6+rrUwE25u
oBehKv6qILxLRs1guAnx44Vi63p1lT3fjJpJCUrkFLW/R+Bl9TS3scBpER3zc/6B
DhPSllI6hGnFxUHMJtjkHqAHl5+o4j9r7U/jTa0ThZSDDP3wpBvYXKNtHvtDCMWE
adygpxSnLaIHXHkcoqsmGAgoqhsIesSHxO+U8vm8Q0YBeHmvN2IrlSE7BGYqbLgz
JvpJkHKbk0yuErdN7E+FzGt2SviVoExhIiLFt9kXJ8H0rYy4fvpv0+6IJaxhT/7Q
swd3xuQ0tzwlOz4CsG10O274IRaOeP2zHrnDN8/DQBxfzlAMJW7Tkm1Ep4sMDVjY
r0ft7WGv198Uh+y3CdtIbp43MyCGQs+gkJOYzo8rJuXncmaFyaUq4i8VblZOFbs9
kdmmCx27SKTkfufZuUkzYkYZJh3uAb4zJ9x4NQVTHGWtXqzZCfuhau1owM0krVOX
oWdBbCnpC4OhHIQ04u+9xkAbbu9UKEFctZzP9YXz5YK9tMYPlqccWbqiCooGYFjk
DMuUOMgyH+VJFGDThoc0V2U3UPGPXoMFb8YSWvsgl6+v/HHV0w0gEVLRd+7ORumJ
1vWQA6iHFyX2Xz61o7ucRqysEoj+35LPJl39+wmvdSWCNIv4ke5AQgZETIonmPbZ
QrNCpCaJagep1CVcnjM547PYxOBz4r24JOy1dUnCwo7f1mXaURlbmwVhzupla9Ba
FGpznHrr33xUfYzpmjEgDSls8HVflcuOhHnZlsbpfkSgkKklda9uvD4mR7hc6Pzh
aqm8fUKQ86rNS6CAaFN+ttRTyFOp/NxEpk2Nr5v2/nMUjBIbJgQF/5HZnfAJBD9Q
OcgZrDLUkEj98qOvubfxJ3XoRHTtnFZcGnlU+kA7yNdnknu3w07ap/zcswtyNJeC
WjOq6+bDdZaZvElTS7L4HMwEeSnfrqUjfjJOGBiemE5tjE776/o+HX5A/drbdyzy
oT83jaSfS86hLDTlXlvP5vK7fNKSn7ODX5FXou/feVtqj6bGGMa69uuo0vYJhMRQ
upzcE5MDVl3O/cNBH6oQA8vBrCxgMJ2HJTjrvzKgmDMc1nTFhjS9JIL8I8OEAZen
kCFvxsSAqUpx8b3DBBQLEIB6K8NjltS1pGfXvt+zU6DR1814IC7FhDg2mM8m+TV1
dBctbBdCdmthFimUiKV9Ls57qoqKP7hKQdNi5tKxF+m4f8TzqmgiesOlXRlXslU8
l4CH/6y1waMMhV/A2SSVItXTpIGiDAZILpX4oIaprxvxzSak+OebvdiMoFlkrrFO
H73bbRdbXY4pQrv5Yjifbt9tFWoBt+NqPjPbxe1Ej+KRCt4+prnZr2L3vcjrM7hV
q0Rc3+xgqoZ9m/a+DXaqmglyUaIO33SWMpG51KyG8nEkxrxUxJRtl1k8cuZlWMtq
jke/KOsSO419qSn1N+vC2k+Rl1TesENJFzKJ8bt99um60qYqOHDJWea1k/4rK81k
f9KKNGqO/e2nEYn5MJYawpIAA004DWWcvMleh1n0ClrL1lNm5peOrhQSm10DU7rK
Vw7CXc+MtGX5STx7953PXvI+DmhF7FXGTgMnsQGrZWRTx1tJNS7TJfIlu0la6Wac
f++/1W0Ri5U1Shy9821zJEUJDFjsfo3X0bsLxTNHZRyNRHRemb3XRKujjS1RGy4t
L9XYO8RzUibOApW0HW8ukYgZ/79HnYfrMBst18Fpm5iaDzhIRP3tnoo8hChQ/izW
U8zCB7uHHa3IkEHnkxotH2fXHrV+pdSO7ZIr/ve4B3y4ODyvvOMnj24x9mebcu53
52sIR+T9JSZHXIkaeEWBpmZSHOEhrhaEUrXiDYXBK1fesAhRN+O/x99rBbJBk5dL
TpTvf50dPRRpcqtKphJboWV2+CQzC/mz6kILVP0IE+zkYMO7IhBN2QSsclaQIDPy
gQo2enn440xA+oJgMhrmqYDcghTCuCRN9Z4SpOGvlo+wzSQerUh3t83+okmUA/M8
mBpOM+suf5NuWHTeG8uKBMs1IAQSrRf/VhkHgh1pbA4c9JSFKu1wvVSFht4/4+Xy
hkmzxtX0VVrr49OdaDPc7+MokfXWLUWx2W3KC9+n/y5Kel48adw519PA3PBw2uOA
IdnpGFDHxT/M20kuThciLlgCwcrSpjY1l0gYEwZQYaG9mn08kV2bdZXndT9E1uVO
tSf92GeX0EGRRRMYWEyTj1Y454XSy+vIarG7WdEeV5E17cSPcP+5DySyq84uwUJB
xsJXQIRE2cPC60Amp1u7jxtW015eff3WN+F0tbg8Y9zDXSAlyhIbYW0T6TYfBWbd
dDlxftruYw8zUvJFdTI9lYbt0ju5bIYHC9g+tqwc8PQD315ivzl8bDAzddx7PX5J
tmNYp+dEG3vbHQ2L1anUk/sCWVKfahpLLTdU4phMez1I6uG/vO01ZfHUldthw0Ck
FBUCzploEMSSe/6irxCH2OpVU85NLviGQhkRJWrwGdvec0SppxhWNmZIN+Bdk1OE
VKIEggjJun9Mho6BHbG59vlC5G0uTNANW1jZw90nINvl96LapppDZsNQ0WKmBCG2
zWKS5C5S3lYQpUMjigFXUxJdE3Nr9LSyN1XTApqiN5FZvs7CEwRZHGRY9KFPob+R
oJPNPFsyXt+/TATz01uazq3RAcTvuL6ryNSt8l7upE63PtEMjUP91ZrwfHz9GLhU
0b4RU/i6yqdFqgH6WqN3a4YhnnBQ79bQ3srGAWozPIBtJiYIN6/CfuwWcPS8DzqR
QahmPU1iiNiGpnXKbvK4mkrsWuAa/9fb8RrFNxQOwUNh9uKh4f0J5c38kayaxQkX
BP5Y+lLgnIsY5GsKQERufsX3B/18jbbuxhvb7Qyr6SQ7fvT2TMzl3/6OCyihdOfW
wqaCHgsEh7dESMT3PqYlQIXBHPDo9qYlGPz/6bReji9+yLvJWBNS/DVRvT1ZSGnA
CPnW6R5DoOs90WBZA3rRTQAOJxDmCChFIcErQZUDfQmLORXyt+Ymot8B/cDNB7qG
/zuZN4uy5wrZ3khdItRF6ZjMdPHuSI35unFKAd0bVCyOIC6ZreVt8kQFD2GVcyL1
DvxXbxTc4F22Gc5y8a1HRaLHnXfO3D2M6GHzqCDSMA/q0GgbxZKae//joPOX1uB3
cy6tIcNGCmNHwGRT80uh9Vm5VqF8c0T8ksyqYeF54Qui8WKmIAJbGtXdyp4hrzXs
Zp2cAuJ1QAfDZ7djtk0uh/W3vMrFcJ6Cvg6VhoJnhnmFoLep1t6BhZsLzkrxm/P4
Z9bntZkWwe+Gk+mKb5fwGMtnqqTDTzoKRhH61FH/g19HoR/a84vYzVieCdUznaQ4
z+B4az3b3/Yi3douWursnNE2c/mqfsyVeMV1HFe50CiRYee40YvPttWpXm595oDo
JSnoMCMr1WKI2hgZR38ujhlFfsO7BJydO1qHL9Ol7sryDL6FaCEbxuMKLaZoheFJ
JaCWM6/pSzUHyeXzQeJZlVMxqqwAn1OjZLfWLlFwzTF3Mos31noFo71i8dhAe0Je
fdeL7Fj+bBnGjEw1uvli79iy5vm0KulV44zrqnI/32FSahz4KaUHnGvIK/5hlXea
MIZ7RXBmh2VYpP7kvKi1WZlRs0+mbimpes7D2XZAurrC7LEN6jdV9X4njlecOdZT
m7CEkcWVIjLmZ7N6L2hDJ2unITgJvqwbyCvSoALjeSj9n7E4Oc2srbcKpL/R9imD
1rBC12z3LAZ2gPufMzvEUSlmTiIdsoaDaTUsI3Mg851qOlcmG3CQZHTgGakTL7dJ
5xmi4UxqKlwx8GoIueXpxsXzaKrm4u+YkQdgILByHmOVDyRjHMBuzz5R6xGh1xc1
/uMy36JJKVq8L3lRQo8B4KLHWgMtB5cZuSjaByPBy0U4fOzjjnqF5FlEp8ylJHuF
TU6LD/+yxvJBZHKrJLoOdPLIKeWhvb7NzwFfWbiGxxmiFAPb12BjGfcAARa4QZ49
0rDm/c5CxodJcjdkMh+ixxHjHMd5BWOREtqucHwB402US2EEptUrCXl5yc5ujS1H
DT5a62SWTduObm72837TLOZiPZuGYC/kNIJznNpHmOKR38ogd7o2F4fiGMdzlDwc
ky3Eg0x/ZTRr9AG1U+BtS75MEPidyithmmWqWrnJheurJtnfyVrwriI436I5WBVF
9hs59b7FM3npV9KnfDV91qQjhh2ibcoiYzxlrK1RI8ouKWJEA5rtcCde6UR9D6Jh
418xMPkAit1lyMdTI74LYqwuaGeVxvKFJa2POUVpHZfD7T67hvm2oniZCHrneVsr
ikn8sQUbwcU6X9un3/nkqNLAreVkBifsw+oCcSTJXVitXzk9AGAdDpCAvppNr5eG
bHRzszMKBgMk7ghe9zQeY59KoZLH+nkipF8+JjBxo8eP6BZAmGV0y7UAa1eoKIt1
z/TAGeuezPX/2GZetYJdDiUjM7hC5FOzzIwwCgjd/arb2G8h43VhPO0l9M2KW+vI
o1nrXklqWkcfn/7OxW3DbNM0/sL2D6kftqCxLKWoSqPRh6D7XyD9dgteeFIBSczZ
S+6UOJRzTR0E89Wd8Osi/A4kvSKdtzsiDbG1I5GqKhNb4nppCTd0o/rpd8CbzsyL
SOR3CmS19MCMHbPpZnjeq0YYJ+qZEEi1nAQ7roY4RPv3QmFlZTLYVIwRgCpeybAe
3Qtz1QDywHLRddvpgCSxJKk7ZUZeG/VrByF21rkCdMZOWyehGkmYq+DYcwZJp9Ra
H49YV6bBdDjsc6xSFK+BiOMxeWIJQJAQyBeC84RscRAl2LtV1ewSIVs+jSzGttMi
+AQbhSa9ERdlgfUTwlJBTXVfVjv5h3nxJI5IpXpZnlj1vNjVU7HIsUQyjBWwzSoL
ytdWqjZKle8c5Mg5vyIORTrZggeQWdme2T7CdDJzG6s/VZP5oCwTR/kgXYn/Ij0V
Elv1F43pRDvuB2AibRg80vxW4w57Jmv3O4+jaK6DWDxQZJGe80WUY4De6sZj63ZN
bmiFFfgAqwo5IUJyYQVligM1kYFyXF/vFcMv2sxgG1FOpGlZTt8izxBikkqByEg+
J8NN6Vlc3bDEvBMCPZF2KT34tQBIbTdpWrw9bslDNQisjUeqwlzwgA30VrWQpeLc
n3+ijKKCT81jocuHqFsZlbvgKjKyLob6s8x+5pjjyzGBvCmL5qW42Z9QvYfs58/J
rYrsHKgzAJvmUjjbNsiIKIRnDIDPypM29SKYuvRljaZt8ygmuRkkDE2zUtOBpV0X
5QTRThxQwRKX2NCs1ZkZ2PYBa6cG9Qm/olCCZOv92luXyQMJliHLv1P0+9Fj8liy
GU8eeJII+Cy0dh8RM8eoLodcaFgUYsSuErmASV4OTwp3KlAy1NhcNarnJ7bQlqSy
a6q+8swh/lKgdy8eeDvweacUDCmtsJNFVZztL8BrMdDGxaYv6ptrvNhCJgbH97VW
LD3eT7ILm26xb9a/ncJyCl21bkyZaHkvYq1Uj0JpzB367BYLG4T3yj6FKeUY8Q0Y
aQHIbmoQGRrwF9r46qsTzHx4SCY6JW+AYLUjBEQ8Lv6s0HI2CCPF4iZWagXhKbIc
PT7qt5aUSXswurLAs1/K0xfSaQXYmegNes910XsERxSmvNr2RR6z0XQyW7sYkpLf
dB3uzAEqHxhY9L55lKhw0YeNAwQFhh2cQqAQkYYzwwHDVV61Deh7NJ4VthPef53b
eW4SbhVSOyxdhiW0spDaG6zrTZjQDjOaxYXmTDGYuFrpYToSXpOezzEFugoHCJLN
deBQtn/FydN6jR5HjyGuTztQBMJja4x3h8HUl/Ut5yinW+maUtTkylXbRZtRuZx/
s+Y5IerYEsyZyLCNrK8XeUfZaE2uzlAWBH3WzmmfQAlfB9uAFEvZEZAWkzq5K8PO
P3DUMFXfVRhvcVD4Th84aeuRdn2YQH73ieOMneiTYt7v8/ps4vLS5IzN2/AFF2Qc
TJtQkCfSvLEBHCaH1xQElGB/RsZR9/QeXtXvN7ntFO/CwFS1RHNEvRehLKQYEuBI
DE8mf+cn+idURkiZt35UsS58WUHhBDyBfQ7Qm9s6Xtxcqg2vuiIa9WzKWRvGtC4B
EuU+jfNVKKOV5sRKJNXpRCDcxqUqw4AifDmU+zcJsPoybv7UqDZ2LVGK7B0StYMG
3YIk48rZSrmwUJLe3Dt8YOMf2uiS7rlx+EyrahXF8oXjLbDhbTsSP2dHb+18suYo
gECgzck0WLlfyLidW932b57uhGClgpvbzsqs123s4IBFXBTWzo3BecyEi09Q9tA2
6kT/HtGmMoAT1zzUYhxJlVXQVsQbjkmbVSYYsVoGI56SrSadVYpqAyka9H6LNUya
DQCChOmoQHtZ99QlHe6wX4VFWTmiFAz97ZLgduM5QSvSauESREl0rYykzuAd2Od7
sADKHDW0loJr1Nonrs20bFyq45y7rpY0N5UbDrn+9hpisCEa9F26vX8goZccg5Xj
OK1+1V7DrmKdHRPqMGxLzWDUgNlRrBvzTW8ORL8Mu96wgGOou53FoW6h9caaf/Jr
RAfq9QGehHtt7sEhQsQeIk1LEZ5omMWqLI7cpF+FSmkte93oDyIk6oSCpTflIh0H
ZcLICSYV2ir7c4mIc7RQf9h4gWwWHVfP14WmwelW8kUAnEDszcNWgSSMlYFLZcRb
3e9qtgZZSfM+vz0rkkuMIk8GI6s8Qiy/b5BLR/sxTq+sZ4yQGSbH3QgMTt7kIqUR
LBE2vVsAtj95qeS1wSYkDQP/u4jKNxUoVrzQaNuq+/UPjwlBcy693BxN3hN3ghyt
5lahvSTraCPW1zxM4lAc8lRrNKCyQYD6YqbGOo7bha3Iv404uBLl83NY+EIRzwK1
gtv56Yx8T4HbOj9/RCjcdSIxVhgbcGRrRUP3NOy8dTLD4t3e2mKwnLC+Dkug1gSE
0hgU2uc57Dukp5fb/AtizT6dChPyHlVtdYs/AkFaoxXx8eNI7IwO1zF/+Na1n904
rqjFWmMpmvcjUzj60RZ1AG4zjW6Fub8lYubpzPfu9SKKM6PPb9RHEDnJ1KvJPkiY
/+GVpYn2RqygNDXjHHiXNiyBg7BmkpTvPRvJg9Fg2WHX3T4mrHHl5v3DhBFcOR5w
xZFv9z3mX/dMBZVnREoq4N1EITkZzx2UYWE3KzixlYW2GWoxnJZZxCs8N1oi/sfX
qyGIdB9ygn1Y5nhTIgvkNCJnLb+yYqiGpFyG5MK8k2z9cm0mtNp6bey+px3o0s3p
RNRiYKfnF99mBi7RtWguGk8Ni2aOwPp/h4PQjcc5FnnOLOX/CfpWGuFtsb+ZbYad
ECfSv8yMP7tHtKcJfg0QhOb7cekouaTS3gGcnzwyRk5N/cyu5faj+mjiFLLPoBcU
X3carTyqdp6dpXfYbbjUkMjGL2XTq//XKeWXzyYUs3YqGeplX6Ai7+okSUysJuGD
JirxSozJt5UlCX5G2B/lGPoI5qhXNwSUkPDMOyN1LclFZJPiahLx5w/98FMLtztO
9kydLgxXbi8MY3cRG819eQOJSHh/6NimRHLmN++yNa8EaaOcxN+mCfw4xEflquBn
2mbYx+hlfjzf7JEYnTa29bJXQepNZz9vocpTeuw78WIy/KZxCF6P6yOYST3CNgmR
6Hkuz2CT6sxZr7Q9jJEl7xoIOYBEdvp4mBE85eaRe5LW0fFXjJmflwN3T4UP66S2
5mI7Zjy8iQDkEQkdBjEpGxPATVzBfaZexvCqVXaEEU2YG90sjmfsEG8qPQtdjC61
1rexUnE/u5USQld9kRoDM3lh1tPSWMw9kWYYJmBJphobfvsgmUASBMzh94IM+ET4
AgwwmMFyGrykm7sJKGvcA6b6RQCgos0s6OI1y4rzxFHlwLfaOEhIj3SO/zVOZAXm
z/RUvJNpNXra5/aQpTNNkrRNQJmjhl1aTACrLhMTOf6KSqI8pbhyZHCwyGZlWpyt
tXPhpvohJV5wMDJs/erSpwW7pVoZ2l+2c9WfLg19urACGk99+jax4NaZ/x/3Hi96
O/25PkHPIfHYsbJKpEFh46zpxXQ5p2X51CFRTRPZgB30k+LfZFpzMpZuPcbwl/6y
+ZcF6FIdgJedfo3RRgIbgpHARHtLXzktKuE7eunN1IRL0cNMZSvgcOkoTnBbyaSV
gz0Qdtr6uBEGSc/QOkaX8A2sEdq3SywUJ2WqrqoAAQTUcA6nBVaOQ7cbcXJKjrwn
2hsm4DFj4EMg7C97ZawbLtDdNiMljuWC5Uw0f6ujizHtpuxq2IfikYQTWJjN27qa
4GFim0a6nHmloUXcBK9NGHy7gUpOHLjA+3t6Ft66zSFIqnYFr77guCG4EBoLs5Ev
UolID8UdAPU6a4lbQk1Ah9RXjETqY9eReinez2c4PvdnzkzwPYb0kchxv0+7oPe+
NXoAwgi8uSwxjBalJoX17x7YqXEiIeQnL+VpxLFKpixl3qrYrYpOIp0ZTlfr42nd
u2jyRlA8YmzCiZnYvOHhmUXzbH4HrfJfhemH+62KVOdjI/cKMGIfQXnSdxSJk/cY
9MgMbXeTSXP15Dl6dKbsffTw7b4W/pyFvBDw6hFT8u2mY7CMZzzV/0WFCDz3VMFg
SSKYi8jQC/qg8nn7k0RXayCmIHvTv76WENBPVeNUf2mXEfPjwQzoL6jtxq7vWeMc
8FZuTGOEVnjUCj8yjLPI39cMCSscmO8BzCRixDzCTjfvSn0D1Hnm+uw2WBoYKQkl
3BpULXNptbRVWnLeTrIK/dtWmBXs3sv8rfRkwuhRTb6kGspoVmF6Vk7qnA35CmZZ
nnv14JlOupqilxMv0it6wIi3vfSK7rB5jeA0IUgXQF4R7y4PEkBBLLiuFBn7ZXu8
2Qclt2wppxPIqATIVVmHTmBZ4Rvaz+kBwGbBbOudzNBTA5xRWKvX9QD/TUXH0x6r
Cnn00/d6buK4zBEQUUx34qAisiyD2q03BSsnwdl9/2cD+HZcqgEG/+DVTbwpZ9RK
cJQeIAN9Ws7DBV1cu8AVAdUnsyQfgeAzszTXRMsn6NRUlZHmJct3Snhzeg1s/7/A
nwdXrvGy+JoCD9TnecXjFpYY8vxJ1Di5XqSEclOoYdtk5WPjwOdw9lGIqHS9aTI5
2SKmJ5I9dGuJQQ/jr1a3YARvtcsnnzWzZY0+MV35YDaVYnto6UQx90mcQkpX2SNn
P7cxEQwI+gbYf9jpEgI5pcvdQ5VAfB8WH/o2gOk9Nqn//yIGwdpEblKzThquUcRg
UGtqoNtnWfWR6qJGyfbo5bZBFVGlSMfGHQZdhy34QuJS3c1a9HA728DweXjMjK34
DPF5i6unT229DbcxeDRpjB+TmoqRQoLMDlNVWG99R429vUPrhNT6kUiWASvU55it
l0xty45Io8u6XbubG9nPrq/zh2p5KfAkE7QTnNrgvyh+WF+nZR+fGSK5USZkczf5
boNW0MAq1bORx5KezeLyuV3DzpGHVTzN7LzzU2l+waNM0KdjZMVjv64GdSeImy/p
6yZnWKnEuXPfJ5jws7nJkiekGaFABE7ibamH2cbKi+iNW1/pTwq0+PENHqhrngbg
N9FWhYeUjS+tRJR2n04ke543+xSM39CYJiWlU1sI2hGHjdHp+QRz01/sLjSvnRqb
WLAbIDruXoB0Y81dgPjQgruidf90WKM5rbDJ1iok3TQyrwqzgA8MyRxYvFNR4o8H
9eDZ2rKZAbmpMB5EMtb6srqRMYE8CQHISPrRUK52an+vQ3F8gYot1ymdwbGkls6n
PzwWkSQ/aeA7xXOc9n7X+mlL97DEoediZXM1cftELAygEFEQMnTfDjumyzFrBpYu
0jRB4qgxoE5xPjJbaqsY6wmL5ix0ouCMaLOMUYvutS/s6XiO+TvtoJZB9AlDm1ga
7HIrPadDnZRv9qpbHFrujHqacc5VszRDo4OZrOlHiWuiXPYCgIbPlSVtZ08lW4b3
GeXOMIVMma3q6Q+5IYWGV71YBiN5RumIUe/530y2fzlDDeYr41XTw5e3Uosj/sbX
AkURkVp7gDMxL9IjVBr1Dam2PAEk74CACra2EFG9FjHrO3Bu35mHcdUHlaaZ/e6/
XABqHQRlcD6B692qnDxWBWCjO/auz/U6PvAuXAK7kzGdT8iw3DD3iThwOGNjTa34
P1OEj3kIKiP9k2napiiSEbYXFfMLzTW1KlacP+6OkgXmFE90CD5DWJKe2mSRQzzY
ZeZqdshQxHu1PZDrTN7setXQ4xHYGxZEwwOTEjfsT8itbh/cz3ytUfowfg11ePJY
BSOH+fx4XdQHnWTRci1d7z1GjKepjiVzJ/N8M87UmKFETg90w6Y85Aer3dfDFHdC
byyE3nctrC3/gmDzzUPN9cRVXHQ/VEnFLNcDAb7h8eP3zT2afUuaxwhdnB1gJh/B
DvSoDz+ruxfB521I6bq++uBW5yIteUoKgHv1FBW1MvxDGLjL6AO65QYyzAJ0YT9u
OlhDK4u4gT78hBggry5dMdKe5of6W63cX0GgF+4L9s9cpJacjL14Hdr0+Zuv8xIS
xaglQFJygXDVNkXxqBJCHNwRyaUgW2gJVQDpTqTrLzAzAID1oTrfED3imkF5fTQR
jvuZG2ZwWjFo2Is1uYKA4TYk79CJGnRcGbfuc0AqMvJkD9no3V1YqaWUR8/IqtRo
s/SoTYuQLwvTVTb6dWTBd/ZIOL5l8UQMh9Vgh7dlFZwm33My2WN54UEwF6HPS1EV
GEKXAnjPjBgNbf+8aiXjg+56Em0uGGP0Z08VMQNuRWX4yS8SwkEznj5JJ54tiETV
s81Vwu65NhsNujNXuCB4tlNpPD0QWKZ4jIxQkK9eSz0Htk68jolCDMv+8SKY1FSV
LEfrQ0ui5xRPK8SG8m2swFOc8pOjvYopE0lddHNWIqPW6Wlu7B69qWje9vgtxqTb
/EOz6ARQMMbSapm+81IgKkoMV59Tcd8byiYulsj+mgBzZOrS68sniB3OMeAynO91
MNU0SWJKRpRpv85XEm1znDOekTSWU1TNzI+kiNVfHH0oOE4GLyvqdw2K358bcGa5
JlWI4JdiR4tW7D7+5tGaaD2VH7ztNO8bXANGy26OmB0Ueng7Q0VSFWAsDoGE/zk8
V5j11GiHAHTIXEMFvGzUA3ydHU7a/k3xBbFtEepG+kbAHVJ/vaRIcSjTRpOPb38X
LkZe7VsA94KHivqYIe35t/lTr0yGaQhJ4lSN6HqSqYN4ia7ihe1vjE51m9eFm8u/
HKBcYLdM5d4yjF4RfPi4N6A09pyalz4xGd/APcc0xvkS1p4HkSKS5g/h9CUGzRkD
cr6LF91Bo4niTp6W8apF9zIiy8MUArwfvxbwsrgg/pPbb0uu+p/gA9ToKD6+GSUs
J+zQWAc4+VmoiAEOMhp7HSD03O563GAvFmydLFQkpFQjuuNUYmrJtPW76RBmFZl0
7stNJ85V12Cf4gERRjtmJs4YOjAixVL5MwHpOR7Ih6ubYlPT6riywcqdLhhmgbvI
4KJ/2OQziibdZOxmwr5oBW14BL3EKnUn0WgsfOMjWa4gZRstTuZ/o/dK39suzVH2
0o9C7OSt/THmRt8KSg84PEDCpCZh0d+SHPgmrWjlUDRsBAqqCwyaqiCuV/nlpGMp
RSwEmTB2LfoW5Z9zVY08ySKfZ32kJ/0yQwH+0L0z9veB4trbA2DKxb0kL03zaW25
ZPKl/ohrPlqZS90T82SX1AVJD7S6xWCHeCfCyMXu/xLixf/NvYIfWPKedWdGqzhN
ikYMVX7DA4ew0R56Zg3UJEio8g+/d+PTRZo2UZfreEDvASDVVtK5wjtKWn7u3etS
9D2CWrDDmyOfhv98eOtjy08PbqmkaAT2xT+QdeZ1ncPi01Ga7S3NE/gJnL3Nv5VN
x3/PclSnsOgiVRkHmU2+ULv/mxTv46txysznfwvuDg8gQDrt//GbUDem9j0pD/vj
aq5fhVOrF0W/icQ7wuL2+618ZwNbURrbz9L6hsGSDWomEZJltQafZVCj5uyAxjsi
k8p1WQF1OgWD2YBjxOGsoNuyYgbW4YRvCl5kJiZKLYTzCBgZtRky2I1YYjRKUwyL
thugELif2HZOdv+CfOQxcemXXozTExTUrgebZRtB2m45+/NtacsVninqJlbQAImf
xtjCmn9QQPE22RpK0yI838JjUsDWtLaNxX26mo/j8jMuVV6ugOyWSY7qMXASXKEY
qRTIDDpv7zCp6cllWmjsu30zaQInT+zA0oAo814NPqycENTGe6f8tl5eAc7pfu3L
DluswEsMHDV8sBUL8Q33MvK0yc/s1gp6bIuP+dugFm4h8q/67u1+W0S1+s5M+Z8U
MIOA6NdZ8dq2xkQiEirFhoFZLnw6YhawpJjUja2lqz26aW2b0lPQAvqNYqNF2rp2
xvOBth0R8t4b+F82plMhvakMfXgEFpMcWyeACXrGxGK5Zw70kbvNQ1qD1xFhqFkp
MiDfGhjHdMbUdjrKPglie7dL98TLPy0zuDXWaLwwhTFyBkG+nXXol/V3VYyAY8gw
3E2jEfS/Nn/ho4Nom+11c1htMvWPbJvBtwwvKMjWPcAOZa/K7SLtP5Q09oHRwYM+
y1DCRoadIx6KNQNDvjttY19BX79NuqB7KeJlrGClxW3LcDktqvLb6Q1gX8+NjP9u
2MJcc/vgcho6bE+A4TRM/rT3u09PhfVkks27FdR3Eizo0I3M4oa/6yHfLQQru2o3
8MIB6zKCA0sULo0KK3ax9YceGjHxDY3npvB8983FPfufs/A0G8zCBx7NVhQ5LYsm
iGRQnJqApGR6QkYqaBr9Q4BXcqtz+Zk6Ffrv/auXCwjynHm4e1Yj/8L9RZ611szR
WsMs5q4dgxy3z+xxKL8nG/Vsj3EhW3BWsQhCL6rqe2UFZ8JKe4tGGKl2dFBRweHy
pVqPwLLDZZnDFlGGd5BQMeO55lyOEXfTOQ1p1Fx3swGXbDp0YIqxZIfkotZaDXjp
gEqutjCPjmvQQ24yXyIv05uFBRCyTGo0wQHRE2rPuQlQLpHW+xXAO6F6yBu9fLlY
8NNGPyFKC0CjOJGIrpw6cz2z1AQgchFA9G3CCIGxmKGyxvNymisbu0g10bYRdq69
sy98lJH/FZ79uqw4rerqZZOe29vgRTkwvoQfNMFFyHeD9JjZ0KLwLV/jMvRFmZNh
UNQbZJj3gAAjs90h34RHmyMPLcLdeFl7HZbDdc/UVYCF6CvlUi6YBBah5iI5Kzyv
gEDhzXTEdoycvPUugKgNQ0XR0njvoPI48zSe1VlkvjCeWLEind0SR/tnY/+TWBbR
8LIjO392+ND7QOYei1OFA8Igc8oNaFgdEaNlu+L2Z5GmhE/byvi7rpQ22sTkPwBT
VMn3D5ctFQycGXd1ZiX2V/8+XbkiikyN7Z9iFdbchFs8N2+txFsCY9vbkugVuvJU
+YssONNLf9JD0wdYuQ4asvF+ZzgCCaHch05e2kESh6SWs5Z+rt3mFgv6rGHxdLYG
du5Nwest7gAWDk0d5X0vu4r5EF6Tgc3p27o8j1Df+jeYdgu5TzTWDB/xtdxerzwN
b92rQmvTsYZ2qXKwjxoZiLOZuzE3QdSGXrfknXL82MPmIqjJ8szo4GXBxdLhlNxL
v5+u3drFYdJ0VUysx4KAZoLSEbl0OPUJ+wG7FLbLotHxxBnBd1lVBTjkyJo7cU7C
iCup1sxKFw388d/kBPbRkiY64VJsMTlQ1ulAimneZ+78LPfsXs9b3aX//7gQ1C/E
9MLawlieISQHjo2ftRCZKbsPRkoEyKCl4AECO9ElsSl2K/j7mNxYze1tsNx35Ry+
ZcF9slg5iWplWiAW372Re1OjKsY153fQ7x4nX3rmuj7v7gAAG1wRvZMD9/jSCT/x
9Tw6ezWhxahaJwnYVcWvHW9JkW1KtwjrSV8T4oxctWSTHnYuSa68niZXbj7MtwOP
5ADCU6etj9lVQ5NjZJlXgnFHaqRBFKDPlfBozKBfApcpzPn5kZLyYDf3rRfqXL+T
YX2qgw53Q7fGcLjogCOhFDjfh85HaoUHN6/J6W8NJYgnEeqTK0KkCBGNQ6VEx150
1Kuq1ij6RA0ZxqH9w/hv1xYraZ23wmJ3sS9tjrv/KxMY2OM4TXGwYr1CJQOFRZHq
M5XXHb9FehorDWdbeU2P4udWPESbxSvJFLWregOs5oczj6oKKhz9BM/89RrW+Wz8
V+6L2+M1V7b26GOElkGAp8Hrgl1yMchIZzrVQ8Ii39EQ6EwnOlf8hr+zYOLqV1Bl
4r+WRov7OOo9ijCiLbY+gBNCTUmCL8S3dQDbfOABdOL0p4u1bVtBQaE5y3YH9reR
EfdYaBBZunepUNi519cNjNVrKObNHemWHvkjFpoo9l2pez3MiZJT2+/8EmOCgzaQ
EuRcul9DGCPguyvkr3WiEniELeWq9lEXgXwoo7jXnTPebjrUy5jvs+FU270dR9tX
vY3X4sZkHAtz6rd8UAVvh00RA6FJWByCcri9g39Vycmu01rsfNB4xUZjj27/UAAi
L/4sAc0KgjhJ1COiEkKOoEoULitaGUv69MgpWJHWpMd8CEwKff2yJeeBR10CD3VU
qPzcHMaD7rGh8mtx5sxAd91bRwbj7+4sZB0TBhbmUVbiI5diP9d+1pc3OMf90W7o
xZ/WB40S9e3hR1zOMxERL0ODq9gzRRAVYnIsXOe8WCe4T9vMOFF/oE+bQWII1YdP
3xuQDgI+ZblKYdn5WX+5yHcpgnNlsXN5QPeKVcoYpY7K/KLol7kx4+ruYaGeiDlH
qlf+HNxlRLHSeIDGMYvs6XH7IuNoVGB1RWzpSFcVUECZFnVflTuIC5BIBPyGcP2E
HoDitHHb7RtEp8wX67ydz9fDA2ZaIk+D5VdVLyO45dDCHm98MvSCvY6vIlYtcQJj
ePrthqstQOdjwTYqgLRD9yep85XooFvY8+mRoGRpK2R5okDGhpsLSNIsH92gNj75
AxjMO+MtmIpF/yadYzGduZj+UTl/xo61siVHzcArIHdegZ267RKCPrdwnVl7jyk9
vMiIkHaQBv7oQSxCfMDdn4TknRe1d3fVLpoKQy/nmkys2kGQIk0PIImWRprlt6oI
BTV12jygq4I6BTys+Z5aiggAZJ3IYc9Er6oEgfUhjUhWDsNUOhnht8aDzsfvHvPM
E9gmxm6YB7GsxBiguJPD+x9QdYZ5ZEyMJIHn3TJsZWxX1VeHlGgF6Iehj5s3zYGf
qe3WjMkH4JwrhL9DnFifaE+IV46X2h2YNIaYBEb1TWrePOasAl7ARo0JrWZ0xmjQ
QCblRd+Hp7c8tY3ZO0rLZMcwtjV6bIfV/jx/vyjzed50q9M9Oq9DHZTPn8+Na/Rd
dhPEn98Pwf6xWhWKfxWRqMz2Bd7DteIzb1+62fj0niCxa7Xq8GtvQCJtW2NFp8Fu
79/5idmPH+qufyZgzFkQDRAl0YeBZCNStbVzo+CuPrjGWnVr+ohCrkK/D0TbCs0L
qn9GuBz5F3rFxyrKZlr66vndgPlqT6y6VE5J9xJeP032HvsxGz5uwCo7eS9VmzUq
f7IDGh3GIhEkjNvT/LUzyDYs+8YXdXLLj7oeHqW5f2SSiAfU1t0gpF2ckRhxi/uE
OkBNHKBkcdBYDWT/hWDhlh8BSovNrjeyisUjB76LrEchkkXp47ejq+Vc774YqUPG
cmAmm/26qd6+/AzWU/kNC9urPOwtmQ67d37aY1mr4iKep69tgGks28ma5NWigAjL
OWUyixRMxWtah+RQTvSUFq3lKV2/E1Lfvh143LRrSfJlHiTEv9BNVYwYAuHdVn60
vmLhpCWkiJXUcNXGc4gN1g3Pu9oxZYAieqtq5p/gO/ySANbb50ux55YFmzx+4zJl
KAqiIX2TL4LLIreoBcyoDMABdlQ/QsGcaD/XjEQXGEqtJOTwJbKo/beG7+uCI9Wt
17a+4gKsoAYqepPT+vzoNLiZpIn6Y9WRCSFhCr2sf3WOgPToXnIi3g6WtDSQyjx5
FHj7fHm/0SIcM1uXvidjpmM3vCkoaI5Ha2hcefyprwdKWG+A2MzOo7oj2VMHKFa9
2i3DHQ75jUrqx++BVeVYN7C8CU/kfEpp1exXq9Za5/IqKACxYELss/KrBcdSLdGq
/tdlG7U6YCdoNrkO4RVtwjPmk4jfps66xkGiHUekQ/XlOlo2IQxOhoPNMo8gm3l/
OBEgflo7JvSdw+VPwqiz3LGG/HQlP7A+vqP+2TLab22E2t4DYqJcAqCMHARHXuc2
0js6jBsY3Z52FZsax3xe2GA3MNSOCV4iVj6LIHD7jqJkNpR0jtHFvSrxTxiezo7R
ShkZ+Ky07JPDTMGR3se7o2820RW+CpcT+SzZ8qYgm+9CcZUxE39EiAqbiJWmObVX
J4ZiWLgJ1KynRyFMiOdUxIjFmAqeS9M563XyrEJHuByNPsGCsWlAve932KAwNSVZ
GGEFiPKtnijXW5oqJm6NdL616Yfo28VsHr90yi8zdsdzhzAL8K4iEwtOqoARE+NO
8/HwtyAq4lakHhHYPVIme2RJaUXKLikgdJU+sx1q/FUoHU295MQCYP/jtbuKSm42
atvNdTceM6rcNmoJO24Dp0ATKNlyc9iJst9SJyoxz58AXmR4po/GFkIQVGjNiWPF
eDPs/S3FqrLJh2uhj2xkdR43jRswJCF4ozZCLzscmU+U/CWziK0zORhnw/FUfXAm
C3vzcHZ5zw05fAMDcXR9rxrxlLTgjpHtFcKgUSmGmcFEiN8UDCJ7n5aAuPqscXIS
4nPmAVoCUsmLrIiBWd16drVBEpiVZ9chQhFcENxrjQPdb2MLKywwTBSJ9ffQ3ljr
NG7HZJHUVH+pk4nqjR5FyBTqkYjLW856FqEfWFNIKQXYcc/oGzvzpvE1/nN7ZtcA
eUORXILAz2t6U7WykbrS9vCLJUiJbOMtDAqx1M9iUVqM56Faq859tnddWcdReZ/A
8oN/ifIBHmi+1/zrwKrFgD7xMCL1y8VQXCWl1J7slW5TndOxz5+xemPZ/RGaKL2e
Mqr/PoX8PJcxHtgSin7CJL9NPXFn4jspzfwphbXDNDmaPj+n+D03EmAhApQlpuCJ
6E+dGFzfO7Wo31MKqZqZZFm4f/xlDD+Jaw5LJen9qtYWYacmbnhP2blyKJktHnXv
bJlczjf/h74nte5hpOrwqEQM8rEC9U/Dvpf5yNMkWaur3HoLxNB7CQdDJg6sCtbu
Z8CfixuZnB/0BpfjhE2fZx+ceLM6/Le/9xWZHf3pic7gfQmrMzT4J4pVyZPPE2D/
lmmJEKzDk6hGZV4GshS929+fzVnLLeh/WMu4eeqRu54rOQySiuGUjzGWYVtHYTqf
g4Za7CuZeVY+WW47acIEdMrFBeatClb4YGYyxqHVMo0jOdE/WGAY3gfyyKiHDUn4
pw7nEEImZmncrCzlYsHbyul7bpXkVq9BxoamKGCpSmAQ9sjgtRsDltqzlfI8mTTJ
sckGAV9iQ0mXzLbxoCL03XF8dHrPgYgrRqCkyPModtwHi3Vm3o4M8diJt7wMU5z3
/WQAzhiD9mc85D/I0UsoLVPkN3GU17bg5eza8N3aYC8/KPN6phQkN8vYSqqSni2a
1WaR9u+3ZiqA6tH6WS8jKozqz0ca1f14WOZxCwlqn5XvPIi5MQzfkgxwSda7rk+H
FRwPYe1ohZ5MjDXBPF9KLkOP58ynZCjD5A6O8wG7zbcAEF9+CJcryaXCL6HFscAA
8hIWxmQ/9zlEaTsO8WXrYuVEoGhDF3yU/JsMl9LOLi6p5sg30/BAwO3ON1eMHWtD
o6sjBoyQi1eHgXTX7F8ZEo3NAhkzJL7rsOhNG9DU6BNGI0klDMIgdtMzwmCgOR4d
5fUyXh2l9QSYUgvKbt9hIHI5XOFBcJIO9rnKJYuu6tI+CfZtEXNgQGq0BM1yAca9
Bleko7RYY0RWsB9xnoTTXOwJxDIe/06IbFiYlzH2HYOtLMA1ci+oo+MvQhIznoOr
jo0bN0nfIP1bA934tNRTscoMJeofY+mJAGcRhTLN2J2kk+BJsxJepcLhoQzlxIXh
G7bQrzzAxsLtv5+lG9VAueY9Ty15mQopomzEQ2XZwPuLeRwuLIy0w+o+PgSl8Ji3
1thekuODvOHkgwP5o15JlSyKEc6N4smLLHUKiHdL0hbbLgLqpnquSikIef6wxQJJ
VlZhO4NCxmRd/tL+e5e6lEkpLi8c6YVbwIy7yPFkJF75KFAS9imwtyeBNDd+VMfA
6Uz8wNmpYMGYyOsg6jXm7pWvFB1XfJl5ih7TgMHUFx+k9ye0eHoKYiCEQExKjOX2
6vP/bMzTkeH70ml8ShSGJ63FZ912tCQxk72mBNzxmiBa6jJW84nZNcEKSoNt2o26
grv8AK7a6iK3EetAhwUZ3MLseOP5Y+4YLprAiTXSaMlWtZaUCUKoGWhq4PZLbAFq
jJfrVxJv+5sj0cxbMYQikloqTs7iv5wQKaNXw5TcSo1IaVWgDA9WZbDroIKRifV3
D88jSSH66ed+iHaU3W+g1CJrkDWugC97LtPOhcttwErRH5Q5WgZwqMgUCSBL/0/P
XxQEJMYWLzkwU+2vT+z2Ib8YJ8/yYlo/giESW5Tt8wEUee9JiM36C+mzw1/k4q6y
JfPT6y0jqqBElcJEpF4bXu6tuFfz9GDYv1ZLeBY8HSWttVlC3ntFaC4OalOL7JZM
p4grHM0E+OSGx9k5ngpYbRviG7DfQsecRUCrpXdgOLGHjLhZD/U7QQDGjJc4rkou
VLlxoL4Bgkj9B1cQJP/Llx4MokbQZ2R9MN6MALFT1VhG/Gm3n76O/fI1Cqmb+zet
K7KsuaywxNvwaQClneegtR6icOWfE/2MJ0jq1yJ6aQXqktKicypnYfaIZpyxhj/V
pDaV3wHUYIEOi7+6878bh1YzGkGlhE1CuUFVZrBe3SQSIfL60DshQUErlltbt6/p
hGdz3c7KAnSSFfWEN4LgpgVilZfREoLIhKfCliJuxfDXHHIXc6o1zkmBsESitcgO
xy4hKFFY4XS/A+V4fyw1vagzediFg/s4/Y9u29hd7HY9sgIjGjQQXqpGzB5EnDBp
CnWeX7A4WUgaPvu44wJEU88IF1BPDVBmsqcFhMFmLtcgzSVBCMLm/FQcYGqtjpBt
BxHye4Up/mjcbRJotr4hHVbFLBTmG2pjgDDiYt/8+KLpObU13ysY70XVnf9ppnC/
qePUrQ0bCwkV5hpgdciG6aH9Gs//+prakyBe5dpAgFYQhEVmTQ9AX7A/fybOSQby
5IHkfclbIXlOmyctCXR622RMv/nLh7ZFsK1YRS5mAyf8+5fPJzsWA9pHgt2JSKE1
0/gB+U+ygHRtZADXL4E3i8egIs1oVjQIceiimvKhhDsooNQSYQPv2fb45apIUBzl
cB1xSzdlhFU9RWlqoCP4WwIFVRQkmd5HAJQN2YKSYdrA1PthrhR3EMd6tkCLyFZ9
fKsFlaGGfhQLoB8XeSsYVYbFNAOFd0Ib1AggqNf24oyPwm0lcQkuWiodTboKEXnj
U2HIhFm742BYOeRJj/LwaMNu3BQaghX3s0rjGnzU8gEziMKqGuAdR/dMzqtl1eAI
tBSqX06KG3yU3utQroOdulqnfVW3/obZ0gkBbgDci4irgiANFfU8AxvvytKnxA9q
K5CZsFP+jHDr3zoLSLgtirgm9pkWLu7Vm/AyyIrYIwA0IMnfAWlyjJ8XYVqvLPJf
gC70ZxWNubBsy3CIU38vIITPPW4Z9wGTsxslE3yWtYrt4aqRYSlnH6T15pbuxckG
haU1uGvCDqhJdqpujYU+m88KXxYA137OLOWrlkDbyGHFPF+PTF7CAbtNPSWFu52F
Kdq1Z42VDVvq5cBW8MxhKtvMC7qdBNP2NBS4cMp5GMFAUlBw/NDOlR3SwvYPUhft
29icY0NFpZl4lqONGghvY75y8sv3DWqyiSJ1PnslRp5XVn87Vwl8pu6u4sw2NB/Q
53E1k40BsKF8UZ+Z2Ol1WtzwBnmeme0EaIDhEMCIbWyYtKvgO7Q1+nm05HGb0Roy
IlLWr+DWV9IFoXwtjApTDcrtzNHG9gyE7QuRzkZJXHSr0HNAeTTjr30a+GSPmnVH
4QJ8U5YYRwnmAbuqZzYYIQnGM2oq5cX2s2Swr26dDTDacdiDN3kK/3rcYpgFvbon
AVMlVMAcZy9lIfy1Z1H9zsGF1LZX/YOjnJxO0s8oqaD9uZfQmAIqJyWDhU32xKki
FlxIhnQKLn9Ue2v5uTHVCbqSoPtqzrEYRGCatXegHupVuXS20xYyEFVk0JpB8whH
1+TFvzEWM01/rqraBivc9s13xNgQuEVII5y5Q14dG3T3JRlhICLRZUXLvQxO2H7r
hBVEZmkaRdv91Gb++uDCPuN3N5igcYq+vLb3fcLirfqYsuZKmGLoZlvvg/O84PMq
vmDg/hlL/iNHT60/nViFDnElCb7qxYSoyha5xDXbOr4GjS/+pV3bQd7p7jIImf4A
MjtI4e8UBP4jLVa+YsojyTDzArE0Mx06FdBr6KkfIy6o0jN6wS7D/gNcY8zuZ6Kx
A2wHgnVQiwl7F91ulUpld1A0wKnwdZkaH4wZaZ3Ji25bvK2DxDktedoFSQ5nZOSJ
DIqSe4D6rVicJcL8c9toalHo6WbHI1Ylg1oOO41YAE1qJuPpWIQmOyMEkLeXMzK0
3v2YOZRTVSdLYSuahQogtaUdN5ouX+sh0q5gpWsdOt+2V+iaw4enAXhL9OQEg/Ec
sC3Lxqtmqf8LSaRuwwqYbgyxOI0SS1vuBkwKKBdsBnpl/9/xX26n824M2yE4J+ms
q8HUSLtJxfU+2a3QoouzRP+Zn1yJNAGMNuPWYuGprPEfYRKr6flYwAJy/Axh0/5/
iQqN8TRbxOnCV+JvuCrjPTaJfTZjer98HTUK15ceGVYwcjqdsrGluUaAHTZ/a6Nz
iiQ01eEsJ6YetsoPSDrDQEzORlqikDyhoBXh7RNb6pBiqmYpDIKj54F7GbvwdHjb
7toZC4TKrvGh5UyHucfFt3usQvJ0xsC4W5V0ho5XPHoquwUJPIIRIFX07nLjyXk4
73AkfdXpkoaFzdsijQiHyQMXlxCsXayPd31ciedVfMI91wXqEOBx+dvgLklTBJzs
QVkBc8R/PtzctUmjpPdbVN4X3wNpwgbJ3jj6uB05/t/V14HEkvhjnRWTGJUWK8G+
9HG2VIlX671whZWmGaXhdfN6SLDJJlUZFq8XuNQ+bqxom+fP6IRLWIFsC9XVMiB8
tWVHbURictmGmzXhW9wtCOrcwSh0QMFPM5ieRq/jalA+E335B72logsUOs88s+8D
0R0fAB18mcanwMGer0eE67xjywSrUgan0byU0uG+XIEv3SP4qF6pZmCmUfOPWkI8
bHAYEEkM7Q/ENxwYedNyWYh7ItTNBM7n34jioXNJIegggszjxJ+DVQKzjTeaL0/u
MzKMqYS+11KpAbAm/f98Vte0Pn0LwHAooxSJ+fFnsnTRzFVIrEbTLbqkXgh8BQKv
d1H9sV4O4gOS9WtWpsjpSdjylDuFi9loRFAtNf6T6Jh0ULEkQqU5rZkiMFmXyto/
doeWk8jYZaZ3a+QWPt9vqSzcqCGeP3KUF9zMuKQApi5G+aL+WT2Sr4P/YENKk5cL
2eezskrOra12ZgRzafTosCvpYX8Bx6GDlQKMxX92l17dH0kKPQbj6ez7AQbgmUL5
htYtU6DWDufMS5eKRKA4Tfy6N8tRIogThicIXx6uQcB8VZWL4CBF7gdD1iDwIpkJ
p07FJlhj0oOII/HC+JMq2eL3TXc9vWJmDTury/adVYinNedPlgPlP5uofxA+uSzF
NjiLi9extXrrS3xFtKmpVX5voT6EEDcIVxEVzt/smm2DtGn3Koij4YbDufyNrObb
9JfaXUcgxfoE/tVFDMR8kEPirLxleon7Pki2eOEKYtjBXxMmpcLioHIAgtQJYwTu
AgcSSUAUm6QenWi0R9aRMVijv27EVhwx+vZXCmsDmUjYZx0FykZ1ZzYNuTifDzV3
fMu4RAxskqFaxacIiF7HDSci4JwnlsrXHMes6kUbhWY2bltMBFwx4v+I6bTU7eCZ
bSQWonPJ5UfOO/3AezI51pHJGtHsUk0RcmscypMbvWDIkczw+eqROe2Kek3h2hUV
drRaVFYGtINoeeu1qX+loBXIHxjIzWA8hTBC7n2/NZgXL9W+UjkdUlmICVmRWnmH
l2MFL/hVw30UIMAFAhX/IWPOA7kJg0kWgNX6Elxl5lfEKAn3T1A0HLjhY1Nxpw2Q
NL17bwskOPV1z99vlB4g4o34gUJiv2D55ZU6/WG2EXPn8V20/H4bni8Mf8YadLG4
tEUmiJSzCKxEvJn+w1y6NBVK7cXveJXqMBuhgFMlPaGNrWW8eIkoyOUVKhLTBJys
I/INgE8NfKGkQTxwndkbNsf4qCsSJg9hLESJp85XWp9IRyPWIbQCljEixHewNpRP
/EBFCMa5oOZYeigu9Kr+iQWZYVJJtE0YyyiKHxh7GJ1EuRf9dKL77HlK+xO3wVQK
dbzEDUOqf13IK5Rvgyv6VrItFRoeWetgjTkelbrROMv5aKhw8EPBK75PHAEryKD1
K1bscRTcj24z3qwP+/j0+XL87z3d98CjMIKXC2KMvBg/OQJnG/olRdXR8a0dJe8b
IPMRFpOsKUSO4jJ0mjVQtUjiYMA20/328NXG3dofygOE0ev5ZtSa5lXE7dwV9BtY
dPQWlY4ssa6jETb7BlzM5X1v5yHqqmRTpquRsg4/E3kgUsMZGAIwLrTpm6kMLrAf
9smZuFdyNSA2Lnr009SKDo7+wRyn6hZ+KFv+2p3OYG0xQzIiHdjqE3SGZh7dVHkK
EdG9Fm6aoxde1i65DoXLK609cUFcgTsk9AdHAizVCv5pZR/jLr9sHj1v+H5T4ueA
gBtwUli8GiBJbkaRkulzxYWoC1mcCGDE2xeUiTUYyJCdtI0gqxdECYrIQY6/7iW3
MDZc3qrcwNDiCZqJHsPj3AOoK0LZ+OIqJNK/rfl0rNl6saO0K2JsCiYDWLteFMQ4
sT0Y0l8ZLnjTs5wrWqFx6VtE2qXvfMRuwFBUtcyNM7d+exdKXfaUWOEQ/uFw6hoz
fHqySST8GLN3rCJaBn4zs0bSC86QY7Q65HterGxOYJ9H2/u9zrlLdfRDHKeL1sAU
VMn1mrSbkl7Ms50gZlzSdV0bBMzHYU25/iIghIjNEK5sXdlrkZcy1MX56V9mhn0O
QbhAJAzkBeq6fV+sizVp/yYyUqk9m3yZBlWAt+3PmVlJagDy0y4JtwdGYxnBToLT
1KWzkckjtS6GdkmLtmQz2YTKBaO1iwDFfUwX+FrSTNIinlBLwIYyGPkfyIFLDBbo
RxyPISZD7+9sHb4tIEgxwJZD/kF8lLIrgIyJb9EgiXQPbuctlAnmf0XdC0lSoBHP
+5WAh40r43x6UhVeMXTX2Now+cdbknGQCOjS7mPI8Szn0bFqhsT6kJcOnKBJ6pag
1mVGINNnR134aNMNpgvP9lqkOu00eN46CGU7kz8cXrLtSSoBoU2dt7AZoSXCND8s
9BTZ17/kXJKtz7RMjyKd/mKY6Al1dq6vrNX+BGTHpDWSD6Obq6pAWoi51YQf6RO/
j704YFLIxZX/MRO/RXL+GRvD+B9cPa0hxRyk2r76oLRtw6/n4Cy0ZCWBItlNaNzE
w4EEr1oVRollnRJk6wbZn+Uca3omfO8A7HQo9c7+VGIa/fJOUDOmostUo5QEewMY
RmnhrLrGEEVGCfda6ya3c1WkymAYriHBK8FP99aLd3C9OgGHzePk9qYWyPZBTmNL
eSLM1MT7ZYsbNFmfgZvKVg0plj5C67S1P/tohsUbuiukOhciKpBv71Id7syxlXoV
cXwUU6ciQmWz7wKOGqrXYZFrWypF1kvyPWbJTZpNLE6dq8SHqZoYZtrMXTkcWVY9
Rni5dLc+mGDCXnoHep6IMFJVygQNnuemtnCxO0DcMSTHx32lyFKrjmN9Hd0X5jir
m4Be/sMMiQMe5/c/KGzUqdXl2Fu0Ct1ZGLrrTdC7CgQR7/nJTpGuvi/+hH3F3dF8
gq9Y6G00cZSmzGJQqbFdUK01trrJxVHLp1beLsfPC++pwYpIe6b2c/O9Jwjv5xOl
hPdVciBh7AbS/NP+lxmdZk4+OXoedNZHu+8zq2RaemMUvIJTfz0LKBIJbI9HZxXJ
gMcc99+wpQ0N/bIRlYpaAgU4i1dkM3NiahjJpMs93Ipp0tBVG2WhTWsXXsbjCZ5/
TOHMOiFvBsdJ923If/O4j+7oTsbk3eByY4IUSJwINU5zFAhiFTK0EbbO3I7ShuHA
wlLbFAoIkm9WKVIDCJtiTTd6x/ZId7P7C7A/fVQpJZpEfAS4m+ba/6CRQqnDghEY
k+SXlJ9VOddfPl9pfHYPr20Z1oOU75yfYrTlon4bIKx8uAVF8RlllqmZ70fUruOA
bOtjx440sFeAZGXvxwATmOMCrWLSL3fqppG2XSmuRLrZXoCefsdxKzBW0BOuX1wg
QRVYvJP7i0xrZgBXCxGmau2aBgnqJJitVDSLVb0cEBor4FdZBotAkDdceDI6fMMl
76FYEMWNpUNBQSTD3OlyJhLaZSlO9KKskPn3c1SnK8iq5Gd40/cr1bz4Dzq5p+WH
eN/787/nVNYehVEQ4Wd4vPR+C1JsBbNGup94IXESf9j+4gKhxgvvMl2H5TmTNTb3
jyLFSveJBlN0IPizo2PRe7NjCLnsGpGgIKqSl3pofT1Qkg74opx029PzNkQJ5fx7
ItFUI6IWAG6Lm9MVlKHmR5HciKzk5d85PjYaat7Mr4reH9O60n6GQ+aCbG610rxo
RsMkYbN/paZknZow85C0DfMJL3bPyZyjgK3lmq6XLIsSnCh6N89wfbN9ifaBB7IV
a/t6K/zaOADH9T5VYCZX/qRz4rwh3zbRBEPe6eyLe5nEkvvp/wpVplxkDRVjbCtf
Ba865iQqWwNnFbb7TVeWw9SmWe/cD1N4tFiDPrVFFoOTcEfKTycOsVqGPF/DZhYk
R2OC9GXXDatA65hInH8wZ4UTP0E4E7XLbXuI9cxjZtPK6GsE+pzQzWRCnQfuC+Av
zunx18kXiVCDBPBQgNF52N0dOoBkYnl5as5zVa/t3qu1w+D6+dYZLJUfZgDvFJd6
AWOhZ6fLmfLWSD9LOkxLHSNbhMfp62ZhRF4iZ3XFbkB069hjll4rvCPg8wO75T0E
d3GxVATSUPbUAqYStOGODdsfu05H+zc1ODCbiD6NzJ4/n77ngts6eYeiPnaBMVdZ
eRdSpAP10rS47lPo+ZyNYmvUaCai7eVs+/ZVxGmuNQJBHqK7Uj0MQ/vuisOv20Hx
zUSfugUn7pymN9sDgLk+DZuEnKhLcAJkHiLKldeP+4PEpxrkRxPYSKCqdh/A3297
Zt65MD6x2ssDi0+IYqZx6mkbneUKo1HOPtY2LFY5pVc/0aH3biNnmyKZA6VqP04x
0w+9jF/V0ljx34jf7IuNOB2o78rwR3cD1u1UqlJ24pGk8U9DmEZrDPf24cPOqM7S
MTMFf/FTT2IkSVe2xlHuJfN+1eqV8aBrgun3mrGkA1vfEo372PFV0q3DalJjRe+Q
8j/nBZ6K5AjV/zxbcKKqpzhuJja+/VL3Xi1nYLAlVkSEt/o3xCwc07lWJDdRjtKq
ISpi9XPv6yH1vUsOF10ftuhxxLly3nIzIEhdrUhx0tDLHgX0n7UjlUQheqIJrLEq
QQk3i04JJrA+cxlkPZHKjuuwk6TTNrf3rbiYfKTn4mz9OrWkTkjsEMoapUPFd/67
WNDClTHWlTTJXBink9MixOQBaTANfWOsC37auQEr/CfYnqyfTau0XjSN3iQqvCw1
qrdhhg7NM+KpvxCeXo93AbdRx+hPuLM07thFeTKVAhFI0vcUjRL6nxQr2PQjt5nj
yiVIL5KGLi8PLJsV7/pO1HXqNuSTyD0Lc1A8zRe5z9Bhd2joiw5QweiAc8bMxdSQ
d2QzEl5qk37ofxfZnmhPqVI9pFBnqTUNHVcCr7mYN6xGt1+VS1k0xD7lffF/JaXB
T37ISWsoOgmsCKGSt98cCMliGSGsgBrkF1bKKlM+cbJ1F29VPn7fwwzKbYCo356R
YS9WWx8dN44nA1lp6W8fkC7wPHcjg07yXfZFS3H4CNQb765zGfJ/F8ylx3sPFaG5
/WtZHFy2wIrKMCIEO404aWNfkkXWnOciNoe6L/atN2/Mf886GtlFL+49hl7vmldW
NAORw1qp+k160tcKMGZojTZfMSgh3AR2OdWMYdEVI8ut88tu83Mc1BLArfbxknyF
r/IXAiFrw0gBHOdHJrjIUdyTHMWJ5QIWdvYusBtLVT7hrpjBdxOOru+O0sE7DgzA
JjEQbDy8PfBhi/exuPHkiuOM/5hdQy42qhy04EYw7ujrmrEUVgmkiLQgVhk1XUKO
xJt51LqmZ0DJMPSE9nD93BnXlFgMtk9bP8+qf7zSo9KRmuKeyRI1nWTylmq/RQzu
zbjZshPSQq/S0fMCoDaQKHyMSs8nftXPgyQdFRp7P9ByoRxUXD7nkCFKhjNtbb0d
fxl8psbjwsK4bJv7XQHmgRSmwvrSNJoHUFoahK628zsALxEFoKdzMQ4zdS0kA5UG
Wj9Sefslf9nd21R3O3qd+9X9OT+EilrI178iLTGNn8w247GaYPQbNn+Jk8c0GrAN
pO+3MoKslH8v2tgC+l4lX8XWJ7yv4TQnpPlcrOZhq/Kou0rOoPSkoVLh2BmK1vd9
JJU77Km1UYV1SGQ14riYAL5apuSAch7XSiNLAwyDplIBmnIgsRuok0duNFEFBEju
O4jt/ETN9W0IxK2te4RlN4jBYkobRC6JryMHJOb8q8BXBkMggDc8ogUQ2zAapF7d
rxpjlt/o7YqD8j4uzbH+pQ6EIlmJHQdI6OCrbPZIpPPGicl7inoGGnuAAZsXdGuI
VsUxz/b7w/el+6bJwSxp7LlhhlZu/Wm7Gy0g06edpguYydKk6nsFBoC8jkenoyyX
peHXgxw/vSuIaGDNwpr5DaN55xtOgaWz5OCMP1e2UxK/5KGd+b5Y7gDv2nl4uNLX
rj9zaIhEh9GLnKLOs4bo6oH3VYB8Qo3w7pCkB0cLflICxga4p9IteuxrYEHaOGqk
nxogFHhfiYD0Zzlia9K0LQa/sQugg9Ims8f+ADLI86XsI90dM160M5vjmtLNNE+d
AT3Mo7mmPZAQPHitYWhQgJmUAWSr9hX5B1zucoqD/EjhGPNaDeYWNfKEmFhLa/5s
OrGjsF54IsKHH3fP65Eww//V7hhLyjTKBmeJY2XyoqNyc/b2VEmH0AYX5vaPZuqk
ONuSqMH/SypJCxHLpQ1/rwc7jhOrjQkcDV09MLLdFa7T5WQdwG6o7OWoPF0pNwHj
P0dAAFlLYra4/QxhRKgHfQI8oI8sjugZKBOPfxffOcsGbn+n11rpVzn/+vaOOYs9
ywgHAVsZmOHXrFdWJSCOeygqvgmb0KuKsdB7Lja2lIoLz4MRuYkx+basyGxF7KJ3
qczy1N9YPrvSys0+HFYZhAjky8/YSq5ouINunRiZlIDRNuLTnfNi+8tVejPcWOo1
9ixZa0CZlMvkWYbrXnFHLbld3fUQNa0Nib1BKT5KRfM2BLpTbLQt9PCHP6ZPJxVp
26ZU2xHptguH02zZf+YYsQVccjZ03HePtfzauNfw3NuVdr/Ql/CALl3cV8lMuMNI
U0slc7AyJ7s+GY8iNpdpq6kfZy7Usoi7s3On8LbC9G2XqfUR/DGqz4q1NbWGCinR
VIxBfq9g+yMjq7qhGwHtBqVijLPgAEtG6wdNhy1m0wtWT/wpuoyGt+85RmIPcdCA
C579aktx72P+6x67/Ne0wn9Y/aJOAsQRpMmxTAhHeRGF9nQNBAeVpZLjbXxMYurW
cc7Dqkcq7S28JMPvHEXiIHy5CV1sxC7py+qxTute4k1X5JCJVpi/ZYfEpJVPITbl
el+E7vuJqbnQkBRDa2DrJS3NnHRBVxRy9fyXGMbDh1ENnOG1nsx8+YyUyIU9cicj
j/XLm+t4vNmuxkOYv0A4SsWmZoAyG+rTDYq7gil3SQjTywwVbz0aSwQMApRgbfgv
5WZ67oSHQ8wUFIZtDdK7UsDT2HP5oPfR5pKZ/K5X6Tinio87Fk9kn2kEG2pJLehY
+/4lYNjpyzdWXtphYErp5ZGQAGx4KVNG07dH5gVZaH03A4v9FcsSWwGygdX9RyKL
LF443u1L+8w6y4A0E2GYPRIncXxk3vePBRsdjHYbmF77VYACh4XSij+qRP0pREyn
hXkpHt/0xnBjCRzw9FWeuXexM0i9s4peKOEVpe0UPlYyPQyqlNjDKKdNNyf2XDwJ
PdapkPXKgnd7pKKo25HwhOj8jqzpwLOCUhOlqKtzP1pu0EvMVRdCwU1cVDHb566G
b4MXTcfxXeF8fMxpSyaRI3q3FQbQ/agbJnYl+zBOTS3NxXV3FackLCQhXR9YMgHZ
tjK2MXFB+16MkDvsiTTpLkT6S7pDSXGBCFnf2zg9EkGBGi1dlM7FM2YjmPk7iUbi
uBzEoq3iDtdsJLeluM0rJGW3AJ3wKSVLXPw+SVKTXs1hFpHQ76Sppt51z2SI54Di
aTIE0HOAZc631DnBAV/xatDLXZGw6NvkrzDV2cBaBOqQJUi+4lqun3WV4y9RBV0I
PG/w1YbRvUWYgSwum4lu1rAYeNYIIA2XP+fctiKnIsWq/m/WlSditoe9WjzRKn1d
Ru6u0CY9OVSIkIOHubxaRXag0w346ao3yFu332WRdKt93kGO7Ye+kpL19bcy/ob8
AXUBHPA+gIv9keh36hudgQWuzfoxyeHrKU0g9g3mYV9JiuxYE/WoCAN5sk0+SbDC
8PNbXssEJSRKKtEtoqJoDQbJJREvED2VcMYo9sJiAdDjuSBzU0aIXC+hzuMlKtrF
PatZ3IiE64rfMkkZHXmqv+7D5LyggawwqmQvvUOlKP8/kXXIfpJ5GLzgg0tSnYi6
7ofKxwP73LYovVfwhNOfIatzWEnHhZyBZUrVAhG9T9pgkkhEUv9W9/t0QarBTzwe
2aohv4bqO1aY9/8NBWy19CCcvkTA2d1UWZxpvr+9XtwmNjdxXdj6jLcof0c6j6sD
zw1AK1rm7BBJjL9UeqCQ9U+JMzNKVaj64Nwa/MCUQ8t7lekWUzTNCm0Z6S6pP+tC
M7mN7WebqoBBlsjcAlZXda77FcdlsMBMz3heDYWy0EDyJa8YkWSeqfqghu2SCrM8
oFCeQqvMaZejH5AXbS7bxqZnsy1+8lKV97T6Rglxux2wCeoAziwAxE53DfkxxnBH
27ZWd4l/nQWZh7tyrJuvviJUwbc9IXD5slXZXZ2a6QO7+FEo6+gYAF+hbxU00elw
f5cPOTJ9c2ICmUtdPni/Ffe9KwhEPaPlUKrGKpIj54EqWtdpKyRgY+DkMjl5VaSN
JcKygusegx5DFurz3AC4+bFQv0KY8pH+dGn4rfaKdeCunS8Qf+ihcT08ATq5Y3f1
3DeKGfHwJ1RTr4KkIRTdqpNA1DOrpPZHY2UKNGcB8vfNWRHpdVCZr8uwocWAg1ca
xWCSxXm7HUPjdR1hXClxo7YMjBu5kYRFKIbl937hykovq3PH6f63W4HDH9kv2WGD
TefFrnB8xPEukQ8Gdsozx0Q2hi2YQijDHPzxN90hGVs64ioHSgKjZPlh42YOuKE6
lKck8xVcR2Q0j/Cv9ryZ2KNkNTMISU+8+45+4L0gYQxpWpb7ggdmtz+wQ526keBX
RhDaagwp4lRYgFWqE0q6qQy6sTWCYwoF64BGvjpOWpRk/XaMEl0isU6mowydky3d
jtXd6/WlPIosccrtxLFhAZCXOTxljvoXgLLCU80/fnXAgkBis361vqah8yl8rgD0
n2fRX5yPrX1naZd/xBuOqfbFP01WpsGFYfu7shm5hz9e8KfjpRyJmVzKEWxThq5z
isHOTtb6jt2m8BHc5ajjQgPRFdBbeZMIDB/XV8zFJrdBLxrRD4sM00Ct5XMyZiU4
eyv0llE5iizon83OLKhiDlhVwNufNuy7G7FqbMkIhkBOScB2A1Xxjq39mbxrFNPb
RgTXiyVmo5YPQCqlDSjRdb+nMZvnd0ZV/mmniPmYRBhuHEhxO2ApCsc2w/wiJP0q
ylTFMzv87beJnJj/+vk8jLXWx9fBaQjk3+OXh9AfJAiEAVEg7IVYI9dkKsKxsB/B
M/y4XbOb7xT7/jIeJ3UxuB7xFbL8Ran8lWK3ODLyIgEhdaYXqpctg3AKSDVTgHRv
I0m87tOmPAqnRm12Tu+ZfiLbOOakUw3XMkFnhT6f547AufCrzSGL+PoolbpEMWUX
kj6tIDUqeVgco1FlQTPrN+jAOvnbb4zGLswQyTFF8XTU7BoXQpPEBIxSaHemRQ6w
4CfQaasrl7XUVn0KdbRYDp26cRu0s5i+d4YO3iRgtt8ZXAKOn6dqnv5ofy2VWwms
0SM4+gc+R87EpieQW04Wb/9dCNu8zWCFQTsApjO94D1tewD64ykaFKeiPJ4kyCtT
dTZ6xfgt6EiFhIYaDTUmHsLK4cmjsXlyw1F+E+Lzknr9Z2WVRDLEqCjoGWoJiWRX
hmD8KSxRv97lp3BjQoyMrfU5uCT1AwBjyMYk9pbRIxfX91GA9PSIy8RJFTTOC8Hk
kwBJ3voEO5Ygd+7gfrPmgpXUcfNeuX4X0dTIfJMAcXC3fJGBhuemlm61IUuQs++S
4D5odArz4wvv0fM2roJ1aB1ZRiC+aoz3+7BrEbWHi/vXD/tEoYyp2svmJicu8u8g
yM3Mkf54UZW3YBXreYBQVq64ABXu10gNH6SqSQ8NRIfqU8PPoHaT4RYng2TZZf2w
nmFLdEmphiU591czllSFlW/BcXaOnqHV8oqw+/5uWgM0ZzXdSffeThKG6loDNHrD
YJfmkGEb5xNb8ncdvkHLhBYLSxtfa4PLBuAMm0QKfvrURqNFj1nQ6VJHNLL9ULBv
CmTOBLaCVapZngoewLPYNkWtybMN2BzuPNhSBFtQvXKJdgGoseWi8sHnBvhUTqNh
dEobqSpowWJmjY5l/X4T2meUbE3Gn/gW0x3+PcyqSZsUJfpMNgOBboEzqEzn4K5T
q7vjUeWErA0ZD1Iuwg27/7DOGT9Ru7UmCLmQcSvgUwZCgxf1/OQNVVBtIz8kl7bS
M8/q2Wyg7cra+zamYf+koBx2wtK5JLcgL8p2tdZPmqNualBtt2AxLfcLgKeI/hbn
RvkT6z3sE65DbrcLpc5ZbZfA6jNGdLYlG4FVQzkQYgt95Xdm5KrlPuXA0ccpaYbt
5ICvE31iBvGoVwrnKA2AGStBPAl+yBs5RlDLj8Qdmkx+UIinuDFK50YYsjJDlFcu
D+9yEAJH3/z4n/l8yF+7FxAmlDg6wl/zqmc+hnyMo4fkXNip9IxDcFNoW9SZtn03
K/5N/VaCuIZ1uYGzcJZCSzEE+W7zXJ1wvD5gAiz0O8Bl/rnTuiZ5q1aXRt6a+cUH
lLOsYzEDBPUuBhdWpHNXdn73GmkhLuL1J4hu7aMSGNUw/W52+18cnuhMwr12NM1+
y/D2fYjGJSB2+zHvbKppfiTanCjI4D2isFJbArbNurjzlzNlP7q3p3wrvGt6EzlM
QwEbrl/+p78XUQN71NQ6ki+ooytQ9N1DPBum4ybLCU07Cqc82ps8//XuDnLoMJHH
FIpfm+91creFhT5c1PIR3yobKHysxU3LUL6GSbownSvYM2AICbOfQt95BcmtegWb
aWGo70OnpBQj03WdLX6UVW+oH3FDaZaJ7o3A6dwDmbbABez55jsLhhzNYdkXSy8E
RkKWRC8BYQh/CvCZT39CmZWxZlg5YISSFGy8V+wxk1RypMwDMAV+Xq5HyOS2Ai6x
4Nd8rTAzqoZDKFIYCPogd9vDONiG970UCSbsfIQD1y/qYhylTKnZGiIY7YMXDvGN
MRTbN90mgA5SA689ghA6gMJw5nC6603JrYKclcFbG29m005BLVrGpAfeLeUBTp+j
2zB4dJjT+C/vRaO5iADFoYIuQDZ9Cq+pJ5oFIdBwTa1aR5n4BY9MGhAGZsTgtZF/
e0x1+wU2TfqXJXCE9NH01AFYWDISR50X7iZNrD7g+ElD1aPisYvAsu9X9Tbq1uEA
soILgdLTpTOD1xfz+rnrfLys1/3MGY1zy5R07gFtO02wdC0YhCTdXx1lt1uzl1+9
JcNfu0z+RRplmAL4MfDW5OSsKQN/kW5zTbS5THQwsKTPEr1k1tf62gPG34kXuzGv
KXmQg6TAbK9bCjm2WRBAnh6FleguWk0kXUwoamTFzUtmrs4+B+a1tUXpIqouxRTV
aXvMjpH2APzsNQrRmWiJr4G0FOkcjxDgwo+fryqnIVqw0B+rOLhSBh2OBgu/VO2C
EtMXrxdXwQwEWjasK79oHLTUAa/y2wYZwqv8+W2QpvJMwu8DIGEw49OOIxheqCd1
b2Zk+FZ6YzT+kzDMy1FUvbQyrHmXasdFXAfyHUd8hSgW1BVgAiWFXsNVSYGeqIbj
dlkgMRWrywz/SfZIGZKyMJ1VdPgk7Dd2ivUd7AHAop849Sbr9PwY4rWCDP9oiPjr
cOllJ+JF1OUlraCCLn/bX3fJsuWR4qAeDyXngjKY7tvS8o4QNN9XeKZCz1F29cd3
IIKUZer7kLjcs+E9S2lLAvOGDG4ZEg0LMFhdzdgU5bH1jLFGQPHVD9hC/G6iU43I
e2RqxUwOVlz0au9RPAczkdsuvXIm6OZUFDATKOSzI9JuQuw/8QUrkxPZhmXKKxrr
2vxyUkDFcLKiv1C6b6sxQEXm4lFbq5ZeBRUUU3XVDdzDzksMxY+kvPDD+SnVmG1e
xdqegG5HF3qfsW3G8DNkth2qwhsNmiwgbZQdlq+qlLpp6OKBZSew7p4htCxnYD5G
bbaR3x660IK/JrQreL+6ccLrQKzsmfyjJwn9A+htVQ7/w200cliz7JjPuZj0yja0
6gUqcEgnSjNOz1/85aKon89nGOfyqJVnsFUsKq21NaG68A5AqdGpLV11+StrgZlX
lu+YltPbmhTekjnGN6xm71kLThbIRHRPQVhG/mxpK6kyeJIWCWwhLz53pPO9MVuU
ZHJyLWHD2r2mEzm3TOSFyfI+MdR4D3P2JIVNZykCDAHCKItTmEZH4eg8fQGXJWet
IgguJiYaEaBDKkj0C4Lp350pWP7mxMc/d+cBh/BZxfB7wWD3l4z0dfreN1Z0r6JX
RFdsCMhaIMb0+PpKtctWmmULsyCorfiyMXPb2bL03QKOx+5CCFqOKTNywryG4oQE
zG+NZQodCD5/0778kkfVOwtZFMgnrHKl6gQ9IT2x+M+bcM05iZoM6oqTf+Mkao8O
pjjqkf3fGnszN1fRKJI/qjX0Ou9Q+sbjggdZJF10lly5VlPRsi5xGrjrztbGPvmb
74t7TTZ8BCTYeHewGqYf+g+rmnblVYZ8hhbKSqQsy8v+YH0qi/iHiAj9mlwfa/T0
f0qjGwb/KvE8FA3bEoeMYU+7/SwQCXU6xLfmDsMvh25nJXhguYU0xbiruwqmWscm
mRVl5CLsUsyBTX6H7wIHnOw3EEUKoQ05u7vPsUs6g2dS7MjF0eFQGpC2tFuIBfqE
ZTsIWjbkrUqT2lgeTQNNa6HrBSdKFNwlWSVuxN32q2tFXIj+yWIVqRdI+AbofYAA
4Y6Kcs9Q4+Ln0wPc29H7159RVGeBj5r+7tEyZ0ZNDQo2xUNC/RMe5Dr8zmrBrdUt
sxy8DNSpCg5ACWYhUKn+UlcF2WvlZRXfN6yAbyhhwRgCYUOSPvWpsW7SiCIbWD9J
qf7b4VxIve3RL2IMDZbfaQTCksz2HJe1etrT/HRuQf/7LwsKoiVxxSIKTDT7OQ/A
nT337XCQ8BK9A3UzDmzUBvSsymVR31TrKflnTTgADr6Up5OrRxTXk4kgdTYU0ge3
WpJb0qFGyOLTvsFxWHrOoQAHyU+L8MIkxjghhPXxk2+sOcXzI8c6syLqXa9GC0gP
VUvpAEXnKBElvxe2bbccAXcqeT646MSWck/gaHCCgU2+9odeSRfwOiB0NaJYTzbQ
e518g9rvSzbVsbXRmH4VGuaPXLPCRoPWlOCM5OcrgNbfuWdZ0uX7S0sYO/c22PcT
VhFnsSoVaZZENb1OEo2FRGHIvrFhB4GorX1RQHL1YmK7vOPHJXPd5EuNmiB9ga9+
Kr31aj+pCcTLIFv54OQrQsJDDU28gll9ViAL327Kg7crUYqTmVqOJjpM3jwSLAUG
W4j0bYMJdYUZoizwxvFFZyl9m4S4J5gN2msVyQXq4jH5dnT84cAfMKJUu1ZvDeQH
o4MBU1/uYlMqbofrzcEBE+/LD5hOZPUnVaCQ735dOvof966wE90udhChJKzX353d
2NPIkGY9nvCcxI/C0ZsZ3q06/5gUicwl1ANy3RVC1w8ZstWyCcWpviZMnGMG4eie
WOM5bTHIIcXAILEc/Ixs49/Wzq2AK2Bsxff7bmi6sMFT5YMOga+Cxc2gAlgk60yd
3UJTxn5hTDrEgudVgqfMnvq8KZ4KYrAZqsvgP8f7gmzPmAfnZ820sdfCMQH7JNcL
i3Hy+46CieOem96iV6m3ipMklSsCeJj7BPZOgADBodIvthJ8QTLkbpLRB2AL0tPn
G7dfbbe50QeHsm0LsK08ozfSRWKEMR0xAKGBJwqEjRlCmyFLgnI1+Y9OzMWxFTbR
/c9Ljmzhs18TMX+HLWDy/7gi3sR+V+Xr7hIcLnReqi2HX3ImzLWidwoGEA06Q0oz
x8ZB2j01EFjNNX8JcZcgRChWOMGk6Cg9Tbp0Au0bUN8l3Lzfx28JkojXB4wqjoNT
0q49bkiN2rlv1miZeY/ZANUgPcYDlGSufn3z5XNw6PX9zaEoAp8SXLCgQCv7EBlu
J6Hxdv2dRXaHuN/wb4Q6fNcuQX1S5jtqoE++KXGBi/kT71HnsPvDgupIU/kV0o3A
8izJqN/sbU3/Hfc0sX4D009sOH6aIKj3i/QunL/XBvyw1DM72Tyv3x7zlHW0K2wc
K9kimQqbSs8noV7d5VDreBYR50E5MnJKz1BTQcRd2ynrQa9AB9vQoCshJDVYOaOC
vVEWJvee90IppH2rxr83vh/hd5gxqhsGUz35tivBOjCUny6Xj/BTUw3wJtsYQtlQ
Yavdjt5CRjpiD8HU00QWcQuyThIaiSAU4nv3eitckkk3LpYcMVwNGZ2HqyMrasxn
HUVgVWT4sbfo/j4LVchPqIAWS1LF8herB+VcuLkzRNk68dK64IGh0H5pepyfGfuI
ptuO/Vxsntxt8MEx308fxm0abQX11Ytlf1XPhoRGTsHz/4XHqrZ+VsJSkQnUn0js
Tx6kOL7rWCRQGmQ84+ieUEWwdHKI37U5N4274Fj8NUKzUBGRrTg82oKsMYzf1x9H
GIHWw0kOXgU9RSKOBnagSHN6CLn0tNTlPtDhT604SVJQYIVaDICM2YDkRcVHNqtm
dYLdQSjHTfBhofOJpfhNY8xd9PGmlCtbFtvwcJ6Ess8cckX3nAQTwBR4W2kAllcM
zC15ibGnz+PteWfGZpRNndKv9xKVU1ItQBoZUzicXJm8pp4Ja/ruVKL/Ag1SWnPv
9K1gJhgehyjlvnfwyb1RCRo+TRIwqRpZmstaLaICcyhfM5neL+5TheY+cciSXXKG
1CfR0huCfyaSg8PBjjAdXCoCFiQt9LcPlN1GJ3lPAyrScAMIPnKtRD+ZWFsBDFFM
IPkT6HyWyXOyrp4IyjB4glxi1rDz/cFvCFa5yLjDTxNtpNQVQ/Jd7NuqmwUexOd+
3Yi1lzsYksTreKKxr9F4q3aypihWNbiuVtv2UcS67jTS9LNlHaydx8MqFJfA0+FU
F4iYGSdf/d0uQBm1u3V4/yuLomwvL0CR9M+Q1ANQHy29/9m7DU0uEfggLy2J/Bmk
Sk/dPxvUDNDhY7S9yQW74LP9QvHAfNiO0AA7tOGP4s+ZeomKus3kAPZxkSK2aZxS
eXyaPhk9z4Rt63+q5mTlzqs3Pxw40Y1FoFykXmUEwuHoee2M5mKzOFeZVtLXVenF
vT0itW449cO8CK8ntlSkG6ig+/TJ9qmsc10ZNcLm25wxtk8pAC/RO1FoNsrZvpz8
SZtytXHauYSlifktIUlVI7VxP0tjRA+naD5f6XRU/lKVal0/aI2fpsthhbnzkTuL
D5KoLWNq/OpSio66Gx4aJphzq7B1cT9O+G2tlBMzoZavwhTLl34F9xPj7eD6MxTF
D5LNoMBiHpka9WMLpv0DPJWQtwK3j3ACv0NX25rClt9DsaBuJGErkKUv4N0LvBO/
XvKZi6dXLMmdYSMgUxij1skuzv7fkiVz3bi1UDNgLEBXFhtGqvEbaNR/e5ZKp7wA
lDBlSKIpSfiQ/JMkOQk5fLEcJpOH52o6xVJFJynGKnmBA49xdCeuRqGSweM51D66
UpLq4YVdd/0M/4ApklM6WgAGaDgCyGOsODlA6pPcGnG97Nw59eNm1DMZcGjaJnRb
l7DPMFuh07siDuR2ImY1+qiAwy2X1vHVsVoJqkeY1eFjcDmAmBP6xgX3DCcklvDt
YxdetjUoM3ACYQ9Q7fU8LgREbDwFC7l06qjIZeE1tCGVdAAOBlh0g9AauDxz0bhS
OLW+w96gkZdnkjgBHKhd2iudiqmdvMNr/dQYju3mBoIhm/yxxDMaZ/1kLNY9E8Tq
Ix15FkJ9qiQF7l+JxLEx4fiJylaQEUNGXq9z+S5aDh7ZxNtBUPGiISFfh033G2cQ
0zg/uZ7L+9MxBxIrNbJkfwuqBJx8Y2JskrjO1pi4SWPkGUUPYW1ZOYM0PjS++f3I
i8k0FYJbAnf1nLAcQ20XtNPnSJBjxuhgpoTW8J4RrTAkjyj9mNnbHJrPibvXjXZn
UvWEoNOLuJG04jTf1MOhmGjCAIyW3f159l84qOz2nSwWRkCj6kahnbuBXABmnCY3
fcwa5cgqrts5Qnr4fIQqqhqwqiHxGoc77Z5mgKcC7VE84Gvh+htFN+KHhLxIrAq5
/HY2YYWw1Bhv0j3adf7SMF5ymzfwy4upXi0tru62kC8lw3itpvc7wPgOVfeQWlqz
fyA6RJErq57iHQgz/mxF6MaC2yZNM030eDZgLe+oQlfWF3rj3ekUOruMyZjNJ3Wk
+eUn2XAR62RAI2fnNlUzxjjBBBA0OHvZgKn2Di33OjZU1ZELu6dglEdEPf/RRAgO
YFAJMEMJQo/t7clMe9+l8BelHrT/bpwNFo0UtUP/I7ce16va2YBfGiSgUnFN4CPX
qKRNGQXyQ/I/RhM/QTMT+6UHV7moU2vZcxG4yi11JA7EVGIjnW5LYoQQ7tVmWqne
EFxK6cZM/2EIL4OCYdJCOcI+Gr4kRp1iJUCKIoIIPesi8t/oC7NcvTrQ36SDHQe0
LZuq9bJs0Gjl7OywKGiiroeWaBEqCQ5KPRTyheLbC/yRtE7FOx2HvW7DhtejwdKF
pWzr531vNIOk41/CWZKrMVIPmsJmU7Hx2nP9aCqolGb0XcyKIecZtsniRyhdlNd/
9YQsGcxxSnQq00GxzH7msG+qcCCJzz9RpK+RsYGn+1DLTEZUF0dFmmz7xqglYV/x
AF9b6BpydehtZIjdxx3xJ/qJysYacXQyN2VbIUhk82+F4YqXbdI3LUR92kF2mEwF
7g0xy1kucH6f1JpoktTGJNoFfiNyxtoLRWzGb7cNAsMX8qWbWRIZ4iO3pe89lJLx
pAYTTP2SCGHODdmyFKkKyeieunEE1GpgsgmarExZ0z0GX5a3LaNfq06VJ4q3AwCa
qVAFsLVaUJrw8Zq2SAmuUIFv2uL4n9nkXy5IrcI11J/T4JrYOciulyVSDW8N6f82
7W83tBe8IYUHzx1pSW3DIFEhQawBhWImrwxsSybB2pDGZk4dhGN7yJ7/JyAK8dD6
iEoX9TdjmyNXpEwtV3SNc80lfYWkCGr958XTxrCfzNTViGjyLINilfdVIOI/YxYK
xxgHEHUdKkN6+trMMMCr1MYPoHs9xbVkpj2NnFAwP6Bx1ekNC0Le3A93OWhE8VBc
XdVmM0jVf19GFN7AFs32aapJ2SqbVkS2HZWbMpDoATRmZz8ssafbI4+Z3GOVw1sX
Y92aY1/z2cVgd5Yxk1qPbTlAwNmbRGVcRtRvltYiCSXBKwHADp1lKTNGaWgHUSNo
HnISiaxBhmyWM8YyFh/wE4EkPdt28kuv4wd3RDS7qkImF7lwW65GDDKYk2gxgBJv
GN4e7ciyOW7E3yquP4xca50qa7Xit6oKc7YDi9tu2BemsGpU78YGcD07uGZ4U6B5
grA52o6sk57gTF/4y9ELbtkWef1aoaD/A72TlG5bFoELgLknMKqous/1+BxFmINU
4N7Q828bEth2ocztmD7o1/WZI9E8Qo/8ozj473R3TkjKfdf0zqhkqaRB2Uugxi/l
//Kzc1ID7r+8uCT5UiM3E9cE5RRp3HYclGZdceRcqXnDXSLVoqs7qfcf6NIN68T/
fHfZuInarI8a+UuhKLnGPS12VsFqwYF28PAlda+oWVZbE4A6SqtByVKIySXqkwjf
zFhkoGjdjXeb0BRW13aCXPk9eQVl2Pxev4E8N4xTVsEim6wHspfsZXrabAS3GDcq
pa2BloHFxGKI/hKTqWIydE+/xM2s32bYYWrblDSODxx0WpMiNTsIfLcuVSYllEgt
XUQ0uC7aGC88qVrNMM0r8lU69B7qLu1m8SX5Z+Of1tVJy29SRGGiGcsMIJrQ55xF
7+Tnirym+xlKbFKJtKBGdHKIPfzF76tLLiZhRT0APtr0DFQIzw30APLlQaZMVQqe
Lftv4m6WSDoDUoK6q+He9iznDAlP2WJecovLbprKTy36PGFetJuNrJUP9LutA+Jl
i+YEjEJKe5VNVzmxgsSTlODOGxv34lto9nTBDedhw12RmGkHhdEiV5EgInyFro8M
BHrLaZ9FQt9RIR2tai2k1r9UECng2NaBemLvo9lpGVpRLbJXSvt2Sw3x6DP1irU7
OIyjH0BvuWUWGn/OIMXFrZQPHNhpM8J2RCgjJVy1JZE01h8W5k1ZRBvt9SBTQt/+
KhxR5j29siF33W6bP3gSex3G8FGEjuz5CUGK2Ci4pyVexHdcD4r7LeNhP87pqb0v
M37HLlRfRnszBdbwPKoUZCdMeCUUyeEw/8reOWT9Gr8WAKCHbT80ty6fEqv66pId
MMknMrjylk7fafLrN7x++cE5l5aKki7+tZYy39MPzhQq8551B0e4VUPTJKAdCwC2
MlSsrmO83ohPK87tnzM8p8zYVLEST4Ae3oIXBIaP4dmUTeiCexN0fbSaPcUM8S30
KHRk8e4Uu5HW1YNHJyC0F3929KvyZ01FLlJx1Y2dljzsoDIYpX1ogfGgH2/f3Qbu
yoKC3ByOLsV6nGqIQcPNtxVoiSmGTEiYkaOrxaF1IsH29ZF56I9APztH1duuZpl3
BnJEFGx34wWycO1fZA5go9qcxJ3P4Jt50A3OjHla8zGyLidTHD8GSyRDa5S0JLe8
MbNG1m/20mVffbgz3lm137z7rlx4kNHw1gnl46X7mU2wXJjVW0o3/mqzNqx62Zpn
zLiFeaEd0hyHeNCn3VtsGMfOV807fYc7FH91uuUXA1eLtvQM2o9N23Cig3JR0AQi
Hh1MrlewIkk4B/SXxdajqFScrqW4OoaJ4zdKIUVMngIzMyuvvj5Hlg0Rr9PEDgzD
D4BZrKAPG7zmZ7O6kxnPqPTqLGcvew9mmS0ruSBI0FLbpb11DRaDA2NNkyAc7syd
hoPUz/+G2WZl3JWQy/INfy+NCV8IsqrRCejhyEUFGBkLPUwmFGS80U/21fmXGtnp
Dk6RM1fiwYIzqHYt1N3QeUIL76/5jF0JCZfYleoj2x6vQgOgvGSVty8VpgXo8u29
a+CoQnCqyJG74lcLO0zKX+KfRzqAZMyYi3JePDiw7Wfm9gEKILdSqMLwAuEAWqJa
I6KDBuDiNNCo+C/3waDY43adLZz1a2t/DhRvacf2LgYNvEG//dphGbJaCSrK2lP/
FYrtPgmy+IKQuyx5hgyEdtOh3ySDm677VZOU/9J5luHPxDpfNMyhMaRnbvFhyaKz
wtdFBq5ypFpwRGxTJVDnLUuAusrkowbOmmZQDdnqhSe8NEtCNxitQjq9NPPGgKxy
sjVO7Ea9guu4ooAb5+i9fIXQuhDehjF5wVr7EvDoUXCPSA1kEByKfbUwD+aRXzIf
CqtuxmjuTOfu4Pc2+DBwS94VaLjFCfbpwKvjVTgzkyIXhwLBGHQWC1p1MNa00dz1
Hx5GJ6pmafiJYfoVRrXOciCgPGPWtMbLDlDxLxVC/cGIbEgg030XKvM6lKsTqQcz
jQMI8uPhbOyxLCfLTpVH0Syu0wY3G6FRpANtJw2r7Z8jrzcXMYh5mPLeroyQE27C
+EogIJ5UGJUCLmBDod5HWeoIJQ+LYMsfsHSD+xVuEptucX92Hmn7fjGYJsqXBG5S
10ucLebTsVngChCRtutWQQvDaxM48Bdz1d7nOsQ40XT+1SzQIccv2TgLxHokWGnP
5IE9LzvGjpBvcA40HJOBSoy/8rGnkXUPpA18hLRp/fjgKS0wvC8wA2nszYAICZLA
AsoKG6eOXefnO2jpw6R7asxviEBQuGefarTuol0VIUhY9YTz8r1F+f8DhrR1gxXT
HWa4eKedxXC6T/flfWLqA9e2s2nKQ7KZsmhGyZycBDEQHHwtiD2l9xG3Rq+OmMH7
g7Mhb9YTPx/OkZVmF4QSUVnTWzpWfQQz6DA9EJBGS2QddK/Jvt/ElLJ8FW5jzab0
Neu8JPyb7RK+uQgbXfixiS2QUlxhV89PugbXBShUpY/GAIktnkpA69SZbgE4wd4S
Ul6kpvTYhcT7vpSfC38uKZLaTZkg4IbP7rUtoDpgLHQlO+o/+P/ErHNR9HvOi3fh
IbyErznAL+mnYdiWgi2OHOlxGOuj7nBd80oRHT37rAI37q+CIwAgCZnuuTjInFgj
47IM6v/2PxA2F+Rb5Shxa2McIOF8WfvWu6Lw5Wmesyo6FkNOoOGqu5NgSKxZeZdS
3+Hf37ik630ZVMRqaf1apdF4sxqv2uj+a5PG8qCKthjhHKdJvjK44fHfFBPMZ1eW
wSN8UIyXxheut4OGK6qyRRkUlv7O01JbM1BYkTjxc5TkZ7Btayyr0j14FASbPcNg
VvYtJoY8CA6Yvhn0nLrH5XAAmiIjOFtmiLPgMvRKjqhYJv/BpZbfdUYHHken6QVo
rN2uXtNsoBKE7DDkP0ufxOvdChZrJIgfhxJVOXioGyzMUQ2J0i5vHiBs02IiP/Zw
LshfEqh/fxsMRdNaNyBkQ2I/70ZyRD4IEHo53q2agOVuezapAksew33uNrM+8v3A
ro7J8DSuqSEo1w5FO/BA4fP7kVsOfrS7UnFbUzw5AB9g3ciq5ClJg0N13PAaXS8Z
1iKrWpF0p93ZkYO8avokEBfvsTn5F6PA4wJKqspqVGyh/FJRaRuvwg+4HJbgDJkC
FTwSqdijN7j4X99ZBlN9UnzH5DrhM6F7xPUIxAaEL1fdBSlA72wtvI8L5HMlWBLQ
t5zjeQ+FaeD6hUUsInZ13gDmSXihIOq/pi/fpL+/3kVYWZ09sbnKr+2I6C2owFAz
9USzDoey5hzHl7xsUNxACWUfAoTHXGfcXmkmq7QB8iBNP0jIqhtfLdVwJ/QclA/E
VwQk/fRJ5pEwKpvU0e5O0B37Cc2xvuXs0TlOS9NgxJamJBhAP9yrHEXAMQKJdSet
ZzLgNIb7iGyl52ReueQqEMujWW6rdkZN2N+7ycMEWOfotwtbQSscePp4jIhOG6r6
7yN2Ze/8Cnso8lweWTtoKHfUFwYCpRE2BTKEMDHFcl7H3UOBCJLknseFPK52eF79
CMRRlc7IlL9Vvaedis1pz3rHqFi15AlJra//9bj42jprIni1zI/t/stLZ7HjE2Ny
41hnoX2hajfI6zk04l+xeyVsqFwC6FOil9RFoCvV8MsXWwDCtLYLVdF3s5n3knmo
XgKq3hwYqTLTxl/wjTc1twwGBkLgW90Rco8+L6fJl72qeT993cP7I1/dL8Gr6Amf
Ms7z2fpx4nX8ftEBQYx7a79g6zh9T7IQiXoaTz0JWlNRqufvnNuJt18wBG+3hbvr
B/rypp4dwiHZOV4glzE5CgQHSVJbrRjk2RyGhOQ7NZId0AJ8u1KFohqIbgP0k77w
ibc+l+b2wNJGcGM1xQwUZEC3yYq6fgHOlos+5JsY412tvVXvqERGCe0gPxK+BXv0
hdL++sXc7wNHfaSCTXTGqyZaEZ1gGr3miWKJ7k0LUB4wBrNEr0ixbU+NL+KwYWbW
pVnUf1yZi0pWP6BLan/uODAirW06OtC3MCGcL37AZU5+DbYQDW+kJtutQrCUt1hI
szLzFl3OKOCElxm2jgJ/yL9dBEgcV4HAKqkJ6Ovnexsm2z/6ZZzDrda/zoU6jBsN
COedVNvcCyTRq5VGArv/Jz/NomNjn9B2DXhb52kQA3AQuxJhAebjqoyiFkEinpnW
fZE03r9b0ouvKYUMZ0VMEHaD0GIRq4jezG/3F+DV99mmvh4QJHsLVTt6sUT5qNCU
VzkXs80Rx0mmCPXUyLGU6BDf0ojynTo0bdRL+Vb/Ti4HRTM5l9oGKed1GJKl+7hR
U4y8+Fb1RojN8bl+VtvXIPDZVoO0zfl9pjxBMPCRvtcHQo+PgL+3vBIUAYs9+Jyk
qevTHMZZ9w/5poe30x8iZf4IexOePB9uL0sGwzeI45p7LBHjWDFkKxAljmxxYTke
sBtG5J3Clg8V9LEI4deCjLoqzogHAO5wcdx+1xBUrBLgDJLceXOlV3C3XHy3iLO/
HTzjU9K1ktUlRIHYV3ncZxjjQupuvorybIsxWqBJvTci3DJ4ikV1WFgdS+4+9iS7
PldhwobF0eZiRHrdTlAq3bHXHpzQZUBMIMea9AOMrqE71yjcCNBvJfIagGHi4VFb
XCtUVpUX9OY9IF6fePZaKMd0IjhFXrmjO11tqAdwKsavKVu9CeKzX5Hp3TzZD4cb
6ZyAeQN26qp8zrmrD31BTp9rsnUph3f+PEqmkXbuOKUCStGK0GVv90ElmGEaXHlv
1Eggq8X+oeppy7LsYDN3ZAAKTlbomNi2UDPBWdhl81RCS7y44BSe1qm3k32TJzWj
gQYGlLlclDNmoHtuVwVqiaXzsmS7G1t+Pqk4z4sgZIfYFd2zK906Nf6lEJ0jC+kD
LggP6uS4pOVl+mdjyOR58qSq2658XQTiNkq1GvYQqEdZUqqVN78s05LB0CN8+b6v
g9vR2wup1x2P59sn2t/q+YSYPjoN6IMk/ErxnQckXSGiYdP0N+VIXRe98CnCNaX9
bKAUwQFaoeWr3zU6lwxfaXb+lVeqIWxH4Ns22Rrd2Ht6TlSaOggCdjoXBJAPMtEV
xGWkyjlgKphwd7jzFOdIdxuKL7ljmvbzQkPpDKtQQyrxWg+HpdeC82uX8td7sdX2
Vs9DMFlMGQ0YWG4wfw/d02NKVd03FBcEWcV7AXxAjVUA+Hw9AEJUu8dGQJPkB8r2
gz+KNk8Zz101cKDNkxCNjJfXuln+No1uAo261+glAIvyCknxWcGeeg+s//Aws0QO
EX8U6cYknp2Ux8LD/WD/sQQ//q+Gyvf54ffEMkfmXmaAwC5TEaYODyVr1Tkg3l5d
/7622t0rvhbNcVqGL6A5Jm0Wby9Lk/LjsKTNXLeOuHECAzHcgQoGpBt7/MvyJVQj
svjfPL6dhsXAXT4aa7HzxhjbfAWuWu8Nu2zXgd7l8+4p1FzVoPDGBDCKtcEbReDg
vBbe41VLFNgpk8U8eWrC1W7sTo/fK4njU7TctR3FVmBNzE2Sb+B5av73LvWvb4UL
RcVb2hLdh0ACBvJU+DorKqjJbq1AMJgtzp8Rxbb2RIfn3Yc9jzV8aLB+TBi3kUS1
PHtqoLXu5TriLUysvNa2b2d4YxSU1AwgTcfb2rlK/ePzrEwBaJGFSg1MXYV6M7Yp
I9mv92lBTzoym6wmdJzGU6lT4VBseg71sYJKjkcO7hw64uT/cppz1P/q5EWg1LQQ
z3OOp8ZEsNqIOolAnB4AR0mifIy6WUQ3ckishpHkaUz4yP6spDPr5hdr1Ie5cOl/
bmVNOK69NYO/nKvyWsjYEYZ9SlYyw+6N1RoHK1RqLu1PPxxuPDjAazDugXb0xPBw
h7ljjmjFw2zm7VDM5i5l3iJpLwZDp6ymao44AQayzyl29ZTpprYc2usZBGiNEjyh
E97Rsc6t2/n+sObvpRbR82QZzK9KEhnR5hlB49SHPoaozQ5jOxBOj9zOVuFHFJFy
GzPJlD+fIr7TljDdk6JA3ZbGiz7p6oaZWyJKYQrZoy5GI9I3GKF0depQ0UklV4CS
ieURnyHBSW47jPKyigjfoLY8QIJ/+VUqhEfPVXFE3b+f8sFPRhFWrqJYthCmze2q
K+s8jipi1SqCgTZsbAhsudmvzmsxXiBBJgRIRmdS2FkxWu63enXsk3GXRvJamL6x
xZ/DV/2tY6Ol6izlGqYaEbf27aHklnzVXnVNxSUwhQ2l5NSFepb6IkqX69x++EJa
witlBqUA329+U0XV9Q9/0DG9TtIRIVyR/iR/fL4pK1DCcDWvoKh1U2tBTYRiVTOI
6JCIT8238axJAYhZL9y+xEsmkMZ2/nL+tagbhDj1z3CIBT5KnwZ422HYugkb+NJi
VuBTCJmaA/MpwreEN4S4Cmxb/MZS5VtajB7bSQPEe5pljQUiP+TclkWFMee96DbL
r83YELhIa4Jc5inKDLBHilThVjC535oVqk9i9ab66CDMSqPbnB3+2TvhU2kb2afT
L1/SpM/9Yt29wzY/bXtwQLWHyXgDJgBa3nSrph0E4tkxkamJnBO4WyJkD4u16Ahx
jYGn9p9Obw08Gis2WPIKPlLyWyiWjxXnHy0a27Q9rC7bGKDU05VWEU7AHTPBsYNA
yKzV4Yc3Ke4t5TqdsPcReuOos1fZ6bZMJhqVLHEOWxyInZReWVeEJzri6oqeE/J5
S3Zw3wxxwnkfYPlemTh+7e/S2l69wRAihpAvsqiaZGen/kGSp+B+lvS/f7pZx+md
AWYT1tbs0IidyKGouU/xlLRjs76UkG44MvHle7QT4H6r1vomueYSw6DhM9YZBjN8
jLPe4CLrVlLlhKc+b8Ax9IWXwFySiWp5BrFU8gMjIUZV7QZrtPIRIukLBsQgTtRi
Zp+27CITc3Sh1IVjoh1fLvb/9e1VFmWjwpyb7LYqT5eZmQuB1ysYM/4utKW2shgc
ed0IPCTiTiE/YHRsPXSQF4G59PgoGjScFLDbGQFMA1Ynf4RZiUhqpHcDLxW4JAlf
+RkrSSsKW4CkAT0CQ1d0hK+LUTI/U7rcRE0HmyyoGumiN3DtSko3Ep0Go7gEq2A+
5mSRXfJ+ed0+ko0ew05N5Cb347QlqIvDcxqhLqXP9NggETPy+lEHZkvkXj3kYn4o
njb5ZsOZpvYQNhbQOy1NGIsDllYo0aAEKfWBjc0VPj04no08WFQkhIrZQRYJDOA7
4meVSiOIoXesWNGd0FtHAZwAxsQhUA0JIQYQdIyMNNcTCu7p+wdzXx9daUGd4Fyq
/1EVKKhEDSiwAP8p2zpz6GsP9L6J5fsDmT+K/s91mzvxcmOzGo/OvNxPLF+s1GFl
yOovWtCH6spiUB/CT9jW3ngcxfh6ytbcP/oZFU/5bIyCxCMbE07P/WDUwWlsOHY1
vJAxlBanfOzfcOVRMcd1r11ePsPFDdVMSnhLdu0RBnxliDq+DN5l42n9rkqLd1tx
FGD9sAFiJW5fDiVDXsojkrqMUuHP+JcEZyqb9jKZaj9i8lM2eHH71Bc4wikN10co
Prrz9KNBHEBLjgq3EBqFPBwDGy3mOvUkiTxeEs0AHa89AMGAvNyK49dbEuJale8f
Q62Qb3Oa0UM0ThH/cRfpKHPnmPfVF+h70hpZBpqvdXDsAEo73rXeEt3n2oeR8oN5
9MoMrZH0NKDwC68sey15FPKCYaEvSzoMkxRnSi7ojRxYP+pnk6yG8kkMx+ZNg8Km
XZ8ggCo+GP83d1ZrbiqcPb4rBCeNImvqzrDLUhMJmtBenBIormuxZnDaC6DrDpRe
kHM6tVf9jLjdJD6IqOVWjmTcvZkdoYjF0pNIMwhUoOzpzj7cXNT9drkYc3qnpNv9
24TfEm/UmRnBQGEc1Hpnxz7ag6ZI8ASjMnmKLVT6Tfr5xn5uUV+IoI9ZLHk0kcJq
KQodra0HyJjpd1A0jhViYogSds13qIK+BiQPufdiP3UnCXIarnrXwf7s3iG4JOgJ
ehIAKxpRNekGDZZ6HPhQ1ZfCMOv7LoSO0m2iP9o1WloCWOOod5UvtlC2R9hFYva+
KdIGFFN81X81yW9Yk+wIMcArA8KPcqUrnqq42cXqA0qFDPRIcnYR0KiFbHzp9/Sd
1qDi/czKcD2ghQs9fmCvVKaDFZV1C1hfP0YDfIasEX1rVIjAQjLKlBBv9bL5zPtS
FQYqEdbA/SIUI0K1DhC/dMyMZJ6vSWQOY9Q0goYy3qit71bbsw4xXaBXr2EMVkTM
T35cUvjwIwaq6jZl12mVTgtvhjYeqFfBVLBw4dbpG9fDwtb1ejt1uPytQgSVctGH
FlFy1phLNVeoOC0UDsvO0kxOiqDj08ZyyA1yEEnkDJOYh9h0OZc1ACXxHw6feRY0
iIpzg6w6kUIIi6nTSlib5E/0pY12SBD4UPaRrfcaeM5VEDi5pfazIfz31pwx8dGV
4aNfwnyvzMA10BhMJECHPSeHYKohiYe+eiAf7vaMZ5pQSu1zk4M2+WlIvyoYFdNY
D1lCKChKWFpHjUyy4vgKGCGH/52KOCTInCj85ADb3GWxKHYlGS0VOGtYF3vPJJIr
l5GrboffzfVmX7C2asqrhskX7vvIvjFsIPGHgW3+j4OnZl69Pqm7twBPDiveeP4q
LeYhMjsPhIEqURVeV7LhzHTS970SuAZQIpzuBvZaCbaaW9wbZNFiIZy118rhDJvx
4H8DkRlDtEl0niwHkFjJRqAUpjyGydzWiIEWFQssY9dyuarzhkLf0vEZ5YaNwYO6
0OqzebO4RHMtcv2tPGHALe8fGRBxCjCgi3tKEVNuBH3JqV90r1jdLmPRJviZqkxs
3sG6FLoPkZxyuLCRvQoGJE1RcCCufyT/YSTyCvqNVzxeqBD7Yw//huZFuU60U8nE
4BCVJeBtqz8Gm5L0awtnrr8y52IUtq5U0HmTwe35P4Y81LhEWY7/uUe7z6J83c8S
eDeT9vR7YXIJOBUIAJTZmtNCM1gbyxxaz2p/ntp7e8LXAGUJ6+m6MKd6N+/haw0r
+AEv2hnn3iMtvaN0Bdu2VV65HBrKgYM9phM45aQvKpjZeYa3FordNWLxCF4t3ZIh
Ih83lO4o7HuebbppBL2RE5N0+48iMYqVNt8D5VNGA9pyEocMqB/mzQrpQ1L/wf51
5gBNFIgHIb2Z1em7df5pzix9DMLkGrdYhyImasy2pbiloNb5ShAIKIKOv0xIMTi0
E1lFYYkW3PzLqVnw+MrsgsrJRBTYg3tWRVzfDEh6SPOdbQDvqtqBdRVAhIuGEj6+
+UumFQUYN+1RLq68XCIho9csQ2DJqAubcqULYUs6fhnu5Qt7Pmr11VtWbGicDkkb
+5XyUieI9OAwA5XJw7q5rzQ80kGv/Hg7QHUdTmtAKeF6oO63qx58vYKYmEpPWtJG
o7p+JVpLpaCY6jSXgc7F6HyChzov079MHj214ohlLX+LKkVrpbO5Zeoa+xcyVl6Y
49AscxcRG/3549e4u8VXgfEIPJ4CGJ64AEv2Xvajoip5yzatXFW80SiwMK4hiwDd
AvvBbqGB8SZ129qJBLDzLBeFgD8vinnEpINuyOpfxbQYgOt2OX/m538LJJ3aMogq
P0c6jXXFvgFwYN9Mjt5+CNi3zOa9syjzdzBynbWiL1QYj5OdnC6gc5QrVTJe/e2X
CTB40MlISQ9Fh5dZFTk63n+BLhn7n4fUCUkdEees+ksaFax8d1H9iElkUxTBuSEv
00BofhrpT02Kj2+mVSEcVRd85A23RGakzfDHm/DlJ2ZyGKeMUNyKW7w54B305Mou
iQbCwsOVQfjxwfRXreq4RNXG2F9VmhFbXu4Gx2qGcZ/9s33msednM191SUmpUc1s
kzgMs3hwaTkPYa/tH0OOjWLIXE/AHsbLTPVeOmhTvo5QF3780U8ImnOxNGnldC0C
DJKgLXd75qv+gGlDdj2PFvR/Vu+uPNnNeUn7kl3fbLNP6G9eQpW5bpdAa6t30Hnm
vsIfUW+d0wfuQqgGSyHBWwIANHT61zN0Dap1SGH2tnv3Jl6+HB2ry2GNknc0FKyY
AtefLn0hSLB892dlE9MgaoraKyxoEoyrGOsH6VkkZDL0X/kheTZ24U0QQcuVuKyD
y/Dq0tb1YunxwBSJg456AlrE/yb44CJCrsKiJ6VIdBTloXJHgbA7v/teMbphH3j9
JnCNE0l+izOETHkNHX6gLBVIfjfFyHW2CJ9+P1E5e39MuZW383PFcvOW+LKY3UU9
vwDXE32XngImPvOQyJaaLaXcL3Pi3YL1LdsKIJ6asFPUCXLnaF8a5EDXJYrtkkcv
9bAqwz4RJdamxTgl6SpAbF1dm6r++1vJj4G7sZrTmTkH9uGzgxQaMZhHftYZkaGu
bWJihbRnDIG6j2SPfBUOeqMnHZO0iI9u5GB9OarzWKgc7pBZ75qko/fRFtEJr495
RiVziqHeFB7dkLQHmQeGNVDH22ZC0ijhA8X39HK92JPPkHKyLk9vdAUacQSS+sgg
3Ag3l7YUzowH9bB0NKSmshS9bO0fB8MDovmyFXP6s/MVoVGLvwF6xtg/mvN3rtK8
1H+0yxJJ2jS31f/HjLeHoOtHp1n9bdsZYHLkNYjeFYIveDDDx4ZHf3wMSMJ2GUq/
nmjIcve1P9qsEMEpCU6MMVicbWEOEVrsMtSGNdF/NK+P5IMNopfvu7Nwdr2lBIVg
uD/zye1QbfNcZhwurT7ZX3FH2ph35F+Gvi3KFOWzmkr1b65CYEluHeWonSQhOn/V
tdQE/hL/TuBMZiWDaHPwatI0KKlWle6anP1Z8yqrZzGa6FaC8z1w4NeeW0GD5W9X
9QnH9nQcOdv6scg9pIqmidzVDg06AKBX39/h8Vmj1/DqfbiyODppt/q+SUkdQ3CE
BlUro6PKSAAjTyNU9XKNy8uM1nlt1O13GuFmohXkRkJgOWMZ3GVg+2gts9Kd7jGB
2eDZsRzHIC7aUwhtcLQoGOMzufqmn9CppJ/1/HWgRSFrAnA0/gUhMjGgUez4w55o
dVEvrQuZX5Hm4sNhj8dOM9CmTxeBA2XDu7Yyj+dxP7GarYVMKDMMe1Zy8yY/jiWG
iA/8ft6E5EByBzxZ/+6lvxq66E963n9fI4YLx84LwHBCvmpZlORf9MY8nEPRyT5/
ZYWcFhg2PF6PZ2cqPBmvr/6yuTRWemHXrvRY/j0Nr4iV+ZuShtCzHccATDtJyt5J
vxOOKSyj9kMbBei4q7BN+EDuK4Shi+MD/hgUtCX9/q42LXQBdQGQ1S0Ib5jRVq9+
8TcS2n6hEHxmb9iP1xGJJPnC+iBnnqOR6+I2cWdUW5O4B6xkQND/RRvReMCd9m5S
ahTC6B93EfffyidWjsUemP/VbwxoKTqbGp1qB/Vx+OXkF65bOH7DQLigLQ2xtCHv
vlXQ5O2UqZ2ZsLx/JmjCm89Vt21YRA9aU9/KdzKGdONjcEUiSKNmvqT44SMTp3a4
L8mH96yTbSSNdKzptDoZS/9cG4jXyFZ1zrOWZHXnd6A/VgdUB9+onYs88jrBR9+5
fsdlfN/rCh+vvTZV3VaIjtrrs8Iu37O50HXQnp9Rp4aJipJ6zyoR0aaiQHqyJm9F
bCLLwc293Pwa+JRnmUzutBlFMh4lfwAI9MGvygX1ezc8HPLBo4gN2vpCinhzX+qI
7/HuwUHcXrMOtHHG+BAYJyGmybCk8Xf2JXwjxCmGe7tASU43sTWxTsxqnZMafdOp
ZYk2RDmZMRzHn4hysEJigye7fCx/CZXj1Va4fuF/cg4k0S6JpIa5nJNU3jT/uBrr
w+2UYMu0f55jbiBasIKi66nwlR65JKidrGUgxqU9zZiwcZUyF3l0wnPHkAqyJo3g
FiXXTYZUVoV6LUpoa4fyvJNImQapH2yp1j63ZUSMWT5+CC8tawzFthE7WOgwXg9T
UfTtT8ItYGeuVaZdFqYNG84HVgHVHINU3uJpgmlIjN/ahguBpLu8IZWkGzI3dZQH
llf5Af5vj1/onRQuxMURi73uByknP0BpNjyQc+sciVnghWaEXADD0MJXsbHDFLCf
c92WU5xlbUuRYi0tw5p3vlO9fE40WN5/PDiYFbDQyCsoMkSQISCnr0cZ9iIJ6Vnu
dqpZ8a8FuG7O6LfzHypX8A5FuLxfe0r0L+SEqnVyQn6SMD7cElnnhN2LH0+q22jh
CvJh8OdV0ZwjIks2+nVPx+S7RXDKABAw+RypWLgZp8U4sZ2PDh62N9rvfoido3Fq
q0yALI+45zeGWr0gp+tda+89czRxwt8B9EeEvIKcz96NnunRRS8wosGm+Lc9+Tsd
+K0XPWdRvqkOQOaxfJ2VIqrXF9aJ2+MGLEIKp1Gfz00TL5wcLfO68Xtwkf/mxxj9
m3/bFeX1/GUcEpoMP9kxVwmdYRbKOF1Rrj2w647zG2Zndt9zFeTG1ZwwWGpac6iM
CuN/Xo8e/H0bpdgq3hPNY5SLtNlXNeHH5l5DN45NYFYMpZVOPnW6CbkalXKnJZC0
7JCEE4Pntj07c1PnzpnsMOpimYxynht4lCHNz/MSPKCpi57DvyqWNvfnKc/XUmsZ
cVn/W8DBj8yBcnt9Skdx4CHJxT/DjGjKV0oOmFXwMtBiAqKY84qicrMYFHQEHq9d
QXr1mfMbcOVqv0DlT376Db+psn6oZUPXFKzKRZJMbr77t+YNX+UwjEYZ7mp1XyFM
NtQxpC1QtWdkD7gP1UCAwgGv2jny6QrtG/ntPQz1bzbU1dlzw6ET0OxlMGybmb4H
WLqmo7I4QxTvhsQK+FfuiIZJB/NkNApQSH982nYrKzPYfD8gTS3dReG5gofxY4me
RS1Y1eKySZ6DWG8wA66BoCsJJpH3/28cNRT/gr8NU0EzrGgin3ixQvAOo8dsxzKd
w3SZD1TY6xaYQlJEwLKjt+Ert+Wgu8eQVbTHdFyJY979Y9bnmz37NgBNhez71lZG
ee3vobnQOD8+QRjs8onASXqpnJgEUaI16a0WoVAG6Lra13SppnlR6LipgAdPzywI
Y9QNUpAJ+nH6FzNxGSLpeIbjAdxIe6CucwV9i5fCbfv8MtOLCBGZ0x43SBSgOdey
tNuhWLXYHCzHxlxxtqNFgLi7W25flodurjFxWLfgAY7qEVUC4c6K7WW+tZ7my5dt
rMY2YatbiN1p4T/QKoOG17a+ZkFVDnkdA6N3EZmxXuTQ3QpYVwsjAGVp8PTZID2a
TRKK0WFIb4RUGkn5eifG6+FifLmYuodnzL1wK382szk0jm/kU3PM3HAezMVpYl7r
w4+JcvLVYHSipIpbfjXJq0/C2l/ELiO7QTgyG/nkzvrPMTKNurPbvLbE3A6mSg1G
2jxdwFaJLT1HsrGGpbK4IjpgOoAAmoYIttt6dwK0Tdvkdf8bsmAKOuxv7TJ58oCh
sh/hJYHF9iVvdkKJODYqM++TFWZPIj50cLWWQGPTk0t4RVK4ok9V7TaBqiZGSRpc
owdB/SPiu3JAGJq94vOL9uv1kAkM2+ocOksHGdZRxRDeiUEbhPKVsnugeXXtVH+i
lHR2t4DuQHSnHIARP59gwKK4m315v0ElkUw7mB56dt4MVibcUrou0C8C7RMrL+Nl
E/mTLGop7I0Hd9P6Lyjg+kSAHisPX14QEGnOsp8OhFvwkcYw9oA8QiKYAUl/IiFJ
duliJx71KIP5C1sbmTn345QmumoFNk7mt9RJHNTFu4R8BBHuG4szutfCl8QTvf3A
ihXw/4F/WbBqudeHDSH0+gpqAjFTZTM49HCY9f/upl0VwEJyh49DU1YpVJ+6V0kr
EOCbzMs9zFS0WkUBPcxhBxAcnRMXTM52dlrFVGnhzhb6oeCe9fMpnYg7pzhfnGqB
DWS0nT6TOmsCpbewqzqQJVwIY6q9ZGSn2nrBJ2vR2yC6Y6bwjWk/i6M7GRan4A6L
jbQbEuSuG0M1lmK2PlLVsMuDMtB4nHlnm6iGZJ4YeEmJzKSPG/Mb2Qm/rUiALKJg
TJc2ziYSNrGEc/vHuZ31lJKunE3irEqJ5p2+SCe7Le5cWc1se+BF4ByCqrMEMlG8
EaskkGgURD8MVkdJY0rKBb6jXURViVAmArhSRmCS1laPoRs59tTFMx0AltxhmBev
BrZf4KiPIC1BeD3X0MdgBYARR1guQ1VKLOMcxx7B9n5246j7A6+ae1rwSS6ZVjV+
7aFrfFzmZ2HlObIo2gJd/Nudf6phZ4+PO1GpCUw1n22UQgfP5rS67BekNwcpJs52
usrmyTjQusLn2192jlC8hucaO3gRXGfRaAnu2c2qO3QB5hG3oYiUTkvfXh5C3dIj
jcp5+07oYhOpdkbIxP25pkm2nNwoVK4Z6BiGIr69Uis9STUCo9c3CzQEA8jofSUt
fVDN3wSjxlK87ssYJGwcAii0yLRe9kjafCd39QJBb5lko/c6uTWGmKTf2FEI/d7d
VdvFNlmNFvqtzDGTfQY2pvTGjhbDL04hkVmQHyBTTFaHVGk4cfGo3awsK8Y7gwQU
E3ah0cCAAsb89PzrfYFCYF5M224vnpUN20thZLWYfI8rtZKlCSuueNNx3hTYmDVv
Gt4XzRRWdj0zCmQzGS0iyJ8OVsCVUEaPqgGl0A/sIB8XdIykLmlM5OOJDv24cgFv
yWJ0R9iW0QzaQBV/iMdr3tGPlUk2dQzzWSFuFEktiNd2KDbvAgSlIJk1wyWlEvaX
yyNGfhxDnaPqxl4g+MJBN2wCVRlWY90xkTIYK8ZVadSfn+WXs8N2gf20FnPYVU0N
JPOLb/hinx9zTbYzQQHxs5Yv1Wmv6oLMwM0xAnOpjWcq3q9lFS2A4lUXONbrgj3Z
5hm7kvllFTZitUS81414mO4I/dIrkKgixhJjZ2AWLAplife+UOJshPdAT3+6b4y8
hVGcbm9ai1uOjeevdu4mLm1gvhAyCnJFHrh4bIF9IglkZjfHlD+4UwcUCklo2OIa
ncQKdygDpcxDBCADE3vZTZJmaTSKxU11j3zEU0lFDACOgj4YdzNaWTkVZke8xnyI
zCqLFf4r0O74RgQ+SPQRoj8Iigli5gyK3nPjKlHT/rGpU435t0RzG9ji40dcomGJ
FXD0QZJJYxiuCoKxGATWNPYLjdp2kWrYhKn9bWvYQCsAqXoGeRmXGERRADH0eTY3
jjNRYreWguA+YNSaepQ5VXAbD02rJSW45QfyM4tZX4sxf9kY2O4WYLFT95ym4nvY
tYj7y4ccnO0Ka5YM6Sh2jXfDk+u7Fk1L7aXYD6/KRgyNrAzXZsRPOD/6qQ9Aisj4
UkoZDMWX0jVNXi42/rmX7GaKeXUfymfO3a2LjRMV0Ne9JQTt5QjrofLRQ/GDkVN6
s+blE3BQEKFlRpRXM8odVxxdr+kqln8uvdw16Pyxl/FJNJhfW1TWD+zg5HfNR681
MKZSHUy5RNl7ZFWKUTnHqUfBzG0eLTNfZ4r7Nqqu+uN37KJJDIswZZVH0uokvRpb
v8vPLhuNvdQVlHNXSV70h2pJMK+A4JqUevIC+1+WglwzxJPNTd7Y2NJUlvmNy4co
BW7GO/BvVc8gQeg4xjxnk7bDG30fZ2TH7WheipfKPCYDSFUt9zM6ySubjv/Vh1x0
Ui/NVzWgDlgeE0MEebmRMRpujLowjWrQbcLXr6wQjOUhRg31JtRZKsmuk3I9wgvC
IlJh65grOGUeig/qX5xfts5WeuElekKA8T5IAI/Wer/JWAXV2UPr7Z9IUkpwCB0d
ZExhdxCMRVUS0dsbJVCXPiwZNBdb5RshG4vXahNK56JDgiT0O7E5kKIS8kcc89EA
J/B9XFa22bSdz7g24jwJNb8n310YiB5GOsf1DofRz37FUNbvMHS5CfvOHYOnqH53
vlKx7lIlkqsjVqtmMaWL+fn7VsIr1stIs+08J0cKnJKCO197GLB1LmDnwDaANmp9
G6I0XGa5V6zqgArvaBct0O1LY7mj3JK+//0hyCujN+BQ3q/Hg3uK5prFdBZhXFcL
GFw1rp4zScsaMKfCmAj+VwA5+PoaucWsBUr17qRDlEDIhVJ3flJJeHKt6pj2X3L8
rf0Rnu8EZGrO/usH/9iCn/kDOzPDLU1dXsO7pipcXnheLRxPS4Jq2C8gGV8MCG0R
KSVPcvhXf/tiXbuDRKKLMgXR2tljXugUYsJSDvV/IMLuXsyyJRVfITZCTzXycSaU
qDHWB5SOKxiN3ztBfCHcgyiRR4f8+tZWFCOXZA29MEZx9B7A+JC1nxRVLzQdi482
9QI/90bV9JbRd/Ss6DK86ckVUjG9wNyn2dQ51DWdecGoz2lMwCSt7F8iJuEZwcXC
3GNy/TrGEY0xsKFw9lfdT4F/TcxQQCHwfrMX+OLl/6gYc2qD78QpRbF7rMxCYqQ4
oxtKYa7LiF4vdbT9v/3ETHas6Akp6GfDXmtoq2HQaBGMRP+C8NekwVVhst1Whujm
9pUZsszqf38/BG3BeEkdwHfZqm4QRnY+d5aPjHGc38IN10n5bakTxT8XlmN/L7eR
FP+N7cC3t8RVBHV7hiSGsE2ekDASHvLYn5esYGTaXvntaAKbEm9PFV0wkJJqv2G3
kx+W6rv3ImExac7b2oMlcY3T0PVPl3HjbVYFIdRUbwL82WTkomvNRiCugkrCvwtt
0xGnp2lQ8ZxxW7jasA+s2+jU//590kMY2u+UDYEcZ3xDLE+qnYXc5HqOVtYFAHz9
qBp6Fy8MhRQv2QFCcfXqYL1uWmT3rEqCZHTk52EZlCARAiwz6LuuDRRlM5rMwHpE
zpCkutk2A2M+RQucfhfdGIo4wy8W6jtjWOd45xUyBVM87CivVRr+dXStOdiVtYUd
TQ+u3QUyx0JweM5Ttsc/DpLUQdJf7v9UPYSoVzdhEMkXBGyRMPgDgo83oa9IxMu8
elxMTJzbduRoJkhTDDdAbOJwFGOCv89IydL8NEcf7cCOqO9gclgc0Zl4njGApStE
Pnu1BOTD4X3fPR5gS3Mp5l35ifKTurIJZROKoB44ZL+bxYpSNVWNpe1qXF+6AiBt
3zgq9tY2jY4YcjgDvaDTuAItJf3yte4QAmCd5HiTDKdpvqcSnWTu5ftm9egCo+Sc
dLy+rFH1rhPdTBr/FO3cqJEj+hHQaPTsvkNBYWFE8N0ZLwQqRtfoQaRQvtcFgAQX
FYtuPI4Cfdh3oKzUECtamjay/+8cTp+T9X3+k0n0W9uLIT0PLTwW2+tfwCZHNiMR
v0br7Pjhemz5uOnmd4G73AytJSN5HLqIzUqdk8cw2hY6joaxuqqt872tgnvpUvWA
ACVLRJ05Ifbx9I57Eotw6iYn8EiZK1+joYUg47E0CFISxLSZrS4lDWVPEnqPDrTL
RLnNAT5RQEly4s3yeemDXIfT9wp1O73Am8Xlmr6NKPw+MF3tdBGEp8ldzhgNOAVi
gepBix4yyQlYigwioc3TcG9jYMif8SHm2TfQr4cFaXgDgDZINaUlpWN2OSDeeZUm
qeovwK8B2BeTRwa7tXMvxadIPz8EzI64rFOvE6/nbjmBQQJL+qUanwWatJdDDYhy
W4LNSJ73LEybdJHT7Dn7ghBzQBBINd8qwF6qtBEfpHI5jwO8rrOGtjUxl52oOCMb
ODKBm8zP0VCzzZroRGGWMGUIWBc3rBNDKtxkiR14Na3f2qWySokKccHoqCsJNGJn
2TLPMwqYGjDTKts6cclXXPKb+qbEOf6NmVt2F35j1j6MkzXYoJd/xwg2tW+7J3u7
rEow4l1SHFlyJqSDY6s72twyTl2gEQXPVxcf/dPkd+JIdpMIZZmYQUBqYEC6eHn5
qpym0tpnrs+W0+ROE9q3HKRC17yjyv/TJpkkRCQkrxfYOQYh7idJtl8FxqC0/s5t
/BHDhviU/p3JII5KgFaHrYYUDhvYRJFKXQkf6+eRXxRvd0EMcM/cqMTeGhpkdiH1
L3HE4Uwaf3Bl/n3fVQ/lBbgwZKq4qL6tpmr3XdzAIrQDbLUHR3ISTzk7wafxMG9E
b44EMxbyXfyCgdu/k5bW6w/zEkyclDBsMKJMhdcL1WeCAJG+QRkPXs1EqzkBLKo2
WPc1gEV2ivXvyIVxfRl08gUpZFii2tu0OBlJDmJiSSQ+SxbfRpmz3QeWtKBRwVu5
wEnMFvCIlL9VuXad73itWTX6hNdiVWBnu7BJwViR+kKQ5BLvAF15pp3IUBCHhnIr
DpD8gjr8YEa/WQD6PGMyhunZAuETP9sH7vC3UrAMhfOtjlX+cbT5mW28ddsWDW4T
ji41mw6HXsXI/cgJ0Zyn1AgCWE6cFNRf3HjLjVCx8w3RaJIr5vwqEkYgZDP4tLue
Yf1YaQuuqbvS0wHbpRwx4FJCzXcD7erfKAC7Krnq26215/jq9lWYCMBsJKWGOAjT
PtD6VUqe+gJn6ZzhyeJqWY1WhnHUz2hdNYMxq4aC5PCxL1XEelTKUabPuh1Dfm2e
3r0iCQU64wxtIHLUEJbf3vmV+RqJp5jlIkYgEor9jteTxMTnUtVj9OGMEW5dv54y
Mz6wQdh3H4ZT26w8xXhz27trQDh5cmRIz7AlVoRKVCUXsxwZgWjqSwhPmiWc/AZW
DUIvC3Vhn4WHV1mfuTUC2Bp3gaO1isujTsf+qyD0SZ3eQMPZ35ev3ZA/L4Omj/27
RBQ4LQCQzDYgNV2MLqDFScTDr5IPU7vDYn/xF09T9Zh/4CwGM4wTlpeLKXaK9Xke
kzL4va10dlXvHYr/22coVuTTZR9GBZceaDTJGUxDTG5wQVTTY6XuEhsif3dnC0iI
wRMY2PUnxc7K+5DXkvk94/HxPQf9PxWnb2faFhPESTnkJC60Xyo+Pet3MCmSqgN/
Fwi0GmPrzrK1CwsDPcSi90dkaJ/afdHxFRCvK7tCpAddxmSViI9bcS6x6rtHiEQ4
McE9/+jK8EHhK1A9gBm3ugF4igePcMp8La65/RgzWjjN/5/V9fnC5heKnhDIm2oY
j3zgLqWHEaKmP+lGD7YLkUMsoLJKHjOOO6iUW0STHwLkOerqm4hZAkJZlhKkDnc0
rKkZKr6bn5yHy/UDcYYlvXL2IOTmzKZgCrxnUbupOx2PuYgNkXK6lqX3VsApn7JE
CzZy31ZHJ3KBOFwKhWSyuD1QsWzBUrPZLWVJvSfOlLtID/gsOtFkUz7eoAb4T9wv
TJlClTioIaAmLeZU1gM5jaMoEQHnoIvIxOHw+dPCXxa50NJ/yWPklRMfbYdTvx+C
h3PFvNDELr5zIwrIZjH2M/LIy5G3Vx6TSQrE9Z9gZGVUJjwOKbh9Q4vjVCu8PRd0
Zt9R+rXVGnerD6G75YfC0Cjq9U5WIVUD689PvPXlouFM+fnuv6jHRojbRIU73BKM
qOTKWvzI09yS7Nd/kxSDn8nvndydIyPlDgnlWOFNy1KgX4r1utW/D0WIbJaXxg1/
muE+lxowpVw4hekP/UckUPgeBUEBRhTA7vFPpcoSCEmkA33FTNKrOGBvLE/wqZyg
5tZ0B3JXTVDfV83Q+MRefCQiPJ44+LPSKgjWyPD2t6HMbqukUcqK+DTedlFqe9pB
jfk8jJNXAICPKEnl+ryEmfhjpRCv3/1rbtRS8tX2q+5bTH9fGTY14GIkXTNEiO4F
jKJ/33B2FMJfDl9rWIV2n8Tk9Iin7XspwndbiI2v+VfM5mGHYwNnXmZp8TSSgQC8
e335TfBOzYwFCNN0VS/LF86dfh4pwx+klLZLqKnfncVxF5+ZdbdssVTA8z2MXYJj
xKFZ9ROx9iMqLmIMpzujnI6fk+Y8W9SgydEmKg3Ru9hwlrSkgYWopflsEtztpXSn
/GYs1GF/slIvkmzR22LPGX/qVKhjGhPEijI5kgfW0FuW0BYnocHrWgaB9aHyl4WQ
gbBRJgdwthId9X1B3iL5Jb0N97WqmM2L1R3wGi6VvJhYlbxtAAb3FayHNXQrM6Ri
VSHP+qNO6OfW9Uo+VTjKt99RT9c8nKvIueQvHTk9M8Ux/EdLm22VI2dYy4LwwxxF
aGzjqyVzwaPuNzu7tJEOgqbYzVBkkfGiVKp6aHLKaXF9MKU5YhsuRec2Pdh/XUhB
Z8+3ewZSrRCPLmdUxnWX2n3K2TEVgiBUzStUzaKRZhVAaGe1Jd3VDKqVW/KArrV2
Uvc2L4Zijp+Wn2/UVrjdMP4MFXVC7MuyQGdfcx+CYEczjm3rtR/WCo1K1L5/v4Oo
IWmWP+sFp7oU+ceeIFIiSRdef2/FkG/Pr6hD2ZE+RdFm9qI0QGctIb+cKjlSdjfW
8WYWVNXv5c0eQSN4dX10LMdKud6iI7jIlETvpNkbHawotVjSICAM6Atpp8Tt/69a
R+jBtxZQv1W46aLVj49EFec3C2CoMQd0TYSc1Femq5WxcZQFaYanac2z/iS2Rrh7
iPxBHQp24igKQBV4lTwrw8nJv91Mx4mVBPvcbDCtIy5CjjJGKPZRCoHexmWoTy/u
nQqZKvdbC27Hngc8RVUXGL9olB3Z3+29KFNYA62GaoijC9WSj5T/Dk5GuwneJaj2
+q8hPnCS5T1SBBYse20zIptcuJHiZwnTmAcT50QAIIsnrZx6/lnipCSOv5R3SHS3
PwcDB/j0ZCa7LiqW2kOBKmd94Xr2jZo6/OsmB/6Pn+pehtDyusAUr64Bo5FpyCrL
6K60cTHGZ2oGlJTqqhrtCXEtDQ/xCbAOkWXUVYE1qyR7IphPKF+mZHSd2bPGpe6M
5UqgGItUYw8RfjcP29s92m0hHtWBd5Lkm1N84mDUGg+B+yb2E9XT8DY7bQ9pWWxT
MRPfk8GN3qZF0k49hCiZb+b5rVSp4uYgtScT7gjym+RW9YxIdfyu6DhHJkx7/AUA
6TpteeLrVdRTan/MaFpo2fYR12jBE0b5E75PfBPfQg6lIBdZG7N9DKwErw4XngRu
xM82irSWn4c/PIwxHpIo6Q/xAQ3ss9HwF6Juw4Fy5OAwx0ZMqJNJ67jc9+Vio3JY
ENp83Dm0vMCodwg4iCHJrQj1oSQJFPgpUIrftLsW0eddgylV3wLbcAFI68noASg6
UxM6hIEVGEHl1JTSgP0weTKWAlWCvWFtq3q2hBeYDG+XhdTrC7mYdxK9SyCEEDsP
du8/4EYeSA1HXddxTXVRU8L4Oa2IwipAQpQW1bLUy1tIn/hAhd8oP3x854h4o+Az
vSEKsXrwIGlr5D0Ff5HNfwlZ78x9B6RZCaT+zpGQ82f1BNecCWUkZY1q8LMnFZMR
y4bovP3KJajX8swCOji9FrIhAx72vPS9vWgM07pEMgb6M55HpxV88Fm7Tsl9Q5xU
6AJipgPUyBhRg8wOJu4m9hU/7e0asiTMD4VyKmPkxNDSWt1+8XNGL/YKHKoH+f0d
xc+tzpu+hVsThInxfWSLm9IdoBZX39jh6aFkRXGGYXAPJ4sOcf4B0nXa2n/lZg/5
SDc9DhVSGJQvuuTR8gz68XYW+zmZcfgzUV4eAHhIdrSf86TFim3zHYUZb4Glqful
FB9QXEaf5kk+ijWI8ACDbR4w41PxWcpg1BZMdI7mpTyHeAtF5Z9vDzH7nW9HWX7+
2Qawa/utLzl1jDxn2KMZ9ilZjiemRO3vc4WPMUorTiMfVQIl5sMzJBMzUuRpCHs3
2/7pNRn/jRDUup8Prpj+cHThDZwBh2HBYOhhN0N97NpYAyZ2kn8cUjlEruteGCg4
jRm8rjd8n/fDFCyFCBuHUXxcjZVGuKe623XO4sD9i9vRcC5MPeYM3BYGyP9dVyr7
Awi85SiCeh8KJ7GuvnM65Qi5wVJHtly4mB9Z8S/mnwOj2eW1OG1Ya4HwOcTizz7+
7TXpuP9xzmDaOZOM74TCYDsUWA7DY9FrHOxoVPFX32pLJjsBa9Fjv50ITu+CZXaK
MmAKAMh8tcWYA6mX37FVpAvla5Q1VfdxH/ZFLOzybsCo191gFPjnU+7RwhiM+JjS
XlgRV4Iz40ZQXXJayikd6VfzqbEKyDoxBm7+TK8PXKql6Z0QjpjhH+wcS0hTQckF
muozzZXlYFmd9gxIZVZZ3ecaFW+J3A0IFAtL958cqEDkJ67Aj2HRQK48HDblXnVw
bKDAm4w/8hKZtrJ+Z9w6BGEFCaHlME+47cyr7FvuxzFtj8xVxm1bHGm1wKJITii3
iijad6G/9nhKI4F6lBuYtF41BdwoQtbPWr0l6cjuumFurgo9V+1nKvxUEvY48gHc
gB1z9sZMpN3NKBSl4yKnhNFv3Pxz9GIIVO9DsvYBDW1mfjIRqW/BXc0WxdMZ/MK8
Oe5OlDJI8O4O7Pxaig/ow5kZveJy5VX3J6tFiIKmzGL3SONQ4jsk4KfuWRODsw9h
UDR7hh34lPgYDS3Z9T30VqdFfIUtz19q3wF2xalx759huwOMaeVMxH/Q2KgoO0Ls
BkUmtMUQIIKtfztZonlhwUatZTcfe7B+eYpFk19l/iaPujJfHuVR/y/m7in0EJch
T0xUpJ/XyEEKFAUORhyeis6xFbdN++f6wyTpmvXhr1RkQWSyP+SRpvqkJnEPFFMJ
C9MP4TRuQ6uqpzAbWuQ34qgZY7gv0j6VIBMe086+VDNHtnx6fkv8HVep0f2LnkZ0
ktxULObdRnhfcz760uZ7koNopDdv0luylFnTTgMuphnZvnS6eZBLj6SKI7IX5eL1
OnsP6TAvWpvtkvepn6d95x/V4xaY+YjaXYj0N3jQsbh1Ir+e9zY4mDo65o9fB0Cx
xPCZ2ojWE+291x/K7MoWiXWV9G0KrAew+By2bmD3GdVB/G1jvvdwQSy5bYXiYYOF
mszG617Zbp7o39zXigiAJdSlPO0lTOnCkU2K4cUyeQVJQsXDnO7eQIcOTkzmOkcf
mMPBj86L42vhofxqiRBs902pPH/ht06+hbJIabAIQttvNKhuzGK1qk/m3/mZCr3n
25+r6G+F9KQoeY9Aka8X71D1rfOVKaAGFYGmQ0w8OfXerIzP64TVOteToA31+/3t
raeBi48o7l6a1iTOf4jmoiy1adcaV1l1KRZ6Yh+trJEcG29R9LYqGVG3AAdoHAX2
oVhw6vSSu+NML4ZDfgBjXQO/EJo1cnOWTA5p6anYXYdPY27OGhtYNyu9dKoOILc7
08gzbsne4M/WpRkMzgMYdzQjLFFZQXB3Hefoa/BHHKuOnw5QucZAX9dIcYBBZdAc
3bfFyZogUTpGDdeHba/L88JJ8m5DA+EVko9IFSP4xzypZAMCbiuG3XpSGj40U0Yu
ih9US/KeN9TxB2RtaL4VXJ+qpgUhx+KCqrr37Jtry0dA3rXm8VvO8fZrbAFnE3Tg
l7Q4qzAorcMYBrngcv9urQBYb3ataqTeDfpv6p8V83qqDmmXymFwjeWk2x9NJoeD
+oHr1LUh1+lqWwwXdq9aoQ5Us+uCnNR6CatCI7HgR5VEHYU1Pk7owSaSlIfgA+dt
XjhzxVdgPWHoA0b8WrJfPCs5R+F8OwI9uMQEyXzlL4y5Q+LWbLctGZU0YEPCFjal
I1fodcVZdqkeMregzZC5b0gZ7asupPGJiA2rZ9BsC4DPl52SgfR+TIaNeVxVdTbW
3LfAoSZdXuLa9pAi5MXBiJPxpBZ8A7s+kc8h/qbP68D7Qgv9Rb/x6Gm1CickV3dk
POlTEp2DbJkRARtpAQLohT2TPFxcXGQCzZdm1WzNHMgoAnmVxEVPeCiLKQwYqPR6
VuGnwkDDlfqEbYGDH4er6W28xBTuJIdB5BcbzzlV9JnvOuv2HBvIkR1AxFUdxXYE
ad2qv9pWMAv306YHUTxuhJFY8mh2JpVnmugbRsREv6yTc+botegRDiu5HK+ZLJiZ
jEoZaf7AmWf4i6rwpxO3+wsLn84k/58RM/QMJ8M3kWoSXgN4jTlh2HfRPM1dpRq7
LoqEJlwVTMy30ISi1f1MnVDNhrxslEuTKus5TuoanxbZ448y0+AkuoA1aUhnHFih
kqai1hLaXg/iXq+x/8/1CEtiGi6WuwBKuPWIV3qyzApmZZieMBAPzSQGcetmFIYK
VwU0+AkMO5xcrOLInvESImVc6+pY2IQOuVbtRMHgESY9cqphT8Bk9KDqZTuP4w9Z
lN2f0YIjyqhUUSESrOAa4zW+bhr0eC2ETBC4ntn4KykzYkGaSakxuiN+k86LSquh
osDjoR34Y1Qat8dLCzgjq+ARpC9hfXVV0i0vannIaCzZbY1eDkLhFpD8WEeZRazA
HUAf3wgx2nSznWFsMGbuZ2zAUDOPiHQHnDzinXn4QCNuXG0bPcRV918KiTtiYsPy
MLsp5ITvpjsk9CUsMhLuL5tEivzuE9wQI62ByR/LN8ewwqTQNXb1lkWryqS/FyON
pncnneQDeqhMpF1GjmIHplN1bWVfRFFn6S3tI/r8hgU2+Fb4h97mpwKgiZKYtn3B
8BDX9hs3tePo4wRtm1mgc2U6LZLNEeiHr1ZSxVTHTRE6/qPWUm6jnFJMPdphw6a5
6rKX2ULD/AZWKk65Wj0E3WGw4UO+utvwjnNH6zsJslh9hwdltLGwMujjW5oKZbB2
JaK/uy8aRVP+Pv/pbX8W3108HjAC6tRHUAwai7rVaQRvqcMLWWjnE0eM2g7PfDlb
ZcGfNzlybec/PEf1jc3+tKK+6uW1ian8FbsAvx/YosDFPJO5eodbnYfAiPE7oPRl
5iyOkQLgDdw+uoEYjvt4+zo+TiwLqk6ToBiOHl5OwF04/pKTF2f8xJ7uZe8KIefs
zf2SzdptUZd0mHRSSeWKiXXKzGuDlAa42OgwYjS5dWIMnxsToHx0HoLyf+eEwNBA
VoZvbLl6b+OrIlRtl7Pj/HHmkoXS1rLPGPne7Jw2YVlv+Hm6E63DEi5f2wX3shlE
9ZjcyZsnAX3nU0aHkLioFrgk+oQZXVc6wiUr2NSQ+cQQdcMaep5H8Tj6owZBQkud
APIA6k6mdiyH3wj2XoDbwtR+7zBqfG9BlPGTScZU4oAT1ChjWJeLVLli7y+IYG5T
NPEpP1s41W5YYT2W23OoK94ymIHI5W3oGftIjV2/9UWGozl3Cojud9fTh7oshMy1
4qGvZieKhjOCd7ohi4FMLW5VEyvhoCkzk6P8LUkfKVOBnlf+Jxr9wCH4KrPa9f7F
fVGBq4oEjAbDARM6zzASyGxt1Ft4NFMK1VdcI9Jv7fFqlcDwWIG3QMJv8amFyeFW
3ydwwZjouH3GlO9m7ZYHe549FbeS+UWePjVQ0eVQKfZaDoj7IUarti+465BodAKe
vjM2d79g3VEIGc3LoIYIRgpbGhdHc89sJQBZpML4dtI+ZvXS8aLv5NGoB3B/Ozq5
XkXw3Vwg0sgK+zz3Nj01N8OM++eXhZlfkVs3lwgd4cXtF1Jl+vkzyBWAKVJ9iR5a
DSV7+AVrr0LVDfk9QB1Q8ym8YLC/VM6iTuKSq7tQt5WhA2Zl0nqK0Lv4n9t/XnU9
RZ5en7OBRc6V2G7VegE0Xow6hVsQERrDYjS2qa+5UxrCtRu8ZV1uBlzIEmX2DRyI
i9BXCRd0/RakaV5g6PH7VkP1pLBCcY7ou/ZTydWamTbrDECmpa8Pcr0M+HVkup4i
c2IjhjlIkfpwBsWpK67AQazH+N2bioCyM0Xf/pMXtyuwbBI5XH2vUcW7UL8SrjCq
IQQqWGXZBkCkztqhxIdhImDq0pvpFLuXEyj87Xy/IfEKH6km9ZdErXwCGvvUo1WJ
3o8Ec1rwuLfztVHg2i8mNHQbOyYXpJERRZqpUsZziHRTbA7S89z1sy2lONarkG+q
1xBU848yP8gbPg+tVjZvzKzS9I44+/uEU0TyjFlAExtjxP5SGw1IeMEP0+kL+Xzg
OCXOO495PDuSonjAPQ8cyIRUBbAz+wyo5uTpAlWqPfdWNSNEFHAcsfQ8bDlqhld8
P8Oy1oscotkxPEt5+TNmaRJKmknZUH3dAaosMbbtnS652g6JYAEQnzGcQBxfrHp9
XseIG7L1BezUImQTu3DAi6acyKMGpXNuuJI6/A3X8HwcDZghzbEG3KYYLb649ZdR
XiHippWHw5y0f/lb3b0wOf2uoQTHpqbl31WR7kr5kwJr3Te+G9RzKc5Je6G119lZ
VCc7+wBX6WCyNF3ibncbbPVZ/1pG2dcXUFDY6ajFn84PcX3odTYI7hJfN1bJbXQp
vvTgdg+kvX5qCSTX7KUHtiX1dZO6vXu/XNgzVswNY45QP3IWejN6ub1hs0HLlxLd
RoBtE7sUDAXy3la96CndMDgtL9wcv8NS3oBhoFQubH+vN9cZJPOlr7GNoV6s2a95
oRq9Sndio7WpXTausGP/5Pc0C8QZsUjU1Rctq8nwSTxzscz1Uk8Q5GsQqTdYymbB
GHo/RMCAToBZkgqP0BgMfrEr0GlldZRlJhLMzcTG+VkLZqn5sjfZStbDeka1rJgT
SDtt1HIBm80SZNaEtEwMXivJzQfGAT7V9A9zrheGZ+nXBWjf9Pjel+AGWvt23MHX
T35ZYwZM4WSkhOYGrLpki3ulK9J28lX0uo50fLnLnFbUeWGo+pDbcyc4NBCTmGR6
+5rFXjVj+ICkC7GZONTiBw3nfHj9ewuRRgwkwpymG4s5VaEprr2vWGf2ZGEr7CH2
BssHlPQOF9urd7SjfKNSI/IKxLHdaN2eUnttRdS8RJp4+NCG/2kp3T5PM36+hf8P
6PPP4JJxEWFOw1cztS+qZWNxqWV9v17oKnbAgHvWGQC1f5gA/QJvj4zajGr4ducL
/jSLKhzJ5oN7lDALhZmZPSTHdkh9I4e3crwfVrtaaostauea0ISo6vt59MFczD+4
5+mxqDyo/yudOQgZwfSZukB6eW/fUvBpsBVWhYB3WqAeY/bwDyRr4vCooMzc61YM
fqYtOA73RE8Xh247fa51b+cZXwWvOwNsr78VBw+3SFWwhreMmDOwvjhlWmao+hww
dCBPiMHXe949t4aNQF0qXAO/Lx17lUVEC3Z01My+iCRlTPl0VBDZ7VjLK4ExXG9+
3m5efDZzo8/CKjRua8tNJ5QejwHUTprwZ4dEWNUcdvfx+g0w9BLZdRhWRJX65c9M
+RwGY68BK7y0Gvputhyv/JzBy9NbHhDsApcKb026VpJohqfDawsJ5C4SIt6W8nkd
8DQUVAP41gf1dwdHEV/4NV1vpvXt4dbaGsKEgBJ0YmVZdI6MQyON71x/DfQJCawm
NpucapJfLVGKg29EZajkdI0qe+mqiGs/sKVpcqFAMRy/hpxIv0SYDCQerVcQsf1b
7bChzl3EVAsWBQzMKxrOQXg/YcGdOeantigqvYex/Lff7pVODNtaSNxZR1LvZPNn
rYdyiGOaYTxJBJ7vGOg1MV/I3ISy6m+YQlHoqNWYVGgfacTCZahEGLkfsawshOC7
PSoFuwWjtDKaAbK8H4u/LVLzInN09e9pch79Dtn8m75Lex3v/ANtr5PmJYLKUKN1
S5pJujxzfv7QVS3lKriDfUnY5/1gFlKY3xApVyrqAa6o0fKeFaLhTT/avEFM532O
hperRVHr6LRTYYVirzIks87OKCWRm3ofVvSad9aWIIK/YanMt5MvwRGFEsxLMxSU
3t11wkny0eiuhm7/fKxm50mO8j+pLG/AK3Y6+etI3GIVE49RMW81vBbKMn7+2qhj
UCp6Hw5SGZb5e+d1wq2kKzY4B+dxhKg9dOrG+7cPrTlrjeouSRZDjYxWFLOhbzIR
0UtD0hRy+4WH1PAExwCNb0Iq10aF5MtVlkSs6rWpEb/CF8UdDws8FdIh3diYvqfQ
yQMLR1q0gUJFUbCzj3tdVIj6jeSXT+PeWAHrnda3QsvJWEwxsiU0YTTMWWLyqJ62
DTBzW57iG9jlz4u+Yw0f+3UG82vctJ+2I5r4S6uFWSCh3t3o/rgfS7IXnoIPapnl
Zn/oxJBvByzWjq2aNMAp6aX71lKAam9gb4khNlYOpgZ8LTY6j7V0Q2KCBODgVOG5
+CGC57KvPZqgvDju10bPIjroN6CqrAzmfALO56fiCWP3nCu4KYR5VlECPOjNrUsR
OV+kyV2gRcoPtyLAOpxlHxuUkt8Gna7cT9s0kElqjxFJ721q/iWSf6l040mciZQ4
3OD5BKu4Z5UfUcwNdZCmhBd6hpum1t0GOW89zYswU1SzxnQZ/XH8TjGE1eUqyurZ
udsS/bF33vpaG+8dy58W4KYS8lSiaqel2yFyOZ1WXuHc4ri2uHooD7FPd3e0bjQY
8GrWgDjelsITUbgu/Xhq9o4LBARZru49RIS9gI7HJRlTNg97a9ocuY4hYxFFLTD+
u0BjGtmoEaAvWNOS44IgMHeWUTImRHE2GCS4gqJm/PGgXgNg3e3IMCl6pEKlRt7z
pEZFu01hI6LYNF468r73OR5MOvkaS21sPkgFNvR+AdazQSqjewlK7XTaV31pWvwW
fHW7nqnOG/lgLyJEyj/6tbNuKzqnjIhtg/stdl9+hdYb3b3+pUzmGfcDYCCPskXT
EUTP5UAvLtUuwHZ/jgNepvHv2WT6XAuHZAHgzQmyURm2WTpJU+DC5mpvksZEuMjm
rjErlkSxhf1pLJRIUT4IM9o3fznyX5gvMJjHfcHlGT9BZUc7k+A2sYWntRtXmwAR
Hw5YbTxu7FlINYx9byBwAcM/W+/2vC4klqM8iO52XHB4QRHakPNurVt3ATvvoX5L
6nVJVre8QvoWjZ+WzhoDuznKl1lN2A4oDole9y0EO+cctADuM69+Q2m/RJwqjd9e
sxcATdrdEZYmnLNayNNeSxpNMfN+4Bpc8hztSeZLkEQCc0bBjWzliJZU7F2AwMgZ
wpjlwMqE9sPsxkg9OdsYp/58lLOYLoT46nOQbMMdQAS0Db1LCTzqTZ8FQtb1r4hK
iTgTf6nPBryZaCiGkmuxKiu5T8aQnV7TYrQLGCVi2U2ditxQ00bdtOev+Jng+taN
flqBjJ3S29R9zqRZ0eDxQlpvgB2PXMSLGu/pAPSUTApSLpVu45GSWhlzVK/dV8sy
ACuGqqs0W6KscJnJzlrgH97+E1ErSnLTfzxigBULNlK3Ri5ltAyN5ZT5m7625W8C
L8gG2DHdWeJGsJL6c73xi1XN7tKpV+AymAOTgW6p4Mrqrd5K0J3AXrxqDSicZaY5
dHRyOzXurfX30WgTkvhK62avE7maqq0fb+U8tOficzNAmyFXar5rIEhNstNY1GTS
NNbKVAIzX88N1dQI/ayQibpCOTEqVy0jPaEHx0Oabx4fTrGIgkOLIQZCwAMJhKqN
XkJ2OgUhkxizSFVqcLHrcLS/EwVAXuZM25jT1H91jhiIGkQWybuhAh8xkQdEQHxf
VXnWguXzOBrSyGjStgB8pTmmCgOKRAYrEKfoj72oqKaK6PxnKy9iwBTTeFnG0AHs
9+woEdgmziQWb7wgJPRmjcXdOqVjlPaIhlfELV7iW0Eu7pV+CemwiQiu4bgQVCMc
8xKDtL+BvHQth0acvIPj+MpGKexdE4ckFSnHh9B1aHxDtDOnlwsr4m70tj/wR/tb
YgXF7RiEluv/8e748utQOSu9jD0hfPBYMmmPKfrU9/TPPBCG93U519XjtKkokEBj
myGOfRq4162AyDeYCGHbh+/Mb/aPh6qAZy3Jp1lpwAFm6Uxr5lTCM4M4MaARxkPx
zTDTSpUklOEs1hzYn/oa4tLm+ElKhiA/09awgT5VSU2sJaIg6Uab0Stt94w/gDbW
UVVqdu20Hu91Zq6uMWmv5xNUfJ3yygbe9hzwIAH9rgoZbPM73aGMil8q6dnJEn99
PL//zPSC4ehBfUZRTXwNQ7RV3lifAzdwNc1ZzQioRxI50P8wjr5BMbknpzAqDp9X
yRK0mHfJwNYJJBRPlHDWMaWIlsCO1gTCwljBUaLpb2qruXoymdc+Wx1d5MjrrtH7
8rrRw81rQp8yuR+T4OdnV+zEKZPKyx3ncGMl9NGne2ko3vBKy6JQTs4Gq3aacdnF
d0udU4Zy+3cLSuHzSGdg5tIrwn2nW6qcsfaTWec8QgCNW23wtB5HQNK6spXOlDCX
x4DLLD6ZcAS9p1lmTxAVts4xgvjkIxkrW0K9JPtkyauvBhX+P+5VvC9RXk6QastG
r7DT0BjDrDgb7NDoViDiFsI2QpsbAAtD2HBF5XgWvVhSckAHoFEqtik8p6C7ywUU
8QbUdGRVo2feWR1C+NSb2blywWqK/jfkAubsLuda98JgE9zQrfXH8WXI1Yj7nnH6
Sjbg4YA2rPKN7+XGNo9Yl91sGL41paCh6412mMF/9YxRN7qJIUdXKIZDV9BsrnQw
M/hHPU+HYNFJlAI1GNyEPetbBvM3q2zyYBT/07KAhatrpKV8neRz491nRyQcWoW5
JnM/JMwJf+n2vpU8QrMz6lAy71lV7Rt/ylLb/M4/oJzx2zJTzRULLhyhlmkvu6zh
cFyyK85vedY3lVeUhjpFmIVaxeEv2lZO1nQzUuZsUaMxxgwY6CEPXHZzuumDZEeH
AU1/E+xCdl7q42alL8rRYYymunN/uz+L8B9SGxxRdc1YdLFWe1u3Cyg1Quu/ALSM
ttJFX8ITeGoQXi7F3GNgY8ChPYY6T7VAvuktAgan79IpCgFSFRP9ICtyp3axXiqi
6XiR1SPKKZOd0czXcoGClIVjLWY0lde7eDW0+YT1ZZrx16bZQNtSSdkKK3J1Cw2R
2ND0DcfVpzO24ZCPq70DqjwgW5eCuDbmtIcQ8OoumHblT5vTWa8Nf1r8NO6hVBhi
xzzEUWWOyzg1riS/yMWyoWc12YDbanCRlo62mVk79f60Q2/+d/0BRS+w42+MocwU
1HqT00+1FWMPghYsV0cQSeX88Dpt22f74ZAcbW8bYxR0TxHEAuQFR1Han06yotGN
r+Xb94BpBK8w0AOuwu3XV2UqSBJ5mORBAjt+RnN2fi2YNxOyn/yw2JmXC4+w+UNx
kf9R1G5Ud77pifV9UYO92MowMY75tqUBC93WOid2hvoJM5BHFx/MmZLUFI1TVQH9
3/GEmqwfqQb6jjIDvNs7u7k/OPhMfDehNwmZY74cOL0NJsVC7fgtFoc2zjg3tLHB
G6X9kddVY+hWzHAyvgz2KCkP40Q34aWNYGitLq0nydq9xN7iUbw0It5DF1ONJQYc
69zbXej5aCcMinoIn5ffjZawEHmwF11qfrMnbHlBWaQt/eDALSULWrqLfr2BqQeL
xJJv9WDTaVjtlHkxbkehMQoLa5m618Tjb7Wi48OSVR0nBfyAZ5cdnRiyaHqAJWe/
8zYDVRlF7gTutA35/L/hw+iYYFZg5W1AaK9W7/84X4H44cj67z8CHe7FL8Eaqy4i
ixhxSobL8XklVpBakXeSFk4Vph0JcbEbRQ5iAp7anR8rG2GOSMDXjkM+Y4AZtACh
32fX24vuQhqLM5DuLCsLat2NCe4zy9qTBW6Zac+Mt02OyKzyCst8P4AwlS9aURmb
3wnT72HVF0aes+t+FZhpekair5AoFtdFXQwRugwhGtiJ3SWhFY2rm1+3QZf/Kmyy
NXcbVNGw2SyYKWvmppnwMlvy88Pl/GrukTP7mj3BaD3nNHUYnQfUd3Lp5uuY4bHF
vOrRzH/JulzHbBS34JRWZU1SNqvc5WZ93eNpagwS2N8c18lxp/wiJNDtIAeEpOpq
JV74IiVdP2VrK3Uh4aouNea7enlIBeNBxSZV0hrZ/og4/ZD9SnNy/IHRmWsYvr5L
JXyX9B+sytbWi1KKeXTjY1RBRc5vclf+zLZsj0Vbi6tb/byazHaooJ/Gi5qCk1nl
W3btL4zp73z8GS8RC6RpATp0D0v4F2YbwWrJDIPY6ZJ+LRNSCbPkDpPQ2b6x8hl5
GZwgrp9H9CUNobDc8vjy1kyfu9oa0VVuwiTcO+J8YKHpBg0gIwbOvc1Y5KesK0AZ
HF7s41FQ3HDAlDwHFihktg/4U3flKVT0KI48WIwABTHHW6Zad7Tq58UNbVFxiMlq
/RGUD+edeMN0xsWuzuR4IUypds2vhXAwlL07TMwpGu7XJrhua0LYhef19VtIZC3v
ac+oKzdJ9YKACSX3FuAj2VC6NNIKBLS5IKO/jPYcjn16SkS596n89lBLwAg9fUUc
Uel2aqkfd9tv5Tdaz3l22gfpIc5tI1O7CTieiqtnQJoIc4gTM2BnEMG8Y4xCtnp2
KoLdtz3rXjfrUJcAok/d8KjQ3pITZTbJBkcBeF/elyWh7j9KDZk0Ik3unZu7LDQS
JkwoeEj/deHoo6IL+Ic2g3THzKAMYqc626sEpdN3pMp2xAly/+QxDnCb9HFh+1ci
PQJ1lR5OJ1E6KAGwVwR9tdjMEvFam1m0AlytsYXCZmiSGqlSBnRlM+dkjITyUwVZ
VQWmrqI8zPK5ZoxNrqyj/1Q6fu9mIviYusbAU2pFIefUkrVbTBRGQTumujSIfvIe
s5O3p8M83lqNww6AUuCjVxycDjqM29DhWMriwhOarRiM4zF5EfTav+xSyw5LzaWC
8nc6OMDceaImsC+d7S4I8KbDIh9Z2SITIa1t1Ud2KCPruuQ2qpPOHIqGR8EGdxCW
r39PiGkhBEGGXhYz3WGTrUeCHj+zMakpfSixl3HLivh8JBKMGUextoa7QvCfJjsk
is8W72SIwApKEa+E4s8Cdgfg0/XBlhe2nHPk/JyP1UbakmSiRt1+oVS5N0fcvUuZ
jJd/GKj/iEm78h55CxhxkSbDtf8LtP6gh5WMx6itYbvVp+FkZlH+uJvR4qIGAYXx
4PKkoaOqfkt5KUhkUJ5lcvo2BZcloOseg8O46M7/k1QV3kOlwTWz/rCi6rSEeD1L
WOWOdNVuy0pxgjcMpJRQs1EhwUVjkTvmk+U9Jd8vaU7RyK+mvyakPmZPCxBjQW1o
WQRSRnQgpR6Q5c2sTarnuMCFfQJ332frOYcRrxFtb34uNDHs3KVQzoWD3APnxKwk
4CEE18HWKKmvajvMz4jBhcVsmND4EOdbP2hhgnofHXTVlPf+tBWhLizDu2rgxLHy
fnSEXvdJ3Fn6KLsNmF1TziQUIPWcTIwAzUwUmO4wclSzzgkhhFpVqZfrhLzYT/iE
uoEG8Cv7FIIz+h/4ZHBMjhX1+PrePqh3HHKDDjsHAgGuTa4dHqobVrm0JWPF+mvr
smSaxiTLIcDBhwfq+so5jGBXQACjI9EtUeP4dXf4zoCUdfp+tcXKgxb3ssbwiWE6
MBb9bx8YWNT59befndvLqWRIe5ZaqG0xYiVrQp2sQZ1Ch5Rvflb3Wn/flfCWDVLq
kH5hms1OrzWYemn7DP9wOABLw0Qy/JXJmhthaVtJDJ7ejLerSWVFufEoo9e92vXr
vo6P1DpvqIO0xjXtk1ZcRaeNvK1jvuwmHCZbozha1LNlG7PIorZ6OF+3vfPKzBRv
anOmXr2krDe7J1tgcNB22nNsV+4EHdUu9saHZ5fnMzZdeyezEzmgyTIlEQchnfzK
pMWQpc27LHf9JlbRNR575VoEHG9bFTTIhOgO7womkbqBDxU+1T8tsaP8wWq2zWe8
vomxd7//bYxMVjaHlqhcsvr1mfMTqQA18jXDlvjLiKd2Lp71MRlyoLy4QgExSqlL
OQ6JC5QCwL3hNpE9NIXwqpl4nKHvN0LpFawfzxSoyiWJ5VYyyNqcddXkL+FJC9IK
Ak6BhoUhzrXln2TTZ6TE4Ux9KVChYlttrX9RKrSBuqt63mUOxIsllhuVboRAZaN8
FKc8ZiiWBYIzxnDuD8yCEQ29oYe3YanLe+d2CbrEjMVpDXMmrQy9MEdIcY6/55+l
6VEHvp0zpqHtBPfWNngqpOQa1MlB8qsR7+oQ+E0Xp5IMWAOjq8lvLdoUycLrKLXH
F/hqDyhsg/M+B0OmoFJDRyRbccS+wX6XyM6yXLe//x+gTsbnvrd3mk7vhlG71qX2
4eK/ZamWLM+XjHkHs4a/5BQQ57juzfHLmCMzGgOY5969U7a2pNo79693kqBo1Rz+
+ti4MkKitJVFbUG7ur4VwHPT2oKEqaKAJx0WhouatQNpCASw8JSDAPS6bDUduKRM
00kpsBBIFG97VQsVdtqqzBPCYXuZhXBVa+EAHHVgVUkWfZxRtuCmsqS3RayrV14h
ZkXlIcKzGye6rJfaAv5o6s/jkj/bJeu9f8UfyIkFVJySHSGnxmXeNnCytZZkG1yl
nHY98t13vPBIZuHpF1kU19UVA978q5hZ/uVoCwYLUBI9xOkfG7ELKUXZLlpNCUVI
9bQv3wJfcMEEjGqFx11dhQuT+oa0Pi7Gu2JWHR7hbBFfmL1HCXXNIcG6lA2hPX3k
WN2tZ9+YaFyhnT/yjS+NVF6x5HmvdosZQ3AiwX/vY7GBVvpjl2/cslkPYw5HH7s6
j/QyPoEIM8UpS7WCSS3KrLCgSJe8pKPvfpxwMPKtakXFGMbapDWL5wxVUPRC57xk
2ygCze4mBdhIJga1NBULuusffE4ZtZaw3Uj9yy0yEHUBE2Wp0qyNElJfQIsAB/3k
qPFtLkXBAUVxcRJCBaI6JAh8qql4VZi9xePTuRE/ixtIRbDH5698nRxpbzhBBCDK
/6lbsbKM+EF8/t8t4xbJ2J0C60K5V7EmAgSDP7TPAKH4CFSdc11AmzQEvaErkWoP
xuotlUs3APQBn37vu2+vHT8li/Tw6L/4DHiHoH2R/XH3nRgLQbTQEoFWCUrGRK06
BVVPotZ9O3BZbuGvusvlHsIFCnoav3KmQYJMyqrGxyWwCljBMX7hjbCdzfxSFpHp
usfQsLjCkafx5nipip1ZNqbgZty7A73VJq+GtwYjZ4MDf0SuRhmHpTLXe2AlAHyS
CeZ7so28xxLK9LqdIZXCGXgg04K4o12M+4ff5DNfOITzxDfCekAKIzpJXtUey4JB
/U7jVQO3WRLeVLPQN105FGas8x98ufxcigpEW2Y5KBSvYSTAFJ3KZzGRYreO2i+o
rXBUSWvcZXsgnNJLzH+p1KOJn2ynmUdTs4CQKMCO8zhv3YJF6gE9En0c3GTay8f1
NBhFKaSIocllUuZaV0YHjHwGRJaKB865J/mO4PreUogXpk/EKnCsbXApWur7rVRR
yk2qjUjFK1LJPjhZtVVurhtpt70wYWN5UOVDARoyKJCIWtIp/P2dX6hATtgNDFtP
+zbYQV+u02DJKdnNFRT9wNBO2iW8BgZtvA8mk9MpTreTZy+bmjMC13qMqh5BjOzJ
FE9OdCQIsBcjl0G4QeDj/Vv43OO0t+jjHBisYhtoXfxG7LBsQ0qZ5CJEyU6tHZwQ
TVaJ6OAQUlfJ1HuqqzBvSqrpBjPKMo8cM6366fgXTKsIbcdBHP8vvsTkrST03CPi
pCp/hl+dqwUkS2xcmRD5oXWZ5DmJJiuLhJ0bSQ+sX1KV6cAsTUsd3LBHJhFB9KJm
QeR4XoMNtsl5DGVZTkt14XSnuwLIjeX3BKSTaYXpb40oCsTuMbGFeRL8JnbaIe28
hmUqEeqAWSqlTGZcUOwe0zl7mKNQcDL/e5EO6yJoUUXYmkqO274qMGcesQkA7Z/d
X1sjgd+93RxxA5O8fAwuUsbBliocNBRbWmDCmhvY8PYmORyVw+Ci8uMXQp4wO5vA
6c6wSiwLyCK7sM+l+smKFMlyniCTWtlz4QMBXX+WCgWzpbGXvCNuk90iCr+K0pRO
CKBZ8TR91d9xO/qns0ja89mOT92cKdKHA0iOqaYCf33lMMb0YvWogksCU/1kMnXN
Ss0kcwJ+WXZzXuIsdhtdRRtQmgUMVw/vpv8PqALupuSXpI+6U2MNWLCheNBJd/BE
lm6cI/6AjW3SXOwbFbihkoRNfsVHN+ZID2r2vv1wizbVRdbrYnS/KLQgj0vzlfcS
dFuayDLzorkVTDKFW1kDXTDZVX+nD3GGo9T2isr40Asrl7CucjVScc9MwyRBdfqC
z6joi7TPOOkRL7h32RWg1583Iv2zHwNAAnXYyJBMFjQspBgsxzs5yc+3JfkVlUur
xzl9VuVc1jRPes5OCHCA2IWPVeo2yx50nQ99b105qEvgmeN1K/GNY7xzQhsBF9BJ
UsQ25pVbpcS6xizoqaxwxLSwqwz1LBsXeZwUDxwxACHsRSmLFyxCAWuuik+QIAqd
qu91+NKROLsdvwNQfN0sjfIMIe3QWfDusJJH3LGDmAUM2DCjLitpcgsPDs5145c2
Fz6KmMmbdaiqDQpV0btAlWBYB88E+ct/AYx81xpr5S66PmaXJocr53ZzKUHePJh6
IYYZgF1bR+CcBvYuU1rc93NlnT7Gig1kbpOafo9y04Sm47PRoc88VoUOcFm7CkRj
Q6ldOuhhBZ6b4wv3T5YCMBpxzBhjfE6XdHMh04DX+kaK/QdN10jcaSqo0sRcFs0F
37R+RNGdXOoJsTtVW0Ts6CLTLdavfXhP+KzjXyMG2QEFj6+eKKmMYgapYWdAeEME
kpSK7PNM2d6RC/vg5qnAL0w++WAl0D0eziGVgMagyqSHu+6RKOKx2kkq9GPiOwRk
Th61QA73+ByH9gOCdUkG6DPPTasp2vG9KVXJvSbJHJPIUjyFF8KiS4nFxWwBXv3b
PrfkHFf/E/Anj76mj6Hwv7eU2AT4LnrryUvKO9dlGA18oySxdJvI85NjUtSUrwMM
mtWJrZoCfZ2MkRWUYMYro0MgG4Sh1qt4//oxIz3lo5Z65EsWuUdBs4mapvvK+qgp
C5StIkBcAi/tRR334/Ny1v1F5jE938USruPEXUu/aOkw9FfdbQX/bBSxunNsOp9v
tVnqc7BY0oLZe+wPJO4pnu/FfQAYIfoLdK1HxKpMj8ZCX7hyHWF72CAh+OT2hrth
zwJmEC8lkCz6kDs2QotRKGSDs/XekfgfThQiiAG3HSPb7ySMFGd5mX+9X8fZftNK
amejcAJvjSQ/FakkVYUw4G6PUiEnNSS1Ni0mWsGzyXVaoSl+B8jxmSDZz3xPW/a0
lSorzguJL/3KcD2JGhyORW8Hbh04N6zSjd5rxPZGPQti9h8A+8ZSjt2Ii66HTEIh
QPV+wfYmszRh9gLKgw8I6BfSbJVHEHlbSjtd9qKEepg/QoCcCbdbwfb7jyQROvos
TMOED4BZW0eilnwMiPvZXAf8NN10qSKB+M0fzDH6HsoiDI3c6JYH/RZ1+5b5mqKi
46hkK+MOP8y5N0trVPR4berGk79VQAXQK7ivo/KTKFPN6R4aUL/SRar0idhN4CUB
Qj/+APu6beyVp54JqK9AkmMp72pWHU0ODcIoaToVKhaZrZyG92J8/CJFMJ7ek0ph
x4iVqjTlaaPl2RzsRnhFrzx9rdThU7iLniJ7koG9V8UnVyzxMbU5IfmJHyAR7QnV
Oj6h98Znpg4bc95sG9lMtKH8+TJhw5guC+UKd/QV//U8gDOfORIosOYAkzUQuP+v
Q/u4NQn8xCF3CKRs1BaoPaFRBqRZMXdahkJejVBLBlrnLBcrJP+GJehCRjDhrPj6
MoicTII2GupoIfSP7v/m4i+fDcDfQR57i0j6PQc8HyqWMBhvyDUkc9bvYokXkZro
VJFzd2ZsYu6MmYGh4iuBK6NRTDIFDGwhpVWHEUjX0lAqj4JGDYIPMO2rbzdbeB5u
SNsjmoXtxdiPKd09QBJs63tsaTHf/ZKC1upX5jUEZgSdp5I17MYUHKVD2nQpXw5h
MGqNln4DdXjYMR+P5FUmbG5VxT5AA6dUHBcwEDlY++kwMEOCaFlBq8iUsG44fJ9y
ned5nZyOF7l/V5cJTMl1XTiL0eN9JZRHnsNfYNCevt0A/u3j31JQTBELDEWumE9W
ngSH1MJYRAoAAYUSp9pRwKugpoumfWvGd/MfO7o7FWRxNRoOgf/ZaauSYJMm7a2G
QykwD2WaWxSYsc9hwickWqfKtnbFkRzNC/08+9wCwktXw5gDtDGVU6K+DuNytaXX
VLVONN2WgOE1hWIybONAUAroiUSCdxqYslFvJUboK+72kRttVi72I8ZOFoccSj+u
4UJ+MHRvwdMHaJaNHqJxI3hMG59b5qfWGP1yN9WanbtqF6LwlWzfIkwUXwMCXGcg
SsVMHw+kx7jJ5XzvzKuvFHo5iR7E7IG0Rj5MMyRAZrjJ/h6rQK8XYL87mX3JT/Fm
ReGycAEiYTzOt0+OBA176U4ewNj9hIVKzDubquypzEh44PSlHt68NwGFJ2Z6u75c
3LELwiYypkDwwkg7upyF0YxO06dgzc9Az/Z0XV7VNGyl2vCuLzx8VF9GS7o1eHau
0EnY835PEFSt3UFdfPdoyMY7zNjewmgjGAO0KjQSZ8NygFskOzmXxWNkomgQSsNf
UHWCbM9QOiChLwpRK93ae133oQhCHyELgQaXfcgvU3TZVluOx6IBFXsQpxDmNFy8
FrNyDzLBbLGGPEIstvSnD45I9ND3Xso5P+KselP8hNzJz13k7F6R5ytHDlB1BBDI
De/dbIOVHk1DOdhyUFzWAVF3CETOOHIRWRzAqmtutqqxae9U+gxCodExFZoUs/fA
mLVyt2so90e4CzO3Sb2uMUdIrkotV3TOuvcyrb+3/s/idEGtokbEzUIKEZ75j5Ot
XXfcMkeqk6EgcExRSQYZzgXDWUJkxD7Efwfx212+fYf3IeoGDQgDYgJL1bZKjSyE
QMj5HSkCCC9bm85+ukZrlbkNzDiuMOQxMs+nCMoq0nfhWdG4HaIebYphi0mYygb7
KtzHZjONifoBnWEEGDrBXF7CQA0n0hcjvJqlW+taTaufbnS+llaco9k0GDhUBUUo
EdWdbjLgp4raQtySdLMZ9EgIM1tTQQscEWwEHvMCuxJpvgmaR2BDzOGU9ZaGV2fO
FTJcjKLaJgbKbheuwIsMm/vVWKxOtdMeU+NLBoVfw/mh2rCEA3+eVhtIIzyz8udM
JUYRyDlE3hLgWr2axqFgZUQDF5qpuP9JwF0zN1uAJhINpGAoB2saJVMZCrb7fSmd
bnhv/2FTMI61y+ruSXGeaP+LITatSvY8ougSexf7YC3z+g5bNl0JKZUlPUZ5w8W5
Va5rNIguCzwKR78Qju7QdYtsyEEErOXEXhu11j7agHpFpwITo32tZdt0+rvqj2pw
+lXeacotk+XJmW2uIwXw24wjat+CKQNZbN8pClgiJNntYy9iNozmPXFw85UunN+Z
F+XKrRQNbBXRzI3L6dvuwxbMEg/PLfAqQ49YsmPnGHhxpI2PNMzHg575pnuhOVJX
uik7Zq+60EFQMbNhAkb9a3G2Vn4xXBdWSSKqT12jrRZHtZxVTi8qTgPOHaEIlJaZ
sp+qX77ekzfUFx0+f3svBdYEyHOjLhLu+yUuEvlNpvcxrt6YLl/gtgwKAqjayupi
Q2oCPV+oR9rogarcZpEXm8qoa0DfWtA/QJs2SWCmYdjE8AlW9n81J6Rvlc63Noyz
Wsq+hNXmxsq3JESqEayVEGY8tUur4ytvrzA+YRV71m6RUOqB9HA/KzYn9Im/t3d5
rFivDH+8/zJSlhXFGo60Xr+X/JSGPWUZN8S02zMyIh26NNOVros0GP2u9Bs/3q4c
uSz8Egwi0qwPPAsXOR4bMotoaTiTs4RGliTReyz8B2FUry0AhRbu8DOw6qihGuHC
3HM9wdazdz/MU7S16mt/c+HcX+QTg9tZ89NjxXw4LMiCgWV+Q/2+YyRMPuiY0hpy
fyeWfD4OhLqBrQh1piDqKhfWpmpgry3XQMJ1pNY5E1u7XWq6MA6ysL9foOwrun+1
PDYbrrabyBqYox7K16rvjVyZBu7+24o61YCVXz2lG3rgdVmXB+oDYMJphabC9Mi4
F8eVzu7xzAd7d27eJ5ni+XtQ5k0Vejq5lwV8VRMo5D0ye5X7IeYMnynRbb/5E69+
u8zGYcQdnhOQRWZX+fsMENjzw9i2nqdwUcmhshwDZTpxNfE2B3r/ew/c4bCiytYF
jCwJ2QRtCTd2rFIcB6tyAfa8z7BD3GmDZTL0r+IyV6y1XkoxvOSkl+OCbGgRT2Fv
tAUaumyePOt6g2Vjj6iKhX/b4agcq8ioHmm2FUwM7SbgGdQswW4yoayWqVRvtO5F
g4r2W6pLoAGDp0nI260sF6r2M3zxvgd5sOKffhshX2N3ABRnVa9deErEMxX6nb+o
aHDuJSct5XYR88tFNejt5KWDFioMBOQfu2Rs3IpNiI0/1ktpixGM45j6/BfHU6pE
t9JbRwyX9va/d/hspWqhQe4swcU4uX2j81tDBTPQOZhjDEmTG9IF3//B0Fjg+2Zr
RG2eSm6AL/P0SC0+jWxZ0SydS0AAH7dqwUzsZ2BRlSYoC2ctyrd8/QKLwDeDXHw4
la7eRQK9bMw41g6AUdLDDRoHxvS0aVjPF9LUAWCTDLDwec3EmsoUIrjYiyvxBZ0L
2T3J5JDhhe7p8PUdo4B2fTK67iGvVVWKqy50Fjd6ofBYdXh2nt3lYWiVxjIFt7Jf
ds0uajM/HOinftZV7rNEX0f8Y5RiQV6pt/aVkOYvGK27yMDboCisJ/HsrQRjq9LV
VLo7cqZy41TekGyO6Da7ntdfFt3T8CEXR+O+rMwlHbo03QrnWuqP8JP/qMeo2ny2
M8fbp0oiDU3rpSBnj9vq+RLoTYZXv/fVSV0UpPKp4Qi+X0yo6jUwXxBXfok6/Nxs
iRRgKR4cUUoavO5yKzOviHj36qCxaICNX6LtKmKB2QTyvpoYlS2nSWV31FmwZJgE
nE0J2I826D9PMre810dvnbcmNl2X9CnaQdlLE+6q2luMai5hTzIRWCoWOXj5KCzd
0qA44kwSX+5M/ynlcIop+CNcBZiOE+YlqgaWPVxA93r5zQ/KOuP6IcQSTTRXzQju
rf/qw/6+5LntUC1sSQHPaY7/ZRoAGxbD1wZjpByMr87z4gdTIeEhpN7nEXXso6Iv
EoBfhkH2ZyWR8DiAat4lJSh3rtTPGVDPx30fjqCRPDxiTgHlFAHS3WNSkwfk9/BK
cmhizarZrdG/btpTjPTDBNc8cjWMSM0wTWGLhKr1MNSbVFe8fpo74/wdmQBQRQpm
9LjvM8CXtz60nLbeinEiihYY6r2Fv0jZOJPXk7Vcj9yPce9pssaBSCP6CmDzRcU/
dJLam86oxOW7ncOrDVHyeZYjgxjtJM6dyq1VJkHyYmCEItuTmwbw4x76AcDUlh5x
QekbyJ5V+Rhoq/2/OlKe/nytOs2VpjhJkleTRRj2vr5Wqb9e9z6xCDhbFBclb/nB
QNjvJnxE5kq2/3KMiZqjyXJFDTKxAga0PmzTMMtHa/+Fbu5vg7NtprV0oS1tdgUS
ljQRdHhaPayKtezIS66GBYKERP4FMnrY5FhORekCv0ws51rfdxG96oZHFaeZ2B3r
l9vG/SJWRPhhJmB9ksTkhkeA3BHvSSCYqkCPrEyFf645GCHrdvjMD+uQJYTFCIOQ
Uw0soD4FzXVLbhY8iFp5ezeKxAuAB8HePZmwX3rXj68tLe4pwnbpOu3bPky3gi1r
2sOnvaOBcljIWIspqZk7Nzuz8nB1wG+kA7RjdGC6Aqtq8W5GG3rcObQyi2L0DjQE
HsuQsZpNFCkRT1XscIqcp/rWXqyDqBsQvfo7CPiQQ+mSCfbzV/9/CxErVYmN31V0
5ph68GIfyprVo+lY2D4xYUDi4sM17M4btOBJjndUbjvG6mWZLj+JDeR6VvihFd4B
qCkOTWtjDHFyhWAHQZ+7pwNyTcnqCcdn7WB7QxCmL0cB8UCmwo9f3r3PPPvPJ2G6
vlv+wkdi/g124UaIwnBMD+9u+G1jZVXedxUwzVKJLKs3eUMVw2+A9NNq7qJnkNyV
QfL/ALR4tKdiPuz5OhmNX4FQTHg4tIjHw/pPhVDYUCH6RsOA5GOz3ZyC+v7hJafW
1zJkV3y2QE95fRqVaDxsYbkKYG1w5qjz+nLmMW9lkJ1prBqwErV33N9zEHS3x9R5
TqyXhlK7QYwHxyxtTIAjJn6PEXEJAHUWi4PyQKKKnhekfBBfxjEQhCwJNrZNKjJ/
N/5K1G0SeO52yGsLFe5egDgGoRT9nzzWAW2Y+LmkXDakdZanAYeWx8CgK39Lh5YW
V6YvbWZ8mo/CeeTioDmyO1XJHZXwdbF12v7lDv8185NJIxWvpppm22+ZwRpDLCM5
RklvY06IXOF11d5q/1iqNPMPpUzBq10O4/O2TRndo5Ly/4gPR1Ggrayy/J/B51Hp
WkcgD9DjottD2L5Wtp8W70Perb4EFzz+60gt6yft8h9d9B/0xiWb7qdAIiY7mZ4Q
MyEUsbPte37AnvNFC1o+xlr1jLpAYfvgKOg2Bk1SCGx9s9uhf79xGH448LAjSXdx
dlvlEspbMB4hsESfLgJ590vjpBv/KKEUQqGk9w2ZXvXpdykK+Kqv9xvh+QZi47jV
2oF0HUTc6JuQhD5IpZRMuLnx787ia7Hda5911M1T+nIrfGcEBuSgQ2ybyCxgOALn
Q5q4LXKzXcgtF5njb90pOnj+QfcBEpGRZ3OGHL2crguC7vcdD7X8zcvDEEM/UdAl
iaXHJIOsy0Wnm/2+YNZfXZF2DQXjUDcSHnFvSq9QzYGT0bGXLEODipnNiZEqE+0N
014eqqkplX65W8T/Z9gVJyx8cIlfw88X0uEaLP4LjulBFZpLU/PfbLjTBbox2/eG
M9APuThPNwlTQXbHmdpZTyLqPc8C2imOf5jAAOFY4uSEkf1UF0p5IZc0pgr3g4Uv
9DyshtvAa9Xeu/80C3x3pkbsRjxe2PVJZSZifNWYD4Dbo5ZE58AFI1wMNJ5W/WDx
vXbic+ERDWS9/U6pcm6oGHlEpdYTe4CHhIL2dLYqQwKWPE3MeEZwmmZFSMrNrbHq
XMzolzEDlKT5Moml9XwvARmLgF3U0+YAzwlU68xeg+nM4xBw0k8GNRNjQ2VYYgpP
LTeIHplZTTTnM3fj87HkCYcbTvXvbnF2VlguPeevyV0lfONXXmiPnqJfBimy9b3J
el5DRI+VgCDAQkVVxVsRvWqHE7iJ+qNDmZXb3lzzmN9PTsCbTiJKPNE+OtMdanVk
XhfdrrFm+9/X5yxqMa/Qe5jkttAMTb+/0gJ9hKZp4BypQA1rGTQ/zsqJqJdjWlk8
CuKfMXloZPKlnYJfURU+VONBcRaccqUKDhQdHFX679uSMO5sFgTfcg664CIEGvs6
984GaoW0v4RcuVRxxHaLX9Hz8ZqzKf0fdGf8WieiGxOhcv3HganvaJdaRE5Xmtji
WBMNc8JNQNgWgqLD8tWGwrcgfmAbf/JTSLYE//KfVCKWHGc47U8axHQpqFA4Vbhi
BnSE1eZ868pbthjAuw6fXUYfaRGUywGq+wxaKCvafX903FB/BJ9GFR1BqG2IK5av
5xCNFfstZbzYnwJFegPrLAu7ZbdpCbMslwViVNDfKJOFUKIei1EN3i7SRNUk6pjE
TW96JBB8yy15l3UUvnkWG5blyUtEvdUzpNYOaqCc0kozncBv7AIKExQDCa6FCVec
X8Wf198pQk/SCtNi3MONmj8zjuvctEUnfkn4pc3tTT3z3tdJeOMe8L4d87l1WL1q
yaXFxI+g9TyuOflRlADrAEs8cHPRYHH92z7bS7cswdsIkWfUMYkV/x4lH4rz8R3x
MSkQqj4JccyWOPy/dsog2+KuxEAfx6hcm27NxenmklXQi3rxBL46VLsyYMIPdCtn
c6i7HKyKl3JJUTzp3YFtANlZHAMfH3sAVoclUIgJu7O6AC/vPX80ezMxVQMUsEq4
6M5IfHJ4zbqeIJLroVljcqcFaeD5cJeDVXmMc6iFolCtiXHxbb8JFsdcoM2awx9T
OT0hBVwdYWh3yZQuLfspbqS5ZAISBflQ5Q8aG9xwOON4z5TrNgw3mVGbhiI3UFjZ
DZXjG9s50Sj/IzqgOihnw8Quzii9u5SWOvPYuf3HFa7mxHT214VraESva6S+Zo2+
71t3c/RPUzHVVSI0RhVX7zAgkdUPnsaOAthqBmBT1liV6EZy/f5984VJPrtL7GpU
luzSvXJGAc01z9wKq4dHG2MOPtSFf47P6Zn/FFgoUAXBgMM99rLuk5dFY37irjRz
aJ09GyOiYjdniHl0eLT03OgR6oApMlQBYlFEM/0tTbDk28aOAOKQ50xrXAfT8QsD
TrQk+DCKe2ivaIJ5HMfhyXxMCEqE0MOQ2EZMhRJaChHG9IPjx1TPtpz6XBgtOO/7
lUq9l48gOVQtfqkf8qDTBFy+jzkWotrQsSECI1FkYOWU4m6e+BUDYKXUMl1FKJLB
wqQEoEExNKR+CTPHLBzIzhLYDtgyH+AFP5dQpnIXpJJWk05zJjk4W0vCFmzPKmzA
/xh5fDfaVN0AQoQ90fvi77OmNHGenUdw+e5tVUG+8ecfYpncO/z1rY8/2vzjTTDB
WuGkg248VbEyp0uPvfNN2oRv+5QdiGLgpS90CGP/daEFffs3Zd6enkLz7hS3A4Xg
9I9vysTCTVWEbT5Ql0SQ4+TgZKofByNyBByOP/KHs3ZkZSLbnoT0XFMDlS/BRnRP
FzVvbcGeuyideEzRx82GabOymwW24aPx3nh4LBFmbhurZkpXwTJ3UoXIcpJ3J1fE
GMr2696ABdxshwuUCWm/8kHCCmfwNGFBTU9gIwbEGzKKL4ZpAl5DrjBLGBCfdH7R
oodT6NCGJLCgUw+xv2WFlUBo1UL15FDP4U0nwknYnBxNQ9Bi8Lg1lVqh4BRi27Kf
xDgEd2Ev5yLDQw8WMMj+AmNu5I96PCWDfaVZa5mCFoF+Ef7z5UeU47OZ2T96sYzW
FO9UikkXJMndAkWoul0/BoReLt6wR+mxJXuZAmSb6OmY6iKlwU+6gqggA3zT8XYP
w+kWwDH3I/e42Hc37JmBzLxwsN92HWzeQVsSUJpikrIXoRTkRnMYsI+qXrl+ARtT
AxgRP/mIc9q7tzKXeSIVwoUc/3PGX+jlwEa1v5xffPvtNt0jt7tlHFu26zWSEF7j
1LIVql9RF9LTgY1XJK0qXLNuaKC9atbp7/bTSrQXX5s5fQtmd/0QzKP+1Xp3czmt
GVVWWXjrnj+G+VE9N32DFbeo3rN8L3xjU1GGb8hMbSYhRmzsMmBCEehtNj0338Et
j+U59j+nY2H1QeOBUyziSnxlHXH3kujgr4mAXvo259jLtMMW1zEM4cV9ASanlsCG
Af+RoPobyO2t8m4lzleO5nh6Kms8Modzeui4NRTiEIC0eD2mbGnC1tF+vPF/XyzA
7FEjT6/HaE4ynrHuSSoo/tvZpHGvkgL7y/7v38vtGucgH+1SmBwLIuRNmazJD3kA
xjH6j8KNVAzipKAzDgufODpcPVbo+baf/y8KyBWWgbs83Q8rhNz6Pwonys3qs5i1
Z4R2BB9u1PYw6Ck6f1q0B+IMKb+GeW3UoCr+J9geUwfIw5pgKZgeVNOuwOhfA2uX
lFOl87ARRdxOLKLrCnuvjpSBJBZG1NFZpsIpnbZys8NSBlc3Jbwxz6x6Vp9uw85+
lT0+0MKtOH3WOcYjOp3BHa9Ww/szy0rnNbouV0qEraTwW5DDNQ0WLqhWqnO3htlC
+0xHnZvu1lsPge7MBwBcXx7vMrMUR6IpcboXUpxFW8QsJMEbCy/8C5ZF3Aeen1gS
pCHvmOaCBmaWp2dbvHJUstH9M7qWi/vCbFQo0l0yM/iWVHLeOh59ISKAqygWAL01
fcLjCx2k7YaqqrmzFivKiDtVv+Kc9YtmNZQ768P7fVBmlo8x6Wv+CX7yaUV1Kih3
A8lbA5gAFNcruMqeQreswB+ykxTED5E//7TbasRt9LGp8dG7L1RmtP4C5DnHDYzQ
r5W2RFabw/yKwPiuygaXq9F197Ky1Dq27CvS/hILn490BJHcOlQDGLzdNsZjL8O4
OnNTnzrvFzhSIBJHEhOV7Zn8F35PuudVlP7lhOKnvsW50TfZrwtrp7a+NgwL3B+Z
9Qjvjik3MvM/2mL+lY+wJB51eKBYDrfL+nFhhT6wKaXbYo5/fNqOdth59vt4WGZw
fU1Tv8xXgqZhWrM9JBx4odXeN1+9s/5Z+b8wGyPGIHXsA7LOtC2hMMH5b3S4Zr5y
EJcx4HNeqVi0Ug1abQl4fAVfHgUBHqbWKvGxA2so1QDUfJH/NMgblaNGs1lFCfAk
m106k++DnsqxK7s7czXytH1ND1aW6SSzT0BaNQjkU9lZvr+9SHZDcuQRqOGKgIFw
EVyBJ652wA4aQ+95R/HXeYtkkzejJvKqt3gTX1H3LavwSAXvprFmqF5CNZWVLrWM
yPX0/JA31t8y1HBehAMU8FgJC+EOuokj/Kuh355VYKRQRhlY4SYpj2Ta6OqNTkoi
EcrTYAKW1B1i/RnKs/azaWk8ru4CgWnMxAEVRkHnGSaVKNBfbpa0k6oRBRmCMx3g
eH5lPB3/xA0pRfon2uNt/TbIH0t0CIcxEyM61IaWMlKp1pv7fd3ze+AVxXizf+HO
nBdIFK71n/O6ZlkytJ5awHHSW2/NgQolRtybc137dp6XAN1XYmazV8FJhIO1u1JT
JQa0jZ6fW9LSTWjJxStO6ykE6f3YImTZq+T2HLLtzIKJ6mwOzd6EsCwkU6Ce17s9
2qNsyxR+6LFdhx8kvv4aWcty65az/5ey5rn1Aq5XMu+iisZH0iEfKHN45ySU7DTo
Ai/bYSTmRLyOJ1zjmjgRNAVXDNoZakfo5LZO/AU5+ZKWtUBpvSdwGnWEasc0SvzB
V2ANZBdxRFYQRUQSZsKgQlNbCIo9g0WL36Wp7Gs+dsh79vAgqvoBEFSbEvTrsqWy
hFDC+LXV8ZKrp9lBUzZ8gx+LsriUlr+UaQl6MMwsiOO4/C3KgVA8sgaRNvlbG0dO
q07IGPIJ+Z+ShpCIW+lsR/H2Kqj3B0Mto/Dfz7GNrAn9ZfILO60pl25cmiFRt0Wv
zfbPuT6gYadqQEIxFx3XvcqftncHY09Dl0O2VJSVL3gPsN+JudHivf3RnSrMo8xb
MSDssF6L31/fFR83mmLR4xAgtOP7qr8OFiuHQiuV54JH5g7c3x7tY4G1Dx4YKXzS
skhPXvaVvkVQ7OdUAbMCJ66e+y6CpUZ5LBHxfTaMXUC78tYPqeverieCsqhafqFq
ayefBXtRPVVl1knFCDZSdATCQEPcOmlkr/gPbJZdVnyfK1mlkJehaUWHIH6b0ezh
Tx09UtmloO6aB7qg6SRxOaqB63FO/srCQiWHT8H4i+KRr/CowD4vmYOKTIPcKuUm
Z0oI2LjKQbD1GOi4zCQmcSLqYh5Dx/2UdKu72QiGtKXsojc1vyu2W+e3Wkbhdctw
VVJIVqvIXHu/EMrw4z9u24OospxEn4hyPLnJtcLCM+4iPoNMuppZ5u7Vu8+fih25
NuVpFl/sNKiP+wrzTWZCuu25TUvtftT2VvQrB0Kj3vBKe1OQ6f4HTzvl4j19EgGs
HTK0NVCeuPWudO4FQkmY8SLbHQ09xlHhUmTNQDQZhqorXBww9MsiVl+4ZNOtk8tV
RjlOXyjiGDKMU1hqX8R3kGD8uOezrYIe0FV8c8JBBxHwAW+e35OuROQxQiAJit73
CWP0dBOlN5wolMPUe/EuhixMlYF++s13fuMwAsnKVe/tdqi1yezhfOVUfYsW/uyT
e7i2UmdKjt0vdwZg/O8F9iXO33KPStNr38pcrkxedpRSTyKVjh+8vIsJMXwi7JJs
vUl9bE5Su2Upfx0j8ivAC1jZ+x0uDItM26K6qS1d+wH2jDhHy8Uin8/LyvQDplhV
lVGKNH9Il7yQSebsDcHbzQWCQDu+aE5Y7yCRxbc81pQPRMc/N8RTNHXVOchKBPiu
grRHJK3qkAQZ/DA+DmAfT60fa8bbdT3TkuQcgQ/FaaGCVhIjSaiMA0JKIIDLgWJe
9qbPpxTZ3TKKpwepse2SJjNUFU7TGRRrSmpvyRBWnK4R1nGI8ahWHZ2eDE0FFWg8
XaWLqAGZS5Gw3uZ6o/TEWPX08ZHkBg1jg41QOc6U+gYumb5CD4oAGJ/HAiBneILD
qGpCGc76sVNkW6bZq9a0lI8NCXMipw35BBy2X7xRSkZL3gAbqok9ep/1lkYilbs2
KObf4QIdLshyv8tTZB9M9tasjE6bQ1Zh9BcXNyTLbMgayQA62Q11pnFUvuDgfE99
D7VrV2Iv0i7nbhSAyzy9m9+jpSZ5P6qsFMzj2XFxaBwIqWnEeKjotobhd0nOf0GD
Kpmnudbz1VtoxwynE5yq6XQe0hhOZPpZ4XrXHe8oEnH5qeJ5ht9lLiwJycW/ye+w
ObTrD42wOJwyN7VoUDu/av0LfzJTpjAvAzumikRE47gqt3RnE68BxyXTnS5NO6zF
/qAJbmO+D1GfyxKBc67k60RBHTR1aJsvEeMZzzmmVInPYML+X/ipE/hOlqoCrDW4
Hu3jQPNnvvEZQP/EFwrnfGZC4AMNtdAbHluxpyZ5fKDL7ezvLL3Oy279sA8aI4qn
CwtOeebSXfjvckc2ls68X4imlR22AxGzzdCFF0vOLCO0nmL/ixfdWlgu3hEeQIma
gkaAfm9RQQ8eMSyDODGZCkw47kTB5nIzMX/tmrNTH/yKX3QDr2SSkSiaNXQuj4Fx
X+mI3rvKUjPIayHFFUtmUuVt1OIw7QKD2GhjRcC/xI63ZvFRSaRsc0czeVWF0HES
DafJcudCH9wETvwZB3ddiygsoFLsXmnRgCuuFP9E7gL3pSFlm1D4M+ra+PUrzhvB
qjg9grxgdyPzRrA40rg7dLuR1yZ7sZdSNgUrBtT/ozOrDaYX5ivOeTPjHNx4907G
6CAFAEz3ETVS1VqGyCwD3UYCgcBpDSGClTAd5pJGsDuh17GDDg4+06f/rCAigsor
Aq9EACYEzGnu4rcxK5I5kLb5AcUgcvsHcA9+L2l+4YlYVUtBskRlQRPzRgW50YC0
DULqYyoVH0QtTBJ6t9ELRovrTOssEPgOFNnt0begdXnpavaTM+AqlfPaK/Y0eMcQ
VQmiq5LmGuW9WkOgaKHNDNlYTy5r3oSUAa4bSFhAZO2wnS33dP0Ad0JkVBTsi06Y
ISqEtcLp+7dyb1bfou9gI3o68cI3AcafK1AVFHkUKfJz8PoXsrPV102G76APFkS8
zBEz+kAm/8Gmq/NO4/bLulKgeTWg0nbTiSj+Srf48ZDODqALKcU/Iy6aSOU2HjRn
B9pa/mYjeQ2M2VHOIJsqV3fcB8dqfBLIrPxncC0KZ808ELispPNpyt1OHq4RYEq5
YlraczNeb+UJBS3NOwE+ONP1Elzss062uKYz9jSCu/4NzjxhlAt2PUVrL/K7eJ7S
/6SW9nhNLdA+Tbu5QQVXs+sFHXn1UrrUQS3aYdvad+rg2voUaJ9x6VEhnA3pBR/s
9maB4p9f2dmd1NHFfb1iaDZPSBdq5e5SJ6Eg2Q95P6k/8Eme/tOof/55eUSAY1S3
6h99iFS4R62c6UFuQLw1a27Xb/yqCBBDAxHOYVButevtxagOQxQTp68StikyZtRF
IVpp8g6cVY1uVW2odchRfFx4l5z5lc1dVLR1zG04El+tEFVkcwECj+S0+mJwvLaq
HsiQo2iBaexASkHs/eJt5HT9HBo/HYfzcBOJhMWOYIEGnmTsOoJ856e/icN9dKvm
mxVLzetbPdHOQ+ppl2t6HRDn/JG4NUI77V9ItyAp4pwh2YBKGCEbYLirO+Fa8+6W
Ufi4o325Sa1zT8hrXMKzrO7H96VHkpzUoKlk1Y2k2AFWkX5WOMeM4lNuCGzCNuG+
ikM0t0fv/3DnLTuvQb4+wcV8BrCQ29l3mlVAwnqkvxH4CXooZvfpRRhMASuqg2zO
QBM1syjJ9QrnDA1EHIPo3+g80HMCdGdmP5aA9wLrRsEO0My+Z7tBqRX221ZHsuvK
AsUWPZ6PlmlfAIKsVNVR/ulIwC/PDiqqe59tvRNBROUNoMmdzy94iH7/cU3hKPdJ
sWAWM93n/cfm3XwrZPOmB11Hihn164Um0zCt3CP30Y3LuYRpu5JFutE5wGpOG3pK
P45GjriCK6XLQNZYFZs7t7difkK56JJfG8UqxxXKq6crVLMSZrTKJqTxXG9bZgJZ
rfNfjZNH56mL4T1CbwpSRfQyOpGLuzew8vuek0dh4Vtu6h8C9C/jkalvVtReQB/E
dcARWC9wv4FMt7C3fAwHQUvI5EjYdB2pK8iS1g5+pktvaRlpU10KNJlnveczT8Nk
NRDcIY4WVu75qEsoqW2szVYqmAAPq9uFbtwB0Kym4T84W/td2deKEJnzcDlZt8OI
80I93F/x8BKHSLF4t05lnuMTsyejhnFRROFrkQxm1pKrEvh1vbJ/jnNnlkm22fuw
LJPv3z6wBY6OkXTTYLm+xaFhbHPkob5kL4MEbGbhRXSUvZcjt/DYx2hfOv3vehe0
gEQWyGtW/5bhfcqJSiAfh5Y8w4U06zxzXcMt1WwdIguxV9u8X4zqof7sryzeMZMm
K6YdjIMqtPjhA0Wltbztnq5Lyq2InMQ+/b2vxHI1wOisbqpyj5pSMnCGzmn1T7W3
iGysgAFh1kJEkeL7u0IcjekmPoIuICe1RJI/sr0zdgoOBP5qqulsBzXBkKX8xFXT
6/SgKLMC45bvRY+SKTagGuzjUbejhMs07tvLuDPihTeQiRKppsPFd941ITovEziI
qliLjMlDXRCNMUZUQkFQvWvaUTw6TsiSjJa7bsSMBHFUB6k2aZyidJhstGA9YK2c
6tNO86hDHdkl7vjMM30SW06yg78M2WF1iaKYHrY/zvesBv+lpdbmmMfg/CdD7STM
oXaWH8B8aIAebzAB1rNKSj6mhKGUQ8WPO93BAP8+HSN1GUD7WWhhtMLSdTOdJDeW
sFwlKkrS40TvVSCFjczi3/jey//qEPLb2mT2EhSFJU5S/BHeAJMfeaq/YdyIlz1J
DV0xx4zT2L1WFIbDWoE9gjn37KpGTVEKkd2WtoHZCqHxRzXiVlSqj3Pvwzifknwi
WDPkwbKJh564jrlSvx8GqeYKJKphWYXJmOO3rGHW0MFkmDcn2Qr8jAlJWkTwbQLo
kyG+sh4UYTcN+ZwE9FwXsozCYC3Dwvq1PZuaGSczbt8rrqBsT8on9+3mnCSainIx
7+D1J2FW9FSScGt3SzMWWooFilDoui9K1znQEwA2HkVQbUx3YRInBwMHEgIPAnAb
zYcf61KeWxBxC06ixfc8i/lBfkudVI907xbmWgdF2abIRFuvu0XQWNyU5JY1/Y6c
wST7SdsAkevVLm7RhnXTV5Jbtz2VQ7YydPzJ+A6FYnTB3IMzJ8pFuQajTZBhmNDC
m3Sx2fK1A03JhCv0TIuXLSUiehLDk8EOWKBIgxwECm3892rI6LwbAq5TGT7y0hBh
CTjdPXO3Xuiu3P7ReUqebhmeoR4+VOH13Ij26Msnomwvd7447Sa2MxrNKFPS0Xo3
lWfU9TMzLreyFgtlm2hr0bOg8butPzlXjwFtcVV3F2SIOhprVu6t5E+F0NgKv4DZ
NGSHL4Vn0+vdpipvec6qaOcn2fhAh/EbHdGgl7cIH5I+1PvWk3OmEHnppzjjYnLF
YjTUhf16yBvwjou+qWKhqIHqWhKutDDM3iqoqj1mQpAffvuYutn2RiKp/9D2mrvq
fFYoPvX7y0CUQcoGIaKlVSZQ4kz315sRYHdhANyZKi4bfowXmz9XINqW/e+XP1NY
eep8Q2OroxDYPMLdMdLiYtcWG8nTt/WwqaUA9M33HaqhAGRqlAVgwSltEKRxVlWu
7TMQL2nBFHCM2GsK9fUzFP+6qVpc24O1EBjDQpNO9xya5Qw8MCySk0rX4RwqX3UL
vl2/7uK7i1V7TGaZWLghi7hiIo8dTPWCiEy7ha7631v2+fzRYu76UlHSrxdLgwIY
Y2rwA4kPin6VlrBGIotc2lTMgVFeoOl4T3IEbHkNywjHpy48KwC7ej+PzhTmW/W+
KOn39PZ1SZYf2MikEkpotuYpTDhfWu0lICrXKXx01Ikp85I0MlTnYuc5TXX5e4oF
vHbndQFv+UY7WxcY9sCaPDIlgxly00w2IdUjHa6mszVHLGOHS7YZojuzOhMYZqd2
NJXWu4/aGWukNBxHci2KoBe9DTGFNYR5zPxgFWYdqjb2V3cfwDliMFLozZdpqEbj
FUh8QNJsmfEG4nparoyuwgWtGi4l0XlDeQjDvFWVCsRx6+nO/VeEL4bXMDgFZ3ZV
GbquE08jwtXTL0GOXAgxnKr/fpKLP41AaHtKff4LLXzZOVg+oYSKVg9Za0oXyQF1
WWedi81ssywwDZitUCA97ZvEYAMpUHdKAntaPF0uPnhwfh2GxeDTj1/QyoFawGH3
vvQMjLcLSGR1uYQcY2Ss1CFTZMEQdw9JUw7eOJKDpackFV70T1ZEh8Y7fFl8vort
avYjeuQZakUMS5HkVR09mPO8jFpnT8TvrNYXoAELMDzG7DOErhgdvKiWpAQh2LA6
BLpDogTz1HTPCHhC8KfoRUNPjCK9kFd5IcmZydkbHVDxxPS3pXn5mzey4+Y1giJA
T7w379tI0m5I95/IvuH+SAzROlzjvfa9rkQVAgW9K5Kb5FMcYaYoP8l4apIlQPbb
veeUELMyJvkqpTSS2S8RDE14RCGFCR+jzjhLrl6gzQRV7IUPFi60H9IHpB6Ev4/I
+A1TdMmPgH2SKOsTRiQkX1TdIAWoK8tHaQ88l301/Eq66BOqbJAjWVlWRqbLxlom
EvyAd5l3d+iW0YAd5LNu6rNZltrtvYlZhTfrSZN51rf6Z8igPR1DrQXIoQT1Mrtn
JoJyjmvp0uJsInD9cSF1Xonp9uh6GjulaosbqsoiPZcgK6lEEmUSN3LnmeJSItdx
4dyix9BZZbxHJE2cRtP6/DclDzNDeojmEj+FbM/MxkVQAQ8+ylvYz5SU8TCfvMCz
Q2owGt+bkz7Z1FWlEJvkgyacX2ND2/JdAfNFlSc1Ge4Tm8LgC9Gk08u56d5sxWF7
Shp5aQdJafjf3ImTPobL6E1qmMIXR2rBRmmrTbtAkK4Ya3TqzR4D1j1EWjhjE8pv
jpf5iEUHyrJVKo7Jm5sEv8gnciStEfPV2HLR+uoXpJ5mupCOCnnMM0Ty75Y0UVCr
7jaqsaTqkhrAOsPMz7FSVJWXnNg3qJbXzOEJaN0pVqnqtYlsVTkQW394e/a6IlMh
f7gER2miIFM8sKI4e8mybGqg/s6xNoeDH/oyaq2+20/JQxSr6v3x1Os9c5Q+C2Wo
WG2Sxwe+czIEy1Kg5Dgq77MvauGyEElhotNj8X/2V7WOoYwXFvY+kcbEwcAymWUU
1LVzpZS4f4e3bLqQnw5bw0V32x/pcjfg/OU/gxLvztPLw1tsv0oOfFGppPRo5eff
4RDqfA/WLLOuJaUJR7ZGqZsuagSOb9pjWLSa+qrlMCTrkzlRSugNpeZHP85cJm9x
8CUg2tEp++i2xoEHghoPX/GoBOwoj96mDNqxsaVFTzZV/zO6GVRXyzTpZDtbXXlA
+tSuhK/3ERBc6WVCHSJ+rEA1u4DCuSnEkH2EAECyO0ENdzv2T6TT7XKRi3hkkJqD
6sO35DTz+Xfrk/OIYYeInYeFneHGa0KnP6FKoBHyeZku/BCjlmq2rfT4uogOB3N7
EFn6Ogx61Ai8D7QZTOdh2fFfOe1Q2w9eu/PwbgoyifYLSIfwdXuRZPsTg8Ft8Itd
x5RBKyqjUDNK/Fdv03OPDLSa0lobXU/5MyHcymAe7IYNTjva58X56eE5wOBwbgve
uSoCAqS3QCNNcruLtSd/QO55KktrP8HhuZ3qxuhC6l65DrhotB+6ySwYmHitz7mP
EFbYLhy3BQZQa7uYQJEs04yDBJBy4X26FO7Rh3QORZmoD51UpmcLpyr5oXmFLPCz
8Dl3pS8cRFzwScm8hI1Q/3L8rjwWUr/a4t5NEzTN9svUuPXbki2VHfbkKchVYpDI
XWlvIV9LGRF51ljrvn6tanuj9Qd3r3fPJ9JU0bd6Rj+T/mvSx0inTloy7nQTp4YS
4NNnvJRMovrwrAU+i8rCFqgOJ8thX9meWJXVptqwT0FjCmpwWno+Ta3+wI9CMWN2
CPqhOlHWWwcm24Rafoa2N7c1A0S/zejmvhhTHtyAtadBT0z5F+x/NvAj7tJhrM18
nQYxJVXmRSsxyGvirMTmXn15u0OBVcU6ULS79r6hj556jkdKSRe/frrO77UJqMy9
amSw24ADlgS1kHdUJlOejtYKMv+blMPbbWii1L5YriAiVGZrl4XwU95E4OOPf1Dl
8ioWLN8dhebwKX48zvTwy8T2vW04nOGLpf2oqkUM7NFg/Z3t7XWe2aGWjjFstWlv
D7bXo99fb3T3us16AQrgvDIERIlnoN6Iz2oQREbL3nQCJkO6HoekU2mf4KpfCntv
oMFtGy5gSbiQ08edv0vMh3J74wPLklLilIBda1a03gQgSh1ek4686c1o0319n+DF
TrhYjcGHDh/78dF84zYZmMFDLOipMcbuKWX7hwr9GFbdxvkuqAKiGjcaE36Z+l61
Ww0+qpkWSZ+Lta2VZ6ukRlES6LDiPpMoiqx3aP+Mgps93k8QX+XCkKUa0nbn3Duj
1MqfXsHmRWsfJ23MZSNVaEWOV+QbiyUXXvb3hB+W5iXgl3fHaQlF8DV0DSGTE6qZ
SWzJ5NNgJSv6S0pkYxTc67hn0LWfFNiPL5YQ3dX1ozWcuB35sTvFLiSq4i2fmzvd
bomwWq4GbLW9mgBnSwL8F6EDzMLmSQZyCm4NvQOKv6t7niIVQYGP6E2AUlla0ayT
EKaAMCPrd9RazaP3czUqIil4q16F0WG1Y7kqoIKi/HEO8gV/z1dYGyj7fShgLiYQ
QuZPcukP5UtYAVoKLM/WUXOPoH4qsNZmRjYchZiDragbCf14928yHSpzj8lAHowr
kRULa5sFgMrne6E1330SSSKyUqLcRHqfx3HxvXMOSz4YlfBclYwAMunqK6O2CqXG
kRm7aB+bE4NAYO1ppM92i3NDFzLZTXbmTUDb8muLHhZCOcAu5N9DQkVGWcGRxd/7
Huh8KszhNeNIg7XjD/iVyPCwl3rXJNHT/6kAQ+F39xNrpll+uaccKi4Zjv/cLo8J
nhSld9UjnuoB/ucIO6hjTHbTiHLTy1IJtkW0ESvcwjnk4vxMmARPV3Q4e0UKTOwz
o0IUZxngDWeJLYxk+NBzruWq0eHRK0Ei4YnFpRFT4ABYVyZzbImUFtf4eKoqnTw0
qMkcYZuxbzi/KP/9Z5uYjyRizBqButHz+z6SW3CzzcHekq4bKcg5b1ES/Nac1zJf
EtwZ4sk/Ui7jvQtx1wcIRSkoYGys59w1spsGezX1YG623gZBZndBzobS5Sa1r2yc
AKTjplcr8PzUq/elV3kn+xX9yHEYsjGcLEoCQF4atWIh67sEPbA8ckQ2tPXXuvsC
FB+5kKb+bT4RcTOcbWbXA8+ePC8s8/qD9/NlwF5oFIcWrjFiR6aCv9CDhyxlDsCq
ae1t01DwU7fOEsJt9uSWjexXtXxx3Ddmmd0VsYgH+wdc4lg0oXho6MnZcdZWpVkR
8OiKjJ6YwyMR/vYLGNvkUjA4DOeHeh+uhGeqXFQ9zbouBjxezGEo3FM55gVaVjS3
vHcTXEObwXbrppIb5zxvmvnU/b9ulsmBqf9/d+z7OyljtO7FivsPW1MAuzcLybBv
0vFtjbzLt8g/19wyDWZmkW/HknL3ZPILul7d12D9g+Puo8n6+WpBmTl1NnVg4jxy
Z+Aqq2gosbmtzsKH6A/5zB5KGjknKTUG99YIQx/C6aCkrpVip5TZqjHn2r/qVV3D
e2+0l2FoyDFB6gViu7am0aHk6hxKJywF9Y1fm8LGm++Q+La50LmtmjcTxXuOa5wG
Mh1083v9gXe5ZLJCrcONdu967iNuTTSui2wT0QADCgibwYnoyjtAjRUYjTrl1hqH
gJ4fI7INdZGSyXWUP0gASfFwHaeSVwt2QjGUrU/C6mRt+WxqtGk66uX2RvYIiEIm
sIeW5PJmcYlFs4gHOxCjPyX1fynsYByNZf6jWsMlh0WcqqiXP4jpEvOewSUd0uke
MJVP46lukL7WxOPSXJFaE25H9Gq9fIggqGj9w6XD+H6gjYHVPohHNd2Di/VBWSre
UtMXfkuqYWwUps8EQVmohnoBURhVh2Iui5CnmPGb0zbyp9IUFyyyV1k8BycJM7Ig
gTay/kHLxs+P8q91TYRuv9m/tT/5Ax3JOU8Rs+9RinOJY4uWCyLOogY3eFIjFkeI
A76iXVdyjrRYQ24HTmIeYMLKL0ahgyfyxaJzmsNsB1wJNwnqzN5gbnNGm7WRq/1J
HJTb8sq0M2RCoFrBiEBZle5CZ2OPUQVN1jlBsBkvPN8M6I9d9vJbnw3rYJSPo6vq
Vvlz+kgBoP5rJwXjiYnRhnfl3igxsylNR+CpzWnMAdwdEJVl812dB04SJo+jAHl+
YJa4aiKCpkcg2pE4jM7FJkQXeRZJLeEevoADcUbPfn5h4chv2PsOmF2lfK+lC+8f
4ZLkJKUqoHsPgFmY+x8dmYonBThVgr94FPk7aEtMMp6eS7rpf5IwiaOMKHhayGR7
x8bDhWYXI5soXi4QJ7Lh0grmxzbM1h0WyEeRZST0dwddS15s4XHbbOitbLmwggdj
s/w/jR21b0BL2bRSnI7vmV6TubeHYTkAKgpKiDde+dQDFPgoxr/chbkSMsJ6U//Y
zvwyFpyhGRE22x4lIId3RpcjAq3ogpRQOxQMIGcJg/pMzrerxdxpjvfUhAm/Nz9M
HjxCFCMfIDwnKnKESDc44S8/hVHSaN/BvjSPF7wqqcm0HFk+qrmZTe5PQraSPT8R
eYYK2U5jU1Yf35XdDRqhVWKaRaGz9VYyokvCmdH+fe6hFDWoQGVDll0ASY86xhGM
pgCiKGzXjo/l7hPImHYKSv6Fu8lvUki7ABPT3RZPoSj+Y4wVfrOjloSAoxRGA8rx
/M0cnDftienWEDwiovb0M+aNB2ijz19HSgZwyYVjE8dlXIuo/+EIotuAXeGg/CEM
yGZq741cy3s++rqOBf1bjyKg2htQM4aGJsHg9gCaM4DC4LHQyy9a5qH0DxL+vmIp
edDztA9G+XtmPmIf2RgTgw+uQvsBjuaprG55rsf5f5dG1ICGoxQfJsX4XG5E2xwk
2rta5S8krEYqqN/iji2LG7xufTSuyLikmsB6n5sVWHFD75aWG0fXm/g8p9bUBVdP
Mes4Ilp4S7RhKSmZE9UaGoxgW/Ef6wNIOaMVPv3sLNqAyeCIuCK9y1YpoYGlpHVL
AsimWtcXBgV7PlcEIwGPSLSTZhHM78Y0GmKOo3dEvnrk4NNSO4EGimJ92oAsdorw
pA8H83XcboXnmwGUkwQTqlyWcOemECp4pMT+h+R7jUbiahsClTyMxce0SAzbaodJ
O4Acr2VHgzq0DtEl9kqbKs9ZEaMMJcTx8PCMfHTA7bJerfltpWCbaSi/ftrALmYt
xURdaDqe0sESvhNvzy6ieYIlDZmdN1hkCX+IXgZpsCGRZFt2KLJKfHXCiGi4KGTw
gYaWv8jSSMCfBBkYw0jwm8z/RQXmi7Nv+D0sTVmro3uHpjgLzoPQSQUjEbRRYwXA
7T809dp3GpjhcF33KtGECszF1cfTZLr27aVK54mLyr+/ldTT7D/fSuN7zWukiUj8
DHzcGRZPWiRSRtBqC/D1lRROhfPqTcqnc5Hx4gQgZTKjpJPtqI6uyNfKl9KxyZM3
zOFfvoZZ1HN8MmfZdHqOtgbDbfuyiCIZEbXrQNq8wKeX4ACiY8AW2sYEBNSsVDLz
/L1nN20B/Bllnc8kUiMJgTwt3Hd23AuBoVeCD3eQ/Q6aUmO61jHhJn4SoN0257NZ
Esa78VUgwab1oj+r9TxbcxdwutPRNrRletNiRdhwRR71x+GEP2OJGkhP4CqcdWQz
V8Tw1yzFh9tAe8XRaIU06uYsIRHGFk+OIIPXaGgnFrcccWT6ppt81FU9dkuAyaGA
mwISc5qBvWAD3pletjNznI21bzNfxz0pdDt20IlsfZAdMZzCKNdm85/c7oFCg6Zo
dzuG89cEbxmJJz9ply/4m09/oPCaV3BuTC39eXa7gTqJtkqiUNTRq4yknz1Rl7fK
ZiMYwauuMr4Qg36bPnz5ceZ7ANEprMb9LbVe282ckgZvf3OdbXV4p/XmnmLMXA43
sxY7I4GNg1GIa3W2mKvn29dfs62UgXPQTddyGsDnfXy11UQ6UzfZPGQ55/bjTej9
DhIlooXAzqQw3WEippWEmtdOARZyvjX9aO/7eTWv0xcw6Wf1WHku8uEsZJ3DGalV
Ugrh6TKcjSWOF+0L1CudmlP3J9HS6y3kSFVE45v8QODjVE9e9tGlx5ivOeuoCZbo
OQm3e6eAnsvnXwsi2WRcbJ4194DeB64tuBI+0N8ih9JvHAzZPtDWSkDu/Sf0dryy
JpG99SRsNz71ZzBubspLqjAFaiJOW34TyPMC9h74v2qvatVSO1zZEbkNG+itqWdQ
7o8dI3ToYisE9fcoChJd+AEkFjohCp/f3yqBmMpGE/JkElTR20UoFDw+XazJzqRZ
KdrvNeBQOPzjh+kRlLyBlxFC6Z8DDAZq4C991eh+MibUnoMyb+Nr8ateS4i8iPVp
0er3A6KNG4d2v02ySiPi3sk+hLle6ozTadc06i6JJ4p6wkrGx5uxcx2gv0GtGMHz
4F5mzTcf+ASHEpNZHzf8S4KVvNMavdJW/TxGyIwMEsUQAS+D3Xgcp3wOrtTi4qPX
bcNsl7d1CXQCSRGaMX3udhFIvxsWs4nmNw1yuTKXths6do++9j19boXRBnaUmrEj
Swsv9HjR9UUHCf/mTI1mrwxl1aEF3TMoRNxYnNebc4UehtUjUw6n1yAvYdqnBUvO
6nt84Q12RkNyFv6+qhVb0cWRkMF/XCGzi2njnerEUN327DDIwtc4SDaOymGTs44v
Dld6DCKskhU/Wu3e7yC//okBbvfYg/NMhx5rygQKA58FmmX55Ge0epegELHcEOzM
IaL7M1y9QHUUvbUSCFv6bN7+eXetOqUeW18TzUGNsXwuRJH0FtJWIfcBRgJ3xo+q
MMCtZC40VuB9qkw6kpUjRQFotzsZl8+TLKULDXEo+YyaX6xd/bB92v1EH17b2I5M
FoSStRMA9G9gaXevSIckl049/WQtM/FaGbTZDaWD/BrW6+tPc+Q3oItf7xZtUAuB
uK44Q3CQJfwSGXxQEesoaJ8+E1wsZcwC5O/ok/aHExkTwVmUpxUYNfcXnNIpp6Su
zLytthNa1J98EL4mm9uiuWNxsxpndUjx7cdRN7VxBLvzQeByjJ75J23z+ksuvqVU
jxtjpcW3L+HoJh9QDf6ew5KfikGAQcVeUPDNdX84hwyT2NzEfuroRQadv8fp/MQb
zmSacUoiQ2QdnhNQ2v8PU29n74yngd1MrgT8tSyRd5WOlh58fmQN1v+qKgSCIQ8k
LN+dljUsCz2B2lGkpG3lQg2WEAv2UorbG+RVyZd49bpRRAZu14NzsbnFjbCSgt51
E2GNMNMSdobzYSdoxpRrzoGHwZY04j/clDPlzZvmSw0Rgc1AjwfEYnf/sqRcT3ov
I4U8xRUi1GOwDyW3GVJyuIw2fCzN8HlJnggvEPDDM1Vdc7QeQ+WJnw6QKUoiFOt/
1ZKjsGWF39GP+sAqZIcL8ugM7vk8tCINjVOi5oI7/zB92PowdJNw4M1J/OBGqq6y
v5al9ERJnbs+zvW5N3pdKHPlHQRdnS6m6ehZFu6m+N/fEaeN106a5uaBrJnItonU
cqN15cVjCAU6GIsS7f6QHcCbccvhoM9mqyevthnw9JMLqFwqqUuhetlkTWsnZ5vM
AIsMXXD5Nz67WowVlfHgVsNZ7MW6cYedCbj4f6z95eD/stD1c/Ir/t321fu+RU+j
5zp9sIf1AyRcLGAVgnnXP4TBj/HuimejnYoE6OlyDuX4zlrxo5D7Z8vjTBnA0uOv
VfGWPxO2DeSF5Yl/LIE6onjS3Qkz0K8tWJE1b/Vx3J1513ouunnAU6UBFiItGNLn
OiGduUjO5O1bqDxPcfZdTAU+aLy96MpWqhzWZ6SDZtdXgLGOeADlC8ta7zg7ij+P
OZj5UkA3UjLCIDI+JE0OZq7Fp4rrXDeLvjfZihnymQbSEOHsFvl5dfhc4HeAipfd
rm0dIBnSDjUtjjQji7YPpV3VT83zCErLU41op96P2jIHo2vNYJMrmoS+du4p97aT
Xe+hsQo0EQEUy7MUAd/AUhgP1YacKuP+8uXzkuwcTGQ7B1Eo5AMhDWvlr8niDELR
P6NuOcGbRISEK8nYIBDPuZCBmX244z3/fiyTDxkoooB35g/HBfOlQ+38aDwf6C8m
Qs6NSnmYklYTh+OTF9LAy892leF7BtNQkxg2a82oULzvheaka5wI3ZqZ55SPh4Iw
r6IGu4fnS7j0KeW1fkEjVAF4ITi7Ct/iMST7S+YpUXnS0eby4230fFsyo5F2+OEF
vlWwiSVHzQsVVgADa9iZiJU4me9Epj4dqAKtQibMkpWNKrMMiJ03dzOKFyfxCCRe
YCjTrWRyswWDSVPMn74yr9bKCK7ZDVzD+EpUH5YAnK5yRkzmcZtKUX8L4V6Kotd4
ZAIv9KyxdlvtS9NyENSGqdFkeTCp9ycpRt5/xxLMbM0XjEQ1PNBjcu4wqFy+ORAc
l+rWzzMASjdaxpY/bTGAPn39E6xTF61k91Z7Fek/dNQKeudYZluXGbm63vY+SX6N
JYViH0UOjYeY9dO5A+UeYSXPnbSjbWhTcfUA1s0VkPTfgB10GVGBZYrruwTL+kxi
C0bAjD1cSEH3nBoAkGh9hTj0wNGWftb4OlxNQaiKD4274KaAfWGM17xVls4omNnW
SqCgxtyoL7w8wA8l+165drTJEtkatNMM+1Resi95j4euRx7cPfEWbdCeD1EOA/9b
/MQ8mXa7SoovDKiu54ietuuBAqDKEmb/T6X9Vw86A1xsTfyVSM8rHHpMl2X8vHYl
itNtLSNbTouxmO99Yb519Ztxac+CiH+hNI5YbJoSHHtvJmQxxfVT9R56MlpnC8L6
gBQhtihSehXbWdyNM68yIh++xXuF86az0rI9cZrc83gy4AXpawMxuLgySvuqH9aa
kxpQEG+WKgtxcKwdiYm0fjlEHr2wQM5KamslhU0kt8DZtJGSBq/HErTkhu2ZLyeJ
JVU6nNv2BtuQ9plNP38btTnUrY0fzURiWk0anBH4y2IprVUf4kHfmRRCIvkMWZgp
8ZzvYOLAGK5hXz62/c5nQJqb42f99MlbPWvOSmUuXlsWLusOvG5O1dgtoo4S3WhM
xO7ypY5hQ/1gvRyC5cvIh7OmxM+e+u5ikydXNnlG2J9HiWKn2nrxLf9dXisEPHRY
e9r5hM/ng946uYl4IsiP8VsKpZv5SM7v4jg0ALW5amqEP6G4sVVvesGEJT6zeSuW
qUCoCOksBuOx/sn8Pdbb00eFxflBCREmYhPQ414xk2tTgxwjmiPKoHttj/kYKNVg
jMHSHeOIzInE+Ri9DipnCsfxH1EEr6sZxuy15+YnTZod+vbAZNfw+ndQ6nGIoMeq
e7W2wmC7RMHWm/KE7P4+A+wlnwkfRNsGGyQDG5NbOCtn0oo15UNgY3tyN0Hzf6yN
A8J+wVIatv2qLIrDdh9EPGv8KvAPfAH3X+9XoBzat+HxOfPqT9IXX0W0fWtxXZi8
j+0QB0ha5S6x0y1TK3JzHvSGxxgYUpx5vvAfSGDVZtvGWkOwcEXwaBp4YFAQH/Dc
cXr3ry7KBlz8a4/phLZvjL3OdBceIIJzw6opDRsGRu0O2iXpCeJDY/Mz59q0Ozgn
TB0L5fehoSZZUUW+yOWhl8SQbPUNsjEe0yZg5DeESPRx0mE0G4Njmi7RviEiQaPZ
9RQLkZgZjspfmR4TkbDJhRJKMQTikPZ0uv7Me+TVJu8WkLW2vxHoBSNNW3u3WMA5
yKzd/i2e1nHTnw30I67IzKYkfUKz5bngSZFQgR02cY3emGwyop87IxzkGKegKZCA
yZVvvWL1R5unkboyxj/hIABro5SHFH6w1bKLKxNR/mfZJII/0WqP5Q4CC3Fh6mG3
oD2XLshQtZBKLLPx0yeqnpIG0UrdjT3XHPN51HZh3kelfv+exn18qLnKNLPYHbxm
s+wPws6Me2WpWhBb6eWk+QZ1b3YNDjOBeB9jbqdDl9pY5gROTn4LbZ9DVDkK3Mcf
HTgD6lmbr5ehdMj/jk9DoBBjpFzFsMEDrNLrlPXrhDZYcE9Cp7gIx0Z9rwXoPDBZ
+PnBOqmjz7aem03RSAqu4GG3LUKEgHaFxws2XTJs8A2y/EYj6q3zf0knG2FIavUu
1qEy5rsiDIAyKmCTOs82+oxlS3NMWnECjCNC9gfkxa6ztMDMXxp4Upl48bB+Wni6
tBqOVhGXqZNi9mM4TOhv9knRecibTaLv9a2O+FVPraAsrnOxNFqZ6kqawtCtwFEJ
FUp5K5fGs5IipCuQC1hdsav/0aOj6Rzo2phUdIroSd+WTqRYKi1riCsW67bfhK9k
ZDrV4KokBInr5a7ZM16iXB/wFDbjYSPD61BKUrbi574uyz5e6t2dftmQMShMwhzN
7iiUhTSVtbObdO85JA6Juwd5RJO/ZNR25vzc8OOqXpFprTnsQyaonBDPXh4h3kQB
9USZXRXe7jFue7bQGhuoYAYFyuvLX0xRGiKr4u6dmtiLsZnQJmqegmxCn/OYb5ME
XYYlureutlqX1nAS/5Gr3PNXFaU1VHWFIBrBkeiGLO9uUcHFsY47xyKC660Kg2nS
mPgXXr/zbDxS8CNOZmWLnWGa3s8bWZDlhACO0B4XRww62yScGGInB2fmAU1MQbb0
W9Ko0PlKc7oQkmKAahchvH/5QjgRPTehFyAInrNc/FNKh6t1xAVTeHv0X57tN04N
4DnVS9D2jAPZWuEO8cHR/47i0CXxTwzpuYvsnDs7wx2HOi+72sJgxslwShXLepkE
PBzz9YDh2ftiL6yDUcgXvMPNGdrz4KzX1yJg0vYx01Zx9rdjOd9UgDOLLnHoqHgL
uKexVvwCKLABrmBoQk4S2miyzHNA/DqvCWPwBcpZaj8+hYS9Btg6FDbe9m00IEhI
uYslDzxTV9we8qIr8U/t49leC66KpRR7csNanCbJU+382kA3KNoVahxsLeIhFECS
F7OH60CgTk7PnZLO44y5ra7ev9r8GTYXy1FM22gBg1Eud9J2Xc+DbR20UPWeyGCB
Nd4n2uqDGzPsMhsd5QMCpRK8MwM1P5wUWSl4S1ZrbmA9oIZMSdN336JnF+339z+c
YoomakhlP1di7GodSjj9Xwi/68MI2XoraoQAl2cYiZlhH1J/QHckY4b8NAusH4T2
roxnVVoYX6cJdnSp0sC+1N3vb1hQoOicdBaWsmtwlFmxBkZSZGtilx+sQYg/U40l
0GS4x+1Dnp1B+g9GSHyH+36hrieSc7uRwyjhESckz/StO8APVbSMoPkmX59v0+Fl
othTdQhnRxawQJRo9GYN//dM1iKBR6uGI18r5LQD0DgXrvCph3xbcTNfRpoFBoTL
BlqxGsfiklf/Yu22yKuaXK940BqR4MVVdX/qTvvkfFf8vKsWt/OzMh6v2Kc9lRoN
pxUJa7N8HEZSVjWNKIDCDAvFkVG9M+vcb76SmpOtoirSLZNwdznuPHQ9zjhCWH/L
rTHmpuKMPVeLTkxleCvkX5vJpyU13b4a6O+d/VXC/gBkeKpybP82LQ8ivYlK5Y4y
B9uyS6v1WBJhJ4uQTFkx0UEnAqn7J5nAoQq0zieEdldQRneyMT3Y4eBNd1bBSdNN
Xbz6Rl7e0B+Hzot6DaBkavJLJAuDvuJHESAV77YtSz7CxlrDLnmM4LV/ayiUVj2z
FDyRIimGmyQPJp1xsejRbN8qFg+1vJ+ju1IrRyBncMjHq1W/OkMvZFSMLVRIMKSe
mSq12zWpE1gxBT+ULeCJBLrKtq4CTibmpFEYTEYduTdSTdLhAQnHHJz8l1nAFT2D
WhSedpF0ZYOCrMUmr8MokhiDUkZ5bvsjyV6AnBL/UECFClKZxtZ84UZxR5MA5qcx
idj+ROrUEUEBiFog4xbTuBS90+x4HIwjpYI6Wu2wr7+5rMgBvWW6g6RzB0CxQASo
5BF76ACUCxGwg/1bMJ/YqG1PgiRLjfu8oDCQ//xXrV67VbjSzndetxZ5yVqcFRLl
zOII3lytHwFeGB4jxksBei7M6RWZs8bJxUU52O/Q+xV9VuxSmUtAQrYHP2nUUbe9
d9QERKohFW00vjg6l4C3V1BpVRH44Hv1Pw920mEhNaqaazSaHpIYErnzNCSjx9ow
BUK86EiglyRfaunzaB4S+IUiTUaFzfNLL8sz9yQUaL6FS0YAW4Le8iNJxxy1ywnE
ir0ysQo/90GSbbnj8yLAPMdHT9RrAefDDFo9Dnl9ez+GTcLDvh3nK3Zyg1YelpvW
CHPmAhJEPpd0qrAZE+6xrc9mCz2qAnN63G1dUxpJHApoTWVAUFl6a5/v58ydfaq3
GdlsltKX4ifNl3V5zyOrKupdGSIkdd4vwkgMoI668VCzhe4ygkxdWFXnXe+nYrNZ
/HOzmE30jdWaZbnfwUNY8JHnp7Zf6EN9w2/sAKmQRjDPVSU6/AuCt68rrAMKnAna
x6ifB8f8NLsjzx+F9AqN3bjMmgm7ptRHKhtyHRmFWtSEu+7ud4yz9vTQw9WNm3oF
HTbjEXmw1s43E0viL4D3v051+ozGO/+f2/8x17Vgjti1D4aREFDvsNiOjlbppdYB
jCVCOqSMdJrnzLOonyTAy0plMFyS3iLa6lrKasRHamrveBrl/R944cWD+Zr1ikPZ
yu+CLtDTufQ5S7ypVy8Q9C3EkFuK/Ju1oCLx/BBi6qhEOzPCblVZo0QCOnuWBWc4
qqVuj6gq70f9lz1SQOsa9lrwh2F+kEtkwBMNn6zsdnmLCLtZp8xY52bHMl4KTjbR
bZn6YX+eZ7I7ofID8hkz2ButcliDcVgVX7Ub2wSo9iJFSQfyYtY1wabucM13FVMZ
JXl4swYoBlyYRSDVBDWOQMy08ZHN+zwWnCoYGZmJ+UaOiRL+YNaxAt6hmUSOvYtJ
n5bTC4a/oj06OFRvuUCThhcpLXgsbFTvbTEk+w/hRxWi44iWNdbgvFrhnikG5NAI
l9w35LAQ6Z+vjDFIseHIrBoMWi6EYirBrjfJr+nyz3NJhHOep8YgTE/xhfEtJRvF
0Gxu5S+fJhMz6SpNeTOmtz+6dzY7UxE/GFhLXYYPCTU48rBnF+aHlS4v6ddsYgli
KQd+acDAbQSM8oRfllIPAc2BPBFl6yoakfS9HjVikKaYbuMEt90bQn4/044SVoqr
QZ30gk3vauMHUnldjsZMCUNh526eVRYOcflwsk6MvfrmHRLssSrUZGJaHw0icexL
Od9+neVLRhEA5LgRb8dO3JVf8zNYzu5YWfarmH9lJJQuVJsoVpuNDvfaFWNDw9H/
JDO5sZV+OuutDqQC3YxwPSKm9IydH3Cmsb2nEdA2tc51h3NtGpjUPG8mrVlpkpJW
uPdCfq8enMigtAglaXL//qy4Eaqy1/22H8tZURdChbV6WW+/aYp1F6H5SZY6oHNR
3YTCoIpOZAHAiWqIYjjXC09eB38SiZs1hd0Sfq5AckjEPvu8j9vO3NDgUZmxRZZu
Dgpkg+h8lBgHGMtCPks1+p2i2z82Qyu7SSlRG5tdxPLp78tpx/c9a9EhclNyQzte
90xPvqv3YJBv+gV2qcdLriwCtwuaNFbpLyAJ3WDbGWfiM9fwkN1w8vkSTVh+SN2C
WaKPhHoNUOWa1tTLN/KCd4HvJz+tF4ap4CRkd8kubniE1OFu7kA8zqXIKE49MCwb
PLdC84NUxu/tI46vYrzMRK876agqwFFbw7yGHIEWj4LY4pNfxmQv7kj51A92b0k9
O7dzKhYtowHixBebikAUzIXlYS6dd0T+bdK6/npsjBUoMYT4JT4SmEr+IWcFvWLZ
iczrJtpqd5cpKqXVKE0qbPCrYj+bvb23UEQOyJXWnJp/PxIXxzUiDRbQx3Nksbnk
wBQVAHHSjJS623jy57ckak9gM2avurKE17+e8e8Sk0MqKCbqkcqYRW32gamZvx+c
yJFZEL8nDb1oh9w8BogcQ69Z8/ZD/L43QXDpx2wuZLky+XZcSc0NdSRAO+csfhu5
IwMc94KgB88P4GcgrYiJv+5zTPdsRw+pLmFfthoUilUGjisodEQr4u8qDqCFj39e
bF1MkpcViMOeZez/V8uElgB5usVbfQaP+iS3tyd6YReOiGRJdPrEiH5obyotWeqU
o/S9ZUUrM40afhjBtY6S3CzIn80wNP4EYSu0T4ROXxoph3ulQeGpj6sCwabw5b+h
sLQ14eoOwYONd+Nhul3r+sLifCLdqWQralw57FJRCaz72E0e/peisuKjIzVFapbU
Y+tHzduy9IgTOcN4BL6L4YoDKPxk9ePzaYcAerITgQIcOObkFnHkxUJ00IREBMjO
hFz2Wwl18G+D7n5Ss4nJ0NarqNwSVn8qXJ0rYqfytP69HubOq5PEVZxYB4+WbQq5
dgtuKyWvNSHmIzHNqz8cJf4J4YYUQLlk59EEF0zGpSMYtR71l6TcLZkr2N5do1xh
ckKS61I9Dq7GZhuiLrLRED2FObu/C/H3cSDR8g/ACfz0P3fAthLlrfnzMYsCbjl6
bSz55hBu9ujG7ZcA4Nfvm1n4aAPxuciLHzvp6vxFzPh92MQjGcWddWjX3XznLqaI
Vrin5aRO1OjvhdwlYgljwJ3jaTbrDAC/Ffg41apDcmACvSD3qsnWE/SkanU2V0mx
jS8MBqGP18adBwUUKygd2jHTb11XdQiZM3+EV5/Lqryrj0fscKf/HiU7tYeh77wg
z5WHjvK2p5M2MiN8kRkCahUI4A4rVHwGDS62MkGo5rqU0R3ymbZnzaw2h8jRr8bl
VQPcBPotclOwFcTkvLsluLSKkfACIoyflEZaxrcBPuQfwXVoDlY6M5noQaX2wejj
h+h4iMGStB5P7Xsdi8Rz495yLWu7VW9Eqsdr+BRDxQawggf9VQN1wE+OfjFY/+Pp
XXvtsFeFFNnJWeM7T2pVNGLP6PNSjNKxKMwyFoRLTDeFOCJp50vkqn8I1sYkw+mq
edtNT+5Rha8k7AaE/LCHyYsgKXUUlnOREgi32p2oPuIHD7i0J9PI2xyTRc8+VaTI
/+PYLPvbZCo8CZbJQxdYeIGDzJuUjNJ8xgCqcjRvlsYYCPelRjnjgPkaAUe8tXjC
Do4+NoSClAQoIzw1dik6PgJAuZzzkibP5KbFHn6i/tR6nKFTghi4cfosGOFtQwKV
X7AaZL4WsK2pWhh+UrtusedgFK35PMyyK1tqjz71a1Ee6MUMDqPz29nSGqu5S1Wa
S0JJTA+hfeS3shs+BIf7jO7UFmX3JV4ABNn5zT6TB8133zfLyMKRkiYNtCT2C4LA
P1QKk6IZk0ImlZeeOx/vCud7BQv4S0HO8SRZnebU/9OUkmssgGa+yHg6uI1qTTYO
cRpKj93VwKt8fwqVNQ0QzUvKrDJVWRLfZIfFOzF6mz4u6NdSUZMljLODb6dK2Us7
5GNNfuViVqY9dGYMjywVBvwilsewHKSQjCoMgoNwhBE9qeA9YhnVNOKZZQZxCo+y
igKvm/NY/URHb/93NORoQUdblSoC/9tBQGIiW4pFq6sfzgMe4P9xXw4kp4o17kkb
AG4wEgKTbvHN6rD9dQpl9u0a1zQcLKG6aAv1dk8hPkWZVfdmRiwFNKoOthtFFxcy
obgDwwLPLVFICC1yLOO4NLWC4cXz02NWgEqseVQPpuZqA+xQkJNWfWU8qxjaQAgX
dHnSolu47dLPCWgKs3VmK5CAltIiMZEXQ3eIJoit3uitcyI6qo26DDtfZlItENT4
PwnUOC7AVd+H1/RFXSdC0Jhsf00yERMgH2LJGyXAcVMAxrZEYMsb6jStijO8SLl8
J+fRIfhQq53tdj+WwZS4Qj276t/RZTmTtAjtBm5ONKJ/0tt2wVoTxUAxjEwE1efx
oz6rMr6iUcnkKD7vn31xdv9hl/tjuR/VDHRgLHG7XDc2mVTEgeIOTNrtM7RJiyK7
/6RZRnbglQtPS5TVKlnGlp+mQM7/baOiEAXmKPO9DgvF73siSuW/hQukWAcNX9p1
9H7Vtw1p3Hz4LRi3ytC9b0+5Qn11nbORvEnxeOiGAcR8U/jNx3JBZvyKNnNI9/fs
jMdIUKs0M+aMWJ/fkwCo18hTV86EWySrVF9JLFyot4tEQEDCnRh01WVdmaxNOx5z
Tk1b4ssNBqt3VcFBLoDNcsc1T/j7iXrRmQt2DWWH40G1rC/zls8zI8Itzm5jo/4o
68buKa3g6Bx9adK+IMs1CKvqW5ZYt1diHBTesmf5xCdGqEiQBZt+dAdRRQ5CYUAb
nIs7TKKsh0h+FfWmNCyRQydfXaNGDnLiKrHDFLqa2v8xUR2xbbCDIfS1p57X/y4C
V7NpQollJNBQQGHG1d0cwoEe7j2oOWlUMhotxmTbP7veHZiQlQFmkwDxhWzqTskQ
Se29ZM9GwmNYN4WTEU4dKJ+5LYOrOVrU85zJEbIosJN7vu5xKpAuIac5bOUHqHhq
c5zzIlqedExXpxAnVCgW/Lg5KxS34wnhSkVB176oYR80NrL6Gff6NzkkFhZP3gb4
A3gMWh/KmEG31CvKNkCG9YkIBhpA57w6V9YLgzRduLTvQjOi44vxqoj09ZoMnESy
rWsOxS7KWEuy6IOvU+3jcBN6DdG1/qCk1fO7qofybtqtLATSOz03x3BZwCcsBNNO
PSkw2NAPIbyuP7fR5uCFvBQDLyNQbGJ/s1Xty2W15b0rEk6qUau8J2AdcqYtPlVk
+7Fv638vG07w5ymVpLqvjcnP1Pdk+/n4NGblLFE6TpsDyVt3sbUz2exZ5aATre6g
tDIBsLTZUWIdr9FDLBetFTj+2GDoNJtZ3+R/hBKIz2xnZMYwrVsmeK4duLB+EUhG
3Z89NRFMOWxsG7Lvg125JrZLOnylfYENrhIyZap6YlO2DYbqBXvU3ng4RTeWJn/A
JjIt5PLVqRravC02nI5KnjHP5t0ihpKzvxMuS62vJY9GmRU0ZtVbL4Hpu6ymWBrY
wJX/4l0dVZEOIryZz7wfb43m13VLS0JKF5QtBm8QfRAw9zck4LVjdsz7CBWRPf3m
227YQGSybXIFts2w8UhQhEncl5R26L4qgLlGGzBiEjB9RWtGMtE4SGTJMcYRaPiK
EQmUytGnLnhBnjum7C28C+cG9ANjWKOTLqdeLw8e70sJtlcmQi32HdxRgNlIIkDR
ZdpWdnNFtrRciRiVuYv1UVPTCIN+HxB6NSjNc7OUKOuW87tW9u4cgvdr60kzroTH
gIqNN9GVI51UJNWyLIkcKBG3aA3Sm87TEou8IrkqhBvOXghjCodC5xIZx1w5Zj71
A7rtdRROJ+eDyKlhsrQDgPnocPyG6JCqmeAzmBUrWPoygb9FBgYBNvJAo9fhMPkl
kuei2moaNgtWLExdmzFjTUR6OqDCHARHrFIKRn4vWJDTgM4bst9X6zZB0uBA7Hj4
I2ECd785c30h28ntnsU9Q73SMI7kT3wY7a+aQS8Q2KMTum/mNPWuuGfeL8xkXJKH
RncQ0f2piv+27OB+rnFlZZ7VEuzPNe9tRK8WVyeZsBHczHU5vOBAYynIeqMgtl6O
k4xXIoqwFX4/HTeWgm/9GWxbVNGJU+5yWLuwmDwOi9pw1ghcnMlIEDUdJXpUYOav
BoonFWj08JyTUFLsjsiUn6p8Iu0jqEOwhGhE86AxtHyARypQtOmX4THvTenBJTKo
1y7CtZLv+METLRvvIPWFLU08s+1loU5+MtWDW2SnaVMx/6FFHL84IIRMWlgcpQ++
LviT4d+e79nhUP1ahbXs/RzgVzNbRFZVQbDJXmnzFOoLmIrHq3/j4p2/qXG5XIi2
XbcDBx3wgFBPkp9o3O7gkh+4EF/BayWpAw/pJmFi0BjjXjdSokrIe9Q/ceA+CaXm
VtOL6qoKjgtJvehrHzTJyPlD+yP5awjHMjfDNPBf4bAOp9g9j/UWxu6H1oRRq7nW
q2+eajt8b3rQ23+Xk53+eUuniuYkUdhVdtqwVe+L7EBE03Cv71mQLy8H/9R1Xwx0
A5CxTgqXlI/oUedPTwPZ6SVesXDr25WxdfnLysrfTMda57ND4Bwfwn2EE2b98fnT
EouvdESVDNzDoGulJjXbBuBwiwd72M7TNPRR8l+idoXHZpi4zY7P2u0DQc/vM0j5
+VyCcyRGTf7DZEe1FBd3RLIOip2K4DG1d5CrC8Jepg81pVsgHqFZ3qfi2weyn4N0
JnwbTCchDyMBU5AqsC+vM/Lt6xO9rKEqxUAjm4zQsapMDG8ThBCu+Ziw0JpokmbC
GM5eDBJ8ubOY4qccn3lG9xGr/YztVMoJ481zUQUcs8h38tJwaB0SUupOXapU+Q87
wCq+LBDkCa9rWLw41MGi0gJeKW5YxPc7/HTMr4GjdW6Hxs1Y8IvM5PBLnYCKuZHT
kv96S+VEHeAfMZ1URJntcZKpyUxkEGl50K9ptKEsK9bbOlRH/6wJ5Cm8vHwXNVTe
HHeFk0mw4PmdrqjdDnr11wRXLFckI/adN+4HdpU/PO3p715A8guo97BGJre2d6Wd
8jdIFU7gvt9reiNSjYgDmnSC3p4S4nQcFge6KEmPxWuTNaQ2G//Ni/J7xltVpzxu
0Cps21OSP5zJNd7Z0uqUCC1hjlt3kiMcx/6rvSmiZB1e95JYMylS+OgZlU7nys1n
YaMorraeNX4ZaTLs0r+z1acQER7RfYr2CQ25LqhHiNjL8ZpDHxVSYUjz+vdBFXr+
tFzMWElBe/dG/UTZH5GfZ6I/Z6oD3dQzRPgomXUTNolVQu2LcCSKAfk8thF09Dcp
kFysvG4SxY0z999pJaEwtRZl7ZutB20YGw3BD/jhYkqKgTxQGDvAgXXmslGTrvzV
4hNKvt2CIPbcI4BedGUT6mlbEcEuvAz7+vupV4xupcIPUfHq9AhG9Kisnnv0nMdZ
U2QgviQo0voOaSfF0j0O1LqQx34HQGUCkuXEwlnUpCn/FO8z4MYKBBBjNPQUlFgb
8vyhpfyX7k6hr+o6viXJOWw6EPdxVnO61UlFZcKxd193R6wvrG8pRgRqv2NK1Juc
ZMUzjsGoJe0tf+yua5yzJ8icPRdt48x/7oQeHPGHgw8I05BWyfQ+W4vdFBUkwG3O
bdfS3OTqNzcG0CXYMQaV/GCwCrjNfvqlyebjSJbGl1bBRwyzyFPMr6Ifht44get4
WOwW/ANenH0DfvBsjrmidCus1+gn1aSUmxys5coOwXGylaUZVLVtiuzG2CrDUChv
Q/u45gYkyaQA7RMmkNRD59Ey6e417o3PfalORE1DUI1RLZjr/j5QZwXU3O6cQIo/
Zh/UyKjK5vTI5FVpMSnL6AkvmGyi8GLKQj9vwNTFTGTA0EoFzj+/WIAcbsc6PsaX
EJ1J3c8MPr2oammaH1Ok7LRTnM2BF15MQuQ6eBDPlwomvHXHbalNXpLtyxIAWqrR
Oqw62dI5qInDdxeE+7kKx0sCQUMIxGeF39wAv9lxeCoX1krfsavv9HSgWdF009tN
yqizFGSMbfBQi8VJe0bebKAh68Im9W1qCVwOU90j1g0HskUsnRMH273w4WMiB7OH
TqVQtG+PmlCq3S2Jr1GQYieqnbix9jwx+govaRtg8HaSoJweHCRUxV6KEV7cP2gL
sa4tNRlXFbdS4IlQF/+vGgh7RkkhZBhehrlLb0f1CKmk1OJvMktWIcKmQj2rUW0y
t6vs1DAwP33mMp7w42YNeDzpXoBbWU/FBX+igRaN+6yG6RwqE/ElofYSN/Esq3EE
CNLFoJE4sASTiDsxFAKn+CTd6NflLJ9JMu6yY1+BgxDPkENLyf+w+FbHP9NQK+HB
Emtl+T4ujQ7OdOHByu1uXkQdUWfTIbQv7bvR0SMASb4YRVa6RyP+xMpLn0zfgEJw
bbsyVgvfh049wtmvfnvfcBounFDNyZ5+TO1Kb6M5C88bRqz5E6DzjO/pZTLwk2Zs
FCiOCw2miH12I/z4+k2Bu3amfpHwuXa17bCbcyUwCIKd2js7iizGU7WrUEHlU1Fq
0Dyo6ifvLgGujNOqMmgJRHqej1oUMb03Wqm+04PGmqyCwuHCOpu8kEtLvG2/MtSW
lFs9gZJNykY7fP8l0oVJKnj463SFrchvCnnBi6Y8vJukyNGFxxMKr1KrvIj/C9Wq
A2vx/QH7otIpk4b7hHTBxTjmJ+UCswyhWnE2ouIDriiGEazv8+wHS6Q4CzYKlHDD
bvVugZuLl04CQd+QmJLGH1AuMAgUfQzy5GQnSWTxG87Y2a20WpBk9RUekU6erSrE
87BkS0I4ctMfN2LsauWjgRWb3Fl8c/2DDgzMp/1f9pRm/qd1f3HPLIGAvyRfBNfa
zTzCCOXd7fnwKq8rQR57oLz+WER8S5M0PKt0jI7yr8Jh2xrKhPy8KuIewk//fSfN
TC+bnxbC9OwtyHP5G/EckASOm6zsOEroz+MVJSZ49ahUBV7lvQPCiXWvpMyIJobQ
P4NG/tYrR8sAA5agYhxC8df8+RM4pKoWy4Sns68BMWqUAO471diiFE0D+TuOL1tm
/YGyyOLNBFdp9YlMuHo6FEuv1YDwl1fCLW9exMxAI/vuu3gHtV2Gd9d5OzAMYggq
RZ4+0yb3CQMi1ftkcR3Q/uqHHXTF2YIqON8SAHhvLO2YxC7TKAZg9tufhcnJESqD
zAyEGWn+HIEXTxktj02b3saTXyCywb0HoVtAl7tzZHKzrsDy8RepRO+l3q2nJoTd
9I58/WuAqQylXaRcZPrR5LSyqE2eRDmomZFp7v/QWLPRkl7rDgj0DZOxT6AGSkeQ
OlbaxvAsCMa3MTqkM7F4RTR4oq0no0RXMykfF1BBieD24eX7TXzEtALluOZVu7rK
FMMWDC4/lLQSLOdJh0AQ/AYqWpAW08N4s0UPIVvHDYAXbhrNKZymkK5ZhsvgNOY0
+1cAuhhjjIjXwhq9qp82XBDBkq3c8dik/eFvgwQ1X/czkzUwlLvXA9Z8ZUkwqGAW
CCysSvJtLdupxP6Bx90T+ol3Bip6H0q+3jLXLA7TeNTfjGxOtFrz1xrY4ILqH4rf
fhcsVTJR69vaMW6ioDFOMqbavt4ORftAroNjEepwkqL0BGAbTgxJClYdAXQZjjnu
cM6ddqNAGzC515O3fPM+ElqnkXKED1vvDel8JRTCzzmoK7F3yGROtq1sMEO4zuuy
x2vZ0yT0oFgfaYeg7lJfVAU5/iNMJaj6uyc9Ni5ccdgppTJNVhIPMAs2Mh59wuj9
25dzg+0sG/jbcUzpuCTFA26KwtkaTl2htiqWbJyq8l0titmcX02x4Q80DuyoYNII
w+RauBxoRES+cAxWrKzRg4VvF8pG2qedDa33EvfPomi6/2LuLp48rc14LbTPP4YS
h2PLpNI+H2KFwa3S/Cr6uB/lhAv0tMk9CZhr/KiPxfqaQHtUnYeHfuX83FCULHbH
emdplLGxHzT/YdzWU5g1Xi4xLliJFwAC7My1vUEJ4vn8Ce0uY/ddcmISRKrFH90e
pKgcxha6nRIsMiD5k4jjOBe3Q3oRpCx0d1rWVGpbW/H8qB5dwus2JAwdlAuNVcf2
P2fZ+xFb2fM9HH9pkkY2YEmEzrHe4scBhYCXkJYo1ZUfRBoMuxZENLhrQ/6HMrng
mkkc8TKgfo7F3QypYNEZOZdkqR5tG3wu4TgtVx0t1DI64/ZKbo7CQcbYMJL20JBk
YtMHlg+iFHro4WpMuJ2d5LGJ6RfsNOEUJ8+03DYy8A4GjOmB1djMzERsLVI5QN7S
jVOwDRzpwd2RnZECysyjYq3CryA/g7OHjdhJMKTo2X/azcNjp+VVHNW73ftutXaa
yOu5oe5S7iG7ObW14e+2c/GUqxyzoXWPOqKgMQDTfP1Q3x+Efa3CUlJ01cNZ4Vs4
O9AEgTGAS7jlE2EuFI8JDRD9kTxr9Nf2FEtVSt04ySv7OZTVeE4DgYryVqUvwduC
24hxxjjJFw3EqEdJOCs6dj+V2kVTAI08AB6etGfDLs/REGUnhPQKcWJ62xXTo3k3
fNlEqgNi5I21AzGrGlMdAuTaPVlBkohCNIGOw2/YpLSFd+JiC9SogMTm9/D3ZcCy
dyBBmAvHpYO33kIA52q4sXFBJ0r0OiVLm7OHGzwGlKVMnYVamNs7y2GmRSwsx3st
kr34Xa6PiJOMUuqAo0dKOtodCRyyzfmgHy9a2EyElXxdV/5P65LFMUPwscFgUwgH
yPlAGtv0Z9FP36iBA6dOrrCbC7nVoU3iqGv//1RTOmy8IkoRJNIX/dzdmB7xBRez
cFp2FampjZgdvWQTIX4TQuA1H2CI8pMTOD2bTzYR2UYrYqfnzjztw8siQnu1mjFQ
W/ZNyUJRkh9ObrhxEkbTrFLQWbX5kLfY4HfXwa9GYYf5M6NWSJxASy6K9BySR1mM
SwrlUkxMJaxSeI8CaxNGsOlyuOmV6g9p3HFAI9KriAUjXHu9OMdtYI8ODPph53Il
d6YhMBanN6JYbpOJdnAOinO2QHkZ4NPQPDlFDyN6igiRxy3wMzMlWgavs4+MUOdq
zUmndnfGMEH5OWnkHrdS+Upkm9SamuBtouVX1C3BUAHmbTGYi42FN5I7uf09vbnR
mTL1g+ry+GkGvyFdmXZPFGcyu6kTS1SebNCKWHoOZUBd8PBZQXQ3QSlVKy6LgiTs
MmML6CKY5szLWXUQJ3jPctnma5gvn8JPFEkDqE2V1B50Vuvlbqimg36n65iJUf6n
W9pw6B030M4KnurvY/qtOqnVce78Q6KRGTnAvuCgu+ySbYuJKScHQpcPBtTLuF0h
UdyRhARDkyxKwO33JcY/j7kD9NmiijvIosjtu8aXFqzv5BogDc0gVisZ8iZnoMe3
8sgIjISQkt6yzCRFp58SyBCa3KkE1/ThYU5DSuPwUJClaAm2yOGV67+f6QZhUDsz
dqCcHKpsWxajI/Ql7TQs82taeYSvZvPTyyQtacyymgFqtLTuw7iUpCApOIaeUk4a
lBLcS983RGxIp1Pc4rDH0WCb42IfEBa9h0XGCbVhq3D6nV5nCWbhUvzLhUCDE65K
yZufTHpEtdJh8opTg48L8Y3QaR4AgWrWsjNo/PNO4b/xiNnoq0LezDtw9WCFATWM
QqNCqpAJ8z+mfqAo0CgZ2fMviOUHg3mGFHjtrM55WWGOdKiwJf0jgjqvbK8Y+amG
u9F6c8DrwaQOTaEr0UnqR5OMoi6RdKjyee2Pg/14dN/bhsinnEE5JnfBla6CEMbf
Ota9pRje1HD4FkJvq2egNFPihdX1tJ6xciaEPdQmJDYKFW5yMq6q9sR3IDbts0B0
nZ/YMWsSZ2ea5P52K1dIK6BJoqOiicRdT7PhZzeHlQLF3wo+DUHAIMq3egOMaGPe
CGPujQ+ezkFgPzhccN+jVVOuDmQ8Y5AsKspk4132kRW14fyWLsP1CIhqtxb1N4ok
hpMjTc36tsSVIbIlkLBDYKSA6jN6MNJ/tTPQbRyYlELWKtV0S8wP0Ei7UBWVEyLU
90pQXgnlztaxJm3P63Ey/NlMDIctSicAeprkFZhQIvNwK9ice0p3y//zRm/wuMui
Yhh9nHI+IitbaTUPmIdY5RsKcXvNX+cETxWd/uXcqw8egYQdDJXuSOkN8YAX2jQV
wP/Q3zlUeIDvN9LmdDxvnCYdn27cSKjmb8XQGHM+gv99Vo6j3pO3tIAC+XtSY2aF
ympaxgYyPoGx41Oi3t1URf6lMm9U2Bbin89de+UCoSpGP3pSfQYTUT/XSwDqAVnb
0YROOYt//D9dleeipmai5bNO1xbELCWw+8eSx9GOvRKvNKn9C17rl24VkMlUn3zG
4vEOjEP51dZcF8nXNY+UGjrJjOy8+j/qC4mT7z1WJFuQ2VQ3Pg/0CZYYTyqsHb+e
by0EVsAeCIdMM8cZaoiOcgGyCFhpTX791m33eaPkKl7bP6IC1s6fSdZLZDzax2Jw
2tyGDniiP17O7RxIvnhy/KDJ4Tr2nFx/FG+m2DW+kfu9sF8Jaf0AmoXW3Ji1VzaV
tFWU6kQomL3X7+/2sp2aqGuQnOc8fxoKqwjIoVSvln3rCYoZ5xGsS9J6IXiBYpsk
59YcAqTVyLQmQ8vKUM/9YBOQrG8MITeSCgoIht+jAiQo1UDMJrsVcJXiMw+oZb8B
kPFcA/FTlv7GVa2cPD0thAJjgkEpyXUNk/QfsoDe/7OfB4+xBf7XQP38dxF5Q9Tw
O/ZUNQ7hW5TEUV4UQtV85mIqrA08fMHXzXmqA2Cmza01Yd4NktvydpP9FjpJMTAl
zYdmGQWtc65jlHSNPGlxGjOpAHw3hP67S7g/rzhGll020PPLPgoHEOHcOiN2vwN5
opPCUsNztZPhUDcWY1psNk5EzUr6PUQZqIo7RZciqDDpOCbtxlC22VZ4lr7BSe3S
wqs0h6ZjxuV9F/RQfqrMlBfOsdotnIYEdcqvf1oMNVvhMPyQhogPMDam6ZtkFi/L
eB9NQeuSQ6fYyXUQ1NdEl8YZHLsWAP/XgORgRl7FuA6AO59CnK4mQcbCSVWu/U9M
k2J8b+BuZlhN8B5JrgpaObN6OtG81PcKOL20sFAUW6F5Hhah6WJkL9UsouSAixnC
Dk+jcddg6QB7g5+4rwjuWudo/k5JotB9D5QPTx4CkkeNC36KzvUElRgkWV8tSHYp
PfEoab+tvoo5eiLtph55lyNbeYvYXVP6lJdz/Xyk5gWS7W3KUc40eMxrRv+4Cys1
l+1Ep5sTIHlS4QMLsDzVuqyojeglOk485Tun4JDW7L0X8nasz2tyFS2caPTYtv1/
IC7YerhX+Kjs8vDii4E9Ayd8XgPrr5LKu2FulHVJxjTiPaDAkKbT7jxZ0/xhkvdV
eNYIzUo+zPpMkrLzResew1htp3vBUK9Es6Bu2Mti9SiV+axtX75ucojGacuM1N47
Al9Xx6nGH2I+CMM3WUPwqKZ9FrKWFJtuIWrV9x6MpuPumUpnTvc9Vdr8ScldmHjg
hgNZ8mgF+YOeiSKLcEjjrO/kdpWdGsuuTcD5sxQJv4SEKkutlzM66BoAWPZoAD2i
D538gHOILaTkFJZf1zkuXAZphhIUdXbzFRUpU0tQdk7Rt4xYP8qqsuOE7zx806/i
xxGxGgzInCS3nt6PHAWeUv0T6eQW0Jj/rd02O5sm2zphadpTHFwI7sZ0KSu08WGo
3Oacb+lK0/V6LlSJ63+QSxv0JijdRgYHZUKo9wdiOK60qQU/MW0pZHl5WaYcl0EE
2m4aHVzshObepMvA78Np+7VzPSA41b7MvmpCUA/29hvzp/pe3unGUybjgyZ/skjt
x2Ogv1JQOQgei78vO6psEY64sEjDO3oHVo7mxfEDYhh27d+wuq0yYes9MmKbfe/d
5aD5v11heoHU85nGLpXI9nb0OGRwsvrk1lZCuEHpHsPGhrwNlu0AQHMJaDBxDyuH
WarmAJh6+HnvvxNJ881fPQJCGXzIx+XFNoIXqrt7xgJeUWjYXGU1ja9cK5topmWv
75LBggq3NYEkqqGleT1qLqx0r/CAMhq1kzS3onwKp5lbrakhu+dd1puMNVCj/CkT
rjjJj2OJrLGuS4YeOYrPCjt9HnZdLNm0WCt/dXVJeWms3DZpWCvTEJiEKgPJMHgY
7nBjKqIsRiuN9Wi7dGz6Zr4U1AGBaM1ncGB4/pN9Yj6wlBgw4h09BHyVWtrixSat
qaAQZ8ITmyhRQTlmKjlcvSIBCMBP9F/MfQPwMFmBWfGzNiluDpPVURNkojntGaXD
l90tTNAlaYnVhpAtoxOmXdFRgx6ik0HeroSW8s1+bw9ZU8PMWROR9FoTXmlVIYCO
PHU/11KTq6pl2vSEmWxB2Xv+wS8wxJ+3BtSt/0odqHjrh2MFpeE4Osl1qu1+9C1B
upShd/CZckPA9HHCebJV+5k3lpWqasJJCqfUhocynT3Q6sWwSiuOyJy7W001fiPF
c/5G+4TzHOcnCBtPg2X6mziiJPKD7RQhyTn7K/XKq3DZ4OKiSYsZBcgQALiDa8VK
+CVaNqZsKZ3nKFuZ9upUK1Bq36GfblarD2h/mSzSpE87l+uR4OlpLD/bxkSFnqQd
ekxorngINmk2LpDAyakfb+8/4oLgRn9kCAhsk+vDZY6x0RXtJFpIDQ6tB4dY6qTN
dIpFXZcV8L3TMRwlcZSsodWxwoQxnLoM7IUAoORlxwgSgy43Q64xWMOZa/2R4LNM
ULs87V1m9vWFOpxZwWGpjN3M3Ut6D6MPhUZomTER04rX7JkX0HFKeIdTS52WXBU/
iCq2UhBWgIEKaeJmIzIySxJWSV60L0VQwHXMqO8mmxq4J6BiL6bkQryX087RThMO
H4joSwu1IGSjxqN4NChc4oWvmX2tnpn5eAwmUZPKWCuwuxjGs0BeL9GEVMd7vHQa
nOdMTSW0dQli5XXa7SYK8A06foGVbnktaTbyidURpvXJEzf5jHm1Kgwono3HJSOQ
fgEet4b/PygjJU5ek5M2xkAtQe+nfw8DG9xTBbJ2zAfsphUNjU8zHM8gdJT/0j3g
VdXg9/i2nZZGB4DGrStvRSSK9EYFzWlnfvKvLTEtY5bVmWB5wQ/Ngd9IREYa3pxx
bn9r/aZTxvicNv3S/pphLVvgdavuEWcsmYKhCnBNsD4D2tvePLRBPUWLmd5YEvEX
QWggGy+ZjcZvPEgzoUFnD/oRfAmUuJsfZPVX5gWsOkIcZitV8br5baCb277hr2fS
qmiGjJ3YfdesCPqSh3uUWqLjE78JP2RA0rwqmJ9fDozqg9O6Uc/RPN1M9A66RGER
MXqiOPygArPJK2mkQEbg/Tr/0MYpPC7VZQPU7ruaaUWtmrNEB/q8GwzXP0AMXuaU
B1Q5a0fQbx8/UoEIlOyMtP+Rwk3/GU7stiTPHlsM9ApoIefVp2U4BV+JQSA/TwNV
lXkfRdiseSLaCQXnoNBLOCyeMxGVepGcXdZfMmtLW2M0OYHdOvot5HtbAVlY23JA
zpGQB/DQMSZBluICsiSgW7pOQB1HoceTmnVS4pWO9yUjZjeEMo89HwQMoyBhCt6O
+3Pqg1n9SozXxf7cR/qNvNHlTacLi0NKosQLeDikZfrg1ks4iaL6FgPbwYrNUh6l
YPp6aNBIJMiP/9cw92m+4uwbbeA1nuf1K461NwhZgFJaTM1vU4UE/K6lI4UwvDcK
vWrzdeXQWMcx6vDk/93kjQgB5nw/TZOev+QlDCwCTPO8eFbmfRs9ZAO4hzf0TsMx
v0SSZhWcBXVVWVbiiuqQK4cMNhyPSzqK3PcmZMt7NXNaWWQUWq6dzrVZZsl5Jsex
LotktnF2HpDZiqArwoELqGRK/RmK3FcA9XvNjjwVdxSEPn1BcXb65h/j33EResxw
FAHbsVbOVsu+M8WgaRXxpiiZ0Jc332iCtovOxvxBCK4cifd7KbfFf5X3EOvFPa02
tbhD6WpMik6R3HoYXLNQ+GbPED3yTeqx3THTYT6K1IHYDmQic21dIYC1TauCWUrz
aXFxJUlpyXFnKsKg+HURn66iklGyUyeMGK5SunTyVxNs2zjweiBU90dH5t3SjbpS
WtUC4HPiFfoxoLVWlC04ZdFjsapyW/yjpJzMWzwhbYHo9ea2JLQTf0z4UfARU7uq
KhHkxx4URBbtedH3bkZVH1Wgwc+3GncBPUcDaoYwOmFTCmRNTyaXhd4uGY7vBkjc
QE42FTjs+/dT+f14iy1H4sV4BQnueL4p6S8fGzjqqVoPfnq1CdohekB5YyvzXU4Z
LC5kv91SE7RWLYBm2eUfe6uNf3P8Dr6kfdBvtTywK9kaLGwxvwCUq+fpTiMe6Ull
eNXKaoE4hzW0j+wo48QgFhg9+DDqf15c4N+OBD7NOq2j3BJwYrgS5sT8y/JYYZ6h
6XN+WWrImUZBTnLG/S3zh4GZD2/6HmY2yA7brij6yIkXdNNTirAAENNWUkw4X3jg
3YS5d7xPn0RHd8gpBevbZjDIZIJcmvjgyAHMB3Mk1/sq2cgSENSt1eIc+Hke8AEC
hQO0pxQ66Fuiv8e6PaUH+OHllEH0/jtGBKOegHKZAHF0yNj7YGzLY6rpYAwYyUHE
AoUbH9dopzrjF81TjtHu3rZ4aYSVGODz3NbRXTV90BenIaG/KhUDGm7LRMlo2GxM
Sk+iRxtItpgzlrL9wQDdHZomp3hJ8sKba6dZ2oiFc3zRdTglYedX87Hz7MPX/an9
ysqrgO99GzqpFLZfZSUFSQdX4LEFeKv964ngnqgtTuIwuXIADscSmNGk9yErEfNX
Uw4GqqFfOeqWQCBsesBo8Ul1L3dgTyIr2yPMO4cPsPA3JVnxC+Ca9eAlbZol97f5
k04J47KFnKEf9pCZG5irmjuyBTa7XzY6EdlDwtB91vNFBh9C/29ubYWcPMYgZCdk
cVmECIiGd2NiSSkvbkM15tICIy1KJlMRHOdGst3VIvJGVBupHcEYE4Jm0/jGVbpv
ohPUs4YtGqiM12aDexjCpXVogPDVa5NZChhUKsaj/JH9mh0ElJN0AW6LCI579hKo
Q2dp/C3HIFiGNWEJuBJ5Gv9ch7HzgFFbqCztcmoGwBtWQze4fhIBPONI4kPz1Qlw
OtqpkzuT597VG9Jbo311hLexSying9CBjVpMGh6PQtaQFI/vRllIbuE1EIf0KGpG
WKubYadyXtQFXjhS1FBw/Kq8b4L56uY9YSM8g9MOBiC8OHjh3efeBWbj+KGZOtbd
K1FjhrIXM7sP+mxDW80CjvNpyLqb87NrC29gfeVyJCrBYZO0SsjINXYEHqesCHvZ
4Yl+BV+LSiYvxKIZOzX3oiKhEIN+NVgyRjhGBJvnMnapATVgJvA5U7pdWj51YDLL
V38YMTY45eqXOh2EKt8VhzCDFk/nclQL32GekLONVBe2SdkjMHh+VQ9+38Hpyt+S
L6lk4HNgN7KjqmpMI1OWqEfJ5DVrYYagehknVnJFFVZlVpgjc8jqxXLr8h897xQo
bTzvnXN0i1ZrSnP5qHlb7Brebk+pd02MKUKNOtF/cl8+uRUDxiQOE2eFUk7RrfD1
TXSF2KGCIOFZk2nOz714gogKgnwumyJtD92qwURy50Qt2RRBdhOi+IFWAPmQoYaF
P/XFoaEGf43pmirN5BelD8yNmIhEG84qqad5i8tLg6VJp2ArlfFT38zaIs/cndIW
tFjQfHPhi7scyIcdacaPc3LLcLNSlqg75re/d/14SjRHKII5cp711QkfVYjhkywF
iVJeVzRj1fIhn0R3URtJnytnR33ZzYxuebqt2cF56l5ZHAxXQkvBBYC+UYzVFBb3
FreCgrDJxlHRwdhKgKBCeIltqePikar5PinO4BAEnFG8rFrxUUhx5uG+BDE4ZVtw
Qxfz/Vuz6fu4wXMtqAMCh0NOrDYWmN+BvSfaUDdB4Lo4rPyK4XWDEYEc7U+FzGse
rfIQF2DPnAXU1Qx567kbnE/pUE/xgfKplVdIhHMqO/aeeBCoacOoAzwq13sRXpx1
aHRrgg4AeuEIgfhG0hWu277FZXQc6JLPVMrMgtHQgCkwWNbLUoy/1c7d5sArkAfx
3S0Po2MtLfQOOyv7cNjpib+TsHHZbZV15EAEn0/ltIO2yE6sfbBvz68eFPsVg0Fj
iOJxUfpfYU1aZnckMAVL/9nuQvFpKjycQfsl1eFDXFUh34+F3Zunbz8q+f1iA+iz
VZfKcEhdCbkOX0npD0C7cbRKgBFF31NmRpV9A/1tRDFcxSgEf3058nTxmZXFbqRn
JwymjqbqlbWiRthaNtBRP4FoG6HcdAZuGrIxvqWR7L9FIMYDBmG4qq/jQ9xNhE9e
lh+YsFGazdr8qbNj+8Ca8fOLAMyrZbxJD0xVAWvlaq0ESzZUQXTrnNqb8gMqR+p7
Oc/725PgT3wmU6IIjONIYtp82errnluw/Jomi4bLQBWxvOmbpG6oc/XWS1SjL9AP
M0Q6AemIc3BZGcefeW66N5XDwXai2qB8kFlsriQPz9czNWO55EvSgVPC9gT4tQp+
JeO8SH3IwTiBMv6N/SRMcjECWTumO1b24rBThvExyZZRfXc6X42wG4DcqKieXsg0
UQHgee8t0jx4uL84Pf1RvzA0ZQJ4Yk0EqiGEsHQLJcDIzr+JaW/IxvlVwqHIAMg3
FZBuR96rF8kKdWmiHEyFYwlRKTLaEN1ouNsmfASNA9RI2MlQ8GTswGE3KNc/YS08
m1v6/wLyYa99mdeDdLtTOpfTAAfkRotsksRb1Fp2QOMefujOJ9CroHsaTfnoSYD4
7YoUNi/j+MTIZB53LP42+MQNvAqN8QbmCEBAu+//HlpGMfYbJZQTatWC+lD2ryOS
/WlfY7BoXTBoDWODg9K0CembPoGjl96OEArTl3l8DdxnMw3bmqiy+pZENdufqxeV
0GMoD/KctJoSe1HxZI/ILyouzef0/nMkCBzeLuEwf/etX4j7Oet71u4jxiT2iekT
tX+zS7RvZ7vAyo0e8lRlcUTz7ddZibvm0uerCOwEF780BubjJd3yafJeHSO/K5GP
1Y6c94l22EGc2SLc0Efpqd4SaX596lDoZi4AyE+QxKRNTB67bDRqUut58NNFxyk0
wRaloya6AvFgQvUjWT3n0LIqdQF9YpjA4BcC5p2cD/KqS5VdanFhSog6ZHq84/gV
SOhcFmIutDnfL2jUbGSU1HBajEtI1XJ6FQhrNgEbYJrONXsKp5seInCoWmSFztIM
ZiZ32B2ySXrpe4ZADqZZQyL0ISxCJIq2RE+dQE6nzP6DYVmLuBrN5WBZ01g65bgK
w8c1kqJnyhQ/kOKNp1gAPMuCR5PQ2CvL82p6mZul6di7n/9bSmpwkiBVzy9fL1/j
UJnqqFaZWb4uTxp4vES5JlZOPcObONxxZseWaZi/v7Yfi8UZzjz/m+y5/ZA0x1mz
9wus4+VYkU7NW9DQGrVwMDrUnDpuPxmtjHatcyNEtiwSjIVrW83hgjl4Xb1P8wK/
w58aTMwjewLB9f3y7hu17Tt5G1bQE9oGQU+7WCMBGlETjXN3pdp0J7m6wEs7W9g1
ndYt7u2NbJxKyZSGxzk/l4lA3TKO0OWvXk7VEdCxd/LO9kImX9DBfwyBpQumqSB7
lQuSLCFMsp5arICSBUeRPaPfAbCZ6QijWgwblo2O7RqsSq64ru3/CpwXB3jREypk
G2f0KqE5VK+GSmUEX41u0DN8ncVWPvgqQn+WG15a4t+mR11sD+iPxf3dD5uMr6NZ
SgLde3bK3R8/Y+SIz4hY1TxOpiBk8l4BvK0rHFeRZ0I5R0TG3Kas83HQDfOOoejU
JKtjzGCGu4lptOetsXhTlnmm2VNG5z0NBqvw/A07v3sNNCzlemuqIFSdHDIhIBoD
FmDn3xwLD99eDchUHfIgs+pp9rtw7i+Hxl0tmCFOBc9GQl5s8Ui6oxltndEg7OA9
8aWpwlx8JY77LpRMfE+9PcZ2Nst8WgEV0sumoUrojd1Gf7ECut3Vr0aQQfafqcRL
SJSC4Dl715co8QO/TbG3ViZqK3pWZDgmewjVnlGrlbjBicQpvTsmWgN372EVITA/
oORf6DDHeRIkThLsSRbBnXy4Pfi+9vWDpxB3+8ylvtRS/V6UvWWzktPiUwofhQe2
Ia3elK2MCri/uvlhPt5Jw3Bsc6qno9DM2NMPaCO6dOWhvmwIi8Pet8rYk1cs7J88
XYkSMonKanLBIiXR2y2FzkG9owfXa6E3iCu0Wuayxlt1xdb9MVI8umSJpyKJ3k5o
J6YWg/czt71QaUpYrt5Y2k7WFfdK9H9jAG16SB20h2u5aoYhgXx7HhHXjbjQu9J8
bQ/EQpOo/CxbXTiH5Ea+hfGDAYrA2fs1fv338+OWRF31WzhX3EjMF6Pc3A4Gkjpi
1lIBLbqGabVZhe7AZFGoRRLoEH9v30pK/SPHtmuyKibdHmbs5pHgJ1GGfzDv+1DB
qBVPoGOEneL55EReV6ncFxrwMxn3VouU7tM04IYyB5xCy0qop0tGj5sJ+WTj+DQS
6uJcMltFWERvq7WPPrkW7zkkv7t+S2jLsJ7fIBTU3K/I9x68nfoPz1Urm46A3C4S
nUk+ml+wGzL9kWKV2h0we/qxLqO/z/pXIZ5hGyNXZUQNrvxFTRDI1a6EotCokLf4
mBi+TmguYbT0AM3Pz3W+S9FmGUuHrMeSaez6ooDmZ8IwlyhB5XyCcscUsRH7Yj+E
Fo86ojzNYLvYGgcCWG2m8uS87tqrahAORhi6DVPrKAm6aeMtLqJDQTR01Ehg4zWL
TwruHNZ4tOMNNsReAIXQr+TQZC9wE12mACW/W8E45mgwG8MfGVGnjRtwau/4oVFd
mYoZFyi9FrQKTUls3mUKynTmZ1I3fq5bn7HU92GjgCB7GstP15MdDQJmf5LaUa4e
+uhAlLbqWIrSyEBUcnwxQ59SYvhLRDHhK+NGbNgk/7IrA3S2hUnw9TweLu6abNhY
w0BhdPXXXZJ9tRLPkN0Wxw8moSKXo/DQNC4H/Uo1PFmWJanul1tI+BPgIZqCcflK
XVvTMlN7n4zWbztZoUn8nK6/rYCpevhQLds9DgTp1N9+C23IDQ4CgeGAb6j6ePi4
1P2fzr8i3AhcXTyrYbzRcoQ2+mXN2Md6Ato9ejP/ZFENVWGB8iTSpxVdOKB4Tb/9
6npSdNX4DY/a0l0M/vKeOky6L02m8ywlMPJJr5plwgMcw2VYSLi+cKwnMy65ZN7b
YtBStTcmPaV6g0SsQxK3YQX7+6xaxaFcglSbRICX9p6tUsMNrP1fHsl0Ii3txTkg
aS+41vO3yC5mtitqRJl9VECKfBS5MAWlsswAU281LwHYveMOYLEkuRRRMkZRwIll
OiYWtrv9bnD3Pp2kjN+kBoWAe5LYYwstwWbPN5nqCSMGAH30J6ac3Hx5x7oIBKPa
hXF6SFyeOtWrckkqwjF4v5SAHRTWuPRmRzi+7ojpslKSNpewsnIe9clfPflUcZOM
z3gJofiFnotvos0yyONFUhKq8oocMI5UweHAi9KXG5efYWiwvGZxkN39b8vH2VzG
BX5m7XAag1Pigv6DF3TnjrIQy1k3lTsecz83VAHerFu7JwHiAzclmvzxBZXl/U79
V/vF1vdsD3Ng/xmzONaYBs+0klBxBSi3NxWCER8fikHDYK1iBH3BRLcYQf/+sb0e
fL2ScoKaDgZYCsFZPO74PTohr0lIgp+wCNWDgK7ji8zu2oP4Hc42WUo4xUPMJSJ2
/kuWw/FXxDr8lI0GgKaLKLLIKcBlTlasqNQzkJsqsLS6nCD6OquCLx0csv3IxmDZ
PqaKvoLDsIGlpMlV9rJzx8Nol+rafWSWjWHwHCFSx6bge+vu2uq1MitPNcT+pBHv
iUPLRVYFiQ8cD+e7OnD2oviC+f7XT6YrlXQOEojTknqlfqXRUdtqMwmug6QuuEF/
kdqnOCl3dTd8Izt1RTylZr9fOCcQHXnU9HsRYznfOuQR0QInocjWhqnyug7ah8oF
Jp++Ar+mU9qJH8sx1e3HPQgmb+AGS2inbFhlUE2Fo7gQKtIBnT2UOzjUWsSyDX9e
9cXus7s8SvA+j3af7U6LEaszYJV2CjMshOBRVyQ1xr7Qi2miowO1bmld5IdAH8gU
9cY2fWWajFEuBmebV9ENqfyGA+tlZftxqeOedf7ihr/Cni0Qy5yx9WM49N19YjTe
Ei0AoOuYWbdM6PbjkBJKT67i5hrDz894yekz3Y4wanFF15O/BVDGrzg+iEGreCM/
R5JfNxn6StuT97foXYcxLid9Kz/e2pp2a09WFIlpte3bbPeml9YCkkJCTS4QHd0r
AQeVQrFv66EMhXh2vgkqrZuJIlzNZyj8Yj04PEgZec61GjbDYS6ZrPy6hRNpCFUa
xNJ6a5tu4EJLTE6EvETDoIuFNAAEfgg+7rO3BIGl4MM5aAzFyA4tAD98m4/huCzA
G8dbzKO7IMZzq3Ri5Ts7TzSJUOxxPlP7FesWA56uC+vrxXD+XM4py4D3izYCa2XM
BiVauDRQHcbITEvCNXrfDS9JNfL9suLbeWHpoZ5A0hODYSZ+Fmc7a/1tYhATdey+
kYW7CDIxLJ1MKDyQo5DN/1TmeqnEjH9y1BeWSuWGpwmRTVM/1nWUkbES45/r9VV4
booXWPHnDIxfJrE3LhlyC7G3JRcgymS0X+shM19lteTGbHpa9A9CvS/FiWyRoLAn
eewRYRaFo727cKHIuNtwG4GVF5YURQyV8Rgbif4/EfWnBP/oTm4b4nIkRTjNArUn
HqA83nkMBVYU/xjSqYtegYuTzvBTFQgmTE5H7flNE+iek1kF7+xCIP84YxSfwqHO
7Gtoi7ORA8sJm5H4b34oOMEbY61ETLw2VHgnTH1areENyJfp8RiuKuOucsmAfcLz
R6735JI0APvN9DUs7UzxgJezUZ6PuTxmrJzsQUCVizqP1T4sZzRNtzZzgHmHnodN
xRe58u+6m4FTZtnuhCPWX8BwJQrKyOlo4HM/QZtp+Sf/rE7q2WfDm+gd2xfWIvge
Q8N68Q5gS6Lk54gVeNpd5d8pHY/Y3uonMH90qYpZA+nnORTgZbtnsm6GxdVDzySW
XSB4wY5M7umxQYOAbiw0DGo/w0Q3yBWIgmNVXLNQj63TnYBbbbenSxvCXGY+eS/U
D0oA/uPxkG5ZLMr3IWO9jxHjMRcwTIeDc4ogGmDqNnGE61NEljBSfOleqVMzttRL
iclPWqqIl7XfsTOI6lJIjDGDcGpbALg+RfdOOX/8XgqAAbJGY8Lxx8Z5rbjXV5Ch
hTIrcVQ7ISUYtkAaKEFlK0C8k0rmH5IVSaQ01F9Ne2W/Ib9hBI6+gEWs4vt7AbCJ
4k5X+xfx9In3biPd1NHLwMNRPfERHszz/FKYzfElaLqzVKFMQP7du8bHd1x6Gf5C
T/tSEDRK13dejs6y4NMERA7NRFJL8fqOuYToLyqrgOatgKgdCjjjsxTy1x99y0Xu
OqyEoD44WYaYxROoMRlPENvDCR0yfnxEZokYffXLAgflSxoapgw/ugj/zWS5Z7Wy
6sc9yK+IuTBQb9Uxw8KWS1fuXbDcNj97XjtSt6TRlVmpq3JOQeYjZIo1ysNsJxo/
wbafhbmKaFkcv1QjfVzQk9CMtP0P/jEv8vw92O4xI4jXDI6Zm0Ub3RFTpAUtyGrI
BLQ4FgYSPPrj4ErMPLDjUFVrG0GF+q8CwBAEeKDdMSqe0otKKdL90boWqk9Qjzfs
AGm+9U4cmfgtBmZ82PevSeMqtZe5O4HbPl4jcrGkn0HTqzgKhtgVOuAk3vNpfsi+
0D2zSDHhKtzlt+gJqFCrYnoe1ReiI2iZt82inxCf3qmcaW6UAK5djC24cdZz/EuP
FhoRZr4M9joqMmJgH6bCKG5h9m191BikNfvOKhMCS45nbrJW4Ua1WnNnPmh8+FdY
3Wtv63U+1RiBDjTH6pMz6GbyQB4gC+8ofGbY7dy2su1w4fEJtDkpcSC7d0zvXOSX
P4KF1kKCYY3l+ngUn7jiAJ6uTWNKQN9AWE3Q02ffo7ZEYsgAkXBFyC7fWQWlzEfA
KLySBBuwSR/z+gETxtx8rkHeOUs8DRhYN7M6ZvKhDUtUCU0zo40NGDoTtuii/4+5
2sQXCV7fW4X868NCE3to9G/Vx5MrTLWaRTNNhSKfJf5CPN9Nu8i32OOU0gWxjTc8
JO5rhjhwXPgVlo3VEYJg9bGxyAnkt1fFgIv3yLI6pZXTomk0/Q4uBqAqKkNBDYOo
vQPvy3XqrOm/u6m6s6jXuLuaLZhOoz/FlaEDVd9lnJKc6oSVV/KhG50n2Aw2iMDA
w+MWDfIToI33c0Wq81GIPUTRbvEQpbdvbA1FSmSjbzeB/dzo0p/GNTX9aSJFox7W
wxhcAo0Oq1lS+/rK/o8TMZsNZENFtWHXQCaF8CuVeAm3RYCjvgFndDWKEsm8b18M
FTeaq2Y7on1V6z+9C1yeKRN1/8wX03LF1WzKMOezFasM4AjMK6E3eYADmMhZ+1Vx
tGywrOJfw0J49Olyb9IAPjX39BDUpJSM0YA+ognu025fek1JhymPYLljQCyCOXYu
f8xUpeci9hcBdfb32vAVT5cF/H+CuXdw+HMPjLAW2ql12OtlUWzcbA3vFuQtRnju
5QVjYRfCoOHhXVvJUi7Uo3g8OgjymxUkQ6MCdnbcusXCRxsTDpNAFS3y050vqF6h
AWMYtRpHQGzpH9XjC32B3f8VfQDslUt4llrXSBpwfl5tVK7ZPmylrkmwLArdJ3Oc
z8d0BohkiYkABmnTWmYBDKnPrYG8Tsrw8XkGN2NOFTs7oDwf3CcHjaFI9QwE30YC
J6C+U2/DTNTvb4CIuZ3EXCqOBIOUiLpgKTbkQTAL85NBAn8hP1HnruFAE/kWWesA
yXj5FyhRyYFlO5+B6M4P4z5XMwkeTtH+wcY09Rr3U9mjoHZ7rRY2GF3jIEn+GWdN
6GY4rdnW/ea0BEhy7DIFEYKPGLuFJR3syLwG38hWLJlCPeSSO5w6+HYLuslRpU16
pjm1rK49YMBAvFekKOj4lyLw+t4KAwZ8K+vauu+Q2mKw+vEvgaSxgofriyvasJFo
DAwz8SOe7AA9rSs8YLHaAQgIP1LmP+z0BfvXWKlz/6IbvT99t9f+2Z39crbintP5
+MEpr4f6ZJvQIN31a131vBGHhZG6p8TY8DWYmeDHM5M5ZYOwEuGNipbixDB7bVER
91iz/WNlgqBv0cRkja0u/7lC/jzMwfbqP0zvgqW8t1O7aI4rPcpeDLPA7azonpbA
T9gBt8c6eAgzvM/c2l1HXwkfL8ZEhE4zlUS2laHbS7vNe2p28cclPwEEcENTuYLc
REaL6Y5L2CKdxg2dr2+1Vrff1aZqy++2GQs8PCzHdwYptRWV9ycirA6CikfqCzfV
mKgpww6elG2ljoVn0tRIQp+uLW0NBFermR5glAGsbx8XKe0anvHEpkqvEsC3s5WE
wov6EhtAsLS7bNGYpE8pjulrXPH2sDd/S1zc0EW8xdxuP7j2yFkdCIrEI0UabgIK
UlDzvqlJpX25y9lO9mB8Ffo4/qj8Nsw/3KZwgNB5GlUyGnttqnuMXpqfMM1MzAn0
YpzvCAAH2XIEPt8FNFcLkbQuVmN2miJH9JcPDVJPWQLsBILpIO6HZTSO1fNoXhD0
se8yGDvkAnx6L/HE17Mnt+iU7gQp4DjfXxJFWS8W9wDewHXNPqyYC/7JKPmy9Tir
w0eGN5lrf/jgK/etqmIm7BUidu5TMGfN8w1fh1KJDe1NmvfdPxT3NCOCxrPViUyp
60zp40u4+EYjU/TCPyVTgzn86Pbr4wzuqDt+d3YZ8MY20AUCv7PBjM/3rV1eosmR
3laXT9XG+D5UVOP53HZ0ibn9IlbNqxJDtnzlRGdSfE7/l1+Qfy7+Uee7yo1tZzuH
Luf8BEIR5+XsQxA6cJ8cjYnFRUDM4wNpiTGvVs92/i1pQkA6pc6kUyQmn7jLORu7
RaZoOdeWz5p0OTCnDaA+jfpzHyw9o9e/bO/FLlfvFW8jpS1Rm35NX5B0pW6fX1U6
QJWDVLqZ/Brmmj4LpVCsJeoeB/pNEJ+gQCuTEeF2BtUAHaCH8N4WZmSaJ+/MIbZ7
M+J9Id215x3/yAWtKyClF7fUHc5Nem5ZOZM2f9JJZUPpD6b7acDfRiilnBGz5wXv
N7fR4vU9GJXtG7BMyFua6D1pge17meYHLCb+Vt26GLwKvigGdpMT5T4Bs27lm6u4
jQX30Zi3msJ3RmlG9jWcx5Vkk5gdAHSX+HoW28v4vccEu+QHfA8qCLJziceKfJXY
kkyS8JVYs2ifJKSA5geV915KyyArKI61owdR+acWrtwJvZEv9/YPE8fHsknnP12P
dj2xwVqCYN/Boy9NfIIDjFExa2K/E2VHlO5LhBN7Rc9hCUFx4Py+7f0h5VNZIEMn
KqsVw7OkirvRRVmKEqD71ir5IVog65Wtaufues0jHWWBqVbxAwvOigZDCSQJON6S
fajz/YzJKt+byKU+pZ4FKW1hqnxZGa7CmrgVM/CGwWftDgRpf3uwRfSBH4hvBY42
nFtCD/oOPTTr08L9WKNp2ThAjQooeD3eYzu+Bt6Hji1zkNAGbjoFyFl0aIUAoJFK
IJgR/APOGz0ikS3s2oNb8wcNZKQHSTcVeSf4oPQK+Te/YQbsEjStvw0Nj1ThOhrG
/ziLfQC6rwl2CfuHGnCa1iTDeMKMnjlI1kjQmQBGBy+0DRLa9aFev7uUjJimKJFy
VBBbp1LfCcuEwaYEtNE0eCGkrGuywcHfF+/cOQZqe0s8EnP26jg1asNnsd9iKtMN
zpkOnEdVsWoY4FHIyDTnHjwlezuC3j5smGdO7LhFHrrCmvJtZDdvo3Z7VvsMbMWx
i2Q2uqHnoWzZ2rVykbc6o35aAy3nWX4H3Fo03HirTcbuSvmXYKpN69tS3PvRs2gp
rzSNBW8AjH6W+2b89VkW/vB6KDL6zMeTDnOAalwPnq7Jhcf2nw18bJUE4Byp6PXq
4QbbS1Aj/bmrYI8vy8ATx3ax5MFr9FgNHq+7bA2x1Rpyd6+0v2HW7MDj59MABWZJ
LVXfT1dzVbzVnDPROMLbo6WKAFAiEZHzl4rnYSTjOSlVrYrmWsPJXHVkPHcPC7qv
4UrRAhrYDiL83CosWfcw1WxvaEb0Xu55Ja7aswZeXY38JPRfYDi/AFl4tTCmJjs9
sT1gdKxjdYYr45PEiNOAkFzbrMPn7YQAMe0e0JOzliOhg0LaMmMpu7wXF4KPk9N2
SQu9g+yMXwUf4nLDeBqfufcawCNq5oVeoDTgak367FPbsTlIXkUftQQpHxI90Ovg
sa8djnF5vB2iuomPrM4xU8TKVOCgg0iuqZNLg2Ig2SxQAG17qj++hpR9ennteMpv
/CVa88iHytxbOpmUedCsci2zWxcd08UieVk+NuGDxFD0oZEk639DwKoiIArT3qii
Jyw2cGnvjz8ge9e0InKJkGXChtBg/atdlUxoaNvnyhX/9OF+lcOySKbF1VtWMSd4
LmPCapKwnmS534Gu3sjjoVSe28NqgybD4pDZkhtL+opsPDhNJPXOJkNA56xAFG5V
v5Jg5Y7e6gf0vpY4QZMR5KK/ul/mmlFkT7cXD7XmAPOPvIQtHNm+7/8Nt6qmqF5n
VCC9LBhfSfiYQZe3D7YkZ76hBf30hBcAxXmeoj2mgiaeMo8JPDhecK8wgeOc+50t
dshKB+3E3xGbZM9UCGZCQ1N6VNFSLzuDax9CVpQBZGPcygPhpugkBFgCJV9PE8g6
yE2U9cMCe6GCmMo4gf3MPwRgkiPbCw7Adqx4vaUIPKQCsLBa6uKZfpiK+EZWyMhA
gMmFZzAYxw3Xq9so3342fDwunX3Q8s4Yhe7MVIhPImmuG0VY/f0wOuhrdNVaG555
EtMT+PHVOImMJU8B8jFGYBXlsoHledpoesghAFB3T05CW09IjYCBxYT7ZU4Gqftc
LnKLOE5RVdGY8irafCofHITF9hM33M6hMvQctnLdoKbaBqCwOR+91Ez/xo2RSKSV
BdFW/RD+uNturZ3XNCQoJlg6E63mtPTtecuIAArfyELBIWVvgnIN8OpuZccozfup
R7MGWxBFueZBRTVJnVNfUzoaOtu+Lll2pIHKIkpxbUdofxC+caBOjuwpaNmbsYMD
PzZSAFTtKnlRQoWZQmZ1XvKi9cNfXsMTc1H1KyRsFZKOqpXwhKvOPMHWU/bTjmXD
vi1rGwCbAo5KhMYkmtOIXVhXQtCyQnSWodWoGEfYklsrHBiWLxQVjdD/baAsQn6q
uH4mA3d9m4BOs4jxrnLdXTfXDvwCQ2SN/3QOlVft5SCuDtT6eBFLmWayOpRBDJMp
9osM/4aMFQrHWEfRXtmT7inn1fvnjJ3uSlxtp9Ue4ODs1xny+lgZFDl90716mMrF
RixYSJ+/fvzlGe9ofyV4N6Lk97TxVyXuRIAiPAuxRtHycOCNS03wD2riAKJ9r8YZ
v8iKOfOVTV7LHAnILKs3Fn4CsnvdXgZLDJug+CtUD93Bb2308QqUW/5W9zqrJCQY
hiZ+oWN/cKG3GcS4lMacwCIkXe5HBnt8oNn86fqcVmMi5Pw3BxEAUZeHYPzjH4OQ
Zyv5/y/qK4kIyZXa7LdSCayG1muCMNVPLSITPVi9Njd8WF6/Q7aNbVHAvn6qvl1U
6/s2NwK4Zxxt5tMBGXzGbZib4p29SSMF6+2AAe22WR3KrhoYd+BjvwAXw2bJLH8p
3XAkZjaanDJnoEfQHltgQ81Tkto726hhut3aqohdZkIb6/Inr6/eRPrwFYsoHoBe
cuK8EjiznAioQrQIRFe2tTDQ4P/u/yNyYKbtGd/yOCPFELqykvhMM+xltxdAyVWa
+0akXjNjpdlQU4CiEw3qy4xoGaIjkY19ufT0Dt94EfSZbiDgKdbTqoo5yLaOqRn0
MKUEKNUe+SBHm5I1G53zJXt2ckIgTNOlqw1m0kSYq0QqW+LcO71NAQw6fmdfZN1Y
aE0BnY3aa85Q1fwwwZXUJW0NRZhNufFuboduDFUDyxIaTTyItCthbLtvI11yhkQQ
fdnpbciedbCJrtoXYUPrJ0geHBx52HTCAzQY7LUwdaQKZbnfVJhdcOLy4zuMQuPr
cYKKHoC7SXsySqWSE+c7QWYtmcfGWUYBXjrSTYKQODK9kARadn5Ioeye8ZWd6jeJ
Il9xXukDSjiawuvAerdZLp0cPVvyQ4DxxwlljctcDNVeTgLvDp5NxqK6UwtaOpXW
IU6TSihaNx3ZyYX27JLbulknhG56ikC87TbN3aZVocNHDvlkmqH1PJXYvId1BtER
HzTDKyfW0aE84oT2sAE2hsCYmhBS0NfYTUmANyQEHzG1uqTd0Pmm4LD48Iisb2x6
0SlAZBTXJDo7mMoCsZvPhpW9X7bz6/1+9Vpcp/57KfqCZoBrtSUwBQD/cztdsk+v
ruogrdWy3/A6TrNazUPpIaDZZLKAXa3y51i63aNYdV6IktM3b4o/zcDg862tywib
er79P+AgS1qN+hMfdZOHmFoGQ+ieaaAalkrWwHntBVav7d9kvScYkJr2lvgJ10ok
7ePh9PlcaoJN6cRSBoK3lkObrwT3r5Knq6x04yMR5F7FvgabRiV3PGzogf7jujUm
fLjI/E8Xt3tgmz/yQ/F15izdhngwB5vQ9uWFFRH0qpIC25U9Dd0fLrw1ONGlxMtG
GQ966tsFgERlO6VP9TYl8EZsDqKl92Yo3DvAOxWx88pOFXZ96yj6y7nXmQOUBSfE
6BmuONDPCR7fM+l9R7zk4cP+RYIvYlZc9AQSYSc2lGJLy5ccL4Y/0tEpd7GG7M7X
AraSx3C8FZjPLEkXDs/77gQObE/WuotSm+jPc+cR4ANGnxMwwnuK9SEkqsh87cTD
TOfK0o/BCJBu1YyYazHM96Ntr0yPgYc0NqeA2awUnHk2HJU8af+lXeNBTdUgsYWy
jpJQ7qU8t3e2U/IOkevuzE2mq6OXyXmdhNhWBMFOLPZm0zyDd2MN7F+/d2hYeR9K
xmej5c3E6MGaaENzrRAToMrbg/mL6HnC3zFk2OEFKGKhPjXL4xGtmBUOEjcDORz/
pjMWpq71p24R8o6teHLW6zT5IZuPYtMIwgVzfjwyLQ8NSVIwXdBb4oRst9/qapoa
5MdzgTSJLACzcvzwdYVwTEva/8jfAiCGDZsOGN3L2W63t0udTKK/onzRmc0BN6f3
/071icnEurV4xtrK38cCWJT70vSw5yax8/w8xcuB2YY4lFowqPHtUmLfU6pY2ToO
fvdiKKw1sMmkbyH4aUH+Wru3pSUlRESF+L/SnfZ51MYHKGX/m3X3Tr7hFR7dXqrw
rF+2gz4U56EGEUBROLY4W+jlVYva2MTA/UTiLscrHLBOtnBj63VV8Yai12EeVylI
wQ5RRkpVEYxQM8b0vqceSJPtyoPT8Cq1r5UcjNHr2HQdrOqmRf4aEA/xHW0pbMIm
6zZdGrhhXZGL4ys1ItHqUVkNrrDX8MrK+8hGIJLmueMxYNIMNroSxDVKlxEuLBuE
cZ5+Q85GYF+AlXxKTRWlPdY99+wujTkzZ0qkiXmdhS2o7kd4VK7XoItos7G0dkHv
YfYbIvD+TCfCsejpwN4TA7WBZZbaeOcT6SArZD8vo890oBdOlOpusN/b+jOdwHUD
OvNyq066GlShmenQ60+rilHYBeEq1UPB2TL2p3IC00Epc9w0Jby+x5a0E1zYxtrk
cmDtUpPX9Mmo6KoxuJ8IvJEGK36F5zaVvwmm0eJvol0eoIS88JdPTGb4ChcC42Xv
iYyfVv2GjNogij3BQZEO/wpZbJtVqUwz4HvaLbZ+8SBq6Kc3+1Va18ROqIB5ZNia
KlLw1TCYxXBVeBWeCJWAeK3WgaDhWZlVLestxv6iPQPJQuDUWoky6z3dx4hTTUhf
lu5IbGGlOGpBM0WHjuGcjYh87RkS1Oz+DsdraA8HVDoavi4Q7lzY5Bts9C2S2Xp7
EAVKRnHpb8Xwx32YG1GW2jQWp288AV284OFpK8585FxUZUYFl3A1qscX0v4TLgse
qb0k5bW2ei1XV0zL0aIEmWhC3mBdWuI+HFDMM8T5rt8Pco6bAbn5QlRHwhrt3sic
0yQp/RCKuCatzZk7bisQdFTVluayclRk8MrQHxd3dr12SIJEmkcuzxGjWrkmw8zL
1XITv6P94r71uYp7IkE8wEfCfNzt+u2WlSR4G9Bfnp3eIIcqXftlJVNc1NdOqTAw
xCxf/VBRYv9fjCcxpQ77uIpRMTqthbnD5JcTbpnq4xlL3qfVlXZx8E+8ZCzJDEpS
urHSCj87GLrl1k+d21N3WnJp+1ockCXVS3cEiRuzZ5+cSxJ26qJYUL8iAqpIthD4
qWuI7+IA+Xns56MoZXXwiSHoQp2cDuzZ99n7181YmBE9sZ4ejiMEUm1sIIx0GY+e
dNcbJVI2pQ9yp9m9MDklMdA6s4JSyDA22iR4L32cuze/qD7yPbZpr5Gr61j2BGdw
vUC8r/zR4bhhhi1d40Uo5Cl+R7GpSzdDQXCuJjp5iZYEl8kkzTT5p2Wj24faqIgy
Co0XoJ5HMMX8siWWa8goD36BLF/1fxZVXF9v0SKatQk2HWdLGswAZKOfK4ojL12V
h4FPsWxKruobNoFPKMD7Cq7OAHBFO037SPJixAdy7BMOvypE2uhAgRXgkJIklY2J
NCGQ6FNHYxi9GLrlFGd5CKnHdERX8QT3vVA50VmlytIDagY354TyUXIm+cAc1o5S
I5PZ/hsJ0kzoyiLwXXfbtAGqhvgq6cdwZ4+AvnioAlVTtp5ucIf4+o8M1Bm/fByW
CQ7pSesUaGVuIJxmh3JBICXc090W8975X7N6SyRJpRACReMJtSiEFcKLo5tD5eP8
wDlJnwTqND2zDH3okdlYfrL14cnx42ouTK/0O/wjfUs9Jnb1dASFPv51spPkVB2X
AWirlQkdtTsMQPYV7ezxQ6UP4hsolgPDfZm9b6wL23bd7b+iUFDR+fkqsuRlK6WN
H9jBSo4/blTtFg6NFdQDYNlde3yUpP0Ipx2fv83YfPkYYoUeNKNRudEpk/IOsn2M
xx0ryDxeOIECmWZthSunlghWgoTEz1DBhLL4V4kNuKyLAw9VoKFjV81g0C630hTf
XyskKwtk7EUlrgh4VdzyeP0sZiwUNR4VVccu5eSIaWboBHjIjSbBcOrv/O+0aA9C
c9XSdshN5Tc+nCMCftjvWHKJRrYxFdHWF5EG98TRCv4m3gkhCuxGppWAy304PrSc
8ZOhnuHo7hPxuJ/Wkhj9aHmN5UYru5MbZWyU30+jrytDjtjY+fIZ4kv8YOuI6moN
VhM7qwHd5JieYhH7gVRrDXJdoCp81yvFRehDc45laW2YBhvWPirhRrAJGtaldVRl
YeT8hLbk+S47dCzBL0r3SGbXOsm6NeECHBFa74CdSci4GGuT+Funo6ENZtEcg7zn
DRosN5stDVcE/S5UoEAKQ/GZThd1P6ZUKszKu9rmJZEIGBT5fKX8jkuSp1LTQ8gH
X+VClnhC+1iY9r1iwQUv73NXrSv9KUSoWY195GgAwmLvfopcmiAjWVi7Pf/SWDHW
Ddg/Ln9O6ebk4dnS2Vv2XwnDe2KRkMmKldhv2p+RVLsrYXCx+vsNy50DsZq4gAiC
or0+VHGIkCpWY/bv+AtY88p9SdEJ7pMrzGc0v4u18zntmp917Bxk8VM8hoshKGpI
sWajW+OKKh98ckXOa3LY+ceetG6/wh4GE+Bq0oue1YkSbr3lZQFSb77NvcDvbbL0
fQbTOrxuVdeLjDcFUwJGLEgWSs4RhPtzlfGmn2BycMTXazC0/NpT6cLyyIuNEZdQ
ZHDR8NfsubigTmeiovvmMO3RWeKx2GbwhWEzwGqhwXb9lSpBRG9BK8X+NepnJp/x
H6YvKYR9Xel7QarStSLB86Z/beOFLK94Z7O5ttC4I5YDV2OCuQffmvgnYV8TMg1d
rs516q7nTc0oLzztwoQAKY5G/klIDtunM5KI/SGgF1S4BudM8vl0rD3wfOJm1v7c
oadcS7rDnch8pUTkJlC6M0+NnXoyCdAnZUZmfsBBvbzXulvw6IrwKDQT8n9oQDaa
UjGEt3e9z9bWHfguBO8DC8VmgZ0X04ypPEZTTAYSzuhYfKY5Md1lzkrLDnp9j84b
ULCX86rNn7ghx0R0RnSluliCfQL2G3Rs7b8aKywvQqvDwsJ6Ecsn3PFIhrgVZ2+V
o/Lwr4y5LlCQN2Kdg0zr8vdd4wUrCQ96QaVaU7jfIhX4VFDCNo72eINvi3tqlqqu
nr9AdHP/O047Vxf7rY6cEJZPWJAuLa2ej3Y3rd0Wyzk9gdtz7LHlcpLcTMeu5+lh
iS3v3GeoAXbJafXa6rPxwBRgR7d4zKJdvrb6Lf1RIMwwtKpXoM3JePqBfSoA+fa8
rsiSVFXJsK90YIrmVP17S4MBk6DgaKsYaGDQGqmLq/f/qICYtnILAVbO8Ahdrne8
1Po2nnRZOlosroBD3VXbXxqPvWQQbQ/T4jcMiJ442R1bglFOWkjE5L1STPNlWcB5
xL778/HxWdJsjZTe5535uGgbt+u1wWSgMR2BbqIBPXS8Z/TTcdv91m/Icc2VZmzx
4KIspvwhnkHT8lVkwZaETbSDl/6Q2/1ys1Bv6d7/JrQGeV2g1Ff3E9LYXafsCTsq
/ZLqr+WH+dadtR9ZqU9CURjNU7DduD1SQtShloba7MouDJ7c38eCXIRiqkFDSP3J
lsz2aNoFB0wsrmuEFkcVd4t6raOL2vBFc8MbkvoceuqcU7cCHaBZJGzctmdTsXG7
GNqOPGa5ijH9rP5BSMoCJJCjiElvthfA3h9I17K8Y9fvj1A2daClpDH8c0kdo9js
mJg1wkEgefPsQDc9DFb/Te7exxAUbzrxKN2vWEJfx4A9O9eOzq7o41FIHOh8MgrO
MGWC6SaCxdsyw3Ixrdt1ZWW6V8NADPeZqt3GpUzEfb6cmT7np9dhOaExmmKbekze
Z1sLgM7l5gYhFPwleebwrOyvYg2/oEEdeNjfe35eoRqLqnx9YYJIrq49dMjMtQgl
RQKeYSvhGR6P2d1dQZ0/lqXX0E+1wM7IzPN3oP0kHzMZIxap2el+oaNOehcNrSyK
uIgQ6NfrXv7Rr66HCJAUcFUbc4uSPRzrs/kF2vJwCY0//067prIXfy2Lkwy+Al7x
dAtHMBKVM8CwKvVflt8OyvNdAI3SkvkCtdt+zIwEOJDp35yr+nuRb7VPaSt6ReGw
FHXqH25zXJLRE1909R99vUM7Bcb4ujXLu7XBxdYeP7r1PfN8VX87GbMILtxh3bMg
injA422nCX+AuFGNAhvI61BVM75h+FsUFugf4l/ze9mHDysnKOvFBx5sISSK96a1
/Y7QcZjRtyf9iAc5ajV1fVFVS09ZxVSFKhyd/DRQ9E3mV1ki+ob/jbau65SmNRoO
WQYpSPCZrbNSl3UjnKIkFii8F6oXoZzqESnmxqKF9+4vsSj7wsZNzzCyVPXnsdqo
acmHU2pWK2wLYSH8puyJDIMk7T99U6VONJYv2eG94uw432GWNeynbiRvEKs7avsF
5Em/UV5Stv08Behd0FufCtBD2RNJ+1anbQfBrCWzggLL1/pjPdG9BESovdv5iq6r
W5ndwM+chzHqLWWZkhK91Rb3AzgjPal19Vy9p5jrK1GO2gjDMlCIAlBy0qjw8ojc
7NXJgbnkGXPZ6ofjKKW8DYFeNB03LettwkygTQzpez+cd82AeHzy1kDlbMxH9xtm
BzhqYHNvG6Mwt0ZpEAfMrAdXjfQPoIykn2KPjHh81WjddNS31IR9DFr8I8H/N8YN
+buVaoOXPyS73jXBl8egB4b4y1eprI4VXdddTV90AI/IaP+fKXjmSj66xvA1u2Zf
w9AtBCgDI82xMe87ukJvdZRbj+gIpHmCkDB3gqPD2EmvRoF/aXSlT+t3z2FHlop2
cPSOeG/Jgnvausvto29Q3ADUNAtH807Bw3wl+nHLRejTn4dGJOXytU1QE7oDBSrd
amzaCyjALWsep6WCpFQI/PR6MB8h+FkzEvUW9RiB9VPfmEZnv84EKFOGKbRxe6JB
67uGAmabvlP/vbVwQat8nCxsKD1X4Mnc12DIUaIM/x3NWjb6/d80ivBsNV/9cR/J
5KEeC3xpvHOe9Q2Qt+uXbw8ybBvkwh8cm8Qll6Sz+9zGILvrbviJBw0uOzES6vRH
64PsXkS8eZR4kadFKUXwgWEgiaP73YHc3bB2XyqAegcl0Rm3e4B9V25kmLXgiehH
yv2oiw050hoOkzFll5z9lGNZmf4oInhuEuxXZX1xXIzzoSw+3JaK9Q8ph+zGH1t6
exaB1LSHSFcP9V565d0kH2IawGP9Sn5oCIl76hAfUb4SD5UwWqYfsFhwz7vRibjR
Cm8DkO4M2ERC4/qQdF054SWKXzCvCD4U6N08r5lvAPm/EEkUXX3CFV51nVc55RhV
RlbZ6tz+lOanJHl/mMWk4cJat0d27p65Vu2HwOT14tYM88gnpVHIiAi2Ttka1/NS
xyy001lQAjsr+1hAqlYeyiaTSFxjQPI3L8V/Wpsk/n7yY0JCtcQKT7ti1QnEoqVj
MrCxJHY7H735e5sScOxA+Qwa2lw0/flreGaX007ityi0nQ4YzHGWezSSMnnkdg2k
ADPSDROqgjNbmbT3F9bUMsj/OJFYnrzmKgpWsdxMzCFeqfCA+HiiBncePjHaw3Pp
gAyOgLRemOZoj0q8FQoNSUaQRNaILNLLxsv6ytsETpWcDUoihKOG0EsNR/Qw/2IN
QMrpbgs07wnvFZhspwQD/r6kb/yYGU8MpktekZxkRSUZjOFqxo8j0/3WJYa3KeKK
RWfU5l3lZDr4LoyNlEKWchMTNzxZhNoOq/8G6TY1REZXye77wSUPC17N8qHOEmsr
oNi9xq2XMLv45oN8AELBX42TA+qLSM/3Zrw5U+GNSM0jMp4/an5eNffvAF7/W+fM
WSIiM7WiiW0KaajSsci3SyywihMKiyf2u/hUHnilewTGJLn6zKXI/bVCeGSvTaii
+55ZCcwW7Cdi0l2jZ2H/qUMfCdJkqoT/xU0l7hb0jrpVRgd5+xlCAsUPi55TAQTk
GLi6zA+iT7DDc/NevId3ZWE+oECDpreH48/60RWgDNLJqIggm2Eyf+oVteC0+RY0
hVifMyYHGvUAgmKHkYx1hnKiwFXi0O4MOJc7rsgRzUQQUKSSYO49Qo4/A2x3lWT7
2QbmmmOASOM3WBuVqBq1ccFPTqljOti23YH5XaxuEaKIAxTJWv/1vnmjOCYeb2k8
XIs50HlYZWtZ8C4hb7mjenoNf3fSrgMI3MCLswpV/9uHibLFR3dKEZvYeVvHJl6L
I8gl/iyBXcbXbv49XujeKQxOIinoD4OAxpxOIPunaLK93uw+3IV+D/81bPCAymsQ
t7WS5DMvghmfIOywSstUSKHI3Bgg4gaVVjir69sO2oobWNe5DnIRGV0cjEHbcd39
RtLbWhx6t+JQXIezXsLCO6LWDqxbkXnz4Q4CX0m7K0p17XVvkcgWT6YMOCBoJcfA
3rQ3XxlzSRXdw/0FIA3FUiz+psC1kF3t3lryHLBa4DjsDw/erhCASBODtw4+jCkC
AGjdRp8Rr+gNbT/csephzASvYbDTC/mB/xf0Yjauj8ESDa9ogYGfnI+gtnFuA41B
OYtECts1/iJrNnkQD+l5l+mUJdIVMHd/FATVMhpWnt3PiZI0/oyh9zF4MYW9WiGU
RFe0QJdV2phNcSa+CKs6tDovoxq2HOV2a64Y8KjfJLBj8jaEcnB+Q0CPJ1Sv/4uw
+5xT8mMhAQnLe26iVX5elYJ4wnY62P5kPurBttdmXijauzKklqVuoe3H/5bBfeww
pHtqtZ2hcqOqS5QXzYHgpT+JEY33nP/Evsjg27WGg+qkIJd9zGiBhTyGKfGa0x1v
22rXgOsK+dZG8wtJDXCH23eDcw76Eu3jlumJ0uJ54ScUdA+2oG24LV462c65Ql2U
gYu07cu8sK1bXVorQiWF5iCKPrBu0S0nAbovC6UUMRlO9Ja2Pxstv76LGB7UNsBo
D2tzW/WO5b2GzpFfDTFswBKLthqbwseRucUeIq7e5uQaqnAGKDkEe9zVjGKwbvnM
GBaWenGdlX31HgllPjD/ftMCX8Z9w5yOUxAZmHkLBPtPyQZI3LCjq1fPl2rYHal0
uqsnZUbDXhg3HBOCpK2CZQUgJOkYi+mzUPVuPSqS+jkcp3z+5TgfmRvqLr81vRst
6ZCggxbWZHEABpJ4vHJ4ouLTD3+ZI3ry4n2JP3RIY1TqQsQuqj2pUWxqtecYqnxR
3ZgVuOfhNpOYVGymdCU5M1KDsR1YfrnqiA5SrBAYKWbTfvhMJ1kw0yTwSxm0NyyG
JHpP0QIRgeVhPEKyDY5j4FejzpjwDrgbiYb0yjz6ZRSAiGQQcZN/EEY04xMOQz+o
74gOglxKuBTRF6DYmMWsup8UOSKDSnKzTlZjNXJ67/pXO4gXPyP0Y7IGkQm5fGFt
vVmd4BTGApYp64J5kISNbydNQbxcrZ8+bJQHprQeUKg4OPw62Ofh+yX6+w/A6oZn
NDOYRUjsDhmS1iBSGKNrBqBz0t+LIno6itR8mqWKc+Eb1bats0scIXEW3yHpVIlX
BCfhTeFoBsizZSbBaWl8r//FJoH/vmp+uPLUtH77OANRgRbMBl/4ihi55jij6bEE
bdmzdXN8Ywo4a2K77h79SsWCMJWaMLWOyqgLBstARUnfejbMjM7nOW++qdKAgixm
5MTKcPIr3SyCQDepLu5ixEDP4Xu2MrJL3PKa+2cTTUuAaHdVXLMMDs4OWKjsI677
01R6M0SFBeyl4Kcy0Rq3KblE6JtpdSa7DgJb9Xsb88vkFFOrQCJQU+HnDIEOrDA4
YA/tX6HeWHlV2+vx1xBpL/MFvNnfBoZdX7bYfoF8upB0qXIDaQbg1iOKVMF3m2Hf
6SFXvVZ466Xk0feGrYsPAsWb/S4mMrefhvLl8paBjodwlqakDzZWrwtCQ8KGBnpg
wGRIJj35gvW7+CZx8Ri7HhIgcvhMP778YGVVABvmu1zdVckVjmRdO77gIBxj7XLP
IwWSPb7hLm6LnlPv9NoORkjLSf8PGNiFbkSyYg1K30YJ8Ogs6FQZjrb9e9vpQj6K
8cia8QbeFe2Q5ZDktrIGKHWx0ULi5DUtp+WYGkdfFL+0fC8ThXrBHh/5PgP4h58u
jc/Pcnj+iDo3n/YTSv5iOlYTzztyHJfcz/aBTOftArO7x57v3SoPGO9LTsieDTPT
LwZV9vLVE906kwssEq15hdI5yMjXDqjQeOrsQGawi3j0/t3BUnUYsDW+/v6uKr08
0lRMyKzB7lwXW30KSPftqHkHq9aJI948+gKW69L2En+X6ETtloY4oN78HH0Ryy3J
9xxt+lydNQCWqNQ/rheYoZw7Nljiz8EMCl8zZrx8rChkgtRaxu83IzjNIm63DNzT
nEUlHgxc5yX9Y6faOHKaG8tDV66J2aisQAGnCx7gSdRCpRviYJ4nIKR2Ue+xnGLX
EIWIOc9XJdlq/k9u7RyqHSJBagQ93ryLkG9+t72hYrXdJaXC80j/Ivkz2fSJif+f
3RHnyTDSdjgQ89HU5zxm3pSFTSoEypVMuYQA0I0TKREYu0s/9VBU+FDZAq6WANYj
0uswi9egDBF72sWIdOnRhNuIs/L7X0+DeNNc2N+UhMv0IF7PTkU2a/omi/5CzJeZ
ddeIOGAjtivqu75vmmzByezTWBVIgIiHoXE7qT6zseGJfCh2wTV4rI1JhxDy3Ljg
JYf8qkompkX5zLfDIm2//uPZTwzY4Q0zsa9C+Y+91Bm5nBvWFElOAkN5q5JFMD2Z
G1GQXyNwKcTxhmXRL96wOCLB/Xmah4uY6Kj2cVlWSt73lnB8ugI8ULvDz4TRgNoE
Bc9DRNSOL2paIg61h4IODoI8pJKPXY8As29LgJ8uZdz3VhQdhV65xzxkiwmzcvu8
87Fz5TvWR21kQFYaXkco+T9wChVsRufCsupY5D+nBVlpu+wAd3YeFUYeP5xMFTXH
1gIAJ7kVxIZ3J7z3LTNJKLtJMmuzhVgZFKHd+FiAdTJKJDCrtn5s8DVrIFA50RK6
lVq00MD7hJD6t9pabTk51ryXmP3A6moRoESXBWndX5JzbZ5LcCyeO7sRX4ahLPOM
cWqIfXWp6FolBkqbL7iu+plxT3lyCUlwmFQFek0NqviFk0a3Oba9XDQ6Suh5hD2Q
+syaQGHYIpH/5QiUW6IKmSm1mI8RlOoOAFrhXqUvinMOddH4xL/VWN0KoAC23jrz
A8XhKNMv/pKn/dV9ZCO9MXY2uDIeM3hqdFa7ynRGXy/8Vv5w/inSYk9JUqgAakct
FzFFG18fAY+lUVNnNuCi/qhPgLkJ193emVWi4ZOlx5e5byf7f2sB7cZIP9mkOR+y
6B57eU2oW1q8Tv7u0diP6abVtgNTpfZ5Csfd51SHmSzrSDdXvh5G9jI39+ZrmPmS
N3BpQWtW2WjGksEsDldKjMnfNzPtd4khbE2ROEon/n6qUOnFxJxAWIWBKDQeQKmp
FQjvJS4JNpy21KWI3tJaLVZLPVuOSxAoZcYkq+zJiFua9lS8KpE+VBT5twJIrBHQ
3csj5CTnOkCX/yKATwz5sE3tE1I4BRhcZOFiLOJhPFNfpEiCm/daVXoW5stMlMTz
yT4OZ8Mpvo+ZZLQWwsXCO2IUUBlgWkrpobvzdAkCn8E+jsU/I4IRRrqfwy1GFa3R
tZVkA32+zFDpbs56NZUna4asWS9Nn3phXMO6JUXW8h5BmBacHjAxi2SphTbqij8k
zgImYR9O+PEU+uM+bfcltM382SOsXc3zvrKRxSermAqkeulzVpRZQ9v6lLvsLAY6
0p0oruR1GVfkZnTfvbTWoM0hf1JBwlB5A04EIX7feHavLbRJWKHtVWWnRTDVnU4t
KZXKblYdbNk3rzBpI5Rgrwxw7FbZYhhMpxM4qsYlMw6wHCC2Qo8gFaV7tOKjYnyZ
pg4RWy6I3Hoa6GuO+/r8HSYZ5/OnMVEAwzDb5sbZ+9lHs5FjWwaCYbVarJ8gQpZv
nJciXwCZolGWWEEcwhApvPTlVIftBN1HCWKQOb45mtZ4+JMpaTsJ3ZQLtEZqBQop
UfWHspMZMLd8JOy8ywWQZqJq9BD7xQeZ5dTGQaODn/iKajVUqQn/mfZ9WkfNULRu
0S0XndHh72/vyk+iGKwa5iyh2aR5ziT4ju1ntPJeMLl17y+Tl8Vjp988IDsOfOCZ
+falG/8z1iehYn+gYkdrz+SewWY/Q0wWeg3i5WjY6GClwRJxzjvk2yw8xBC8p70Q
OA9f6Q36MZL3Bl86i9CSZrdb0IQLjMP/LHVVf51N5pFJM74ZC2AiLOZ8t0FOHoyC
zudtteBgH3MHk+kjPuqYN6vfnwWpZE/eAq9F5PpUOogOCH7qsuOIprm1r+JrxhOj
aHV9RixNPkGJ+YIIsVYKo8hfQO0vv05v4tz6wrwcZ2+dmDs8RI/uJ8BdAy94JieF
o2Mn/AxMk9+jE54vJRRVtrVpZY5Z5sCrCXNGrBfqsnZtbjBTXoGUMoh0GEi5fdU8
OJL/UlDmoEYPZD55Im8yKpEcA5GswvUOLe86KgNizTkHqlGn0dW0+GLaXttGgzTg
Ufmkx91a+3+SrYaL2EIcBR4wn0H6HSss35eVQHGxXoGERp9GyiVvhCg74894J578
vo1AbfTcfmmPKaqMwWs38O34iumBkF0CquFAq1UJA9DVifn5yUL8fc/VZtxcPj9Z
55Z606i/hfbZeiexMbe99LmOnVXvqjTUP/lBT4Xcz39VHE2AYRgw/17LcyUNt3+J
e7XdGdu8KT3hyDIJJWxNEvJ1uPVHmirzHEQsZspJB9ToNOfz0PIau6y20klKhSCi
lhQ5HdXU8MKRyPzNk0RLi23lkvdZpI33RwIcB0Lw6wHJRd4N0IVibxG3LVEPqFOU
XNqfla7M4rW7ihGD56BmUOZYvqb9SNTETaxRIxTFvEsAV9Y8mbtHAkT2haqhXncC
vIpFYiPwvMgKTKQw/NvwSsUHq/P15TA2KkC4dI+YvyHukTvnduJEqNP+6t7b7Nzz
qqCf2ZMgE8LVRJYX/e5kK89BfZ1/GgA0yiz0ASz6nugbbdbj3KKv26OesmGW2ehR
QHoGC29HTbA9eeSbaJz/iPcjR2DTw8X94XWbMhviMLmz3si2Q850m5ZTydneHtaX
CRrCEXmJwD6M8+kbqYySL8y/WnRJJ6r6QcxdNRa8zk0jZoV1QfTHgUUpqr/yIYdH
i6a+fBP77ouxvy2BfkbiAYuqRhLax2EZYSlgXTPE30Fzn24r+5W6TCr9OdMXni4p
6SHaGSlFJTAWmIRoAcoLsaH87Sef0uJeHUEhKhFxMOM8GsCZcxOtsnLL6bQT7sXY
GA50SwnTj1BY5kLLMa3uQ+GlyBV0MULBg9G2gHrxYnUhYVNSxueP8oHMY/+W8PNl
YzPeQXaAtyIiTZfE/EWcbGC8wb2ceLfr/YVzuaPbJ/qvqHNe/Q45W5yVS/q6ItCp
Os1hTuOSR5mWtuKJsDtu/d/8A0jSI0VPkG5vJMUkehuc6nOrwk22es2jQn0ScC04
PZyo8ZCJZg4XuT4VYGcD2iCGSrJwKNMqJRHZkPtrFwaPJDl52c1mJITkB1mptkfs
zY5tpEdbNfmKhQKP6xz7SIJSR0Gh2BuGXtObg/mA4bYDxmhrcu1J3X6u5E0G2f7F
559WX4tP1oI6ur8G3KVe6EzI0BWkI+ops5TUY8oW2J/LD6ZxtCmMJE7kq5R/WChC
V3oU6C254hekl9FUS7HhzzVkS/hwZ90UHA4yGWjwepQAa1z+ojy/RiXNyHlErOZU
TBNWpCjnt8rBwezpZSE/OyghnxgpGwb6GWKauEnm7uskw1P25+DPUPdHdDW7CXr4
SUpDfXUXE2u1ZgjTbrrrQeKgI8RCJ0Cj63r5okDCS3o6gNxahAMhjiGKR8wkKOtn
iB5ATxGFMkTX6K79c34ORb03dXODYfEDktRI98fVHZlLadxaRRcUUYMy9TTkd4y+
xmL44o4T86l7F2TpYlydViie7i+KtAkXHHgHLJV91LaTIkso4TRrdhjLKS/vSQdw
8BBDoCPdRe0DfTNXE7iGZskyENmArwRgraNeZUmv0oZHnWyPQqoRFZlTpEXFReKs
kDJqnRB2eaEhtxWcqHGTT/0CQDIIkTYyIR7dXgbCAWx6AIxr+SlNcFsLqWBtyJtG
6e23YXGom27CCa03UjFOXopAzcM/H/e0EBAYf4IyVpeN5mabwQEdV2a1CSxBIz7V
bZQFpK3NuyXOZk4orhyguhzWw/pkL9+Y3JTNvLQvMqJQX45N+LTSNfpmQFhA0Uc8
a+3lHdF/m+vf5E344jgLBCWsdFpPPLSxUXrfd8Ua1PtCCAiYYew+f8RZ8Go5Tb2T
ZMdEV2iifpoWtxobS/Ttu6B3oOSEqjdAe4C1Ag3YZyK9fODLzOLfk7DPW7muyjlq
VtsxITIaKIDfoMRrkpE1WFHE4Yhtjfg4q/hOL1XrlaBDkIa5UyPMgvaNdFkiHs/8
HBgeTxwuiwL4GLBsf6nnAwPq3ZILi7DqOHGFSlsJwT+l/llbkBzQNNlQ3jC/bMDO
Ws+K7AN7o/pP51Fv4ZmyWILB02foMkPUt60TTrewNypMPHVmJ7dTEpVyFq67MLR5
xgVrwuut8lI9wrfJdTTfr+km1KlrjffUkLeXbBViW6tbB+esNeSMixUu4hOGWbzb
qSD3roEXVh7WORrRcHjbl/9w5ur6ehaP4DpT5R1kGigEDv+4FVNlSV4vPzYZR7xF
HL6nRQobHCKW/ztzOV+r1lW7wMMb3FXTp0hfhiljzT6qxdbk/QK23JPNAPWq+xhy
yGosmXgxQjt1T9AsvxR8VnVdUjCvJSGCYRq3WixwlG83S4pb+OxjEppG8Qhx6DUD
lOj7Qasi9+cr62ZHHOaBAcpN+RkkELYhvtRZYbaGqhtdCG3Pn2CBGJ0j97meu3Gd
p6Zho/Gfr3hxDgRbN54MWe8HoLYIvIMUR3orkg6Ctw3A7Z+jvVTbdVnjQ+zf9V6M
K7BuG3RiEtq+mkkrzmar+jHaPWEWNFCpFeO/8C8796nS6FpvGYGV+YkBQAfA52Qe
4bDHArcjid/2VpThAA1SDyKAparJUE3tX9NZor4IAGg8HzHgL/A0xiNXnqs9U6rY
k1ONL7E9om3vsVb7pdghn8XbMKVswuvau3crKJWaTK8d0Bn8BX+nH0SQ5vD2KUha
XBUXptu27QFjoL64eEOqWlwRLnW4AHoCkrF70O2TRaG3lvTpTUNWVhQMM2NdRfPn
HpkV1kVAuC1u7QTd8OOwQwexAg5pHbEOBjPYWAaFxueTw/NUBpCFgGv7PK5y1Zkb
bjemcPrJKiSdZyWxMaRY644I7C4F5MH3pnHzBYgYnMkLQvLgQy/l3SRnFSsYHHaB
QPIWQMbIciuGWgAcPn6d9m7oHAIEf6geV35SV+KROVPVZdXkuNitnfnyJE2T8NgP
ZdLDbkmW1o35eH2chDTymLxbRshynJZYjmQRAEgPQIa49i2rtPd85A3tKonb8+z0
S1N9PsIfqiQmXoXDKSuGZX2EXGHBdomjvwWb0JA5eAKzGVwxhGy0A3dEC2AQqNhT
eliOlpj2CKPPbgetIR7x6prNJzQY6ujlYSvSc3bSy1yCWC/xSRkF7g6NPwAA46h8
csqPahnSSWHxZjHpaxbn0FaiPXtzn/GTE2wrfFYTLwGu3hr555oE/y2EBXu13QN3
XBFn0iP23Lbs6Wfgw3V5/u/KwyXAP0+DZRMCH7ijEQ7oBJRBGeUFeiaX3UYiit39
HuWFpjIhY8FLRnMuTECN0LH/tGDbq8YC6WMji+nV41SiaX4CZalYttSWepHSmC73
s4hXYhUdMzf/f4gjyicsHVhzAK+H4mxjBPosqsOGbbRv65BlkzFjn0TBpnDG9nwE
mUQ9s0EF+PrSGDarvbqSggT1jceqi9Xvg6en5wiZUXYmIE/iXq6PZKp/z4zVMIMm
QWKCAd8DiYCyNTrdWr9/VpikaDpwF0+ca8kACXl9h+qLiUTq+IqJO1Dyx2zS2yK3
K5xk2zSnsxoQxUenvVsXi0uE9N1ttwMq/O+dzhpLN4AAcjqhtgIFcvbZHascDrNB
3htGjijWTeeI90fG2rtnC0H3bnPbuzr+dqRYFCk9LE37imBXgQTRRepauQQd0mia
PnS8Nl7sLS4Q6QQFtICash339lJfphlPMVltr2DT61WGnHkOBNTzTCJ+gVQOx9v3
GWUMrwneclprOtn+2Ve9wPQxUd7Rqrmyheouy2m6i6aJ2fW/xaqvzLDXXtt1/mWz
loJkHesdi7pd50YMtmoALY1/fiPPM4yO10YCaeTGyIm++YsZVwKZ6RMMVM9jnYZH
9xN4oRjvczLHodoYxyWjEapaW+35kLoDA13aslnW1UqRBjvrfMkrocr6HRzxZvXj
cvWk3kZd10dPWfLHggeQDFj2ZyhiT9be/ioAnPzC6uy+2R0Dfr43E8HQolmTCmFV
RpXPEF8dgbatgeqLVxwIHuAre+1x0q+8PA9AOO2hm5C5+mbF+ys+G8GQb56Hhjsq
yKgHYHO530muvvX/mvqtgY+i11hZKjnOhHZYAw2NGsOpqYI6H0JORLJQcqTz/T3x
cjIzO5JAsmL0UdwO7cooyikPPAbX3E8ox0yg/Sy3pzM4fdSQaj92LY7f9pY30nJC
a9kH8LRCkHku2Fwgob3MYAnjP2m8Gx2k90TQ9Xbe9DjPslOkoP6rrI59EWIhKr24
mEogrBz5TLHKK1UgoRwfAz+kRP8XyuK7uC1dnuA4pcfV7ajPo7LnpR7DaLJvZGZV
KYZvhfPnJDPV1bQ6AOkMCA9POqlmWRZWrbm6EAFHF4D2aCD+cTummvTUo2z5Lul8
mawBakVdYfjI14X3P8WlRJVT3qR6SNbjQJUkWRQZ1JYU8OBkc5lGc0WxOXLISTNY
I/qTfI8mBn3zPS4Fs/t1JA3WX2m7uJ4bK2U+0iujzyigAKofz3JlLSqaW0ffv9SH
rjS5ZSk+0UdZuXyvt7kJaCzNPMTg3OCwuihMD12CLPr7AkOgkkgOre/cGNLX/E83
FOhYPiZOXBVLwcSNBd16opL92ywcpSm65Ytor+CgWrLNxWnfDw1IgnVo1W84sU/9
CURBW//aYGBZJ9IeLDHBUj0QaSAiLtDVEPJ+YBdBqX8/lUuOBpt4X0kEmGhDEpLk
oiNVL8YQMc6vPzfgW0i+8cx+x+aXaOb9VyVnzxRoyu5vGOGv40qYKB7Uj5939SPP
SP5Xv6AaectQ633OylrgsqeWSy6lSZifrwnUxWz8lJ/jp38cfrkNTrY5MWfPR+Jm
6jFrSAxNSZnOqe1dMLh6FQe9kjtYnzODESBPAyzVAN13CLSd2yGv2i6cqghqcYIm
1pP+1z1odu/LuYiymdnuJtKN15YrLL89cq1Xxx12txGdU4haTAS6Gs+3G/HL7pO5
g+26UzErfwBT6LmeayK4ONWvw0244JUwcha+5sr2IYZN1eW60mekeIl75/66E7Mr
y49HDtZeoYgsYIoO9r5PZ5o0XzrL4C98TxpPcPunllzk7T3YqR7DAQEt4gywDquv
EbqpDjzo4JB1snlu2MLa3KSKxVhNOWYmtRfVCZXWcXhNkujT+lxCzmDAa8l80Fz/
nZzRfkbmkF4xcVwSbwnmRHAAcEx+cPqkPs8qapYwjr07BJCbbRxQ+BvrAP2wsjsI
d/uJP9bu3L1gq1OvytYkmVYVooDNWr/hzDWBlo8mRMMY6/GOaE86shsqse+QyAG/
9SzDvnAL25h1Kjn6o8Lh0tdLXKznBQHHwDO0+TvcY+G+h4Gq8R76g6ffL3dZX/B8
Mvho1VzD572xnWytZMtA1QvzzsSkTmdzWsXv8GMexYyxeL78Udx4tor4AK4GnMIX
dSd4odSdM5R4KEVx5H9vuCS5nt2iKCv87tPZ9+EhZbZSHhgR2rTQ0ThcoJO3aDiy
MoCpKBhu3k7KgyxwhMmOtcj7jF4rGzEU2e9ghUDQFl2/zbe/7GZ90ifL++R1dudF
bKWrRlm40yRJs07NXeZIjKaKqh0l82BMDaUFsjA9YlBMQfayXCx7972f8OtVkQNO
SrOJxCCMKjZ6vnJlNsHIwwnIYpJQPJP7HFBWPGI4tnbNoM9jGfWRrXtS6Ogi7xUj
MjWKEpykLTI6mSTBHA9kd50InubhCYdRldf/Zs0ROWhh7L6H6Jx3YBulIsbEYY30
+52ZbUaX7hh5qoYHpVFsjAbfRVKapi3iTLxBP5aWUtPCmIypQDxUhN3T+X7+ep0P
NCqQeXku9ZyDbOY76WzFhUudufw7JXAQPeuT8i4JIxQhhq8gLQTCYGZbLui3hJ5x
YDiRmz8A3WNqGGN+dFPrayzvTtqovUDhzQ5IBJAWbm8Yh6A/j/RI4wvGpnD+W3+V
7BM2Ju8LyjZ9Y+X9Czd7qqPLYH6exUOAQ4YjcwvQVeB89sc0ZcfLhKnL/A2IiF4T
DTUdiCquOjKAztnL/6uSpWILWNJCGm5kWyQ4eUNobjxFQsX464fD4/WQ+H1210uN
RhUyr7ZK5w+VYiI9XooIqaDRFQZk2IU3E3LDYWH8ykN0HWDw35TXoyzTt5Mu7P4t
TY8mEB1/z8G61BAZoHZ46pqzfUa6ncuG8oCe8Q1b21KwhWdSrQdWQL1aZ3lrJRVx
2+Q0B7w/q94IR8WlyYS5xn8nretKz0Xvk/2+2tfCU+ia1vAFy9GSYd94kyjLLqHX
dycweXDRnp+tFFvDNKCAMQ8EU8sk7NlQSmand3tYvsVn/IzDhILGn5/uxeWTH/AI
Z9/oizYU5xRgyWrXXbnXUSRE7NgxPIfnQlCzZ17YLXTIueeSdmdpqtbHbzA7tixo
2fXZ1GxkPTYStbxF0BQsSRIURtMgVxhNcoly1/XGM44auc13jbWDhvJGNefrlqr/
ymnliQZ9axXoSUfln+N2DVZEIJG2hOstOwu7OW5AOFsBhKSBE5WzFei3ub41J072
locY+rhlpT0mABn/0SB+O6q0rMryC7NJIrVhT6QCQJFWpmuSw0J7vcSHFJVBXvK3
3Dbp5AfRp/geBZGqDdBbBn9heWyjClTbRjEzq342Wobf1TkfiPgx/vCded82ZtV4
q3eb2P4J4VNRYGc16P2odGP7fd5fIPH8PX7GtoOn16rLZFLrPOCCN7eLQweDQzxM
DOZ9ug6iJVSaM0avgeN9EwgSmk6YqO4rhPzBPxklDTtwZRLimXsKmOJuyhnMzglU
IbwVCMdHwb6KPcd5hnTxHKWeBaZxKVP9ZCQqOeF2TWNlVorRd31m8h+aBFT5vTzp
UPym9/L7Yt+q62fciu0O3h7S9dGojMdp7GiJGad8QXxpXse3pQ/J0ocZAWg4QqZr
U3OFpZduy2xLrNjTHv4/OX4AUFEJqeNq9Yc5BMr/RYchivOAMGHU8Y0Nmm77ArSW
TJol08nm9kK4lwiK3bKN2flu8D6CiKGYqnaFeDgDUJv/iNrFJELDNjQ9M64hiui4
QUSPZ9YY8ItPgbl6d993Cz/chxkXQOG4AUzlgCHFlC0vHQvaKtIfemOBlu7wa8lQ
LuW/6iDYo6qWD/dyfZNkPO1SCn2qAQa/24neosR7QoUFtAh4xPAG7lRvrPVZdLqG
XR+NBOz1k5fJG1iuRRLun/miqIoQ5eSgbO8uGortAWKbu+R5sVSiTRu0wEXL/gbQ
d9GPbWK6UNgyzV+s1Q+/qQcuWMlhyd9t1+T+jZAZKB8ymIrz2O0Q8xk4xBN5H87O
EAeRVcPcoWeFrfNzsfKTv3Y+haUYQZFIUlIoZvDAbegWPnwoaPntw3VkTSA1I1Xl
1tnD29Ic29URr3kIf0hg2oaDJ8huS/omIgCYNOdSHgPQh1D4PfFzS7LmA9rNOTOV
tef7t8a82VDC8Zs3gjKrD+hfYhBz6Nhmd7Km1ntwUW2w8Oji+mBQIQXAcu2qBNl+
I+Gv0+iD6f++1e+JXIdw0uHTEHkNGNMH/bdcEeWiG0lSdwYEqE4hMZ2MDLi8Krci
mek+Ad/runfZcPB+86MdS5/VTuomKn83NWouCQFveTIIr+fFI+uuruY3q58iWupi
nN5Gz/QM4pDeyKcauJkQ6UNREM8WQCuVmcJlOZjDmwSxElhCajWzb/ItvaXcnYWx
Qk7IkUZ2m7db0z2fIPCyBdiVIp3HFXe5F+S1nkkwaVqV2Wa8y+aNGX59iMuxkOla
72SpE0ZBgY2XFGtuS5OhtmbCi3HH4B3ITCw7gyU/ap79NS22LzfPilE5FrbHzOCK
b4WfWZHD3tf3olAEG0raS8tAV4j8mqkuok3bsVv/SsxmlCZue1jRNyLZWik6zkdG
yhb0XrlOtGdaBsTRv/T2+fLWOC9517+/E73mSwgr4uppRLU6GlVlMfE2viDwWE+C
24iOcDLlXtNB1l5QBBPM2se5PzvHaZc+xhVYrMlhs/pvb/+QrtpuZKx8GD9CDPNO
pDDOU/n/c5HHHh4+o1nDQAiZxzxemhYSQBTbb0T4ZEtSENDAmIvThkQs+lQtHnZV
bF6LWeS98b8W1xJ3+oglxjnuAZ5vnJ3Pvjx5W30Jn/luoZA+nVnGJ1lcIOIc7eAE
X4HFR/aHGt/mV09wjHskVx+0OdnGOf6xXVvGTnCKI8oG0PICtp1rwiRiioaQQcR/
Hu7WxyW1aar8JpFd41FIi1v0pr8el6A9WFTeJSM4vohUO9NL4PqsUrDh75w9/YgJ
o/1WDq5Uf0D3ZJRdp4Bb7cfwX+fjnx2/u/8p6e2oBNeSg7CMxkWD1jQ+G5pvSU97
nTmX7lxQLHA6rYexcRAGVLzMRUqw79WfrOJ41XxlkMcl1CI26G6IYqJqZFbTlINu
caTXqRvUEYcP+Ju5GPzNBxsDs8rPmfzZ+4k5imdRjKfg/5n4nEPTUml+OL/vueDs
Hh4mK8N9JeSRwb4u2QUPi2AQ/PTRPHIIOsWwKneIwzYdw0g3+qUzHZ9tAp2INN6C
4ol7MFEeLC7CMsD0GErHGN36+vkfvAeXRdVeWQTgzEGMOk8W/jq0k8M8Sl9DlADx
pNqZ2Ryujpy/Y2PLeiZnDulfC4MkEW90WCBOHC7AvU0J8Q6DKzIVZWZ2lSEpAtFa
+8dA18cMnvjM4D5tjiSpMYxWh3Pa8ekWkEg3wTnKNFLS0kZqk1dkfEUEYklkU5dr
JvZ+pl74Iov2wAkNrG2yuVI728MFC7po7Aen76uVhwu/gkssZ2tgIBgZJbHXwNQ6
lCVKBO0GrrCycoMaCwK1/XxbPz+ipGqPpZynDN+cb+CHcWr6yjKF2pc5gv/2KJpT
XgCNxO/DG7Zm9xeemp+itNfblwHaMsFIDkPtN1RI5hkADLBEqnGynNo4vvWmsqMP
DkDDhDaUIkX2HwXXZj0TnOzpNYzYb35PCLu3OiVEZWiqga4AQYVa86DSYnOy+qL9
zG80ZN7RSxXAT8eLZr/qsV8xqnueK6S1F8dyu+ZyzIEbyqc/vf4A9nLiTf04TJKX
em23fr95c4JKwRVEVp4vrt1Nrv1zWmu7SyelxEnjxeh9aojGKuN30pNjmw6RWJgc
VzkBLCm1VRiCZtPAA0MqP/TbaOdC9/M+bls4Pdxmp0SMI6bQ4V7M0bGO1XEDkClk
2DkOmSRQavxxBgdSY1Whk8VvHXNMwzOA5TgssGySndfd76rAXcM+r/p7UC3TC+Bh
TUdTIj5OSuUdbv1VMAB0XJ4bmIFl4s+2ny4C0WnpKznhrRPFyUayJp1AmtAiZ5ry
bfurg8Wbljo7i0zLBSdUSavqF8uxKbSXex0lgVbmRUreN+k7xif74LW9B8fTRvNq
hJgKr7tBdRfYtXEB8K8FpE9prFVluKBgiDozmbInPWj6B4jOhutV/fHQgntv5Xja
/tR9f3Nby5XpOFI08GNLlVeyLDJBakzph86gIcuImMsoyW60/dL0hKmu4l5FGXpl
KVL2kDXkDRzbfkplys3Mftymz2eLluRucOcU2VQ73qR4qCjO75Mx65YYaXxva7hx
jRchrwFRWHaFvjMTsxH8njTTXOcANefd5rF1OfaKVrDIkicGzZK/WgzH0XVq36Cd
/75Abvpb5mhDkwLVWOWskAZ3KlY84u45GBQn8gXdfHoorqraG3zf7+O7y3GZPpMU
CNbIV9R0j4vDeymX/NPbOmdF+D3MvFRNkH1/L8TBOLAPbiPIPpqWgLnkFnE8dD8H
7ZboebV/rPG/Ot2paw/81L9+9vbKdzi2lb+Ug0Y9liyt+n4FGja60u/iwhFcRjIV
mIv8Td61ru8U7ULRaCbmiKG1+yGc+0cLg97q1oxJ4407Bg1VFRvApGL5haSYAIzd
b4WI5+JVcsW4+svWVFg/b1dKJC5CeU/slkw2fFQf/N063KHFqlnZfj+BS6njgisn
m1KsiQ1cPQcs3SM6cGdVACpcNjxBgBoeAwH1B0A8ApyRBbFOwic+iLBkLYWWcatp
icz3AOZ5e6z7rFyTAbY0h0B5dLfZ3SIeqKYKRbP/Zd78KHJ8YpEYr2CwhZafYR2n
77lSpV0tlMp8UG4H57iFV15njy9EqZ6/lkNIjExlUw+vVC0cn9bhUl69GG92FWzn
8bZ8i6gYlh8a0/oMDMkSLmt7dAJFfmIdg5iS+FcSCncrwomi427re7LIrrIgrhNm
4W2rPmk+eDPIr+A6NVIbrTXIbD8+vHSduwqkglus6KS3rqSTaOQXpytkrX1UuuZs
k1TfONbbklzQH6I/3FI8CSG/tWuigTqxASK6OrS+j9phINBZZswH1k32F/JFg5bl
WF5/LjVgq+0bsvRF3v2NTsTD5nu8cZKxlZsmz5csbUI1WIxNLTdtZwJIbrl7rT8b
qeghoTILORz7F/E+oknp4ZgDNpeDM7GaofDc2iocCVAcLYg8AfeKH6m0cYNYXuBg
nH9JMoIgr22Rs1LAI5KX+ihy0NYCjwv+4nSzqQDpsM0Ud7qvOPmn2EzhsGUe90Dg
wWK3DwU+V9gXimveDd20Yfkbvz5Q5YVZi8SeA9+3ldRK3YHUrTl1TIhL+l4sXU+X
Te0D28NKm/+JNYAbCCFRAdP12bzi0JQeCL6qw0AqWZnOUSMkc1YYIvJd1m0TxSmD
f+/NFevyVxINJ6QGnthhHS31vLL/zyqwWAkYeWQrewKC5Qu2HBcauxA1locNy3U7
G/lmo36wneA4Qf371sJENXomlgeN9iYPYJoRY/kWBoI8vy0zf6W9KqI7MYLJgfRv
a/07oDynVdnEbAcfyFEEAg/gFRXomPIV/+FLWoneVmCT0EBNsRzjTYPQGcLFED/2
wx6DfkT6dMRJzcQTgm7c9W4tNPgWtxWgayCEdXlpvtmymwdJ4EauDzWjTdzwlOGw
u/kN3YAj3iRkjOrSTl325OnS7j0P0cCHLwWLIyQ67JaHsBsdWAp/fk4upfA5+T9Z
1mV885XfDCDH8/LL/Kvk7oCwl1BEfzZLOQLYnrByIW350DbJLoprJ4XhK3Sc9+Sp
0rkwKG0saoqsUamSRpn6v6WmRuLzE4MCLtPFVj0XCImbuVCyHBGdBaDimMiNNYDT
YosfH2exag01ca56WQSxPNIb3Uz+x5DBvFP5PwenltpD+yhSpvfLOt4Yf44Ovx+K
Pd4tmjKGh5icAv7moNScnllSgrt6diZCExG5FoHoA9LgTZIsI7+XaYNo6/Y0gcUF
BZd2et6fIM3LxKOu9gWPnGM2dVDUsPVbcoZWSGjmbAtP3Pp2AF/aXZutSfjQ8ck0
pB6V7SW+3TFJacDuVYgqgDnH2XeuxMNRELZS5hLK2H8g981Z1BmHVxdlUu4Nd4vM
aBs2RWJDwr+qcu+D3X8DXTHlJoi+oUMVtgO/QXxuR6co/vIO8fWagp0SRQUQmxb5
n9CQLHFbDPyPmhDC/SwM25FhtFepzrAWwOUSutVNB36dJb/xBkmarjDhrHS0s3p3
MBAxntUnDgxnUjcRtMwDS766IaBjpBCTwoZt0ssASKrwjmGvvbJK1FjZX4Xk5foj
6VNfwXvASHxY9mWWtM9Px2YCTwy6WxUsnes2KkzwdXCMPEEEjbEkEASYQtfzjjC/
CezEQFgpcsB3el+oTsA6Vkof0vv/q9lJZa8gK8G88GXOmvPPGFrM9KDMHp09U+KJ
YL/CwdLftMBTn+GVG0SeE9PS3OLz8mEO0xGYhiYJpjl8AXDvBGUNaqvyloqnvE0F
vLq844znwn/YXisAUNnJvW38RJTbmIX+AWc3gny9tex8E55/BZqm5Smr0lh2ikJv
Arqs2EikfdZbQvX9Gzik64/iZ8Jtv9VPRF6/nkPkfV2x0BVguek+sPl9+SvSr12j
/w4DQLdPzEiAYANoi7PVczyIaQU2SsaSlzwxhiJ7gaHbQMI14dkNsEM7iIkZV5+G
A1Q1qCSkcq6L9P7zP0cfFLQTV+Glpfg2huzLzA+YuzWOqFMe7zHXAsCMbNschi2U
38wFgRw/M3fvv9av5/0mWkoPHXjs9Xy8gU7RVeeQxYZxfa9VWpd1JRuHrU9Hdh/Q
+IfxjPvGSyO0B9Jxg279fWuX3revFsoj6YfhsdCh7j3RAveZKoDA8kClZ2KVpkRU
78Fagv0IpDZ0/kZhoC5sKcocZBVMd0QC7xLeVc8j0RhMIBnTGIhy/8JGQgXAsVcU
i7qDt6dMvMx0HgmKlkh2FFaMCGvvJrCwZ9wSDDd6lORHOgD60JUfEjF4VAQH+hrZ
+Tp4QSF9DnjQNHb5SSFfEjd8TX5Y4Zb/oZh5Zn8Z0qNEWqFsgFSdgn89nvskXI5T
UClf1DZzgQ8S8hIDJrdCisdpYpQQ2qwOg5J8My+hWkdRdZMnmfvjei5EE0WrsYyG
v9AcVW9xf7rsJvockNfqnncO4IafL0gCz3KoeW3zJN8jJzOGQ32V+HOOwNCUMdr1
vjH/DuR63RfsVnyrBeLRpjSYsWtG1O8JQlgmTaebwvxvkVqnV81EkCvxlNdpQaFn
R00aUuEDusF3LRVziyNvGCBjZV4Zp7OnNjcNBWEEqUq3hXJtLc1OjKQnBeraFLPY
nR8Kz2QFuFjlUrCRW/1fHKwgQpTgcp6fyOgoy6bSqqtTwgVRFU2is0SuH5mVfzR7
mC5ih7AoaS7EgXXfH7s4qhqXWsCmf2SdJEpjNepnWPq0Wh3/5aKP93/kz+KjHObj
7ixuV6zN5fd9IV6LsWBm5N3sc3Tm4YJw5CCTS/vSd0m8ffhTHwNNw6v7Nmuutd+8
BtcLPha3+CuGnAtFAd6A0Pb2/h0A1laqgJr9YIc0deMipTjDWwxOOWYvxwtxGsy7
xlSQ+31xOxNvcaqe5P2dfIwpNn55VTsKNXwsxpyemt9m+T1P0VqMwoGyT7Qqt0iE
Z1JN3+NST2aruCO3P7zoj0m9hFPGn9mjIg1vk+h7Gd488rC49YuKiUbyKoLuLKMm
TCAimWN4y+VkRXnCdDsenHO2KEf1Jklqf5wJ2SbBnfRMNSzYD7MVyguBAdJp5UJU
ftlsomqGfnAzVgf0k2ETidskDbw2eAUVjn/BTjWGHItMNmlFS3og2Z6T90wGyWW9
n8Cbs7O78A5rUape24Vl0s+39H51mw6QHSv3gN9P8mVTvWESOvE+67kEG04tkKOl
VU+750HDMzhe3GRBv85mDsEQQlXIcXy6kfeoswhD+U7ztuk3DrxwdX9kutg5a0/J
mvG/kePTvI3xY3WFJqWGxvwPSBAVqXVacvOM4o5/E3Jv9XP3O2nnSTkmwWu2xcMn
xHUokgpKYbDwHgApvLjsTmA4b7wdvA21moYPCkkFifK/9pO0KPBV8d6cveSBtAzm
MxNR3P9MUT+hX36xPYXui1+HGXbivGFUw9w7XltKEm1krrolcCZpjiRRnE2sxFXI
udUGDEkpywVnMEZLYayE0jrszGPCyUfzL3P4ZJeHGobFzQ/JzVrrALxPOgXM2e2I
WWidKfchBi5kWyv3VntyVxy0ptKjp7AB9sg4Tmt1c9GHfGzGyJCWe+XJvUnTmEpZ
SwFT9SxL1y/E8uVRsnNPeqqOuo9zL/70Ty8mGzGZl4UwHZZTCv3pE1eR+IY7AztW
Cnonf0mlx539oDPnk/o8XJ7yoKh72uNERIJe84lhG2Dm+1k2plAFhZG+Ld0PpnGN
9NPxJ2b7hB0S/cEkKxtBvbtalhzcdu0OCd/IJPYRTspxN85CvlUukdCFVjZ3ROO2
EasV/UK9NcuT6s5FT5siiHbfAoX1QfYFl0x70NRdZ/3oMF5pVoJ5C47IwesOLoqB
8lgHQaSzMIF04ItlqJbt2xx0D2M6Vhctxb+FNyjtyIcCraC9fibIZDGT6AMkwBlI
uOqc28Zw7QzVj1vACIkTynnFqsspASYiOVaW494QHJm9VTy7wcEC/u1fErRlOHvX
GuqeOuepeQnUUmQFxhJgDCR3HvuT+9Mkt76dO77nCdkJHojRm8mLfc04OOpo+HjN
GPx9pgDrNeJtrsuKimwFDDAdPQn4oOuYHJubnm3VnmMJFFl0lo9ApHuhjzho1Rq9
o8dv9M1h8uW5kqpZjQ+R59n0Pm/xpA459LtTdfOw9Ybg3C73bvGdqglLhJyC1VF8
EdzLQttwxKqEQ37x2GPGNMjg/wlRGEGB4MN3eWPXAYmKVDP1a6FuS6I1UQs0VLzp
MlleeBmFKsvmKu1kNkZBI9Eek7pMEfzBKaLQbfT5qzB+Os7p/YkoEDPYpiun2Lfm
nptHmajcWmTS+cwCEqScjd8tUMngx5NdQROI1OZJRDgWwq5bq0GtZS2iHVgBVIs9
8vabxnZdBmxVPq5FHLZjwszITFbWxzv9KJAZ/1C3Gck2NLxdpNklKl+DHVra1bd2
wbNPSGeLljxn3z+LZIoh5eJs3Y3T0sFsOnN307bdkBxIrjCYjEODRYbL4hTqs7yM
umaCUxgIWX+QestbdDqOTXTfNCF2K3t2WfkETRgzFHgEfUMYF+b96xr3gkQXQxXV
vutvQh+E7K6aeByLO0k3s7KLilsgL4aqhfm34KAxz3TckEQ9TUocrFN1YRgzUZMH
lRwuZdihxOog3s4+I6WFc2Dr50ChRL4OACxiddSPCqYZzj3zIG6bu9EN3hbVQz+h
PGeckftSKJIrWrs/3JSjUeb60nc/Me2cP2JZh9dimV/C09I5+KoW64vKUtaWtnkC
zZSAAnqZX3sdXrm3fjuXSdEuc0ErD1FPuMNN6YVf4rOlFVuyEz5RmE5apBvbmYRx
TWXCyoKI4BnTrGLsWZChiRcoLdmm7ZxDPVJnhdLNmBRXSZvhEsRRf+kEMJm/f1Ot
k689PV7L1GirV3Um4jH7QfcOK+kQRV3axxf2WrBHIQcERWFro3fKYuvU38h6qwkO
RnF8hrx/aURIa5AhBUYfK9XUbYPxAFSZVWTSDmEcTJUZMCRw6KJ73UXih2T5iJxa
MyY8G2skgmxn0kvmruo/77x7TmTKGhFe4BrgauTGKWZO17IeJ6MO/pZsOQd6Tfa/
VorM1H/UXU3BIuBJJ101xdxKwWs76c5VEBDYS5Ik0RH0arTq9RbG9727Pz7YFt3q
L8wprDfvlA65MRGaMrxVOiCf0DPoPebUTYUj2Ziv3n6ShTElfFMcDIWtk9CLbChC
3pIZg8lAHI4LT6iU7ZnLsWoq2r7kwOzPn6d+QXw3U6NNubyb8Akdof0fgeMqkt4a
2XpsBqE1/mqc2ZlRQv6SeKprPjPrfRnC3jFsd16rSx+Wy4L3eNgpgj247sVu5tnf
Uk3EIl5evc3Eo4FhFlKG058d28cM1PVDs52Xez7sg3/3LSgfEO6Y+KsLqlfeAOK9
jWv4BjXNhLQiLOjqgxYMib8GM46eZUnnw5sy2r/ttC9hCJf5KZ7v14cn4q5jx5Ue
epHHZt1ZlwbRDpdjZdT2k/sP4HKQA3ivEiCO8WXVbDCNj2dGVBGNLV1ynCMdWDuB
HBrkncbe4P+XDs2l3n3bq53R8x4z+3V5KFkO5LKgIZBTymkLw8EZtnrnAUXa05Nt
8bRpcAA/pMxbA++tKb+teIDwHmifw1sFdaSzyRCBgeTUgiVEuDLcjuSMA4HCFAnb
8A2NMbIIKGz05RGBqlb3E0IdBcL4hDgUo9jYNR3YA8LTKiMh2j8q3SYrfCdUsK7y
vNPM4l+qFmHGbwMeM+T5Tn/VqMbwhTEhyV1s6FjBFkzpinFq7yRLoLPwPUDpAbae
P0WCjN5Fscxo3umS3ISVCEZHxNn6lLx/Mp9VAsPUwTeECjWw0VgxTnP07tTR1e0Z
/isqmyRuh1/aHu2hbrfjNaIEP8rzV8oNnsf14ID5h8UD04D4HbrDhq5Ns4m6CWDI
rIzXleI5RQ0zfwmx8DeGqyY+1HQR29Sv12GMqlvm9+zt4hI8OBNzE82D+riwU2Av
NEDi9R1VrZ9n9xayrCLDLcCXxOE0cJ3YMj35yHZCqP3xtendnZWytyK0Kasz45EM
pNrkTGnku7yhzMZQxqaEg2yA8yPGGP0+bDBn1GH/U9blBHop81GOMR/wLkEhvIJi
soUtcj0lwe6l6AvCFuSgvDBRs+oSBXBOdAaNQ+8qlCAvG243H/89apCa8AugUKqi
vVRRTKcelHqY35TgN8gz4VeFd3vZkj37jA1Jiu0+Myu7OjnxYu0I23KwImoPrBz8
SQl57X8Z3P3Gp14EUwrWL9fUfrA4L1eJGphSjfp/L9fdxZEZM2G/ixlh5u1QtMbc
/px5719AypZPsUSczv1tmKIJJSTbfRGDuPTWrHsU68HKAp3dZlXSdndP+ZLqV4hE
XyWZoI09FKV1os77/EZgd3ua4JPuUvkwGIPKe8EuNE4qPbcXt248vVrewVHkKenC
fYGMy/WDCD2Yahm12ESeokxfWQp5oyD7HF71f4eQ7LmIAZI3I1H/wUW8BiY+M3/C
a1janEqAdDQ6Y2vGAiI1z+TF8khPRncO0L+IXLSgNj5gogV8Znjh2/Ufwp2WUNSh
293UpW4c3JTw1wSK8AE1SzOUl3Jx/Ui9+lrmdhfDow3doQPdd+YOOSwJQdFvT3eI
XF/w9XLDtsCrBQq29tgM/0HtOIUIyNP/IC+s8MpXFm9g6pFhmcBzRlD5+yMaVYjo
gjB02NkuqL4zVgQXsLZVUwXY95eHZyY5V6+VQhUaLM6A2Fd/aQBqODnHKNor0Pl0
xK92OD/7Hk8OxmXusHIAWJ4N/8CM1DZaY9Wb5bVM5DkItrzaDrYTGXBrHsEMIt5P
Lm7RV+Zf0rctsutxp38QQ3+NVSeWPfA+n8+4H6X646OrDAnbmInrg8VdyO8KIiH6
D3fkd+qoqqGS9iR5bfyXP1nb6ao3YK5DUu5BQSs57dwzVs2xUIVYOhdGr1HQq8uq
NHarkCjpNl288ZCliAmn2Nxrizm8DjQiw449av2RYfMisj6Vuch9d1lzQPox/XAh
KMi2R8wXbKzxB9eF2rTlp7eLI45dGr8E6UySXGAwupbA8p8EIpu38ao0ZhhmMbHw
yTk1H3XeTkiCGejEgpZ/ShPTDsVq/A7G9D52v64tUpEswHT8MgNZWwJOqrC0FpKX
nwj06bpwX7mW54lZGdIanjtojX+sH1YCcY0U7Ift1NtFBo35JPPzcsnZbKVzFZQe
JrnoJaOKFjprf2Z7HAG6w5gZ4xWdgyF5ojpHHoTsemulROQA8XuzhYuEOxXccJOI
M7Lv8oP1zczSxie/eu9Pdz48XGjd338PaF5WtJbusNKb0qg6aFmslXpYQayAxOPS
HEG26lbrxvby/aEo35vMfLc11BoORpZOXMHSbXp/qzLAwO/VpardtdBz1jzftkLu
w1e2nj8kWtrBJEZXIYT3aFra8FJDUvaNt0TJThyC2Q9TL/Lvnww2/K3k6c+uk+o/
sUESi+0DBRGWOTLeLxWspY2J8bGjSQ7MqQG/jPvc3R5J2d0K+YORpm3xZ9ZrJhXI
d1vAtIC/PLwuWXiB0ZZ0UQwnxM2SfV74rMYybTSFTIwRZ4they1epQ/UK4UTJe82
YPZbaQV3RlXCY6D7aFysreZnlzghiE48/qkIIpJlbMcsxGE2sFJFaT3kTG8DiQtf
P5/W8coJx+buAaWxgyVkeNu+ZdCItsxGMdppR0qym9RQVj2Z+1Rtz/y9hTZ4HPz/
QXOcI3HENqyQ/0DAq7oA3NO0VINm56wHmmW825tdroR5rrFCr7ob4owkCVjp2+wH
B9RQdw21w4S48ps0Oj/BBxNBSU4O0ygGC8a0X6BeulZefGH90gmxsWm0jjTw2u+f
R6bc0cWlwjTcpjycEQrNPOS+halT/jFuPVG1TalU/66OtA8irHJ0ExZD2RzodPz7
vkMLyjRjnSMujqN2uJRkDeqAEH2o0XMLJPBaR6SH3n910MPk1VA5nSVM9A3jpFPj
rgrNLRnkISydN/2HaSJZEgaoiS9zmK//VufUlIniITD0YWH2i3VHCv5L6YeiT/sO
JkKTWqWrutHpz5VeuUp1N3s04H67PYBvYgdQqVQ014IdNr2D0mpumYJ/n1QgiQMe
MsnrqHZXgXKw4WLCTVu9TLQnD8GhvD7yIzbbMjalE6uXVrnNDbtphW5VFL12kw6K
KUSv80L4mtR8Gs70LBmsNVULcmVIu2JPbtgSMGAUuy40DU+UsFtuGH1RgHM4QQX5
Ha05M1z2fESJt/C5+0qsmWENVRGnps4vI3frWeOL/dSlghspNrGABXK0w9MUbxEu
Mtd1uBRbBu0bF0jLBhTErU3s/RfxzYXufvfXMepQm79OLsv6EFSGe9pALcMoGmJ2
EqLqu8lP5OdLj4zEo9ZCaGdILLq2aHAXxcvAjJvQBVOj2bqXRdP5uD5MylPq+ZZX
j4cd45D9h7gnTNGi7a92Cn5N1nZsET6ngU8Su2uVv24v8IgOLOG/IXujTFZvsvR5
tgOknSyDFF9WLFtJ9fErxkNwU0cRqxVEobYqsFsYJA69OXBd8MDZkAmsj+CLX430
ihbSbzrMhSQbHt3Bi47arE+yOIH4OnF6JBbr5qAom/02+ul+qGFm8gkiJvWcrvku
KMwku9Zsf6frpvNN5sRH/FknFU+ApZsImrpRlwflDnLi1Ga24ZvCeCW6WbnOxTeM
1n/pAYhlIKdXWZ33PlSgLGn5w2gNvMB5HBiehBuR/fcURPHRpCNq/L4ijmRMLfxg
W/wO9zv0g6ps4mgs+KBPpkD/2LAGr/GnAX9Y8XdUMPb7IqoRRZ75NY2gLgD+gtgn
S04vTLZtljfs4Z7t5+Ly44HNdr21HHTJyfL98r6VYtKAntR1RxMK7aqCGN1nPmHh
6dJBlgyhbt8JHpO1b1TvPPq+HjTBfNLT0DQaoM6Mn24vm8WIoktvhhrgqYLZVSvX
j73/6gXU/19uhSgVrJ/8EclpK7Mcjh4c1qfyfxNU2dxhhK8boCwjgyrk0leOfQ/w
WhIyUIQFVUsLddPfHlA6CG1RHzZ1UZgB/PFnOU+4eo3HRhF6Ocg5vGZoXkX5QI6N
QfDFp+x6Ajo5ZDhSoXIuxMbPRNnSpkFMQEsHiowZLJxB8MZFSvDPhozDpOhyfzAe
Yxsf79M9Epn42RMNKhvbnSdoAiEXDW+DW1ia3m31FyOAFCuNiCP2DAP6b15HGovW
H+h6s3PTxzGWZtlo9NjzM6BMNx+HNNW9pHCErYhlXkG5qwMjECGYHUx6+wM7UiML
Mh60/aVRjUc9f0GQldioeNGsYgdWHjHmqiSOCk62TytU6pRhdStwHJGEAyhEUrO+
x5xNd2Q0Sk7g3k1Jp3zvlcS0ojZpOzajjkh/0DQrMKq2P7LYDuI7kuqvqwXfRf4M
XdnbPqDug24ZNvfuvL0hnZXaxF8xClqY8KNrdMsPZg1xr92VwGlY5tDdKOlPnzMM
Lqh0+NT23A2T5KDqH+9cn3wkQ7rnrvwnH7tRyhi+0RNWq3GieH4AeZl+1UStRZVA
coJZOg/+9g0uGk+T16s1YF/n6onlCm/zPBvn4fXbG39RZ3/NeU27PbT73mi+umLz
ciLzqGAoMTkYMyxVWdo1YQg0VYwmxzhBzEi5Ei1MAavOkMxAes5HbqR1X7jvMMAA
sJsgdPnNXxcqBLognMpGpK26wLabyv4IkLgSMuE0gn6Gm1vpJ9vreLKtic0aFMBy
Q8Mm+NMCjLXd8vG6+56m5zsczF/hgMSuUvPpKoOBxeCgfNfXoOgNBJnwen9ISnVo
S36AwyUge+ebdgvb5YhVIuk2ABqw27OCmy31vsjSm8uFHJaq90YKX0BLJOpv1QTw
zDs55FPLM49x2/AeQxlvAK+qmIdEbCPzclKU8Dy4/rEl84uuoR4bfPwp/1mSrQ5e
85egGtavSPjgVjn/Hlm+1Oq4yN6cFprVSd0YShf5/wgbdkXdKF+bIqb6OXdvYK1P
xSZgw/Wjue8JRb1MRJ0OK1eyDMY6yCbvI6u37lcPYXH3gUcTNPv2vTDhzVkpprAo
ld+AOMtGz3n89HSwiUliFk8vx70682q206/asY2QR5AcOgAfuQvEydxEnpHuMaCQ
uKIw6wPYN1OLCTU42pEMsRz70nDsI1DGkHmr1uYb+UBe9PbACYJjCVVS08W2wCAg
l5vR3znKbRRO2DVmrSLjHGj7VOWU8i9kLkXyN1qk9396I2jGoBmHhV/E/UBX3kag
spP9Exqg5JhQSw8a4TpiUJBybFd7U+zj7k34NgeRGUjwgO5ArLfmCX3SS3aNRTR9
mrzGHRkeLNAxsc50p0IqCBHs34oEM3jfbtEcYGgnyEh4AV2bAi3rj7jjRro+4GIS
N0YNraqQiWtHdbBigf74qKo2yQ2JNmTKr/p9tSsmAVQVZPlur0ybVvogJdBtIRaI
cBgqebcUMV1mcpNF0PhoupvLSJyPCmIbCDsnnQTzJukFxV753AIR5tWoIHgB29BJ
kIcdINGLUnNNvPo5qhgV/0A8NzqC9x++PVuj58UXdBoscxrDyrqg9ZnwAEysLXqG
S63BFVAo19VLesHnPPjA4QW+PWKpWZZPDYCdO8OoMl4gEkfX3XyCm8rbsBU4B14B
dCUlneX8nCp7Rl+yUIX0MV3rFkrEBh+QlVHhl/T4ykp6E4jHczgQ0V7ad7bbdl/2
l2r3SNoAfHNjZwtQUWJYlpsX/q5JgcGcH4d99TmesRG46iObHKMnMqYFWABjIuii
eEjA77ep4avKdRXOkIvae4hmhYNSUkN2Qn/CzD+1+Qpu7v+ZQ1s56IZWSiKL4iaC
KiA+jQ282bvbhE5MJaX4Di2NccGPXMfxRkKwQFuXJNktrhTyECqHPgTIGJRna6Sl
sVNkf3hJc+KWItzv84iZjXqU9mG9xVAL4NEF/9tBaDPj4CXPCIbT277asJ7CyKpL
/9Z0cp+P/NyVA855pjX23Vw8pplmCTCOPK6meniROt3yhjKHp1kzuEwW4ghtVCQn
PPdTCKXe1RsN7jpAgA4FzZuTAToP5yCCVTrV7JCh7lVSbCCj09eQ7Tt11UkYqL/N
Ub1FnWF3AahU3bNrp5USpxA/IKSSw5MZyv3ENKn/OgtQYNBo3YhqIv8FIzfZGFfg
Hpg/7kaYMNxBhthA95dKlKwQljAFAqYbxlbKZ1THQpS+4pb8KI+HXT3C0vEmd1VM
KIBl8pBfkpTdrV8krvTYc5qtnBCiNoAihSyGA3nXPS8rmeXcpHj1Q0TjRGnMZ0C3
BZzvF0LCn0R5oS/0UYlea05zXW7wiPoiENvNffy93Q24oTCXiu0f2agOnCgDlr/w
Oc78Uh1qtF9jskfKi53nkj1PELUIGVdlJ7f6eY1KKqyeSGEWyxRzKjrtCCx1ayhD
Q+GD3HmWQMVqx/S+CBaZnrrAwNEx6xkSrNfvXDw4nOkOPrLZIBQkylc1eGwvGrjo
dHsb59cs5dVw96g2yk2BLkTaFImmf8WKR6SyibwkGtBRzJ/qvTUuDaD+cwFJnTVw
cYND6POefyDcjBY9bT4oZw9D7cb/VCfqs6LzhgKtgYpMZVPGC9HWyEcLxD9aA7p+
BvmAYevY1oGeaSsTIOnGhoJTu+BbdmRneVj/rLqxYMwHjnM36ZZhOs3NgWEVAMYD
kFoHLCIFyJnm6LQzdeca/u2o1q2kFtLPse2bYojNnWv+025D7bcHBjdilmhE5En6
ZeCxIrqiyeEjDdzkrxP7KCItMMwfAtKKoezgaSSnVkB8uwqtU4KYN6vY4NBJY3Ro
AwLlDTmp+RXgOoULKnGqoV+V9Pc7wvdOxu87bhcstVVjYK02qNMsONi7RlcNgBN8
0W22UtFzruQpiFHg91nU0vOjojcApKZFxQYb5Km/Ud2fFBCMO75JfdIbRBptz5XS
6yKLnCjPfyHWEOx5B0+fbUJ1LXABuamAbjSAFSSePq/E0vEe8PvMzP/T5RWHmIEi
cL9Sc/gfcvpR7NEPzzGQDuIPsH8wTYb+DX7Wuw96KKBHAVoZNc5OkelAy52GAroi
Lqd0SUcdIftRGsvaxvwJ4aC3QSf8mrb02tNWPQljTrJ1xiaQcHMUrozy2d23SRsR
VOhCR5JJmHmwGorqwYXJxRrUBoFEEBW5iKzR1jr2MIFZGxx269ubUh8m8SC9yWwp
lsie1usNlfw8cpKr3ay17s56UUwGQUUzfbaum6ktZOegzICytog5Enlc5P3cp2uV
Va2bZJaB8wr9hG3MFKb+AkK8lMEej6Gqd88pkkMIv1loK77JtOI4adzWnvZedrSB
XxjGd5njvwpNjKAzCoZah3mGBlUGDpPuEh02/1MMwwq5iaFd9OPaNxuEsE8rwxP7
zap2SWQp1opdnSxqbY68PteaOEvENnhlfXeQsQAnyeG7UEz8t7/6lirFpRQbCO//
T9j/sYZuaFdNxp+0V4eNi1oJhD04HFM8KVeyoeDz7hvEDGMH0PD+hNMIajhdwNZ4
15PT0frqcSNkotWgk2wTCtl0kIOI4uL10caGtLn2fvNj7K+8xEPZGO20P9SCn+gT
mYVTRGnPleFRhRCBW1ntsTLrJAZ70zQohwS11PUkL9lmTTfmCvfHmrcofWEmbnlC
eQ8jviq7oNav/xtOpCdPaXcGCdRe/sBjgombCAUpER0KKDcQYhq6NafF6ReoSD6N
PI+cRKL3jXMAw2wEz6hCfgJzD/DV0WUeOCQ2iu7+WC4zplZBUcuuDi84DdvaiTD8
VCr+IchLbRVv8eja4TC8LSUeVB/U8qWLI68yJiYUOQ2rD+lVpYp7ouSSnW0zgqBj
cldTulGPdFJpav3reweVlG4Z1ExnJsd7eoB78/X554xBdK/o7pCU6ZxfxqlgCo60
FtYlAkXb4qX6RXGxNaF6r6Y1e8G8I3XeMzgPBHuvbTI4zIPt5dMa/TvpqPoD11nY
I15z9RqBYllTjBzfj8foFnGj04zcPzPE4qZgdEg0GW/sHeoAnCW5Upc1ZLyyW1iD
pyaEQuj4WcLi+AFdKnNbBULTYrNXu7zRipscwAhPHXI5d5/8oOipt0snC3PboIkI
wgHLkmISE0meS5vLJjMo4y5+gLhI5U1wAW5PJeuj76+stPOEVk++4hEqPoAbnU+h
OvN95lNTHNJReSYW60waiIVY2DxtSKQZM4xux3aD2H0+I3WjN28ErxxyPDfxZaOv
S8gzdjbCYLy27bMr7jkH0vYy+ToWH+Tdy0RviQp5tLbeIchvyRLSoUYv/OgbZMPw
pvCEHb0H8EqKpCQeWlkj4jGrNutah0EcO4RsuEJjIWP++pzmgzRHUbXQFDDllQ+b
ut84Ws5yD9CwEtNBFbJetydez2PUm9syManhTEcp8iZfpzq9kAJGQgNfs/A8pO4Y
lmDoL40ACA0dOiTcI6qOPbR3fXkbVwSVmSAGsdni0eSer/0BucKE4FFshWKCX/mg
5X1B/k0RCZOnKwJIJuOcNADnRxlmwn8hRraM/7EG51w7Rkgj0Eg1FLJx9P9trefV
A4HaiUQzv9k6FEPoUKxLp0gZNgqM2X2HUaKMiMH2I95SXjQzDiVTrGT9pLrms8ED
OKYbgPEeVFCnF9KS7CVHziBJuHAs2x7Zp5fU2j/3wF0ZfQVDlWmybo4MzXtUBgPu
HTwefUDcMo0y8zrBBW/D6OQSqV08CuANKXpcq0iPTCsbvjGqdhcailhRTCHz49Ih
AVC7XAjK1CEYZrexV5GamouW/1sWhzZZ1wyFM6YaeyXAbNY71C3Pshgt7/sGDcaz
QORIVPQhscWdo+PPfC60P5ewQD/wXtYjtfc1lz/0I+KTQMJSHr8P4yFBycaCDops
CPKofeyCSJ88GvZWGY3/5mz298tjUROLm1R9mtXbD39I2DsJxffnachuTDwVvgSe
Tfo/WeMKnFh3ZDMCtmvcj0fIh45mkJEPvn/PqVPl0ClV6DHWk0HsTXPvF9zVjoWI
gzUddSQWjR0SBPu/Z2gIgAYf2iPKYjQ/me+URFaOEZENzMcy/k5z+4WYqBttSr1s
7sQ/lo19Ym9BIECqxSv11YbmYATCMv7Ww4g19bdqizaxsqYshyCPEGu3ulEeYW/o
NmNPyTPCFPn20KM/IoNqYfAVN40B7JWM3OZOm0v6Gk7WHPD0+7EXztqmZZ0z2Zaz
Kc+wMo2KG/mFAwB3eOr4Vwd5O4s7L5Q+xiY1BB/lB7b23nFaflUjHG1acd7PL0Lx
bmir9seAFsf2vrPtoYd26AB3OlgiS3xOlDN/f5UweNirqqgSEYNmVNRksKWP9H1Q
hAPSzsVDnq8rkAgCEXJDdI3Xo5vCYouw+TGsZqH6U9zMG+yznMIq9b/M0Q1qWzaP
8Nbs6ewBv9EvDW0tQpBpZ5mi9n+T4c6ERQNyLCR3glpU5NKS9QWNmKgfWVDO8Fdk
j1gST5/uZ9L9IZT49gZMaUlfasLcjabAxjnWQqNFSO+0WkWGOTXwmrgE5TyOfPFw
re8W04B2RZbD7twOjBAftJNKaz+sAfq5vNClKwdIbFvRkwdvyzXe8uVdUmEtOcDd
vqm3L/mJygzPG8dazmHYDT/sn+xth1ZJjLocryJ4PpHlgvjLxSbvNHky3IR9dXBt
sM21Kpc3ut7EB/WYchc++5LrgNnfkUb6ZzRtd/gd51ZtXR67qgjdA4I2gpLeGsol
dV80qMXv5R6Fyoju3CQ+B9sBLUOidNg3IjrRSkiJ4yjM/kCZ+qoHegPG5980G/F8
Ew6+wS529KJ/U1TPpg+EUdtai3mb8HkrrLPptLD28s+cRBBoJTH6kxYEkhgO8Z1z
m29PlT7mnE1q5pQ5yMcKpvZ9owxw3stDz3pD/SD2p4vwCfUU0WUYsJjeCLXfbTeG
g3qxa4UDbMqvChjrTzUtATVPRQluohxPsgy4ngjoo0owIka2V4SmVxp58gWh7kWA
NE4tqZj+cn3PQDNH7FkWvg9bObt5JpUNCUq7FmRheV8btNQfZQ8yyjVvbfxc6ryT
UWR24+ES7AdEVCouMKCkCP4yzM8hEcPVZJlKu88d37MxAk0oatE8md+F742B/KIY
ojrjcE4fWAFTZ8svpygEaxiRH3Yz326I4Jv770RjpwQUhTsfEf5nb9tYy4nO3gUs
78oaHH5l5GDKh+IvchTnVf/hNmDSN/ReMpI3Rx+WQyoPeou5rzGrnpiHdus3j2M7
IBXcULVdRjeMFHWve31/GzsMeLhjHvoqWDmCdT/Of43U2lTK7L8UZEEa6fyEf4AE
pGiN3xI7XST07NEsw6qRthjTiJ3XuGQMjsdx4rEG9PC9eiOrCah+R4hLxCln7u6Z
bsU4obId3R9oVRO3nFXWTj7Fop2g8ZUz6Xm06wrFlvPu8sc4kiJo5lXCptvC+C2b
EPrIjdopGy5v9/TPTYqTok4MTveluQ49ixOPA8+S1GOiOkjRTjY3IqfI4/r0rrXs
Zec+uJm2DbOn+czmdpSjS4V2THPa/Ov272TbYLYzG8aHSJ5H9IJB8DpO/9spmaKW
6JrYmTX1m9A0/vyFiKx4EWdggxMYddsHrTx4YJIYQ+IyKH0rH6z8PsEOouPA7KSb
QssW+SMy/hnZsxHIASdh8nd3MgD0tHnb92AL+p3sAMptLueyUn2lRcdLCeSaeYyN
7FPsRE0tLj1+EZHNzTVEuRFntN/ip3RY9r65ZCYJ2Qe8b2T5U3HTuKtbVhFjfpFB
v2AjIvw505jAyZaSxpJAaNRfqUwDtx0vZhaUnEyKWqGS1ZHhQSxMXodYIBXCaZfA
G0pDGI2CLxBOh02tBM954vzOr6IxgXJaPhBIOqIV3LTBC16whugoQxxSj+S1hU9D
eihCcuQi5Nm1l+Z4xKmGdljRfIjegjwYClEQSMpBiZZsuA3AlXtgV3pupIZo/9TE
FjBEo08b83iogs07TQwzzuIf6lWIaQZWkqBQK7x0LVeIiR8mfLEWVqxS+hm8Tvsb
gUUPx5G+Lx+dqlOW2qVL+HsKs7OTs3qBrVYKEmTxBCLhquJy01BSb6trKd7wpcS0
9b6umdBMDqKk9urAXgviWAfaIOXKXTNgTHjdFsNcF0b9G5l56fNvGHW6m8Rq4sxm
Uzz1LEOyBtqSI9EMnsQdkdYS6PPEYRYWWmC0owZppM967qP8VVWPLnte86GfnYwD
5JF+/dx6oPdaQWIgSzLOI61HDytbJhslu7xP6SLSjurri3VNlfB5QPoqv3ZmzQuA
lM7rM0W38jppF9OSUnslObenAHjcn7IxIpwE3YQJPDUxV+VivJ2XkNT72rclHibP
JhH54kuXFtqPE8eq6g5eOcYd7nYZ5yHw7M4y2/BU+9Ltwt+9h3tzQf6rRjcsa95S
rdgeDFRUK4uq3yYmdGw00vLRf468VYqEhYyVvS01ALhmjHUFugLvdYIEXjstvsvk
9Ecz8TiZlRwdunJEMITxwWErkBbzWFczdppSgFYJm3JyniFZIsQgPt9aFw8df/C3
EzYb2fLaCKCVm6T4iAcewDYFjLvKHClYLOxGOXdWeWIpaOkTpvVRFYJ481Kduzx2
vZH9k1ijD6OCYYxUdnbfAA2CNhQ8he/7sD1NWxta+AH9mgGZiMsU0hj5wa3Ol0xG
L8zzhOVhDYgOc4zoFtGRXRENyfrKd40XITU/7650tVhTop33ZW0KG2Tq44HMVcUw
vvAxgCraxuHiPO1ovGXxrUhWtLCJHtMBYYzwJr923yLJnRJPqw2qRs+daG42hAtM
+GKUDgmd5x4b2Ed5sKnA3vIu+f40u7hoGu9SdgwVIHbhzuhcperpZPvoNFgTxQi0
oLh6D+s2Gpxn3zr5iLZSgU7/EVsLYzpgKoC9hbtUTvIcMuHh3CrdAnD8ZTk2N2OM
udHCR39VPUFfWiMrNK5b5721eyy6bXf497yCUpHQxCxVwcfsh2zSC9byFGB0+9lG
Qk9x5Ki2eRAtDibJoB06+C2zsAemG4rVOmUonWHouWoK36e3TPY1hHsfHwR9f0mX
DQVU0fy5M5jP6fo1XADTP1tEaKpfVL3kh9EqlqrYFohtPIv/5QQoZ5viluInlQUq
MHUaPGFsOAyIYIHR9o4bLG62v0YGZ0FClEfuJJx39Fumz+9pfD0pP6LMzj++a8Q9
p2VpkrGAq+mDnm7oof6d/J+eko3iiKt8Luralc22l5RHrr7H54klBcyQIKIQTO0X
TC746qQdg0+5Ig8KqZ1fW5JueJApPiPZTcnEAza9p8wwwoTRAvIPQsGAevV8kw7v
oSV4YNi6BGAHTRRshsSz+0aYwl1HF3M+BNXXYT6sGMB28PXT9c8m84ye0pJMGgDm
eFQg6J4FQIVFkL2/7wRarZ7L7uB7JCTbAXlNYUdIXTdJHVqFWC1WV+xIinbIcRaA
hbyB3Gr7tNQ1r7kbRiI03VXr9Y+/emYhdRZ2xC3IBVXZsIQGk8FIjPDoKyKnIVoA
giRAiIejcSxU7ZwJTonUVErI0rBP0HHOCSyLvvhR2IpjdFU+XnGKkOOD7CDEN7ga
wy+tBuYjps9QGlTo5Q7CLcnTEySTRMnEuCyYqydL8bIaXKI1OBHpj2ESVCm7dZ8Z
5qdZH+qIqWbuZnLU3AaHHH1EkwPFq+EX3YzYxvxJQMyKmkvJiNKeHH6MB7KgYgcc
VOM/0mJINOhR4pI4Ibq6buE4vnWYRF7cfus2tMKhWdrVTALlcb1GQ5ff4iftLbGb
SvxOwzNAY6By6P2jlVioAFqeh5Qil/dgtdF/5aAGwHqcwcSdqg6QQ4BauDFKN+gl
R+EPaiFmfc6KgzEPHdbnLcXjw7xQZj0C9iSn4EIKKKGEMce7lGdiG3lMRp45KU9x
9KHA4K4wkFZGGBE2PG7YGxltw/kAO+qYXRuSdgwd+Rz3sNk2Tvrz1azEcHbFCag7
dE1/AJ/2B7VMjsOWpnoZeESzQMYMEVuUWcyrEONivouanu0wUVgPwIaIO2Chp9me
hlEcnyMGRcg8iMYpmyQ3HnHwi7MELiHnCCz+Ijum7f4D6bzIfc2k3eTtoiC5WPI2
zHk8m2uv3LFrv9ABMOMvSnMgBpCj6XfKU94t6ve1V9Z+LXxixZ5BiNmJPUKbH1GV
ij5BdI64V/fR3xCx8j/OvZV4lzxDNklLb3dAZfkJks5VWAhEA9ceOUXMJ5TIhYlm
i+4AqQDILKjzJ8lUrkFIldGxFR3Y3ev9ziWJom+xOBzQfMRraWAGsmjzDfQfaqwC
8zCMQBKY+7rpX7yAJ6c2S/HkSIxXearfoWlwGcvVyfLzg6sMPNJ5rWDT2+zY3fYh
YuXvxCtixeRZKD0vxIlPZT1mV6Mnu9kxE7+UwWsg5q14C9J2E2Z4J+bDH7/Z3zF0
WVvro1stClefkO+O6V5J7lsHJLl8K67zxKlm2gO+T6T2Tdkszzx39yL32I69ByaZ
Ay+/XQ/QaHNM0YRpMwbaszYNkYAyHP4yEU5gCbuaNFvKpcnXY4jNEVXSV61+HYWJ
TYzWE1q++2jfwI6Hv94k/bGIRHOCakDB2QrRSQ4Ldzvatp6JCyIlznlgL8kwqhs+
gVGOCImZbuqEOjxt7suyP5hQ9XskichT6kVT6g4HpLdZNoRZhU7+LFJWveVxyK12
HQzjLP0rG/sxuwfiUlEPQECbQzPiDdqYkLsoGDZGn1mgzGuYK7a9wkxls0RrpWkj
t+8ta++gYmqCbphPUQi642hKrDIEyeGDutE7TCytJfwopiY+Pv+/6Lu5kPft6pbj
tvXdBOAEhr/Gsnih/QNBGBqM8i3Ubgm4fFGf8Bg1TrbiUfKXGkjA1dqsRah3nDUe
AkRF6dtvU0slHTJ9Kd6fRcMykhQWEI6QFW48jGD5+gcuY22a9ETX+X2tSjqVKRsi
fzM3H+WmodZRvnrD4ibQAbkiqeW/icf6G7dFK8kTXJH50rUmfp26lMQ0hODgp3/J
bkcD61YHm5fRvjX7Nar//HIMf9S2uAt7zgBgeYqKVxzYprMU3CtRRx1iQ3SeA+RI
jGtkMdDyidXOfXlIoPOrXwISKnjwdu/TfPkRy5s2ivVCmuQhXitxpAz4FmWHFBk9
iF9ls9yODnUMW2W5RSaJ9tjMQL5JbTiDFvwOSjB/vBokr7hqYCzyl3GoH3fwRVU5
35FrBBCcQ4ZPd5E/rgdnEyBYpU3/XlWI8eLuzFUwtnUtebCky57uOs3Pgp1+1Fc8
QeHwhQKOqDcl+uWHDvEvWxpp1ThA6DDZsXtSZk7bSUdU60pBQ9J/iJx/pAy2/neB
DNSGLyf9S/sNYzruKIJh/GAditk3D0c7VabtbNE1+REIm3NC2drBIG4R2wYimtEe
d1Qs7FNmW2Eq4HDAFkKY6kPF97037ijoHRY2v9Ebqu65tU5mBoWS7VtXpRmM5xoH
v3falIHkU9YzIH1ucDiJQTod3mxunoUHYEDElkNhYc4xNESEJse9+uDu1+/mg6jT
u4YEVcE4JggjeB/g5rWJIsjray5uVzWN27BnVVACTWnsUWcvr2swhYHWluGu3Fit
stlk4imt+hKCv19OpxJP4uVz7KErFXW/1AVYRH5MCD8J9M4KbA4GGwjzHn7FLdJp
j0obsHsJsvpyj/E7ag5MK8kGggUnRntRnRTxjRDh/PCZuptTmtgGWRrwf7a+ljio
4HT/j87LHdehuHikbPrO8sBCGR8eHD+Pw7uTyOxEFVe42svLLekh9LcB5wF3QxuG
N25rMe4p7F3d3sA38Z+BNhQgLJ8Gi1hOk8HGlXX7UQQ38swHWaa0pQ2qFquPSaud
PS362xNjhpmg8eWqNr6h8Y8SmA/LHzPqhdD37yT3DwyyUEH58PRAfINeU5JgzywO
yOuNfTrB33khV/Mtqnc3fANjutPdMYFSGwS7ofDF7qlOSQQzNddAOwM8vlYQLh9J
GdlucIIYyQRaFKpsXh3XnxnYDoLLx1d4gGk0T12FqWsPezpZH5c+AuhSqvDbJoSo
YBV0wWn/kBou2EimaV0URZGIZmWnifLh6KCvrhYGI9kNBizf7IfhrVMlyS55CJVH
0CSv+Przp1KAiAsQLIZ4toJzZyLnhhKd1ZBo6ec/Q4ZsSwkY4TvH3ZfbRzpAJCe8
X7uWw6v26Htkq3i56w/H+dVyrBMzME9415jniRpXtaHpxJEJAYcQUQntf52raVLc
hv8RrJ3Z1T3I2iBDoBaNG5YMqPaXN4tapYhw3RajeaeZnL2+VFNyps0arm7tJQg1
QgnIYoMqLdcSmd/k0a79UMZBTWX/sI3jTyW6tUkazEMnf2t9EAlxLkfzEfPpLmn+
+QuGcFcjtVhN7enXo/DpSO6Iwx9xWaTgnskI0BhBHw5torXoca5WvvA2ZDZlh6lf
DTS5+vTbwsqKZF3kIhi04ckQVMayZdZjJjgm8OuofNi7LtDbPJhLQ4Md6SdVxNU1
yGkboDKroNzE1D6HgaMd3A1tqo11U+zvaVeiLaEAzFxJ13gVCF85AU1Wh/J8T4pn
lnSfH3mMX0q9UdsCQqMSO5TcZ1MAd3Tn/tE3MX9zw2aFuYTKH1zN1v2KHxix4NJ8
2k9A9DcF+zu+TuLnXQBomvzQONLM11P6YrkdIbiWQA6d7POHQY4z2+LF5iVfOGZK
Pl1hr9drI9dpZvoZuulB8DLCF8U9hD7xKKpkihGzt12IaaGTrkGrMX+etuLUMeb7
i+tCgJppbhshN4oIcLPInfeccPkw6xc1RUj4M30b1w1V9vz01BAl/rCFQZVBe7QI
vqRBXZnRewAqWfLBU2BWL0Tql7aHqx565Br+5qio/fshh25orxZ3W1Hp+9AckD6V
HSHUUvqKbAMpnQD2b2vlWAzBm2JfKrtmg//g6aZK7HRp8giLxs+eqmhcVStoVkug
v2vlUavVotR76BDpzRzFK9qJYpe5QLJOHJKu7ib5caMg3J2l20RWPasWY5Rayb2P
odw+ami/C02moXC+4sFDtx8Cp+8Ghq/NS6t1eyKQoBMjGCHj96bbLnrn6XrUKvAX
+u7JukCrFP/pK3CkyY0EuuPBo75xPcaflyHKjfN88gcZ7JS9U3vlZJQil7R8MMq0
92Igaujk5m0N3Uqn3HfF4iubi3+V+WCY5UKfNhWKC/ETcxJjhO3ImjcwZbRWJ/JO
PAh20gTqGUurZt75uZnhhYSEsrxyh4nsVn1aWwmJEOEHxGN7IGUvETu3I9Q1/4fo
en1AT60s+6yyIyM/YPZncJOvpFeHUK4VFAGkX25gzPrBHzzIFRMM2IVSeAtt1YLs
OugwoLkUkrhV3ImpmgdJ04fwArLAnRNg89zj5Clsj41JqvjUlXEfF1tnxdl1q460
II4dm6GqR0kop8eFhWEPULsQW+NE/U4tU/yO41IwLVeR5IxFCkEpZ13uYTabAr/Y
IWXgDPZLm7b3rNRYnoUJCvOzIj+z2jl/xtvR28ZwY04VFPcBTOhV0YAazKxwRMYg
OTaZwK4dCHEaypbFRUmf1iR0jKd83ecFApxjPLLQVSbwHTrzFgGG5PE9gE8cDxIN
jV6M6gtfwtlKBekZc20G+mcRr4RJt2sSc/K8Q7FCbzFDiA9tFWjD3OMSXjfpKYwu
aDdhDDAL2gYH+aL44ubvO0yAyUIF0vMCJQ43TOT+SaR6Ql05QzeVAoubBeHSkITn
1owwQERnRlnWvWE2ae2fqQsBonZmET/GN3Amrd16xG8HkO8U1sD7qvAV2P8JBut7
CLA/fBe7rMVJxHpgHAVQSfGuB1S1JaAYfzGcTHnJ4DFB4OXBFwBW9NYhgtETtIqj
rLarvccszLi2Fr17jC7eVuJpCZP6SD5yM9pN5QtbiU7X2R277xX65dkw5AAtjXT5
ZbU+VvdEBU67GmUIgisCikQccr4ist118DX6jX90ISG3FSRQ3meKfsO5v/FXeUHg
E89gZh5QfAkVCOLJiKozybUl81AnHmEDiEmlbiJJxmBuo6F4Hz4QyQ2rLmKiJgnB
k93WBDLFOuhQIk+sKXZe0IPCRLhOYw7zC9Eu90aG5GDO3zyCqZNK/01ARI3FQlyP
oPpWYH/1W8QP/cn0lO8x/bbXjxiXByIeOFf0nJN+3HDkfDSXaX79iot+XrLHOILH
cXC78y2Bl9eM/lfkdETTrDt3X+tTyk1ezyI3GOCrkeAGwzrlrJEbTBo2SWbjSPjg
wrq9JqmNePW8jJEShIyIVeC1Crk6bHqkXXnWmij5eeD3LpIVLYlZGxVdM6IVSiWG
3eUDlKn1Pk/lyiWRnwGFP2an9G3imUW+Qy1Jqt7y278QB5ozUI1vBvOPI/PKHXxa
cQGXOgYw9CzZIqIAg1d4SyX9CZc+Yb8+h42mFM1BpLyWy+xran1oKWSNXYncB0HI
S8j9uzhrEt4Q0msUrHpTS5gRf3F4+I8rUe2g/4rChwv5WD/yhb0KjG1/XCfyZWXW
mwxsNH+MqBMDq6fuyQ4nL5ePwI7Lh5+UX35FgdSaWZ7r1WzWx1H+k37GbQCZ4RMS
S/IBpCF0lrRxGY8uTNP/fV0k9wzmhVUfY3/n/U1W2zQXC4RHD9v6mDbWClGDcTU1
NeU2NbBZKlnAWZqruASPSZoKKRpUzt4j9JIGNBjmaAiJCwMkY8BMAsrp5uNmirxN
6Ljtzb9yeHFMZIBftXmN8epkNF9InhS5vn94iMnRZcfluPaG0EcRxhVHbAQzcJAz
lk3eisUcquZQiHMpMq5i00gGrdUbR5ZSLzhtCOQNS/+5V1TngORLPFNfwJkz7aMO
RnULEEz+W2792GyObChN1/GmWynSVbjC30B9GY0Tu8rokeXsRa/dGjQXW1n9BwXi
n8aLBMjmB5ylbiOV2MP3/lq1+86RY78E9madURcaear+PDSvJ6XEtX0F1kukeNRD
S1BtnOk+DVAaw7ELwqfpKFoWbhE8VfrqQSSAhhi+QI7SE6d6H2uQKKktZ8JeGmaU
tqCUf+6MgCcBxT5kHf/tUmkfZI+B7ZpAM2AyHWyIGj0dLr5b7AAUlv84qaU7x396
FPjivmDFmChHtJQ282r2HbUsomVGEDfT3M1bXZ46D4t2RgpDdYxGIaiMAXUqS7pi
bd7h/v+cgnNYWmYV/reVCI+bg2uYKuE6cHgOjDl3gvMURIWYOJk7JHvD+yoDTfZW
Gr4WJ6dJyu783LMJSU2VimKH5+Ci0LMouRON1dzs0fOxtgUmVpD54pywcF6FGghj
YE00Q7bCQsk/LcgircV9qYqY4Nk9cIiVXV1sFda1GIGeGuFD0peZgOC2yti3VLQW
vdXgMVEaxhCsDBAtu6tCmF78e6vdkRk3kpK64l5cewuEYBkxoBBWZmDUbT5qU9+s
bONedcCkqjuO018bff8EjRF095Xc17KFuHAQmajWhEXeMAczYXXIYqTdKwQN+Rp6
fyLsomk0wxeKKpMbCw78ZZkIa2GKupg0w9dxQm67GFnSgdEKe6xzc474u7yqwHRA
KaJruzwgwzg8YQsC+c6S41KSwEt9VUrp5dbwe/xs55zZq+jA0sttN3hp+Qfn5sT/
sUoIK9teI11l8HnVEcEtEynEraYxvNGLIxzsVLHCgoeM58j4iQMUxtmIBmNorgmZ
WWrBo6Z3d74GNJR2ULK0a2MdhTXnunRHIDZxb0jT+k9MsHr9DnDO1SgEeIB3uq9z
Bt3Mz20fG5mgW6DqA6jc14KuQBl0K7qoT+aj4i9T7vDyqJrrd3ciUHAj9IjioK5Y
nyuTk/YMPga8wq/wo2JKOsElhCMk4Aqy1ZdAXX0f/IgicMFjLoXMeYW7oLOT6uhn
DqO4w1Oifg9cWqsDkbAso81dPAijRCBM//RkEOL+aEwJYlP8WasFtiy3PI0ekcoF
GwIRjtbIbGWSecZ2Y4EKokqZT1NaOPZ6IiS9kHwhiyFv6ZobU7jDAJYPy+tXUuWH
2/FGjdAT/GsX2d/cC4fVCgzv9sSZavfAlopDnzAUIoDsBQ/TnsIUFUJDsA9JUPNk
biqx5n3tKq8HMPaukWjHLAfyMtP4qcpwvcDKnIxhiWbPtJcOvibUf4nSBWFvRBue
+ctLhLwjMKHYldvBf6ewXGEzypFakc1iBYAXZd1oQpNm6v6lQbFQtykr5pJCN7l7
5+HbVyesidQPkRe546+5ue2PVI5alEWrgaWE9q5xnmCWug/uDdKgZWNEkGzIPEkz
vXiNx6wb4n+yyIKZNSfQyf5QJIbym35Re0rY/ieSK/PtJffRyx1iS2CM4mT46Bmx
itGD+heP4ayuncYlWl2ao7BEfxYxUrxnOr5NBlPLfbNx3Kj6JiMGlG3o645Ty5TG
uTg8ibVnWQRpnmPpWTaynaQxU9UdSSG3k9G6bqcZlRp4bH1caRW3CtK4ldAzX+9/
0rDBQOVExzNocYz7Ly20tdKR+YLRAxqejPDRosONGfqaO96qgPQVpVkt5AWAhRXE
nekUAfMdxNXBdvTp2NgtTG7BIlztC9FFkLDhgBMEZFNdbjjxWu2ze4OLAIwwHk6f
gGq0UYRZ6SE4igNH8z77sRdpgtaCKMYYzxIHLNvsmDXfVJhQfPY73vZFT+GvFONI
kAvuJ2wf9i7ERJqWsTSBtwZHJL9+OkBcxMhU3b9waOghr8esbd/jRBT+pijKoJav
0gWnfH7pM/sfH0/ebhnAWKalOUYc+rRirirP9CuLF6i5CBEeTQ47YcSK/iahdzZB
DgMEMI4ZtkHnAf2TsENXTo/QLsW4PxzH8yOYRHXSEHadfrL5qrLJhehmo2NFbJZR
Aiao8Qu5ZlILDd0GtQzYFt6ihXxrL2Q22j5/yszHk80kJa6C6Q/82N9ZqsZIiVLt
Ke/SLnL8A6JkwsB8oYU40deTvQm2DG+aVp3DtQ0Qq6wr0fVdjbQ45ukvo5ZztBYr
qWflQVHi8tMWr6GhinCBIy6A+e59bJdE+3htoODQ86pxm/cR+XIhuRE7hoRGpMTP
ZfHOsRQcgtF3I4oYviHcglKBaKrMzcJfckylm/jLqiv6bOTyu6orDyUeyhemXwVR
KwKpzEVCymGqWJkDP4zd3XvT+rOzAubo6PAvJdKKJsf/6OT62gTfKea+Brm5z5bS
k8FVJLtcudp3EOFv9gN+dE+bANIuScffOqbKkMfV35+6QETLE1E2r8JWbMnmqNDF
2zYZyCLYroOYL1azYIvBt469XeVemH90KwKvmwVljXtnVG3sytZJGkMgV8NHqXSX
6XmTsCJvAN9VUQLiUFa86UotuxrcQlV0Z1tz+CkRNCF/BdFwiWFyvA2FDwPg6xbo
ZUFc+MQy3mBl4QFOKGPFh6yw45HG+WoiTodtl1ACWQl2ZQxRQznoo+7GuWGHNH7z
wqRw3wY0hTaj/B5CgGytF4axHeCm2UuiK6XnLZEu42D8faf2TXoXjWA8OiZZYEyR
Cn31xrlf5GBeShfW8sdLnIxjnbwPVCZpFIDCzRq3ECbIosDUJe+5HQefVr1+53EI
RlJyFi1T7TVwn4lj40KTC7pErnGs+sf35PNrv9wLYnKTz/y4TBj6yj5nwBpsjehj
66K9eO7Z7SblRlxJ1BO1/vZhSDT7wC07WGYguknjbV260Y4vrZR6nVfGOiwWkShi
fNktO5AQ1n/wRJV9C5z3FLKXL59/4/Sp4kvGa2guyzilBbTXSEXYjCW7KcaIJ28U
tXqqOSRC1HmQ5ALJvNWW66qnVB3lVZNuelue/S6rkZbFIwjG+sgJ5CnfOsGRKpVW
ApUe5D0poBo4Q0SfVOBR7Y2yYiVKo5w5n0KAKsNih1/8We+4e5ud+y+xY9o0vAnL
6foupQTkOVpNBB8vx9q3zVJqFnI5z7ndHulyqdoEMEHJQVJlO8CnCBMz+WPbtWmf
oC6ePfo0RdQiFIZRlXOba9tH0EB8eNFDQTSUJjJY1KIjOeZu9gI6PCXV5hZ1qY3H
xgnhLokYo9b0q4VqPqYJ5Ow6PDaK48ue9C7XLVKcisC4Qu7LHfLj1bbz6G4PlIOM
Bjom9ZhNhC03y0HP8yR3d9zMlcxuyq2w0J/uAC8QSyqqMbnXUTts289tAJTwfINE
fVnuah9PjYueKIuzgi8hE9g5j6qAVDd61Ry+ymQ0nUQRKeiBnwFAg+dx8kCzJi7c
Nps8U1BYbe8V6jZlcn9ZJI9eaVdpM0iz5DLxK6cp1Lh2EyVbH9VsRMCZqn8aWpkx
1qu1fFk7ey/AjF6grnXNsYdZNhLuNjlPWTB7GubU1YqSh4R93WL4niSS3qb9LXyx
c++ZkkhODSZPU7uo0MJ0g7OeOsuXhDivKhj6kI7w7PU8qEcVCk8aLyDe4TQ4hgUM
n3FB8lxK9m0eghXlbYfAdoefefjveWBXg7ArMYInvpLojh9bKL68V/uralIRFMpR
JRFRcOzKabGwg2oaRILxlcWgqX71ZUQgqeD+blr5ZO4QAdSJjKq1ky2xOMop59S6
bj1nzb5PRGKzZVMT3lnxhnbEMOCjH8TjL75fwVwHNeVCgqaW3lckoSbiYtxT6Ou1
6SvYmGOZ4d7fbIreAti0K7x0ux4P/jJAMUNW1CXAlFEyI/Qc4O4CAm6ZCEURm8az
jvFiUjsAFnKHexIh26M9jGCTS9XsyhyJq3ZbQ+ks2qAaZVUvWR05Nm4QViFz8MUW
9Pvu2H/fOaunbI0Of7A/xJTIJ+Y049icXyolHubniItZLcVb34g+jwQCZw3LTYF0
O9rPVURk9dnoojpe1CbVfWuNbwOS4GwRR0+oDTQPcmtwcCz+CUZ3Suqr9uLzT7eQ
QVA1vOBI+C2jnRXg6TteCQ/p+HFEdXbD7WSs+Dj9vaung/ote4Z8E2mdeCDJuOV4
7BijZ4efhAM5Km1KdvAlgl8iA5w3McuKgaQWdTUGOpi+Aerhv1d8EhyD7RtYqXQ4
ofSG4G5U354yuv57NgbY0jiPUHALF2joERotB6PcGWtRWsXkBd9XnW15I6ZNHPU3
XtyGunxy+VX3QL0SBdf4IndFZmOAZDApKQCCWJq9BwrHRSPOG5HqGFTLC55yqVr1
2jTTBxUQnx/8rDF2uEgHCnLiy3jhMBci4w5Vix2Q5FVLD7uZ+/avDpz7YJ70OSZc
hYWX9sCJ1OR9wkGKNQwb71n1erRNpJ/vr3IaM9WzyZ8ClDKoHJY/Zbf+3Jfmevqp
/bv4JnXRvFawVoZAS3mDFtJObfNncUZ4IhOcbLQqOUmu0bqot9yTxpbnXWFKuO4D
vbCSW5cO1dE8VaMnCbmC6/pgfcM0MdUDt79sI2V5zeZcP1uyYQ+ggBSSSOWrAWpD
oAbyydm1xNMV+8VXBxAJFMTnHRXEfd4KUM/Wzn88xxorcR5E2CWENPZoCIdx+vMi
AxHwG5OcsGihNLFfUFrg66maqJOcYiQI1JMqpUptoBQk7EL/NVSUEIyIVWmkuDq0
retKz3fougBrNvmgp5rSQDLK6rpazJU2zuNgQ36gMojhPYwhaNhZt4i2hRHDVt/2
zysNRnWcX4p8KFe9YImlno7iRyyy+2SQqDAPDEd345MLWpZvtE95oYcYSVIfPP9f
7QAhBhmM9kIfNvCs48v6/JkjlEGNpk9fKFaFBqJSuJq1tqdGClDqlqpZq8NwFC/+
VAUP0Fak4py8vmvJUdDi2qooyhXweosiy/0XSp9EQi5zUSyJHbe16D8cunuyX+3a
2y0HMzzRIlDUpvl71DQhLtV3RJpnYKc/h3NFXy29xwRELcD93P7fjxiJulOpcJuN
TTyeKQREogQ+tQEfzmLhDxH39x1Bqqr1cXxt3BYpeDptm68ppdgQT6JKmpkLXNWa
UmlhAGJaVZb7Xr9JbDZs1AjuSQfglR4r/CWBUITQE1g+++nOkPFF4VbcUftdgnhM
ejE36iBGCEgn53GLDV5KUy9SM5lYU9nZLBfSYOVnja4CQ/IvzDWCmm0rtRYCW96Z
Gu9Imjpq24V7K+ZYGSqN50l3s4PViM6/v8/GnW71blayUoNK+yvRM8y/Q9lo5BIk
wbMiyMVW7YSGNbVrWL7ZHUYnkzO1m5QkTpEmDbuoxftLVzhkVusBhxacToo1rpXU
wWc+RAaSxgYmHOLgTSCPIAhnMo+WfSI3G7sCxC6wM1UwouyGq6SiWU2LuxmW6VqN
HB1MRrKL8TgcHM9BkqeTcyPXO8pWYoeGSnLjaFfpLfc16D/Sguy/vDslItuo/ikx
2BhOHFz6qOvgFKgg+qDK3z9Ayg8ElSLcNhWmLrFMt6nbgLZdF3gYFNSeN1To/Riz
zgVYH0i85pul3urm6SDfdtS3FL5S/s1pzNtoOJOXTrtOBIp0v2xYsMll7HfSCdeG
T42gqGub9e6iqbe4WBDFzzMdFEu7v/y1bVnUE2sCan66VBOO4/yqNpk2m4Q0eJiQ
5a0m57Fr8dEIYxABMxxkHIhtTW4BYBXugCDpMwpodz1Fwh40YztYH/xJeD2Fi2rY
2ijDu/UBI0khSOMxIiZ8ww5rvnH7FVCCMad23aeq4D1Wa3ZAq09vgvEtZDOjf1rt
7mt3OrCKgAeKP/Df0gYjwaXumpDlbG2iSzDoW77ToRTNcz/ESqEtlGUYt7V2Xzej
6/CZlnsu6g9+uGJ04DYWLkZ9aRe/MBBBkoajYj6oN0yRs0kRFWqKjiTRc8sVAAjq
nsO0YFr5l81F4c73T9XizyTBYaVP10Qg1eht+h7z1+qeFNscH2DxM49FpWpBZu8/
lQT2BIb24HE1Ix/mY35y1L0ZCYwuGuM6qJxT2F3AMQI30H6r748VEMa4DsZaYe/X
W9dfRPtpPvrVJKHmI4IEveBaea5wabKjKpT/9QgZ1OpuEZ7l8m/Pw4NuDP5txaN7
YbEJVPAZp1ghaBtLMKdSoJ2hvcXNINi6nW1vbXlHEHiJSL1OZeknujIkIaDG0B4K
ZE6aO3Gv8ePiIlu+uAv0tx5D9V/SQp/rEHBZpOdfLTmXNH2VUvMoMkDGHG0VLESN
iWDa4x+eEKpYidDnsh85DiKR4EbBESXex8vpjbQyRrp1A8ppDGhxwQFQj1VYW43s
6TWOVxB9HrjiqafoozH4dT4+kH5k/flPTQBwCLHOoghJRXLVYZSRGqekCOJpaQ4G
LdIG6mn33e83gOyL2vvNZUMucItXderosDEDGFPTWCdgUmpRDy/5UufeJAz/H71D
/eEVvRhcqQZywH3WWoy3WKimn+rkfPQYIPgMthD5p1DDUqT6HULRcapn3Xt3F/qf
HBaAZK4sRAl1Em+ewtXaUZ/M/rN3YbfFbHKLYU28F5LQcd/IYKymqOrBhVXjDClp
PxdBlSYx+ZtYj2AS7uOAWBH9O33GbeHutIrYH/RjeDda4pWsflPuFMFFFXoiP5BF
zZPt+yo3aBCgW5jJe93T3NstJVKIW+ZCJHUYO69h5nNhEw+JwEQupTYrorNT7sEu
ZQaGTBlWaJ1UCMEZ1+O42O5v3NDhuxA+r2AFPjpSdjbv64F/uz8XNVeUAjFBGcHI
u9Z27iJVsAoKHDuLd0yQVQ+FFJ/zZDOQ1eFeGOLA4/4JmMryDPqIo1hKDIDvR/aA
n2dwa5ElBzeox/nhJymMYCn+9bzTifcKeQCtMvf4VbevRE08rWwlHrtjlo5SEgYv
fvTSlqT7N9A/MA6cQEUoyjzbLlMP+eVLFjvYCkZaYiGqkHUYESTGU2JiEQlX3hR3
9w4xIxiS/HduBEru8G97w9m1j4a2s3OrCDaHTKRYKclBAO4vvXH1da34PpSCn+Vx
sG1eoF8l8NYVyy92ImvpaRnLYDXa37UcJ5zLcMLNElwKxGvl8wVFCQITZKyEsh2z
nZ67N26FSDnV/1Oh6ROsIr1Ib5AlZm0RX/l1adMHPdwYN01ZO+MDOLUSUhvGnokQ
gvf9T0c5EPc2dFd8TotdMPUdP8Qi4c7Y7xrhUlz84Hv9gDNMRyaJiiR9Miys/TKe
IIVWTJSqd4X9G1fmW7lbBOxsbWVE3DRsUNgfmQ/6xKjrzt0i+W/J/0q2w7nIqdeu
nRDc1NfDfLve4Te5BmAAPeoiUd2bzsBh7jbrfC3zizYyr8L0+1xNkz8S7tcEG+TJ
iPepRIhctlWw/bXRVrMShniSjcP/xrxc9untGOe6Gx4BvTkbPtAIcfaxSzKiznB6
kzJYNbe9KAQmWEz1mEXpCfq77GxZfhQaqMGuPR5mnd9CrgC5ELjtS5DgmMz+KN7y
N5vvOCgFQfdEOJs7hX5iHVirryWpzldTNR35v0atnSMMK/Hae77aTn9UK8i/5p19
Gp5NSrjbnG4W6t4yUoDdq/8L4N22fup8q37gzIknTA/RN7tlTnQBYHFQS9zneGNV
TAbv6nE2d/30IJWopBREL1pwEZu4nUXWnByK05znU8BVR151sq2Dfs2KJUhX/8fb
aSTl/fgRDfoCe2Nw5/TsbRO1M1ottqssPyO2bXacBPDcZc7yY9bovruzPq99qMS9
gOdmzADjmKywGStS6bnDixSKSmuOLge7OPAen7VYLzDvVFQ8HB/5eR63HM70M0t3
T74CTb9Eox49yu29+2CM/z/RMvwfzgRq1DxXiLXPIzrqnRV75z9NI9pkU7QlXZ9I
ko3j5THAzYsCI9dVvmMJdBNJQ2z3ctdRoMVDs8FBDjpK5fTmUT5WxbUjm6MB0zRs
PQFmSUOIdFXc8FWYL0PquAxcXLrohs4HM3vNecDSt809e3faaz5gnPoY1uTmApos
f2SfZ/lfGmaQHC0JkR0mm/KLvSOhoo0dZCQcMp5nbnmUuKsyWhNIpcaW/wghnl23
5QWfqXxn5sWvFt9wQ++1ZaDyCpV/Ae/wPTQufcnx+BJggbOdxKCmd0sgQAsCj2Rt
7kNX1v8NWNcu8SQWYM5dtHUa7i1IyySAByJkZBbEWhwZ2fVXzCTIZHG9ob6RClHJ
m0naHcBClNlJetpEzuKuMtHlqtAiC5yNaYEjV7SO3/+1h4vMIRHwuzpfDdtAXxBw
AonkkVQ+yuOR+zd7UwYwOqg/CZrPZdDFbH+4MeD49NEOU1xjEHlgpJvSWjnOcHzg
sHS9srxJnQe/qTB61zu8+da+DVy3GnNxpP2EbgbUUj/vxC6hwlalaReQ+HuJ46ae
C/rmsRZ2FMvJfsKfDyy2W9xie2ftdJ9q3dhp/SZj0k95Q4VmzUkvYr204ELePbh0
AsbeDRB6nysNlngWyO4OrhzZ3ybPyNFc1/RjhrjGYt6OQldAbkfryI8cR8KRg6MP
ZqbJdOWtARQ2zAj0WJRyITnJMKHzwBa+uQWqEO6Y14j9iDi4JVlPaLS7NSJkq+oe
Wh7iAARow+f84ZDfLs9CJsXC8zpzsPvCIndItm5NMj9Q3rRwcfamkIB0jkf07VHX
60H7gJ4Qekhlb8zi/i7qD3y7NTq3d9wTMnrk7qS1NYAIO5kL0B6fKVLnwGM4heQ9
d9NwEYRtPoCn0NWpwYiJtpNBMZO4Paf6VqJcHBbJlaSW2ukpIoSBoMBbh7uXRK+x
UHXGop57h0+mGAgJkZkrKCEksIxh/fPKndftkw9Oux5RWtJU7Bbfomwvc8GC21c2
UtKz9Gq648hBNC/owYYLSugueetkER1wq3iy06faYnmZ2FK75YA/Eky3ZbM9BGl6
NCWISamQAr5BmQgS9vSBD5t5DlrCvCU/ioR8fG2gfFnpjrBnGv78m0e69CQ4M9Sm
UlxpYDXM0FrninL/yqNxduMjNuDraAjZgq/DulNWMr7ygcEWVdjxt8VGyhmjcTUA
PE/in+zP7/fX2sNYEmts8xhSlvpFWZkAcoRVPSUBwWkPapz7ZU3nCtGs5MDdG12S
jmVQnzgzUfKYnUMjgzTbPxgewmCqTwnOfH1G5V/283hKwj6NezwRQiIfZPtgzvEr
nvhd/sf6iaVIxkanWkHvd4Bf32Zls57SfmlETl0gSu2CfiYl4PZgdBdwoX8Upjft
8tjPS9t01mnWnvMZ42eI1ibCCfMqAh+PQIUad3n7jNSpcVxnv/LyRDvos4bgxqGy
hu/DUmVP2fgvbZ9ZZ0YPrByv+En4vgR07TLqIamGijYnMf7pKuZpA7Z3j/H1WL/i
ei8o6mWUjXTHrq/BiBC/2MoB3YHOgJegKkgZik5Rwwl3JlyYM6umr3Bo9dd9Zsmn
FM+Axf0jm4Yy7JvHFGGelAYtsXaJHrOyYmnybHlNVlXG8+FTLgy1Z8QSm+vbZbvN
IrHXRCwcwsWDTGwmEXpqhtld42mFINFMSKSLumDcK0ObwpvY4YWCtcqkzfzvRmja
hdxysm12tuNk6fP4/uk03WiKptQiSt6ZFEtN1sbeogrCEh3Qjz4X7TFh51zA7NKi
Vng/5W4wZpWK4NRrZNgS4tPNjuT3uEu0SomF6tsGd7NNaFMXBPJlSB/0OyH8M4xr
e2L9lmd16Jx5CzBMepmQoYeHvrH3ypMAKopjuSOoPmC5lh65vDmKmp9JcmZK6q7Z
b3y4cA3OmKsVaxJtEtWnzAHmLvNkjnZKyW0v++nNQNiBTj4/NU5BA074P+Cu+KBm
3FNsQrydMJul0R/nm49ki0RRFZO6N5SenvPJuNV0KbWSsgExhzCDNh8M+ejceHQA
C6cO/F35Eh7ESLrOTuftjD2G+1OqZte6Tluv515dp3bID6836xFtl3C9udPLymgC
HnxoiSwvmbAsQtOk9lOcQwsW9Up/ir9kFweU55y/zpyMWN/8RZEUkXfzlZqShYLS
V9Qq9auKK5oEz79AdWle/rOkL/el38x/X33e8ZcJC/vY4EEovnc4vwQV29088AaH
8OjQbha+x0sydF6bCNabVeLn0oz0+dTfabK6UBATD0wM35IAU7GwcXGUI4TOmDkr
uMQS4+N7Bn5PED+1+BhDw/lz8Ex895+pJTMsQKW3vWDEikexLH1Ha0kc7Lifm7MR
pNsGWsQ7HUOw90GpXuqKeERQx7rU/7QGdfltGBdKARF9D/DRbkPr7Ib0UAauypbp
GjIiLtVdG6P8/3qjLq/9FXvPBrG7njrBOOSL6h6q9Jz7e3yV1fu37n3B8HoVcGqT
MS8a5MUvm6PSYL+wXprnc8JEYF6nMqjaQBOYMGtuA0xdnt34ujgQ/Bwe6mfdl4sq
ccxQJwUCUh1pozwW1iDimMCnjk3BOtfP59mPiIboFROzzf/slXvLzZqmzLD9FsEa
xNeVea15UgCKbePGjgTFOFR2Jwlak0zR6X+bMuCqDJVpnsjFGd48hUQoKHZUiMKy
csQDSXBdyxewjZnf/U42Dp/uAaT/p0WRJOr+dIjQ3/T+2LbUpqWGc70zaJMvqUkw
4bWBBvrC7+QP6zwKOR18ScHT2Ua+e5dONGe6xREpntYP5IpX5+YtZnnG/tzMOpVx
40pqKeiO9R4TR++6G9LqK+VBnMhRgLtfJx/mvTUOu//U4oDlnc4h2uGkMzQztAC4
W+PCjlFkyrvEFzSdI26h8J9rqVZ6DiStFhuLNxuWqtqCEnwNn4j4jd6AmJwH0yNO
nw9V9qvv90xxGoDCiCTdHOS2TJRd1nwXE0MTvrpzZUB7ww38xu39uh0j6j6CUw0W
Nd7OD0PE5COxwUMZOPEfPAG82wYESmQG9qB7n2gHbuh8IabHctcPIJSYXXNzT6KT
Gj+QeYcqoyaePEu6KMP7ZfzJpkxQ3k2wX3Nitb72CDsLMvvPbL4NohvnfE8mGr2+
l/TsrYnXdVM7OrixjWJcuHu1P4/w2exU4fGziuWXJFACXin+/TJORxsksdSDy0ex
CBCMXmi9BRRwVtKzBsmHf5z2FDjg29TVFh/TIb7n471XqiwY0N/BxM+vLLaIe/wz
PxfmwXyDFuWGlNMbgff5SucrkD1umzVaLv/d1/xSTXVliR12NOJ+blnSSwI65fI8
zf5EAx2CKIhx9fcdJ/0hMmnCsBE8mc3E9DbWIhs9LSAm+6pjyQyelQG1KRRGetDH
jroZIHBbqOZ8gZlw+VsPrTGnBJHQYccdljMduxOIkBmG9hpVZ/NrjcsYlMtczwHj
Fpzinwa80Bnd3EanTKH0zasD/wgi6ZGswucDPxBbpm7ZoiNdVjnxCrW1ZlzxSoXi
HaHWsdwocoGHak/7lOjmyMaucozZhUc7IL0whKrcd2x2nEPzbXWhbPGshgfbOL7+
TJijPgPfIWBb9g0VRh529twgl7Le9Ry37z+Nx+wUsydZoWYzjSkEm2AiKRlgGgeD
wqWKwhyHc7fCcLCk37FvIYMoughRgI6rPact+M30id8++wmd2t79xWkVAGQewEDz
KJWvdR1bul3NGg3AmwHeLh+4saStx/qwmJZ5BI/vOoWfJgdkqPISXpx32SCXmnZl
ML0th+iyjUn5e2uMYQsKibvYdbFT++K+yLOtRBP7ezZRQrtyoSPPSg/SAnAXvifZ
4u+6N5n6JBvwUfjlsQoc0DDWHq2hRAhmD40Gtwq4k+AUO2TPURvCAv1wUM+BcdPY
V7KWeAW9py22SPSEHiZGvx/IbKS6DP0aNkHm5tLdFg4sK0lCA42hMH0XCO2Vhhzu
75V+Kvq1CcNUguJeCjxrA3L6arsppaLVG9bhmQpyRop9aap/caXB8Dd0V149ilnE
x2WfZnyrL8wvBxtmRP7/9hRIOniD3JXa51NcuUxi/ZOQU2HphIbYgMqoj/cSyk93
F97Iisix8yiz3e/aE+crV6elR2c8VOrIUygup8poFi49GlhbezXkcS9esuKoKdlu
/GOuWrT8bM8azYXHB49NQikdbaOHYnfvo3UHBa2WALnjGzec3SLtZm/FUe/bP6tD
FG2BCrgC6eQlWIz4M1ce4/brs4g2bN8CClYDOhGk/IR3jL3Q/hhsrcAMu0LTmOIM
LBv7PA5iS/w4giE43LsSF5jlbHnYgjTG1KVwVH6Jl6F+LtR0rbSV2W/AHkO7t+cl
5gLedptDrBEBwVgh37DHTMkcaXUgpA+ctk715vEG+kQ7TQ6n3RV+d+Itl12POYZ1
ZW/sQJpTaSL02uqPIlcqYPP965A3FZkQu4a/8g5D0wpEz5IzOOUJycrElH3GPUCr
RBKrfSW0GRpJ6uUwXJzen6JiD2kD3Uqy7uprX6FKkOnqKs7QmSya7lA1TAEIlUSz
Vsnr0SLLGP2RT0dI3wrr++Sb0R7YmvEnqGHA4rBDzT5ISx/p6Kq1Zv+zLlgVuWXB
UsZWjHFDa1QNykZ7vKGgCl2RuVK/ydZb/gx8rJoLgeef4OPLfxrHABpCZzM+xqgu
ijBfTXsv9LV6XmHPqccjinDsP1ny3/TeN5v6N59WZilwGVSJ/DIlPRd1V805bD3x
JaKBaGA1VOGuNFZbkrGau/klZCNIMXsdTfWUBH03JUn3ySVAchSp33QerTiqgZiV
ZwfSIlUNXYgLektq6P8YigMpmdElepyZHYJUElXMI6XS3OLgan/JqVzSh7/DI9PB
ag/PgI/ftLwxpm3/JRQb2yHj6V+0fPxeuBkeY8nzt7+2DUkxZcJuf1LQrqs+Wb99
2G8nDa9rRqgzvFsrrvTARu5euv17Jw0q7rXT+lQgbt5XPhLtTZVhkPfl5GecYCNa
DDvV040XsizNGRRopLLMyOtZAwMb0LnJjss0ubBQAtkKmh5WZ6CqRE0zwkA6+pjv
r291/ylLaP9xgDt+hP+tWH7BBkNnHPisWOd9EyPT4dVlZRuHEXuHh2GCgqDbdwl7
pffxQzNYY2EKcQfQiOtVg3Vis+rNOGxTa0Qtw6b46anWGr+11zpVKT3HIMFv4loo
/d6AqyvrIBlWudyIrOxZJlwFz0S5+WGjwfWuMrH+dN4twGeSDyaVCDfBa9In9SAd
VU17U7M98G8gF4Rec1XykGboeSjdOSXW4sweoEkwWjoSBrA6QXPMrnrAH8yL0dON
v4MNLp9/Zhu2AQwxdWsB0rUP+5qKKY0a/BLdYRRE4ZZM0AVT+k93kQcZup6+KCPB
LVytjN1x3bA4IHGAiaa10TCrUsmMaHsAH2/UWRxykijk6Wtbdf/7+zNI+aIVX60h
tp0wb6aL8VnM/9Tax/9fz4iJbskvyRKLjKL+9kb4ZNpzHrN2q6pWp383+NjGA+lz
QlxhRNBgIv7+CsrpYOZ/4WyGa5Un509ssZpHQLsGuT2qp5kg1xRkLsIqc/i7d28p
jEU0VIilUEFbliGEAxvZlME6eU0ofl9CRbnxZH3JUFzb/JNDA9izmt6zVlgoQ/Q0
NOCGxvC/WbIA6N7sRFlJe0Hob2lpZnYL+FyFUkDChQphxo8Q336e9mAAkFN4t8jK
Nts/IrtxA5Q1U7yZXLwAWRKfnDmmbL+O8grmaCTgPViVAin3/miLO+cuPWJOIQ8O
XmUn0UPCTAJKye3M4+p7u/KVbljKpNbMdCvyI9ulNiz7WP0k0jl2hZFCoeg/zUD6
0ycrimm8NtC8lssQNFemXSSj24xGqEkxozXT5VrdR0zdTdLphHh6H/uUNoefGoHd
M8rcX/QVuOCevoBeEBcBuDf9p2iz7UAJUZ4PbmafAVeitBa63BM2kzFXqkdsNK36
rnN5dXwUctB8M+sd1FYUdb+YaQy2bk7hOvcR28g7FnANOF/SS8i1cRVaHnoQ8FWw
CQfd5TZV5tnPxW2ZNM0xUC9Cb4WPpf6UBFy46aq8+8ExyrTwIVGrecJlwD0prYi8
zUALoBb8sVzjy2B4XAr5QaFaDPVZXBotBuz9W+0PnoPzCM0k6kVPxzsPmHn22Icj
+PZYJy7Y+5z2pdLc4bnrcJPwbQl4hADTi7n0wTCYBIyYTOV+h1X/MDnbjZsrEQNF
fPy7CGXkVzQYo3zzTCILlgYnC07wQ08f/U4sEAXhsSGtLCYXtE0xjVip+7FUJPsv
2hP60kidrfMsvNRLhk7s4QRg6hnLi/RM8HrQV5XrlhKJssq2VyuYsi3t/gsXH6yq
ADUlpoqLmWpNd3AKqA3iwUlpmIOg8NCdY2EtUJVHVqTBGkXm/vOlQY9SZCaK88pU
yPxWHoUO7zRG3zfhbJWStpFW80FNb77UkepYI0MYwweYz9+JN6nPkzKhafotNmfA
p//s+VLP9X0Hyfwv8EKfgCJytDmVlwM3JMIwRdFNTNel2j6r/y2wQmlIdcApdlDV
IKFpnLAJFFiRs4qP3WLmpjaOUOu6NutYNc6At3v+B1ah3qo6FLXGLPT4ZfsOp95s
0yKrjxsfyHWt2YTV0ABPTu6M9kk0TCZtStM3iDVS7WCwYej1xmateHYEfGQJX11b
iqUeK49d/COydGRnoFjDVc5sd9BbPiZ3YE+mJfnspJD1x+r3l/kjEJ/Bc50JwZEB
0nQrK9FIwXwzg73/k8RDImOqVQuYW+N6nb+sMrYr22Rs04ikeeqfGWGqCHTWOgs5
qzkrRpxl7WPhDY86UDZrbcivyrPxK8whF78mUMJPbLNhxnhpJ/2+my2USoU5qOrX
JdLDM6K7VwTV+aUW77WNmgHg7y4ITVdRVNeDflB87iHDCe6pnAVVAWfI5eZCF97O
VXDrrkWbT1P7r4yOZpj9r+b78i6S9Rz31yHQhX4loN6tYq6ahLFFVN+OA4Xt+w8S
yj4HgxzPXjtsWbwa+YVVxvbw+dR/kuUFoCWOoC7a991XvHCVmbPMkUyITBzoFrQd
BvCXqljWVyBGBPP4ItcS/F2LuK6KfEte4GpT+9kbg2aP1DMljy49/Ky/pSXuN8Ny
DqjfvRzTgzkEog7yF+yLlekdMopVo3OlC0ws1xYjlt9r7idWcHH1i+PAt2ARQVEM
gP7bzlTR4LmFjz4+nYA82BUMuGEXbasVnN1yLfKKN1+3e2Y1glgYXvtzo/s15m7w
Sqz4UcgqfegMdk+Hww9MJ+W3RLSJIBMeTo0h/m04wB7NTQAo/xP/nKBX0j+Iy+dl
rvJ/Wsk79iabLH1LI6poaNBIhNGgVV/YD4A/b/A4BRDcAZR9efyLaTNG0ysLk4nI
dUlgXJMI9cNpm0QYxU9jdIZF9ZNoXJsuXu/g5majCX6WFN3Z5hHsUV7RyI0ALxKH
lrLlHLpmTfwS1kum29u1+aF9JZ6t+UqRjGg1hVnVi0/ebdBAFuE7Q7pfEq+J3KvG
0rysWiA36IzTIPeQKrZ4EfJ3Xwv+COuOYWobG/cskjlevAEerYmdmth8zHUyORLN
/XvH8C/LBc7FPxRYig8SoPJFLcxAfagusxuS5zq1V8Hf0gO6dVlOwq3ieO1nwVWm
lMqDwinZ17cYivoApsRqGz6/jPFSmxZs2ldh7efSLj8zv0WXxheHFm1m4WAplrPN
58bV7DBfJ7p/jBJkp22P1BSaUfUehHNHkjKUb7MsdAlaZw4aX9ZZbXicsNtV3MHS
F44D6yXdovqO8IQ82XFnbbQNr4PeTmJL7BS8IJv4lpA9xm/dcb3Y8vFH+j0+tZXh
arED6oD7o+GtX25l60qz4wj1692I1u0uCm8bvBcws6Ts0PT4nuGArFPRUeYuupWP
9egFB+yVd8q2tNROSQjfgPiwcDxLAI+mRlwQ8SRHWiqZpmaxVh+58ml2IBmrNNvD
sbsoNnwWTuG+xxjp93Eoz2/k+N5tGSFmdfn+mJLZ/odbh1puCW5d82QZ6VVqXYq5
OHRVNl1fFp8L82WsMqTLltRoUGd6mRhhMk/m50pDanGx2qNR6jl3Tl5vEu1kZYv6
VQszfoTfkKP9meUbkGIwp+hKzPD9DsL656veJFKHlIrgfN4qpwgQTtEQpMmrTN9g
xfCVYpcSFR8Lp3jeTpjxaMdp26ertd7w+0AoALs6Q+80e4Hw8ZZol9Ae4TGPbgMj
Ou0CkHuY7PX7b2ggvr0OY5C2cI66DPTriASRrz5+5X5CD4ZUEMS/SubA1J4FyHi0
JDDc+4krRFky4314GxBCylUJLfVQpIInm+8m6OQ8CMrqZlGYKmAjGTTeVYs0AhTs
lVp5duQuf8g9wJhDcoieqBOibDGWXAFV+yQgSRc0+TQEPQhPClTT4XlpaRoxY1wD
M4njFJCBAuKY0C4b5uTYW5RPhQZtNUkec3Re2aOdzKbyfuDazYl4qIb9oRlgWy4I
1QkYT7Vq52v6tsHxSXlsDqgMJgS+8SvH37u4FCyry2a+xBayP/+f0/Du5T2pflIc
TErLfvizxDTbmJf0T6AaMukO0fc0xkv+GGfrhqMWGuKF0ubUjYIvWlqJ2TQyxRxP
VDFZUiDTE3hn1OFHiXccnUHLecR2e1pWDVpZbK4QEM/vgXTmU0j3k35KeQUpPCjl
oEg/ONTWMmIe8zfqliQO82aK6teHE7HEbS6b8I0RX/lYStGjoYPJ6SqRddfbOGpi
A5dUaaxzzlU/nBRpkPRg2PVaRdYjXJ6FMymKn+jptGVkf4qkiSXf7y92eBqS3xnZ
90B4cJgap/ykvdbPSjF4RglIO5Edqingm1/QspQvWwpv0m/rtgFtLpVIdceIXDti
j5N53aD5A7e80JyBqsTO7KeDCuhDGrN8Pt9xYibSueJnUNsxyUgSLwRV6XmWo8ht
EdAZfhS8+Y5mKiKgzuzbGLrTgODuDlqgcIAvfNnDRZGGkYo7LIIWLE2lHJJXcjyZ
AeCNAwfVuz93Zqmkj0uoRt7I8DUQWmeyl9i9edv4W1dcOIFGtRADjU4bJcY5w6G6
mzb6MwvLBuzXwWxRLZNjovRSWIBtBBztlglKLzoQqrc2EarHHMNy830VDjiNMGid
ZTGtWTWL7Wnfx8wbZLICLazS1wSzYL+ORgGOAGwLVoT+ZqdigBGVI6QxqCd9fF/J
jeqY7ab3lJ8ywIJ6+qmjrj2p+whVNECMe12WJfkpVAN9W0quSc9s74eYBMtHps8D
emnu0Kl4EpqkGwdTV3Bg1FY422BiC54vif3mb6O+Am+lUgD0yANERL/AB/PTYHiF
9E1RbSN+P3t4GYV8B0ulHyQv4fXLgV3v4bwa+jCKNcZOBwdmUTwuE/+oU1SLcNmS
og4b2CsIf9xtBH+MRPmDoa9smayPSkvhjDSVMW7WquJ4vIYsugqG0z21alla97rX
mqhlj/n+gVrCQTDPcjt5FbKFowYmxCxhvqJd17wXr21aAtrKwpetrMdSjrN8YLzN
v6IjSnWB+mXLMphj6xMv+jJ+rXWTo7S7JSsQmeE/o71SiGJYFRL7mAMqodqVexPN
ARp9REvp30PIZHwjL+mqQLV/VxOKOvBC/ydoZOPHQgrUPN6q7HyoJ7b8P7Lec9Jy
wCeLmcNz38570fnodegvEFk5zgrgUGT8aX/gOH4fPh92UYST7Jg6SCZ9/vAf+nsp
da9tTrCgt2Pgoc0vDEz7+pqddFQrL8xXkmTlSr9yi5OyHTIKiY/zcBJz6E+EGll4
TjNuYn0tt2Fk/1fKroBEpdKeF9xT3KrRfNIWIrrkmIxH0rRSQnrBAx+j1NqI3xof
qHC3t3cK3SKZ2hGKVT1z+kYSs78qscHrPUHX3X+zIccPprqPUscb1FxtTPjj/GlE
4VqHEGsQA7c9h1baaFqD7NBTxyQ8u5X+78XVwayGe5uYzLVE9LwFu9lzruLGB1ZE
rC3g4ibSov+9NmKeYFH3wKO3wtKBALPWMg9zGw9+NGMsLSS6SDwmxWFABgvyQxL0
cQBWIN36LS55eMGbjDRulcpiWPbPMIA896/AEBMNzmNTpuq0GTg/IHu3RMs181mr
MuA3K9cwRpe3sgacd5y/w8/g+CwUwDLAKL3yoOQERQrhmOhED70jQeXz25jMpwS1
Fjd6jqQ57oIlXm8XT3QEJOQiA+HWF6keu+YPrmsfVwJMr/QwIyN1zdbH39N+J7Zp
XCsjfuaemmgaNM4b28rlp6rRdLSONyuBm3iueFAOgNMUKgqdfCKbg7Vi7U98ZmIb
3CJqzd8cM3zy1+oYZMM9kTHWna1WmQFOOWpf4aBRwx2ahDxFaIFlixfM5e0sdq2J
78hPh4X2705I+GMO6otGh4SX4Cvb2Tw7PDGXPUX3/NFmG62As4PT+kZh973Z+qbx
vKueghJsUsVdrkD7dmnqJGCQ6OVci2DFP8es/tVfTB3/2sieNAXj4rUcr2Y6visP
OqngkGJag1IwrHBh8UGxnnV/99EM9/pWG7bI7rrZUKkDdEwdOIIcLv6mhelfQTUo
AIFqeNb0cxpauGDrXCeBwF/kFqXIz4H161/Wh/ct20Q8YpcV0FHJMnmRZDmWidyN
DA/jIMkx4Ow86PKFQylb4Qv9KIarxT+nOoOz9WJNQ9ztIUfuIMWQXuS+rhFTkTva
UzE0OajkXAHNErw31WRmWIfbncz7GLSXLZg81F2v6kUOkKbUngD7nuEJPlqDbg7T
iCF7n6KXJgo3aPVQnJkFIOR0xBFZBx4FpzIjr+DvmhujlFbVjKykhHHl6G7gdR7x
gRQozr+t7vH+vGcTZPjoQyzSDa+G8UCVH9qNEueSX8f0dH5rQJgIypX5/OSAlaAL
EwbyyGvOmZ/t0W/MHRrrBVUcbvicT4AsLXV4UMy5x8ZYv1zYxVxtz4VpVc59Sf+f
THpSP826A+axQpH6ObLJuWo6HHCbpbBj22pzofvf7D+YFHoex4VQqJskPpiqWW8G
4lEzeegvApyhu+UPsZ21lBGenjOFTtrL011To4fNLkinGc+VMO719pbCYD/kki5Z
4M7P0gXMtX2Sa6yu/ReKRVstQEEhM05RX66lTSsA67jiAqR+mLHwQWMgufrWf1ju
9jZJmWQVTn9fdAsbxFMlEoPE9HKlaHlC/aRaKeHqFgkD71gnYyqpnNp5Aig95S4I
PUeUN6OVxVoEc6VyFsYHT9ocspubEuCx0lb430+WHPDiAvfFJfGXZa6weG+sgz0C
i60GlyfFY0rVJnmdSuKCzMPBpCSDH8nXNKRs3ydZd23uIE2gUcrxsFjK8HZOeH4C
dZILumgmFmdQlopwXP3gb9IBGjdmDcWsHI9baHCCOEk2PLH7nG8F5mUhZSYaIDG5
VdAcwpHgZhjlRijFGa+fqvrcDOFzYUL8BAQkBWtdCJcdgN2c36oT5cRXvzwOMlqV
lJO/46R6thmVmELGVM3L55rwxnGftOqsJnycGPeR6ZE84CFjAH4HombjozwGtf2A
ILPFm0zEWSN+oFFWiIK79+9p5otedth1nOHUjRtXWYcmDoSD1m+2F/3IRfCL63W/
66dwamocJFUdrg+zolXNNHBOxRvZfITqbGzEdDeAgAevt19yAUj9bljF6i7Fk8IG
TzvxZdkgor5ItcRXsP+D2ERVnvfSroYwCUMPwj/sQ6FbCyTkWhBo2d3rY0Qu6TD5
+2VVD67wA4FXgMRDqYY66y5DGzr2CUFgOU0d6Yov812F0xyBKQZxXruBqIfA+u05
oF33eUH7oxFqdlMKGTUxcsf0SrAcXTLTn8u9TVmvIQubGDefKv7VmvDhQ1G2yFdj
BJateK/toZIoKa8WtLyArwPQModNtmi98fmngVggEpsW20m0BYatQAKhvyOjm0bA
+rbG05jD0QwWhvIR3zkFXgKWPFZGs7QM3BUJP+lwhoZ60U8hADbFJ5AhnZR+XcJn
gcafud84creQC77ucJOOJAV6/Osk/qFrSqcIcXDpDwB0M1weKNNgI47idwPuXYYy
S3B1LhJcTfyp5Hl0JMLQ++T3do/oHFMG/5tFSOZOr0ZrI+ZZPZGwJWTPJ67eNKbc
/2sry/Jhxj6E/RXy/CWTHNXCw24CisvzI7E4KA42Ky/jGsuUCCmv7kRYiFppLLSx
qYQUy9FR5z6vjqDDO5GzqWhXQjSmjMD442hSGJMSR7+VUPh5AJH+4LgVgI1JW4XA
gb3EhquOichSNhTV+7CJt1SgWmt1PrbJl45/RFYLAwCoOkoQdTcYrupTs+Krwv9J
5c8ZVa8U6FrPF0KRkx3p2sLTqfWGNzCTyVVSJ45BJSp/b5Ht2h2gFkkFsVqrgNqz
F3KtZ8h2QIe3AoLIoqCPFeGJ1jX9t5stKNXVQPQ5/sK5MfVof1jKdYJhjq2ObbUg
ilx5qtrBthkyrZkvTCVzZ+c9ul1GVVtRcdh9l/FyN1TEjO4jh3X5mpVpBmFp3odi
a6seeCxUV5LyoinlDKeAUhkg65ImZJDrN5AT+lobUJdGQxl7qMOBO32Pt9oPoarq
l9Lnm1z191f7IUP5XfaVvPPEuRR3JjTwmO4TqpKcvnJOwq8DleHduJOtUsvn97MV
DuW73+Q8c9WwZrIBGIQhWAPqXd1ujgAlqAMAB+F5kiBX1RPe2a6RclzlfC5XsiYb
XCSxT56P0Zbry49PVg+81LBJA+o5iOW4UlHe+trlHi5KjdQqSM7IK7uipUm7qd/l
oqTQuCfT5QJE8gB4Z4rg4KMuqM9jOKHWmUpPo5nGAZJ+TLjig3cJY4Xh6sPf9I9N
ptfhG9KzWXx/1lts4zRBHkjJVntZ0TiGyghiwoCUuNjSvT4Km/0jCU6G//cNAVut
2v8niMf7GLMiknhDgx/AeJa5I7wrzImvWFY57j+8Xll/KsTKz2QIGQZY939Ll7Hl
zGO8EBu6QP2gD0ZzJ1fe1YKndPd1bF8uLzY7fpw7XWpYO90sTSHxr7Fu+0vQHUsl
LVXb9LJumJpmR1UVxv0wfpmCUYLVGxq3RsFT5zEE3vDEjbaMa/LPCHkRHb00JxSg
OicoqVcTdtbw7YHEuvejCLuR4gWdmUM4MmORBn12Tfq/c9Jz6TysTGO8FsSymSbz
paHTHa09yskfvQzL6VN2GEp5kfWBg9YcpgXqxs9+r6fERyTLLwBI7357udn3JoHt
r0RnQg4/GknL6OuuKt82JMJQUOdNwuX8szxRkRpH1RZnxxMwPTQBqYCkggbEsSX+
C5Ke07AaToUQwrYpLBeZvkwFVTQ05UUwRzobfaHKd86lhxbh0CtKFmI7y8UWBycs
8KwMYwA7LudFgb6wI8B2EHvIk38C24XfPofaFGf62QOgstm1otnKUMP+zAD53WxA
5qzRc/ptIwGOFbZlxVlsLL5cRjOVniu/c4B98LWvtbVV0BYwFMKiv1Y8wjSj3B3k
JfyZVKM0s88dKbEXQV/UchTNqeh8/crwiA9x1yvU+Efv1Cq4YYOe3otnzVI3Jb17
e1hEBj+vlGrOISJhEemYjKyDfdncovbrZj386k10qPYEUljJjClblnpTNF98ifs8
1KF5oDF1/QIJFFezsFnxqONJZa7SN3pzKmBiaY9JBV8tWUgaSM7XSzoOd119l00C
ex4+88f1/5V5vgHdYxWtGNcninEQVIL5St4w/LFgU9WN+VV5/h02Wkd6Pav7Vl6E
1Qdh8sGz+3Q5dcmGnbHXjUqCozGRfBsdXPMjt4R5QaBIpXS9uyMh/VwAJqLozr/F
envxuyPfC4qEIRcGg9EvwAz1wL8iPc/hWPk7nMO7QlZuQJVqPxkrKfMnXBIukgMH
7C5y3bDl4b2B93IaMeB16aPjOdBptx5fAjyz/wLLh5/2oD0DLVLmdIrmwIjYLxNK
Hq2OfgYPD80lwtVn+lNyDQlVyTpRh5TMY+kaLzOZyMBwoNsdhqcNiLc8qao+HEY2
TuLzeWSi/ffLCOY+8b+UwWgjIcZX2qPPa6jGEbx7uINcBdYyf6zTaPi6upFSNoZM
Bsfrdl6wgjH69MZz/3vcuWokCDNcPCZNSQAQZLhU4k8UsyJBGdFkmTGf/vM6u1U3
W90GJmstbo+PMpAYaOl/GrhGCYnZvBAC1zWlsSyOq8Cwhj9+Rwjq1MPWeHNYN2ZQ
3Ux6lvNk0vpxVHJgCuLQ/xlHSvyOLzU7q+ODEYKTn357lyebe7YJH0jZH8ba3OTk
nxLZwSP5Xk1i/kA9DINiiFhfSB5ACrLghvkj+WV0mGbfJNvosXmKjLVuoVkGEJ3t
GebpymRqflSTRo+iCxiEGfmXnsiQvRdjzKMH29c8oGlmDOWxyxw/Z7eE3ZLjkry5
EDJ0z8JBGYGB8fVQb9sSAEJtDNufZVKX8tVRyLMuDzvAr7ffeJlR+qcniryP3P9+
HTvTsnti5j/KNdAWln+TbNfH4PRZGZf9kbxTstrfQejLtjyioFp5C7alFS25pLnP
X0R+n5MmkPh5nM7OqAtLsRoTkVe2FWH0WS/Y0O9CqBZ2QV3p3hXrNq78A72lgpiP
g0iPZ9TGwY9ACzzbTuUVw1fFwMI39OqT0QQVEr/7pgBIVnngWz/fxCZ5oka69qqa
HBlDUTP92NGk2xAvqwh7BcDBpb64phhnebFZmREu7AoXSO+B6jMD22Kx9L46dXY+
LVkfabi6lQZbQ/jtHWYEIjQS+YcsEAYIhlYTVFMVzaoXStxLqnrpOm0brM6mcWpz
WRIvKJ9U1Zu7ian47Iw5tIGeuLTiUf8ben0E+y7NOyZBDWYwimGzGs5cD7fFW73j
ODqmzAc7gsgub3zvEZxql1q9ia2aLVp1DxOw5Pu1kEp2HS2UMo25rtbI7qIPnNDJ
qeB/3HCCp3msTV4MXMxg9WrrY6tkyB2pzf4LpLVhAx3qYn2of7OVuhq76u8221Zf
7jtxcHoupQp138Bg/5BPxvuvIWhm108sV94eAO87D7Eylztohtxez80grGaDSZrL
etnxg4FzyPcmmYGkzgKsxESauQQaaKmA9CTNg5RDc8jSTwceOm3ocQeUSdXAdRaZ
h62Ud+saVw/6+CGWyu4Ox7qUM3A0QWywG+zbUwZwevGwxd5EBLTHA6PrnpTjx6Ry
bVhHtPPzNI+jCaJuL9wZOqblnsjhRTKnLj1ioDQaV2F2eAn18M7/UHh0bJ1iQJbF
VJFNXxhXeEClEKlvY8OZ2C07Qj80k45ZXceF7c9CdWMj71gg5SaN3ZNIDgUGA+TT
nIbiIBTOHKi+bSdTztR30TG8uIFL5r1/GtMdyhGZItybyNXxcjRNl9DJQWRCbInV
s4aX11fmrwh/oXWzdhc5uO2ICGxFR5Gb0mkKmT9P5G6D23RhXSqlsGsdNbafots1
t5v8H/S/Nodw9e+YpBK/dOwZ3piRYPjnYXt2klErda3Pqz71bH7GvGN/zgOqcOX+
L3M7xza8HCTfCVivobFI/TbTZVTDLGp1pHi0EJBIRCoJSPfIIB7x4ClBqEPNQCc5
1WF6HLOAXp6oZM2ot9J592rN1qT41xbtDP+TVLPKIdwbmABghsuVSe/yLC6YEYZq
mfKDw/++UccbQaykfqsWu9QF8HSUXt4XMf1zWrgAPKLusOhzPEgBFB4K1jIfwrYO
kpAN1oLa64EW2OoXn1pDFYe6NUD4WX8Q2VJxslxnl5KL3G9v5/KnuPghK8Xzm55s
H/OWmBwHGIUD/gRZTmXpIb3HU6cxh8ZlUPF3wiZ39xH0yoDPypwuDYainTFwGurr
Tidw5yUj/4K8aAKyJoA+K8MyMBZvJD4jAig44b9ctkyZGsCDfHi9xFS2+rBhj0NJ
IJ/k2osUPRFf9z5HibOM5c13TEJ0VqUDbq4Ent8V5q0ziTuCmqAtKJ7QPpevNyKc
9lqhfGPpwGoktdgyZ0KtuA5Vo4Jsu/C9KAxeLBc78nVhQEdvTcHfbtlvg+j4cgx5
FssnVnAz1T4+M1clnmuqqi+v3b7NQ4E9C9UwaQKPqFHH1GCI93cR66VLynV77C46
pI9aM5tsronMsjiIwOoMtxhiTQJbshGA4sB965SRavUTR8GhBJVzrYX19z92XlYB
jw3JjRJrtEeiFKHh3iTuli+Hg77pMe653xtsU4qby5ugi9TEyOKMpcGPVULN/k64
y+TGzF70t+QPGklVZEx/gJhlM0A7DL6keSup7Novnvo7zgeMlRVH88yMAscTOemI
oVvyiWYoI9KpahostcVD3vvp5pomDY8JikH/I2EJFQkVoYMcxxYxDkn2x4HNs2yk
Hs7M3PBkocdA1uZ0Rzck7FjlPahmz7/8JqZVfeM36DgjYSGS3WtdRObT+wiY21eS
FapiWAj/WiHy+MqrMEdYAUhUTzKFof3eR7oKVu7pgNoIefN5jXc6b56pUbpvTnIO
Z7DMSnP0wvfoOWg2JTdQLj3DqcZJ5i46tm8KVWnJN21bI89UewrGAlkmU+hv/D/l
ji9l514BVtsxZkywnw9MxRLpre5IVgTVMTLEUIEXMSDJEp1iDfrbybJqwt4PhbQK
mmufp4sUC1j48DdmW5sPtXcH06m/f1WaLBrFLgySgOsxWL+wAk5SuWzBRP/K6CAs
Dq7IhrXZIUzKe++XKee8n7crm6JEsCXJsQOq6EU7L6X9GcRlMLCT8fi1s2FqJfNL
XsScGRqK7zzAPHdXlg3WDi5xD0mkCyCfrBIAMD2QBLhoo7YTVXX3Ng0c+v8aCn9d
pJaOFgb6efULqiDN3qhPalODzYPtwKYGdVoYRuVMf5GArOd2omI9/UgMlHkicXqD
z7KSYmTbSLVyC1UZP04xPgJah941G8cDQORTNJsagxHwKHIQ599MXvq2kZvz/BWM
+GNbNwZZi3VMbtxKadaplo29Qz7Chtl7tXpO+GojWEtjUpPhtw8hRUI7Fo1Lk6u0
pmaTadB5mngFifBD2zmeyKaFxUgivPoWeYqgWJzBZr0SDsiDjl1Pa9W0BvZMSxbd
Ba6dsFRbonGIBajyoN9P4bUMLzT4ISbFnXLQ9j8R43GNXWsMHf6ypN8AEvOj1ih0
iLWr8Qn9/zexNRQC4mhqcoCkBtv6W3k5fbUFJwfHdOvSACNTpZZGwJo7oRQMOodX
w60KBNJ+RRs3YUmZlC9D4UNQngXaTEet98v0QR8I6uFGv4ODJwnRXi2VvI+Fs5+l
FtUymoaYqiB+iqDAffQWFnw2C6MY0a5jw58Uuv1mqcYO5fvFtHTGmZDCd+bUlUqX
kOjTa8i7TmACpq3mDPHUHjopCV79/hrn2FSAtt+VM/drm/I/BEbELhvKOtbTeuFh
H10wc4vUzDBhochR5P/9S6QRrWuziDGTfZqdqjz0XL8tYNHjkGARu7xhh3Fxetan
r9X0KOF1851lBoS8UmYwPX5rWPfkNEb+mjhd9EYTf32hEzMTa+vlkVqHhPNs5u+z
ZshXAhO9zK6qO3GMkuJAtiJLL6PQu7RyjUVbS49SwMF1bprx8UqKdDrG+gJyOWcQ
JwrjCjRnXY6CtBboU8r2q3L/MN4mJtEsSwBDz9ijazyS19w/e6wBCrJRGyJ/t6jL
C9D5w17uUHCzHYt+KEbiXpd8xvTXokpp6gtuDALSHTyB4VabHDZYDyu5B3Z+TDF7
A2F8+PilXuMAjTCWsP2hZ4tfqSeY7n4CnC6t6JeHuT5d+y4W6w/00DNGaOMa/gHX
OdxNY1b4N8i/MX0P03Zv2cbUgiC+ZUY8KIZEJ6DjEJdNEFWib9zgD+gFNGgHRxUH
K8tBLvFYa3q9D+UXEyrSGVbpq/lfziRFhncSUHLIK9FCTxT8AIxDCEmIrZNz0tbK
gw7PobBsmyPyGCF3QZxj0d82ZVeNBmpVsm5yJRu4CO5D5+Fg86eJ0aj0N3zTTvFQ
kGStPUcadK9Ongj/m5Ml6tm4ycZ2T8/YWXfBypOySc2UhoB7FCtPHgziR46C0l+u
NMxyS4Rfv29g1h4canwSVvLfR9OiB/dBrs2kxmJXi+teHCie2nnoifYODxn8tVgY
Y5Llz0BsFufGCx85u4UFUiIFqFUzDKL9pTsBIdj+qD8kLhJVOWZ65F/DTCUu/Hal
85PZohViVtpBAfwyZb6tRjbzOaXX3PLflruNeQJLweDk4ektRLV+o5rC8a88X5FH
LzvvPLsTko0FU5zcEaTsJQJWbq3eQ4hn5mDCRGI2O3yiPxqgLCdxLEJWbXNp1SVt
IwKtnhMlLoDX+BS1yQAY2GwgawlFyuNf0gU05bckQNLsQDwG3ApXd+EZb95pYQAS
PzhYG3gnQFOgXQywUU1Zp0kgXQ0Wqfx+tk00PVKFNU+OXmoOZbL0Luvcd51nE03X
xZeS2p37rdWVAITao8bvNmAezLKTvBp7OlRTbVfI3JQ+C6FY1e1NKrgGzgYCQTlA
NTTvU880vbYx0Djv92T3XjDwuBApIwwJsyUZlwY5HIBt+AnMqEaMZg8JnoxekNKL
wpfTlWoRk40QffXc/J0mBscXARnsHoik1Pv2toEtkTa/gAo0bROB0VBR2saH/jhS
oR8yoXsJ5c79B92uSui1A0abcgMfH3W35SDfquLcw4YMsAkP3mc6Czh2NW4ZUsAm
Is5Om0zYBmrfXF35DkKU8ueVGuyQRGrssyGU/xnxWByM5f3PvCuM4mVqtjw6d8xR
9i7luLu0uvqk2MLa/VM7h4Kx3nCwhhe+V/MsGpnbzap2pjeG9JobxlUo4WCSmT9m
G+2WFSphfRSzOmDvn3ktZEjNLCX9ItzSu+uxKorI4glTqvtz8p82w98xWVWsGah+
X7vO8PLUYkqEyyE6GZ/VDDhTiH+wbZyAZP9wi1U3DfunEJspp27X6I6hK0i2AQB0
6iM8fPOj4folGE8DYpIpw5kItmcs+4H9FLhMoIrJiHtwERS/NziwZ5fKpV3bxZfz
8cOEq63W62jrl89bbkFnoBDyIUnxzh+hymKVkUb4FNnD9RkoppWFI8Rs61WlHfsk
I2Yb7EdKVpP8OTipDhb2Y1vp0n6w98nG7du0fppp60RUqyfPoeeb1pTX0Bb6j6JG
CK1sC/ny/+dn1X33KlCn5BorJWccbEJz8PEDWg/LsOlrmVOEunaruqwt8v215EjT
dRqbeK7Bl6DALP0eytDHK9TNqy7azGC4NaZ6Nb7PcSJyzKdXzUXswOux0HyE6lwD
xvi5mycAaKE/QeVU5Tg71SxwUEnXMPyJn0EO88EgkMIHeoOW47Th0dfuZ0AqL0/f
TlggSNAIk6un3jE3xwaRhVcThNKomxd+wRUEE3QOtIOXqXG9bfEjAnPBLpWPtofq
lmK42dYSd9pd3AZeAT6qH44jiZqVoZ6L6hG6q/D9aauMTp2YjtlhE6fKtSeYALC5
qLpMkUkfYcV+tR8NlEDwF/HJ8tcacqNPM7VmR3mrcLpcQEgyjbaQJJCON8dp7zv/
8z3COc0ePq9XjOizu9foYJWUI4ZKIy20ae6CYp5jClqWjf94HwuZKUACRut7Hl2a
S3wYSE0GrKKaQYPRFm3a0uqO7PpU0Ow6FEL25upk9yI3rr9NvTnDkPXfiemKRe86
Rj4kRpj7pk5unWixIgRsoz//sjnLE1kBjxOiMCLNrewgyovW3zs/95yitzFtY2fO
e+xm4/TUdi1Z7Eo2xIj6GX5mn81Xjork1lMv+Tz9NDEePhCa9zSy5ThvJ87iyBMe
UEZAxXmlVnQBgbDRVwXWzkZ9cc7rTKk51cbwHz7BoB0LoVg/lJeYMo43sr+XZp/+
8Fprd35CRzDcgc6J704qIMU7bfEdFp5ewbl5KJfX5lqbBIFJUsjUZ263uzKYCca8
IB/NE7vhWZIdWHCv+DkJRxwtyv1NouXcpQ4gMr4Omacz7Enh2+IZEDFj53DDFyX2
mhmJFq31LwQANu+8KeyKc9Rs3zuxxIDypDrllVVQbwahohdDGKLE5iohTFcAL8v6
450xJHXGinnldnJsY7L/e2DR4SMpWOyp8czFLoDCQAII2KP8q+gRL4ea8oDrasUu
/ed9v81vko5t9B+iJH9FiEgqsaw/762mzJgnIKsrFSRzFHPGEhfgYZvsiVBxOeSc
SrTMhgJSUu1/t3c3CK/3KvZ2p7QN+a5ySRLAmm00W7C2XzIUq/NpxEqG6BNchmFF
Ok7JHt1+AgnSYmPTEHRHU+5vSEGP62oQ/VF3sRFU4h0Dptzxxp5aUOSyr5k5/U0+
5LHd7fj2vO4UestJROb0ubBA45G25ohg6F4I/yVTJ0IsiOGcy61sSOUJcu80nQJq
BNqUtuI33je8TeIKbZAtnDl8kp/juYSYUolnFN9CgQliaN9w+q+MgnnppB5byk+N
Z7yUVQftfEnvGyHDTa98YXAUUnyxKBQNHYYAlgE5cm2IXayguehiUJ0uUTLJbKPe
BgZeUKaeo5VvT3KtUfRmWCKe4B5o1okHG8fGnHyAI0TFYFEtlGdpPG0vMlS2lRSs
4FkKuK6Nu/akJyaC2KNibg84DItznCNFwNHpPq6LPY53M96+x2a8X5b3ARohC4xI
35zwh1RqUgMv+eHc/Rdk/dC9pii5FZHQ7hA/slc5O7y7Nc9W1gebIjflRDvj1GfY
46mlefFSYJmQ8dWcuiG+0W+p4TftoyGLGLYDtZRfsu8rJXvSBSC4vqXS+dqTaHAm
KKRAxp/tYuLgLgseZ8gpaMtzB+YyT+/O+ebsPBmfrKyrMNwegY62+Hm8Vehi3gpA
jZ7oQNi9OuyZv4XG0g9IBeU7QyforQI368JQV80X3PkD3nQsauPgGx1zr8Y8U6rh
9kFCAYs4xJLPzMuqKctvoDphA5oEnKJ7By2uyr30vVL4jH1AemwsA6QSk3qKOnrb
sEX3yi0Oo7yeX5ZPeyRhFCoYeZPvgGmtpJ+xmFGBJXmavdncFtSAsEdvw5DR1sLF
RNfUaRp2Snpg5CX+YLWnhp16CoKzTheYUMElZAQP4vW4W3ITOqTnTaVCXFfHDou2
/acFO6+p76hxzp+FSnGm0jU4qbR6pAFmKcDAhjTOYGZUPS0gS8g+IX49AIR+OV8j
gJdb33Xa7pA0qqNIn+CmLTj3pLv5rmuMBbhDGLuh6dbLf6AhvRfrdPy3DbXf+PrR
GNFyq8N+UUw4a4zrzArpX1mf1ZFbOL2+4OWw0Hn4xqw7uJydN4MiRgNtTRl+BCLp
HmD7gLhqiZ+MwriOYyE5vV6n5juf8EFRcR6Q3gzuQVdXURq0uhMX2lqfdzDSnXAw
ucS+n75ASexzZwQOZBIuB6aK87WRE82y+i6RnREJ/qj8WBrWT2Xmjke2oI+rict0
lfU9loI3WMj5EIOMArXXhx6CWHxLTWq25tZJ0Y6DKU9yre88AwoCCdj5cIJiLmYX
ek8KkajVVbWSGcmIppuD8Gh3ViVCUxieleesJjNOxscGri40aRkFu+CfkBuX56/a
S5w/vypPLSI/xH/Oh23Uv58CLSfo5jqup7VLeOd4aiygc8t7ANvD0REEZ4o+cbxu
cLh71OvbbH9oNb7i8NqyJ000QJOi+yQ68recoVr7fEkC8bu0I4XFw+yCNe8gwCdq
tYpx6sbAqWQxV2ewlBU5YinZACe1xDJ0BElBbq+pwX5JU5leaW8LQK4cdcRFkxfK
8FDdpf9/5pLZqZpUYf4n4DBmdhXsUb3ihFFEMSfGqx52jkw4O696wA69lBndfBWD
6Czg9Dd/z2k46YzoF6SzMYLojgJSVquKTKGnO0WhgKFjn1lyV4uuVE7ktV/u2dz8
O30R22h8kYUF+B1j3I9epAsv29GAW15wdYmUNEWo4U8Uibw0GQRs71+TEJ/8T4vM
elWLygJ586bpow008JOTDK9XvM0tAZu/YA9e/1/yVoCJlK1FLYVR9TA4ItBYjZ02
bFmTlRW6KdHFu5NA0B1pRLsytqoF88ocJ5p226r8hUODTtK22hs3CG1jmpQklcee
UeyorwRFHxuGpIBT9BnRrOJfZ5Ga1Tm5g3yg+xk7B5SoH9G//JzKxWYEWMW4ZFHB
SkW4Bazmj118GYRNfRqjTWfiquglBM2tS18t1C1bJl/wZYjD/33hmgYx8raAqYWF
ij3d3q+zammGvfQzR9bwMlU3ZiQoo2fRRxmjMfXCzKN3m17x5HebS/OgTRpNHqSD
F6SCx5RvbYckPb/3Fu4GxzQotylkvJiQxkJTnnYiVxgH4O7EMcIHmCMBV2rsFYrp
+kAKQzqfyB/ohMmSi0QwgiVqaMWFGrniMjZbFJGhYhv5s1xgNUwqTAdGjHHNPNSQ
bUC6IPpj4FbF1S8XZi6bHCOl/fQ9M07H8i+NH7xbSYi1fVL8qFpm+VmTK9Ia0Cph
yNZSNHzQPW8zSGIWlqehqNNh1TEv/kzdtI1DJNsDX2jFvK/gH813fEMr/TExe225
w0Qn59H7LMgQovhLSHmO3KLn5u0SOh+u4QW6hfdlxWJFY4VuTwoRmHAc70waJoJ1
OqUNMZxpukifof4QNzMnbXhmmkoAGfPMnXc3387bTOz83ndv1b2RKDAAI4lEa+9C
vG68Iipv38Lica0qRyInI8etnYfsLgTNPosTCkXTtUF1icBZOgkgV1Eu4TdfrnFp
M8tRRvjCtPnEXNhkJHjl0SNPC83CwdhPUe43lR9lVRR9/arJuktzH5WnoSgBZrkg
t5k2uApFVKj8f2YX6uIgBUDETkxC/clDLPGXmGEfQHdPRNoe341v/8b7B+3jYy8J
R+3uS1joVNZkfCNS8Z+oGkzXu2DTbcuisog65M/uPyJ2NaB1QyQzIGjhm61VTuC0
2DPf8L3sGoZKrzUEAYlUCzFBedRjw5Bl59TA4xLQqsVSm8XEeEGTTscSXxyMYm2T
Maket2alSE+WisRr76Roi0HY8s1ePkO25XyyH0vslok+HDKiRY8Lz+CPPqy938uU
7sGqJEuf2nrX4HxryzpMdln3LpMFxt8UqeV9Q5XijOPr11J99Xp3M/pFRs6ZVryQ
EYW5YnKpAX0Sll6fyUlJBODL0fo15v1qLJaBNu4sqzq0x6T/jV+ZS4mr0Ynmh3Ak
omA82usaHv6/Twh++AmZ8ltn3d4F5iMwoHrtlNzwOyWIxzPr8ulftByNVwgtqeYU
K9mrNHgQmGa3rT2mZfFxZLKkhBi5IL9toQnfr70i0dkVI2MA8hsjNeAMokeVZmaw
xmHGImFuZWaJyi1nvC1tvQYHuVQk5A8I4k1JMOu0Bi7xSdFaXwslwttgd1eddmFR
W98Z4Zpzza2H/jVskDHGKXm+8ZUv42ekJjqrxRjJzmWaYZg1mCxz1O116twTsep8
hqHGw2ZMluonaydnrwpNIlJL86laK54Y23e3wG4Tt4Sn9LJAjAYbPOYHViWzaqca
7EBYi9FCvvuZ0Ef5Rs/TC1J8uEGh3Xfr8uuJFjQASvqOLMgIvZnCHHnDtbAVgZ+U
Xan9TqgnO+SsW9dR/m3AWwwvZFNgebickgeaz0hsgOwh0CHjFEqqaaicYvUKfrYA
NT0usDjwSbdcv5NvNcSLGSaxdD2/IDYa9AEwrhZdDQsY29I1gaytea+kiWfPWPfT
pwZFDIZ5cYBu6IdxDGiVyEKue0csNRrhtDKb/9YS6jXtiPsAnalLgm9zDNIft29z
I28LrpmTPj/rpObmrIwSRzP8EWu+doXzSapjohQVP50gjy5KrfR4gcRmjOPlL3sx
WE876ENA9uv/KbFNzCfCM1mW/dIsfu8ZFb7pqf6jWT2oq4irV97I+XIazEvRF5Nn
257JhW5QCoNKpDe5H8/tU16TNrKRF6JxbsV/v8wPqcmvYYtUaC1YYcaRvrq7IPBF
7G4tDZ5uXR9QTF1oQtuklbJhzOS4tpI+Hc9qJdN8zxkKWGZ/M8vwLnfwoD53m2nx
HSd2MOGmJOY2KS6ghSKzCPelwoBvl0KoX2vmaChguu6Ub0JMi5lzRWkFWrAmtV0O
LbQQPYaeFmxbuvOz0XFx/KlL51n8Qy96y12sFSoq0Z10ch3Z+04C+H+YEymBUggz
q+eWaKEXxW5OWDW0eKqyj/QKCGv9aW/kIqYfLX+Ezc1LQoOx+L+D+HolJtjXhb+6
F0bngemm/zo3wMoEJ1nG7tod/FUigI5FXq9iVzcESZS/UzwOcN/F7XrGDFqj6FE7
mgXotm/3G5Fg2jTfeiL8FzEqabkDr9hY5SzqV588Yhe83M8tphfdO8WuxjV/dYBk
urTpQCvgRHGeoSaXi67xWdPaN58dpTKwSnNbiWb1Tq89Y+JDTxKLF3DOLaPJE2ak
IHGBgDRwAWkNNiUfLIHGXPL+qR8mBC0E/yAZvfM+0Ka8lEF8QBatmPIjW8dlZNuJ
++1MmZkuwGe07zKQGDt061+sAOQejLcTm//4UYBNV9CvhdnQ0Ul2s0oEmZtrRH0B
6tkbHjNN+lpm+RdGdYuxAXe9fVSk3gFZkrFkPuBhHzLWPa/rOYtjc7Vh+IBAenoy
LKMi7MpTEGsyv2uhoVFvo948P06yIsf9jUgSUUTtGIgVtVpaODgo7aRVR+xzpvCY
dsEG2kL89TjB0cMd5DfmxLvirICeXU/JHSucK9bbGJ9TArrDGC7PEcwxmOkf6jhe
+5EaphhizFxny35XA7uqKjMXIofR79jHMMFaJRLbBbo0x4Pt76sOrfSLkNvWOmoW
wtp3nmeTSkM0BZV8TEvjP69bk63+QC2vm6lE7qILFiNUQTkP3TRpgmCvXxE3Ykl0
kzblnSaTSRUWfgwW4ZVOGQF0JnAWmmgwBavea5MfXOi+neawjGy/86dFvNAIRliA
h8Ir5Bc+JhkEjgRKm9GFCvaHFzWnWiY0+qIW5rY7WbyPNmRKwbH8fM/OMLfOFQwV
b66Q/UY3OfxhknjY3RLBoBRHNFqoubYRyLpBVyVQK+RzU2gusmpMBMvc8niKsQkf
pvVTYP6G7P9vo/AYDawPGlb3mQnS7H7d8+Vsvu5uDQAlG8u3TzdVKi6rBp0V6uJk
w3hYEHb0Tysj0YUoJGqvHqX4kiPtmUTNUQfzP6F5TthYzPJnKWO68jVhIR3kJ64D
m9L1BUTo2DRh2ff5cQ4Rf5IUn3BHLKftwL/M037h3i3wYXSlM4QbcpvPferELWlL
CAASN8bMUI5Z1c4D0vsGiL3O3HA9J2rmb06IW2PPZuPoOCedmwIELXXDEGVjgQ5J
EYkc76KvfJLii9/zHigOGr/q7GipefD1kSStJN92OKU4AqpH/pBU7jEoep6oaOcU
CNErUM9NDfi56niniECyg6h6q5h2pK1wyCGnhEJK2yNNbx//zs1pEvzrUki0JJ2V
ajKWGx34UmD9LfQMd9cwCfkc2haSrEBbicxf1NqzP+FttRShgBPwCCpvPgjJIZ6O
whceTX0eICeIrhVtPjCOwi3QNmWgBllZOZkapfxhV+wCqKwXRwL92093WJlTvM1s
UQLD1xeU6aSWyn7/Sk1bYW1U2Z4bjhMd2tsl+z7P4+uC5o0v4Ezx4JzubpQPir7I
0BczEie2pxtpc9C3gvLZPq4o2xxGZ5R2GwA4L/ufk0Sksq9QORIXehftecGaFaxG
4MIK/L6qg6v1D3nWwy9N4Vgrl4It/PDetoIGihIUAZaUk4784ImIqSAGX9jRUuev
Wuwe2+Ad1YSBl1Z7TRXi9IKmqtfZAoA0cN5an+b56qeGeg935edYimyLlOg5LdC7
FKd7Xep1FgIw9SHcTwv8qEqYhIAHmzAK2vaWmq+fe8sEIyMJ2QueorerA0IJjMP2
uGbgzctZ86wGKy1WuDsAjo8Sezp4adBLjW6XZ9VP3XsFaxoOMJRVqdZ77BR3NRoh
YZDPkuU9QaZQUGiEoIPF9h5Mtg0k7nrNowb6k0GMqiVJholo+Nby/mZqcoJfDUgn
BW3HF+DPawMdbc61A+nCNPkk3lqpxpfOBsZ9ummyk7UPNTa2jZ6/FlhANqNabslf
/bR/fOPRXzMIhA/9mUOpLWytMGqu2WWIaWZr6YAYkZWiDTeat8wgGEj5QHwBd/KX
6ldMvSTOJOlW8oebCuuoANuri23b6GjrOupAXErEmg8FQApfuoVnS17FEBDAngY/
/tCp3NdHs4rjgxm2NHrKgZmIRL9xD0KYv4CVSMUgjIKm26ET23YOWzuJJ3bGMdo6
HctU6uLbsxoMuJ5YULNd9AuoIXL2HYsJxqYQx3Jvqd2qvzr6nLRREr1FY43LBKcT
QIvIGSX2kb9L/i/JOb/Iz4N+0KWaM9vOcLh14Ul3BC8fv2qEERUJJcBsXUYsKhFF
dsVaFXXbS3A/q4/U/SH1TvuhHBFnLP3btojpxaCcChnSDws/o8w3J7my8zn8/G/d
crmVrry8/lqJ9cjsJGylGr4akqCo+VK/25S2lRCK8sdDR4sHMFow23sTy3KSbv92
a3U1VJAnfwD7mVpI4sRypoYD75A4NcdF+14AN048DCWJCPee5DRCJjzamvvEjckK
BTWtM0PrA1NXw2FzNsGycyD3JTd8WDva+QP9VZnrikVYSf9+s3xd2AEl4e7C1mZV
CavNElk02yxsxrb6Rp9bEOVLaU0YT7WzTmxCufnMGf5aNpHh5JtCGzPOfQZ6hZ6B
BP+98ZlwisFZUun41qBmuswtLwZh2wBIgYpexx97NYo4RogG616pqb/izUYpjOLR
lrjhUWjmyoZdPCWWuQk3tR4wbrUrnGzsIdiTcME07IzHFPInuAN5PPcv0Kmmjdb1
PZFShu0hReNUmD2TRiMv5J+o8A2l05J5GdNn3QhUIiMvs7mBzR8x9Vx6Y1LySMUW
tMV2IT25a5jlX6wyXaJtM9RM3HphiS8S6Aa75DEpok+GfjGOZkPqq4v8mGWDskvI
p9HFzZzZzI77ZRWOw1gkgKDjzaNK+kxrvh5dtIyQnlksaAciuQPf7rHKyDrt44oW
KTQJSWX0hX2ksyiOEsceZYMi+qCJRiGCKIZ0i2rLMFDnuYITfi4xxwGNAkn6NafG
fULD1j6+TiQKE2Du3VVgevSDJD0+V6jnMiCkgEiyLQTEoooOSPjjJuW64zfbw3bJ
OTZaPVld8/30/Qbj/czh2jY3S5jg2M9d48EYXQ4TS/M/eA7pQh86nC9X//zSCC3s
YP8LYPxG4tpjAj6B/yh52okSWNjjpcol/BUexQLI0DsFqOYjKaJlUWcXUjZwQf/O
z4758kozK6xHM+VNnldPOexE17ejfL+TL/2BtMjsv3IVmzVOlsHHnmwIAPTdhp5T
OfaqtpcIfp4f1jCaiBQgrHzLXykRXGaEq/SwDqyJvPZ5Mu+xtwcfm3dUt1VyD7Sl
dIrzE+FikY8MKIO05xvNYOaeV6h8bXskRCCUq+PV3yhtzsf1VorpR6DUyqY0lGlu
En8sLejv29TvYRPdzNhfKLqVF5ZNv8bIG7pQ34KHORQ6TvgzHDXQ9aDNm/fEU3PY
EGinVOZOm9sebcFuKmH/kkFVkj38AiOFQVi0Kg4bFqWnutd1lI+eVsS6otFdk2vA
Q3g//x8oAP2ZcvnI1p/U/iWHwmuFVl96m7VqM1bD/eqZQdjC8hE87qJ/nNHn3pT4
juOq+V0tNHiqMYKGElvBKEVJGvSlMh9Y6Re7I9XT/xyqv0QbhDvEGa6i2zlNGkOz
SAVcegWahdt7oNgdwbTWz2jL3v1Op9/U9qY2Uj/SMatsoKONPrdngXwsLsGE24Pb
L4tNwulJgmn8KPE8nU8IDxzQzI3n3SnrgaABrjeIEilA/YUMdftHORAh1q1s6zxS
6b8PsdkMmYzpIUv2Q8zMhP+hQ12kLUfWxH/RZCsydq1VerlLYWubKQ+uaqoILw4E
2ckmh8J3LuYRDvMw51I/FafPbaTybiGVsRauSrQ8hEAAu+mLY424c12QqT52PmS2
AnzNa5qnDnr0FsAoalC7uwt02dLZ/ZQq1TeKBkepWCRS4o427Y4Ie+7jDMWc7jdh
kp4e8ArCGZloCWyX1ePJ+0GHKOQO+H2eMx5/bzCjCe3C9D1NbJFR6g9EVJP17101
aDYmGsYOGyU92WxZ+SvapdQcKLIO0M4CfcYhoS3Qajuiv9ZXULHCVdN7qSzcxPky
HuPRcIMv/2exrUTIJb5oWPjefc12h8h8//uLUrS1Fof8ydTohvjjs7ZQ1N/Q49Hy
r7VsnUwjdr0HgUyFE03YqEFZ3M0Umm7J5y1shYreL5tARlhji/snTociV8rit21w
i+M1VUM45ZuMxZqAtOWr0MApIBIBT6RP7cQiAxWsEtK3nH3KO03tTqQfVkq/qzA5
/UcTRqYrollskGi8BFxmL+EJBh2swtb6gLoYUmHaMt7Pq8rN4v25H9XV8HsNMeUg
9Kk+ArNZRtkqq6gvtsKCnZ1V+7ntVXpnozDXMH1hONsNpNqp619mZwIbV8Yg4VS2
3WEegKLV+vC3NLm6lbucYuR2NAt2ZziEyzVD6ryG5Q3qxl+GnSMqec8M2rpxsUtU
cLK5kw6A72R7lwVUAZzB6Z2OlnEZuQ+4Tj+bGVtFXrjjUyqGmURFtyVW8dMbV8Qm
fc90Psbn5w3/AEcS2We8Zcy0WplY8iZHE/L1Mvz8Gk1kn2Cuy0cPoWZdUaHLT/0I
nJKuRsZOKz+vcrYWv3crZhCUiIGVfh1X1Tp5714VqdCiHXEQt4Bn0sSA1p4xn9wZ
KnmLF8bLoIrO5ERlMKLdvqaCRyQQb2W2PXaJmwB4M/k5mu7kFvN2HzoykVn9nl4r
QTKlamPeCXWZV55xW0VZ/ZrU6vXIhRhmVf7Wq6+oyPpJFM5dpcjPCPr2fwfKuv9Q
hEGYft2ZTqcgt/q1++JTiSWqwwQYiT9p+n3wx+4SebOXcfr/F6KnHLEVhelQHQ2E
0BLU6PIalK4VbJLy67eWPKn8i2136CmDai3gRqCB5HqEDBdpXiSQ2/DHV2C+Oz6c
pzYpABfBk3dVxyuQ2rUVcsWlYrRKZ9oXn3D05BbpyjbfnnSEDAI3HITjcYiyUeyN
av8rnmukcV01XAaRTogVPo4yGLWkBdOoWwfeFePcfyRMEBB8+/odNk61YVntUUA1
PtvpZzguWjPQR8i4pJwc6r/UUV6RZlgqd57D2JJu56YKNhyuTIyne1npIDI+GRmy
0+YE6eVURXB4fv1eldw5RZ8eX5Q7MeoFTtUfj23DFMUsTq3zFvQ38jorpodv0eI2
CD0EkegGx2ENQ3oRm4AS79g0j6LZFN71EkiUS9g7Y4YFINSmiKXBZiGfJ/0gW7Hd
FHhgOukiQP6/Kz3di+YkmAXeoY0QGQjvJ+8cH0YOlz2DEO2Li9unHYfJ3phdpACt
4MxYaRpOclSd1GkigKVnNfjPdTj2AkliYuYZWTRT5/bknUe3TZkNxOkrdJ0LvA/F
nJaCRpFTqEC7YXb10utqhc+EpckPevpgux2926Z7/xM3soDPYk08WQfbo8UNBtsD
rO1TJ5DRsmoLE0j7DaQwHbdqqfQ+3VI7wE4SND5DRTIeeqL62qmL41dq4Rnd3i9W
/Bj0c+6smiol7cBMgeb49R2BYukWYEK2HTKfos166D20yPkVgAijvMYRpMkejW9n
bDzE9eriZ/Ib9WtqHPw/UlJJ9WWQvwZE5m4mSZqiCVFU5lfb3DTE3A1j/wbQHnHu
zEgryKOv55fvvM2EVOfKS19+E9yL9vwZkmlHmDzQEzrHWxlVqFFNCRSynkrPic9E
PYHn/8LH2pdlLg+hIyWu8nM4Dt0dm0DQL9Jqq1uDSRj+5B0xkHxQ7foXfJhQSe9q
2H9czIr0dgt5cSATSmpbMtvoiNTbb05v277PlmxSXjL+31SXY4MeZuVi/WgIFAMA
ygUyvBhUQyX2SMPfCX9dQc350QwY3J1UDDeYaPIct66+g9Sg0FK6dACoxleFCrQp
BstKynpC4Mcr+9w2suGrKtQ7X/1A0yutaxMyXIlF3IwQcVbQjQFWoVgovOEOMhOO
4uM3h7j1QFeEzh7I4ZR8W+LYiFWLyTOFdfOcz2uR/7aL23WBd/bfyhmma9GRkq9S
tBzdo7m72yFrZ3x0D9GP8YPdOUr6ie6JRpCx23RxccFXCQaBDSRq7nQzylriOCkq
h3UXbovkXNgcXbcOLGCx6LZi6JqUvkwNafPgyOSwLqgfmtBXltwy8bqrwUNm02cw
KEOrpZ6tHp8319gkhOdaQphgJQsX1YrRi1RwH5lFBHCYQr7W/pFCzjr2hskggGMD
Ro5E8qN4Ow+v1rtfL9XOuUUMFxZMcoWg99PD1xBb6PAKBnhD23o1w5D5kYIyFxWV
FcUBYTnt7PunyxStTjWQobRuY5PU9Qyf73vK5iQdXzRKYrl0iQuDZXAPJpH9SWQ+
gYZqDiRGHHMlnklldcA0H40ihxugjEZQRZZodUgZuUU7Gs3qyVWrCT01e0nc2zeF
9TcYlAfAqahOhFIIdxyEz2QwIcOpNuO7LLEZvL0KV7mz1g1I1Pv7EkCjbJA33tae
t3Zuoyxs8eVL8dwmvkLoAh1WaOe/cJ2izhrTb069xXbaCXR5HHIz/GCBfSgMmfWC
fhXnazvxsYfPhcxR5fPWT8IejrVIU9pxoy6dgyOunZeUpgPHZd5qB0a4o9IQQ0ju
XtyxTL6W+dqWEOuPXhvO8K2htlS9inq3Z5CUuLXaouDbpV7hceDDBwxn5OrjNbri
1v2n6BMZRNTiFPRGvqchZ38WnzyJCJntvSUNG/RsXsdwecgcCaH1MopQw7XAGKRU
6OGHnBVcK2SIxoRjslN9g2RHOUBRTAyhEGDFPP3W31I0sjknqkcYT1Gbcks8QGCE
WhC0UJSoSV7YtlioGiC0aEgb2fo5TDgIrg9d+Jjcc5NZJ9dvwfRmL10pEe0EspED
l748q7LhJzU7D8MahZpMHwOZMiRDbbIxF7vouCCjkiK1Jg6eLAZCrmF+i4Nx1/A8
89hz+/mFMjwy+lSKVx+SZ8BNlUF3odDF4hgjtMQi2nPZwTmTVc5/8qPgaLoeh0JZ
YG6iEFl3x69ifFtO66+KNsHIv2CVMPI3xn05kZSH64+lYAC1Nbm277efo+amsPg2
izWpcW8Hl0cfU0FCHWdCndt3ZrmfgAXWCuOGV7kZ5phacn5x8zYZslwasWP+9FNa
MudAmBtWq2EdIsol0iYDsc86Vw4hvRkPyRgkvFc/GM26pU+IswmLh/RJFu1+Vyr5
CB1H5CutNtkpoiNHDimNfbjOlrARSyBYVgb9kfrBewoo9R3Dag3exteNwOpZLX5u
XPwlTW8whF4xyttEF0VxAVuRTXdrR29P4imnfDxyYH7AHF8jUck+TUFBpp97fPsi
DlBaZJ/VZR53PF5lQMCfrMK/tinu+te+dI/rvfeZjKxm/KQVVSydkFegk+o1uH2p
+9Ztac9sCFicRSw3DqCUyFqE0LB+7Jq+edwwFaQ+/1scuyL5v6eoxlt09hEus4TB
zQnFB/jEQu3AVk1nCZuuGziG3AC03dBZxbYNwkjjBOxKpyyuOCb3aaF6nN+0suSZ
Fq8wu78sVFxjVZks9cpuhd9lseSFQdc51u6YonoWjJsYrTBl8FBoA7D5m2MEDitj
RFrT/rBGprmkQ9J0nJKfIveyu5Mm6Z9suNhE10JB/Q6Vb2wlhqM37cm9VCh0QRFi
4XnGVjhm5PiIGGZiVY3G1Pp7kGh9yf4Jww6+BZe7pknsvheJVWbBLSKsTGJ5jkvV
HzPwUZVpnwv0xizD642DDFxCez9aLkhg5vrygEdGmrLY650KSnXUsnwLHWJQAaIc
lP9Kcob6SPXaSrKHyx80zaJo3uJuK0jcGFIwWt9KmokeNdJsbrQIALFfn5iTYDs3
pisv37QeBreIxsQXr6dwM0yN/AMMBC7B/mGPAT/LUGEoLWRxEGvlT6ytVjHWnlFX
u2nu9/jZT/rpzFvQuNuV8vPQEl0a0Vh7UoHoup3I/Ld7e+MCBK5fdzdgiDsfdMvl
PlEPOzv8WJPUCDyz41b26EcnB+5CX3FsKUwzZbdYPAte4wH2hbGht49widw3hA0C
MiSC9sR3BWkQExC9nSHqXIva+Y4jW8J3G7l5Nrf40fdUf0QpakVTdzKvzf/wtGck
ilMcMlpvzN/FocaMm2Xl4UW7UST63CLQPtHnxbvLZZ+pxaduTXBAM+oGZtz9vu17
mFW9H+ZBUEamz5049bW92G46MinPuZkiKQUVri/zh2oY5qNzNvelpe+36dOVcB83
D+2w0oJOBzYhpNu0P97ihrmZAjR6pY9pMWV4dvywpu+Tij2O6tNInq4ZqACLScvE
NfLsragKs1KmcSHmFyCY2AQgk0ohy7voIBO/Q7GTxRruxkKpPN5buLcjsJzEw9U0
egit02+Y6MitSvalZuDukaxEnzCpRYwGjneesDe7dZ1+RQQMrW5qZfnBQ7mZSRwa
zp+F0FYTov9ngvp73LrbtpThBPTPA9J4sHpZcgt3Mu+3SuFeFb/kfStCILe7ddym
HRWlSEZSoAMiFmjFLSANRY7jKsM6TVDAcD8xzEXBMHzfZMn2cmA9lC7QzRsXpoep
fvV4msk9RpVAjvUB7+zTUv/5rOXCIChWNESq5owDBpEA0TZOherUaHiCM1He6OVJ
aJJ31i+J7UN92cGNOBPYp72p2NkRmPqeeIDrS4PA5rjNmaDXoi09+UuL0YUZiIIp
Lcl85PzgR2Cki5E0f9SgQvm1dNJaFWs5lz5s2VADW7PDqG++fjyuUEYJSS2HQzvg
X4PRJJfdIDYzCHac4gy0YXse2QjxaC74de1Z6j/kyA7I30lpfBL5aG5iJ9FsSstL
QyrCdDci/6QkiQgAY8HlQdVsmxp6/As2nlFaVlNEL/AZCBvMdu6oVrj9ACMXWK44
VpAJ5j0tUSQKHMnreSNh0G8ufqkDXlkIkBAutitnBa/qkyfycqkTHx+wp6uN1PWH
Hz+cRM0ZwaDBLyGSrK8lFcN0UNLMNU2AhhelrMre0BFeY4gltMWkDd7N1IPzVa7J
XcEaj52AzYWK7i0c3FzRPqm430kYoEM16HeMyWQrG2UQD618C+Y6iRg1clOvtloS
+vDZPHXxAK1Ev7BHE9w6stzvIWnAnL5sbDHHV1m0CHpK/zzLpdQmrj6iP020SRSz
je1UIXLdj4+adQe7ybhafOBW0PjmxFjIi2mIAQJlXpUE7niaJRep0jEfZ173/xz4
cbVEU2BLKcdhWi9VWP06L6HgwXp0TzbrGKv2Ev66exh/m6+YRy0SCvV6Fb80ECMA
jxPSuZofnWyb0n+BX90/cHScSt9SmMJVaRndCESyO9Ky3Xle9k+Y8fSWr64EoyoI
oKOEMd9yloHsYiHLGrpdFi1xtma81hhWFfgIhUJbDY1SmG2Wt4H0+YORIhawOnhB
oNHRl/bYCjTh1Eb5P8+vv0prjqZcCN/CW+0cbQ7fZ1Hd7G4VE9mvgKWAuWmPdmgn
RA68UsDnxkRUVRhazt6S6BmFVgwflhPiYcMLa7lIl/Ku+D+FXl1jmiSXePmpe9k6
KmJTe/S8b75qsENbjA8wuaFfXHg4oaeZogd0txpxHTV8dtugLx/N4Qftq933WEWD
+bRoXKhWDYXOVtgKvzvMFuAl+whngUgnLVgDIwz/Q0/ZxiFHowQYIAgOLGSP7kP8
6i4iImMLt80ELQrCiP4mZBEYvKcRJJDjU95kYCON99LK1aZaWmS3lWhRfJQJLa56
jNL4o4oTKaAQeyNIjWhXMHZtZhEB7EDm9AxTdRrmd+tZpTRADxz0P+mEGDt5kovo
txgjaLYkU3hiJYmsjxAXTyUc2mJcuA35IdMeRgOOtd0KgjxoBDsfYkmim6/j8Ur+
lEX5rednbZ1OMwZyP3RjPKdQFpe4Jv7EboWaM/aLkuG7QgH7XLDAvwTG4TZJJiy7
/DtVlpF+g54FR7hR72GQVDx5+1VJZHu7yhzJStvNX6hS8oJkiUYNEexwxyi6Rxug
gtOyCDe9TefPhQvJcrqSyu6fsKeG/gbnMAaIQBlw3F8K4fT98R77Ry3ERKP81Olu
WD+abhhfOtWHUYBkIeD6O9lSZahzyjdDdltR1AfKovolMO4Y9EheOyDrOP8nMxZB
gRXfKDfQubyBjVahrSdB2IlNaiKcPyik/gOKVj5SowLX1YCPbbfW7zDCLThYAZNg
DQ2DrDlxrOJ+ImJwgD75OMXQVZdrDfbtCIRm+myF88T9dP2AJFLpkaEalKqbmlpd
fUHBMrN98YZ4h5yx0gfNxqcopIPkVExTtfnAmeqoClRNSrKdS7R4ygzrcGeyiQPv
cXfinpxLLsVDkWB7z1S5iB0etwWaMvmnZl3SAyhUTPZ3gfSGEUmXJTA/dv4HceCD
JYpEXs3LxHS4A0e3O4qFtKpXq506JCduRYdZKUZqYpK3RUZbijlFZieAs2cvBEtj
eglOnWD8KjPUv2zDw3KJH9aPiMgC8XMNQBW+e1itPTZofUxNXbmUK3uob1E2roCb
H/WM2lupEj/+SjQhqb+syzZ0SG0hkDSu0rZfMAeuJwcdYl0uIl15zd9eW2NzTB6n
vsnTiqG5cdlsZnbpQW17QyYMsa/ddNunGmjq3U+I6n83R0jyC/bpH9sms2MFdo1E
UqsVmioxUU+Zah8i1nhNQt8jlCERWqj0K93KSEaaaCJ0DGd07P1BOz8bg2BlCnlS
CAY1i0l4wC8iN1lIOpDWbTR/D9HPSmH5gqhKB3lfQF5RD2vl4m5XluOVocvQbihY
c4yw5JNa2D0fiyS4n7BDFiTLcs4kYAmeEEJAmu+IWUq1Td/Y4OZatNxmPztignwa
EHXW6ip6bGzjYLEHTibSyeKhLS50vSQslJ8nM+JnMcbxl5tQX4iDv/0UptDVLVZo
USZLVQ8FZEodCLM439uZApi+8vViUJ7FDzIQ29n/2h+9m0fFxSkCfG6MXvxOEHT9
8waSsXqpYKN5gPIgUohYdZvssnrTJrawX3qgb4YS4Evkiba/SmZ8Jw75aGLuxQVm
QrtnCfoSClE/o/V799MmQBQQNsWTvONLwP0DmiVpbLfUvA0ApsYdpdtv0PNxIxD2
eegRu7Keb9ETJdyEmJ0x8Z3ZuYe+htOIKV1lO0f7teCX5bsqKxetM05uCKUzFcOb
hCI2V3rP5N8GOaCxQBPCg1RMoLwGlvIIKH6wNQ/T7oxzB2EoMK0s9oSK0w8fFV5/
UMb81LwLCB/aPtRUEb6w1Lza+CgT0MkCg+FS/lnUEyhLdIAzBB92SM5vgueCSma5
DnacwNen0D/sw9quAcR6vYp6SpJlWMaD+loWut8ZlKqVJQyQKc3EaE//0aSXpmvi
HQcWUTYYJo9jsb9KN+06RYz3u8DSY6TgObQdhXv/hqmY1qvfoLhdDAmOfkWKzD82
t4FBoCbe/bCjdj+JkXr3Ta2mkA2unhBeNyNADmO5rOhCRqHfbBZMyOeKOALIK3Rx
tMOSdek0bcgmxZZVuDQ1L49Z4i+qvM9dmkD2C1L7BvlRVdCwYPc5Rm0aGlgJKE3Q
DpHl6cVMfKcUG3VGIwcAdPHCQiOgdrQX+NMOfxU1oKCAh6CXHTOEAmG7HZrKm3nU
wynSQsOyCkeBHiRAs7FhDb4Am7I9Qvm5u/kBbXZDDU2UpyrvPKAb6ZfDxSEy0oGK
u/gQ3dRtcrUBoVgvg+H/rjKRZ2r1dNqIC6qhXODng5QjQm+mG+t/uVD6b1el9MaX
dsTxo0trmMHZzK4/DS6G/uysXQMY0WgDvPMYxW1wMp6vwWS9IL5Kp9Rjqjx1XmbB
JrEG6elaJfueep99oBQR7vyOKOeRGje7MwZT7ZCqg2xk+lcMZFNPezRFiS1biPXa
nCTh6SSukxd3DK+xr4lLH1TuDsQtpnPJcosXh8LIgPvASiaZ1LWMMdox7FWQ7AUw
kgqWUrbKsLQDk19ndPu3fOgu4Xj+CTDRz1EvH846Xpidz5FhlQ1VPIxlh8r5vXdf
687n05J6vk0MBztG986WBpypVsI/nzt66XAqocqbPbHm8l2DRlfbb4F4s+oj9dFz
tTBAtTQ9z5KfVM/Rja8hbb1chZqbYxV97yqaCEDtOSFnb24RWVcmQDfi0PahYtqw
yvFF5WY5bGjZvC7cRpHtnwBFR2wl5pHLM1ES2NyBF4BoAyvU548eC0HQJ5rj4eH1
htCLwR7jBF3rBbrX7rac6AJdo31Oq55FhEqgnAAoNyzOxV/Zi9Kvnsl9s81job7f
vsDN7B9Q/LBSv4f8qwPWWOqi6BXLmN4HUO4ZRR4Y0Ofo6vEaUosNM7344fgAajIp
uf/OyaatXDgopwNlJtSoGzFVJ1X49+xaUksXs77Q7cOB3zVsHd2OCZ2UdduXyFyo
0nj/YjnJPsTHY68bUtdBMytL62NufxaiWleOacqNr3qb+t+tmuduEnLdIV1ECY8W
+mzDPcpbUY8IdFd+PHeCtobrugXOY/q6cy6B+GxCyWPzHi3qPS0Xcct0h6TTKmEz
6cBOXsUa9KH9/Vv7FZpMgB/3EdUsxiKBbsQc8DfY7BSXigQeDRR3YWdKRkbzl1y7
hpb8+q6Wgo2i75XuumQJpS9PLk/6c52iS0drR3Lb8v0rz01O6KE0Ygwu9zdRBaNx
XzhlKm09T4CQXAtl7TbBLSrmIfGw3Rbd6veWGyi/tEKfuI49wVPIrsYC6ZqTQMUl
AMnumUQEWJzrKYbjsJooyi4sz3hsJOfIuXWiTqLNTc7eeCFu+hNd9qWTAr3FCkpK
s2LdZZRhL0pxR+RX3v5noMN2V9npzdPG1S+YJZ/s/fesO4GkN93UNqcdOdLHT9+7
XbPGV9WxFYIxHiS6q7xlCv276lrFFezzg+1xEbKaS4ktJT/rVRSqpEHy3VTkIvA7
BEGbQlaOhOigZSLY+UkJ4LIgMtQzrGfxHo4LUhyYrxt99ZzJ20V8J1/+3dPuzvmX
nbgQJuTQfHCUkjEoWaijAi2lMZtVpODPTnBabSwwrKUSf3c5JdcyOHvlwoFWT9HT
bJPMFeJETIpwuQ/MaaO69XPGhyADQT/Q66XcBZy5bX2ctF1nM+p9zqt5BMT0Cwm0
rrp17Y8C10w5DQWAgvSPa0EgxWg+3rHLwahu5gm7Rn+q9e8v4JGBXW5rj6a7g8Qs
02Bozulv+H4hDXGbGA+9z3+bxTyZ2l1oIj20WWlU0F5RgNlxxSy5XgHB31gAb6wK
BoT1F37NLQmIDPFbRGzGuQmUqdCxYFWCQttGUj2DxNrhgE2TMUmjJPNFMPRupjzx
kPS12W1WC08RHnGMFFUv51fgbMqloIOlwAa5WgrSXE2Dtyhv0sMV7knYDoihaf9n
hMY1gW3F1svefrsbEXdR3JVDavG6rH5wNAVe6W8FGBgzw0T5fB5Z8Z+jEQGwY6fu
18JCb7YmnqLJU5OSPOXjCFc17FF6Ts+MUdDBww3SkV0AYHXJ9l70M85Cg3TumaAI
d6NOkQJdXvYc28N8jbpepcDLbi0ORU1LPIW95PF2n54Qo05GNvzTR2EGRwl4JYzH
rzP5g7yN+zmPkx0cFQcx/3b9/aTDUchx6pCL4xE9MnrzoWNMQT9gb+JwZpKv7Pp/
plMlGHMbzZWxNmjc4nhYj60wfI0j/xHkxizVEruro244MUR53qWaJRjpBPTKc6Dv
IdkzrY+133dqzuzN45DxtGppMKiL5G3xMjmqVDK9zjLS9xjbBApPSeZQ81l4F4zQ
H+xMCK5yxx6J2gs6OGo0g3je0lNFKAcsC51JdPGqCcP+U6LDWkA3m55C7hfcNPa1
0OhVDFLT01kCegfBX0YmB2rpa7hZgg+aKnhQsUdMTV99nRcD9WS0T08yeaNdffHz
OWUa0FtKWmTTiUV9augM/Rvgd0ReudT2ZEnuCQXq9b4hV1coS9znzxTfM2SQw4de
kkDNok2FpLyV8SgQkSMDksAYMU+p/oUzABtbg83mCjj5mBc84tpkr74s5S7XOw8Y
VcEoSb8TVYUeATqSvu8cul2jUQQ/Js/s536ulEz2HHyXGvRuECBPel1VtPwHO3K5
nCM0A2gz23W2R+M9QMDjlWcZDEwK0458aU2/xPJ27yhyqOn1PQefXwQqVMBlL6Wu
n3Vo4kAkICzTHGy9rLGkMXh96ZC223aJgNC46KVw8OOER6Ty0oZUCED6CqArEGXh
1+gOUe6fFQJbGb7cWHY+zC8+4cttVR7vnbeFwwvrPKSn+6eVqwwHaylNGhd1POPW
FjdoMHlDb9bVaTTb5zjOX2ff8q8iC7e7gkmw511Rm//TR3nINoL3YOOOGVFeLLFv
dBHRk3vsrqrkHglnoqE/Ne6dECswIkKcHWEY5X5O3zvtJS0NcugMtaHI8Yn9dyCd
FTYYvVMDBGz7vYsSOxUXyzkGQHnNJVmriZoexzRDjF/l/eOD+L7o9xgh+7oTT3Q+
eIWUguyftd3UojEy9hskOnBjZf30SnTrO48GczDmBsWBTo+mv5ar8UgRrR7sK66u
vg2OaigCezp1c0YgBDp5a8726WNixCb7uanCArxqIl7U/jwya59X1MCw2VFX3lYP
RkjJ5cDcLDM1PgCRDTiu7a8B7RHyZOo89Yu5Woz/eB/TptmX+DGCL8qW0a1I3VnX
9Qbq7gRM1H4HywqfXzInN9f5IDUv+4+Ei7G1ZpqbL8zvyTQ1hTN/X7H1rIEBKsOz
WUas/4mhg+3NNYrSqrH/dfbJYj5ukAOmZjn4GWHPz7v1qpYJYnZQ/nGN3hiWGNV3
pfElHEQPSNAP2U/JcJ/Byyy1balQdu87XWvf0Cesaw4R+rkXkNZ1bglMRd+CjM3C
QUmra6FRlTHu70jCVpeIxoPJpPeMKhs+naiDkqXgKNrYtS2Sqc4UHkbU+CyP7aMx
Qi1Ykp9+5MJYmvx/pfEccqmD1QEejRX0FQllz98stptnP1sSJEuNQkQV3BlUFyIO
yKgL/Ou1ITFDMnQOugMdOllfnWmd85bVd1RemwN/btHg5jd9Dsvpk0MHH/mRkWJ1
FdnZNteEhKFbOM7clphxNrf1+BVADxUTvC623SJcq9PSK/Mgl6A+TIrK/+EGM3WQ
uzeDjIPdBOWUH0sbLlNUQL5ldJV04T3FuhazbBEkRekDBPLd/pzbvIutLTYIa67b
yh6LuV52+IwG31JBngAD5XRzeggXz1UO95zCFTyJiFTPrcMUf6WpFQ+NQfy2DzyL
Yi9gRYjxiAmbrjrSuHEVkrSOYDAJsbBrW9Vb+6A7a2TP16qq7d7KSlp57iOXdIlJ
ScuuGehn3/Dsz1peFFq2iwAFm7et61t3hcQq0rjJRjz/3wYKwm52Tfw+d90OeMwh
VEZ9AZAqbPfVu8Bx0ft+tkkOGWhvrLNWtwk0G91DWFuE32ycEC1UBGI2ry4u+eX7
ed3yW582ye8s5ySqdAp60yxmpqMMAH+VUFD0c/7SByDe9tOm2XUqOUHCYd3zyOWz
UUPXjwDwnZtvudOTilBkQBSQILCuXX7yRBT12LasC0SmAam1kXFultn5z4CeV2li
Y/Ose9BYF55eA5bwpEB03n4UJCeOWqMmdJ2Au8VOy6P6JmorEsyw6v9Ty5xtI2FO
ZtSQM3xmhMV/BsdA5ao3eBS2sKRq83B+LCjt0Avp2Ak4YqRHDD8EvMJiCWrO6u37
nQAe4nF9/iFhd8hkY/UmLK965pJHT6ztnpXgS9Xu0uAfvf/P4vpSVTNLVgNBah8I
T78sDSqQcUsInvQ+5NMkLtD06Gw1CL6ygNE9mICsppyjd0wnV4gK/rbI3ve6aET1
j49Fpy64Y4ujjCQQ+y98UtjTcoviahXivHm3+FHHyRgl37cPTzNAxbRWqaJpE65+
531Bg5qdzOUbi3b5DSCnj2j2CZFKZsyxZ0NzqmIMHYi1D7DJTwudGsMdRQcB9TTI
vE1WTE3BwqZpBoWWpbHMHHx5QFx3JIjqmTvxm5L2x6atrY5VScB27l7TFIAE1T4G
lxlCoQLB0GXexn83Y0Vc/9brXv4lWxq1K6aBs+BbITJFx9RyIQIuCJX/epG2HZgS
g/E2lWSJYcwcrH6JarPmlcdwm5envL8t0jqh6XalV9zX5ZsS17EKeHbXUOd5TB/0
05pBtL8UdiISsFDTyQwMEJ+JnxdfNkDgO6Arx1MEEPYh/2B3FkGgII+DvlpX8/4h
/JhDRzZBbfbxg6s+n+cW7Bg56BwFcteZkDfsV3cu3KJBqr2fTVjYrxyHXlfB5CZX
zjAXzz6tVtTbmb93XvBUKfP9SxX4l6aypcSLHl9HTOPZXYzzTRbwZ+sK6TIwDsW1
DoiB/nX3anOoHaR+zC17SQFeUl0z6uNEeT+lGURMJpGQ9W8iUGG4UMQGJayiE6tz
lkVdzL8A9NOttEPyk1cv6lqOktQXA9Y9+dvKlcIlkvm7M+pGSYEdz8frkkaCWNV/
SsObbdZDM6Oqw2CYQsHuVwdgH5oYwmL/PqqxMtZ/Ir+DPGA2T3hmHuxhctcx4Uom
s7wWaI5nh8dVDaq9yJ1gEweK0c4dqYhJRUVgqMN/kjHwxUrKM98FtjmEIDsw6nGX
W4LxqWnZRgYX7KWuUk6PRyILRJtVfxiCBm3T/CQge7C4uS8o2J4705Qf+DR2i4Ui
Q5thFLsyaf6/55iz39vRqEafeE+GMNZMjkdhDXMuoYc83Rp9+DRO9nHOODfpZZZW
1Nh+UNGIcrt4+AJL5E77TbMHeDv6P6iK/WAdfO+IbxZOR1rwXGS0tvVMuFmnE54r
TcctNpQJwUNTi7f4Agygf4HrprrzU+voWIawdMv4gEgotNNtpPDWOg2wzPLDS+l1
DdzN7rhQ8Z1GPKERQNm89I9wd7RGDG2hm3C1X9SP26vl5oR5oFbu9M4X5aZqMxr6
FScIko5VpW6vDhFilqduyB/uj/68fdeHP3JBoTWHHLdAe+mAbXx3SqkkJmPSlRIo
JQYQLW0Zq1tI2b30ZQQnl2VyWikM25c/bFnBOmXChOBj5vtV6yR6Q+45JQ8chw1v
+e9KBjnrLZL8p3Zs1F1SoUXjzLk/fkE3WYuz29N7XXxAtAtATd8G5q8I/QMV0lI3
ghbUnJkgaKRoNgLF6X3lGCyESBdXwT6x9N15XbOSXs0IyOjMY0bNc6xvpfjvTIAB
n8XwMaoOWGNWy2c305x2j6D9hZ9u+NTCyfuPO585/rYivRYj0s29bPIVUIH+IXbw
oBxYZEgcJZV22loCLh5zwoce3+bSbxYj4mOVIW2vfSmVleqUjgWsQ14oll0Q/ioq
GTniwscCpGF3Zuw43xmxStwG7/zMUFJr+Qpztz2Gl2+Aziono2nm0uMo/rF8aB9O
lKNgpQqrQUHgdbXB359PNnxTbo2wOHlcdDAdt1thIXjI948CtHabJaUFLHL+CcMk
Zy6oRNAK5176LykYMddtqKfctk9U3QVY7RsWaxQpr7DHV+bZoavlbPFG0pZ7wiNw
YaNB1NG9JKwIQWoy+9PyxK72yIphddlVZ5wA7mgKUeCaqFTTjPkkmlKGm+iT+c+K
oy/7Qti8tosxP+GpHE15Wy+aZD82R37LtGBqPjfVUSW/LNxGYt/otPprJAJUvHIa
nMUjs3A6mdaiSUyRVaL/O+tCuHDwkzr3+c5j8ZMn1zQOrSEnWfuDJeav+AnAm80m
8+Jw6fSYi3NzaDvuknkgcxBAbDY2JwNvXiYBIki2wm/Mf1ToTdU+HZC7gdNojkLe
cu3KtYo34Z9sJw24TnLh+X3WLNtV0RjEwt1/Yvov8HZuKBjiksHojYpLKcUJe6MG
piC5ayb4bjDLWgt0lv/pe8F+UOV5ZpaS28okaGXZ5wSMeTODuanG8hYuc9wZtJW/
RHrhRDUpVeQQDvA4FkUf05Izhp5G3biKvZnAXBsg8mbB1JAb3T9u2+Nqdlernfga
lDySW9OdBVZIQagUhaSK9VvH3qiP28mG4w3O2zWnTUHOHlZGJYQWPpvWCnNPh+5u
O2LWDv5agxWSQ59KmUrPPpREccjJcIoSmFn36eoO8zDZHs0jIu65BxG/7P5mM1BJ
HRnR7uzybGhiY2inx7s+wBfvWvBvAo+kpX20hqv49+ictgvc5+dktm9qALr4sfFV
C/qHbTubsWaTc0cBDvwPeSjKsDbaeahy83lQYAX54tlJrFJckfQmJYO1Cjtak2Zb
6d84B/DCHbHppj64mgRj8FCTF2rSyFnpCyf6+Z6gcB4gInLOybAQCvJS2HXtzD7b
IT+MNKBPxHUEWekoJ9+1CwADrcHt1w1gVJJjPzMt5hS4790HPh9V4cVJHG2R0cEk
slUr9TwyT3X7S/gwWIYRLw+MICk6nPsOIkaZ4OU+1Bb5PXYk0yBE4tI82QOn2mbD
maXgYcoYgcwGVtGglbPRit+/FuHuRknN1fx04oXauoKX7scqiYLB4el7RBYOn7BH
sZXsovSIeI498IRer+yWRVVL4a6T6waBJKHzLrjnFdhgUGJOA70+nynyLRc5fsDx
hL0CTi5xSeQf/M9UFha6H/bU4vThShJHjx0G7KCzmw0+KhB/vNfmYR4+MlsN9Y8g
DdunLiRyfXp9QxIk0EKRPEX7uE3SP3ec7Urzs6DEPi/pjdzgG7jAOUKoQjb3mKLr
lehl2E4CrL0QFG1eVh/YcyAEPZ1QsgXDHlaMiPUAzGYxRVrI0E7fLsQjnzYvSjDo
voLF/SleAwT1oJw3sJJHQA4bqDfF/FL25xACmRrlR6eW/5NbnGnbdg1+heUyki3h
dSPMs2+CT7HcQqck/aGYUme1hCwntpCITMZxY+7+YuQ4cdsGxABiZp0ffpReEoQv
V7IaYhukMNb3Svr+7xbLP9YUffT/fOMICqcT0649ohK5fcUXEtwkgjVYHrSZ2fpg
SQ8V8t9ROb2U05nXeYxGUDE7dS7xEQcUgTbi45Y4Pm2uKLf0puSB6ZL8jNPgW8TA
U4oPFY/BgYH/HkFzIfK+X0q3JSqcpVREWpEhu3P5RF3H14jZ6pLJqteTl/2VcDF2
fqWAzz1yKxz0ETRF1YA3sUWaAuitS65TGyAEVDOxgCXlw7EWWcd4ZpkfWq7lumFu
3huUinCN14ihuQXtgKre7x6m2+QNiC6bSXiU2QEN/6x9h2U4s9mzHXFH72vInA5r
UvOcshAj+flFWUVDBYVWyJ909GL82/o3iA63vGiF6vxYUYNvwlqJMqW4nHNtXfSl
5xtfz1MfYKztM4XgRz3EWsr2BirA+3fJId6YtUv1D1l3ZtramRWAHX/bh8jtouM/
b0Yk7oT9dCH7sbNUE4lC1IEH8DQ2ArhWUqsjHoLtA8jGKNedhHgn55Sql3N+fV4T
eMPi5VOEEZ5lgyfBoJpgDeelmr9uiIeVI/9wlahCmRPi7Sm+ezMdqyHXVas1a8KQ
vjnAmUQoBOK7P223WSdEbQ74AylUXrUVvDKHIo5nMVxWrquPo2GqpEAXbr0VaCNI
SGUY8bGxp9tft0i3AJp6Y5QcQxZM4eWJO6mdsqZN2Bnw3WrlDb1Xrfxee862EQuu
qCIaR4k+5f6Do6xlJ6Y3y+QuFEzUuRDrBLAfdeVVVXTABcooukTeDkdgvf02WBSP
w5jdus91JlGn0wD6+jwkQ/9xonnIftFe57PmQKB0FIAJO0XUejYU6lTUln7doAkw
EfgL8ovxqKgJG44WyGNHJjdfgXwXNfffP8bikZIwh9EIusF9GRnlvuA91YUB02dG
Jj7d+mOgwwrAAr+vEXq5W3+We5MXt5LaXiHjGf3j/OLXAKB9S1DMmLPLcFNoIatr
NLOkrm+KLBMsN2TSgtF8BvJQGWiCDDJZCjlcxT0K+hzLPsEcFmQsg/QFQAO13QJ8
dK3oGtElM0qu8zOD1At3CBgBVLVASfWqv3Hp29D4R76GSChkV1dgegDC4xRH116n
/VOW8WnF/Sy3kDaK/ZiHpMYgG7/3ML6ZUr70cnU3TGrDlyLsevkLppmPLoD6kF9R
Azav94P5gz1V06+9gQJx07IabZLLKjvi2lRbURFEnskZZ5lFABhtLIt3NZ3LF193
zy9Iay/cmhge5BZVm2aPc9Ei7A3dgH82YA760SlxysVYFZfvKBfu4NVW706M3mw1
rCMvZbnRX4NNwf2srPlV8v+sGTOHZ/+b4TmouQ6Jnl+9JAFbFAIHzDnCiIW+pVFD
GVpErn6kqLZBW3Nf9v4ciWX45l1HOcnEVM/hbF6i1fIArzWDna81BezPFjrFeECY
vFPZlsp11bmJHrrnDObwHvqlNA07CR017n72V0Peq4tKDIxqjPeVDRZTtAwAE4mM
C1SGGNSCydk6PKS/WOBarXoEchvkX3jjTcac5W5YW27ZTydqTk/7l3XK4RRYDRuA
fvG8LlChKzcnfaCFBTKl5pnd+hxG9lMrqHOpUu5RwGsB7YRLLhePI7fJURBlZVYj
3TeOsDF+Pgv9j/m9B1DIpFH+8TXfDHXu6Rluagc7PIl40HdS9JoQ5svgC51TR/+3
+0Fp51A7c282NaIskEmdIFISGU/m/x8oLP0u1BJg7FhhVbRVhbxSdnIrKpN9nZiR
e9wawsBWMuupoJSQQ0mbk/h8xYsYJ6x9EIjgdDkgbkoimISvCDaaI+Y0ypkIzSXM
WqJyAJdCnkZ0+LfqZla5SjDsmKpNt/KhW06DEuqcqXAmuWv0BOMDcHFl2Kg2BgoY
Sd0uKmyBQAhZUm3eTNmS9TtLi+TwHvHYN3s213iRZ0H6ZTWpI14YhEMOTDA2iBCk
+OwVC+dMuZvjsGiR7szO/I+8evD7Ap+8udcZwMQK2EIZolSjWDA8lJz6AViHek0i
4FsTwhdtCI7PsHFCKsSk1VYZ9QQdDe/bLV0tYgGRy4EbOUSKs7aIAbi07s78hcO1
Dzl89V+7qJIajaH/9q0PDsgos8HGf6ol5S6e9KOlXIF30l/6bAzRyS9QzfmgVo2V
YNQb0QMWmvxvAJTgM3G+Dcgiwqkrk797sQqXaDh72p2Aoa3UAMJYo+ZmahG2zgJd
Fb5wbIqPQhx2RtgV6GbHBLcyE+CuDkgMvYsCZxdrj4ukE6uOrwkI0Egajlm/sdlI
l7s4dbCM6+jGBkrvmLixdUmlfWenDHuQut2F0fUZrAuN6dgJ+BNsnv6pLGt3W5Lj
HuGj/2MVfl5quVPRyKXHpKhxhFv2v1OVE3OpBeknKR2KBM7OCEFkwqphWu396/Wx
48iO7oJLSTVupNGDkw0YtGNC3uuWOa9ffcMJiLYSugEd+IT/9mRYT4zfawFSo4hI
T+0mC3KnLK8b1LxmgcAMxEm+fykdrD4w3FFe6JHTyGnth5H0T6KxYzNyLIm+QNpa
Ji5BqludooFHuX+ZCbX5pGv9ARY6W/nvjTRyHq4UL/t0U7Wsn4jqdBNUKiCZdofa
mQret7yFaBOqCa5PqpjTdGdDV1ZNifQ7TSa6Gyee2VP1lCaRhN5vcYGhxdXbLb69
djhJAXm64JosqCQ6k6IeYrNIfAXhtRCb9fKJRcPL6dKKbaMcFUba6xVm1Yn5Ndf1
nj0NeZ76gso1PKhEDjC5DstXd6h+8grNbcpEWKNZxbA90/BGAr8OZjLvRerOvzWu
poq3/JerbXDq1P9en6IhMxUpv041+nc3PbZC2n11tWH1CN85vmFP/6n1ebd3vgMZ
vAx8Ft0y2HsArbcBufyCY9byv8Dez39UTKmoNq7tjsNOrb6+2gdIZUYLgm/OEa+t
eqjoOIP+B2ElYgrJ0de1FOHMWuFuCwlfoTZsqj36SOxbPPXpfg0N3R6VcGcAxCyO
PSnI2OsA8pCatNFH0gQhNYril6rtDc2NUe+OIinie25Ov33kz2wNAqf874nVp83K
zrZF2E3eWWgktnxQwAT5B6SL9nWIeXdfjbsuoR39IW6BatbE4oZSTag5e1zU77ud
XUqTXi2+5KKvzMx5tZUmGPgVXXmNkCaXnDc8JzUS7VEeh5nbzX8yKnwcvX4fcO6l
gCJ1wINkp4HByULpOb8k+eRE8Ojw8U0vXanpUZ823/jqyfe7leQeSTT3iErgJYIW
8Wniy7mPKSfKzRZqEOJc7Dr6ILImgN46PFU4b1uPr4PkwjxCuREWFVtW+HyhfAeD
0zEQkoF6sZmdJP0lrKxEAzrhpzO3N/LwNxenaxf9syWP5y1YUToC3DooLfDcdmvZ
dlHhRV0O2cwjfxUYB1BPUnKIwVRtVlXZW6HLDio8/32ai0l/ohzto8uqBvLEBSkc
idtrNoPXrL3lnZwOp47wEr5QuzvS2rkMiXBVzrkz3AiC8PwIfes2aE8ctbuqcbSi
1VzEUnDIrv+hLxdCmp4vYVgxZSU8nLbWc34VBomgrEVN/CBAgwsKh76gWwNEK7IB
4y71fZ/CjH0HCVED1+WhXl5TUPcNhSivEjqa4g4YhctoF81eMK0lDwfNWRG8uoVO
VcDLC10ft2e2EO+8DLqYmrpKTDwMRciggWDb+GMrTuKZSLMzKPaSF6X3+Fvfkw2o
Uq8zwAaax3YoGhoBRCdBHAHlyjY5q8Cy3gj06YHRkC2CGtZhA8wecE6kQrwN8LWu
wu0b783W0jkP5oT5mMF1Wz8aDSYDlFgNU3ZsEMdDhNfgbgtwxYessHqLHCgLykSw
tziFgcgtASmF+MmiFDWui9vRZWVEBHs45h33L3ABdqrhvALhPog3PVm/PlKLI4uQ
+SbvniV5uV646yiIONajGwKBzuJ38x3+R9VWUB49m8bHfJbfVlcB1MXJ4TwMoXKQ
YHXligpWsZpbRaBxeUOQ4hLJkfCsJuAgxOZBFtz00r2PY8hkpL7U0j+1ePBgJAbz
s3hDDIUUYjeWu8gNeL88hNkBNXnLKAYdAI5FtbS4LpeBHcp6qPAHc98V4TafYJ+a
xKnSX9kmW0jv/VWpOoLi/nfeKLHQe0eLoGcg18wAtdvGjqgMh0koL20KvpbAUKjv
/aTYRTZh04l3SwFjTcfoa4mjbXXnwnlC5U4O4kIisBt5BEPdldKcRuGuh6Bn/Anx
I0CgKaTmnSKpL6UN7U7UsFoA9q87yz0hLGxuwxzTJEElTW4icxbqEEEGnKx+PaQq
BbSsSppsS0FtYFyBkfJIjV0DfuDqBjRSkUWjN/A2ThdJ89QF/M5RKhWVozpRb5lk
glfv5JOaRuMarUP5JVWMsVSCn1nuLLFjbGeIlTBeS1nY0WqSDcC9AwDONE8nsX9B
91EvmEeT3SnCKK6j9rVym+lnIMKiKrq328MzWSIC/Wa60phdyBGc89bar5L5VILY
NP0c1lG5+1eZ4Js4CTp3jNgKduh3+ftVskS9wFcTU6PBpZ4WM82S7lkd1Dv424g9
/IMpISJKNWR5/hezXXvJ4Eurp7DxdWLsjAPIPB8jG8WLsKPsdoSf3nP8+7rwScxy
oQX1KcC1hAAUaVMFDije+mJeHWCNNVSNGN3bWbtyJo4vRWDAAyS9SBzn2cqzj8gf
+yE3NAqTbqQ/TFqAwN/pIczD8ba80Z03NDDUfFEUZAChRusA+uW1bcvhpf5Xe4eP
1G4OZBISonuWpUIxkTCqLvl+jXOQLLNtSdZGI31MFIPeGoPGrwBbq0i2MP6UGtol
EG/Fh3gImR6qBBsRHqrkNDEFggYzZmdY0rXAGYyaz5tLweT91a77p/j+y6irzUCf
uJRXsHz+ciqAIKY82sf2C1BpxlAUZjEZyvfr7VkT4TQzwiBv0rqmRucEz7D/r/Ul
tcv4VGQLRBValmHowrGTZrJeSwg/+zoD1VSJNPBk45Hf0Qr/vn3ADmqmO1ln5uGj
P4wjYu/S4frsFMUt9tNxjevxCfwmwmy2LsUEW5utSBKNOX8+9S3GsnAmBrn/PYHk
VeETEHlHbvJNMRWG6dgcpWamQrD900IBnfZpARV/U07+0NFfOV21qpVpqVWJTqm+
Iis8cskFxCCL40uhIF7FtUbZowRhQfQZIUNTn6cFRcOnoyrOzWHIhVNkr7HdczlV
7USejpy5A8RfvG9t8lXrM/YlEz64SYJtJbDspPDSygeXDDJytxLHxTBK14zD0i8Z
dfduX/P4f6qUsUToxm4iSKV8T4MTv7t1NFdDmuDYuqnfWACJu7P4JBv+5QcXyFxg
0TUA7Kj41jkwHnYUmtl2B344Zc2Xi7CscHMJ4sYOXPEyqorFsGN3g0Eae6RkLgvh
LD7GhTbyykByCHaj8WmGSJl+fJAgJlPLj8E4B/aP9QuIqlIkNyNi9K873PwTnIlR
r/OuOs+lrguwuutbzrGTjRKH6mhwb4zLBeY6r3/j/csJ97C7LlkRd4bbl66AtRwB
oT+7PJ6H03xIIF5aCinDk7ZUGRQnp/HycqoBrS/gL62JfmgjcDXmANbc1e9ChRvY
P8q0TGq+H+M26VJfAzdyxkEEIwb9IZc0pdoZO+s6L4sbk+0MhscOVML8gKfHgg2F
OuBt016d4lAreKPr0mN9IlxACn0pjrGrVuPRzhl2D+souUy9CL8t7tkxQKJ2tquS
AiOkA0eE33WcLOmn+sE3Wpke7X1JbSRrAoW9Ov1W7J0nMHevXE5gDLc2cUvI0jOQ
4ieFLlmHGrpkDew25Rs88EdVsq7LKqqc7iuLH+5ncEcXaGxcglgszMydsXVDHv2+
FbHIaCGu3eASU4NOQ90virtekEiRejgmvKFQtdoJ8zzpltHy0G1LwIoH9kkpCsVh
cP2dab8E5kCmy4z/EWrKIyXXVVu95hOteoqbL6mOC0GUBzJVrlLfuCimyLcGDn2G
3Ravoz88xsVITYhoQIIRyxJfETNVH4Z+ppDn8xSxW95vLpa/il30TPYn2iG/RxBW
2GvyZ1TtpLlsX1WyNq4MV5h4IpI9Ja+VzosEiWqkww+b1kB1ZR7jYKXD+XZ+PqJ4
d1LZhzGOZa64A2RvcJa4pvsJCKa8CzbWzygoQEMhNIk9HVY51C7GPuIuFit4ZOHU
R7Yu4yDfnSl/udfqtit0TxCX7+Iltvt+/s6ZtsHf0s+w3CfE54DA0fpnTM0w9cEz
phqdrFYXhKxD+311KLnCB8kxgtjEbbHepFkXa2yfkBDUDFL0+5sKwhddrsqdLV13
2kUq0t2XxSEvGfK1GIVFrkkKwyw90UgjbE+xz8NmyIz8H4lHoIjEpUY84njytp78
ykCz/+jYcYlO9nXN1h90Nph32Kfgn5qBidAc37c86z/PP6cXUQM+kKuYuPd7pUvk
HRnw9NZOPmtffOH4QqVHl4idamirrTZzN22I7K2BnuXuYCHU53HGjhEf8QSER65c
/x3v/OciWr+QU0i4Ur2ewBmjL0rsn/GZojOjHB7UgH4b+mzpc4Bry7lBEDtaadup
fm+MOHGa70qT7XZQzjT/O2LdbBIodPfX5CLpW6zo0kGxhfGakP0l3WpFcGdrQaLb
atGLt73w4waewGO2db1HDPeB7YihLZVwtb6VZYOLHsqjcm3hAXvV16T9kAuNVc4S
dGkd1kwYWx3rY+fIMkmwKfEkQvg37eceLFkjWfzo0GHC1NTdb2Vh4SAeNtDmD4AQ
Y+GPBhR/+Ce6I0u3oykm4ApZf0jCOghIIX1E8bQQxo+zXf8jMks4VglTH6o2FH4D
tnKRFs7rwJbmH0hHi6IlzGg1+rMFKXaDLmreMUmZHmb6DNqvNmHW600Tfq4VJn4Z
QH/Tg3GWcD8zWHmUkEjkYW0oZBXRRagx1byZRkpPKm7REBSkeoNYHW9qn7wAPTV5
ZmYr8Gyt2TZGL/GEZpOscRzJ1uFr7lhBN0kn+sxRVkyt1h7pingMju9jjEh0HYH7
kVo/Csqy+fi1ZvNLWYD0UkC5w8qbccU67O71ueS2jGT624mIeTOynFDRBvfeMLT7
GWSZNM1o8bfpuIsMc8zFFmzZPRl3e35IODQfV5kZUMwh3FOE7SFGoanMaNLjsrQQ
TZkDA5KVdf4BGSmB1srJuwK4mxwzk0W7xaPazrF/rnBDGMncUKFiM0KgBrk173pj
vqDOeZkH1SnT7YN/ObXsC10vpNF5UccIUIg3Cnn0ObdLqg+tTC94G0t5HEoa2WR2
msk/Zn50gfzH9b6WrpkD6ora6sw0daFlQBM8Pd6iylnxLzTrC2IC2rW62Q2eGF4n
LtB5L6iHF3oMiwGdBBMgLYbJAgm6DRnBmTFl06qsqKVn6ECA5mz/VZ85bPeMUTrY
h2LepSeUjKW6Gs8Hbs+eT7yFdQd0GJWrJvXKAr3jXQFlfVJtLBH4JMLtieKtFNRx
9xIiQnqSsqsbd+yM7tpU/ZXmrcjbJFd2W2QYlPyS6FhLp5DUBrseDqj+r4eRan/W
lo0cNRfrWWUVQhXe440WOFPBVClynjh+emYCEQi7/dPE2hngxL99kRLsi1ld3Cf/
KIQ1gbaDTb8We9AbGJkJKuwAglBiVlQFLwAX5uQTHvX+BxLprkDNeIBlJHOEtQGf
wrFS8bQYhsaCP6SGgBTKCVvJ9sWM3Aj/8WneMVejfNQwnzKNBMdgWDZpYBKub6jX
1pIcuEHjxZ6Ul6oW1cfVrsgilpbpy24TVyhg+nyCJJUO7Jd032ab9qIjsUcOiIAT
RGzghPcQcoPHWSkRecMC1wk2uY2wXRK/0MwdH3NghHNURovbNAyRv3ldFTfWcr+x
IhMpp7zTw/QVxaKcmAf8mK45DrdmgOS9EMPeBJvQaLo/bGctkXt8F12S/UsSdcsi
tO44LNtAk4R9meWgXD2NkIuOOKSqqXRyyrB4fj7BNRiOxZwqotwso04w9RlpbJqA
eWD1/8UdihPAvq/ctqthP7Fp14XIgVKgE5+8rbX9CqON7ZhqyIr3V0l1fw75qjqq
VkdSYCCPMp2sZ8M7B6RZu5Nj01PcUxiysjIPhHciMOMds+EbW19DBnhr6cBjH05d
HRhLpuNmfhILI+hli8+nR8XLm9ofTnhtXjFxPyNHq0vpeMzk0mqn0ZC8lHavr+dp
vC1eamiq0m3TQwyYhzZpCEC1DyrgZLahHOoPmpfc9uykIyABCbxo/3O8pDFXitVn
7tJgcvKzEdXz6OL2lewkuGC+vGUl4thEdTVldfP7rZcyDG3r7PN6kgwsQyn/+UxM
QopjKzdSfSWDFPCfOh3J3VPmh69BLjWECrhj00uRop+uTK8yi3MKmYq+GwTe/2AF
ifYeCqnR+cY+eFIMdy6frYoYW4iDttpUbleXtiBaiywi0LI4VMt2nhszDDeyC0DL
/PYdy+g282FtqsEY4kVC0xBw0mgQi7i5/CnLs3Pi/pIa+hY1z9cNHhlhUqWIW2V1
HCTfFgXDrc8hi4MdhmVausvJo7Dkuh0svfqmb0ZTvTfcJPPNb8OKVNbPuGO53tdV
pyNXhnr0A1H3JJ8FhhAohJePLaQSXr/LAnEeOYSmG/nAleK9lKjY/PFKkLdYmYlH
2UhbFlEn7SXqT8ml0G21tS7bE4xZAeCrPDN8nlebhKbtSJDSG2fhTHXE7VjsoilH
8Hh+7wWsX0dyIDdD25w3UsDZRcg/GzyMxY2t9NYJrm1QLUVoYbK6/cKqx5iIZ2GC
esCVFTiBNU/Fj11SeIFwmr+pLRHkeBmti1EgbXE+eCybvy5KSAtsnLTHOdIobtGs
/nDUGJc/+yYaaMQoEpoMRrlG/cTm4STExsKo+ArZBwvf4dKLR0wfwQoxk6ynTRRm
LdNdBmdvm7xqn5yBB6w0DYckfYYOaRRMTgOzkTI+H0a7PpzqP1iNB0xdXCl16NW0
yXO2LNf+gIEECMghYhOuve5eUIS94JY6QkRY+xmyn3p0nOKychfu9yA6oPcNECMY
PqdJ65MuPN97PgHG9L6creMPSXksLXBdMEUXhIkMXUue/U4RAa8DhxESVZrTg8Kp
+gmX5yCD7GsHvkAy96g3r7PoIWOt2PFfdCzWQu2bOUdNKx0RDgLZUgudOw1H9BDk
tBQ04zmQlYBbjebCDaaFoeJJ3BYjDRXCszERlap+GnTyHvzMxz6O1oabNMz81jGv
p9vhwIYHnOJpyz2Vulbd9maXzroRQuNKW+d3z6I4xSowL798LS+EzQCkQjqTGB6p
j9aWqXFgVOnxcx+1Z2mLrMnPWwyfLf9LKRC5PRlJRPtpqoQUhtJDxYDSQXlWl3hP
63byahO1qXqgDH7bXuh6+ML1Cdd0GwsDxa1NjMb4MtCYekRxbc+C3cz7Q9sLiADM
tNIcBzKNuXau+NXMI7yPuI1ml2bu0YbZHlNLo9ENEuqyZJ83DkGxApeISF+oA3HO
vAeroIlqYyVaimDis+jWFzyNfiHzEVrukE3Eeewd7/Hlyg5oyoDecZZkue0/rkAb
81xuszuSG2xdFd2l96v/o0XCMmzLlM01kDOgNl0kCO0OkQxZ3IGH+XMxFk3JbVSi
vzESBMbeeX9kjqwlB2YK67zNIwMeaHIfYcZHhTJrEZ2RJznQFbtuX/VS26Jdfikz
wwJTgHYWan96hHdPPnPEIcjffiHQa/z7DdwKbQuotGnGFdOMgm0LKhziZeTN1Qtg
38y+aeummqUlLIviV84FkwFkZ4CTxfijghY7SfSAVlz8sWzavG4zRnPzq1DZ7tTS
NHDQs1Reo5RW5iBAqLvnAtgUMnQuZWuz1tDlnJuc1PEM7BBY2ppF3iBDzh9MKKX3
wRZfWwMklZaj5mosZSyBtkUTFyN5jywGtuFkbYbttdeV/HAqdP1E/5LJXcB+YZm7
meRBuV7xxrkmTF0Ujuhvg4ALt1qn6H+HPKAwvf85hgm6GOZZH7nVrgkLTBAPwH2b
/apDyqXI+QucfR1ftiJtnFO+0MmgVqLr4Gv97HMrNTUEoddYf+01mANdKHCN0YQV
ScJq03JcAPZ39/g7yzsSzbDtIKxRBMYcTknfM05zwR/K9XpFEnztVIVFgCE5mnmP
DMKewKN/7ZlFPXP7j8v+cpxnaJs0sM3fWqD6yJlfaI1ttqlslCRJpVWVq1zdlmOb
OHOhae8ZOUWbq4YSoRPj9jm4aCwV+wXAyKNSNqyD6u9SPNVDXhMaaXYN5OAY7jJh
QBVCcbjTKTin2RlOzP1LY1+nMMRKOmv1o1Kf/Q+peLb7lZPPtB0HfguL8sgxr54f
QUSjB4jbAfAi/Iozftimdhmc9sW3pMtDEXYPpb9mLX09/R5UdzBLQX8/HnC6zt/3
ShWL3+rURarwceKlb4QUiA6WTokwVi2krWQFZopkjXc3EiN9VbnwWjvm+iWOm2XV
YHnK9vmc76uX08b1idHPT9ZwB6XARl4McJL3/cEh6laPzDR2ar8qrtaUu3Rk9ce4
5869QlKcfJro/YHkW35i5Ep3ZrH7EsV4aHGpsRQ4d9JiLdvlcQGnJKcNtEWS4Ol9
fWA/GE3bu8iO0y2COWzE/oPZpxPaH/XgBwJcHcUr/HJGDBMdUiPJnpkcJ3B1W7le
OwGFZpUMmbhIB22Vut9GSq8P0d+ueNwt2jXj4P4v/+/hFi4G8xkRe0H+yJm/1oID
n5/+vU517yHTTedxSaYi61XwDfhuFSh8QozA+abzzHDkj4tkBjFIOxd3VfbP2PRA
IC1jJ7xJn1c3YpRiSvGxGTF+FYZPToq9Ukx58EbD2INNkcmF0ZJ7jfbgA7c4JVEg
I4vT9/9FMiSDdMZDteIi1Wpwl93uPpKktVob7N/eLHp8vBuI8d2/A9DkhvYXYUL4
S6BGvV1k5lKEO7N1ZAcXB1PDOKXRjnUYABaTn0bhKtzcvSBgBCtsPqru6nObS+S6
DXKE4a41Rdzy7JabBmSLT012WZ/P19p33oketYp0Y63Hiq+YEKlBtsY9wMwUuK5d
iPR8T4bN3H6RmZy0c2aIOX45NSXrM86zKdcrRQqQQd9x0RScA9TtXiBJE4swDNj6
Pob/37GWmQEeeseJIuLbA84fKAdf8VQEbYB5a8bHUkAUFTLNBB8piwbghOLuBS85
qqoBZk2tAOrjLHJ13MbNp0jlO7n+7HU09HkIZ6VJxYp57P5AS5cw0plrYC1RvC86
UpYEiQttfhY9P8IYzSTogYdkTNjEIzJXB7PzKh+iwsRlGwMq7nwN1QXY2Tl59jGY
63WTGDQJJXnPiNTZaPhCt0TVwJO76E+YNAPcIHzfnnNotPBHdMn4OZXBhye5diq8
li6Dl816JI2Ch4UEfilP5T6WwpA7vsEvFuHPkuhvwnBLuopbifFOsxbAKuJtUbYQ
spzYzCrK5wToLGrqY9Vq90YjASbN6ztFwLFDKAePle2SyVEl1d9KBWnKlTjUstxu
Mn7jv+SxY2IxcePH/ILch/iWOcwOW5twHorrqHvp5cj48YBBuBojl63lzQ2Y1slZ
qQV4ge/RwkZKwQTzmR9wLcFZITJiT5ippUtBDV3eAtDqMUOZA1aMAb587iT9JA7j
ckMVj1AMhzhgVREfatu60iggB//BWYZwZRDcSjHB6FCYuloyBJaGWfejf3TvqN8E
+S7ozz6OPRw8C+tRCyrIxTaBXkG9A20RcvZ94DDu7vPk2eq5xGFFmVEZCAL3s76f
uuhcdyxFr1k14HXGssr9k4MPcT8eq0WiKGwc+BaKsLsjhypyknexm8aRnTfpeqxt
A3PlxDwX+wjPqrV9p46FxdWrnusOvj/K628O+/E1BBdllt/uXh02eI16SaqVkaA7
Rv7HNY9L4KdK1yvcWxUjaK/a64crNuUmZ9TI54fIK5sUC4xV0iWzOJDMYKUS53cN
ZOEWodd9lSmyktnjAHOjWg049H0km4O2rKmrIMhZWDGpr6AGwhNekx3hTExUnKhy
L48SfYQYB+ZWVHNDz8Qz1tJYjc9ix9dl3a945NO2GqpoDiOacPnU9SyssAepJckK
P9g5wW17VV5qLOk8IWNJGHlJw5MvRtDArOvLuyp0Y/8sRYts81wAIk8sYR/FaN3j
GEsAkK9c67C1KiibGF/EaeR6rykl6bpafdQpZWiVAma/2cYLGQEuXP1hk0rBxZLO
ok6fCS0JY7A/YUVP3+knAyMWd6CHO0vOf6x9huaa5cC8mqKQYrh7/aWYRxdcFGVB
MUV4rru/TU2TCfv/Vq3FAOo5ujBxMrK/3eGl/yNZURgGLjjpqmPlJGi7+KDhEWQm
ytyH5Ms0K6qVEp7TP9oiLIX3+kGM4eFXVRxtls96uAXV0Yoadf84zqMW0v8FFrl3
s4U75VotrItOK3lR1V7AlN4SesIOAORNuw8oc8k+4ev+PjtvaqNd1xdarpC8hWXR
ThwBeraN7LFqghsHIdUpQF53X2hoRndyVHyOiaame4UdEwTK8MLjtnyw446SxuWU
mIz9p4xnJB8fWLXjAeXUbGvh0r6c0LgqyUWBjI+xLLWfE+ZWdRNQKU85TWfWz46a
MKFu0JxfMfDY6rBsWDSW/MZ/7hg7EH2dCvb6GW+ALYmV9ggsRVOqWSVSqUmjRqjk
0P2NyVzFon6XfyKLhxwAbtRRiJnXEw+5lO3Z7P+NQp+sGKWSjC7ZMerEXC6xdAaJ
65ApVcbVoV2Smg0f4IK/ZmeVYpzy69msV82ySJbXPftFi/Odrrdg1t6z/3HQ0JDt
h50usnjDY5vcGtf9xNCWzFLDf2n2nA9jkfOUo7pVog4AnYJmYCeSShB5jTuwZI1z
u1rbyVTQ6QumZcirfXyRenegGxXc7tYDTEVi9rVz1IXFoXfgUlpBwJzf2020nPvv
aMTb+lXgMt3XMXWMwCgRw/8meaWB136PnqFCJ2C7VLPjGvG8hwC2Jiqn1/bFH4zj
HlGvpmUQoKNB9+jchqpSPtINp6/xPDFvvo8LMXFrqM6VxJPZV1jG202DFSZaSgcF
kjOS3T8jGeqBIdTaNsfKO6FUDSgzyYGnLqzurFWakuFkqVvWo2+iAftsLDCfxZS1
+t/xAujTC53goIRfknBElgrSNFdphAe2IGy5HIXXLqApzN1TS9Zp3hUQcUjTESww
byuFk3gJ709GsuM5UU8sa45eFFyJXHBHnoZh2agnUhfKDrOdFr5/qF9M/uAavnKW
7+UAEMU8lgDMU5W1v487ZJS4qKUEywgAoT2VuWuJnmN+N99rIp5gnex0snoS+vFd
8hfAI+jlVBYjkRGfiYrdYPDm/CUT1ySzC4kwprE9TazswaoidfCn4sFm+JKlAzhy
/aoXL7uXXV6vqNNDiPY6tdViwx1hcfNI4kGf7OUGjeMe4OV6dcDUgKZAH4Kw8fS8
tesJGg0r1WcnrwtGNoVVveMbtQNg6TUpqyaCKYMEhiCk2rEAUX3hs3SCO6U0MGIB
yHpvJ13vS/Xm0DWQqPtoOJFml+MEEwgU2AVJ1tD1T21HtWM2Zv2aUsrvbotcrGox
LioHkNvFvX2bq+qfrIWMyp6iIyRY/KsoB4yHMtCuMAq3XkTBJ7EsIV+5IYgDtcmx
Kfr+EQ7Z46ZhUMZeyOsAYYSOXVkrlN1IWZWDQZq+Vho26b+/9XGO9hludQQL0w4Q
zpHdaRsdfQrLk1wJLnaRzH/TIc73YzEHvtsU+yARgFap6c0RvJVzyEsjFTAIzYzU
A+YRiM1WVIabBgr5oPsQqxuvCOWpAWRYpKGsk3o5kFcZEB7F0LiIuhOGV/LW7jIq
P7o8td6gFGkMRRE0ODs/Sfzyc9g6g3Lx199qsSXbGIjwWYz0Gu+5fjmNniW42J20
K5CpYEDHPvsFmp6nTE/UlX1hYrrURf4XPi/I1UCfjs9CNivnPpZJGZw0F2/n31Wg
JUebjIAjEpdKVaYlyFFNpnoIH12GkME3YRr+lJ+m3olGvoICkLUfRITIIB0a4MjR
P+ePGSoO6AtAWoyFirNeYP7fVXGxZXEsgtdQMlznm0jcUgCUXRjke7asEjYqn/WT
6lQIjlN1XL8q/TozHmkwItxF8dgx7OvsTrq0o5cb52CTKzQcEZ0hE0Vwr6LOKWa/
4Vyqsj6cbo1n/m0ZnHpOZeUgvO/xbaI296z+4xau00n9bmpI7w16wejHERF+XJO1
t/3q/D5xU2gIt22V8BErpKoEqFDbePnCm+Q9wyKzmCorygiQmTsOGqOT7X25Yq0h
81fCAX7lJsM+DjsACfigQkJOczHIyIei5bOMq3gjbkZfzD8vQwtgBy0F7Q8ZYGtT
UaKhKi6wj/V6mgupZ7lzhFRNSwL8SziUjkVzb9mZDxeXj9VWX82/xT7kTY+RlFcA
pfzJbqQzNIUqsqn7Q6lXLheJXhuxGL0zca2Qwlcx5rKbM3xOxd9uXq18x8DuRw3x
eSfZHIgIqQD+qWNrTs+VE4+xBQoyzAM/P/bklIGLiUynE96fuWq45DCG5faT1a7m
5+b4bcvDnYnCmXgIApiPYPEF07RG98bBCubrmjlf62oz4K0m10GlsF+BWe1Ih28g
2tr2dUamrrP0wIvGH6JljQNNRqqp8cyqP8TA1NYxM5JTGznDO/ZCAh3n89IXnQ5Z
PAJg6nlPCKOpZ6c7LZaUf01ee880NOPIIMBhYNgqFv/23EILTzbBVlv9myUXF2tc
dfQikwOujCy0nYEnFmFPD5wFP/SSw9QwKb6Y1Jd2RA5IIGzWyQwBRXJJgK+h7Wm4
Y3Oh5JZMe9ejLKRHkG+A+ZaEuH2nZxQ8PibMI60X5NnFJ1N0bBvEQovnkdWaC11P
Mha5HroW9Ewz/qPq2OSwlGtOcLg6gAkDq2tDR43mwnlssC3U13QVUKiTw80ARcjb
5+2gT3fzXFfmEeg0KZcxvfbm/OS0yaJAkCGbtJsObSDIHgj4ojq71crBAspWd7Ca
PDQmOywlbwdJx3Ng7CfnIUSWvBFo6j2rp2JamaIqoc5Eo98okviHyFXxW6jt//za
M86gaIGziF0H0rZEsr5SYHZTb8DcSaN7MIB9zzjEXHihmFinV1t9ClyWlCgSjnIh
/gz4iR9POD9na9eeZn+mP5Q4uvcOELkJpq+j2XWNb3Gx9YayW2zY1OjeGYI2gOeR
mgeD0pT7jdyt0ixZIzM9JzWuZTMu9l1DOZ2VfBbbpuB6nVY5lEl8oSlt1GSYS3+T
Qs5qWq7UPH7bqvT0Z4YNXPbWyaU0Cmm5Ez+C5SeYWuK/1ZWKv3yYcjHwjkK+unY5
ZbCp8/oNAGmuFDg+rc6uxCq5VdU9gDbN0UhO1E2YBXd0/O8Jqpih+6udLvLfv2rz
z+XmGyvuJtg7lIL/AwtJFzCoQymyCLI2LkUGru0e2w+tOxk/vKx4kKGQ4RtJ/j7P
9skOPYLis53XynlLumrOTqsNx3bvACHIsLx1iKRNMHnuzH0BVS668jmz5pxNXtzr
gFuaSeaQpnBfL6lG+8pucuC8BJ3Uy4viqc6MnsNAViOwSxy2rKB3Q5z0AF+mnfSh
N4e+wor+zN4S9pc3xl3iq6a5d0XIlHV+uxF83EuAjJRzalqD03qjOp5DrzaTQeRM
HjKF7QD11J4aBmdxFUYgL1v1KmPbBbQANQ/buuqQwilVqSflZ59sw8Wwof3VFCU7
y2ik0RB6Dfra4gj71z8IWKktg9kBPu5cVBs7JWQlxJfiMw/5dpah2A/wqjIcGssp
ey5Ujcx/UzEJDeeupUezNqhAmYPou6x9LjalAi+Ugag+zkikCTUwjzm3s5ysPa45
AY8BXEMTH3PvanIQBUe6XQHztXPjIgkyICoOILCmD3kk0kkmB2vyooU12SrMkNa9
rRMnDirLvrio5t9M5qr0ald7GOIg8IL6Z2LSnHr4zInUNRJdvKXf08RUzAVfz+PS
Gx9kaaOa9nV9yEGRjRE5K/UvMa7syBbmwU7myyTJbPRCmZOpX616LnKYRPFPb2lP
my+EASqHCnUMvv0FusLZe0ifPzRLhPLZ9iDzhptf/qHuVx/U1U3X/vPiuCu+d7Ym
mY9qerx0HmUnDTWOpCHvcNF5Jzd6Yz6omh+gxXFRGmplrvicxw9Dr4Lx5S3U7jN3
vEv6th4eDwTDb0N42sslj+h0KL8UtAzpz8UR8MMrwlKJP5YgbCq1SLDOtVdnQRDO
tVno4gLNy/FtRYRDuc+9AomCm3OORUW5lDnVpMKqWTg3QAdda9pSHog47d15c0zy
/KWQw8r6OEBLc9HS+X1itbOvLyTohT2ZHv2WNiVRmO72ppusxttjAK3tAbCB5Cug
ngIDYbl5Ng/OxnDdTQkqM6hYHhweC8huA5/PAs2gtMznDil3KPZrUKLjUZofDiHX
eme8fHRgsBbh2CT3BQuOWVVUkbyCTbyi8xIjEXcwNqIrV3fnDsx7FdPDsZt1AaCc
o34qJSs0bCYB420DoIP0gWiCzKS1/nwvzEWksD97FpH/toIq/9n3nV55LmQ8KwFe
4w52enj7o3ZTukY7NRtNLZnilc5Id3tCuvUl9IOwLjEJN8eKCMK5pUQrGKlcS5K4
Atozq2E+GEpN6/tiJiHtosye+hIpVgDQv1Nk0eXz3T4dki+I+x6b12DDaFfdFGWw
JSvjEAqxRW2/VE/zvMzeR2MzVhAgPjTEUN+Tt4awkpMOjJ2orHlKjFgbT9Dm5BCk
yCUO4d7PHevI/xHyA27Ejs8DDvaVeEPBl0YrNaGINgf7EgaHXaxx4wdB06x0iqDM
l6I/inuPyZzoCrAXTLz2Y0v5K5ovhgNQTtB2M2JZNroBUfKmcZ5SX8kNumg3Ce+5
6iblwiIAFYx5QVIAueQO/EBN0OysObIxh2UHDPwwdrLswo0H0gpXwA8qsCf6n7Pc
tY/CK7okZwju7MnF2zfAHrhmcSjnUQBMb9ZdKcX0FPKPF6msi6A0PpnGDc1xGJAQ
dpqTlFw+JTgXxoBQI3LXp62FSweHMkbK+mkzsVhxJerjbG4wYI5i7LzA5eE/hi//
a1vA/rY7mj1mQWZ4ZL4pJ+cThDxDAXwALWqBSF7dG2zoHf7t+UnX/LqEipVxvuWI
gFUQHy585JxCxAcm1hYSO8HWHoelBeo7F2Dr6D40q6pI6QuqjW0OiHdBN9IZb0+H
A3rKV07Z1Z9XKYxL6nDKUAhFZJHYmcyLt/3uKZgOgUjLaMjI5O8uZLVJD2qmjHuP
hP45LJj+wweSbj2PdQPh42JB04CDUqDzOw2wmcxnyChsqbSLuih8w++RAdSdfOPh
MLukFGs8IKMGKuQmXoaMJHgYGWZdw59v+oBGyKjYi0AlEOW54/fuvcOa/wL+FdRu
mYpj8aKqIDni0bXsjPlxUp8tVORpJXo2sBfSTRhYhfJhYtpoV6RVqfRF9wFPf45f
Qoh89dREJ+Y5P/HUIK7JDdn9rBjDVbhNGM9ptg/ooPTAKP+G4/YhUywzBoCtMQHR
Q4ysvB2eOquTl6szhBLiKm/uyhdrH04OBEPtbboL3pWzhwSoXDYpSoJjQYzqBYK9
kVWhgkVjUDFZSnEL1vjRTD294xzFNfx/TjHxZuoNA8qLa5OSMEZhAWwlJ5kOuVSR
06bp0BznWnpBnY9HruLpOzaahTqkzlU4yn/5KVxGIGPrCYdhth7JS05z9+sAXjJj
zItVeHsEiYfoDX061nOXfmwj+DNyiaG9M14hcMAgowG2M7e5cffFQu9xDXgKSbkZ
iyH/1Ld4v6aibpIVtvhURHlHYIUsxXxX3Smc94tAXKx0XtRWGvYjGf1UawIJFuCk
Wb6LkFH9UG96cbNMcFtL4A0Q1dtQwg3MsN2cpshSAaRlLsKM53/1VYQkFcZ3Odxl
IwnmWwq7xaSDcw6SVxIssvXaiGqxqcyj/mBg+y5Peq8PdPlD2EZ57dLhsTeQFQre
ysK07R0VwfutBKT0t+7YhLy7Yl3z3wjsSewDRvcNTUIEawbM+3pNwEaWRG7atTMb
OgBhoqXK/zeYiPw9dh6q7k9WwUcXYxJ5BO1vntKpnwImFHZXJIEtA5mFoQ09xozN
Yz4nH6QmDTjQloDtiWyVy91LUeubTiNhXZz1bFRmTShC8qMSlPEjLCUqo3c8EBFB
NHGDmhFpX8pPZ6t7DBqS4+IkBtu9MCNi63JfTV77wHgf55riZ74GXcA57bFQFBH5
ugKS66bfeES2VN6f6OfMMzGYgUGpJr4QQRnA42ZdBnZcDXjV755da/k9b5ZBgQVE
4E0/932Y7wenhViuVraiHSHXOqf6L4Dv0A5M/1htiL3L2mjAgGZ+sQ0keeGoUn+/
SX63lViUfHPvXj3XTEcMaprqXaOXIxY9xfWfLmrjwX3nFWvYWytjb17KSBDNwxbg
eFKOaXx6J5s9T+WPGIguo4KT2J/PNeffLkZcfZGC93XzRrIhl0GZkNFZwoHbFtpu
JzCISEtr+zuoONLjlDJXP6h25eJpAyQ0WCIkjLgHsZivHVtcDb6Yi4bwEbar2qPH
i7HotvqUdhWVke6HjtkccAQZ3Ld9OFbhozP2Ksu8gy4Sh3V1BobzXMIQj3JCKeVK
MHOodhlyVpkwyfztc83rLWbAS0V2dR4pzRJjd28W9Jh1JP+R0ZMSpibEbJI00Rov
C0UjaZAnBg2DEP5qOed2kJaxlKtNJndcmZpT6U4edSQGXU24ZMMHWEdegtMuCZlg
RujFA5U3xK9YSCD3WqvwkN/qxpiGgj+VKAwlj1W2UDIWvxvQinUaPNoi1VEUmKpk
GfOYL9YsBH68YIc2eR44SW0pUlGs5jBTlIRAI5H5KUF9XMPkVzB7eiask5IEq8bC
gyZdyIIeH2TxE5WSrTPk3IQ2hBML/ykdDsUWHhGwmWw0C+5TqGOccxEJjc99K3an
/exmssnGACzRfLbPtR6OYLvb0Qxin96SJURLMgvRfuzuTB2iRSWsGSDRy9HHsASQ
vpTPA5DuPWOw5SrhJ8LJHJmacV9NvMGXwa0w5gIedWR74bq8FnCYC/puIGmANPt+
gxhe1QiI1q+VqSgbv428cq7B4fXvSx7BaSwyy6PMSvhtas8vyUQwLJvvPmjC6OPd
RuggOI6nPfCWGxxpAu/0sRbwdCW4Cywz+fbwH5oU8UICbh6/6X8L8Y+1x95y45fh
J3eK/DeSdeJ/SlQM/JGo2qJi/wxoHZT2oFVJLyiPvs6wJJ43JdYwDMgIqlHI4WLT
buXEjbhp+QG3SYeWta8LnBguSSLmNz17gnHj7eiiS7vSgs8mp/4nq8qFlhXgJSh2
woNmnCk8BEiOWAsJVd23mc+T7VkfqAowOQnIMUtKB6WA0Epl+v/6iShZNlH8ViCn
1O1fB/8HogADu1DaVwgF6O372G5cQA2qBIrtkiAyvyrP5KsBR44UIj+Md6H1aXgk
30xXI1j38wT2SRKtaNmjPWDKKgihShKv/j9FsKBSeMOCNRDcji4h8uaT1A8OT7dV
uyaLqX2W9lahnZszOm550SICQX3+DTR79EM7K+HPKSsHxzm3pR98yGZdncQeAOBC
+fr7Mr/9imak0HGO5u6Tm2Div+BGPCj0nXaiovOe91t8uhn51myUiL3c1ysHhIF+
v3v+w4maeai0+6TwY8UHo2nY5k5cp55OcvtLqggHpH3T4vwcYsJI7zN7lvVoRwsQ
E8eNM3Bp4CJlNH51S1J6WzrhsrjkDf5zgQkroHGZPwRSMTV6th/mzQejuMAVwyp1
BcuGue3KUqNe9My0CQl5gvtxxz1zKh1p3Wp7kqpanU+xW963vEQRopQ2kbtvIsoA
NYx+/kMFbhrVjyKYfyCTUJj2c+jlh/kI4lZEJzbTjketPw0E1HzCosa0rumzzg1F
j1OD8/aN5v3a4UX2OeIbqVgkHYiHooQA+IkmcDoAvg+oi1441yKt6pzqc5V9u6V1
4AaxHUSgNOeeurM0NMaitvV8CWkGSB9zObCUETmBV7NdnpGyQoqfZxnqa6+Zv+uu
0Poc3WukRzl3XpzgjXsv+PzsxFecw5BAC4SVjWRLwpQo6C1QmU+WwFUAcucrmnRa
0FomNLdxrf80CQrtc8HWU/du/2+IYGizQbPum9xmd0Pq+Fy9kf5upH0gfT9qb8lF
PJeukBKwN6zk7BtT6Yu02Yh/NPenC8xyd7bMxghsyz47n+p1oFUT7J1A2mH5rNqJ
NtE5t/VCutibuE09lEo3GFk1cHG9mOE87jLuAvedb0ggEjNYx5H/xe8BSJ6tD7zo
WW+30YmugKuFn/oMgNXqczerAEerE1Bu4UAnx3AX/7ixOXKUVQ9avAVCD7anO8wJ
kgfskHl2k2oko+BjSTWafNmtAPJOWs1q1ugqicNcV4FthAWnyVw3Eb/msjXhFXG4
yYQrbHyiLIyzUDojJvUb6CYXx0knCvL4alqpXYW1DF7U2s3SaWBj3ihTU9YzhaHq
02HwkvFXYwreYI1foOKPmxzQ2Z/JqcpVc8iey7Lo2JynJcHYWrjt/CwXB+3F0njw
GKEVtNwDi3irQLUXcz5Nj/YkvdKjlLsrzEWyjGPHvPoTOJF1/OJ69uPcGULSAiVm
Qkf2QqGAyZUBjCMMcYmnBFnLMreXaUJwADGlNdpfAi2CcOU7IoPq+hEkmbYDHylA
ks2/3y+Im9IiGopMVj0WtnR0XSzm8551gEJVq3Uaszc5FgejJ6POS4zB5K5ipiWt
JG2nldOKA1wqjFSCbkd5HoKfGitBLcYGb84BwyFunQ3q2q9VhK+Ee3U4q1qAOdvS
+u8xrDzuLON0GH1w6XQWKDUOq6b39bamp3xkl+rfR+IHdCpQXTTGSi4m5ZE08GBg
coqwkZpBJnfDXahFmSpFGRt+CbCRwgu+4BxwjsUnVjOLyqT6IGavos1Wj7/BF3hM
9MCVLek/GIxOyVEUJRtQMpM19G1i+2EnXh1FBEEbc70BnALnAg85NPGxiXvCGhfw
md24oqj0AZAAoTb+hWvNe/dLzvgZg/2j+Cbg9hbOtQtNF/BDT7fymFHJJYNpdOsC
ym8KBYXXItqyp0L2WdlAISGh0iCN1JvQeBoikNnIVA1WBX1rOeyiuJhxmDVjucyw
+3blZZ5Lg0gBZk3tC853yfvwNFu49mbCPNsE7rHdn5fAlCQ4cUBxW29TkGBf8Kr9
8vQNO9CPnfcp6KDMx+kyILWQE58nxs8SJx2DNs390LOT46c48TJ4BKNMkCAVF1ju
7hykT1jRkVI3WTD1PlncZgteKneMOMC/163ULJ8v3PFfKmmo/ciU/2g3ocfghPAz
y6nAr5YBbXYrY9hAX2YxcoshSa/cCu+X1N4G4GDVfP9+aTlkSuuoUqO+HGtB1JWA
TOYwjtqs8onPjA+aUFz4TngtnfQQZXkpvt2TjLGoQSXxVIy8uoeKITt5TIveZDrE
eUqWjiVnZ0fdS1qWTNWHcibGUgvzYULUBEQkto4hL1+A7OHxOUQOaI8c1rm+20KP
000zEnqUR4ieIafN6pnYUrjkH6eW7FZuNj3j/BEURV4LQVvh79NRrLonRsex/lih
KgsIbS6ydX9on82HyDhCcM5ebHFOp7OyTwV560WTIPuvhcNW/mHB+9UExafA1P8c
fFpIMZS6/lPa6xgRgk7i3D9VauSIVcZlnOdls3mPIZnX/5kexiMDOQXSv5GHPK5b
aMqG1SNCi2i036AMivW5eKnZo9slChRBKdEZieR6tojQ8thtd3cRIZtvMnuU/JLF
hUdnHQPaaDZgeg4wRnqfwlXDdv26L1QuHspew9qVqWIsT46RO9t6NE+wvcQhMEAX
vwiH4pUtzhsvC2UXQ08DuUFtnvhKsoG6PToZ3db0pI36e8WiHoHXAjxiayC2wAb4
tzjfhw/XqOVOAhGzEuc325fBtLUpAjWpP4MuIwthvkTcdEQPqrP8+zxIlYFUa78m
jJpjYS6bTsh5JQo4UsRbucdAfS6T75bildpDThNoPz2FWqzyMuB9wm5f7XRpxGO0
crGCygJgcm16JJxr2Fg7XCDDL9v/q6evI9ZnnmbeLRfQAn4nvfoHErgUbPG5UJky
yHgtCiC1EfbQdsyMqupt2Zx/8p2BQtcDHgnnCD5t+xhIjH0pYJjW20bgQDi3WYFe
5gzKlchrDPYSiGY3H7NFJ8NXKYB6Go1KJlXoj4Td32NgNkS8bacpfLxxl5pykSLw
SEY+zJbb/6iVmfUQYeQI12pWK+ov+CoVgCkN3ASTu8IRito5xvJn0Rf+eWvhZ5Oy
KCkYEtPR2+vIYo0p09Fs1wyilH1Fi+6MyLjymYm8+0b+RFInOc0uH8XtAcjHZO8F
/QnH+TplRw+sNbS5Anx62hbS//Yim6gEtEmJocFKwS1Oc8KkwXOYd1ZcCLo2yZy1
bR+S+iEB1C3ZfFgG6qz9s/K8+I0f2vK498fUYD7Q/kPOgQDW441o3dNW0fOVgr6V
2rQhSNetTbROIhyN1ftu1eCT+3AZYc1SqU4ekI9pTw4BAjsJdo07G2MMHtXh1tB4
GnGXzghsyFccEvzGhdx3ULVCDxjCT61KeaqcLYsu8mUex8P7AdTd4kfM01ElpAoy
UHanBnflQcrAeophZqHAEyBd+mza5E+oSsJTR9ERGH6BWec5ns1ldMDwjgThtSd2
imJ6yZ6UNljEcQ3VXb+BGunum0wzvhzW3X0SIdvweBnqEwqsQ3rAzmZd1uXy8hON
7aaNcLDyU1Jgq+fm7wSpo0Oac/sqKhx2ESgzs/8tfDdGegXY9SXANCli72YtJJi7
KCP+9WneE7MJQ73jFDQE6Ph96Gl3MjMj3O0M4m0DYynFgztVIiiKB6b8AGq4sK2O
8Hww1F9j9tgfmupU/IsmIz4QHPP9ftvOTejWkc/O+xV1UYhQf1VCu/8AILjCGJm7
HMnBTNueeXRf15rEQlsgOQkjImXRqZJgqdHJFUYDrzvrBuTqPNDH4/agxDo2MMjS
H806c8d0PEhX9dlRnpwgezLiATpsjTjn+TcbhH63Ph8sOdbNt3npxdPqoz8fMtTM
YZq5SHmVojGo59NITA3d8zHIDt3nhAsCSET+qHtbDYXMS3MCs4mh3MqegRPFNelA
Yliyz7tnjkrs7t20jO3P+ZO4kRwNPkP1S7/9h6+fdT095AZ/wYXTmygNOGkVNz2e
0rCe7VwsgMbx4VaWe+NPqsN3az4aB3cAkmm/h+AolCkS2+IVCS3VAVoV4CBoa+OQ
NkAR/W9IzoUXTVhul1LeMjFJKYwny7akPY5WcQXIoP1DoztwXU8sP5Cb+2Y+soso
+FxBnVp0fGPdT6Ed45KKqA+Bo8KL40PlVgi7J2N0eKxfRvtvCYbfhZnqzNZH0uRu
EZ3StA1FQgH4k0LsrvPrNL/F2beIABK/Pgk0XxCbKiMym6QkZn4XgC57aSnMvAeO
8j3BkIU8Nug1jN3gvWf+h7jNiKMhCXWM5B3MGxjIUbd1GHK3VLqrghooqRGwBOTv
foLWvi+AO7Jv7czv2pzx7uq/Hv7oWdZfgBEFQ8whsABxM0U/21RT4EqXRdIcXjL5
w0GfrPTdcjz9+MktEw14BvZY1dgHtjLV3rubcuFh7jAcyM9hqCCnMIcJCEBZjrse
o/Vm38mgAzzEeXieZdEqzAsoYETcLxWkv+P/Om6tOjbd0OVRzfUciTUaidIwlQy3
pZi3yGAcWvOXFZ6NdJW7Gcn1+p3DjQRyYTCUiqPXtgk6p7wWXXqk6jAE/+zpLupG
MbRP3YiXTO/XIYPflypRxyW/5+yFn7640s9EnaXfngtheF47sIIkYe3GtHGU//97
Qfq/Ginf7Pu3q3GHjVjE1pEZno1d+ljsGQzyYD0svZn3xMpMFHNVwWq6Ni3DDkN6
TIb0u4HjVpKtIOI4y3T2QNLGFjF0ZySQhcB/WDmic3jMsGpthCB6v03ZupRhhKhr
C+QirMLJo+B8X5ORr8UOw6RRx0QfYkU9Qurfhm0DT1jLirjYdn3v7188fyiP4Y2Z
uV1dCQIfi+9bEdqhaAPsGKjR6ebbFwgNQQenBWrprrRHBxgf8EQuyAmDTdSpWhas
pfy9xOOzpx+pOJvmebre1EwmfHmF14FXWozcHvJ1PQfRwimphGh9nmqXCxW8HaZX
FZMztIM3oqP7Lkxo5p+muJ2iHAK/lzG1sJqVGGNNinHuCV/QiSz+bMIN8cpfDsZn
pftJtJJ4H7PzKPK5PKq3PWJw4K3aRmZHoL9FRhCHb4NGhs9nfsoMRCM18LQYbH6N
x7Xw2zF0+B8FtZGiKPibxRJvuxiC4c+Bd6iT7Pwqm1k+3gIRt/1rJpqoZj2oG2DH
nYIW90fngZVNVPQSdMMbHOeOJgP2JkTkXmvyYImsYZa+FZIgohl4qX5fm/YvDZzL
ZbpmKiqjqhtEGzIrqKsWz2aBH1wafpclAOd1vWbGdFQAc2NsCjDMCBQiao1pMZOY
nj13g5z4lTOX6B18LlaJKeR+n/linUGCSrnA0xbYx2pHaB/o2i24ilAWiak11V30
Gb2JkdRuK1pX6Ocjyvtm2YFPwwfrv2+7g+R+mAkNAIqYP7KEv1cG1H+AmRyHOqmx
tYKrvevCuHk5Kokb11AUyKlqfspGxMFu/W01QlU4Z64H66TJic8lTj6HUdCDBwCG
UAHxYe/38Xkru3SoxszkISlhx5nBM/tDJOgeGSgqWqJdqR4oxHFRKrsr58dg1IJL
/CtGxq2H4k3UgtrM9N5X9v77di3MPEnOaZVCMIwdzD4rZYk2PjHK4SU0rQ+qSa3N
ZuTywHGaHbS7jPpMQylJU8x1mfIlOZj7B2YoAaUnK9/G3S0H/fTjVDIM91Z8S+h2
ejbSQHurzi+dy8gBrXPO+oExzayUX4aBTRWiTOxWRhnzhMKMdXilbs6ANtcLInKx
kZ7zczm6TJN9BRvmr8SK+I3h/bcJ5c1Z+wpY579zHTz0YsWOfJPachwPhF+TaBk/
IEk98W1i7vEzUsSKmT9hP+K8HPlqqpGqzWtAT9OF8ok94xnSxVoHN9ROm+zR0hX9
0UdtdCbrGV2fzpZKo3e2R4Z86nQk680QA3dpR7a/LS2lb/4Zj0nMDIuAKi0lFoR8
FAo4CDlSwYXPEiWuuF5p2BnwnD1Rvy0Gv9rh/GnJev1VwkLip67xhN5juGSYXLRJ
llzQGJx/Nd8Pmrp3nDJ3h/3QBHxF7bR2F3vrDUXv6mbjBOl0yWjG5Axfao0Ckxbz
h4fX2S66M1mnevEarmBxCRxhxC38BAjApSzPwkk/9JVAcqC8gPVrt+O8Ji0My5DH
VFpUE8PtzlXJdQjlXNwQdueaeOZl32st1u7FJVOVhhlLgmC49cHL2e0mRk4xB/39
7yOQA9OBqSeFC69udDwSiyvdOYOrBkAJKb0Byz5cZU18kTIlcy+L5zNr6sPJjIOG
jWg+vsPfeR0ouikFPeAE0+wczUm+BoN/2ApHxU7Zb2+doMePtr3i/RLmdoNMJLXW
lKokh0y59CgOfU8T8Rkhkhbv4r/oneV4MGSBcBNLOcJnTYfdEXMDdvkpk3nLRri8
v8ldjOA2lvhmuqGFg4nfrutGEA6j614/FaK2W511wqoczw9+KePAe/uNV9vHm/41
dFVRc+SueRN7Ps2LqZMnaeJpuAE5jlm98oP+zwfP4o4AnfLNEMNsbvhXAYCNunb4
1Bangmk9rJ9c7c83clZk6GYnAFZn54/I9tD+hkawYF7ktu77vfBnPBiiTiWx/4dw
yHXzPDr7lZUMSOdkPhQkC1Q9d59pUkvg4yqNRhWI2q7WBlbsRYwQfq6AguZiOSlA
fJSP3xXrtzqtlWbdnEnK7e5Ap6BOsoO+2nGlrUxXFThced3J+nV/fl+qh4ZA3Gy1
w19ivOX1Syjdu6/yVx53ie6X/hpwQlh4W/r5oDFgkq02b2PaBzProoF7QOvsICDg
tmRjBDoFY2NnituzfAebA4aZ7lBXLasZbZyKws1uKuZbq9qRQjYbyIklH+lX2H+i
uS70SqzCzbCrgKiY4rNuAU+yUylwhY9jEddqM7warO79QJgU6zln/QAy78R8KZZG
rKNFZjIJJ29dvL4laRLXrOQ5DemAVuwAqW4AtT7SxUe5QRT6UoABmomA0JvVrPsf
jwVnYHiK1GgSr4twmWZDcNHJT4YI4TjCeKTssiqMpzhr0RSHwfvr0uC7PEArdK73
Hr333fetvPzmcfzKhpm5Zoivnp4n5XaXv7flwrCKezR6sszRrLNGKIYbHzL7IpeR
OQkGZ1CFU0um9uRCcfuPoxDAMBn3NfYJiT2AJckWUpksLvYdiBsuLJLRitCXLxAH
yZpmLMfrudFEd0WR/hiouXzUfdS2bryJvTpmKKTd/7vCAw4K7QsOyKwgnmtiGwiw
uicJBuaBAwP8SsfMG5K9UkN1ycLvacYWvQymbXxnl4W0KXUY6cUrMjp6VLzh46xB
H5CgwFqMhY/qZV9SIVsqNswoWKV6sPWPESWNCrlXXWOJocCgJvEJvOvNkU/gTJ3x
EW0R9YdZfprKDX8d/VZLUwCyWbmYu+yo6qWhdwvQuAhyKa/c6aN4cDdk/ZJ419Ox
I98OhnWbsSS66uCfTKpCGoqfEgk6m2YcPkEQZmJS4onu/oFjOF7eT4lVLdoAlyTU
8hgGLijWlQMCY3VVKoimMLxxhiiZRKjbaSMaCGJthG85xiaFUTn1mqLBC3DK/adA
16duFrobNqIn1ou1Us+00VDKLd30tdZIXc9gU7KIwhiJaBUE5TLIPuPGnKDLJ/dL
ldSerC4942AHTJPud0xz1Ma8FTxBEoOUxiBJfa6Fv8q0Iux9Ha+6S2QmaBZEJN38
/XzCYOxiogVDhoAt6r76OpZSssaE4jQ1NcEu3wymNUErtbAFBdpx6joSVJQC+grW
M9kvG6bJ/tmRrQMFb6LwS/KfF6pHmCuvEz9PE2aUVetb63hrUn2+vdy8Fl2hIn9h
DOrloho2I+yx3gIacqD6KU5rnHO1qfMSSQ1cVs2dKBsmCYashvmUMuMyQMIC18e6
AbehlKQApxchmFzBWubx7gdQyjLp3RlS+Gc1XCP3lhAIfdj22hfWiOCMKTVxz5jb
jWro3QBAD9O327QwZQsGB44FM72O5HNkfwxIcn58vWeDJQ0Cmm10IN6gltaWziKT
CN1aPUpGR/bda/s/8R9NNOeZfgvzec3kUOVTdeDFiwpFWEQio4qR824YGfEi1wEV
FDNFzk49c2JLMvp3zXfBulsjUR1ENqtk75N65yxT3+I61CmMfSDKK2z361QGUl37
18Vig9OsHscYggi87LTYkzXVxy96WdlAGRbRFPilsWOdSzXFQIWZaXw8wm7aDFuW
fCbowPXDMyhAzusQc1/v0LiH2X1tqztUyiYq1yo/fDbMG14m5d4+PYVH1qn/WzRH
Hjb8CZZ0W3G+++plum+qiFi1vWIEpGYHuY1g1UaFcrOO77bwfaiEV/Sz/LC736PS
QQitSsWH3lv0uxrJIPZ0G889BHai2Bkm5vKe6/YThQ37lDZOe20pBjX3vbPh2Atc
dNEYmLDVvSswqA+WHISon6p+ytqbdZpeZMShSSj+r5U2sn14Sxhok9i7cUetNGIB
4MKcvakjWwwzl4N8YrnFZZTWv0LysVe+cydbW33TYtm7myVF8cgbrE+kkhvdlrtp
HL+6D2V9auUy7iGzmx1ahCWxRgbVC91kLnaEZr+USxed0m6Nb7/fDnT5XzNljcfY
y7P4bwMlS4YqWHZYNubte5q7hBqy5zWnXEcQeb7i5mnHP3OVBytK1EKb21LVTnY4
1XCMCwcRvluY/M1OqfEJwF8x7gekpx3/6dakqNrkgcZ2bub4MH6nchAbTVMsUbgv
4m5N6nIiKTfixj1t9zUaw1vzvgHIIjGi0L1xxDXn56xTDdJ7YleuTW/rH1SFt53S
E+Auefipo4EYLzb5Yl0xzBGy8hHcm9CDGr8SO8LhDn3EFTc8yWW5k5iU1oxv780o
NFZKKzXq6RhTkCd/rdz8ezRdt3Amks50wsOLOe20vvuksUGrbCbElrZkumYP99LN
Hiccnvd7L4d20dvsL/Di8rzZkHWDSDWi6Lt8QzuIoIduzSIeN23UhwF7yndHxVPH
i67ums6SAuUYSrBHL5T3CXO4MpqK3Z4POYH8bw5n3Bz101niDji/+EcbP/6E35xo
2byMGo4qIDumEflB0mRFnBj0XXF4B5klMwMoMzq1YfKF5eX9moueF5ccVijkjygk
zeRymaKrO8PFAEHVzEghMONWoGZk9somPgR0HKxQHSgsM1ou9HawPP7KXfKkwG2D
hNoxJl2AJU8qkliiH5oGX257+vd+NgAFVxwVCYV+tgbyWN55wGOCR4xLAeVAney+
gQvl41Uy2KyxGLsCV018WULZMQzX667eivkS7ST0Foc830V7g6vZudHLVbh5LOR7
1iuUkNseo5YC4j6jW+FdyBMmXCnsm8A11zF6M1V/ye3ZrKNLvv0UT8LCPd0pWL7n
ElqgIGNqYPQe1sWrn3ERp/93x5w5lRaCxkaU5joA/6YamumqutpUwPNbmbErHkY5
VDgtuRw8AcHMOggsSSFpCLHjvj+CH6cX7MyPm1iqggkh3Qi8FfMgwrZ0orb0/jPo
GYIP/UhVfjrnPKUFDcFm3KtKVrdcn6K3cI8uKTNim3zAAeqn1vuHEfbFuvu1tO12
3/12+zIVtIyMk1qveKrrhuBJFqNqgeunvZWvDIgYf+CgBNDhhcSvN8QD5WzLlhgv
2/uWKTRGEmQ3ShdFUmb2D2q7+rG3tmcUDRtoWwp5gZ0CzRpGvU1ubiGtWVro/7Nd
Mhaa5ks2OfKaannREPEsTDVlDVgA/KkkbvA/ukh3ZADY0BTx//Rlbp2zEhOHlbXo
yLwb1j5VeFIb8bIRv8giw0A7qzGFMeU77R8N+MvV2XUJ0+jJ2GR3ynnz0zsS4VKs
WqMe2QrfedOxYrMHB5ID0rGsm++u5xom7zFFLtv0rknM3EFdkS7A9qyQjqoVYdTZ
/a6r1Y3MQ9dPJ4hJ6gRsGXndto2SdgOsluIIQo8WfmsxIsyKJy/sRb0jUZ71Enfh
M8U58DlIHPDRADLaiJ4yKRGnG/R7EjXxkXXTqJXaQGezdDhv24SLiTsIPNu24Q4V
ZxFwhZtSV5qkSW5r+TIG+MWC3OYXqQP4W8wBxzUV6xYAXD/7SMe/1qIGzzmvlPqd
GgrsAN0Zy3qln1FEFg6coPB+Bq/vfoAsxQc+L5UqLXSnUIqOtvxBlclOtuZgrfqx
YZRG5BpvndxykoAtxPW+FL9O6o78GN/VOltlNgArfmN6eTwxGAFvUs+4GJH+v8C1
XKg3a0Wy3ZzHAbJkn+bxweD392j5EiCI2l680yekaud0zAYvGW5JF1zQ/PgIaZvh
okFxhWFzEAO4ncwrse1P/GXOxOCVbhSxhrGVgCioE0J51gWZc2PuTeFu0cELF/1h
2zy6h9uyxbR3UIxKexD3CBQQjlcPfHd8FGlmqUVlurAHNeCOdPsaQzTvaWO9vLXc
5QTyxonZGV+D9PPddQhxF+yUDfWNIUf2jbK22pn7/TPMBCDY19joVrnuwP1lt4mA
eXOjEOJ+Rr/ntlhdtul0IDHUaJDCupm9UpSZTIeZxqw/PDBlxr7cJNujC7I+PtqC
ghkoRxgIk8ByMIxN3lNVit28OlVxbX+Hwhk0yyMW5ZrGkZcEoUb4mznGulbuk338
KDGuXdCecNU1/QSTtFwGKvvSgvboJaNZgtCWeraoFEwDvyyQhgcYcwEEc6m5PsKD
ogqNySXfWvLhrcKZnkXQ+c/z8t12o+PDnJhdNjSfe5qhPXIwZBsnKSBU2bDJxOl5
94QG1mhS3dvxIlgdC+9Cy07KRj7RkpgVe5xM6kSafd6d40imyayulo9o65ybx4I3
rjJ5TNwzwAsIBit0+/OE2q9b3DNRFGne/TefMhbNpw5Oem6AxvlhKzUL1b0f5GrG
54mzZsPIwfHigljcZOvLJ4mq//Go8qDTpmSjXKEUo/VTGStOfUplpZhdtQjLbaZF
3E0S/W8cdgQGbK9Vqwv0bCt/84zSj/bOK7id6ClCV9Bu2unPswWd9yDJSU6lEy7D
jcsQAbNtN4dkhbOC+AGX+HSle6gxwjXvI3j3gyRnILVbQvZXm+LMukhkd7/wXxO+
HVD/g8ETojk93egvdRg6IIRNVvLw22+8GP4W2zfseD8UnWppaDC5pjnV5yXcXU4N
8oa/q6LUQNEhArcrPl4USSEe15v5y9ctiAbow9fmqlZ86qf79pluY+vjs0lxkRYx
rPLf8cw4v9pz6CmzZjjnyUlUhP3+73HA0/2ch9p4Av+UtQLl5oujXth1yHD7ehxb
1sUeISZL4XYYTRMscB5pyru3YH/S0p0ayf2myQWYSh0YWdZSk+YWvFfnGiCj+F4D
UY4WctsG3B1kjFoIKfC99UFVjNCt+d5DC1zLxkKgUcTLTvZFDyMXe/UiAaNPSj0e
XPRVP5gVTJ+U/rKxikuq03Cyeqf1vN6XlpiUtEGJl4LQqMyw73jwdkRYvWllWjbU
U9uV2uQikfD4+W5Bf/Dgc1gLMZ6+UOvw8Vmdcsxz7SbWelIH+lUieDMhrWvmmuUW
o0vMnDudJUoMzgN/OtML/nN8+ygIQ78GO5w9yiPmXrX/AQ43Q++rXzNDQa7UmtmO
Ic6yeRTQMAJxSNwKNCO2R9MUs5M4fZ7lAaqwmXajkQwvknk9BWV5vzslABa73Ehk
/kTYk7IyGbztjzW2WVvKaKXoVK94J06vUwykqDDxbGchPBa7VupPVa+EJquFvkvr
2E5O/fSYPqjtyZKxAPcO59f3L6qPUMbo7zd7o2NE9u9RTyGd7PJe+iClQI8JgeBs
RUpptRMAJX6XeKFOkUHhnzmxCEaENk903/iy1hTma5iUXjwlcTvo/QeYFIkB4b1Z
UK/G7uJaIFkh1Y7t/IvUpqbAnJiixtgB4Q7GkY5dz39Oa2LRCeGDbgimm67FuvZG
Y8P4x7ejo0Nj9W6xCu6UlfC9c5Laf2McPN9yfMXWN1m6IT0GckrwFWatkjXXEhT7
4EXBAF0zRABkC3JNZESdh/NhMiNG9bepbWRcFWvvU2nD/aT+AGOOYO+211tw4hIV
V74rPYgt1+kiutgqAt2BgpMJsaYYvRhxh+Z6AdbeWGI1J+p3D6LSp5WkfF7HJfQl
hEwjpC+FBLNq6kWrPqOmD/kZjVfkvth0O72S1t/SqaXqE2GQnSskXAbUOkZ0SrmB
rcOVFz4F9dOFtXvrzRgX0I3lIKA/Lv/d3FtcEbPYHMgwhhNjjNO5Z6aJkiwPncD+
+G0/Gm17IcTfHe790ddGn15VuFiRao63JXJCjsjV9tt4Hdk3QZTFdmUolBrokojw
Zb+EwuYRIW6QKE58XT8MsQmnYRieknbOtM9NGOha+h6GjyqXcrLkj6yy5KMW04AH
yQto1bRC/pelB5I0XdoSNfvXMB7wqZ52OtY4ivFUDBAFhRKfv77QbUHlMI49klAC
rZyiSpeQKrWKb72BKkkwhJRK+PHgnBNZk7ua7KNf/GbP3ZK7tl2e6lRmNQcPSAK9
IuMpGt9z1cuHOqHcqV+kzKq4mypRfO0BYTHwBre42t6O+i18AWDlde5xhnKFRx4b
9ceOEcVsAN8p0M9ZlX1aT5oU0Reo3Uo+hLfJFZZm4znwBUH6aZZv+PyoZ9i3bE65
SU/obXRG28YJun2uwv+wXiZR6kUJungN3HR41SraS3agR2jpEtItBNJQRyVWfUbd
SnNN8eW24fJPnjGvtVSGKeKOIXypEFXtf6/xfz0R2uvKUQEUh0MSoa/4b2lKD4tJ
kuDbXzyLYqDc0nGD+I7jO5yt9i8F3XyIMQQdX5D9sV3VXJQGgMebW1QciqOUu5Bb
DMEkuLeCMOQdETM0f+g5Kgqi1iHDZM4YfotGtYs27f5ErFuOyyM91ur+aVAiibue
RJ2gqyUVutxH9lsMRuD2zW/3NVGjjR+NAsiho/T1RJQ/E6Tho5JdsyeoM0TTySCi
z1M0/edCI32SdvlbZ9kATxTRl4zZuqz+AsyYNtUqO1B3VIIKkXEaJPP8LhYBfeN8
w+XIs0I90zwyyqB3KaFDNhOllX66/Oriu/mzLsPSFyg2FJy11viSq0ewnHFsiJf6
n4PE8TgE2YxcilDcprv+H9xZh0XqdjqnDF9ijezzfNq7gAvOLcKrtjea+lWI4/Xw
w1NWbZxvt4lkrf+GSCoWxaCjqb5t2zEwCRxzA1w0ywmFWKiq5kkf2YWxd5op8FcI
dycyWJ3Up4dasi6piGelLK7gVa10opTWGnbuM5I5WYDj9KMrdYxdqJ1ptveYyCfb
b/MAVcRdNMbixiy6QvGcs3CyWahlmd0cBwAHOwGDxFqN7I3nDOYDweatUJtRUCF1
THazRWhFBOK2OU52BII3xqGtojitJHbB6DT/Aqnn6iK8ICbAdQc1Fhsjl/cUstoK
rMzp6QaibiGjZ+87ZhOISS19c3FUJ3y5ya+cFVPqAibtxR14QTi/Q4JN5q6vxNrB
Ylv4xmH1nosmOK1A+mDiMzQdXKgmowsKT2MWNekZ9bPBgHgs+xhsnYnyj1zYQ6WG
vwF5glMOTa2WUVKulfdNRsexFwkfLqoUPjzqkNztoq/OrtLWIG+iDYbRJRX+8Ylr
nOzTpldBZ4Q7iTzRQee/qHKxKIY0S3p3H1OdGEyNVteHC6RHGW3GQ0ZCiy+QpR9F
PPn7xQCgIy1a5WeDaikSBW8/Q5Bd/TfM7WABCjZK43v/n4Lf9WKzbOoy0dpbbkFG
N1P49Pwxs1yJmIsyuV6zonzqHsyIQcHG/nK/IHKcYrE7C9M2+eopHAreVJmG5LRq
rsjejTwh5Ch2yCObnhC/vnSReuzhpne3LwCOAP0liwwernIYx8mPVYQgLiAnd/WJ
kwyWBi+w/dqefYUd8XbelB+rE0zr/nPrgzVbTTc2NXqXsI/iNbQg9vwRislU6Ib5
Abpwz70QIWKGAgAHI7zYINmASSq5ctED9aDBo9y9O/nl2odlfghzWl6dl2SBrGo8
sMa2xU/iO+XechFEcnK+0IWNQWzscdfuPaw5wF+0Dpz0oEH40srTufNevlgR/Mho
PmODqQo/x7r3bL7b5ti9Bd/aDceWUrYQesxrwlcccGqTJ6xdb4U6LDBeQo3VH/+O
+g5TyAMcyAmAUrhBnQRlXryYzNceqQNDDVO7futvm8moqjJ9dHYBMehR2Lt1ke1k
suDtImLOOML34S5yY/eVueTLty/BNFbqog47QXrL4046lNNefwiG6RObjPPG2IPW
hf1bqcjeIvd2SrY+7KDBYgGkz9OfX7dO393Ll6YQtIEn6gjpKeM34xvgelrnbaU5
c38+xc1OWKFiQnuwIJ7bjHU5V4QoUL36e760wga5fJYFkJdN1mcPDPuy8VSRMqtw
j3by8C+YDygY+S+yRD9hlD74MfxRd2gxjdmU/7wEUiwc3XQPFtuymK1sGvtm5Xon
l+c+x4JT3RnDWJkU0uryvMB/vppzozW8+SuT5sQkDUOUo2w1pfXReGHDbE27ZAbJ
7kKP6c/PrQ2OVO2Pi/lHVqZVZ6OiEbMcfmTL/213FIQHB1Egw44hCSTITjH5MS5y
Q49VmSzBtqhNL04E90UgkM3ng+nt8J8Xqc76yj2hN9ehQrGxYDCWn+ECFsI8muzG
UepUAYqe7dioqpUtXZ8dY/eWmu60PWHaDtKwubSax/OYal1yL3gTf0SM38Us8Uc3
TeZJqm7swncNuYPBCkzIvTpTb2XUN9d9eNWX2YMg5FML8zHzM+tr1DkiACafTdO9
U/+mdyvLg23v2o+eZNN4hINkIyj5wGAzseo6L556Il3d2/C/VV9s3n7YeRb1WvnF
RXRa/+JCyFwS+UgY7vAGm4eCNJSH4fxLMx6wSiLNQdqY2E7ZhvLUwi5/4b6bIzd/
KYN0TBLcpIcC2nDm5sUgHafOt1g2LmIp5V0Nl0CUlXR5otLSNjbWVrmJo9ePXztj
NhkWLhQ5kpdMUhuJ3qk6W6MNRYhY/vtLLhZfP0nhJPF9Om/N1EqwBKwbDrW14/Ft
K+NEf2Bbdjcu/oW5sIq89hvbAK6K23nbsmG8+xDFzNyD8povRPxPrcMb4PavcQ1r
qw78aAjj6kAKXsrIC6W75kj1HjJpx+w/7XUCwNf2fKPT42vlH9dVp00Cn1ahkeCc
I2/Z+lk0QscEDtRIq83DOCeP6ZlXGS9Q3SpCH/5OGQNBtgrh5lzbquW9yLRWsbe4
bWyci934Bf95HCxAhTR9tQW1BNwGQM9MWQiz31HDFgi89a+gB3qiHOviT9lznKW6
gv7sTD3Vef16GMNt1mUwlvkeXH+U10L7IM9QMuNyJne+5rk+YY42wTpXAxAve33L
p7YIF3EjoxxzohZvEx2arOyVNG2cx2C8ps7r7hlzSzwdi6SXm1hB9YJn0CMPZEUi
DylkxifGniKVsKAa46TTPP2dTkjdC3ZxVgGc0Uqof3lxta8Ci/O+kagoNHWtU2EP
qxvr0XoWojYwyuUouNydBDGo9bLi8VjPNeMwTaUvZMwpn5uml4O21Hj1eDgzIucJ
iUZeslg/L8w/CCCOv5BTeKcMhcZ40gDdRC3K4ipJ2A0G6unLanEqUCD+Cah96SxY
gkzK0EZdevnhSX20qR5MgbhQXzg3uWb9KUvOrby7x0uQbgK5qdkdZ74YNqvM+HrL
goreY69r04N9R16Kr8kkvsFcVy1XwU2shKPBquiEgRbpzD7hULLrrgh2l5kjo4Ck
I8IsWlQtcSn3GYw7vyPu+jOh06qZ6Vgf4jjACB4YHlj3has9c48JgiZk6kXNdKts
m2aSM4/jDgp4Yt+89Xvf2FGHtXXNP6qUGZWc7C5rf9SDorKLEA+gDrbdXQ/3JPKT
MbP1spR37983Ok9L+jJzZO+M8zUDNbOJftrSbyS2BWD4XXy2/3N55M+4xnU7xnpF
sL0W3mB8WxUUBQ5dQ7lEVwzMXY33d60+EI/ztSo6VLpDI2ZAd+gaVdp7kmzyon4P
wWAfe/IT6Ljo3Pq+6e8tmikOZsgw4vpeoJwePZHz6nNMWFWgqv+cI4s6vB87aMti
jTeT6HKjYeLpEeuNiwOP/k4b+SbPAtxsic94Bzo24xC5puX0kmlVKvjYIBTx7bQQ
UQTbi2Sp9O1Xi3cMb3vTuJUw8zNRy1Ch3BwafY21O4XlADxenSoxMq4c8zrb26TG
AB0mmBEzFE2Z66n1xNXHrvPUuMVigUjCqVtJIiPMtBdRqk2kYDoeAOuWV78KknPo
Xf7cFTu7uczLK1Ldr+1AMjRVBMatGGdK4Xe5BRaVAn/eJ2Yb4DSoVblbZxB8igD6
EzzhihzGwHA9f9izOqgjOue63BKS7iH9btSCbIWALGds7G7DMdtzE+iFuAT6OqYI
xgB2x14PF5rRi+oUM8Zujiq1GLPQaP5eAYWtm+ueKkGcTS7nIh649gzXWyFVWCZs
z0p44+a5Vna30lnlKImtWsVHlP/EuO5KC0P2nvI7dgrUjOsgZRLZfwLlqlh5q74x
bud1M3uT6byfwLs7Lljgg8JsGQURkqUsCs8vLacs7JMwvOnQFW/wQSisjHHFmZ3R
CF3ImwqVd94OjhBaQ1z0i3mlppi3X4fooDqgr+G+FBM4F0OqMKT0/GRkftsui2wf
uCmXCAF0j0qpChwEh9FaNrz7q4HUNXeqkX3F9LRuaw3rYrFJZNy7LLJ5W6F6y3C5
/TK3BS6w382Z2hmRWtODMjym8zBSXU95NsptSFi287uUtIo05nKfw1KNwHtw9i+c
5GoBe/MqnQPm6wPJ6S9H2lIgQt5zPSgrjYpDWeUxHS9ryv8zK2r7xY4jW/OOOqy/
CWpIF6GANaC8+0eYNvl7emfFuL5ESJtwGE/NZHGeEkYM7cN96afaHLIKtap5KUge
rHM0gwx5UkoXsBkx5qxhn6b0GFL1uAOHzy4HOu7/PHajIzNtVfsKE0aPRWCxp/Vc
N2BaFjoO6XrP1e7UsTiOalmgQDwiVpj1c/YDzEvyAOhDMXtWk7uqVreorYN8n/T9
zc9yLOBzzbtZWzQomeNymJLSnR/pjmu4aG7jmALJlLJUEcjJcpgF1M3Z43z92DYL
+ZLf19V4ml49ar/Xkv7PNoqMjIM22jy9cEEqmyBzD7lySQrCzCZ19a0kWA38cLus
bjes/Z58jZ8lllqQ0c/pmP2tUGruhVBqUXsWIXhFGA7eiCVzcvgj78AVLtK+TR6O
8HRVibNZ94HyPG77fA5sIOPT8+q0iQLeJu3lltR3qfPidGNmBGWMTKjBBfOhte7r
poJGleBfvfs3LvOpTHFHPMAWjAhgfnElKMotdbFpLk5N/8wRx+h49PjlNJxpJiYd
02PvFManCT6Ysd9H0M5Uq2Z9SLOPTB8/2Vd+WHrln4+HSvHpnBDpBDNck8vdsvNa
762/ktXlLaj/kMYt7CDBv95Yxv/Fj5WZj2jzPksHS74uTyp1EheTncItZ6Zbg6zJ
xeDaqAgE+EVIFC5KaT8yB1++B+ckImMqJ5KDA4XIthyRYOisZv6NKq3+puPtP5Ld
QIBlfBgH6O3Ltp6BCjykK2pNjLiItQ7S9TD3LMUF0x8lnvuke0Qfr06ULKCDAhWM
YIXSwhLawEa8lEBB6/Rwf1B9ylS0R9gHwbKwad8in36h+Pm00ufP0Use9YA0xe64
jHmN+1Di+vCDwRgOLtyqbBAZlmiOLPzmkl9Do84YmgMBOfTvoR01Q91nrCo3J967
lsjCnqi27RMGGqhSPFEblDySrGZMmuVevspde96Y1hAqkdT/7jhDVwa/bdVDgkkS
aiaz1ATYvQVPbiGOK2mT4BP31gFsnb8qtpHRy1D3dpE9fEO6jHD1ZexZACBqpxGg
f7cccoAS8sCcOKZJITxwMPNYzFLrEueY2E1eU8a2kqYrfWsmPC6wgE553uQ7Gtqm
QHZB1A3uhAHghEMJ45UnS83TFmgwwoaiY7dsCR1Fjfpt45s04O9A35VP4QoTpLwC
W3zRDivO5CpaKwUQnH4F6Mzy36y2E10rIGLhL9LK/VwyudpqtN/pZuWO4+3bOVaj
nj/SQlT7Nv8o54E7uaeVBJFnTltsL8nExK6d4kbMwF1z9OV33CV8uspOOPpRmnhD
AixNtQiaMXrg6gtGx7NWK6gAfI1F1fLK9kPmt+aw1G/h/l11UEwca08u1LRuLHjq
LODZ4cDmjYxSxFqNOUFUCRD86ZwCWDERq4wndIg6mPVFNBpJEcc01LQvsoi7PQxS
UNxMrS00A+XHlP9sRNJcOXKtxEp3bx3DjZ7hyaKvD9dT11Ls47rn/pfBz8i03bGR
uQCp7UEU7jqvg5vzpxDfplmrZ5AUloYDDzqny0awIEzz477feUVV9BMBW9DlPkGt
u8SNpC2kmtPsqnchObOg+t1p+eSr7F+ilA8ipNPNh6vLC/HzKg8Jv8MJWo+Eq9r3
U9W5lqeJ4zbTbMx8w0/RZD3yisADJ47GZKqhtkQzRG7JRRi26SncUIWUfi7uOHkb
Evt6fgtaK58bWhVL8MeqMZj4h9k7RgEl9/aaK2En6W2Xgbrm8qyFTvV7T55QM9Fy
Fl5ohbKJsudfAfGNc2wCHuJSNKFb4HZ5ZvTWP4Tiw8+JS893mAgm46GaeMiaTUqy
K8Ix8Bme23MVwVHREPlczWwo4RvLItQo0GwhpDIFgyl5kDrauePK26ZLprGsIqIO
sM/RVJbiExX8GEZw7x6Y6X/z9f8n/sTe4l/HlsGP6O2B1Zwt//nSsq+7gdXFsz5i
525oW30e850d0Sde8EtILQNQ3ASbi6o4PV5JKGWBd4jPudoEVj/9E0XboanDD1Y5
+pknF6BUqKvop2VXRhjSLDaK/WxdG6wkj1bhpMoAPPfJeMiviM3vQZmq2IsUSgnU
AxPk2NUYlxY/vDng/UgJYfewxkzW2Qyfiq+CS2xGI+1ZVcoWnGydb2303SfEEd+w
mvhpt7Au6ALIKT8xskxx91Sxt59TVVXy91Fpsx7b3DEQEvG4eNr7XvbbBcTuqYtR
lfjTc+7nkzroxsGPcsIBMZ5KRKPSN6lOpkUUHtD8ne1huces7ZvL/WBds0ct8PWE
8BglA20HsjU22it8iDtEfTyNxTVcUiZ+libApWli1sdwKJ4gRD19r5pFNFK7tnHu
njTsNQGC2rDHYs07khm2FB5B5JLG3aw6mtwuWBQa2KXoW/wqcK2WhEQtsL8z4GgJ
hIeOd/vfEz4jecnRRY+0U+8mBIjCPf/XR3bkxrHam8QBHIGk73eHhatPpskisHPY
CPcM6JJ+NDSEo69OVwbaLrptmngsvyD8BVQAJmQQRJ6ecDSux2GXHT+QoX3EXeh1
mOuAdPZNVB8IFRcvMMj56WzwvthRXTmE2u+TFEF068NmPgOxeH4tlAMrSdAlbRTj
YVJNWxAo8erslDAwog2Dxs5gJIbYJZIX26pM14hYb3uwxRydZa7CNAJyC6kfDLKc
aJl2By7hsDlp6XVJ6Ez8BK6JyWAvLdtCCdr6cnDbZ/VJbTG6yf/kGbMuxho6riQC
QIhmpWi/BeHyvLoLCycg4QmP4t6nFANRRQyBW3Z9375lXcbw9F94DWMzt74zwr3i
vcpzgo0J76C+Au9ED4XxBOM9UZKkUF5wtzkp2S8gFjGRNs/PKxjrruJkv6I7dCnq
AfF5XFGwwuD+2pGhj4Xaw9vdJ4NP76Jz6AUu6iL9Hb0A9FB1DYjEnbWlrnKod3nZ
Vdw6UXorRFsEaD7SrAiYxaR3/ZImObISeRJXOka12nlVoM4CkQ7diGJn2GF+uJmZ
zXDZYsi3++AvzBJ/1yf/LHEjseTYLERL0P7XcGp3Cb7mjTR2tpQ20IvIlH+jn6Sk
8Gtz0oDbqxR46G6MLlbkoOlg7LuhU7vke4v3VK9ySeYHt530NObxNeTstbwlzbxW
Q58bGv1hSk9tahMX+ImpbSzwBQj038RdI7plCK7A99jHBBwm5i218I/qDEfGj00s
r39F0m1E80s2P/kc10p0WOVMWqnxw9krY1qQN2eETW6EakfUurK5VD82k7VREpvY
wpnM0e1y061JPscHKBR4UpwasZ7Xqk2DEE2EkaHbQcBo6yxP5u6P2vyJmtko82qy
009fbN3GRqFuQn50ukW8wCQ07Nt1/wpbCV6dzdtDA/B24ef/5/nnu6v9qWoYJsWd
Fzh/JFZtSUWP7HINnsAw4lXrgVWh9yj0LVxz2XfTCxwWLH8nOhinLJU1q4GD6zC9
A6q8YVufyocqbFw5PZ0IxyItZQisTCWafHRo1lc2UJX8FcfB8L6VzcluyqrEOi6B
qTlPcVP73zuxDaCZcm2fgYwRwxAbKFlemyoEsZ46GRw20o5s1fAvlltN7BKqiyUx
GSmbxifzn4J9hlyQQXVccv+I2avsxtYbWsFmDYyt3lr9HDM26wlC5+wjaJb3wDq1
LfyHfmDnef/GeeLaNRCCX+XXFWGR0DI1kBKC2xK5Wz91XFG44nGinrtq8gb/DitZ
BbUCtpQ23uw7WM47LJDF/8kAqiBvXu33TPSKS8fRbfuwaSt7Sotno5ZKhM7oCMR2
uO89nK3ug9cO4Rt6039bmcjwj2LJCxqoSUXW/VuRgBi/ml/7Pqr1t3jn+8qmHUzL
N6VbMWPGqDro2VgXqD+lTJ4euyLEMBSLlYQUVuwetk/bLtpyFEedsabeQweRjYxJ
1YzBRahS8UbTQG7+b3eMptjESqmNfa2/bbwScxhdgqtGy/aa/AfqOWAqRgs663FS
XWLLj1nbLL9S5qaJo2laA5a3jXm1ZBHYEBEsVwEoyw0OUermc/gD/hYcgFdf5ZGr
Rxp91olXhjmXK0W4DcNzJJ4OUodZpmfaz0NPcBSWnmzywTH7SXC1V8BAPHGal8ef
shAmK0tkYQkEXFn+nu5PLYSbeL5FxEmR/kIpelRaO3fo/cI9FrlschiJTzllB27S
TYciNQikV0Z90r7roVD4LRibnm8HFyaNDBZl2HTuV4EGYFg3yXQ92qi0lap5z22U
RJU8mTG3MOupxjfQEwEIr7utwOe/W1nyNoEzsJmVpC/8rYHNw5zLLwKamvtXsC27
zYadQNGbKUkiCSoQhBPltDMUpxek0+U6rsQFWhgXQpuf94qI+r08N1FxXmzwS9kL
TkrV5tt9hQTdkUR/pXsaJY06Imc4YGMHks0OY4xgPtStlYpHWIeR8Gs3CogXLgbJ
a8Uz2s4BHSg2RidEkKJrc8f4SFsh2YX+Jb8CqaljsEh3BEkHCNy3YkEZsLS6reIa
53UxSihNF2rlfHv4tsvDsHLuYorZ17/NZRFpToGqk5PjYFp6lpZpTiau/sag4sVZ
8+kGvQXzb/4H8ACK+LFxWo8+iDZ4rNZZ+ZwlBG/21DnOVDZvHVss0G4Dp6lpc+ZD
KL9OxRdbQFsdulh6kFKezuIND8P7VSNXOWc6CCmAkD1E6KjOofqhnBv1JiOJnd6x
y2mOaBCLMN263/R3iMRzD3GwTpIG8+ixLG42Kq/Ud2QpFpjr9vcz4uNnRbBPHqWt
VaHP0BcEdxTBm6jhRlQ3YXSea6y2OIj1aDcxOJK2FMcTw3IjvtmXOyTTRS1Bbemz
eP0Zp8aMc7C3joHbEGOiFHuXcLafT9c2+v9wIw5+B3cXxc3AHjnQ5aoXWxtZTlrr
rscKSuqEcpTLHkjfH4Rev7qhW3w0ly042ljkfl1HqjUMrLNJrJ7iIlIxddP+Od/t
UNAl7BlQvpJyOpOnyukTxtfxgT2Hj6nVQZG8nQCY4ChfLmACpPVoP+YIJroBkduo
5M0YzNhU8wgdiOWAtjK799kXQLAuoECRdL7Ft24eisXKnwjmRorlFlmgS3/u9k7G
J1NBS80JWjAqmNrz9ech1PtkA5Cc1Q77ixcqJHqGPUBzAaKWHA/4tWPw+7KakGwT
DT5eHApgOwySZpjjPK8E9HMiSO09w2WKR6dViukING7sbRjVYiBfqFrMNxEMaR+X
7BYcCggrBgpg5h6CcJuF7bg7CabLom1QCfUQyyhC09C0FnNF6UsHu0OD84sPYzmY
edmTE/khAp2cbUim4S0UaQlqnkn8b1IuguEeDll+jn1YN/MvITYrJq6om8TnPJmk
YPm2l7q9kOylAFupeFOKIa4QwWuqTW9SOR+HOvKka7AVKMtQ9s6YP2DC3+yZyv/O
JiqtMiWn3GwIv1UbLmZ8qTGGVCm5xZxAT+Ava1mTIqykJjZIv7DGCnKr5xjp5mwL
Ao1NBPlEfDPdVGoStOerWwVkTtevYqgMBbrLtJVAvpVT317BQQcnU15Tes5auXHE
PKwICq8fIFItQQfCZOWykHmG7NDwcCjKbcEwI+6nifNaHwoW5BdGBQ7ibYw6OQzo
YtvJfY6zBSUXWgAU+tZeT4OZrkXmPnFRyacxFhU0YW83eE/MjGQtyPashUDeGC+P
Ynk9x1JiHzNrSfcznPDqQc3lsLtxkwIyuZMRKsbCpRuMysJXXsL1AqaJGKtLstA+
Y68RQP1SJHA77tmxyZL5030z2kXm7lVmsU4zJWRavOE/5RwA9yMSEuMKUs3rYIDq
u+n6YGnF9uhRdybfMIzinfVQdUgl47K2t5eimL7DeYi3Bg4OWk/7IvDu7E/xHrNk
+HD45GfKNo4OG5RvSY5mNZ0A/KHF7d8UhinOovYReRS5Hh6w0ygl8YJCfMo6PtK6
P3kiIf400welAL7NZRKe08YeLH3f1ZOYUS04NO2WSJK5OkFHc2J6WG3B9Nn5nCMZ
5+Z2BwaGCH8m9G1icE3vLiAuK/iQMUAHBI/WIRDSHrv6H6AwB6M3r7NKgTikvG0M
liKZlD77o4Q2tOrvzpH5kGxT0nwHXDBnrh3AmgW9q2h47m4ErLitMevJd+JlFp9j
mS1t9YqzdXsUNleqyMoJHmCIQctdwTXCKIoCuWDTy62/gqneppZKIb3n7Iph+POa
Oc3i4sDiQvDKyNPPprxS5WRrm/4jCiY3lO4SoFSmMm2DWAqptDUA7v2uPqcteYEY
n4qPR2l8LkHNDnxs0wHoIg9YjzQZ6X2Oqy2LHGplemP5rqGwxlDEiwK+AtCIZu3I
ZFDSwY5NTL650QR8VvITaR0BkN25cLH66QzLQ5gfQ9GuqWxmiaj4EoZqs8/DutaB
n6XEpfgP/o9KB19tMXM1teCZmU7zvqxZjfAsgTMAwXc7eKb02uhJGtj/+jXO/emi
G52FbuHuxqMHcHkkxIG3qrlJmT7lhtGfTedikw+gUr37Kgsyn3F9LGtSGB13qEi3
Uj1MRdwre5nkXrZ0TyFNi2KBAjZShpgXuHnTy5F4iwA9AAV3YCUhnN7O88LnIOHg
+edew+0kbiYRnzNRTZyj6f+EpEhQN+PzSaZJMET42vUKhO/DQHhZXZxkRRN85S1A
ClL80ypo95waYXCC0ChceXg6mcvSaoAMPDR2kb9ZXhsylCpItJ5cNAzC3h4OLwve
hPZYW0REWIojrfK8VoQo3RbfR3mxzViZ3ghGhCxzb8BI+GP/i+kQY9AvGZlJfM3F
3+1jDpSrsjjxFEdGX/9MQnCm6vLx92V/JgPS/6cRRAltZskHF1nWCy/P6cHSSwB0
lk1td8Y+2vXhMmMCf+KED1Xu1scPpX5Y/yh8R/bqFyPxbJhXgea3uF2hXrxRSLks
hiUvPpJ/TkNBCsy4o/2EDwuyqHYSKyIhYJ7vSxFXYigCty4Xm9tzxNq/9+ankwYe
MSbmA+kislDS0fj1Q7xO1TzJJSVHI6UYHyTqOlqGFEKRM9EKd99JWwwMBo6YzFC4
bbe1t7dSpivSGq7zOQ+wzF+YZy22YpmuO3naQjYMixPJvSt4oK10QmKKdnO1gmWO
LAm3ohh8EDbvOyvrKr2M9HfV1ZIX1rux5+OJ6cuex6EYHzI3ArQVvTyaIHA/3iEo
JIr2OzS3NoxM3rEDg9Q7dqvFdTm/QhTyFZNR+rhTBXT7VeTusY7C9HcY3koCc+dt
IhWSg8zpc5e8D+/O8mmDTagR99fInjQHFIxK/67NeH6oi6+0k8PnTBPHf9i0Yp3a
tn73bWBq3bTicKeIULDhRKnUQrpvahGLodeliENI+zrNDqIPmr3a0JQ/Nar5dgps
bEFW0e5h0x2o2xn0nTLa/18XpHFysmKpAhJNB7DV3kVlLA6ahGnH0ngaoycDa8GS
JuLbn+DbiTEh9yB1eQpUP2ZgRSd9Sp71Xirqs4PuSHLHIL3R2bwJaLGGbUQGFFpq
TBmMLMAHW6mOtl61YYXwTG/yHCLSm1NFA1Fp3tkizXNYr2Oyk/Zhdtd7liTxBZdg
Tj6v73ra8ZgrBrZ6mL+4WeOcEEMUP0MC2g0Gbpn/NUAq3QGv7qE4S0eNIqBKWFF1
N/L3kGLweDHhq38cLLLQ5hjc5cWqedTXqfVchEk7+V44LUZFlDnsRQ5ZRJ5O7sVR
e4pe5fRvXyKgj2MhbWBOaC/nD2as1QYvRbTq5kO4UZRCSZhXCw4WLQV6TvFTOzmw
CHcJx62uCGHvAoGJELCtPwfgMLKDSvJTMJcNMGU1TbvZIuvNdZxJ/Dmg9j89iUKq
xZCpzyX0LBzdsMhK0NSR/jo6nKd127c11DNFx0uP400ZKsZlZnvd6ITJgc2VU2X7
7XP8nKghll1wbbmWxnwmYkTssltnmaBNHhMcvmv3EILx6XbeHaOexf0zFfYADPfj
uq9nSxuVM573dyN5jTEump+17d9vC/JUTWmQ1lglLxAoseu/xvjeH1J2IVpR7kan
4K8WMkaIuUMTJ5waBcxUQs+kUjQhZfc7DLvD+r+KS9XF7uY0bOrNuHAfz/pq8uF9
7LVZLoIbspOKEqTKV5zDko9H5K5kIClMAddpTVhd9xoUpCmpj2bJcVrd6vEuAFTA
UmN2KwnXkOg6QQitkp+Ytte1dzfr7+vfY7UKAyEYtV6pOo3niKksygAvN/9eV0gi
YRR2FTLegVW2lc4rAuU1Hek1NF9vR2je9h1MtL1huce1zRNNhbka9tu6yzHeK719
peuRDxXqaBGo3bEhvCqPJuuNiFqp/9v2EFOImOlqhNRXSO78/YR/Z3w+Oq7AZiZX
yWST7jUjTBEQP9EXdBDD4YyZZDeMsHzFDTWn3APYzYvZXcrdK3YCmLWN7sJ1NBJL
CDFiGGwJfmvpRLbLzDrJsQrPWBQ5FT1Lf5hz9dMKPV6BNbIV7Za4fDW4JMElK546
+qjpx24MkqNESmMmNb+/s6ecHhCWUcLjKPK74W5lbJ6aLAiTz2pU1M460qZ8/rt7
2+/ILuYboQNLlj0L5QikovdYB+M8MIJ84eQNdzRl4/HnJriNe5sjyupbbdw1k6QL
+vzHhVxG1iwBpxRBopIlnaPDE1V1nuJ++kfQ8RcBSidOnaRFbVcaZHQ0PFqqEBtr
YBOWZl1tfeHYo/y2lhT9B0VWGC/qjP2jWnDnQpJ7qdwNAZfbqm9wlVvGaeXrc3ZC
EFNUoG/yyj0hPDnsg1Z5dGl2LuVJMesEPRyFbXaRnNEOvfyJLNjGtZXxYsC7leLC
w+a9P2VTRZDUVf7f++4ys4th0EbQG4nIc/2MNtxojsuw4BdxG88MQo/FPGcaumHQ
NtNjzzlp+UqNsrdZHDlEw7/Z8A5gXrF0T3V4Pr94VKK5XjQiWTKVW0XyPGoP94Ej
/MzE4NahqXSpOjKI5Y46yiyOkLg5eaaPsgLOUVGDjqLYlDH4Mdqoo03HAl1dfeOP
RGKqyU+K/sFKXZKyieyMXpx8X+ho2M9RKsIfAqmABtrz7NDXCYiQmx9cMJs02B5y
Y0kdQZkeI1cPVTaifS+MG2tWy9Fgad0LmWXTJ4CbALzTzzkENYnBruCIyUBu0oq8
icg+G82pAYAuFcz7yrAI1+rkk/HzxbG9vOKgSrLRIAuS2w2POWfRReVGcSvFPnwK
HLyFvvUIDEjR9K+nJSs5JXDle0VjvZ2yyLEHUBcl3AZRbs/bMCStciHK8Irou6JH
oGU1e1Qdze8lPuSuYqXZ7osjNjY2LDtZIlBjYX1c9v4GmLgUrz0Fj97qczDGb0Io
7H0+xihTY1DxvhlUztn6VBUv/RJKRpP5YKp/A0sFvToewu3ZYiDg4NAmEHCcIFH7
aJGFk2pSRhpXDKpCODDtt2YtGBUyyulO+/Omqsn9dmiXBfiR6wguuOMkM3SAsgsp
aYSoTq60ARHHR9GrIIwwSXItuUbS2RBjBQtoe+RktGFQ+2L28CTO6JclN0z/jgrL
AEu2PvrUF2dLMSlhYGBkEXV+X4x29eXxsYtNhsR9MvgvbHsmy6SUe01BiK2xe0c2
dKFEnlpp280wrtcy4awGAbMY7N3GPwePuoZSoKBb3xex1wfIhesA7lTdplFjAxAh
SLt7nWBgkxMgkmznrnYeQv9dXf3jLI4IkO4bJ/8crTO4JJNB6efN1fPRdI58evwl
CUJor0zA2lntEYXjpMys2/g0ZAMM/Sfbwe1Oc7hpgiJWPPLLB1qvJU9Rvle9U6lo
itq9VRt4tyyB2gFekHOddWrP9qCHeXBHrbnMz5TcLfi26QZZQM7hvDcBh1EfPfbl
rdn+jOI8z/HvuqT+f2+xeOxbu/qkUfBTBkCTvZSSD6BaJn0ZHNAwgLD9DoltUD7W
i6fJJXmYsbu1JdkjEwhrey63axCCPq6Xri2bsO4b5kH+AE18nf/AxEk9vpbJWG8K
lNTf0fe3UfNKmIE4ek7WrsRMBpOyRlM74PW41RG/bBwroau/37wV0n4k31E66Jag
EPkn5Rx0dxqRwXBfqONyVRdI4Zv96srN4hzwh9T1Vqkq97Do6MQQhM2fkw9PM864
Uo/eCBNCk2zYxBqSsUiSurGq5b+nF9NQvPB5rbCNrMuFfpRKHGmZmf8gyNVWNjMm
+m60vVvpXjND9k7NEdmqABdk5HrTEYSRytkaAoej6uYCQEdv/tYahWTBVQsyh1EW
FB7mOozvN5MLmoWOmWzdmVRFfr9jOQ3L2RLqFa9m5yfwnMso4cOQz7jX55KCi8+/
lH68Ca0geolqVXAEaW2fTkukkmHF+XTdBBiRmaMH0ehV3HWoKMoi96Prumea1YZe
Z8ZMz7f9t1pGwEySZcIeJLx0Jqf5M/BV0PZdgeEvKFuXfn+5nxe0n0UNjMfrZa1S
2Yu7yOX7xnyRAfAuFLiocZDuilZmpwzDg1zUxECVBAtwfhh0+yDg+HgY3BIg0NhB
oR4Vw3uGt90eCxEI7QJU9NqN63L6gXlPF03mwZHvi+udrqXDccNOvrQuf7MNcRga
zoLWgUhQDKyJH/JMjmByQT4iICpzSpCZs2GjoJasz5+2y3wIDq+Ts/sEUBaiIn19
6uOuUGUKfsTcoI82X8pubXqfGa+sa5xnzr9oWnPhJTs3vNKNCa946kiBtk4dxsKQ
+rmcD+0nx5KAuw0Wn8SMcfuYzCX/eNkv1S6LKzTpYUL6BaXx7BxGn4na9rpD/pE4
xjZc/Y28kKZAu4CRc6Fmtdo+W479/x5EeXRkD2aqoICmsWZ2wOuuF4TtOYVr9hA2
mJ2EjldLhqqDm62+CNJwUFjFG30Edpt5S9OB69qvMHHo8BPZs9EBUCDS7WklDw3V
hn4j8i2a8qDNHas20gQZh38Y+Enxw4SfP0hzYRl+A9lZ6odCI7PNi9hl0R3t03bK
Em+czMqYf+UxiLB1koOPymlnf4uruhVTsPH0zuR0NZ+o2q6gIF917N/sfKD9Z6Qe
KPwgOXlDHT+FCl57T9Da4HJEX7PMpKLsmodIUUdVB1xOAHroifbaoIZK9GXmFaeJ
w9l1bZRu+vZPaxIocqWSfVmIJra3fKCllRfh20X1nnQ50FL18UZxZU0+yxGHh3Cr
OLH0rIja00Cslp9N8s5IsaqDtbwG8EUw0a5U0jM3YiSX8hSxZslh55RMjqJlPwAo
t81QxAyqd6N6gZQ0M0SPxKowZ2KMJAt6BgmEK+7JVfToxoGN/lIa8BRbd2WJnpXu
Itz/5N1VLbQJtJYbv68rGpvFrV8O9DsijLnxFhWeBDYSMOmb7HRCErdKFOMyI1kw
0KlPOHnOUYjXsT8vT2ZBIic8bhHBcAzdkseqhFNJKoVoRtoNyuIs0larOVCoD8UN
TVFxvEyUbIU9ZQxNUa1pc073l6kigZeWSB4rQUtpbJL4aVHMlXKRDtGlUi9liz8B
M7FkTClNdArbQxajPanTSDXTwWPGcq6C6QuBk0fD9iA7gPzpC5mmWCN9LwxAnt5y
oHIlyuMiycjQfTVVnsfh6vctZ/3ICpjQj2MaZUjJKmVPARDkp+wG+dEZMQvgOzRr
NPLXwvkjnGhXiXmvKogjSrt5fa0Ub1wmHWTKncWyAFyA/FmIDEWWJ7Qqq451s+HD
EKCERbAu4q4PFzjEaC/gkeP2R+n8lXCU2uL2Oc3w0iWRed29UkY2UnhyS0MMPwk2
xxQjnVkOpwW2MQwLHelY4A3MYq11I8LAbDz+ekuZoCO44v5knbeLzd8LTDQJozxg
Bp1IkXoEthmfVok0zAg0h43MTnFBNPIjFr/cNVOEssZe6zatEWSkue9GwZ393o6D
QwCeDHQOAMwjA6IGL7FkhbpK+hdVbNhDb0DzM57hMNnWx25sidbv9OVKXER1m9GL
FeCM/Uio/qv4YKAFiVptCkFeD43MRSLFVeCacGhy++RrUfb2s71VezMhKgOyt+j+
aSJA8ZH6TXROWBUFV1N4AUL980J4nYYQ/p4kxYPpxOmjeE43qmaKOovLaAoFTMuh
puPnePPxXEWG0K2oAQQhur6Fq7uwPdQliy4DEf6GFa97rndNFqxmG8iVl6PidwkX
aiDV30tQkqFm8navdGWrWcDUWCSzSCDClTT5reMzU1DMHrObXS6/HhiCojmcIcTU
NioQlI96YAvRYbfd30bFV67fm1qFBfGBhB/YyYbywIIqAZ2jWrQHJO8njXoxDivn
zdW1JFFnP+7gLO/wLSBNcwBL3Tfzr4/KiMoy5Vr0qZ6jPDhGywB+rGQBX0WbqwS6
TVtxl6PzuWj9/TEr/jNBcYnIEhbME+hLC6/XsD8IESiSSfgPzk4n0zjzTqOKkVcW
RdyqHhWKRK7ndSs6IJd/gImwgMYnrhqvZRMQX2N4jDvRFxOBY8BtUb039fi4RFuM
CrUp4yMbmCKTE9golGSNL6u2IMWyDs5UnYMMkXLE5CDK4H2N1u/Fpe7YCCkA80ty
ZN4d5lRrhkpKaW+1cSOlz34oRCEPWib878/FsNkmHNJFajYYFaCCjDidtnxA0zHa
rTgC2QgGXOoWWLOBY933ut46FINB3xJ3VYyNSgjm+z2+KTcp7xIFCiT0ZrT8DH9x
ou791SMCrPlYKw/6DdqPqE50t934bVQIFvV2jo5t+nu5ffznOoMd75czusLco6Mc
UAUQQeJq700bw1Jg/w0lzJO6OtldtkQFSGCQ6NI9c6d5FaME8N260vKJFZBkHKoe
DF1rAUXYHF+ABAKWlqacKVZrmNz/7PxeQezVxZ9Dlc47DxmWk2WN1gFz0qmDer+E
0tcX1MVBp1972XIvpiZsgTmvzFgrBWbBLOszzVozMAxL98FP1BJStySTnb76pnOy
+s50YvJVXJ7SKzMcGhRHaxoxCG7b5WvUFACR5oTWyQGM7BKQhAEcZEaHwHrTXMXU
nGTyOjbZb1K674XVKMuzoqt74gqPEBEncpTK/pOVls4KgNEW9eWAMloqRhG4mezB
lGysx+zl4j7Vymnxg01+PY8CV6KCn+6H0Mzm4OF0Rndcw7O0d2DFT05LOa3o4n3y
rR11ADJIjn/96jGxYwJmGXt1+1s6h5yX1BHOmwfPwsQbb2Sy6RdRlj0ayj86cOdu
MP83vdlb4TeztEllWYlYr9XqYdcbTLuxHb7PI17k7CvT5uX91X9RHlrcgR4JZG0X
KA2JPjB72eAXNlJVJQOOEiSsbmuaieVNnU4Vu76MudmQ1j9zJilMHFOynT1nqyWg
9VRb5IShlj2x6JPTqjApbaJ8pr2BVzcpucGYr2vJfgZ2EVe4zjQkuxRfi1jdM8Fj
dXX3vRX5+cTx98/2LTUzKt3ToY+crbVRhJqjxpmp/7jJrk4qloEjUVUuhxdjX9SV
icH8Zh/dSa0vELHg9ZJ/URtgC1l/Lnin1xMxUVBwZ2nxvHNw1pIlBVm1tC8ixabE
1cwJdi+gc/wLz/63vizj3pkvtXM+gWUSbjU+NofIXNtUZ7LmSEKK2hnnZq7KvpQ5
+Fh/mLLh+HeWx62u+OZvCjLm8bCO3+XPZdx3DI15MTw24/iu0OeEyBBXQAO9Dw1T
iL1tC8cv7cl0cwegEZAAAGiLb3E0qWNW0qWFrJeocwMijXm8TCt/Nqv4FF6oXmbU
FPijiz3rWQA47q4YrJkd39KMjOqtbpt2P8Y8VdwvyJCcLyg2FH2IpAJ+4uU0hEl3
C5eMGygspgrqqGZID12/9tmY1giUCHv8zlQAgjb9Q5VgncFatyrbM23gt9yDe9Kp
PU3ltP2XUDLcUCVKmCXZpF0RZ14dmNLbWsYQw7FUUBXKslhyif9bTDBB7+zQcYfT
NUO38Dd0mY8acCfsovsitKNlUKNnvhileL0bPdbG57KlOMS7u/zImg8j7Q6Qi69a
XO04KyyE7Pd2kmCC8XMrZ+fo+O+Td1ONjbdXTia7nz83oFBCiU2X9Cufay7qX6DX
H3j8cCgVzR4dapO5BLu6c44X7LEGmCz0R8+STvswB2JqEGc08E63LpAoq84y2e8T
idKySSci16zMOEtDEwY5gx5Tw5rof5o6uXo1TsV7taL4IkU3jaR6kw1Y5ioJxZzC
sXrhU2myr4A3Hz56PblEZkyP5WNmyR/aBcbUhE0ReWccWh5MSGG2ZW7dlJbEDvU/
8IJQxOIriLjyhyQK1iSzKfsgD7yZdEa2ymiTLiHkUcthU/d8acHcjJECQrt6ESzW
/quO46URn+VjJQnRMOGpc0ZPMvQNAc2NdVGU9wkukDsT1aynt6sQ7mfM3QxVoXdg
w0qJpeZnrWJD5QNXVTJtR//qRiXxItRIPeZihVDDm7zogSbpMDMOdfbHbbIfu/vP
wCkxiTsHY5/ITFN8/0hDCOiwoJ2hCMJmvIivmtVpIt8ttZyX+VfxhhslpArjVef0
OJbez73gJxa51lyVL1OkzwmY0XB+gi/R0kZvNWuw6mNYm4d4FOVU/i5EZkcYaPLA
/RqKS0YoCsKg6ml9E9lNTmicN/qGvIjQ1BNM8KF01JJZNe4SXSNhRcrAw4WD5aim
K+Fp+QxwH4UXsWIYjy2MTXwhY8TnpeIgfUh3NmZmLpzDOlaFuFBThQWercqBKoHc
gVZr+dxMPqe8a5S21lnd8xT/HA4/cntnQEIPuVS7xMXpyEC2BZZQEICdLiNWE3bo
3wdK2nfhXa+0aSZEqnMnEawvXExwfKH2S7uCBcdXYvdLJRiMrZjwI3Io7esD9iMG
p4TA91kMe7Jn0+jAvDrMnV8bVhdQGU/9ruwDK1wUV2HDM/VrQyxBJoJJ/jPKZwKX
zKbA6a9Od2qeAtbxAwsfcwjz57YZWJG4h0R71tUHCSEUx285s4cQ5sEAUsNiT+c/
jugbUO8l89sUmL6VH8jpNSVDI/EqgqqONarLtrK+7C1Cke3194WRxTSlDO/Oa5X+
FAXWgyyjTF49otrPxNcqD1jSCWnHWDa6tPUGpX7LINlTu/8BI8Dz6qFFh5yukwVI
WrQCu+KNT9I/7iceqtNYZ4yfWPUpZxDuPx9eCUknRmdG2ToKkLUkvVpNEmQ4O68B
PNwUzJka29pnkYX+10b4pI9EFL1TqsqXnznJ/n5OYks/rT8E+EnAVaPrk2x0J6Xv
H6BpEPxBaaJJGjp9RiveJpWR4eV2NsGrx77WvC1/G8QtDKRcX7A6RahbodohBQmH
RBGOYhoxki95OVqhFd6t5Ho1m6fQN4ShL+3fmDDzQp3578Pp3auUl4FPbk8CYZU4
xZ3kiTSLstOCx/9Reiu28a0X13U+FFnOA0At/swuPuAs9XYURCZRivKXDXSbS0KF
lB+1voogbW+ZLVkF27mBLtJjvjQpxOCyE9LjAK4X6f2TEs2ybYRqefMKAYKjamSW
M/rvL7xlXXU2habPZbTyXUtW2du+T1cz+wXi/RW4HTIzRrmp4RfUdsTdwWunboa5
xaCHt3Wc5M8UmnLyh7RS8Q70/oBDBJvrB5YkLWi/xzZqeZAdzf+hFkDMdYLXgV9y
pmFg2r2dGBx8EERk0MA8xKfiN/Jv9vxuC5rr1PkGMtaSTZrKV/W2t52zEE2USGDv
ua4W8cOlCPL5nss8fchdX0+sucYHRptQEg4Sc3MhgDzSDgyR5cctXc3TM50ju1ae
D7eYTgklLpdaAZbT3nFP4nmQSI7Q4JtspfIGyJF+SQv62boyUT7jX3Z+bI+enImX
H3jy/CP/mtTpJbPtGaLndw/cp0hKRc+JKI+GA0mmXIUM1uJc2jbDM7ThdIkbN9bj
oVO9sBVXJFFN1ZQDF6RtDR6FzFsJegkHfRI8+X0CLgz3r4HEHdp+dLjM3QL4rgbv
V+wiCWoWk2Aw5HVB5PvZXQJaOXUXMU9vprCBlMkfIyJCZPr3iheWdJC3Za5papBj
lnPVMsNA5Db39+ZdH7pXY2zIN8n097vBEO7RI/tgqKLxfkTw0AyRVwOEG8tCM+V1
cxQRlyfPK586zXrHTuWj6LhV+kdJdaqEAAPePMLQchEumFD7TllZfLunnSHBHTb+
iVRYlM8+T4Q9fPs8/rZtT08FUBn+Xa88rJw//9KRggxkcJDFn+wu3OA6gJHj5l1o
NqWHMb5cqy+VXkBYFNMfwgcaa34QxOFBx6VBSM2ketuCaR8qyRx7wXAYGz2AC47j
I/hgXdrbo6xiNUbPT+jymDIawLFXFleae8L5/bHT+34Xyk1waCNhGPJ4ujGAQrQy
av2bFd8lV1cAbZV6dWAjod9ZQqvxSw0LqxNT3RVhTWP117z9Zb1J0ox9+NDBigBM
B7xjbY8+duomCB21Jmf+WR7LvJjSjLD6TyPpO8fDivxzeYQ1wrCLSYCW+oWw86aZ
ZRANYDS1l90+WjAFWdaQJCA+GYwGTAAWck9ioIr2o0Z7RfBKc3zazhH+m/yvIBaZ
7zJJ+oDfq8BE9qRcBgquyXWLDQAQLx/9dKSJctgfdowkFd0c8DllYaDZ7tMxAA0w
30x1iQ/hvKsfVwxIbA3VPXZHyOMXUQTz6aHzxvFcWhFXLm2x2V9dcpIgSS3b/lDH
PPHMAfOgOdWtRMdZyvvdCc/ll7c2ez1n4VD3eYuPNN6frDpGj5Mxd04nGgEcYh+7
IYYil/ETqqmH9oa2kToLSLdqqQ/3jMWvyY1ffbyFRwtBeNlvB9VdqVSeKcaS3WGz
ErPofJarP5kKV8sSUCJxGI8KJwZnror+Ga5BrcbZYKWcWChRvPZ7H7laJO1x03tv
SMeJtUYGRdeFbh02nLAhSSDsGp/Y5IZwhRYEJDNW09xeWoAoUTd8uouRJL1YrRoh
uXzNNrMADYsgCzxVqBXkKgQ6vuJBZUdRm/1mp3/sgYeg9TNQ3MrB+VtGw5z/wBiN
A5KNeeZ94Z6p3/078iId+PIqbnKmytaH4m02A7i18+m1umIWJw15/CbZbLVH3FKd
O+VlvwoL2kCW/yf/8nmWgo6EDY6qyp1QeHUe2n1WFu2RVsh8K499N9ro5KEOqgDf
P2qA/Gfx2m9lHGqTMi6rgSje5tMXQTl47AhChUwNd5VUH+NCEmRz5qi9coyNAAtb
Jn0Oke1HZwFVJy53RefEsR4RCTNUhHQV9b1acHozh/Dtxak1wT6367IgF/x6/iEJ
GA7CS89CTBKMbuM2Hc6g6vcQwqFDDqBNXj7UeqyJD8lUw4GpMQIjMo/xaedFgg7s
koLgCB4GYbk/r025g1Nz7JPF7zq0bBX2/Ky++GZE0quQviFmcD6egbsAUnoPUy5a
fCvUy6HyU5ocz6M5CjWPAPhFJ8ysIjOYronR9/j+yP1wzxpAPwPbGCEsJw9VG03l
8ufYzVKexbHkOIvxz2Mx2ilgv39avi69/lfEL+3b5BAcNrddqh92TjlOzUesycfo
BBl5SrOydGYRzKTSO58+w71FH8y3JRegCgkQ0eLzdRgjWKtWF9wcPkhkUzMrwA3J
/w3qHkIjWlY63VWU74a0stDsqyOK0IPw6E4pgEdrmTTvd9U51gtGUESgBXd/dJb4
o5tN2MZkgpwpDlOLSI0vvqN5G4/jv8OZKl9NO9SybYVttkMiDRbVXYvHoqaZBiVp
RS8wo/AaQjHKQhiPvvbhvjUPTfyMZN6IIK+dA2aYu5HmO8wJgwt8W6L14M9OWcTW
ww6zmshqWqslCUNQ1h/RSXB/FUKJ5A+nt6+j4L2tG5ZKCcNmgG9W0t8aSXkpe3BA
5c3Lc7X75zC4dNmRVdUTgrMJjC5XefrztgcUn8ijVR4CoSLMGX7ngGGFYIwd0VtV
blWKv8pgo8IyHFQ5d9bpSBnMx215ZQs0pPJb8H1c4+wgedOUGv+RSIT5aS8f8J3H
MVdBiEOOPsNv5ZBEAGaOpYU+Km+kOpV99J1ebNTZ2dm/tQ7uNWDVHjGcQtDSzk0q
9Bc87WMcCTQzzonCaIMse/3lL+iSkIkfxxW19mHRkVNId9lM1+zr8qluEI4M+B2w
UTOiGmw6Ft/bCPa+VfiZ5ZU9+VlU0EFWeQuzXDBHH6X7cH/mfy20s0tO1kAuccV2
oWe4dliOtuG2RjkiFrTSrM0TWoqjhG8c4fkULm0E/NdZ6PJzzhGLFXyGsdUAYXa/
v6aY2B972QzVvJpbiktpUD95GCdE4w3YwZ20uFW7CeZioGNH187Epc4ao4AdhLEG
RDP/lVuJDrBq5trLhlEDoCO1xQn0V4XFwaGtOrmI+GSV5v8XJD2m6RvQtUd8Sy0g
MgDFcGXoW0uUysxdrc+OnpoZ8eC0n4IDCmbFsckaOT0QzBQtA3S7TW/8yQSELZs3
KMLbB0tp0DYHJS5KNhg6Vho2k3FCWxXbnJ/H66YOM0DLaBOnSA5HWchhxolGuLLq
68n2qnN2mveKJakq6oCdOixZHOLfxAKTS+MkiPTI656/NnqTpTw07wifNaVIE844
uiX130sCYMLC8jVOj57ryxKyGPpmkpOr6MU5KgmBt0FC6TAk0OQmMQuoqFPCIPL3
lOHwh40yZXWyf42yFu6bcLw5e0m4dzzKsxGrk6aZJb5k7DCQBDSYLQ+Rq2/NS1ox
VeIIYDeTswg+lA0Pid0A1HrnIG6XQ7R391ie1ucR0GyKmTW/tft+07yPtYeIfLBP
pgSkiFZ4x/+WQn5wqGvPAQa0Ds2XAAgzqHXB/JxHNKU1EVjKdJ7vJF+JJnKsBN9v
S6F7wMaU9mFHeaxANtO4UuFgaBPfWbFTjvODCfniBFuX0kXph14vxkf6L1ka9hm+
qxIsL12HeghreoBFm09vlEUvL1pVXetjxWEDKFgLgaRK1AHSp8OcrmMsZEdGiNlo
XvXTufz9Fh6JgYyM6Adt6LEUX9FR6zDOPaS7KdTPzNMTXuLAPCZQzWpWwj9X77Jw
Cu2RoXN5sLvGKZI1jPQjIQbRVttE3PbMqYnZg4N4bQMz8MMuNj9sM8XFEAl9m0ue
9UWCEYMt6hby57AUy/JGoqwbGv87IVx5iC+PxA7LpiI5B39nShftx4At3YD8pJiv
cGYNM5A2SRHzNXuDasa5PdjxWETh5DpLGCIVqCgl8/w5TWc+4TYNLEW25LEbFiSM
QLDDH4sDOyQ3LN4165rWPZB8lbOvetmj9yEcQv9TazboacHGvR95XhC5dIpVC+6j
LvaV0SIfHnMUc9M7XVW4+Wf5E18sByQxumOkox9nYCHr0BzPEu5lO8B6zm+l4Bg2
LBwbRQ/Gq6uwn+dx6Du2FlypLWx1JQdKspUXoCYov9UeB93DFQcCS1EJ6e7/0KrA
BMSZih43MACb34garqoAFz5A48wSya7vDBp4FrUKvS9yxyXttRfyjdP3bpCKgGht
JszIHLt57IT4B+8s+LTg4B95A9p8vNS+kGQnMaQ5Idgz3kjUWALGXgcX93oFhkYM
emBq5azfTTNv8shDngoI9T148JhiveEnCNS8Szv7+BKlZkAY1hBJP9IBZ0SECb7p
16gWDJJrN4NUYr9fKNGDu6z2qGLrtcZo5xN92qortQbz3AsKliAkF1IXByTIvB04
J63ISH69ya21SeJFBTxjvR9Li6ALHb+D15g+tRBzlmiQJMErMnjAY2Ay59L8qJI4
R4FLdJ5msPAhIqKXEWrzEbJuTt9zZzEZnr8K9hAUCpvUbcteIk15q+muVQgd0X02
GVaO2HoqdTRnfdBZWOBjOY8wc7LSPb4ZH+EtfwNCHWbEBWDtv7WZmRdnZ+YvQ7XE
C9JsQPKKpp+g16xX1iI5VIjz1sR5WPG57FjvrRihXMUiRXYfb9D4qG0W0C3IGgVi
OGlGdmOKDKJxfjutmNT4tzfaotw3MMm5K8Y4zBXPYrDEhITTOaa0MsKX+7dq5yUY
JVuI7y/M1FRhdYTre+W5XKXqsjjhX2oV9eqBQP33m7vIcSHlUl5unfkZo5Rkz+tD
qpaATvIQgTWN1hKHu5CeoqYEUK7sdt5vzh3vwDLHTe+XW/joJqRM/Ncj+2irMZXs
fEL0RAtY/E65EZuCF6Xa3dnxYOea98JaQT6hAsPQy74IPl0W+nOax7U73SdlmWgn
DqunVZIQolpxgacpDQ42LUYPn83i/6Y8iawClLBzjUEmBIsn3bVlJq00G0uLvWi3
/w9reCKu47OfE/NAM3T3SP4/1QEl8GAN9+DOp1Tt67ciV5KB7jH+cofeBL20JiEg
ybSiZL66N4D8x0HyGUVrrgY86LpSsctDPBSvC8YLpnsFZcxrMZIGVQxtnXYeytiQ
iLjnAYl0BT90aCSSOYrvvyCqALHbREj8KVGiGmxAgEz1m+owYJoKegRoafzHZkt9
yWK1Rh7IrnLQ3HJVrmDJaVWMo7+IrxhBNd7S4qDoouTqYcoXqNJr+xoI/JbaTwv0
JbjdsPtT0VYDreuBDcjiIcKtUSmgXXVCMJlQ1E1eS/llK7EX7wp5+ti4+KFmSr5S
zMDrzIjlTdV0rEjxxUIP/y4OFDLFKFeHoOxyrmsGdaDOo9JpDaGR+uTW7wrxORnC
tzP5R04d8ohes5xhvq81oQX6pBka7D+E14n1nW/i94rg10A3/y/ot0pzYh/t05Xo
+sAnaJu3ueQrjSYZTBX0QbW+y1C2npxF4XfYQVZQcCTzDtct8Zs0M/6lEXjwv6/e
fzh6WyoNn1k+Z/r6GfoKFQvMOaz8C9by9VMkyt1io+7B5OcNyY/2KR1qQdxTGDn+
c/XbIsBbXyOJo4lLrCTphjzZR2PXX/R6k9+/DEZrTTTJ1E9pw+LxkhtjQ7Bx3ND4
6BVqe3r89LwsrMCuDlX3RivEAqwB7XGFbLihb1QZBLRikRo5qTNSQLNmsKIM9IA/
aY7Wfxu+WInOC46HGoSaR+L2Ydg3QqELKu+IsB6RoL/DbBfzlkynihIX9IdCJcZA
+V5Bb56DhYsAPHSD16TeurvPyAU0ZQRybeBkgFubigTzUEMM6s6Bl7FYVABs/+Lv
mxPUgzky7OOdAiqFYisvQvtbyPzwMMhsbf1Bf50FxiAApaBpKgUyi6i6DCyx30uS
d3XaK3k5hMOSP2Nr9Efvza1MzX0o4Wk8rJcBBwbVkUfjUX8pmyma93lDLHmVOIfi
H8fumIMnvg+p7G+pAizePLW5GO4jXA+6RE8m/JBjCyTRUMogD5lt4a4Htm+eBj17
jbcxZmuGlsQuTxTi1LuSpBZId0n4KOftHBX0/ce2iVuGDgPlQutEP5rUlj7itqyi
NqNhUpn3hcRoxklHIuYCEA026DXqU9ekaHfaTKFAhBF35MJWFw5Fg70Ym1YV+fNW
isaNC9EdawUPaSTb0LZvRkfWJN9jWkqVk7ahlWKDzMYCQkTCloEjYhHXlklF7a/H
DkRwuc4UWZBO0aPpnooW072Ffnbxl2Au+XDYCiDG7a7p70x99LeKv13Nr6p05Sz+
eZ6u6NdkaG1BEVIMrDbc7/ukTd5+BXGRd/CgBR3fUWDwGsoBnOv4EXCImREl1YOJ
A+7T9FlG/m2lGtAhR+1OG7moydXsSPsnAkqQ9+9yLZaRkZPoS78kCRSaCDX/m9FJ
b74hiujd9qONTIAR8OIIWZTcJWQx49lt0oH/K1Oo4rp+fc3Z1ZjRgRYxE/xVNCas
HIU85hlYK2AS1HVMI3tXET6e3VJsATEQzcqPcAvxnNQjVdU+8HsCp5BWSfWSfurF
r0p7z6BHdQxh/HgPKQNQubWmiJbSbSw1kPF8/z044Znk7ukYfEiKucbdp2/ACeDk
ETmRRBIj9rXr5BKhEApBkLIQLor0VTHWp/oQF6RrhwFsp8IW/hNtUc0mBRO3pnT+
xp9mKuwBP74NG9wvicdhJ8BJUcjPTm5b06AOI+mT6dDaIjlD9ukLVBWic6TpqDIs
WprEXFoOOnPGtu6O9YnT8RUpCEQzKc5NTMTGgt4nUJ5d7jmr4xijy7J6jknn0fOL
onEb2Nt7uYD7HATX9T/C5Dmu1ywnUkXMwOq5A9vqEGfuLfu4GNIYG/zOiCC+u4+K
N1rimK/pkXKPTThjt89S8oQn7Rd2qEhBObIiIAKjSQXCQ3hQJZ1zvnr1K/Qi3pxQ
53DyOXnAripIWM8JObjBRPKUt8FnqJFyGjn727/fJFSmmEj7E5AufkHjWXfXvLt9
iVX3bOZBWb4E2+EK2UkwBL6akug4gzjkRE6IqQ9DCKSrFu0y9Lr4iWpw1Ylwg/XY
BChII5iTxeJbRNkn8EpAAcdLRhJ6DKHdtn5TX2vq10Ic/PbjhhuTFYKUiszTzaFl
SDUlpTyJCDhanfezlG7gXghp8HwR0dmjvG+xbudU0w71iyAGsf36GWjXSeqcEx+C
q7ig+klOMwPm+G+4weNfl+wH2U6ZHJcAZtqruri3IT60VRx7xp+Qbphc5R452WWK
E3JFu8+G8pioL3Q2KsGaysmNH6r9fGv1bVbNma7lJebfzzwoN7egkYn0Wa0Bhlg/
YRVjcDAS1k73flAPFX4RCYsvRgy0PqYYIstNDbjQvWnklrivdrgdofbrMGkJLsvp
7txg51EzDECgkFxevTokboPLQAWgYc6YWD2iMLEUfUFATqab0n0ZecdLu+lVCq/h
GDoJyKUJApoFu0IP9n55lw0ny3Q/CTqBOzIpy3aTzJ2TPog7f9pQcEvcOFeu7Irg
fO5POUhxbwgZlHRMbc7bLtFEOrj0fMd4ev6zAttq1yJSKF7/6XQyHGCLrbL/TjE+
1PfsXiZ5a9e+vk5ECnkShD7XmBWeDVrQ0N6oYs10kbiZm1+XL86oCoDxPDcTQiQM
+gR65qSEZgLqiy3MYtlGK5MAA4aFidMJwvyyGHIJ80iSPE/DAeUoynH+nN6wSQgf
ZFrKI8kggC0KVH6EuJ4UfqUS+R2ikWq3ykiPjPI300GIZYX2zjEIGdOZOB6hZO5j
o1Kc0IZRQlmhtxUKS5pmFf68kfCtNbfbOysaoe+w76p+gSrskypZv75xojTb7n69
LE3qfgltn6fUhQeNSrRzA1jrkqkaY4xW9Da1x2anDv2JVC4mB7bmrfV2NShBcU0C
9cWQEUJ0ImyhJH+3AGImSSNSdiaRRgGp5I6U8o2dnISQKfufreSp3VkJfeKJf1TV
2xgT3G2Qv2O8vj7BK4gbLbjjBu+uId/fA3JgrdwEjv0jE8MIWhTjfYbtdFFHTzd7
ryW4vEVwOGR0TLiPQ8w7/ik4zNEtgNmLPrb32+Cu7TCzCj+uZh6GuAwjxSWtpagf
dnaBMg4G8eQVlYWynYP/quvK/DA87Ja1BGcns+FAcYo/wyCTlEnKIe9B23N916fI
DxsMv5L4uN6wb1W1Hwp5sG9jHkm9BsCMNW7oe1Uu4uEpK+gKieYDVF4eF0v7zOBd
JiJy5ccGW4lwbmwr2XD/+0hlDFzb4ydhej0ikmMX9DQKChQ8jCngbslkwexfIYbG
3cpYITaCp0B/4malZY67spdM4aWANnXZXTFdJBDfeEmKcKrC3fn/D/3FeNdRCaRY
Lx47cQiigHMnZi8J51h0Bhf07n5rwPaeBoV0H4+PBpO2TJwzMsAYemD1aJ2NYp41
zhqoHI7FZVvv8jo4rmUZjHnJrrXxptFPodh/Hn5I/Y1lxxjOlPeWQUgdzOvQd5rR
9R7aOK0Os+R1zRKzSmX5gFdEpREHirrJbKg9a9eREyzokNwm7oQOom8Oy+lNZpzg
5dhX0UM602MjdaopJaJkqdiaiuBqQYWNY88XqCUJBjGNz4zv2nnr+PbdOfdNF23I
WnWs7/9cSgZLNg7Gq+zdBxdiYrqeiCDGW45PL314rryHabIBp08UXzxbPp8oFzu9
QLUya5q0Tb/6zmjWPOB2eQlssoN5HX9BOeeWG7mCHK0Xzl0aRBCytge3jlTqQRcl
TX2nEPBNwzBMn1IQZ3s/ivfBNWWGkdhvAcFFDVVKt2YYgzjdghVrYnLXYhgoMs59
SWlufTjrp3AbFH/jql6vUK7uadOgRA0oVGoV7lF14GjBvE8vDjvGaxQzCEH0ZbSG
zKpfKvwJjTr1PJR7vOZQXwvhOxefGAqy4oXJtE137l0RmJtbMAecjyAnoqGcmP7p
meXCAud40U7jqZcT/DQEbLnwwDfRZ7RKd7jN9yEQ0RYDl63S3d2GUfj17ZxZbSwm
ZLQ8mh/vxepvjTTsbu5h7/81y05gloN/OXZEczWYvx9irGVfNVAsxAz7psJlLFVs
zeuk9IXYxaxRIZ0C9/f81EXuUlXh65bdCOoKZREhvM8uJwkP4/gYRkKKXY3mPNpB
Ye6740hf0tczgVJa51XCe/PRrAzI9XOKaTw6nqcTHTC+qanC3y0W7rUenKz34Rc5
5nK2ijnsoiJ5wSfGk2C7Ak4fA/QDIgFLa8cvbg4GiH+HsvDQGyxjhhe4OJQ4M73I
BoB3MLK2irx7E4k73dhOYRxMrsyMpdaiB2OTV6RawbENd3ij0iFq2JBIjpThjT0O
RiKwd87IDN7w44bgOM8fe86pItqNa/vjj134Efc2CfMi798fkumMA/AXv3Jw0yM9
kQiWt0pjq9ASA6oidatMKtJop6yz5rJx23PPXcAjMOSni04AoLFb9p+sXF3Ie0k3
AV8OWGd3VdaEhca1pZ3djtN5RPk9n8KVPCnr+K/YB8ZQPvcP/7c7B5l/nlJoatp6
vB8IKB6nLmcaVzwDff1Z8nhyvk7ZGoF96kzdksA93qsnq8AiJjE5eP2vQdFg0xBC
GzrFQ4xW22/5UevZeilpADbMumyUBPbdxW9sr38PqZkpAcmlmHmM6+xJo/cityKe
7ZrukUoeU5G6LK2V0/LF05nwg6wZcY5qNL7JTJaoxnZ96MDp8OkngUoupgQWOHGE
jZZD4/FeU5RIfUBMpRdJKnZWpknSz1nw6TuTs5IbIOKHRawYtkL+JOYkLE7gAbE2
NsQiVERLk9InR9EqBbGrcvepC4oBVel5BkETS7EcC8Qym+D513xNF0SWmWRfBkPN
+Ts7nuyD1Z0Enw6xeP86PHQt7OAIFstp3jT5yQvyUVFETGa4pTyb7Y+HNPxB1D3c
0ia0L8b2++4L1WLTE5Q1WWBd1yXaw28DMx7A0prdVafUOlqviZRpamCescBgycEi
Odmg06JhWmn/Isfa5BLWbH8c3j01FvGbrNHFjU34sCCAkvGvL5kMgX07ritz0fzc
QMwqh4Vjp2ejC2pL6BXzLk/rB37tyLoHib+6Iro6DtfHJQJWbzaD7bWHOlg0cpeW
322M44a7q0wK/LfIDXIzR2eDXrRpCsk7UGm6Ji7rKD7ZFZ3YjXmM4oJQihno2hsx
a5o6inMOZIyg41AXuL77iZknPTipZZChxYcvrkTpCuoLAdfm1L1kQtRsI0/qnkJb
Oh509wxPJbXWsh87/9oNAb7NUcRNmgbldtKzoH3rlB3k0NOSLg+jqh1Oa8YdUEA4
A9+hswWxM/R5EhIvB5gFhAB0kNopkQW1UNe1nTps4kmH+McC1oDl45x+V2Yy68mV
Jj2uYkHnyk3u1Y02OIhhQj1NO0hSl3osrudkFOa6WNsS2yr/hBqtTYuqOkrv3YAK
rnkNOOUhaBE95AF7tRkZGsGHmoVo9e+Flp3EaVFkR0J3zb2x3bOUU1LX18Jqv01d
rqA+dcedrcPrK6PZGxeBRCH8DYJj5CYVfsvllAmzHSwx7DewWQ8qMECIBs17k9g0
LEGvyku9EZy4BcsGaPNDx8FPAhInMZhfuZltvDqxECJqgx6K6gK2F5FfK8V6DT6F
Af2G56kWARnstS0imya4u8QOjtNHisSbfasuU25EPoG8X+BR/5+0ZYP1VxAiPYup
E7uUvVErLnmu8GCibfclyoYLC0JLCaTOMuTNHqyMf9C0LlzCY5C/5KVjfYtfSYp/
8iycX7pgnR6WxEpq8L2NqMvJV/aAh2Isrlts4moCjImEzdGOQwmQryOF2NkcUB8F
zQzkwMVnXCjHqNfHVBIJarZxys3QC23VJcdCtsvknQSwMEY3QQAPWmDIdr74MNS0
Ir+hCW962s3mvcKICfSrHvH3GFt162whUiTPfL9ohcui1D71HdPyXLTGhuU29d8s
xCdJSLi3FE/4jyp2xz/yrzu70n/jFhW9T0RCigfYgyXgc1Mbgb2AMQVEd6a19Fz1
vYAX0qOhC3VaW16SdwX28JYBDg4zTDwrnKqLt+9DnSGQEc/5aj/aFXM9YKx436ne
4YHA3WJhW4ILarLBjWY2tc7+EIEzVcN09/I+NEVCGMfx94Ac4xDoe1UNSTyxMm4v
8K5d3aq8GbbKQ6Z+4gfh1fsRwlapLAznsoTH76Tdvn9iP8QvW+Z9PM0h4WJvG/HQ
kTRNEDSSzpvUVWNr8rNHo76FMTgH3EoqvfTRkH52qZRHzFxLxXzg1fNIaPpsh0+C
q7ZEJMo/87wMolWs1wQBDnxhOPIy3kelwtEv4EegkJG1wVPefKvGSJQbt4MXI8Fe
g5eOFeGdFIxTlQLH+mKettnN3rzcHAu2RcL7liv57yn1MqAP0Biansh6qSCYm0a4
rOZa5R2IAolDnYUVh9x7nNSwu/4+Cn18KLJL3gUzq/L2rWPPFpHgZwUMzi8h6+LH
V1keujpsI3Rq8dee2fIWE7PgfEboJ/HqVje41D70Qtxx94UUnMUodsNWZ8HMiIwR
LhNQC6do+hwBIi/qVvc1PAbB/XPs3F8yh2zVehhGktzdXMU/FZyo1ysjJcM2RW3S
J8Gx31/27+ueIQTLHGnJjM06QXF1PZHMZIraC3sk9EHqiKOja5y78vjRBZ0z3jo7
jtQWBvNlAPk1y4nXXgGSYfOUZ3MR6cqzkDfwhxzLEMPLRBd2PnAxnAGzHyK3c1hY
KoN/Nyk0YKoOMB/WAEDCY4wOaeTrNI9PiRltarpjuqiM95jHbrnHJVtdg/qTgZ72
80CMJlaE0US5sp2N/xqOn1KoE04hLvHlDdYmXrTX/eP0vVMArTmpSdNmdwhOTkfQ
C+nVtvqWzZItBCXoF7BqVTgwxhGd5tLudACcpuYia1BdOzceAfEL5awFrMxuEUlk
YcJ86+vhR644/MUpwREmAvgBjL5HP4LfcoDvAAbI2f6uLQwA5pdrHJw3xlK7hdMB
1Z2kfkLffq2aGpmeK5oc74f9WE+T78i3yU2T7SFyAp1LV6XujKrG2CPuPqRxOi5l
wHF6oeVJeSGNbJnL27INJI7NkaIRecOutQf9M+70EhoFGqPX7V2CMdwp15OAuLV6
m8mWgogEw5dYQSfcxMJ+dE7h6Sgqejl7mF5wyWmejENkCK0igx6gihVCgj7D/hXo
wuoBPWS4XakLBS6HOA214f2DoknPvA6Jh+QowxuRugvuPFagoWS4FXUkYUYL84K7
5WAUUluXB8pED3NXFiJtbwUTWgqgH0lEcWZC581MyHHORCnDIgR/4Cgq3dq6gASI
qPehqERVYxGBluMJy0DFSDoZHbENOmrikECrvSo98eoKDUEVlh7pX5wCWDSV5tW9
jrHC7DoSsuiK5bFCcJIpF1TQHcvXyLdSR9BWsoLH/zFMopdPFpQj9V/wroRToy2D
6AlDLcGmBgAIxXPfofg01yqzcjFZ1f3K8EcuwLIjU2HhfX0JaKc3+sEot0AdGuHQ
Qqa8Yz84A+qSx2hOtjX/e+xwjO3rexLcconXOojcnOSn91Ypp3dctAnR2//0kBb4
q5+aLoS59hnatvyuyMvgVNu4Pp63XqA2dNtJVhjaSoApqvNvvWkWEKysPvJWQZ6k
ooABDeiLzo9T873Ppd7AxsXpwDoXDYTCP6sdxI/MdpWhrU26/jnrLFXyHRAq7672
Y64x7G5AB5M3G4u9ivN3h+3PdSNvQFq0H1a34y3arO2ousdtTPfX/dzfYLcAlgv4
+6ocpxuoFDIzDSEGcKyhchrVw94FdV2gENQ/NBwYFhFPIZoaPTh28svZ5ZejcxGI
PuOlaj9FDGuRTCVdq9k9f1vXkc5VPt852E6rR+9uHwz1hjzrbgeOtiF6j6oaPPGw
vvrA6gjz3K+im/kRjcP+Y5gsUaxCLc7aMCZZPF17VPP8KTBTOjbPcTk35GEUu49o
9DkHR7bptyh9Vhd231xsmXXtLHmvclYc8lmo4grzQF8RV6LItroLRokm4sQ6HY+S
aidHqVXuwY/AXSmNqCx6WclD8Gy6eeyezKwOdm+MWu3M2mEaZ1l2mVuOvK6wBmVc
kmA7xsgvCNcHP2bJj+6hLCrWu+nVy//mUoYyMEURRFwbZvNAMyC5/aLyruVBX6fh
XAqnw25FRpjweM6222LkOVn/KtwNxg7aX0/f5KAl1B0xJTpThlCNTJ6L9oHID4lA
P6El5ErZhiIhz4uzDdsroylwQ6tAFRpsx52Y0JdnhDHpM0B+1SBXLyhY5dbnTXkl
SrNdLpWMyaG65T746/7MAL6KUFMKS0tjdtFWZi5Zxbhs51qj1vvdxS3g7mPriswZ
TgZIv9gtuKGlSUEfnCM1Qtlo4QXl3ojQDRfgf4ag6NZyTq9Eg9g26ap6Jal5e/Kw
aEjAjI4TThVZDDR1MCbVzO+B+8+4HDAF7L44QyqCYx8osq9xC5TqDdED6fBZ5T5v
jvNJwGtvPkXNf0zvl3VgjzeJQiiMKnlmtmDC6ShwASE2lL4be3hyPS4AuWR/OEIG
bF+yH6/+Auc15Bsv/z5Yyhhbkiv5GpAdR5INQELbnr9X0AR6agO0hMVVCjKKo6ew
HcUep2GGXe73is7SK0jSrXZihfA15dtnoRk/XrhKsMhONGOE9YGdD3NbHDFbsGOR
QUd+So7gHRR8Mcowbjhf7h566f1nNr4mBQWkJjr0UbrOxvpuMvQ6S3ZfAfRF/RxX
V/Vlsw43XNKPbsoJNKPsZxR5O0lIk0hujsBxHroaW4vfv/wDG/K1g0xvPYEnvPtb
CArh/96zZZK0CrcYsUdpq9QcMa0EJ0/RMeIlaWBPl2Tmv9zPaEPmRKnXf8f2No2f
Gsc3Ujdab7qtK6wZoJwI7Ve5T1RdHkuvXyOcW5T8fOmMnnSY9LGzwK5Uh64kR4F1
80T+0ZMRYTvwuRBhl+7+4ql8IrVfGJw/Jeg2yRCsq/zy+/EstSlNF9qlPX/6N2tJ
GIuOTKITrtWuPl5QN3RMv53HHdzMA9GlQQF7YiT37tn3ln4grrXHHc0GdtVOdJuE
2WYr6Zy1mbq0F+6xfzYlx6ybWP9gt4zrIEMrUZbTYIMci0sN4x5qySinf/6Og0tm
48nqFSVDSvLmLieAXEvcoMl0ubnDnx810nr04tWAlj6IbxMwL0o9O9xkpSrATq4R
uSRCkUoNbpJVnMhs7WpDEfx+V0B3IlSzHygxlzOVzXvG0RGJl0PSh0uf+2oR4iDf
6POHVuVlzpmr3d/cQe0Sk7Cx9cpSRp/xCHyfUGJNH/NHD52EUMComtgrKAmIHovx
aK0kjDuppXGv2YiuW7SUY9MKdGBvLT1Lwo4x5YJAtDQkIp5Fqd4PpLMqDZzsTI7M
TV5OYcwx6lHgEbsB3fbJeL9hX9Wys25DDKTF+/CNqAeB6UBkrOeYXh8uF67SZm+H
ZeFkUbgkRbndezGJ16alNPATaus4+FMaPcbBuPYgZVE+6JArztl+JaPO2533bH/P
OeuuxNYC2/3Hpi+KCIbdsecp7qW61HqNM2bq7qP2o5xmqrjbzhJNvZ2kTsqQyfkT
EoYoqwsJiv8bWImG9/e1t1Y9uy6M8v6+f2AUc4jmYJ0kRzYielzqmRGvns8Wnpf+
q9sBbtrPYHBEPMVrHVixEIwxoZGEpbMqe3iMlTkaOlXv/s87lSyhLbrKEnBNNYhI
f9hhwJfERyQYqtcqA2EVGo+5EAe9buQke0G9Gh+X9hckCa8XU4ioYaFNq+pXN3Z0
PRrx4J2+lzU+7Z3w6pvSpmaAX7uYoeMSVOgfR0U2i/RZ+CpE3NWiuoy/LKEofz2Z
+iTC54X8iyyynoKbMo+Cs3dKUJYrfZrsEo5c1VCCY7DEdfEepMGv70wjCQDNFUEF
r3/7kHT0uC60ck4ESbuIGcXggEgcNNv7pZPy6or/6xxICWTZaS+aYfAhwMBnf4Ec
AGzDkHj9MwgwaA2Fv/pR7PknmLs2/H9jmljCOumFrpapFnsP0sUoylCv0G9FQoDf
GFiSeZRBS92+L0fl52FvsIxmev/vN3K4ytntLnKbjJIx1jB452zqUMw14AFtdvq0
5eHrGiWHmc+Q+foddiTeRCjLpUP7yGBSHNwHfTgru09t9tUya30oRnc2yjCjcyIf
v+GUFDgC3V0semMWKOnJCk0wuun77N3/M/ISeHZXjxx+Vw0r7P1Q7YifqcgsEuUQ
PupJpNS9mUf6osamH7gHVhPJ5TsVhst/QutvJUQTV7B9lBuQnCjx4EhSnduyH3su
We7qJbNhMVGIU+F230zQjIBrFm3uIV/0qmTJBKik8mHh3nbmb/o9BR5HudcdEUBh
x5VDzK6cireiZ2CVKerRgdVde8i2sM/fRJ/M94ghnj8K1jrcz2KlGrrAN7xacuRi
CwdwcDd7x0MREamDfQlXqFQ0qhjqwaHirU7XULj3nqP51GsL/qtEFN9QjBIvHL89
d3in10YO0/zqldwConLx1Nl/Mv3ISJZPag0Aa1A9d5P8j7RQ19OgbY6C1mhSVJkw
Qybvf01EcIFHsJRFBfcuGQmCCQLjcgkVQ0c5LF9b3sV45+blBR7dYqPPT+OdIqb7
BN+zkLUVkvIM7Eh83uCwHb5fPuXlA/h3gywG8ZUOVuL5kQPN5iql2HGkbNHfSe67
riI+FRZ/oabRCY1TpCbCBkSDLWmK2eS+yoVITwZmPonUez2RhpsStsisTIEEliY9
H4aTDMP7eB6uwGX5s1X+fM++Gbb8EH0b2NBBxmGwJx/NAiAlbB+uHDN1gX+2WePX
nI2KP7V+dF7yJD55rQtm2e8JKZRKWcce6IWzT7CyVKX20wjipecE4hB4vrGv8GeT
N85X4mQyI7P4b7JlQF41mZUckeRoHfPL5RuUsU2Aai8Fw+l3RhF0rZgZw6ZdtxcV
nIQwHZ2C3wywy93Nm/keIN6gHEeH9kXFp8doaXGTvczzo6VoOAK6Pb3wBf3CKgu+
28OXjfKeuma6Uta11gzSvGraD1J2HZzuRj/f7eO+2OcuAjHHtWuGeSZoGWmwI07/
dPG60kxlN3Y0Rc1vfPqDL+FRgr7PGi7/2j3oDnsVcXTWKQhNYWAVclVgIaHmmgDF
wjIJZ11tCOl1sciSGDVgHEDNEBtUUkO/bmX5AaCtuXl9kFAi+fxG8fBeKm/sxRpI
nc9MCWFe1elMwXXh3FrlrR3Kgr1slWFFj8adW8GhSmEBlLfKl5cT+GTxsDrPZleD
jbEdZ/jUnToINbqWG0S2HfR2MICDeygr7C97vvNWtbi8Sj02KvZQovkrS6v2xCTU
kiNjFglcsljTBrk+G0mYXJ3N/dX1grSDbX9JnQgmF3UwZxhWZDv/WO5Nxv8iDwzI
n+X7UedUEhC7bLy/EI56dSRL99yG7vqMEAC3GUOcdGOSQuh6aL8RxyObcQPOGU+H
KmwBO0EdoSkAw0KbHzvT4iPmjz4Akec1HkIHvbyy8DotT0GlFqZRGZDP80TBKpxl
pmkbCNTuKtRf/Sd+jNI11HXMySU3aS9XftmM+WfZKJ9vbXyp2qOwn8ebY6nqX9ng
j8l3HrwSaKykYpfDMDryEzOHFH3ywdMKr+Z/Z9Q+mIjHd81Dz/1srZFoR1OFnb0n
9q42XgZpHXqjdfQq5GOM5iYFX6pNVt4mL1L68V+BPBdlSSnAP8FF0YGjLJ4eyz8I
/jsEgC6Y6SPlBo96SSE7jdf+qdr1cjFLZ5qTb2/Il4xyDh+1Q5QHkjUCDsC1A9qZ
aIVNHDx+VukLO4CZmRejh7KICinmQGxnpKvY6YeyuU6Zu16kjDsMZLxHHWaivLXz
Jj9ZKA2txCYCehzkFvJ1d7Q3a7YSPCJEDg2f+/VRkl9MePm+tP9mvLBFr5eQL7aW
v5wHD7pJ+xD3M2mv7wGbtz1aqebNwVjZcIMwGR4sMEDyQoaf3xDcRwJ64odkqkaf
rZAskzYfMj+9bSKzzK7NftUa6K9oj9fVNvgYvj4yh3KDJquVFwv3CDqgli7MOsdX
wASPA+BtYgelu1H9hEHy9F4or6UZnSOXjvXgVGtaVX0oEx8Q7kU7tkslErvrv5az
Cwwmx0tab4EOrv4orAb53X9gflQcixaJ3QfD+taBhBMvYxYumcSjF9C4U0ZvWgmr
law1vVNqJLZ6xq7G36yD0BVusYoUPVrHPYfOWRB/duxqN/eftIp1gjOcMIEfpo4Y
9ExSNRIbeSffwRndK7dK0tcD2YDzzijFJ6V+Xu2Vw429ieLQYtncv2Gv6ZzIl9M9
tYSc2h8/tVasQPIYggevUVuJEiU5sjjsHPy16xDXL8HzxSi+VUNVUm7JPd8YK1n9
IKaqhSMsmKMVq8dtyAcecO3UEWDnRjBhrfEm8qT4sSChBZz4DncJ0di1LeL7kNsy
SRRqENNpdRr5Z/LsnX9rc3jqb8CSb+zljS+3Dr5LMl6doBFk0Fpm4r286gG0qcuh
Z3qJChGW+xd/NLkAwxNm0N3BACCUnRzjT1dUkb9eH2tYum0BEBxBLY7xUDLQ+X1u
7ILCD2ZIpKJvLeQqHBGdmTot+1v3gYWla6FdH/S6m6HMFpTjxu6o/XMf3j/cqOel
FxasaDpNvjWqFYYdw1W4dOMeeZlMR0/nizRPb1FtjN/J6OXKblvm+ajFsjhtoqs8
iUMCzaEey30qANXLdd8+GWVi7u8kvf9nEn0AIpz6q1xEqPhBvbkqaao/olXYEYxI
+TiOQyLgdZ6yGe8b3u0E4PwBs/1sUs/lluqQIn/Jv441hoTjTgzTt3suFiZiyS19
A63d9mqECUgt3bqv+C0cIIhzc6cpeemagfGREf/Pp+dkw7teBdOSV3Ob7hRPYSZK
KipA5ufGeUvVgiWSSgYPGSmFvx8VcgTZc75pecydA1emUZohc1cgyYdywDNRXeWA
fkMqhXOepKqLsvh7e04tgDypH8v99YX4zz6PHChVVeaTNcN1GlLsUXTuHrJoGYcN
Gd3uHWYVuj15CYs5pDhkugZRD6QDKwMkMZmA+DIe5Jb4BJpFjkGK0/Vjl120/P7a
td0DIsa6rGzSaFVKvdD1+v3CmFLhMto1BF/tSwqT0iBF+cI4hAUDZJmXS7smJ7UF
zyjfai00wn8b0Vw9G1eZGuQyvaC2nkAf+rLEw3PjxbY4X6DscLpG6Th+qVlCiqbt
nmTf1aXRiUO0agiXrbGMuuyBliOoEgZff80h/vud92eYb+YRw2s+D9o9Ktue6Sff
8QU5C+G+KhHtnKjXcHhG3MR8oP0uPQ2X4j4oowgh1QgqpnTj3yjSlN3VBiKty5EG
fopL+v4eXZEoT8c2P4D65z0SRsrzxNc0Mq+/WSDeW2sHwm6FNw1OfAHE7IpPlbXt
ggJK/Hsy2IOuFR0dLhjtmXCtVNoWUG0jgdnQjOjM1VJL4+/oyn2zBI5bD/0ayZTd
8HJ9VsakvEKXnl7tl4nlqGSFGoJFYSm1eoxYcnssLrgORxHk+uciEgMqAPJmmFg0
zct2sogs41lUFCqdOvkWj/6aSF+Jsbz9W11hqUj4NwJs/cw/xPOF3DezACJHifrx
cW651ggLQE41q1aJ/84HiEnaHGWrLvjOD6yU+ja/URVUDdq2cdayeo3xWpc+38c/
ZHvMPF2AsCDctdGgssJygOoSLeNO4KoT9qjAxIkKxnPOg0FZkMWuz+xDR2j7Bdno
XwHnKmIz8x1cPDbhDw6gnc5Bw0MQbeakxN3fyRw9uAhoI4UKrAn1GrFubpjNW5En
icHMpO2fDv6wr1N0cGcehQe+89gHjkrcrwUYSYHKV1IKnvJ5iDWK0gsTOtchFusi
po6XuxXnqONji234jzw/4LoVuNrxwpu+kDsteOsNzOFGgYi1h3H5kKK4GN9gjtG+
y53bQBs7coG1pJ5xmMqZ0l9hPr/ZvsNQXqPJuXYvr5au4DtFI+IrjgIzGYjqMTH3
0YD6CrSAb76Dp23tnSrXMLlk2dT54K6Ak28zSOZyPFwEE4G2sVBW71BHyqY/NDk+
1kY13xq2tVCkW7126zb4ZZCYHTNiCwMDi3y43zKjhE2vj6bwmgDVKNl6CZpwj2Fm
6eiUQSb88ZohaBnpYUHoQB5nFgudGM0z9qaH2qJO3QmBcDCzn8t4JdfWeIuFMxoW
Ah85sY6EYxFITIhwUpyT7uARjLo4192JQl+JzfTXicPizmkg4htlYwOJSYIPaiO0
xKICHEBoSy9AgWcSqClKI9tG9MdZ/k6kH761d6GhnpFSq/K297LivsTlQ2vs6GqW
hERLUeH1pKjBtw6PamuXhhfRd6tM7W9KGkfcFSoxmPLEn4a0K/5thULWVoWsUuu5
QYYCg8lQ8dNUmbkcrmLaMKVuwSD1/aL7jRLiwuvzIr9hm7YKU9+rNkpDsnK13oym
GsLEfEqZqkyXPw60xvawTKyI50m1l9QQTS5T3cVGu/UQJtZqHg1Iq+VMF2GA1ijy
qBwcAZfHQy5eF6R6TRgSlE2LCsIv+yn565oPzw5qaNRl2LebupgNBpkvSIEC5pdO
60mx8KgcpvR9BsnTPONxl4B2V0kFI8gOe1o617l1+ZVfzI3/RRd3FehP/yP7sdYN
rh08z81kzwSRe7ylczaht7HYMNCYttsckbgARhf8acjAh0h6zS0BwD37ouhGwuce
OWtpNbuU1YA6DN0dj0MRv80/in8pArlsjej0AMiGdRapHJeOofqmq0JW5ud6jGq+
f1VEyOJXNhMtCbq1JJ/9jboq0mvsuxf0jicrtWwDDGtgNTHTo9UnxzFqFGBMq0Ei
uLD4JwRG5MSpQGBnhAiimsZNeqvyjbEacPokNyB94KuBkJPz4BOmhLK009vU7L4L
HFE6wmHJXZqPnq+94jC8hCrKtmzx14IVkHkRILb7o0sqFRIbego8RjEWW0fqyqwp
Hv5ejrbA80UMVtpk7seBs6GR6ZR6kTQL7jFxBJCSomMom1UXmQ42GJIKfrGvOJOd
g7gp8qkw707IXkmwk7urjsaNlWiMg5G+LkXb6fcw9ntCiGDYJbOK7nNl8nxiWExH
VcF/uuj/9qMCQMHzAY7nG45k7S5Gmf+PtafFH1wKP3WhPcwB8Pvgo8xAZ/zlQxtr
AfocF50ec1l6UFnYyzyYESy5m928JVk31XkyeJEUfccv5QPX3nM41cowj1fC3sQY
mNDRyqDQ0WSJB+pkxX48coDqgm7t58dBGQ/m/M1+LXR0Vw7Fpcu4POzlcu7kxc2+
yMZgWbmLAfPRGy8rnTLjOi8+w+URNnI0YzA6htDE7UXujr7Ori7+J/7AxRyTWVM1
8lfbGjQ5Z5Njt15ttXkHCqIDSeU7X6fYHmEVQHhjxAjrBjj+bAXPf2AS5GSPJCaM
YwR/Naqm8YSUvhQlzz9PAxRun2id6Dr7pTEDb72T02Rm5+q7AqMzYYBjdLg+rDiN
Mw1nN/U6TpVLLDOhWZB3f3t/aTc+G2fMSggD2ekuXcMU2O6MzCE1UeJrEtg7+19y
Rye67gv7lZdv4cszeRiU08j6fKSYCtGNDS0xtIh6icK5CdPnDcksTR1imuit984o
0Dfem0ExcrNDvSa9Go4XKi+0p5pOQdc1LeihpjfOTN5O/gxmgGJf9Dn5ZXMmCwjV
zC01J+om7FnJ+WzjpkLCz44ag5L2lyMUItoohuiR6iYTovSXjkxOnSWpIE3JvNOp
2msm5KSLjqiI0AKC+6PIhf8ZfOFckbJZ+VcPsuDD/A8xZKGu6kET1UKwODrJcfLv
abDsX9HgzWUa6S/Flu6jG1BvoX7YR6m5amfCtMSCXKDzaq+26NC6wH9vzVFEJvLV
v7YansybG6ErH4ByhVsTYW1MJORROY5aPc8g9/Km7t73JXlYnYtWSouubn2Ew1iU
oF/IIRexMFwr/0Pug3Sn5q0Jlpb7ZbvhiQMfUQQsujqozciBm0swbe7/LydhQU4S
wAmfXa6Rl2lYnYHXE3Upy5v0MNAWx1FTLN23u4nJBhUIegmEzZsqaKkjRI67Prhz
w0D1Hp+JmWbbOzKs9sldI1sM54trDuBQPp8c9fo1dujVXaC257U4SEldtTO0W70o
JGWNG4M0n7qOf7oyrJQNJzf/NxR320NKDxuGNrfWlkuaR8ydFGb4oL5TB6GvHVQu
8KrAEt9cLyWcwCRZ/Hvjy2XTOwmhTG5F1GVXfwRr+0p6Phj2g1EYyanJY7tH8T1U
y2KuXJAoOMFtiK3/1xGAE3x4jh+J5CEWWipBDo7ppE9Zt5abBxTwll44QYtEFLCM
R/XiZ+n/5OiiXbBHZ89II9Kkz5C++YGvDfC5lK2ZOA8utDe5Of1wMsvQN20/jE9z
nnZXcQgp4cRlQ5x34mTBBj9kyXY9uJpFpBAPWvbFy+WKUmuaxh46KAohEPTUKLpA
OjEsW6C4D6gBJLRsIJiShB85PJeSjMBLEohJjRbjx1FrWUThE0PtfPSwc/sGqp17
lPLZwKsE5CV0gZEOueEn3NCFIgKTT0JMLcfsX088Oa8e9o12OdSWXZtD9F/klhCz
h7XXaUczGO35dCIokZOltSSsmOVM7/KVaS+JUCENrfEc7cORuuKTwoHfYXtcqmen
fQYVQN5BhaI6BXuwbHh/qnjaSDUuKFg/oIlPHLY7qJ4N9tf3xjVbj7Lna0N5CR19
andtTnLZVoIK1hCslTAkF1nh2oe+IxMzZvLpb3wzVYCV2HlX2jqoMfNAz3aHv1Jy
kiD0oXE67uvg4opSNrKfim+HwWGGMPEwVt2aowWzsJH5/Bt9+AcVMtPNHehc06IX
IwhUeUKePJd98tMFmGrU2Rlyh6cLzTSf4lQcXMdNkNEJ1hnpCTSPc0nZPvtza8y5
a70RxMT793oJ2WCV7DU+rYs9jo7KdiJLrSBE87gcAitpYE3rl22g/fIL26ocXGwZ
qt7gPi1iYxZJlihyXM1x359a5xlrTO4fjvnOgvWeCR3qu01v8AF+7X0ujp5xW6Jk
rNGqT7T0/+CUah+UairWOnVbJZvUVWnnnsKIHj6GgMp/GvguwOcQRmGnfD4GJX22
cLm79jI/v46Gh+VreVzDJx9t1bTX85qO4ZfTmS7aAfZONxnXpKH5x89PtHsoBkcj
TQ5L4XuqpbKKU9oZ8d1dO73xwhKpG3n5WcT7jxc8pv5h7RJPF2YvBdH9z5sdHkIu
yQq2/o2feXIVJhd17YSt4v5gqBfGH3HlYm6cDvUH3lwIrNVZezL48OxMpSGPioDI
8SgXU7MnKuQy7zD3rao8nPjXyaUDCvhF2artbW0WTUdPpxOVZqR5xIBwlw2UCWll
qc+N79ZdFQkcoUSCWpKm+Nl9JkUwh6mETYmIue72vr51EabsFNit+XDEo0kZHsSc
eE4ZfLvzdS3P8d2nuHGMd3FFozPUzAHp0iv/TghFO8uf6vtu+hBJ0p+/PQMIGV2F
xamhhnUXsJhRLFdcGcXVrP/RNU7JVyj87hGZhUcwu1G9RQSc8iMWfpqXToJg595M
PxC/2iKHWqEbkE/LAgmlk4Zm/A8Bp1pBz7zvz2KG/MfexGh3Qkic3PIuSl3Ai/Eu
wHQEmsepPnUNCxrVA6nX5U9n4tzR4R73zDdsoaRNkNEwxX8Hq711+H0QwhjUrtQb
6q0GmLgnitQ3MSfrMK5p4/BG7aYXpLpXapIJ4BKYjPrLBm8OPNp+K9ooZp3qaRk6
5MldSpOj7do9G3rktO02oQ5i2G1Z2AFuZ196sc3Luj6p4hUkhL4bixCfcyQxuQ/c
wI49PAcCdFt+q0tv6h8p0BzCsL8jlYgfkt+nXAAhCP53g8U85PRqSwPGE+mrCyOX
nBVH8XuFlDNSRd01ugfnZEFUVl82KW3LoPNcdrszoTCJ5czq7KlhOgp4DSGOPrOA
0vFkeXIqXw2eq9O8WUq2U/NtdFNtraQeReqvDmnuQsLZb7dvIB4S+qzJXsK8NGcX
bfKowji7UrzEBVFfBGrPfMKMObLhE6iZ2lFYRi0aiyNeU4v3438iLyGENyL3PUBA
v/buBMZKSmwQO1M6c8MvQ3OvnYEKQkIxpV8rsi2q8yLSW8Ilk9rTK9qZcOH+38IO
cG1iTaLVHKkVGiI/rIkUpqE0NCHLF0kadfq/rv9Mcms7eXuHRDuRS+LPphYcbj9Z
R4cHmTo/3a/GAWJYUsSIc1iESd6iuDGHJYbYikv7LVw/YgMOuqSogPKxRtZvfVKK
ieTC5EdK5cLuL43+Zm7CNy6ovt5sYMQyrOMCbWEG+jOtJboj93aS+2DDoQ5wsSiy
NHa+MG0JK9VjE1VMIFioVPN1xxMOBLcU/jLpt280b+xhKmsv2pn6jPMAuD28jE63
zTYyboJViQQmY4Jg/hWxh0xCV8/pPrmfpxwaEZGpJ6ncqoPyiN5FUBOf6mmWU+5x
rT9/3Gw4HxSud3N+2O7u2LcBoy07XOWOvQfd13IYNFnUelefN+vQJIR/++cRSFe7
8AZhFAL/Xj8bBRnc2faS1bQxuwR/Ep7PEYrK35rU1vPyAihf2Ux72UCygYvh5TJr
vmqpSndO7BVPM0aAz80cdMsC1q0qriN6nD255Bq63MYYgAaYHR13oER+TzAi+tcs
gN7v7J3HD7px5TDaUocwAjG6VZigAgDOvES588oIQYjJvPwu4q08MXzDATMe72B4
CMUxp2O8DxNJDrRR/8y6MDk2HDC2bVelQywklboFYwNUe7DZA6NRIIIA3PE7Z/Pd
gJe7EcIOZTi3LIgTuJtiMJOwOtKz+63RgyyOo9mBlGL9uMpxAYWbwD+GUDKIQvO9
PfCdUTdcjSwD+J2kcnuJZ1sIWRRd93Crg3/GDRg0RqbCXHZv0GUVPwsE3QvR+2cz
BAXL3en3JmLIulkSgVyXweh8U4ofb3ALK78K7PXcMIaWbNLnWf9K388zjvlGZcgt
5szbL7dJ/CSY4DQYEW17uERvU/Tls/u5LEaSp6BI4PiBFWgBivEHf9dsDEy8Ccfq
weF878odmeRSD8eS8a/TbWd6Pd7zZqnFXYh9H/GdJRi4hNZuf9yxHreJTKBOWuNI
0RPFx0B9EJINz/76NX7GVx5we+mMgmIcx1y/Rb5OX3f5eE+gDDuYnZfFUNYQWa7o
hqS2zmH6pWQoCBiboFHIyq7CdVzFJO3vquVu6p2t4sDqJ18ErqEbLxSdXf0gKeuE
dNo8qKA/+3VK7QD8eipPdtX6UYWVfIe9FHQKnZTQd1l6YYX62dJPIOZql7lOTCsY
S06FweU9IKC7Kz1EVuoJXNhDJ6xm0CbY9E+OZLU0kAq2n4Bu3AtnK1owNkaM06DR
JmFIp5jlLtZ2AvedPt9nHF7db8mQEEta8ymU6Pa//cZvZ9cNYGz5Wg1dJSbxvLdG
BCDIlegFvfRhfY4vHue47H1KfKdrgiPVb7xAKMlEbrzHvwLlMvpzHQgPBkAGIrzK
+oZyJTT6aEQqM4Yl/C2bgKVDK4PA7YAPQ1CE39iaiDhi50b9oD1wZhQSXj5dwXor
iW6w0DY699nDp4zMxvi285AFEH6Ks7fIyRnALSCtMnyg/cyft4fzAYsOnsMFwfRb
HZXbctRqQuxzg9rVi98vf+KTdMQJb55QWmsfTKwfjEJGMS5D+CVLsWtEYQg9vr8P
13MbBOLCEQVsTWWY58G0RKtaBcjctY+FSU+64Id5PxI3qVPeCFb8DhRPi/ikpvFv
ILQX5AfMT4xeR8NU/9NlU7XpPsdRkmcQnU0S+M2NcV4v4DLkS6klrfBKImAW5FQM
RzJv+ABwUFspt1DRMSy/VpgZKI18q4PfYuXZQEQQbh0/nxaCNtUO2OM79bGfSxNp
7C8wtGhySBNma5Q4u3tWGms04jujxLF3PTeDjU8NBUPMZt7iQ/i8cLkKx0lTNHav
b2qxCyGcQRAlJLAA8m307Gxw+OF7bKIVgAOjfDhy+OV6GzWI3SrhUATpKWpRrnU8
4m149Spqy3tZZ1HisDGdGuiUqp/2Nl6duEt4XVtUhu16TXO7VwrgNCFerxcpZdqF
Ie9k4mn2VYJCxO5CEnjVaY84uIiXxQCsifjyWRiTUMHyf5EtzkrG2hs9D7JHuqXC
UGDkEF+m7h9Q4+vjogfv6d7KLE+0O6xl/NJ+xMBmnw5Ub+5nhJyyx8PIA9Gst3KI
889aGmMwDGEOZcAXkptKTkMvG92dyZQyTf2pVZ+RZkErcydnZZahcbYknLmBxjPT
nlpm7VxWWw1uckprCXb99TVIvcRIlcx+Qz15D+E57t92xdTdncUBd/1WCYqO+5AY
NRRE4eGj009HniYmZAiaYMH3cNpm2md9ZFVThwPMGgdzp+DasyfV/jOdamFjWlCe
kt7RtoL8ELy9qmDUmv18VQx0IUEdGxbEpQ9sPsTUz2wB/8qvMt6gNY5hftbCUD+u
JJ8ENHlcLERCkKA/nhUpsiA0OEAMrv+SzcVP0kdo8IGA5p10wxsVsCo3U+xY+0J/
r/U4ZDPowIR97BgypWnv8dzZ42jl5OR3ZNxQaAvpiR0t5PVZDVC0xbrFSvjl9ekM
7SrMbCteWeoWNe27ieNEDPdXfklHOzB3En9A/wEPZu94SZFJumcj0dvUC2yQrA3k
aeQIF0Rp+99I1UAarHSwr9bPJPI59pkmtAVWvqhTus8O6hueCH78+fiLXks5AcwQ
trpLSLqTzjQuwDmDRk3COZyg7fEBJDTIjNN+hehN0dLbh1WQjOd1Y0A0m1vHHzte
zUUaZvYgaDGU08OvXKTpC+Ck81bEMk5TTxBVNWlMr+acD+INTNPA0PW607CVCjBn
UaMTVsPzvRsEUBbFLFeBx/cmqLv6UfDnfDZxjG/5J9d1diqBKjXVpuZ9Ka32+8g2
SzMIksW9dRAy/SnvVlOt1OkFTVaNwsPR6xeMRuW0ff7ncFlmdseYODJnb1XNvrdK
9ZVpnqV+9u1gig5HfeCcr700whs/oERr5/6c11iyrh46Tgw4OVtMBEWaE06SKu6h
pi7yiz12mJOD1VOHeIE9JHWQQ62nQho43P14KioQe74uxxuoOpEpURKK+K/VMeVz
h64+hh3+SxNSJ785CbNCSCdHtu7gEH7XBLg0l8s91qpZYRefaPKjGDjEuDFIEmVs
QwhF4Yg20vornah0hb6kFKQn1/bgU++iBhxaPC5HBhel+b+7ljpRUxvb6dH9hcO+
sGoXS+h6VmMeBcgf0zFi/mvB1V3W4ZhdcQiiA6F1DygPcqk8Ldj4I8Cyj67gEHhK
N/IIRLQisYhbxFAvhUR6JUA9XNtAXSozVSiM2Phx+/uwWQspD+qHY67vEDh90vpl
ddxQntkgyLwtALudPHkRKXEZVDRIAHrR5MyK5VHIakDcnMI2VMzTFABePrZIGhWk
0wydQDcluEjxlLMF0QLWYMbd2CUeazFQFpr/hq6qBybmL+tFkoczMjMdzN+PEI8t
lpIWQhME5zpzIv+mm2Nzw1qrImQGrluqcWx+N/B3PQl8M+a/zCk8/BZIkUlOM8no
2x5WMCM8USAMC/ZCHbLK2w1U4DWXOiKNLqCJ08Ck9Eh9CW/pc74GInLWC2jEPg+9
yw7yL/frMVf+1zTEazyesIyS5x9R1Jywi+vIwwu9+n8ihq3t+9oPT4cSMEmDguek
a9LnKm9YVqJ6NfZHGGu/I2JlLsGzJQtzrQF5rEunY/tH8LSdU8vagH6tW1wpz23l
21CeqTRdmJc5Ygh1JNds/MjE6diwgd9kAzZj24fdyp7vLo46MrbJV7VCpXaPPUy/
VCPsyIlOLU7tobczTJPBonRyJLYQIaCFwju2jzcEjM2AX78N/NcR6aabhoNq/0J7
g+28OAbnLxdgEmthvJ/P9AhtqVvYCMdNMT3RzDJJ/Y01jDCrMU2dvWGyaPl77YpB
o8au7PIH9Yv/arljVZxgZNk9/LLuJg94hpAnhyYvSQbu3uw10fpKXj3u9utN1ZgN
9T4xhZ3vJIYKHSdQnFIoEt2N7zsEDa5FbcOYwYMdIA4EVVnC+i6Zg8UP6JuA0Ff7
4LHD9H/djb9F7O10mw8N0WSXIUKUfJOwMfSInWyFLBtnXDBBNHHyFaLyw0hm0qOm
Snzf9tJ3ju+uUHc4LRhHaZL6THZ2OUuQdu1Pw0HZQRaRUZp0HLV58S0HOq2ClRtR
ecQyYHf7nAxf78ygFfUB2eiD88Z5Ja/ARBPqLxJyt5SdMpf4b0YLZUy1zYwHpRzL
ylWis60I+Z7lP+E18Y0IEOjJUkDhrXw0JptEbSU3CccV0aYm+BYVepYR6EGq3b3w
13jRbk5B73iDu7n/wuE2hSBUeqGW4KWovFWyts2F0/wHRo8k4KMmCoM+mnuICUw9
3a2PmijyPQKBYNmfo+am//djAG+vneLN4G0dpflJCgjnLG369ucKtabghs9ktmGv
ewCTdLZhddxpfrT+krfYCCaBXxnYVOYJdBOX/Qpe+vAo6aUDKT+oxXg3f1JM1tD9
vwYGHF02tdo3FQnfcY3f7nHZtm4l2RkUIvdcNKnUdVTk51ldhUvpwZBzPRKfsJiM
9vn9zPLo+w4WTMlWzRLvrctDAV5NwSPgsbJLNoW+oLShvBZ7fO936fdV0do3Xq7G
rSG3lNNWpZGp+k9vhk5z5zHuVOTncL6cFlIoCC53WhRzetFTg+rGMj575J/+4no0
JRcNAqNtKXx/Yrl8Xo+68xJ9lkh14b9SgsRRJfyG1kaQMx9+qWOW9FEwE3k9SNAj
X3cAJSJoVkBPSaA/3VUkxSgfNRQExlijC9HRQRA62xK7EpZ4k/JIz0HdOxDNdDo5
BH1Vv5himIgUU3vWk61VOFvUzW6Zu9cD8SDfZOxN7oe/LYn8O2hsQ4UTonTHbYgm
8Q71eHEyA3in6dWPscxhhTACn9XhEjU5NeNtm5kgzDYfKGiX0U7tkgS9w0hgUER/
rk4ujOOCwoSt+CWd2G7B0CkgI/kSupFZmRNO+FdeQnHQVI7gphPbwOzaf6/cLxSN
wchyiiPFIDeBE3iunxR0b/xe80a8dhz4zDoW8C1J2+oYt/WO7abTqfqNgGpFZT72
Yrf57zOlppEWSMo3ExUuCC49L2aR4ToRNcOHHGKD7FKFeOPErbwCKNSG+LkDmWng
Rf6Uyps6HyQc14eRioRZX/nIks8NY9A9bg3hW2hxclZemaZjvR3RdSKj9RnSVVWH
lUwJDiKmPFpBpZuULwzrH9PhY4ovHoW+//+7hEcUEwUI/UtiIDNqssw4NS08X4J+
cHRFL1KDdl0Ha9xrmh16HIJQsMDLurGHEI2MrViaVwRMErJGHOGY/7o9Zm2tSWNs
6zE3ylCO8CZ+232MxqhLhY4aqBJRW2p7WMstUYnLPZ7FUJNaHJAFWv9xzcm4zVRz
2AvcnuIbORstLKsjuYX32Vgcg5CiQ/gzYOOMKA4mabC8PaZAb8V9KTocXRQs1u2U
kTIpQg51ZQaXipUEduu+3mTCexSxLmeKhQqXFzP0qKqqixNcvdhjZasN+d4nqI6W
elTcLQd1welb5yyk3M6ZO8k8YJnXZnJCkVUqx460XZ5isniaE7+oHIuvTGDufrIz
B6Ke1X2EeepZGWppUm0lf1Fiz0AerZZ0dLvTCYgQ6K5m3Z2ytaNLbPg6rivOICvE
N+1eiTNxE4nlSuhhUuCXMai85pgr975P9ReL/TIYWAnKak6gvLk20VcGLoTcAF3G
mH/qtUwUW4Wg2cCRCh+N6SC0tEh5Hl1d7Y+UO2mSpgCosoQGg+lWTgivayv+DR7P
Wjsy+jUwDb6+Wq0r9t5+rFIGsU5/mmFSlmxu7WD/UdtEgdRYA/x6AUNohk7J5G/8
ZS6TDOjorNB+LO59NvlY3NkNwX6x2WEX4ursBKxf8+uxIk3K084vdblMgIreKJgv
t8uaxRg3YDb0XCrgcwLVk0qj6RJD3REg57PIcDiFs/24ZBbyC+hcRkh31tSvNVEm
PPpv8/lRar8AHvkLqazIlN19R+sseNxzaBPUEMzAHU8Tw8uvvsREGCEH28GIxOck
1Ji+eclQ8a3LSDyaTeMFIunqKOXkdAWPMKn9caC4s248FDaASUc1pbh/qo2K6kcU
EejMtTpHraX/+ZCXSWD8KWRMSOpj0wUqUCwzxPd/AOY9wuQl3WPHcwGzSUynJ0BU
Tqx0nJH+9zPLt514Ca14teTlposbdSzo57PKy+fYXHiNOa7ioHWaHHboZcdY/3NB
KK1rRNj+mdELE6Tjuhdbvr7C5JGs4boAY8k41bovBV74vE1D8J2clX27zBPVRo+o
/JdixMHBveOuI1DpVuQk+B6K7Wcu9nMqEMWwG5xU7r+3jZzGfIvu947jCDMZ0Aw2
5zzRNSLLA+4lqwxmGjocBP6nWp/hr0E4h0M4Wg9VvuQYQi5s4Gz1wxoLTvCktRS0
glq4YAbYdfggmRnzZYvqVEMmxIKHQPObTFu4S4q9lSSBAXFAU7a80RbOSNCXOKUI
zyyMF/2GRVZONeJW2xI675hR4tufIbK76UnbqkXWXvePgAcSyDU0Au5x4rfyA4v3
f08yABVI5hf6S+XwG8CZq2Dy4Vb5SvkC+CBxp6AY1o3iIhuxaQ301ySOOY5dz7LY
LNX99vclLcj7Pli5ZkXDxJ90hAVuERvcKummys8rVs0w5vMP77l07nKgEvWF4N3R
7I4xLNPafteuB3RBqUIQ391REp7p3JCIcMG5S744zBudwWtw/jXIKcbnDGzlwSff
3sOfZdF7BcSiWYb9Ec1FrrV1boAT22h4IWOFgJ8whTuYX3CtpAEoQtBa70j8D5Zp
SXo36Bn5vn2uqWV6vlyuSLROinc2/za+hxAyzcGHCnlx+nop88lX3np73rL+KaUx
DxmMbdGHIdyVujYuo1/Gn03ME4WILf/fuBesb5ZhsepTWhdVdbV0imdaaxVYfrur
Vbv9l8jqlifzDdQHeHuosXXtIzv6B+NjrwvNzInXwWdYe7Sokh5GHNS6DXNgHl2W
IheqbFbH+xGb1r5be9GZGqf/8P5DDaKFO06sAijUibya9SfW37z+pCwLITUQffab
7CmFbIam8usStvGy9wnRDY9HYpL8rCreUnChknpYcCX7C+lGUVf6KAQn5yLMyqpK
g4EA/E82i1T/P677t3WKa7TKh9m0ypipbKuG8ItUh/HnTTp4iOMN37LexmsL4TeC
UZtGfmcuPAXp1dkpNVrVAuId0G1T/WVph7xNqoLTUNu4OUVucbU4ozP2TwMIZUIO
YiNT9YWsvYK+lqjeG6YW/7mXjGMpDtlZEptPXS5wRixo30o8ZoOdCAypMH2VsqB+
fgLJYKAOesUKoiM0A0Ywq6Qp7BwG0tOR/0iSpLJaH1nhuo+fzeUiYLpHqfeFwB4t
Wtr0z1v0dbHLiTvM2Q7l7TWfI8EqrkXQ2vxL7F1wsPL0JcGsm9ppm9htyeq211YM
eIsdtF1NGJg99KH8GEiYsNkiXPCj8ScbMguY4mP/mAMG1MO1iSxgL5owhIAe5f2x
9Lzv2FfLjWins99cNmE07FuoZOOVX7odnkYzKZ3SzflNwmTT2zApnymyNYIfuBuT
zyfujQZd4BptKsdgNFFT4AjhxAcEZQVKzZnoT3OHKYvxpQZ+s4io/leY1/OI4CWX
hs2vpwH7FNmIW2oWkzOCJQ+yw8tIU4Wj2SsCwnvLc5uoCsAJBNM0jeFhlvznNBfZ
veHd59SoLwsUYXhCPW9c3yElFQdiOCUYVOTsVSjlIbLhidIVSuMJGR+bTp+hAtry
FoSeOBFf8UtL+fYQ/yZOGOwoO17smV1gRt82IuUL1GUHnFX4xANmqfOqWF0JWoaT
1W2o3FOpRYJnihzKVRHJkquxzh/CBaa6FtyCn23s9lEwS5vX2N2bmAejuEY3VOiE
OChkka9TjeRpx5PKp32mhDOwiEp5yLeG3f/Gnm8T90dBoJrW1HNmd5IW5sj6usOy
PStIbTXaWl4M2t0qjKnW0Jurm4gb4wgvU4musPj+PK748r0tFpuN4VEZj6uODDYz
NNZqNpI0PWsAtwuikYaFqczCqC/ONyRvOdvL0cUmlKm0bUbZrp4xFQuaOi7Ym6o9
oLlynk3BR4AhElEN3sXk7GYve2K3YyjmksRyVlIJUl9w1KEPf7PJ8VZ/kKZ52krx
VoAmiurHG1gzFCS58LnGQdFAKA+m+Sgo4LWO0zEvcLd1BYOFdyWNH6tPZJlc/z0D
fOf4VGZpFBdDwmNT314daQoMSYWymZ96QUhdtfxO31PGxpdr3MyGaOwyMg7L8bs0
d+I7ZY60mOySaAoCq6+k7Q6jlfveNZVaRThlnoobyuAmeKGqDNhwfUwofgarooxE
/nPtnC5GTYczs8WjOJl1ZgErXg/10A/ufJPeQnuKD+qHm3gzRnm6HUjlvzEIEMdn
LePHunldi3/fy+s+HuJPtm0+BsRNCvwhZmjvcw6+3Ki0TwFsFjptzO8XPYEzY8Jn
hYVIde8kGsJYUO6/099gwBAVrmPFGQPLu3Fjm1H9L5aFw0csvLeh+Y1o3+6JyNwz
9nafezRKKSbQLrTtJWouAqTf8EX3Ay6YcQAqfLy1EFMEMAWRyIJpjaoYmzsT17YL
UFnAa0RvnEVuhtUXb7Au6uxJFl7G/JPcwJcqUwPPG5Ls8JBtdwxVF4CHRo0YfFOb
/YNGMLzN7W17MeoO4VaWJoDo9CvWtdFFVco+tmhFquj9+lsDS8qyQZRHxcGM+992
jyG7qy9r/bpdDI4poMxZmL4/yczGy3AFhj+06Q5aMIeCUTLX91aBA4ThzZyp9kES
bdmuzgHGHnw8YKgGynlYlL2zle8bxo76n0ynrBRFgd8nJDHJ+3PNUEPhyCkedKHz
aGOlfqhLIykmm62KlgKMFBJUAk4sD/Hl3tC+BN9q3uL0I8hO+SmiaIPkNM05WRcG
2NCXFdwEk0SrfgfDcGQy/q72EIOQDyXzmRqS/rBtt5RzFurddNGHLg+tABWm/KeC
/CHIpe9kQBGWGttR+JBqsd86uMCHfQkPUMgp8yO7gmbNokdba8JzpVb6NjkfpQTx
RlbogPSe6wpEgK1VIs9Bdd8uHN2pXNNVH9Qxn9m4n4eJZ7slMy0bwS0Ugw6vXG6S
IySxLzRBu3WaZ5/eH3y1zq7ozxklJsK01R6veImZqNk3dCIJ4T5tb+GElUht+Q7Z
pBT7RtsJ5fJqm6Ozcc/v5Gbg1g+DsTVvanYsjBgg9SFN17WFVLgYJOr5L12pVgJ0
ssJSys3M7vpsN946F6VC3zLVSx1MQDRyIzV3Ueir5egChZe6XFh5K+v9hnuxY2t6
4GyqH9iHsnphF483g0hpQpnmHkrlBJoKPLeiKLu6A2gAAOInYKSSDKosNYoaL6B7
37dKE5/StF7+oEo3f5rRPs79/CFq02gJeH8MNtC5kQ6svTxOcllymGm0o7MsilMo
cggIhHDJZorflc482qj8+gC0ENVvTt0QddxDj+avke24r/WZX8YsIl+QXEM+hHkT
cF3ksK75ViPYadjX1oqHPXulWTz5m47+3fDomiyy9p3MPS7wcpJrxvnMkFF/yDNr
yfMeVuJR0YZWdqNY0kOo7eAoqbjiq1ST6/S9iVpyHAvKFLJzemFtz+MNLfTZbOqc
1kFm/WzRWYe7tSwPFxZ+OZgJep69e/oEK+afn2P2OCwOoAr53w/dMuGs8PD//60l
OV5v6wQNpsfLT4Bked7BLHo7B0Ftmvua8aFaf4uVQpt3dvehAPhyG/W8p8OrEw/z
sLr5ayq0HwadPUMgKEyxgaAX1ns336bAzWwx4z2P5CzCD2zyZ7gZYwO1bbP4zHSp
bc2QRbbgPNpIvgCX25zK1HB1dQQdW1dxim4flKZcM7Jmydz4/2p5wOyqg2YF81GM
eI8FMQp+prEsaxaEa4yYLhNRlv7n7xnerCIcy1niw++T83bmwT+pjh+dMmxBTkRw
NvTFuHrBVei8Kiw9AT7E9rG64KNhEz/2pnPaiSnkKJC31qpKl5KARxhI/WeVfwhf
vGMhsWT+fWhGxeS5D7LSwElbUgyifMyfg9ef+XsdRVfa13Ntn18L5qQxf54PlFUv
oSGIdMISKBJvYv3rpyQ/g01t1DEiUg37f8Hz9b4QqfUjql4oKTibQFRgfv9/SO/J
+p4v0F9cc/hb/W08kgnsgE5nU7HgTaR7p4oisBDdgBwwMNW0kdQja8fSaHo4rvZh
WP/bWKS5sEYNrY1cWCRW+J06Zp8BcEZbiTokaS+LghVKawiujF6RdSzqyZ8Mk+1g
XNt1qJTkq/O2Yl33+t4gL7pf6Gf8T/QQkpe3IybrVhnv2CoG0M+LA3uQCa5daZlL
VjOqj5JGexcoP9+B0qppWVgh92c28JNZY/mRhPEVrb35iHk5QYEmPfZ7/w7CtoJa
aZzVE79HhKvDi6F7326AHgVYjcggwSI1tPDq97S3itRE0cFFYnmJvapia/AcSOVd
EQT4phApppA1kofSxJ6TL1UAWB4t05FrMO4iS4sNcke47SUv6dzkyzzCn5P9ASTb
5MHrMP0bHwJ/bOVF2MA7JzBUMm1CKvNs/R5sh7GBLExbjNweNRJ1AOYAfO9JGNlh
Yu4/ZQ+yyJ2xkTi/oR88KdCtR80MkErPGTEpgYgGRN50WLkf/vmsI7xZfq8k62OQ
vuwwgfqxBF5ieBqrSIOmxWK/+BpW8axg49jTy1urGK3L9dar2juI/7P72EILKGUE
e86dtpAomcgDuplHWE1fhMOzL7w4w6dF6HWypKuB1TYMbWGRJcPaHmSUn4KUFuip
m2ymgIQdcLF0lPQxM1Ota8WZu1WZz6U79aVLXCf16nHH3BPW/I1tEomToUg53w+s
N9XjBCHrZ/tkLeravoKfQDaVGX8xkPnqY4FzSTPKSQhbB9vrWVcb77FSqjIUdVWk
a2pdg6HNo/2mXh0gUlicDQxHAFocTDnIzXTUJnPAwT1ZQYEhPeI8JNxsS7+ts8rw
eRCSKg/ovg1TRYrINeoFwzcsVN/+NwAblGbhiYjTNEknLk/cVh3iC64xuSr97hnv
R2d9ACQ7Q7QgcY3gzmBc7a9I953SgcghyN4CITGwKpg5IEuGcTuktB2h0j+O83hB
t7FPYeGc3fEWYgdJr9q2xdKMm1wy1OvYcRd/BZog/sBPlskRl9U5L3SenJ/NJAzl
kn+dEESVKBvDTp3SDMdGPyvNdeW7xEBmc1YD1r33+Wnd1A/V6oKFvBqszghkFdgb
D5qMnS74YwCmu8dEpEr0AZhSsKQl3I29E+bwQs1p2B4OiX2TLmDqGeUL+tr6qN9p
uUYpS3LPunOg/nQ0SmYtbTFSjVZwqByyBWi7U43gER1yxwM71EjwbvLf/HG+AVDa
bGpa6/nTiSJpJ2Hh9zvyFC59RXuS6Zkn1zhCghU5oQvljov1ZDQ/OxMT7RNk6TYf
5mCVfkrTXh+ZNVN7d2IUSuADVE2VFACq4pqpQk8o6ZThx9K7h27ewRRw1nX/p0uE
jOPOFoDD2uzXJXQbF3pRSiXvml7vZPR1cDp+F24jMpwGg1eeSo/QiPR9lgwUZzFw
hn214LiN9H+71ZISyE3W0HqAsQk1Mo44FXEB/ZHZApcK5iwXR/6cmHT3vdBzrseC
ZRZx1JtTKPbyNJ0Wnh/xSsVfosCoz59BgQqvhTTsf4/rb94LiOYGymCns38pzuwW
iZ2Z6ugV8Nr4TO7RLodEJ3HwgxrDTMizm4zQKd9dmjUyxWBRmLMjqlZgBCtRU2/j
wjIhLJlAf1yf15wGGzgbTH1mscELPyAPzVcdkSiW8QbW0BZDGKS0E2SNmgVioeLn
AJmYd5YC9HkQFbTmpOcoHBioL/j8ywd1bMsaPsH1IkJ+RcLQe7frtEiKhEERPlLX
58Nagf9PBtNa4gRVak2DS1KIYoUO9y9axGDPahmN5QdAWRMEeIjkFCvo5iYLeKL0
ePmJAk89YBKjwAkXxa9B/G7ApMhozrJj6kHrwf4Bu3GnyZyQVwd1HesKfUNvm+fB
0rAhBTFGg4ihcHJKUqcMw8Gxg2BJa4nU361UqkzhSkm/G6R10J9wQdqNVjk+99ua
vLWign1oMwq43pHn38NVhshyA0VRTjJyKf3ocWzFPZBoKlygGYllD5QdJ/vlUIfq
kCH/p+9K9H5wWvpoVhGp2/vFE/MoftGh62Vz+h6QHIyOENWn1fIkyLdvrpOX16cX
7meX6LirgD+IGrNJczDT2htw6c/BlEu0cQJlaABMBzpAcghkoKGWAOa9HMgIEjUs
ON2Ie6TiQ3Ps9UTnHY/b3YvCEGpjuFN2V4YpkgXe+XNw3i1kwu0g7642w1mhFsR5
pafZFXlGXXT9YnhF7VyxaF52q7pzXaZBKn2nnzOpEdwX19iUciVyI1kHqSGlzUWl
xwwC15uU05gC+fhjzJpk6dJ3/lsGuOMtthf/SYlMxNd7H5mT4vCLF3rHOU2lpsBy
5XqzWSRNBmlauL7bXFDwQbclSREBZuZGnMVXJSXGQwXOkQoQZyKqF81hqKAYq6Jd
aNynSyU0dIBsrKI53UhGciDFGjY92p1S0tErBzygjCMIXdkoBqHGx4VSXUbLlWKl
8EoPQuydgYpextx0fHYzWM4pVkcmqZO0NXOF5v0eP4L4upFKrWwv9LneSyyD1QWc
jIyByzhSEIAOCt2G4mNvpwxGq4Z3CioncPnuOmRG8fy8Jk44XePgSHeyccjPgiX0
3w/TEQCNX36UlcpC+b0IxefqgdxRB2VKl7HgK9m1y9HgARZM6KWBAip+wLv1sKLP
gVOsVVj4XGh0DkdcAl7ofEkzheyl7OZoZCeSfAITtBTy6dDKxonKwdGVe1AUiiTj
9BsmWlyLd4MJOrmWXTWhSQytePfZbWB1D8gmhbZCEMGnkmtsUMpNGj9ljpkm70za
3sme6r6/q0PSnMSs/zTr0Cs7ZbsErimF9doR/gUQm+owhNmzgGmBiT31ailgkAwH
R1Vtp6VJszyiWeRhkctOwemZcBhJb14RLeu74Ii+BmYdvGorq/vzKaUvWCdDjbf2
Wku1qQ6A2lbQbLMOIw7V5m5U0jpBd6+SmnYeZsOpa/tvfinFgdGHF8un3g6pqUxW
01Drekm3BjHs0KimfxMVJDCJRW7w+WGjP5pmwyrSm7iFK0jt7/mnIJ5TLqCvAH4R
b3M4N782uJFle4hWl/PIuwkZEdE5r3IfINlTs3z8smxOsR+WG0tzpTOR+m+GO8ZW
D0EVsAaXJtCJO6cjBN0TXeJ3k40QZguDRFmi0eQ1RgcLuYmx/KDASm6TA6ZqOVgo
+2dewcVymmP3mujSJ+GQL60XpcVe/KriGXAM3PTKc/0lgxB7xy75lAzUhqDkgpCC
FkCmnKbEGM+nCw/OXtc7JYvWvbsDpsPKRWdyiJ2waPChqrotdVEKRMF5/pK0qKSa
qz05D2CTiV/n1vHUbH5lbG8YpUFbJGOixgm31NA1O3D2s5cWI1C33HIJV/s/4PkZ
OfwSXT9sNFSmsLuUPtO75DG+m2Fr72uhAwq7v+fAG6OPl9nF4bHdRDGrMowW6/Mx
xtBCmkfxgGM58XLHo4exioM5uK3xP4CsuUwyIk6lYkcVwCmJwPFgq1GgSG1PmKHS
tcJXicAXUpr8ro9mXGTdiJn7Y7Chia2NdeA2wRDZTYVDIq2YMx9a0t4hyAUvQHzs
zQ7SKMfMpl4TG2OF/R9+JkbMNews+0CLfPmYS2Sk3OWNZP+jYVQ2BnyOLW/7MkHG
XOBOTQjn8EHmhMSnTGXnuQY3rXoUtkEPKocKG6crhD5p1SbNiBwS6fytgyXn1taV
uhPA54T/PShaeJq6nvyi04X1FZTUwI1F7Oe05168dSH9IrQgzlCwkXlpM28zxJH9
Ar8hLyBQJERyol46IYYCzxSQJCRtiPa3mycsUNoPkI2jDrhWaP7u+Znug1e3i7YV
r5evXXMtCU/5gRNBZIL3bzEGtUFy040YWN095TCUlEOn4SZKNqHIu5ll0rRS82fM
+atQh8ghHCuhwn0MRjKMRfVDtttsrlh/pf5dnFJi2JA1pWtQ7GOw/m9wpCkrHxPP
1dBbnk1HFLpnJ6U/bkE+K4+m1tMSXy9Ubl6Y1cWc8Gfcx37P1cu2LzzEkS+XVn9F
ycoIviL3E0rA0wVW9jcqsSPfLgrfCZAN91J/m3VB5St7MHdpI3U78PdTDwwoQ0Mb
p/SIdeqr0wRXR866FNmI/lW+Qgixo9B+wMJ7Ty2ndCh46F243QX2opdtX5WxPXKw
5zyKkDVEyLvWGBYaRo5q4tJcFmJ42JqJmgcRUH9CrjBM2AdW4ZL9i8jJeTIMnfuq
3FAlzTqubv7s2i0qeaLJeUa0lGQHUVYSqDomKB7D8I/pCp5G9x4HW5kqMuXUKdHp
aBvnPPVUtlPQl+GWinMA+InvDqt22uH8rP8uI/dDRh+njZUIcPZqW5tvLinWrKgK
hMIdFwa4m7E+uZ3lzNpD99GXekuwnREQkOD9W053dnBF+zyjeXOiD82q2/Ne3TbS
7YxtpuqRQJCKxcosPa7oBHoPujwCIWQuq1VktjYiIOK1jYYoOkhUvsCuXH91Kraz
F0lxl7ACP+4tCXVYEHQkR/L0BDjfixfQKMprJsY6QNHU1LQ+OdGBRInxA6/l0XrR
dmEAJ/T3VjObGMp1HI4+HZB//Hd/ePAGR8QDbvjpFFzJD3mdOOfMv/YXzTEFFswF
aFphahrZ13iy6iqxnrJ924+PP/IJoiKV0+sA9wXDPx+almd2uIL1Q1uIwzIxqYQ+
wth1LFkxwUMbY5Y+kQe523AQIsJtZOJWE29tR1K+4V5v9yBgM+j9AlYvzThXg3s8
yriiQBs8m/kRlj+vYiki/pjglKoSgOeBA7umLm5GdHZG974xPwjvYXg7UjCQ6XIg
g2J+EnwQz7A2HBQqhPXEln7bKTP3OIddzr7xe16RYcdfRnrpeqAlfdYvabmy8a57
zPBwfTXANEAwTDEBAY2Pd1jtjNvNyDehWYh3mSIklk4nIVTLzOdpwXUbAaJ2lkmM
a19m9BHoWw7dAzmYO7g0TrUGNgp/luMfIc9S9wqic0KnqdN6zHAxKtLHqwPryrNA
W/3b3vxyk4HX/lktWnyahGCxMYe5jqtEW1AijniS8k8QgG1uEzSZECw3iIfuD3WL
bXI8a4cwdFvXGxUn3beMFYbcMmDsyJuZwB16q4wUKrB3S+ZnN4noiH++aBG07kYt
U40JqEwu9crL2E3FAD4CblXoeq+FvUOpXUGXqxR4emzFr6uVC5gX3W4exLbPeKnn
wF4rNFLyLKyif37jww4YdmkffbZlVr2RBx2xx/5OrvMgVm2q30KAyuFGitYDZLVp
FpKKmbxnBL7ARVQr8SsI2dE3GuWF5f0l+q5npEBUnd31nFguX88sryLqZniGF0ag
qx0Vhr3P65KmiXRClX8I/Uh51l7nYoW0NXTQa4IBXOjPaumThXofpZnv+BMw1+Bd
YVWXRCqj54kGWKHK2tt3BmDQOvzxjbaX5Zu8QOoDz2piTlLnn8/2x4cKEAleFf9f
FIEDYQCUOHEvSVetnIVM/v2p2QEHPTp8TjEnk1TCaGdaFNMWwFMRlAsGo60inL1C
VaZKj1kZeXKWdZtjCjfdSccWyVZwmBvzk51FUUbqPiaeOiLea1yZBES068m0lyFx
qjWcjeH+mc4IBlCVpE2GhVBpZJsuQsK3kgkN6zGEWIZRz1T6uh3X9S4NhxEjBvaN
9jf+OGS0E7eOlL7OGztVDsN+FBHBdS/m0zcnzeheB+4oxZzFibwK2riOmVrbni/b
ESlrZyjTS5QTH5k2R7L91uwEeSzfuvZpG2RKN0gsva3z4QiPFcO9DgtP2mptocW2
SXDcy0ii3v7MSyihmHPyGUEHv1LoXs1UExcRgG2eN9GLSgp1fTWLxiXTKGp0cN1y
GgR4ZZ6g+hP7ApKhBvSfbpbaHGCYIw5CzHNbcsTs1SQbrk4SAopGCkjJMFKCiKwQ
esrCu8F+fGn58k8rZ2LmxCP3k7ev7QWP1aMF7MWFnDMrR25nQFEvJRa06JC7O1pK
3/jND4mHrLwLy7kUV6chCrKRH+Ah5Y9QF5kGfpkEBfzli0m/gNmu86WqWXhxzeUy
NJtSSTTZEI5TGLCLo+nvlaSxyFsIqbtNk6DJFjyOMjClkG2x4ZJj8cfitjhKMpRu
3Y5cBaIm10gtkruqboafvDjqgVG4px8ciIYQJDnKHIxnqVfhvLEYqON3U/HPW3X8
/z03cP0jMxYRRuTh/2S5DNUTGpZhBz3fMKCfzhmZ5Neg2Uxcxepmg7KczpixOA5j
k8pQxKHBjjNOj1yjHGYPQgGzs3GbkUMJ57PJ0W+I1sy5nu3OgDKt7RqjxO8fVhqE
PwzgYngeJ7JvAXk6fEpOe94xxLz/GN6m7w3AAunxlv2JLpnogIuB924jYl3Y6XXD
mzosrN5hldpMKX/Hu2ReI1mlZRwDzxUMpJxM/y96gWjWUv3quG+AOFY9e9GCQ5QD
D/1Su/LVFaQZ85C9/QfML0vILnflpM5J6ej3O8DPJrNGTJsfvLWuVWRfYJKtjgsL
8Orvby+8knKabJoOVvL2DurJpbqsCJVUGYzb0vzB9TVmISjHP4o8x4p7LCHvFjiZ
5GjHwnSSIx91g1C/JqNe2o14vefyVTOYj3zbzonP4xSkX2Ok7dgmi4F9FfILEKeM
4f8n6Bbw+wIq+98uVeqj9orVMP/C4ykac/anUL/tTm5oz57lFBjVmBREPBoodir3
/yoy3pN+pa3LU4zaRwW/vr1KAD07Y5CuoeoyfI6gfrIPJ7VhlGk3ebkYD3/7uDlG
t3aAf6Y8EDfA9EBHc98WH0oJrJIflxx3htFOkQBQG8ACw0eRg4akvk68NpL39P8c
ZQzvZAR47FDA8hadGTtquprkL+RGBRqh9ujuI+RVB+dwRk6KwclQNlB865rPK8Qk
T0rGFIHBPpUifyMqxm1ma5K4k+OACJufBdDSFKcjYjBfhPYOg91l9ms5wEaZ0BNi
3aMFKZfk1gczLT7rEnuBD4xYLQWpWSI5HgOeYyNwy27QihyO+j0ruto0borOaz9p
2zm5+TO9X/gfhDNm38Yk+gaP1pYFDIWLGe27yFgupfQ1/27qQfPq4KthBGFPFjMu
E7AEDd53/Lq0+dGmsZJd1ZIUWs7GLK2wpoL+VlCQEwDcQHMfjbiEJ76i/flbavCC
K7ci9nxDb56nlWqNJ8NWra8W+z8LfkWHmMR6FNaxNFoi//0QBwTY38hXkMnEx7bK
TL6tdjytgbPIk3WSkGTcT99qUOcNJjlWJzniqmlIsXxU60UziUEdpXkeAC18Pphh
IpHDBnRSdzDHRvo7BrY6urFBe4R22dx4iSXBDg8UoOZh+53Va8GD6oRoC5hIURmE
//8kW9sojRXXlWDdz9jQAmcbHCkAd6Qy2KWmjGlvsguDuKCjDPh6aWJxj2p2ft/N
CKRNBdkZYdLKis7CkPteolPstjZVpkFwGIsyUy6WtC7+twUYG+cLWE1aUKWaBrv1
gw9WQDm8vCk0tcwzHfE0vRqRrYd3VcDVeGBp4jLj6nuumbLFft96JTri2XESuB98
RncB6KjsOnLSGX5kwnew8TnzKgiF2l+3R+KFqTUoAdrc+S2Xw22oNN/5Mr8LjtJO
3KhgJ6GIujbq8CDAG+glayNq73/Jud9zZKksAo8vSakepR655FT7/lHTIE5Ypt5b
Rc3jQul0fECqg5sCVoS5cIDNmmJ2qERvoPVwtVMdBZFsZjbzRw7cxalTm9zFZgmu
trpj6IFfyxDCdS3QQngWujE+Pz4Y2CsOHDkZT9iA87e+mG0mtcuoff9mOmxsv1Yw
J1rWM3wd2mdeTB2/eRkdALOmp9DJN05TOjZ8kFhn0Z+ed84Fg3HOcjN/A27tE5HC
jkQlJZwS1OurDgLvyNh0JuUnEvnqk+RLm/eumIoDdGt2bYsrf+BgmFKCiugIrkCs
Ad/k4SRQE/dyowBpGPLcrr77fTK8Ix4KjJrhInUgy7/SYuLjCNQZph98xVJpbNyf
LQEUhYX3uBe0TyhKKTfV9RgjppXOTbB++zNF6CYAgO7IKzAhUxLAxq0Wv6dtdHqq
6ikhixtncSvYZ7ATIt8F6/La3gpqGcWDQUPtGHQ3NQ4BLXDjdCltOB2fTkqIVLN4
6N9aryr2O1BPAyE3DfDoUvtT1pFSf235JUKLuRrjUfGM60h7Hkdq6y8s/4Rqo+c+
Q8AOgUTTsl+s4JqE+uLpjQxaFpdE9h7uiAilWVGyV5PStgTAjzM4ERUrbT1mqBgm
BHNvGWBlEDcUBNBpGG6YUr9C63+iyNDzOJOVjGmmOeROUprNv0/kquhw1zuY+hNZ
GGHJvsHqWIGylztLachV4PvVyXrfDaJvsf+vSBJhQvYtEesygZH+x9R2YTawmgaW
Fv9Cr6tWfsomMApWj1+9Rvnl7jQbZe1z2K80eGdS6ErA7uBeaEB8YRmWO0swK9in
3LDpBRSPpwE+XBtOAhVF8yAF93CTLl/YQX3PYc7TMTkQ992/EM1lLXC3L2no2oxu
ZgoF3IUrpOT5zUu1WoeUajWNRozfWXxL1KKlBFV2ZtS21gvnyeZtPGqbx0BPgm3i
edbLVOkWRbIbtmTE5obgAdhr0foMT4M2zbtW2UZB5nzBvGsFDh5KVGFoC3JOHt4O
a7WSYBSaZMADqqAXa7BMZR7oYn45dqInzoDqq1GVJHYEvanf25UBpXQNLKrI/oKL
1DWrIOwwsqNHkRFW+KWV9QIIiKP1FQdaYZVAoYm2XgEXtVshzWN8M3gkRWU7q4/i
1CFsI0rI0ApB2rn22H4PYEc/lanSsvGjuuLncjRHeawhHpVlHwAFaKb0V5atGuvD
H6mECGzvKBF4H411xaf1wX3CEL70MM9/vxGFfBUEwaVcEWB5ittPgqR2Dhqa697L
TBxqikOdM2gt0ZtIEy/zYILZQ113U78pf61rkk4JU7E4Attmn2uJstWMBZ16gCUR
5gdz8f9SU3p95Vv4Mp9MYohVe8T3WdFmJa9T50ggFYEonv9y7xieym0++0rQqcpp
oOqTUSFFek2bLR/TPTNnc6WNLGeMNl5smirZ4zjKF9BmzpZxhj6ppk8YEdoouikf
MHWFRl3JxIh31gvVQIIvJBuFavtuBoExptYUV9l5SXbkr4a/BHkJBZHXPABwKNJY
7M2aRPt9Gl9bYmk6KA3gdwtg5mWnxyUmWqwQj9mysTjEcX6fqib3nIHoeSJrECcF
+Wd7VDQgq0tGOk4mdP6kDisqNEkggxLWchWCjMqg74rvWcuQkQPVS4WPf42CuXRh
wL5tK891vJ4XWWl6BY9pyIRfda73hc0wB/MidRkClPpGaQvamrYMJsrmsb1SMH98
79irc+yaWPlw0yvrYLB0AoUiBrZp91R/YFfp0kkOSlMN5iBvpxsXNnXnJFzzOHsc
CwGeZwNyZ50W0tDt4rVjrWMz0/ATyzzwr7icaYmmgrLjvjeY+urhVa7Ee8csH5W2
KLM7g/ZsfDDoEO6iaHdJdQgEpLo8JTy0UFlZclp12jR7+P0/C6NFUkwJvQgS0NDa
0kGyM2plqWBWqQpjKEbwD/z04GS2sjx4ovXRFS+lhmqCYHOSs0eVSIBumA4BJse6
CkkhwDDeekR2NrMc2MSgFdP6J9cJOCJ/G8lQ4eM8uKjS8gx3hqdzv7nykTilMnyq
m+I8PuJgo/8jPZndgvi0FViESyTRjPIFTehLfm9OxOtioiGHO2FGiD3DYjxdn6sF
4uSonvb2VcFeGzuV4m59ASaFieWkMYL+jiBd6Gh+dvNwpBLMncGWGWphOvdYVglM
5nyPcaYONSTFjihQjUR0i/sZvFCOACXS8QckQNNu6Un8KCZWcKiiEey3i1j84EVA
zgqv/iwkjeSzJJjwxRUbzDxnGkLmBZJeROL9JWMgoyJQ1gQKZF2atQ3DMNbdl1J6
44mMZt4IkX/miEdpiGMtCBdu2+Uw0Hl3Tb+I8mEU4fOm5ko4QVLcTWXn64Sb2do/
SKRYTWy8KwkITeCm238+NflBa6Jorxlj3oTQKfxmLZbVf2J4v8E7cl0JzqAOI5do
ujq4MA8/cjAJXUxrcEj8UbcbkB6UkWpXH7yOpzoOic18jeXmVg5t6fPNRhVuJf3w
d6KYT3NEqqrWd1xCGT31ev0Z8fanGLWdOFAUaJFYnqXKaU3htzAzcIBc3kyjSr4e
eKLKuHdE25N6a7S9BKXab91MtCx54XOP2oRpWGoZz9ww79sPcVMxojwhdiWFsGAh
6k7iaqw/yhW/n22XOaA9iVkzPXCOBSdzMd0ICZ6+Rd9t3JFBRNvcz+HUTKTEKewU
4QBpTV4mI/KK8aROcqSiGE/CGM1OX1RaLHpK10yhX68xyiNTDfo2dVtrTY6Wp+LU
K6fJ3RmFH7woCGJzCy2kvpogpq8FyHIbrAVYqN5NFnhh3mZFmMhFwMTwdXOKk/hb
IMAvcWSESsshU6EmJHlpF3SpwUVYKco9bdoufLxSFhd61l2bm1K6S54hl6u8aHI7
jc1Z5rxfbec3aRJMlfkPwD2CWLLrYJGn7RGW0A0gDY6f4R18lG1fT5jk4SBls4s7
LxLac9Bdb/Kvwn/F7/z/MQ+/wLcCYGMZ1Lk6ZolITsPReORhx9ZJBD+ZhY/JjVJo
oSPyHmLYKZ/++KJ0hqWlbmAX60gVv9Ln+djI80lTYODl8iFODIVGGPzD+JAoJxEL
/cU0m/IH53w8wQXYdelkCmwlN33EvdyOT3VXAamYkKoE2yaxbiDqQ5APsT6BZ8z+
dBHVDVKRANcOzRG6GV9MtyWMZ8koCfpgCOpBa5wkzM048eSAeh5Ey5t1FiQ0p4EW
MYyVOkqYNYuM71SIHqnq7qfMVNYVpoi+g5fuSkMs2rIezSlPshiy+o22h5SEMazp
ISDCmFlYv3afS6ZQwRmEUr23rY3WuRBjAhFSBBkAIFKhB56UhfZ+uuUxPp+FdxRq
ZuXetuGTMZjDSVM3KYGEa0m84FfoRpupjUMOvLg4mTzTbg8hoIIhBc4koHiPzyL5
XdzkqMFawQoUd0n8USCkSqwIcHnp5U0Sf8zy6vm9Tt0pfpG2rTG0UpURL/PsuvRV
hkzZ/Pwf/BSm4gZiFVqA6bDlmfuiqFCs3REc6lWB2y9fbAhIEhtJWva8F2i2iMsC
q3fW+3DQtxXpBKVYx/iPmbOtjFRgZ7og87NMprPtHqi/iDXnnhfeGSe/y0MA055n
RbLIPPmHshNrDNPNMz221aDH/DSvEn3cVNZa/FHQYjCrQ7RKioLTjz/FbqagmGJ3
YI4fPMSJSkPUcMH+HvJOOmi8Z1PuxkwJ27U4NAFiolgWlwZOJlPQj9fHXMqv8FYC
xLhvamHCn260cXafpaauE/HVxLsEiEBInlnJonx/rKdetPvCuM32ZAVwd5FE27LT
qLlTtMkrpebUw0z5V81uA8lY3Vu1VdyTbIAMuV/qwGH8tz2XXNoJLoxmcHHaT8ug
dmC9hUeVbS+Ors1pSmdtOJ/At79vC/eTq1X6i4a3EduAvbpWWh98rv4QCNZzQqCF
Owqf0mZ/n5Lt5OsT1nPt+X4ORUn/DtLpGiFtaq7dYhffEBXmW6hkUtkStpHghgD3
RtUf3boP/kqv5wyQa/z+CqLFSLw2eXnfcgvt5ebjJ6ApU/TnSA8som+uA1WCNF1M
VkoZZCTojNTVCAbBFlvqlrEkMM7sGa4TzCUPSWWjEpIQXUHlmh+O/RF3pLBHcMeC
D9dhacn5QJyCydoG4Y5QQwWu2Xox7h4B80I13L9PstWYg2TMg/sbF2xAO8T0/uuz
BYNwEA16mqkRvR04/NJrClUTXGyIu0oBlwCT4daufmr4AhYaVROiF7JO8+DC2lBR
owUWqBlhVY6IUlpdQYpV9jOCwnZ4tfwvSmR5owHn9Tvt2+OiS+FvwE1NmwmfUTuu
adZ3eeNB7jeydvWyLiZWJQv3CzoGvJFjrlwkBPqtmmWPOeiVzeHPiIQDCCCyNnz5
W8JbR1ErdIxUKsLVrtF8bm5EjbwUU79is8Jj4S1B0clXR8f/+cMVlHqO60F3r1BO
d0mPtcv8OofUNphdnxlSO/cOKTyENg+7vQ/hLo662Mf8xofd4oIbsTAXRxNL+Mmb
s5SOOJ045xqxY8mXEuO9xwGD+/zlGdSrcsesNXF9+oj7Y0kE8E3CKXZgcnWFgrKT
zxvn8CCe8bkyXBYw1kCR4txfOds62FWdT2K0efxkrx8K7ziIwR0jkJm4tbKdAlLj
GJoNskhdwh07SbIQ6NQ5nj3iadCe9saTtXi1PwYzMDiFFcDJlJdIpaNGG8gYLwx/
jhQPbTaaesunPpJJf/19rTdwUAJdM2/wobKNO2QWRsER77dmZZ8t3KxfquuRJMYK
lFchgzvJmQtN2sU1t9uwwV5hChn1UqOh3FpNJtXZzprKeDAs9r89QLY5IkR1jZ2M
H8635ma0jumpcNEROJxC/m5XRGF7lMky4IGN0+FPS/KRn15mXUjDDsK/F9Iz8GOv
2V2QknzcvdRM9qzFkbIhHmtts0obywHbf2TPSlf7i/4wItbOrothikWH7RcW9cvn
asdHfF0sxwCf0G5dOENQPvXDjBkxMn8afK+ZxiQT4B/QY1kQ5D3jI1F+46P/6vxl
zL+V0v8CMW0iwsACwxbHZovjZxWFYBF8MIvaIsi0hPK/JXpm7qZL00S4ApPJE69I
eedGUIGYDB7trGJQKvbIcX5tfky6pnXBdi/e/kz7k133uP8fehuhx7HGUOcAs8d/
vHBsZunjdpw+2TQnjfB1unWXjnwSSc/nCnoHHUPYWXW/l4lBwrswxIw1wXmHXGof
3pjKl7aSPrfAoDnTE9v3n+5FFdtrXfwont/VajDZ/RhSOOjK4W5UDQtl4KXkCd1s
5VAJMtGKFboHan88GnG3LV2UldEhGyrqRuavrLseumL22be2CMiCFwexFp8hZaC3
vJTPZQrPNJ1aj9AWXaELJFNfvutc45Xd9Z0IVma/44iCxsW0wSdp7uXx2+kjdmfH
4rZOE3enE78cEGoquiM+D4KiqaY94Br9Wa3BkFUmdTmqjkmdBEqW0YhgZtKNR+Kf
XzXNhYVuGeO58ZE7o3wwowJMCKukflYaFzrrV1iyhsYPYL34h/h21BaI1jqKpxyv
YnC4sTj1W3BN7O0K6zYvkJF1nk3x22fmISHiqzzceciWPmcdq37maOrGMy2W6FRq
v+JhzJDMHuvDAVkWBMPOv5ZGsQpf5YDHTeNmfCfk4Lo4RNFVQl5m+ayi7krjwBTy
AslzxGhlWnyWTrsZeIHTVvxVYzQGBe7MfPpIBLBCWQPRm9HUeSfwBNOBFZfODoa8
z47B35p+7exQ4XXgIt1AnJsyhciuzDrGKrdTs25BGv2vSLqflalBS5ZA9QRZKYwJ
NKXRbWBfpCJvtH4PAgjpig+k5satzQCHf0HsNq0+av/ImH7oXQDcoDtGMZ6qlg4M
rvVwC1QNEwQI/h6F1viTmOuEGKh2Rq1pSiiH6K1BHi0e9JtWX/BDJsMF0c5GbF9o
4DoQlurq8gziVRYq1a47Q8M1O9xXXSVn97WnI1PkiIpou6/Vd/eiLv7HeifjqzYg
OowlaRtvKFGOOaEKjronylObQS/OA9h5TeW6oH7qwnnOS24Pkp6EvWNtJhkQ2mOH
o9REbNgpKYSDV9dvmw8a22P/Ivzx21JHXTw9r/lXySr3CN3hZw/gTR0SPHkGHMgT
FfvOVS0I8OnAIz0Jl4124W6aS7r0/disU1eczr/FvsPeXF1nZZK3ccEoxtqSdiaQ
tCDHWAm2esx1z5zVjfgSAoMTWpwjg4AsspC5D7m3wIEJYQLjs277gBWdkL/HX3Zg
VMS52cEH94n45P8douZUarWOVwMkizDAIZZNIh/ubgjxpc+LuBjL1PiVQMmH2BMo
sn+WYus4oDTCru2k4gyA8r6Da5juMedOJooBvznz96nUITJ8duZeVve6QzWp4OdC
xx8IBM59flpC90MmOTi3/nnNKpzso1CLwgiQQq3OdYNgrcSn942mskDixt17qVP+
xrknrT+mX0wt4oFHcr0UtI5PbwBda0dRP7zhzdPBNOQM7fSC/mQ0gPobYumvjYWP
5/KmbGVqdvXU9gLBsLEoqAwJYY/coLqtcauf891fhG/8rfEpwxZEmNzascjDaCa3
QL2hkoyFzViNwYXbxfQHFYd0lRxZgIzUAifapRSBOLjCu9cY3fvdL37n7ImAxZFg
RZ2y/UUECXBvsXrvD4bdkPcasoMNbRZDw+xK1pZ6vA53U+deC6i7iT0KiWUsJZxO
d0zslpIvx8jMShfmLJYQt9QH45Fa3CYjEIuOrE90nZy7Jb/CVKc3Utox1sl+jjbX
qIbGOX42VHi41C892g7yBxLgQHr//v6JzfWtxnnXpjXIatNoKha+/Lni9ifUSSdQ
x/mg+uKhCVF0+ZaZu5auDJOEpizV31l8cgLTxAHIACFNWI8WyXvO8HxgOJeOA/Uy
MJVCLro6D14+RaUMh8ux0RahBb0wOOFg6nwlfUS3lO/RoVJl8tgSN+vAVlOvbPyb
W4tzb3Vllf2zEnBxDvTNQbYFCK0Fth2lSSizCQDSCay7e0MAPAVm1e7ST5C6pmeY
tiGEWW88KXyp2RLbXHgvDCYtpAk8liYegWI1fZu5Mbkc3igh2XQ/IquPXdxV7X3q
+08Lqcdu4JrZKI5blLtJfPiW5tbVmQWDcKwPHluEIOP9ZFcbosXhhzcxCi76mqeR
7kC2pknQV64ikieEROG1CQTDhEnakkadIpjR/bcjS7lD39knwP1/HkGlsmnIrI1z
f7n3tcO2HExuQ/bJfZn4kEDNCLoZNeI07jHhU82vxO0UVSS/CGTBOeA7RnPJGX6Y
l1L4tVb45vsy2d2ovCdKg+JuXsfInkeum3YAjUyJMQDirKywOMms8xPTcHq3IG2F
eXc0w9l1yuO2SyDHmBmjJn5n1vt/+dQpwVQJfxQJf8QUE8kI2vpqn+j68j+G1ZQF
mNkxk20lQidgfThtVaSSp9YdShpUWC3hrQ4RyHuuLjQWvsitEHuHJNtr378RlvaX
ytAvJhZmED//oN11C8TpQRO4fK0oIU/kD00WQ+rydGQ5DWFfh/PS203ZR2i+SYFr
LzOWf0vqaISAenAaVs81a81IaMdrl2qmslAezeorf9Hy0k93LSQOHyYoe3q9vfyh
byuAxZVepwCrYula19n6AnG8AnybmmjlADhIVjKKRYIb01eKJRhFMObAkz275Y/5
mqpcm+DUHytWHdlJsBW97W3R6si+iBSTqc4fEDGu5oQyvyKDdGdPi8/OR4E+W2U5
Qf48reFILgm6qhY6Q1KW2Ez9XG96ziaIt+IAQBNK+VM0O/er/8fzVvwSb8hALmbh
Y9SUquzQiW4nZHG+NnD7nisrHQggXyMfJEfIR8v7czYIYjXQByOcMXx/qYfl6wl4
N2PVXwe3Cju+dLepGwjrP6V/RbUO8xGkF7PnEIf/3ZyYqP86gisttfIA5+2JsCKr
Mxa9cvGI9z+trajiZ8Z0Vq1CFs+B6keJEYe+Hm/9UgpOfetEtGp94CkXb3t5pdr4
M+yrzlJx340478NUAx/7L3GzNW6fY9833LDrTZr6Ceq3F7cMPZCfIDtvKF422a8O
PH/06L8tV/fv8LVM0cFsdyAmc995vId6Cjn+8foXPqIT2BvJulicVSHbrx0oaC1N
GSq84Sr0/h46DtQ2Y7pay54QgVKxq8vQ7yKSwvd2UeptJW5GFAZn7EfBMEwjBVxV
tIUJ6T1GtdbNLhtoxo4Ed653Mwb6hqyXi2JB/rs+HqhxyKdwykE/oth1ANSM9mz6
b8ba6O2oE/NQ75OngBzhCXYmtahCPXVGCC46rO2rB8IGlzepds5Hm4SIc00PhuzJ
CHNm9MsLdrh/6fsq8eqmzDlunltu6pWzpr3oqj7O9ZgKIDLrPXU5llmJU7Su65rx
nQ9fFRBvcVd/HA8EGn25b3HsSnGQTRNy0y+28/2wo3+0Jw1giz4K3QTSBej0OHCq
/V6Hj92oHJ3S9WVLNz4P/UgKuDoUzxWZoAyteDiUdVVOVsUpPmcLVJMXEQF1Rr3m
W/p7CYTqVsYsHlkTNgM/38qKTarYJXFq/HhZc5ho5KhSXcYy3idC8XM5boN5bOpr
brut4REldPqWHp3gbZqUGGj1rk4KjQoWHEl5dFwDQLn7vwRSE7r+f4uANCt9B1/U
FfPoPBVOHJ4DgAUHW1sm+3k5ofagDaG81l6NVQiRXB6pMBjOVoOMp16o5GCvsedZ
flnLsmWKzWwbOYYwXJdZG+e72IZflL2Cu8ux3MvYqGXnQOWj//qn7KLcd9Z76Q4O
tLn1X06rjvdcDkunvm4k+cWY6E5hFVPBoJHWg6ROzxta7Kid1FYcpzrCLK/qQ2ID
fgmcnZdJ45fl2rgQN26kVJ7W/VTKkQvxxxE1SeQ6LOYjUF+ETmDviv7P6xGPbwVA
sQ7rnRBgY2nJBGHKRk+w7WJIY5ah/JwAeQoM62mT0G3p+t+eZESZJBHPCH0Aw2WF
tkxWVSR7LU7uJQ31kGhZOJY3vOpHaMNCiHqMU5PVNkIYHMESAPeytz1oJmI3RwaX
SdoPkpdvwG9o3CHGH+ImvLXrS5E14ZmUI7GHE+xuCCdDZQmJ+DkgEQoA5A5WCRVZ
6JZbUHhxYqwsW2vKRpwcF4Yfi6nnhxjIhJcjd+84B72qHdt7UR27ogGKSkS3/7l+
HfOAtQ4AR3YCifK4E7H3mYykqoifrSJ1ocwq6LPm+/uq05HTuS0wgliYhRIrSfBV
AUIFwbKFx/vpz2aR2htacVgzuLGIWS/nfNyupCq8SRQCUVBvFA7UOmwwoROswvXr
7kQVNFFAmJz7MB/LaVQ65EDz6vNi9+SQJFxa0Pzz9Vuiy8d6+1aZ8Aul2uxTbS6l
6QVbYW/sWJyW1xI15c0UYAs+eRUyP2zRTdyQmzivNujkIevnMyftYmiUf6EduNCb
KuUzHbd9odQery+rQOGJk8S1eDPWn2mqcS+lE/x/LBvVZMn/eUN8IlUxdoyQI1Jw
2UrHMnP66hm/b4NQtXndtym0wLyMFfDHgaidlHR+YynHndI8t07c9BvKAEXlYtmU
wSdmx+L1NVIxCHZ+g4cDNnUUPPfKN6jZarq+e2tZD0G7zwG99cLNRJjGovNFsx09
7tQ/ZBzuYS63yl2c5dO91mAVpZxK5pbC7XWp2dcKy4gvhtIGVAhBhNVjMUb8c/5G
jKbixkNFWdT8UlG08Vo9NNt9lrNExsJ7+6XjqFbBvj4PRPTTIyR8eJcAYLYjP5qY
LUDF0ojaWE/C/iK3cB4RwYV8twGm4Bn98sE1rNVdW3uqsBAD1Y8F5oXqK29yFOMg
piQEfOZoNLplMhxoB7w//ztEvuoDde4ymiHvF07Npwbq6RFinfFbc1Y9JBwHIjat
n5l+WBTEhDfqjH5+mkEXGTDXGS3i9qHdELc59t9RN2O1aSoloFmTQrdgi/IDTh4b
aQ0MLskWJHmVoDfsYVZXY5yGmUdD3m1IOY/HYsFIIZRvD5Z992O6dQx5P+hgz2kw
56iw+hESP2lLus5RBl4AU4rw73g3+I8jsa/LGK4rlI75WQgUoMguwdtMbhut1BjU
fVeQmlUNC1TUnaWzHID2dCUkCMWdPdA8Nmb4T2uWJuPtmIKGepmc0ljbInJKiktD
GasL89IzbOYkuKLvO6Q2Md+Ppeofs9SsF0/OFhciDvtZliovOunys6984cnXQ7z6
/da7n2nOTIV64EzcM1eIKzsdzPqxIHqFJ4sSE6I+Uy6OQWr0Ze1Fm39YE648QVQK
cs++8074yqswxgd2bQnn3dckf2/xyhB6AUy2M1njry3ExAKh/qq+tKdtJZ1KdP72
q5HHKIB2V81UDX3Y9klg/rMkGe22AqGls/r4hDY9IzRPU9gELwTpPJNwl+kz+4yH
JwPlJcbQMpsasHtpf6Qv5s1dsdHzERC267Me9yEvSPc5PEb+HHeXXafVwX0B5l4b
UWOdka00vK+128pKUQQ9nRtkTsVj+UI2iz6oqLSbr8htdjtLEqvHVaB2DvoXrp54
tWyfxjsDb4N2iV5pQ5JUrIuJt8RbXR43AKN2WUA1op9ZyHIloLGhpO8D+AcP+kPS
Qy8VDVLmuXkfnfNff++YpHpQG1oxaOinm+jJ+MBgP03cdiO912ehJdUZTCnKAr8W
UzdZ1IN+cY+FP2+nbFAv4ejj7F3oUS/gnhH8HF+IQORt2UtqHCXv81fVERV8Fvgm
QiaZ7Mx4kYKzJ1HG2djzklJt/SOY45hftR9VMI127z1m2OaZtwxNzBXXzvQ18LTA
2GsgqO1i03E83mFdf12rHVueO4ZkaclYMPY3fOqh1LY5PkeqQEZ1NPjZeQQO6h01
IILCdNXO6d7i9WdHVKzrXNGN0T518DN4/DuDyyMVjUS/qSNz8bVWjy+molL9Xj9O
O4MOdSA7y6rfttcwrvusDQ6AfystNhd8i43yO1nHk74607bTZ3g8GeCpnRLDOM2U
fOpYQhtmiJw8MdpaFHtwYe3GQc5oU9CG2hTIm37sN62Ekd2X8UhBkLzfrQifAdO4
TnKbootJSddlppD2WFzSiP4X2oN6GaOgJ2LnonWfmE7L+vLSQfnbvEDXMAYH8ZeJ
WSinbi8smoerrJBuHok22rYkacQ00wT6Yn9f9HDnedKaTXKmS5W1zu+8f/I6NsMi
TuNl6tXk61SKWCDWLqpyCjvo88M7ldU17qepTs+sy5tXoVWXXc0CZUxKwQ6ZqyUx
PTwVtxK4NRyAlNHqXgKcwVU/aECgKt9NvABqUv3RYWluXeYe3bGnB8jzUIP7QFKv
qVU+fg4GM3Li8dTLN9Q9/LjXDgD1mjEVg6IofmL41fDVk1SXWOZljERcuLPx7Xnv
AzHgwVNwxM4tzrsSOtx5QM/xhF5jJE2a4b1VX+9ithQJ+V1uBmQ1UR40b398sOhD
IU/doJZ08hNtmhXK6uMeff1GknAZHJ6hmm1I0DSfv2tqZdkfyUBTw9BZsn9ZzzPX
eJlSVKlOjX2u9q1W6CidK+BV60GrKWIf/NAi9T7TVveWWpAp9AczPeaSyE0/ZBKO
GL1YbT/YFnfN7+HsVjcq7dzG8+DZLykrAT04oI0iv1U7sW8e21UaSidA36DLit2O
ElTOLqWZP+PVvGfdX/Ql3QbIW7Iww+w5rA6EMWtDcymQocNno0dUFKb1Q6VwAJ7y
Tz7m75qobhAOec83ot9WzryMa/V5XbPr6pAaM0FWLlVrn5lOvz0vV/RCi2Oa97fF
0yPrUQl3ym27tZkJoroCBKZtS0rbNdN9+KtxuSH+gsDIai2816ptszP0q+Rx6lTP
vpRtXR14gm5D+dzy64Ti2ZpJ3gzmHWOvgXrdqWUYWlwVbssdHjpRdeBTwitxG2TL
sqvJqDljUS+TBLvnFjrYhqHnFFzV72ekWICaR10feO+4BYe6oJfdQWocbb/T3ltd
5J99fBNxp7AvpXJk7qc5AALlrAyPzv8IqO0rl/V5Jktvi5w3v8Nvhmr6jABgQ4UQ
6lSK7EJoxrFC+gFPwbfzyx+i0o2Jco4GOpvkb77MK+vZgGy1bxYRfxwkGuIS0yoR
YCjaygzYfAqwCHJ0rdcbIptIteWGKByl+3IZRh/gU9C79S4CLpwsd65UVr8Ke271
sHs+/iKYomM1hKMdE6jLgMKUzJ9kPaz3/ljueRpKA4UnOsSHmt9OKk76KmezTAL1
nugX3pYtQmwSxyqZ2ioHLpEPz4OR8TtjDRof3I9t2bv3aabpwTjPWtB7UhTsNQI+
gudCztd84GO/L0DquSbh0h3hO8f/rWSuKZIPvE/FUPSUqKjJLXlL9Z/UA4caNkrh
Y+/m4mcaWmMsSQMSYi5OiIwTlZSmHJrfuCKXhHHFW/1Cg76VfGrXASjYA6+dLDxo
Rd2wvQcmriaE7mW22htwXmEjpgQbeSFYPwQCoptY1iGCiAx6z3MIRxC/5RSUDm3r
pXllQ6vTN5+/Nv8OLI7qRnxteToqJgolZK/zd78P4xUt+qdxKioLQebUbjfz+OLc
/z/znhTwU79FiVBHtB3FYbL3zEqILzHcTjAVAs8yTN607l0n/Pdr+HpY24EVv8gB
9ZCYIc38RvikuKTsjzHETfawg+Mt4Hxt1Zcykyq94mMeIl3bVelZVPRrae1hwPhQ
Lk/NRPyIAYX4TqMdcJ3ve8yGMLV6Un5no0oTy4X2ccDBtGxaYo8nAOJpHxZAb34r
XdFzH/f68HdLZKR0+sphbOu3j1ANnaAgdEjHvlVwlzEantPmGbAlAAlTYw9TENv3
YDccXLS3ExLfccoO6RT9RpD+lknh1uRZgXzQW98em9Osj/QqClQzm6mvOKrZXppL
qFETm3MnW09QCj/csd4CyquHzh+3B+StcetOc8MJ4/+7/BhgyZqmw1EvzV/owvS6
NKLsyhhBRQ2fQ0bsOFtnbmaVJdpUtxO89X/BFTgHRKm7OwMMGfyN8FCIlT3OL4FW
Wxo4hUeNcc1Ef799HsBO4Xtf61tyJ846Ry+E57PB9yvsMS3KM0CJKvtsCZjLC3Ze
mzQ2DHysa96ccMCt0Nt5CEb+M4bjCniuIOavf5IClVwcbdJQHMww53Qai45bvMNx
xtb7zYiUfC0xN8/L0MtmSwk4b52620A5WMlohL7wCBimnejbCEZUtuU3S5el2tK6
gRDiyBSfX+uvmCuXYM95g29aRnnMi+20pT2uaukIJfRGw+Pd3UIqTMQMR9iVX/ar
dnicg/BYKxPE52U67zszw+V1Fi85yO8LPfQauzHLRA21zkz9zPl6EWOzuQE89Eoq
PTr/VIJdTnlqJBvz9giNKrItHtHlGvexIPCDD8bkKLlStkhkeVxHgw7kJq6YYtGw
EIrxUwrmgJfVzEo/xGzzbNVY17s0vkr1zeW9zEnwsd1R3Rg8ppDHrKc87FD+ol9I
Pf60mcAhribpnBv4U9sP+7t6znLGLOXf0WPfEOF2R5yFTPaToR2mrziD52LOWNyY
gjAyW3lcMasE1OYO/uHcz+TO0K10pZ7lYquQ9bTpLjTs+yCbUsry4N0AODF066Ot
PWpv3+LzAOOLrSDllRKxdEnMRwaD+i5L+Ve/LmHSWdrtke7HpHilaIW6lKUvpr5B
kPkAMNFPm+a2csKiSDm3twn2AXRRTNFZSFKqr51TsEQOzMy+qicq+n+cxgO3iXwV
nxIoxO9FRRejiCQ2DnwpYJRRHqekPd3YG1CL20H8BYXV8iqlD6ajnrMiqqFMFOng
B5XKjDa2YEQtmD7eQdG+VoN4n77EdzA9aNMzIk0RxFBq9YFCGZbhXpN7kNqzIqcz
brHcYcwQn5MIfxM7NlyCGr/easLqnVk9r4Ax9X6nsojvdKYggCNH1gN4j0L34IjC
EbpfR8XlMSe5VxvyPcOEFZnvopkC1wqZRvZ4NffkZmr/A69+i9+pi3BTv3zWPCQT
ICiuupUBk6LyVumZKhTbJpnhpr3d9r5u0vkQn6tV80sPReMLXCAdSPRL7lzPzD6o
+S9v8p3tBCzBxcrsvT1D0eIb6vYVOhTiqcz80yY8zQR38S8Te1uhC43gw0nRZ7Pz
4Zq5KhKqaMWzOut2X5bSf5AzAqPEItmc/ob+4ghpKsfiKO3/2htvDH9aWaTp61rw
/tRgD+pfTGrWBpa1482SwGkzp51uUO3i4mzQn9PG4KKKK3zh4G7eGwOq1Eazm4wl
Uv1aZpo402meqezttH56aUJfpn21ZQAaM2YGgTR2dI0353WXoevjhIKuabldBBu0
GcFNyVHhVIOHRzFurC2G75y8dI4FMVDRk4wCj/wg6+GNXf7XNquUbEW7In4JweSu
1VCmPyzCxJmS2BddRHU6/PpAPoFCZD9B6BY6zUC6NXcVAwdkpzOE6FxFwKxg9ouD
Bek3n/OTrVc6TxbOxg0nBTaHXlWA/5LtqKEfox4n2kWNeWeUrO6+FRwwOvCP4GwL
CYplbsfvy0vqxMVyEdwVYnurN9qcN19NS1OFv/f2j3g1MpD/YJkc+fL6xu35ZJUd
cAp/by7+Boqir2A6rxpoqoo1wOhB/I+fYFWEgBWFhdpwhX4jfYYjutDLtlS00zkx
BUV4KUF2Plg32nVI1Ek5QgarV50L4y7gsyfgCBaidu8nstNdVJGBODZLzZottial
5DmP4dGGpZKQrrULL/6OBCYVq8f6LmxQO5ZfYrF/7KYiHyp5Ft0fGOdjEXg2q3wW
JFqphHxibwzqe366bgrBxTvZFuIegW2rqABU7l82zRHQH4hna0g3Bgvg5QdwG/gT
58lkWqbmjjalXnLLilOU2jFwRQbrHAtDxETL4naFIVisd2FcZA8ADF1w5uj/EyNL
JcC27a3LeYffXh7gL1arlCSDE4rrvuKAJpDWsttFqJomP6ApHQfv4Y5/OwBUq0KQ
CMhPGygfuLNzo5/cCrXjG1g8aK0NcD4c/tl6eLDB0MvOx8jPd5RObJ+gu8yX0I5o
sDTXhPuURTWRjUdXLYUUlypX1xMD1Jv8KwyxE48XwVFbhfCdeNLDb3wFVVIYBkbH
SbjAmN9w389rTZayABIVyF6pyhSRumBE+DcSUJGZv6aRAL0Jvxy288hZ5yh0Fqqr
TmfBOA7uEht2ETGibzIXLuTcpq6d8AnCroKXGBlDH7KBCj6Pu+x/OieT7gdIhxjc
hx1YO9hIXBgGU08GNMlg+L7UJXQevm5K5zqe2CM3gbpVE+mk8V/zV9PteQ3UtJp0
hOkY5WV2oSrRlfqg/oL2A3B52JQkKmlzqmGmFRNHRTWlYVIXl74YzzTuNcaP3Xyy
BqwmTZ6Yh4+xwhRiA1nw9FxIKU1j7nXd3KAYkTwvEzNq69c+qJLhJfrmyC0YHyUR
vHdxkGJwsyz5QXt3P/MuwSVoI8zY1vQbV/0aBI6XsLDFwQaqpUVA0wJjVfRxN8YI
cWykri6TGSIEwkSheARQkZ6292X4m0vjaaTrMQicKtBToAeC8oeWil29BWn4B6vE
Gptb+6uXs/p8IUeiEjBBSqismZ0jamHlXV/oMDGcr+YMjlHb8pKGuBqGK2vTSTT9
swoR/x4McgT0zZKLm1sTslU0qU+MN52rCUF+iLi3SY/f8PQEIDoGuK4WFWQjA4Ef
83ZllhmhVS0kgs9uhSwSwLzs7YrGiFuropxWFdiZ0uEvSdfp4BLN9ra50yNGS/DP
xzijwn/kuAu0ybIigj4o4Q7sMf8ubfch1hxmVuGiC5J2Xh614Nuh9NIQzb/NnwYT
Skty3dXNADM/72dG2LMVZEDn4Bb3S+kTUTp0KdRUDHBpKnJH20OS7GNy7CEDVmeg
lc+pOseRkrpwRzrfWaQrv7oZwFCSbnowR3e+0BExIe30GIOWedLVJV98pF0MciMp
Z0mlSbOAtJzaqqd6NyEfovDIu/C5xrH7d6r9gJdlpX7MH3PqjkndqaWVsOz17oNW
XX+BHQkHXCheDkvp2O9OS8UZBuX3j9w7uGzOzxJTRdwwf5sW2kBbw6aNgJ3wQSd1
qD/SyQkouaFXt2QOup7vAoUdd72qhv5qnxyAvaUkeHihf7fchpQjxXoQGH2owGqf
BCTV2Os0oyki9vh/fjA/3uLZ2h2bE+LYxOsNpmuhS2wolkQ3Es8jwbUFo80Me0h/
Fd+XJ863YqjHOT/mIx/O4XNeB3lJypHOOKGv06VdOLSuIDvhCHFtdtcds8np1p7x
wObd59isWHbRotkxP/SINVe+iMFwehGwwP82V10MOji33Nza60ou1pHWoW8kr0Dx
QNHw4pDHp4YBHYDVmbQ8VjC5zIUj3WZizDzLuWBX+kKHV/PDCJQCqw6p/u+mcQeE
u42X/kCjWDT76Jv8hr852VkL7QUmxYE1zL1QMYx3Nr2c+8dkKhVcFVzjqR8w1sw/
Bu5kbFTb1HHv9pS7/XW1r5IH7E6XpfIBg4tq9fnDg/roco0XCw3XXOHvxuYNSBte
FyaTKjkbhc/7OE3BkrbBqdj90wtki4uip7ID1J3tUAK8EzQGqZwT2NKDCcVltjUK
Pmhcn+8zZrhMqF3wmi9wYxSyrszo+DR6+OYY6eDGNRtWOG7bO3TrYeFmjklfFk16
mQwszBKUwUWAXDr2TnoUco3ZRebc9m7L7ont/3s2gy/fz9ts/tCnU1EB/5NtcOJ1
J7ikCWWLJl7D2PA1ObCFTbRczhmsdH/WlHbpgHB2aysQtvALBYKWIrFbfcmIItqK
TpAWxuhhe9AxFgxbqMdQTuE5N/hJE/ebNU8lhwqVRnk1d2CQ1NSkqX6umW7aNq11
sR6xAtRLNACzPQL6LFWOIuW/2kXTIUttZnprTpVIT9CV5mR5jyAo1EFhQOl4/1un
NuII9ypszHN/hkK7bwqBobMmAKt3Jr8KA8uRat6nYoZ5XJJFSucDohxEd0HMf3E9
B2MYwXf+7RnUkuBe3xL1NT4Mtvny9SsAuBfzWD6VZku4dtjyg+cMX/dfNClW6fyp
Clqs1I2SSGF6Gmtv4i22SSzj7almVrhe2sQiLeFXUV58vys1ZVm0uQfqDx1VU/kL
BXs6kyhOaQlJFQe/Wop+mHlC7mkockq0PIHCDjkp5X08NrGYsaUxkUiB8x3/CyrO
JIULfls+QH97QjM1LkEiYrKfCWhaqbGNP8p9tUOu1lyYMT58UTYqM2ELPkqJarxs
jJXGT4uRU6ZC5gKfQfa6BgwNWtjT20aCCm+gEJA+DVIOT+Knsml7w5l5bbMsfK/E
nVxbj2N0o9DX32yqac4AHVqVhFWKRQAJV0RprtfKU3pdRkn7Z1rkl3vW+ZcpD7rk
0NFavJNwIkx3eT8rGM55MaNF8s39cC2kOZE3qw3kAeHQ9CBNZesCA2qSC3Sf9LIK
DEqR6Z/cuVu5R3VW2xLBM1XZGXiT+mcoHd1+BfhKGDb6CQkzf9k+SLmfH8R758qA
wfLZXmerDf63yO8pccpgesWvvRjl+Y6oEIMlbLzOHmJmjyS6QdTlsIc1Y1GIWKQ1
cJPvABRrVZgy4uH0Gmxo79bTITwcmNebUsy8dWYKP8w3m6JUaTd5lRrNKxfvyg1H
VY0E63RhL1T2A29edwPm32M8WdppRhhJ2i1R6//2ieMycl3BR2vsJYZ/cZyZEqTf
+JREzQ7BPCZfcFxz0J7cSeuXG/lUM2+Y1w/FVvrtiII+x7U15oXszINleU3Iq7Mq
ifmFzx7krnmD5X0QQSCtJ5d52bCPYKj209K2pVmkkaBlaZ/3f+F0BT8VYHbOv7GV
TEQ8Mr1j1qgza8A2rD5470ADIb/0qE86iwgvc7FIKX8BAU9YndkUoUtScvaGvEXU
P/7dyioWeS5rSuGsHpG7A56pW/GQ7kL5jhBNcHeAAkoqNytAwjQfvdTnIyiwLcH+
G9GiYtaZv8zhSLiSwlHP2K/v7VpKEZEYUvxyGYQGvJRcEtUan/BHC5pltVL9fEa4
9sBYMhxNkF071ODyVHaTDrbH250Dk8cVgQzZ7YdEttjvxSzpIh9NjXCjyP+YSEzc
Br/AEAMMMBp3tMZBk1rWUcLzRlPV2qA407fTq5XtQrXDeFIHtc6VSpGKiorlBwa6
Bh7f2sdvSrlKZtvPlrWwzP6lAUgAsfoH6NQCVNhJQCkPEdEeoSoON4g3pAs3MFr1
q+yLNA8cJZ15xz2zqtm8QjrBHRRmT1W4gXd5ssgWtUHwXX1BviUWcsNp6RQdIxNN
zNf/K6h8FJLmtDKhuQcPTVe0wacMtTsXm2tGQWQ5CotO9myXcb34gdY1whewpV2k
VmQyxSOzN2Y/6hhp5h8eZi5q/4X+DMyT3liDIoCErDhXitfflSiQBnXbcu3lkdme
8deCjJ+1e2D1CUeLDBONw91jFgq5DejqZO4BefzaIpoOMCLOjjxFEW94tgrPmR85
SRfx71U+65b56OE23KG+4wPJN/FWoGkOJqTb0y+kkZLezjkM9GDpxhw8o8plKPrT
2S7oiu4xtlP45Eu3vsZ6WL/dGMKOT03CggOe62ezI5VIzHED55/yx/IPJ6iKKT+x
06klSc+gLbckCCyln8OBz6ddCfH6FkebX+V6gS7M4Qbi3QvdRVYYLV51cNXQGkho
wTztw7vArYdUFtWayqFctFCfzRuuAMGaDIDl52icBz50trthYbYVW2TfcE9Y/AFG
gLP0qP7NM7EzrLEze82Zm9YRNzFQi6hfWybDsZeTctdY07hNNJyPDqyO0UpdTX6Q
ZcT8qscNIwV99Ef1fkbhsJNDVO9OM0Jnrdz1OWr+2Mf6ivQapiSO1+TaQ1Qy4uc0
W+ZyHJjHQw0HtdnwXUiRQXPifMTS2cGfsMI2RowoqGYovDA3K6qK6YMbuUg+F2pL
sXjA0CPgsIjDSyBSMTPn0P49lAssn2rB95omUU6kp+FV1MWXys84TA7a4MWYoAUP
YUk8ahQpO3iDoT7nEkso/kjKB9knIfy/Ir0lBpOQ/8yMPz9R5HxBl/deNUqonrsT
x9vbXy7glAWlddBUBuU1bQksrpOXjpHuBOJIPTYtd2X9J+X0bTyJip3GEJZygWe4
QoUM2dmaIAmmgHbAW2SW5SJlVfOKj0KIIxAKecsYwQSU1BzaB5ZqSWoY1565qtTo
Ob8jjuRBOk3kfS59BxxuzcWd/CQik+86C+dbZpTD9QIYo9a/ubQeyPJaV+rCWmsF
PrtNLKqUOEQwIMjIQM/jvcnTGx5bVd/7VkJwKulhOB/giYavHxHzmlOfwqPxKhY7
4d3U7skrnGN1nwcQbiWWd5SLOJiHlJ0y/+SggBBdwAfI4uE14IQ0fAv4A+r9kLoA
ZwDURg4VYbwAFGX5cqbONanb6RovUnwMd9ONhUk0qx1u34sK3JbAo1xh/UuU5Xmo
cDEsoJ5Z31HbGyfw2sd6meb1IIVHpJm2A0xo+ks/1MzPFtPB/8jM5PKCSszpyoqM
b6jXVA2WQsILYRveD0rVS5kaLepiUDxYK11UqT9lID4eumTX5w6xV0Y3CV+6Yr0K
/NirEHRJnljsZDlamRE1S7HtNA7jNW4YmySYEh9jcv/sJZ/0JW2YbTp5HVn30tIY
e7tFcVJnaOCZfwJbQfxAlUtTXjb0eDslQ5UFOUQz/kd0JUahXmGWr+idSRGS+LAj
Glt4qb5ZK/IEengWKW3oHVXTnuK5MZRDVrfQV9BbWiApR5fDDfAR7MUaT9xBK2sQ
9vDuTI0TdX/tRIeXe9fHFEIIiJoLZsPWzB5R1V6x6cKP/iokr3Hblv4SEHb0JU7N
5eBTnynT+LC9+vHlDbHCXu1cEcFvZ+wYRqpsKhY1FGDJE6G7k0HrFzNEGdT3z4sg
hfSdMDtWHg7iJg16fcKoOx47jopJ6EbNlfGf6bYf+oBB1aWEt06Qkj99CSuzLnZa
488AC+tqGHb+pr/PKiUo+vQHSgnWHmrQUOxBstjM0BXG2XAUc8OSmej3HUDa3k6N
X1mWYIFUjuTtAZtp8jYJTn/E3RBzMbhXA/JvZFunSeFkhT293l7Jk4msIgAuH4/P
3JD0xILmOiqQ8dJhlir7lNfB03NvGHGpz1lluztCr1tsmfhhGwBxGykoxbsW3dnr
of4w+xN5m9QDQg/+HZRiDQ2mBUF73qGdq9hks0qGaPKuSfYFgBkBkU2Y4NCDquI+
BnzYAmnfwdAp99W79APu/wyojIv56kiHD+9B0Cz896MYT+WgqgViu4wXruqIoPFd
Qlz7C5wLtbWKesSI8yufNHTQn4lV0Ahe7qHaozzUFCSk+wdCOAAdBlsH7WZEiWr3
zW9vcGjW7nizdQovDSM8paQrHAZhft+0McerK90DyZNKDCIEHo7nHVpeURxLN9Ng
LpBEEhGl7CFrTKDccPU9VXZ93ZpSgsRMgMASfGDSrMrExJEiDC5ZJpqf+x3uodPu
IC4GjVmE4FcDsL90Uer8alMOJLMhjoInbOBXU6JsY6xtzlDWkzxJckBuKtWXcJEN
tAGWavYQyxfWMa8kTk3oXtU/m7vbMuw/C3VG2JUZ5enpsG0/hr2z22bWLLJw9gvR
Cpj1RAOuBMEfdIC1D/ycQh+KiN9MtTD2Swp5I8zaA3AyMTEGUAF2ar0KG5eMZpwe
kQ5c/rxtYGY6CalT8qWSVMaEJFh6gVMNYTt4hXQ1pqGc86z78/pdZqt6L0efBO40
Jl3LTfVEp5sQhabJ5EgQrn3Z3ZvOVsNMYVG//KPVAoqmNlbS+A7qkX3KznSpYTmc
IK196PTZJ+SL62F2lcyFIKmiQNRbhDwikQ62n7trZ+jFdPVwqKm1RmCSk7UeNSdx
dxCzFTFRrI7qEW5NeGQh1wGjZLMGJ1OgfCi/AF7pft8WR9nna11CrzJJHYJtJOMJ
f1J9Et984VfTYtSXEQf6fBVXuksz2RLTPYkJS44VDl5MHEWm7Wq/rkR/g12FOl8+
93IQxj16Dt4dU8wH8hT032A7dn1B2TQ4LhZAEUP73w/5RZ48/l7tjkLs6wxY0nct
ij4yeW0urd0zXi8mjfdStx8yWG9yM6xlBNPWI1v+FDJ0pFZ0M2GlZA7ataDECCjh
cD9g2PUbeSDasZwQS4oT8CLBzt9uaZu7sjnErKpfbs2VcLxDEXMZwlII3+IKXcWy
Ek1Fo6WP5kd2g8DGUI+Mx3OfAqOxWbMucZkft5HGKhInoxlFpKVduCkAKHDeODhN
PQhtYjfMIeWfpEAzzT5f761QO+bGY9KsoVvJRasonscfn6yoZXgeAdzcb3Nd9eqX
hfeE4ypafOqLaGvEAL9MpmhdM7dYu0TxTK1Q79Hc8uHScj7F2wqDciYldL6bPndf
hHI+YtAca1ARDodID7+I7AKvXmxxseM7L9li3zE9dLgU3qdUbTYgb1eowGQUTfD4
gpXvFRfsVGSKfAj7y5I53KmNUkvRHa5QtKP/Z4Ukl/SE+nJn+FG0gEQ1BQz6ct05
YHLeOJLx57+awXKIOEVd3FBJiI9Du4PUKVAPzTvS1YqaS85WP/ZJXw+pymmYKEvq
eqqYhyhHLgSXvigi6CNfS8WTVtMTR3lAv5gIF+WNf5XfwFewKG8v6AR2uNIID2dr
ZI4GkbcoWmC+WJhRqOFQVho6DTqa/m8ee25Q0EfkLqm1uskIgd4BIl7tObaz8hlj
UgvEEMEnAUzQoAyb3XI2SaVHQ5s0y184N6ZxOXbU5DVvHcxftK55eVFC8vss3FfJ
ijAeumZs4XW5MVDB4tbcqEFHIPYu5RDwu5sb+Wyphy+lWGH84oEOw0KmQYDKUUb2
Fg194gGJDkwsstltuk2Y9BtVxvOdLCkjg7j9SkZnJpeczKL2MvfevT84m2hnFpQI
FAbanhjzKQgMCQlUVhXfYsDlX/FCR25gK+gQnBfIgTt1+0EHpLvOTmQ0rAHYDXHe
X+IpDzzg6etTcBIELEwGLdsS0S8RwC1sT+PMdItpXBwK6VaSWrXLHRx9bdk3JTpD
LuAxtlqY5CDH3WJ+uMvr7bu9DG+J4z7UfCyh2HGmo+oP0xZBIk6xqIjvWBW2kXbm
V+VvA22jm+iHqXNKVsXkNn3Xxnw+ri899J89CjbLSmNhiZrj9rx7hfGyr9r5doIs
lK75vKOUZvaycdjp8h9mU7CEL0cZWUuC7sD1nNC7DcFSzUVo7T+2mWJiYEYE1j+D
7pxBfCNS824v/eIc0Z25BzZ6i1CDMzbe98dZASirnvgTuAo0J5YOAGSmMyo8F82P
+FC7pb73ogfz8C8W1Rw2hb+l7R13H+HxwteujMoRcil4J6eItAMrkKWem+BV1GsZ
kJulW4ALBGfD7A3/OYerC7d2tnBYfXbBWjJPYFVgYv1qtdj4o+8eYZwCAUqS5WJU
xIb8abqw5oYoSX0R+FhhRnRDAYPEt04fbK1SAj6dDKh0xm6TXe0AYF2OWqyb8p95
UbOhOA+fo/4ShvY5MzoNtX06hPVVJ0cEqCxzOcyCpPkFgh2ucRwltiugTDWJ/47P
NhH1WIhmvy7ASX2VbhUU0ETCVoIEoNC8O1bP0cA9Xkmd5EyqNpVi128xhMU56TEJ
lneo9qYB2sn8H3gvwELN5TF45N5kmOdpXJMRjeA3HGG7x0wBFpAqDaF2niMGDU89
zGWHabf7bh6rC1PxCJs2ySLMss9dyKVYbazb7f+BpgmRkvVW92ra61Et8P/F8Ggp
h+0avfxhu6wstART2wvVQ83ulmpjK+6vuzXLGUsGqpW5EgamvsnDt98+sY7o0glN
gu6zOPxhge27KXdmpOE6DkTGIEWvaPRxiNZVnG2lpghGaqj/+sChZYO2lc7VXKIG
6ECEKcZqwwtEuLAiYICwRtlV39TikEbHS3hbaDx24u4ejpLdUXneX441bQKDfTJT
x0irjeabkFSbzRfLG25jj8ZPpo9WekYBqa70jXv8KBlurvfllqGvMn1RHMD0O8bh
NFmGO0j8ckVP6a9qgo/i9OsWQ+Lr29to5kDjE2NycFYJ5AUJIwSKLCrQInc2IZZQ
AwN1ZXndELgr/p5sh6jqqgpyEXsf0D7X0L8TSHV1MiaoI82QfD4qXtLwy6+NPFGD
9fF42ERsLCMJM2drQrk7+18+pwMUDTP/AE9hSpubSTI57zPOyXQZySIfnkelvayb
bPPfAwz8zrB4ufx4WPcYZWvFzQ/5UWDviIxNcp7ulWhXCxjLUjNrojsKS0NypfpS
UWlSFHjepW/+dLpMSeTrZUTkcjrHdpcHdn/3/5YvlJAjXF1DRt2h8GMdzsjtxN4d
kiMGkoPMUPRwnePVq2JbsRhWOULModppbECzke8VszTpMQWJjpSwqGp7tz2wljMy
o7wRhm+zLBh8Gt6ZdCB4YoNU8RdiKrLOQSakkmlF0b8KYhIFYZzUmu4Q6iHRvdjM
zKznjxf16V1d1ZwDJK5CW9iWuwTP5HKt/Rlm1ZTIGnT0mRlwmdddNwuhu+glrqOk
0q8BLtQaOTyMcpDcX/iALyE5mvIAdT7X6evlkpmDDCb18Ub8tLQnCpYVKnRYSSd0
3SOCoRGV/tCjqDgaIw2Thm3MYBPp4R1StXY6hhl3SURRHeg8dCfdywQ1euQjJ4HX
05sFeEv5Ejk/LFBYAW42MrLpbTfB1IJKXcsaRkahAPl36TGyX3V2GqEBMBbwoqm0
RpLTP7QztV1YYOoKlYOUHeZCViFuVTvIOasrl57H9RqSrosMf+ilsjt80PQo72/A
TiGVaJrnQviO+Mckk5NwMs39tAoQPMqeYtHECdt2uHe1oeAad26w6K4mp6TWIO4o
jG1l124OVD/3KaI3KzP+XEm8k59gYJi3MnnUvJjhfRjb3wTLfMcqcaZb55MZM8UJ
peyjhHg9qOGyURMZN0WKrtkR5JA/NJXmuL4X6o4Oy4EJTEmzGZRsAZhRzd42hrHv
cfTjCeSwMzukUXsOGOOkUIqOl6/5xVkzR8mnYgc0+Qmv7XjC4mtMxWI0ZOtIPibb
RI3o0CV36w/P/QmbtQSVYn75uLo6N4C8l+BiChRYX9ESlmL84FddlGTMMAUDHfzu
Em+y72n3gra37kZZOiwVcvtWq0zkWR/dXTtUWu00QugMgeOKZjxg3GlgZSAXmNzd
S3KprSPJiAWhv56BhUC0jYn7oHL3rqU3nKOWOxHdIed1CAeGvJXmbsGid6TOvJ6j
4ISEFQH5or7RCCKPl7JLbDKcSQWah11UmMI+26i2iVeJblv5FrHkyH7cQJZRCRJQ
zYg+iVDoeZJ/JdhYbSfRf0lBjW9nOZthhxnUeZIUmBdd116TMvX/ddX1Ug3ARNH3
PdiIiRGY1gUCgFmBVTtJLAr5DU0LkYEUupz96k2tcEbIoowa5ncgVtSKwBcLne2m
YmbEzNbzw4F2gfq9Ej1JxFjXrTeHFgGqStuVdUAcs5MQRKvgwzXRzGXFrmA3RKoe
sbzUV2JCwZTU/+IJvRkCsksEdkfSGuuXwMOyFHBjY7s4GoiNZtfCclndbFEJWDJh
0AT2FWM4gsHO2QuiG8KdPn3PG/vonrc2k578LmK6NSfJhJyyiTc9xF7gI203DWrk
qAH993dCg8psNdV62Tt3b4yaz+9SbS0YBKb7XCANa5bZiDZ0D/HanPYf23w5pQUG
YB4/2iIhwEvjUcb2hQTzFeCi24nnI5vtMOIkW7Dah1ZUswNcYgclny819CTkOIEq
tr/l2KW96lpHK+7opCzauff7ijkManhNfS9VjOeKQRyLS5DPiX7Z1B+Lm+TYPlzD
oSfARrbYcRQNLtjkzplPv6kCVRIvJG7C5qrenOQueYO6/ooT6ItfV0YTnkmkjLVh
d7rx6EeWEcF2VAYMuVq2X9z5LqgA3MSOKzUcW9UYzYTT/SVxIuFYX1IAEM3BBlx/
CWFDpTlCLEBfoZN6/xs0XHCIInWnDRm2VgzInnWSqyQ3Tn1rNhkkHlWEm8PyP0kL
IntFDswL8kfh5BOY5hzho43H0YUEYLZ3DVg7B1UmZvIVga63zsH9QU1UWHz8/CeX
x6rSpjJzGrA/VVj9u1ejmUunicY3eJGTiQItRmp3JEG+4FnNJ4+kz8y0HlLH7JK6
98drH7PFBqgOUPZ6z2CeA+FTkPNxzNgLXSl9phE9+5d6Sr6vbb2R3JAwG3beGuX/
Vx5fPdyMQXzmrWfPRe8cAW73cwM1Jur2lyaJ/XNT+vk5ZRI7jsFQ+QT9wtQL4eoD
ut6AxM8vDiYog53EeQ/esEGVUfyv2LTt0SRcoNRgVl0obRkYhbBNv16cIxfLMLQu
70YhqODZjk+RJYpMqj3Nf6Es/WQ1tZV9MPd7bP27l4FOVwCskRBN9B88sYHP5W9/
JFlbJgervaRBiFANdMWkoIhSydZqZnrLFS11Sd5UgDnJuTpMcvue8Z7reE9FlXrN
b2VccSIUBpbhTW+/flW1uS+5ZnsbpKLpKZrrPs+fbWXlrQH5kujNwN+RSkgBjdQQ
D/ZVyvTAGZSlKf4gAmD9U2SStQF+j9KZlrAMLXpqaicxAptwDijYaTOHGYreYOnp
+AAHmgytTd+W1Fo+L9rsl7CxuLyB1L3/3O4NRoOCBDXsU/XGFCL2EWZAVfb0YUEh
TZPfXXsLQhN/7rA59mvXqp2GkAFZk2SOh9vwDstpxIP4BUgCgyidM2jrAXK8exz4
plBvgoNdGNA55uY7iqkoJPFK4cayrxU1f/7jv64ZiZ/aNm2k0pkoydTtN7mGJ7B1
X66H2vkr+5KmdLovRSWvYRdg4jdE+JHVwKCG5xh3Ox04Urqoojm0UCNJev0SJcg5
+l3ffLzirY7ORiOgdxxv1XOyE+MMCnkkcbaxbgRf/n2/Ze/HiYCVdypW1kNN6U+h
7AKen0iHhVcS4EmcluaZkJZXMobNEGb0wDhkTigmWUjMW6VVET1d88V65wLaq0P4
p0PhtKDTVqDKvqaBX+9JGXcvaaWJ3NJ4wvgBVV4vzA+GEio9l1pwHVt7w8/KR1+q
BsvLu227hTlcVI81Yd5d6j+34dUzo6VDm0yoptI3EbUbkcGleJsogXbYnEzeYuP2
T62ov7U6Nznfgjbqjq/dDVCL0VRwiwzsF/t6tvyVUlTlR6M98xC0pwDXl464H+HD
KPUYRJOjFxgBnSmiqGCBemQWUp28cyfCMXB/8gmRaIHFWmD7LEW41XM2qWmmCaic
oAq9YwcQJ9F8BB+GLBfS9jlXOnepFo+Xy5Ni5WHNWlNzofXG0KfNHYN/suI/KJaY
pvz9FT11Vbl00TQBK75bn55IwVU3OnTQAPfPoLlin2zwVDOBKk5VUshSYs79ORaE
7BdGHPK5WsX2ERSyJhW/c/aXQoxuZtKIP89/fAJRtKdIacc84ovTOghy/0ABW3Fi
8mRfgxnQasJrMnAf4QNtbA0LHQTh2faDyusOE93TpLmyZraWfd1p3fY92XtPaO5P
zqL2rBHkSzHhj1WDYcAjAVxHewc7aM1z+Eqxvm5zELPA14vyVggyTVLk1q3AE0qI
UD+UiuhQc92XeIY4253Y1g5M0s5KMeTSgm1tKdkje1WCtMHSAqqTEGRvyj2gG/0S
M7ua3MIJOFr440l9k2KwSK5HC5TRWv0x6knXjI4INaZpsycgiGp5qqeXziMeaXW6
LozON2wTNdE8nv2yPN6GOqsc+t3h/RJGvMcfzOYGxDoHGDnVZ7CBgbixn2gcw4nZ
AKnRJ2VkTorms4u6qUoZ6ZNbbB2TjtuAIPh8isdMuU8ArvxV7632mhop64Cpzpd/
8txuePt6AfXcYel+Yty4hjkdfJhZysYl0emVjz9mY//FaWt9l41T8kzVQXCjv1u4
VzxgrCjzlGLiJJCZrndhLOgJ/m9FTwVJHYbzIynYjjIvwF0kjfjVLpGlQyItoCyo
LSC94rvC/DyJevm/mHjTZBeoUvJfTfYrsG3tgbnXW1C9EUjmjI723zfa9Qfa733E
6eRPKRILGWvtpYKoRhkHmEmWx+qvuo27oruISs3OfJ/kp5KsQYXuha/Cn+DcCgkp
E0grpUZWY8ErENT7idNeKs1yrJuSgWAn7Zfjotpjy6feK6LkXVanWJigcz8ljrVY
Tmha6/14ARPFcCZNMEW51j7W7HDH1CKL2PMQfVlM6KhOPjC8SCVsgIa1h8JHebrO
CuF3tvFn8KNY8aa0zszjYhqytGGfedYpn7ajZs9rz3ZqUUKj+BijgNOdQNUix3h+
4CmKm+OtzEt1JPAvP87WdKWn5Hk54OQbqx4bSTwsZlI6uP3crdyvfJyyE31hb5yv
PWj7oeJrI38I/od3UBMd/4i9tfqER2GlMszY6NLhhJDL8yndN0HypgDyi/ZsE2Ox
O+hbd7feQ1FagrR8dkA5TOIvF6E+1rAxuWA33ej8eyADFVg4c5kwjJ+knbb6uxIy
DOqlYUsbKMuYXUYi5Yzowrjq2BsU13xfIy7r75XsW6DvwAHZ384IRa1Q/Yo8rRjY
r4u9T/TkeYj/SG9uourSmVBSXPAQZMAXu7ma5zfmB8tLJdsxDThOrEczvEehCsUf
fwA4nW9CYXi0CuTwyemPRmHf6oVSNBptppmzIbsV2YWHozO3Ptfx6qGMEh4MGR74
m7Ti5b3Uf0H+jPNnjEjUrwZqxoTvW9HDU88P2GpHMpoc2c42ijpTMLgbBHWtJbNu
ZvjwdAQmq5IQUgRU/stPeonRqYzQwRrXEbVuN8FtIFY2j4ZjuJazOT2aCIbK0jJM
QFjM1xMo6Tpv2FN0iJapxlk9DfmRIdCa2xkRRlXZyxRBUXrAEhQjl6YLF0qk0Y/z
wcldE9zsn0xBzomsOq02kyHqR3srTYFvco0uBNIMYfnNQJ1A6wHXlkMNhmQvXhxm
yykpXAAthu3Bq9ptmxmx3PTFRz7i4oIcsCs8zeyszsYygSUOj0PPNitZUW+/gWPd
JGm2JObgIypDw5c/k7smvW5ZXNBCOvms+9I5KFQgKaGS4HxvBsN6wBkMxg13Ntki
F/aBSD1JfVNGJkGtPmQ13XFTxw+dbg8dl7wEV9Zv0/WZO3aPcA102IbNX3iYkFAI
fX8o3qykzqK0pDC+f1j1O2saGyV1k3okHHSgqUclzvrgoUYe2E3ObZe2vHrHFS2i
4/c9E6pyPkaAjQtGjYM7p2SHkPlOP4izTk+8qTgDXY0si1liY4aKtFEgUL52k9x5
EqG2z6JIn44t4uvYtOsdkQfdB+5cK2eNlKm3fstjMoR+97NnBcX0j4ZFT8uyAJuv
eRjrblCRUZRn1hu4G37bOhTudMATeHpYZYuYmekItDLs8g5ASzNqDBlQhzgb/Fqw
pu4RhfVkr1r/P7Q8ieJG16reisqgquI881HJe2NWGvQp6uf5fkIrGtGGrU8IVtCF
tNIbEFSPiAZTeY6j0VWWtkTJD0YVb/z8voDKHmFff4O7Y0zGsuoBqIIEsMCrHjRJ
o29MFy1kpxUvMcpMRNmLVxHpuJ2bkf9bH2kRfUExcQrPfNLN07G3wBxlmDOT42q7
qSvXWAEdZgseC8bfZ4nDGOxRc8Zxl01Wg7fPk4Z9PMFXwwymKP2k23OeJkpSPaKJ
dh/J21PVovEMukgsxi+k4RVVRC+M3y7WilsCmlEsNZlO2cMzPS4NqAJH54aqu72l
8vkM6jAiZMNMShV4isJT240oG4QXIkY642IaS/AlrbDVCZOt9B6mkZ/W9rM6bjeu
WqNxGyOkKgI19wjVl0L7vQkP0rF9x2USSGOM0o/cYIqsZ3Xkz3aBdJNCH0Db3w3T
oEoQTx/+LyphHhyuG43KlaXAXK5zC/Vgw2bwv9rrLIxM8ie6gtqEzROupz8sTNxy
52eY6ILaZ9ZiISBa5Bj75SqC3CHjgTmT5cJ3nUbSDeJF5C+8syDr5LQ/o1Nygf1f
1jNQwihMQ88lLlZgcye51AqTNlYfjKJ8Z5j6G25UJ1QuNvPKsAhwwJE75e8czH4S
NY0mIagWIl8Upqs3fIkjfJniIIO0st6IUA6jggZjtoHU+JYjyyx6shjx/CepCGpN
14ku0y9wS+QxvJX1q3YoVnQ6qtLN9/v9YLawhwyzum7u7ma48g33C7XyDP26elmR
sdV1+0mp21+bfUX7yU5S5BkIrHbVI7/i4VAGgtkSrU961PIcdmYkGuDHv8dtX8NJ
+90PZit0Vbg1nkXVlg7inmVmeB5stbxN47nakO60GM491LlS61+Lq2iLGoP95lV6
iqGhOsm/No/ymbu4uoA5McNNu56pp1mWCTfpnRi4YoNBKzwuvwQKEwzWzsD6q6Za
732NlOaEXT9UCo5nBEMpYQQTapr77kZp0DMBd+z6x1Gy8R5jaFSyD6RUfPNNYauz
YkVrAuDK2NhDT+AszUD+tuRVCe+NjCpH2/YzKmGm4AI8UtJp4t6IlwyxKZcjKfRX
h3vM+sKbWHZVBH7TnSONvQibfkBsi68fo2sz8Xi4EWZUHhNzZDoVfeJck3j9kVwP
SdqpYCkvBU19mWXXr2ZnaCZBhrtvpvlxB5Mo5r04RZCQ8bF5qFcAQjA52BLtrcWf
PNYTq2RyUiO8G1/o2NRK+EwgDfZ9R+R5NdUliv1pBuJshGEf5xQr+QIojlYDxrIp
AUbRO58wgAwPxkWjmIC8KWo8H53aPCnP5HfiVDwKfHSsChR3iWFh1BnvemOnkie3
MKkZqRvyzoaNcvbr/0VHzZ4kRdzoWwJEUdvkUdy3w3+gYe5Zmkw8POPSBzSh3yFg
bquReP4Z2BsY6p7qoYGfctMM/AmH7V8mAejKzBxGGqCESL5U2n8EnUBo6kyoJlmw
YJql7bEF15NrvE+xR51eRxCwQ3mvAygf7bAttk0nc0spKaVC0mgn+gGffAVNfYFw
tC2Ch4cYrh2INfflsxV1cpwb9e0oWSA5PvlmC9OukMcQoCPGYXAZOoBhcB6v2cGk
a23mIQZrHh2274V0swnfon9+1eCC6N+ixmQTTClZs5nr8baJkC5qoqK3a2bonlgG
/mEM5OpdoLqNELiSUTeyk3FnJH7SbaJfRd3e6QeERkXUE5u8846es1zaC0kmeGgK
Ui/Ypenl01ispN+vsnvVHScLpRzu/RIujC3MJgTZ0tUTqtsycH2jiGwq2od6fN+b
MXvfv8FwhGT2zlSiCSvlXbIPD3OeqntKRTXKB0ZgPVizyZhEWolQVX+Ti3uNg7Vh
yyzOc1PrLeJguUnqWhm+ITZ/TT1JOzPfPkbLHNNXbgkG+x8QUARBXzvRkeBlZzlj
/A+MhIwI+mpjHTLW8LxoufJEpZUK32wwkL54dB67d3bmjIjj80B3TQfYZQH0SXI9
UYgYs8fvOdkaBe0mypC5QRVmKDognjX3ral1zkHbsgogD4jPLoqlxf+N9yxl2xS7
Cbq+M3ounrbl8X7ukMowyLPXZlnAEgK3ZGHwXVnLO6u8z3VGa/W0Gl04P5r2skr3
rsXmwXEkIf/j5TCXc0c3Wfuim0Y71fpQw/vv/YMpyhXGy9GitqAqtDSKRy5t68Q1
knaIXtMhzy58GHuU9YmuxcBUUDzN/wNO1V+AGD2zRmQPlxNgN3PJxy6TWSl+EscZ
oi5IvE3TFnmoAHqZtdgz4KdrZKs2UheThSAfIwi2JIXGNniREtolUZG1vEexWvhW
MoCWzNrK9zSoaK03FhKLOZDr8YFB20U+MCJ6OVmawk6e2AxP7ljK/wMGtZc9rTuW
JEXXIkdyyW68FNs/pnhbi6+PU3awIIflzsyIJy59AY26L7jRwGGtLx4jEkTYnaZT
QlHLcAG/XSZpA35tMn/LPd277t+kXdSg/ilVymp6LQ0w1RRZC3VjWj++hlnbIvMI
wH7Sn8YrB35gt9jdlE5Ipy0YXMZ1DwC+Cgyo8H7DIdmAmOOPGl0q2z6rap5bgco0
0+zbhjKF0kfHvm/NkC3saBCoSYtc/+kUOPcV1NnPIvsyKAVT1kCHoyAePvCycJWi
AjqmpCvJ099HQXlrkGP+w2Lf1j7j0RKNzUPnuYTJ8fkcNaFyzgTqFrjBmcFr46GR
E//3VqJHIlav4VZ2XZEfEEfcDBA2eepIetdGkwSgK1AXXZAmH9g7NwYcLQzH9dLp
moal0b3JvMLseaNgeKNSQNAoxMVcNKaAdVJnRzEKy7t9EfFnjax9PDJB6iNH8pc+
O6gI1mm5B/FVZaM+w7tHmSbohyU/kkUWFWG1qvfLFXWiZyP23AiB5brhUz2tBNfO
2e4gVgmvmbyZk/wnBcGpd8C/B9FVc1zUNiBgDeBuuzhGfxvKdyqXOeoHU2rSqKKE
GCFuKhQDcC/TR3JBoFEgFs2qDfusqey2fyS+uVx7rfx9iJDqywTJJ7uJ8SRTA0xj
WfjeJng5Epn0/rW1swkD52U/ScJ8+POXf8FKGHkPYnrU9beVQEx4EoTz45hS7fFu
UhNjRwhf3KH7g2O5bLvIYIIO16rmjYo6ZudNpxfpv4jDcc+mG9nOwEps4Jb1IJI8
Rfw3/Ksnhcck3qmxOAzSXEIKq6PGq5Hxy5dh+Lqz/Mm3zzaSfTbFdqDuXvsoCtOJ
ZaY0czSsoZ26MRqAf4xDwJYgFiNwLt2pu6B3f68uq6crLfiLszc3G3BFnbD0XFVu
3JWyjcdfSoxw5YWlghh/j85oBmrwEJ3B69LIrOurZxgRJL8gIBxdtmZUapTGvz+Z
RNNu9eoc1+0ui5UhAQUzrKyBiYcBz5n1822HCcougiJ225WaY8Z0+DaWxO2GaNCU
cKyH2h5ZyxKxNyZaLlSllDCgAW/FvNjNHO7j0Yu+TkZc3cHDLff5070ifp6K1v80
VAF14bk9b6HhWyOrKHPlDJf4p+VZAyXtWl1GM0wqMf0AVziEufplrPmRzJAi8hat
j0NibuBT3wM2JiEHfq7NPogQikX+eHvT+UE5elyCXvyELmWlOWfoqfZnZ65VBNP1
aeuV+EAV6/0LB4dN8GJCtJ/hLTLm1B0NiZotoeBGrcFXlq+oqgueeW/uhTtXG4l2
Hp8MuC+URvuW0EMhGxmMEAPhTbthOwnA9+veBLEsKq3l9V7UDl3MGlg2tyg+iM+q
O7b4QFXHD+wooqo2pr/R389vdm4qgJS8UxS0j+Hejmh0zsCyLVdLve9olfagmTZk
bMmhYjxxpoeIjGXVW/CIpTNrqf5HNz7XsEJfRzKwDADe+ywKeNyCAA2EXRwvhExA
JFcPxpT1YLxdAEURIkcgvgHfJmUxv5ZbnPOOlI4qKns/V7YO0TtfeCDnKzx36e0s
TaH8VplVCWU0jqZCdFZBXQ2bRwCYQ0rvrXChMS12c2HhXUw337Kyi7NqADUjF9Pq
Lg5/90dImkrOkT03V6Wqyizzlhs+iS6QPv7kC/fxo/3I71k1BSO/GCUU/s1cnKTf
kwMXP/Vxw8R2RFB0kZ5JHWh+RXLBWbOv4HteIPcEhkX6iWn4JHfei7JDHZlAAWMl
5Fg/gYhcNt2CpoQCbUbQ3gb60dzRUFiJcZ9FOWOXgooacNL4qv6GcK8FACV8v9I3
rFJ1a7NotCvyfkuSfa0/bfv5XFjkQULT75k3Dsf87cMnDBddjaj6uSZKvrd+OQwl
fwGEecx0vKd/HWhK3IPpTVSAUUv6K5Vgd3Dpf+ShiDRvwylq3nT+gpNMfzW4sU50
kEcJKJW2u0LZ5hcrsClyC7UHlcAoGlBhIi7iJz8+pDBOiELoYnin/JeVS+gWf4DE
xzFJbjvSxam1nYQo6auyrOdTF3M7ssUW35bNvWoj2935PCXRk/HZk+eVQcjnd57+
tJLrEODnLSHVFeuArvjm45hySEPS0+2QFJ/ojs7968b12UF7PBxOlWT3KOMA+r99
Icp99BroexWSJUmyjwNOMOlTPg7JIrhIdv/CDyNvOq/n6J/UuGgRqGkdC5MqyUu4
nA5TY+TIXpBxk70Chdq5uEZ9xq1MbMaxivOrEJD/ZcP51KlRf57QKYa3kOWlHz5f
7N5Y+Wd75e2/naak5EUFPqjL+XS10o+DPH88kqI8SPCQ7qi8/KtBbqzfyR0uhDey
B5HK0ktZQ8Dt8m5whGbEw2QJ50IzXSHZj45zgiDvADHWpR/4KJmDS0MWM30dBebh
7BOcv99YxkQjADbFQYUgGYybHG9pN/Sd83eUGtm8+do9dFOX5WUf21mzzKEfpTRr
XCOYPyJgvymxNDgAgw8PXbxlV0RnxAuIApcQTqEGD6MjNaOkCDISrhAmajfb4UBR
H0RWhFvuGIVqIHllL0E6YI2X7TikMn/E1Bldw1ngFeT1cCvDampg4XR/LQTOTPs3
j87GVKOuoiuS9kfEPIt6bVWa2qW3/CJc+lj/f4ngf0ew7KaeLovuGfqSPBXHZ2yO
WvfP13tQytMSJSQXfm+Cyg6bTxmCZ11y5speZ/NMQ26jFuMIrNo7/GnUZ24qW+vY
2TteyXJdWZhiGcnFGB3mFz7c8Om/biwhce5jvYb8jZpIHK+Xi2DLQCLWGFD9+0+C
Z626ycBaHHxxpGzojDah5mhJ43Sg2FaQ3BJpbhKsLzaBREyfeKSJHtizJJYb7Pdp
fJAQtEEl+M0yuxMWyeZtz0ecatOUN2yzbxFEgYvIDY/vrZiD2l3QORxe3xEp2tfc
Rd0GULLT1QDCcndvkwGHrhhREx0lqaoxK18BN9kqgieNikd8i69Gf6B1o7ovD6q0
kt8CKf9LtA/J9CifyCFqTDMYsA/FvfjIzWjXVHv9dTmgLEtlqEsDOwdWSq2PZpu8
6TfusY4imLu51dYhNQmK8cNY5Boh6OR2IC7Kh/eB8SEyuctSpGMkJwnYr5cPhCmZ
wUHnT49khIMLSf6ZHKR8pisyDStw7SQAUq1/ioqb1UUdOw43ZscCGU95UUF9WaEV
XAFcXX4yv0vBZKOe5DrTZy//VMFDyoyTTniGBylA1cFkC8uiK42bRastBSLprpoZ
kFcu7lOIt+dv1bVLZD2rIeh+b/yr6lJWVrJiBiUzH6CMiC5hXruQY+c5BQqfS+51
BVWPjo5sRbaNGum5Lqi24xFbtOas9EKkuV5eEIea9Jad0L/tq4uUYRlhOcW/SuCH
vzBWUpLK1E8jwg5ZQdvQrRRYZYU4SzDJmd1vsuYRVTiOaFUNjxysUPX/MbbdY7Mf
11WqHdD464je3OJWgdL+Y39f57RHND7R/ydDKzG/cDo50WmeOPCSPWxmvNopIN2R
A5MPzi9+jRX6Tg4JD8c/SvDYfFMKhQmTrjuOigpAee9Oa1Nqh2+3YxBnjWSx94/Z
vVlT4V20ii4TxNAS8eruIvDsB+aqpiASdt245fxjMgSsfSeeDCvupp2+EpB79tVY
OVm2bs4oj4Ft5zeJzmHsAq8cGU+iZMp5SJYDkTjXuGxRgBVgVE9X3OR2m77sZ/ST
nAUbCDW0uJhjkUPZzk/InWBA27fcuI6bkCVEjcOdIGsIgV1DHvGUyrhWbKaTENZV
I1mTGWfE1ILgpzwgfCDFsCp9muBH2bxcOTrPImejwBOACbiI0L6Rej34ym2REVza
zF2WWhczHgD9o/2RgaxbJzKPMN/k0Av52ijy6UkI+6+6LJSvi6b0KtTmqLuL3nUF
ZL5Gh0FVbPf3zl1V/JqZYwZcB39Pc12s3H1mHee13R8i0/h2SAsjT0mrOz2WqoUE
RdS78qlca4pm8bGcJGS6pw1IPnBBUYZcPwLosu+oAQ/MFeOQ6n5VSkHldrs4vMm6
YalJ6mGFqimj71brp+WWMLF1nBUahRyqv+2gwQVC9h1z7jtX23KGHTLx5Y7l+Vos
swhAlXtui/Fttt8oLYGEE+3advLAMc9gp+ns+UGHbWxJun174PrqdhKTbppIBzZF
g8plKFJCCRWS6Awk5G+iTwgoS9Lpx7qjLT+8R/Uai2LMvhSLpScyC+6XsoIzBEXm
5hy9gvOtQagfkz6UK7zFjdQgmKrHik8n0NxGDCXH+MsUsSwsqgCRIq5wrIUBAStZ
EbHikFOjVHa3alNRVQyePHxtWtRUQogeoYu0BYSHlnWRpZc0qwfj1vGP0d8MxZ/r
QysP0laF2TY4Nre+VT0AG/e/HHYOWX5+snv0LtyK0rYlUpWomg8v5oUDPArvMHvN
tuPtS8rwtwTO2KbvPlgPOUS6cZyrh7+9sH59V4h4m09NvPtadWc6FCXv8rqofAOV
uhPRJfL3PFw9xOi/g9Y4T6VDL80HyFTcuL5nuc6dYDA1qtfuy5xKj8dPxlBiJAbK
xtN3Mf5Mg6HfXUI8W6yvGctLttIdax4oBCdCBRbHhwsemeTW4boacvi3NVBqOszj
SNbd7/E1qQ67DVyB3Nq7TuTMPLPi1EH0LdErXbzKSSqoqyvI5X0YwdCLeTp5GJv4
vouEmt9Qm8GK0LTfjXFYKEOBhhaPNjc5+dlOYh5DG2e48GxX3l0lo6XVX4HXrnvO
9yN/82ATlKTWdISiaT0c34SQR2/BZXrcr4mLN3JL/Y5Q4HTSwjfS6N4rxjNJsIf2
XEjU/PSu/I7TPmN9n4A/mZ1q7reOh+7BEAwAM9N4V3q9yP/Cccx2qb2zZIAYPxF+
ynxfFDAbiKMY1Vc7tFVPTMm2hRnqpioVNy8YIGSgqiu9m52fZTgkJEdBGzjedImr
ITKP/P226A+SKwnPn81S6b0WUu374BjtcNsXcsrdVChnaCZtIXmPdCQzByaYsnkZ
NmQcYGibEFfj+Jcy/mPHj0LO6ChXiB8/PTDwGX0gCe3bxVh/F7s+aGRsaDmsjnz2
p47vcqtnqeNfWKkwcIa9QdHI+z/kPw0NwhH4P5w3+MZ8PGJJX7qYQafbr8fxG1ue
41L2luXrhK5YhiaD82RZW0PzvKSO6B/5tvtjTOTJxWbxpbonS1qwTn6SBdQ6Gm45
MnE1Iul3vGREZaTx9m87hoO47ES44T67lsozgMmHb5cUQ6n7pWXo+I2D/HtWO2m9
0UzSoRQrunpektzUBLEiHr1OAnxZLImWO5tSIWevJMahI28l+FEV/gTPhsACZbaq
313EKb7ePCR0Lyz67oETQLH+u27WOvaVJ/xKdsAtpRNJDA1D7pR56yaRYNYTarjV
CntPPYZtO09oCBb2QWJLQr0/QTAqAD75hNPYiz+cv9Or6HxM5VttjOt246qT/1YM
Ciz7KImkBsoWFag7dMxslJv9TaoWMfuzhtHl2c7vid2rVJ5IDy4c9i4yk1PBFTat
JyLctGuPhUO5V6Gsxd2/Usc289t9Gmk99meiZUl92yh03djkC6B3Yko+qKrgWT5u
oYmQXv43ntvoKMonoxAQaPbcsQzN2FQHdJsk/rYlhaFdxxAzFMeIsZnX1nPoCCYu
Fkd8/domlAfQGmVzb3TTPOFTiChOazM/pu1UTXdZr3jD52O8df9rScIdj1QHhG6c
BHJRAn/0wGXKM0RnH02AmlnXVdDXIiU5doVvFiaJp+hcz5t0909Qi4t2b4KqoGYK
bvoOA+kx5ZCnLB7Uk/jnAUOnxAlP1NXR7JY8GGwPoGFHt74A/j2od3Hz7cE3cxnW
WQusHVHr9fwHdjpmbfixrxWumX2G2uuZ5W1KnidUTq08M/YxmNNYX3765fkHJPr/
XdM+uXFzmj1H95s06FDDgd7lwlvuJKqr2oWMaJn2c4itl40b7mrKJTg5bIB4JQmC
R5Ew1VMVwPfwU6Sjubh8k71p5Zey0WZG1a+VJmrtVwWxPPUBJpoeHYy4AlcVCWb4
9on8IixDuUkGeeqQi3inyDoZfi5oMttJhtSP09pYvDlZgk08W+uy0hWy+Roar9wN
ylJEHC5bkMZppuEuGVDCOChl9m/fwHzZE/MQ3qsPsN4MxxaXvcalNUJbR6PEHBSM
YWcld/58aNB1J6bGfRcAjjpB+C9ZowZ4NOdFQ1ymFvkmIUkqJu/qQQheOZFOlbHj
ImlaTnEMe4eGUa6f+dUEy4GuXA5GWMlF6mVSvye+A+8FrYciXhRFCTLoiPi9N0Gt
BEGhnINF3vvMgLsQYrKQLE8Gy5OgFclH5U+Ngou1zlmSnEwpr6KpmLqHkAoV1wUo
Pt1bBjfhTicrYLhFGwhMURjRltfhytyAsSAd5dYiTiHoh6ZugsbV2WH+02F3/pDH
waWKJ2ONvF3FuBhkkB01fCCberSU3LLD19N7jRkd7VQ1LbRHrF79Vm+tDI0UhmZk
WIvLi/xgnF7k5/4D97Q5jZBOAu2QP6UKlkoMRN7X4gVaGxYmwf28L/hlgYuTmADU
QfS671T5ySj75m4hJcgcTo5RjHd2q9V3oulZOcdlmq4CJa9gTePHZpZecCVJqOEE
pjcR8wrV9XBO8D4HoCewVmQJRNyUlPXY4kIFSXce/0x0P1R2tlBxjNSPQuSYbKqc
sVvM3Rq5v3Dohv1yG1kuTUMFACbo1ifdwkubIByrlGLBjIWmGqTxx6NnGE+79+Da
LRzbW2rXaA5U/wLQfNgpx6kAsXWoAzWOc39z7JeXKqCZJxqxtdqmFBZoFDhyHch3
yAmJ1QpKEjWgNuhHIUdj0IO22ECpXdB3LY49yXv17IE5cNFpkSHczNS8uMg82fc0
YcVmNzEVnyX36veNC7Ac4Oa9JSUDEtkh/8kYaLd2CKCiqIbZAnxexWZ8HH/CuWMl
WWEr9Em5EHFBe/NtEOVF9Cz3P1gSl1oXofU+Lz8gd08/UG30filMCH/ZTxlZhj6t
Opv+yNiq6obPJ6wf16F7ccDHmSfkqYPHh6mj5ebFEerlOcXoTrWw6tFo5eG057j+
gk8PfDtkJVS63YnELDSvPuqN2TGSP3W/lSRonCN7OmwPjIbEIt8yqdVxB1cAK6dw
6r2x3X17d/ogJtT4Z+RpNDaUwqhbG2gwmDszu8h/D/jXZ+ix22uAJ8Nhp3wKC6LJ
0Gs/+ula+jiKwZSyPif4mv70Vw1NzLiy6CXstb7kLOnBKMw0WO55EVURzX3M3/An
Z2p8BVd34AlevKTI9hSaIIt+McYD/+aJikZhF8OdEUWLA61G5LS1e2QKHGdknA54
geE4ZRa0gagiDBSHKtT7PZ97QRj3BXATdYAouGx7f1bSYss5Z82JkAEt2IaPnyuf
8N2sjV8WVO/aiecOxYHMQTX8bnSaLBoeHlhY1rdplBNzBogh1SUbXT0ZNRTtcfhw
pxk1jpTha0jaGEKoeoQkLFRHYRRQWL5CQSXy4/xUdX34GsveC+Nz6iJBtLCQOrBM
BaoVzo2MLItoh2+vvZzRTOsgCiso6vnA8EiJA/hk/CdeZgbg94L4XnzySwTGuUp2
2W9qR1Llxh0PDhKlBOVXUbzZmAWugfVs6Y2P4wZDCAMKMm26sDH/ZT/3f8WVKm7q
bfJhEsDfsc0fVqevaPLPkaVyTyV+C1ro47SaFD0/G5pPQOHJP1KVXctVX41zDgN6
PfNROdd1wOXEquPAuIxrzlCyYudzzD1YIXy6X1E0q+OnPV7RiqjsrwVRQXa4zVSJ
mOE98tGrQ0K7NlDkE2uAnLcMfkH7T5CjoApw7D6z9Bj0gRDuPI39QxhdU/r1ZvGZ
bzeCtRWbHIEm1CGg5E+nOt9Lf+xcRprO4XxVkXzzau8mtIOijQ89geqLsnoPUzuY
reDRZoCGC/FzaGrDmJR9y/MBrvE6Dg3IsZFMZm7AvDeh5Cwo3jjQMIh/IMFlDsRf
xa2Nh3+zEnxdrkteLP4vhWacgfGPF9Winx3ah+X4wyjhW43fLABcN+fZu41b3CaF
tf3Oou3l/CXfSBWRjdI9gk2gRSS0PSpoTGVO8Y1+QVbNrXXkVOx0Ta7S7eBCdjzW
ey1L+OpLi5m8Z6e+e+nU64A4+CGgmem7PdsomXl8V3MXXnfP8/TQukNOilPqRtEa
NoARcb5428n3YAd7Q8mL4Nn5nYj0yZzFdUaFvvNKU/Q3zf7ZiG8XZsMA8Mnlgsj3
118IdhsK0C5pCIX5UjIHYd3BJK33Jx64G0nEL4Fc/edSsOkaDZV3zsSWulUbCFTZ
BWF4AWJnn+gIip5Z3m3RbiWWoJeAc2fsVeFHRalVhVCjkl8+gVWmpQyPfTzglVuQ
13qFdrK5nP7mEGs/jOfgdXg2ftUjJCTBjYuqq2sDpy+JNjGyH/f0cRFpno/41Lrx
iUZq72df3qC2mWszpD3tEPFvlC4+zTlnhqI+K3mMKRnZKT482l3OM2QCf6Yrpck3
2W8/SwyPexsPkB4vn56npQo2IxPFTDM5jyH37olWbyGViVmyfTa1hHFXsSnnmoJ8
UG07TOaX8Sn3Glm5l/m/lt/U3A+L/EjBQzyWhzEF1l6HifY9vFUTyn9/j9qTYwqZ
cQJb0JTif6pxP6U1DDLVtJIsh6PRXyXy8OtpPdMUethY7w1ZialgooFvucXDu5bf
n4FOSwWuq6HAl8EIzQdrA6DEF/bhZGVgin1qwhxoJ3Ax3TequXJjeL3hKqPUu6SL
q/kD6EmYo/je9+4dDqIPDM4X0WLtyarHrjqa5klVz7rDWA5wS1WQYi0ycUXjbYvd
OZMTl3a/r/SxuEK4s1hDV2sHgqZ6J7Ny96BZqpWDNLtKeachqMOqxJwVxK8TDdV0
ihk+QQEAtQqOBB8GKobuZaorBmDPgERzv734LhlTvLjKdgwTSVlP/tkGlxh8igc9
l1//18YLZB0sWnUdgr5VRj7HwNCKndmJ8hCLeAH1Z9bsvUfHwraGxWEbi8ZBsqPl
Hf+iKPyt+rSNOqlW9vXixxSKw4bMzrIiMzuw5ZvEPD77lk6E1SSfVx6LzaIjls47
vN3vVmWO+357GMZTAW21Olm93S/hONWaoua6Mmxgu+g0WzWHuFjtPNTxTyrw0lzF
yB3t+nNYvjNaPr7bfWywm6Hg1dJPHNH/d8prnHpJa0rrljY4FZa7DI7Z6PVLfXMS
eR7DXkpj/C3JkypprdjWF5Ej5YuiF8K1pCqMpxzdBPGHCoPE07Sb4S7w0zP8fJTi
/S2N8ezfCDIFTnAVqG1iUAGS4wxx+uJNKAd3cYlxo7Ur2yl9pbqwb0H6dwDKwbh9
fJCmZW7v5AcP8oteEM7KJsBQPHy6fuuo6nNZQcdVCoZHj8+yjB0pVXYFwAsIexio
UqCmirH+AbZ3d4U6jM+vd4durIh1etKqI6hSavOCksgcqjlI037zy6NsddsIwiKv
CxGaPUXFRPZI/sDHsdQ2RRxY2qKaj0sd3xwz1C0iBbPeNLHEw+NLiWLoUgcDagq3
Yl07EAUfzRB2fTvi/+wsi5DaWcA1UdHiSHyLcAZagx4LB4Wi211s9HnnjHBNCWGM
s06hK+MIiW6OuIQSWZTqxNgSvCC0R4jIutqiSU9QRSskY7KUkc7VmBWcLDp8yOYj
I6gn5K+TiqhYbAevb0alUjUSazN1KnXKEEpR9Q3UNMIkNhFWTy6XJ8/0tPumpuBP
ziIOULBuHNRMWUjTODFVhoUE/RS1j8PcMm88xmJfYhXEvJ1j9vgdrIFdBHx/EEId
z7Z7bwkLYmrJ4OP415xBhXBCdf3l0l9GPoSbDo+ctNODtVQ31OTM8HkTh9ixBSI+
g+AJS3/VkXERpQRlZtgV/V7GJSE4ZJkjg0L7YnrIbeTn9MxTkFHCfdIDgeOINWie
Zhx0ddePykW2o2uBDoZg8V1VaTXdHl7cpJz4SCLb5lbGzS+sGjtdBUD4EYtoJQKH
/srAQbiJUXjk/d9ZgNNutLMtKi1shrmfH07jYTueNWwMB6X4880UEAQCns4lE81t
uf7amEW0L6+H1qNZiqIMDG41YBOVDHMcWYYP+TLxw22fjOWo65BUSOmZJk0ijZE4
apAL+SpB8O6xZHYXen/W03CGMgxvjGft6O7C9No6m8NDu2EEBFZZrLkM0HNRH/oo
gkLgxIbe30EAl/Slj62spLHLZUJesz84HXecyCRin1FTD/0ead9mxCgLkK8FMLv1
HJWbHbxW20oJEZQBRlSq1dP8FDhmQmEkUayLODlT2GIudAy0DAfZH+Um2i/8TnNc
5vW+1zK/fNGYAieLJtrEWD9IN9ImHBZs9J++SkX+V33/eONkdDQDxHZRxOUaO0T1
BJymFTgRu6adTrj0aVubaLHHwoAamHb6aTziiPFnVpjJgMNDGh/bBvCjRQTNSNde
k/vMXUSf5lDwbLukNnSFBq+SyKXmyQEaA6FbZm1TEbBWuJoGKjQ024Al1WLfjyWR
IVkkHEY18NjoV8G8U9wCgKRDkTlAcLAbX+tDh0mJy0890vGm3hc8YfLy1cBlODaj
Tf9n9MmRzTZtFAJyTfdfTYRnxRnPo/cR64AjNRKYvMgfKqnIMctZAZ5DU6ULrZng
fjmgqb5BUMqJTkGl887Sm8bCDGvYmyF+6oVEnTnnxWpouHft9AU5j98jbqYSkK3f
as9gpdBnetw2gQN2XmsKoWiPYS8bVmowsOhA5FBy8AfZj8MKBVcrvlqW+H/XB2gq
x/4PGoaFDFEvRSlZnsClvPftiHtgcJbdg8ywGm6AdUvdAw6ZJzSCNa2dvxVgYj4J
TtT3jnaLLfryvky9qrqpndZGjqyrtZPGihFBrhqPJKSLatThDXPFyl9XeLsXv08d
cIvbFfCu2IvvsG81iNzrCpZy2D+GsmtMjjHco9ey8yWC1osfyaWmkkXf4LVroTN7
DbytNFxQIZE48p4h7/srwhbIJ2jqJuwtNhlac6pV7L6LW7lmbRAFgHKiJMOm5ez2
c8IO15bXwV5k4XzI3ev/I2/bt+EMetRwG8IlaVAw7+OiZVhNs6I+FUXK0/u7hOdp
04lscq4VqE4mskqxwTZH2/WGppb9miCIt/krLZ4p/FRVErqbXpf07XIM4bd4n3lY
IFSUp11b5YT0DDk4tH6ENbc1EpM/qWJ1LG9zmJ8d8HB1xrYL+5reTik0eKRd+Q6j
jr2yQtbRcUvDqFINonX9ZOvLhcSS/6WoEkY0fuqx9eLX87FvUKx+DyjcsWXtlzqT
P1gzXxWBqKGYMunkyI2hniAhl3494WNnimUR5isSXAOSEDWAdZtU4S2CkoayZBAQ
HnQQSZhEzPu9xq/o9QlfdDW71G73JE42g02ICn3I3fQ8UYlnr8AmxQmLsrxpXW/o
Es0Q1B/9R06ELe5dPSejRvPcw5+LY6i0nMKYzj9B3KuxcPzoAgaBRkIlVf5VX2jY
4m8FyqOBVMtokjIcSOwm3UmlyPCreBR4zk8pWk6QxzUcv9BmRwSggQCXN52TGYlp
0D8IDf1KP0ZxlvDGyDcJb9OpQmWzsojdQ0OFz1GsURZE39xUS/clOfJeE00ugXh4
Novg5EdiyRRzbqwV54+Y6TA53LjuJjgBcnYL6eG+kU1EuodhcdKBNloVrBLF3wR0
lkuJ7EsgWIFCmxhgrHH8+RVVt4q1JciV0rgjc1Uan1jaZ1u6PViZU0CufUj9DKBo
5MKS82p6p7Tu+ixFxX8j9d4YEvM4kl5Ag4bQdUDwPmIa2LzPwF4mUGVFwbT4tCW6
ktHq3/wyF87h6vrt49Q2wz8WtIGfW7tcfYL+zrPtGOw5NRAPXATcmpNdIBGe+GZC
3wR+UhgeB73PQEuEoKgBlthV5/IuFyjciAUCFE4seFPfY/cW55N9s7FW5KMWQbBf
kYQ3koOLiq5hcMIOh+vepvwEy2qp10klJorDimP7/yqkDUQZSRLg07a+lKlJ37QH
eo2SpJkDJox2P/E3VcP02XKiEUneo6nlxDFc0M99rOvkgK/WK78WkCZfZObUUumY
/etpKjNLUdG+CDnAIaCGg3SCkSPDU0R80yqgvlx1BwsxKw2p1fHxASHLy7D/HpzY
WuJ9L0qYIRBRMZnlAwQ5m2w/APwziG1UG/N7abcafkh4Bp5003IpXREKpoUl86XH
L1YT0Szw93MFGFmRbB11drXmA5kpe+4J3NymAluJyQojVAgpe0Ri9SvBwcbZJ/v9
DPrwkDZauMZsQgBhBa5jnzBoHubGvDaKiBS+cMVzOmDutoIGe45mwbHTin6PCIbg
SBe3OlQTZKy/xnCqMUR2zMmesnWO4okpb8GugkdrBY41BX1Zq0zJCUIDUrqDwHEn
oTgpkvR0kEjQXtkMPjFqQrQwUkxbPE6W2WuZaNWeooRt4xVbU3fW2SB0Xr9GgZUr
yMj049LoXV3Bbxqj8V+8dTVad0klHlMYvxQ9uE0rTComvjKAs1q3cmVmJkh1Clv7
0VDhald5h4XFNVBebzseRHGkjoisTTTkqLckZ3uOoEE1yGMhUQuvYjIxECAWYal2
UWA4LGNuESEtszOWWLt2ekt6QuRHOZHqWwiatEeswmj7504CMx4LBQgoK+SIagHe
6GaqfLefuGPXKIfNv5e5HjRrfQ64ktD7OEk5btx8IsCo+CjuB5ryUEillvy+fFPF
J7hEOOBO4wBs/VSlrCbz78lgyYRainqspS6G+Bssu2k0V82YOHgtz3RroEudCe5+
42oyq/unV4xl9Md1264dL6n58qAFtOT0g7cRrypbu24gkK41i/uY52sizmU6MzUQ
xbUgOgB7KU7D1eGIsgkmPdYUMcSuu3DJbf7fTX7qw8SFgk88hgq5XZmaeUj3tc3U
ppTeQc0vebiAEN6jVlluHrqckcoVtb2MKC6JsSV5RC4r3A+P4C0Zs/bR3La0bZlX
zy3tNmOUCQZUdWCkmrjJkJzzUqdFg0Xb50j4ChwZYtnLGEJKOWP4SB/VPZZPLt8u
izNjOLU+Rf0gxhzJrJRzGOMBMQxO9AutSa7zhBJtzvWA9UKd4ERCqE6H0iZOXqkE
8FexQauMW4ZtWfnj+wVGfqCUgN2XVL5ZmKbMuEIzSUgQTMjkPyHOCorBJAZ1vQqw
+kfoDlpo09sSg/oihGEQ1ea4MJrHrIxayRTeR5+EfaJttqtzTaciP4WRY5oenyp5
yrzZ7FOboUrMdezHB/qw4LywwXCMlrlipORUKJk5FGjyPawPQgCJVqXPpvFRDS6d
3B1Keb7/OTsDyPjDlj1jI4xUi6fCGSygsyvlapaw3/4rCQCCbcbQcsLSn+s6qT3n
STa6h4fXSQurR/EhAIQOdIy+iT893ArSfUiVGoNhVm8PRBNoh7uJjCCMw3gh4K7v
I1RKV8FdnCxyfjAgcZjhERqPh6nVrHXXPTIovrQ6pitWsii5FR8so2d0ytemj7RM
Jv23BIZnaK7Ci21kbwxUY4jFQyh07qSUw0wk1GruptYP7YwaOrfAEzlgEeQyQLU4
NRcaG2sQrkmIhNSRaezfIerDNSZwbSgFV5mA1dQvZdLHqOgufOlofZK0s5Kb/dUz
iBDbDuuah7NhL7lGVQq5tyexgbQwVf0T7w9K8jt4gmNYi3ZrZutGKSKMzyqADEUB
QVpe1nFfgSyo73rc3ionJAU0UcMkSpKX/tP9HxjLPIHrIKU+2ActHhND5V+BaOn3
uWQ7KwChkdP6i0AMxoTb91oamu3HBAfTTiobBVa7mtizJLS1rlfEhN5SV3XJiUdy
lyIZNtR198RAkNhi/RliFdT42VlSzNWAa0V3wMqt3EKIumfzF3ndw2NJHDkI3OHT
rlRHcUbWmJOj2GChk0kz6ix+Nl5qOmYYesFgF67g34wnXz+QLW4JF9oMZzVb/MYt
RxFquh//HXknGNrjd4V3RkYgV7AUeVcgB86nddcDF7Vm5AkRV+rYlFgSqVFDNrk6
+eTd9F3mxAYZFotJRh5j6McrUkw3gGn/79zEXU5gv5+4EOwX6YdBE0/u7r7DSEoX
g1meH8iO3RUY4XPQiVDgnkgPHJf1IcNX/OOcpVEFimIg8k/A/jvRyfEX9seFf/xD
rUcBEb2RoCXqhe6jpA18pdkAAyl73uBWAl7AOh3o+rLS1ExOMRWNRWliEc/C2TcD
JKdcFb+VMBqo3tVJTolFJ6kHjLVOJSVSlsJS0VPll9aLMh3c6xJ/sEDuyf0lMstb
xkYkBctvMeyo2Ox9KK9rBjTkJdbRnmewXuagMybF80vDtJMZV51Emn114tjuJULi
6iDRzge+KEB0SgRwM5bOy7Ui/DPjjb8gbutwBH6/HufvmMJCuNoSEC1O7kfB7C6v
zUXWHDwwp53hW91EmHwGbemSlrPBJZ1nnEc671ZG5ODQTqfmEMlP8uMJ7ujW47Us
5D5gJ55jXoQX/4ZpV3dKBPCzz4XAlT1UGQZVvBOlYTaBPv1bncodnt1OcpbkKQkh
i2DaIK8BM3rxvQNMyR2MLgOQV4IVDo2yf1hAQNKIjiyEUe+TGTJpLal12TAtVgV0
70o+SqTFJoCuRU1EXlHWeWaXBRiMREsBpRiA8T63ih/X9pSTVqs/lxxY8/r4Ionm
3P0iGO1KIukHIN0NDtWqc1lLDOACBgGaGEgnmUxyj9oa7Ve8HF/qmCOuHt1vr8PG
1wLdpX3uVfweTKr+6Gboy0XBVAO256wTPJu6Undd9gJoCYcwhqpoHszDJQw1dtNt
5pY3L4M1QaAJu21whRLmvOECmNvd3Gj0pWZJ0667LNnAGBprDwD2ClhcS3k6yk35
a6mkuSW5YL03STFdGf9dKRViibmCBscOtF4e46nZRERXoEnuR+tYudQkOm/zU3Dx
bUdhivsvCXDdEtd//xj7QBRPGgSZtNMvF6FAGoo9sXwXXIj0RIo7bumN+mVogk0e
cdmLD+jsZNBaDgOUhqf6Yiknhso3lFtznpt1Lfk7sW4Kb7pI+uI3tJ9B7Lsx+3TG
irehwk9v3CI5HEQXZoSYFoOgp2jkGW/vWgfMctaGT9E8XPeVdp/6TUiZuOFjG5BV
5ZIded1rNdc2IV/CYL9CiGZAA8vjXtduonEr2FgwVy+05/VAfTGmT7Gmy/8hPZwu
NE6WCeiCtlAYEFCUiAP8RvG3RkZVFbDdZnEnRSe2LmCcdH1UXTBHaA5zN4vbIlzY
mNYr7EF2+iALbosKsp1jtva8SmK27CjlQOUdEXjvc+WhKLCbM4OvRIqiBdMOGpOH
XV/av3OlOoXhZ4F9yTfi3MFGlbLIKYhXJ5qt3KSoRZAtIfNSu6QMqoeEnKti5kjJ
ssS83xZfQw0ME/hzIWSwC1CaZp7C5QkzmftbMVy1e7bXPxVcBIjtKCbdfzP/8OaF
KwvTL3Yub7R6Lv011utSkrRE9vDO+RAbFhZMLwnVbtlmej2RrpRt8HBG6Eq4oyp6
DYFm9JefVx4vDzXmIznTZCfUHGm/SY1jAvhfHrQ1Wag42cSYertgJBN19vyum72U
DD3Fd+mHjKVzYLFj8CzXLEninslyCdMD13SRrUT7EfIg2Vvbub7nCjdVq2SlyjTA
EIQHKVDN/X0YAJivszISpjIi8o4X0Rn4JVgXwWlSjawtYklg+2ap2Ss8paa6XzZu
dONyrSFjkqT3ODDTwjaY/tLN9NDqOyslPxVwiLgfrGLB2Kz9u7DmWQNxnb2nx74v
Ds6r43H4saCuQ6Lvd5KeKGC0PZfgej4InVAqLiFw/p+aOv82gv6yMw6zTfyRM7MP
2IQRKDaIUfgg/l29hsedCOUVyy1EskhtnxGRpniNesn5oFzjhK5y4629oEmamGWx
dNIpnv/UmkM0+iYaTXm0+F6um1wl7ptzrpWjcanMVIi1mWVq9eFGVciMA/Vw/uJw
8v9i0CG/6NGS8CD0dOapCL3eNRaN4wTpyu8BN5dazpgnppwo90N+70iL65qxmV26
G5Xa6FYQlXtjAen3SVCUgdD8tdh1rUTAWNCaRGPwNF554m/fdb46nYmUHm05B3ip
Lxi6Kp2q+wkvHNYcP6O6XaV6kZH+WWbNhMVNsaxWDYNj4TrRhrY63ZxNXaIp2HWl
1xozM97wvHnWNL7afw+l8byi5dD1PA/cx2JNqQ74nUeC5ECRJ/dmmQA9BVzG706+
h4EU14nTOgvDbUA5qhzrQu5JQZ5OUBL9lh771gqYx6vDz8zlM62zKionMqTSmITa
OqSyFUaZ9tDxGYLK4StTfzT40UicBuO5UZQFQXpaL/1u8Ie1+sUlXOhN+P8lp6IE
2Qgu0YB80D1wlo3seb7Btrj9fJwsPuSrEeVfZDqktxd3CYxxYeuHSnHB6Gtgtx+i
ajX160qRk6RmXb34RKFJSL1VNk6CiX/HZ4Qq8XR+AGMdDhFU4JJJkJpT30rdq5OI
j87lBoMOP4lOkQbYPNWB83gJ/2ubB2f/WDOE7kWOzJRd5Bqsc/rrewtvbHOw5HTg
pJys8aXsmpRRKAibCFk2ol3CWdHH11YvzHlrbU7C5C12H6wUlOh0So51IX32RVj5
u8RRQNfB5gKKcb0CaS2YUwubXn7IfUG2S6id+/Lj0hYTXlib4OVfTIUGHm+9UEPs
5mG1pXGmcESF4TlFpUJTY88rPm1WYOHeVtSfQdRBYL9PJBJ6Rl7NzLsmKkhrAeAi
kCUgw1HNiZwddx+WSjoiwILELU0xA3+5dg0A62/bDRDuALxOaHJSx9mLEItuX+BZ
1WjPUxlVCBLQP3JuehhtVItFVFUWxdRS+wQGLygmOMPFMMACwvX1cgTHk2eIPCi4
w1IIhH7f5PtBrgiHcKxzrYkAALYYRMPYZDLnaYnFffFhZncjfAqqhRdDoKp9y3vP
d3sbQnwKzq+iWsL+UIn4gVlc9bKiA7gZtJ0odLKSLW8rJ0RQqGDD/pQ0P7wDCyrI
fqdsNVlDECqKUvfSAbcO2Txa5MoaZVfJdhknAvPmit2PDwU1rxMVnYCalTkas4Mx
2hRhX3W8wdIenjT1r0HwZjkiAy/Zvz6afHNwnHXkKmiGUkr6eAuVfPkeBCJKbOBc
wMLFTx2zbjeKo5vbExJWwnP2IYCpzH6/7YlaM+mOjcjW9YGu9BWODo7cCo5ADpKT
3KwxBSaq0Apwdt5eHsSttnQ5kihR77ufeZEczWhmyIrN/gL3Y2z4kzaJ2m67N4oi
yKkF8tt2O5hUqphUfMCzE+JBmqO716YDuKXgIONlhIoZlWabeUCZ3snOkkEOEnh6
k6Y5R4zu94wZ9pd+EARdHoPP0ey0k18lnNim7yF+57TAhatcmljABhHBMxH7eaex
6VvP41+458U0KECIy54h4BEiESVGCKxwp3jWaM9n0RiZLiQHVSAIrEDF2V/IZpZy
v3wfAjAin4NwyGQzqzz5GfUWzVwNaHhalT180f8GRBjlpjecozkrk+muanw3FDVN
QoZMQ6eR7xKt6aMAJ+ntcg346iAVFgbNfDKfvqHdu3yHGH4HXOdboVSIKXg60JLE
T9iK4f5Hxh19GYIELsS6mL4qioeRkBOBLuXAWLdJZn1I3JNjMjtW5wKizqfwoAGC
OtnuSDmc7feBjmRmBj+SqpIuUfX8khd7iygnj+rxT89XFeAMRROD+VZahPVwQzB1
eH2i1FG8jLH8GRi1szG34VBH85+hlXDDaAaDCf2gVPPxEwYAwzf8MpOeRdhywU/T
cf67sn+6Q9GK1MHY97kNs7X4Xf8geiFRztz4s0L56GJaelNoz0k9pi8/0m61kX7t
A15tBWrcLz06nvxGKEKFnQnTBJbzq62yqfqvJ8HN8EN3LkoY/rUMKLgeUqWI1GLG
2XBHdbE79Sk1UpG49dSS8cqEOaetOljvBYEag715WSE/dDUWVvYylK0XJyXz3nbb
APb/fyAtKXCxPP1Ua5bN1d/+9IMJfIkb2xAtNfOxIex6yzn72k5+HCMGja28fcVB
Ks6IN3SHME/JAgp4dc3AhRTk7KmspMPz02bJaLNKJ6MGLr5c18QZmouqiaDDHnY7
6uRcpKVESAdXiCMq8yZEymjMaV7KA0/zW1uOF/RWSLkAoWNqB+vewvRrDQKUiFuO
YDZ/SxoJoqGsvfhg3eDFxtrq98h0atbNLFQgknyPsqunoNFWIg7903HmyH4rAxMn
rDbU6JOCuBt1+EUNERfO1v5QMb8itYwyTIk+X1tysbW9SN3X0HAFVhpRD7GSz1XW
+Y9ZQRFB05fpupRyXjLfrAKyOr9vXGyB+/bPV+XQE1Ia9npvpgZQ9tDB/ApXpI48
Usmjh3zMuS08vBeyqFYxzlCRaR9OLNkPnpaYvN2R2FXC4ycUe8IxhjmB1ruwA6dG
HZ1NZ7/7ZulP4n87DA9A1Q8TkF43OVS7bnLALsxTIDCiv4lKY/HLJIT6W2aJtIGU
/zPnCRnmqHSLpujBkYjTBZN3cT3Gv/sJVWams5EXLUEEnM6YJk9T95/NYV9bTeq3
4iSoI5R+4oKYh9tNCI072sKQn/kONsxWBTMvprMPuZgep81aGvfQxUSmYuZu+jfc
FifWkO0hxVtIciPgDeDVoCALoKcVEx8QUjjanD736ZaBFcTeXsRu1+X9QIcO1yyh
X86MLxA8qJy2Duqh1NIswZamFeB87i2O3NqOVWx+SA/CPuDaZy5yxs0GynlJUmrX
V1ifGyY9FtbCzPFc1Md/j98TfG0+NLhgZ4FgpOHEeDK2oIXwdElv4Ku9TanDi90j
8nRjCdN93sO26Uf3oAQ2OuuRLcfTNSvus98BL9esenf2h69NN2vpc2LeKKcobxJS
e5HY08uLbIQVcHPfIkQqXpESghlKZMK5SBYS54GSgY4/lVtO2BxpA9TzayKnHIvY
lSjlvWEf3NNc4hK6CaT1LbOyP8ZpcRIBE7F6PdlXYbWbMiOTLplf+WXzck7Yegg5
410LMCJJRgTVaWah350njRCIg1sLdYsmsAwpSdVPFzZ/dlciDI25LE9mK1NhUiAR
Jje504xaJv4YQpUkqpsmmzyaR9NSSzpZt13RKDrLlWZK8FCCi2R3R1ryB1Aecb4o
EwCbUFzKW4En8wIDduG2ns3S+8WNiUIiivy5yDjvsSVKk3qs5byqLd+1YZu4mXF6
anptnlpQF7s40MBLk1h3ulaoD18ksxYHn3mU2s8zPrcaAb+Spl497MugJboSzUQr
cwiUx25+DaDjQEJPxxfe9TB4OQNMngu1FkmDHft/b72NLwP5iT4+WngHAn0EhtEX
TQ7UmOz68v7QESwFlJ+vcCTAy0B+QYzzabbeENQpCGN4Pc+RJ6qEbTvvTkjvmRKi
fZB1uk6LItLuWWE9gSdFiH4RY1algJJFeN8R320wGasJ8/xuKXrjEmq8xi29fyua
+La+CPS95K8w6W9hOakurI+Y9VXj0G72/7+3o1c9ZBj/zHalQRVSF6TP4Hb9RpIU
zX5oaWHahEsVRgzBdRvxSNtIgLbVSzAWTh/F7WLHALsXELL3t2r0P2XTr8rY+i/U
VRsNPpdCLwe4U9H/HlIOHn/lsL9r1N24viwTCcVThes5baMSYK9dzWlB1zuYx7lS
Ni6MwpKvqzvqgeI9t8M1EJ4OB5JbLWc/HwMyUmHu0Qwnc8HWstvrogYoGrZbkMeq
oXSuZBiijpOwkmi5eWmTUYhHJsQ7wErkJmbb1DHUTw+lOegXLw26D5AycnsmIs1t
2bEZDd34cSsXL3V9EAbCAvA9BDuF1exjYm7lPzZXtFbGAM5YkhOYuEYs95wLx5wR
JS6lE8CZVHeI7lTrkwTFqDYTdfmcSIhbEOMMrX7IvJY/gKyNSowYLfd/cicDdvtE
yYbCXN48PkvtMkTcFqWygEcjcAJWVPxi5sV1T6NA3uEyTsq5r24oBPnkYJ5yyyQ2
7XBHPJVIRDy3HTgc/iVTJFgWME3bEPOdy15lvzvxtMXXHeN3vJD5tJD81v6SZIXn
RK2YRgs+MpOwQSvt55tuMo6d0hmfOu1UzcCk7HsXWbvmNegYcad6K9VlYP/045C/
WiHrIvYdOeLIue2XSeRxvI/j3yCn5cRDcAL+uMd/aFyEQCzRuTNnwIhw9TNOq9Q6
MgvOfpxphYUVlHlWkjlwq37VCz5f3pCZ6rRewCR37wfwGc8MdRdKAdLYHLhetFBB
ygDIW9FM3/6yAoLAZu4XqJXsTzbvptockubnZy5B0hvq0NmFiraoQwLFT6vaPIDH
4KVKX5I59vk2+/IImfvArNONMXWqVAo+2DRyguC5xEmI/zU0mMhXcQ3CwWyA6cD/
+AxLh1l57ERyzp7knXnjkfvW2z1g6lvI9do4nbVgErAJfTE9FDX4gX0rWEFlRxX/
IlKiyS47aoYPFT7Rs/TqYMu1ZU52unhum1WrUNBvaG4uUMDixTaHc+aP3HXiLsC1
zi8d8IZ5zYRqt3tc5scT/YjPuvV59OJRE9DB+7+8rQE0pExeVGp5C4dtKi59s8hP
6XnDov2Y5wMyXVA6Cwr0fSE0XpEzmN9Zcm8GC6hdoGMII0kWyYsgWHbS9ebqVwav
3N51/7oPbfZ9N23c4qIfQG/r3yeH7oshD2D+IlMQTNKCLUd8pcjac9bpIKnH+xoZ
dfD9RGE5Cl6z0hP+xnsiE0Pw3F4L6cLR5Al1Dbviwzj0xYl7RVNysn5Yu0FzMfEO
uQzuksRPEMvbk7LkUr+ZKY8GxkaY6psAFeYRsL5XO9A+yRnXdNDjH7pqIrAlWzas
9CuC1UQmFIrB9IE6IixJS/cHy61S6qeVW8n5gWupcVWhM2WVhhjsmQHZ8qcq4dol
eyxNnxtbDO3p6eZPwd5EQ6Q3m1AYlvTX5PHyHburhaP2rwY8kFhe4hzo1Q3Qf9s/
SFehqK8tDRwKiFSvTd6h2EJR8j/RzS81f1vXfEKYneJ3qq0ck8PbqUWfl+cbG+aF
/yKMps/3eL3rnn2yup0AZ4eD5PeFAWwGxantyArWwV4s5Lp42VsSRrSnssCmENRg
s++7P7Qv9q52FcKj/UhFBr4HRPLE4zxeZ8OijnFRkaIzCwJB+7nq8Sn+eIqA5Hjf
u+0YhLhUeO73fVBvIId5s/v4KjRgxahkYoi0BnbjRUKLYp/UWel1N6bXP1ZYr+fT
UyPKFv7W72LgoSXfQvLak3nn7CWwMILOSu8U4iklVVq/dogAdaW37U034ik9V7cJ
lLkoiTAEnYf4tKGemOkPuTt5fDWY6BQtBJ8F4iYfSbf6plEqZpH5N8U18pu2bDgY
FcelGN7pZUtXoadZTObJDaepLW/6fIxQfr2Yt08JfzZB87IbmEYBEPGcXrPE0jTT
W6zAtvCY5dQTER3oD6UgbN1EQt3FOr2+ygXqnfXMOxJ6/vT3gXDRFCfehldWRcOn
PA0rdtBu7bRde+JmPJGTvZeQ1sFkYHLJQ9RcqIOZMqVB9Xbl+IFKbULOFbwlqxUo
lLfENyHw/u8qUCHFHiklWDHdTQeQ4I5vretRY6UbBPGGj+404k3hCKTJZIaE5B5T
xV36DtaceJ/F1C6VMpn2zVSE1liAUK098kF+nEw9GQEnqQtp5C9KFcsuF2CalODh
09aAcQBRyI1XNjoYutByfHcr3FIExjWBVXlUKITDtjByI6wiv0BCXjBhAIVmwzIL
nWaqWkjZsxjWulbs3W1ONVDXITJdy6MBoSH+4ubaImoEThBdLuoGlCgCpFS4qfVb
lr8IsyJdLBUjMMgW/ew9+kyg1/eDnvRxy8226z5l7dQPCZf5DaAwNsd7ROfY3pqe
0yaBYCCB0QlB1lIOJg3geCPORwtCj7U2yPz+ZTGEOMoy56nFevN/3NLTuvAy18E+
+aPla0cWwF/8BdZFReqRap5solldC/lfKD4p25Eiv6u1OZ7xbZpFU7BEiFrwRHCN
3cnUZHJJSl49jxQmsu+HC9HygQK1n61+9v2fL3syVnxmjxXsJEPyYCFXrjrjofTn
TmCxIGvhMJpPS4V1OlLWyvGKz/KxxfTN29Cyv9ee7g3+V8WKWkW1uhooahM4TwPg
yZZ1/12t3uskTS9w3vQnSkttrnOTPzVzHljZduVCjUtlPlOwNknO9Vg9yUk7Wo3f
VZcYMKCCl9pPEbnC8xnzNEiGvoHotpyCAq34v5ImLw/o79v0y0xVJO2Gm8axyK86
ASJhw9yfSXu3/enOM1Q8HrVRDTv+cje204u2Ut7EFblJwXoTWZybvA18C+1Jk4Om
u99AyPIQ/AQ66ddNmn//ItTG035TTiCl8SlvZ0pZRFa+BnWyY/9WNFDWNaveIFRw
7REW6hccLrwEtWOLJassLj6l6yWL+LRsYJew6MAndtk0yzCIkAEjpPfU1ffWSpIw
Y3yrDFJBkcU9wDfinXXivnxYmQTAIfg1IP+Ov5a/y95vVnYPe7lJiyv0IeDV02A4
QvoHmo7Zdp2IfCwPxKSg0glaDvZqk1snmtBhLDizURjJeoko/zWi402VleZdWWjX
sih8lPMqMGsiZPEn3xd7oMLPekFBPBVDrGuc16JBi+l848nAOGMERVVR7WuSbZyO
4EY4Hdl7kLNoohxFLE7P5MkswmzzjA9OcqAKFYyOCFNDshrwZs8W7T93NRfZja9D
ZFBLecx92nVBmyaTZIyBAmZzBIzDj4o8RRsEBEnedxOz4z+tV7gpbcu5NTLL69Xh
j53nF21qHenHf0zqSkhVOOUzUirXlHEIWuhzJnxjN0k179fYXqmeljNRT0uBS2zk
sxDenmYGDkp6FNkBh22WhM9j0zSM6Ttfa/+gfx+ii8QW/c+dwR5utcsXzhkZzqWe
IFHeg/6IXhKbl8HiBNTDarPu8wu547KnmO8+7bYeTMgrx5I1Nd54rtSa4w9hKBtE
SMgW+QhmBnze7WuYU+GYew6RXAD4jAZFHODJAHDsH9VUV9oMMGMvZNj64bkjjCBF
K6bkUK01KSrOZBIT657o/imxbWSW6+khh9BCQfBKXyF43PPh+LqQl4U2t2DLXHrq
SuSdoXZ6DDLwGKSap8+L+8nSBcawqIslHESqTqtS/MsrISuNkt9jS0J5K0ljQ9Bq
hRb98LhTD/FGZ3QZ2wgxYNtuGlACqbPIjun/8S6hogZ9DvTZZdKVj7clEqd0X1YE
iyeKOgsOF15qHt35OCOt2VbSTmWsk/zmYXiBYgcLUDTlT78VJlASdiLKlsyaiCdh
DbuM4SBht124t0EPLDC3mYw457Kv7+7t6pLzbGUELMGf/b/DX/wDR5XLcr3zYaKy
+fpu9vl+i/KP1SXcRZg8Cj9g5XU+WaurmpTLFuZg1WocQL7co+Is1CH6UFV/xesX
q6nQyvbbzQvjs5+lI89WkOyaBn2SIUYppDKPxpt6aZalkOwXzRD4NCOLOyWz9uKa
GPenl+PZHNZOzvdWsMWrlWmYFc5S+FdeIbUJ7a789L9/KISmBZyjzWMbMmSUNXbq
7Lrkzw4LKvSo2c7AhQySXj9z9Tx8Rop7TE+Ee+aVaZcJlanMUPtcFQzo0P8vFIiY
xorqt7REVQmnxKlSi+5ymqcmclW6kkI4KyynowSqk3jjAQyMeTB1tTtGovxiY3yf
ohruidrQNzq1yq7Dpx2Mf4m52wBSHzM99Cau1MHOuILM92GjpSd7fbElaBGhHGPR
xha1Xs7gz6s9UIM51Wgm0ncCKKxpcdISUzqD/bmEsQ6BFclgensWG7SWzJnZFFRV
M/Q1A8HINWFWqVWJOy/sKzcYpQNXH2KeWzNrpsHKtyRw5EFcrJA+GDJ5+IXjVG0/
PkgTlVuk6T8p++/enWaw1KpTAPiDsX80XlVlRKUFqXsReJKQhtq33S0o0quTFu6b
ge7trj8C5kkpZ78Z10NkjZK8RAQxqKUtEwgl4wCNPe7lZDYfV1YdSbYmfj5wuIBr
wlXuFAtuGNIS6g5QbCi9MfbUB3z5VXNaTLi8YKLfiktPwY8jno2XUeZk/5cNPfyu
dIaqk036ZfZa3WYot0ta0JLwMS46BrQDScjUlRH4PtlG6cYb5BCyHnA7SIGgQNqr
q08bKF5AEJnGhnMuWbfRPXVuncjTDGzXr/l8srWkvdNNRbXO8MBfdh2S/ycfjwqL
yd5vzZWuv9lnc4624LqY0Mh6u8jdIcHLbWolIwXw63hnf63O5Fov9blZTQtWpPrs
gq8et3iYTfJe5k6KgCjTZOXMEgKdR1S1zHe8w87oKH2t/efdqPCE2KkcMa0jAwqB
kE6rXf9k08HePGc6xc2EeUPi6yRBrmaNMdZbo95j1twSS+iZv+oQJH7mUmIBTvqr
bTxewp9fUTqIfBjkLDLKm85sRYzaWUZAYuaSClVbkBjV9ymxiRJ/G7fBgk00ZBnJ
NfkR4RQPVaRv2uo+Mma8m4tXgVYDrjahEFr7yaC6vcFfqg0UNF/NpwGRXtOa3qqV
lpqFqQNk3ATGuibNTFkenSdCVxV/SIyUKoqcAeNwR898Ib1XymHHH/kdZ/MBfMco
Dvcb+9nNnHmFRZkOvykFQLjmeOy6aQmWnxesTGIgx5ngwxFitrlrIRsNFGqtotgT
2w00RJLGINO0OpO6NooKchSdRlybasyEWyn8hbvpBGJZL1YV8KDpmiyrlpA4ELWy
N6jxuucYKSoM7gKoFxwknON9O5fsYU7jUDpHLqT6d429yCmar4gtdOoK3ftFb1yW
Z/qi7fAu7qmm3tmNARDUiT2co6wCIiyCt5f9BzeIEiyhRjHjekL24WaUVyqZYrdP
YOVZr079IK7rktL4vaHJMNVh/YezLjOmepXW11PzMhznT9ySgRGKFgPRMZygPJgD
DQdkyM9Gc4jm0ElU9Gr19KCodtFR/7LvCvw6j603wFJHCWzOCyCZ0RWMRoxOK9+I
AHBdT5BLlnIlkxq9idzbaIZgfJrtEIADHZMgpNXifLznY39OlzzXsa/CAR57sTmz
5p8WLxrdFZ1RoiVyQM8PKbH3IWmdMmRANr8HhnLIZP87mD5xBEnfzeGnOYhcFbpf
CAkkBu3eb7FTZRrcz6NeJjKdSzYbWb9N0STxZjInje8ckcVaCfEvMunTGU6wMCqH
tRLK2fOfnLYnrt94yaJRNS37ZVaafL32ZCMM/I1br2+xw+NrgTZIBfUpFI95mF9E
qnqE158+v/9vrKT6hgHJcCDW1t9RelqY8Q9zRFd/2WghMaTwoDZxqeUbfBIi2CV/
1/Lgn1TORI/Q5i8rsCSo7ELFG3Xo5TY5+oSKU+cFs5R7rFnEhbVq2/y/63vrjL+g
jcVYRN0M25BrUId8kKnrTRE3Ct+z9zoj3z/liG6bGe/OyYHMRd8S2oCr516FU04H
/Erfb97LAAFwAbn68wjwqH8QNFPcp5qXoCdGncLFQcBsEuTrVmWWpyZVQkQNhchU
qOMRmkjyOwuTKLm0EUseXsOGoqjUryAozBiDpf132mCpwXAj6n+pQOwCp0Zuc2Jv
24Z7xjI65Pj5syl5elzL49MFVT0eNSi93RnmC+CcB38E2+/eBnDxSszo5OkCe+J+
Nq96EvIEuuRPG1XhhHmgb6DP280Wf++ADn06YnALz7KkXAXAdNc2a9Vnvp5nNKXv
BaoR8tocwshSrQBJJxFC1+ccDnZ/y4/RGuxB18LPZbq5qJL1/skpk7X2EcqFO4VQ
FvnUD0/qSkZ7ILqxoo/Ca9P21MoQMLJW3B0nePadSF5fV+K1n42wGSf/fwgYtr/M
ntQv8ogn/Xf9Cf60pjzX+gtFrzr4s9kpiSZ0ONKjcA7wnMElQ/uNt8gSBEYQF4+B
7t/SJQ8My46IC3uLthyjHQNPpRhjiDOLltp+5Db+umpJ9A5qYmLpznbGsBZbnzbR
ZzM5NxUm0Fc0taMp0RhScqiqYWoodpDcXBaV1nMbFnyt4GhnDIsH9V3oW+bNO/Pd
Z9bxUf7U/SOvt7Se9NS2E10MNzpV4jIjezRIa9oWwyRbZa+mAfm9qaTs1XAgj4pL
UsZGhR/jJgsvCzFdRG23FXucPuiMW7pFYeH4FC9ICF9zZdP3blMpar98UXOCptQl
8EVrXKudpNy+O2EcipNgfI9xOet5m3v2o37P2EeW/4dnIbzRGQCRMN26W7Gt9lAx
gWBL4SCpuo0bQY2F4O66Hz0DeMRCwGLLsC+Q/Q8Ot3SO4UW4FQB/8stV1nEPHweT
00vdJAzgZQgRLI96e+depuP5SSHC5QW15EHmox6cKlbGLnrWJ+5SQ7n6s0c8pXrE
wgoyGF+W2LRQOn8TDldCPi5aIMFEyF7wMAO6uQUedhLgJlgeEFURJAx1yB73f/GL
rQENJ7XVC2cyoSOTpHZFst2cGa2+jkBfTgk3RUbEYZ2rhtSZTqhbxXocH3Am55wK
oQR7t3iHeb0AgwBsAnnjvRDfl99GdtFLvtD7pvjRK8IqWbjR5Jj+yCqRUZZtfsSa
yGkMDA8Lg3MhqPr4agl2hSF56SHtxYH6BZjYr5wigJGzamf/8xlrNwvkdlA3YEX4
XTo92W9Yq8WRX4obKw+R4hahgq+puSxey1+Of5cZ7+4c4RpXQ5L19wSI39Qiokn+
5iegYVeWplI/SfquK5tDm+DjOyQwF81LdmgCaMtqRZXYcaJIj/2LetqZ5/9FGWc1
dzJfmm//1Oqfy7GFq+7DjjVMzBo6YZ0SeAZLe1/UTVc3auT+5e+ZFJ/R8is+Q2nh
hBThRpk2DG8ARY/VSXgXUDfZjL/fJxfMbkNWwTI5QQelbFVQMkRNMTbrnwM6dnn4
vQaNkCNfwO6uQIlFcgW0GEes7qAyqouu2tJfYiqoKkiTxtgfJmc0iV2fmIGB5ZAo
9SkxEulAy7xmDW9SVkNRE1tW0zapxu8/2KmeGsi5OHbMEIv0t0FfdJs8bqBvr7qz
6Qa11bC4hUIN2dY0nEgwZvQVMzTgh/NAuZARoUVP3IuRhup3VBdIHv9GvLB0fgoh
ZcK5AVKWGuzbqkunxYZ0wVWRudC1Wr+YwaIN1UdzrQjwEhYYxGdHghx/leMRzJEi
vK903r58HAY5i8HDOz6K3Jc9niSHR/CJIZ+I1hgbG7dk5f/0wl3LhTT2ytIc5Y4V
rcCX6Tb4eZ4Z8dHxpgGtgtWSN7HpCmdODtmNteuUmM7Mzhnfu05hdXtCXQ6Cd/Bz
nk+7ljF7fIC/rf7Gq4OxjHm/1vOxjCF1xtj50EHDAFomymK2g0sP0i3x61TZDfqd
lMUOODBhxZBiVWv+o+uCI9NAWWWH7P3UFIk//5Q7htZMbcn1rKJpRor/aPeAGYgt
M7wICEuvRkhgXXIVP5HgeJriLifORx046ZFM1hhE+SikEirOkTYZlRkNyrRSTtPG
jHC7RGbqr9XzD6t9n5v81faPFLzo3RO0EFqlX4jZMcQMqHPTcDPoMJyykGAOeoqm
ERevOUpKWSRY58kT9uhVTfYlV53/WfLmU1HukrJwmZLug5oONkjqlwgsu3nZ31xr
FQ+a91wXjn4rtA2FZrE/ED7BYATDNyNZSSdQlGhKN/F1wuU5ZkHVYXMzjQkwt73A
BU5wIODTPeaqRfeTTa+f8r0gHaALommZMqPcjts9+hrEsnTMmAFJkOCKdZXVzMg0
QVSi68iOrIexz4R5AQgVwsm2cAuz0r5O+ZtpdyyX+xZVf001ejaGjTZHS35scJLA
VEwJPxcfujvxR4DhmpNPNaJ6VLDT9oIbdDZWmxb31utTdCB6Rye87lDaAXuP1JxE
kM5aMv3n0HZjWFaHFajXKGKwvE/Y6Dz0OGOeIYWXCkCqaMYNe4EIP03VTCXf6r7P
2MwFTY25W62319znbtxiwVwG4rJQJ+7boegDC3ssGxKOWtme5Rv/ApG/Byp0GDQS
5N05YS3JxyO5VXeqe9SvLnGTz93KsZ3OZ5xp99mQtI6E5osgbdWLwbsxeAzuRmE+
gzfauNpAeuDFdojjE6XELFzHr7hbHYK8mYdKUhIeKCAl0Qx1WHkg+FdmaUDMhZsd
OeQZ7zMVoxhu2Fujn9XpfDKnjq7y5WE33r9M8/0lgX7hwh9benVL+5bWivvZOMpH
8j7HfQQsgohpEspwSkZgtldL5raAm/Pz8RtZdYNm7cZodmdfpN1GCw8NK49Mnz2C
8Y172b8HnwXqd4UheRrUGOPZaMlnW8MG1DRaLwFB00Lr5sCexI/5REK/ij0itE3O
GcdqxUZ5crrW4LryffzAADeq9+M37vvoGaoZlwQYckw93pBZ0jf96fWqMVmnTMmv
k9oOp5hvkMyeqoWTF9Z94d4G85iNedyDsEB5UDj763TVqN/ScQdSspQYUdAVN+ZC
ystUlRwUO5Wmv4df7Ej9GH/KaO3tcd9W+gD+UFalSyabV5YU+YUIu7+P/jWzJDJO
d46aI0UaFnpDUGSROY5L4LZsjGPQAn1zqrj5bjRD/aSw2/hGVgVwJagt8Uj1x2Hj
UEOtajNk6OCdZYQVWNrQk4fB0i6lDRUo10oqt/vn/urHYC8wSjoGi4CXNtu7Rxoa
tiBxMupbk3HUQm9wax1QIw6JwFa0y3VFbB3AQB9miWvD2wRi2mSjStsMVkDyyD2c
KtRGLoXEm7ejw4PnJNl2UHidJOuVXejDsuyYUyPwCm+Tsxbq4VyXuk0YGWvn+3JW
wvHVE9cMpPiTGJKQLU93veDQyBR6VqhtuTnxdHbpWaB9wMvKfc65S8C2YcJxMhSf
2z2zW9BLgaTGmSZ77HMCtlO0SUgKYe2Wy1icGEm21GM5mE6yOYK9MVbpqSGHFOGO
6Mya/w440P8wJC4vLXYpSBTKSpzS3Ts4K8qYjkbreBBBip15H2qU5mvJU6KcqfcS
6gmFmyDZzlH3Wsb82v/ewiGz7jQUvtrktMQClJmTLPya0tVUXRKneIyLH1FOlxlW
jY0HYr4nf65CKR0nnkXzeLWduwpRzgEkRrGoKG8/qlnGjbI5bm7LNuxfB+68yTnG
MpjOKrxtsifIZR7nf9EZyGW7N4vmNR+GP0HugUz3kN2expGljFpeN/8Ez8rrgsMd
eQRoHhGHSx+buc5gAoqZ3fPtBg+x+ONs2DaeSfOiRsEvX0heOMZPYvzaRqoqKO3G
QAo8wqP+onX7Y9RQNA2PNHeQRRtqACYclmO/H85/RgLLQhoz4TDBUgYY14wvhbdn
r8Diqp5d9Ms6uREIYjIuP8iLgE8mM/sX1mPyGDOpdFUDMg+WD1R98woWl9WSsKD1
O0xLpPRMafDC2dIyoG9y7bERSGCQ1xd5ulb0ETE1CEbiVYHPZRHY813L0os21WBP
6AmqeBv7nxCLLdH1w+p6DPyJm3DX7KmYecLFyJ+73nkmMJfh1AkKaE1BRTLQmszB
QVHLIcSiFnzkoINpZJncZsrzOKHbUoivd9VJEwXn7+ShRR2ou+lkAV36WARWMqPD
NcPtaws0W1gGmI3+h6duWj68CdFDWF8Hrom2NACKPA4DuJRjNWItzDlVsVETEIWO
xe1brGRiosXCHSE6X2L70snNYiyivvxKKDvtq32l/fFWHcpqJMwQrjnnAZcr3Ahm
EXw18A/puvrjFyP1drETOv1d/j7bkcgbI1SLkadR9UzCsHDcQCBxXj4iEoIzDhuL
fUdYDf04Mk6LNRt2FitF9l8SKDwcjlyKi8pPTbqI5eBxBv/4D3wglvB2FRLhzrvk
3FXieYaiuIkLTomvGfN4oOCCE4csrRXSyNUo8H9MZVzUYQZ8qKN86+0lPkG8hw/R
pYzuFJW/JeUJ+XSjw7FpJp2lN8Zh/bd3s3HJp32xwAs8UXgT5swmA/5w/mbGaKhI
tT2aXRP65W16pf/62xWgVIZfUbeVmvrQnyAr6lZEMPpjMup+8B/oDRIi4XwUFpNs
E7JdjbB1RElo/77fDCaBfrYw/i9rqPzrtXPWqFUDtO6lYU9+fGPePPPxS5didIYI
x9EJQygx7e9xeK1K5r1DFJ0LTC8Xn8NwJGhSlBbi4IaDRkmvpG6PmrdWJnppZRmk
Q0GQKFWUFFojt+cSfXzWci0ZKybrIOecYyHaGiLqbPnxNXabhW951GAApPRZa8i/
RDn13fr0hYahlK+kd9cztWdzteA+vUPJLgD5ME6ZbUDFRnfLE6OMNBI+mJxDufYT
5qGP0jnc9pwgT8MtpRiEYgcar0abrnyy34gdatOEJZ/G1RFsw9Lll26adYsHwQ03
cczC4wVItrsTA2ILphD8SSQfCq1Yauj1ZxnWF4ZRBq2g/bzFQxHarGOFtBWfNZ6h
/cPUd7zs8tQ9Cd9OPnu40MiVCx1xnccV5BVCdfUUkZ/UhvhY/2kVnStaF9SnId+D
vJZ5xxaCHshtzeAUkTVrTKTlZ2fB288MbwOHVFVaf0Z989ZAlwKBHPFxSYql4EHx
AFeyTmAQBDxvPR4ALfIk/hMXiS2LDd09haa/qB/fbw2FLLiqrubAv0Tw9fnOkSHr
0FQxF3gMwsNrvF+dwQdoMh+YReEPfFaOolSdPnVO17zIxajNxHrtySX/8YbuDp+Z
3BSh4WL/KYsfNoSUm+Wo9IcqaVC6EFqwwFnVeoiEc1M82BzIN3Ry4ecxKuWC0K2k
1dZaBUFyCTvaEuwfYxXncXpPRxhe1vZL4xWeLfoQrq9K3lFmkvLx1GrOO6qQFW1J
Fz3aRLG89LGPH6JSGr5LSAjiVLfZradIkBCe47p8OYmoQihavDzUA/HRkO/OEZFI
Ck4OdkapsEPCbjoPNltWq1FlULPwsHEKQ9g1yUCbKcfciNuPqVp9Uf5yrjo6KsUI
G052g9Eas69d/aKOp6r+IGbARHQwlJLSc8Lcc1PstTV1pksTsc+BfLVO07QfSVUV
reUKwPmTw/Q0C4bu4cXotZImRG8XXEg29tPUUgDiNfAzwv2nrNJUtFEaAw2gXRbE
My85D2gazkjAPFSHznm3HHK28YtAjXQOmVS7ZVdi19wI12d0CaT832ip2RmtbcES
akBHLCcHMFhayMxKzBy/id7pu+CeJzPRfCT6SHKI031HVMOfBmkxaIH/TTUh2nRr
OpphNjR1owX/MVBAbQuKXWT5cm3JZItmczepbQs0xcCkuNXQ5XFwkB3j/mPsQ2kV
LcHp4QK3+UmseLfYlRLDTzUcouXoiKxXMPbPCzbOv5LXNAS57kLqhroHe5q9344W
BMcIqI0IlSoEyYR6CFClhYV/hC+8fOGiMcXQYvRLnl9/1szftpBf7j2/wp7vxvR1
hhcZtDAeCHdoYsosRhpj8ywpBwYUy+7HF4Qj3+zTSZicGxm3waINbUAshZIrcLkK
HMzJcw817idNi3n1ohTny7tfsT7O/uw/FNAfxU4Yn/KchGsAUz7VxF5wE4pRCU2g
slQ29swCfS+85efsjMs/5hfvCMbZJcLlCXc0A6rUXug9bqdWTn8TSd5sEPFX0Vg9
jzHRHLCqGZlg0GTjysxm/z0ZGv2bjVroQK9u+uZ+O6CFPk3JkzWEBtfDF0SoFpnB
j99M6CSzHpZoL41vXvcdYvcoJni7pepfRLSZF00dGp6ySk/zYBxvJ9MndIZIP7mP
tnhu9bLGiZk00znhD8mbZ1lMwY3ENTxDGPDs60E8qO+lLvdnlRaTXpOlxhe6T0vo
kaVm6xRdRpQ+d0lCLCWLWuPsjFt4jS3ttcIUHJrN3s/82eXUVWlwzdSQFyQARHcW
DPQli6rx5yR1/D+qrcgkGR6QSeLGT2J+pgN82jtxwpqEquM8Bts8V8JuPjnzYOts
gj0AJX2u947354rFeFgRkGLrwvoTHZDVAQcEz8AKQD6nY+nB0eyB8T8Tx6TN9f92
mxS39FrcdqFkgc/noXhqMVYvTVenoCuBHiHRdrII8gQDEcwoFTcAsfPJMN9gf0kB
/YHv17/V/j/ifaUekPaAzI/TfKY1tXpsFgW2/fZrO7uLxIcydmZs2EJdoIwSP6W0
lZY9cYnLWaGUQ8b9ZCoboCrxbHJPGRwzpFk+be+Y4pPHEHq/NKMmWgmImJ22k+ff
LvoPQ6asHCGmmJgGmyopSRgLo7ck2Wz9Jfi8jeEs4dKeAZDbKJMjserHh65rsu0t
XKR+/56qraOSA/79PLg7NWbokMllUdpbKx97kL1Ul6mnicPrC5xnxdJBoYswctrL
OOrxEtgWlI+o2yx161c41tQ3wtGJsTs7f6B24dDys+NCBp3g01liHqP2e2i7Vscy
NtwpCdsd9bEiah8ZRwX+zpe4I+jVwbxdCfjlfAZ/Ubz7g5QmC/WJjpQv68nHKN5l
Irk+I9QCMUa3lVK9qZ/oXhPE394FFzie/scP88d/xAM7XSdRAJzrvh/JFvyZigUq
gDrSZWmievYsiUcWbbxh5Sq7L5z7veOS+fpP02aZfKgrbh1Ng9fO0C69TdQ5Zy+1
vvEiZfb3NrSUFe/+sHc1wEfD9OsFdmy7wTExRpxY7D/88fctX1rDfNfWM/2bT3vt
UDHri8HjuHjga5Q6c4Ec6uHikU/vOCs/QiPjMp8rMrPatDk8/eY2M3LeKO6pSmu2
HairZz+NuVBQ4gFQREproGruE2VAL4X4vJqmYPNBNj6jtrKImSz/sLanbl/qzpuS
Hm9Q150WBBoQvoJtpSXFwsCDpoD2bPS/MkS44n0FDsJd/TyH7nTaDc+oTrAdJ/V7
NsLeoMr+8BRILf1sWpRbgJb2MXyYnt0n7eWuG02KKgov57U1vlKp4LTggxCJslxJ
6IHnh2fBnlNYZVrFSdty+Kvsgj6kK0J//1ZwN2VOIgk5XR2Eqq9d56E2XQ41Kjbz
/rj36WI+RJh07rYVPZtdk3fFN+oyN7UDX6oClbYP0qcgEL+WpnpBkr89wsAzhKEb
lCK97Vkfto1syZ6DNZHE0W20SOh2vYIZCGg2olTcYFgpPWF4XLPNXX+N8c+qKLdZ
vR9TGZlk/5bSpE5adsGDfYJfSq48f3trDEj8tFWndtz1QA4f12xBoWE+90KiExyg
OlsO0CPZkyUn+v7b7SO4lbYXH4FIev4rIhBUu6t3eMOWLI5Pklui7EZKuzLUQ4n6
ONm3lTHbOeMpGiX+OaDJEJAPXcVoX2AsPwN4Ge4KBSVI9yMts/HndDHxfDA8A/ZJ
YbLzIYx1Mpts8n9dWqUwyfMqUTmDsih6uNTMCLP/DTTq+eetwpu9QXV1BHo2eFKI
WCnnJt/+DFoU6UeYvdPYh+9IwF4EUkkYPB9kIyIKft27tamffSSDdVAY0IHSPov2
+SvmmhyuipdmzYV67m8mzlN30IF7nXSzuC1jeZ+3EoDX4RnLLzepux39HVVL8rRi
KTVyZxG8GIpKAS7dfw17fgarPvORzLPbfP+cjMF9atumJ/lvVh9LQweQfVbU81dn
9a7ZP2c42oVFNOJ5qyT/M4URzPNKEnUlPoTnDWeHB8fYx1zygStyjJ+pk5Hq+Cc/
42synMV0HjWOv5XY8WaLAJzYqHJdItPHhMM+1iMEcCqtYED6+aiIveaw1VS6CnIb
Z8cZA37Dq1DfdX+8vu79et918rsxZ0dSeFGeyqJ8xoTbDTqjltXPqiJNXT8m0ANb
vq0HoqIYbNoN7JJsGXL8slQI60mYMknxaH4yQ2pERG1lAMn0cTF6NoKTbkWRwicL
E2j/rPEePdAb1cWfzxM7xqnGTvOqAa5aSgWOI631hiuL4xfBAEv+60EHaXCxTISx
BckoGKkJMvqdgYzK5M01kQQij8VNkG72ZodeM+IhP9YfFBd7tnaNWbyRNQ8hIBLu
RoIQxFxNJPyJxnvnAZ0quCpiBD/8/R8O6uqmQnz8fG1FNqN95wu9iG3TEvA3pNMz
5wkFVc5QoZtx8vTpLu2Bi1a/mz7XxoVlvU1xxvA7l6MvxgWvrYWInycmuS4crtxr
QeQR/FmZZgtzzfZNW2hs9fluBnSfuhBOwxDMPgQeo+Tp/tKUlsZkyMpxybYp6Ytl
KcYAeEft+833Sx8FqPEgte5YDhcZAFFV5ZJA54KsG6pxxWc00UH1XLxZ5A1YGFke
NYKMXreUWHIJxSKcgpjbAVthovLujh9ZEXotRsAze5+pM2WAXlbJtSIfV7NzO3TG
q3yhmQ+e6WJy+7cO/l206Ds4rNKJ76ClgemO7xsOBDfWDemSKRP0fXakp2K579PL
1W9NQadtWcv0v2f+AFfdTVYrWRx/Z7HiW88WvTGDRFtiOYvoMWdm/qpeoZV3x4n/
gStlSemFTJkJdq/4UIbu+0KzsEpF2bY5jgwyNxRdE0L61fKYDrCsNt082ZMXS9Du
r+foN/2EyDRQ3EeAl3WdW0O946vYIbA0RQv3+5p/6QFhfacNRFr+uhWEMm4wTjYo
Eim7+nnE6rY0iLOBjR19QOUeTFR/ikIUK3XDMy8mUNfACCtVAiVHptcXmlX00x01
NG0YbyCz9fKk3wl3feyX+bu9cjfwVXxljoy5HRk833p2B4MTsGqug6s/bBkGIEky
BvHstHHmzy9Rzk2Ve0qbKjQ+YMtPRmHnqQja1z/hRah6no5noIfown4yE96aK9x8
Cd488YNm+i864I2/zeW+IAp6+7so259G1+n8BuElI1i0UrVG6wNB/IYAHecslwqa
xICb8lcuHVKent9h1nYSnWLsPvvaLhURDqf3zt07sfdlqV/vmFIBBtHi3PGXIiGO
mW0ulMsBSiQK9r4ZBtgfnLAQqrJSUbQQJjIjRN4KqJEekrEKPoDPWgUQ+e0hcU2b
Z4fh/oXPd8oYffg5YBxUXKqpGgkJZfEojHndOcbJ3xX9DUr5NkQnhyPBuZ2fNcNi
pXmBsbDtu48cf8+Bb5kqS5Va+Ru3kEC6Kr8u78iW9JWcON8oo8qhfdvQYOGSi9MB
SSKbnImbt6deNTvNRJP8yAm96TbZaQIJyYBdtP9nJEdMJ957lvPHbA0CK+0vi6LY
lIn4F1EHeY6HX+pn9+eUfV06Pka6EcbTInJBM45UuB8GFJEjP0/Cyq89UG9O/7K4
Z8oiQ2W5lHsDkVKUOf/iUPzWiNWyDjTzIgcCDd4mWyTmp9A8MCd4vI2Bep/3ID8W
bVrrebmTr5YiFhTDTrTuuxCn1eHKEmXjw1rhrVgtaChmQZ3Dh9ZnUfMnFjl55E+M
nuqMelSNGo8VTrhQxtoH3ucoI+otf8Ci/sAMg+k2lH8BrINhNvvfa5s46wI77ctU
SyXlf/pVAvgxTxSkqWGLzw93dHfhOiiSyJtn+FssZ9F7PNEM6/aYMcK5Q9XKS2wr
b1evSZ6YaMzkR2wyY3hpyWjRD02vO1GvxCDRzK5kMs9246HAj6V29DWMgneUluWG
XzKTqR2xyntp4D1LFr3lQOI1bK5c1hZp7JKcLf0puJvmy3FXl/XXxvIgyEIEzLKI
7G1NlwrUIutJtwIMP/CyqHmqQeEKJCUthuTyp2dIFcUySioB79ADEcIgr7jS+1RW
Wxdr5MOOGxBSA4nrnBZNjpL+NeGlr/FPTJ07CHcuuhExwYtrBnDq1gIfZaFo+BJi
l3gIKiDnkD9bfUQ4rGnqG3w29c0rwdeKJjWdpcfPn8EE0DwSE1UwpiNC4p076qed
512wybkhUQBqyShHXQpI633+r/86Bc/bSz+DgnX5xfts9hMRLW+pWC8UHAd70g5R
G1M4TEILePZ/8WkEH/WUj9+A8KnIw30LPLL7wI6bUg8dxsx/+psd78FYeGDrJ/QR
ViOgQq+Hu7QrlAYRudZE1RkX92Tu2CzWXcVd+Pb3aem03HodszEbdP5+e0NmEy1s
cLnPucW+f2LkoUeTaVeOIZccbmBvBoUa0rsm6OP74G6IOZ8AtxbqoPh3YknBJO5D
5Y0tBJ3h+o9iCX3LPEzJamkXoSXzm8Z7qySdnXvSarG5T1ZFNSvEwaVO8kcUNMHO
BRxb4XwagbK9yZt/k0w0dUhDLGrH7RVCWIKIWLykxNL/4PCjm588/EjRvTd+nx8p
lt/iWZw1Bo5VJyUZbcz0A2IBu2I+Um3IFJZfwW6vBP5V5rE86nCrrsoRw6eEuIQF
aWNws499hPNlajMir8N4oN6VXy3kC6oUdqjZ8+woZMnLRko10oQC+1C9zwEm1SzP
RkQ++GMTw953lFcGxe9+fLhpgyocKakkPPubmu77b5Es+HldvSQD/zeV0oRFaXG+
tRgeMqf3T32gt54KohRaoTFZltZOvSp3X8wwvqgugB9/toFtrO7ig7k80lEUJowW
sQudGZfsbXCdpMSR/I6nSeTT95RVCo6C756nNQUShTl1hF94ZBLxn1BSN27S1eIh
momAoxy6Qce0ySPU7GsC3cVmR1TjYbWmKl9xGJWZH+ZwwaKfR3zhEb43XdOj1OLe
SCiyw45qS9oouVHJuC+mJKlkHAQh1xPlJaXUn165rvhwRStiROShB4lQ8Vy5ddMo
D2w/fcIXH51/9y6FoKqR+LLu8cv35BwK+S/zjE8PLs7THBnUww49S4nwOXzdyyys
rSjlz/nNa2CjTCpAD5D8V7vRz72GCfI5uy7u2xUnm3BPvANuJYVblQreF3ud+bhh
TFMrDDYpS5xB9tTRHjCeD75w5AuxUbis23qhDHz4gcZQbOeDB6SLrAJQF2XY/spI
7Ydec1XJxYolZc57/8e44Gb+k830sGtQyxN3AWa2camXgDzibWz4DAI+Z06AARGX
IxyaWiePoZPPNFpBcSnMJug+L0WjxW4t9sITuU+xuJ53/QJOjoucg37xiTlyLdq3
vuZf31IQ8+n3drBAawIo3LawADK4G3FLLDgnzk/Vv2PcYsgjo8tUO0kCeZjoHJzg
rpMJpLGehEIDc0PcFRFiq+N6//RxXCKhQgC04bsjg37PA8hf7kLT4TS6mI1oxhWI
ytZO4vYwnkSqR33kGjk1liIHitaivk4Mspp2oYZG21xOfa92gi+FHQQ7Ao5mMtrO
fUloOFOPc4aM5IXSAmYMSqRzjstu7RVoouaDsMvTbqRsNzZpJxYNxLZ3Ilx0oK9P
k0QsbxLA55TF+uDPyz79C3k52iWCwXpLtw9DzoEfM6slz4BHKaejyf2AL8rnIDqQ
a/PycG7H1oXQe3Y/ZBXw1wrlt931cEL13sCguTxXkLuBIapEYcGTIJ1wJ+Sm/1Wz
syI2ITQt+rsZnEGtrsBaVWDXaslWFgNaqhvvtl1lwTUkmdQaBoCvEDCaj0Dh6yu9
ROGtsk3LnzXmIhcfSoFUxkHljt//owpAjUfmIxkdElyKns32oHIm/A6CKDBkhbRN
UPWvs6JbS0uNnM7QgabN595T8/p7Z6+IzCAc2XBQXYhhoD97YQ/4ih+X5fnVcwpT
XBWhurl+9Eyj3AC/vZqtHaIo14bpr5pqeS/dqWbK0Yl80KchGQAkLhQ7R1GKw7vT
J3uaBSqMjaoHjp2fkaBvSwSuF0l2di7a85l77FRyNkO8DfH65TPJ25/NZCOp9ZIB
NHsL1y4E0IrPDu2cNw3GUsdYyN4gw44ZPxeGEgfz+Q3njKhTLguTXrYWbe0XCI+v
wc0H5+GkPr8IS2zb2zsyPC58ePJG1s1zTDsoVOer+zaT7rTZcnfDCV+qCqdlbXYV
q7gXcxjtuAFL9Vt374NXuwCy0qrwHSgvxa/ni9Dm5H6TtXmdTWDVhJiIPOaFbJXR
N5Wc2OUBTgX0jGpT8FlnfU1RZIly0fVbTlNg4eni+K9gQ7JYbtqMK170WLYcp6jU
IUmns0F5RbkoCUpFjv+oX81X8LaTltrq6MKtSECwjxjm8R0lMB8gcoQOa/kaLwDx
dlWJpuWBGWHlCi1GFdpDtCz4x+/HJ2e9rvQtD+TDOJOMpZJdmUmXS4eyGPb62jNV
9og8rn5Af5EBgdFL33eUzRX/kKkNesj2Vz4pWEnF/f8Z5DoYgpLGLSr6UqggZDgu
YvwssDQlkIhMfVMVdl0XLI6VloLq2UllGariKTP7PN4ry+SX7Qw1C+yT1b1dEF00
SHK7dJJj6rShRoFTtkieEfy8rAzYyTaOBTrvsQ6ceUh9QaVReKrxYAu6ZNnRYwSs
tl9dOy+QXS+Ow+jKqi16+/DL9A0qGFt/VFDGpPINbQh3TsNXfOECFC/PuKwPOHx0
8yf05VM0rNqajbXs/QfvgmOxcIbhGNeJpuujDFrNljbAT1hXrU7M8nQx/JuxcsmU
EMqX+VCuQoLsDXBeA89UYu8Jco8omKgjjREtoTET7vMCTYd1dGmujCsMDTktUOYn
+Nyhe0vRq8FiK6SJCuWQsPic6ybP7Teu2ARPUBwVejMl/TkxS91omzxfRN52Ujo7
sC84zsMLggiv6RZmKVAaPrEZFG1MFvADZc596oEhqM+p9iJ7C62YsfCY99PS5BcP
fRxBRF1QjBrXiBtnIQd0StjTyfzuKNkykOFGtrDaRiXvQG4+O9aE3Io/lVGsBu4K
1Ex4WI8sJ6ysTO7PRbqKH3+Lwf3ts1BoV4Egye3/fLA6Xu071qOzsdOjHJwjmBHc
uUhw+9pENWJfJtoO4Ok6y8MhzU8lzlsTDWg8b8Sr4i0RRWx47iUQYvzgWGUvV2Jy
xvdO/k0k8a8b8OID5xRIu5DR0HmH6VMEeKckaWhNnG7+39eGqb3uy+z8AMCBbS9R
UEUTn3BM3YcZkLdh4jWYHqVHPiCkuwoXsGypuxbQi9YUYGG3erZ8MxUAsRhEYSHj
IoOM0IrQ+cBujP3q2pB20nPPSRX/1lePccDF4K6UVa8Ub3y9oror31Iui8aBXHKD
7RSI2D2b+xkO7SC2+CcpIWK6kChuTInv1VtZF81RBEG3cMMuiC5n0ODZ4snQ+dh9
k58jyiUb0hPavWX5xjNcC1mSRWi8hM7JREDy94BfsKTMKj8j/XS/z3nes17GGTqA
wXbauXpOxutR1SjrrAq8n+qNekPkxpMAtR87wYAEclzsM2Y9TznhinHfLwZ+d5Dm
fa352BqjMvIXlAD2BiXhMlhIEy+klvzZQaEguX3aFu5YpZN/zL0hMCP5fXFqFusl
7rIc0UF7apaLTLpE4/oZSP54B1i3mXE0EJn/Js902reBYuspeDApujp5EnoOU4co
jqTU30ekpItJHwt67RMGWC62KYQikldOgGDr52L8HNxwdx/T8LibU51C27L0Ugta
mRWG4Ewqp44rhHXpFyX0cHLVRj5sbP5idrJeSwQd1jnkc4/5ocOqzXg/jEvyg2Y3
xg5OeYL+7VUID14flgQWfIqaxpVvQPXkTdynXCvrAqMwkOUEAKrkCc6n16Yhm2Re
molOly2dLBYYhK++Nb8K9g3cwWaS/HwXuVQ2aDh1caM70sA3axyUiD59y/LNtUld
e4qw3ifQy7RjKGd+j0CSVt88AIF+4qJbGO5pPm45O6kaPvkOZ57srryU6h1CQloy
NBq9H0TTcBoUGiwP3/RPsLpLolTGJy80c8UYRoNe+Ly++ndfRd+40uP4q9rrZA/Q
N7OCS5m9HQoW/N4lsEKg2TDgXAWaxqRCtoblR2/29wXhoqRGAbRhYvvvrmWiYeRy
b3deLuKrnhFMByijbgdy9o7Z9kGP6Be6gYoGFrO2NgO10wsWczKLSlFlzbapkcT8
l0Co6nz2rw0dKvLToEemqQQUg19+sIgokwL8ivVd12PeV2lN6UFQKVZ3X6zwq8S2
gV/BzRcpB8S6SltBMi3DbSV9/HPH1yy6gGH6PMOJfKrR7qQCVLMOkJjq+4bxof+V
vB4q8fWhAmPrbMCHyiD/DcD+WZKY8E8G3N7MailVYlGDo5PUDm+yeNrDiG2XnVj4
WS446gYcFZ9HPSYS4a5AaehAeF2h9Qf0eyJy1JHFRQhe81/rzWsUzPrLva3a7l0t
n/fV0E/o+Wx0EXGqZBpznClTi9MRTcB7pgpREOf708wgo+eMgD24qY014v5et12T
x6gRynxhgWbVewp9XBiDYMVTlklTJKzk7FRB2ZA+imgaH0RF/vX5GVhZ18EYtBzr
muWSMTe1LYzT4n4d+ZgEymzKs7jSelRgBTMBqoS/UP9a++zDBL/LmjJt3v8aEmsv
/gZBlsUo1UL65Z10jwEzR6eUGZnRLmTBQZ1W9mMDDQyXfpN6kShp6JVziO8RVBV9
JTzPw2o/4XFDhhi5om/7SeiDGw2w+eNUB47enGUuDmjQz7XYDKPTuI9zQwiHmZEr
oNCrisPB819E92c+HLFmOVrryqNOIg1V84yYeZPzywHBcfMratyTJ4tP4PzWMwVf
f0eddLfNfEy9xnO0cHHpf2z8OTLiX6zZQyT6fqBhNiLSinpNAHpMmQFcpxUoE9j6
UrQu4+gh5pZjZV3HbwnY/dze3dnfWDzjgZrdvFPMoB7tRKX6BPX4RLykmtHCfdI+
o3pb4ciA4PC6r/eMeQ0c2H++UDxETxdyvVSEdX/2NgptV/ebuhgvtfDf35ELQQ62
3I4Px7OCTqnuwcLWqID+Njsis2cD2qxtyD3t3TSWUQ2oyogP7NG88TDpHdo8Kls5
Dt4chKwcKPN1VbA9pnZVt2M8CXVDu7RKZC32FY2bOP/uZ4LATFWr175uyz2m1Rta
KfdPwFi72YzT+fg3yP+cCSqHbL7EpDgLWZuBZQHus9UfQUyyEPJWjiv4QerQcTCF
q2F0WegCkB/rzhLasbvUGKVvYZNCAx7KKYGzE19Rw4WtSnK7/u2ZydcpqhMqlU9T
6MaBM6BqAWXEMM3O60MRMwrn5mlcJyat/jQxSm8VAUBFH2zLEBs+P9BRQA/lKS5q
a/ibY3k3r3TvZv2NewB/Trf5hwmJ3cbL6aQN7V0mSJX/wICKWqn93z2HtHVmGx9i
WpooQbV2JfoJ9miXqOHxKmO7Hdlb6pUgsb3EEcBX7//AXV5HgrF2UcTBGPG2ohTF
kvCs2RCYGe+2Ln8x0T9ASNXkHguK0Tc+wjlhJOfrNMYXNaJvi57AYkczWM+GHi37
313zHfYYsi5+mcUJl+U29RVuwdUjmbYAASaA8LtR1O+bm8G150uPTaxsDTAXgzNB
FEGErrihOjUi9m0sQVepCFGeLe1+1Ur1ezLbpkQICY56UQKwROgGje4jnU3VHiyU
7js9U6D4oQt56zU3IEyl9NiLqgUwpgCBw+be61lu85My8CRurz2GGT2lTKhbxJzF
4yltevaVP+of9XrNvwXuzodZ2ggf2DSBDokjp+E2AaG2YqFfMdcWSqj+sK5roRfZ
gH/lc9HR2D594jdFTYhm/JqGrpg8ah32cRvBCoN24K5uec6weE+QQHhS+JNvivoB
KFIMOv1eUnF1o2eqetk79iziHbSWC/RQc0rQhBV+t3h2FJVHTE1ddt46fQu5XHjg
Dv39jEML85RPOOnbgoXQH4HifgxS/Q4U1mYJDQ+1Oo+yTngY3HRWPdvSCAYUayT1
/pNburWoTuLDzKUA2Jo7w+qSaMgWeV/gSySvN7g3gAmpIsID4DH1iXFSyh4MknAl
d0Zk5KkEUHl1rpjJCMAU0enR46DzjrERImUlfnvA8CORET+GbD3z0GKpBehHZj9e
BuUtCYsKFa2Tz9uBlPkPK4SURP21k1z9VD1NDHaKTvItXCFZJeg6le/knmKNmWFn
Wu40pIVo8Ay2z6Q7gb1K0dDA5BVqN00u2EUtJBJ/260vUBIESwAtS6acG/9Dc/dM
7SHSlcPr4SKHWbFycC1mciUPGHfoh8afSMrCCj95CSJd7hBvLouJSnoxNc8yPWhr
8zy0UrslS8hD6/FUKP+ajar21NW5CxMER+2FGgj3zvqm729VMNwB+xvKEEGab2z3
qNGlQbiOshMh9mfLCXY3uu2E3do6vj9jgyzymhtmonohPXHKbm/W1syn8w/VGbJ4
uGij/aYNuwyDG4747luPJl2/95MevbXMGmnwvmU4CnjjtkuEAG/WEdVrh7ICGu78
7T0SIxLOjk/7UWqTFAdUIH3g+w6O2a20gTnJeBlG5oSlL7DzxrY3FcooKaIQwwpK
EetG7QResGJRvX0T1cu8gRMXuWO2TEpwYQqSt2lb6LJcEp/DBytFLvRdYtJC5Z0f
9lVsZpYxRZ6IONsDYpNAOXkdf1FR1fvrdw1UmDZBrD0Z+GjnN6qPWFURT6Zim495
DzWw47XOpRqqiZBASIlSIbrO+7FQDzxBSBtrtkWnlktiz9N7sRdNX+/QOjqMJC1F
bumvXjVca5EQgRcZqoV2azhWPyIA8nJ7srezzXGAxYKfg+6KYNT1RzOqr/GXKMYC
CNUV0UzQwISErzkAePdwgC9Yj1Iyu8a2TCVo1j7cx0N3aDRHueky1OLKuUd8iUPS
vMGad3hyMaGIYB9ypohnwAN123X0SgHUvZDs1cxaLA9IblHiuanruRwwe4fq0BVg
Vqf6mD0NDqygAU6DuXGXql1lDJW+pNhFuEn9o1V2zs4seAwPI02DLgjDmYh5ADLj
rV5Tk3C5pk/W5FZKEH6ZTYfp5xdv3bHg3a5nqJrbEO63gzZMbeRMVdcbCFIkkJ7P
ca4dvCiDb32uuiaJThS4/dglcECAp6M5fP8BCNXwzhgWO5sV7hQz+pLVY80HBiov
+yU5t7sl1qbpv6h5itDZG+Nny1tjhC/9eQnTQaHsg+F/ir5vhAjlNqaN0IC++5mT
lfKN0PHOJvBvq3E6ls2C8cRCIZhqzuGRkCTC5t/d5FsI30dzuywsnwGaZKrOROcs
7PCecq768TL5aQ6V97/QnFWFrHQub3eoJI/K3rrV/KCOC0Nwp4yhT89vndINB8tB
uu61dG3W6GA/BSdH6oiKEv/gq+FaekFHLS2Rwgbbms19wkYCFSaW4TuAhKoah+es
5FEF9qLKHC3ElEWwZIthbCw7jYFHKUeW1UcjKR7kEPdBTkcjrfJs7txZrrISTkXY
alp1/NBlatvl/Z1NzTCOtdfLeTn97PSKkhj0c90XZmrZ7nbZvx0nF6LhEDny8cuZ
EfZjV9zBY3xWi9s6gP3LfUGbD7FshgdqEHkBAa20UqpEIT2wFSuPojnngMPPnvKi
sZVCq6IJEoU/vsPeDMqMbwhqrJsqqAq6ii121GZWBCaHS/dgp1GmzzIvFabEpsiL
UAY1eDrcHuwjTBO9vbgTPfmOQ+DzDIEpmLRzp8U1/9NiJy1kRiwKW2OAr8FDwev7
oEgzE3lKESXrNBQf2f/bB8yv3OFPeI8uziely5cJ0j/NSRrkjUwcISe7ckSVDCfp
o1tTDKXWiQTmJafpTDFOS7s6Bd+LMAp6/R9Q9AGd5gzUZN3t/ZoqYThiDqHo954E
JhZ4eo/U2ZrQ4XR8L9aDUVJTOxkvnC/VBFjXyaWlHGOFzxLf3WGwoMzYw9IqUXkS
kXID5umHpwAVc6oXgO8sdSAv31lK0VVxTMEZZHjNaF+9eSwmN5VS1OAwiLs0tyw6
Ia8AVhmDcHr4ZscY5x/+etUQW3oYUfPR+P+WyP7BGmqViTU49Wzvyw2obKAHQwSx
W+M0urrKzQ2WxxFgwEYE3trLBYSaSjTHIl0ba2bcya0KXe1Idp211VOwxabmuynz
KwKmEsfJztwC0dewTPFvMNnXaoZlHsyatlJidO0OngpjyhARdXOmw9ftd87kuCzB
9ZM6YIZ1kO/JH+FfC7OmBiL59AGY9fuwKGwGzYfw/rIlGmV/NNhrgqG03lBX2aoy
n7u90GS1KBuy3B7ZCkBrGBGELQoqklHgKSsk1chEU0BdrPS4WHL0h7bp+YJlKqyr
8O9H2uhjTX3DL6o+G+7VfmfDxyQ2cYWXRTkTB4vF9Q4f5eO80N+0L/5VpWvkOik6
Gaxd0yWBudBP8in8uzB95H/koLN9pRWlRM8mOv51QVptPeYCX5HMqbGMUzUENAz9
DGX0QFcS7NgXzelNYhtsrY69UgpWCMcTpcXB+uMPP0XbhA/5oI+1N5t4a8DDfm5z
/RI4I/bleT/thoZ087iysbqBm0ICRYl/yPZ/oMY2uzMzCsVuYKU7liAcGu7qSmNy
ldKauS2mx1GdkZrGBTpT+Dst1EFjksCPnjstC4yBaQxrfACfCkrUen2mBNj3JaMO
bN5IHnVTEhdO6Eq+hun1epzdm/wPkRfBQfIekkpxRG1yYHHU4VMZuC6GM38ClJV7
A26wCVFslZAek0D1kUNr33Ud3QKLYbemkDUyp9kw1UK2L7HCJOT4R+0AnC6vChi+
4iTCa5M8ib2zpU/C6vMIVGmhC73irBEZUMTo5KGVcYG/BeBB9ppD0PVJYU66bFNW
4IwEXKbHAGTBC3h0FSZtMt/6RWrGfZSPUFHNISxIsult/RgKJA7ntHhzxenNtNc6
Fvn6jPxI8iLlw9QFNLn6ybOUrwAYpOR1XIEvHvh2kyFPdtEwqErsMAfNy27Vpb3L
iONp/qr/KDX3vn4jp//0BZHedQhdun+gWoVtXtPHl6wTslgxmK7iFa9L2Wi1AVbc
vDEaSzlS/J5QoaEst6VSuBIe68xlZXzYXe58Ct2CFBeFtxGNcfNjzKE9W7uB1Sgc
YfAZLK7aq8w11tKZk5I+UGZcaguU37Ytjj6OVS29XOTjcC8QZWSZDg1YmNrOQpgM
KOCo8cCZwHcMUV08uY1nmSr6CQtAJ0Cglp2dHvgDtbTCjZst08UVRZLF/uauqiOr
IuxxBGKIqnxnMzJf7YMcfX/fkm9MyqpPzYu/q/AleyHDm64Eu7qYQSC08pzIdr91
kL6R7nuoWLhLj8Cu494WThbnT+dxX6x1V4m6E2bZh43UteZ/LjSGWs5zrZi66dEG
qs5JrlKnrK09EjMERL2Z3L8uDo/jf73O8z53PUptzEG1nxN9n43NyCXrPxaUirpv
srCsADrJIh4Lz5gQonnXa2tkhpoHcaLcdRvizx3xVmhh49QZ3KSnMhns3FfmetyU
yqQ4077YyqOwDLoO9ytOb6wIGrKbZ9id94R5AbxAh8etomhP64dRSowqNKJZEwpt
65B3RG5OTDHjaAslqr6TB2qJsgeBKFptudr9rzkg4wyg4Vb/taF/6sqG0hzPmFFy
IuyFU4guWJ5VQexF+tO0YPv/v9hdFWWRlKFbmpoLtDCMuURZ4r7aHxTBoTOErkX7
bNoM6BLTmkmz7kLrAPAx+g4aIG/iRLj9npYY1gb6q6GCNbbYUcNxcv/7azvB/ejv
F081kfGqiTaWZpiqWCZJ/VNaaPbHiMhQalp1+9ogCB0w8sUg69D9diGjb05Bz4Hr
RdWXopgzkVQfjP216jEJapBFUEzJ4KMeAv3VqIVJVVyAMkUIbdkbzeFcDHnJc+sG
meKo2IirYQEq3vpt2dXCTOKFrky2jnjLDjQ/54cv0CUcLvVoE9sac0eFNRuBZf0r
P4SybMU1xEyB4oaEy+VfA0XKyvnbnEq8/u+GFhyCdIqG4ug7MukUOQqPDqfEqVYH
pKEEhjENk6k3akq7lQCKNhiYyVtjqEsB2pmv7uAGRAMNXt28LDAeZ8HVdFLw5HCI
4Nq1chCJIxHiSUbBOKlf2xomYeFEyxaAoEeGcJSdVzUh4QurW5y2c8KL2UagILj5
YqpJyoI9ncEqKklz7/jDY6ZgN62TsRouazP+Jpxru6IOjiIw783cGieh0eGlBLFe
w563xmfo6xv331fyn5PK+RwMufVmlBVoL+K7u88Wpw6EswPyDDD2ZiHj4iTYyJmd
ZQOC+lJwwYh/hBGKZleUwPDqicFoCLQe9I06OSvjPd8nniznAZ6P1JwNOoafWoqz
dGO09wxzrPGVPs/dcmPo0beYjVBaoVz4O5r4bVTBIw1TGSI/My/HbyeIzieIu185
m60oFtaVqGGF+oP84Lmk+du5Pmk4CgPghpUFbeBJpNWtHoRuPJBDJb0N6PPMzaUQ
r4TNiLZKrEifuJox2ivGKF3kkvS3fKzl7i7m1fJPyrB45KrkPT23UxolVMg5kP/Z
DmcRnoctJJi0IHCAhCwcxL+IiZe0ivIKvgH+n2a08pUFhNBkAOXPN1a+0trnrOfI
4pnQxRiM+zYibh957Laz/gsVlBRA6Aqw68fJJbEmWEaM1EDFx/tJqSw3MSwV1DiG
oiroh3K8lK7StaGZsqRgLw8kqk8QR7ciwIeflsnUZoqdeiWJ3f6S5U1Se4VMOwPt
YfcTlxFcxBV4CtAx2F0flGeWXEWNqhxF2IeFjmYgVKyppoGIx2EqkwzI0M7xJk85
whWDdcb6MtVKAsPDdsYBYVu32s7QGsaGYSYpMTqezNMPYo05sBCyG6ypW6Z+2cZa
+INveF7GnrVLhzvu4pdqoQp5NrAwu8YxUxEDbh9OQrMIqOlExWxG8wWgpTRwSs4u
wKd0BtYkmUPeaOkpeR6mo/g0mVS1desVM3mFUocaKN04GQfCaI/dCW8iSdHIYpKu
m7QndjPNPvY5OiexdEm8ZK2ffz5dYpPy2cD0jRdeStpouwPV6slzxctMeJba2oA4
Fo7pahxc3YudXqovEXwANBgT/DF8KxI7m8PLxt9OmRjstwK51cDBzvcwDsT5d9r9
E1o/0E0WGuq5savYWrt/lIIJELmJ9SrOhQt8/zXyPlrZyZk1SW8f2WOQGa+5iaPH
ceQtxLWuk2FJ1EwykvGVCs11Lv8BBGsCehbU565r6b5H1o2rCrWLVzvQPT2uRv4B
i/70Nhjmx79VkqljNl6xFDuiR0Ap4hLXeWwYjOXR0X0883eu1vEkFQmIhq1frgEC
4g9HSH9jDc4hHojUDcSgEDwkstHGRqt9DMJTSH3ybL19ZzrO/i5Y3sZ7mSkO9wYx
wZLfs2YsZ2dZ4TcRyyoa9VXAXzeeFk6c9SEhw3jIVa3G41qvT/KHQlZY0rj4i78i
3roiKFAlvnLHrfPYTK2v8DTCpzIZuZFFDbSfe21xpktEfnW4iRjo577OkhmmZLqg
CZcsX+EexTFAb7/iEfa2kSeAHZHzjIRMT9qCMglivb9PA+6udpkNkoah7OCBuNYO
TGENaCDZJ0mukCHXxVld/rqnI/glZy8YkpAde4chL6Fjtq5X6eeZqqtlqGCxqKbB
IaBwsscu6r0q4rUBPo5AAxklcD5R0CLqM8dx34wyyanjKgLXPzKDoPszvP5eaEdy
DVf+ZYXerKG+qTklqELofZtj+yVw22YbWruFI07yDaXU2zqm/X1sqiu8qpyCQoD1
zyNYMAOEQ/B2nMaeC+6Zb9/UB4rgB03vLYPoaJtVWSq04qJXoEETp2F3c5AFvSem
Cry9/PQfUT+AIN1/BZYkw2gIJrBgXKnVj3hdVNPNbXWe/jF4vuobtfAICSi4UQ1V
bdOEu231Bxho1nwt6Qkxoj/j9zWR9XOt/DdTuFOBBvnFimWwZlfzmPXM9KZ58yLp
NmVHQtpIEqvIdEbdRQQN4PAjL+UEYgwqRYPYK7tUS15/4IpGWBU72rkLKycBFf2D
2zEF1QWVGWUF8d5dhsrVHee8vDCDBL9sQYGEyC9GtRX6DL99Gzbs09f2XFW09RPZ
ygM8dlOvwjwkg9TbKf/uUbDPC/qNWuyO91+3RtzJTSTMXvZ6mNdpC3va9v3F5dp+
dYoADt5BXsUsiz1X+5u4jpEDFezFvxTa0jecaHNrWmpL5vCWnBvPQBURGdGjT94M
Rb1Ygr0O2PJeLiouI+porYkTyCrL2ORSfpbcHGBry0egbQoK9bh/UJeaaJdbbdE+
5GVX3oT8rgoEAweGAe5pUxk6tAhZDTOJgWm8VE8MmYULKxViatSwY2/R5OfrIx66
ifLhz3nPpIqxk8WS1tflRHe4OK51AzSSUsU5nmuKltVjTKR4FF3FIc8Bbz2u6KcL
FMm8SEnCpEJ1Q/E5ynkR4JXYoSQmF2v+yfpR2vajKvXCINF8Px71983QU3H5rbCY
vytSy+wYZ4pTyRvKUmdsLbZjZiCXy9URYZOlQXh9n690CxXekFmaI6q0HbvUyNuR
Pw+PwRj/MD8CPcD+GvVneO5iBMWUidHqkJJMFs2rRGejYwl9A4RaFd7mBNHpCDW8
W10efhKaWRbrN6R7vOcWHngK/WkQYVv1RHvu10J49b0b4aUKXAFdjYAFkPaCeA3k
u24LbnINSvn3S5jBZ4ECbC1G68+VuP0o1XV+RRX6rSN7IQNlerDrC9J9EltWV1H5
PUINAoDxpsTOn0U+pjisbRclTULsaF7kwj9ctzxUqDvrm9L9zP4Eio3VGKRlpYE8
BZ46ExtOM4hPIHr60pFwcPy2y3YwqiYxYQ86PPvBrmUi2+SzsQu9DAcSQjPpniPJ
UhLGYwbPtw5c3ZE+Sc8YRBjZGvSsozw9VJKFfue92MJJFNyI2tY1Ex72nWSjOTxD
k2g/nzWD6kIBjG/3+lv/bAZZBDWm587p4RJFbE9/bkvHPGkXWRyp1na6Pb/qmOab
R8ITyhSWolcKm5zaUm2IBnTCMSJpygf6AyXfdr048g6MGtm/91JB8j2ZhUteJUtp
4hX/tvIbCJ/8HgS9ZOBHFGmWnY446SkCDHSMiEXx1PPix4aYy68J++vGArIxYnVL
qyj+vnay4j67nGM1qqMTcAXUWGoW6St0ifnCeRCB9/bjiHsjlUEMLWicbvKFoCih
X3mcdmzyusOeUDs2Dnr9Yjv+c9tJzk6VacJ0jHmepS/wU9AM4E/A7lqCq5Wd42Wl
N8TkU3Gq4MSSxZUK2drmcclp6wr5ZkAcBCbyk/TVEwqjG3ZkNnCnppWWNXywbBA0
zPQLir9PK6jD0OC7h9gJ5fucrbyq64M3A88GuPkAoi5d1xgoIjaBZBKA+ysZhztY
Yqpp0Qw/d3XVktN3ScTAvbjvhgNu3JoyTX9X+NWXNWo3G0XsYxpLTPdMnjKKBe6r
O0c3caJhNRaZEVPGH7Gn9/2Rz6GqJyHwi2OS7J5BFsG1sqiAhxrX9S+EFobgfZbI
mcD3W5lDxrj80lvToqrani9XKQiYggZNmdypAI4gNTUxpYoLNzBP9iFW+6b6vpyq
0Mh3tN8KY/RpimNVz4psbQvR6UlNWa2T0ahGoQoXi5fBShjo5JKnvgT4OjMNDt3T
bZUbPqtTA2ZvE0UKb5PygeulvI5An5+P0hAtm/EtgBv8FML2xRxK+UyrNafwV8fL
sQS6WSt673nGAWPyJby0RSU3qXdHgDsXt4uDSdlTjE3fraAllhXEjPjvEsRdNx9e
O829g7sM81fCpJk7uq/PIlXHktSiRkWOwgln0mu3CGFJ2yg0LmcKYJXMRRmwo51v
fGkG0J6y6033PhvSM2QByK0LbxwMUN7QLgmyqgXVlX3OJrwLAVsEcx1/H4wN1mzd
5LfhPcXyS8oUkfd8gmTNVohOd++jDTfvgGi+iwy9EcdjgLWY2I1IYkVZyo4Uckji
nutzKH53T9/BlliyM1aMWtD5PD/vRo/kxllyvqqmScJrTwLuxJnHLZ9j96xYceG2
Ts/AZjU+wMfRcbiHA3kNtB1JJMbytny7V1I2mciKPTFNz9PJC4NY7VaTIIu1ZPbC
y0Q5NNlGJrW5wifx8EGD1vvPcFu2elnTsLriHpS+lt1K+w2nrlSR5YUj4Rr3lBJq
hJvMlvV2VTedX5Imy57IMC8nUKq0VxvpEkrleduxvHD9sef4zvDi009hCsyOnyVG
y9fABaIKo+nQBnKl3rG1EZ2CSVdCn7gfxXePinkgEa6QR+aXl4D9YEe77ro2lKBv
miCOf/vMMxuFjvsA/++eyElGCe9PQNb93PRX41gUzE8x/wpNnjsZfcEs4kXYphRm
6QGoFZqtwSuvvqqM9UVrTsaAL5m+l3swAb6+nr7S3FdLGmEntL91E86AUDY7ELPn
LJjyYl0czy29gYgD/ieNt1paxhBojrjY/h3JkLMUobIR1eqMi7lNPP2Hb0wxTpMi
jiwC1tP+7q/IQLulhfWi+mXrBBozZpajGNKolKwe+1aCrPnQatCTm4yUUpzo2DKc
x7OS1rm5tFPBxTZW8vCkITO+Ebh2hoptACzddBeM3xxsA9fu23PgKdh+lKt9e7Wn
XA0zg+/XhY7k6enzXfin/aUZUJs4iGaJrV2dBXfPePq6g8meL6KJQrCAggvNrwxB
KdHBUEoyNnlH4V9qMUVQMHzoLJS57sJgc/TjeTMGSwVU3gANpzdZ4BZAnJTxU0Eu
j5P2CsFtkh3YNLsMQ+Wlx6z1VkDfW480ir11pyfQQcvU/VSFjqFw3scSwll1wn7U
7hDnOMpQXxLdSagSTlY9yGccRJsdN4nwG9p6QgCK5YXj/Q+7TAPYo/hKrvPi6aeh
AbeBrwH7uuX7wHAX6h5VUoA+R/t7t96NKSsags2rxfpsQz70a35ieNGIktXTD45/
hm6hhvGgS4X20N4inQFfsW/213pOyyYEJIiSnZIrEHqe9gcwE9vibgkjDkfs4Ffz
ngTeaCKdd5xAVatVUHhEQgUdQ2iGnAwTM47uDn3YwosfXXmsJODfsyED58lyKbZh
2cI+rs0t2Fn0dEbzQ6Xc9IAtFvEPJjk2i2PvbIMRnoGKbdo5DIIYflF1nw9bnCK7
BLs1s1DwVfgIVqQ/LhS+HyC8hNUc51lZFkUaNM0s5EKQOvg3uSiulm67U8xER4Ri
dC6mi7izFS03RROVT1HuzY7OJMnDZMXGmwJMx7miyvkchokGwKqnVJoQ/IOJDnev
Ydf1/B8NUUnyttSugFtQRRp2Wd0VGShWxUOiLbwtXC77uo5GOhNtIXk8XU5P+8Cc
1w+xHnOOA8y2yGp88eHXrmHn2gHI+HCicL/Y0CAA5TNgXQoRwsGhYrbasyFxG1th
ibQKsCiZqXqswCeWcZ+tTSq04XoJEasbQ7eXVhmt62e9cteykzQfGJxHdM1qMJNX
WDHdH035y3J63MkPgKsAoFavDvtrdyMhHOmhUliJfDnxSqOgJRrzuLv8YsUY8iHK
zQSUqvTINtarDSMgp9D0cy2IMiRnIJhfkNpvla9yWXGPtRHJQwMnVo1LU8oIQoOV
bfQ83zHBZrffyQn21L66QaY/9vSUrxImjAeLtCp8uqqyt1t0860Brpwy+U+Q0YsY
WSlVYGy+vJX/fUultAoKg/oOD2wI/ym7mqNT4SbRzhvr5NYvci/H1y2iIvhxxk1H
nXorHybv9D5DGQ/d/gsLK6yA6NNgG+TDUmZWbNDPk1FA3M+exhtNSgQL/14lP1f9
dCIX78fG1Jm4O9lDicNVine78EdiKzgj6HkSXDwsssD71hgX5tUA9FrdJ9mVu9Mr
gnzGTh4K5ZP2m/yS3/H85+yJNmONsrbK4X1d+Tz9K6KRPCfavLPi0//XcYVwPWi4
mGq9hJbDdMrxxYcnQ41m47JVcJ0ZKyRAx9yf0eA+OaixLNdwsFXRp/Mi+hXEYkuo
oZ581y05N4B33VPCOav9PKkhboivTJtJmaZlCilcHwaX0rl/snGWp9ypKAyKRb78
1HpUXElAoi7Zc7jSAr3Hu6CwwAUMGugIq2vncfhnHyKmYDyaBStyvJ9EC5Ujn/hQ
+FXkFgCOqCknNbx5EpRII7pivOlZS21Ip43/WAoZ4bS72/GisrNl7c4Ebihqxqaa
Joxe8IafWQ3S8yqm959mXYpTCi1YYg46gZ/trGrOErKiMhfua+qqFAtmE6WwQSf/
v/6am3Fe4xqWwqEzVHezpXZz6epR3BjqRBpjrbOelWGz9i+/QtXFH2ZrIuZc/ZDB
SIo1Rs0jfE/z8HK1N91vkfT3vwBz31hTN16FEr2r41Rv79j2daJAD/lYm0ZU2y3b
rN7gO5hNsJvYm6o7MIub9xiwbC0FCsXUznmD0D/PZPCpskhAvhQx3wMocDBYinYd
ggTkokB/iOISaFTaxJdXB356zCGCp3tDFHvJ+ky3OJKW2cGSMWSN2AEKe+oftmUR
iJ9ztoMZcGWjRnwdcZbbS22TYzFUoP9fMnYCUELVljoe6bvba9ISZtn9LGf67tzO
bR1DiO3DNlb4GtogkiyQsCmN4/iq91lmdr2LugoQodDz7lTj1wv/SK/CyWT6+hBi
jm9m3XlXkJc2NsbvCRKmJBpsQ3708MA/zME33uWeLd1twcafcA0F2mXCaeqAl7k2
eJ2FDR7q0SyTWD5qewLncYNS/AapfjZEGMesBL10b91/5eg365txy61Avy/ElLg1
fobSbtheLyrUkTKqozI8tXAw145wIskdoRY9Ez0o2Qn0DLqLY4m9HoW8mV1wqkrl
uCDpaSIe7hHJubSdGYNoT6Od4SWCE5yUDUTJCEpZ+0FAy+IE5CJyQw9oyN/c0+GT
zeWbVk7uPf2dMGO3ek0+dcuQjY8HzP5yVCQl4Ng4EZ9rDXoOQLpaQ2IQmgc91Kkt
DUPM2uhVF3hcOyiDez06QL7p3V8nx0dYosQAa1c+G8E91QWUCxp+ZsI1PZ7SA1n6
NN8T5cXGx5jocMSHsNziPxaOT+UO+6k+QcAd3rlWfWH6HZwLkNXwFeSZaTg8eRXP
1UdAVsYEV8BXBTFoOfOqOQGyAWPavaMau/Q3LYjk6FSa4p32yyGdum/3l41bXRA8
Z3i4QR3vIuJDEhFIelxBiQegspuxp8dsqhX1Z07/k92E3Pljw1aye8tJMOLv2kXY
dTS8DV6N4VXVJluV90PWVz9flpjPJXkskUjBvpu73SZhSvowuP0ggD80gTkiTVB9
VmCLSMfuXDsxg+IPnJ6oztvdTi8JsH8BZjy2kebko1SjJLejS4Y19Vq7zkWDsCvx
qeSx1/34ETYr5JyZtvNwHLhzNN5K3vR/IC/A8d80oIeXfNz/rdmIIAF9d+OPOcAO
z9ZQCASdEg5vbH2gaYOurAIiuy/M/kXON5FKX0IhpiefVo5L+wHdKpPdkNoX+I83
+9Mwv0I6U8X9xgfbcqLKgZ2WX+fjsc94+43Uxbz0mt9olohBEWujssfr/P3loT2V
OjmfkPFtASl08hNeYSa2LyINEtxJmu77435tFvhAb1ChYCQPXeK2ZMkZyqyhXXWZ
cop2qhjigg9z9e9Mm16iampNHI2WOvtrYkoaV0rYLlkiJJNe5mHfDf/cPq15/H3Y
RrIiF7dC8bDm2fltQ00D9sbQ06fHFQHH6mJudnPKJrp/hAmqvav+NjxCzu+N1fWb
yKCTfX7q1FAKPhfPzgrhGSpzn5lNbj54o7vsvhitpgepdVgXaW6gvqo+7kPlqTrd
RtS4JHda0lMW4J2COJUnbEBHDWrnoCHrbwA/bAgmVnDS3nMzGSHSIgahvbYI7AQi
jKjIxdaqRi0H2X8lxsIHxN2HR0KlYoEZLb8/egLxolg9wLLUbHcCRvg/lyS5h8Uo
h4JztWOPLLR1SfPQsN5JDiCunT70N7hPyPlIuRil/7gWhEurNj8u+F/hr6E8xqC2
SEVn53se6o0bv8sGwvufiJ5BlXx6tOPF/+T2CZhZXuT7KfdqFngirJaBPE2QHrTN
tccWGtnxWGfByRX7Q48Et5A+0Z1MqMU82YSFlpXDm7fn5zAnhPOCGgKxCna+kDUq
QTnpYsv/61tvdUq7rVa6oFNVSDWLbFy/icJAyE/0HR42CAJmuwvHF0O7Z4T15JNU
JaoBkLa57pLxNrVYFDlGXv2LfVAI8Isvl8VSLtW5EzvbSpNUjbbXS/0gENkOUJl2
BgTud7n+xpxv9JZKfjaqww2Ls7LdYZMjZg4pX40ZJ4ZqGeEEpzjP6uWQSAW+wpLn
wTl8I7ASe2HCCKd61531SV6Mo+xBhij9hGkj7J6YgkrIKdhrxGw/z4JHpMbA+UCL
zzGIFDVpfLN3bQe7kJQ0W1H8UakF3M2qUYwlGh7kQ3flGe+BBMPTEdd+LGcIePEx
PobPZ/FfCxdNH75qhc2SDdAuCzPsPujnJnLPgq9HQINI/yu+x5AZKc4qrxevcHrO
YxysAsrMTXXxz28PAKSrmc5VMB5vzlRRza16Wr2AbC33nco6/YDXuy21kk5l40Wg
g+snf6RMa/TME9dz/ZI7QUrv28ZjbK5K0PXx07iySTWbJKXqW+GQvEGXOTVjGZ7p
gVvIZUB8RoCE3nasmNMKlhwF471e8RnLgYjPoxtv2LLlfUywnXxnJqSSdztHo8he
hSzgG5rgX2onL9gxk5SnlAAChZj8XrShV/qLBHRkw4yoN8haLou929yJKcGXXfUq
/xZcpgRQhE1K8D3RqKaFsEYjHJQrtYHKtPgDg+h/KUcQVHMO4ljUBXNtoHSs+/ba
hgbk8OpLnvjxBZso84TULWadPODBarFlH/sNarI5n70/bitb6mdQUNSb7hRZbzzM
oQMCDKFfMfJmBZoMpJx/DbPgmXgJS3F23tfXMEEJwRRRFx8SMGU+1VnVjpM8hSTa
pvLmMGdBde/rkmqgymbmGugYoFemW0/szYwsHn1CjlmYCutXes+ZVWGW4pcypjQt
DwgIUcu1LzYcrGH9+ymjDOh+BC+cQoUB9yDAkcE3a/tA9LLSV7IwLZAozJV1tyDv
AN5MjTL/yVUGABqfcjWQeN1xPsO2UOUenckK3whW79FOHP5SXMHc0sM7Fjsm3nNO
awhMiFIUiMI9PkoFSHeaj81MBw41rkOTbhGdGkko1eIgx6eGYtuEl7ThrhxixzCG
YgUodddXNkPwGl+EOLzJrqjY13X9Zra7x+qRH9g01t8BU+bcUctlGEqsWBd5qsun
tTGQBpjiwEy56KCC1UHC2+aNBGlumGBCgE36Hf6rRqg0TesD82u74xNRrUhcOZFJ
Xu+sfDPBjtU/lN9jnLgoCdPGNQV3Xg9d7fOKnZR8K/eHQZ3l4VdTu1qIZvIiivPN
x8af+47clFZApINZoJJFhDCooSooA7aogOM2bMgLdVz31MQ0PoSQ3Plrf2bdiowK
nkwv1SxzDUxTqvUeZnpeo1guI9qw3HpgW6iQ3EildEaAKD67wq0FGLyYGsPCVpXm
3u8fT6bMRgIOdGJ/C2kN4c9iugu47hN46TP1chStZ/FDecRg4s9U19yehTbp67/C
wveWhbjMVnK689F9ixQNcHiUl0yJRbaKKeldPYbV/AhLRwSfmVF1vliBST4dk7Qh
pRfxzRZZE5rkTKWa6CaGEZQ32++J6mOTdgwZAoODQoJUUnW/z/poFpNtAuBgC0zr
ruNflHK97ZoUCnByrVZJuAA8WoBPMntRrB/s5Fiqe4gbwDXmwqd2nfr6BErP5+hC
jI4my1YB/+cUvYbQ/d5blYrHIy1bB/UCUT13W4cD/MvVz3LDKpAS1B9CL/hmt8Y9
OH/Xl6XCCggvpv8N0CjQ4mCh+b/ChSR12rlWPcDc2cejai82gJFAwYIfo4J1GJly
w22MZ3ECWCNaB0Qc/atU/3i/oL8hTJggLVXGkrEFIhGphm97ehXda+A1DS8FNoeM
nhtfsxtmZ/1EWV1N3QTWdIZZUBLRy4SB8uNDexWSvOECRBXmMUWFIzqV3Q6FYVzN
mavTfgW7KPtOgJHaC+4wz9UYdC3OwS2pMTRJjVx8lVoUc6X0IWUBHymIPjzaRCBQ
pj6cZUbZiUyPuBv6J13Py5TBp/sArrX+P3WI7QMKpt8saC42mU9tfds2T8iWwmmD
BI8n420feTvO1sjCeIHxyA9TX9t+Ae8Vo/+sYJ75osAIn6CFVrYgs321foBKneY/
RAimbX0z9q/ir8CNy7Rt4a3E4UIYcWgDejAbOaqDHNSPa75EqPYWiEOiOI5XM6YK
/JQAx2F8qLXe2TBepAUa0hE29SjbjmP9Jt6HPWSP3ICJ7ujqjWYCeFCdWd7Z1g8B
nMuvVm/+sYTo9fk4WzOekKmo5bD4jjfgAQd7INyx+RdPyR5vMQhciFirzI3xQqdV
XdgWIXOH3WAeZTSPzLY7BIMSbRi8ZAeDLPxp9acpob/oSt59f1K1Hj3JokKxK1Ug
tBNpt6BrJWmyCHRyS971vzKNBBmHI/a99DxrCG5lCn/uam1BQ8IPIcGh7PE2cf2y
2H96qjv0FqekJ7IdIXpQ99cOg65YJWtBUgR9NWccrAT3wVNjmI0ssRWl3WLzbY8S
eFE+7MWBWDeMcL9CEZch+nmI2YmYOfuqTdTP5YqGSFQmgVpFstQoeNOUExoZnPz0
iRKV8gbCiesqf8b4UAa3/OdJAyqgC//BrXTnyraC/GHixSbfV6X3iD7icXt3jTu/
rJsIhh5RtxdDiw2VayjfhNUavbBJqjfGce5gBlJVGqDcDSRrIyUUCLfifegsWsya
F4eB65zXdsAwQsZvvf9J72aUom/fupetL0eVNdpHX+3Bg2sFDaVb8O75DgbgvF2w
6SuEGFzhNB3dclUYT76OMajNfI+ietD8BHVCl2krCIR8TIt2CLysPJS2EFsYaXtZ
OsVPEZ2Rq3TbrAfbJfoLBpzMIKyiG2UX6ShHlAWbm54ZP0USpL0Ad668vufQV1dM
QQzVTG7deIPh6Yqu/mnpAgZeJU43qcWrNFaqJ1K26mpTOfmMQ54W44VBvDbmSnfB
l3oG8jK4domIEj9w8471yRo9aN5WL9LRrHiFMTDyQ9yEW1uuqui+knUyKe/nMbwy
FOqq1h9BAsgfNVGfAYuil/juwonoRVgi2gBv2/nmju0UOuFjmb39001ioZOXJ58F
Ak8Xw50osiZOiJjCgiBO1I132AUPipo3+MvoTdZqRBJ78Z1tPma8YILoGEl4TNL/
8NVQptPDGhIXE+gZDN4bm2dbrt6B55NBsBBxwriNyFeK4cTwF6xlAJHCOceCOwhs
DrlskzubIMQVONSA22QBgqiLznvCnSzFTAJDZuo/N6T5DOSTh6FFnYOzfYG/XD5F
x4ET20/H0yPELEMLkk0k6z5/miqTZvDXthMbbfLcJyxSyl/Bn1FrHBjr8n88WlsX
cn3V+YgOKuKG7bUzuLW5wuCUdpIKnLNQl4lnrkKyrz9Fw/u3O48IwcxqiHqDDe2h
g3flBl83TWL3uKPY1Ins5ZrCCUTg1v3dR+7chmlKNXTHU/xB5RphX/u37+59GO8g
CBilM/3vStNEGaoYi1alNhKCAc/LD5m3sv7bSjl8Lo7W0NlLA0jKo5dnFOb5JUsK
hvSUY8iAa4Gj7dLOWicZsbqO9a7BFLEsP7fMOjs7eZIcWvPRQEfbVDAMfOvOlYx1
ZtlGGxhnx76RBKkpetG20XH3/9s73QRv/vvnHgiBHX7W/SpX23u5pWOv76t7MJ+o
xc6BgNb5IWJmkJ/Oxh8OBpXj6N/dKqzmoC77ayB7wm4T0EFBY/bwq/I/Tv1kWZ5G
f4lC5UjGjJ0utr4gbVp+K16usZOt3bK3tMLQqkGbtaVZ8BP4Eaa/AIwbBE2D0hEm
odfes+JkT6euxfoRRAfmPUcw9NihZwcVtLZlDDGYZvS0J4aj8Z5fNprCWFzqoqhz
HOGm+Se4b2Q/K4NH98nMK9IKfeXSDEbvb+R7WXlRN4dGkEuk2ZCaK1O/uUnAPRcd
iXFzkdHBZTr7ZzMHxNhwIpO+TKdYLQvgeSNDcvF/rTjbEYgaQBUbqWOJgJzvaMhJ
q2lmLBoE+8YXtTgi5qASL2Cl4H5kjTTktr8uZZqbGjUrOgujJw+aarHpyutcXOr8
NaLsU4CaCNJAy+u3jR3gFoctGhBGkNPFOzwq0hjlt/LDk6Y+rZyhRHwDM8F3p84F
b6ceevlkYUyE3MLi5GC3YvhLvDxWyrnET1c+9KcoXrin/HDN9DeJ80qeIMOGm70i
5PRXKWg6Ul2HwtSy/K55zYaxeAa/RFI3+mJiO4A1V2MNRgmmgFgVty2tGPYHOuca
Lc+Om84IaCuYmCM9a8pZh/057fwVQePlavmgPx8tDd25Rfgj5vDnnFsK06Zqg4rX
e1TKrnQxa0CJZevbGnExv88XVZUwLubT88210yDPBDdU3rAQbvfja1UC3FbgENyW
i+ckknq9GNeueJ/rWRQMCaALUZeBpLKNfGQlWEFAwpGbxiZd8ShmQMw4afyqeLms
6myjooPFAfduz2UN8DBw/xZeq5Lfje4iZMmeH+q39J5ezaZlsgT7RcGiWJyuEjjq
NJqZae68hlJsA7Yiq7lXPfBj05o7ssjcFJ8CbcxaOrpKSyVblAgjv2oOW7Sr3Ysa
MidtOYyL0MNV9FA+++xqbcQ/X72TsxJQM1+ov6FtIwa75tNvfE3kbhl2JeJEj8zT
eKe30Y3X9kMABiQop/FF9JHAztfsamk7vv7vHT9B8hTice74jzFlVF/3hyFOC+76
AYVEUak26eS7SMUF5UCyz/Zjt1/2Ndv1p+0qS5wES/sG6GZYBoYQpNJYC55hPmF5
6Mm9fiITXyTwLC5Mu9h8fOF/zmVfz2Pz9zQzRqpFlzZYO5ciPP0IcfcjA1HQUf+W
E5B0Tace4GlDwpuO++vn1nPOwp9p7lWzt0qXjEKA1LRaSoGCrt0XYsQFYU18ISz3
alRSuJrDvRNnfIckTt3U9tMl9OBxPmXXU3VUtMgZcEJygH/hP414lQqweJknkDEv
Zt1nw0tuy1Ksko/btiYtK4Gp7ycPdeuayrOWZ/Kw9x6R4jAraKEBIXDimGqWzVuC
3VpDtS76eGmywczJ1zKST912hVHg+DgR71VjYOwj+BafQEoLp10cjINaTRKdwtfF
QeClpa9WzUCfqkI5Z4C2uxzGDOAmIgc7e2PqUW5Fu9VxWuXHjgbS+xxQg0GMMYtr
iq1FI/BIWZmDwIGTEGoggdd5ijVYCYI+7/edSO6f65mgbD+PV1ZfUs/V9YmsxVDV
kYZrtrgZloLGl7nrcca1qv+iJFekuibSoiDJiKn9nmkbIo9i5VEwhF6T4JAoCJTK
/HH34/xAZWcCToI1k8BGcdaUdOuUwzMGaEdzAvxMiO2TOYnB8a/kgG8yPiLTlCBc
p1pnjwv30qt+Jgfo0kNi//HlpJPg9uG3eANVxKcrpl28aP38pT9g6Ezisxw4ThQo
N6eB6LpTMk1P6SlKSqsjUU/3NnVAZOXOKl1ihilZlXvyaociK5cQ3y2GkqhPhhXG
BJumZqa1l3TJzLZ1VcrnqC6868z4zW8WhA0Hw6dL5ywPFitArYDGu47rcOybt19r
uEjwdP6ZVgRFOqYfWPN95zHg8jxUq1M3QMEKb6uWYGLWlyAVUCv/MDVf7Zc0k1mh
dt3NNxs2k5nTS6tGYehcIc2uEndApvcRlE6LwzLyQ7tyt0yV3kaq6ikr7ApqQ0+h
QMqiY5toAbjyoWILQstIQxEyxButwkkoXcePLa4gvVnFh5l48NJu0enbqd1hQGt5
qlDmyF6QxcTQ5XRV4cCF3tQ2FiRFHSO7P9qOrtGv9FTokDt/kpaFctXD0yzBcddt
Zi3Kw8jKUo01fsXaSl9TSF702i7QVgz1aEeWWHLYOIalqKu27+QbxzLCqKkmAhPp
y83Dr3qcm1xzdMFiVWEyDxLmUqCY0b449UnYDsAPRie16kClk2NI3n6ygwzBJ2w1
TQ+bi9m3k900fT5jgawsK3EzLXtUbThmz+lkmZWnnse5qi98wFgWrY0UIcveRR4O
cqHyGRFII0UIUpW3r82wwDGzvXFVqUEKIEIA4bepVJkl1EEy3bqq5NdEm8FsTyzf
0JVoLoEEzevmfJ0LF86K4wKsSSpuWstJ12te6XaHXmbNU5HOX6icGqe6K+QMjsQp
j6JwZf5sNlIuTKBzeqFubacvXy+we1Eo5Ra9ToO/QCk04Q8PvkqRQY/qHEcpGqW1
BqjiChvd6BMOc2FE2lZw+H7dbSdAgcqAmB+J3CPv2tEmU5PSoe5YB3ja3y4UukN8
6aIh7IU7tvdZaHxjStR9UQJo7jNb+6eVHuDUo+ikgDwoflkgdHl8hHPm3973RRHy
MlTwy5AdAjscpmr3/LERKsOE+FjwiyV9GVD3oi/QmOf9kgcsX98ufovojNlYgsZf
IkCp1fflG95BbXIHoGbMnmsWwOjeoR6GK2z+zymx8fvn//Z/QdlpZ0R9hhHA4sJx
0LS2HvsozEjoJ/s901J9rzK8Z1oU9gu7a/Vk25Trv2+1sMVJr6YMgc6YqaCf5LuG
Udgts8M/qT0K7HEWn2chSEcWoBPpSKbdlpy5qh1B/JJynlnIddIENBl7vVvWCAmu
S3TCtNtNDuvyymmorZ2nScz+Kiqnx5o+reRwOnplNFTdvan8jxlGhEMaKJJrIS9a
t9YX8RpaGQvMOyDejKKoeWIhVjowy3i42PtkW8OxEtJrzTOOmAWqAkBCkVQgSymc
T1T/5P0CuC9K9QBpqeLCPTZgEAA+T8PeO9j2Rup3dfUTKpvy8uecOR//9mm5lqYF
41ukN0JxKd20s4q/43WWCHybQra3uuOcaP53BJaHMn/JBWRbMhEbbMiNifMTO5eP
4TK+wuehcSgH/MM0DyBxIUpO+iQViybwjwnkaxATcGGMH0KVjCDxjKj74DShEwoi
MyYs26XCrE34K6cWU+7orHgk/69XNp9FOrxRcsbaYtw4Fw970HPQqsQk2JepteaF
SZZHxkYoNrrrRyl+CWdkrAqpAWtx5kUcQQLhEH5/uk8mJqhneHiJYnOMHr7aWeOZ
4q+nggC+JukrnP3mvhVfEMZRGVG5S5iYI13ceeuXvp8YTtGFWCAvjix2fL/VGXdu
wAA6+XX7n6A9oQ6bQ0q49w2tLx6bFr8uFoejKz/YzOVsKRm1uXVTSk5YLfDwcmMr
2L4oVidaRIgpFqx23bxZ6z77FW67DRgQ8q8TZXte9M9JSsefL0J99luqd9cBBINw
p/w2C/hjmeeyt+WmKSUU6n1QbzpxWCz8vLsfqvQeUU6sUmUqkZ1siLulsjXnnSxQ
huBvai3J1Qkw5NzquGYsIYhh7IbmJycEyvvsHVErS7jQMQ64Y1bJWPShIBoI7fkd
2vaZ2oASbzFmEeh2xMxqMViobkv8/WquhMryK9PrrQsf1n33KeizD6jViNT5QzdT
JM5P4Onhq3P1BXa/BxTH3X4lSZFpPGjQtUYdp/4TRkN57uusu2vwl52TAPLRuZp8
dxDNWWS61UeBih7Mv5xX82ehsm4h17ccyKgN4lMKnJNxo5MHW92RM1Is/3LCDpM/
/u0o4HW4T0MWqZDjMGnDuoSmGszeGjvLJJH/Q0vHIfy2uWYSidx2EWqa6gHq7Piw
bVbsThw7Smgm6SnL8deoWCzgxzPtdnfFDI7pEMz0FcDf2kO5gh6obRWmmR23mEBg
2y0h5D/9tJrLEp4whUSDdK6DchGwuFSh2fpHcUUkYBunS8JBwrnF5DgJ3Q9a984I
qI+m+9Uyn4OuoODrrujpGgQ2ELMXOjUThEVHpq6kRQGItje5LJdZeeMvlvh0CNJb
5I/TsgqpasUJXf5EYkezOVvzfZRWKEMbG+L+amcSwJ01hRwUEJxpdEs7avvfT5bc
7ByPzdLvCvQo5uhjMpzmoDQr4FxLDZZZO2cHW89+d7MAftOjQbuuxeOEZuk3BFZ5
lFFFBfpJq0pS6lmRuuehDDl9z7g2UBi5sOivrMoQ5ba9Wj6fkr85/ngoFzGlK0ge
tvqW9OpTaSdCORPbK4+KmCg295J9iybOfpdpQ5k/ECPabIqWqhQ6jpUgOkHzUvSQ
cHB7jueb+Wtl3W1xlBeBqcQs7gXdAb/cukKbV2IEINAtw1sRRKTxXBbyVZU7zyAN
qwKjjHCtzbzZ1wZScKbdIur9uGFs6IlBKdMgJdVuxwDVqVfRbWW0I/lH51M29yJH
/euovHrGeReA8bwbR5GOlzHRFK+jCU8ped2PQtpqKDiTLBHYFYMMdjKy/bXvHJf8
ZQyrBueL/YZB4K0j2XIW7M7VOIbddP4l4l0PsOC/i0uRVoWcJFiqJj8TIK7y4TnX
CPWibpsKWdzAh7MP4GYJeVaMN92YWmED/9mByV3KaLRqnQycDke10EbHWLszNapB
chMDQI/R2cpkQZRF13Af7kO7507ZGBNrXRlHYYnw5buVNlxFDXgmx3YDBllo1mSP
IULhPu5qliKaF4nvLtWiEYNoX9sto3tMyD1F7zfHCl2F9WZ/jkn+QhmAh05+hFGL
t63u2cARBNV2/CfevZF3a47P/7gDpLoySDKGYwL3MSrBiVEds/Im6JSEkKCRx0Rn
9aBMwwJzKaUTXIQ+3v559FFIeYwCV6iQWaTr0ONsChiK9dl0xiNll652smpN+MfC
OeVJkeYstrhsUKUpa4ZFkVknSCti85m25aUdFGIup32Qh1J9lDsulKAyuOi6DZC0
AcBXb+X9nOpJooB81zd6yyX1AUVRzDt6R2o/OCAz8O+DRM3MAke4q+b5DJ9l+fFD
oUOljBerE6/6s+yO/XP7GpWZWZj9sbpnOdzCJ1ykLrEWudAwNXCoxgvJHJEGwCJM
YwHR9QOrrwy5vcbogIOgHYkxNJeHklWflKWwJCoaGuRgLMCtumHK0DfrI6sESBKJ
seJdiEvLev6ORaMO+gT6gXPATG3p8UN5q7S+xdZIhtisk1gcp8o0PYvCv8mp3Ov9
T2BkfIHRLy4wqBmPS8MvdrUThu/t7hmXYwODijVJpNxhIg9x2pLGKMYvQAnMh667
WQIWuBTG6O52vAzayU+IjsGEAbeehj0hdd6S/YOnfSVbxcfKAwM3Yp4+iUkAwySE
lyctrpyAY6RK1tj3UY14fUzNQGJYTXYfC72+XVjggf8IyyvMuDLm6EId0XG9xM8o
gEVfmchSFL3DfEwckuLncBVwEpG3EeeqS66erPeYS4X2Qz/iF1lwn7GOtCJSNdY+
WMpRc78/X0KLITA7UKd1S+ogdN2e/Myl7iI27nqPQoffdX7y8W07a8SVmKRH/ohO
CFjLAgXW6s+o2T271oTLL51l136hGQFhBSwNUDYvT3M+nwkR0Rr53jD0Fv62KH5T
+sonTovrfdhhuVY572FTZc85h61b+bRa6O+qDts0AmAk3QkeahblmlqmLySNcWhW
Vi03lFA8wFj2/JD6tUSl17rNllvKiR3F/o1z7vveW4qnSd7Aw+SYRnUlQjMC/0Xr
PYIek3fq/Kje1ZDaCs04wsBoUyi0O43nTVCQYpl1JpKskQr0/tYaceKM58Erc7BY
wKbT4RfQHWrLslY+lBBq0lJcw2tiQSTa43BHe+AWHzjucMBd4LN5y14KipSqph7j
bCr5sUqwV61eq98CK5Exh55ukEejZWlHWK20QbkkLd5hfDpDqT2X/ikWKXxJy81y
shc4cNG/ppnW/Lpu5C4Dmfwtt6OsU8xxtpKm9mAjIxm6zCvI/ip5TiHMWVhJKqxg
6R30HofGHpzZ7yYGSXDSgcaaPIa3IrHuidqNWHebg8rDfh7WAPd7Rr5DTZMfD+aK
ao4r5s+wef8TboqNfvciEs+jLZR6bxooAlF+SUXwfVX/y/86uhgZlm8j6hemaRMC
N4AjT+2hl3kBT+SA2MnxLvtOVkQ3rBN8LEbGZ/y4bDTxy0rzHkEcJcE51u7oPBfN
Tlg/qf8X+y3O+ClsQ2EVsYFVyS8f9DUxRg+CHLwH2094O4UntMMaV2mOmeG3wAbA
ML1StB3WXgEHy2KMeyJoyMbN3XTOi4fkVpxjEyNToxhqkJ3sxDfQ7avtw57Xkdoz
ezMk13epuQIFLi7+dPmCdmSSMUSx+qhwmf6qZwvVspR605vsVfiypAIt8B1Tjj81
U/9ZQ14oMOEpXM4tnIxkUc2UVmDJErn0VxFo+KCzWTL/q1xS2tHCTt98OtqZkjr5
9JhrJxSsj4cjdcBiAlweTxivc7+MOQ8nQUmPyZeQau8upV9yT5BvPjDLKiaJZqRy
jfUAcQXDVz5K8MCn76PoOiS+gVsTMlrPeyoJM8ncAb3QOH93xNJsP2am7ifjzex1
1dfNLXmxKtRd+l5yL1weIlR4cCx1S3XLYibLJLeGB71kQ09cMvho4hGTjKRWaxJL
+NVGYOtLoqfttB0/A+pD/h4E2AghqTgXcElNe1/HgVR0cw3rD24pMaqPkrr3lmoH
ak1MPp4NPBDzA9mmQ7uL6WKENAIdFflHW0VaFIYLWmW0kNADEqA1nslsaE2qBYU+
RAcRrbTc5M1YAOl/6N/5jznS3qHbrgfHAG+wIYFbBnVqSSV30tR67JqTQYwp2nTa
1xuxiKlw+RbzTFVOvL8oy8FyaLC1Tq1IAw1yRYwtgFGNXMzw5mVSh9gnqourhC66
dN0/Z9XtB/IGhBg9BQDaFgn0S8tRQni3hPfk6E5oxumLlEOh0LWTIUmS4/UphK4O
464RbQEHweCDMjqrZ6jmM9e1QcAdA3DhBYjiImGlma158AEXZqD4lfaG5F+WvCi+
J99ade7Oi6jfV+7gaP/4RzkiH5wHiTr2NXkzaWnrszcUPwfjqFyDld8CUsATh2Ow
e5HtOY4z586MazwByurQrrQZF4VvOI6GRltjpSQVJ5fJYVYUBSRx0CysrXINvo5w
CoIMdm6QQGQB//gE1iup+uE/7cZyCA3d6b7GGYxDcoNcAhgNtxHoytZKaey4hsLY
L6QyrNPIgG7slLUjyIkEJgo3fqGxpJ8qVdIlGxrcF2+wpxdzu1cXBCq6blFpTJ/K
VdLniQfj5Pbf4c4poTqk93yT1cd4643sIu8waNeibYZ67M9wHrVmIzt+p/Z81JkF
ofjRU3YDyMnfdFa5Up/iM6G1D+eisicDqcqLAJAHzz0LJitgF2lU6ERGmOVnbg55
ZnOdledEuaj0PhNHc7f1H2f3sVL/PiKRCPwLdkEEsjmMpaKBgCTOkkFBkCsYwVBh
QXn2SIQNmOUfwhxu/kVYrWUtSSyCVgkhsJMY8hzyTwC2nq/9cxXVBf3x8X6IMNb5
r/CRuScpROgVXOINwlUPMu5oP3SlOyBevnfECTo1gVuyAPiDq1fchN+8AyhzWB8W
fHdEzaFq3YWJG4UYfOYtSkNmlCn08xFfTfOBvLSoskC1nRg9yBVwAr3/NVhNyRbx
oIQVZP0NcfcWRbXb+XEHb+3cQq5DMO1hQFx1gK1zOqpE6igEP4KBBV+StMYw5VkU
k6hKJWpK5ouUtWGQx2BtmnvLurp3DLI7e975fD9Gtpwp7JtY0gzMueB4FgPaQyos
8Fm1SOXGnFdrjjYk5fGGLoncMb0jGWq0x5ESWbaCrzd0uBfoTjvO9jO590TGwNlP
e2tzy5cbw3ELKESGUd289jENLIU0uSm0WGWIEVx0Y5emiYVFy1kGZexLM1KAFdvM
WbFjRLcdqoiu9734/hSZgntYefUbETo9/dzp3oGNkGc+GxOHWOMWxTS7AEX/n3pA
lTAiKTWR9p+dpF3crl5LiLt8ng0uFjeR9sNwfbwRME/qUa3KPY+LDNYemfvr6UTT
JyX1XDrtq2NsWS08raThavV41ZV56VPS1f70SZ6y/G7aNu1IH+UP/EY7GInyh5GO
C7nW02DXdiEXqKMRANCiYHOS8sHlPYykJNW/blLux2pGe00XxdGW5GIeWS2Ow4F2
hxBZB5Euuv5B2/LXNYQviex9f2oWRc06qYVQhuu0YvImY2F0Y2yuPSGCTh19sJ/a
33RwLMauo/7e5Hf6YE6sUGBTcDiJXcSTadwRqrC7RFCTy8WfiP8dg5uagjUByeEv
ZgFvBwB+je5wtUDiFhfgrj2V85wyP5ZjYLXeBwe9rBz8TF7cjmAV2sV0gc8hibFz
vhRvldadGm+PZwStM/lg2dgc4uKY7lz28oEBYzkivdGNoMa0xlzFoyZTalYMUPRK
Vc75rkzau5v2O2cusvDUgFboo1zFEbThFcIvg5q8D8s3t1nnR234vyth1yRsmPLG
5+mHFA0/l8ivSG3sJRjPkQXQ45cHriuawQWJ476U/yra45wUhxGfw8k6Kt136LU8
0IalUtsx+XRHhSyEdSaPbZlwbsESyJBUp7Vy6V7luwbPUtG4sGxdrXCA9b6APW/p
zbaRd7ONDlslPvDrF2TXGcd2Uivw+tDm/5yOtHBMfoVq5UumZ45ZS0w/Er7RaEXT
WYkJ1jA/XrwkYiHWYfjjyqi6TLdW5RLrfu1FgSb8WbFVqn2EDFO5XbFOSWVGErjH
GIHSHOJJmfodLR/GmV+QsCXumizT+hZf6F2kz/ZkWGofyd3YLxSi8ufac8gIuAhj
a7Lh5yz5ObswmXfo5rXsAEe8qi1c+hUUftkMCgA6iKgI3bd2+GDK25c/bA840MLp
1QfC2Hoo6AQ1s9faMtcQzT2dwH+oC+MTSQO/3k99FNzQlMSwoGXHDULh6afVDhAQ
jN2SR8MgO/Sim6Ta+BXgUEpLzSSlQglzc5YEH6Ijxo0zKoTuIoqt6Gmi75NL7TAd
pH6eKoWKh9b0IOuOAl0mNuqYOPuv6V4o/B4Oc1x512+OQ2vU3LtPza5xD/VQcBOc
FRu1Nw5Hm5BisHcY4axz5ITyyBkxlCeq4vEbufOlzcfpRbqLjpqW3xLtBbjmhhnN
W49HI7NeF2JsSpW9Nu4UgjmJ9u8DF1H5RzhkBvA++crIsjG5XxyyK+Q5akNkYRjC
XG4A3kb8zo5oM6lYVrz+Agwf2VUlLdQf99Nj1znIBFTvxRm4ZCmhDm3qqX9U8xvq
qlfynztd3pthhjfkj7Cd2pvLqkCs/qu7j/rE+3PWH31b3iiZs/QW0RH0SXdV4Pyy
PeZanC74pRhUmiM1U5HA1v/G7rGV8oOoBEVc/sjs+GiaiVL086seJ1ruanPUwEcK
3aWbHUmr0Ilg0YbMnzR1dbiZPq3UImLE2hx19LR4e9aQEqw2GS4XVLfZZp0SjozT
fNYjjEC1TxW8ymF2uvI92JhIUlEfpBRWbBhr5Ibn/DD/umjVqkH+EPenKCtJY+8N
sLAcbDl/B0OHiuYPMJ39y6Hpd+wvNFPK8ExfUSBOTIDQc8aGQeFUulqbbnhKbXPS
Dp+J9QROA20GtBPNVt89RmTwVBCI9ihLC6dk6pDLZMkS90fvGb3z2+Xv6XZCKdXr
xJjdhE6egETeVn8qcRp7xb8JLg+VC0x8juY8PT3QnChpMmXbFTNg3SbPjVnYxYdX
p/708tKY0jXbPqbXaWbHThtQ0V7BLmR3P4QuLFE1pfHKWlix7YjDmkIcFqhlss9h
H2ervew7CXdfAHy2mpg9YXu7usuWGCcV7Al6lqB7gK6eH0riMrH38RWxlaRjYGa5
3xijGM8HfJ//4Mr9XbWt5J8jtmqwgx+jqF0BGNnZzMP0GrdPkcP/fbPApDH4N8+l
BPqn+WWmEeamQRSQHj2W32VHVbgbLmnuyXQ2rGiUXzlFPCjbGccp9VXqKbpysbFo
CR5fZbvnvvRfo5HF1qnoh6c8RRYDUrb7jzcVZypMvZLbJj6kHmf+dH6QQjQWu6Qk
7LCrnIWzNZZkgkg/PK++OT5NcNt01DXwifjXtA6Dr5+YiGJQe85veL/pAkuvpx1H
5FrrTvJ2r+hu11042ZAF+i83yUfMkn7bfo2X6EeyKQjM/kSMCE7V16a1rM4jF9uL
YtJOTjXTkvGmJkCol2n5U2R3IU/v3hWz/EyKLMku1txhJccS8f8wAJAuQpI8A16F
6UX3PdvRo/+Ti24vc5Wg90ntTg3IArmgY/iyREJHPNGQDO+l8eFkRCIVkWSGcm4y
Ot/cgk6lpoqlhyM6GRja7LuDJxlvaRpFuXWcuN1uJKZHgsYJ+17qYGi06pyYSBaG
9V3VYRWtCzK5gsMzNEmoWKRtvVXi5Onf1EjOVE3qxvEBsh6KEfow4WCl6Me0ntf/
tMmRC8ouh03mieOgqnhr8Hyig2OzZ/yLsfVRdBacO2rrgrRIKzu0DRtv0kJIOUQr
BUWiJw23K0HdXkoyMNGbwSquQFk4F3ApSRtIWzcCHWaZdWy0Py+59cfPw4/sdi4a
d+diuNalTRhgEc1dLWcM0C6v2EUZ/AKHSXkt7OxrhejHplfsg4kierdZVLRHjwj4
K2HB/VM/ytgZKJdUa9C+DtbRtuZjoFF0bxku0EVsDaN0SWh96Iz6X3uOtXdxjOnK
18HvaUUsQIDEkpnlBu3ZgBPzS7w7y5HCIWt8MLQRqu5k1eXWqgwcUO5GrQEPfs0r
GO1LSS6/gVx1FeNDnItY9wMp/nXLOBtBQ+Zf4U0arQn4uneZFKYJsL33FLd+/Xhp
mZZviLdYMNDT+WqFJvj7c2FzQMgxujf/l6GgwOLjWSAN5K8vp6UtDpt6j/LK/FZ9
70gmM8IGmAtkYLd/8EJKReaCLSYpua6Px6SGN19bMPEiuDzVWdc5YCfI8ByxlwbK
Y8zBmVWDmwlb1Ed+dHqKPwlVN6QasrJNxIM7PmkBKfaXIAjwxjxFkZzpc2Lo/mrt
T1t6JFtN+n0IWrBhCwNArJAG+AE/QihXNwvDnTVSelxYVY8DYa59zRFwqLZk5/Sn
KhxgfUJc2EhJm/OyRmLtTWj9zSSbToxoY7+hnTZTHf4xYPYY/HcACQ1m162MsG1z
1+JEXFgCUNRy4zPrVJTlgCIsVlJronR30yQ+Oh0xjVDWDheNX3xV/eLiEJRqBSVB
UHu9P/XYlXJk5fPXFGA1TEmf+70CuCa7VDFSB2cYI/Tc3H4zCAfhKYYCOu6yjD5X
u599/HiN7Qf/JZpDs0Fg7jppmZ6jeKcCuQEdJPBL8HGlNUfHRYD84IzXvBAsrjcT
BKr8Nv4M0uU42iQitivqljyzXFXwkVbOslRpCh2SFxlDrAM2CSrlX2wm8CgeXUJc
J6bPpv8hrRwiuZc0vY2djTo5d/rDpwScfK1BrQJSm6+CpQtZEGp7GisODlajmuiI
4cL9VuCaqk8nCcfPcR1RKAEe0OaEt6zKFK5ynsyZdP8zIxUWojLL9Eza9rjFtCpB
eCSSwvfzLM5EJl72lkybP8yKcR7/W2QE+tdmqj8R2JEjp6akzgGF1UyMUe7a5Rgg
BC5PNOOSVhoYotbwkQkCzvkXpaKdUb/9RMYMg9lPpYCg9ae4GzFvw1gyK2oO6FCP
ocGfaJK5JnZQidhJ6lImV4joCKClw9foCXtDyHLw9P/TKLXnHb+9NJUynqZLamQE
GoLwfzL7+UD9OGDEzfbSGfu+QAXk2LvnrAXLW2djmcNOhxZu8V875cY6bgmoBVQG
AUPVCy+vvfTursrDuwA4/YU4ibKHokDJRFBREi3JZISc8UH9br1t+lphTCCVTK+v
jTbGURvtVoAilVbxnfd8v6JYbsjIKWfZCSVMrxmEPAkoEh6exFxkPR5AL4u3pvyH
C/rJPuH6pm2cVLsc9X/LDmikc1zMIk58uBOkhAtMGrEYA9HiXpegsviHBVvFRS54
iRx7FhVN31w7KW3awU3TPG+4YPFNcYNp5enqsVoj1q+Psa70PkBxMZ9TOuh41pwG
TUU4pvFQcVYlroPJEbzs7kVD56e/SuMto67QQDUXTbO2YT1kTB8SSARkTJUIWFWb
5c1oZEz2U7IriAtZcshJYyZzuKVVZMLEmnIGYfOLGSvpXIS+PbqT8EHCG0ZBWaSn
Ihgr40JqH8rZONl+zg32LovWQRby6H5urXBzxWDHUQ4SI5A/78X4OotShUnRw2+e
Mpc0W87qNcuI2/n6NHymTDvanZlaYOXTxFuptQmnVJSB+kYVH9CgAaeJCsWStK6j
2mqVLnHq9vYL5cYHtgtMCzItOHUcRC0qY2AgV1sj4hfDX6jpwVPo0OM1k5vHz2/x
4vFIXU3gLXL+TdvOeGgXeynWHHxbXdjyon4EZh1Cng8FyOzJjtpKQ1X1jEb7JBTV
7gZ5Jop4axsnTcy7vJi86RqXY9bfH/21dRW1SWCMzILPkT0FIdCnrSHd7NFEaX/I
9T97/n8JLtIOwZLvNurnNeYa3VRkRbD7RlDW6lQnd8ythrMjq3iKxXVrHA91dz2P
bKbsNOSQN2KciulAcXuSQJWHEtJDee92IQzG/GzAIlvwOZWnIk2EjScJEqqO3s1g
WhaYiOo1fFAxHDojnD770bQolc8CUKl8zVOb53wN5jqHVB6bE4attVt9KTcO/a7g
7AluygNc3nT6bm9E9YOg3EfDU2yyEN2izUr3hWAtF7Q/kF5oi8HVyb1Rsz0mZmkW
CKmC6W3hXjnMbLkJroaOsqDOMH00+BZNmXLPP/7D4STl0dGJI0rHlA8lHMIKGnSk
ShwlH+k9cPIZ06eC8KsGYnelDnI5jRe2rRQc83vjy1MUJTSSEHBKQHtVh00t2JAX
4zNCZbA9JjynHlmlCHPLjlXXhFaZaS3Qi2WN65yzVLIeC+zNwbFg7HxPCuWEO2iW
26pZ/he2Dhy2YuUMw3CRIAKT1ByWvhgGf06rcINOHZXoY0V+gFXBDHL+h+d8i9kQ
L2SKLwiJhC1sXovByfAV/M1J4N4fYw1VheOWxXT1kmdtHMX4DCdE+5HU9v5np9z8
F9LDsNpoUK+hoPdfyZe8ZBtInuH4yeUvwXKjk3OGe7RUxQalH8JScFfTtW7peO3a
Ig8iZiNgFUkBeeOR2yCdkvO7HVzhMNluOQ979UIJWtRJy9CM3VeNrMAlzrxVhjvP
HZ7kDfEp/76xef6NphR3ZRARVlkZTuFVxicxYv4mx5E71DdAq1tXT5Cy3xG00G1j
GSAfqVYaRqzUZesxZ88hBeXC7bbOnujsGZmwgostBepN8x4fbkNwe/RX8+9+67Ea
wY2w3A+Icf5frLbNSE9i2eQ9+f/KmafUARW6lncoa9oXKBGbRTaz0JEJovZBOLZH
96IcsAYY98rgCYXmD7wO3NeByPMtMYEhqw0NhtZ2q6kPTre0P67zGDPR4ycJ5JkY
dF3AMA3dHAXqR82omBqFlCwmwQd8ljfXvHFdIxxl0hZqAoJdbtpr8eBK03Y0nDLP
/HjxnGQPpoxMFOyIxjsjyzzvGT9cuRTQZQNKAbIqCZEfUoGOGHMOURD7FHYtOJq7
DbrnzrnbasYV9X7KFtzVarXzK7/U9uPTed5sQektNNQSj4M9P4xlhUBdqQmlhMxY
/x8UPHSyWRc2tE8D34fZyWjbUshvO/QUvc/Tj6XhOPNTRsPMcPC6K175UT2ipNUe
zjCbs+wMMgfEArti21VWpQIVyrrEdwcGnvtBw5JKHv4r52blSEssqwFnpcU1OZSk
TluV8NKvheUWLkYWsxiZ65mwYlxtiATcW1OyIZ6MCaKh1kVPQ44iodOTUgQbCttn
xrDK60HzSI79HEUdgkUqPYkUZegFHUIVQMlgXxJ0y7360l4uyXqGNs0Ub+dWru/q
Q6dDYQnKLskJcGJ6ZBPskF8oLiVnAzx72ji++ClN/OT4rxtoNo6CSp1ALxmvzigR
6twaEaV7RK7RCgS3uIa23xzm+zcYjpD7ja7RnkrYHKt22LEOTFpVE3nmvAkkEkgE
Gs/5ZZ0POsCXoWRtfE8Ga4qF0zqr22rNV0x07IAE7OPzajbsHt0Wa3+tjETwhi8/
QPAfPtktT7xbU2xRgCr/Er0JJWsrZi1XhEWDwCoTcqejdeG5q7wm12Wh0H/QK6UA
5srlxye7tNG+Nu/Rd47pFAI6yIUXao1JnIdnCxE2UDH1lFyfR7TRhSlKN0SFtqBk
aRQB1GykHBV28fJ4ClbSM45osxI1LwwNWQHHVU+nnb39p8f/TMp9S1cYFETol0cq
kTqblu+x2dhw+tEwD237GECBgzJIoT/8GZt2NW7GWeLZWpYrdtFJBZoCX+WRi3xC
rHZ++AyALvJHncheFwQnwkcNiRfPJzMXX4UQCq/AxsIuyR5o6jhJV2T7ZwxbhAEq
ztGx0fHlYOB7upMdFUQYKVaUkuPeWB9FeIXFZx1tlA73PBUoKSK7DmOnGgtIkUr2
YXDRbvmX/hSQP3yo/9ahwyHe3F+Bb2PHjlsu0Avm+qqmrBU+sc+4pEv5vPIHd85B
lMhT8u6Tbvx8o3hQh+bw4pQ2bi2vVzaiwKCfy9bsSnUMlFEq+90t7bPMcE/AsX34
o8wG8XD76uisaOrV8T08vMPr96nhNxfL1OY11ncEaaBzhVMrpyJaGFvUNhf1xeR3
OOAhvXJ4VPmJ9zVGl+UHTjeirQdKyDMMY94NTJmP5LI4Er76GzHfZwang36rNJ3F
Y69WFz4ZxOpDz+L1wtONJn2R4V2NzbHSMeaG2XuCdbvVRm8VTd/7qnM1FfwId4T2
Mn5WsWPhzMsfWayHPZSO8h8O0+uIEzpfSSrYQrKyKwTpf51xn6ACdSf0dNlykBkV
E0wV4WiQhhCkF9LrLnwV/vjgC+nCpvQH1BtSZGGB99W+WVD612enQCeJWmo9upLf
gxQP9ASr82T4D69vuwoGmU5GhDY9AcNprlfTpaEpFxM8CbL40PerI84KM8lMaUvc
FHRn659uYAPzxv/xOMESCbSkZD02ouCujsCZxm318k7FUkn4BEyeSd6S4uTjqFlk
3y7vg9RHHbzvrvrPfRrsrspFfxGys+bW0LX/lYwAV6G43oSf76qtlUI7pTZtrxvu
mTMGJ1pqCvB1qPsQluDG1aXnxOAnzdFJB0T/rWQIC/7c/jC1aWg8LrP4XXSJ8jEO
/ARS020WzVBY1EcHgeVGG/pfmiOyNj9itjJu+0sTZ0T4jrETAGfGn+HE0rdkWmwa
TH1cYhU5KIhi3Qzx+qxEw6BUHGcWlbHuHmQ8/ufs1IQz6lfKOjW2K6XBokSwkMBg
uGJAGblMo5tou9l/V2fiKs2A41k3tlTFIMAol+Pw7HaqwxgHiDEd2TPoOaj5h4dE
DXhFTRRaPqxtfjyOg932lofEpVcRSuu/nGakAmLotSoVo0vKBfS+S50x3UMQiRiM
fu4bAiOKRnCVeGo53hgAIEvr5xRST0wPUeBD5n2CxgoQ3gFyMZsDf1LyUV2ptlxV
AlrCzgEAPn8+rto8ADO3LYzzXeMEfkNbmix2VQdOSqq4e4nU4O+VxPToKjlG5OCI
EpxQ47MlN4C0UtZ1qhyEyogz64+xMhpEFriDp8WDGl66hcOwTqe/PeufMoN0m60r
TTtBx7yU/WBp6rXN1SN0r5isk2k+NZ8K7xaGBorfDqQDXF/HYFharqaeYhMdGr4E
HifhXunz1CmA3HNTP4aTXK951lYaLZpycMBxRcmRvq+waHXEDCRQO3msbdVoB20S
QIglodwvf5muOF/FX0tymrSKRedaqDtdepQNh9RJR6A9vVqZDTbYi/pY/m4gnE6n
JhisQTgUfcrzwOL5UNNyenDn61OJpR+yTN1r2xL+51zp6XpAOE3wUZNC0LAZjTPW
xpsDAd+owvb4uN7vs3FrS+0GznEGmcGi3tnv6UCUsoQjBQUIAvRN0HYZcvuNKour
rnb8PR8eKJ/1zVm6f8l6D84Ws/OPhNiKApDLdi3YRlYzgIjCBQP5uHFb9ihZDMHl
bwefR9Wdl0/0vtnNHgA12NL8H+S01l7ZyBpCgClKg3hzk5bSTsdt2EALNPlCuLBi
PhdWZ2xgsJUxT/Kw10CMkifPajshrhuPK4sf2qTH8EaOvplEmBUdwNpYHPQEBYpW
YHoXbYz5XPkr6jjyEjZUQfrY0kh3K0rwoZ1JXt0GDAtbHgp6+6+Ltm9nF9jTJU6P
yGx8KxGPjcuA7l5n2h+tp1UASgo2M9vJiWDQZNpZqhYHUOZTJnGgJL77JRS6oD/G
UW4tf2o8M9si8zD4EpjiItw/wJ2wcd2v7a7nCGUPzYYwvSAqtmxmRtXougKI0HF7
ytBH0NOpJCKRsIWZnqxw0d8B/i8Wz0rCGXkSpWKaREe9C981OkaYXR4Aww/6KIZ2
Ov1cmawTApHOK6EuaodU6tP+ibSdV80yfFXrtnqUCRWk3tkXmh3tpszitLShmLyY
iLHwFV3xT2PGulSUEuWf9WnZ2w7uXjxkodpsEPSJtq7LGFWYlHSy1qBBzYx/S0/s
oTjHZlfIyOv+LAnMKUA0BEsxGYONW013Q/z39wAt2YB6rFnFNEBFOyzCIeoXv6Ua
U1z+rO2xOXw6WKIBjg/fzQ8tncraDbuTbHCd+EpFYs4RIAMKSaTX3DUc9t2CUdYA
7HE5ATSSo5lznRSnbj2x4ZAuxWvvuPWeoPqQnbb+wueQ8InvIwNlVrL6WD9KwUcE
HO62c65NOB044lmB6UGio05JmQ2PI+rc4hHDxDK201hlu4oBRvh9pENimCpUIK+W
DXUq85UEsr2Dqx0MHLcxbaQO+fGB99Hv7fCj4t3Gdv/SYaWdHBArNHVB3Cu9IH+5
xZgsD2DsQjyWrBgKW6U50ZQ055zsklm8BFqpzoOVvcjDCxofJAqkkwiK8d0BxCZL
YP2oYoqEimI/LaPIUPVx7raCZtkDD3zYErbhqvmenuIuzTRwb5ybhgJxDURv4cqZ
ebHA8ThInxTJiUlBGeoelm+BOdf7cX1czcix+daiIjQ8og0majRMpTnsr+nAQn89
z93UYI5BTCfX72U5A6joKOWfHE6574EQZWIiKVW1CAaTnNKbuFnezhC+9XIvIrr2
mLTVytVKl8cvILJ3NJzXdtKzFFI2ehiHUUVWkz3wEeSVofjSy3cGKHQr5pxFet7t
uJqTHCy+vGGVFt4BMVEYFx6LJ3tD9zUycLlZQHxPwNRzIzH3D2WFhOJW7lWJHImz
Z90j6jgILW2tBiDtXNTFZnuoRnuLGQ698Zz6uuKJFqGB2KotWpQpEZ9mtys8a3Cb
uKql4cOPkqD1FMUrnfDjkh1a6QINLllYnoXTSgkDGbtNkNVwAFB7f7HY0Hl2Ga1l
fJuv3gpCWDAh92y+SwDRqAm+9qrBNbchb/mXCKCnMbMB5lXfevSZyjFWHJRwskWw
k+O2fiwoS41owlnIsmcy6CjUG1Q7Ssj+UaKPI6Pbc63XdlqiPRaTfhtQVcNKzvIa
WnCj96XHn6t2+IxVnCYI1jVF49j84Kotjz+Er+39N3PY8WesbJC/Z0csiNnmmuAf
eKVlkn1xO11KOuqfvWrO/jqLGkeRet5qaBeZ7clwM1237XPpqF22LzfLC7RKarMc
p5oetF6ann/PB5krOKGtRvRTKFLuRxxVj0GBhH3lqxl2E5OEEX1xRqx2xNnfYts1
M3Dk5mZ4RAPTPfPFLTmqd1cSacX6hWhN385p2Xs+qEwh9jFcSsPpxF7UZYGd8x0S
K73HtQoHV1ofwXpWhzvPkjQ7JYckm2b+41qZG6OUtq//IDVJwTPToYdDcaCOMzBT
jAJAWGJ/3YucM/9kDcF9vItTRtXix7dv0xuowaXgHh+IyjmhRP6gd/8mRiJsk53A
uPnR0kXXeBIkfOJGsp0nobcgMw/ZctyDajIB1d0mBAijLZBXaGTeJtQLGibcw3La
PfHD0khp50FQqq0FUqxWvmAmlX95R7l3YwAPti55pSaGB7AQhkX3H2Jd8Ks/Fc7s
iBHjX04te9L0WumSevbP6EX4Xw8eTrcWA91oBfV+rwaYPFru1HshiBuCFQKlPTRs
zq13XAMt7OJRFEwSYt5FUORUsRv3iqjDO1Zw4+fQ0xVT6n35Hptsq/bsqEU81nAr
i7aXJPUs8D/DeRjgFEAFD2MvMJy9kGyIMeIYfo1GGXtmPIdX0p0tNS4T7boJUz5C
SqWPXi6Wk0T0speQqwgHMzWkay9EYJnmr27SNqPpIo/LDgIRmNGghNotIO39cH0Q
SITxL2X1QKN0Qe3wcEun2eGxoJk8kYKWwrchuMkY14bMDrlOgSQB8w72sDzrgGI4
jFGED8NNSasEbx85UnG4ZNfunpoVArF0JMLYK0uEYPLcgtKRwaPnVB5MIjwAtTq7
hL903RKK/JwUdzmt6VqgSmlBLPcWPRriHY6N6uoL157TlN5OiVEN+rOy3hppT7fz
BhlIjAupcVCluDCv/+23oSrjWg9HtPHTivogY7jos8osuOli26koSQ7E1FUvvCUM
ooAVtJ6zMoRisGFPNABqOUVAPpvpsM5aFLeZPtJZZfIi3WQewwGNhkWIrn3zjmHN
PLVpHrAotSloit0Du4YH336gPJO/cv21CuV5LxMkHbtdQ+ifEo2KN+XMqJP7ODob
OKpxjnb1ayHNaHPpzb2Tqpvpxf3tcF9WIEon6RCDFHqFtPKmEMqFzkVWhHpJ7UQr
t0P/X9+KaFrSWZeqD7j7ylZxBpJ74GLyeOAP34UBbf+2OI+o93Jz8yluaFk1emRq
MT7DcGNifiSiHjA5Okyx7EIv2sp94k2Y0wCshe4cFmqPL+znmBuSq97v7OOWxvu3
8p8fWoVIUbm8XA0JYknByqUaT+Tde91mb43de0sE1j7+PR3kJRGtaRYdhmK6XUcP
KObDfJfxu8AUwXqRq85vhfRA54SWQyNkmTCEun08phXtPZJ6x3TlsSKmlEDw94wo
k16uMtSeRDvR+pJp9UrxKzzzEphVRtcpYBdk1nqDLAR1evv9z2u8h8sD7EZX8B2K
rp3Rb3viQb15zBPR5tW9C682SGpsRYPdvQQ6SXVneI5zctXyxorlVpFR5N+TAfTg
EmZEBnSmaUE81fga89fsh9ZVVZAWlLsE9maMvCZyNlU1uy0oSftbSwEHfHEVKxSZ
TTGyPJ3BGjWevgzqa2d+zw6+acaFJzxGjF7jtfFUsB2LSUIt7SReVE0qmPRoig9e
yY1s6MpbUrsnsiUTpmiSn2r+daCB5CkWTsF4zSolofgsQ79lpblokHo/vkhupTGw
RgPRSNmODmRS5777qWD+qIuVqgqGERdgnMcR2tM759qeY8TfATNvYLaNkvjoQJMi
vtJyIBV9rZmqZNpj9Oh8y1kd8x/JxeBukyGb6zarXNMabgKUIUOYoo8DgSLiEMBw
TcEHS6rPExhh+rwgtEWBFnVpYDmJJwGgDELUsOls8K0+9aY0ff319bElL5TrCACK
xRxjYKb+k/e7Q3wldRCOblkyDi1tIsRw6gWFB1h34WyLkFCHoJwZHHSIA/xZ5P9W
IIvqrtyUKtyBsANq3AYITGBxLlUn5KvrMIkQlxhnIcphPl3mPI7teVkMXvm3yAV9
odEeOfcgBGMoTQPLU0QiF5oeXJ7o+jimuEtxkmPYqFrkQ6F8vRmV5gr0nSA5vpzF
IHfQSjxiV/VdLQqjAPjF/zwEEMjR4rvrguTip58ehlHlSB56KpEWUppbthxw8WUG
Wdn38jjg/6K8hpCY4P2iIXGewiYiifaTHdaTKRAZILyLzdR7SrhgnK/zX292YZor
+NI/WJ2Q5oiH2tzdcdNkgQx0gMuMCNrqu/8c8FIS9xKWjhLgXzVMbd9NFHdeyXc+
HQfk3ORbwCBNeiAOgEJak0nmb0KzSqJ0DDY2ETbS3ldpve3SwjWl2C1PK/jc3hAW
YrSsy89/47ZV36ayUFzfIdAcSfWprfpq9dw07yCVT85ioFq8XtdDyLB33Sdp0HqV
dd6UzNAUwEjWSM6RqAvPwrcZwYK5EyOlFwVLGlwgHqvXyneiQPvb5NaeOBOb7+Dz
A9rk/eYftmMb7O6y+YwtJj/tBWhqNgoYmJ1bC2L+hX2htBAw5//B+u4Tn7kBtT/Q
PGldjaDzHTy8jiu8Gn2cz9GdlqfV8pUVMvq5ArPTlaZ4lWlleFSLDbuLw5HAgTMG
HZJBsXQg/2pjX5hoWyQeEQWbBu96qIMW3QVmFGWdpnJ5/DuJUkko0nmvcE5wKIAC
b/MaUwmwYzExbOMzRcs5CTS8sP64i68jNLAyHGMwU2yBHFl3jYf0bH2hR9tXwXpl
xnjsW5xtxnNdkgzNBaVjPwwd6qxqE7J5cT6oQmYJ2h356DieOFQ/jzsOSE4ogWa2
494bGNWteGd96hAzGiEGVSWIvsfI+LPsP6H5CT9gfj5pRKWItWC9a7mkYUVpmizQ
8jXc7/uQQp+BjscGhi+J8h58WOhne3YOkwlbxVfxr/6obsfBkjnioYtP7tUi2HFD
yrvhvAz2FuhVuQJYSvR6RYfCrahrOnBm6z8LWSVkyQ2/xrginsiflFS5OFHnqE7E
+1UsxmL2SJBZV6IylAAmFZtYbeDGQVIxvvOPV3+km0+QAGsV7XXijzL0GZsJ7pB/
a32ZYAn3grbzSNA7GWmZ/x9s4eMTWIT6mCu7q2VYqqaE0FcPn1Kfs/EIyBLEHrgG
d3OzlkZSM1YGYuJxpS6/OJXEmRZeh/yre1SMG+OeZv9fO6M0DcJj+BIc9TdciFIc
3JZC5Ifb2jx6BILw2nyJps3yrMMOcQ//Thqmaq84rR4QepqHzgSPDwhk731bHr4F
YVXYx5gvor/HKSJwWWCDsIwS++PqThBNE1skoC6pPtveJ/dy93f/VyB9b1z+eDvW
a2FUiAAq6cH9tHYxMV0oL+Mnr8SukDO4GIps6xnfiW2WdGIoLy/pOrk2aZO9Tlb6
D14RiSJ0t4ct2DJRSXSH5ep4IQHDMFNZ3w7rIiYTVs+YZ9AgWL/bIKxyZGRbpRNY
wzGRamcV7XJPm6hhmVM2ZqAqAg2YAD3kDYBB2G67NqLQoR/WKvbWiT7Biika9OyS
JSXM4hUgchd37cuU79pyDm8UM/RrlNmC1r987GKINr1zJjse2afhGsVR9XAJJ8+C
lsPT036D9078xeksZakhnhTC1VS8SGGgJFchiaIhV8Z0W24RsmGUaoLeajMiQmuj
yn8yTGOyG3lSkPnshw05pFGkEkq7qio5HdsWbF4o/KRrwhGFk/HQiL4rJMTuBast
klNv9Za4AebjQGsf7FnB+cNiBvIVfatZ8LifAByf2gxKMztgC8oH2q2FejQF3nCe
jAvwat6/N+mY0jhVtN//1Vwu48YQtjxwZivJdJUHZespUZK4H9X1PxndqFOp1/uy
Yq0iuFEcOJ65O9Hsybxr6A8Z0TFJw0WhaMGJkDXS3I+h6Q2ocQc9ivA5tQnETY5G
2ZQO+Ox3t9sFsz5gdFcLAy1d8JXcktwx+yIcgGIIjyBs6H0E3v9/F566nwbP1WmU
ard8nH8pahwKINq5ej3cGKsc+o8GxeCloSecmLqZKTuXUEPXc/lh2ttae/72drNv
P9ZbkVVZn1+2qopOoFaDe8Q5hkR4UzWrBBCvYV+1pJ2FuYD3BtHAHgFbdhtHJLZe
X8kddhj8m+A0zYWBMBrNDMndOt10pQFkaIBE0o1ZF+Z8/VvpYDnwGVxSTWR8iHQf
iqHLs22LmousJgaoONBUe+NqrW1VX9L/saBOmiecx7JKh7gAuBnQ3Iuh9BnVFbPu
iwCTv+MRlFIrX2gS0qxgrLDUTulkugJllCesRQ+i87Iy2H1QBcqANRcgccv+nOlt
KciPWYz5tEO6qLee93xAWggefXOWRHrWdAwwFhUWRUhJpC6g+I+jlSLJghJVXA9k
aixNHkcicJ6Aka2uS/REKecXVjLWIoEDPSIOcB0Ckv20/VikGN4kdwd6C2adc3cJ
oyEfylsStmGovQxlCJ4a16z3tIVD0ySObbN0Jn/j55selb81GwHPgk3Bjv7xncpk
/56No3kDR8zwZjGs3aeJ5Dw3TgXHehDbC0/tQziaImgyRbxrgWj+CiVAD8LsH7BQ
tOrGO/ALNILqYNss0GrtBNNbDrulhJYlk2te8cn50hfJSiJ7kFMIWxWBZn7uBGIR
mkUUNre4hMeLwvXhML1T7MQ/qAkK3jf8/2XgtL9T4vugtEWQwstA/gYaYeLm7b/l
gFsAxCUv1eMB8rphTtbZXX2SsK3gtkY1ltG/xF2RjPUGIyBo8xqG5Niz0bqY73WI
MZscfwziUWvyuBeiWIlruDn0XCZXkX976nnqgAhzDs4ad/A2E3LSYu1XYYnA817Z
P8UDWHMwMBO04p5Y9Vm1VKJjU7+GqC49jRH2NhKHcRYQbmJplw2rkaAe+dourcb5
I9pGzJstaxczLGiOt/jnWfpm7vGmo3BKtWlyZ2H82svDAKMRjjrPzAyYROOghSTu
SafKIJAzgO8Hvp/h0mn//YS02Gl1XMoHXt7QXI3OHb0ACC7LWaazVo1eECHyUPDI
q5MiPApkU4lxLYhE2qlLvTSKPfqys5GF5l/aR4NM6Bogf0ps+FJawBsa8q0oIZ43
gDpuDLgz5stDTXTI1hJt2k0EBYtZIlCAWeJfJHtwRFJK5UYJFBdfwIdArwLXyVC0
3dOYALdgCkR4grYikYw7OpWTBVvublXgt9OzhUkt/+bO+N41naDu0UdM1iC5+bQ/
IwZ2ir8yQe11mJ2qhBBFZHg4I0WzzCtRgqv0jXUhIN8ttr9oRx0ufMzBb8VrNnNq
IVchKR8Sip3rcemri+qDyc85jxZJREBFLdyT8GA7KzHQAcoMjBIrq84gZWI7O6Mg
F5Rc5G8aBNnxIEs0nQzPH0r2AKQqNbL+imhbrx1hyMWCJXjnZ00GGku6uEmo2E1/
NkkWiVXltLTR9uCVe09awJEApTCUsYEuEMqiKODKAn04n/Q63UpiEFJxyyfdp9bC
zOVH1rg5LwFxrh0OH+OiTnKnO7W3frVt9gma0CCIihG910fTZfygdAHrjai9UVvy
nnRdaGTdbDJpa2feowldlhatf6jWjdfMWcDlYKaSsKb4RIFwk1sq1incrC9ECxsS
CCkKAkWFD9yK/ELkUagCZmHfrmKX3OMS2Di37KtcQwcByNZFSGDkHqsnMyOaxu3c
mKwoB+4SFaUje8Yoh0cY78imrMQ2OO588rAFQl7C3MLGw17tiXbAFwdfDgrK76sm
y/Ct+/MoOfJ6vLTR19nE8coFjKvBLz2VGkEIvA9M7+QGz+vJIqSSyFikYL4I7SsW
DONROBD8Vv25PNBa+ZYQRRK/QoB1i4HlDHS1qlDFH4tdtBmkHcEj87zJbs3M/X/X
HTYLdna4XjdYCVFxOtPjZO5m65Gb9oUoQU++omXgM+HpbfkEPTY3VCBJ3zkNIUa6
flXdvSrNaWk470oTu6xxl3pmMJuQkMFhchUQyzYd0t3at5gtqjz9EklQpFxMdaxo
U9hEeZG/gWP2KniNpXShHph0AYP9afXs+Hxi7VD3Qb19/oaycMEbDudFAZYuulNN
IYT6LbRwaIry9Mzt+iObO1pLCI86Ec9j3XG3QXtlBxrxUc4Ri7JU+4ZezmhycQST
8zUweoTAHeAe83RJ61HDwoQHjVRqsDsE+wIv7MO8DS9G3Z1HeBizohw7OjkkgLm8
Hgy37jML0aHNqP4BtVezooTZMGD/DhrvwYl5XAgVhbwGTt3mURNOHvls8ApFdCny
lm7k4wkE7Ln8fj9mI4cy7LjSGgEX435Ax1unNmTrKgL+MNadqIcRt3p23UHwVh17
v0VW/H0Gx4JkPvbRbKOxRraPDjy05Nd8GHrAbTYzRRQ4XUvUKoXTQj75lK1BSoI+
dfymYO5hevuOFxW6b23fOKtOpfAu7TivWX/lC4Das2RGrwOwPZizApqgerW3P47S
L7ksY8JHJuieb/fmxtEDyFfLTzW98AFoaecRZBWpwsnXEBxE/Ml/He6oo2YQSL/3
tSrVEQr/34DgZm+YkWgePOiOI+fTI+qg1MO0qz72cbBge9UcinfrsA3F188U+9Rq
UOJYmRDQJCykKluWg2Fc7R2Nn+2jYKqJvy8YeYY95uNnMZ/zod09AogpeDZVS31A
ext1HTVt1oJSVUBnCwCPqup7mIQnxoO4vfihnRu3Tt3gGWrRR1sPLAkZMH8ELoaj
W+V5mphjsHVr516eybHLG0O05QU/md0xX2KmvvUNSbLJ1nqR4kFr4L/SCSBGlRjZ
jRiDmKxXmY+mXoJGTguYUaKQ+BJcNfvlfPt1x0nBQ/SVIuVOLuhmzJwwnolFvLc4
Hn2t2RQBYomOZQg+VawZsT9M8yADB8PMj8+VD3hgT8Np/qKdmG1ChFCYSPttcgNt
9ZWPGZNrKCKk46mgJrWgWUyDbe3TwkRNzdoiu1haGypHgmEzevgeWuenYPa0bRmv
ZURdivX+5ZfKLWNbNP+AQ/4CfCsYqEP9d+w1jeWhXE4JbAf7gFvKFdqmMwbCYNSl
EL1R8x42zEoFMlur52QGNzmyBcRhhkPTM0A0DQjBvDA+0RYbO+7et8kZPlCs6Cb7
wXZ7ubyZK/YKompMMmHDtToCsAKrAyaKHjgkIZN6jbiD3Y4DCxTlgzaO6a/cOUxJ
IB+PpC603dlMHjNzsmrRB0v7kDj8yPBKISq15vVs5+nQUiLhALQaRXc+P0QhQfwz
3Y2NxM3bqjujAS/mnOzm+E83P3biRP0QtViznMjdKQQM2v4rs90tcfYriXkpfoDR
d9XjBouCh5lcHl6gsjtc9skeM5u7EtshOZYDpU7HODuVfWFKbyFjaV55pF14UMoS
0iZdGgKSTb0SPhw/gBD4mmeGjb4VxSCTiG7clqnFKNM5XbMjt++j0XYoCX8iZoSK
QBeRuL+rTYHnDG5wIA/5wZ/3CrKrMcuq3MBrIhZlnm1+Qtk4uViEfKYHFCfZipOa
uUptsrnpw1jHlG+GUIYtWid/y0NQvmT8HMyr5KVi/TwZjiPOPxXsSMpGO2NQ3zFg
Qbc/uRyoP/vZd4skWazRHN/+qkhIy2ePS7psHgJuNqa0a70QpBLXaKRklB49UsfU
oiDn+DhHkh+EgoY2bAJ7r/YfoBiwspXo8fK3Kpm+Gox3arRYNSjXX5LPr7qkCjPj
sIT6AZKPAJFH+V1RRVGoLLB1DYSF85BxOxX/CMOhZUIFMn5lscECs8MPU69HD5VM
fWl/l9YYRWUySiO+5VQ/LuPZBrGKl4WOj3SnvVAKZ3AsQ00FgJPHrJxY8+anBPBL
7QiJxUdtXmCwmi8EJg1PBz555LILtpT8acZcAJalpSkksKsXBEH+P9dvC4629y4J
SfDKAqJLVYjhSco0YypYNMJOcWvDk7tY85h9tcxOzVghnu41GW/TCRRqP+5KIfqv
gxBjTvNPXmdX1IF8cLIR1j7tSHTYulz81KoDN/tpLLSR0uCdJNsdi1VBrdt3s8YF
Ca6hJlhh8FIwbkDZtPF4YbhdJD8ykIZr2CI7yydXxNOMMiSZb4e+b8EpM20UErZ+
rUibxdgXoqex+nwXx80JYV9/t4G6nx3ZnyKnccXuu67ehYdNydYJzb2X2M7bUil3
NxXqesU/lwJ0sw83dt7rAoUCpnfctDJGzZgFm6glfLSJBWlzb35jHZlQlfk4w7TT
pXk1QFYsjdUY9MfQd+ZtwsNLXzZDn25J5x9VNsBwigq+SteOhmhb0OoGRUhW8jM2
sxzXtJzBVAYuESAWoIA0BNgVrFOBSGpzLyLxFj1tAchZl0p2XMrlR/ezJ9PJDN/y
8k8yVloafJTuGSU8K5rCGtPlMCV0fH9TKQeuksm/s8xvzHzJie3y22Kf/RcKhN4w
LmzMfJTAoFnbOXqjrQFYHXtoyuF4YCjeFsk0nH0DbHofW+vMVANXr1ArhmwCwriq
U0jst/onwBczhcLMvR+hPf9AI3IeIl0oBwtnQFT1lUMWAPL+tzHBfF9JuZXPAoBb
c7OFtTayAZ6LSZKG5iWwTlIqBVjPzBpY7ywTzyIqK7cBkvMoqKJDB+VUUDY+5odj
ubQrB+2hMKqzzJQlGSjqoKn3DWaQZkw6Gire2zqJy9gjjG/oLCYNo1uxOwd2KYag
k0SRaXkmcUWYWqPrlcmwBzUGUyqnFDkwgV3FK6Kvv+9o8aYj9HKjWqU5FIpqEU+1
S5xJ1VPFcO0eN4waiM37zberleIqK0vYEKPasW8iW4RwxpT/VdbjA5Zv+9z0ggGg
bz/WOVroACgTRWGNrMN3dT01xmcXqKCNzLFerk8bQ/hU1MDcclIDAoNyBMa7RnPi
lLT9Ocohsqxlky8W8zg7dZINtE5CHBV+ICUQHh7ZfmISmgLJYFXnKn0HZrm3QPiF
sSeu7WP/if+qPDeeuqa3xorkOdUEI9ot3I0rAaFtMjkWJo6wYoxqMDPFre+3dSNu
zAeqWipHrfikSPTKpL/xPUtpcFysiG1opY772avE5bhXlAcT3Lrt0ATdxwJtbwOy
ERzgNvgWlzZZWCaZUwq8BYKY713YwcYUmp/TvxFy3Qy5dB87OcZCIjsGxSTqQg9Q
HYskUZDZOWVeovXKYOWUe23JAmCvP/IjXlgg8QJPAM7nQtulG8KFd81mx+7ryOZW
hq08dUcUbSbMJ8t3ZaoUhwoiE1hwymgfBiO9AHDs2mIhdYN6B7UJ93QmvFzSz1XT
X+nthxJOZzccRpWS7DsgLT9MnpXMlF0b3cO8MCOlzbZaPjj+zAZrkUBa9X5EvH/N
D6Psdj9oNtsvKQ1S9gucijgpA1N9Awa6o6mVcb3OQxB/X4pjQC0LLVjfsXU7xQKh
/WlwX1Q73bNvCaLwqPFtw0B0S34Go+EdWzFNscPsqijC0y1dvEmUt+Vi/ThuUXPd
Kjfwsv8G+M9FbrHCmnCqt0IEvKctNGvOgqzWjrK1c6SnuftuwbqRQ73hMm/Mv6ik
4RTjOYjC/3dgRGXLFCFh6UyKdQsg7toRll6rhGIfTLeWNVqKDqEEbo+59cb67uVj
4JzGm/eLp03nTPYNQrDV69jAm0foVW8YfZAlh04/UKb0SnjJimBR1qXc8vbXDOzd
Kf+FmqcAMtkCm3qEbcVOn1hJriYVbg4ErRPXJJTSNRRyGcuc5W6XYwUtFobPylW4
7V1z/MBR3/DxKC3AlFcQBqRgCqtllQiJq76g6KaiCozYIeHfsZofMyp4i6hLKggz
zIG04XmjoIXora/J2VQOTdLPWAf8vSX7BqVQiBKBwmpjyJjyUUobqNXyjyaYPUuD
EZXb/dz+CwTqneW5MlrpSksf404H+OQI2WarLnD/HyARJK6t902DtfA/vKFojyvL
lc1Ddb5rswQtYsNiraWPG2dTwB9eolzrZ3kGxrtFJCFnMl1CykjINawfNZOJKtk0
nB4L4ECe0wNQCfnEzwqJkmZLJZpgCIvjoISmagtWs+nZB5xQnvJzkUHjnAGEXtUP
Ty6DFoz0uVHg/1n/e/5G01xiN6LcOzW9bEEpjyQeJ8/NBS9dRQAu5iHHzhURqOwd
5aGmCwAZeeC/y3HokTSGr4rgF7iNAitPWigExhYMFSUvP354aQuibKDujIwVe0Cm
/6bJgiYbJbXbYxv2u6UE9utH61AICUnkHv9Ucd/q+wrAnH1r07iCoIpg2AP3QNpp
ytyxkH7H2mWrR6IPKPPCUXLMdR+0h6p1/Uy35Z/VHE7pAQnJbIFsMD8O2kxhH93U
WX22C+svJdBNGkj9GOfPffNxb1PcJA17Slt8j5uKePHTtmijY6biUVlcmiYZ535M
/ih4Ugczv/azxcYRAvORqYC2tL90ZNnEmvNEwRYESF5usQTvfor6VyuXbpD5RPwz
hTpd9Sgq4KGe6aRfPKI1Zr7wBruziF6p+OJjoCWigtLXsDy91l4fnOSppqTQepqe
haosa3kR75z4V/v7ATsS/UT85mipjXfLs7qWytCKtuwMR6BO+RmYaoT060edF7QQ
jWipjkmEEcpz3Z7Xj0giUDGt82hl3hOnOWqC1DWY7aabhEj918yUpeaZmnqcvDH/
RQwCcTcTLKWFu4trzP+XO4ecW/2CIrAOtUoOLo5RQ6K/E3SELfsYpZu5yGrYcydc
iLNAvI4SVE+2UPnMksqtagtDItp1tG6qJ4uY5pPdXtAvz/SCxFIP9rr4Ti4koFNB
qKH/6qjcm7ENauLRsPUTewVNLvni2hQ3hsbNWdjmG7jIhHyes2MmF5mtYAzQ4mMv
e5UAzQtDyE5CrTVVyQxBw2/G4PcouXapCGkoBaRCPxqSXAxYyFXanlxd1Ydaf826
f2WO9LoS5sGjyoeVdO101iBjvbH7jnJXbg3GEGnuJJ4qouJvzazrzIA0de4u1PKM
WDPoTtLtThvigICW9eOIEenxLF7M95mgwOOsj9CBUJlPcolEJN1K4eJiFF0lWz4u
m3K9/js5ZIt3Qf18f+eSmnpAGXR3MMd96FKs/atb4FCfjbrPHqv6qqVHkVAKsxoI
s/SrwTma8RufJYnjv2OPzGWyHqpR2Qh7t8DbmJfUKDUSnd+WWqSQZOOmBxN/LTcK
CsiGMMroyBntA4wo6MEuODXbIAJ87fHWVPqq2IuLGUCKcPGh6jLF6Z7Ur35tV/Ml
HBJwVkOf/CTNoUAcdFwRrayqIz2C6pjIOINvdWKtaWf0hCAz268BygEbx6lQhUXk
XtInYJs3xK8ywGWzibP/QHwtFfReGJpjCkT4MX1ty+ZKVd9BTn06n7pVQccqrkWS
Z4MiBt60l1SCx6NMqxiLFudmNnRlQEOKsqxC4orZ4GQU+vYs1KDE7cmAbty7tKez
n4Z5iXTh+IZBZzIb+M+kQfgsWpvNCSs+1P0j1L9J5hiIbAerJQtTP0+FwRXIcG8i
ibvlJUnYmCMNePaQw71LFEYOFdVGeNdtW8p/UMOZaq51c+ywAOCoafJoNG32U5R2
HWim7IMvPGx3pcwtEMuf622DZAhL5CgGsqQ3LR1fmbqCAZJZwDcnieykyeDarxlT
HmyDqsLF2iQ/EM9mmAwawiGULYEdau+41KRmRVFCFLXi4hCgsQ+coYsgdH3VZeFV
iKLK91biBFug10I7R5cRPX0He6FPt63srGhwioFaQGDbNOYZ2gesvohS3mNQlT+j
01ThksW+phsclnMa+tdZ6ZWpTlrcLI+f0nlLpymAZjdSPtznT2ns2ctgCbikJd9w
klTnO9MBn90Eqsym/+sy3ldQ0wT9cpnOD9LsflDWHyV0ryusT89ZDcOJ4V/1gRKQ
nvq9lelSoQqzcJPoxlXk8EXfdvwkNpb69BElOBxtk/IISzsV8+aUzdViFP7CR7mf
gkrw6QsSIQP782acgGfc8gvcoGg1jnIazDtce9Zu6CHEo+Kqtm1Jqhjeb6q8xLrO
HuIavtkLIPIG1O+7iZxDe8JoFERNgxrdbe1TOla8GEYJ9vpyVllXIhVdl0ocz+76
RALJnswr+K4bXIVa1ukcrq2r48GTBxjwk0emCrHcr/Y0bPd78qqr3CECY7k6gNw2
sCrwDR8wG8KuJczliUhOED31i7bJ9s1/kydgOlgChM5phIcYoC3KotXzya7m1zZ4
UftWKGHRhXBVuHGazaMiQrdCszMhwaXjx9cfRuFQq+lZlrDBF+L5ryTpBpRrCPyc
Tro3V9ZrHEKzJk7d6eCNRIDHrQvV2jT+8gaXDdzCU/r+M4nucdLewJ9Zkk3p5YYz
uAwL+br1WZ1ADMYH7YL9BU5tCHUXDHzyD8LfMSro4jgmCCF8v/tpT/knxDFcZQUT
xnUNp/B1012yi6x5xxWG/vEI2yIk9zYyRVOleNH5pRujsCjdGGIoPAbyw0ZlS4Ov
eJrTR7706G/ij9T1jEjeyin34CVcTE+tGBoCBSgxcPKmizgV342xabr2Rp20sR2g
KPVWRtKeMLG+4johNWC3lmpiLddZlu5HGe3HwnJ3x1NLDm3b1ABeTo0+5dDDS6O7
g+yxQ/gNpBNeOqbchXTpbZtb+qTmm2ButqV8CK4nm1qC5rHFTD7lW5zQLgRK+6Nb
e7sh0NuKLu0Gn+xt8EXAbMSogKWqW2/W3rKewCmyNn1riU+fbYUMqdBeg+me+XS0
vqkcsaY0GtkW34x4iCRDqKubQlIVVPzJbgrmUN4pTZP9k0oMklc69Ygi5HxZl9v5
7avbhEwqEuQbDPGGvAubboV86a8fbctNiPF4TBjI/Q7itTr5lWyd4oeh+IDbLNyJ
/Fpoqxx6GbIewqt+o6zldMUgKvcIxZHbUnExT78gTCoZlVZidKN+IoOJLkE0ttDT
kw+WWZYIgQ8TgLseeGUNeBL1NQcqt7ivlwtXKwQsrClTYT86agW7ndnikiLcA1WX
wtwLjrrNLKikSbVE8m3qY2wF1JXyQp+tHI56iOugaa/bKS6258cdEVzgaqm8Sgfh
Ry9mdOmJIfVG2cT3FoRSC22KPIWTnmkujKgOTmoOsHfBTtxi2ZrKqs3+BOnYBrvi
IYYbzhb6yZRdUZslRF+CPM7dalcPeTYT0HeniTkCyJYRU9h3x6vf47tTevyA+bcS
Nk6u8NV006EdzSgbSKjpFtW6qpTx8ORjnSTIYk3qZHLL4cSakRg0XA5umRNhBcGJ
06csL/lIjAcsqLSmK9vnOK5uFF0a0GeTu2bKGp0VfR2DtzxXw85VeT2f6FHwWIrm
LLrza4iJt4LgP1/Qi4hhkKERyGnviN23yTAhxTUzvwWSrB8+1EPFBBQi7EklvPRt
5nUifr5CKixYcpS7ID4JO4qd1djMc2EaUjSy21lfxSvLCZhiLkJeMjy0PxfukUo7
vMHsUYCWAy+7F0m9cqG8Lo2nKo2GGqjLYpssC8Ak8ouO3dxQKO/JZCad0Bkm2eom
cHqUm9cin6xr8heMq1+XcaYqixKId/FpjCywknywQsEZf9JyCmBHx9WMTI5ylmB3
bMip1ZDLRnFOThgmdH/EFqQHdPGYxsMyCp9vjqWxjiPTWEadsIXZZJETRcaxcVn2
XihfzCmPkH4/olXAJEc8cdpnyvjU8EWBWJLM28+RzFSVAC86eQIZSL66xNYmX3uN
nZtaj7x9Do/eBAuH2EA+uWQFEgBfj2BEjeoWK+wSFL2b/hjiYfsH5VR5tVg98nD3
/SZJNNwT1XQvaUVTZ8uc1X2ZZUyTsw/Ci0MSrFcDwkpq+SO6vtEevkF8Txmycv1j
x3K2a7MJBg4MPt+X7/PodXRXVF/EBWIgCuFWyjcY61LZd4B03jdnytJOYjwQZMkC
BEHIEswZ7QY9LLzezgRvpVG9nxPPde9zqxJcE8gVEmhZgLfc4+gI3hfv7jGBp/Ru
ka0dqeLK/X2P6GWInB1zKNEWfcrNrXtC+gVlL/p1l8E//faGmxDjhPVjGTOBmxKx
tbkxx6JnADdJP8Sp8HFr0Kpq0SFvBjoopEBQRtxzllD2j7E1X0DN5dt+zAaTWz/6
0zhXaUleRqu1EbJ2Q17aBIF2Ev89E4ip+ZHISkl7JwuSW7NVB1IDUiqadLSDPr6a
4WN+4GaDjpqmohez2Aa3u/r3It4EzAdL3Xc8RDNBDEpEXzFSkwrEs+qhdWYYsQMh
l5cjUsY752aOHSTxjMDc2SQzJGh2w/BccSDoDUDmmunmmZrtbEYE4Arwwcte6p90
9m9pc5xo1kLyX7zMR4hr/k178bf7nhRNlyfkGmHmxs1RUNvOWCH82lTZXS23iDOa
Q2EO4GLJ9X791cIeyUQw8mhUzKy+OGWUY+o64ab8y64dgEK5qR7jcCO1+dV8cmZq
AS6lCXWzBNogJVWfEcBAH0OSnP3irFlpAGg94NOvgT3k4h9hKuk+R8dssGviI8s/
CiyJD8rOlcQGtmw1HRxPQznxsD/HcpBoS+X9LK2X5V0zmQL4a692bxll9NnpUjQg
IFGqO33rpl+qaWlL+ub/Hjr6tjPcrMbVgFn3cxnCblq1L6YVkuFATmYC97oJzPyS
nZjjo0BYsv2GCPU9XTbGaNKNDxTrRaSDzT0vF9HSmaMyCFXGjzijOHCK1wLaq4vg
o5X7VXfzkfEOneIE5P74vAIEuDGN17Q5hnoATK1xzCwAnwk+qZhhs48F6ay2XkSX
/gNkGGqI8k8+JkBrA4ylQvv7uoA8oGVYBEqzdSx2OAZkuBGXkxsEC0QttD7IaD7I
8iZuC1Cl9WTjM8YRsXXidg2bpCtgC0qbXDplVXy+w6as7psqn2gFzhJq/tF2ausC
SSmKzSLfsxE3WeabO85xx+kasf3W/YCIhK7xSgnf91tPDZ6Dgk4Vzt3Il0RAXK8P
FRFz6gnoYEp8L3Om24Niaa3VaBr/+RRmurv1Da/zG7Ib/A7IjZDc6DAEaR4slX86
9Zu8mJDlYplgrwx/tyGZdOaOKAswD1zC124fMfLvCIdiB8KuKgR7M02gksh3plMG
1aA/7XgMqE4+wyfoeOsHcihAiB1o5UzTs8vohoqYai5x4DQH6sIitvQrK5Gdx5Ai
uC0oy1SwWJuHcEkg6fL+8AQzvwrLlTS7gsFSEFYHIbd2i9ja2n2NYnug80hshfO0
+ZMhCXToxIA2GYoDgii0S5eXSPssHJyo98V/pkuNGdQvWfLCD9xvOMZ7StW6ZseI
SWtcbAWFXrtkGdGCKouPE1gm8rbEI4hIxODqRCCzyn+T+PKcjfwXJeRvzV6h+JMh
zS+piks/Mi0rq8NqX36XT3yBg75EH7i5ZG3AadVsXpct1QEEa6kA22ojS3gFY3sT
HlS3ahd89WVftsqsUbAtCf7A+pe4njR+DrTrUyXJXyiYXfLCakHYk722lHSf0qUM
zdLycSGstoB/IP+uz5UeNRmGLD61uUKMiU9eP36sCBvpzuT/x52EuluxYmUysKU7
CYU4qW69EmHk+3BQH1PuglTpIy7g/uFBlmVKqBblNdjOdXLjZ+ojt/nNabcnAqUz
Na+PWb0qfgJrCncJz1K68/pBrgBhTZFTpowHkybIzg8ZdWPHVLXwNI6fKfg//4R1
MCEQMVKE68XDlJvd8KYwoSW4OUjslblSdf0y0YkPkpOXWQMLZ8LU0omzNv3Uvx7j
RctlmFmUghh+HTsBQZAwKAa0MkowQmf2C4JZkWnoxk6ZI/XNIJ31DH+AXxrq+6DQ
RURk4Tw2YZPY+NwKJ1P7B024pFWLvMLvQpTXbkSZXtGed5kdyaNS+BqPq6OVxjJ2
5H510tUmpn7tcUkZEq+H3L2zo7MNCExD4Uh0sAR29ObSgDq3IDCUO9b6BaAAGvum
D/Um+5cysaeRbw5jV6vHSxWFugFvXin1H/uevFxe0BypHcyp+xqqNjvP06ttFDub
oIbufefo0FLX/XxX+PqQf/SmblKvHQ0Oy/Wwmq9fj9uYo2k2EudAkaxMx7tP5Gjw
xam6HKphY/WYiHvrUgbWcJZpLKBy2nqfcZ/B1z2HF+hgQ9l8PplukGbOYruMFHi6
bl+ZQlKgzGuytr6bRDSd52Yhi5ikvvtaIi3ppxVeFBAuE09rXz5sBhDGLDOFpk2S
buKhYSkp+stTjji4W8/hcrz7PNiXIpQuJL7GNw3nBmcY4rQdQrs2fZAfdCOoBVnn
JtmDrDrzQtmaPsWpnGvTJpZfyBuwXErFQ40lkvHkjiHnnOPPZAM4d8Xff3ceNdGB
O6r2lHO52ocsk+FJRxRMRR2F7YYFzJ9jdM/xToBKPxRzNvmU5gtGPknlF3z7TIk7
4We/J/6A1gRjRQNSJq/iFz3SDbEn/483TCSXJwSdxpA5NUwe5tVwHTUQAvvbPhNp
bp96NsyjuBeOoI6gLfjcLIW8VAIboMtDX627q5Ea6AK16AIKsFIKOu68puMIyyh0
68AkIPQaYAO20hvhM3QWFNCL01xwiYhfyMhf4x6TfTaSyKq3PSTaNWlVI9dLGPMP
SQKpzGtsyRceL3Vmm7P2SGvaJVq1+gEBoxvLXgmHuvlDKqQCEdwsYAK2/lkZYZcP
ANqB20/bcDPIewMELUgupruuIWdspzJKCB4cmr99i5oL2w5dVK9rAHn+pgphSI3E
57QzduFfg5sErslIkRFqhYhcsy8SwKQ30cKO+i2rwvbsyetGRYZorKdHKgfDdSI1
WNbl9j6JLy+cQPfQqUA16+aNg3YEP0+w0yM8dC2OTshhn1ipmSw7yGiotii5HhYh
1yoqmwnYbW/QC0/BWm6b7JzgGDgyPSYbFY0nzk5mgimlJpToOVrffeTOkAOtQwei
Js6iaDupYHN6k5zWrJfSkHWARx+4v9OANhktoHNdSB8/yw3wK8pDzqjraDmR4ZXN
r//jEX8a2sK7QLU8Nk8sI2VXtD6mfC5n4cqZaUSUAu26qlBgYKKS0+WobAJb8IXd
VmT9/rzqLQ6TTGoGIeASSlTzP+0rJeewadaojGKA5k/3q5Upfjnm+LIyoCw7odv0
oqf3eO1ZnK4H/39r5dVY88wrziyFVT9OWWPEHUvtSy5ZPt1sM7Uj/mvutf4WmwTu
T7TwavMPkmVRk6xDfIepOAKso8o+N7+omUizkDmZYMcud3kjPY0mAWFrzhFsnDu7
RBwBcehKfA9QX6qHH8KCmMgeQvHW2g2g42F6Z/hN9CDfYceolKht0Sb85xUrbjb/
bXR8/JqHkxoy3LaCSzn7EQu8T7wbgecIukqx8wHn/r+u0dRJt2JWrmdGv7NNmShL
cO9VKI9AqYhChm/6+CxR/w3gI3pJ5i43iYZfGNINqMNZoEIrQtJdP6z5R0dLZraO
CQYYABTVLYPYMC/2glwS/IlRay0WPYZJpQT1An/+Ula1ZHNQVMMr6sOZ4Jfmrv7Q
8HVN9hli8td1pD/BXiTgg8gmpfhKYexXg/bPNkpu5m96mt75b42iyhFRR4TC083U
8ypaNvzzJbbvDNecBmbHQy6VnEoi0PDaep75Msu7dz7Iot9u3PqG6YZcM2w6ojUg
pwMr+VR2yYAU2MhLWu4AqlKwh3M+PlIfG4F3rDB3LfEtN625TWMrni2StthHXD3N
DfvGfm6KLAPqqWbWxB3l810+H1eqi5GVv+729fLGJ+X6jfQtOoKd5DYLbWx1zxmO
nRClD4rkxnOqG9PIgWri/o0qD4qeVyEDxe7ecQ+4G7A++tatd4Sa9vPlhMyPBsTy
k0w8ijvQ0ge1fgM0MHiqs7hXBNlu/zVGI31Ge0BaWnSo7erAw9OO4JXCyXp6x8Bc
xdmtsBL1VwgDh6iHDXPo9jBQbQIJMuvmXeamXeD1x0WX+HomItrU4DQQd1QqYL2o
RXq9+O3bGQn99vYKfn3oIc+s6SFEAhbQlBBQpxTqK4R/BVZqihHp/sIxhQMR4hf7
YjpVPJTuZnd9P4NkHXwS89d82UHVU+PhF/oYUY/yGrU0/uX+HjxblDLRhnPOH+Cr
OONWgXe9hNnsyYjNgmgESvKNEmO0yNjq58gaJynHfgUXBSrELAQObGRPa91yO3wz
r2JlU2g5nof6ZsNM8/TiHhW/8JI84St1adupH2EQHILZH0s6vEAErp8r6aQ4mFHq
4QCd+cUi3BuZ63JXKki5eQuDuyIhYz7WJloJzkh4vM37Qg9FyML07yr89XygToXF
i1sHY2G59qAGm2dps8N9WeyFVY2amXHdQYUjU7PSsSyjZzaGpm/3ZrWEg4bE9qoK
eEPzoJTmMhuLYCJPK7wHeetA/UwYYMkXYm9gJzmeylXvUJxDCtj2RUzB+Z8pJlEB
x0pejZNxztiIqxG6cPeOfM+m32u3/iRSvmOuOZYn6PNJN+ask9YEihVKxlTTiyJY
7v0Agkzv9OqbrYvHbNlm1kqb9XVOuJb41KvLkTPk2+T5tq5KYHJ8zpclFrDqS0q1
pOIC0bVYZ6pxSWjjWk6dRRcXOD5eInMlAd4qrradEHyo/babhsYD6BhAftGwMZlR
AyK/hzTKyfY+ybB9gmgtlA1tMz9AwRoDD38H51uomaLy8M5SOEeHi3CSz7Eb8tR5
8ipSZt2MENoUkf1tYn7S4j7bzGROnz3/oOnXT/IUu364/VmWLEc7CUeo5z9kCZEY
ucHcinbyUJ9Zm+sGv/qMPzLKj7Yeoz8YEH2x0W+Fz1gDVCymR+5wbPTiRfTlHKMz
/55nJLIqnyvRXdVYver04cdGKuW71pC9BAbvQrn3e0LV8sRn1R6Doj7oAnBgOfu5
EUYV9UQ5b9cQGCW6zXs+wb9TArgLEiRLWaf7qdnR2zBdzTEtC+YeX9TSlmQk9xlz
Mnuq8tIfmZZnKc5AS7qpRzB6pu1+GWITtlibOz2TQAKDgSoOAWYvyNuP5BbBPkC4
xYJYYnyhSNVBj3MMLRtyjAPJKd4NDp85QPY8ZqfnsUg2lPeKxwcXs/br1gFpe91p
96IaTU4YaXhxj6jd8Bn16TJpCQM9I9Y/4X70KkCmQ5A4/ScsoNxhPP2C6w9UyigJ
oLbpFQ4/iJKjTGy1L9qTQ1yEnSYmC+0inShi127R1Q/W0vfYUWXAvvJGixFQfO47
Lsxx2gdqhYEdnD8SO7ZFqc8jggw+mjGx0z2m86invIGyUw1xLCGFG9Lb05zn1dM1
ibl0Ts4OTuwwOWSuDlJeK+t7wAcAD+pxDQ5cmMOetUkBMgz2WYy5a5Ax2WL/IyVU
FXyw/xhb8ELtzuQ2MeOy3hxpGoqi+E0z888oOd6q7fxzwnc8/Kfsg4Mgzv/m/St6
bR//HBZ+QjkZvB2sYO+67BS1Fadu1Yv6a0rVoqqd4oX20cYB8C8ZVQ4TQ2L7e5oi
jWkTSlXQuQubZMhiCdfWs+20i8eD6S5vFCSdbdLzQIHMRz7i1y6Qq+x1q/kWBFIs
lQns84QDpCIDE9U/H7PZfNR3lTKDs1MVVuekk4CBSZeiOaPApWu/WrISFPauPkn7
APUyOIJBMiDtNjC9uqaKrbneGzUQPQyvDylXfY9g/WucU6QAANn95vepYFllTnI/
E4OKTzBilBhKENLgNmZ6MOc0/2hsj49ROHl0wFKzxN+Uonzg1v7Ujg9JIGnmNptr
3DnwYg1+9Ls3sQo2CpqkMdY5KVmN3PWHxYjPq+jgJOGsLX5t0ZraE35mw9k4dqZH
EGr4FLP9PZPN6rjbwKLd7kK7Ltwv2MmdsmJI8E1BLsSWeYjZiFOfrbBqX1tvQGQm
nDe/ziLUMPRr5OmWrxc/SxGGzBj1lkUszmMgEAA96ugfA6e5HG0y7t1fvgKXq+sA
WOyrLe+oDVKQHhi0QKRPAHmn1o3hEQHE7p3LGv32vENHccZCnEVZmk5peciDUNBA
kNfbAcXlPDANZFZ0jSZd41Sot1P9AGekaPaBqGzIkNOTgU7gO0tFy0639jU9Tg07
ltedtOWtL2iu52gOcMJj3gdqyelW3kskdj+rXrKxwoEeOOp8vvH+BWDjb+KGP5Wi
eBTcmt5s4IvElC+zfnOFWYZUDNxEyDZoLUrSmtEKkzAVwUwEF/t5nI1tl8rfQpl8
aPhM3sFmdNekFC9nLOVmjx/HHkEZDV6DwgWPoPJt8OavR1ojbPRiT04H6Eni6Hm+
+FFS7LQJyc4u4dqqvrQcU4unsC3jJkO9KYnMlZQJYhNSSZ5q1G9KejK2Fax7uxI6
959gucnTs0bunQ2It2ElvVHAY/VDGBmenOuwURKvUJ4fnffhYhjqxMjkj3iyKrno
/BGkPbSb+mVVLN9S04VVHzNhD+x8dFp3Cqx4DTXQ4Dgb/TEVH5t7de+bZS7BC8NV
/0I7VNIEBpuXXY1/BIDeqMrRrTGHDiG2CNUs4UTZcDjS+TbTb5IPFAis5E4LD9k1
GYpANTIlsDMIpMpzXx8Av2mxRnueM1X3HqIPhvnPaIQ7D5cFnivrW9RB8Xxqchuu
Db7Fb178y7W3hqnXNd6YXwxu2mX+J+hKAignUhn+UZrwH2ixjEn5f6E3RDdS06pq
caveeK0Brxf6fUlx1F2pygkgvPV8eedLzN1RxXW+1KDJuIDe+DSqJS1YU/c1XgyF
F8aqk97VZV657LUOiaXOgFsAhazWi03w/bs7CW35vaNC7+zf8NkjDkT5lsAsfD/O
8f7Y36GRf+MJqkDbqB23RIGlWg48PkG142S8imYCF7Fzv42ggQKfHoqFH2+EtHAx
gfI9bmglKPMXebRDG3IJ+9Q2lEV/mALQcPSbhuEzT09AqZamLpOC/GYuExxRIcBM
rF6bpxsIUWmOm2L+yEHPKGggrUxdInyf4JPZlrxZt3bT3ij02koQegGjsi6nXP2C
F8hr4g9iX6kxpTFhyDHtBl3OWgon2sGxK8CgvuuDB47m9OwNJnIVv6hNMkjFX4R0
w9REOJlpjsCaiaoOQCZPJZmEl7L5oICrJCPKe4eSXHb32xFiZ08ty4PMIaB14iyH
/jvwZdmm4oE/i0VURPy++hLKbeKD5UFKTK3a57SWHmwDAPbhciSZKETNOKPMsHwa
noNHvPtEwugrR2oLvQhGHu3lMQxjp2IRXUOdIhXek8mSavMVJ6usZQSZJmg2QuxD
d5tuU2zpgQvn1jXefOpEXX0KN0abO+OFHRcHvH7a9yGKnPYKHjWcgfr1Tsp6zgd/
qUA4Kbfm/CVCUcHEA8ecyumBK+I2E/aMHxIalUwEb0nhk8XrvkKpRAi8iumpA27j
J8qKMjECFHQlwpfEVt1LDAWV3OfaqLGX04/xjAF1+i86oZIubxa6mgChlrEUl2y/
srB3SkG45KgEr+dmAkSFDPJZ2plGbFfC3LvuAOJtgejz4xSLEMCd2x/2ovqU/oHl
jhXbDVRHy3Fgd3z+6mFp92iAqZi3QQFRqr20SnCQ6BiYLssEgnIsd+VK6CqZ7bhl
wPql+qcNb6tezzaeobc9VbgjNAiXQAVcgNQn6ImOZDuzzrd17mVhw/rXjl5O8ZGJ
v0qLs1PpQYR3h94OtVDaORmAHa9rIQA33GQHUX1vHm05Yqt6f4kNVh5yBYm5DKKj
faKvUqdrejWqiah1kBqxfyq/FSTjj+otxg9/M3y8oiXeio17kpzN1byeC5hZKsZm
SYPaY2/04BliWMn1/zcCqItrXEO1cySNoFBRzbHyBbzpl2fw4e2J6YaN6sjLHmk9
P3K+XleAlfJa054z2yaJi5Ox524TT9noEptNRKGhbEQZfBTHYI4YSm4SVTmRbsC/
UHj3CXLtxtGBrSvL9RCqrIj+tl9WBdzmmlfu6kRhs6JHJu5yhGZTCjufgDWNA+V4
0eg7jOpd16CqASS1lI0e0Erpo3RB++1YttEUgnV2SAnsqHx13f0lWlSlOyg25iFm
kxATX7Sin9gSKt86r6LumsBuOInSOB2mCl4vIUIfMhTBwoahD8Gbe7JQs/IXjLFK
+rDRVHkjpiff+rnHxY8K9Yj4OALWl6ZOP4Sb+6kMfHTQ3KxB08mjxsVcPMwiqQd9
rvzwpXh8ZHby3qbMm++kWtTeEsgF2A4OcQ6MIDUUZ9067BACUn7kP2ZGyvxmzrFJ
JhqtfOGHvCyG51KkZUVrKK0EmEY1f03xGya8FO7J+o1XXKZxnQeNitEP/r1AwoV6
YFZ7p/qf+s0QA/mzsxgAkrkq0OHJ4BHDU0glK2PNzMGRLw/0DL+KXTKNXd92IDxy
fiIASbCiKpXOGQoanoytFOwiO6+d5FTZVQanpZQWX29rnWROwn/Xb9jypy1tOa4k
svFnNR1PaGZ7vfvuuMn/aecqmXr2faY3PzSC2Bju7L5I4VlqfMEqWxWv0av2mYE/
cMv3qyOoHvsFckqXQ+nhgpz6nyPKMi/HzjVEa3T0h6VcOxTcFz+OoeEufyrfKmDM
0Dpg4kD2XHywy69uB6lZLfuZKsH+Yk6Ali2yApGcQLaHcoZNX2nPGAIhTR3XIKgv
/S5OhXEUegtf0dIpVq+OuYEeeE47o6AX0oBCeMOOM3zUhUQOwV2qai0l1LjT0AKb
Te+eDjSuyAr7aZOXN4VHrilUlEQgRdKL2bafoNJTiQf0UmHD0gJb/LbnWcHCwfNn
7lC+RNJDpQ6QxBlU1zFepX+BWFfRUKhN+BWLIeb8sW5BxUY1IzKUsxA8Ctk5akSf
gzvxx0Za+At7dkEG1qsojmgOoQ6eB4XWHGskZoDRP6x4aH7W/fwT3ix85qP/Z66f
Zfx+Libytm3PklIaM4c1p1Z075FhsGl+/e+jGS+AWYe2xdQlnxsTRgdNRTJ1FWm0
7BWrUWiLOCVMg5P4TdRRV4sbmNNf1Fy6rPsEs66X+a9d1aYM0E4Bg1+NwPuofill
v5E++0ylNRrB10+3B07hKCzQfPD0N/m9ECm2la7aISgFW3OfIlyifJg1T791Lo7w
Il7VKmAxCBZsc0NVE2fZHM5dDxFt301Sz0HOrDNyyfBL3x4p9nuBDn10q72GwcZG
pBVJTYTzJiDQ1Ffokt0Ys3zbQ4PzmFB+zlbY6ltV9AdRSGrwCe4OqGZbmAQ79zZA
EfpvY6xcGgJSHVNlpGZlE+33DA77kNhlkHJD72lbpRGkoQZy4Z6MLVc+NyGmed3U
HwlT5BsB7zTn41Fnj+Ta+dJwpQh0RQCOcP4ASIO9waA4cxhld9T2OgPmJRQqTEgi
qzvnF1h2Zo2+ylLR4JGXa4Fpc6L2AuiBMX007+QVg2reL6Cv2n5TUIdsG+hCQPc2
0935jRr3cX0J41/04W4vqYnXrNL6a8e4zlfFYoHR9x7R/QM2Fx8DEfGIxZD5g+Sv
w+CRe0FuHCDxJJM4ZkQno5RoGyv3CqwJh1hKQgIWEXhW21r8Pu6rOK85zjh0ULDu
B2hTFpYz2gd7nRCha08ZVhukyEvzNxKOPdw9eYIuPWaR3BrwVn7Y1DAJwgQqEInz
euLz8F9HDd2dcibNwTDVaXHAwS7YFRwvvG3fqLfpTCEIiCrj07yuRKySM6XwmcI4
Td2qmpavzGIQEcZDyReM9LF/gZpfYPjDdTai0LE2+Y2RWfzw1PkJbGnXQ/CmMRqK
UwtM5cJrkPGglpxcJQvjb3AeZeu3d3ASehjUjsJ8QNEH5OCg+TOo3pf4IpwjjvBR
RobeAv5yYz9lScxcFGMF+3+3x+j+LLRb3tCtLBGYTXgmnYhr6G9LEECgR7NDQDDj
2WF3lB5vhtGMe7cWQTTEt2GxSAompVTVaOLuThoQUuKI6d0BgIXV6x8yMgFxbtyv
LA4AKGgdQB5pmiVOWV/nfPG0prlfFz+3E84aEnXR/LbvMAjhbkYg2/deqnjx2dTc
7l3mnyfPlEZBzoLxtOzFF5rpGxTddHvzIyifDqCdL6v7AnJ7LIRRSI/aacRuaot5
hKW4fiBrBgSlC2Rb37ME4kYQvS8Rbwayd/74cJ2RTrg3vmngLIgvWZaHEGyIzWJI
6+Gfs25rARmj5185PRI58UXE6QyiTO+PbTBQ291ityx30/OKG1SIgSVbF3TC7SCm
9e3pePgJ3fZwteXwOd0EYoSMXQieD4UKL4fK/T52ZQrJyEXagd7LeVI/vuPYFMSH
cKlpWJ//FW855qiwS8oZgWqK5KLCZkFSn6wZn0yqsNbZqt2N3eIySLMDMhD21u98
o1h69UPqfJd3OKlrp3/CDegNI/ft9Yv6pnZTRhiesy3EEShmMVjH3WWe/q8NDzRv
AULg1ii+RNTZ38V0SotJnaAnNF6A5ygiu1SAHU1FTd3PeYN7S70CdpTPMJ8yAerE
FbkOcqYWiP3MwFFZi2zjMWHXUDJ/S3f5r9OHNQHEaVmyOUjcZQ1SzCIHM+uTVWWu
ODlLJ2Cug/KlhEIGdUbljCMmmwstNS9+tgqIMkoYCZMaLdIf0+asbbwwS9nALSW3
wjpA46vkN1UDBeyNbr6oA72RPIWtReqVK6n2FVc7HPxG/t3xYcs70SXD+mJuIf4N
+2QmAGgbjRRZ7rSGLF17AbUrjWsoTugxGiDNvnRAbo8QpxsV1RmkSF/O2WCOOHO8
hVfrGQ1K8XGcUG/bnuAXXPMw2tXZk6n7Di/4aGf16zN2lGOrlz1NW0DfEjjyOe0o
mbrlaOJpoDDRvSDzvjsK5UPYN/7q7X7n7HwQrA5HC44VucdhB+YEZYd06JiJUM69
CS6w2XUDBkbBkaKR3HeYonf0bo+ym7Y9YFRhrB+ENubeiVhTUwYE18BgFzXJmhQG
+pd+zsJpO5z0wYSDxy7mPp0w8S4rSKbAccz4i0MoYThGSHJ9eh4h8ktbmnSpSuZY
8cVFSzamBL80AGxtaTk3qiOLWAkilYebWQeSfTUNTBRkEZTvPWpWH71Uty/ObatV
bNwO7I6ftngl8UUbm0LMFo+XtA6Fg+EyDV+6pAKKmKBUaLZf3tygf9LMO8ohmMuT
HNcmLG4UfgIkr+lyoj31c7e+pDKlyGpM9e1ctRB8QAVBzuevYXEC9HAH4kpyjkfO
3/cSZFkRtUw4xLTRcjI1yJwIpBjTqImjSBO7s4UCPxHXAFPoq2q0yyT1yp46u8LG
03jQugoEpP8ti9sFwwxYhmrnRDn0xcF/6TQYjCr96vDFbXiX4qRMHSRMOcJeW43S
5PRdq/ua3OiqDQscYWtbmjAK5amVLTdxi0cwMicNbLZmIpOHViSDuCL1/HOyKRvf
cQ+XViJOjfQh0eh8b0As8M1DqynZQtWSaXoNAZEUVa4W6tdHUICiqe/CjC4cSSET
+0vL8hrjSDR1B7lP7NJEusaUENtZXG/A5EEtBMlShcERmbAgwOTW+kREl+WLwtFT
NQE7nGe5nn7bYS9bDtuWUXe2lAENMUSgJ0wYtZ6ULgqt6MGQHafd2f4gzfmPXmR1
cZJhFqF25Npl/KGHXoZsAIo5ltYHsQMR2SSQuGgBr+0pLC8OA6Mued07D+gjSu4M
BQLNI3PYqVpDjP8cUx1buQsnJ9n7bWFSZ/vMIaGwiW0gg5ZQpzj3kOfUWpm1E6OE
RFiFBZZQ7Gd8b2zvzPA03Iox3lGEFoopGH2iij69iLzNabYIkRPUSVKjkuS33R0l
ymG2c25RcfLj2AMNPUFcAWU2uYnSTLfsTg8c7rGWz1KkobTVRHriX8Gq3Ux+1FFh
MBq0DfdlR8IDvUBNcpePcoZsnM2LIbmk+Z5uXpB82G8TA4L0arm5hMyeghRXGnk0
92hdPtU2pDlV6MO6An1t10Fe7F4L0k8s2wJpGLyi4lgWUBoVfymDtGRfwDAqSbxH
VADyJTDGqvyPSuO/skAc/nNvHpyydbR9+s8iWV5Vs3djzPipjHpqG+JwvZjZjGpw
0dMwLsuzvu9fUmOQTGKsfd1GiiYtvh4BfznrvlveW3Z3lsQ6vJicMkWq8us2zwHV
LvFdZnX8Wi20OV2rKOi2FzfRHAtqU2YvBT/xyESO88RLeV1nj+78tzvYUVnjaTad
8vrCpN7CNzTu8QV6PkgMiz19/vmA92+TE8x/W38i3oclTelZ0qSXJjxX0/naPKDE
W2wGbj/Ig6hmCis2X9rm/WQCXt+yPDDjG3VOpxS1ezOSoGZbf5XXUhIfigtJX+hh
+imUSOiunolVdwkzwUurAtO2774AgAXIm5pCRm8Vetmp8a7hQi1GrPBn4o71Ssgb
AkyZFDPNTNurofedcNvnS7NwHiKme2ql5Hs2RmhwQ/YyqcrZqCppmDmcNJo/6O7d
hLUrt2emK+iYsSdzfYoaRmSFJ3HZyOPcUWv8AX3y6naBUgri28RjY5AO4/WUaSNM
Re59ZtkuZEN+gt1Y5xC+eQKlvyXfVWuDX21KXGzkx8BWfvnomI1uQrla89Gkm/Q+
H9RcR3O351w1oKWcTmhucULXG0HV9TiKXnHfEBgaDaHypI0X63oNLs/Z/95ZkcWg
lQwy4KYjjfVaM7cDTGjJa+CczZmuQ41V0cnhM/l7Hq9/lybTCFayH3+FvyypxlHw
ecJ+6CyD2+NbES6KRc9ON/R7FLwUuG8TxQ5WwzIkcSZCCNxRIvlJ8dauRYMbqcTI
LC9p3iJNj43STlEn91POJOb/heegoTHKffPqPzPzvvpN1d5u6HyQdsYob0W5OTdI
peFjkZubKujlbXMhK793O2g3Fs/4k+ifVaccNFWqXi2gqwTH+yqgv8gDTknWQl9L
MPd5VI4p/iZlul4bivDi8rkUme4UMnIiO7ELR4Lx38/aBkGrOEUqDOnE9RVGlmFk
SxT0R5asKtFG7TgT2/q/jOnez+BccKLM2hVm+GhibbRA2EXnSoBLCZfu8vzdC4ro
1WXMW1Ld/7YmO3JJiRrMl7H1nljZxHt2ZVfLwJuIMrpDhnXdsXrL0RKVt53Vu1VE
THdAneimYo42Tv5DHVtOpS3snR+dgpx3S4T1AVbalnsfSWUl3I9gyH30VviH7fdp
kbi7ikBV3rq+N9ZwwLz8F41eq5vdocAt5AgbDGakxMwD4Y/RwMFnUVSIVk4qcbof
0QrTngS8mhu6u2BM2h31TdE9ZD7WuPoCuhVZ1HMN2O87mFUHpPR4mhdrqVJ8iwbm
o5wV0qqCze27VUrbP/o1fZDtxnbadNaNLBSbY2KWBVw8fZHr/7TsJimcdCzebVyW
7mUswElOPbm+84EtEQvkXf0gMCteRqvdW6p54MOarueM2wj2DgqmPizXBHVD1Mh2
sVNUFfW6F5c59cZpUIYsBiZxAs+/k4z+qPUlL9QWp3hrUkzwpYFz47t7WWMxgJw3
Lp1z5+NJMG+zYk8fwn60pCBSWyQWEhYH2Y+n3pxz9jyGHIHkZAt8Wsi+o+LL9jH3
QKc+2SuhXQme1M766UUcsUn2caVBWYWTSWnBNR92cy/lScQ7P92v/E8rLILEhILK
q6dxIe5DB+UkBJLWJCYUbt9tqJ2g/d7AU5TKr4XA9n6BRN87dSwd1MrpiPfCulFW
3Vr2Z6k1FveQJtz/6MoNEiFp9YR5mRaGRn6nBFh5Gxhm3wmzRHtuSH9tslxNYV87
yOnHvBh0eJlY6vAXkRCbD9Cng9Ys7rmNGTyHplZQmOicBW/xd7Q62rEBjXzEEqhq
5d/Hg7TXDDWArdKYQl95KInB1EM5l/7iGOQHw5fh8l8dmBmXmWfHJwi9XMgR2U7g
It3efZp/tgSgRvT+FV01LSf0JJwoyObeZF/2U8PX4Z1iX0g3CmY8zMNTWK1XocDN
nKZes1Lw9ICHVy+ZvDSlaOhLpmYGS1DKZaXV5uUzs8j88miMRfxMzwoRNLvQWdt0
VQkmfXGBpSidk9OUsKnir4l2ZcI+SfW3abWXQiPMbCJ+R1Rqb/eTVCAEa5g11T0t
xnnDgD1q9TzVY9kfUxQX1C9ppC8Nrk4l/xYG7m3c/HB0AscxVJM3SGxUuJFKUabr
AvWCk7nNNIAC+dvxnYxV+hORoQJcnYiqEEVkNeAqqwUT1BHpoONfWCb8WvuuFSUN
G5MkneDuucoNlpwy0BwYTo4VHI75IwpnHQ1sG4xr6gDeL+dcfBXOXFnYibsoQeYE
c5Uvc6zS/oo41R4f9HvJ5FAn4WMMMoHM5udCmbFyHLJcB9dOiSchisdoFni6Np/c
1oVrictxLEHsfgphlD/bZ/dH3++ebR0WgkGfsBrGTUPpr7bROcEbB3CqP7VeETNG
rqwT7nD473YCDW9rg6LnWfULGh9icIMgQjKvxZ0XRjSBpi9PSKfgzYoFN8sWADw1
bq//v2cchVB2FQi8O59q8t6Ar7GDyJ/kCAvS+aatEqouzXtgYL0W2KkeHoWJWhkf
xuUv9sdoePKnPXrV/ZQh3pZgI6PBexVRNqkPLPZLyIEWVdEYH/Crlo6MRjywxxqk
AvlEtWqV+lzaM+R00vMW5VDg9PF2F6xiezTrQf+cV3Hm31nRfd5UUpsR8iF3e37E
hj92J3N2xRkg6vax47R3fcSvjzKaJkLeYtR7tGOBQdcksTyD+7/BQ4f7ljN/7UDf
wOIYX/tuhjghgoWJNOCKTl+fdi7HZni/3732g+7el8PBaDQ6vwNuSJ3kHaSmluvl
IEUapPdmognBMyvu/MV5/iUUAhZCwB3ibI5U7NsK9kHh7Gi7weieudTaOZaRwTqN
FYkA3v/8V0yAoV34BA02XFWQSnQHRT1J9UUzNXzrRUHmVHDuFdBsXtNiHxjUT+7h
k+seFIVy2g/50mqNSrvc4Nl6CwA3nNTZTk19lc9DCrm+lr0Sy0CjOxmz82wK7iu5
hWp/izXEJoOvHQFbMZz6GTUYuVeTlf++fIYE2A0YLOn4uD+kbFPPckh9/QVmciOO
7KPzPx9f7uY1G6wKeadOM74ZEPqGRdfspn0hA6+my3VZ4797g/NlAf4ValdA1WHu
erz0Ztz/EPSDD7b9khw/xJFFpGr16cCfN1Eu2hqNvQ2lvh5Nxqzjh2sNKh+Pm5fw
ynls4LdlgABiK6FsxGOZSu4K1B4KTHo1DByexuOdRm6ggqYbgnQP+4r2KozWax0H
9gKM1hVP6hGroAhEUbOCcYh5Rtsv2sGapWr8qRnGtJyWv6LxInp+L7T/kCq+7ENW
epBsLfBzQYW2Kddyd4xyZMnKYzVQV6vyXt7xjSi7jeHTk4aD3v6t7o9brVpQ2RfO
BQD2VWqj2gun0WGUCtqkoTcL5QM1JDSD02rM/BKkLm0QkOUnpoBVLJkgk9pm8XRQ
gfqOrgqsyXnsaEg9+z7S53J9HBzJ5QCC7aHK+/dEah46ICHmwuO5Ma8YxyGm6ihG
K+927hx6HKc2EC87cY0lmtfbOVpRg5VOxtCtNtbr65wf61cP9JbTRXMlKwZSr66v
d3TjLT1dZUfG0vQuZB6ldlKzAM52Dy7Qp73kG5Tiks+Y1oJocC9OfUx5yr24hom/
do4pybVjfWEOqHBuAKsUA2xP5fAji5EQ3UOneAW52CuZsjwjdh5l7iqv4iE+3SXH
NQqbqjbqt/7H1bJPXehEI5GIwpSiB9HlC+EwK647P+1VmHtiK6c1QkXSafidGgqY
gddm1VsqFz6QlvN/S7Nagbh1bbn12rMvrRh2eBItRLXijUbBJqohnPpd+geiPbp/
uybt8rV8GZp79Kzx5v/Qu1bHbJ8QC3DMLcJ9yRIhnw4dfKqkjxYTMkuX05taJnGg
5z6iY6AXoNHNYPXiSdXj3p6DkMI1XY56adhCyucWcLhgMHXBVBjLfedsdLpryIAp
BhoKGR3jo8l8HiwVcLg8D6w89dD0EP0gSRPn73YRQEW4FHTBhZXR6L4amriK9rbM
XqSlxhLPUMndTmOKJbfLgYUGWrYLV9pd6k3I+UtTQtoGWqeFpVDHChaIICz/egKb
XZTdzHagTkCChAOf7chDKna7P9ajf1WnSVm7m2NwL2rppyNeb0lfz8cPX77vfhBT
tIgRl4AsxzBzSF6Xx44jsuvFjghYz/RLVtfvUY+MhWcnV94AvaGPazz8EiNo2+SW
YUftFSnXbyU7p/zu1esszO6MmASLTecJMTAvZdbIBbLTnOL1PC6QwwmXk/pNFC5n
6+cCapUtIv1zmgcAAP0Exx0p/exiize6LvCa//CR1EyZGwvpC6jSrhMZarqm2bT/
BFmbPW/lPYcidcR+CEC5W5JcfQ9l2S8tkCBThOZ0sV9HcQ9XcSd8CAot/W7Bymmm
irjeAeBt+XkK706l73utSSBZoGA5AYPeDQ0J/dlHyObUlye9yfSSJG7C0GkXioOE
8X0BEW6N3GQLt4d17An3tVMXLWGTq/maocxLQZfcn3nVK+GdvkLXyTQJRnG+8SMJ
Yb7sGyMpaHlv6WeQfLs0GCV1pPmBiIg1TrzQvIN2zj4SGRoVMp/6+HnSlM2I1den
MZi3GUGKJVgxO3/+inxZB17FMFXTPQWUDgNOw/Gs3iMY8mjICX/AUtIg6ktlzDru
mM56MuOT4T5hOinAgGBJexuRtFe4aqkQgrrzwQrlnyzj5JRrP2rPr9ANQ8mUogAC
M9uWQYa6P7kHkpnPezax355N3HTFbdW75NyYFm4kegTa0VwLUYPx+bTGSjCi6zya
ieP3c01KzzCepnCZPbTRYu4lXG+7szJC002kRXnpoGabA8j1RSvyyzl3LUXVrPnl
KlusxbtIosdnT9Iya3AbFBzlStdA582wpPcvCu3Vqi6OubQzxJOKiDmwJfiCQbBS
wa+CAQnyah87sqZleA/A3mAeYa+cF+IZgDrroYwpR7Naqfb6dJLMPoFW03/YvuJY
4B1BsfdUMLDZCG9snC3Vi/qUpm8seVFRzVqnhEglCT1+3U1pc58SOSRtrgVu+dCj
tNj7bnN0XqOqpJdJGMH/dOeKDH/pFouyhudaOQmB9FmLWN7yhrnXCLexaICuaK+2
h0gHRT7FpY9mMrqy1P9z2LlPSEVGujDTNoBI7ttOVd3Y1zshx79PBHV0YTNuGR7W
JqWGQPoRHH7Rte/8nDoZLLaJ0H957sceQ5qo2Qm+OJK7e6mUUHTNwdkcz72Ppn3/
ymolEpZOYotOmlendcstFQgcLSMduW6X63DcvhY1w7t3AM602hD0cQ+oLRFBFKzM
aurLQj+b4n89Q6VmyWVcqNe1hKdF5m7fi7YnI8x+EsBag4B5d7B6us045vhh7sJg
rZYwXmTDNtD4sGpgv+mP2/8EJBv7kXq2HAqdL4/IyAVO0QeDMb9eBVUg4pVOiN4C
IEyysTWw7DE840xlXV/7l+TGX7kSdXYNfxHbxBP9/neW2ee6rAxqUV2V2Vr6d/rN
C+7ISlQsUSZZecjDvaeKXzxEVF4KAiRvhK0S63Oeo6QG7Ug5kf3GROYCD7H1yuNK
GwfuD4j3tw7lGuar+9AX+B4J7vPgXDm4WiiAff6s88ZOVF/P6OFhqLZZ3lNZj6yA
7xQ2BDalgxO/R0D0xiw1cbf2e9CGJOth2UfvudHNXDNNbCQH9zPw/y+jWjJ0MI0k
QUDBqnskf/rUohlf1SuQsSRJZ0J0e66hhlswjNnjUyHglI87mS9GNb2R40BKnTHo
REjbJY0gZ+7OO4f9H0C9I5d72Onb4RRGe36tLKRdhi8CkFao1C/euECwiIV1gXCG
h10Bhz+LdrH8sB0N+gyisC/xSzRq56LKuOjIrmwEFeBxx7eUxjVt08O06ZH1HGGQ
U+cJWHLCXzfDAioNGZvgbObr9Zkz1HoGlMVH+GXbWcO3spdVmUSxKOjog49bLONm
/yxVq0HySnHqada6dFnKXDXdy5dctKCJs3VXWnTkCIwGHcUPhWp6kKNtOWlxdgX+
qy9uL+++kREBdY4VOzie/V3vMzHd1eOYp3+obYdkxU/CeNxcbQfjnS6OhcZAPNfW
Nkx/9ka4LN399EmkTziMuZPezqesu6D/RAGAYqYtOpRm2y4Zr5n00U0ZFKlctXW3
1ZCa4eq31RHGKrEcsPAKfzt9uz5Eo1sUgbVj99LZnMrWtxt+N4KWF+H8qkwREPqf
dEPh8TCfezIqjgpLTfkzYRfdL1VI3rAD6NXdpIacNjw8YusZkHQ/CDFSUy1eELk3
YT2uN+OYIu1bgltjuphJwzKd0w130BaNNHu82MDc1REbjvMt8syVsKPaymbTvgT5
6cbqu9yWvTiAsAAVbmwnCUPy8xIToJvRANBs1MnhCDynQPxsTT8cHvlMPxJQiBib
d80Un/0GeSIDOhyNvVnepr4w2j4aUAl+RnObkB9RhYDpXJd3mc/IaKlyyCzY0DEp
w8+Ueq3RQRQXkfWsIhsn86U8gM/EL3aMMHz2sVWDQ+p8yNZoJVqGr1uEILYXxzEf
K0BL3uL+/p6bzh3/TAYvNO2O+X1RePOesNCpSHzmxxu6ti2/+oDVWeaFXPuQu7Hl
kBJw4kh0zhmIF9iWmMmBtD10G73dE3pyV3PpKOcFMq2/MWHIXfKcBJ5/pXz1UpXw
JJAraKN/Zg38d4/24UoUyMOOPSJ3hxwLx7Ekdqg+AiKvbOqt7gBw1VNGf2b31G2b
VR17k2mg8i0VD3LnVNQcY2Ty91eJGWEs91A4EGRFhYxdSY2YLt89j88iB6pxkARz
z9vPo/x6x2O2t89uULH097F7aGsplspCcuvIk0m9kRVLvgnWmtf4N4XMc3iwn7yx
bgLRn3hvifA85RFFF1SNbYjn62V5puVW4w392+O8lZ6mEF1lSPqvYl8hatdocxh0
aMdxCa35q5bX60VeZ/VIo3cSNYV2ZIUUjGPUK7Z4bLCVlk2HYqQj0WJmQUhlmWUG
mk5FFNbdM0JOU/EfMy5H4/nlkx5VLUHpuZbr9f17iYdN1THOeaGYiV7UrnSctyW3
IqRGvNLtV0y23Op7uOuJgTtIZHgS6kqI8ileZRJrMgUbHe9KcoM2pOVLMN7JF2As
0ETddjauEQFNDge4jJYL5gi6PVch207KnPbpwa/1sJNVYjYr/hbO/FtgNEm+TbeI
zCAud/r4TbEAlReMj7Omv5aF/bUjZG+YTcRPfT/+iIEn/lls8X/QdBvA4EzxAL/g
yjo6QxTBMBZhVTKMzi7r/9mJDGtsbwAsZeMTGAXPZKbwg+T3Afp0bFbDHvKhBDYC
XNtcdFBnQN9yb0zlR65xGMqE59eYCkS1oo7xL03NraaHtpZDarujhJQ7koeEwc4i
EEkQ75EFdXLdlCDVKJUs3OoBO7FZGAL3K97DZOu5KyFuz+kf9wZGPwTKC/dYAYF1
9Q8KoI+mDFds9E1UIcYmCoYJAEyekeJ316JdBJo7Ya1yW1dEOBnuK5jC+ETrh4ME
twD1EsuG7rOxmWOsidOvZ9X/h5dKlhKrp2HHHsbBoQZFJL7/iJobDFvqmLFNb3mS
tAX5dDMn/cMmRO1HHv9Akp4O6JvXzsADWgA0vcbId4rn9wF2IngQ2ufXYntZb2ob
AifXjVDx3qKh+ZDrUeFrfORTZAPowF3Ivo1eTVaIeElz3WLhtN50dVorPZpRtNrw
oTvf15BG/OyrX6yIK1k4i+/IBEBkzGpTNs3AnKvSYeiLnyl+8nlF44N/gWVXX7Yt
CmPKFq7bxtRf+sasMt+jMryzgc3vvRC9MpCOk2S5N91Ed86FUafZv+W7jLGf4QtO
5ehOD7E1P2VT0Vl2I/k8HnpeHutMZoDzKEyelv3x/8JloK2ZxYB0nL8Y8ajsUvN7
Qph3RC88CkMgTIyEXJF/jkjrlXgc9rTgLdoK1uvIsrjAXtxg4f+gekJ5pNth24G9
sB/QgcuenqayINEeNw9kG1Ni40n1im+9BpRW8vA3YCFnoF3i+KTCJ9MmVDlbeZ/l
dFgr/VETUvMLsNYM9tdKtaAAM6G3/FRxOMsMXY3lxRV/kaLXjPf4OnxF9Uc6ENgo
u7R95K/QDR3Nz6Sjbh6n9N0KWfeqvtvrHHnydiZfh+T7JV+fi/tXqLKFgF4sl8ir
3TVD3glLxpo0jZMAUh0si4syOf5A45Hh1C945ksb84Pp9R/iBSss9Qpk/5n6R44g
DJ0LDEy2GlXaAptVkduOP+qLpJjTl/eu1Pfn5hgmtmBreO+dBlhwwsCU66Ipofrm
SiX/DuO3mayT8TW6/OrA2TAjFDUreJACzaoXtRfvHKwY2xMov0PEPKg2iUXmOyXa
T4NrMKJJ82UYgqKq5DNyiKpUiR3v/KpdjBdTZNADOqYQYh+Sfy/l30fc5MvNwdCD
izjQuT2KVHJN31SCYwFtRllCjKVtsFIjuBN3yBGp6Y7ye7rBmq3jjh0EZ3JmivUs
Wsyjm4MlMJa01529jGXkyiEFGvtBDTJdjKZbAcmLjjWFR2urM52TMjteKS2GM8+o
0XCQgVhf9Y5stVcJZEEam6ajHETAkUupIA+loC3Xa15Ws1mCuPuksbnNO8vqnN/9
8ZdNFERM50RQ+AtHs/bEx8OMaZP07mIVSuDTq9lmQjt+stLnBbRbC4dv4sal1Tlf
cN5vyDZJmP5wu8D1IJOC/5DuT1vu7Hjl4elrM6aAMMyg2DNVY4VBcPbopwlNUKV+
g9V+coiKOcm6cWOoVm1X/F97hiYZKbPjbqyr3vY15ebe2FOFs9TsgcBKYO7kRLfo
vWKbN14WpIM65GT/S9TCUjm4/Psn3tobG+cLGnXyPMPLGGfN0rX6qmFUKRPLU9Xh
XL056HDnL7sJDzcIvTvTb+SdhlsT29aQyBevlpn5bwg5qzWv3ceYdFJIq/p1M6cW
K+Zf0xr3rlt2QuIaeZp8P4sx/Zdoh9DqssklB9qNwJWkP+96KqFWvPldVVz6YTQS
O33+60srntehYMlNLR19SrtbJhoe+Srz/0kT1kvjKo82qw4T5pCS/XYbb2FI/AoH
9gQClm19CLvB30cIbvDqhIh5d0/ALyRo+poQAXVzhC4z2RUZtEY+LPomtxN0LrsI
qsXoZtsCoDdojA7GeHkW9un85olP12P0BFUKAlIyAveHxViEe7dgELFKPtVHDX6g
BLjybpl+es/mS73v5KxNgVNvG+g/sEJShtxjsXzMwfcECMoTInOvu86YetvNQ6aK
Mnn3jcLrGWP8MtGeXO5t1QQSjYvBrt61zAknhf948vz59lFCyhtRMgz+VWI7ND8z
IPzmFFwCYkyiA3UylthoEw/j6TEJ/fe4AmHQs1Idd95LbzkFfX9zDyg2cBrpG8Gn
KsVyPqtdYGoxlWhSLz8e4D6oqnqA1GjjFRj8e76+8Cm4BWutzqdK3w+35CAF2XZJ
1qI4Gtb0ajY7OIv+hrCl9H6EVeb2fOOTR4Dn+NfBPSS14JnZztfgkv+gGFur5dEM
aB8dfxytrLXTv+HiVyq/ADCrmk4WPoFrn63PT7T1ipQ29DRJt4vqj1B2S9IbecU4
jIwHLfgx76MTfQ8RGOOfQaJtV6yJpmml5rOWip7hmOw++z+BMnDybr7pJIQ/4ZUj
oWXCKTPnqzP47VZwGHAqbN9RvDxTYd0069VJ9/BnfKja1nK4dQSWuLXzS1vucAK0
/Wj241ol5aMXlf3pHD3hgQ2/M+wd1C4Gnl/EDnwt1UJyPBNSSdE6l1hEupf22g24
sRzMqomJE8Yk03HDyuW52+mLDguo/Tg9FzRCw3QN0HCKRyAWMTM2pBPwfwStygNi
rJ7VEhuQc6jiPZTdaD5VRztpNqCPsh+2ukV99KwVt/1JoVa3MD+uPQoAKtkLI2ZP
uRhrkiMNNGTZiUuLWP8fe/RByCG71HAt1GdwhK7QbBz3Www9rCrT9uVOc1ibghgY
uRWNr7LdFCxUuCJaG7eHcyqwDSLPRfOTTyt633LUzoupJLDnRrfR+LCzgelOHBkB
XXSNp3NC1zpaVtA3FmzmKZTFvVRvjETO7aHVTZW5ZGSjIt0aikLYVjnY9+dL6KNx
fV7SrNlsVOJyaOVqTh5Rc7//fL4fqL2M647yYDuLia3VykLl82tgP25QB82G/Kr3
gUVsaUgoKvCJxqPVX46WbzQlFDwCQQ8TK57UL0IGCsSt/I8YFMgWu1FbUWVIZ2iA
kBwQbQQYVlOrQHeOTDEn35LgLyUi6o50HaJ09hR4MuyR8npMa+nX9fnpnU0ffvCm
g5NOq71faY2pCwHfhCeqXQFmqh6GTj+NqTxV+n8sIRb0WcJc9gGExbyymoU2Pfde
gGSOBCFwVMqpyIFG0nT72vg3FowC7yGoHwhlD222v5LoIOiP7adkwqCletrth05P
BEiFOd+49wvkvE+QRrm8UkfN7Z1Qg2VtHLF0XtsMXAL9UFkL/2AEwNtM9+YrxZDz
POOB3xaLMm5FSgY2K76jKuMNXqKOppezlOKIpqhfxe5Vo/fO4jdAd3R7tKfmed6K
MWqwCcAjEACQiq1wjaKPdRlY7OtsywjQQvtJurna4/Fxn/xoVz6nByAcsf1TEiXZ
+hvjGbBT2tUagtddIgxh58aM3s0OUx+/ZYhdGw6xivCR1GgKX5KpxMTYWDc0Vs6/
oEBpQi4jqGQm8GYBYK6Qf5qvVIc+vv82TomxZQwCPJDpAI39vv+gDsvCRElQHj7Q
/pLcGM0GSkldoML8hQ8a9GmhZ2lByhaOb8pWpCmPJGXXcB/9DUJUes82f+O+HTm2
uQT19uxgZWxkWxX/iWmV8dn91P4opDA2+2rF28EPPCxChzkxvh+jsiJExrOj6XOM
RMQZ2cdp9CggYHv9tkCPb8VP79LKO4htzMBbNmTv5Ap9jheLGWdWIIasa6w78++4
vun0Rm3Iffs2rvRjAak3m8n2y6JrbZ9BVwg145O1yAKoJl68waQRxzEVzhLPGGlg
0ss75Rbv6DMXgczyWbfjAyXodDaxHCA6ktj/04yM2WVbnEn49kWf5lrkGx5aDzQw
c5Nlcy+dbyA24ULOWuWXmAruQRJ2m7o5mFtO5lPYDfNJhxBTyMDHrUBo5GkdW7H7
JaEKTIFuOiA/X7yAqpksEQiBIrG7KDRnNgtMdURZSsC+MK67Rd+4o0I/cmuvmIFj
1kN3D6MqAwKQwLZFSpomxn+rUHdOW4ERzZC9EB7o2QMXumonXdkUb5cMPXUOco2k
esPH8qP66B8+osbEkg/p7Bpi/aF0PNFx6Y808tyEta+MW15RE4iA+mwpvJCeT+L1
lwp5Z13nE0lz8F9liucUYQTBh0+b3YBAb55RNbttUEA5hVAb0l8MhaudZY0CPW9d
QRYxrhGAEUEbOgzzzW4ax2dBzitMmeXqnpG5qA9oZpF1lS/wj88BXjNAlh66ztUw
4c5VUcia+gLrErJF1pFnqs6I0CqdhUbS0PnqFujbxyaEls3YvEDRCGy7Ne7bPHU3
heCuRQju1Msub8f4ND3zixe2b3AOoc99mQpTuF9MZus4TNV8iACKkbcnz4iD5Mc8
d790dJih0OHUr5QAv14esMzfaSfzPVaC98lZkyBUAIqj74H3ivA61XCbFiweGbrX
H2jslycWYCUoEGnlZNnOmEZWEvwOsQtmQ2rkEONhAgszsrvM09Cy82ho1iNNPTLc
G21QQrpilHJLScLh9E39liYOm9Rcqd0PykcYWGgz8dJG65bisY/aBt9QIgotknsB
XVbDCsjMKs4GbreA6if7yl9No8KK5SNcap8xXpribAlMfI7wCMCBglvN0TZW7YN8
+XPS37yJ0jHlgU/DPc3M6wUjlDeAROhTWlggB+3gt+9KXJ4wFyqrdLRb7wnZfns+
Xyx2lt14Fq8B80onR+e3Ya9uEQGp1oTqZAA6PDTObJVYjX1PRrpqc1/AT7uTiRfS
aNUk+jiz/z6XyqSp7kz/lZVlGcuFkEYZ3wPFwy4kJx7ZGPAH3ltjusrXGzChaMDa
q5yoTCttiz46ylDzlHtIvIndma8iiRMO5S1sB7Wigi0XLpVj6lQPuj6XkGlaWnM/
QacS7xcXAxIiT1AkZnShmDmqzmUyZ33Tlsy3X+oj9Aw1bcGHOxUb93y51FY9tTaS
H0dQLsrOzyr7b7JLABx9GmLDFMpvad91QyoMaqiAlMDi5ud/TDpeK7BeSnqNL4VP
OwCGD3IssQaYKvVhSQqYcT+JHBuOx5AHqi9WCHniBcWjjyQhpNbNsZ+in/vr65sa
NGSvMZwz1p3l6hkQ317SMcE6ccQoXWyoDxZKh+haNAYoak871iwBXlHpoIt5++Up
IaHsxEiT1d2DFyAJA+HOR7epYIDY1tpja+rjPMfEK7dqfDGV8d+G/++6lEPmTtze
PgHPwyOU9TFHETmWHNdDHBNULOB57Q3ITzA9RWGKLpNdLsekGKDlv29Wb9Td5g7i
nFxqB8b8zCIHJTfFgiULMfOAgbEE+s+7n3b0PstoAp6xZ0l+dWhWCKBZZVW9VnVv
Q6XIeafVyyZX/pN24pgR/K9cBZU78LOFpMHzzPio2S7dm8x2hZoIG4+QYEb29Imf
VJ6BhXlQ8ZuZeSHb94+UozJGA3OJdylC3v/+WAQ/tgfrvLkrYipsIrvx793K2Hkc
eK6FCwNqDTl45l8mqFfDs+DK/gEqR9umBgGvRhqilutAkD/Xrq+hsuu9zL07dqTr
1Ro/62MKq1dljmFy8FgN7U0hce7F73ctOSZK1K/MLNjJwvJh+OGCNx3ORbf2P3AQ
5c3iaA+YFu0Xe01APQbDGmK7VNP5r8RgIBBVVlNK62tEN16GDWNl1+nl8UH2sK6L
QzprwIuYK/BfFPkkzHLiuPPnPblk4/ntTjcAllav6f6tkuq1pImgk2CCrekED0ob
iY+8urjyld2raVLhULJxcCKtoDPdh8jR9ghbUeNwjdSNDu5+Vwa3UkJC9LsoYZLd
QAjdUFY2AT7Juq6Uajre/MlkcrhhabeVu1Zw/qQ0oYpIysV2U+1qserrjGaaaR46
GW3SuOE/RGVzf97TiJS7IjcQIHGn9kMN1kihci7oEuPRmdX1pJlJ+NgQKJrnMF3Q
poUVbY3N51BttkMlVOLoQYOcxkkfOPTK7WAhpNkcIqTnC8uijKExP3NZq43EpoF2
fWSquHBP1odY74UTKWTjVCuJWyU+8c2QKAVcEAQrK92fLW2DX4UvlXKUidhvCU80
nGah6RhKUv5At0bqmR/gTZTR+73elYb3s6Z3Y3TJnG9gbPOrEAewc6gZ/tsSe3uG
zRdcMkC1x1jBAHsxabRZorRz9Eu1OdDuOWqRq5xi+lR3oDPM9ABqZnYig7juB71j
ciqaqFj8PA4iWkwf96KlT7jTdl0YGPyIVGn09Sx1yKjHBE4T4uTQhQk+tNY0Q0QY
QiO+QhSsziW+GRxreRzspxTAtK3kptTRRgpJ2mxkn3xi3XfmiYDqkVYtD2w35iYR
zkK4LnOfBil3IXpQLQDhQ4wFuJJWr/Z+8ZpG47D33AvtuDsUoqtmD4Z7tmMYhasZ
N1HrcrU0HeapbJKhV6q4/uP5Ag8a7CIpcxofMmD8WxjJMZ0HhEu7WYWUJ8aRNBl1
5UEyHp3OCgSmA7OA8djiaG6as3SgQURoJXQyULKw/SSP7WwYH2/0rVPTrwi0lfQl
ZERUtu7/gCXWVwDnFSkBsI3SDeGzQL0aX5Be9IQRUEgs3Eb/eEz1rgwTvSwLPH/J
tIXeKplnAvT4J1ZYjI+1WcLT5fi0w42BnaARX2jwg9rZEpbovVrzjLhkN0Rr2WWH
xG//x/VnstGsBF+W3ED9l4+b3TVrqTxMSnAeo8ptkVHaSlpn+k1Hyc+nfOZPWCcI
gvlokhhtQYXZZhUbsIrmkxTWv7bQefft4QGfprZyhgqSKnh2WMCUJj6SaMWbE1uY
xrVHxjx6Yx5SrWRsErKsYG6GPnbSPc9Ww5/qKB7eQVLVrx1SzJ3qCH/Um5/od3zN
xSTXbSAAoCsbe8crVvs6sKTcy8/GJKR6cMIlkLEOgJfLpWlHbS+gEkqmurOJuRas
M+Sm5HsfeSK86uDnGonJbQDbGwX77LLGb1vZDuLeXlA65RF48MCmM9cvf3Z8Ra/R
Q1NnZnNCf/+4IJaeRXwvfpIS0KiwdZRAoetUXhDg8c21RdFBJv9mnJaIw6pHqSTU
N6AAWmHk3PKlMdcMHfMI1X8jKPyZke7MeO+sflQWVlf7Oi1oE4aZxFOp4YGWnRh0
cVIXo/da8LOyp7w5kqM3Yl8bGMTp1zKGh0y4KDdGPCWFlQUpPCCVDhCZsLBtka3I
MAIdoZFK5mMOk5w1divezmL4cbsJi/AsGyDYelmYZBJ1A3e98HMbc92InwUe4WBQ
x21NU1MleSZp3lEmX2NSCLnmEwld8CYOKZR7AZ5PK5H7LwNVutmX577ephfTWd7T
dtEckApkxSx+ita9rkYr5hplLkQp+0DAjhzL+8g9WuNoMsNAdGhqzXd1O7DxrNeR
mePdBRILmOSBE4IeTpUJMWJE2t01/7jTLhOO1SH47uQzJ6w0vur2E0wb5SaIikbj
uyaeAcUwGXGDR+46FYfv89b6oLEIxiUGcRTvyaiwz7QQ5bTb96S5x0qwsJZu3+Fi
dTqGlX058ZQuQLB+u1oZWloo7QJ9LOXsohbI2ZLuUFdj+U17FxQXXT1xUzBI8nWp
8tV9+23k1+C2NxsRNdc+2RbPqFPg/b42+Gl5LfgcLPRW9SZK3WtF2JhpoiU5Gifs
v6sd5aLmHg+aaXkIUs5FGNh1VeSSCLqu1bHOn5eYo2tOZMc3B+MSoP8vvg224JjG
dl3awjUJioxAmAcSFomO8THzokLfanoRZ5OE2zVihKbHjnT4H01unpYwA4ZduAKD
sJC/fg7Z05sIjWWPBtzDqA5xRd5jqFKiVsTyXxNSuOVVmDMkQHzgRTr9Z133cHDU
vdHKoPSiX1ajcSqr/TI0ibjbvvXiP+04tiiAyqnYjAF/UkYAumgYz0l6Mq6QMQVe
XAey8BQKWyDM/9WCq9CY6l9Vctnc/VQglZGvdvGHGdPPFtJSVVS/k0xI9X5MFSMb
HwoVyDgfRIWUsZSRYu5TiLhP6Fj5uvwkkIVMHW/5cDPTg11ypqWCSj2lY3uJKBNC
kdtDdODQnoALcH+d10ooOsbdlvtAitV+iXkxiCMJoLcZiGbsmhWvf/OYbpJJhenb
oV9DHqlyOaas14DXqAcrnKdrcifvZaF3clJkYEbEKGEZDmKYSypsSthkq7lLpY1J
w/Nu1Rg1kr9cdfilblLs/glWBBRQN+QKZNUQHpTivTP6W78RDZRUSkZAv4huTJp3
J8vBdqEurgq/fvMhzNlfCp5Mg22+U6OAae1f20XZ2thzG7kPxIa+sTT/ItFZgfUP
r6tsu8nd9KZxXIlGYYujDMFLevSWYt8jxv0ZT0Sg2QifPN2Fp0S5gwqEpR98UYBG
RsFlzwbqwVVlWA7/wmVqFYwB41qVMHfBeiE3sAlMkPN3eVEMSLTDwFzJQRAP6ICj
qwWq7nhfaHXWjKVT+OvyYV1cteoAvAb+GJyB1mPcVMx/i86WZfh1qSamY+jawsoV
zqJuzeXWHgLJPp92moLqjNxPvlDsebWSsjGouVfj75Tln/8iXWZT+UXOeTY576t/
p1/HYRt9kKRYsVvWHtRxXI4llOuDyBboRZuW9sSkXDzqsdzqBfPifHw5pAkjU2lQ
2kXEJU1WCbej7DQ0MGnI+U+iVs1r8dM87vb02bgnur6Ff8tKlTcoluI7XDS03Uns
UOQc6RU85ji8n+SXCzfjLpDPFKM9TZekBx07Jmlek6/gJ4JCvblrvJ6fcJy5Fz9Z
vqzfBntXaOWK58NxXJf1PN39HyqDxJiQ8tApy6iZzvArmWBPwFw+Oa8VeSCgAGvs
CWIXtCGAmQ/veyHi6vU4GlYfEFG8edZJapQF1EpF2jzEvAUWEXoBSgr0gUhTpsiW
JhX8NmnwxxYjqN025T5xmDSpfpfMLR4sF5fcNzB78/U2j6wBVrpL/aArcPTgt/4L
1biZWpYO4HC/UkhFn+JGAssxcbadYmImeKImVZg25dXn1ujV4KqguwHURtpONr4H
3PcHB4COM9P3+YnioQxavp19u6ssBAoCVD9ilm8/MRrmxTg8IqJDLPsYi+Mm73Ov
em79k7mwZHPyQy9fXZdeu7h8IGM2c7NHW1v3X4QUJzeGd45/AMLrTGyt258VuxrE
ZrcEeHsG09f+w7pamBmLbvl7yzHbFXyL3sWkW0hRLgKR/5w+LqMizhLU73wMYYok
HZ+tffAW4iLh3H6HoYzuY5gPQb1ueM1s3qU4Lmj1oit/aCiMqDIstD5o65j3x0n3
OA7PdmOR2zm0MvPqO5W303TQJG8zTRSTaiIawmJT+RYfIXnZNg6DBmQSHjTRreqh
wE2dAyOji9rNDMWZqKI74n1D7wEIi1bSk75o5S8esFiAjZN5QfCEVMwAjU3dUN06
x5KUK3gbxx/Sd2QEDue9rCNP0jMyEgc+JDTgYu2kW2Rcx/2qr49ZRKUs+q+3MzK+
nAFJ6qeUsR26yYXcc5H6UUWQOUJ3f/Ad/NfOwbC8Gln2AkChCzptDCdT4Fs1yGMt
4ynqlVmyUmyy0+wlSqQeIqudCGPwN6lyxCtl3yimNtbSIkzYGge5g2GoT1PW7Lj1
YCJaLT11RGLZHygOhGeThA9hl4+AZ3I5t3qOA7u94FAhnpQnoJ7bvt0l0aQz+G9c
pXkUyjrRwTy9abjmFr9S7ojVxA50KMC8ySAH96P6xDalRgmYQdRNVepaomsizmuD
ouBizoA1dCxVS27UewS++sqt1uj+5Pvb5CH4luI4Z5il8dVVSISnlDV33h48MRb9
8nZ44zzw1tu8lZKoDL1INS5JftbrOOFwZg+6CdPAwJ76+oLVNvEl1NX2wfa9RSJj
D9m3ufTIkCyQufnvaaciQejAyqqjtc2dvBcDEPxleY2LJoIS7hiw5YYAzX02ScrO
ROY+z1JAtE66cLHaoPpGbtI1wfQqxypFjE/ZDd9SFJFznpDmMgZH2EvBZLtr7Q3J
2miZND8wx/eE4aDxdAwcxk6uWmxQh86+eh9tvUNT9/DzSW8wNINXNKspCVC/3hJw
CXT9gKkdo2zGvMkvcs5rRG9yHx3l+GuVuJ9mUaRdQ2rvtX4HUjf59Zm+EA91z0X+
4OAU/7Ej0CAQ+QM8yBwI4RvFVjSFFleLpGrktMzK9D25lzUx5ryN3lAIVImKYCEi
Xs7yLt09zX8J1TEfA5E8KvM0kRJmY6XBagMqmGJbM3KJqiHojFLxLkcwJJPxxECd
H633ZlqYl7Wphnz0gqBbSQ2SHjusR9uwOz1e+NWluIpC2MrkwtpikKNcHqIGr1m1
G+ZyH7Inn+EiKRyjxbWbQl7sminndsH0eKvBbqRmkfT76PHiyf7sfIdWVShc4bSg
eLDnAcFoOtqwirRKy4qSJCdyRxB3rkIyBDO+/8Jlvbitir2uuBt6/KfpTvwsCHTT
FO/f5ASzRebgZhuPzq65aKYMyjtReOkLepclv9sB7YqPWk5UOh03SmwF/slIqO0g
lOzAeFjgdn4rbuv6IY1bWUiET8yBmov93SNFet+1NOLSzrLpBETj6ILjoSwyVV9y
NhA2fQyTPob2YHd7qhpkpvg3TaRk9+Uvu97A/qJhqgkPzmETDpIhcj3Mp9WGr9My
2RAYORa6qgU2Q53epqsmNa0luksmcaojNG+QShEl/v/md9Gn4Z9H3kjyvBE2yzA6
IvHBFh1JFyiFRBv8AB6JRixCrUGmfPtkcoZdfInhmP2xJ4dFRztRf1EPcQ9Lkpv7
XQexU+N0bEGhSgjGS/NbXJiTGArASjSTNrVsSiS3ZKHy4d65TV5RxjGcAEurTuiq
R/fa4peLAuwh70qtbqfDwd8nBIIE0F1P09kyv6+tzw2hf1qwMxcERUpfR+3+W8F0
xxb750dV8OMjtOgHk562Qy06NnQDHwisu02YYxkf/1MkeTuqSw1qHd5hahYZbJzU
JyCYlYX5+xOC8LEAd79Sfq+9LvT/uk51aHJGVQ6rP5TfszCKBZErrnMB5kKSUffu
UAgY7nI0zIPjrbmJtkAJZ1Lg5EzNeuhWrHEh9sTEq5M6IHMYB30Mtbc4Vel8qS8Q
C8ez/iwXKagHOrgTcytdQLq6rAKuY5CldaiiFlK2RhbOhjXchTPuGq0W5KE5e0Jl
YTfgvAlOqZmq/c8rk01xvSh+BjwnkoOWL+PJk/DeTg/WmOq+sgNoiOpnGETVWDAU
B0z39sarnyxmpXuM3v37bLQGXyjiVisN/56+BR/nupP/TSd5ajkoJsWU8f2/SYkb
cJw70dHhfPJtBnY0tufXODPe+lblUvdAH8Zko8pF3X3E8biYHndTLYpgJAGu8aUc
ic6gs6wCD0m6Rr05TYdyD6rovVWdvc1A9Wt3m7kObaQMxO68Beiywvok5asF9Wiw
lbaSIxbvbEWySVjTG75vOS0b+CHUiebMwMflPkPpk7cJr//QLKtIhJn8eiebnDwP
vCuHZUl4Uh+caw6ERXztaw9+Ky59c7LW4aCaUNff/aOqgGFtx6blLXd4HajQzept
haC1xSLdLxbKTE2e89YTUzzWf3nV/ocQNlrJnswvOStU261G95RXNv2RlzM7S4ru
QPPnV1hl21+NryCbY8+leK7tfzi27y75AIynCPw8WxmmgQHWzM172l5QPViCPwX1
ko4jIOe2wYq/Muemjl+vsIazNsGYzqAY/z7QqexMyrnSzm4Dk5KCIKLitr4CkoPH
wcW8gFHlL0Sbb8oQ/RxrGZdLEUev/GgmU7IvmduwT/fi7mNETye78kcHfLrKiV9G
gQV3e4ZV5wOe6Ft06FF2jmOdNmZUlgnFDqgS1Qb5LZo0mmaRttpfSVAhBx0yKldY
exAMu4jDtP6SM0Kiu7mlv3i5V5q+cBKpEXf/xrU7KVmlWMy0VUTVdM3o6lmm26g9
+ywme4CmC19IT1YYmRr0IZoRtSuwUqv9X7V76dFMep5zZRm2t6xfovOD6WQnvi5i
iE4PTD9a83KvagsaaG1AQJ1ahF1V7dQwNbidC7RZ2Q5vYxM3YtGODPO9KkY+F0gO
CTeAcfgeJIiyh2mMznBYCBXYo84awBZl/mrErca3O0ZVWuQKSZRLUZ7HlnK1lEQw
dav3OJSqGIhjOoZ1uhjPePO3D6mGqWkLVipPTLcRvfg+5RkXKFXKvdLuprtMIsLN
pgB8u5A2xm+5MkJm/WS/g/cGc2X2tckDdR/tjSQi27CcOTBh0YVVGGnIXyUSup6k
Kidt+BIFZoPfR8sgFTQFQ1lhuXHKQ+nHCeyfIcbASiTv9XIDL/9L07c0gOZuCv0c
8kEeNmnG+tMlD1SXDKOgxbC/2cg/m5AYycqBCA6gxMYvN9h2v0IVAht9cGnp/GnU
vbyt6MH2SVHCp6p5qFI0gtKclt8UIT2C9JXlD8JzFTqDDevcWqlQCpdElfqp8Auq
QLugt/ZY7Qh6B2GfXnkmS8dKZ1mpV3LohAqyt+B2QhCBD7hbFGISQ7Mu5+nE2d9b
bh1/Ba0e2aHaeRnu+HHdWV7zcQXKrGxpCE/l0iWR67clgplbWVbIP5Y7GC9jmypu
QznYGaTkgzpDOFh/j5SQ3JHjOYzC8nneh1FGmFc9cmHP7lKfRWaO7LRdT8O8ctvR
nErmM7ujt0/pDldRpljxl/Ly+kWNMO3yWSB8KLfEdnHRNuKb1NfIrcLSGLLt8blK
MUSdbRU6oKFmkKOQIKS1/7MqW9auCEC3Uk0dL+eYTAjiB/+854zF7OteFMAL/HmV
DIYoHZTD/XtPq8Qrf5n8TLzRhJH7OtY82NgTwwSgzI/1GeWmXniAC6qB8bd3eckg
TwQTNS1peFGloROSnvR/8hm3eVyIlROVgUchjDlZ9YXcK8MLdq8+4Vapf9fwDKAu
vb2BJ7K7Uvbsz9bSSu+jhK9VS5Kibm6LtxCUa4amLLV7McFrMDfJ1OM/r6V+CsOC
ujgEkanjPoHyax5PVipMy2h6NqBVcIZvK9qOOBrtBgHvLW0oUlabJuVXXnp1Uigy
cm4gPczOswBqvLDHvrGK+ZOjpsJKnfnZzclhq+5hRiXSheUmJyaE9v7YnHYMlWG/
2U86CJUyBIF7SfeyMa4Gm7IoH+6YAZPL56OKTG1FwLN/UQwgFFfyT9LiJlY75kXv
33hA18cA88eIrXL6mYQK/cdWAaO/Noq6ZT2Zqz731nHVshkxNW2wr21LJnhffmOo
AyHx54zNeLQzFw6YdP8WNUkIhekU1PAOUJcIwQyHuSdvS1izOXYqxELl8i5QFERc
Y1afYRZ4uYxhxpNWFFx4kIlKCfAVWTaqI1OTwCKpeae55bm6tBTINN8RJOICLIT3
eCIq7iZArRiLbXW62YKIeeUoSIhv1kAdHU0566pDj79M/76PjCAgxtW6CKhk1+H3
nHQmMb3vmV9djb0qcPKo8EOeVR4/+SEY3vkCm8CR4KC+Z4vaHTUuatjz7u7w6QmN
YdRn6U2bKTiDGEvBXERH6x7Fk1MrEMSzvjLLePpSk0oaptwD3jJtpQ0UFCr1Ii1D
Ri7KP+xEFoXi5MJgAZ/g8ozkilwZb3YOxRmwjiv8JoPmQg60X/9Jxujd5DQ7T6Ul
TWH2RglAs6eMJWw1xWHyzAtgMqRsV4IrP7VM7FRDe8rIcpA8p8pUQdZ3fDad6qSR
a6wQydmFPMaUv7wtzjgGV1tiE6cnhbx7aPr1qcYjZehcey9qaz9MuMXpQv7Lbh42
fQoV95gDpbWk9BmlWdlBUc9//FxB75YqtKgsjm/hADPKXtee/LoeSri00RLTIWwD
A9TMHgqHjT/1D9t2hTU5K3fkVSHF75CzJTr9q1kcAWbQb6SxV8vdVemKl+H50/q0
kM7Oy0IKBPqpHh7AlfSSqDKsYOis5vDobUNiv37Zsf89AyMouCH7T/US6UqT15mN
F3yWHnXg+L9BIpfX2XK/Uo/sPTvxvOVsl3J2qo712CQ40385nfNi41dEKxOlPV8J
KkwNF2DxzsImlaLA8FPHAPNTS3wBoIoJ9QbKuXbHeN+N7lgmUa2bkYZf824TLgYK
ICuGk4S1uN/zf6f/Gul/KgEzAjRL4dityLNwMixdk95Ze1xNpRwEB983hWFI1EPp
2i9yDDcFsE+K5E8YKAiZUSGicgA3MCsvBOA5oprqxXva9lix112vHPF23ac8ilhn
y9bUMOpWY37V7WA7hR7aFlRKsPjm4r4ZJa2oAzAqLdkgIOIt2t6qu9Henc3fDZUO
Qp0UszidrKpdGdhwL64GNQRLNMjSoIy9P22n8imCJPA2V8CrY3LI9l4/viQxSQ9y
yxBcpY1jJ654nt/gqqIAdct5/GOwkYQ/4RzE1NVmykOW5ezf8V5sFiJOls+36coz
nqI8iQlKNGgBTIu+ohXzMtirfRyOiUvHbI6yiUyfbtLergqDOQ92d26CqjXlN+6B
EcdmqGIXovSdk5RfrAt0V14g/xST6GvkWKJgt9x2UZ860ewtFvZnAyGfpJj75oix
gkj6evPwRy3ZP6e2fVcgUoxsv8/Wx9jBGmZLqy62L552z8ez1KeRUDHvQbNSot+Q
MTERNIxcFn8zqlCK0NfKtvFrniZIoCrPR6h3eBPFIP1jbYbppYnNsk+AfK0Bdscb
eL4Ibg8V00rpTKYP+S+89aL4dSyjNOFJAzFdF2dEcVFEZiPhRkKkpcV7rK1ia5fW
EoN/kb8zyQl2sS7a/60TH3SvOkUPE2psSMZJqGwPLaa5e/p7R6kQpY43HaQn0BGu
4nFRSV7HtVEFo8BhuntHKvVAlvta2SxRxzz8GKyK/TEKc/n2vCGmMVWRRlsZgkpa
9tuCL/yLhTalCkHy2qgg0saZxY1CfqI/yBzRXXBORGidnTuBvOqxhH8FA0vN83Oh
ZNjvtYqDaitPQ2sJu4Bo5dH8jUsdUtJnEBGKPZI92OwxeSLXDGXxDnRLWTz911JJ
aVobpnCqGb3feHBGOE5yDsxaQl5KYbYblBdT3/RVIkX8yULIWFhBXnXjb5ydOX/8
zDexw0FpScYhvDqJBuMvMf8eGbjuPZQgk+5o80A3GMbgWoBqha+DPQqdA3rpV6e3
PdbvYw1ZC04OSx03pu+VgvqDDy3lqsvtra5JAsQain552jBmW9Jl35JjBUf2AaKV
TMbRPoVoS2AUrwnZB0GuyFV0giFwjbamzP2Un39DWAgeUVlNp3lSV6SXhS5vtL2N
3JNLDp+Yf/Yhy2Dn+JI8fOVp0W0l5l4E5DmOCR9XrwqXsb5YChhbruy1YfC+JoNV
UsNqQ4BVR9KNMxDc89pxQpJb6XIp2bfm5ZTAxR+URznIwZmzKmDz1eQxGHcZrNGq
X/saNckxNiZr3cb0eOXKx61WhJJsrbWAz1DVT3nDe+XgTSlh5mUCLKX1+P7Jz6tV
Z8qa03qlDGwBbRWopiF750Ffnei5fkWy8Rx663v0lcIqB6Ik5I1wE7f6zHYouVLI
2r9usK9S+Y5ymqs07qGO9XSpoTqvxuCUAlRpQpuSDk1qlIY5E4wkjkZrCVwVizkC
9l5MmeUBhJdzddXuWR2aEpsE0XRGBrYm+k9SULmyNLMJ27mgJMHDjiuEMSvQnTGB
P/UfRTcQQoQ5fBJRd1GfMnTORDdJn2QFLkraeNrQsA80i0XQEvFHEbtwrXrOegPQ
w8UqIisRAd0F4ZYt4uXuI4/WBi7wHYrTt3QV6jen85GtBgFpWCi9W/UZqwh56Rah
Luo6kSYsjFOQnoY3ghAS2r+ot3+fCVUXbW5EaWQhfnf4Ci+UF+Um1pZsAAsUGakv
ND2+lNDW+eu8hahKj71LrOwheDPo8TVDWabD1r6qwYy5D//AGxs2ziVDUEzuN9RN
W0Xl3DPH2JGiRaaAdGnASnqwX8rjwhvk0pE1hmtWs8Etq+hdayM+JVucxtpZuG6N
o+PR2LtIGhvCdu/HuettI/nTgfic0IbF8YFRBRXMzhqbJhFt35RG5xe4hQiYJwZR
g+9/kz1pwRf3sK5lXVPfVb3LYlYjjNHZeC6AV9G1uT5PybMzHBcu8HAz3AVMau9H
uduAq+i9MHa2uhnfs4mReUJyN7ZyL/HDHx34vKuDzAwxJkKQ4/+upu8IK1OE7Vq8
L7HdnSZlpJ12KhIqOk0IITaTQKJHVz4vJ2dttLbqWpnwl7UxhTy1aWh/xj1I6eBa
niA38fI0ulC54J4q8fROVjnkELOJJIIl/TMmM6s+rxKyMXZfSYlWm5vVbblCmPug
k2M0cbObNjSFO98fuQjs+fFJbTBb7Q1z6fFDnZrC+vQypO9vZ+ilNBsuyb3g48lh
EFgjUrNTOAmZmp9+8mtXV+i1vCYH2kHPmxAB7XvBSvSdrjbCpJysaOxKSA66qZHB
R78xCSix63KkiFe5GTNthmE0qsAYJjyRi87Cw73wjuZmvOCkCVEnMNq0Top6j/C2
UXZt3KQ/AlOdq2HqKMVMlSi9xFaadm7gfZsrKOGZ9ZNRzbbcyfOTmhzxgpVnhXI+
a6NjlaQk8Q5urxIf/utqIRJcQhMnJHMUe7vMxIYR4ojBuHjjJnhbcAsIi0LPqXiT
3HMrtUBCnrvRrSfOvTC884spE8z0myARBginjlr7QYhFeQ3XTLgy2Kqxfg2G0MUI
FNcNCvWTipeYlUg6p+RXzn69OUZ+3yyLVRbkHF1A/isnIpA9sJ46jnR4/1rhTKHX
iGyZ+adC+MGXlBmHiRRPr650OTZ6vCrsWAbrXHYTfkTvWxhhPEMPDEsk+yXdZkFt
x9/n23DkOqEeGYj9TdGt/iNmBmCkJmag8UVTNzITaKpgRHN9D+MuHslmUkORSTK/
euQX0E2mtarXHcVGCR2uvTrOUjBtPnPjrmJPVqthXZ4k5jmn6mwTQfsn55Jei99i
6j8dkCRD46xVO/g2fwhqk/NrhdCratJzWTFO6qv1KHR1Euyt3CIYC3BC332HReju
EmgFFq5ljm40/zQKTrFxnmyI72OMNUmtpj6XOO6w8RUhJjhKHbd9RroSC+4o+yHm
VJN5Mcqaas906JvaBk5wKp1sB8gTkmsiTR7CztBkFPIJVfQq3V24VCfs1lvkxdgs
JhuqG4SPNzmrKfyFKYwUQzIod8cGCF2lrr7Omn3S6toDWwTUE9BIkujysa52MOZy
jMD/GEjs3b0np7PucRvLmGDwzsUyo8H3oHqX3ai+OwM/TRchqbMWrN8/TY7oa74/
x9NC2yaPWaFXpkZioT3Gv/fI6OOaFR2axF1HrHzKyjJ4/FSlK09y8BepfB3OGAGz
lhXQtJX2yKhweYBJF5nksE0bFnRpffAX2LEue/U/yzjIZ+zucsOuKLGi52EvfNX2
ysX68ZbXmeFzWfqquhTEhWho9ZlpCZdNBgjGAEIKSB+hMuEB2U1mPrIRfzeKzFi5
v+2oTkF0bXpfm8pe0tBQtEwzz1MXAhJHIZ2/vEgGU8+YmMc33Ym6V6AhUIaqTIgq
upk3rJFGr1ZnPgJKFx+G6gYfU+szmmTR9ZzAUfXAeWDl3JBIHp2fCG1Oqnx+kkQ2
gUG0QloGRsy9+kpNnJ/RbbL3D4tMD4SJloIiqjqV1xVxFoSvHku8YxF4FTQRNhNU
qsBwWTCvSN3p3JbqEMOhpuiM1PFneoO5Lu4Kc+sCeGp52XNX7kLACDIuA7PkMXrO
kTOKkDJFHG9c2Pl1nHi2NfKHoy0Un26ouLMd3OHYWfA10vmUbGludyVoD87ZRcCo
nMUKC+G6rAF9JpVDubYrMPYlqvQO3YXi2pvgLE5FaNA2QE3BqQ3qiCFCY68ydsHC
MCdoPIs8VDpRuExRzrXbMNRrMgtI0S0b7xQZ7EnrXCbS3HKmD226kSWSHZBjA4af
RLUz4eOa1OPxLxkU0ruNi0PCtZC6aqCeC2mVA+W5XV634Kt7FB1d/jgsC+fo1yoX
YZx8NG/NCKn3gZ8tkmtOsqwLgBGDpZXVPU64F28KEEXkfFqZZXqDwo01P7sNYL/D
cg6uWWoQJN9s9EKCwsahRajFQCi7WZ281587F6d0YWA6DfWZcdEdF4NYPoXNn+R7
TJChYbeUKXwxMZQqSYYISOvfIrmn6mMhh2VdYXvWq2dHc7fW+FApQ/JBpyKHkZ1h
rbXmPeC91uLGuS8CK91b6RpFHkb7VnJOX0CBQx3QQqLu8ftg8oQck4AazIUiZ78Q
gYeEzvGhmKLIr1vkIlEDb1eGqPslAW/LicGF4Uv9E3fnS3WFt1f/+nNaQeC0PuWv
0Vqr30jiIBXcl81by0GZv9o/jjF7Jbc5N9ucArTNtd2t5ntuKJ0cdCXJt2h2sdi4
JTXH9nwkRLDmsAtK2PCKxLT7qPhdPI22arZjQezt1OiFP0+yiCBI04E0kRZPx9qk
rCh6iqWU0GsG+tnevBItK0N6YzlEjFpVgHYkx8uSknzqq0+JPuOtRMe6hmqNLmP4
Wbe59Mk9qo4Ab6fov0ZLo9uHqYeg90d9kTjvmLY4/Ka/BGNJFStP7tmgveA2nFTD
VB1vUV7hR5xsIMwsKE9nnSAJWuB1ZF8yb6UjNXDIwG/XuU7TDwhFI0oD/HRw4HO2
IUhHxAxx5pwjnsuGkvn/y6GhnBGZiLagZkm37upC8X4/z5WLzaauFr3/u+Os4ctL
pPH2qqO4ddelXv7YF7UHv8V1V5DqxWtFv1SYBZa8RmRptvNTefLw7zAsCYbdnuyH
7JSn7MHHpql07UkP0OsOyETevWxVLXuCsNgWv58lDSZW5zydWmJfmadma/YYrTVj
xrXPhW4tVx2pPoXgumSGAnsdPrtnZrJ9CppA0Lsoe37nQmHroxNr+I8SEqiR4JKP
2v7BQwb3kK+s6PK4+IhyLTLWdrgjy+NAx87pW0BsoMOoWzgPF4MuODol9iJWGSkk
go6F0FmIQcwZ5lHvzSCq3kNluHup7NHRbEOPC+V/s+Ie7yiuBz58XoGpamROZYdU
TWiIlE1xdZEEyb2yEdXbXMY8805Jt5g5AWJx+QRei4vMtFYV+3V/yJrDBW+tYFly
Lc0d0QxbLqYtSfr3Z9TpKA5VvGqavg4ZcRYGtPrHwUL5kmLpYtkhurKiEAiPRFe2
F3HeeHGKXl0fdjTS5dsW2ojxltepKC3FNspEvGOfgoy89Vpej1BBXgk2LQbzbuRW
U8Rv64e1Flu+uvbs7ZTcYm8mQxVuWV8ByAiyJlxHdcyF1HJX9aDHV7iUScY1iB8C
cOS2nwM4JQHeFaMgR53uqrc5n5lfrsayfJb+q0bezdMA834AalLZW31QBLb7365o
EyIb/CUqkh0Q44pD7JQ+YuS5qxoL9a6tNuscy0IuzBgzacCo90qrwtJzYrRGVDWx
Pe5ZF7VsZz5BxUdy+tTgGD9jBefGnN9P3Q83lzjtP2MhJR1z3lzVr1120xdJjEFZ
U4ipmN7OXvIg5/z5xLxriU/TT7aDUfjzVXyO3NLwPWzBlMF2xUmrVNAq0a+jBFeY
cdvqIGmX/q6DhXQTsRO2EB3Og03RfDLyLg0Wq942e7vvmYY1mRgfcFX1lPDMzLQW
q2zE4s8KnMnzOMNlpi2eN1EpTK0ycjIxLTvppLV8l21kOmvoitr4A+Lt1yGCeead
nuiwi1xMvGX+peRTYO46BZ3ih/7KW5w2A0XyAcBtjECZJaGVSHXq0oPzMAWiJ8/w
rGOPz7XJ+RtY094m1temwdxXvj9Hn8SfoC7kyleOoQsu5mz9ClSSHheOBUSvtfE4
UfmnJHWH6Z5oJHKMmK/NKvaqbH49xMzFRGHhHuSCXwFgHGAjaMVOfE0yGmKerKuc
L2F2mgG+bkfkFaR9TFCcFTETT3bo0AlDDRsZQFFKAJpTrgG5EUuVDMFCfwtN09XD
BKsM9NqEneWvjBhMMWdB3/1JnauV+djq3CtHFY+M2sY4JaV2vW6W0q+MXJrV9Nl2
yWVfSoRopNTk5xdNDdqxPCeXM4EjzylABKN3oSzb+pYsqykQnGE89gt70s5oWUDV
MuW9MW0GC2+2cAahQ5rc9i6JuTgoImlwM10K9lJzjozjBCznsn2y8z6jA0RofNs3
FK6/mIkC1XI7Sv5Mrs8BU7BsTehYgQHO2UqwO5Lvf+z9QTwv58NlYPYqilRnIOUV
31HtSmE1yrBRiHrFiL3Cx5HZDyRfn50xJHzSQn11M2NDr34IFc2E+4qsID8W4fTy
XGK9jnNmaH0bzZVoRD8u3T+KlAargD3RrWtUlgK7YrVtBaofXlWlKdfowjbM2oQ4
ouUKTq9oHEex5flJFmw+vhDciqx18A19rftDxLMM0O0kdaBBU79knBK6YNl8/gdP
yYZYyLL0aKkrr3QNMpqlyZRvt7pSe7guPrc3kx5K+K8bpgG9tYQrlel/TiAiTKsg
OdbJooItPo768eGvDbJzUd32aUH2Yu+9DCaDcLC48NqnAyyaYYX9rcjMTWjjVgMo
Q9cWRtJi/9L1Eq4MXLXKvdAT20ex0hyoDw783H0YND3TWlfqpLNjvmJeHaOG+t5O
e42qCZV0iPxP5RPmeVWLaQc0q7dkxdduUVa1ggrFA8WegWfHGs70WRsiIf7OHGQq
csE1J5P67WWdnFDScbbGN9QyrxQe1lBH4gIk/bbf+GGIU897AHnMIJJaTHGPTDu7
cSA6adRJuHR34tLDD7grsIalRtJiPyWuFpKByR1Mnvg2wpidx3+4XpbFNCq1Ot+L
BrS8tjWTaCrcWDZwAGqRV7wCc3u8QccTJbJ1TCklJEMvtExfjy9LmmeirETmpWL9
8NB4SKNTV/aFlfy38bAN+EcHb9dD6kwFfAJa73aW3YXde6ectfrRYcX2QyrCtuKp
YVUkQOj1n4N3UE2i9gGuWY+uVkvxmnViebzHS5M4e3XDAap/yLkxvi0fViuAlLEL
Wjd/lLCQysWp2vsmHXQpOQtvHEYhr7oLFfig5QlpzaKs0IbdlAVskOHdgzqVqtpv
SbsiOdIsASmGKirFAoJJ4ne6fIfH0sXkq2xCpmICyT47ZemcOrY6+A5GVSuhVo2L
PYd+bRKh3FJvPCdj/ZZeIBQjKt6i1aXWWR35dh6/IKBbDWxyqEk55DNsytJau4Cm
H/et9sIuuYfTuNUY84rj3M8Sag1P/Gh2g3SthFFBR0HvQ13p3A5I9yAQENcGdyRs
AG+4z2G0MRc1lyI0W/nrnvBwpzOomIZVwP8riVlwrOSo6JHri5huYutXfMTTb79L
9n8ZXsqxxTV+w1At++TJpGCioSZz+6XcYiuXhHMyG2xUsU2I+tvMZ3gZnS8WqOJ0
qIaSA0WaP92STWxaI/nZvUJGNWqSBwT5LUL8W/97DkcaIF1ra0UsKlTuhP4cu7IS
kvn3XldEbirAkLfSNSHDtTrg6kYeRz8t5ZjZDyQ3FLk4JB74VEOpDIRBNL/v/nCM
7fWzy4gwoacVnQx5lTESwXBkrXwSeLCAcfmQx7vn3opqUpsHTEWW7gs1niRZQx+0
5urC53TG9Cgo+hZNHrB0Bf4tN/7Jo45M7Ajuiy3qZPxBTvZzLR7L9Wig5/u/wdg9
ZKnlJSyCi449ylzK5RFKXpwOADlTMfnAhz6h3vBzEDkF/lPwDxh/x69n69hWddwB
HkU6QlPNNyIuYOKYJALgI5l0Ep3feIq+5DmV0RgOrZLJCNpnPXBUBwXF+s4sYquS
NHrDqW7XaJpKYaYDCH1ak8yq+ok0jIEzUBjRqwg49MtEvfeqWtOX9MgkFyRNv0lR
qHmfvkGuQno9quFxi8QVdnG/ve1mOV1MDUFCkYH9TTJdQCjAXcs/3Fj+NyS2/HTE
hjdRzLgE8VVthu3l80s8D3w+roFC2s6fJpRqWnAk90ZpRIMJ6maBujL5UeTf/1bi
Qwhm0x+a9XNJDDToM/CsTySYvXW/jhDxnUaYmiRAf6JrO2+SRk7TIg+9X8XX25Fu
7FnB/w4QuE+1jgAMTPEfR3EvTYoH9yOm3lkjIQC8aruq6TJ4xs4K9nEyVnSl6313
76As4O8NBT+1PjHu/+sUzNYoGPJdgsX4Ay9L0NeLS+a50C3/ltrALVEYhJCSer9V
+KwRU48gqIHbeLKI7EXQ6B7yMRmEZ/xOuqsuFqM9v/7H2HCPjRIhLppcGe6PBS0Z
gGSfrfvmxaYy1/QqML0t1LGJtmD+5Cy0UCmenDuoN9YJQMtDByllR9tVz19nr1uE
NPclUBHwtJzeM2PZa6qlCPzbhKyy07CYU+cpumgOUgqh5bJRRHyLK86ukliYA9rF
nIqZuyMfeex00R/V6h/4BmTTCA7cjwX2utHfCXEBT07fMVf5PrmRE9qthS4HwdY5
c8WvyfwTq03JqjAFzkBm0AnFVCRlwCOvJsl1CNv6d5ygvPecGhBPUM2qurRkYvH5
r7/3YRJ8Zmau8rDJEEBBdJvAduY4CII3jCbFK2NYXXeLkXfMDa48a2pE/7dv5ZGc
Sjaa45gbBSuaxdViwN1zKLJ9+dhFpi84sfYpSVB9Eu87t7fdvJerw6hQDv0UC7/C
aRFS2KKfjsxW9XYERlV/m7zj+jGCqDfCN8LqYnuMtL/sGQDcanE+wLy7WhwBvg87
plKrhBY8kHheOCZruxhFnFfEkW+Xy9iC5ev3ue/+mdSPYE+JJI/FDoyHq+3IFpxH
D1/v2Go2/FLvN6aRstM42gjnlc/yJa6iDAaZozshtbgNsDcRk/y+1kS4DpRPuqha
xZ8wjb7ObQStx8TBNuyC7DLlRrchQIcqtNX2SrsmIQ9Uo9o0gqFzYUPKY55DD2gW
sWXn47emJHS+vFUxreU49eYegKE8RYDNNy+lTGzZkJq8xmCmaJoJLB439vfV6MnZ
8R2OMiA5m8iIpOg2ZUL84Vi1K2iPtAH3RzGg2H0glPjPWc3thhMTq/jbOpLvgBuX
I3bE1N6NwS/UIXPuoWni92Ol4tLLcTJnh8SA8Qbygwma3Oj+RNlQf+nsfV+RzsPe
vdd4TlKwEskcuDr7OIdGDhJZzlqMiKnZmGAIItnr1mPot6sG4wYuEQ42Uq0LUC22
1KJrWynUvVRtQaE/mTVCt61wPHE4ERmxVR14kz+3BmhpjxCy+5qfXNq33VBOSaHc
Jzx9o8OcUtPK+KDXI2/nim8/HQEX8NVoZ9GA/RTDNl3D6SFQKa0akJtn7X7Q+lLJ
hhlHfAgZPXwdkSLos6KZoKjJQ9Vg53CdYf+QiF3eu+dGii53Rd3OyyFqECbkyNtE
aeGE8M0N9wjuBXBoBR3/kSCrSpLhR/SenPDqKPa5SFTprDLGPSA3TZC9t+3P0WpT
byi4VgXFvH/882WIUgaWCRdRk2MfKkueRizZZJhOuGmS8G/Mpyr+SXG2yjnbwO9A
LxKq5yTYrB1uPxmzYBGeJzkbE98cMdVF+YnUDC4+fanYjsYjC6UHwG+bXTRsgs9B
MPH84iAPvnp2r/kabUD/gK01f2hzsPi5slWCnRZwoyOE9dgN9BAKU2ggJF3susl0
RSUKTlU+2PgbPHw1oXrPaI0No8bxuQ0KcTStVyl/aLPQMASimmMk4TIiq5aWRhyB
QZ3xushG15xx9K0o97ZUJyXcbk4JFdFDoFCVuEeC954morJFwMgPYPpY4nKtKjM1
OzIxfDraxArGhru7swGcWupkMClsHQ8N/GkHoWGSt9Hay/nFCBsPS0Cnn+19wk1I
NuK/HOeaLAa0llb1IuQKI4r6e3ryFmfSQ/dA/7UxtaAqPKzSswFvprz6hgj9XhU5
wiGlHjjumyO1hdyHQEI9y5M6FNt9uCeJjQiBiPJeakyv2qJ9M+BR5GnS6pbRgMGh
dg2GcbYfP/WaUe82E2nD9YjiSmw4W7o2qyCqkajDWkMeLHrKP1p892vjpnt+fjN4
7r1mWphzxOET0CmvNztCd2y4jiwMWoQUcM9/Q0ic2eNOVKhaciWxlqUEjkLcwowc
/onTFLj68/2Pn6pnctnzge69hWZsqEB1e1fAI/Yi4AoCrZ2QAG/JGKyXh//5gsts
DCI9o3M76MMeC3+hzY89dFbyAQd7c6eMOnfAkJEFol90ZOywhFU1YFT9jlJ97LMG
FvYG9xzebmM9htyxHozNm1puGBnF4TumgzWQiHKvFTzR1uZN2GEw/gPd9bjgdflk
eoKjwVpKy84XfjK4Z75Pmodo87bbKhJMVDtraz5EnBzEP7V/Z6VvvJtBldWV6OUb
q8m0Qlz6ji7MUvzWjvAYeqrmKtTUoFg3RHd0KMHJOChLTL2r5NpTl5/gsxS047nF
gNocoasNHMzYEncUs1dzDM0jbEIGs5IvqSigym9CzjEW0s/gW4H6BCMljumSuhtJ
MMKWFbNf0FKXMvxKzyyhJBpOpnkpqZZRX5JvHbEihSsKUyeijzYBLGLh49nlliwI
UFGekmlP21VsbiSeaignvGRrkwNBXDO3lykbROeurBc6VjC3zZG9NLMaKjBj8VaR
9DP+J73tCFA4qQpGbX5IpXvAObTFNqGG7OtYiTVL1yB+PtFgIfga6HQD7P2/q3VQ
5o3I7TegBDXfk0KdQN5jSx7E9WRqH57bMEHLQcjG6YY8GGGKH/z3uGFaZVGyhKb0
UQbj2lL7Iky6V7kx4yPtZ5wrWrNtTIYxlXB+ExBI4wN3rMPNfDvX6BpUq7sf+i/s
EzmqofkfaevTpIyoJJBEXMysJde3j3ljMFyXSNnj1ad6/lU13wqZqRljcejyXyXx
eI4JlwroJ567n5QR098tpHFyqMMEiXLhoDJ7tytonwHwD3ITq1fFmYwj6uQX5jDY
Awk4gRNnwxBZkw2lPiw7n70veCz9rYuw6MpxnGEHjEUqacI1z+aMA0rOqPX3Eg04
w8s8JvwLnf7JWqqj18Ol+J99Oa9vdbUDuR6S0NdFSejtfmKzIRnbHFooTf0lywXT
RxGZIEYnQ6xNdpTwHmHAImMv6Y/6tF4ta2jTrl6tKz8GUeSByLZ8m/SfEMqLCm/C
w+u3ReR2g04rbZv4GFCViZnOPeIEbNuMQVWYdPQSVWY7VOGvPaTbxOHWOCpLfZ46
k08OdzlymhEWIbErLVLKWkQeFuqy+s01aIKIyxsNlsmJdckNdQHp4PuXd8A87ukE
5z2GGEoFGhcT/DZGBJAf4JqYSwPviTmEbTOmV64cpMglehJLWQDgFomunJZgmABw
Qmei/242hMj3hclE0Imp9NS92YcQPWATDggD4u4kZcf3ZIxyHA7uKGTB2+z5xtrS
Fbg+IKacFRVNi0naux9XJH8G+VQeiM2AVhyxpJapw/w6Msr8TExXSnz2SNkZ9/54
lZekX5b41PrNeFgFJh+L1QNyGoq2o+7/TORLjgwhy2iupIGeBPAnkwYMaxh0zo+i
5fJAFIbFS4wzBH9ZHEeh3ZdjfCFax7KxHTO7aQDIdAdr6yNHqSJSy146MUZjD0no
OWpSu51WKps5jBYScYKmYcRJmys4mJT8XYORxfEXO51ydtyLxlYCRhFMZM7+Chi9
ZRg/OBaLu1tt3ox2fi9uReBqIFRzottnimJhrlvlVup4jxDecg1OEzBI4g7QU427
6+e1kn6HLw6JNLo4+iIYi8RG+kmRUpTCx7KRfUd5BKycPj5YSeAJjl0w9zhzVH5L
Lwxiezu04zso42iQj1mnV9vT8ihv4Y0sBAlw+HEg/Udq6SdCfqMSaMc1DRu9WZ32
97ocsfRFoAuN2WSQ//ueRM9mKoZYsDjskBTFxWx+Zl/coQr6gj5LPKdAxBeVYuUx
zmjn7IUzHS9u9WgiP2seWxPRd38h6HJ/g1V7TGy/eVuoxTkucw7bXzgQe7Gc+S00
ZDeIvqFcTFasP5+tc3clFlMjAas54PPbfAN7VhKLh+Ljdx0jZdh5PQ4Sm1Ineqhl
D2TU9ZX9Vdz17j2DAd04FesXUSbO70/l9sXWmoNI/i9lhDsLRy/JYb71BEm355cf
6cYbhHWcTOq1mAFwF7ZP2a+nEwS/dq29w83/sjJxZyQxSOkqDYwRH+rNAsrWojh5
rvrkMnFpzEq9ox5ro2k0euUxOIDQrYLO4CGZVEBvd8KqmAdVeF8Xq+dTwiybv8wi
ReSGOxnzUNrgYd1QrlqnFPk8QXVkwguQuO/gDXdPRtky4uwPr63+fc4mcdz2/fHP
hVktRHjsOqPdxnAgUDXhK5uzlN86Iocq8rzxKEuLNqVMIBQLQZA5IAN03KISbzvP
sXb39K0pnsqFOSbQ+hV2ZimgovgHmyEQn9gMmFwNbbD+FZpXUaeB2wcK8w8byj9U
/LJQGiCb8kdf5b8/UwTpfz9DuaVXx8nrqeGUHH2UxtkVWkCOYhm1N78GpgoMtrNh
cE0lyBf8HikaDpvBohK2RKI3vITWUsLgI7SvIFXM8EFuv/TEb1H3HYK+rJNI2EjX
nR7XmrYMyS86VRlcFKXzjUTbJF9nzD4jx7jEGgmEU59SSP5jb7IHB+OM1taOInU5
Gy05kfD2v4tmd4pc1Bw96Xmp9n0NleLneRoqLeiNO4e9swV95d7umN9/ixhEl7/5
fNUDGxwetzKR0EC5Sch2d2ONwvhgGyB0AnwFjmJ1NiLBtWVv8k60SbyzwDTfLtn/
V5dNUO7M4ZRBnFEvVJczxnuw8HCAyojhBdw8NS2go/Ja92vUPCE/I2voESA8aJon
DXruOROObHMY7rqWWtOopJkp46YXyLFQYeg/yrHE1CvWqrnT6Ju1Qkk1bW3Gf3ir
Fm4SKSjzxePoNVeH7Ep1xajQDdDLpJX7qtoLIjR9MTagi6tgUIGhqcIErqDM80gl
efeKjqzJwxia947c6zbSJgaKPBEeRZ6epnFLT9uhMgwMFMYvMT59tZG0FD9h6nxs
bYWtAa8txnRyKQzTSU0rnH2lf42x83ranNFNXefpk8OZBf5u6xvFfcwA9Twvz9d2
CLbMvuLXdXXHwoo6+QKU2CkMlJRCMwlWFXMo7FzZi51b71ka5Mp2PWevkHnDtWtI
O4wN1C49/7ExJv/+h4mpqJbsFRn5OF02hhB5Pb7gQKtzlD/fnvtYKKGrtBei+VRX
IZmNDC8VwVKI/1I0Go9pXAz95GXYiPCggH0rZyeJ+BjPKP1frU7SG9PnqSqBjKBD
Hw4pgrQhbaS9Sz4hAu2W9IvX7hRT28HFWo872pr/3oAHTCRAZm/Smq16oJGhQvm+
kGJ9QKXbskycz9jYqsgykgzbHMPCeAJxvfx/RC+ipvHOcrjxMPWnATTFE4wG/NYu
xjxHfRAaOQ6jlX+YCKIet1b04SEhNgfmDFPYQupgrN9h11ut6ulu17XRct6hpvAb
+x5/dBBi3Bca2Gqs+KEPb+GfEm0YHfWR1QR2ZIMTAEDgPYdxRJgv1HhxHO9p+LSq
rOodZK33XgNacTc3GvVPCR3BqbIxR5tdOQ4QOid5z0HXDLzlC/hrShtcQH7dTlMT
CeB7lauvjU3mxWbvMJMLLjokwfPHAOg/990cfrN42Q+kzOCTKgw9hNmfS0JTcaq4
1QMZV2ou23B9XXBHIYZ9dixRQRsnppVFkpN7wVPdLyNUUXZeM8pbIPWvNxN5X9R/
Af02HcqI/yUkSwE9eT8MZbJXJJYIfU3jYZ0dSnd2CQYP6cYbIuO303Ctbbx3txog
ZEG19sbSBdgSyk41xd7q2b23RohIieLulLbWV4t/hHdkwVQTgg/9w5ygQjJvQhRN
DyqItnqrWTOTzc8WBYEYT4W/mFpGXnfgOLLCm07rridHlEM33tkUSt62zde59Bf/
Y4Pk6AzsNNo5ulnWVkbCoMIiwBsfxfcT4p5LlPl/K85SH7A/BMa1qwDFFY3i0NQw
rvoWOy7WOT/WuZyMAT622988NpTfa9EmAqx8hiR5nOfRM/420FXK2ULjGWLs9Cz4
9pMPS1WfOEDLRq+YXqjympywrMoMS/TmgLZ4s8stqKVFC3sV9DDlrdIVBwbfJRKI
FsdRII/WtWgzu8VkhDhpzCS6Fs6geIK2WEuklKJE4EJ7jW5rvm36lck2op/USHKe
zNBcLTO6+ZbXaxPYHLZcGSFMwYwzGYCEDWJslh8DFDSqZ5Cpb1kn0YPUVbcyLM9f
728hY0t5dA9oGBJLFjwpzchnwob63rcWIXV/H7SsaLiK3WxzNql7mA1cYSENxUSj
61ou/1hrenz+pEThUJKnivasN9TiNU9/OGOvSfi3SLPzGKJYVC0onxVlTV1If/Bs
d9V0fbHnW3qgwEO6hFllHi3wYYM/yB2opEwdY78W6vcoNjBAK5yRqC+Yx5o0UEiL
2jAvr2bCkNYfYxuZXfhVFlHVHqKeoKnrhg713sv/O9ev0O1iRNuzjmXGxCzS4a4U
Jb+hx4ps5BKNwZ3uiDkbLhLdqEf9khowmLD8zGQ34mEAJQGoEDvnUXUbDh7mDAEs
M3o6tP0ZJUrxGXW3m5gXWvb2xi0/Sarp/SfxbcLkdjw9gnJVDJkgiXaqQyyMO0tW
gtJxmOWXUHucnBlbs6XrNP745b8kiE1IkMkReT9bVYLNyJHAuvbyPnL/dDo1b6do
gKkJWDeWAJ/+RPe9TXLzEysYziXlu/FaUYzefV9km1L4+kzsLZXG0v9ROtxL5g4a
LlKaw0fitHtcM25jZa4EUicJb0pSDFPH4HLg3dXP86jdgDnsqP7wz9l9Trp1KJWo
G5A6Y8afqdCRyKlTaWDgnjNiGzC+fno0hjaFOkr6Ix6+sTZ4Xej4nWdxnzB8amfi
YoaQCsFedw+qu4rGdOD4jvmGsMPr7q7crcYwKBvAQ+Ot7y0EczOldHboe/sHUl4/
n9yHf7S0R0/tYTpEaQEF48Lcm8HvUPRbGNRf9qPcjAzE8uEjj07MUPXEbJY4eD9+
e49RWZuStsgTYRL+kV0wYFmnyzBCplENQavRWSTKpNskRySymACiUA+Zk1z4mOI4
tdxdMpUeXxhEwYIpbBOmr1h/Mbss1RbT3ZVK5CYDCzJ7Vx0ccJhbvVjiG/W/a/+z
Ogp4StfzyQgQ8GjlgcT0wQW7b0Ww4EdlPEVlze49HEUl/gZcP/EGVl9erSpDDnIm
bl1WzF5JBBX6VIx1R2a1Bz05tiLbjDQ9I6KJqkhVQhfV/MZBDsQ0QW9VUtS0sNF/
B99KX56kf+ZmqMiGQMCfH+T5z+fw+QIpEKVL2yZO0Pg3Z63pFhMg5cGSLkd6jJFH
0+B5dnhV/LtZjmIJsQ7Y9kJ9l75quLVLvBibqAnJ/IRV2QiUMPTjBbWkmgTXOoE9
WeTeds4B/Ky2Cc4gyn7FZbhCaLwGKvfubzC7LMpdiKf0VF0MaeNyHU+NTiINF3LB
1isQCNFeYRN47m6kHIy6OPu0P+Xsza4ULBnV2rvTVcFtZ7vxghINEL0EOGFpBYOl
4SjywdQudfxjvHHBYe+KfWKiUvnRvCwgxIMfC+eEBRNJ9o+dHCIJbaiDthgyxHlm
o2mj79EZOshg9wK70DvFoOw0Yw1k+EgPkbL9ow1qtzyFgOyjG9E7lXLbOCMnVhA/
AkzrQdNNszNvWzogWCFEImmkrvh41jJVJGpFkGHuZIXZomreYPv20bC8/w0D8fIK
zgXD8Se+SnnS8ZVxUVQAGW2eqR1tJLEJPjxGXIzdwR+bA8ts3VfN8gg7y0bZYZpC
n6Or4GIZmkr9Aqe5xIzAg9ekv3P6uPBS9HOgdba9vO1FZJXAV892R5Ka7nbOkBU1
9kpX0v7wPm0x6GzKKGmgOh8h32TlIdQMIgExZBv9+qBNOlESjJ0CpJzSw87sYzYP
oIWnvXTjZ0YmD3lwAc6Q0cP01uWGhs3kCBicnjHyJnojjJ8LeT0cwuTJuLOTSBEd
F1C6KjqJ7AT7RDWUdOS/IFxFqI8/FFPqi9JzO8Cr3udrsigHugBo7TfsswjKXBz6
oJ6JVnSWjCVEm2kqHu3gYTJNP80652sw0smNK0JXWI2+azz4tur6bfjDJQPNKJ4k
tENFMFl1C7pSRM5DKjvH/zbRpDRi+XVnuzIdDQMwoQUWnB9boZjT7zuhHCWzWIBb
0vsnpJTknYNJOJSRHdpFNaKKcKgwfDm7IwmVf1jidxUaBeWuqCtUiiGLqM1hFqFK
L4iV/gcLuTWDZzJ4IpOQ0gY9ATnBzvWm8HmWDt1r7CcLOOc5q5ui/n3dk8LLSLOZ
eaWsDiBYWysNnJCICXE1nnhD4/X3ZvU0drb7IKcbj0S8/OYVUcGynvtRGArb7FDx
8LKp+ehF2E0xD5U08XFZy9r7IjOQeyBwFyMdlGzjp9PhMmwc8hS3Y+637/O59CTj
vxvfmN6g/6w88L6hG7LTlGmOR4z0sZPETGajr2QQVUGL0PTd/Z0faa/26JBqJGcC
GzfzhcB/uRwi8bgcF7dsewnt+WfiZdFJ14hj1wWOwNbfwDBeQhHYFz2iegs4fkvO
nFKHW0Urrux97qEWyiBjixa7kqdFPGfPy4Xmgbc0wREM7qnmSq4x0iXmQialFQr/
WHzdYYNKnd9pFQSAc3hObLnSBPPmmDPQ2FdfItPpykz61z5f/9VazIuEXJqAETw4
q7VlKYwCB791wCBd5ZlOHyOnz4x32LWeJOAdyMqKT4du8v+DdPeDUHUuRt6oHLeM
rGyvFHI5SyMnWibk3dozt/0Ji5cXnlizjMJMqZVsOXHfIim9IgA9/QXaEXF9ZJaU
d5A5cTdqXnsIJ0/OQPmZ5zmtFgMMURr+aK95GnDnQfqkB0/U0UG9XPO+VsXfdC5H
Hb5+X7jS/p37+pxftQD7ZylghaDEBpw2nksCHSuHcNdazL3aFt2kP8d0s/gETsSF
QSyndRwMbXJkhZ8JECc4OTt4BCRNbuvOaL8bOMzDoaxFlvYUikrXNNBjis4oMxMY
CiJW4BaEnVJMikrO9Dn5Q/oM+5eP9NH3ZhXpsoqv20siviLH/Jplz49NhzIQKaq0
gqFt+VE86m+Svxx67Sr6MObXAdjMsPRkonwUoJZpgSKmKqB19NfuIdAtTVTTDxjD
wEZNIHo+Ir+aL7a+LObJRTTu+SororCv+X7MkgcNsA8mtbZItbB4eJ+o3l3w5Gii
3di2A+If6vQMROV/VaNp6f415OyIt7r/D0PhTUVjOR8XvCxdk6g2CZMPnejouTNF
zb09cegR1fTodokqpB/v5cuyK3b4IFhS+WPpK4nuIIYnjM36ruh2jtmUQ0HcZH9Q
kLvVZypz1EBS0KHx7fawc1NRbZBMD4UEx+MKt4aUxKrWblDLX2Ackita5881IAnw
HfNChporaMfv9BaRs5VjnlpA9Z1in5qjZ/jBiUzYUgPNraqNNOri5Hlts4dbGuD9
GrGNJQCvkzcMLzzByslv3pBe6wxTQPMIfdpNClK1096upr1PZ7FwO+Ua6KsVNnzA
2/rtVtNDqeBnsdmVEW7srar2yjyw51XCjTTcX3AlopsBWfz6lhNij+BDTEjxH5t6
nEfVY/kvWTg3IlTMpUQah/1EmZN4W7YEXXy8xmX/1DgHpzpWjosAmb4s9sDRTAY/
YAvXGBlwUrHKtJGSIVK9hxHGcZGhvgs0CO7GypuznLuXcYTF6JaNluNKGDuHfTIY
F4qqXRm7uPdCdkIdqkYKt3Bvm2zejCTkPTo2E2WdNZwe4LmJXc2+QlWpmO6kXXkb
iOqQRNQVZJhc86bZSacKOlFxyAca14iZnswIkmuHdjvFmroUQpbfpabE1aJM/K+M
88I5ECYCrDzA3xdljuXRfYu8GHOpcPF5lekwfWdx4ib+Zy4ntE16FO9TFFElyGwZ
+NwRI2xgSdzwTLqPXeGTHdLdwqvOPfgryrtxGyx9RR127XSD0tBafrlY+KVoHkrG
Kck2INQYKRZm9VGo2thCYHrDKqtT3nSCPBmQdtHamrC0KG/OR+s6t/LH/2Ko7Xlf
QoluR8X8Gusrg5xaG8M9tNTyS4dEAd9/y+O0UfR356SMhrNjwFHC+NHw5OMQVTQd
7fOi67mCGDI7Yljuv+WqQQDKkuLJqEshzmZdT7YrL1pj2B/ZY7EIrjxoVA0OlVY7
AyK0ovi7AQXizMAKUhKpLye5e50yo9x1PVdzJyZ957f1A4ExL2VpWrzZn7cnex+I
l2savQfQShGmc3bbBHxvjapAH/h98MRUr87k+46ODP7yIQMEkvQ60l4xOQAqIOPi
20bjTDB5bjto8XLYxrsJ3v1T/3BhO8wmmK6QjMKFRNL/eYxbsSw7xQWCVILQjhcX
UVGOGGKODWlKrV/IrkimyWH9CVpy1JCo+Qlg0qQWUiuYZfqYM1eZdb4JBkLXEMCe
fEbTEteDONF4goDY+Mht9Q/jol/aTIU82JzZSLR+whbDWclKnLWb5Vt7sbuhgjik
1qSqDX0JqCvYTC/j3XGjNzybiC37w/TrbU1CWEzLIrFTRL43moeu22avP132A8h2
0lQVVjKGVC833E5ZYYf+JOWkSGMn003TFBoMO77/gH25anDU6Mw1ntGKGCkFMlh7
tjOkv4GyinTg3CkYphbejAHEVDS0eWMgyTM/5r9PyZ+1viuMIPbUGjU2YsocIg7v
WH4ca/OIl6T7QSECej3MoMA5QSHrMgJZvqFhLYjHvzXzM2Og3nweZaxemFap4Lvc
/44RXNszKEGyUEXyPg9EG549pddsTcb9Cvic2sYYwnm+gvYcUnioEAjoHQSRO+Ai
He3hDyg49rRKlKAcg3OAvhQaD/F0SPp+FVLa+PJ9C0XJsjDP0A+CQ4G/EgflJe8u
noLrVn5aZrg7efk3W8bqWoix2tk/kCPE3AtAeSXSk/xtm0ZCJgoShp4fPIP7faP2
VMsjcYUgAHbs6T8vx8wgoBvSj4Fl0yraStiyqAeDmVoLVQjdkRSx/WQFb1Kqx1R9
NIGlfLKFgUnzVAvfrEZHdjRQxOt1lrKx8fagq5ix94S3B9zAj0WFZy9ZX/cmPM0z
+f7lpVM/5tZgE5iOBd6W49tn5d6O2kI6Of9u+2pjQu8U1tWsW8Wk8yLBl7v61EMi
+o4JIBYuiuQN4jF7SK7OqK3UKPyteNxjz5BCWlNZH3n0ObXzwz3B8lvGUP2Mp/4o
7JlKi6s99v9PBDGW50DhgTRr0NTK6PIJibKjl8iaQlHWgdys8gLfq3BQIJH/Boz9
ECLMB7tsk3uIZdCeVSgFBRl/FCc/5WAEGzW4olxUhXNrAlPls2/kEJjf2qTxFYts
+GdblZRXtTrNB8JEWzeUkJ0sBfl2xXZ4qi1LdU+0Vt10IMUVehlIXOYRbreU7GAu
LSfNzv4DtVuaf6io57zjug5sV6zA1NN7VGi4VhAjposw6Eh5BaigEX1zwKsSMjgs
ppm0wB4SvTYSkAoHzhSc0HEnXBGLlg6wuBuCcqSs2t/b3pDJ2TLD9TxNnRSozLb8
UU7CJNw/SrRlVRAwRtf5aQapv1M6taeoczklmrMd+gYNXvbLMh8KmqIvLRwKWtTg
iMq/Zik/DDYRgd3yxn52Pnxhprp2652w3O9T+EVUFOhjI6UUb9i16YI/yVUKbxRL
dAx1N7p8xa0iUc8PcoKw1ZOjll04rzx2vMz9QL8F35SpHM9Pwm59ev/J5XylZZSE
bouxppg5OXEKNJV1XwO4cUJkG+F1VnuHbdWyA5JIpEM/wSFldWTFSXg/uYWU9SFt
2pPv6rKuLk2ZbH4t4Rf3Q7LLI+/RXkAuzGnzkhQqzZPmhSZPT8HPCIc/pay+g1Ra
0szaZDoH00JfH9Y4ENfLdyb4t3Yijvzk7tLsu79Tz1HNtGV6qDZQ/eRfsT26sn+N
7gj2ZcXqXYlE6/QwSTDdU/a6AvFN135qK6TKPt6TkN/4Xl10t4RHTlI5j6WKn0pW
DxHyArMjVezcZoiKzZFdeuenbWJQqfnC7xmFfdtbQZWAUfTejCNVnz1B1cWXyJtU
xRbhknHTpAxG7pvB3qPul0o9Zh18NAYrtkP3mM19Po7CmvtGg72Oym8GdswWPiTn
qCFoZseKS0etXsxBmnsF7q0tLl8SM0/ocDgRuIYIvjrCcqz1b47eaUiJf+XTinYQ
AGnWnuK+E6Wg0onpem4LmMTJnYTDMZTEgtAV+ktnDlDpbxKgKBappYn5jOpYcpI2
1psvrhINC3XoWJ8Rqm7f+aund1zu3BSvrgawlmEX7D/4clCQEzQd+f2ozuWbdM2K
ZVKpiwjXovkEnyxobJ4Yc0tr7LnX417B2oI+oE9SQIBli9bQlNDKrgSNgt/38MZg
s5KhIki1s6Gz6UfUvHjhOZb25XKKieX6udLCJkKQzhj50T+vfeHscHXJqEiFHoEj
x7tb8XXAT1G9A0MofmWnWGAlnplJnBykUuhxipt3JNABWMC38NEN80MB0mR3GQ1w
r2GoTym9oIfnKpcUx2HupbdgmO4Vi1D4o6Fmq8belEEkSfePQr9V+1YQTaYWLqh8
harVOk6uzNpeZUWRP+gthUcaiV6NEI/t4nt53feA9Pp0XWhI7GWIepuSLTA7iXrR
bDGLykSvqV8KOHXTafUK2/C0Dn9FNm7ISYU86A+V7A2UO4nfNrZ5InQsTuCe6tXt
rHa6zLrd5mBxCeK7kO1RxsfShW2STWxZUgPHnyLDSmqnjDnMSYZLUpOY3ZzngSd3
+C4Y6Tf1fBmXQ7ZnDuaFVqBimJ9ViVxsbyJSg7QYTm0wYGfYxF6K6g+eSM1nU2iE
L+apHsbM1TmZLRgqggU8CcuUAh6h8J0B1+7wrkjK1UlxS75UhMnO3xNrOYw4gckf
mC91ZGT/uYQfX2jAReXiLFwBvq+MC1I0JhmUnS7FSDLEbyVjc8uOMpRYPSnONQ61
EczRAqBcrA+25ZL1e7yZyeMWSQ13Okc1VNiHMCP3uCeKeSpq3Np1HteEsTKjTTbE
QrmX69W6SfrfiT6degR+z1cmkCBY9REdRyGev8DnQTzI4O3tNwYVPmUjs3aPgO4c
V5/ymgcVmdncU6gv/iWJlOUrXm9KcinAPkdK+TM7a44Q3y8qAdlJuEvXh8kL2fr6
Ro7Ynwh9sx2AlEGbOsETqqJtoFc84PlLVIFSnJ4kpktDtWZIiPotZNltFC7kTB0N
Yd6Gt+yDVHTBc8dl7w7vpTOpGYTj+e2P5TerdCdFtQn6nOfiOuinIgGZuPODtbuL
BKOBFBCdOFapuzlDswYng1Xx9QVBjaThK73z6Lb8HAF/JMj+DbYjA0qJ8HfwbvPU
6806sOKgKrTQrbKI5TPDnhUbDe79Ntq2y99sav4zXgXCOOpLHh7WdA/JK8VYp4ae
uZujHLW2itJugfSm0kz/relLgNwKoXW2FoQXvlcxauxyBu1Skn0H8H2akg5kmm+l
s+ML0VlSEeEE/1n9xnQAqOGpnz0HkeuUKnuSr59jEgsDZuSDYY0eeFqSd/74NIsy
JU/q9p6iRNBQrTD3O+HrVe5AwVAQG30hp1S8aDULXbI1JjD/tESd/sJy6bvFlCCs
76yjxTLYJ6c/QaHCGm6uxfGLoknYl7qOyoDal4VfD9FYfAy4QdWzFSGAr6oWBIfy
x6RXJi8K6dCh2Z/Vs+GWpkWTQCpmdpU6TZXvr6JF6izn4VcaumzKgNjJYAjkSuvO
azdIRwZBxt8i+sbc2HCfpdZoWvlZtq9r4zvGusdNC9uOjO7NfrZpZM4PXMp90Kol
enYkkP6n2yMfkgFtUnVIPGLZVoA66OY/Jg45+VJpHNRMiceREpbh/4TiPgPYWWnM
+wCqx9mjyenq1+MUOVrzMo5ik5VPbyidtjO2pgE6HOLnF0NCkQZ//cNrZE0FdutJ
NsumENeIVj06OGhOLjxjSls4MnDEK0DYwHt96KVHG/f2OY+r73Q9DPqU7WNWd4rv
nUBE2TAkxTELErIOZGFhq0TLJBAL2zYwXTk1BAkgYceTrFjsSaztR5Ph5dhe1fHq
RatM6owmx+ZB1qVVvEWo3mPEwNa6xQwgn+YP62r5O9Gh6+mxzndDEaTaeFqRJR4B
E51h6zoodDPFalKSRNtG3rQOCouXBUylThaJE5N61w5SpmdEhyw3GOJdAtYlT8WQ
sNYBf7gb8HerJ4TPbRafJ6iel3aWOa8/JVSrpl2w1dwnfxUxqwcULpKM+olpxgF1
TWvYRRuc78FL+JZ+4KqSA8/2HBDoX4EKqDrtMbMkQ1ipvvK45OfvteUl/3UZjQXW
7fDs6OwTClOra2HKxpH+yyMQh/CCBPaXQrNmkK55C/xmc48mh4gSA6MJ9aFY7vN6
OZ+aCSuNELZUmA4s7WmeBz4KzyhfMaaiXWwDnAc/FoIHexLPpTmtw8qk7fMjaGq+
zFSPilVtzHeIHnn3/HiolWdqhltf1LSPmDtyKspdD/ZoqOrMGVqeHFgCx0F2u+v/
89afDjXPgZoAo9Hn07MT8mMhmgvD4YUh1cyXG21ViE062MrBxX4whjYdeuV6Bxn/
KCnCjMBCSA1AESJ8wLwLCNnDhJAtsgpqmZXTudlw++LIVDBixCFgumH2jmtNw6a5
gvmySfSpGSJL8zX/tzTd6NDN5zaDt7r4hAydsNTht0TMbQjuCj+mesS/kE3Q9e/l
wNDCB/vCOxq18w0o202YS5CwGGbLZ4yCaUUaM03B7LNe/wau6Od2GwXGjUfxaOrB
5l7Savv/CX96BZLIIqrji5NdGUrJxqTIvNPsHWy4wZYBGuV0moxtxYuLWa61JGiO
YxBLxZn0ydm/zshDVgsZoi96s2J64Q0aErnmxbiuRVSvJyF3ZxbnBIRjCRQuZ9mF
9h+dQaOCY/2HIjrb8NmMeawY8XfcjLxjiGIPRBca2uzzwNDCS7sFo39chmSXuc2Y
TAUTImwC/vu5WfHrfgQfzI+idwk+hm4FiuAm4b/lByslPTacyzyECtrSoUdFlYh4
WFUA8C/aZWSYT+PW7CyWt8knbF2WC4k9e58BPVDhGRIcZsWJDkRLPj4ubW1CkS7c
LJx6jGed6aqsuh/WWva2Oh8DqopUDQH+lhzMLnDVBBmTlOcCwj4qDZjNFYD2uctZ
qzMyPG7VkxLum1/Ji3SEjtGHBUm+4hs9avij7zN7h2UeaZPZe1rT60w2uuBb6l5y
gCFh6S/CpzmBYMv/lyHUvbVvjfhmxU5n+K0W9HjGmrntoQ7ZSPEh/yjsDtqcNNrZ
fJ0wSBB3Jh5INCt6f381k74m0nlH7r43kG7yweaaMk+wzKFwEVHxbOnZTHp18NlQ
HUVg5V4U8McS/t3HpqmJ8eeiMABUAmdR1Rp+spGShl+kjjWCu+IILf7khZFJE0j0
zDdzjdrKz866/2/K5Rp8K12dcDjW3Cdhgy8jvxQxtQC0wTWzotjf6bRDpBoy6cl4
lvxRStLqIMnjSixA1zYNumkjFTqOkuZw/Xg93CYHobkh6alk96qMG5INMLOTNgl7
+x/pydkT1ZCbzgcNaBu+rEBx/q2hkXB7fHiMsE598SQlXdgBW6PbU1pyIi1H7GcL
jKasHKaGqv5duquCL2UME9GhTG6mFNcGhSBtILInnGtgnjhw4xbbfNhrldAOX6bF
imqh8rm7u9Hnva1BgJWvFqN6GbugVLXVfl5PfQnfHCnXtU6UZhgrvaQQM9QC+W8N
RV2IDOp8JyiAZUyUd3v0qemg2e7uuUcPUDpp2AEaksrMYWqkysUAgbEEjZ7gQkwr
NMfWduAqfVt0MvlKmi10+0VY2B/QphOHLvFOmLATq0rJ8DQekTb4HBeRnLN5ccNA
i/p5U117Fcnrc6YTI9jqgpaXsXKel8rbg1vnpsLgc29+DgAD5ZRIMDMVJ3Z9dsXc
AOdZvEVT7wzKLlBuqXmn91v2KB8uj+KVGhmW0bsx7RkpnYti1za3EzZn1Dl3BxLs
MIDUurawGzqM7NHhBuY59zJfD9mD6C/Xds3TkyNvv8ibGSZTnCDmf1KSKwQJB4mW
AJAdahp/jBDGjjHU5qPgHgfvonsdDHynjwjd0CTbUnDh3kIHoXXdjsXjvXpi2z3q
43qsjXFIY51zfhJ0boClSxdIU8Ioo1nzXGz0zAPIKdAEzbWJIITIiBGUy9Qlekjk
nl1cRtRKgAShsD6Qq0xC6ljlLf2I6NQzyn4HtXYINoov2YKBb0tQiEJJ5MznA0Ss
5TuKIALnuyABUhNZE0Fs4UBgjteuAiBRSEgMx3VqPZtTeCv2yypiPT4de9MHyV2A
FQrXpIlwVH64sc2JEmXhid03n142Nk8bIJOz0MtAXHmwoIyegjhJBTnOPUirPGdF
eYZ4QfHxUMFDC8fosWj1maYes1RT/SzCsMVQBrOwUu9KlggqKu19RR4itQDDW5oP
xS/A91bBJJbten5AHFgIRRXTuFwXEyt8eADIQQxaUDXKJrprX9VeBp9iANzS/CET
EQ+TyGcIB7L4piDl8V201SkOKB9sUfsumyPrxbfH5JmiXd7+DdtBn2P2gQD1UJ03
gWDldocjGfkyduTdg3JEvaAiZ6IhBqPga9XYkNPXr4TOGM/UAGy0gtnIyo4ZBx95
FxrtGKj1lhDKEYv21Bmenby/qRXmbikSfWUTtqSo1OOB7mLyekhKA0j9k9GQRKt6
F+MVEmwv7fevEZ19Z81gKKgimNPv1WoUiMjGpoyfHLANg55/rsO97+vVNGkgOgn5
e9AK5HPTymK8hoisD3+i8NRgg+On6wOezsRbA+G0HFM3zWrL0Pg5Mdggk0iVvdUi
6KzUyJQ0swpVhb0zR9zKXy7JlWANTXpVbnZ33qSef3Vs/PHHT94sFkz7xVo2yK+g
HWcobvd0RHGGjtoaNpPE+vLEeoqUvVb41ckAKMvscWK5AKAG0hTm31fPJn6yvA96
PqrsW+eIlotk6GtkLcWFUaiR2Gy2qgI60Gmez+SlNPkJAzBukVulk5Pp36y9auFb
VURAqMhJ24y7tdVWdwfwn6q3jNyli3FH5T53eW0ZFL/Q//iG0UnVUIPBCMcN0uHx
p4w/NQrnbPBsnhOYIjVeqYTNXr9NarwqSNcQo61PsRUfodNUDyk6NawEPWyW2LP7
aT1Bz3UbkM58W4fM5zEctUSWy+Hq+9mRVchLBuEA+TJ7sPw3WK/tBSGfLMYZLBtZ
6YB+R+fAhxJRgQVO0IiNJ63i9YDp1HsFFij3OmrZmIoxuZ+N2cTtOcZcgcrVpAWD
Qa80Crm9ZCSj8C/wSo6pEYIdzM9bbqqjtoIXAWgXJujrbNZ6Pa3Mm4m0s6TJpZpW
gKzTl5pdOgLLjM18w9EH1ZGauygOZ0ZZXLuJE1r8TY/3DkXEGThm3t4HNkMx2HOF
K8f9wT5pjf7kR0srdU4ObqWd2iosDlDqCGP1MKFpHoeFJJQHU4m123fRs3/t3BGj
7XUp+S1SAfgvCfHmcacI1V9lje63GCWFZ6FfbpYyKY/sFctDbXvuKhEXHuUozHpC
BTA18iM/3wnFzuz61TqtzsRfZE5mc9vO/UqQYL8U9INrIZ+/siPTSoBuwRlcv6nO
43ZvBrHAQfdWofOMK8f+ZPdW9h27dz4pSeDFIPmhyLNPdv7fXrJd+T59dD8ltJZp
gL9KWjjE2G/IcgrDh9vxasSDItz4/4AazVT80SpLKMrzJslR6jffIbJzVcWFkZaH
L1L4cm0l9tRquLLvjDOj7ECITlQKnkcmm7yR40GcAye/jKg8OpdlWjZ0rsFHRo8w
Nv8cAd6PLkybOwXc3XZZ5A+O5D8CSMzBnPVtc3WRUTuedyAHNrJong9j4zhgOj1K
jX82aZylWI/GjDnV5W/T8A7EyJbJ7ReZR+NpdT+DGL0Y18BlIALnOSgoQddiFo4P
HW1bBP6yk3TYQ0+uBjtL9796mRFHrhzAY27ECguDO1+jqELCLhaRg3IIuyy3Txa6
0g7vqe1xeJDbdgZ8nlibUMUGuKr1k8RpsjhA4EXaapzm/FrL17dGD1rKq36hEmgu
hJQq2MfU5qNVwNTg0IBQSFtRBWb21td0I9s9aSdHAAcV9F+9SISbrg8X7akroy43
s2x5d4wsQ2tOUi+YXDneWzaYz1g1kqW0cfdQSViR3m3wnyCyYm3RWJcgv3L9Muow
RjUmpVmsP88vRqMyzOwa7vYl4sNBZ4/OzXBcatSqZY/BYwRYtG0R4lXj+Sr0Vh6T
9bmB26XoWQUJlrfG0CI6X1Y9Aph/Xb11DPNzad7n+ZqYzvZaKlGIxoLDPmPmwxUn
vBr+MltRsKcqcOewZpLyKrVTO0FwSaiBabM1zFC8L/SVYhpbf/lzlVFvd7k5RFMn
fgZAFGiUeSKewzU2WzZikc+3pVT31lFRD/+aWeWOOeD1AiGsAB1UVviKO3TzAsj5
C8yirCpLkCMwnisjkPb7RNFK9Q5o3CoPFcGfxY7Lr+yZxSSjQ/PzwMZZEaxtrJml
0JchHpuoSBOZHpHQLbqXxkpa1alO/ZpAvYcM30Z44DIkKEEDwSipiQIe/wPSPTlz
gWdE36BlmnklODGEXu0sTXmSdUOVNJx9P8yp1obkQTKsEghPVo8xT2EaRzUhZ0Vp
UxOETAhFY94NP2lTncY7jtPb2cNuSoguqU8gg78lfKIKHLtDONDuhKInlB+Pm5Pp
+ZI2UuocejVP1EJL7SKEYhNQRm8ut+qwgDFH1/outbBAjSd9vEPVD6/BEEoW+b3i
d8SMJqLx1qT5dv1kISHT0BP1zTrzHnn+oNvDHt18dMBDlqhI/TqtEDSLV1kV24jy
nFzokaoY+jE9q/k9KMtIoQPQcSAt6JAB0sY+aouCZelI23KZP8BCwMdtOgfNh3+2
KuwrRGFLKZh7Zl9vQ7W1j0Or+rE/NpO0s2kinWj6kqT9jKLRPgp7uIGI8KmlrKs8
rB4R9Aj+jnHrO7KdUDPQNBQCgzLXqiWZyx0Xo9k6HgMuSpbQoVH76AoM1CZUACIZ
3XJfzEI0Rs2wGXbqt+m4ayar9hhZPROUFzP8jQnst2GAVY7wJWPTuwaYvaqs5n0e
XoYSyBRl7cziFo/2/xNESQmojYOMjOoOd0DMIZpxwuvCSqMUmA7QbbzLRlivve8m
vH3pSYkEK2PfXYZVHPNdoWFkogAu1fAUroAv5OiSqtnr7xeQd6ssdpWAJG45FrH2
CIDzx4fd1H4dVzs5dnUSder+R/kI7ea67/K40N973JVVt9YaMRCXWYbagJM49kn6
u7U8K0GdGUOdZwObVs8Z9FykjpArbEWmN7yv6m7D/7P+HCI9Jvnuc4pBx3IjtAEr
OJiHuMAoKfhXGtf0oUl5SgGHBhZZKP1XvLA2YimOJ3kfgPFYFpF4TAwNE/JZnDxD
XgJ2JgL8+b2/dfUMpDvwd4AsOLi3MWZLNEAkKhy0NlfmEdwJyOQG5D/PzswIwmF1
1FRr+hF//CobczupB5PHJsS7qJahIymdu9L4HqEf+t72Y5nkcvwhB6n1n+N1/XsE
SwU6Rbj5D9mAlsXI/bWPh2LKPhl8Kjfl9cd24Ol4mY6a2JsRPjaubOhpl1smMXgP
ROTUAv6R2qkpouOpUu17Pw0lEEx0YxcrG6Jc5ror1vzTBV7rGcnhf50cr3uX/yap
9Kva9BEbMPv6+77mw06D+uHqxFqKuv5f1y8G6e9Sypa0AHiMm0kWSRWMFf7g4Orc
q4VKMfQGlV5y0S70DrhXWd+kJiFIL/VXaGVRZKNcaNiKhbRL+JzZNvnZfkY+4l3u
pynGM3MoXLPx0+c81jV3EA6w3WpJguIWXmOID/ZUcb8uTr9TGFWUdHlLPcvu8GPi
pjOt/4RD9n4Ct13RcLeC59w3nE5C9JhgjVLeB0lKs6C3nXtkUJ9u8yp3yBgNUG5S
2ncfQE9xcvyZ1Tg4wabIHtIc9R4OKMeNSFJVAK6ZzD48SUyld3oQSbIBm1cy1pzs
616fTl/vi2GlV4LStTTdUKyZlCMYJGQXj0qK9/gmdJigswV+onDY4UOazcBO2fK9
HcsFTPGJYxXze3OKOfmDmYoUm9jikqW+itBq04Xf3pVIIa1NgZiMpMQpqJlVvEbb
07/5075BBF5NhDBwkWbPtVTmiMyOTVEVJu+cUBGf1nfVoLDuZAHbhOnMCi+OPKIo
Q9GHG6aSgUkHij/r6TIt8ePWYMABJr73FVtV9ihpVwfs3VytCExOTQGHYDRTUaE/
cpE3Vev7lpYtIvTZ3W5nKROFr4B3OxKSKh3Mxm8t0ho915Q13FukAjvYs6nJrUF7
Y0LnPh6zruONZYk0Ps5YzUYdtyo1YCEvH3+RgkSih+L+mCocOuHKz20zju6nx7tx
VFHD9kC7WfDUPYnpgooNf3dhBEEAcdvg0yp0YIJfbKVJErI+455bNja0aULObFAt
JeFHmuxCLoj010JrDoyblD+woIcPsM8QORF4BZuKzDPaQ/uh40hHk7WAm1z9Mdro
owZz3nzawxWQcgyj8SeWoD9IAAuKTzjx7pxQnzJvHJkEQHNWGzTrqNg4NaQwQD5p
ZHdEom/D/G+5yWcvfRdraFh+xrT3LG3DPS/5SMWhUOfVqDjUeScH81Ql3GAZ12WU
m2ITyIpM6ugkcIcPTUBQ+e6sCKLSnzf6JEbT21tOE3m/PEwyen7X6zrwop4x1V8W
8wTQS/GlinX8BQbqigU9JCjnLJRCJnplIqdQFT2UggFhSAQKmno1jY8HfzgZuiFh
Z2LJdbn2xZq/ts+t6EF6/wTPTCDi0UobZMuqYBmCCHhtDqWl2PsUpDVpYFP0yCnO
t3goLiaByhN7ubJ8JxXXotSfY1qFIdDJF+luKF+c4y59Yv/EbSUMOrNy9qbEX36b
ztd+mWZWqJabvBotRIPGkZDfn5lTorqBZN6oLUNMacNCevjgfy59lhIOTR6up3fQ
gznsgglmkZkQ6q6Q76sHyv3mFtsoqNo3UgnIyTBHlRiRYAFFiM+rFBVbaUiHhahQ
HYGfgHrMbA0+tkgKBRcIM2Hsr27ILmQGqbxHt9xgYlnoIDUBZXo+FHTZY+rpiK64
j6N5SULeSCTc3b5xr43JdG1/F4rl7X7YY974RjanN6TTnA3nmcSvcsBhDiCdw9CY
GV/XzOIFb6hn57hdhEzglownV/JWAwQlVXwPZ5r4RvjYIJksUTUaPkSK7jUrOpQr
Ze9R9Nri61cmOvJqFlelYTvzcchewOoFXaL4vRXHsUti+/Xd0sge7oujaKo1qQJr
sYV4y2VZI30qU68825nYBtX580FhKIJEOu/PyknUqJNeoKt7o66HUKj2TBp/QZbK
Vae/ofZlb0fKhB4t2JMdfstoyYzL82VYwzSHTNMJWs08AbkZM1RPq7krLjkFpb5B
xfZzMMXggLT6STZKyRB0EwprzQXZGJhqo7SztE4q706+jfCIq4OfQJoyFr1bh/sf
WW5GeJQZXXyCf0WJLPEADu+ftRaUlGDsvUZcMkIBmQR/emiteTRxuLXTwKMS12Wk
PyBuoWyUmv1nyqBvxcR2Qnz9bLbtYGq353H5/K0RHn/7IifGGlFxvf87NieY4ZaC
tgio4bqSplkoK19HHxu6nvsL5kqrvjdkaj+9i4gsVcDBsc77A9iD+0dPVcflKIGP
pof5LCJ+HobCXj78gfY0RXYPDE8mrffA4NnDl74wuDbieCdyjFXxyH0D6gANt4Y5
wMrTsu3l0C6SUyPZTIYEYGRcNQs5fsWAcpwcajcLOMm5T2JuxSJOzMSqUT2/vK4R
he9LrFmk1hDJrPfLMVkqUQnKNIqvICEWJVA6e/oXxNfkuUSqxopMKLsI8BtHOwAr
utAY0kOxP2u7epq19Sq/diFF6CVNu+0OBoUDyTYUw2/Z3urpiY48OMDJpx3Cj8SQ
OlPAM1GrFdnpmaJ94VrUsENMjDku+Y8G9j9hTYd6Ul4s5e/4p+EytH4HQQ6O1Iy6
mXRNaWvXuJdyKWEpiwyGiiQ0178Ne3AQzbqShxXyu1MfXF/WZbGmTfRTXbnLnOlV
Mhz1UeclkI7vguB3Wkk3mpQrQ+Ej3qZF8VuzeKyfvMGDaseOAAvjJ5OeadoRn2gM
wZ+ZZ4fn1riU3LK5gtDuJHxdEPYqaq9cAYng4BPW43b5lZ4WlB0lFNnLsD4uJ79d
7UBNvdtkCEXQsZ8l0+xhZ7LCRveAXCxv1TIhOgQ/P4PDRiBXFGHNP4kxBehujyi1
JyNZWgxtyALqYjS5Ujtdzf0/vd9vv7333L8c2XqkzGaIyZN6qaVIDzdyLCBifT10
DOyGizkeYShR8KgK9bTcz6D/lgAfVnAY1hrGDYstgV+sH+1WCTCV4wz+aOYlsSjI
yz8DWXpbQjcHSFaVPDOehDiFIenMGx/y8T/DVSndw7gjJAY9QOyPH3mMPxH3qtTQ
VVJWYFySBW68dJTw5y+AzmrwAn45e5MLGCuLhd1ZbLWaM8HSpnnxs7s+LtDLgTPu
Lpz0APH8i3joX2yYR2xy0qZtsb+w+ZD5CYgOBslCdUaYsIzaVkJHfVFhBgZO/fzy
7CSfV9iKG+iSEcOiMNkLXOtTg0WY7YpE/YDU6eL07RmJ41eZogmWyE5Iwl/tjc6j
hDgkkNUSAajaC1HOgAdGKOUayG3VjKKaC6xbCESbiVeVLmL9pAUJSvENXePWAxFe
cjYgHkDgKjnPT3metWWH7yVgAYQW5FNGXkguYkqMfZ7V3sZaoivepSUOVKfNfxH/
3RjHG0qHv4LXow7bD6FFtFlEIWXyaLnPyvkrr7XQeZoeGXmM7iAGQp3rE9/FY4o0
m28xv8OqongJx5YKrPCyytPu0a0VDjFy6jS1bDeO2ZjzWvzDDhLp0NLT6CyMRzaD
mM8drheMsBcv+SDO/bAd94Wtp0XGYO6kOX5mmomU71VKhY72kAg77O5ZWk0QMxt+
8GgflmyZaZeJUm3QFz+5i/Ar7h2fIxVQRuhqKIRvLXK0yTR2jaOZKmEMv0fBUP60
r4AgNpP/5Q9ISC0FbDlov69v6IMR5vhyfvsHRCP7jGhFSOQwd/aCDLqy9X3lVT27
OrL8ikWwlC6IMRXc3SkTv2dt8F2aLfywwQ5SqCSoJKcFD9Hrj/UX6JbCpZtl1tqi
UfAZuK3YIYI2OzO47uHKagpg40DRuLO4rC7QlJrXEE+mHPbOWU6xeVnR6XWKgooq
BrEOLJZzJ88ZsrPhMP37jGFjzG5xEnWQgCJoVvx28WMzzRBdDbif4Gi7lk86A5rD
UvI2UE/aJs3ABCqKOT9WmJdh2hNOQeesZlAOlLC+PrNn7oJba0W0gM6bDJ0fYdmv
gH2zJZ1uLnGNTaykjnwiztbap6jmRMKYRz7vPW17L5tXWG/XgxTxNGm3lv9glCzg
g1RQA4Lykj6TWJ29nHVianex+v4MBEMrQwC61gUquDNyqxEd51uwg/2mnzXgKE5q
RmgtLhbsGMYSRubCUE49zKz4ABvev8oMrc62TpO1Y+QGQUI2GfC3OIsFy1ACzmqC
O6g2b7k1wSk5u22mFXoJgnExdHAFqp1RQJYHebtI4bpvpv8Fo7hA21ffumDfx4KG
fElnAeLrQfJkblRqu15PdmmR/05WReH61wQme53z2fbnNEy2rCnn8E/GjFrGz+22
u3fcYKRnwW3ZmGI7tELDHH0EQJYxWrgMzl/w6PXCvyKlpGvjJxG+UC1I0Pe2gIuQ
RmZMhYoDrorLy9kA6JFQe3JFJXbDgCy6ueByYuAHViTjQPNrJoeSt2eLz2ONAsIg
Bs6A62TD+/7uUBoqYaw4+jhKiaBv4bAOKv6XU+QceQAmbSYCNvxqS+nf2B97DNCx
+TYNf2gg6L3CAmRGM7zXK+em5PINDwrvLI2aIJxR5zwFnIZPdOwmEJ3sbZlRU3wu
iN17x72TXxmvAw3t6tf/M1MY/gJgYoztEhSZYfCwyaVLd+TaXDTpQ5yP9HsI+CJA
4ErOboqTBbBkR3jHnTC4ScmOGjfg/NrPbHr8iruCw3tix0edqUtS3BqnpaPG1Xaf
vEv+fmShYsY+k8pJHW5tU8L/94zL1r+3TRC+iJrH5zCDGBsn19mgBVJPy7Jls1xL
h2LURqg6oTWNhOvltjldB4Vqshsc1nWA1SiIORhQM94Yrcy3eNJ/DI8rd/1Vgzsn
ZlYxWfBqMC3s5Amgem+z9I1LlC1fTSeNL3txmtNcvoRa9o6cDV4cGXM6z55xq1uO
pW4o4PxIaLnp7rY0cOuwiOj1xykUGEzMggeFWf0p/+vVXXX0XaK+lFEUIw7qgsfX
BS1LAgT4TUEZCE/APmfg4HM4FTZDwX5gmFduF63lb5pr5+ymRyn5O8XZHAdwErNc
a01tGEgN3oTDiQEuxvnikkOtOE2K1zhy89W130miJZf9MlR18QvmkX3vSzepriYi
s/GGx/guo5TDKGsqYwTPs7aXbQ1GZUgHA2S/7TskY6nU+8IfehSkejHqRBvfqRuS
9T+26CPrldgo54Koz/9lAdGU64XHpoS0A0Ssh2GT07LsgfX2/55zsIDeGUtiEBaq
UZsn4/7EdzJGX/cwY4TXJhZHmtQY5Asa8EEdmduC0r2b06ajztZx5CC1Z1IOTDi6
3Ev/FOWYEwoSA7Q282/tcLHtyIg8nLf770jMnQVSMXsBp9vDT6oLOsRIp9zq5a66
2DhdKxs4dWLJA4i/HKRUcViByGbt12kcVwGsLM7TXjnRRsQIRDs79feciKj49wYC
1WVauctgDKTdoG60MzqPWW5dIJp+Lt99OxWiT+q6LFYRtRi/D6n95M/QkhnAQzgH
iT1bKXinpOMWZcXTszpdXVs3DNywUQ/N0Lty8zCZ7FdOmykVax/0PHzHpvb09oLi
TBn7cvI9AnjuJuCM7AY7nBaD6pwWwfm3X6XIrcD4T8WPwYQCc1bXWqHthm2C+KKI
oUvmG9Giro0wLq5NBHQlOSfmQRFaC9lx2uNHptOzXjGomTEBj/RY8kDa3Eh+rSn0
Qxt5fySabxeO7y+6dUH5eoIVcEzDF3IhAMb96oTT7R7uBhx0D0JysZjin0ASgvos
GPF+l+tOccBQ1SO2zl839ujzLWSM5Z1jrAPS0SdQblDtpVOPWnKOX8V0fQ+6j6dj
YDc9t2HPJZzUAlJ4HYrJBpP3i2yvTfd/A4aBGGkC2P7y2h1NlHMAYV4/DPrvoPgK
VkfCWwj41PI84UrGKn9CAnOqE1zRPyRQE7m0tpibU5lUPCNlMxW9rD0G19Mk/yVt
eqQhag4F9lxWxiiH0PjprjiuL0JchG6TRqEWsq533f1Ilq5anV6cZO+hQwySxz0X
KZD0YMpWo7Jt7art1lW8CsM0o/XrSmJGo6cEKZvVqmvS9icKo4GC4ScRNwlBhIBf
LKz1bf3RPOKex0Wj1tC7akDRVJW52i6uILON9aoMOJyRWEistrF2s9GwZr3Q7UjB
UFHq9D2TxCq0wN6lUdEfeB1bfQb5fS0nGhPlSMyrIBNxIgeWdbkJAKC0mK7PhPfJ
X0SNqhzHww7bF/d7ivOLFT1nhZfDaV27bWj7yXzj89CSmS5bI0BPUBo4R4+94hZG
0YlvK/EzABooxjQRpfit/rtsQEWFz+lO6K/4ibcc3NbkQ+Yro9PAP3+jI07QpFe8
3+yoMKAnCwKzjik5AbNY6BuZ6fi0KQjiZ3opxaAU3Z8q1cJfuzY4fcivNC0oOzII
/yU6zFxuqEZk18fYcbwsOZRBCu9QHbuRKKjDHJkuTnmxN4VivIFyeFRR3Rr01K0T
ysC88zQVLEX1F1f0zBM1rtaLcVw2lzB56aqDZDyjVV1f69z+pmKR7MvM/tnAb15w
7+NZdmRtP7WNsANYwQtQGtDn47Y6aaH4nKy5C9zqmOIYh51/uGsv9iB3c4LL4YMU
fZC2laBA9EGv/tXWlWRTAqJn0SWQ4/uyqBKM9YoTHPbrLB2SOR/Rf+C5vdAXWx+a
wMua/FzQmDK62mMC0Ss7V2aAL81RRB7dD6Jl+yhGOl90Sy4N6QUx4CU8qG9Id5oB
i/pusp0tlgPRm1o/72ov8R1R9E2UQgVlYnuLXXP/JHrAiCQ/DZaX+6Bjmp5SxAGn
1ZamSryZlxz2f5Ss8SZitTpA5k9DcY+h7kVSkewdrlYbCJ8vczQebMtpx2K5nHEk
7WQCAFS4zSvRt0y65ilv0OLtkdY+VbmEqonQ5z7Qu9W96Gf/mivXg0d5a2cy6SAl
6Cm4Z3XgtZr67jKCQO+I+s0hmxVlhrBvKuFlRXc1MkyTjdWbRUQbnX4kLvPVMLB6
nu4+/CKHkigZEgc/vnn92v7NLR2seLbMdIut1JgANBSa/ycCdpdC6NJuI5oelGem
cFTCPHCWbqZ7A96HReliwxItdTHlBFCV2JVhb65WIlvcIT+A5ZRVZc+/DxoxZens
7yOdu14e7Lw7QDvrKXASUUo/uwLkosus/YBFdD9KbSbLXTSk5TV3sWOR/Fffvg9D
6hONbdW1sH/AjFUOgL2RhleoePKBAehuiyx7NdN/qBNKClRq2lYyZaGS6bha+k3H
sDOogCnaV8CqbhS/ws6wIqHTDzaSImWjfAvnkkPporGYpGVBEnHMuQGxbq0Pw5UU
29n2YOQ7OeqFQOEkFGLKvd3puOn9inhDmtfq4WRR4SRV205HlTCq7zwsEey0scoE
QJFs6U8vpKq/WMiw54nyepdAWDJV21pvfpJQDPSGcmkG5RJKcMBCa2t7Ddhoevd7
Cmo9i7BJt21Nv5C7a14SE9naKBAmhvelWKss1OG9tjcxOC0EyKmu3BLX8XrGiM2n
Aug/yOdUYMazwsO8PduZj22VOny5CFf5eCRD7LzY4gfZqgoWVBZUuZsu454Whoqb
TIwEQoyvAYf13zIp+9ongg7kUwBirpTGizMw6ROiLWXrR/UMePQfFVCAD3DfaW8s
d8TZjHNh/Mi6UW4KckEkzqJhz02U8AE2AJ/bAIwHcTX3Tqvhfaq6KTfMgVvbbQaa
Y8k6t9oAnF0LPgCgtr6eix8WXDUx/bGtFSoZzecJY6gOxtFXSCIx2zGDDdWadmEU
AuCaV/pNOfbb53TMZ5OP7upx6iWrUB57+yaPO4HzAaJYso76dpdS+HTroVeqYnfU
Q1r85X0gN0IaKVetsHackyJrwjE3vTgETYZjP6HLp4aaXenw+InFVob7y+uKGbqs
MmSa+OTct4c3LbqlF+xtId7H43DF4CQ4yVjt1iprYg38hGenb8RvOoS1cTZRH5Sr
eLyaF+GMhsCF7Ol3m0gYWUy7IdLPtAY9oxiaeb7uwbxwvThLxwHYWNrMlrjUzmhM
kiNbTfTYkfxLPBR3EYz9Tu9antVQSUW2jYbA1FKEjGDq1k8PbPikaN3FdxAO5EVu
yfuZQEyzY3fYiatGX+I9lGW3LbXMWIMPCZPEuOgl9RFOC9fMex+HKFQE6F3QszI/
vC0akH2hY/Q3HhN4xoVYY+/eOe+fNuGmjyb32cHhKSzuZTCpfAVPEq72CfrD6McL
vH1p5dLeZf7IAuEkzHxI4X7hSslRD/lGH+4RU53+rELimY93qddnBLaGRHB/Ktqg
224MS/GARzcGHXyHJwZWcTKr7TesPe5jUG82YxZuDbQSmihvYyVunmzcrY99Xbse
bS+WxXuNrwJ1sJ8v9YN9pTfPd7Rt7IdcSkyRWon6Gd0RZBekStmOxjiqxaypxCkr
nUWdhi5F5lCG54J0Xp2Rr5X3jWhBQ8SelAcvjBueUr0D3avIkyP6fSW1gsKythmR
Fz+1diCUYhKleBljpe+4LBNXLHFLUzMI3dt8n3Gd22nfb1AfPxr+95Y8W4+DILGq
hw/dBVAlUAl1qiK3n5ggfKdGh13Ds69xpA3PO6R5xWpOzaIb082ZZpjTNMkq9DFr
pZT0Kxd4MwuE4NyAjpl1xWfvCyEZz/bnb6P8PxAiyJaGWodYPiXCNcrrOFUqnBwe
+7Iz7SfymZ+t/13rAdc0N2lFqjzCvpvfeohtK6H1xjG1+xWhRNE5U+/EkxS/s+dv
P3wnRzKOf6KocsGBwdxVs0T2vvXyisRBzfX83a+d6PdglopHC/3Yy7RQc66B9zc9
H+b6Ls8DOQ1Pdow47D50DKdVLS7dxXAWI62Zze06cDEqx/jWc8Hb9c8lp21+ni3G
L8pyK0nZqZ9Uw31TH7z9NWpaf/UkEmS1vkrtox/ORhXp+mj5c9bG077tx5V3xlR0
GMKs8iB5R+h3I7AVL+l5o7u6YSn+F4kSk50eC/btupGIdqG+LzPTsWucWBruHRBH
XGPZNwwv4z/R162S6CZX7x7vXx64t8wKnG+HlE+I62Hc88Vme7PnE4eJZzsLrraz
mtoRcU98LDW1b0BUzGG8IqaRmdx+TgWIN5jCR6Lrae/cZL78p/w6ylHaz5YTSHoc
FU1fpi0e7c+am44vByrnrk4rWMii0Ku0CZSAXJN/ZMIuSB02CIbTMUUuDts7XF7O
0cAe5QaJFzLxNv/4gc5AzeJNjoic7HyG4YwkN1BU0RzT1gIcCN5Iiiq1ItaUvhjw
DLGKXS9/RWI36H8zkNEacNdG7w1Fr4QQfxoo0QbMfmC/YyWeEENkkDRCkFUh6hbq
wYJFZgQGgolzifLIPikhGeXZlG8oqwWMXKvdiv9IZ1smdb4gFfpCafy/nVMWnpYJ
RNXGdwvUfgVMFsrLd0RN0JQe6I7NzcZn6AC+8Cx01k1++CSmMALG6JmO/k7WZnGi
2mV6OSt0QVZ6t3CXqL9tUgkWkz23PaXwz9xpVbg/XAodUfwWKORT+5wUefs2V/r+
+fRO0PTr/RhYp9hociAFSViZu+caBDvNDh2PbX5KDpbPgh394OyYb8z3OK77+tFX
Lh6KtDoM4ixAJ4jA+9sQogVI4ULvClfY4X1NVoLo16Iv2gMqb75zTFXHYP/l7EgA
7vGKnY9JriRXQ1ArwMTKqjUx80TWKDxtaJ82PYJSvvc/v0ia1434cN4GTsSlUIkn
+RZ4u94MAnSKkWorgtYTqeOOG9+/E45AkoLNLQxP4GtlAoPbMXLewuPJC/7/2Hq6
OmbddG3dffumqYSUqkGezlpuadyA9fjdRDk1RffxiI6covLPVnEYa8oVl1QK5ocu
iEJGaINi2IS4yjkJlV/buaNHczHtd2FYh4stDCduKphEIUzMlnmFw0HF6UJKxbFw
RUyuZgOIQu0NAR7dQNla+y6E/hy3w2tvPHwyJzZWY/LRy8ht1/Ek60Pwvm86etKj
PxTKrO0m87mr7cWqHTCkk99dpKpRpc2+ZpT7mt+WsO8Yl7lxC5aXH0E+h41UwBVQ
GbUgDChu+/8TsHc4MCFchyA/lHOvhmPIOEaP/KFwp/HmQpfXdWq3wjB8Jx6D/onz
6z0VHp8XqRuadxwuF6DFtrwG8LZWwWZFvSTtYK/iyiOSKDqChRvap0KtfQpekk1e
VwMPooFyck04jXD7yaCRCewlzP3V/zQGvrKUBZp6VU/EXzTTVL1TLe+sSlJDPu2z
IHoVEdACvPHeqLx6ZlOisEkPYCRU7bgSPOH47QlHZLZ+3USc69HGmST875uWbzbl
PLczmXW/dHhFHNnlBrUoKWuYGhhpBom2OWLjJBS/7znr7mqOKumj8Fj0Z9986XrT
9PyWgYnvLkiJiy3qXaZfviXO6cAoY+M552zhSpqy86bNWMjeFPlguOgQMei6x6K/
xqdd3Dlmy95hVnw0/CCTsWkKA5B3xWfESS0kycO67RVcZJgLxKmNgvvBPVu7l388
hbSjYln7NtidqfY3D7IXj1tG6D6ettQKKkynSyN0Ag55touJQXEm3EGAb4z25xGv
LbXOeIsqSR0yP5SN7G/j81c1DI8x4cFcoNlryyltKLHwRU5/B7SLqxA2Bfbfh4jK
e8f/tkTYkL3il7f3d6SCwTogN4aNtaS8/ijEoO9jWeiYD0Q92EXmDQxjyXcJz4cV
RYKj/jrRMNzvBecEkqoZpw0if/zMY0jN1sucPa9EOMGg9Qffhrq6TKGUK3PpQWcn
jIIdevsRs5MWvTuHUrXRd7Zpa/fDJeUNCTZLOZVRqa0qdRIOYI0d7+cO6jHqNpHi
Z5ROqnXOm0k7lkJAamnS2SC1Ll5wT1n/cImKMJ3UjaHZK07IKyd4PbhLOrDnsYlB
u+lVm29Y7EerbN4Vu9aEM54mUE2LYylWtiJqWMqzBtGwlB4hUjOOp4iQmewteAAB
2piOt8Gu54w7pFBT0c+KVwI4YoFZ0F0SvZiBth6hPr29aSocsuJtMlyvw8tH+dJl
tFK/7lM4HeNEDiu8fEhO8ip+it5hI9FYqDtvNKCZbcvhiMSu+5rvpSDUvPkawCqd
KLy6MPuht6Mt/egwyBckT61m8Z8ZsAtMvR999wxMbpBwHFuFAch4o85B+CVZhIsQ
15ylunZywv013QcsMH4CGOwjolilDfI7BHDHbJ96c29alpJgtYc9kojy3PqQi1Ws
xHYZ6FRkeS6hLB+PoNPNCsON5kZQLXJ2GNQmIgIv2BvsWIxcw65VwNp0iviUxxAe
l0hbpxmLYa14BhzoNYDOMJ2HhGalxw8vrcaNVYD8XBw6/jBlfmevMDZF9JeAwgMO
1mETpX6GAv5i7C6QgAKkS5nxX5qypid8BUSLpRTE0/9g20W9V0l4OHTHJgIHCfVC
Ei15Saf3oFE8LdUzJmLhy/KRo/FHjRB+5uYYbbdLygKpVFaITtXQaBMKVjhpIxWD
knbH5Ea7E2G16FAJkdaa4zpyYzscqcQfEezmKYYjioeujTAV+fJa5TE7HYDXVpqJ
U7AibmThmx+chZ2xV69fSklAOfM0u4LAknPCddqyF6xPLc+tVoaCInQuzF0DNkJv
Ecs/IZqkKZyY7TeODYy+swkUtE39j2s1ZyyRjt1DlFpyZNsK1g3fAsGd5DoqzEnT
pZBCQ6c2+YqnViB0yKN5TKeJauJRzaPyPw+41FXTKEAO6mhVg4lGrNJtWf9ZxIFw
mdno4p9Xuv9+sZdcE8UyqXdJyteMT4MFYE6ZRX1dmrudWmd2Uph/FxV7cB+yF4FN
Mmg6nIzGW9fjedz+nM1xkBreN7EfqLxOLxIiVo0XJ8nVvrkDQzwsgQ1QLz/EGgBc
P3Bv0RAe770gnjThn0Upw4bj2JDnsZv46iNkHyzXhhXZ/6PEhprNGZWNaq80hOaM
P3B2Hx7kX5wZyZi5pdA2U5fqfxt64aTCU05trnZIZNlfZ0WatQQQe22cgzou3/Lg
y3uL0jkRHhdWRB5X61MxAb6rgBeIAruJbXZnJbeqhlypv1809wf28+oR63iVEN4d
945KgHyQd08dnmO7b3w4Nf3D2r4WOrM6NWZqhhNYEQTkE6OqoLe4tSBpXWpdhDB1
3YjdzNnxa2EZXzxaVaK+EriswJqLifbvZC8MWKdmtRHnAcJnuH8CV6GT4sDgw40I
yezFnWqWk3qM26MQNpPF94PtIPcnmsHmdHCHbsZHxA7cmcYwpWRyOQyR+V8CQYvb
xSx7igpJieVTcPSNjWthWo2r0X3ol3pRhfz+6DYzb/pRni6fel/Fs+MDACpy/25i
54b0K11hccEFlgo0YQin6qBxxJT+OhNdMXDcNswU03OVhLSGeHupDGHfaHeyRGJv
g8B+6iDJxNiPmats19TQWPMSPfjAddputYSod3Ifvjvp0TDa5uw15qWTdYwABKkc
UMB9glnGdJlbFec8Jr4wf+i1utMvS0sQD6NpDBgqcmGooQph8Zqf+V/fzORFKkgv
Ad2kfU1tR2CpmcpP1jNmQfCKpndnbvlD5FzslwGvwp993oGuIFXUeLo0aU8JS5ak
RDXkLVqmQK0XclB3/1UQSHyNNStMctHAI/lf1JuMKhfpqL5UaMLuYbuVP7VsQ5NV
GwwfdzGkq++4yf+ehuSSJQjH5xTQdy5b6TWP1mjunOyUCN4umbnaL5K8kmeg/vDz
J4I6LQTYzzlUIPYE5N03Hluok7GL/dgrX0pOintY/uF2GlrwhxmToYx42tmG+cIz
ep2cE44dwzb2az1q06BaMD2sJgD5hn9LQ3MbqlnR5c0kiX4C908coyt2OdIogQ8n
bD4CeED2bio0lcuBm2CxukDqV36VUStR6/ZzJMyIHZdCjpdXFj0nWcRIi09mpoFt
Jvb0lfmNUKB6Z5Nf1c18Ai5qHeBvLAQD5Tc66xiFy93LXTU+orTNI+0kOcxV7L5x
hezftAmmUUSAXzom5paylasz5uzNboYtDcSG2zKuY3O9+X53s3AynAT0rMYjGd88
2rpbHCIt49AKgdU8UbTKxYQOcuOYcjakxM73tXT9BGfWn47Lu+G6G8Liij3QjsxO
yz+EiS5MHdNcJf1D8GOWiwq1ymNFYP6mxYq3nOar5hR0K+Ai2pYAQ4t9AF04WiHa
rxlOkvxXzaTGzazycU/ILBt0Wq/BLuw9walXCWTXasOj9uSGWWEfAJ3o1eY2DqBr
1LLuBsz5Wf9dQ0ik/XysqJqgSUHx19SiddanIIRcvrd7yz32T680BkZ2MTbwma5M
4LOikz2Y9Jd7nH+eWQ033Mhci8Rjp8Yy6K2F9kCRZuCdy89Bzg9v9S/SQSBYCrJO
y402zWa9JzJzZj5P2US0lYaAi2stA1Gq0VwMZKa5rLgrhidLQTZA56OefmV7vvcj
fVqvMB+dNLEspS7b5ge9Atnoy7+gs/xgTreuGpYQLQzTLDvy9apCblkisB+hEJvv
wjwrZtE15T35jt0DrF5wfaUZiiV+3iaM6+bz9kcPN1ZceimcO9p+BkSaU9sYaHkg
uzXr5OvgpPjPiW8vNqldy1a6/u/2Hq+VyNDvT9tVFcVsvBBH++HJOTrnGNarAT78
/Pg08Zsmb3HwacfeiN0zXBr1zvRszEymw6GtEwpKm7YJZy3yr+GxpFgA7KUTMZQg
oZQOWy9hLZg2sn+afRPc8tKZShsTIT/t4EqMM3njxROzl0aZbSasOuujfdAqK8nB
kOU0cnl+ThWO18ykWpL0SpM9oKKTfnD64RQplkwVKPDcOWMuk+bBvlFxI4GNjvRN
SdkfWzda/YCTcWoTNLyeOtT2Upr31NgP4n4YbHMN47tJ4boEII8QXV4mLjgPFXj3
Gii5sAwGKyJl1P42xSItvVaUAHxoo/dAm4zh6vV8rfbgDY6a3X/ZUcaT532+Obv0
0LKJa9aeuiqamN1yeHJJyhEkjI7buSZNAF5hSludsfvwKj0enGU0m/lS2wELF34K
FPTeIAQtCYjvTbQhltpIkAg/vO4p19N//xsWeM9Ay9VS2HmKTCFrHwHv0wWDSCcd
UO771NuQp44a5zpLXN8jSCIU7aotxKaMTe1xjia5xsLgHqgP0Mzb5+zNdDyjuxr2
6bf7v29CZWPqTG3GfKsFz/7na/RIZrCkPvkc1AgjnB0o9giE28FbEuR9HtidIOo3
rU73zpG7nGhulIG/HJcF2m3BKG3o4lVShyr3SNrY3HogYcM3dUOhlfskYVGXPCAS
cQhd8pjgfjg0Nr/oWGlRzH8h5OofivtuBQL6IqVdxoIeFOPM9ybdvxGTsyD4vmEi
eKVFE5/rh73gUtEuo/UEQjmom2IY4eJWP17d4xNH7I7UyYQ+wLaeX4H4OYwQGxSb
/bdEkGluD8iVl2rxdtUb7nXUNavoiBrsJFz7D2Jwn1nNO36PihIXVPdsBue7mmKS
lI1qKpcoQfmGBpKpjcygLPQA2vRo62Hsy7lKmh3vzLqUIN+geJxBO50alMXMwqx8
zel0c8y5tju1jUMGPeZ09yxsnSR3ZfVBwaPDgwufIjNM/QqJCgqQI1H6512iHmwS
b81DmW7o9NCWKTI0oGaiZfozbInmqqHzjACRlv6T6oWHQjOacKujJYhDpjy2/OP+
vmEgONIyhS5PNLu98HBPRTNloeetkn5hstrStavwiNOXYPC4kPwy7PgooJM3fJMr
F4otLrQwZp1v6s4IztiHJfB6ZOpCORV1jy7W5hnRf6vRLKMoECOd2S/CsHTMu3hr
OInA5ftyBvYHIpTdV1Esi+2KHUFf7COUuGASPC/V6kVeSK8xRc0aJ2eoGpOMvlcP
oo2WNaDzHsgeEqJt3KvzDDYCNXxh3YpWgqf49XuabMvnJ6bX8E8B8fZul4Sw5q7i
BXW1au2nOcDruGyPWbfi8QnELT27gYBt2HLdsdPIWTsGNk4tbLT3SIgG8soOgxhC
yTQqiD05enCjMv/7kq001nTWyuOKAxNFFTCLlCr0W6ZJkBRTUwec0AWtVmdvKlQH
qO7D0Vxa5LD4LgTKxIJqcIj84jmdZFcIXuQfOwPex71EfrNuCHYyCTGvpJbms8a3
azFnN9wHchL7GEOqPzUt5yAX6FIc3RN5uwB+VAZpArxuE38pENVnalcq9G1z6TuJ
NwS89qxfN/hDffwIT1YGDGULzLDHj87TwaHxtduj+AAGSXpOVe0et7eT5DuvXtmK
btusTScR/3YDKFaS+k3rSJNOSNHOHqyF/nRf7f39/9LN0hv7iiupRxerFiF2n3os
OPUPghVwHe55MpDnhvZLIdGB8GAhP0xJ9qYW/cuS9XGkRGvPFqV3LiCZnyRgA8ir
ON+21V0l7f/5Odu5BYKeCN8WB9IfGvWmiSadfpnh08V67lmwjVJaRkJRb40Aft2s
1jNPGaz9ywuQ23HqKsXRjkrprIFa6tZohO7WLr6NbRoYEnpWBz9syQKO2SFbVwje
4k8LnnWSRvDHz7IIhxJfMxfTufyRaQHedn0vZaH1bSdMQrKW4qzEcrufa7pbqcBg
ROjYPCBhWChSv/UUg9Gt1ThLhAp2+siFp5Fg5sw1ybC8wWHI1BScZCEkUeauKdTw
ogYKu4ZKURiV770MotPemdGA253esZYqr5+ElyER75rcCADRkZy0gKdtX5ieacgw
xHemWbGj9qzU2uwlVFvCBvJ7/j7oGbvqu13BQMyxER15K6Rt0bOvGsGspUWMtIuk
E5rrH7yfg+wajsRRukzUB8Jp3rW58PEfhEJNNssn/o0ZVz871N8yteLso8D7ibTn
Y6BGWfZ83UXH4YGr6ZA36QHqq8pkgKyeFWIKWQ7vqhShcP40U03DeUEWKXkFoby6
pY3+cJlg11sQDsuztyfeNToFwvXiFlQK1yw2trZC4pUcMJ3CR0UBiEq4HryIqmd8
JxzudsQtJyjg+BTaIi0oNXL6A+3mlKXCOCElkPwLfucuQ/RquyR3QzbM6nyT9vSx
u7qSY7lPsfYoi0dLIZnx1yQCW7GCYdQcwMdWqtkM1VU6Wu6M9b7VPP3EQFho4IwL
U4jf+Wl6107s7iR1PUmJWIU3oGfdCxaq6AbuSxebCUlEhnSxjX/q3lf3TwXD23mM
qPkEATG0jg/DTLWX3a2mZ3JC4fVrJs++2vdL8MvL626fxKHdj2zDF4bqGxow4Fl0
3Od5cVm06rzJTD6gYGS5EWN86H7zSmJ02Ey8mh+5FQWR2Hcqf20TAvcVi5KcN0k+
IAuP3awtIJLxwc3KA24ObqvRZZN6crZoTkeLGA+zf2YsSh38T5H2nlpeoq+X35MD
eBARdXL7m/2Mbkskgyf8UFsti1oNiG2PlJpnnZORYXW0NA5UWFv8LAWRoAd+vrPU
6ea1PIKkXI9i+2aZTpz4afOGHcAaMuIxVZ4ihBviKCgeFBoVh1q1rRq08dpVhYaF
CzVSZLrJKdKv7XRXINriUk/N0EoOQqCJG3pdc0d8E8fBScsWHGdC9H0PybsXV1gd
h7RckEoS6VTS9PwQPNbsAUlDDjqDIV1KWUclWBshDKXoubszS79TvvlCssP9xgJS
KCwWU66ys84xTmqlqBsnV581bpJqBHW+8Ef1dA2khxTwZ/UzMpnvcmUCBiyARnM0
pWu7Cmokz8TXyI33SmxFik9Fwwvoh8c2AkyBR6O3jdQO+o7p/2XZLc4wGq7MD9KU
XVO9wQMPv69LD4J8soZJrLKGQCSDTcz/+GrJVodhQWB7RT9NCwwsXH+GWbQp6nJp
ioNWwXb30UpGWHtijP34ShaGyVVz7joL8Sy44hfVGZgWvfpqTRo9kzmsyWnZwkgg
a3bp7U9BHS3gb+a4TKsVzslFu1XdCsdKFEKdviChqjNzzv4itE4VjU3rUlcyUN4G
h1BJv8HkgWNfAMdtgjFLJhvcZFpAUWZ+qhnJEs0GyhnKg5aSTyPEs7v1DbO/zcjL
2HDTEUoCETf9ybX1Wt0SmQKrrDkl4MAQ3fj6s0AeLxMnG6634+snUix9eClJAGyY
jkYEIG0rsXV1/7UvNKJuM6Z9W/VU5smt+Lp9jAffGG4hOSBnn0LReO5mUm9udfjs
GKwcb21Oh74zRml4WNu0W6J0g1Py9Z1zep18JnNmHpkMgn6jv3sLMkmC05pHDwim
/xPVfrrMgxvbj/gdvwOygQ864L2yb3MQ+RHEbgCT7Qq234rH1bWq2vTjfYqzACiw
ccx/YV7glsGwvsjOv0r1ksaEg2rC1sZCk4PiwfGEQugv7KKGBAQU9z81kivwuCbd
52TTj+04vruzXpTBlMb2UslaKjxgf3jMqZHN3MJjTnLDlFFiIfoGweRJie7/Y4yQ
0/kDH+kd+BRPUzu4xdnAlcNxA5FIAblM0D7uxIE9N5mrYM7685Y+am/TzZFegyu/
aki8etaHP2EzZHQ2eneyk9UgWV6Z3UchTNOMdOvGpgT3zOhgHlWyIekzj4PVADeW
6WbeI85EiY4sPn/bONkWvMjouBNw2F2YI/Sny1Q9RVE+2mEZbBexDXEcuouXTs7e
MWMU3hVvZUmARGJDbPXU6vi+z64ptFRiZJ3c5cWcEXcDGG1ADRwTgDA7Z3gHltbq
Nhq9VycAjRpCyEufn5WnxUMqAzKCZ73y96ZYFYfY2HDpBWupzkOaQBoVjoxJY/sY
LdHhnY6GTcKW8e4i5LlIgL2WFhm6JlYQTnPVy7VB9CErfbKKIcU4b0416yemi+Il
HZmUoVkamxLFfCt93b9oBIYdROux46kQ7Ba+ka5YqnDDGVHf12agbLEjgZv4qCCb
w4C1XCk9ezwgVN/vAtepyFX7bylNgS13mOxYHdw1UdYAfin8etYr+LAD0ni9YDfY
Dt5lFfSGc8FVIsvFSyQQPLmMnazCvm07IzPYQkmU5h6LoSn/q0gGb+SVtWlg37Jl
wk1+lmrEgdP3nsq23fCrI538DgzMIudL7IUVnYxKT+WFRfuS1I0UoCoUV9pF/yDn
pMFJ6x1VIdaLv8x9EnGzO/FrRkPBBeKU6ueCuEtjnqOuLaBFEji3T6rFr/zuESRW
io2khal9AOQqLp5gf1UF23z08ctWOxuUHDxyuI+WlXouw/DZpgn5Q7bI9241y6bI
mTnW5p08Ir2X30vdVHYBOUmH8PEl8D79r1LKsnTSiVKLOcvX/khMIevB0TYECnEd
wuIYyU1ON2HMHlVL1NFs3IQ45pEUYune67PSA2qBoky6h9dKsJ9rWxqXlvEZd18Z
G3nACTrashsgnl1BXNffUzfFRCamhKHyCtoaJN/mAevImW/XyCiJcN8nBQHtKFkV
/7ivIGr+USWem5hjkKXdB018OMSVx6EDOyWcKhdm9wmclBUS4ak/ACFAzeSNFoPA
jVtp0dcn7WkxFJoyRL2g56ogg24ppl1Wl08fqs4oHV8oZW/lJCoeRajP8xA8cn0A
Fdfn+kYYo0wN/q8A713dnELN5zUr8IGlaIIP+JLTb6ceCiQs66ofCgHMlytZNKb/
1YVimkPBMfThV8GADBGGS4GxN4nTNb9QyL9GM16QhR/y0WZh4gZghxhviabvEvoH
J1ugtNTX9suWyxzkNTaYk6LExLs4fAiku5dpWieTiWTFD3LsI1exOLCoqxSqKePW
6lnRXiH6ISYtjtHFg+rJJfG/N+OBaGEaiOLH3m9opP0/sB6b4DRzl//Rqx0ITfso
O3PL0uUIZhti6wJ5ciZMKz856xi7JEEql7mSas2/J3ltBXSvGVjrWDUXtsOAyxn2
M4sYv6J3SVgEEyhnmK/RNby+BWXLdXQE3heEaNwurbzVY9kXlL4EnZr5TRmYTqMO
wltDjRWiqxoVgm3uVhsYuIemxTrhreYUMR+VZHBIFM0zpAJEF/h9D95JnuBG+I9t
cRnTDzBbXn2gzns2xn4L15Cgam+Vmfy+4Omg3BKYLlGbnYxkhK59I7Xt59LBFs8e
L8zjdKSUhmjTnJQnOCztZrFT5V+2ydHBg1Opug6s1XKDRwJNDAYx+HcmojAlyg67
wVnB5pQarKEjkhJIvyrHvviaDg0dwseCoc0wECxpBPM4OtOgwnabG6foUWrzsAFk
OGtau7cHfxPCQCLvtJzHm/+kP/FFhpqBT/4NR4ay6vTRM/CYd117PU82No06mrKI
nJ+3TIDehliO8WFqu5A9AK+QaqifI3syTi6uxktIB19eMgALSwbmVLzyeyb4Z+3F
K9B2g2ZAAAV59YY17o2prOlmUlytcVYaeElwPKV5AtXjV0VotGKPTHfzgW659ImG
o7a+UlgzNkcFKt8boJU3T95+cciUl5cBA97MQ2q0FuOf76vdr/8OWtnPmROpd3z4
+3UL+dclX2WOGQNKvAzc/uIpsCt55BIz4KIkGDqGRDxYvhWWIjtpHQP0roDPKTOM
QO99XCQIbRl2xum6lr4RtFg4PQH02gNdfx1QYLZBrcaP9ZhEhG2tj4c0d12z3Iue
Bd8OouTbmq5vwCfdqUsee6mdyIgVIzmkeorRHQrkPAMzT8Iq0aVv5jrliC7X7CcA
xEeV/Lc2R9nTxa0oyQhTRMSfNhaffNY3FC6L6vKxbTk9/DDsLKRz0yr49Nm9t4pK
b5PD+i4fbYK1fydtGtNJevzNlqBbVeIwrxyHCc8XHAw6lAwN2bjqxNJ4lXBPoAMd
MZXguBMIu/Fn7dPKtJbzarCjaer32kY6kjwaA11bYO5dZGqdIBU/vfsiP6MOTJa6
XmowIJWWmopEEyniYf2W+8UFNqmHxFLlYsvu/s6w9JOWkfrgaIyNkam1surIRBKn
/4+tRBmiPo0Et5NcFJMoI9OUq8Rc9jw0kAB45bkdtMK2SgW/vNNsDHManvraWfpG
p/Kwnp8YtLN7mjCsNVzMZ3ss6EbaPF5q2ALiX4xc/nHdPT8vDsD5iR23+qOov2Hy
b3PtbKMCZztwCvcsaDn3lZeDmoBMZ5Fjv9UpP+F2Kp7OGK5YsnwB3D9+2DJIbbwd
oNnprIcxQJe4fwoy2KnoYV9ZxkmuIy1/qWGXDUryXPQEOEz/yS4OpflT4ZFz8t63
B88Yl6FvArB5jVr9bg/IQSoLGU249d/YSxCPC/CXoRlr64jv4e9u1uXrnHRmLin5
cEOCdVvJCi4l2iTjZIfdqdqeZf9KpYTTFWFKvKwrrh+2sUxEjOO+Fw3H29ZTJIb5
x3Vyv/i6bM1v4qXLn8tRLBcyIb6TluohhyMx6oPpLXkUB3OzLV4WWciPYSC6sA0N
TyCUO6OCpJtJrCshEVvkwzlq2lIiduzdhKNReJgP2wBcFPSO5qqAKnAGDUeD+PAj
dLhqwftiu4F8q4++aMPRoEMPl8UCZ4B5yaliSesZ4d9EOU50Txs5UoN/2cKhUts+
9AM8D0YqH9Wvcw+k3vBzhn79zQYvmQJS7FclDbDXT6Us8kxrnEa1vO4acTde938J
0w2mn3X4eTsNluZtdFRpKDaX6wQ/jCT0BcvgP3+u6hVyPg7qDGD6d3tkBVApEhvc
XzMRneAFOQS+PeFkatHfO6+oBDUaDAV9FMemNeLU06o0PUh/H0Z66ntgCm63tJgu
HOgc3lIwK2+MbVp9KWjWBw34oGKWk5nIwhWOpw1PDvvlmyrzFry6PhHLGptlo3x+
OlUQNyhVUqEi+tZ15VSV9QrFHUIVd8LsXG785w8cwwaIam+9fhxG1EEYhO7hJX7+
9vkfc1b7PJkkEA/xiU75+NvbtWEx526AyGojopv75ouQYOzqRAsjUH6lGNo0oYxO
6fcRwivqzo+o+2X8WXwL0Co/bPOaXSSrPXQ9S5yhj8xSqWQvkP4BKFIBWQMlddNG
t9NKfEj4hE74IirN4UaevPyzwl9XrqyUgkO0XtnRaLxtSUfk0goHBjJXQo11YiIX
QkqkojByvJaWvBBLC1w/i3e1yd1cR6OEXfrQBagp+yHUGLbka+6Qe2zLDQ0E2E/u
KnJ8Kn5wnxChtBb7G1348TywBWrpSyWrExRW2AFuOuAmUjKG0A2gRfzT27MoUzR3
MEPqC8TUC2VkWdcIEphcmaZ60RgxkfM2e3SphlpzDy9MklkRqY5UwH7cEhPKUHc3
c3+PYEp3IS71XwxDWHXpPOl+Ir7VaglQ/LlIfXjR0n/m667lK2D/sau6gLTBqewi
g/WzdfOdOaYOrB9dzqWJbb8wRYyZMY8Yc3rq7yequFg3TB0LdkWyEEpkKbRbdbAS
Ja64Nr6S66ZiBeq1ls2NEpom7F5gGJsaqjrx5bYsNOS/sqx0Omdys301U60WSoum
bdRfmZa48yUmaw3VFInRFyPk6TEpKegrbVSg3a3NIbhZepG7LrdYjitCNwW5iMxL
rsC89JPN5hVIUI1txFk0TEajcUGEfrYYCnP7Wd32hEn29e7aReyzUCoMLmB+sKPP
y2fxgqiS4DDJ6c2PvZhgMo7cyMPrvXFCbZ1k/VcLM0EGkuiVJWO6MtiZG5R3bjHw
W3rJxEDYYehzc4YkG96LFss5wiBOSE4y1k949UWRlQb9qkzlEv8sf3C6YkjUvo8u
MhHc5aSJyjLMygkNFvQKwboKD1PX8DS3sU9/esWojHD9RW7ZHIFm3ZU2m1eR/Muq
se7ehZbcDx8NqkoC0ZYRNJfJ/LIfs2obYTUIK9AJwHN2Vj2NbgsfqRJPSiDed3MH
WR4ibAMRD2kISD19tTnLiLDQqoyrm91srk2Q97BKTvpFiGSSJvp6sgEaHgARugRQ
EPYRI3g8Z5OIh5QFNSSV9/AoKUpsBrg2j9Ohj0hBaAfBI968KCyPBetjx9Q5X2YN
2o88azJZK+zzj1+nXFxPNYlK/+5JU489UEif8ClvLcsqYaK9aulSQYFDdEltu3dw
5+FotVeHcqo7nsDHH1VRsI49mgIuLb1cYbCtg/4ERAdJAmMHR2pl45HDQpadLJxE
03VQ5hXKy9HJ+jAhKEJMYlg0AYbccZ60VnkJcdBo+kPVtz3i62zs5ztaNroVxs34
P0PLTylxQ/Vm7fC/qM568zda0zR+YW+IwWyKjnb9UfnMHPQKAr5CcP0r4DYHtLDT
RByYJpXUgDD6e2kV1CpvwTXAtn35ARrIdbVMY8YtI9D/y0lgeb+uFs+R9aal/a5z
J55Wre16ulOwvL4eFORN4J7/wCSjbup6iVTdN6QvhikZJ4lziTDq2D9hCIvswdlz
Dqba1eoI2MnxxMX6Gud+2xI5sKlui5fqe08+3NuGQ1k3mfBOTmx/kM1LtmSMI134
Tok5zavre12U+yXhaiIfkEjXl0g9RFjPjyawpOJjgQ9slNljucnUmotutGBpsxxz
9qej4UIGL8x/87m5X9tbbezdC+T/aAM4spYvvpzSrAArYR6ZJ7NP9SgGDhBwHvUa
FX6JroQ9Po8Q+JQ2yYkjkHAp9ID0KP8tNX8rUTc1jnvuz+DxdHIqRAYGs/NXVurH
KSIVoV76n+A5krTZcB5/R6o9ciZ01ugt4UnFPyv40uu+mquy8Vst1W079Ag5Ybdl
xSQvbBb5o8c5GwHz1D7GbrmIKpe7wF+7cRqCJKoXGx0L6gzES8Q7TBfN7W+iXhZP
P9o3kHaHBwXLg34kgMwiZjJR7Yo6lOuPKaM9mjf366Qa2Csx/4aNgomCJG8RLZoi
aJteVgrCMjxqmttlb8ggFVBl8K0LepsZUUjDKedRPxdE0u8k7MYU9lENzdhaTFjh
YLBpAqjInddDGeHQZo6WJindLmVeRIKDrZ/Sc15O/YpVnc1hJABrNOc5XSOAQ5W8
PcQ8apvkZf6YgzK/akT8fTiHRi2/v0GAuvcBYqDG7PwMU4uaTUmO8WrMU/dYXDH9
AN7oKf0vrgoLAmaV1kM0Qvbv/KIApvkoPnzP97cePZwVnvgWVfluxQzI8vnGKp7X
hF1mQWSj1I7R1w17pfAZLe+hvM6SJmZBeIfvBX8zQVCssTSjW9DY3MXRt6HkkHHt
xRmTrBMEIkQXU3z0VdGCAYnSJ7U+VupC3KkiNWxyRT+N4pD6SN8z/1S9GPFuJDpI
G1b6DLq7uOc+VMj4wiw3wJL6GB1/QbqmAdYeURnDXV5A6pBh05CPaNq/bOxKbzsw
c+2V9WkgQ8up99YHMDEOo8k0XxrEfIi4eTbfD7zpQ0oSqpU96IrGraGN1ewEG1j9
hfsu83j5VP/KuiKXAiKp/DKdzOM0FIK7BLgSGpoJqkoLhRwPaZDneKnlLl0Jybtv
xPyG2GyrPmNT8FVEnc0fERnb59R8Pug1ohJ3UbNc0II+K9htWTBMEjOFBeADmaH6
o3o1o9DZQ/ZBraKtF1hWrsSMW48Snkn9nx+0l6XkyQm/sYL/DVCoWE25lcmuTDzC
tdqSlbReidR7lj1+cSRV4oXYUFECJisH9AVFG67X0TOpuqtLUVll0GKa/Rv0hYw4
wp/M+ojV/lECkOL2ko5GmKjGOg6FxPkBYUx1qpm3x+xYi8S+Js//Ya0WJBG7REW+
rVU/SI+bCoIR02JYOBYNUJZ0jmbXUBzh2PeUHkgnVC7K9VPNgQE+/WCAKqdTJCBG
LfVg0dxfSN9/RnNEXF37sWEUR03bDKkOPb1b0okP2SEBa8ruCKqFQDjFm/0dyt7/
fq3f/cCwolLPeRGTPzHYHapIlo3zUq8YILnLZt18L2P0/GwJucrjrGlJn2sZshVH
heAZHw7FsLo4LQrwqjq5K/ZREyCVTqolDAfIz0/Y9UZy05/xVleBpgt4AFw8LJtK
CwpKhPzxYav0+JsmYdlAWM9rsvkuvwS+Dz0bm+ZQuk+ZL54/1iBFOJUBaCoNeWmw
DwmJk3wjh+85aYaf2hLLivHJ79i4r4MKeqHu6svZZntnu4AvZRSMdBYr1XGS7EH4
qk6egna1overN7MBwSJu03Mfxy1n+9FURjfTz8Fyurcz7r/fjAEFIQyCcD+FInaT
mgMnmCY3vWDIf1IEzurHIJVQnI5Q3CXqKf6F/NNJnSnPOjqlS1bPekp0UbAfZskN
zsT+YNljjTOtTIP3vERqpt8RlU5pH7jt4evaPlv4NmvbsakuMqGRkqJoY8DCFBEl
C1k5efW8Keu9FdobMgaR39U0we8VeQakyl9bXgToGrBPSpSJF/J4qGNvvMhpvOCX
izP0aLkiHe9jThRwESfizJ3VB4B+Qx5RcXyXLPgH/kihXXM5Ie76kAYLBOYta8EA
+L4CG21HB1jPP8bamXbuY6YnEGtVuEEOpLbUtQFwWkT/o3+n4yz5UcbjUfgi/Wmk
tj54x7Nzgm2qh6DcfVRM/92DTHHbAXLUOpeVy1kwNbUdIwVYKfMVBNLqv+BGvQEf
dckV/VvcypT4dskLKSqz7ium+fP6veimICbv1G0nnld56Z0MnZIDh19If+7CrGiY
4UwnIZaFg5THBaQrFl1GTvjr8SZlNl1DmbV9CNyICjS6OExsp6ZVEeaDwDULoJij
nNd0gMwMNdJ5XJUbpMIRJkXEXAYImPFw0h3Z8e57fFSBYcUqekDykrzyWHTXMLB2
mvH2cO5haBQj3W+pbaraq+Xl16cTYlKtcLsDC9hPtSoWCpBK32icXfjAZBCE9Fof
VFMLWrZcIkDAXAmOg9H3ycXKAK56YQN3nRBGcNE9yNppZoEOEj0q9uoalTUcfd/6
p9Fm/QE1zmws1vn03NKEaPQoT/mzhkVt/NoCthE4j9jvqVlBj+Rx3a1dXylFOEMY
GEyfAjygEH+ppW4wW69udinhW9tIkorwI2Z8aUrh92J9fXkkZjN9BlPHm7l9Gl1f
br6UZVJiOsem3gEcW4G8Pt+cBhSx9edYFLuPSDfxOKpwramU+OZbcUZvCRvb1zlY
OuEh1jLNb5NO36fkxWj4qeTIhpmS2Ig3nkmqCDwKJjYhDz5EPUPqhywtjrcb7L6b
dmm/BPsvJD1DZ5W6U95bmA8hxCWtza13+7xPwfydQbESft5V59Qs9z4E/nAPPO3w
eiRHn+300tWthlPDGwfFafYpz+a+R/PgQYneHISfBMwGZWOMt3NNhTirv78mLl15
qyaq8TvmRUKEV9ARsfazl68hOvyZgHhvyM1k7M5p9g66U7aJXGZkGw7EtbHZ9Njv
ZR0RVC2iGBlPTMHGXbmMALVGab+GpLdg1MGz0V++DRxZUTLu+TmXMYwsBVQ0dyUJ
vd6X2LGFmCxoaSOM62t8X3raBbBzwAH8k45Ydxa5EzePUDtqeY8LVV7i5IhTf+gO
arcO8D3UT+ZgRZ3xONDFOWpwFqiDlQVLvHpqZ9w28llV1nurJxxNiIBxi/vEEkyP
H43W0arrRJTwgwD8tdjpZV+2uqWUkOd8t/xuFQIdHEQpNoEEV7TeUO/wh21g/oow
DDJX42J6O1QZfapt/rusd/oHTCnX0p7pToqfpn82JjXUyjhPe4puSNowZr9BjvFF
hO56rcQU8hIAmZVCXmH8HHMGjSbrimEt6AMh2z2i/df3RbwyIyBu5rDZ9m2xz8D8
kt/BLYYfJk4/iUyoH03XeSX292wPKdN8xvZU7tMXuCWWvc8BYjPcrEjqYimq6A5f
OxQHfPea/rE12plttxJgJ+423P1KgneE4JutWf6lopzFn/66fRuZQhbf6wHpkg+L
HaFudNztCR2wP4ISGaeGeV3ThJnOOe/MXj7qoZ80x3dImeiazWzlnZcbKcfrSD3m
7RGb2APnpWEhjh+Pj4p59kyMtbUVZNuj5eulp1DnLYtDJkNbZ2xgMj34+nOKzuRy
raHwhFBhVfKWS0FaxQcPH9JC+JsCx6UiWykJ6m8CKVSA2becV7aOaX16VGQPCiRL
3I/8l7X+6U1lBB7H6ihkBaHxewZKAAksjpNXe6KGJGNJHA9mgbPsZtuK8biyOAAk
ztzE8yVOtEJNn2oHUNck880poC9xwZ4sA2yivUTu8RFfddevF2DeJ3bexYqwfj4G
BSaeigZy0vbWUI9JfkgYcIie8/ME0jvDKddTYMQhk2lBYBvmL3wzi2VCHjgpNOhY
aesLcNcY4zY6GtblLpH37+kZ6k1E40bJ4j+PEwktEGMDgFAjZyF2MjZ+ZEJsegIO
5B5Q8/ryg94HdnbFxAw42zIBFYm0+Wthmh7k4XhD/2diWvWmrwcq/rCQ++aqadc+
9DVGjsNeHxW9pIWWEmHHTspOdCXJzoU97VqxC01ogw37vkrAqhulJ7Y7y75WlBOS
Ax5i73YbkknU1rfXV5WXW1Fm618bj7HLxZVNvexAQCpko04iY/iGGA5AkWYuEjlL
FpfcR8s98DjeSakZywrZq5wMkIwhxfm2vQrtsI6inLgbuFJx3X8IIV8j4FDHgqEE
tGe/nGq9LQASq9SdUZCnBDDVc0eWidbuI5VI+UoqL8JKFk5tJvlx3JQ8YaQMoPuf
qXO/KjY4a0gi1MVBnnLeOAGVWaBtMpl0w+/yqN/Lmfo3aCMJF+LksGY6C+VkfZev
1tYxjAmbHX7Uh4kJnwekZ8d8ktVjTDFVgkz6oF7NcYN9UfU5Me4rlG3jfj3UMAOS
W4ZHFdj8DKm66eAnQwMhARwPoe0r0rXfzEj+vYpiLLOrkYKFUOyX/R+oPJrsawN7
ZY+vpboPw0zKjH69NAbe5heG5c9lwDAlbtAX5mx33e7Dr9jCegjrKpedqeZEgXhc
dbHidnEGLuMPhQq55sJommJk9Pqrh2Q+rUXMSbL8+Gp6m3Gl5NLwIaN0VL3Z8mQQ
ZgghVw2u5ObocAzw8rbUSi/71/CrFkzIcU+FKWo1nBSq6xYKVwQh0bakzaTxP0lR
H2t6j7lsbe5kSGuDTZ4UJGv3ruXyrkUbNjUcdOZFO79LXRGCIWKGorFP7vMZRJiN
vrvZv8TvCMwDiCPG3mh+yZhs+VlxwrePi551bPJWaZYkFGAMkk/Xz5rjxIA920nx
fXtdGSWha5muXteB5MH3dSl6n4lPRmNKwZnvWgQE2d+DoKFRiLPogYb1jDb9NK2Q
mDN/BhgGvWUwsRTuIhwsDn52xkczc6jaGfDuQuKgH/JGKNMg6CUzd93sMC/ftKaJ
QrEHLZpOUVtTaPHG7ZNQzo1JNiwXYdO01zGvvJKfJukFfDvH7UPhYemC7PWcC7ec
YAEiS+5lNeGAtRqObuHSfFYPwX1GsX6+XhELv3nc2veOPdIASwKDW4lwJz+VzsWe
diDpSd/vMGNXCZxZuMKCmCUMpJjlTa4BGMku38KBscoSvODiOFfyOoHk+9W1eEva
jWGJvatRJlFiT5EcPsvEx+WfwQ4gnZclm6dlWWhSAmyLfEsOFNsHiqSXHsD9C3tg
kFFPVSnuh5tpLAexKSQr/QcdUaB6fSbHBDdndkityEttPhh7EonU7SOUrK/xIw4a
iSfzwjie7GyiyqZQgYXvYdT9cCEtHwSuIOhIJzJft81DW6pI33tdxej1TBNt7cqZ
//o9wh8ahOD/6gsYYxYrdBv36SFyq1rmmMSfVE6AYqTISTPlFvitpexbu+o3wZVS
YLfagigDQ5/ZflMoOy2mQw+6I4T3yWncDEaR1QKTtqRlIDJnGf2CjdwRXuodZlqP
I1w6G8QGl1xck89UP0E0dNJuh9JvvhvTYxvbDw75OejImMNL0yYzUZi6qYJVYiTa
PllexjeSr7u7CowENXPbnTsqVz/bTzkzLiJMvPfE3Y/B3IE/ZdN8cgPyhN1gX3nD
XGG1JvTYb8gm7ym3HPPzrniMqzyEVl3Wk5dGW3u022NTxuGjO9PDbS9Dyh2Ai6p8
t19W9k6IhCdXSLWaFGGqtbo/pq5wl5FsAXKf6jXhsEURwamiKDxexCuOlUUlBJp1
DRtH18XRAw0cKohWiPN1onRNEh4FIlR9aYQO2LenHZ35mpDeEOCb0sf9GsVXQm2b
aLLlrEUlU74qrv3j3hz5BaHG+itfgoFT9jpeWumKo2libcrdUv4XLSg+/ruxNcrg
Ne6duhyHaEkSLVNDIyg889eOb1b2hnNgUq/TqL7/c4sioL3glrypUbG81OF1hwit
s7E2MimpAOv1qMxCnSehRjZahQc9pf5jIscDKDeVtQy94v4JfZ6AaQpLsinrmMrS
yjqGnJ0aVJI6Z89I4nZXcfuK2fncNyXQ4A7PPV+erUC70GPNBi+QlK1ObP/OQ+IW
0ck6RNRes0VM1KcoOyZ4siQoLgbzKhsnWVRHlrc82e89KB82YR04bOyYqHKUbBTJ
xRECppKtZh6/DQKiopiOhuNusG7VfkJCVi6nAYAYu79tMa+hf7MG64TsOBIp6cZ5
C8gZpCVsCEse2PGi93fmS82xflVa2J0tBZdiM4pbTDp/jnZXlb4O9AdWolOabyDG
tAZz0s10d12cCP26mQOEeeMFjAFfRVuaq6sevnRZMcqgbdA6QGyhVQp/652ATUc2
xnnJVqvnqIIuQQjiFIazerz7fHro68yiLRZHwyEzwzW7SnBzLaC7ecpxy+bM0NUM
HXKUG+m/xKfAv1+P0ZGiDiQWFzY2iqFOlZ9EmtrdlvD4+/8N+MpeDXWoKiNNLTvR
utPOgDu+FL1gMSRSenhqS+djUbNxRYNdhOLue5zRQKFTt8M5brNHod0uiLeEbM1i
I2JVad44+j3HU1lznXr3H5FI6FR3ajp7dPUc1bqAAbb/b2egc90fc9Q99MRQMnn5
i00OS1MnrzQq3yzg24wJdVYVFKXDxL8QBH0L5nJKiiFATwc0nPKmoNNGlwS2ERRn
0QbaHkYt9SsyVHk1IOGlh30rKOXvBOMaixsuZMUJ02nDxNl20XZUwCXcTBRqr1pX
ta4QUdnXHSTTqDmBhwo+Im739KeXBktZUWgtcTrfKw7MzUSY0ZvaYY6fn/7gxXJJ
FSkXuMfpjua5uL6QHtr+4XFNfJ/HaedSY+afvAaf+H669oYCmgvZd+jdM1Yx3kki
w1xpfB0GQEXcP6O+SISqopL7XVcRtaCO9+j4AAKLPoQLadiPeSK8Y7eKdY4RqlgW
P3BpOWb2xCnV9AE4UiozXxtvJFTXNV3ogi9mhotIH03DCJmwYZHM/gkJkm7Az+PO
zBNW3KsSs5IEcrBYDNg1SzEgRIOm9sRpQTuMP6PcJpeAlxjKPoZIT+3jyayA9Pmi
YC9VZ9Gp5HY4YgdbKM9AM60/wg0C8r213bVwQFzMhyvC7xQmKbGikhNMNBZnqmk6
JyocMwmQgcwH17mDVvMpfw9ZkVj21cHG14viyvxnDkO1SDEzNNWIyXYlybHMjGDA
/fi9IDNChbvRROv8lm7ODLvFx9CSuEy5oBfssUno3Mx01lsDjbH0V+A39IoccNGa
7cd1zrulw2VCKVAWWAtetl6NFJrG/HQW+rzMTl3XXhSZkz3jxG6RK4VTi1YxB6Bl
afqilbeQ44/2t5mglUvASOQUHOH34kto9EBcyMvTTQZgMCJe2jT0MB4Eud30r6xe
lnLGjp28L/P6DNjbUYnt8bfkKt8YRXevIyF1UddekDMZQIZ1pXEwa+gCCOlSekAB
/smDL/ygp+GA07r11ptkpK0eHRbaKNuJMskmP5rzc1I9UJiXL1fXKj1Dk0DWuPnY
UojIdRZ1o820ooK6aAuRfugtSIzr23Nm6KdI2aTh2w7XwIHKIbH9OqF2LXFIzaSe
RwMzSeK1+2mh0bScHXqSyp9r5vo1vJi330E+oGyzTBqgU8nEZLzszVlSDqiDd/J4
8whlEpx4T8wJhfC9Ci6m4D6QmB2hb9lvO+wdd0iSyGHdbqk9fvOYZBCOvoljrnmu
Ck+Xwze/qdeCvul+CyYpRfXKnZgHMVbxN8wNbIrW7Ev+xjyRjMdRlnnpvaKGa10y
LEsuSOqgMFlJgyodj1XiW1cydA48+h9BxEs8sbXV7+m1zu9OZcuwXOyv7jwcyTVL
4QfTuqAB2RE7MFyIVESYX5fc2ENEgj60yKPop4FnGmFbFGK0inIFsjePkAGsfpun
xw+n7zp7YZahoFQHkJnqSx+7838e8/mYtBIr+A2REXkiG4WGHsbj70euqi4FPKOw
EarlEXJSpVq5U0OTAu0raqPnbS3ny9dUrHNSooSe8e5bsgcNpr5Qo0z4yTIEZvf6
ifKgbwp++pI/oWS+T8IraugyKPoAtx/WftWF314cHVifbVGnQRVlqbiW/2tSgf/m
oEXDWppkJ6iDrfp5tahWI9fDwF4LpvmSS+aIPA4nABIjbhehAFsM5cFgj0V2iAYH
lcYULJRA+YAfMiLM0ZJUxN+U7sjnfYDg4AuJcPtsLq/bxxiiThDsDxXIWehsZtdQ
/LApMrGNjSgZjLarD9PkMgqOxfMPeKUKTnaRIJxr9T4ADOukhebJ9YRNGB4G7Jsd
VwngAv65FzFbi8wfQAXI5qZ3ppiaME1nGNPene2lcF0gBh1QHQOnFyf6i8uUrJ65
Ky6j8HvzQZF5HezNhqS35xNExWewsb9bONdyg8Bq0z46yd5NLq9eE93JHZbJdDL9
yLrNJDwG7+iqrB3CIDRW7bMJHbSfk9T0wTLWGx7cvKL324nIcH9cwYa+vThXKT5A
KzG32Mrtq4bVKmc7AtDcwdyFK5p5pQDv6bBNaF02uWN5vpMCbJZ7kXTGLCjvmGg/
cdPgAVuxAweYtWneW2zqSJeSXvN8lLS8W8HPvxMEaR3pBQickLhYFos8rIIj+FoU
/t3tkO6BNXZiCIZPK/60/KSvGdHNs5QLdwIULRvJP1fvPXO4M/nm4AI3SlHiFIhd
heM0sbE63qKfQZySjGQIHqs9d4ntZMYdp17TJ6PZdhgA00NclSYq6HugVR6C++uj
dFahKTbcgWHQUq3z43jf0uUqB8Nofdq65MTdd6HMiICx9qDzQB0g+e60MogPfEUs
GG9y/rIlvjobd2rQwFcKpta5r1MIZ/zHh9t7iAB9odNsNCP7nwTlgitLEOBD7HRL
22jYOH+3KHBWkmmCOHFfvcDFVFnJyR0cbcZulYibhDRvMIKYcR7/g0ph0fpNj4W6
5LH++I45v2LgbSWw2RYj1iC3XUoDYVPurP/4GXpOt3tLuF6du0KwWvrpLWi1zdOG
H3rz5FS1/KSfPFXPXFdQrBaZ2wuJh5yEj4/xW6EdiNb8uHDXerCBNV0wXVTDgAEX
VoC3S1azWC8nREMfwugwG3fMIs9LSBFVBpxLBFrYNtzxoyCTq6SSS5zJfElsvGiT
VCV4y/zVofQkOg4H26jhXOY+lBiANyHbOZHMUfmQw85HAcDqNFbCEyohIdjXag12
NNdy5g3RHCRoxQWv83w0Gp9FVI8l5YtYS+vWBYbUl5kLR+8ZAbSElIo9vlduMWZJ
Uk5dVP6nTNNXCrCkhG67kZE6xCWRLTFI6o1DMbPa2mbboyqdJibF0G2rszBMVtnY
no2K2bwHWxihQFwJ83eQhmoWCV3uhxLbushzioX94UGPoriSJTttSJs4AB7MMO6H
yAFbFUVLsSrcbyKb9pJ7GMffpZxzWYf+Og7lJM4FG8CzvGgDDs+m9M6x782f98NK
b+3XoKS+eJrdmrjl+OnNjBqm92VjryVWtpjsWH5A/esb6U5BGkq9ozM21MA0EjlP
BoUlVh8q6YbsKr2uyDYG6mO8ZO4Kdf0AQ2qNw3T9Y9HPmjZNeJZxJkCGxOVhOlN0
EWPb3IQoIDdkFZthmWOuF6bpK1ZmxTekrza6qK4Zxnnf0VBW3+sSUHC1wEjxcdP4
2jUdfMEhfrK+JiUfPHOysrt/QCO8XUeDjLoLJoLvT5+gfqSrL8uxEH9FbTk4Dynu
knzYrM+/hmHuwvb3U76JVa3cVvXNMY3qgU7rlD5wajb5jqZBo2IKqQ57+v7XATZS
OL70np9klo4UHh5C5jH6316cYqFny97bG09VMIP9HNXIrmqGbMU9x9UiG5YxU1eh
0CRjXMFHP6CHzjah/e+E5czbn61l49VGhSCBPfjwraVwATmjfXbIORtHTOALRa0p
MMB6O80tZiGyqzNAGEqPp4i+bNcPBgx4i2h4IvXkL/ZUQK1G0JUxx+2PnEOqFeN9
AtabEl7QAsrBeaDhuRX0n51JRAitp+FWx6dJMcgV29rnaYxa5OFNxzBMnfuHZrGf
FXeNwCAHLw9g+HSUXzXqRtS1CJET3oFzKvRf//ZrPY9B5fFCP9zGwDDSvUJnqum4
fWtpzp5VO8ogaFV0GLnNhRP3jyKz5UjVoXpBJBesHAj/dP9umWovyEJxF6PWAYIp
bemOywntKXfr27D3Q2sxbc27SicZhwM5w+JgJQX5SWDofhYiap6PQ4bSbI2tXJNH
ft6SWt0LmZ6d9G44iAJ6WbsYzXY90e9wuAM2dgR/T+4h1Wy9soS8v3A3wV0vBfCK
8UHBOhJwu1pCEEmdYObTBIi92WCJBuVCh58/uz2w2CMK7lPDUb0eFlakE97uxUF4
2Psa01R4jUtSNzG0RUpjLF6J8dw5KIsCsEHcbmWKV+yhFmfKpSEvD5aPqoILnilQ
tns+UQQm0PxsClXvx2mYDaJ3TV9raqjIai1VcVqkv9bCT0WOIYrIyj2BMkOeRj7O
iYEhqfZtVyZhIYqqkPpxD3fItecSK+KhwGfIRWpMBNX/0enK4edbXrRLt1bbJ+wP
9P/sEEKbPF5+l+Vf5ymo7Ie5xgaKC1uscWjhzmc9T0atJHYQm4z+2zHwjupLonnR
94lF/KUO0HMdcMoiICXjHs4b0TpXNntZsD25z0PGtBOplbhjInu7Mo4HMujOqffX
6ZkNJ5wLYDLri77iIPhMf378D+eUn1SLavaOlP/awMOGJUk4N8anQ2I+L2rqiYq5
P7++lPEFmD4O2OF30G6Ekq8aUKc4wOIvvdQDLI2vcCHa+Y7TS9m4MKx+fN+WHV2j
vnnQi0Xe7fwPIUaykhBMEJnbqFMTvQ0PPvRGlJaIjU2s2fkHuDBYcudB8xW7aI1I
5YOlzASUMpq98QbW5fzkf3F97TuykdUhHMW5c/4VBZ55/w/qGvrWUOmuNXD25YSs
r16Ua7A2+N8aWWYHL7ePcT9zuHp+/cTDmNvPvPWLkvOz6mV+Ra+6wx8Q+BFKJkQL
Ubnwc7QGpI+eh1lm6pe/m7RT7jY5HyoaQbsUZ3XjU5Leg6IBf1fQfw+zw7kjO0iq
ObTXdXPqvlc+3QDqDGvOMxdEciITPEYSkjlIu5NFta/YXFxYP7MzSbMMXu4Wo3cs
4ku4fOPAFVupkCvJOrTcZVfxOWU4v36I2xbK7gtcy2xb7IkyrejIlBeCU3PbUB0F
a7J8kdzq0G5bZ6nUZUqoZ6VeCueajeD4Y9a0GJI/xhKFZHCHrgJ7psu5+cPVXROr
f7IL1mBorDPhTUIhASLxSJ5R0ZysByd9e8d7/QTmXczS0c1VzE0y2kmq1YewCef8
F9u2AzBsXVWHec4CMeZI+XD1B9VlSTY5fu7nLa/qUWu9QZBXBwToHI/LujOeKw5i
K9JB4lxd9HuU061p+VmS7th17C8XmMUBnG5SXZA4vc6MZtM16UEMUiS81/XidgkE
j+rZD9ZcR2H3umcafYLqX9qTnE0jCaFr70q4RHXm+jJ4I2a4aLulUPqK2XG4LJpo
gKIESznz5UuKk5BqdHK/wcJqM2vypO3KnWI30mlbEd7mxVbyrue4U3rl1Ofxgg2h
WDenRMgTIk7r7FTThAo7GnaHnrGcQdqm9Gk7fmeieYg5JJQE8C84f043TgPlq1An
12BqMueuMEaPkzzzmWF7mVp3RfwcuIg18nTq0i7ypbpxpG+a2sMfDNRR0lTX49et
w3i5yNRFshqovQp/DTTRlk39lDpoHUJPPGeMVrCQXgKxLDI2vOYW8r4YKr6Kxc57
7SUFsjkY7qfR3aeFYlTPI6fkYbeEyorNkO3QX+d2adIbTu96iDOd6JtCYczHPJLV
foobQvbwYOPhn09CxGoO6jm2joS2+HI79pAeuyqXDdQN0FRwzwXsr9Ktbpu3PdaA
apsbJUvj567kiENcKtiMvOARdIbzTJ3juEcEIgVWzPNvvYEf3DVeNkLjP/RKyl1n
cUcao5cNr8NSMds+zvAhGtiKgLRMv9idWwMFLn28HoQD1msbXzErrBo0KrIFJSZ1
A/cifGTmfxQ6dUSujuMmY6JLHoJafS5ZNccYyod6i7MXoVpNWclY3VT+h0RKEcGm
RWO3+/EJR/qGXn+aGe+2YH5ybc4tywda+OCG0CYAsNJIScNW9haIvoJhRczf1Da+
7mdlE8BvR9WtRw28s71GsjFfMRlGm/Os8HlGyEAEQXcEkskSStULa6F3IJIQhkeL
HClMeJv/1QxZT6GanBi5eH/XtopjG5H4peeVjD4ms8Ul55jIkzVfDTLVVcf+J5JO
/RQf8cBiqKOdiREmoM/p3Z4UKlNJOHPWzdIcABz8zRlxZyRhRdOmL5X8KxrNqubr
gZz7q+9EjutF9y6fgd9RLp746t6zmQQKBcatn9uJND3tX2rucu11qY5ovFWFPA47
V31fpm+KbSeBjzJuh3hcIqi3MaLVYrXXdl4J9+STXLfYqpLrft6a7jmbqs8ZlN7o
YpMqo9/LWWO/Yzrs0fYul6yqcFe7VT7S8hlAnVxbTRfz8rXqi3jbMcunAC+gJbxs
SZp7NdqJcBHHFkmPZ7pFIgEZfCNM8vJ9XJQ4ODXlG64K9Ns5cxTFBu5v/+JLy8Zj
QAO5S2cE5Dqeb3klzHEnYZxa+nqiVbhs1WvMUJtNIkRpbfwQQlKwA7esJy6ijrmx
2fO2m0vbKxdmhxfUA8az+2piayMtDlxMuCpmRUx2XxZq+b/XBJ7VWYQEYHsgJCzR
Vvg/Aq7irM5FJicjy3ELwaM5LGlyVi9GG/vC7c9Sjcuolm1GBWl0fI5InrB455HU
/g1C3vEwIknUlDMy5NH5YJkxR/BAyyh7fVoM1QIw50TmyDaGf2fGife6HOaN+bzI
kl0f81fI5dSdlNFjjF12t4X4SvjXjlwqGlG55KlxeVzy/SyODtKHmVa20fwcCZsl
mJGbq6KxNHGI/dGKdri2iF8XvHsko9CON8SybBlqNSRg0iWGXM/aZEerqBV4qSRw
o4V3rzJvZk4LvUeN06Cuk3tiEfl3/B16SsZIRekelDykEjExlI3sIMwKxK+54f6w
73gKD59ePMNRqRUEhJzC9IBghpP8rMR9r34n18rnrT/HHGVt8HF468cBU/Vfv1iy
eFdXxsfIuOmp/TGOGlSqxG4SnO/FjWBk5PJ7MHBzoDqSBJDQX/HzVNoFqYRr3uDe
6x3szi27uraF6LvvCfeXFo36eTeaMV/2dpCn4+oa954zYVGcHNl2HAaZTC1NYypG
lYziknSkdMDE8VIj4s+mlXohxnSTDTXHLwT1XHMy1bxZbaLNcbvMoL/fdnwrI4ka
4Hb2dlT8aLdktwIMDMYAlouw5AYuI1wUc5u5iYk2a9wQXUMK2i+kZo5v0V5pNHVN
vysToGcuIAqjqeSCzKV5v1s4outhq7iKokVrB3ZOyHA6sTxn3l89EPNmm1keAeB+
59Oz+ysjFh/X+icP/TxvoFqagqKb15QCEMXrxzOfvKFyOmXjHwOut5qoqsK4tqUv
jD+VSbSwCagdk2Xfvg28GHpKR5KzZ6WP8QuDizGwNQbuMXVk4mNMEcq52mRC4WkJ
47+Axcz+ddulDmI4wPRKuMxWsVnKo1VrC74sp2XeHiAzUdVgZwDSziNxOwXzWmph
XVI43duzze8Qd48qiwo2vNwJanBWX/qIE/f+CH8Jz8bnQU8HDz10DgsvOS3LDjKl
fFmGA0V3MPcKvvkO1KFzbX+vWA7onTYCy+Y56gt7uMtTR26R2zTJQERNVIxdJqVR
oMigBDFikEsdDFlVAY4/ZUfD9QWiCi6iXmHkmGURSokNm2iHnDi84RpkYTMUT4lR
Qur/IH3tXTiO9dKGBZq2yC08UeHxdnpX1zTVGUBIV5Fb66g7wqI6nhsF3y+tztKl
Zn/tYGT63k2UzSnBoX2HQOWEEQbxcV57vyl622C8ZPTcx85GQwGnIm30iYzMYpAq
mL/yfTFCMIVgLGagzupNna9iSrm/54h1h62PqbS6gHtbKiXI+OMcLz7qIFr5pRqq
03J1qNVmdgbqrQOsYyWNbZ7V89tbipXueksxQRb/XEsieGIXquwJ8gC7/IcOqDyS
GaPs9DcbKGcL5M9LKMph7WBeZZVnpO+zdvfAGvj17rCWFa6uZgdKE51Lkqile73K
Bp6Es+nMIKBB+TYq+lOHDNU6iimpKaC+NVUu14FklWgly0+bgQ0lPCNm5OoDTmdt
8YL9tRhfD1/LubLVcRSadJyow0N2O2f/7SqwEjFpnNu4/esxq2eTq76lqC3zlL14
66YdY9Aqg7oiKOpxZwa/84Ols/mavKWAKghE6ustWgz5ycMJ43+3kTM4hFAl7UdJ
jMXj6yVPbLgB5i6A9rdEjftA/J3iOg+8vjRTpeq30NDCdPsEzITkcYfDr0Jokmi9
mSHkuwls4RTZsvK6tv7R1QslE4zXdrhTh07s5AaXEnnybYNGhKvFvFgB87wAlymO
Ffek59Gq4kQVT+M9QVYQimXAWOK0Z743qEQCRW7V2qN7D5nuOS3tH0Fe7BseaKcf
hueikA/9ObuhbfsC2SZR7ycdbv3tok8dcf80iSbvDvmS2QHv7v38Dc3pMKepAl3I
p6rl+rVb1pqAe0baPLActaa5Sa8KQF9oDIiHEC5MdA1L/FrNZiHvr5YceMjsKXL+
CZfSihJ35zMykY3r0zMs6Ca6kR7i4LTe5ZSiZ4C7C5/ohCoEvAkKDHkYg1dj/eZt
SS+UapWjIE0LQP+pvdOyNMyiuKpDHEtCGEk3DmQDrwZsmu+q2FB1MEeawJb7qxDx
3BMCXQWe+SBXU5K0fgxWQ954eeGLLHs20aIjeRBghNv9EZgu6r5F3vZRO2teL1Dk
oMJ/HxXJlkC5K7DQwzArxPxb6Z2uCiEWD0F9Fd99uPUUP78CW+HpGROi3515Gtc/
LrX5cTSBWy9ihaqqlG0H5PcZPk4cfP58uONyoCMgzQ95vwvm6AvgrmCWQlQZdfDm
JWUEvdmB6Gm/Df4SiWzDuGkz35DN0nblcSIPakb6uT3bDsaxKMYW/+mKcjo/kejR
ytNF1ECmPK1kB7v3/r6OaXR8I5XGvOdWaF0yxiCkmsIVpaDJ3GMkKIbkA3On/z5l
2MAsUAaScMb1Paj6J0GdZcVyk5g2EL+SHmW/SqROAiCc5+jJFgzsclyamexgt73I
QcijzVl4uIreMcM3Rq/RZ0zn4/OZ48HgiQg3Cy+qxq3rvrJzgrFt/6YYWC9oUXT4
tYEmYXyxrTKUKT7r4S8wV1kohCVItrOXcxeTZ/P3IOs5zgK9nETQMpoQvqjqRfVC
A4Ih35LPcnD93uqkHZ6z65tGKpYidVRznR7IY8wnloewD9URGSD6WhnbJnA+EyWp
9UWksx+jktQA9ajvT6y6ZgCBP1Linlx+22QHcHVoJ5hyTUsz8JEbji99Y0lPjHpr
FZFj463F24e33DoLvLriHbzE5lJ3NetA2hX7voQ9fpsg2KCQX8+9gWlo/OhX45pQ
iK+hXNZ2zIzjM2qx0iebY+oPdvFoxtcrIFdDZaOp/oTHkTPWI840uDTirbMnhXC1
FCzemMDjYixh7WSTVmppkvBQJ7ARrPr/PwuBxjfuBtAT36BIS2JajCrQ3SGQeThx
dT+WQTZXwFaVdIALvIQno4qAn6KeIymRH/CBGKOgI1a+gE1csVALMdHHDq9I0UAR
F0drH87dfiu/inYNx+otMjXyX5d2xOuQFofz24DkVM/tYueK+U22BW2yIid5lchu
cM1iYoMhBqrlMmMRBPo6aTynKfcEENakfOW0PSHh9r/wqG2/iIO/mxhBXSR+hPEv
YVJvRh1FK4hRd4Y/Dcs1S/oE+uAG3zsyAw0/Frvh5CV+hebdG0dWJyR+7jUa+bTg
HwRPqaZxAMi1q2R6WXkFRZIV/F7acm8iLz51/sURT+yLsbqy7xeljvASVS3HGVWs
UhaO5x9Po7bQwXFTPcLU6qOpywzPuWvtE7YZ+8VypfHhXWhXeEnssr2vW4qXeohW
6DC7GpqpGPAaMO6aJ9ZRdTPEAuOEb3z1kH4fbt4s1yMUZ8Gd8gGcNkUP+CZMozfA
wkEPvqSQdx1lIRHnodBXv+6dS2oDCiyyi+kKweDFAQIq5G8e47b1wL2b8IqvJEO/
oYSjrFDYMm8GrMhn5D4HdkjwiOGDsfmWfpyG6Pgoqk4ttIk+p+MZNX38T8gfygkb
mqA7FJzZn+1kyx57eUM+uW5vveqy0e0THQRgzIGumWgZ1xSW41wTOI08DQacgF9h
yNO+y+pb8NbMaFd+paNCCkebNSJ8AXpknb0y6jDbr4GeGahs0vBgdoX2/Tc1caQa
gEx3vmsnVBCc4HuTsHxd9vCnMcXwwLWOQEOBs9LrjGK6VVYouiUaAYkTL5SVTaDh
dInzb30WO8zMMqClXr4T/3EuFelLo9q75VEiY1NxXTZZPJxxxs6KIDKL8Ysi8sGG
WgkilKOkq14uFBQx93ghLl5Tqi6mZsqDPIpXq+3bAMcUZfspUwo+2ExCIjtXGUCv
RANCp5RG1XKJ0dLHZtKIowSKu0I8w21aehcQJQmkBQqyPqyvfZY2yCJBrzMbP76/
3F9w2EDIlVKFV88HjWPtMBAOILIfPwfQHQBVQGSybda/n2Cn0iUtL1yCBOO+mw+C
1ScMScSPOXQ9GDs4147k4UuoqRQbVxTyDj8xdz7ghx+1okT/GfWtrzYwWFFv+7v6
tuJaYFBqI3tJHp7s4BMArrmNBYtDv0VLxZFQKL5vE9DMV7DdNbMoQiosXFCZVbus
cT4ASZd9ec1qIt9WnzUhY8k3UiVjc9EEGgeqy6L0dGBjgW2RqfWlgPnQBhM+9FCU
7WtcCxyZJaZHMVvPBMik+Ja2zVBjDGNYGWQmuDJfpVolNmBiyrgsUIIFTj69r8Dw
DSuqOjSCFTOiuTyi/+Rtg/708FEDPPhXClROLN9CWuCqEnPSPcs4q2NVm3IukerW
9Ywwe7BIm2p8wzAxPD1Vzm1v/pxuywYggpUQgtatlQ9zNfxsNUcU8lkhRVB6c5d1
gOMEBz4a9NTkFstFRxj/0i/opqqjP5FszCA7GIAQ6oasIjgcSJlcw2xBlGYf2Gqf
2zBLU2gIwM38LU54xLX0qaWnN+usWp1bx2BE+3sA2iyYPUCJDFNSfOxhFLmp48nW
bNEsAlLHbxPL6WglQZX7HHB7EKdzD8PzzWWFhtT+VG5znhF+FENUc0+ToZR9bm9v
1IPitb2KfSJ6MLtfZjhV2IqTBIh3T4prqJyH5TdfUm9S6wLYjEIzwOTSW4wUQvZy
n9MFdm1HLeBLlYbDR6cDKg6LPggk6Ph+9rSPylfcZInRFiRmNCI3w7TM82Apkwjk
ma1i5WitqYnXxUaE1AX374T7MLIkxrBQqzS5z92LjCUqndKeZ25fDz4RVoSQuRvw
3SDY5/tJCsvW27Jz9ghy7JHQljvp0VDBygq5oNzTcUr4jD0bHeN+s3ziLxcIsml2
oRb5xSGQ+01HQVwQrCrld8SQDGh8ADDDnuoKNSoo8AtGgKaabdesCKOCbkGJWMWu
EUj8NzC3vV31wSHmCXdSch5B3X+FNoAiDtNiCMLFOl+C/Qu3LRXvArhUoQJkl2jW
atg75PcwaAhjwA1su7OzgJeyPtA1UhIH26GP/t+zmn2G5gnRlWbDigwqlZzCIopK
r85gc89FRRA7bTc/KxGZqJVOo0uO6khk/00Wv0GgGnuv7AU/yNNz99TMUVWY2R6H
3FONcycZIw8PWco0QN9vbYk/f7/RXooAJq+fpKc3+/zuuZWMzSqAkYPRwLPzqsCv
xbQxede+7Z5pJCOMYX5IfdkRfOtGvzUaK6VNO6PlL81k7PR6LNVgpC7i2swfv1JU
jEoX0dFVP/QlN29NidEOVFwBIpZHeXzgTU12CFcQ0U5p1C/YbeXcq0gBf77Ic9zZ
xKHcs06QP2KJV/lQtHfBI+gOU5MEPbFt5ZZSDNutDFguEvNFVelJi+cqg1oEuV0t
W+OnCc83bYh8esdE/ZY/cTOoxOW6dWlNR3KxRrJbE17/GqANRk0sTp4he9A+dO1D
i279y8iZ4UXvYfFxepQBvNiVW9A7AaP9aO+G6MyF0UIejeKOAWiFJaOfNR9z8Ya5
gKbAhPNTyDtiinkHjLKSSYSeiaUxYHWpM3LSEb+M4valUFMJb6I+HfWDnd5hSOP8
J8TJv6KgHp76OTD+1P3PM/TUNDexAMkcHRGkxF0/8V3PdzyQZ8AFNHPj1DJZEmkT
H3XrkWoU2XhfuM/0OxhI2kI3efGMZ/eg76SL4R8xTZSSQwkMeNsdcjAq7oQMV5Rx
fUE8kK+OQtV+b522Z/9UH3xiCXof5wpivg58gI0p54/sK+j2tSQJVQsZs7h9Glax
ijUmAHSsn6nAhugYv0yRG2Ohmb6yzA1Z5AUuFff98g9owHxbVug50a1CI+lz/Y+t
L9+TPBgVvscoGaR4aiNq7N0zAWy0bFGV1ds03js5jTn8LkhWVE5fg1E2ElxDWdxK
A9/IUJIfk+lYKOE/8eoOu7/Upaf3GlO05W3d/Eu23EOpgMjXx7n3+FKTJFQ5pyHc
YtEwmoHYkih61E0FGW5yhGzK24eUlJfFc0VqpEnWwVM2JRgE1QIzP/6vB6+XcWSF
jews/RxRfOkKar/6C4ZNSo4J+W4ZCzT+zid319VKIu0EEGlsu5Ba5V1VuGe6WGcF
96AYNMettC+KQupvX1q3K4/+f0SPqEbo8E8682KZVP8OE/HrbDZ6mjXsPKjHiqRl
RptUQa8K/FQFf7Ra0zo391CGcVtOm2BiQSi/YmTGIeL9GevCdKXkWSERXnaLJlm8
uBSTr0kILex9rWbNusWro2U8sKiuGrXS8hZOZOvR9gxd+ZiyhPY7gA4a4H4fK7nu
2o3+zRkqMnoiWBjbex4ShgxQXUPmJDC3Rva9MnpVqCxJEzgH32bAHLg56MNTFsD7
1rgBqKlNB49w/7DgmK4TijsDE2z6xJi+Gm5o0OOT3Y5Ut01qKI2lJrjMscs2+/Wl
n76f8O63o+Ql8CUxp0/yWKKgc/VPK6OTkb4u1o9o4JEAd79X2+34NIz45DMQTeys
qO1zuyLrtOCPggTo1rvAQdyuO50gAFllvGJBNUOxYb5E4Wvt4p9LZjLmUTKI+EyN
2LDQs0aKVWd19uciu6uLtzUCUl/c6TeHpZwk/xrvwC9i3PgKODRkNQtaxpHucMaK
stHBxqcVOdi4qC7D/DV7RucpdFOJeGB8K/4XtyQMVEyq2NZfwllzZo+p4vhhaSMW
Qa4CD+GH+R5ukm+/xrIzoWqHDfyJo2FVI9TNi1i8apQTD2+4NQ1RHXgDPcd3wpv8
dcThPApNLpqKAIv+c210YDeyJPOBHnh61kqPknTM9pWRGzw5jdgcij28R23sVBNw
i5UCcNaJ2KHnvw0TeN4ofQPzw5ibGuIa9aEFy3BVEYuiuWm65swLOqYhxoW/QoH2
usnXnKmJfMAvEUbA4kHT/QRRwMaTPtfkKQaQZJBILQg9FDv7Bk+3pvsdizxTQ0y+
5NqqII3baEMNZElp4jrTZrjvZKyqWsGy209Bmh7OIMYMYn33Yrv340iY4n88zrW3
ce2d+2mhX6OUjDrYYTVLvCrjT4SmKkmN5JVDNNViggsUWkHkhi1dI+hvgcBoeR3s
5ee+AvM3k4SjoB2L2Qu3pR1LlplxqPGP+Anegl6ydna99SROjzGNrV+UdBDFuZZA
HmLihLIoyyvg0BmJLM6dCBaRkNxaUTjvYGnUl/GZaKLgldSakxprZlq1beXTi2Qs
8uOARjzcJ2py+z1M4rvd2R9ZieGIqAUquoH+KM6sIDbwAkIxzVGe2FqJPzBtcgtL
4iuJaVf4yn8Gqqkyn5ofVsNz1PCDP6aXUDi4nE8Ma0HKmho3n5WChOtVwskmDXxi
6HCWto9umofA87yfCLyDJrok965doloty3VOM9dCPS1WWfqYaeHwyriM/QWtyNKe
13Pwzf9orG67ZYmFrQm414A0mdiCZ7L8+peWiHOCOxAeHgY+BWfB7RM35wrdlmoa
P22OEbFsn09H55+B6ngDOjLMQfF5jMKljF34gpsj6AqkHgbFMDTEEyVG4EWglA5o
wh24KAx9Iu57FrEOojgfDMz+ZAWj74GRyPbvQOdScACY2SX8soR0EdsGH32xHlPa
+/nTWO6QIhotDTasyDU3MsrWqnVX0ZxmBbgbDb/iLoxK+lNQ4vqx4YdYBQYpJiPF
0xhZI2VnL3y7m7nP1F8/6zZZ81nahYi22ZAB9Glxa37rI5KjPpOoRyN2tVhVJOq3
fDuiz5TVtAVi7YVuL5OaOSPQd17KhlXN9Gd0q9lUH5qhf5sGfnuk0GBbzcy02VFJ
sgKEHd4E1uxTB4CDo2DLwiSLEXzEVvnQDM6cE3HR1GJ/zvPjRC4cFzpzvWPrQYIg
rhtAtFmA5DZ8biMyonLrADrRCh1jcf44XyT8mbCY8JHVVPb6Td5hUXwGrDCV1SV3
On/J5gAgbkZDF4BSXtoHLm+QO2+wTCZqjeYWRKnyqFUScnEOqO8XbGeMmARYVvQZ
80SOPbtdGy4i4J8uYWTV91kWmQd/wb92m3mHyaTy6TH66sHyH6zKSYeQiko4RXQV
3B2yoF9ycSpWdHsNyTy9/3WYlEaeVGzN2dSeZIupSotmHmiJexe4fpmVV5L6j9Iv
qgO2QDm2IANApZYbF6+gq8j/tr+NXH41Xa4cPObizwefgCI67rROzz5nvMoyZ0Cf
1GqBxy1ev7sLC6OftHhNPwnUMiHAkhfiLR+knf9uaWFy6Y5rnMykjmXPgtSXJDRe
DRBvUbdWnQoIFGJUQ8SlZf37wmgln2DWwQ21zgulgJw3tst3MQi53dQiSIi/Xq5q
XxKDMwkfl+6FSphmwdpYTZQZFclEQE9vB9sdtqXucFHw4F3mTjD9TxTgejsi06C3
tbpETXobU3mcgosFhcshtrMCs3MrdLR9TysWxvYhQQzH3GOOtXVVrG+IRnbpW61a
NVsdwDv5IyY/lGzsJ5KTkCneLDLkFReMDU0nS2LITtoftsixq2H48y04ITe2kQrV
g8xXgZpinOAzuKD6b3y3I+rHkfqYwQDLvC7adMB7HEYBfGXTRNIL6+y8llzb8P5E
linWtPsH/xck5lMzQcTtjpzbXKfMVMeGciKO6x5hQt1meJ9zPw7OxgyeIsUUVqCo
ltHcH00Uf8I8TIqGRYbCqE2w1ouoHaze9FQWknjEKx7mDGDSLj7v8B7hxWLB2E3R
w4L7OD/5rWsUt19YijRYiS26EDd4mnDveREUMWj35mr9hJWJFBUA+6KRYqAcGTKP
t5Th6z/JA+Ve5OXdRkjTo77x/BU4krHuJkzZSGk9ufisS7R0Bd5qOG0t3Vrujqml
pvW/vRUKBGBZIZmCe7u/cO77yHGTbhbSZqS2A2zanJP5TGxZhPfw4FrJdyHOHKwq
WFUhxJa2rmJ/BV4RiZmyZ2HHALy3VHwGNV/bjLPvgzyUrn//c9URACTsERxxx4Zv
Ky6QSXR8nHd20yiwOOr57RpCxcM/bMyueJfkEX4d58DetXb0F7pqwRfOl5mXoMyF
rIt+bYoPAXCSZORRsOUp72FpRIE3DuyONyPJmh+F60ISOJVuxleYdEhfacP+df/m
mPClGtyjjuydfjTHcDUUCYiXnRC4Aw0zjbt/+HHIwv7IC28gkQv6KGOr7zhAofmD
BJFG3O47K4LvRXQD1QMF5mLs803tCoIq1giMp/B7Fzyu7rfE1z8LZ79f50G7Z983
2Hj4MUk4H7gBxkUbBe9JowLVf5em/bfNCI7aCzqOM6+0RIS3tT5LVY5MHbwSUCBX
3/YuAnAoAV77UtRXxLclNQRDXsJ3nJQE6sNTvJyjhQM1Up0STn/x3htcAoUZoBqF
0BteCJW9dmNUjuS/Zx1sKarf1B4pEOkiQdybrVab5EQ2q3o48kuEa70LTyCe5or1
JB+7p10hbOvrXwMCWXd8T00YbICtmV9u70VcX7b6J/3ZsJEPeqFQrrsfi3Ajr4LD
lX5LftUZpN3rmv1k4Jwp8JkQ9JMcQS5Lvffs4VL/aMJ01qpHuB+GoRcoyKWit05C
oiVaj8Ck621gvxrn53wZIcJofgfKRQsXfk5DC3UZ7o3L9LUm52hZOxBx5NNF7MiV
aUv+PejlKP1eYjBPFP8y+dnlX8xyxUlylj9T9BqG7pMNKYMh4YIsgXR7fDB27kQc
BAV1uRBsV3aCitSTI+Vu6rL+mA59JLG0iwYDr8jlugKXSElrHMhEvCIOBr0AWyoP
ye0BbhpOB/N8QATLVEyAd4lwdAhe3Ty0E1WGtBYRulEOg2cqP6PArVjktZLNDAHH
z+vEx2QYlevYUqqRBMEXyjLV2v9VhJb0mqSFQsFXh1SLNr1Q2OGz1uXqwMpGxFdj
4U1xWf0ulaP3SD61MlzVQIk1nAh1ozPgQSoxW6OWvnxoWGMMh6U1do8kyXQMrBM1
t0mhyDKf0IS2abDUUcWnPmrjbYDwotJINOvRN6cpnRx7Gwzd8kmCt0UNsaX94Yub
CY0dCNiM7eMZmkM4PxS54BcVCmzC7L17aWiZCnMdSkQ/Lu3Ro8cSnbEzcoKmsmi7
WNumH29dh4jgDVwVJh3DnoQuDjwfSZjgne8gtQ7u+ERXYrTJIpp1LPYM59dHBVtT
uBM0sYYC1mgH6lTDWca8KmcUZE8ObzgR9WXCNoaTuY0Ua1CwLsH8aRduGCtiDzsp
wPfn/HKFesP3vBWtEKFfklBlu48K0bHla/pAuWztAw/yiSPkIWcoUNeuhaBiKK4J
Ll664kmwPb5m5ApyVu5NlH+E7mO2lk6qRU8Nvc4PDVP9d0hsksa5V3vy7gHQ8GC4
rtTY9gBuHaxvV/efQQ043CUNxOCyubKddOkwL8FiQDfYMKzEvYnagG4QTe6Npgof
OJW7JDc+av1rThCvNTP2pkiuQB9pT2S65tTasq0NseEhDsMtKc9X6dBed9jE9lT2
7hM/R1uf/6M+t6tLqJSo84FHDEKcB6h60tzf2vVGzS3espF1Km9b3RRoZK0hX9WK
VCCrehMT+mSrsB1PjvMHMsLGvP7B5oupCc0vSR46WqsQFy5lrfPHpfQ8sklXvlzh
oq7NvWE1Wn3tcwg9vL+KybFEHy4JFzyPCrN4OR5cKaOiEtLKOnX4Px8owdOIkgt2
+xM3NLHDbO1nmLB2B+x/cRs6gkQRxfBCNIgw9iRvy2qaeaL9wJNRJbfBLnAJq5ig
f8y1HysTFPjx3gXc03awNKEqLDM9V2Cv637xtmgrswYKGXDtCBtX+RaFxdKDmqoW
b88q3tXljAztLG2MC7p9dCpTiJ0btAu3OGhqfeNP8XC8iCNFkCF65q+xPBn++b3Y
FJgUnRT1D4nxTRBlN4TpjvO0yYIWZ/3t/95y+K08PmxTClKlO5/EdlgFQ6FdLyf0
IyDKY29ymkNgE6P+LX8ksZczRT5+q8Oi01lXbtP5QbHDA96lH8IY1VSYBrIEN4tu
+bgPhfzBjt0a1kyxDlxdiPFmtTrlGIzj6Z29yKtUfFfiwNAIx7QrGfRPGOOtck/9
3j/gr+CQE47P2nAD3Xm9/5MmL4tTDAT/pGICNxb/9KtItBXRVlWISmb3QopvfU4Q
3ls/1X+JabMBGyDzoTsXuliuNosdabDar4ogVEYrrlzxRAwOuHrxlYwXQVdfQb2w
bYnB0youo2+jjcPB6aR2gP8uMzDsuTlaxnlAVmMj59o2IR2Hp0kym2mJi5qCaw4V
TotVyMWFiEgDO2j7bZwSOS1nqNsztAvrzGq9stkeKejrgEi2ZWEYrgUtBohtE+GH
oDKlnCRFBmgSkMwG0EFbN1aK402OkKM+AntXJbikepajClet3rD4LjUOnLYEIrgE
b8Hxh/pZNxW5F8gKXoIQxGEHUl41xfEFnW0UUO2KROSWKbzJVc39wwAyazuSIDtN
tni1NrZIOsDtZO7b58CSyYmCYBdTr+tkM8H34EONUHYzxyuTig6Jnm1dwDOnuGj0
tYnQTQTA1XtwCeLXyrHmnR+1u4E1LrjxqVHy2EoxQ/G7ws3WDz3COFWkMGkMiacW
5cpQEF8TNQxLAZdNVkI+fbMcx4ZOAJsOdxkeWjkbkd/at5cRFdkxoyb5K7I0ABDP
d/lUgiR7wKCkw0JcCpiEtXg+clmpT/pgDTCkSL2kj+woP8I9t65oeqhfKG8xdNdy
3tyKl41iyGGAqS8MbUUtZahDtI9CpjBUK9AlURaG281RhpRxiUdJY33RET7QJDYk
GOQ8PPXqTNgeWSp1J5C8LpwlEyvJCsNSoFx31tNOUexIyaoJjEBDJ07zEjvfPQYK
TkxHeo+Z/qqCkuBWI2KgFza90lPWHS31TAZR6Ln2G+XsyzYZ94gaYY4mUp9RJPcE
sKLsge/FrLlNXvGRib0XhrRhnZnWmdahJGwapB3yF+kKIkAcJQ9CwUB4oVzOxyr4
7S8zcACyOw2Uj7+ZvZiYJI7Id8MsEeZlt+uWO5nU54Dg9x3CgzAFJBJq9RO/SC84
v75LV2gUPHPmkAVsGGwnhxac3rYAm/nQjLJ/jrn24kDxYs89HWGGPAYxJa9jCNAv
WkScYyogqD8LlLXbNnL174Trs5fN2XvDptIHqvDw71vrgLamGF/7X4Rx8hmxIORr
D3XN5j/ACPfJgogNrd9IZkbY+QVwtz7SkxUKypthPJwJzQBBTrgTsvQCbbpsCmre
N0NSz3L7h6Mc6nl79cBBT1ZQ1cVD66iX0LK0tD0dZPvnV+YGgG6tsHfhviPVIutC
zoB4j4P+bkZATMM7+H26+kuZ2rcxizir9eD5t5fpzORv0G+ZXjnGBYXdKq7uEVrO
CXqpSIoULW1oMLAl+TRCFqVeg2oqPw7VBaoorrDtU0zUFEdJag1yOn6N0IpCNoFK
Vx9FtrNFxx68CQO5w3Jwa/3d9pa/DBaMtIMeUKE0P4Ai6qi5SFOKleuv3bMERkhM
VRBXhedY04IpIEBrSwRkEBZCRcxBxyC47oB5ueOIslLggl2+WXlGTiqyzoIRCCP7
YIDOOsjALJbL716rrwN6NpaP3wapfCKlg037vObV35KmyvQiryH5FQxSNEUGX+rN
BZ3Uk7cemW8NvTkjsUxCs7l/QEWWGS/9KdHokVMqjJORLmzuGPvYSkbGOzQHvBqT
f14Y3zxt4y+ZfX56Xpv1JiZlO9D34PvyqW5ScjPJu1IopNmcLFVeZN+2BjpBGsS9
89qNX8AJdcobtGv5BPWyxufdbxIMEEK0xNLFAvGe7uHIGeGFw97wEs1vUKNVj4zH
PdYCuhg+rZ8GYfWW8um0yaAoQH+G0T2pbjYJ3SjDjnOBmHSA4hWeaWaTFI8yBRy8
S9Y/LVdSCINYW6g2dcyhwyzRbOxuEsJeZ92sAB0qlervEnd3Y6XQZA+4qn4mQtfj
Wy2FPork06cWqQUHXVFqoTMAXjsgSNBmP5xCGjmrWL2R+7ZffVI4rDBSkER5DOy5
81NRwo11vZJiGkn7GxKPzvC4DvTqZguIOCm3719ecYAYj9zx/arfud/cEZz4eWG/
p6KvjZP13dH09TqRrcl7b9+7yrdpVk4QoKB+r7Ix4rml4YTJX4yqe5YZv/UcrgUg
m8zcdqbH1tzm+Z7sWFeYEy1o9+uWqkG8sQnlkurgfxVp12AJE0GBXV5/uscOzFGl
GXVkM/Qx6AU0Sq9jj5Xi9YqzVP7vuSEZfVFump8wrmor0WrbR8Yf/33PXn9+IZ30
/naqsFRlaE20ACIrNLNaLXKtVYJuqMe+sW7wjDDrmhk1feIHarxsZTo13HTiKN5X
7P01S7420Su2i1vWq7KOemKdjx2hjkqqK7bPFvf7o1exAL+3WgUzwxQ2acrm3KBJ
LU6HH/LqCcqQZGEs1COYwGewigHZVKvnDGL3YE3okrL+bdryD7nQI0jvMdpbtPSi
xqH+qVbnVH75YtBed50EKcM9ITEeZlklEGFigJNgyf+p1rjViqi77PClPOMNBdui
XT/iqfkdM+hn/O8xQ2pxPJ+Vb0L0BL2ClEbC1ElFjN4YLJR+a8mPkJ+cpLJpGsVT
5Q85TREXcDUkeD3/KXVXlYBgWZJxT8gfLbjdSSKKH5YQ2CQfqNIyTrd5HU392tuS
Qu4MBq+zuhFoSte9xsAyAGatPfrKpOjxrtWdyIXEyMDbIkTgKNhbsi1nIHhubs/2
ylfWixB8YZTE4XmZkFSCrPmMAV+JEO6VPe4HVFxqru5bz5jhS5B5Tu1sHdz8rlL2
9z4vNCuffSFY4oQ6BZIlh1knDv0hTntiMwSrOcAk5ceSw8o9sk1aMOKBjGL//jHS
I3BLlmqLiLZXWyLRv1rlTVp1OB5c9YR+RVpdUT7/XgpN9SxJJSuNITxJAy2XG8/O
8jcPdLYEcfNe2rx5gahgUJ/14MVLYaankuztZyuNoS0aPrqyOKUJZg20rzVYrxcM
fyHDvwpRIgA1t+AC+z350ukykU51klFe0JAoRwQ0i8UszPdhV8iwjevNueG4IVWo
sO5ZjHn2cPDg0KxoYw0pk+i5Zjj1GhkDV3iEGvZQxUDcfA13YK6CQos0IXQKtRWi
73EaWDMAt4woZ9DqvLb34CDGHCcmGg2g2RugjoOBBbsXa/1K0qxMxtFSl0gm/VPz
QE5a02gQtIjfr76f+dOEtDAW3vI4845I8Z3Q24rW8AUvmyruKN8oZYorzq/2hEoL
rZG8LwK6vq9lnpL66saTqCECEvcNHa3uURyWDklqzAP1BfrOlzu/yo7uHEaFae32
OpvwxRaOoKQ5IFyfKkf8dIgJ0GFgzwmNXiUrOnM266Y+ugpPZPkliEiEUZShjjNu
DUMBX5lAZQmLETIfEzb1BKaNZyjRnvsGo6hsVOQIt8ecQwGXVZs3q2KI4j3raMDn
5OwL1/z6nT/Bse0IcJLIneRDp3izPB0EhLJOUcDRApW0Z/Kltf4uVG1nP/WXER0u
hoO/rHUAZa0/AVmC3pVyXcBjq1BoMkTxMJydZeSYs5GSHZKaLFdka4mohiZ648Bc
R49ZlL/d9REO2gGvWo52i9ogPpgEJ2vBimi7VAPOLLrJCEs7fEYQ40FyWhnhJWEG
An8m9OLfS0mJziDb91K8//L8eQXTrrfzpu14/BwKofbsAqoING3jgF3JGIw2hQuU
+4QPS7VFk7Ba7q3TxBi+uftmYFKGudM8o0IhgFSxQS7elXTdbj4IlAMnAL2py7rN
kovTuaGTNry1ezruhE6FKOas+Vcaqu2p7l7rqNGjc3NRS89oGsYhGlTX0fHCELll
xGl5VZYAOXrQEr/h91l0PleUK/Mqn5ZJB2O0zQT1nH+eBEWriziMpG5hwt1ayF1H
i0Jk5U8/+o0pfO86SOSfGGNwvLCAXqWEyYO7W/Ct+hz35CZ788Ptv5TdOOqqKq8p
e5YXZX+85cts0oiD6vs0A4NvXHI9rXbiZ9FjSOsqKl28HRjcbiehfSIofdcBk5dz
oNrVc2pAIcDnKRjI/GTJGCp8y6QTJojA0hc69v2yH/j/taqmkx0FvtCqMjcIQOTw
gcxwCxkVyS2dBYGPK9rjOT123wiENL6wSRC8AZaXeI4txoXL3YWevYU91dxECOKA
I9vV8Q7CVKx0n3tEFeFub8YDRX9jSjpfulitEs7Z/2w9CKA0MCqyV8fQL6X/7R+o
ggsU1S2S/AOg0nbWHe+UTndAmBEXSk4T/aY4ny9VroAo5FztIa6EkSNnWv7g8M2g
pZKjrr1nVFoRq3CpqeyCKcPAMeczwA3xDHExVQLQ7jK5Ha05i9wS3/fvrM6LnvQp
pnZxTrrC5HKDNHPMTVqASI2ASgSd4iVXuU/56EnzRWeFS/1mNXHusOPlOPWThTur
Y3g4Z/v/LRanmKp2YKdurezyd2VeBGQ8//CijugeFwJhQm6iEFnJmxie53LCLzYp
ZbE7G+kzvD7MJSyeTF8HyyAPMtT1E7FznvfeiN4/lJgFGM0RB1VdcU3j8AozUh7t
KEfpzOD81RUzZMcR8lAwxbES7myWQs8tzoyud9+GP2yK/bWE6m0/zkBiZjL2GFH1
qFAsgjgxyh3UfWJ0I5Z3bXMZHws6F9N/zd3krliRLd928pOYqi5CeXbJorkk0X43
JyYOD0yhNICgalJKByVUudmqoPc83Ob899LkhQ/HJYBeUnbsR+tN+43+MbR8FQWK
0guFLAKcc3RkNMQoVWB8vUIjXQk09OgCtfRAtxRBfXUefloLH4AcsqHPpScjmrZV
id4a8wo7ldMUOVLiRZGFvrxBqMGoTcCRTFL33h80iWBUYtbW8+OsZUktPOgCvGUN
WA7R1cR9jL0QFCqgXNW5EA09dCjUH9GTRlwHce5mHVmPi2d4X4IRShyU+PzXMe+H
kCFJmkgEudR9BmmfIyif8kTeEJw99TLJ21+3np+F6sZn8X6GwaNocHT5CaNdU7v7
6+kRNW14b7nt93yFnOAaj7WHyLVpED0qfbvCBK8YdLb8ufZjMS5ShruGU215n66j
cVG/B7MN4pniDGQHEbYmKa0dEVweouLkt03rZMbIX/rmYydSmqQffgyEwaYpYHhY
0hV707PW+Xy9n0VsLGx8Yc5sR6lXqALYAd868YW/036jKSp4HFZIji3q1c9tawrZ
6aeY1EDvteTXd/+fTzyGJzgA4sr3DKwI5rlafIBUDbQDxgYknoT8iqFN6kwGAWfk
eE6WLKCC+A1undXvWa2A1nJV0hyVlUUUfBDtjtPa3/HaQuuqf4uABugUa/0A+V9j
daANDlL44lOR+8jnhe7+FcX5v0QZUkpzq6LFeNeKMvyYT5yEXBacClnV75PLGMbo
dSJ4adFtsMOzgV0UBYvAeN0MK0nOyRXfPRJ9WYPeahArQttf+qPGnSV14WnvIu74
+s2cebUsjy6p+jF/5ht9UngprFgTvoR5la2heuw7DVKxCvVEZKLdLAaV9Pb9UyiV
Ly3N3oKTLO1YnP1IIUWZoNfJ3FFsVWR3anVSb056FWDf16qGmaKlzdVtVi/XmsBC
alUwCBc546UK14oyP8CLWYF7PRRchL7YHGwSWvYTcsOqwkg0KlA1qKpuUh4AYMKD
j39AzfH7mbRJh/4XhnO9vSGZERCZTxEvgT63QGFbskGBVs7lO2+QqRhW2Gxi6r2H
JKHRE3CHWi7b+WqHoR8spswBE+dAbJ8L3R2B2Gp0mCT9eMrtE5jIN48Y4qXhV/IG
6xRCykLjW5NPeCYXoViIKBj7RCmB/Pv7QbFOeR1rfCtyK1rkfGR/YX+HSdj/hSmM
xmnKEWqMEy6lJZlJIEqYYMtAaz1QwK+DoMpNLh7/W3M/TRO/qnu0bil4GQy5N2FD
W7aHR/8DyqWLNBHOHMl0AffqgJXwyMzFETQzNbGdYZG0bCk5kCHv/hBOqk53UN4j
sOisIzIGwbjXKPRk91XrVu1rWehsMSaGCqhXs56z03/rV4ouaoexTK0lhmw6fw4G
Blsf2Bf70a6wqYN5W5iHfhp1+/ZQnz/CGx5ckZhf2VhsNIVyBAgydLFwb1Vm10+y
mF421kxntZIMR8OX/e05M0BeowPXDMcdJtGF2EAAMzkrMutc2HPnb0VVmA5sqJB8
msrosnH5QuRfG81leqi0uJ56giExyRFLeiJFWMr/6G3EP9npMpz+Be7lioCXb0eY
JaCgkSGbxpF/gygGcqZ2wa980nezlv1rnKdZsIJQPcedMb3rzYgHF+GMf5eQCdRK
opmiujKK5D9324rR1aSzr0PJqPQELUtPGO5ULTVlRLeIlVLN0CIQBrGdFuSF0q1L
ldo8HGUfdSo169EqqHy4G0OT/QSxY/T0ig0G3QJR+xJS1+Feh3dVUNNLdCFtbk9F
kk8D/ukJcz7T/QJ6itCNieUKAoFsqjPcTBd27dv+3Ish4wKXDbrElJPjsf3V7rVq
Dxq+yl7EtDwzhazhvVaToistuskaVYHiotgxkWxWCBRY4uslwb20pT/+qBbqD9KE
IQDESUpcuXxT5+KadntfBBGnZQeJe9jWGtjE0K0noPPMUh2dclWZBtrOxBql6Kl9
9pKcJX3nMZimXPphRf2LtfitLDK8Rq8OuiCxsiFA+VFqbLVUHnouGMeVgW8dCUP6
gGyp1agBucYRo6yrCF4MC67q/WWxMorJbwAl+lOJXAyxkwuy9vklL8uo7lBqh6GR
dtehJCCcT3NhE3Jst2z8HCKkoFTOQimGJaru8FatxsMHCfepFqG4e9InKY324x4g
E3CIis5K8LGllFbwghsvhwzBBHJeDxK8pWhmOCiPAV7svdFF+q+Fyovx96M3MWZ8
CjxiVuCPUx3a5Pw6Uz1j4Ek4axZeyZqogH8W9xj9UPej/cWc1aKAqdHXFw2S3UZ6
P2QzFBTb+/oHwBj50V93oRFveUqpmpNjJLANRl48H8TeDEh+wQzaEcvUikBSfE/R
qTCpcSH/FnmdoKpVCQWmcpjykxCsIplweTHZGCT0OEPk/dWp9PWfGwAj/Qs6t1Fx
dtD2zxoGbhyeGvPluPBy4IjhSkjCFa2SYJ4wC7m2oJwheW45pxLHJqd+jWQ5/5bv
kwmDBYP/almHtaskdnbwnuxA6TXHFL09c0I0EQLUFc9nzxNc9k7/KdZMjXtnPUpC
7iykDm8nxkWs5br6h+kYiFuveezc7SnBoJu5iIn7CPKh1h6Y7b6IXwOr0RvfOPfy
42mRhx2n5riARxW4vbJsyIVfUZ3ARROgjPPR9D3x0WqxA5wW/KSTWzGc7hjzi5Ld
N5X/EuKoX9QXcd8nmZXaRylwPccMF3cWdc+8jN07qN8Ia9A1Iz4PB3nnW3GeIIEF
tJqNyqaW9bepfKkzQ53WolRtNFBdcmKLELvlr1vW1ndjMR1EGalzdMDlhz0ru4bZ
e1QAdsrfmU4Q5kdTiV+jUdcwd1EjWC4d25RVdxcnglg8fo7RqEqPqXmEW+tFyeBO
ZolaGp778vEecKzCaBoFe0JASq6q1FgXDC6fSv0KBPmIv5tibtrB5HwW/4W+5kd5
tRDpfPidFoCqEl6M9eicafT8c/H1JdgoOmNpsjYm2i3xUSk9g3jrV5DIembeU1b6
Xf9Hz3/RvqC8KGYGy0zBf6Nw8cWyKWmAt2adkQuHgnYofAUNIWZG97skIuWBEwGg
2r71yBtCJYqVAtqNAsi8LGsJqaLEaX74XYWWk5gdl1+HAYsZCM+egIcY5Ncg2eGs
Yf0NSaCVyq0QXlKcx2fOQixM2U93P3BxZNDov90RyLpG8xX3qW0yERZafN8b7HjO
5LxeLef4DuvxDVI2INvC8qPjg3Rbbi/U4fYz+LwkEzVG6Xvokd0dvcUZoi8cJ0Zk
iQn2IipHlDjD9aPW5YaPh0esFaifwQ/zMNSC/qFS1YvRqxDS6DFEE2i5P2y31SIG
42aE/qTPFJ7WsfJcJsMo5yGYXEVlYR4hJHepfb3F/7AUZS4i286zsj20XV2D074o
1QOJyCtLbb8J7ZVxi4S1dI0bmMtOPoPW67foKeVtUWkP3JTbi8111fpYDJlK5ghk
XnIdX6YAESVAAI1jusLs8MhK4lpS7xljdoOGWyX3wPHdCxHrxfYP898oKqipdvjW
6JlHXErDufP/GCpNtbwYtbl2WoHiaET5gONL1rylFL42h4bTDX43mqlymgtyvXiR
sf9fS8n+5Len5pllWV4ulOEVzzh0+ImlCuQEeolnrEdT76w5Ne2rd2CtMvi2iJ74
7+u3CrJldfD8G41ZO8mGl8odFXVxkAX90/X6rKp+pcsdeH6RISvpuIIK047FOxSw
WQHgYQvrfEHKud3MYgEecR1XVnNvFCxvRVbXAQu8GFfCeGyDO0eyXQOXe6w4c888
s+zPP1nWJ0WIxfMmoKR6b8JpfIP+xloT6+J1DREyGoSBcSBlwccNbeawV1AEPJBl
5AhnnMMgwqztOZZzlbsvfQgYe4y1nbVYt+oWh2Xzg7FStxoHR4cDokwsIxnfrdtw
WvRdy/EMVZwhlKL8G48mUm+KrSldCUn9061HUz8Jw3sykTCt77VwKl2iqAbx8WEz
zLixCE86bXq0FeBrXUKCo1OktYFtmN81b3tDF4uYB6TlejBat1p30iC9myLzgVhL
L1CKTWHnZyOxYD+RwQFSEyjBypUc4fAuT+UER2IesgIwVDnlQESxNM/gDIVz2azX
3llQOp4Rkp2YuP2hjMwz2+TBtdWdhxTvdH5utiao54oizqA1IfK9YKRA65Me4FNA
+LlGBEJXCBsgj0Ll7x4NnxUlrxsX2mMskJRBL2fSJlFl0+F56quMQA1aR7F5N5BH
rjtAnTbKdS0eLv7b5FxzPXyr3antAO+90/fC6UA46eykXJHUvsHe62DcaWbOhzK4
NllAJmlobIun0P7Zp3Bs24iN+Wm5XWL+2KsiS17FU+zp86QAgsE6179WkGRDIU7h
sP50+xOMdQBUzSi9C2RaECe/jL989+devg81Wa4RIba7vYPg/iLseQ/tq4Ay53tg
YuQFcjlrjukStRGqrly8W6iI9Qhf0zn/2pssz0xFe0IAg9eUO6vpigJnm3Iut5Ef
3rwRRF522SYOxFInXFG4XlD4o/nbhJG/8qqpnOUuSkiHkf7wtIahjXg+t91Jn6d7
IlroTmB3hesHwVBXVsXsI+23kCZNS9AG6CKsDdUnFtM0YyDF690Cp2kOz4O9noIA
RiuUEDjWRo7NsBHqaEcXh4DrtDCXWoekcvIhzoq59R4pk5N2fi1+elEkwo4ThsNI
IjOTyFoWSdNS9em/3NlbqtudioqCvyxs3ItFacQwLjPzogGlgDIaBGw8T3rZX27r
ZItzfxnfe5S7PVzXCoR8SPeu4I4AYhAHFneT5JR5ZGX+ggeeAV7rZQF079veuuS/
vi0U3hDcyPeTpwDcHugVp07/Fb3IZcdnhUyMFqSdVnNKVFEcqVz5icwbE804NQK2
M2jy6YOwK3o9CinP5EvWmZcF8ssZk0bJYbbB5b1GWvGnGLo7bSYEgvYlDO22Y5hz
SqkF1lLC/NOSE18S4tuovvKNl1WB0sWi1vbdpaBBcvu7zM4/Emn3XSICXnWKx+B+
vE7PdGWZT9I690AB0pnea8+2lAUOVPL8vUVVgrmziA4BXTVhMQoXl/bWkbI0LI6P
c3gbNndljhDb1OqBiFG5hV39M1GiiI9oPaCHStL71bUhhJYusfHkyWcEfdI46LfP
S5cfWnfVqx2SqAgmuALf7JTQ7OoYdNe3pzEsnWW/D5okz0JlD3IuNciJlTeBIEqI
E5gfm6OxbhE5E5JEE6SBQKLGcN/xAzNv/auGqEe2TZVswTN8L+WVi+sMeKsEKCEX
81s7XZfMmbBFKD7Y68SIypivAZxPMVxNDjwA+R3Cp0SODhz9fAJhj1oiLO5PhFSB
tnmT+UZrF0RjhnKufY0/zGYXhZi7pbBh9nKV3i4dDfkGMzj5gZOryVM8WEHOD1UW
CoshY1gXw2feJ/+Xda7fgqwriZoF49MKRgNLrBRJ808/pYetxP/axRfNY2bxc5zn
aWRjc72AvFyUVXb7qnvU+OZpzXGofBXr8e6X2D2vPV2t9zPBXr2x8TXqypK2Sekw
qAfEaXf5wjQEG8uQ6cb7DRVEyF65YBTKmi6J89D2/2VNNhyn9KEFPZPH1fMfdEgj
G0NWh8NI4imz9oK2sQwe3urYNMMJMJZ07vEBMh0i/MsuTHoIkK7J9qngXmGshwZh
FNlPNAN1u/Xd6gj10Wjst4xyB70xGyDo+T5kQl03YowSsqkrWQ02fzJ7hQxM6JKr
1HoRvRn3iR5vN6D/NB/26+em8w53ZGyG3kwNVss0/zqhzksUcZNHNsMXxYFZw1LK
2j0aQskMb1BYzO40Qqg0WXebCSa1ICt6dGh6Bm/q5U52BWhndwke58lb4AOPoPgP
19A1Bqw4J8vccUjlsvXQPuilIbjjpBZtt8DlVkF13n183R/of7cLCyTWyZbS2Zzc
YLIwBQu3ZWv4M4nV+FEIskWjVdBxoP/KWN3ULIHi9HLoUKWCo4OPY69qdEYdYpzQ
bjARkdln6HC28JJg6fLTULXSxPc5zCwweay3mVGeBjuIqgMH7RVdiJlW6l7OatTa
qOHUXGdXc6a58Mxz+d80nak9pXIEyB7VEL7OvQXuiIXSXjYlYyyzzRcLHo1LDH1Z
h56tTwMtqyHBmnTLvIh/lWFTYB3floM2pw8JEGz+P4MkoSPVyfHJQvCcjKjOgR/w
SonjfZGCwX8XRAUBFodX3N3D2B4C+lhCwVielfixZifQdhvWB4N8V550EJdNz16q
5CXuV/wJRmssMC3meCQFQoN7OwW+LRVJHjPB6pLtHb7RN50hjSKVPZAzO48SI195
iDpVq+bWi/rL2DO8fCwaK3dnVvQQphiYPg5mpfptPpsdPl9yPBhE95dL/916a1aP
BpYYd5/UPGLfH06eta4tcTs9rMgvfINkx6vWqX8mDIv5WnHuJOhcg519/3bqkYrk
7x6koXWmLozgPfeBRZ6hL3oLWFn9WYI1LBY8LPk43Houkg8BaKnM+ufEHnDuZ98d
hm/jW/ikU6Vg1OaZr3ZxCdnXUkNLmKq5iK47CkZQe4r64F2GqylWnJnEYZSmVicZ
JGaNg2CK/V/5Hy3KQ2lTi5IJjhuRIxFEvn6OwnaMFTC+M2X98C8lamZb7unJSaZb
KwEWBK7C5swRmuTfl5/Tyx8q/U2gElXtjJwiV4Xao05nqUqNjOVK5LOiUliNbHn2
baSKrChuCdRoGbqeVSAy9tyiRC9hS0IGnyhjsTLPxtqQm4PFID1A9O4Uj6vMhblr
O1g3sA9/BBU8eZmpKRdYvl91dHI+TWXdIYbJWwW0u/67z5gFQXEvFXMWbJxKtoAH
3Ce14zoghAY7rUFTgeh7w9vCEXXve3w6L7PwSTDW/xwzOuxGn4i4LoFoXMxPiJWb
8yITtsI/RRZ7juBnJ4rwrHIKIzJkMPtF8H9or/3Hgl2JtoL+VAQpwLbekMiR34q2
S8nWsfT+Pk6zr/3+PsIVphzyMvDlIc2EC/auKvnynFZ6iWrhZmokSrOJ8+Az9FgB
OW47k38RrFzppyyC70l5QR4Q3JFQAWX4z+C0pFJy05422mAhVYrSqlAg97NgFRUa
1Kex0ph0DEatefcthofWvUmBWwwR5LM2kvpv4v/Z2xXtfyjUm6zNuHuPxaGWXYvm
57G1HuaQ+0uYZJqNSur6cWkDTXUZve9wxhAqCzU09tkgJE4/Dns2tXRwCfT70fb5
yTGKV5AuZ1tQta5W+LOERcLKaEJjvVUPVR+evqmUDYahbWuokctzvHlyd2hxxUpK
qovWOMbcI2RTZsklzny3znUmZx2USKoXZ/C7ajoTmcmcAwg3FMayE6Oh1d2bBRhY
o4bvU2X+tNp03I/6tazqeN0OROGa0av+gQIq9TYVp2haT/4dVB2EGbNaCG2oiifu
6Z6XZ2X9SnlITgIvRA+YI+VrSi/WUc2Pd0Qol0Kj9/epSNXzvLPWKuYOqGMIS8Dq
PB1hTJ/U4uzHx1xfGFYzZGyKrIuNBm7Q11TxBv7Ou8QW/EIRYMrEz9I+qg3m0aTa
J9N9EXQnMvO8CA+coW+qBD5vwyBIRV4XKcOFsRgB7DrWA4U3V+uCMra1wjc5GNvZ
5ZWdDEwC9dY6sNQ6HuhENWnRWFacNRHXvaMUIrJujWMYZQwhJ26RJpmQga6NH4No
0dZ2zlYzoNrUkIm68I/wAc+/PAOesmV5FuiLkG9gBCFxL3Jo5SEzPpFk4os+1JLQ
zOpi/5BIshhQDFEE1UbV3edG4zUK2ZK3Qw+e+8oK3YM+nh8KL+B2ZihLAB3pIBcn
yQx4+ddXci/A/lOXvzORITO9CEhflJjsSMCSofZQZIulEdCNbg2zvEjk1lQo5uhi
4mAA9FXYnrhbhsG8bdFoZ+AYHkkTDGOQtKsYP2e33zJ+3CvIVzgkNh/ixugA8z+C
68+LM98ZKhqmfKfvmXaVptQ3eSdNFCnXxSSYF+mMvoWGazytU5U1Nz5cuOrzjJCU
1dhfSY9FsY3LET/uc17++MIHkeMK3sFRBlCUTx0/uBgCQ2ekkm1dYW1pkpW8Z6f9
eK/0SjUsSUjLxjU7OOxn70MxH/4yR1e9Ed0PM73kgI8yj7xOOhevWXzHdD2oLb8d
rAZLzF9OkhpTZQPLlBJig82SyvHSlNuMSzmG35EhBVT2M4CWLe9QJJ3ysVAbvTS+
qscdONg3jDRL2K1mDxLChaedH7ZNVK3yNyAw8/dE7VMWRS2akpZ3fWkc2sABikrH
XviQviQsLB19qLJNdVf1Ows9oP7qHrc0uALa7G/60LU0yM9yEnWlXpKc/akxvu37
Y48gaWPJgafl3SgAJOnmyZuXX8bO2Bx6alwLIXhlJT3naKGoHhiU3vfy3vkGMG+X
112KBmfKjFVWFOOwIHcfHze95mRvIrxh4muFQT6GYITgKD5WJkkBomVnt7iLTNft
DA20TogsDk86fugHmirF1RjmN5DcCAUn63669cU9/dr/naYWOME2McQajfYPfTiV
w97+cRYkcbBbEVwMZwSwaYRg+ieQb9OuEnaVFTD5BZz6NgU1w+EiZT3nu4eODIDG
i0/ulFezpWPBsOUWfyxIjdIGqwgd3eREX8sSV4QUGMEQLveZEzfWaupZP+eWVNXl
xlK3uELg9a7Nfz7dxG2O57TL856qvV6Vm0HXQptAGiVSoLFi0vcVJPJdh7eNQPG7
l1OiCq/2X1Fvqjxijy9ftCI++LDF9ZFqQYtrtGD799uw3Vcwm1Ob2nPY9lxoGWrh
TpA0SmAOU5KrJRUN1FENWDLXKtTGt36PZttxKlvK2tWEQoMyF1ucbbHcqHxgirjY
eipUMJA6JRWgsikQTpDCBgvopBSjX3tzhKP3IEzzxgQEn8K0LWKWCHaAAUve/Rh3
6X1u+WYlVNNuYC4baA5X4Pl78nsjfZ9ghe5xkBaV9uVg+uA8LsCVordhn9YU0tp2
jlLJSVDKN5Buf1l1pNADeDDhnqd7ezlgTwJJ3KE6saLksDO5kyYWc1RJg+AV12Qp
clTT3dzLJqRzyxmC8luMOQu2E2qcm6refvb+Hnjxn1xvtQzb1HscKcYC8SruvbbX
0MmWjx6KKgZsLggR9vGXCDKPvR0Iih8+a+RjkCYXyVCnkUd36UdZx6ekqCnZi7h1
8FiX5hDWMUQYT02aoqiQQobXcbK0VvHJtKcShnfeVvItFCOGSBXvmxTiihkNdZrP
GR/EphORupjNa2FcN6ho983qj2OT6pckrUWKfnb/7z1CqDGqXcTmdjq2OVSKM6AK
xvY9IvbQNfV4FmpB47Mpvuf2jEqkUQvRcRiBneiikD5xGD2h/bnzUQhJcz/wDhLs
3BxkbAGqW3QM5BHs70yYHNwlSgbkoYiENCeAHKCja3ZPX664ny+MquwV8tjwRr8y
ZVffjO0HCG+kVmn2UbR5S22TS1s7lg63nG6PUF5gJj2kCHicCd55X0XJIrkIR9R5
oETLlfBr+EPqYFCAtYJ/+CCs1IfofrQZXiWteYl6uI1gpNzMJcjeO+X4emO8+G6e
t5FRdAHOt8pWR2CIIKgj2eRrma5nM2DXQH3uwZa48TFhqNNg3j/LvyTWVpKrse3K
NEtfwigHY/3OI3jPZdNjjkjUANR3VyqhAB08gNTdD74PN5HSWy5wVoIhXuXLu/4X
kbAfqxrQKezK12xNYlOVA5NYTZVmk8tXStOM2zQlOFky+UtwlNJZ1ow5JSRvz36d
fVOouYnBQ8q5+0YQrDNFYKtZKV1mcA9IzEksN+rRQ34S+7KtFls4+CpJARgReFqa
hg6MuZCOcQoDhR7TW0OYEOzXAvo2N1K3RRgGs6j+M/gQV2ePgftwhOBYRNW8c1EE
Bp+PNmjnC4sosc13DtdRV0zVoNd6qmTmexM59Uf+unNjI7HCipHCquzckwSUanFy
ujjh8FRBcL/mdpQI/qNTN6nRPsSIEbOukpPreWmdV0+6upSWcD+BoRli1BPl9dmm
FrSFVNzXVu87LppOp+ESseVYCSTGjQFzAtRQetcFHBT+4Hyupfn2nBAcEP+ztUj1
6YiYDhvRaDT1gmmXD5U0lmWdbeX+xpNDWnLfsgXZvTqt91RB2jel3RiIdiZiWS0a
YWS9andWdnsjQK4B3kramxaXAt9P+hv3weWQCCn+8NO/jhXsOZtxhG1UtmFgsTAh
tSUF0qptxkxgZGbDdnjH3qGcr/pvGLYlgEdpr/F8vQojBgOEOkBg1rVSk7ATVw2Y
VaKubaUVOky23T3PRtFexMQJSjlsiRZ/TvY/hEmJII4//0GuP2HWhhienNjPdDqV
Kyi0hL+Q3EKk6hKurPxoUmtBwHnJyKsHU3UiXFvLpKlhH1MOQKqXC3V98cypueBo
qJTE8ZOJm+RcqB3eFfOB9EDtzKbvweuRR6lsQ3GkOyWZgIwLfz6CeklYioMJ6etS
jy+1dAw2Wp0hTvXoz72+gBeRCMWsaxQ27taA8YkAKM8LIH34JLy6uE6i+KDQjc8f
L8LCH/mIYG4b0iWM679Kr+4a13tV6FX5CoYClNvjU+8VPTXbZk+LIEH8kr+tSztW
VnIxz1dr9tmY6glqfUhpr78zRou1wGZZzJkyau6g+t8GEaPeOHMX3Lu/dqQhbBsE
MA64/ECnJpDLtDnf/LNDlC8WlZiXzwH+gM/G/CdM6IdcyU09bG91vU5XiU9hBIRA
8GHWCgF0GR5sC/35hs+7fjaWJAWEiwadOUn9MEeaQfW+lJnopytO1T0pdy5mWnht
XT+CYynQcTu0LcXnJSRJLnwyyvzqtsUQGgACeutB8LeHNQ1XQS33ECsC1NfN7/mA
re8y3Z/cb3IkTMwbdO1z2RG1hsZh1BdbozwfWn8OmQg4Bx293ZSKdA+LLep88Abh
+LLWUW4OlIee07CHU+isIQFoyiHM7iopuLpqCWK7yyE9r3TPQ/KgjWX0qiglc9jt
TXoYIDYHZrmkO929BBRzeiXguUXR/Qs4HnGzVAuQRIsOBsQo/Kut0dLog5VxemRp
4kXBEb4jOA6RKCIzp8zLQT61G6mtbijcv/u0kIBulsiBygVxb1AilUyv0+3VDhBq
QOYPIpLHokKAiv308Lmxd3so/pcD6eemX5hihxXQrtfdHmoMy0jVFemmKSfBmS70
XPykvC4xh1deYblyR8wtqXi6omjrmcC7sPzl4aDWGG8N1v2Vq/qS5hkpEUgqvS0z
8kEvqHC6Rm5pVhRORfwy54MJZdAb+Z5IasA2NtmyrNOyqXulN2g5Xk10Vl21lyIS
A36AYjekScUwPQ6sRmarECI4cCA9ZUQX556lbmHbA0sXdjLUYStmREWFTWnnIkPK
EgfNHm9f2VxmxAuh58LQWyc9jLiy8WdwjXcLgZyJijYu78iffSIE2QSTwoqmjx5q
fK2M/hMBrjrzqLew1V4oo9l+ZvSjpHMM/XwcLm8+u2/9THAtaiDsBeFe5rfqQ+c6
3+pWB/i7tnYblPckhVLMiN5eg3LpGpjrb2awSPvoLrNLfJ017RLIH4hviMeVvoVG
4dpK+B9dwFg4SrNRFIk75mUrPfr9+/FvR8wh4I2s8Quec4ahA3hASVyWwtZGhXOn
ru0BpuVoSVXBsGb6DQTlzOnTGstj/hAtc57cgRifqcyNGs30SlrgILeaDN4kNXG1
C5OcmkotL8Ge14F9Xg0fPFaYhYkWo8swABUps/AE5KafsSsO5BN0a/9TqZdlO/IT
Yqkd4e5cJudx2yVOOZchYvho59Dc0/qeV85BjM2UUuzOTcrtw9fRbtOWAZUC1ETt
tshB6xY7KapOPPwR6HWHmChrQaKttQVGjCOYnqOMB1cqB1GY/9tnjPiIdlFe5B3E
YUwoTMQtGTY1FvpFUzuEHEs08fLW90eJf2EK22oOmZFoJiYmnbZqml5mtJCKo7bL
//ErcOkI2rsJGLo8KtlSZC/FVtKJOt+e51IUcvEJJYjxja5QA8uWFA4beF8oHkFj
sNGXutccwmBt9biCRkYjOHTlYycxzoKLZ8zEZew/BF3kRFLSCE6vyulXTyXy/n88
4+XAaPrIkxRw9IYphb2aElOzUzqDydX4lv9vEDJM/IFUc9fjlAwT8MNAPTDpUEqs
TyYnoiAPHUiMJF1uxnkj4SbnIJBj8BNQCQiQrFb03FJfALgd6upTiqk12NIXANpT
qHUu3+vb2ssTCGsV0TJU7nv3Le92dF54B2xuD+LyFeHnHynCO84Ivqf/5h1YtnyG
WkfNECPpkyrH+MNnUOD/MKH+Lvwp93pC3mIfCSwG97RZTvc6TduLw1dWqIzYL7Ge
CTKg3spU683XzBzAPY0my02K1bvj8EvCRJXCYGjIppCRoXv4CL9YLdvnK905+y2G
Ytnz6li3mEpf3L2cKwi6pFamXYkzjm9TtOrRhnc/4Qpzw6+nUj89t/y63Oel+TwR
g32Th4kQ39QFM15J+Y6XRXT6eHK0KSGSM6sa22Ne+LAtxemKrdjTiEyRgoCuK5O9
HZhRF1P7nvpu9FMOlTKoWxwtRyPbjxNAorHK43BgKWc2Y7PHF+VmYGcd/6mMHEGt
PdLBPqoYUPQfdidslwL0aTVXQPXtwxNtBt4M3JMWt1vvL13VaCSzLYWvMBCUAtEN
55j/pLV0JRXaHc89wT4wjfYfldbzSal6rBssKDsHMGN+QSZr0xj2T21MhoQ1xNt2
Fz89hbA8Apx5obDjZczTrRxgzPZ8HfzAIdLwDN21dV+68Ldy/7dCp8rpiDDpzycr
l91587celslKqF6NBpkwMCGV7FxVxKtvtAWqjynu3gqQpLs3KoI79YqtNEuvoVn6
LINGjvqd66dyVx5GJzdqBgmYVjq0n3jEeKW9zBHnZfHmGQ77ZaBEo4EQVbhyIPhk
1TONUN0earSHH55+ssksWI9bDSpTtm/xPR35KJDUJSBI0xzmVs9xFH+/WjMfdZCp
GvsFJwrwhBmFB7jRLOqy9vcLEmDHFGhoEH8Bdl1MJB87JaMN9q/3mvvBBpO3ShZP
Z7CqYs7qioiV/ZjmKnSOJlgxplK983CyvSTSHbMRcJ5eQZKwN3W2pbj3SX/CA2N+
/nsiZj/Y/C2z9zQ6hyzeKqj4jlKFKQB5YAJOORItNvni/6ADtTXDQLhDeFb5pfXK
kWB5bLk6KKGtWRyGQI3S/7FNQ6Lzi2+jK9qJfVXGvbAgVcyD7Y4wu5RIRKHs2Jyy
PoV9kxt7YbhRsERT/xHYhGO4PBX1rjwybbhfSYDfrS+pB9fAPVX8ABTKZ18APE+t
K5CGVVa3sP2CkUhkWYURiZT1sJkXPpoyjsb2ca5T1OjR+bJ7/BYaF7rmCzOE46LI
ti7fwvomaFY5my4Y77qzqku7YBTuFyQVsHKr0KVUVHUuMGHcyt6QQCYt+noB5mD0
8r0obFZWm1wL2oe5zJQAik+3E/l9iEzbiAaOJ7NBGnpbAeumXMCzxOIDR0QzWQQV
SEpX3mkVVSkroQYilc07B5AtFSQXH/yZa/WP1MBKZ75en6GRRkQQeqz2QavVBYVK
FCuwcOJXpDa/Zby/PTPWGDV91g91KvmAlEF7KXofoznepTtj62N2lyFxC1sd+u/C
BEGE6BqsYEKdMG4d6XJeuuIyTCFEltHtXqYx/PjvCJYesQJtqEhtj1ZNdgmWQAhF
mUUqLCG8ShpM+KZx04lrBgzsqBf753FQK7QHk/akUnXuRZ98MYhpgUaCzlfaKLeL
8/946Hg3cf5pkIhJdHJJ9y1JH3F/NJ2HrtALnl7tRGRebWz8AY5EUCEomRTbbAYb
791/BjwxF/jCCXp5gbTS+OU2ycQlg4q3TJMuo2XkxGK8koYeMAUdMm7dNHIc9SO6
6p6eL9fKgR7BYyfpQYAU5xbjYN3WUvwsmbs80KT1LpHz+xj51mjE0sXXjCTlUzWS
Uih8gQIRO3EtFlqoJ56jMEM51YC8rBPQl3KltxPxpSVHaVMJUw+rlTT5prX7+fw3
MegMPpg/+aaoiGP6px3qhckO3FgjCTQvQ1/pnE3fcazdlWMge6YXsCp13XOQ2Doj
TimERkLw8yk/MmLzxuGzcH7hgGY+Gy9ZYs9fjjIK8eDYqhc4jY2EhNSfJ3s8ey5X
aSxRYNL9Mw9VoyJP1CjW8CWRyUz+7q2ohx6peIcSiIX+XUuBHPmN+I/Do5wPwzpk
DxkTP2A5lMlMV+DZEQPo08Ax2dlXE5+QETdplXtwlBN+czwBqrMgC7KYQvmAybol
6A9XAsbWItpWz+ZSBzrq6PHGVe25D8HJ3WY9p8uEOQUGMT2zviw80qwvo1n+A5VC
fZ18wV7EexvD7U/Oji0v6mYMQ/OOxhHiUnjxlcZ/X0L2xOoLhXhGmlvRMzFQ6pvg
Q0Q++jceTL6kZUkqcCD+K1E70LOyP/FQqThpom8BGEeZsyD1HXBQJl5rOBrfSVxq
gvi0DMfwECSta7VliaxY0CCUOiIwDn5ogGldLBGw/U3vPaPM37TORTmv2Tt6icwk
laNAILXlJZElLFcYLp70AXSTAFmKAqx7eK6uIOYaHceuv1asWxkLQc+QS6OPuc/v
Qt9brdZBApTVSow/Jn7pXl4fGQrcuSDyGGgA4IO7uMJIO8XII7rsf80wP5nMExQY
c4NtIfEm2jULzUYPu8YpFakRfR24T4iuidglXPtP1OO9+Ttu5zRaVdNEI3VzOq27
gDfBmdYBOyRR2XwRmSJF/2At6shw6boGcFKaC98X0vN4/DwpYVQH74jrWeqiXj7p
sZMNwdZHydg0MIrimxA8iWhFI3zNroUyoxuQX3rS0KHyX1yab14EXWoiElkSdbim
b2FhXSjd1uHALTA/e5MSA8pxHNJMWrSpJFudF7q3Tx27RcO7G7VUcyjBNUNUggyv
cm73LUG7pkQLIMWHcw6oLEMj+bTRloQjp9cIRI56XOg0pLWD3uX3Q1l1wG1rqTFS
U8sO1l3RIWFSVgPSRw0JN7/a7rXmZ7oVC7YfWoDIi2iGK03o7i66IVGpXxjB2jqf
It9WO1G14iu10c8rrvOtFChz15HfbOqGhhwGjS9/uoagp0lHHIMonZvMyvRSyPVo
2Vzz2fSM8Lx4828NhpIV+ntgxd2u+ie1v5sqgKymV3qn+9+X7/ZZJtkLquO4D6f8
3vztBi1YAUc6sHWS3mMezHAKsitam5aZi+patHqBhLG/ZpgtDnulwS6g8wg6hlu1
O26b7wapuQaGvsQCRPJkrwba5ijSKPSLJFk9cDBCk/69wihNBRXlMntKmXw3nSg5
wtDmKesB2KLWwey/Fs+JuRswiQgsuWXRMcBs+SS6lKNis3beFDFdqmdsfXkW63Hq
GAmAMbRCqqEhPZDP6UVEaSksNstkxie/5CEmXSPo/iUNtnjz7vT5//s1aFaFMfLW
6o1eA1S5+mcMlND5YVSDJFVgoxOaA4PjmwmDq+JKm/gkOGNYNg4wLBME7mQ0eEMG
Crf5LG5kHen8PYDcKLxLzXiSh7tBPro9cESVHvf67gp9HMYMp1maDDZgbeI7V6ek
m7JOQa49y8pcl9jwCF+Hiu8mGLWwDO6PR1KeQENusO4drhQXU50bRw3sdgRb/M04
iNUoJvE6CkJJA7m2hmg0YOuZOppROJJFGHpeOdI3y9spyQL7mGl+mfc1N7vPLW+F
bjxgZxH+BB7Hw/7Tm2FcIDVvp/Lw0Yuy2MEA2ncsKBqWRcsHJ7gccEhz6FZ2b/r4
z3Xk+oTBO1KJ24ngUhoAQgv2msIeAQmJD56+1RpjrgOxD2VjCCQGVYdo1wHDAD3+
b8tnZHBGFB+Gz9NZKfxSOc4zkZUzXNFc1QRgm1OTyOYFt/tfZVJifno9lLaiCcv4
z/Nd6lXD8kFe5eYh00Au9HUcBg3l+FJjmS5hk7RYafMt99fR68ZG9rHBCQZoksIQ
SPNVhjPD/kSSD45nEuTMo91SKNHAehLux7/VAhkSFUUx+VjqdmfnJOgCQeF2tEP1
Oq+x5slBTcKyFA/+T8bhSk6QHstzu0h8X0EgHLKEabEq6Fb1eS7PMCOs8fPxGN6i
b5DB2v4fzOhDix9+DK71zWHQn+1+a3rdDEoZ6b6UEHQDHEo+h/sexAmIn+0xi0Gu
ekmfk3dco2LmrX1Me0+kCFejV8x6HvOdPtlTCsgj7frtraYqjkk63Dm5EvHXuT6t
04U6kHdxTS7Ezo+bf9V1TwofAZ5o+F6Yk2sprfXww1BYXUnowShCTnsmDAmR6Qfi
RoKXwlqpyhhmyiN5DANz7YBtRKtX6o6+kfrWAtoD0UIYOKQ5Ddkt9/+INH1hed9F
BnZfaHici5GVhLUpBQw1pO3KNfSDtwU0VPpj33vlXLdNIBDWkPNaPaUxEuJUN/M/
yK8A2uGS3nLWRymujQGQh3NL8uk1vww6YDK1Nv39v0k0/jvLyMF3NnLCrZyl6owc
xucpgBaM54FkTq6Ws3lTMHUK9RCdjRhu/scIH4YusUYhsVo0JCT272ZunQuxJ2pg
6U5MiqzSY8CVxAjQVVVXRxoK2lHh0RvJG1QQtxbYOwTjxviY44Vb8hAp0q9RTC34
sbRrKVBCAv1K/VSFEzDlUiTgyFJDEBtPpBFdHYQJm5lZlDnD6jnX9XRSLZ4ybMNi
52KiSotPtOW5fCnS10vO77qOYyQ+dqw62YXX0DYxbDYWo55JawHN8/o6NcOkNmbz
0YIkaT6oa+KWxM0HgAHIyEDHLcezcV1cgFiyPsZ52qYiJhqIeZrlD8ViSfg9+kws
y8cuou6hHbZEyQj/65N6NDylno+DchdkPzg4ozMqbggK3ofU658fugPkNXv+97+O
+bxf9dNNpirKAHIhz/oxcdB+xJs5SmqJY3hfsUjt+gnfZzt+Voe1yKVQSmJZzbas
WEZkSdCzfZSo4d7gTevUOdtPXywvcBq6HxYdneAIfk8zs/TNRYchDSWT77pPMdvT
9KmSQ735VvHTp0q43Zewm1760q+l7kwK/1/oqwaPIbZvJjFiGBdvNvJjjD4bWzhC
OOxkw2EZFKKkJvIG3nGT1Nzkb3slk3B2K1Cq3UOYwkMewFSRQoGrzJ4ZNWvpGk6I
7jRodjIvPY/d3vMwcvw7Di+BixlBxzimBok7vI0BqZ4S6AvWEPA8xoI3LYoPr3n+
lXwfnliZV6iSSa1eJIo5PVe27tHA+DUrKyWUtMs5ICMCnbLgeKE84/7CG4elObdB
lXiRgdkvFzBqZeA8QdUW4uH1nAz/r/BpCAVHgnWJKGLCrcAxgvVOO+eda8PCs4HE
cwdpZPS0SDK5XYDngxk0iAt51xjEqg/LZZzuWXraluAUAzPkh+TymTjhqWJuNNGR
6Z1X+YmShwJ9z/kTJRicoyPDwl9T9I8um7Nzq38B7eNkny9pvFzJXvvWESlLPgTc
y1JlNzFksiDmqq517tksTIgebtNkvTs9kXpcCRt1vClit/LAq+DVhI+Axij6YBIu
b/Gs4KDXQRWOoMV2WlqH8gmJztDiY6xZrGHam+yefkeTdzhHeEyxtdWyk6OLo8t6
6VTu96MjHDLj/alz9LMgTpOWWcvA1KB0AgVct0Ui1mTIBY1lkuu/lNyZesgHCQHd
xgCd5cN5YRcVPXeKxr2tkMeLC4MA+rBeCP+eg/gJonDjemnLZrU9LrB06igpnIYv
pQRaNoxpCG77LKlBEe/P6M9+6jKa3KgORB5qmIOWpz1ucNjRcjTEG6zbRC3TTdC5
YidUChJv6drhC3WIVBDjtlDIA/NUmkQjjYTNfJgJ/0Moputpk86ug34YpYzt05GQ
y0Wzm9Lof7HfHX3rdVwbxHXDLyntA/xVhDzmel9mgFaeg14CF4dstvON9WpfXFf8
H5bNWG3xm82PLGAvjjnH4qCTFSUQir9VGs1T2tL2Z7eXjsbbyfsFvQkBqtEse4RW
jzX0Jez9OqJS7UYXQqtcobKZ6wwM+gsLI0U42rgstXo+GwoPAg8zTk5cLnes2s8/
BzpCZj3piuzioFyAMBOscSEJ090N+6JHDd81HWxLdT1v8VTKkgzL/U40Dm77emYO
veCXx89ucNqknYH5Te8ufbD5C6oBvR3YYZHRTkGkK+mmtrU4X1TiXaoQpOcKcyG0
xATgJXQYPKPTOugdWb2GNx4RBQdu/HABPnidlH2S8oLwcKiE9ev0h4sE9+sFDqgV
nLSRNuDdgWdekUHmsnnXyun/nXcUhU42MOEeO2zKQ4E6t+JLjld6VzMTwbgG+7L0
Y+w5OB95nRPecwjiy39jS/DGWs5l4MN7E457XmzmNfKnJIEWf5WHwcZYJUod/yq6
FG8l09I79kuW4qm3d+9g1i6DKlzqBG01kOiHneVp+DmoLybWy74UCNwwgxDLckCb
D7DVDxjIC0vMe1QHqj+IOfm/f0QK3b/0B9inQFbXpGOd3qKHsQR70JFgLO1TlGV4
AO1ixIWErOe3ftXZnD8XHkgOcrab1t0qHTbVHux4cfTogO0dgqBvwf9qCyl531VX
VOlQH7313KV2Wz8GfKzHCJcX86DkD5FbeJPYIk6piG5YJlYUnMgsx7HJGuwUhrUv
yPe7ZdYWOsDdKMKNqqX2Y4TnTUoXLpMimdbosOAhiwzu0FFpqv+CLfRRg0y1nNmO
ViYqR+SwShGZRlpdQ6kQVikKP9w/HBD6LHqhGZeTwzNMNIn+mI6w7rrUkAf18wVG
EvN5++lMr/aFdipsvs49YHHwHSZizDAiKwZz3T1jyz8ZgaNBOdtTt85kkB6ioHHs
DKv+pysDmd2M2usWD1ozqahvfH9SsG6eXLraE7v2PHcocAqiuHGKIOtTae4XH5VE
bUv1JiCgbTDTwGAgABF+NR1xW9n9svvxU9TWkQFM6oS2GA6g38XNLBNBEEGiI5TD
pKg9MxarGmPZidCKM9XFuv5onwsRy+G+XBOb/OtIxp+ZcjgcrwXg2rywblydcLcN
NW9P5dF+9AaldpoKxJDISYEF+4HmoVw4q1gJEeRRP2G8gmCXQb8/mFiEHX/SF/o9
CQy/uAoQCAwmy4tk6PudcnFWY8fNw+GuXw6T4JoSejV7J83FRfGJ2zH+rDNudY46
MK4vSrOxUtVrW7EN4D6Y9xfD6bPuem/KG6eyxF2hiRF+oJBJTwMzdsp/DoyltrdZ
ISN8AK6Haeey7CQzHw87njF372SLm7AHbfU2q/GHmS1UlXA7evOA9WZMP7psNUec
ma+xGt1RUFX/vPTYhCkyWCo/MxbRlnuq4QMLXKo8uZJ3MuO/xe52DRKUx8hkQP3I
Zt/TAK+Ytiph0fiThUguHsEtbR1MaxBmzQUOBy9adwBgHnLFTM871IGdPnmRr9Vm
/Gdc1UbAiFb7Kexdan9uKP4UrT9SMiW6PJrg1IB03shJ4+/0i1H0M7yAl9s+KU3A
bDrIMhaCVDsMiqokfQGEYiZTH1yRNFU6MeOG7LR/vCpLhby5Vs7V8X6xIGI8fJEf
+mHARl/zcJ7hZLLhsBCz1xWdalzHIakW/hiE3cTWNXBv17dV45GiJlZ/I91jbLJm
CItt9h7jxlXOPCz/KTTjH7XyR+5TQFewGlRDr7GVIJTL3gVfSHG0WCt7/8Jfl4ot
cvlJvUfpOpWYNXDrlAMC9iFEQ38eYOYeUl6/hvfUuX++UP+ruDD4BmbMW5IWc2u8
BuHx3gaa+QJ6jatxJSBljFIQo7JEaklYDmJ+uAgW02gC4DQJv13/HgqQNq0VRPd3
V/7JxhfMV5WfUyiHf70sywYHKE8CfMGnp1IX9xzyae5f0RlbPrlJtGj2W1Xuhjud
+13TECljc89k8WtG1Ggd3lPcJ8piswel9+iHk6ageUc4LnUJMw4gbTjSyxEGjbHy
yJ2MmkY8+JXXGJmOJmlquhI42c3cM7crBO/Qj1G3wbaeRqw54y5V4isTKqOq1fvB
Pj/UPRgFF5M+YodDTT9lkA8KxYPsJZewyBd25hD5SSPQiRUU/EcqF/bw5cGoiUpd
bXKSXsdtQHw046kbB2iQL8xaoBPdIsiv6AciHWem5l30lPOeietpsqefkEVkiOhM
cXB8nOop2rDfHfoeVHmXWpXkd4E7nszVUJWwjL5uGIn6Z/OC/HbJPwCnHSKuGBN2
wKUELvoHaJ9WFrYQGbhOGfD+nXbFE4fzqdB1lJSI9qWwEaegmkf+fM0H1nOSvybP
lqbGMKOESP/zlgTi0IPeMfawbmvl64Sn6ZKVHbkdl79aJbB2voVazpDZW623AZZ5
MdFNepumDNkJO1Lba4CJ07TiCZT0wYzVb64HQ/X2vW8FRI1RKvLl1BueoLQ1jnz9
HPWMjEZLzkFdCjBg8Zwa+A7TW/8oiJ1n/UFDaQaglHKKD796TfZH9WeL7HJKg75S
XymWwA1Z+4M/LWgG1CxGp8RDtckFPASN7448JNWxpZORFIRAVUXtuqK3j4lDRiNc
SkT5XePndAB8cZ9pmg8hE8Rkzu7Thq7CxhSdP/MllmzNnOaRQ3dr0Pv7EynYrlis
622UqYJu87eVW165KxlXPBtiIXB24bNdEFSovqlXnC0cdB2Ar++SbaY10piWDvy/
jQ64lCVkQ9+IkHaVkW7MxHcpuPfnUSRa85a4oB+DYkNk20wKXJJDw4dvyV1I1T4V
VZsOr/87JUGEPygp7ljJ5GC2sGvwcG/1nH5ff+ulYexkvS5J5OHw4JImnuLBkqDU
+D5SR1ajl1zqhz5stgzt80ZSn/VqGcPm4A7pgQJFiQVJaWfWFVHzz7LHKsB6rlaG
KJF1n/wR8gaQQLrIkuSeNYf+6DoCNRUPq+jlVZzrwTjIsV5RtmxWnbCFftot5f2B
Z+YQtmhK3SaXHvqNId5GKdCxjzQtiRbHfnYROEGmzE5pAE4mYErkwivTZy8BSOXf
NvF7dbo4NrMnLZ97WQDYfZc+eL1QqlasaghbaLfyUvCL8FY5T9IADlcxaWegsG1x
z1O1zhgfCwQJpx3fjYyG6S7arW/7/51xzq4uvfrEjQHF6MsJPB3Sd3aWl+x0+Mc2
3cBPjrcKtC0lIUKDikjxYVR3KzoSbJ04buxdSG0ZuG0CL/8O2E92WFe6yk/8AeU2
chQFxW/+hqtoKH9mw5sqBw+S4iRiTzIoHq0PJtb0+NF1/DeTmrjrR3OqRwQD2xC1
Y8/CnjxEEwx4yWSyC3Gig7HXyBZ0vdznkn1ARVrGHHt3vYR4+qhvsOyYN17So1XV
P1Ig3Pz2lGYskh4ujXpcEU7rpOXyOX9pK5sUGA7A/6XfsUsTHrTJtPgFzlZKJOAG
tPuVzOxYqZwd+1cPrgwjqb6PqncALKKeGS/AjSHoMW83yxD1Jor5GGjCmAX9GDHE
nDbtxfei4QxhnnekIuT601Uy03Od+gqBMDH43mvHF8w+EB/MD5t9OWURSEdUbz1l
rNnWgYi3J1SKlseZ+IcEU4I5VKMzLOgHlY1Yx37CAgp8MlskyoGVGbRxCEop/WZc
WOO48/jRgiwqSVvhyKAni0+b4kUGLXNCqxJM8LOgjxQVabngr1gGXByGLhNTW6OA
BuBlptBSiN7ss8c5+U8ErPnt/0vaCVhwAZVxq7JhdMCuTO9H29V6CQWfj7bauiJl
5l/4duj+SIjiF4K25pHOBA02oKq5fFIsK1NYciS+upQJ0Lf21dKpYCMtE+qj5Oxu
L/EKZTeHPiX03d6eDerSh6cm1pTFT0ic5BZ+xV1yj/hERAcdeiQfY2L9cLmjJBGP
P6CDn3dlsvIg8FU0vFI56C3YLRrmlf7NbgYkf5Nk3QOlMgH2u0W2VLPQqXYrFKax
q5N/aTZ7nsHO/oGP5p1i64VUSDrUjUyaJLjG9UIzJwLLRUV3tPOAalLpM2FLOZuP
17UaiJthOc9p/wkQMRJzZANIuvvXHobQ4hmbjKEhy+gxBs94ehu0KwkkoP9CBN8f
Vqpq7sBEKCo8nvxwjS69v4HbjLuIgQwB80KU8fU+ZaFyQxQzrpwews7t92njc7+0
s6JzE3XrfNFPqkt9rkLp1xnPV+Hu7iUybMZgLwkiQouf15ylnkCcw26ujY/q2d6R
zGQ1JgW5XO6qYOh73Cm/4BJ5UwLTjyirHyRH28k5QRvhX/sKxSEOt2nUPq1iLc6H
2oFjtHlyEvVg/eEEh/mELogtvY4YJxDnxHeRTdkkaIZttnFny/PzKv5j5iT9OlMU
05oJWGt/QUP8WMyxXLFERD+LVD4zsdHXak6usQ6QjrgcQ2FN0L1cFYGQNQ5hpM+b
X0aqX4KyoAsmvi4iLunaKBGPyvrtRt3B75BIvzLfcvtC7+K1+Ni31ZxCf2JumvHB
oaYyN13cFOXEEikMvHulbDJ9PnedTdel3fRowKAswzvMjJdFOvad67rXacJC/K4w
MEygwZ4LDMQlrZs+BKAa+EK5YfNovsJcmtzryLBoWJPrmVVg4xE7t5QK0cG1H89x
EEl+KPGGsNzAe64XQ65q2LlKUpk7LK/zKa1SRvsyR8KYkmFdQklZGuVWYKEfy2gJ
ZY5ntDSmOJZpmHQe7QDZNd3fo50PcrkaY4qh6/daqH/mP/H+OX710Q1F1TWHUcWf
CX8FWrv1ZJwzoxn3RmENXNYgvOlMSs2ypOYHadTVRppgO0n51tiOuBTmM9n0OsW3
RxY+3CKboX6BGG1NM/XWR8weLExNZv5uqFwyIc5Qt5ujIIPUs9P7omBmnwRnS91n
mIUucyH5GOn2YnAkkI2I3vEwdamHRCMlb89kgysgb+wLUJDqkgbktn5wf4NRfxd5
R/VhGIdRpLuxjBFIRZiINMX8XlV7fj0R6EntgPRCcmWkrK+n37l0WdqLZxNuV+Lc
MJlgU7mkkqoD8FRjhUWd6bL0pFherSdJ6pF/SCRvu/193Kcnks6ZaTFPJf+evDc1
pnWyLJYkiAJV6SQslFunnna29bpeewwDkS2DeD1Wq1Vu1IjAUBkj5ajsuvPb53Bh
7KTvhEWjkO3CIzmHSAdaOvgLsv8ltmBPll1PmA9qqFowrqosW06CJr2YOpraq9dN
/mU0ThLHlqHoMrysV7jktCZlYnL84WIEMGKR2nAMON6D35mGJMjLMqte43yM53J7
otmTtG+wYMwOv18xs9rPzt3SxDvLvPSrIlxP2R4yNSQ7APQ5QhUcFaRhVUtHsopZ
LVbxUYRbaztO7IARD1HHiNTx2kL0SsjQC1tqzqa+lxbJA1/vYMQlTtZ6ufB7/9rL
MOGtlHybwhjYTlyjxrFR2/JaiadBf2EL0Nh8z0Jp/HB+y/gIjABQa6najqR6oeNf
ioF/pAkFOhH+F8cJTPCaiPUugdqsdyr1Aiogt9FOI1bbHx3GjIZAGibG8j8+FSuS
PWV1y8oAMe7jC6XIKRsyrK2qKvVQPJ6BOg/UUJ7nDO2yJmU391a21Q19JLwP9C0h
a3S0nsjsjUU9hHodpb4aZSh9gLehj5fO3+6Xw1MCVZzbLq5JjDk6h6oLfQQ+HQ5k
G9hlGdisbvYcCmd3vS+BJNgj8jvDL6o94Z8R9VCvrE27l2m9ULWir9WO1/Haa5ij
GtHFjo8sCKPHUiHrIq6kr6y5y3a56ursP0l3+UR4YfI0Lj02opANo2+Y+JO/C9EM
1zLpcVzegSAYxpVjxHF6E/2FOr3ks8TwyPO6T0GA1fBgYyM06dEt4J1u5leHSWjG
/K1f7wkpn1bYZHEVROMSCyXHTZQ2WXuPUPHpJwaN3uiSqIDII9kMIGUwDT7E7O/B
LUfO+x02BfAh6c+zcOtwFL0OQVe7zbMdv/TNZ041Jaufp5h3ZwQvsr1Q9RPyc9pp
RmhUMz1dh0+IiFuh4wVWVmg7CyB4InCwpWuT1rbBcrRTCeH6fCxJCM0IcA5lO2V6
fZ7Pt330PtcWixctRyuQTe+fu1mtxrb7cnVBzHdg/mfYN20DqPtI2mWvWAp6P+xX
P5tjc9OwXsn0U4epfgYaNSm0t0pRTKQs3AyBw5kOe33jbUp3j2UodlAgjZ1itw84
1gZuq0uXm9AAeP3TtHJBYddO6SaV24WZr8EgI5puCw2B8ipctgyEuT7HWikR7vi1
DAA4OLPFUWB8o1b+kxzFUb2CQI88nN2vTLvWYwTh5IBhweXKbznPP64Ziv/2I+BH
cJqMmmLkRpCR/QyMWIXkf4+U6vawF3TvE61p8Q+NlWoyscRts7HwcxofJby/4jRR
WmnNx3CKqgCBAXmPDS7eEuTAnPV81Bz1ETDY1QCXf33lQJIAfQZds1wK5eoR58OW
5u0JFkLCrpTIabSpb6+BB8bTZA13yGmwryazAZfa51h1twcfjrZy+7C4/zFxGgfh
9K5ZRawUaIMIfAIaFOCc3aOhKhYOWlvoCsXOtGyurMroZVH4Mv/vjXvSOgBgsKXV
NXDdd9PjIxLyX8bon6onF4ZT+o+FBofsfdlPHG6f3y4V4G7TeKEUR9Uud8S+j6j4
z1VSVWHHrhyM7D4Ghazfh0bg79QXJNjw4iAw1XnArs7sNBfLn4E90qjI/jOKJB83
VfqMbxIzwraJQT/Zr8J1lZiCpJCZlR7VcMb3P5rqvqHf5vzrdtj5+O8rp+yp8HKO
c4JlC9YdKYeEjtdFJKD6ThYAZoY6fsA4O7gd+Khmn/LpHzHyTDulYlvM1o/WU+GT
yATPJ3YEsySmpZoK9cKgQD9XK6YUJrj1BOcPrPDvae326qSdsOWzRyy1LCPoM6cV
1q+fZgkCJUddVCYiAQL/Y4AIKrGk0HvwICI3uQ8QxZXen7TMNj8gcCXeSPdWmZAs
X2Xq2XOSToWMjrm6OPOcVy8qx8tSl+cizTk9VJ43uFTMX3xW9/iJhr6Zz633l6EG
FCNtOF9QTtTl2buw3Z7d9pzDDqZNxA3TpYs4DI6AUdSH1OsjL7rmGx2jjuSE5Ebm
EkDUsScliGRAsGTf1hZYs3BMiDuawiXzPV6f/1it85r3+lH8xc/LHHZ87gYndqUL
Q6j37BmQouLrY+4H4COrIYYkYW5ihhJAgZ3alcrWhIyY71aox7Nzycleypxd/W0E
RPjhtgPOWiYbt1GQpPXPQv/HzizayF+JElty8DdmCK4r4C+g62h+OhqhBIxIFxYB
XVgVJ2ftMofV65VTMe3sui5WpqugQr6tT8ZSDNvQaYYe5KUXpPxVOWGV1DFhK/iB
PhnlwArUSTNYPLPzvy2rjvCaBwDMn9BgrzTnab5NjZNnr2IrfzIB98Zk+gaKalkd
D9VhmjQ1vRWaNp32ONUUWfBdIt/s/khCQUAWWI01BlciS7ojGOIUYJB8XFM6BgDg
2UqnxtFJrWvYxgzVUpWu/hyNU2lvY9lLi5bZLQFJHb3/xgkZ5U2osObysHiwH9u4
TVGHwiyLbRzRLPcLgObw9BbMRFVr24oHuJxxFMe//RR+Na9PjiN5xOxH2/kETNX8
xaCYTJYD4irt0/3r3rT3Kul/kUkgz6GnFATmDlChrQ83nIyGs0vYFt+q0s7+pokw
Jfnd3CbT0FRObvgmp5tPwLnPb7MnMdwyrn19zR3jBL2yb0UheYJ3OlPqFyE5y9Ae
P1DVSe49mt0EPbdDRI9KrdBT0/pk37yKs1D0dZS6uIeCRyT26jSCHjMfpV0bZa3Q
anutv7njzXIxZnHpzMMWyBg6Wgz6bwZmu/Nu48so5yw6fZVDrehBj+bfAdYL18AL
VtEnxtzr+9xNg113DwBi0+aNNYR+1goKXl3QIcP+1UP3gglXYeLD6fLrT/S/vXR7
fgfT1L8dWo4vFBnseQhb8Lb0j2WoyEaWlX9U7oUeYiOjPsBaJXVJzt+ptfyVSlZK
7RQD80QBX3zyf33fbbewAiRY2TN0BX2e9RSQeFlg5RZRfMs6JlVYvA/detj5ZEDU
biBdA7Lgjo8DiyTHn6JkYu7wYDLxoCxNWOANQHoNl1Au0Tnc2zmzeOuhW+bPsOME
7JOnPSR1sVC3TwHljgGgYmKxZHmFqwtJiu8Hox1STUNqeil6khsBO0yh61m69iRO
g3Pa8177KJQFluUhSJ9Ah7k6sL3Z8wfsFWBuNvw8RSyvnP1rzBvNLDlewSKLzMgM
Drx6C0LlHeEPGYh01AOujOrC0zL7Pl71FlrBqd6Zdt09W5B6C9mdqEXe1SbKVY2o
3lfET5D2Vomlff6IJtr195TLirLWs61OLvwgjpjz+oZmGas97nK++bhduh7NymFX
ulV88MzPP+FeSAPvITLOZ4YUNktYmivkxPU3QPA9Piq8yPozdL66mD4Uvp1Q0P2S
D1XvM9Sv6uVukQtWzs9PXBnH1DeCy047FAnG/o5pYCiFUG1de9zEMDQvfap+VB5D
u/S8yQbz8tXXevfGUrJNhqNBLw8BIvTdi4SomcDq558R6rU/tQ4GsuvkxQTJ+K4J
m1DI9Ko2ZKIzLD0UlJ0/IHKvQDfMk1Qbj+TWPlxNhZdQEQT3txAe8/Q+j1XT7WQl
ReQ3i5IqBkW+W0d5wq5Q99FM4Yhr7N1sMhoDw+5q8zbLzN+LVWy46xt+6YWYzSo4
uMjQcWnuHn+2e8dBbJlU1uNKi45ZGU1V1wFLb3CKlgRLOL+3GbUJOTrJtIm1e+Vp
rLb8x1J5Ug2lpT8dKJhwUntA4vK/KeBdcQorP6EfvGgu24ijzx51syuJZXeQA1Vr
h7TKP+9RcAUBA0jLLCtcxV1cR6CHEhsqwi0FR+wnOhqUHlZ/DHePnNUtvh7aO4WZ
X3w3ZD1DWh/Kg/GOWyaCU4+eLlKqmR5LwVzjAOlsRbi/K1FueJxzpKrzSPOYNaE6
F8E3R2gejOV2iYrdVztc2uZHv8w0yvqpmCZS5mmbqIrrvnnesQxbZUdPZf0zyFyy
/RDREa2OPJG/wlrJTVkn3jWNBIWB/2cvhe61Zpq9AktCisfjQ0HBQT6elwM5mBge
mlCc3j6GxIUleiPCsbFiK/ajFi6TwXtb9mINNt6E0XHR+wTNON0ZqVkqiKKVtXCp
xpSLt398/65UkiI8k+62alkPtjSRn0YbcCxDijFkUTp0l6bGmr/Vu0jUpOGuJlet
auHY9Bbq162JRSlXmswifXeU3TgYfDMvtnPQ7q7eecCIi2hcwLuPY1TObhmJvcLF
mJ5ZBG9Gm1AJ2BCcgKkkx9sXORrVYPP2CvgyZSvX2o3SW0FkC7F22nb4xI4MTyTh
+y/qi6wQ1VmjOdyV6UR+LBWJvaFw5RmKRrmL0STDUTLZCfUXjFZAR7bjFafS7n38
FXjtMxp0vqAqejeYX3zcY7oSxtYcXo65+GmfoZpvcI2QCvUgL11ttTQ3mnjBo+lh
eiHlX0+Q1RzXLPLNzEdCf7bn8Djyvb1jIFwxKUGLiEtxKXypc+CqDO1idh/H2P/3
Xvdf5GwvgzPSJ/wn1M0j9MKJZrJKCXrUMMyizWtyiY/5AKjEXWuzgexEwx9pnXV8
r1UTrsbieryvNDyZNzexCJvuXRdUXAUXOv/eq0fdbNFA3RTa1nMu45NGw6axqI5C
JmWRusX0QXUgcUzSgUvotLHq9zXYyFtMPMq/COCsj4jY5MRMa9GKuHW9+oW8uh3w
fd9zZmvsEdC8UEq84ZTp8/OjTh5qmEx10lFxLKCXW4dYJVqT/rQ6b0w5WoUonvE4
l5BLpA+v88+gx9df/6FM+QqG8fInsXZbKsP9K93yc0dEqBkIjnA2A0QcPOkTmPD/
PrYyTl8QKUbUI8d+ga0+rKYYOOZdkbAXwjW8WqVD2c6z88MKUZQwxlrNnvnDCo6Z
AR5+6Cpmkvw6eHxF+xI/OaYylSXOShAI8jd29n4c4zhgI6lVOEUhHdMj2bxWyb5b
y2jWW8U13GyWHSlUVqvl2Y6FJ4UTakHvmgGhEYzPqFsAM0cTPg2DmK5J/yLqXJsD
uyNiZDPvhvNEZdRqsU0S6yjrEwbxOfEJFxIMOeq2zBLwwmrlUMrovtMsQlMwkNxT
ec56slLMHRmpPoWb13YBr310xePZ/6AljTB54UFQJTJUwb94f9Oi0EvEUN4yGtxw
lflVTSKU+WF+q2btdaq/gvNCOZWF4DaNfg8who7ieAhoViSbCHEWgB/8ADa+T+Rb
+ElogXWJEczzs2Hz+x8C05RVLVuPi165Jpd0H2BUNppNPhr+YvgBr/URR5Sm/LGL
hyq7Cl0y0ZuEzh2QqxLehBL1tAgzM7nW+pJjpJsLWi9P7q6dG+3EXj9/AWgWMTSM
BvadSIQYz4yXf9rmYWl2ZAGwXlwPIPNquTFQGTejBpPDBC/nfEdePdGQMMRxOMXY
OOkh0dHBBgdHacgQ5XVV1HMENVYjo9zTDBBPbVBZb7a2Geys6eQnu+q4od2f6h60
e/x4NCDWAbM2QSdQf6sJLvP3ug/baQIsnkMEnRRFhZNsg5EklKEVRlXy+V9TPNQE
jcNDz3pkoLPqjuanRx+Yi5RJSCmynZDES/6wLdD022Z2t1pJOPhjqF5IvYNCwHaw
EaA2FLsjhwOFiVVRb24QgfTIIHr36o2AB6hE7JkGYNAIyyiBTIVKW7/xBh7923Ur
WmlVQ16ZJSWXNicgmtWR7yh5Ts+BZdfUqrknSSBxx4L4O9ps+u5tAv2AWknRlfzj
inuf3cZPECkQHCtN1KR0LbP3Xcu3Oa9MSLbtM6RTmVHOUKYlbYOeF4UmaUz5xP+Y
DfTNf6FsyxOLfrtuyrQZlDKL0VZiuSWCC0BKHqVlDPt50rwqoj3WZ1DIyxaCzKzV
C9QCwZnhmPQ13BecmeFwj0QV/iEfroXCQwt7XPSvp9pIpF6Y4yIdkW3SNTxmcbOE
++Gx+2UrXOAtdWa1XGh2MysRxuRdSGrxzScN818hppex6biDPCKiIZ8jLDMAlg7s
Z1qPieGl0UHNrWDZPKSfqY2UsmuAKr08AeUMd35XsbqecVmbBENx27dMUYex8iMv
ldM1MPysO1fQ/Yca+EltEyfZGns7Dm5D2zFYMssqq/RbMIv02ps6JpnB8BaTmIPl
Io93th9cJBVox/+Wt3ZTtDPQP/HF13B/4k2w4B0wNi8KH3TAWukCay9JdLj4qqcz
KYxXvmEpB8BE4uU98Ow+7I/zOmnKDzB8cuBueRlqVbYeuSRrHfn/Z7A2wuqy+6UV
F84K4GhERQ0G9CTB62XbMyrekcUGpLUmD5aS23YpAi3D62kUD5dl6WzIbu6MpDww
Rw3ty2TfXdIfV99MjwKGYqNdujd5+sd52G9pXnNJi5pOCngZPaLSCn46hjSxY7fz
lT/y/czTBwUg2kFjFj2lKBDHsqgyqM/x1fpG2mvpX1gTm/BNOpFiwUFul4OA0GMY
uHIjy8hFRVg9uEZk0+kb5chAlcqTPXT2XrHqSAmFYQws+Jc/7ryyJ60W7eQAnFzX
eS35CqykXgxWdpnfPGIPga5R9EUlpDC7g0nIDY/8B1vZ+E1SS+V64w0ZAu8Vta9G
xbK6hVqF9dlFj7FY38pl/rH7gLrV20rfZdbjhxWk4FUasPk0mPtD4Y6B1zYGUubb
YLBcaN/H4SQF4ci4S47SB4bM2/QTj/oRnZRyO5Ttjopszp/Gex0hq/f2nZB6rRAG
1VJ1EPQVw8NTgOEOZI/ktTassNI6RXztyTbo1vBcwDs2E3MGUkPC2bHEw9Kx3enj
cKrxwoldP5Rm9G0o7YSX8IeUw9SZ3/GS4jFFTUDHO0JNdlA8OI0XOwlF+1zuWc01
cI9QJraloCb2+GJ9NWRfeS3IXgsCupuR40PYXRwfjtz/TTG76/Ot4Dl1dgZCu/K+
k0DRSHMe74f8ZVC8ZBnjtCNsj9ErxcgE6sn28DiTfV299h8ZlSIsGXMJKE3TpPCf
skho61Wny2GPlWnCWlJ3+egVAL0nRjNwZWmmCfOWy1VYY+6fqzpsH6fBHLmZfKPF
oZthIcTfjCRnc1OHLJt1lJScOE+N1R4D4AfGmof2f7G/DpXReFki4ppiipZ+kjCk
m/hmSrG04EOJYIYHD0LdsYJDLERoM+qbsblXKXLA9sIl0bRjuKlum9KT5pKAB8jh
gfSSfUlAlArMmh5oOTVEPjCuoyzhEepcRcyDB6rbaOgIYnqYSfWVt7y3i+iMW0Md
GeSVcBm9xpy9CkHiXO4SkWGCa2k6z7csg9OVfl2edyJRUe2JQ/YyHv6OHegzD5Jg
Om0hTtB5mPgy8JMDqDfsmLt0HzaCeNemWqVTDJ9OSKkn92mZ4RcGs+iEVcmTH7KN
5RLOFtSpJRotHioupHVEFQsLGrPoFy7TWj4ppsy/KNR8VYy1/3AW1W2IYDVTywp9
HSL0NvGGMMwRbPT94gGp3SI31tgfpQHMOho6h/oYE46Dw87OjpMDGhc5VZRb948M
E3vwAOYb1UOhbMGGrtQ+GoTykm2ZJYwZy/nUEHQH55bT80Tc7xhZfVsXK6zcCpnG
tJ8rJPxMN55IlzXm8CZInDbs267BqboShvJ0LNAKQy5AysrCvUJcCpDvJK6wVDvE
1+K8zie7j7KG355jFpqBleBTOHAev3n/109gsJv9JxjYgDKmWxsSwr4km1q3RgLF
ZDEV21Fmdj+OQhw3QVwDsjtVb9MNeQU2nk4x0wcgGGf9QPVJEZanBK4YpbR16WuT
5+9XhRrERYvYmCLHrPc7R2Zd+5HLQBXbahF2SOYTo9G1k7pCmPT77hYskNgk2gSb
0KCnnmb8+kaLjbmK+iTNoS71BFzcKyhyxXEe2p6tDxBbJEVbrXHz2Enl5z/Pk/q+
XMXbcrOZgeNxt35GYQqOKwmvPTwLuGLpHl623rKE+4e3mtJDeiJhJ0yZnM8mIugR
a+ms5OUKqvd2DoDwPFlWiFet6Q3+bZzfheA/O18mCRW7gBb1sgSJCls4d8us4ahi
tbHWMeE51F3mWg40Ldw+rrzW5eJRJ/OeJONY4cMCrZEi9RgjIjL66HOLaX3FJgyd
aYhwvVnISiodXbXLeTJ/vjuWfufXWIC0rxD0Zcq75sab0L0u70Ka1aGfoedHJw3V
2drblfch5lFdHkSN6cHE14zn7Q8uXDRckznXUuiON3gbplMFUKPNtPShI2f8kN+9
LKzcd4h/DXmyOBBFxYiQ2vPDrcPelgTBKChVYpQP9I4Na9wFa2EM41SVurQan03Q
yppW9J0I4bRFjdOvTNiuzdGHREmSbumGAD+dKukJuHXTTcxbdvm96nXl2o59B9DO
on8xo0UUkdgtLzOwMNLZqMiVUpJkQg6UABtvwDDmRh217dZF7lc5fyMY1E3dtNTb
8722CE2Xwoi6Nx7Tmbxb5PTP4NxENR83KcPC3GjVU09WnyX/PzvZelg2m57ouKWY
pM9qUwjCvG2Nxtces0ET/V9osY4swVNMRfZYWGzCOaeT4/bVGKYSE6ujBt1s4FPW
mGVUjWWN2tI3gcfmXYjKAQiAzUdNt1i+yD5aKamgYDPeqPybMhD0vzaAmOBtC/d1
DMGknhVuXYcdqwZxMtKpUyFMUACNT3z6bL32aJTyooUfcoUgFjYI8hMRRnPt3aPM
co7TeEQYpgP13+mgNuKJ2am1WeFVCXCZAxrmYm1SOYAelTy+uZG4zgOGPBTJkLYC
/vvSq3tbACa7FCu7Ih2uMGlbD6/5lbZ9pIcoewZJfQXQnQ9kEKImVmyHBEjAiYQL
fj8mY5OEXJYkkoMeSMVxTbKChBq4WnygDs1/tf9WgWkm0Ks3LCYUfGVjNJRuH6ED
ioKEtcfPSKKRC4h4heCjMXWwRYndXDtMZ7hIUiuB9oDbXOuxDwPbM/KimIunFCmE
TxGpSySYbvuEHie1bcN33+Hkl9qtD4EVI8pHC+aEqtpcQL2SQo8K55u4Soy10//K
Mx5h+b1AnpfEjfRhhEyBe+/Rl6fTsY8EcNi8oSfbb8sBvRyiogrgBGGcqhTgB/8a
U/5EdRZegFv/hOcXAvG8D7liBl4w0gHnnsek2knuRHcojOt6JBCEovrApHEFRbCQ
YviIhra8T+saaFyUxCsNgRUJKY4aAQ2La72qA1mO7MYR4lvlU5enS7Xc26jNf/Jt
pgqECsKfCl6MB5GJcExQ70qPJXZVkaFf5xEODzDhkFw3svn8BT31l5gwCu+kEUxC
apep7WeljLmAh++ngxBwvV+w1Q8jgbZ9sF9+JFZurG00HkbstmmAbvyM+YQCFWll
cEwgRChFLu9xxVOU+K5F4oClzJzEiz5WWtqT4jYyizj6ShnLWcnzixdMCLbG13JR
67R+fHYEiNt0DvG52ulwqi+VC9u1E9dsLNHLsvlcHAx9/EjH/CDk86ATYy843Pc+
jE/UuZTNCS97vdJn1S2ssw==
`pragma protect end_protected
