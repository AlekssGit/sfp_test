// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
JwQVwkK+J6tZMC5w+BudKYQ6Qw+79hd4biGBLlWTsd+nRbH7HQsnV0JbHzaa4Gm6
3lIqoMN6Z+vKVfdJkc0Kq1YVMpetAfhz2qwbxbgIIIZ+K6X0nyhJpIFOAZyiSTCx
DpowikgjtCfrQM1hcnyvg2B8yA2+d9YZBORZ6pIgoNQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5232 )
`pragma protect data_block
QJ5UIecA0t9tTGSai+aZlrTo+LtRr57rMb97KToGLBlSN6qhc8/nqeQCA1TlHP8p
BPhDrPZBCxZNF8rJOhTyTCMgh1GcFrlHhK7qso/kLMY7P2FUvDulNJtSTz1UkhiQ
s9qw2R4FwK2fMLdt3is6N2FJhzRQGXkqXrT8i9uxIv8s+WI72BzDWSr5H4Dr87FB
Kw1yxJeNJv+I8Nei2AxkSZantfwxKlzO8dMHBZBNyQWeTzgFKsRQtlp43MxwhDP/
o1kdL3DMX72eI6Rhw+FvsS4CuIMYN0B/xzxziWen4oPgiy9+UKlEGw5uZfmh68ku
mgeuA1F8nWGOSV7m5dgcSHdcZ4jh2/aVtKGFYj18dUhjNJHC+WpU/rQ2YiwBU89g
F35+o000NHsOH+LCc/8WSB5g3eI7IhQv40BywYmzoFRSAZSrgV48xeCgVfgFhbxx
G4d5MrZDCW0ZI1n7Lw7ImjC2PvmOHhYvsr1L623EcWRic7drVImwMulGgPKl4xCe
/r1dPlax6Sh7mCYWhUnJxJBDAyFgrlQi2FcozaYEGCuEKMvBRuz2eE40pzelYQVp
fyBEOMrXIOYYoysdq4r1joJZsXKN3h8y2YjYjf8H9ZXqiyvdg5MqyQLUy3ZfQ0fm
cdTTvLwFRULbVLj54gVr32DFE7mQPQ0A9LZSvF/uRfOcrRH2EQyQI0eZrS2DXjLS
M1lvXTqq7owmE5xVg7Vx+ZsP3d0qf40is9CEkqYJhYsMmG3oj9KWeKRb240HtkRX
XPjaQYBzCOK10R7eSDTiec08fv/bRI6gjXYNpn/S5cMu3p8UsNazTSNkqLocUiGn
1tVgdrRrL3NVj763dph2SaDqCctlrCyXPCMNEDxOFqrCNWNOtfb94qp/I1NXVVyq
l2NLEY1C1rkr24tg+HFAQR4ns7nA68RXYo/1rdahUJkFNJxwBT3ayfk59v6vx7Hb
d2wN3mr/BmiIivfkhO8+HXq0bS4ZpD8uuz/F+iG1JnV1ecAqerSJRkw+BrsOYrON
XEbZJLWhrASGhScqrHCcmuxTEcM/DuFK/dZiAGlCcdK5whdN+SErUW9fzPMeto2m
zBsCVKhOefpw3MMyp6omZc1ppktuLK/LlTx9eKZb4G/kpoxNp7+eyqbkaQVgbU80
a4Y/017OWo4wj6U9kyUcdFnc2Hraa3nf0mtaJ3ZG/wUkEvFqAxncxc40JJVBxOTz
UxADH0D1n0khDJVnTNf0IyMBYC/oNlXzn7MlZAL2AL37wg5ksOet//BZabuAodgc
SPZnhHUFar2R+cKgh+17gkB1WW0vkrxBdlHkWo1YJ+3wH9OXUGJW4LWxtjK/uqda
/0VE8AcP5HnI5/mN7yUGhypI/HCDBQ1CTwYAhMN/qEsv4EmzQsivRvC7Dfh8QaPv
2oNzX8YWLkfi1a242dxLDDo/v4JZhefRk4bQOEUYm7u5l1uH31qR+iotM0RkMf1k
ieI7ZW3qQtFAkSqdQDNsZDQn1+ZFUrmcLmdhM2z+qwYjseWw4FNMW9URQLUgeq+j
x0WQA8QndjWozpkQ4qxY1vMJyX+3i6azuaMAeOiCHGnD4CgYal5ZLGiWwlN6dEdS
h+Bn5/Alckpt/ocpD4hXY45v766GZ6UV9Csm0Nk+8QzDT1C53TT0eiEZTNJUV8fZ
mUHMO7odAOf7sUo09Wn7R9qLonQpAGk765hBjyVEAkXzAOejTMxsxxepw+419HeD
E8aMGUtdEIM98e6C+Lpp8CKtJ++egHYLFxUe1xKDINnO/uoTvARPaa7ok3ph70mM
9A6EdPHIxDcocQC5PQpVd0LmJB1ajJc/K3pojDow1/V2lBXMadIxL19dUQHuwlly
0d+vZADx7b4OnYcdaO5dc9pCfwZnUMbBy+qOo+sedlKSa7EyFYPRJ9eVyE0Ki3bI
YRAj7seHs5jaKnGUQmdO3aHSumUS4oO7oYO9ZhKjMS9SCl1MHvBmqZJoEz7iRj/N
Obm5AuyfEgzgbbEpGHkUSlB69OEzXLqfFak8N2UZD/p3+CiLIa54scxXV0n4tvTx
V+lMqIHmzezDcJOYMZMD275uQ8tUtNtdwoHIKC3VOJPy48YbCPlv+EqFZPaSDHoS
Bo4n3LRPdbHdZuCsQ5b1KhBVMVvWRXF8940ziTkl8PSDinvH0wWrk9vWw+M5rA0M
fDyZ1wkxpH1CqXN1zCOibvf4RXNu4JcNtuNzjteCuV8EwskUIWUMU6Zho4SNbSey
wmITzu2pGX+PjyX037oNojK8VA859uKl/rjODS5oRGcdO+8ldAvvSrscoa0rNtyh
J+PGGbVdnHMp1vJjHkzcMV1TXFA4775B+o5Td9OWF6cFQjkTdJ4DYM5s/QN+R+uh
Wiz/3I+SRmFxcg0sFt24yYPERaJgOFWVKLa6+A+ItmwARNkS8fCnd5Uy8P6EEaAt
jVw8O5JosHg0uVyEQLmcyFoAIxRRZWBEA7kCZ/FWQSAH3t4HfKJr0Xxn20O2DiL6
bMJ45VMk/+niJ/xjKIDRLTwuf/k78kg85jEimxEhjJ5XVGaLCtawUusWnL292/7C
PXYilxz+ZaI/e5PbK3Cp7cGg9tokJ7EeOyvpMcyvOfKvxDroB6vjsGYvq5yaqOA2
iD48OJcqOHNpHtZZStdxnR0R7kGp8PT3OzwO51mequRjiP97KH9gWKez9U3eP5xo
lD12kiOf70iVWomv4Ho6/re77zqTmVLiVrCAriHREagygGXEdZ9LhbuGK/MXjoCv
wcmpO9Xuoh+5sWx9hQjTY+k3n1jH2V5iaKRTY04i2WkA4DGLppFQhkEyM2EgV1nP
2KHOlrWZsrtFpBLh0dJbSxgaMuHUjhhPyjhCvVeo7LATdf7bTRoD5dZDiVyrD6qT
YkOcw1GcgOQKpLxB36Q5rbQYZ9UuAPMMqmvx+iF3iYCH9l2tXQbc9rB6G/QhJ3ku
CqC59Gr3Kqfe5bM9QCq12tj21jBP3Tou9hsi6pIgpaXVZylryA1m0Exo0IuV9jc3
EZqIk/z2yD2KlZ8KoQZA2IKLC6rquGii+WM3NlzQKez7wq6/ScAXsDVl+PJi8ZjB
K4t06At/24lpayfEePtzfeVO2md3dIb/wg1mUJBIw2EOFi/HVoZAPC4Ibs9nknle
mdHlDaf4yJee5Cl+QG1HM8C1VZHJHbYxqullhAivpgWsb6guVSGZYUl5J1nl6+d2
xHoQOd9QlYZ9jNyq4Vy1TZk4vVeNwkjgeRN40/bow39uogG92/pVWEnFZBNe70Tx
PWFfyguFhwGfsOvI/saBvjQkieygJzlw1Sg1KJiLSQAfAaWSLCNfceaaDaU8SL6W
B21SprcTGm3OjZ76fxBOhqolCIm4Gy0uMpOMwRqBi0bK+s7T2h/vfqKPScevqgnE
FT5JgqaIp40miKC4/8H6NozkcFTi/adbds4aPCZ8JDo4P1AJuozbw3bsZu6gzSzP
BXy8Zkb4wjjC/JAT/KZW/zksaNJl2Mg92g5AI2/AY+130DnR4BFSNYK10i1QSchj
G4+rVEpLNn3t3NCgaFTWooEeul7XjqH7Bel2s+OeyJKPeO/mSSmm3p/QY45iaItu
Pf3w4osBDEYbBhGeQx3+/vig0rWC95/gSz1tY2Zj7K9Wd3n4Luj8B2FF3eqqFMRQ
nNDaW3Rm8XPQevoQ1X0nlMKX/dVO9GrS45xYqkKKBZEaziT4JRc5sHqbpIMG3fDw
ShwAuQRh728oINIdg0gJGmu7eR9WZiuzekO16JKO3kcHEneTnmgR2cjZ9UAF/b8c
JlHoiFQ8X6Al1YVobZPICPmhKWvHvrikR21CyGGUIVl6m2eQRbvJxQ1foESAWkNw
NmGrLOC+k9DirH4NQNGcZTOESgQJkbaNbzJVX107zt9eF+XicepRu2G8sMG42aYD
b5FLqmCyXADSMHrAixCmzYc6+JEW0N55lKWBeTSoT2g83Z6UChvpdz606ktR4K9Z
Ng1x3H0YwTEx4tNiEwyXeBhtSWnoigLCQSP1tFTeAenbz+JZEk2Y9C6YFVbmQlzb
KKc1QtpypkzBEbw3XCkyDX1zG73eYgAgwfLFZlkTdo5pjobej2ZVLhsQ0RaqHSAo
imS3J0uwS6BCmVLOW72wCLANaxwph+vZP2VpVLEmGBskPR61QPce5fQf6cbg3ZAb
z3WwVFb8gt55x05Ld1b1p8hoVqdsmofdhlw43BcOL/3PnKqLTBjomzv1malziFdl
j5b3/q2SWdQ3bg2x2h/9Z1X+zcK2eJAVf2GW5Frads59TgvXIFi3UhBIDVi/5dp9
OR8VVOjrfw1QNGDtMHO2wjKk4Q9+s4SYtG3hfeipPkmwifQm6gj3FovEZHwOaTjx
1NGJJUKLZ1RAcc6YEkbPnXC2zdK3Tyl91wSYMIrf21U2Pn4n+WjuxNwMwPvMKdF/
ma5E/cH3+soJWj6R/hv6zfbWXpoduCgMyGTp0o6HfXzKvTS0e4lkYPjtjlcV9eke
UIjtNs8B0wqvJzVyvQTB0JOD/CnPeNdnCnpU/WqLWpeA4qq1TpRsWu9dAVs6QxWu
nXcGWHoOOQrTe6WYf/qCdcb/U57daccRuKBqRVAFuJSK+MMX1vftT3uCTuLmduNF
LQ7UfMkAgV2jjcNi98dAdB4h1PkHBa9V9Cq464D99TIqZSMdAJ+yJqTmtuZIKKsZ
eeKOP/KzDDnEKWThPzrDSZ8zWlFtAoFR00ZKZgyQN7a9MAQ8FKb/eGTun75Rji+N
V3KCUAx+Can71QTo1aSEK9WIEKD9mBZ4CeG/Iplf9+Twp7+0j3kME3aCxZjOPWw3
q/UjH2IJfxz+SrkiDakZ2dCvnmtojylt09rC8B8Wg+hJaPrQ5ZEraIJWlDEAWxDR
aA8p/E/sPRCyN5Zqnxf/tzYM68Te4SUJ0+EmOa6QEL9fcFeofvHsjkcqJieokasj
5sawyS+LqNJtRHLc4gIeu1V9Xc0Xl4KhZCi9NJl4csxs+0dzDqr8Ky71Fvn0EO5t
KuTGplLvP9Xi2gTg/JvaGaIoL9MSDo9hmhCaEzGOrja50KHuVvHJ/jAOxKUT4zuz
vZK/1AJPvBMqm8iOSoMSo5d4sYl94iDHIPXIuD4c5B+fDv3vbnbyLyeCmrJkL6IF
SFSvp4vT098D3Mo2cG1pPhSYAW6/3Y9A9BvhXyNw6/B2RUY0WyymAotPfdaRNxwY
jdUgj6dLQKwtG61AK3mTf9E0Cwfyh5EqE39qGzCt54nAQTGFLwjvuQ0QWu2MEct2
H/Qgq0mt0qKAqzYdV2731lA5jsojPGYaLG9aleoEIkWSnSv3+rQArCEgWbDmxRvj
9r7p9cRE3o2nSa2R5w65Bal4WtCsPqyQpXsZM3FebNyOoGIhQkkyEApxzQm2EEh6
y7SxnHdESbqa3R5S+QX/Lcs4WBCfllkuQd/LYsRq6OnWa3NC/7y9gLdpaod1TeMK
WWQCxsa9T+BWdbVcdGCxqPOpfOlT0I1xiYsE17v9447P4tMUbAQd6V8RL24QD4G3
me6CeBM5eljV9O7NcmXKPv5tYc55ZpWW7/xO/qbPhb2g3K8BJ8tQXgpbEhJWl0EQ
BI0XOBK62jZ4J40CAPIT2SWVR42AAgSRZJHL+6iYlN0GcqwaHI8k+IvUxqo3f5Ke
i/XN92waWY9VXR5HFBQ3oGsr+Y7lBIORJpFiSi23U63wB4Ctoof+0UIUE4740yp0
xia/8cZ9wv2kpkZCbfV2q+2Pw9F9o1SmzG+SMfQ71TwqR8EB2HMY5F4+XiQUCCXe
YgkAfBs+V9oxhZoBVFXZPolveoZV5H5DKyJajEgXz3jWUF6eaXAyV8hWuHwpsKqr
dvKaqMC62ezrHyI7DPpYGK2JEjK/6YTwx8tq7JQ9DODm4KObBO7UdJcM6NZf0GzL
IJs7DXM6gaKr1+NGigZTujRBp3O+aTFNQ2BtPuqpmgxsDqDGPqK86vf8luX73o4Q
GI9ouaRGuLcnobmA19oBAVMRZdk+cDDdeS36rgOAHbiSG7Ght0MXuTWUlLGN8i6/
yWAVQkQiVGxftKJvHI2YexssK6Tx0dVywfmHe4xXwbOm/3zSkwuP1MZz8e/ku4g0
b3gRhCWbxmGQeRtR9l5hNdqMpfGIcE7r2SKSyyHL1kgv1mr3iwunRMnLjOAP1g2s
gLg0ebREkRVfn+FwrxcYqnByhnojJoWZXlG7vIZs3A2Q3kVM+gOEcBWHkj8Lomqb
KF//TNbuMhwQUkYHPwucH+u3bxBbzSB4WzeHiJwSbxB0KzTeYwsGJxRdLT1dZ3Mm
s82MquCkucqQgAbT4IeDFIO8USaS05fM1SCDvYW82/rWVO0NPE3RQpCzJaVbYVzU
g7V223NCtwbGH3IIiKew8JtC4ZcRC+w43GD2RMwlZFp/sutUB3swvdHv9G0hrI6H
p9Q9ahqBZ0ft+fAqCMuTvcMIhJOL7Tl+P95mMgXwS87dWPTZfScFVVINZSAMVx/q
BASObfu1BOVukjcZjdBEWfE+8V9bsQ/C7IwRcNspk+hRk6UZ7Iay6GhkqOrhlgaq
A54oQc90IdiS2CM089SpR7pqGspjz9VabK0navx6NopptzLjUFBhc2hFaUBf08Hn
+v31Ku1pQ8nuQZDCWovXb805vEddJd4dt3kSy+BeHQVcqJoqcxrvfw1PRdGxs5SB
eWl9c06nVXPzBluC7uChUOdc+npvupqJZD/2qqMleXE41XOswjQQ//8CiH5+VgVj
XAGIx9Ic2HYJi7cyHWnaYl4YxHNP+dDEQKaW058fodA9pIK5DiuCJ9ZSNuhYLnz1
hHzvU1V3wAszkXrLH3tafdQzvpSAdsf7/6hUG8re3dYf9J1RpCDWhxqUOh8IBOna
CyS2z7/apDAY04Okbwm0STI5pVKCnWdjR4pfkyPrTJ6CBTBjiYWsZYdov0h6qiYi
pOlxxDknETnH5/Q5HkHKAtADVTEGN7yZbnl21NU9wCV1ExZAF4JIN0DM19xCTy5T

`pragma protect end_protected
