`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
QbN1fxlmPrtabHiH9PvjPLWLoPjshsDKB95/3Vg1hxMabMicgPzf/ZtJXd30lWz5
HW1yfr+EHkt8bx3QwE152PNxR1RHzUIMsC0hbAOfrNwDxCoTyMhaT8NwzkMJ0ISg
bGnpaGi32OHFIn+h+ileNj0Etx9LvvQ+qZNDrwiFZ0A=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 9344), data_block
VirN0WJZXLDB7p0Tq8N5eOXIiH/1T5EQKSCKF3ThsvYeYNH31ThfDwC9dw7hhfn7
4oOJR2r1gyv78uCOwJFtlkbBMJokzILwmCaseEDH95GSGaa1QbDd4m4CtvRid/sr
s4RhpR3kTG3+DWRMI5yOOyc+OEu/dmRYSUvBNbQDPlggBzbch4NAzfDzWMcgKd++
96+iz7VOMo3i1Bn+Ka6AbYNLUoRW/N55R6I3se5eIfWIRkmXciUVTxc1bk1U8u+p
8YMS8EgM0x5cUjttC6uv8IfoKiPRvpSAhRMwxB1CmPb+ymaO0l/v8H06CmKAvPYj
bhTpW6znY1CA132VcL/WoHvYye8a2TvU/l8MqSdXi64xjAJ5W0sSf+BD+4UN0raq
95dJQzeUC4MJv/OuL5YIrpkKJ9SXLpNrfeHXzVoPAu5STR9ODsib687ge6Jolosw
+vqB9xhvQnGqxUYp2yMlpDJbv1FAQBwsif7uWYhwk3RL17b9dOPOJeMeoQbRON7A
zXD9ye4ZWkeZJZyqFVaFSgDcVjRAeUToWhgmt/I1YE00RXn/pyk9jLxT43RMUmUN
RYlAL7A1U0sONyTjFf9BUiW8h4XsgMfqcBtdEVhF+y+1YSPAsUtHn6USgYmBmh53
gDHv92W56bwx9L7reluVvTwPCx1lSk3epRh3gxSugVPD17kqVx/76cze4CoxrKRc
u6NSdAZkuNyA5oTawTMDUzkP9xVT6PDNefuKO/liA+POH3d5Q9a98RIQhEN/bz9R
Tq4q61kOqcJGbwHgWziK0IEZVq5IMR84554ahVqGvK2lWNcEgILm7+23idouaVQC
C1QioSr6CY2VPlGwkBLYY7BFRmTlx1wgPeg57RfvaB5J2syK0/75I+MsnZ2oeFNx
eB7g7Dy1K784U7yEs258N5dbsMMQNPmPH5PYf/B8+i9dAC5JDvs/Wmi0ZemPUK5t
yJCdbNrT7UXDxbMvcIT2djRQaAaNvTeEFKo/HXwFvoIOFLjXaqwNJm/Px3m3U26U
w/0W821ktua2ilwM+M963Q38BIWlozaJP9WQrJr5L4AIURtF93ayv/4RaR8inYSe
b5l4kQgLEjOliz4n6OXieHI9EcLnkOHeMKpV4hycFr5gPgFI0Oqrgy8IUTzvVdGa
5/292Zxvgzq/k+NgX6ea963kvPvrGLSpwI/LPqikSaFp7Yw+NUyxGhgm0L+Di+wC
mWc2F/ap13zYLX8EwmWLnx1U517tfv4Kav5pXlkqG8a/5Ra329Cj+cVu/7zpJLln
HHlCsFXDjF0iGve3b8OGi051tsyVxlTfD+WfDd8HhdBAwRqid+RhDCc/YX4b/apc
Qxn622vyiNYfSeRcaHttIGBKIGyW4F7rlWJuxpGxR9II2JEThxoVI4M5dI7O9/T9
zh+T01owy93E/Vu2Rxk8aKd3eEpMuPCIcp1a6UWfIRxtkeo5KdWIhdUfzrWTPlIe
wSaHTHznW4Ea498RLo79SEVgJg1aSqsoLETr4AsFxoNOxtktJmydgxHvnYt2aj6i
Ho3CrmzRhVPKyP0EM6lBWPjFPl7l/ZocTg+WzkDSbnvbHK4MjFh1EtYurmjMl2SM
QO3e3x4HtkUQyiYFCcSnZK/6vbF5QK/mnWplVMLTu3X0lrYoOQwSXegIDZST8I53
l6O2C74+k2ocOnAvmg65rARf1ebN1h40J8Zei2yQGJZC156HumW+wmuLoWle2GVW
UD2odKMLnvc3SjC5QiKYfJBAnoza1y8NN3g7cNpWdio2GAQH/gCSMGjrx1HX5pNo
CyQ6ugFruPScGEGNcwHh8ZdrHOe3tPGkG7mssguDGeyGKk9O9eJyE4Vzhd8ZLwEu
nzhVrtgsozzsjO5gE59GWTBRiJ2/MAhNR7VLI2mamfwJea33KnBzionL49cyRs1h
YFHIsrETfiAN3LnttEhtTmRaNluutxDH94f6p06E8EYlpxugtDE+4BG4LmQB+Ctp
f7staE0MfJf7e+mBo3DgYjZ15hL9j9bNweFHpYEtKl0+Jqv7aUVviwbSaHhpLKX2
sPIykMaMpUG9MsISlQ2EwgeB1TyIA+mT8+KYZ1wwmGd1WRpoNQDboL0kS+o4Z9NM
wQdbTVawzPIa7eMLGzXQkBNzqqKlDeyi2Tj/8RUcP93SSRYTUbxpPfyOdseaEdMD
r8uqDoJ2fFe9QRAZg3BxQ7s+oHBo2AeY0iArIhJ26XRaPb3h2MSZBSP/DZ7mGE6p
ZsbkM7VpspQckieDXNP+Ebh3JNpifXivGGkRp+B8WMmRojwWdGFffq7RxAp8ufbG
1WOSrLCuSAnAzjiiu82XLMaVf51p5ZRqkWAVTN22lTWvPetnGTXf0bYt4e4XRMSl
hp2zSXYmJubzBYfn8u7AP3esHYnWYTkCaENlW4aT8gM19q2NX81bfMf7/AroirXZ
7ykqfDjUbH4gxa0iMr/5aTdojy4Rb2DxQnF1SZKfbvVH8rjbzu47vW9z4wEObFP0
6yAwA53/W6xTyKc2ysoO1IoCOlI0jKmHUm8RYIDEk+t7sLrva/e3W2FYmy6TrJqN
iKNLZCPtATY1sNHiog2+qGIiBoQ/gX3PiNHOqCfWsF1w3Kflb7g+u3UgsMhzbNmO
vEKcwQJIbzP7zeLqF6QOwRHGNWzvD7ClOaMLIaAZRasxNEQQlE7gs9IfeLAweBU+
pfjHkHIZ4+3nBsbq1yoWKLCqNEQUqpND787X/OGQDztKVcDY/7dxCW9e/Lh9iGWc
3TGg2A30LQ02Wgvy8sNZnMNHchdKpGP5eDzI3ef1Jb4D5nDIGhGA/+JAHKKoz73y
Yz73gyrlLzcklJYDGELn/uedO4A44m7BCrPJTN3XFp133Vs54CX1qj7ceS9PfjPQ
SL2Yws/tMcl3lC9RwGEvgqCMYDDIfcxePgtOarkltMXzIrTwZkSVP8Sabqq7O4kl
GRtqT+XEJzEHTmJi8fw0/p7Mhthi7RPi22Am/r+qiPYuL410xkHgcUAocTsGyd/Q
DWFX31QgpgyawRM6XvxeETn55crsZqihmsoqRhfrviN1ZNNZgf/HCvNyR5F/n8t1
Q+B4CEjSjmkHzQNoqBMWlVxVG9MxIJjRKz7b2YfZDxAJHIMkErlxx3fi5Jx/nK0q
VTaOw0biefWyqTA7ZcTArqJ7Sk0vI6umHFZkJS5seFTDwfo8/emggF+jALdKfApG
QlooV+nyl1h0lF8uIcAjETptJZkxPX9kX0bD+GGfpi68zJsiMVrMoICqejTF2xny
sFlJFEqBmtITsb6JU2c5HzpZ4tLdbcU9UT1IkoWLaTO1fm7hcyp5gQSMN896Il7E
6omqNI5NSUyrTtJmtcvGXO0OhWPLVR9DpyF+52qAbr4BFuE1oeMRO17V0GK0eShT
GD5LEJm3IM9YE4lYQBq9LP2yag+lrJdGHp4DFYwH9aPUFDd9K9rzJSdJiMy1giGY
V8nVbaoXWxkkvL0pGf1MiBOneagFN1+ki5xgrl34MOUqVFLXmhlN7h0KJNjNbjqQ
6yZxCutRA0pAsVIA6CXnpZlNaDNU0uFCb5ByU/nG3/TRBBdGag+p5cGf5xoWgcD6
SFbhWWUVXp7TXqXDxsdQ7QlrrfIEMy3XPDLzzy2ABnRdMFG7ReOCLNv05afK+VOi
nyVgT4n5CLQG47xwsevNGZzdnFLwRHXaf4dRvUFTmR/pKqp+iE9SQIMfJCt4XCOR
npggta5heZHA6GfaDfGcQBL7teo3oLTm2ZhloWJ6rWhIkdc1xi2Zav85RMbPLBRM
Krui+juPClPwF0pwMLsnyNEVzXwL3vT3YDDGArVdIgAEEd0yPe6yTgw59cbplQqO
/fQAIv4Nr/Ld+N2q4816WuZVjEVbXfcAZCuCGTf7oyWHx52hZB69PQr1wJk6xeuf
ijImfaqI0UjkvZdkWB6vb0HnHIVvzgq6FYPTrqnQYR/73r6QopD7ZLHJeoIG9nHD
ZeFQApI9LTzmaWtC1axOzYj7o2B0ua/i5pKW4MJ/zkWJkfz1c+1kHU5QFRUAPSQH
LDGw9p0rgivNO4D54i+qVXhTjBn4ZYlQfE1ELZhAVhyOqRm+lL8jqyplMrvCekK0
JmTVWXTE5ID9SkRJ0a9oDCbFVltUK/63TyF14c2KX/T6qi/svbMF4UAxN0Fz+AVH
3+rUXPLGZpGvy9hVIx0Akyg0YR05BlBahpdf0IzZZ0vDzEq2obbmeeDCnnU8WbJs
8UjCjOcHyoVFs8nqldljCUnM14/7G7XHUcsjpBRxikYDgy2nrtMzcy2B8CgkrO0v
WmUPKEclCbnn800z5+2bjHx8okMEuFGKWUtPgil7qNnW2wal/vNzVZMXtQE/9dnz
iE76yvj+AdI8a0A07DsF6fAG35sBGPBMmjI1emzY3VijsZFncZW+xR5uor/itnOi
3MM7bnzb6XQu35U5gvsUR2qESpPOXypg00t5ztwg9kxPFgp1+uR9nIOFw3ZM11zG
mtqsn9NytGZyghOu5+EzWbsHesbqMOSFOXUal82qwXGSFz9PX/AR4Qv0MI9i60wj
Y5pVzV3OOcOEwbrD1skXyCytBdz8O6ekx+FalCjdyo5vWr1gfdl3LxJ/TJMwVMfV
NYI4HgQT4DlqwcnvItaSUEx1ClhfuhKiY7gXtOa59u10xJfrnLmPzikwo4lst6GN
xf16aJ5C6zKe/MQ4QiV5qkBbwqPYl+9ZbFvAwFYx24nS/yymLJRv5ghGUYsESDfc
p6lwXVUTnofHhKP6DS82QSNrvS91VIkfW04HXIgMYiMSsFtWHC2hOdruEnTK/Y6F
G/G8/S/PraNbG+1ZaAPHZRviwFc+5KA+/3fUH+d8dUgXNvO6N+AjgakRzkxdKfr8
xqTAoMcng/x67Q7ksNiktxi2/2eX9REUVYs52xJpYgxc+69NZ+R27rAqUwOaBzBs
K8xFgdrxdfrnr8AtSiD1XgCHOUVBWK/mko2Lp9jQxz82Mq+530BwDe4Yaobl1t7M
cMuTFtJSUlS/UsaQqvbQxvLTkbKYIkssyrncSAb9qcBJKGhU4aKrq8yGADpl1W7J
eRiYS42lem1xg++X/E+b/n5gJlcbNqzrTgOBLEqb3TqXdmdKJmiRm9KcNlKX7M4c
Nsunt4O3NhEUHuqySN42tGgCysa+lWBik9QQg7vmbROxVsDEJ2CRzOoIXKYn4n+6
fvTGpiYrBJ00Rd939SjqUxi2EVZui3GWhxmT9wlRu2UMbjF0Kja7orFo0nHgXJNw
ESRtirGRPKgPXo426H6yi3IzRPNuF3L9GNXATw+gTD4hsclbM1I6EbQuPAR5JUqa
BqKRBOfTJGv7rM2StXXvuVzQyax71S7b88cFpagL1Y5MiL//nJO1zT+J6nias2Rg
iBDZGj5MfDZjTQDt5TJSiNzCKDxzE7ODZ7AnLwQHr3/DmMVctls8hEr266b7IoJ0
WQrkv64AgHpHTXfbt4JN4h1OQxal6oXWvtWsR5nl6ZFn5jLsi0w2ZbEB69n9/Zhc
CxuO70a0x3zfemYdv29KbUxg5etbFnpso5HjWPsFTQYd8Z0vVWceVBuOgU7mJCGm
m+8SM0AEU7m/Ufv/jF6csQ/n+dlmYCbtle0+tptkXLVitUTTR2xwhvRKaCzqH4xL
nX2GUaX5DBODYqu1QgCJ3kgJH+inWVYWGXzoavmsZ+YO10gmp7JsmJhQ7os37G3a
aDdSW4h84VAm3VMuMg9JInvcDltSeLkbk8jfzB1nk5fmc5ZtXaFJJx9FDivOrqqD
BuT2tM/bkE03RHYx15qD5nrI7FXmVsdVCoRmOefIL8E3HPgMOl5YUdEK+ypdzi0x
c/UhNp1Lkc679zz0QLkk7yikc/haDcu1pkh3xB2nj9gZ1j/doN8W7U8iRn+y9G2h
0U6dmDBSu6vdx2nao9hnLv5qEg4fw4I271mo5nnfqXpKjgEF4olhYTBjrIANgJJ6
hvJZKMzgXnwPEwtXe8ce1ly+BN207O+x05831t+SB4gdZffocUH12E+UiYVR+E/G
xHPzPj27R8PRppAEYem4w2EY7QdK4KxqPP9zUBDy+479uFl5Zu5g5sEPsdi19mB0
4uHE6xBTTaPnOB2BV+F3FUZU2P11mx6urIlidSTThD920jt/m4bq37YWOntYTYY1
SgX71JlVpWOMMOXxdJ0dSIDAswNRaDtBxhkZamUEVdhGlYQBCa2Y37l/W3BQSl+1
FTmRH3BYW2utBmei/mf44JMybghaBCi7OnLMHNp/x7zio0vxGTP5D7o1EnM+D0au
WcnCTbtl+Rs1jkMiykj9TcOxopGCkY/7YgJJgTJXrFXlI8tGDQlJ3khcIelwPdVq
EXQWy367sJAI1yUM+fbzV+9PkEHgW8/BQsz1yuKPSVcrq707PpUBp9qvwNsDMTBY
27cxHyMm19ut8tvShorFccr9aV5Enn1o3pwLvNbe4L9A2Iu9p5XH9UR+4HVqk3E+
RsKTirw8nnM0IGntVjjNeflK4sgCC5p02r7hGdL53nQaC4DKM6QLa1W/+nu3L3sJ
LlaCBIBBLlp21+HAKfHAiCQA/w+kYFHrc+ZP/FSHG6VTopVQGbabwaxdkvV6pDF4
4MgDwEVVxrDuIpywn0piRhjjzljVEMWgYYKAj87DyLQyUCU27ZtPqiUh7zvapQj0
TQ7mbUuaGiovPpk7/idj2LP1jUO5G8NSAAsqd92CjvmRgXs6836NXluI/QJz8pv3
VvG9CLLVO1Z1wVqKaBGYupka8cIiTtTm/94cZ8Ro+4exQKT12fyRWOuUJ9MZJuoL
a0Urgm8AqLGtIfMgpoLQ53eOen/C8vwcIecxNbaa3u6Li4uMGEfX7etnu22IwTrN
Q/Jn7haa+pQlQe3w/jtBQL2QWmM5TL00XOzNMH40bma/FHsJY3VkuFFNs5Ya16VU
RmmaylYsBfRLfQGngxVvSjbrgOZHkJ17lAytIIO6kpEyuK9QzDgKcCYEqeivRImw
O2xg7OkURdvvVUW1nY2YbJHuPaqD0ononWFfhQIEfRhoww5EPJjOwOLOQLBnPCZn
JbiwT1yhjPvujWBa79k/6uOwvIEfxM8NAp1NEFqQmwmYh651JMlPdlZtItCF0a4Z
N4yKP09l0ZeZ3O++259I7LnEQ+OP636ArN2JYYxzUhL95okRtBcrVnn/cWlWm863
I30lhjsteNoHKrbg3HH5ONg0KXE+6091TrzQd9krNNOkSzM6Q4UTstdRM1024L7n
HXDNoXVip2xv9TdMojt/UllaILrdP4eKhH/ws1qV3NM5LPJID6tUJ1C6u6CtEVr3
/diDngWPIGYu9o/2dHXEkPFG8gqiiGGJjKX+7Rhlis4ZogyiMq/VjLfO19dMZjfr
WlaUxfBa8onssVZsBtrh44uQOyvc3ARKczWjdGM1oblJ+zr743xgyYYZfHS1GZ+g
QpUHjDV6S3Q0ZiRzSKDsLA95vHEj7keptsSjLrpHDnh9cQXdoqsnl8yve8jvn2YI
KM4aFOUHvwy6sLUYQvn5HxYY+6wujSoTBfFRTGDX66QUuEn3t+xVhIcTyFrjtq5V
pm4+F8yfF+F4TtH4X9FX7juyG3SNkp1CxC8t3WWhJTjH3YLaVIsOLFuCPEpRdjRA
A1jcsa5Fos85ePq/upsdRz2AxpqORi3GDMsAHwxQj8DBigSWfDhi/LMQYfVY4Xzv
6vo8EPpY1W2dhLITDzBMGDSSmQp5Ob/mOKSviYb98bFY1kLv++luAfBznyN+X/vA
AeoRYS3/9p9iZM8cnEExJeOYxXmXj6PSLj4OodH58TRpUMpcXWZhZa7YOpY8RXwK
MBut07m7QFdZugEfFiTdpxq3TirWBv4Q48rm0wT1OtbGi2P2Ka0q8h+/Sy0Hj0uY
4s2Ot87/txerTl3m9Q/YvXlSVCp4FNGDgvh9dZFzvUtXot8sxVl/oqlVcJmJeBHC
DtjMs8EpP9ZOVmgfOb+sbDyBoxIp7YFgVaF9s1YhhSbPGZ0Nqt1CHZ9avYSoHBsA
cUNDNv3SUgnsy4Hlx0YAigfGS+AHVqiuxUpDYM6RtwbhLu47L0fnppSbOAtyPs5s
uhD4Vd/iJupFHHchb83ln9t/OXVpJCBJKd/AUrrMwB0mgBPDuOlocCXSiwklWL8f
ruJFTtbNGJ4syJU7vNKKjEsw3if0tfOzsj//apDW9MsGf/CSkpKGC+KsDzFwtamS
ZivXe119Rc5EWIWSS8Fuzx2wWAdbCHdYaejkmW1jRqVcPxWb1AfEB1CvXoq8sUF7
ebmlWIcTlQJGQdzsTxzQH5d5F7vKeaIlSfffi7EzK+/ZYjkbz+0EnU1MwtpnL+iw
ppaZtCv9wITqKimX+xSPnz5h1kcmZV90s/UCWCDnapcFWlM681gEJFcJOde4WPNk
GzX/heFZlzvGBW4PkBMXU01Z4N7lGGEj5qnMWJm+f4Yfx+lRXf/l5T708m5TxXCO
Xo7QqvMExCy2aLoFenkREtrKWar7FHbYSo2ifsUI1VX5j6dRqlbhpTZjunngMXO7
L5gpovbtADYotmAmDnwxoz9W7cU8TP3MhT6IPXgoQLJldGkCKzte8aNME3eD9y/O
U3E/MasXjyTbgfvXcGz2+6ewFN3T/apbHPBLrzmbS5vXz/xH1GPLEvic+mMuYSO6
4tqXMUenxf1IcHFzpoDRQkXp1rLa4LgTbtvRz2CoxCT4MNlxr321sMxTtKOkzrXS
S1e1q/nGxtLQ35gAbped7YezGTk0cLZo8IhiX1XmenXkHrMSszbgUDJtfgWQI0ye
HSessZ0kMEmjfHs113qB14MCZyhNgazspi+8spTG1oxZM2sgngZ5r1f2uuq53zWN
xLhHPk9YGSqRSuUZZr50EC9OzzsIwPLjQv38vAwiU5a16/MS5fa0wQTzPuBBi7bf
Qy2YQZQFqENBBio3WQBmlWRlDUwU6t/Ch8mAWrHyaRx/PX1r7fw1/rWuF9Li5WTX
1AMwQ7T33mi/mzgt7WWmBPduu+MKoUWMIEAqDZ94ZJBna8yTyzc9HSWmPkCwh0UP
uwHRtszPdm1+bWTGlum5oPw0rEjaMwhGL/YiKCMbW5Kr2qP5WHgzvnGVbl0q6B7u
NnueHCuKEx29zMeCbKG0fnTkB3df2/IDRFezbZc1TWJJV+miXcGsD8QbW13uWUcL
2bR91xNN7E0wdFBc5hGbvWMUyzcvMOQQnrVSdArstQlkLyR6jd4JEA2NPh9zAqHs
IrN1fnVSvpLzitg29iykQlXGsGIkXfpFlG6Ov9uoXNrshK9dw//jJblJYP1CRuos
eJ0ZZlAs4lnDhZCwauJJJd0NvLCeFdHpkFgm75mPNRq1Y4V+h8QvevUgaUCieQ+V
1helIJrT/pHh5jpAsr2mr5n7H/3cLgJA1YzT21BUdu+pu6Xgt4bfl5BHsqJFKAsK
SNxYxcDs9YrCA2QFlNDnn+ifOwuHDOnv4a+zRyqQSqOuGJHVbY0Zzq4v06agxmw+
+YOYPxr+Tv9vBr7mhX+rmAlBSwAVhOEsd/4/yUOddcTbYaUBcJ4CSSy/AG511kbt
xqreV8pcD4PjfNrCbp4K/WHTDv/A1JIfkvEu970dlPiSvmkr/2O/rYkT87ev+gED
2e6zz1cxaQEKlHnqDcG/yuOBFv6pcqldrRU9DkmMVu9MNH5lFCHu8a1A+x1f2lmq
GEis4C0GPfiPu4hy/28P4N2F6G8zkD4INgxoK3v7DZxi9T3GiFqHR2V7f0J7ewlS
lHnYtf77AirlH3Rulklg18OIYj1R0hsibpEDah3L49yBHRV8YNX5T1ZJmYgz1brG
7I6cZloCy9i9zx8Tsc4kXNlIr76xCaiZnwzAlRwzXKv/0h/FcW37JnpEqAeexNMC
+QvKC6iiSnLNrhxqV68+ym8aD2KPSwQNMhzGZCAEDCS8mkSF/ojW/zjoSrRpv+z5
sdeBcUIf/wJjJj+uvO/GXwbdnQ1vThrispWGdfZf0TVWUv8vAx0gAMwhLB8gm7mu
nistuqfsnGIxSw3Aw0mJbVvWF6FU4fKqn2zHYXr+ey53h61j//PT39rkuif1IVGw
rUrqbxH2jCOPUuEuxCV79QNRBeov6MweDDjYQXBBlfT3gQK7JJvl7E+ixv2IZQK7
7BZeYhHeg32zRRvbi1rGfk1B3OR/sj9/jdp4levoddO5UIaAv/Fmkf9K5pwLODgP
ybOnqpZG1iZMdBkBBfnlYgPOypNAyJVfKCpyq00/+FjQUjlyzAiGP5cX1rnzT9yK
InyfRrah1MB2HEp+KEd/0ziqVyrKGIPEqWnwJftsCd3M0fVUs4VCWxAOp87e5GrP
TwuntEEeb/6R7D7Ank4/H93eXDeLbBh46mKh7TABQxWX8B8Yeq9UjtUlVQh8yU5k
tONmxp3T6oadPCG9YyqT9PZPrB5cYrNFaeV+k8mqxQ4bMnc5dbrMoGhDyiGLddyb
kNnEuBAryRtXWh6XEOLKb4xCIC01YSpFPjS/QKWIserCpBXLi/cnDLT4wGBofQi4
AOll8mJr0tjZZWds1F2gksxxDI3qM23b0MoYYz4JWzlSI4PYSOJfXZInwDHwlrIb
/Vmg1qqWwX6d1XCCpBO9cQ/2XGv6XpBZF5CoM/Fs54DfejYbaDC7DVWQbPkflpHb
JOl4JzLOV+8pnEEn/1UNCiEQEqHMAXESwpm4FakNQZKC0v1aGNYE4wRvKe4bY5l7
UVzLXM1rn6mDCrnMGaSczMZVVR8YRi9u9A+M+G/0YUG44g0epzctT4b3U+Uk9Cqc
ZVi9S+NtQ7pEXKA4/KuLDAO+HtKyTVeYFFxoYrDYAbQnjdaCZdg7esIUbGLZ0Zt5
i7i9LcPpUIlEeZ0B3KKNU5AdrV+DCOz5jWrB3Gn1BBQtYk+evbmgJfsPePspBJtl
L3ID5STatsRea5p01jFR3t2uEH0M2Jmc4etSeVr5tFrX17NsVdcqeuAKvD8/qG1J
szcRHGv0RI04aWix7KgJrfxlTOWHIVR4f0TkrvvPhgi55Fci7Alg4xLAW68WiLpU
WENaOEvGMvVdzP2HrmvQ+H64t7/wfukuING9qs/vyIarkoRZT8u0dkukFbYCDoHL
eixy1tYNopnmIKHtv3exm1yvfBfpFUVRR+eTmIk03h3snp0+kbiXrKHej0oN0/A9
iuZbNhXFl5gmD2Kb41e9CleWKUsmwcAV6wM37TScvC1uaUzwgL42PVkE/2CdLXpA
VcuXqn0VY/r4H665gpSEFhxyHfKIPF5A6hXNOabZlmzJQC5miIet8E1gUVTrVvEt
t7mHwwg2FUmhshzat7aVh6+uVdPidHJ1pu1Gyr22asFJp7/WyrvjAQHeoF0qHI8I
yNqK7C+w28897pljLSs8BsFgm+Vbyr+vE2x7TFzbR/v0K1v0xL7DDwfaEN0p38J/
LSb2PttDOJsF9RgeauqRWvIfxnInYCtdReJ2DpOy511nNfXDXpu1Dv4FoAB/HQQk
LgLb0V9yaxAJeBtpnuyu4uMF3FELUpBPKe8ioDl4WfmLI79jHNFFynhuneFkQjR5
gAKZjXMmNNBFrriS70jq6jeV5x848b5YAsB47PeaQvurZzBUAC0o45DDfpYlOaV6
MWSAXEi7L8q3fjqmrJQFaXdS/XDTQmAi4D41J/o7Hd4M9tRIvY7gDJp8MqKx2Z1D
XhmAfVXmeT/eKjddz7S7h/yduve5TK0FKwqvR0vk7q9mst2acTM0oCY9Lfy4CKXE
jcTDz80LpJ04S4xEKM+5gurOSGkeXET1tBoKmKxhCPdzAuqAWhevVNFwkYI7rhKq
RK3V60CHRadsE/UMwkV3x4heZzPWW+aPAxuN2/by2O8ix7RtgKMh4oWQPXZuvAdv
lhjp3BH8uWN7np3vkj3WGiHY5861u421wXpnUVdr+iMZdazBZK4sW5xYsUxYMXzH
14uaILo++/DmfMSbHOFx9Un6kpmMnKbLxHUQY8uTb7+4v4QERpyOwOlvgjXeAI6E
M5kXs8dn2pPBVntMKim1yIzaYSGaf7Go+Grc51pGmw/brF79WuS2CMkf+m3omdRn
eg477hBQhia/mERDC4/BtKDwsXKLZWf2/5o1+zyeqRfXt8wHHJVqhmm9qDzlXhpA
KEDM6BMhgyLmvdXUDAxYIDB3U6aq3AQbTCRZrNU35FbG3G4UGN9FBTpYUFP75TfL
AzlBdLxNvojd0TkZLVDVXWZol1GtPnvPvH1aVcH3ooPTBMzNXav7sKAG6/JmiZmV
1Ykr4ZrVHY8DjRN97B2sqV9Hn5XIBSnO8mCHA/9mMtHK0+B7URsPj8KhZ+B5jfBz
wXl1y+DLp54IyrS2SHWDuGmt3b9gfVD1TK8aRavUlDI2kXqSTTPAW8u/FxPTLW1+
scTNTo71y1FRiNm3JAuwGtE90LTqJRvheARrBt/Ty4CkNyFb5qjJMXye7QwpzDc5
r13+uTFt+TCyBLrl+zkLO+EBGBLJ4r+g/bsOI1CvQPE=
`pragma protect end_protected
