`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
iRZQyfzytS5pL7zVhPW/95Q7oExEE9OM4Ay8bCFCeWS+EmIAMB6tM7si3kYFCI7U
0hlBlK/O9dWcW29B8y/zE7J+CZhQERq4eEPIWSeaLfBOl1MnLzPNaihESktdQ9GB
x1riZHHRlPkRd/76obhGBkDIYmqVAUuUA7JkHuxQ/Cg=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2992), data_block
zeyFPGU1/T7ChQIq/1BjmL5JPu+WOIH+h/MCWNTJpXXoORm+0QbV/M/CbKPAPMo8
wgizF840nDuYm1GgiwS4W9hvKc4UbekTAIrDIc4w2EOlVZnNry2hX2PQAmYYs2RA
o7ZKfa7DjHNZ8A8avpjp2Yb5cSK59fXQIrDGTQccroS2N2Y3tqU5MQgJ3NqI5Q4J
tlEiupuhXjkgPqfg1/4L/3/stOe0pYuDlLOumMK+pvWUX+kGUilkAgNwOEY2lmup
RwGglGXo3ALaDQfCpy+sU1y3Y/YRqDjK45cT9icJk4BLvUcwzlOamNLZ0jFEfy77
oS2WYJctmnrsMtHjMFR1WsfJSiZJPlLGN0dMS4RXomoGjozj3NkWmDKN2ypNIHCB
UJ2VqQHJOCkON9j7uC96LZRdFpXDWo7+K+lumHh0ZU8v4zCDzAYzhMcIsciL9f0R
kF0QWNYV/X/0sA6jJMxjkPpvi5MCTX+eRvmxHEJobYCJPmlH+C3U4MQCVz7ySGMm
0FoBw2BDBY2c1cSzMuzksTpbRQKqW+Gnbtwz+uTM1tD7dS/gnJ6nPbhkdksR8hh4
BR8Z6XBO+mxc1260W41waeXk2yWYSK7wTJIxMD52wAdGzRy4ytdzGAH7Okal/93l
LVq/IqIpD02DDGPebCufQCRqehMCukYnxPR2fQ07bhRLoD/pKv5xHHQ1gyyAc/Bd
02+utlAEqTstf594gdCypf4gcikkKvLR5mXir+PolxdwJ0UlcGzGixl6bVXiHf7H
6MMXQD4IKsbi0eK44A20E6cWNPl54v1/glAktSl9rnv6NcckGmvqt8yk/b2ECXR7
ApRyVThp4Q3rY+keSThxpY56Im759jieqiQyDjgRCSN8sqxO0wpp3Ez7h2aiyugG
wgMl0nf/KC9/OXoKf9XUUm7Hmb5TbF7qhFVWErGgCkDJYSD0fs9bSY3/9et3gult
MlBgbQRLwg4FHHrLB8+gx24vRrMx8SzR/v2/l1SvUzVKNuwuOJMnpiTG7056fuJC
apKSa6TuW80gjp2oL7MwKLFYWrdxWkVOt0L8K23GmD9RTLgljecj4+MKs6rd/Agn
L+JB01f2ZPo6QF8ZY/VE3DMAJGfATK73DovFgpxH9r4RMkkE9r3QgVQdytXwUqkE
6DMBatiK13wvd0rKz78VPt7oN0vcz1UvHez1FicA+ZGvDAXzF4QAASXdXJKWjua2
zI7sIuUsTxwDeFO44A1kFT0bUHg14B9RVgrlJp2zImHz0QzMrQ2bhODB+tZ4y6i8
qj9p/kvoq2lJWTGKERtwIdKv9FfqqdXyMsKlWTwGnNo6E2vIgnMXi0jme16nVYf9
9+dNHYNX2HF4ruH+7hUoYhEzNTL8q0JWe/uWRuMq3Twt4bGDAacJeztmR0TVNHvR
d8pTP3xlgTSa8ApnEd3uzCxwCz/bM83of9VwhaXOFbwyLeBo53nRQy/NmVfUOK0a
h9e3uo5aqGlAQovnNZwD8XF130gCeYfW56G1M69BeW0mRLDWG5sPN+3RfKBssR3v
hB6M4rfPN8sD4TDm8GBPomZFhH5fnTO1wW3xp2G1G3wNeJsn2QZp15s7j1UBssZD
aK2PytHnfZANYNX4uKO8Tw32Uw9z+8+6+osE7AmlUo7lddxjxi+tw5UmlE7v80yq
mNdGJAyg0qcc+7PV53VkwitPkNSr6r2lHW3tZQZZ5KLuTmmeJWctRtOus+6K70hr
IlFF1HoYhRfdjEbDzX4eDmyewEobpKTj+VUZen/eh7NKwmWP9hoLC5g+r88CaoEK
abEWCny71KCPrSMaKmBY5cKQN9ngWwXhQilTNair5tEpbsKMUPSs0bigE8Wv33FN
ncf6TzLxZHw1OvWjy9zeYf8yKGEQU/kw9Q/GBEXj0D/icSrLPa0mdmHzYr8xoeIt
m5UUsOejSLRitcp+TDRaCa3A5DIvGWjvLaLyfrC/Qy6imOniuSzS9+7KzcsWPuan
1+uSGCgqN/ypCCEz5jBzjvlnb35CL8nEgMKWzB67TNudwZIk6+JALagaQHeaM5yt
SnWBYJOFYoFK8OfkzLX4dbykHGelhqH2BCYNE/JTlN8uBwroZGK2yjWIRbMIff0B
GKPTWI/FybyMlRSb5XjWG8DF7aIisYSNkNBP+dgSGsfU+Md9Z4uHT3YXTo9O/CSF
/Wn1VAASuUi1pEbB4t3ytXE5YnmsKUckn8KPbZpQypRNbLiscAcn02Vcd5FUK059
Njujaqiez1eveqQLrz/DpR0+cu+NrDBs1C1Z49gJr3dOQP1MWeixDU5jgR+lVOKC
NkFPe7UFQ6VbFCMKDAuDCBcddV2CNICfcxiavVpFUOP9CZXpqhqopbCpW7eCuxw/
3dMXb/PTF3X3eqG2q+tjuFRBOKwP86gZ3UijPjBb/sl08vLoAl3N7FdcaehvtZVB
TnDhMud2kHPcFefmgRuzMGLO7XRwvdFCXHNpDTyWkjUlBotINLR/VL8KS9zEUNKQ
T9L9MOV8zfH9mkZ8/jOIoE63qa+/toZ3+LgAIb+XlZiO61op5mQ7W4uWLT0Jnv3n
xXVZTtAG5GrRtmR/xFEF1CtkSgdG1w0qAmn4tzciBvA/yTUCVGHqurq+0qoQeZAM
G949RPEm2PKSMofQs6MBtfL4Ng7dVqw4aASoeNVmoSyLLt7PhmihG7Bznk9Xa+E8
qWwjJH5t3/6CA0fJZh1Wm6ErfzVlviD1IX2zEadhqB5D2abNFmQo5wpQ9Qmw+p99
FKv4/IR+Qxnl8HPS2y90ByiGCi4aB7dS1Xn47WfOFan+zpDgby76C6cXa5SZov5/
0WCK566xVGJ58pLoaOYRbBOv7jQycnTOZjTqUg/KRPXBQJPAkmhqc49rydn4enH0
ztv3Z9FKyCfIUUmNFhdPHCh3nR9MJPd7NdV59jNXrUXdCWuN/UoyQviQp6B/WLSG
GBQ3CBORCkqMNgwyYn7ven23nRi8XMG9KkiAn6bgo/4GHRZhYiqo68sD5vMdeiHu
5V+1gupS4mW7MGEQP1DVRyVgjrQYgvTUuN1Unj9xT61a2OYcXIfAesR0Yq3VhA22
dHaVwtqHmInUh8FenG6+LauREVP2NUd2RMhe/Qf/MNhojCcn4mfD+187MHjQm3fB
YIjk/94wi4H/SFc0XpX+XEuBNrMmHeeVns4HM7r1mRC7ifEjqehgz47mChUmL1g7
riWbSa2LRdLVvL0RfS9StdTq/rSCk4Yt42tOfTkOFurmuS9yOp3ZD2u6itw58i2N
Y7Bz6p3Plk29hCae+3rqFYybt2ayhip/9fJrhYmV8FBrD4C5VWdBaA3t1L801g+R
pRpBbAQWuBG2Ufu3zAn3qwwaIWqFpNyBE7yFuUK20Ge4JruNfYyvnr4Vl4vyUyJ9
csSViQ0CFmmRVfxtTQsqbqtcCfgKdOlmTJCrlbLSAga4FO4rCJeapcWZpGvJY7Sp
gcfWKz4m3e8LoC+K8YJ+TMOIxhGVODAG0QqjS8W8KbLS6grmYZsWaW5m2b6CqRtr
T3pNLHTcaBmB8ykGOqxEA045VZFPXFDb2L7MZ78V33kvCfJPCP/NFjP87eSjx5gB
wUe4nBBNvfgEO0U6blDQt6WysKmnV+WhJeO1Xgp9GDWC60N4PgfIFyRuDV3g90zC
h+vp0p4aLDjiIBzlFCGrOkPpuVP1+NsLC2vCJBu0nzWFhjnovPedhxGIhtxcjZZN
8kTnWB+h/od2/ximlUcMXd2DrPsNtuK2RTbzavjcTU6EYF1PH1GTqWn7b0uWrglp
JxmmWv4pF06OQ2RSxZr0J2vScc++V6GgpZ7dw0RURKOxgjnv4zRaJxarhbpAd2l1
vdmG8ihqemOFEyesGZE77niPlan5qBcl+h/jJ5bxztiAS4lM8Ywysv+N5P/9xEfC
nMtRMZxbts79jcaCic+keLJ8tdO12Umb4tlN1k7ke4dAWbur62KrBKc8UICm81hg
Y1wbYnNWi2959p/VoWlvAw==
`pragma protect end_protected
