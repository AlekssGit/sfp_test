`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Jqn2R0hyYE3OpY4pzO6rK/spsgmjE4rJ1s9UrGTyXNC6OhTVnpZpdNQbCiYu+8dj
zM1aCUg2ojQJacIH0SzzGnPk3mRFTsuiVIdzq0qSOCk7UEHKSNx4tehNDU1lf6YL
T5xyE9AbCmiTossSI6FgZ1wnPhS7PXj2hknbMzY6RMA=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2452544), data_block
5jhjIVm7DkUhm+3xoKtpHJ6sG7LmTT9XYgnDzlgdSn4JvfdLQY0yHuvvWu4oivmD
t5kK0IL0qAI4uKP7qHBcYPk+ovpR+RoJEh7TycNeW3c+fV4TYp+u60sRJCpMmvx3
YkuDT4AL21NvkTwJZQfW9sTnueVwP0kN8j/JFBxWopw0EXjUKyUoZ7kC37/3LY87
FtEV6MR1CKwlFsZCtwpHJx/6DJOvDRIUFtmC5M1uL4p1uFLFNO+flya96I0tGXLv
tVoBwdz91aNfe46gjYII1GoBl0B/Qe4ayRUAFFUTsSh+Q+Iit7ZO/jUPctuXy7MI
ke6DCJD2VH6CHX1ea6fod3fieX2TeOscVHp/bRDUnNVuGkBRfgrdqBzuXfDPaa7D
lfRJvvV3YioZUprTYsjzZhftQXI0ByXKCMv0mglzvmbP8sGgF/Y0uvEkwfw3G9y9
zT0LJsaeABwaKE0EcwhaPLJmHuuPKG2ek3Gp1MW375NYNT12IWRaIt+HNj0Ja+sD
UCThZdHrMuJw4Lk/E/CIkTGaVHTPDTnE6Cxs6FZeNCHKFNHaPPvCZd+SlbgGdqGL
Nlwt5yO+gEUWC58VpFYQwXjp69PKn0v+FqPov6cHzOg+iNAslK1ceqOr+sqjBdlU
dmtrvjoBEMNFVCINu1lW3OGYyVCRfec9ObkKPeuO/jt4bH84PId+861IcwZPtGGA
q+6/jYMpmQoiUXEoVqDxWKNWE8ul4TM5UKxSXMonStXxYI+C92PKtSK2IFsKMzHQ
TmpDx5+OokdxM2LDDW9Teh8MwRfTucHKj3j6gTQTY7rqDXGclrgncL0MSEOBLa8c
vseZnp2/pZFgJwG+9Mg3fPMVEru7sIRw1Fppciw07WO3332VuGQ4ErN+HOl93Ld8
hML/S2HDnQzHdjI0eFWwF9sR7YZhP5AJm6O1y2KF13i7KMfyLD3HekOU6VbPvQTR
Ldsb2zKiVLYhTiaH1joZfMnhsnleO9onVjXRpVH/JVl0nKDvLZ7QH7HRg167eAFY
QdL7t1Wm2h13Q/x9nOyo5LdaH/BlEeRASiLHfOxFp+OC8z3y6p2RmdXVECAsIp2/
o8OQqBTF43+8qUKUkZKA3zZl1WOGGiYWtnEdu70d13N5wNtlmZScFCoqPQkkRSSM
ZhkUC6TW+K+gZgCpSQU3k3jbL+UEXpvOMtrcxp2iM5w6YxQ6nri6x9gZDAaxVvtv
9npbqJTcJvfIU63PwV35nyB2sy0eQT34gN+tSBfmncs/LqLA3RJVI2ZsWOlcnFBR
4XmrWCUQ+nAvbgu9Uefj3fHD3bl4Il/y+6TbwAAxIoaZmuNQzBCkLFR8eDBmZ7V1
+ugE1EdDixnmsrBg2CtuXdLo3iYgmT3GuxzeieJlEg+0nS9Jnb5a2dWiuewNxjpS
3ajYhYl7+pyPIasTlddTh5DL2eNHZGAsf0MlV/EsiUq1HhishsxuZqDdW0ivii3C
XZviH91icr4wQnfvxq+LoxtjZ53752K1rjHuT3DeOLrVo3Cg/LqAjS5Vgn2Zj0tF
ayBx8ctnvOJ0X6T41jg5ocwm8YnES8Y+1RClYJCFfhBuwo/dV8FxsN3DTi/bPBgl
tQKLhSgNLvBPdOVB+PTH3ZPiDLysr/AairjBAe4bwBsvQgQ5lXqZZNHzlzeaglyo
X17v5JkXrL+ClJ/FAJH4E7PXNYi4gITWM2Fr9AGJsXUnyAXbwc1OmcnS+BwF5ajW
bZJJcv2GiII0dD7VBOShVCRkBs8W9i2Dbgjv/WhTL0HICCNYUhbBWlBbUbr12bUG
X1DKB44UJHnSfX/CAo8NCMwBqMGfc4Ms+UJNlaD6oI2h55Bh/rjbKrlHFf6zbSNa
IW74K/PkGQPlxseWqNTJvX3p0BUulZZl5YstR/j4abaBbgdEDb8Itl+Uv6eTTE2g
rlp7om0JQ48mn5+QtIX4OTpkI1CtEBxuLElfkcFbVx+ANAK51KHoHLiOUk/2+rOp
PMxG1sRQAcAvoeHaNp9yoPUjEofpYKmANuvHZYu0iZmi1xKnQwnRTK0tMsoCf0mu
O+GKVYuHgvhFjqSmbzl6OMST4yoz0XL1Kihhm4if/i2Zmk2BV7YGz/e3GLzWZlsq
QxhGOEKR6jc3uxcIr+ddGGLXJPvCSKDvUZ9sKLVfirKcVy/wj0Usq9fkQDpgY1jo
e0JmYQstGyJ/1VLgipCqwT/yeuxx+FSY4L/K2tnHpQ5JMZOslbjUFFVmXD5jb7bs
4A2+4cspogQ2cTPwIfCwvfX/Le7iC896I4COCcjjoaBCJhDC3X2/HKWXxEa+71uh
3cmnaq8htyYWbI4EBgoX6GLrpcM4zWOCKsT+wq7mI9gCSONUrQqNPlIOdWaD+7zT
xLH36Am7UdY2DNNz7R4WbxhKoA995vfxYulOdLdazzBAZNgCDFaeJbrj6jMNChV1
gyBmexHOBWZi7qkWGG/4HiuNavxMU1BP7eAFlihVLNLyPybMuzMOYDGAun8o0Wju
NEvaQuzxQn5l38llxBr3OprV6wzJSyYiG/aNrM+ofo1OVVf3HiOj4xl2yfroOFag
Gmhf0P0Gc2qsEBMVoAp1aTZs6ErcdRn2JQ5ZwBGNeLGe6FAe0+sjjE3u8YVIJEFH
0jtsAIcTNZa1UjEOABpe+0oi0tuKxro9MzILIi6OtbZPC7bemxjSEcqblvC6AHTH
XuDS2FyiVVa5LUbpnt8uMlIlpnvYeuaY3DOcg7f+9RGpfK+9PJ4besHCsraKORbp
4RR45swAafSR0Sughbow/ooXuSbsPI20jha3I3f99yHICxeQgGayQmBxCrIEo/vj
+lniJUGQfKb4SpywfkEVEx021oUT4u/EFcrsNY39AOILhmvLnlb38+04txQ4Lnqz
hEEc2p0DcDVLgo5HTPHi9PXakciMzr3YrNM9kvBJD2hoMIeEHdF6oRZA1Vd9QBwO
ye1uAWmYTpwt8nFx4BuvRVts7kxAjPK/NR7bR1sZz1iataInbk2RaLAPNmReZH/e
3cauXNx80i7/5aOmqhGi878eU1L4fQdPkyec8WkOHa6hvK4RRXv2a+GCxgp6Es0n
rzV8wXc45jMXkJXdwXQ60jGyufVhgIZV58no2HH5Me6Sq62ceR2moks/daqcHas+
9JzniNQ7uCbn6xoec4Zo3eGq2CteGq960iDbO5nngFiZlMRAPtdaC1fHsyNdaaa/
HFfX/pFMiA2P97J61wO7uR07raOYu02PaQ3VJwvj/C8aMLMu/HqeY2Evk+zIlP/W
Sa8bZXRGJkqzQoTdWgintqT4pHRBjrPIhMQymscnxJAlQAPLKxKY6RACoZO606wc
alEc10bB2pmn1/Zb7NpQnMYByDhb6JV3Uz9TWzZXwZD0EggHnefWybevAZUztnpm
YispBzfOWS8zg2Ly3fW7rLGE95oIh9Yx2mHPqwgq+JBYsTuyMG5zktspoWZRwV/C
sNkskgrWw5OG9S4Xg0X2a8aLcFVT8A4mF0v8NJbxE06vMntrvj52vAK6k/3Xaz7/
pla6hpmvbK2emWkKQVFdisVFDTGh+7jBB5XnP5f3kjqfmg0wus3qRLk0Jl/PiIwi
1CK20Xz3Brzs+5Blen7hhS5/0HT0saEPTQPFpUOkFu8LxZWkRAtuBGM6pxlb1VO6
mTJAX2prdJ/LCLLpkordL+jBUXK8HWeza2JEmEC6IXsUs1P3a/LwOASEufrIBVqW
cyiEdOMo8YKJzXCFr5yY2G9EULvvh9hi+/RUeht8nVRz0+kyHw6L+FX7lkKXFQ0n
7YfXwvPKfKNCVxL28Od/XmOuUq9+UDP4dBj71Pf4GJ/os4MOqJX1WV5dI8BMIBhY
m+8x7KRKCnd/InFIk/+uS0ZZMFGDSyFUS3/MwyaxR72RlnIsscE2kmIo8ZKJmBx6
FvjnVriuDo+sT1OdkjYD2RCKo11nZqLAQrx4lKCglzft/9BKwnzjK02h5lD/aH2w
vF/n1Icue6NpGzH4vninhfHMPPtbKHhJ0lvhcGMipzIrc08qzQOQC7rqjrZ7HyFi
Vzgqg33enll+eZLGvMRH4vfiD5lPYNK2lvP+bgzuAG6KpjjZPido8Ey8GZSQA9G4
a7MTAbTJsEQtcZLAQBMlrMDNrMha6sqNnNbFSoTx+NV9w7O51M8mpv4pSebcpmFD
dFee9A8Fx7NPCIrZc+Mj2xpv7ACzF+/rlmOwOjgKt1ZDMZdATF+3cwIA86tGHwiF
9ZpxLrgEyrye8sJ7rTncRqqg+3Azz0Xpyk8AtVBKjp7VzT+/5jF69gEKAPg7sYDM
YX8a9RLhMRYQebItECMTbjIa8Yl+5TP3obvDTMSnDzGvxmwrJk3fZXy43xFPwgDx
5XIbvP0+W1Jssjkp7C3UzRAGfLVBf1TzManjj3MaO6x4ZDw3zsETOc1JJnOb1q21
ACtmYGni//V/7S4Aqw9KvGtGzdnmr/iRqLsJIpgjSexQbObHuOqqq4M73RCdRPm4
Z8Pj/3FhBxBUD4KY35elnau6D/Ta9V53eK7Og7RrXS1NUSiEVlEMI6GqS+AHW8ec
2YNxcP8nQAGqj6h2kgKYnTyj7QWN2RbPtf0QdBZueKLflLnIGyde0DFLhHxpa3DH
KjMEvTvdyUiFoAJfGOPIrEZJvnuVi8PX+8J5JsLsWlYmA9+gtkj/AIOOZgYJewUq
+aA8kzAwAKDcf+yfbKKpUmaRpl5xsBvLnbxDNORXG/rXwZo/4y+4jTKqJCx2JshQ
sD1iHrlQ0lzXY2D2dW/7fexBomWvTrRH5tQ5ESwOg8TB0lWAsJHJnNXSxX5VkkHb
o1ztNdOhKvGfu9tbYD7joNR8wofe3cpF+b6UgSP+ZAA24ZriyrcfYVb8JHtGs/bJ
ps1DyWEhGQgF523AcLKAsqZvXwVGAczu2WD7cQ/luO5feZMSGfYgzYg40LizSkvN
Mxsa4RLhBXbov+9Ee50WbRlQxijp24CUaFRjKEdUDDt72FUTHtDhQZ0LnuIqgQDT
4SJ+WNPJbyQp+Nzugdx2kjelcn9DysSqe/xYkwNohWw/+hSnPU+BhfnRbPMIAPFw
b/Xt53f/IpCOYxlxVqAL85qD/RvWMw3Wi0nfQHE6skR3JAPiHHry8Dc7yIJjP9Xp
1iMAt7uAJffs7O/2054JOnGK3fSSNohaeMqgYIl1u8CTgAvKs8Yl79f0iI1y/Of7
2AQMTo8giUl3nPc+phcHaKiqQFwMSWBOr9AvpogyRfER6QA/6HzuU7FJLpbYiGAZ
RFYKJ7n855S0gVTn3hByY/r0HK1gfbIKtcyJ4iXhxPjvl25CQIRtdTK99JzhpK4t
+YtIONs8UCAqbAnANLgR4ahCeoWRNPRDnyk+I8y3NWy1+DOyXDjsGZXpZO0xoHU0
dFAMBAgaFQqzJ5OFvq0q6jXdvKHrG2sCp2QXGnWhnYx13nhjhxSfHtwyjof+YJ8Q
Ff5a9sBxzCWmSzvVWs815lCW6v7+ojeSmn/T9qJnNFdJTfxj5ECkdzj8SyW1+MRY
cHzqqTCilMSmyup/o82HkBD2Zla3ADpWvY8ooxyRIGQciiMlWiFMEc3z4gPn0P4u
PJ8bZbkXEi+tyqhd3YMjBjfmZctg0yQFON5rCRtehqA1qubYjsbMVdCdKAyDkcBW
c4OJY7rbmyZWBSR3yZAW4Q0HWtO/gUMOIhOtBBDVx8f9sUY+umDkdwYCaD11Z2qI
12sQeiTQclcvN2L5XnvPfNIvDUq8XSjaonfrKhamkOIGrTjPDV2SpaZxcVRHlRRZ
mTFJQ+HFKD9NeDLqzjfiN/7n13bgNoPK/d8cp3UASnLGwkrjuCLe5GRCVlVIoI9b
ZzsmEeTK7vhhepvG7ntJmSPVdKdUQcCx693mXwJNxjeHObkaI5JRGK/F+PsAzOG5
I8E69hXWyXJnnKNCDxREswhZ01o9giS7kK444mDqUCxhk9p692CcBCbKDQ2GSPXX
wk6KLnh4H8uT9FLiLjPZe3MZ3ma2nkOH2CeyHJO0/TdiVB6ZG40bTUTMnHRSza78
dYoqMGQIBVczy8SVozUfmGGFV5TAB+22Sz34AhZl9bkcYDgVidPqlsxH7ZNEdIGC
1KVmm+cLRI/04HYzkWiiGmnq2K2R+QF5DFQn+4J/4+Gkclf3UPLnB+8bXmKhQLA9
Gp9eZzS5QKymQbqQAg2NL7PP5P2/eHaEqwBSfW/oumjh8+mKjTud62oNjWOVIpMI
0vKF0F3fMBmJ9r+hcLOxgu6qkjFrnnA4eYs+cjD0P3t5iShuY4O10EsJWe5Uu/lX
69XHZZbUJDLW+p/EhsTyxrT4/FELp7AXijSpiAKAfnT7LG8MCDfwdt2Bnsj5uf00
IVlTBwd1JHuALIIVArUamK5WHrbaQrjJFfNlYfFMnUwI01DJkvzpoLDSoPmazEu4
My3kqk0cgk2ys4V6yptFjiLA/YdqNxcwNPvnIVveUUDSYr3pziio6w52Mq8pZN9F
wGKdc+Qnmil+B6nklDIO+5UeHJCu+3Z0k6t+IdceHyruExrG2R0WyzHSY86j2rDD
uSlyMQ4pSVImhXNXyKI1UdUf8uvy12cyxnOZgOkmamjHNfZnY9SuzpQKM0EVw0Xb
36kJzY0+i+ei95IFBOcvsvl9xwOB7L2kHBwsRPABpsQs2nUPMKk6kL9rYj7CKvLJ
xZ7U6drxqlce70Ck4vG8n+X8HhtPDP64Eydy8pQdyDDH7nXH6vnjlSzkm1oZsK4h
0L49VQ9ViDG3wX+6bEq/sb3Y2TAvmza9n1QjIYGTfgSBA7qS/K0/QnKo+u+0MfTZ
GFlULC2Y819gTFKhZoxsGd1L2FDcFfRWKH9WQNp46k5KZqV0gTO2Usm/8vKRzu5m
rxXY86HPdIe28NsdTiwSriaiY5mijinxWL3aVnr124gGWJM02K4PVkYhB/Gng8Wd
wEAhJsPo1iItWhWLq/fyuAZQHKWoi+pEyWqFti5vTymmNP4oCl+wAHlm35r+Mv4c
BZswXMKkpohaSeR7sxf+k2JwnoJHObKb1UrOQP1/A4p1SQg+BIsHcVrNFiAgB7Dh
HYtBI+jt+hSkUCVX7PXBDAiPDYgVZ/Clb8Sh3dchy7AJC+9bAhgScJu7+qYMjTe5
usuKxjipr4umdweW4K6b3dQb6uXYUJhW78rBYg/ZoLSQw3uJFFrRyfGTZ8J4mLB5
56D7W+3dNVDVeYl4brtU/nlPSm2xsNM8pFxOKSpA6CYyVWfPFY1Ogr7O81ECckXh
UODH9xsVLgE0FN8Gdt9w/2PayFfY8SoFIBfwfxxqO/39+NwFi7RRaRGBeQ7+GALp
exrBeUhGanDJL9bAk7MJ+0CI/UsVCnXdlpgI6g8Xl6oGVfV0LbD9CbwolOdamYT4
JC150EZluW9Y+FjZZ9V7jsk6+CAVG81W0b+IEwpl0b/5wUMvkYbHUiti89r0+v51
0J+7T8b6VJzA9Xuar4/jjIXG9P1/J9elr9H2C3STIQzUL+1nc9lDo51/5xKIPhNK
MX/XBU8LaVPfvuPp3vRhEYbZAfJIZeaMt5l9wP/I6vQP5y3oljUQFjc4L0KXrkLh
5wJ9GERbSjNzSSKTkWqF8mu0pC1p5+cCVi1NIqGF6LAhmLgxDDDPvz1IwC4rfU9Q
NhRxtPzmOny1Gc6Z83NmacMgpKgz8VuoY/F8oS+VQI8bMMjvG7mf3MCuBxXsEQWm
LK99+2SgnyUVeQgXIyTCz1CyVT3L+D+uhc1kNGI6klRVDeRVax5jdCaggZxr7h98
C04NU2Jpk7eA9hwmTcLAa0ebJrH0CMpqDr28o1vcGW23/+5q4r+FZ+7piUprzTyh
YZAfcJB5qVyEFKRHmV7Be7LPuaD76hC5P6JvF3ZvWf7D71IERLGEQhOiaUsnhZ9I
y94nyz/uRp/gSEovSnJM7nDa8HEr7V/rF5H/Cp0c/IRI7BcemTtyU8IMDvOD0DEh
elNqlP7p3BzeDYm3XVcjG6LyFrk/BUcfmlPsXL1YQhBjM/c5rMXrcYF5k2HVU2AH
gpfDKLmgAZQlVvWTA7//hTsogNKqK8fcRNOsFFKzR/7LbgrZSk38XqUA90NrHzdp
/NTxxiAyijaX/CTKgOsKnpqx+GO66RGgVFaZAmFrFjCkuxg2HMq6NdqIdU+fsRj3
M0ZpGVtPD6DCNFRZOzNOH0NvAEEcdHk2GoxOiYecDu4zxgaaPpcz8dmdR7s2vV2p
kEXWvyMqBp6/OgWKaNJYvln687oLuN1fa0Suv8WhFZw1Uky8dFLcbAPnfPfYSKWK
0ccGJoDvQ2LTCOoJ6UXZkYH86Lmucmn72J7r3N4Jwrbw4o5lunmy+JhBIQ5Zzy/G
kaWxq7vjyVEMZWqjmqWJf22zAyheHcLcXfPaaSFWve79yULzFsHY25LPYcrpgkmQ
5RlY9JoO9BqO7FWTrp4/I/QFurt1GzoSD0XkzhlChlSfdTMOmcumcuwwVCbeW69P
VG4JxP13dqXcwydQE/c4oM8FU4JD2R4pFgoesKsTzbplskIKAq58B3+k777VQXt/
miGm2UUBiRB6Bi+qHnnQc3bOi9peKHvpHVOcu7PLBJB1FFzL7RPt2kBcoM0r7ynr
CVLdYBgv5ddoWKLYDAWykpLgIgFxrmna/YMZpGsTiWY6AFj+8njjpm/I7G6T08sm
RvLDXbTs3q8S9YoBJ3Yj01nU0gPNC8Lqo/9aeTBpV4CImeAiPKCSbL7nTtFI2lad
Gal4Zo8bBJ6MpZyocyPPqDJptAV/hqjeFXc0lrwtZU8kY18neWXcGUjKJmX5m28r
VXV5lmIlh4g0ZGjvG0SKvZjJVQCmnZlEA+0t4RXjT+XdASCDb4Z7xunQq6lOilg9
4YxOSEddRNUl55ZrfbccAgqnkg9+Ettp7iA/79tEcZ4WEdtx2zfRK6txA9PUJihu
vpi2UfXptD+tnGGtiYhJRMwHzH4wy0wsvPtirV9X6wOuUYKrSU91iha4gVuj0otP
uPRMIHw2KLNmVIlyrlKxi+juKu5bGtMpEvEiEHFEm08HiF9eGFEt/u9FWoj1PGDK
y8nH0ac+9rUVY9AeT2jNPbZtaOhuPiB5rKvp0Qa0CRXu2UZLQFT2iv9duTVUkkya
nHOq5BTvge6WV04VtPZj05cHy+0ec3NUDVcfkf8Us0h3rYTo0+0AaS7cL8+8l4kL
U6qtTwwqlMFvYyMkqSyE4mE0OEEfWzfb1EsUWbe7T+IpfRGfiOjmoOBzHqZMPaJ8
kcwnwB2298/DVWekkDP63wwRdKagAYoIIqpjiFBs+cCdgRkIi2KU4LsGYU8r+p/d
fif4efbO/GgkahmnFIEI0/2l2eDmc9aILAuvcUEczN0vvy+fY/WL60+dYALaYkU7
zw1vsoHdTceYwSf0fiJH+gEH9tk8k+dclg4tzEsjhl0tR6c+mRy/fjdh7VIvfRvo
4gPpmlaC2OE/11rxFIR/VGVXe0g0VLpreGV1mfy/VqIs3UBOzIpalqHZ5mtegNWQ
XFO1mdz96IgV2LMxhrkaMNnjdkCToI5SPDinx54xNynXSwUIHTKWKUIW+InI3uHj
a0DM7NyjpyYa6ansVFfoPL6TLRtLgpIbtrTH6welf1W2xOxT+LARpkTXmHWum79j
dWxLa6iK3h4qOoQkmdQ1JZHjSfich48glH9J86H0MW9M5k85cSYbE7USY3fqIuu8
PE/nLMWLA2xd3Ig9Ab5kEAy4n8PGzwRVU7ipSWr3weTm44sYpFHosEpHlUku8IeQ
4WHZCmdEESKL0SPISwKc53PEFXZtnsBwzj4nm5OUH48HPP1uhtU4jGmwzRG0pxW/
dbajSpcFAcNK2+UhqHZ3iEefFClxrBrzcGZWnBrmxtc9mE+eX0q5IxE0GxbJFggH
g4OwfoGxLzjkmV1cpEtPU1C4vd850Z5LqHrZgNES+FLuIpuEd8sNNw5Qg92gEseR
6xWU4+DcsLgxxwNc+OPX8tbJ5DVIMMhMU+KFO4iGTRcY/1qYzQBWHJUxgDbEwdoM
rGl2KGMIqiz4zykNIFMfeh5tH7jthlXXg4duEjEpEdhqYuw3nhaIfGo/lvu22dHY
Aid1Dnth6+Eh8pMo5NzNwpHJB7HrZxbwu2H0BMvn6JI35kXKoawzwEriFKRewFKV
bS5DJ6jfM3wypR55wQ/DM+13D9MihdQIBgYWFA8Y77LUfRqfXnfOr6wrTj11RpN3
4p1kb4ksaZulLfTx+6UGmZFjom5bmvPTyaWZ6+HjDf7rdDS1UGc0SD/IQK6f6Y6X
jjQCqctJMppPfrV58IDpvbRkQ11fSYku4hr5U+CWUFrkirbLHJu2M5nGTyhyPpFM
ByorJZvPy0XFFN8X0kDP8bWUm3lxmUuYNObbFzU14Vr2IXdsA0SntMCV9oO/+X0U
TBI/HoNFvUOoj/cg1iQKElCn4RwbdVl24DTtER10chPAcZLgGa2odTioY4PGbxWh
wgaL0ejWd/BLj8epks99QGXppwzb40EqT2d/q3zTp5UQD2Z2vkZuM9NeFdB6AeAg
6WP5sR0uhLUBJm7VppLoDfSDMCtDS/vjfo+kf0yE+CHIjPPqf5yjymY7dBXtcmTh
75YUTnfkVP8SARoR6xoseOWtAZQb3YIbxP5dlxk/fE+cJeRASWs2ne5r0qQhNYZU
cuipiIMwhklulRrnGI8os8SgCgjwDXuJaR977ILa/6rAFFC3eiG6rfFSHycAR2sB
q5eg1YCvp18k2X0pvxrrfw4KhTMG6r319yBlJw1ERknCLVqSxjMoX/DxXttoYBqu
xAM5x7OLzam/3F47zGvHSSUPoXkfe5YUVmZ2RV1AxC+etfxtQ6ZDIBP0yFnEJEPE
ZyOQCs/xqOyjBvajUOckNbUO8LNiXb615ziI95EyP9cYWoiD7vVKu2ltYx6+nwCH
BBgsEcmaeTUiEmDnBrqKt+jwcui0xPifG6qdGJaIHayXkjoRuUY7iCBAY8WESkdD
7JckW6RQBa/NU360XDFo5tKaCyYWrdneWsuloD1CLyWd+zcus+SPI0ntmiDuWcJn
rRMAxiJ2mflxQXwmd0dPXAyLnRLcCYD3w9AnVthVJL5plQGB+taSDu+ySIbyC4RU
WmvK0syRCTk0QGNbj0l6ZJ9vy2A52cnFKyCtXQ6h9YiWSkh9ibRnYHyl/DmXzciH
rPf1GqihWH/2IIbhBqQHg+aRgI4dYDipm+AwBIN+ekUKqfFQGfP/T6WJGfysLgLz
p+6Dc86y/UZnBXeWYYodWjJCMw4lWrh1E1Oz28wE/N82W0Iyvv3t8lkZtr+OgXlT
UXoaat2olx3EOh/GpBE/I2WWOyGwWSxhvm4YgcG85KJJmvWbIRt+LkoSvyp0Lbtl
WO6rV3s/ZNgPwiJ+j40ao+tJu6nF3njZxwPR6g7nKtISx/UNo3m/R1R4RKuFrJ+O
lRouk0Oa65LxDyJ7FwyjGmJga+Hlvo5KAI+8YAI+rknG8/4bdcUd6m0uQsIdiaVF
6l3s2LFcJcu9Kp6Hn5JY3h0hLR+UozXR+uJwQO/OE9Qh7J0YvKArRoIGjM+nmGM5
wso6EVs5z5WAztlQLSdOEspwAPat+fx3xBnOh+qDFnn6vzwAujYJN+Vb55sOJL3F
BhnVLMCQKYY5zy6JLlP1C8s4cTpWA2UElP5bfaZtJMpj0AIkJs/gXV7mDy/mx/W6
UMz4F31v4cqrDS7i/NjPlvmwjh1nwOI8TcMbIq+04kxRfNITRf2YMVnUXbtvPWqX
vda5mz8bHtjLXv/0fvsWbQOoqdWxPqDehPcTZRxVCplWNylVwWIhG0Z3r4U/0NXZ
NNBgej11nZhLkMXFJdQzn6P0PGKRz4Q92xvUAakUf1ISYJ2oRJXsqdYEpJyP8cC6
YRAkj2F6dtrWZC3qG2j8a9YN0WLuPiNdlkmRGaC7TCHHcAF/AlTfHYv5KrmBvRs2
IkdbvKnzEDqmPiVMD7ihRYRtgOXd/PARxCvt8VLLeD3ciEz6pChgUfMrTsp6tAkI
BJt/YFjVa5J4rtTGWFOlsrhjieWy18hwsTcc2UHoZPKN7IyjwEJx6p1JDqWufh8i
JcdxZinPmzr+b4lNbRsrWz/XsnrWiP9Nh6U6ErCOXtTzyPoC/q1O6RievZ9thgc5
q56CbRNMs0CJmIvwE5gqsqni5GeBVukuuMGtwMdetDVxk+Ls0iYOlgP46mHz2c+2
sYKwRcKdObeY+6n1jCKd4TENMB56U3NQ7nOx7K8I3ECd8xoJpP+sGOszbRi0yYUN
jjxVW8+XfDf9zZMr0I5jJgAm83PkEx1ruU9xLf3KeV+/t4Dw7rnULK06cVkOB85Y
4i7RuMh1lByjbSsDGyJPmIzbHW6ajL/kEwg1BnHwsQNwAqZ3ha5GGg//9jMCf/Wy
F4loGRlHzUmEXhvOcKoZPK57CScSH+9UFJAGyV2ZRvv2ORgXJq+zZCHqXdlu4NOP
QOueM9t2jzzwBs3rgmkBOOBWMFHFCTwAm/gWY5fp5v+xMUbCkF5h2S0bbbyx8uKR
eeDEW5HwvinaQ44WplkzfkFg5za3BgO/KesPVtHzWbvb8OuZrnCNYdIJriVVt1si
54AFRhr9O5NVQ5XynyVtE+dxPNeUZLwciydx7gkRivIFETkTdn6vlxVER9eFPsXq
URhHZutB+abK+IPu1TxxIi/7KTzyqpRhWTOEBMJ8CLLXCx8tpbhJn+UcGYcNNArG
3jySufEjx2xDqSQxO4TGEr3JC0zZbHi/06PJUUImUoWmixr7THQeegtY1jx222e7
ofzWoAtWMYNfSnIHoGTr2pmIxRLaNJ0uJKexSnLNJvSWHt/603DG14hHpsCfgysF
vvPx9sdgwGLKZihVRuH9//2pYmrwHZ3shbpjIFVCqMK8OqP2I6G9Ql+b3IA5ff2i
J4LrFLZRuLWMedrpQ2aQ9yZ4Z/USwDiNBe1hcT1zZTJHOFu/HrNcxvEDNkxxNgfy
2aPsKTlSHPbjRbzk8zl4ro4dpTTlc6egGK0ndMl/Rf+GbpXEMY2/r4rUx9CdyLPd
HlR9lPICwehYoicbQtFBJcAB149cxjyFaaJ4UuWTfAA1JX5V/qLDK54oSyEAVTYR
xu9u/DOEFgIQsmWI8y8KfRnGXH3rCEuOI4dih8yTMCRWGF6Q4NNUWpumUj5H+ZDa
aRcjBGZEyeMYSzDC71AbHwOCIWDblrdmUFIdhtIHoO6uOP+RlQUGYl60+SyWQLnd
v4fkKASUr+MRGZ0fOKy3C2rzcUF2TZCVLEc9K3X+Y11p17mlPJS/TN5BqFjznI9j
rLEdA6eiPL84zNf7N6urdSeRL+ViGjBfCgeuceWwJ9BkVtQGkTmH+6FgV/xgqp5C
MrYiaAEwfDp9NdjEVp4eJLehwwKZ/H+T3aBQJ0SzAXx2jjFfRJSEofnOrPGcc+Q/
cxLgHIrsJx9m65H9imC3tHzZ2JL2+f4kB7faMoHsMBtcgOsOaFpomJku+el4Tt2n
giLD8+zQSErciK4oZSIBgNR3kl1Sg6G3o9fDRXKss8sGewEBg5c1cvVHLozWlXpo
lirzZxexSxnc1oSu4DlyTpDo5Uo10vBiUMK5X5lg+eO4BtsCxTPH/9AJ16Hz8+qa
tnpiMpRn1wHMHy3czTGG5MGvjzjNnmJD/LBbaWkxCO2FzQ50TnVj7IPxIygQXyAz
Eq6BImS2f3fv/1Tpqv0nm4WS6JrcE/0efHQa3e12FaIhb7RlG98VqVgCkYx13NXR
uzA8+QL8ozv2l8gzy3PFtdYHZ8iPmB01Q/Bnv76S5crQGaxt8KIbGMBFI79Jq8JQ
/y7I0DHoTVZ6i7BW8CkToEAMa0KXh/eG7S6lCO6iaIaO0Tov5CaZDmBj79mQluBN
9k549A/jP5RVG+u2pUFipa+/03voR08lw2+zVUhYPO2YfKfRgp9UVnftATf6gq/T
aVs8ODTTY04d3D7w16RyYaC/b9TuXwRBpdStzzRHAGk4gQKNMz69qGAP+YIai9J7
OAxF+zN16ZXwxdQUzE0ce8DUKnPpNdDrkDTioK89HnUIU93ItaUxSFnVusFhEOHE
AUXgPCnfrwxhF2APIAEr5ymuYvlp3ORtbG0e/s2eBdY1wU+CZu02Nd6WzaLG3tK1
ofNW3xMC0NV3+0rrElwd2XqSALzivuf2xBPEGBI65BvJRNk/fAAthPcsaLTvbfzC
e2e96wgpN0XUEWLM2StCjxB/sw06j7awrdWTYoaUjn2JGrLQW4oLEF6jXP2p/bWU
Qk6P6kH+AkSGCYpEGhu+QDnn2M38iY/+mvgqu5yW+DhLhumuKzFRVZNGP4BsJjSl
ymmU6vx7kJHihUJSi1jWlCpz9cdVPE8Oi3waUtKvRdbug/9uCiZ/SMElahoM3At4
+Dx6IKXXTGAOULdlTgkcsXb9GuNrqyLxhuwFOvkgp38acyGeyfuUvkhiPxW6bGYG
vIfDlRwAvZNLkrTNSptncXLwgE0QX5j6BTPWke3JCEMHczw2yIfbK1t9TfRa1Sq6
0WCl+PBRwgrVqFjw42VyID4+Hzx5UgjwlYhI4FfxDw6MX5DEe1zpNBaaOqCF9SHl
ZHC7FX3vwoDpjIudkl2MED7daG4xmec10wqhdS7sbWVgTU6TI+2z9T4Nr62ok2Aa
7kww/WJrTs4VbZ7IVXn9Czw/lUwArz6854DE7zMUugS2ZJgQKvHi3FjCmVLnIAFA
ol1odbNHGLK7BUsdFWsxHfnoznI1tQB34FYoRKvmaZLG4DjUzrHYOxzTmm5lQ/Il
v96R5wS0R/pxM/NU0aQEyNdbMJ2TPK2ic44/mO05LeWd6F6q62M+RHtORygSBAzp
UES5tuNiM5iWdgvO7KvrPHFLGNtTJ1pWc2pyUW1s74nDhpg56AqfnmgcaamoEyB9
IxznrKbv5ikyESj1J9kDSXaB103p4noAO5DMMKp2FyCG0js7ZoBzUCFusPNzk2iZ
IscNJJKwO8cWAgWerAU6AfNsAjBXdSYcJSSm7G25/MFO3E9+HtFJ7h6hwjOPkR78
3ViaRl2xNy7bAA7I4W+RxmbFPwHd5lvFhnzyMA1IUQGHmYqIbUe/pRfrwmVIS4SB
oYX7ZPUobUZOqggs4r+NlyMCDtd3p07iYEUjo3s04ZuYFC4zuLSBKPEosXeCiGSX
MGHvVn4/fzX29ZzNwpkqrm/xFE9wk57GuGM9HgUnhPRHYNpYaTmZxtyLHfVRwRfv
f88wmZvZmWbWgO4rxUdDY9RiuEnQkFGCy9maaTsGTLOZGz8DEB5eyKQZU3OH2Hw0
18AemhWegrIKR6bx1GeP8kz9dBe9LWFZqGixkM9gUK+IJhq+ASaXXWFCtwL6HN7F
+WkwEWjrPpXg+3kqt94byMLIq/wAXfktOuNd2NaMOmihmSHz0FC1tuBjT6s+Y1iQ
MmLkAkcR7TXGYAtvTy53e6vvAu4CHFA180eYdg0yt0bYdl5cDlfgiNL9tg8DIDhz
yEHrDVNMvgzEh6PEphTJ7HWPWyfsc8Haa8oZBYmYXIT9jPotkxxUb37cNcJb9enY
9TKwL8M1L+UmoKM9035NeyCQoUOzvbVPVrGseVx2YHhrhSz6UzauwxlYm5+xa0ut
wx8d6YLz4CI9f7SMf1ScXkc8Mfumgopep4aA8Zzm+lO7/oD5zH7AdWwiWmAB86IU
FDWp3D45HSjVjsKRDoG1m85uyoG5I/ZlOS9J5ohlZSimeWzfWDWYSHZOsqGQiECd
G0funIEcE09Ip1AQXkY1cxqDb9j7xrtXgt5HHxh5V6sDa1VA2q8RL+91cWQfUwzU
CrgyxhIczaPVsQmkSjcI1x7RtLfiOwuJRYhjEOIosJT1nSoIA2ubKXXtDntO/Xdx
X1IVWo+jZ2aef70hGIMIxCWHBNaDYozUuuOyhCejQxONM55rlIX3dYsuHzteqvXs
E5fYUDGNgJJ1C2V1xhAjlL7OmVRzxK/jWJB8RO0Ro3RFV2jKkAh6kkBE3Juc9/M9
9qtveDvB2MdqxiCTYlofl9h2kOuyAMclO6qFGgVYd70euBRefSYsmHcq1yXKKt+b
MGXXECyuKRAFq0FS061g+eDKKXTfdXU9CmIE/Z6C6YB2TA7zWZlSlyJY5Vnk2iVU
+pkHjjsuPbP7GZETGx95ab9GxCTQPmMV4Y92KLn4YCv5sd5TduzofOg6Zqgup8MY
iRlnhmdNFw6ibBbJqZM/SzPaDOmSoQC/K14esgIRqVnN+PTHyL9L+dGDkt5PYfRF
LTr3IvSMc90Tu6yTehDmg5ZISiZNmS1JzjyCeapWu+VgTY2cBR9v0eD/XyfqZy7p
ou8FwnEab2qxhEEmi+EIQwqChuq2LMXu0fcSFl0ZHcRy+boPmPEl2B9fCwp9QdSV
KlnBML5LWSlmbR7UqsYviADCnPiLyj2sR7dTijMpXRNZc8vlz6ScfUXBFIq7dj2B
vL6GwrgN2h2VYeckAL35xdXM87RIJOWWF1q5/MiCPvmOnkl2DN18fxAKukw6nZNB
VG8YGv9/8DBfQAzrq1LrsXu96voixR2kRyronl1LH4jEq39mtVGsoEJtK8awbxVw
PlFUK09voT2PbnJr0d3TwCiu+AMJ5yER06CVUAnjxrcndDk9d/xZ9L2U7Y6+amG7
LFl8ZNEsPQvs9L7EhniVIDLXSy9ha76FryQWREOsi+GgZkCi63v6eqeAyOg6Qmno
C1cO5oWdpdoE/BnsUgDJVMc5tOTv/Z1GLi+cEJnk6CZbv5EwNYUhsk8xa0aTOmz2
EUaKxNpmnBbM0rX9Glcwsgbkb4MEjbsxhIGgfXKoEB6sxMdj4xjuci7bmxeyyrY0
zAs4pWE9soJ78N+VWNMOiw92wHVKMjsiq4nw+xLvjq5pnaPDo1sh6yJOdx7tHcUO
ZNxhDMVcPtlfsQs0dqALox/HY/vpsSykcOmnBlwU6rsip57RkEoREPoZktgnyE3L
pgtzfNYVO6qY7Pp1JeaXWyr8GX95EvDccK1ZfokilHzo8JuxXdgzlKj7SifZZiwv
sIJ+lhCX4+Yj9GgdAOvWycOg4/Q5xctO6Y6uC6XCpvmXiZ/6GR4qRFcPqoZlH+2+
ZnB86xmqE+8B2UeftJG5Tw5Ysb6JpXqdIIIJu3PCpH6YeO1ue22SE/1kQ+SNWlb8
sl+VuVjAUuFFXMvP3mjok00NDTihtTmPXW7f8LrDOvB3p9MlIUtujCw3J6B0NzcI
xi3EYpSi+iT+F7RG6/flCxVb5VAsWnZ1yYqKiMyc7qjISk85td65PzBz2qIP8lE5
EAkHkJP+9GahnhNKJ5MUSsVeKahWP8BFpfTh9HRjpe18AVul04fnc6jW71KM3Q+7
CSleMdcnReKukEaSD8axwhxWbk6LXRfj6wj3HJZGCM4keVwldqpdWstG/o35z4hV
0qO2FrLNQYP8rojT1t//07NXn9o1XuAIPe6UdIh6vAkJCpbuIhMf3NRqDBRuxXLj
dzdSMMknaSuHiIZ0BnXbM8E3tBR93vq6BH9eBn6cKNCcpkLmM7Lr6W2fpYO4DG9y
muvusCIUtqY29CEZ+tTVakras2r0GxW8ywDZOleBdPKHJbVPP2dpPcJw1zKaVSpp
HuEgTe8LhlQ7LPSSlPez+NzpB2e9Tl9LBi2YnTFZOriZFOjj5pLpR2aczRuAQn9Q
rBqSW+q8wE1rJV/hzCjkwXhfSBPLhOMavoLk0wpUeoMItMtSzpX+00JLoPLcriKX
//4oEnFdJDrPzvbz8iAq412z9sNmWVS9yeePvKiX+zKaifi64cChouDaW7LYsVKg
HREE2EOTlSnVXycGXAGiLn1Az5Cj3xiTxKczTh7V1xpmVjjYlY7ABiojv0n2AeuV
fEeOoUs7E1cKXLyAjs8qWu35HRg2IWhTBLysxVpna+EBCPmLJWk8ZR4ur18+kNyH
9IT7ehEEaAR1KfCvljwfq1je2QxU18BWP1XNt6F6/eXac9ddEyBeOcfpHjKr44oI
FAPHiA0iHxdHvBL6zaA+p7sXN+5IAOMz2oAV5RVi/Pcl3ZAyCVKiFZtGmN7U6uPw
qF1K5c014c8jM0Bs0xlvXpj0VCSutLHlGo4qLOvSOeCxBM0Hrc4VBbu2WSaAMQr9
LCTJmtkBNd3yAhXbu1M2CvJqoYLrGVFLDF5UKjNo3mQEilAXHvOwQGxjZlnpsAmL
yr2u4nguEeMgVwO0n/dMpO/nxwWy0s78Fdoged8BMTDQ/w4ubk6pV7D/00QXLZBJ
l3Utxb0K+6WC96Md+KpLnA0SFn6rPOwoJzG3rscyOgw0kzoULA0u9EnkbuTJh3oy
SIb9jX40ipT6024gNOARFJM0AiHnoN1JdcRUf33LH4y9ZNYt+m9zynsshgftBjmD
Wf22aW1GsU8lpjcdsQEgpG9rpF9a9XRdirjsaiVp22RMJiKlxJBsJTq+kJQjLMbW
NQw7FlecvN2nPpLpJ2wb4EhjMdFiRJNoQaJVWWYnXDMyOhksG7SahqXTDtNirQB7
fJc9zCH6sgrogy8k3iob+3pb4+SB72a73KySmBFaCiOZnnoqeIU+/oJQjk2EIkmB
6M/UzNhPzBkwwMzSpZfOZGTvxHhoZI4/YREzJuNz9YmOEL0cdZkJabA+W7IbvNyr
SxBIr2IaLrk9modGrWQHHCnx3XM/+jrRuXfad/aOn3Ffa0IvKdbvUR6KsGcEdVBV
YUwSi1kLQZ6xR6czqfOke3p4e4clbA728LKrCoTi/KCubXEra8YGSlBWl45Mk4Eb
xQrQBN0crjGXxLpqPpFphsaR0CwuiUY78+Mq4umKr9WwmP700QbjiYAYCqh+pBTM
1OGIuHYdabY/muzABkKFa9NCGQy362q0HvuIMx29+PTDESCbll8UL4KLsdZzkVGv
1SRsSEAPguIuQ2tcQkEcBfvTG1emobDdulF6ncEe5NXB2Hz2iiBcwSMn28mbIjY8
N1TgQcW57yImixHtNeDrip8F+a2KyzBRf2fOS/wFQ7Xrmf1uqq+3MbN1gSNF8MZ8
HCTHAKnoy9/86edb0oS1gS6jzAEl28Tx/cTZITgo9qo9sG/2wDlhuRVsUL1CaRxK
qcgVw6K7/KEiLKosg++0oyvMn64rRU9/Mxv1jZqbXyNMd7K2QnPX7eFVIQFxIUPb
029zarCtMXPFHcaoB2g/cjTJGrVri59Hx5BR3HVxqqP/f4y17/bmBfTIIYhEJquF
J0I4G0ycZ1/KILpbuFnX2LTDySSPDxQNhAY4vlP9pESCSjCo+bltyv/EXWSigMMK
fcqhqyBV/EySdv/zqSXv1wES9ANikegkfZ/B/n8X98dfN4yyQ/WDlOWo7RsHfPr5
Ce7HizCWgnTc5KLLafBltNGRfumdXX0oXbnZDPdqQH3MbYWz+0X4YAAjhoNTVkmW
iDIrojFPkgUrRAUHUK0x2EUIZdfpFSUBKwCXnwP2OaXHhPyYS4N8L3CT7hgNEhbM
hVs70s4s30XMbrwgG/qT+6k19HaEm/rJQHdHUbJOMEVmHi2UfjYXcnFdWGr+Ni+5
G55/qYeotorAxV7jFMis5OjkOGDNEgb1Fo8xyeGI8d/Nz2xM0fRRN6CjcFndR+cB
h15bcUsfLhtnM9igQ1TiMCwfZz2bU0z84zrQqge3l14jY2rLN7apKezWwyh6k5At
LcmBP2bxgtKZN0AoNRhM40ze3tQ8F4Llv/n/zeH4yI2MZiqchc2N2dOvwzBDFR5B
PcJBnbYa0qOCrJw2nlmonaRO9PKF3CoDLByHH4vYtvUr54NOgoDpSfXidBytbOun
0hwpuU4R+0mGpHRA9fxD+la4yTTtuikbLzr8YB3+WneIhqq6RnmBRBLoAPXEjmXn
Xsi60JKOH6YzROtK6NmDKJR7XQGCbwP4F66//9EdxbtXdAF7tGojgUIh+nULfLKC
OEPM+HP+3ndHJ567Z1bDAu9OyWUovrz7e+yGX2tt63f9czS4Wp0NjW1f2MQcP6l+
MU31mowIdymeenbQdv7dADoV+Vg1we0cQVbl8CvAzB4Nfjxpj6v+ClKxAEWSM23/
WtvKYzq6feIGx8kAcovT9ebgAQN1+Q7+Xc/sqZC33/rGj9eGRFvZTJA3inHZDr+Q
8cKpO92tAyi7r0Ss1m4+nSSxwFD/Bx3cIHAFKfhBOfdrPSP3YLN1c5Euq2qylH00
8qR60kdOwggXOMvOvl+3X/MeZe1imtxBYnJEJxo2lMYbkDkPRNbz/Rr2suUFpiLk
UvOHTbRi3rXgIv69IULfVJX9HUWJqRnVyRLmLvmTC6qL6dJt0d4JKzYEpwbf7eSL
tf/xVsPM//rwo88m1xjYrfEYqoDk6q92bXausefxXVJJpKZH0TCtxO3/kPdJEuLn
8c825jwE77tvjWMFYJfoE+We1T17fOrorATY1iQlIPyuvYEcNJkLsJ3ENi/i8MOy
CxbkwgI1uLnhpeK6Es0UK2TnCyCllu+8nmKupkTF2AClA83Sg6c2Ag9UGHbdpEwJ
U9l36dRLEzN4cBHI77ACD81MEVzn2fgoivQ+6txnHYGOmSxRuFnxlAS8s3lUs8QT
erEicT+aNbs1kdj9613VRDj8T6+h+kaP3LFxQ4allrkWqK6uJNG4NH+w/U7SEq1Z
NgFfGV8zWdhfQDIrFtPehDLmXJLYaDhBcO02BszKnz5nWHXALR777lwYG2PXDJ89
lqOOLiI7tk4yj8N+Op/tnDKux2CUzNyMgkwP/qZeIuBk3oq978sJdSbxX7cicGu1
rMlNY5hFskSTsxdb6vIjNG4tARz5MaoRsWRyDPpgoPuv3X5CRYghKotsIMtlmLQl
no39YOiv0AjxkrRP23Do0MMCIgYTieNlSiRGYzssAnRjcIyxz60NpMhz2sVJirCc
gOZnCRw5R40FCXSPa5gSjaypfALCg6I+zSsf3G696CMPWx5E2p9n9fwsuhMxV1xa
WKsyR4naIQXseaYc9mw2umORwfyH/zE2E9N6YbqBJ/pNcMoorbcxtAe0Bi4bxokk
CSbTC6SjcCTHYNT2jEtaYteFQ9Rt1tCgbI/Ar3VvvutDgCpCg1QYTkWXF8AfXE1n
6X80I81fYukjAMKSu94aAOWeljh2F/CLPt9Idzvjwj2vrgDnO13SzC2GNEouiOdg
zKl4sRiAXO+oEdf//xX5fC+Dpuj/GlY+Te79Tusa2sJTuFyXrkK7uX7Ck9FWDe9T
KkO5IfIvo4XPcTwbo4rNt7N3MK2t+63HdrtcRDBGN4phWXMkPl0ANtGTZ4qHYJh4
r/jrOr27lhNcQAkEt2ptDAdemIafPbWR9z58tv0KdqmR+XdvTK/aNYGuhfVv8IWP
cmGfLnK6etaIsd6HNZQsjUXhMTYbmQC8UIRaUsRmY4rtQah8+c9Wh/WhrbSu9AbP
SqyWWlOzLXSJvTmTPW/Qfpuf1T1h2D+0JPv+5u/EbrPgezDbwRqf44w2S38Qq9X7
p5Q9nIB4jkGOh2xMdQQ3K0cOGVKm6cKfgGXODeAgE/L19D8fCs4aOoT2WoyvxmUJ
FONH4DftpGM5H0HRVsvuUzGK2JaJSX+Vj9Wp9+QQvTFOC3ANshLEfx9+J2XzCfxr
fBs9yZCEzKbXqMGxXMQHKjv9ad7ch2Phc++Dy3PWR5ZFmMT96qQfeeFNA5kgh6VD
vEDPFqVMiOea1v4W/J04uASSnN5lClfEe58UHdxvolSk+FELaaTsG8xC6xgBm050
FE8q71CX60xrMUJszi80I2O2ZoHd/psj6OyslPESb6aDtkQqNNK7XqelBoPnEMNj
vNiRdAjzwm7SD27bfk3e+tO0K2jffndatPiSiqpQoSf9srBPhqsm2Im/sb63K8WI
PzTFWcPSu0Skz7FxwHjPd+fYOjXiyUaDLaMV7lDRJq7NjMd6d+fAGefN1MQx3dog
X50+KFqTk7hWeGWoDy1EAmulj1ovAl0/XrU1so5puw29wlJID2nnl0opX8MpAVJ6
1cDPyzmz7AtwBRFY7g0/nCmeEDUojtpJp+ZTPxJl3SVtVZveJvJi0fW1ZXIQ2ZPi
HLErC3WfMtdLfi8oDR2eSaRTJXO8m74wfNmZ63ps7AXmNAApaNI8vOmEx5fSPlXe
ueWj01SFswXzhvXYiY55gfNyKthphQ/ZGkMghL8iy1gFIybeTWrZZP/aG+GBakME
xAk5jYHniEuGJ+eITLSyDYJhP89e/hBXsy6WyNZCfSgEjp4KqkTlak38ROdaRvrg
PmWXPC5GBtMUNLmWzKGkpr7PI3KCUxqx6JwGvh5qoDu2B90tMSPqqkg9NXQa66vl
5oB945P1jxQhNFmikQc0LDQZuE1Gw5ODmnv81qp/b9+szOfXT2UgbjdvzePhQEg1
10mMqGdoZQNA6IdeNMSm/6lrqK3K8MWixqPQKstekb/OhfFYf08E4fPm8B27jNSg
97hyNJh90UKCBw2c6tTW5w/OxGOp4Kvm5RgCys7dlbt0C5VEduhLbCvzXM9tc5Q7
5DWwiQ10alic0Hmc81yjyizPZa3XSGxrNum3e9Hu2SdI3thRhMUua09cpyAS1WWy
BPPcsxLcKq6V2WGo3tLGY8kpFl3F78p1hJELUqI02kqoObwzyUpG3LLMjsWBajIb
9R8y7Djwfx5qHFJN06Mbc1iwCBiL9rM2CFwAyydWxafCpaAXDWWRp+vL4agR0oYY
CYG7dqArICtDXnKCrLhafZT8rG8hZnSbM+OX0/NIT6/JeofT9vviL66L09+M5/s0
lBuA3Qh7G2JJlMtqs82PRV3WAjGIQWVU2BK9jaBeW5rTYdaooYRoKiivsxMFUHCl
dzY344I4XSef+ANhck3Cq8CXG8LcGHjXifrE97eyGBDHH6W5t1ZhjT+hSUSnaAj6
2uvfdJRaIZJ6dXQr+3zWIGGGjLJPY9wEXR6mPLCL8SrNxcK1Xd+H/2stQTXR4LFg
s6KjGLuo6UbCLk03XMae8n5eUykCcGy1M677DPZtvJYwU6gS/zDCpUMnKVx0Q+rz
KVIF0jQO1Ec44mbOzU170pvu1ZIAEz5T/aUA65Q9rzKZa4NHGNwlbeDNnstElQR3
FZ78ftuz/uuvgzST1DZdmIUyOLbL+/Md7QVP7oxgFcxCNX1bgqZRlxwvSxRxLn8d
6Emj1aXoRgbwPQmZFyEJ8MB7PtTVjAh4beegxr3Y0GH3cl/jq+TF9tJeUkdfFUJ+
rTTx5Olt4QJuOatvFCiI+ebd1yLDeOaQ09UWt+38YmOieW1kFQp3bBcj2T4fUTtR
PB5BlKfAqfFFtrqrddB6Nc9RToC8GTEdTLs22fWQ+hpzpJy0lZy5BzUPc81CMr0I
5pwgJrcl9lWpBbjK/SmQdG+q6+7oDNK9NcUgam3Npaq6viTm9hBCrDzw/ERh4M7j
NTnou61fap9QPyK+aiPwoAXq9kja23EyxOggxGbyCT57JjtJgi/gwOtF28Aoezvg
vJf6f0LlERcNJ7WRYpWRnkAAVuQr+chpqG1ZcSdzdPfv4KHK7gcI2VPsKWJk4/mu
fjr4bvnilO9tzuSGTceGsXp2WCkbsWMnW6MGQ1Nuad1NNLGWBNkfoSKTPF/qzj6F
sHWqGtoxneCLtEI7v8f9KfKlnhjG6DYmqvv7vCPKw7TExdO8pNJCIc2FzSD7hOA2
WuTwETa7Q2U+Ibj7blzROfYvV9TBtGsl3ErqlkbAFGqW9rBGRWLpP9gMg18UNigM
eUQxI92/ZquNHQvfoxYewFmhnFt8TnpNVqbzBgZuGJzhPdFIfdDx8rY9gZhNRRJ+
Z9+KYuMPgvH5BegTizVkht8fG2EoC9ES2euL/Seh7AtBRJyMtjgvKnCJEtH+f8Pg
RpTpOLFyzSzFnTz+USpRAaWzcG/N0yp6PNI2ZYWUQUL37ubFVwD3xlZaku5NN86g
tZf3PnsrxFIDsy9pSQX3ZQtvKUdxViE15KC/5wuQy4/5x5zC9mFfSZ2hRW4uMgJF
eSb2LrCjS1tbN0m85STyWaPcIwJJLMv4S6AxCoPaFNm2w4pkWgcr64ByH3th65xN
BSEQkFhi1YDmOKDVh0JkQZ7PtPxsE0VdqZF9vQitDBnp2NBiFBC3vCUct14g6iSk
a6eE4dEakVlpKh6D3nU05shhkVKI60g4ibZdhvHGAwW/nXUCCAdsJsSZBI6NU5WS
AMK4R9NFtmMSHHf1huLXn9rplHH1FddsXBEsfpz+sscDCQ49AwkRl2P/cOlZeAJ5
UraIfTjVbcMnDNVr9beEaCia7t34if7RaT/NJ5cEKei1LFFxzXM1N1eKbXQcVLoq
7w1SFAHE5Gz5TsuJkgw896fFdcxMV6tITcpAAujipNRItX0tmyEI310Ig+OOEgqr
F2fvBbFoCLIKV/eJckM0ez8vtUG7swqrQywN/sp7spRXO8m1T3M0zeUCa4Suki2K
OJ3ODF85bBfy4uqN19YzekQcgls78yt/gZlB3bxc79/m6zL+OtoiuvNAYdGf4Ifo
JHRyn4BFU9rddcM0RNCUHzK7zuL0xKMFmLfgKoOU2dMWpYpJpGmRLUM1/IZD3oNQ
9j4GVwMudZ/a9ZFQzeAVKFrYyT0cVIPeuZ+eMo3s6II6PxY4G9MKXedk+S97vgmB
v9YNe3c+VnhOSx90U6kpOuUKaji7mm9YGfPxa8gdeHLjVCBR9pxkUWOZM1O5Cgnn
ya+PJkiU2eyoWFhsJkqkN1MD8OMat55kQ95p+nCW9oWU9gWRQ5P0srdATJIeFMXB
sKZHJ0kh8IgEqugeDUBQBhEnhF43N7m13AgB/6iLkhAIajiAQqE45aUs4IGY/RBK
9iY2tukDIkySab2Y/YK974n9ZxbKtiQbn2XSnkHIDPtS30lyL1EylBuRdXqUmSYC
L2whK9Yv3iOewO4TSxO/Vnyf4+bNWponL2klG1Q5MlpN/SYr0HeLwdn63hNrg954
cIX1yW5ITb5S5SgiQC9IbiouYy4v5Y/jgSfd/R7sFztqPGAGimwFRO6D8Jo9lbQF
CSSkyqZZ08Xf+NIOwZROwUGxzHP46FfFrO90Sg9rsRCa/lBj8YFQbDO7AtP+UQFZ
3pToLF/ysUD6r77C2D/m0bRJbTG4DVsjwcpeAqYD0tIq3V3oEn3pQOGVArdgDwna
b65u+vRHiooP/cPI10VAwuU/wz6kSdqOnU5LuamKKrb7Y08xsY32g+EEtkhsV3a+
i1/nkGOK//GO21GCwX8b1rf2dhcTIvMiS1/4p+5qlveaIcP4X8ZhreEvK2Ua6MRZ
8BGHzbK/ukbo+dBCepaQ1TaTqm70tnmQ0Wg7pFyTnGj4b3Ei1LFXdLftGeYHJh+H
Ku8OYZKf5lqSuYE7EVaUWh/PWjTF5jZjSLWQMb4eVPRbGzFtn+DYcq5UaBeXP3Wh
WRSMQDCo6q5CnbnKkv2warsysB0vbfJ12UaMSBguMvZL+wWupQyaafyA5tcSV9Lj
a5pnxN74fOG4rIYfySazpo7wRN2vVpWtyzb9rqLCm/Bp69N/NC01HsaJYlofW0BP
D5ltR9b0LJib9Zrs3uz7yL2RZ60F/tOIYqZIUgJ70VGJZqvcB0vt7UrKaNnQP+TV
qWQq73UCX1rLgOWSKd3VmVqfr1shJQ3YZz/Mf81+Ro3Abksq6aKjSfciQtJKS60p
X5XbgdaPgWCAmqUiisfwg12gzPxTqXbSezJAAfP9iyXIn4eTc7iIHn88AKOR6muG
/17eRxrpV5dHMZJva5EXOyTjijLi7SS6U+7Z6jhfpbq4lidJ/caoeOeloVXRsEJM
VF4wd4MmFs0HjSMZeTsYakxeaNj9izlSJ6Im9eRvTD3qLeprENcbyzVOUOoJy6RO
boB4ctCqmmiXFLZMDUdCAQTy0K/jpV8bROZp9lAypKxaW/GSKFq+f7RxtXD5c9Om
kr9f/zjS8q8J/QjNMxeZNx1xqC4Z4JcsYJzaXrEcatFOdFnIeDzC2oqEWqCv/1gu
mtKvBgw5jBs3kOhIERgr213XuOvLVAdfiC7ffufYcq/b86wgzt63Oq9d5nJ8Gzrx
D/+Hdjkw3dgIIDC585GlzbSQMNVQ8o8yKjazWQX7B/j4PcCYtgNg1nPzpD0c/OvV
MIJDwcHHUr5C2DOWEeEoMA8nqkPzRwEaF2BidLrBdyeBUCzTogLPolAFX37bHdKd
/5qRlSo6ogipdEwIBjGMvuDcXYSS9hPfIh+T9B4XAYF+dTzvIKvtEp5bbfyBXUmO
jIPrMWCEChWZNsIK1HJlSeMw+AAG/ig0MHkOBwfaPpgDZaCd8dwN5hN7e6f5CrnG
v0j4Fl3RteB5XkT1Bbp3HgiBUq0SkWrVeyoDPfZv3HIaiPyH/F5KHW75erbUUedo
qTQo53hjBXmpRasu6R6SplhTTYj2z3/+VQyjzkwRpoWWw2PPKp+Qo+tTY54abe9h
3e2pv2dhc05pGWa1IyHh5rXl2413PLPLmfOQUPi4coSaqwj+3FObprrD9eRsXY8N
5Y3ZclITR9ogSUpj+G+7yVJ+witSx1zSuS9/4qV2r043ubS5qBoLi353/fPUENN3
pJz733KHBvG+Q0i4JE5EX4J5KD5oM19RkEkO7NhvyVUFnpgiI0eJ3D0mjv95mqUP
Ds+bynHx/Nf7dLYG/hOTmGQbea5EDTRjBUhKocqqrRbgcgQbp89BsgnYzqdxMSlE
p7lQbalAIasFULEtgZR2FmO1Jc70nsHeFudYuHlUc+47ofu9njx1Bfdd09ynmFKc
i8dLc+p6JV8YUio+i0R4/irxTtvZ1fZHKZ8/IH3WvcNoclZzYsmX4f564VFmxJTA
QNFsa3SSemoTsK40CQpkp7inzZ75CB/qeqg+ABdS2wJSJQA7xsTYyjwzBYMqS4QU
K4ho7SpwjuFEk6S+i4b93c+/uM5VRfw0ndyYddXOz6GQqzhtu5h3676lRkGY0IZH
ZtqexhVVdC/Z1wD60h20XmXceUVSjGNc33NN18nUmYJrwmRdJ/8PuilltNmYQYVQ
96e2e7D3c+K04suH0OVRT4LbGn6GGl3Qz97snm1OpUOJya4l6O+P69ENt0uh2X34
IF9kkIKr3p22H6dJqt97x/FgZmA9SMp4E7AXlcwXMW4GHEYuMucFSWwrInqICFQJ
WrfQarohEuoW50ApKg7zOWfm3CkapTn0iGSsnOpQPpsrBxtFpA4f1rNtjHgO3oK0
2q2W2lFh67Wt6ifOuLY2KemnKg0eDpo5F4J/9kpmikTHPkrXLdbMeh6Q22KfCJb/
okqwCCO3gJyAD5N5aFHC0Rx0LVhNYLTYubjjtTHMEUuTGe/vWO2KwxVpnAIxGJxE
a8ydJ8L6oMaALorOzHdGyF3D26pCorsgQw6SxuODazWuCAZ57EW0B19Em2UytQ7w
3Mcqbs1ki4Ij9xgeUi4Wb5FJyk9z6KdwA49Up6R1pYslenxEaGNkxFqE2ZFOOzU2
+KNlqYhm46PPfm4OtvhTv7N6MWN+0RNbraU8w/UvRmrbuOhDkAev91KqG0lpk/n7
bv6qZPC0nMVgQ76Wfvn8t0YIXW3jhbOCMm6sJrgfmifhirkr4hghSmL1+ur87Xv4
Rvl/+AM2Mt2HDTPfHrdzaHDw0+Wnc4y2lskv94gc963B6eW0PDcQPZ3kh7Qh7bTA
Q7PG1qEZytR494AZpHjNU7pATA81j//DNtLNqOFtK0SQzsPz4uz8zmqvEG8zEv33
Xucp0L5NTV/SceXjw2Rn0zYGsVQeWsSG07SL8wsEOqK5CeoZG3XMaADl9CdBQE5g
2gZfiZ10ocaUS3YScGbHfaK1Umy39HvpKoPm5m8brUOOU0yXEF0jX9nr6xqWqQ2Q
k/8edR0Wu8H08aNTN36vDyy5TbRSbtCcmKq415Gy7RvjT6O0Rb1UJjBGBajqocQM
4d0RNUx2wn7MW7ySGlFSDSDUVclyKqgBp574A8y8j3Gr7hR2BVvYJk5lmaO/AAUh
MQzVrDG4ixUq7ZMHLatd3frBNGJ8EepGXKyxJbczaSGOCUspr7rA7WidzZ0trEDs
30KpER/zvnbQ/DXnYF1wX5pAhUFbpdafaxhbEoubOXDCs0YNmLKhRblhz8OeNJzY
j6Me3ZF1dMDaAJ/2IOs290a0TtJm4rE57y3PRH9SxWZxGmmWrsd6Rel9vRV2wz5M
vKc51iLUPVmZfMvi6OfOXkmju7aOuqrQ9SH1w9WxP+g7xxdXluC3bzdaLku6pOHJ
EU0fiBMAVGC8m7iXzff0BoemS3D9LdUAWWHfOXu9QzztftXPtX5iCyQWtapp3+i/
zhyuoPPrOT67Nse7V1mA8SvULMnrdIxymwndu0yPuanFQT44QXcSU4k0OJeeHdjv
JAm0L1lmi8QKvMQ3/x+HaBwjuUL1jplX0aegpA/vZkZCEMJx4mCPlVQrEHtCOW3E
QiMIeMBQzQyPGqNsS73g1P8fuv/igY+0LBkGxnZP4d7nVoNIPuMznvTXyG+46w+A
ulBEfkVQUKRRzVHXc6+pjAZDd4qQzk1IkCUwGILSIGICH3uYScSiDnqAroiXZsbW
/HxMR9LLufAtoadEGITVmpWyxg7dtfPl+nK/SLXIISIvM8lzlsH2IHffrVHYGKT7
841QgtKC2FyjL3C1yg6yN5fEkLBu2V+N//fDUCv0LkpmfLEae0pT6bI7BTptEhbQ
0NbFkmdQPQDW1U0xZRBUDpIwUH+jJvwhQnZJEpUjOBR/FzEwSEVb0Jsjhd4Hqq24
8VkPgShKDUzOUpz6Lr0KoP6VG6qPbxi5HYNDf1G+gy4MU+V1FZjQah7vaTqQ8FBs
+cMM+lHJSHvubxUWOaWTdaRvfDALVTFSHdItc+fqZcBK//q5un72hwIJRgA+W8jq
LTE8MezkQQ5deOD8QD720x+B9VF7no2x0XqOCzjFZh0hM2b9kW1/yWoHCqJQK4/Q
m4ChR2uVTjd1kwwBr4fFaxgFPZ6MalbTE6u5li5rxxRYz7tSA8TzoAdOZcwBX3YP
bOr39XVenzTECTujzEuHq6ypvbGDMrmqy0HRbtf7Fyu3JhsVXBfPRfQhKucbs3b5
sWwDbaAW6d+Xy85ctwIvTwSfEVRb6IxVW8d3Nslw/jmOZcslQ8M4CYIz3MBO0o90
NsC3WlAQdErLGvk6StRV9ZNoYW+CSdgnREA9BxC7BzN5ydafl1xlGh71LGYaNyPg
1IXmDMrSv3oyqMYpZf3mwYEKuFhyulJFqf7TgQ/tlVD351LL++7SFDvfeJ+3/rdu
E7JpTqRsy0RwKaNod/nk9TrpT6UCW7I/2svU7JL635ngt0ijIU8oNAQ5e5jqg/bX
T2d0jsG0RN8JLTzx7TQQAsP8LFLdCgYwA0SWyRQj+XVsrP8TbCE0A3zn+RwjRt29
1dbeGNAZKQPygjhgm5esfG1MMgeZuVRXS1MfC9cnxEcP/l0VD2JbF0btnFprsLwX
WJFARwAGVUL8VCasEViozNCGkoXweNUnG3tQ4tMvh1DWkUpE4OooRPubYXzze99h
NPUYGADthxmARSLl/oe9I3CHP3E17DyciCB+iw44xeeduRyyMku/nAwwBn8UCNeJ
dhxJLsAG44mCxLn6V6mbCleof9ilp7ZvTw2ZMjVgGaVTNEiHxtsDpPkOUqjUxmNe
wgxaYpai/131L1T+rjBP4zSbQWk4JUJ5hIm3nYRxuv0j/JyffoBJc0zp8A+2AQ82
Y/F8GYC2q+7FJh2LPGpYTygnJPv8EkgUUYnew0V91mSedGlK2zGhxivskkDWA9J4
Wq1lxgmmb9MH68m+LzeqO7p3DtO0dgTSK+Cqiaq7I708eUnnvGwkts+KHaBDFvXa
8BRnaWI6M5HSeT9vlLgc1bMg/Ni7xTxGc9d3ZPqnXjW2IlSZg4bhrsO25PV4EbMy
FrOaKMdkufBRJNc0mdkekDtfljGKYdgfLohW7rN+hATYKLi4Xoeln1qqZaUkws8J
K7tGrkhcdM06+6Hloy6dRIZvyf0nPI7aBk3UiYU/X0IiyozIAh0OR2iE6pvqMwFy
xinmAe2uFtoppCTy0y8T0wGHAV2HvGznT/p2nR3cMtmb3iWbxhSb/WTQWM9hzZcB
RUL81Qnq3GBoeHcbyYRcvCcrUNbB8J265RkzL6J/ZFw3P1gpog2biQ2rJ9cGn7TH
hoJ7XgBA6x0bH7/PWw8XMJTa5qD+UpoHpRj4KDNwHB25/D+E7DCpaJnmXrWLlKs8
fOY1DXWKxOosKNHfSQ+0jCroTY2raFfhN4DbukJKyhE8WK8j0zjFgkkOWAXAEXJl
Z/plO6k3SHPLOF8maFhJBYvhFc288Y7cGL4R45JYq23CImtunXxct35sv/IRNC8H
ZxSCbPKk65y61+acQKm6PNJwSNa5lDjOGpXCeVwfS2h9WPUMKmrgxujHNYka7Svb
2sglcjYd8Mq0wENQ/FgfcV3JIn+PaeN/uFKPCXLYrRPsLkvlyLfjNyzVUvGVDWIY
EXYRD0pzReGfzVhU/mmvn8wY6v1281XIGg0TXTcIdESbkK4D8Y4T/Urf+6TtjpXl
4ttH2lKX+uUeZi8Q8GxBWywjIano5qPA2ycXlSgeykbkveLn17d3piFWk7Ciu59c
5Kyz4EgMs2+rFia/rqJukhXo81cGS4U3kADmPm43vBhXdqRUVhoHFnAKf89wSHIW
Hsih1KPXUYoyFgGh3SmdwhkWRPGOxVvP81gvausn8mUtjuaYg7lStYsbn6kXzeIb
1UFGIVRoOeb2RUtQZISa4LkXvSwcvbjCroexk/9LqRrOL7CKnMjPQd3/8kUr+pY0
iuPaG6geJgGXnN3Ttp8YY7zlm87GCkNjqheqzRfLK3zDGEbNd0lJSIx1JdKMyeLI
m1yUMlHSaQHqa2rqaoCDRc2AEBYeDiMRLEFYK34OwSG3IazTpV4zZnunCNkDVSVI
mApSKVTFbO1kvJbX9QplD5uNEH5c7Lk0ie2ZZV8LniyFCwohE8xjMRHdM9sFESEz
omY9Sa+g9wnYFeP1tq3koCriSw0oS6581uGRuutFpXo1Hnu923wsrcqy7c+fpsPd
65/82SIqTj4CBkEx+1nogPdvATc6UVeod3L3nZQ5JF96LErxVyhT9onhmNarlg74
ZjolbH53P3G+M0U24uShU+oOChoy9cht848WDjtbo4E1oc57GrLxjz6QgmSL976c
8bdTVVOuOrSMsa+iT5EDINlwVRdJt4hlss1mmn+oOTA+rFJdBHkzYgJoh9F7Gr2U
KIyzo2Yf6N6wECmmAAeOHMYWLuMbNPp0w1xVfMMrHZNGV+tourpBjfdwqCRAjWLm
jFrM8vJz6Nbr/UasLL5hw31ZcKfUnnPsssII1HyRqzZ1ijGFaektylQP/Mop61qJ
vBzqUUvCwV52ubtNGLIuC4mAz2KSrMyfkmU6jmKDUZiuSJjbtYRxLpBRDCKznncG
FNl9zMVCiFgqVetfqbW0cBWa4GaATaFbKCsbCnJQi5qkJH8mhHAcRj367u4EQrSq
uoHWrwyAGQINJWEkunrP1pcrZF3yo15bdeFYwvsMCs2gimC14I0EGSewZ6/RKpWt
+SGbDabKkGQHewwm7+Uixovnt0uKyZZXvMFfhQDCb+YmJMYleK0cZ7T7iHyFbr+Y
ZypQ83IdhyD9DQCGb828t6WvUHnOtn7s4t/ISqRgSrJ8MCO3d/C/fe2B5siCqPAN
nZepHyJ7Mb+Ed0Q5f4uR08nd4Qqh4Cu/s9md2ckm0ann/yC9a4cTKnesHVZMRdS8
qnHndnJTAQD7CNM5KEg1Zu9ovN8IgUY0sEwWq4k6mowUoiI4ey6lzUDBKUKCfU6g
iZ7L/LKhUa3Jwqx4rpzdz+pK//LblkXXiEAqfe+hu07VHLLLWuCydphYrU/E3EBt
TZ1gIjepVnb2X9XXu379xZrWMmTC8VCA9lxxOvn4fsNZUv6gZMKVCdmKurZY9eUM
xQfLTVvJoBssDk96qEX74f41iMFtds/sXFSI6OMLGFkEN3EIJPeL3tAL+2AjmGl1
M+TgWjtjNxqnaQYQLf7mTRZ8PFQAwOFPef/55li6pbo9wjrbUxZ5XEJt5hbq/ask
O5M2tccVt3vyFeAGqtv00/9gOKE+LGwMZqdKud8lpcoyvU8oRpXQhTOJ8RrkyRCD
9rll3S8tuD89RDjANRUmlFhnZ1AE/HgO32LWwOQsA5e+in0G1QZ54tUc20MC9SX6
r6o3LK+MEqqNVwaqYfuIjMCkgiNGe36/z61PTOdtw5uY9gxaAqPLDbyqp0MVsf94
ziJdDMB6ztSLuhgAnedLLS5cK7xm+p4C8q7MP4nP5DuSXy5sYNKtvupQsMI/xdQ3
dUtx49arPghxpSivpsvpXypZlV+14vJp/y5iBn8UdsPmrSuD76sQou2+T/viK9yP
rq94U5/ejtf1z/g9I9fAKI+va1iJaTq/1g6TxfyJTXTMNiQnBFgSIgcClsK6yWfk
b8E9lmG+KBG1Phwm0EomTos6AJ7Vu1cxsIIfsVGjyj1tgP6cZdreYHpZSnBNtw+a
y3oSmEV00p8vZyptWs2BvwUGZJmUTL975NDtMFvU84c1KASVRvqOyNOFSuKt8UN1
VI4er+/o85ASBGEH4jERAUMooG5mOKmibp7Wa0wu1x8XeGCFzZBBlhSTHgxM3DMr
ssUR4fKRVfCeTjapk59WYT0ebhSyKYNSjkixPDRbUY9+RuNa/rVa+cJJeUay613o
t88LsLaeoi/+TjCGM5boM6R62bFwxhspBviKHdUdSMRbyiykXd0GKsRCRyYTrmI3
wdymo/F39C0HLG+BdYWjfzh25F1KFtI7w2oaw4uVocVc2+7a+yNe17irnz5HYQeN
hUWnpOEnwNGkpwc7zvT0ajrpaNT3P3sfg24Ohrdbjw0Ob5L3JeEXZxGCe3SVAOZn
Eq/rQjsYLh+6tpojl6HavhMuUmPGZ4ncCs4LMvgBGiAftLaqk6Is8Z6G55yz5L3V
U8R5vFGv5t12RsPTd0RnmyKmlOAuvkLOV+eInOX02/6doSs+hlM1eD0aBgJJqGfR
JDelNwTJfRMFJRmPGBax7xKnP+8rkPVOAXGU/KiSP9RiG5L0jGTOgQlF98Nz1zYf
nWBH5cD4XV29LlHisTdUrnJEhp4+xFiJm4594o6KoIbjltTv+8PxD1NiWt+2RdL2
Kffi21RrrC40QXzIoQBAfbcO5IkOfAbP7XYlTVlAi0lXFmT3oWRY2ZGpvA+tZdp7
U+ntUaporEa+/gtmwjKHJYjG9Gc4sdCQfbK884CRWFWFqFExu63Yx1ULBH4tpKMz
YFi/rgF857KBg0aJHsRxkdug2EtqRB4Ib+6qZrLEyV1CDiPMnlsAFDUCmDM7t+pR
+zt0GEv2KobaeoF+gYg3mfYjaXt99qU0+WES8q1+gg+l9daWGZF1zmMZxrGeZWZO
cqhnM02hyGerwrsmOw6875YsKcFNcmO3FceplnZDpOn0BfZbvlocCKRsbneK6ztq
uCbpKraLHdJjPYpIHWwib0GjBrI1lnEj3DvcNG6564uGJSrA99KXbXAMJptN1Blm
aZknsd8EoR2r2Th2vVV1VXThnhMfPqv9yvkmswNSoihhvOSZ2aphJovkSeIb2dOd
mQKguEszx75BQff5bMP93QmN6RL05KO8yGZXvUqNlTC5z8+EGXGocAIv2mc9s5xm
WMHWTzOal5ga4100Yk4Ynd4MFKBoPhkPK5/fYzk7nIeWLWEr4UnUYjsS7ZI8m7PX
nuDAH4yGVTm8dBvdcPCRAtuqIt766eXbRzs08Hbh0hAOewDmDZzrt3QQlG+tNDSA
X/VWCD/aMXMCF/8GG7Qy98J6tA20A1b7VDo9zLMALawtHMO5SJAFoApmq7HMOxY3
RZwRI045eeVtlpeXTabkCusKwRdF6mANdfURarSa2s3ZSoyMb1mbE4mYcs+JVbr6
mU8lQDvFhq3QAVa9u0jKMPLKxmNmBPBGIlY4hnP6WwKNGlL8N2WaDl6BxQaWRAHm
hOMsJFl80d00ql+HPog7aSzkjSLnWkY46M1YDXvuf8aeLyu32VuKcWyZSsmD8IXa
hgkkzohlPBve2pcPoYykx3oHLmZS3IhIe40I1+h59bMH8hnttN/GUOY/MZYTmVL2
LNj01MpQodK5ma0ZYZ4yyPeuEsQtzohKjffEZ+0Fer2P4Ll0mqg2tEcsRPPbM7Sd
cIb3+jIY84LMVA5kkQfyOcwtAAW+Q6NC2J0X0EJb2T6B6N5zNXbHFjSeHZkVi2gw
qPaYB6Gc81Wlx7sp1FbhRT5hSBYwM0lm3UVG0TFwAGVC2svKmGw6H3oK0lzr4+zs
M9ED4oA+KyTWBNIXUrMzQ5rS7TSW6JboEVi07GndBYV50rTKnYQMX+eL82CsFDYh
XeBG1i0rGMEWNnaRshea/CqrbMb43PI8kLwRiOUDlTB5UJyyaIyovJveVetNxdHO
3rv933fzTKB23BHC3hGpy44qxlbsPBALMVYma9sHOu1oRJfnBdTNAdfLah2OkChs
rMdPqkK3lFIq2Nr84vuCFxEiwmnQUi0E5+CR+LdOkYBk5zHsPVYJnyUkeOesBY/P
jpkPM+fDGTJxbf15z9QtnEV4qJdbFYTrGK7sja4RdjC6+N18Z3mnuvSJmN4c/tUZ
P/OJCvb/WWzopvV1mh1/9iShHOkwL1dPW2Ax6rxy8BJfINA+TTEdXcGSC9SCTnD2
8aA+prtQRg5k1Yc/pwAKb+lCO0RJ2RtiBAFJ2rm6p0V6f2203UwjD4AONT0vRk+Y
DRbhFH/noInXyBJ8OWpkhjp26bUGkilYVUaFLhrJlWyYyXDJLY4pYqQDrLNV9l5B
lnWlRpj3oPUnfPUyl6/6J8vVlcRpKizIeA9XRCgXtpjpehnTyZRi1ppNiZ/7BlEv
hsgV/6e053AJ5pca6Z8srIT0rzwcRLCcaJHEzUxWicxkYRZxpplDKu1Wv8NwVdYH
mJr395FCRBtB0rKHRTQ5pzRYjnk3jK8P06/U/XFGQOl5DENVHVixXgYrqMNVqr5q
SPF0ByWsX6RR7GhC8njPvBPO21cSjvTmqUDklNICmGwG/nBeL3jkZBaW32cqsWYO
mCUGL/e3tHZchq/hslo/vzQCh6piTIEtD39h7lfXTN5DeJj0KJSID62FxJXPXH2J
QnVLi6n7DvMw75MSIb8/vxS/F3IyL4HSxEPn/fUZ9BPlYiWhwJ3aUo8o8LMErIsY
ovI+PEV4CI/lh5+yF2M0a9sJ1X6DezVCC+WTMmx6Uln8UZ0PmujnRolkwolYHyWS
/YLYndn3pSV/a/04tG5DtB+XePwSlSwwIuy7tpgtfuEw0e+KBDD6whfK3xaZSV81
zynQlH+vUhjwrWp5UbRWgnYMq0L7s2kXkb1gtcNYPLjz1pzL/GNNmgDjImVPJLcO
HuWvgk6+XMc+baAcNrwME6aSC1amsrixy1xgJ8l6mh5PS58W3IPC2iiE0b31s6oZ
JArKt1neNLNhuZxtas6OB8HcZmrgrFIR58o5gMFB9QjF2r+wMYwACd7eBhYYFvDx
z4FRKztDbnbeneKs2jxAniYMhStAwCkGX2fxcEY/UeWRwkrMSRALqqjg8gik82vW
FhicorgifS5aSQXPO92jirI/ZO95rgq3/+UvKS9kgJnUNpVhxNvKKsZCFs2wSpGq
iDQpM9qxKmGqg458Lt75K9rizrp3AUJilK2j/7KUIQdMgHK3Bd82G18Z7D+qdlm7
S3C4obkZCjtpk/oLX2mzsynfP70TEakIsqVuA0GS1+5ot8h8BeJeL4n2ZoXEuo9e
A1UURTfXLzTMpjcYfa+W306V0VO2tiVm2FLz7yzRd4t8jNJAn3xRt/9PWzWQQcyX
5U+b/uL0vk7B2zo4Xx6MySbo3igMFSm9eC3XoBtHqInr4aGs6zPxtJ4p7ytrCUR5
9xFOVFXJvMVSoWWkt1r5nSyO8wwwbWh/RZ8I/6gmiORiwqqByXzibidpT92a/Tlg
wirXXsoUwJltwJqVPrfX2r0qGDanVK1yuiGs/s9gJfxp205LS5hpZLyyUdxRVkwj
JJ/GIonFqFKPcmS9EOAz7qsL/Fu3C6jH/24RWYhZ9+pp1KQWxh15Rdr4EYRSjzwu
r7s/hK43X7Wj2fT2k3jxsaD9pEIGuWWuzZ7bSdfvNh5LopDmFEZuKnFU8J96cic8
rAsRdxQ3VO9BeaeOru/TY1RrVB3xYtuntmt1T3SgptsgJMywxuD0tRDiLZyXLaCJ
GJzq5h5+k28dxpqj4GN28LJ60cQkWf2j2J7ba0OJ0npNOUkyEMnMfUXNe1gudo9S
QslQmTAGsNvV6E25MCXxscLb7XfGgMqTYzj+cxkVA1puV/qmglUFQk4Cb0cSN59f
c1zKk2QBAU50msFSdCUMUMp1zJKZUKK4s5h1YOfyOz4vz9OYsn7ct1XiAx56p+4b
dAAPHilOl5ou4xhDw0i0ofsui0mwHJPGYHO5Gd9IDeRbTwnpez6gZzEOcbn+Magv
0AibF/SLG1lT4QDp6hUPgdmaBhQlK4I/Lafo4tnrzktnffOomUPp8zbGUQOyF3Nz
bItqnQFY1vcC2Oq5DI3WZ2JUFuhfYWluc67KFUqjCk9eKjYdh5+NIclMdam5+XJQ
SeQqzfl15SVn2ZTAPwvB+tshq7OtUMdt4Nysc2oZkpzc5g9rJTVyfuLxdkCXdk+M
5Up8eIGaP78A8i1fl+2sKsjio8MxDsNU5WP0wHizFu7hUdouYvHgP1Fl+yG1/6YC
He9ka/iXyq/QH+sRcwgDygiOCSzD8liPEzrbCrj+trADHez4dVIXszy7DknpyekS
Z95Qf6yTqCg6kz1051ArsB0Bia08Z7IlmvGXdfAo1tltrlX++44zfm4cV+EHfsj1
CKzqT4OtE+pmlmmPVLSBt620UGyof2peGtJ4KJcbzIfwJPcstxwxMG4Nb3ZVAayc
dykVS039tPNfnzZEOsskbKNci3OYoFqyqvGvUUZm9K71HPtA4N5VWOITCcKbNINU
7PC6zawqHXoEpVTspXb1Bwoe5RhjKKb28qNwN5wTPIkJ/YRE0giHYx80IyR7V7e6
Iy4vbq0Hj/nky7ts1ItmFLyc0y23XASmKEGhxJOj6bOaiC6ezvaA/i+tqgo7wkNb
t6zwjPM1kFykPbsOmHU+rF5CxZvVzO/nglifREE8xwgSbaIHZdoY/mf4hjYzuRUy
ULlwGF3f82bne0Km3x7aFcwqcdO3iCmxpdxt9u2lTBBDvYt8T6SPR0jk/8c1JqXV
U5+vJ3QhrGTGRzk/XefnQY8xlEoeSCXjffFaVvyphgxBoanrZmsr7qhoh7tIYalw
xY5t1jJb3YulH2qzaKqdKKOP3OeQ8lxRaAjrZosP+ZG+ONjnY2mIFk+d+QGZ8nYn
4nc7KRmAXyjNsWi9ceCr7bjZi3+o/58EOb8fk+6aEZufhT6xByt209UXR+Wqfxv/
LfVhfN8q8aIUZwFa+eQQHtQuN/8mac8peQSPWjhgYIJf7F3ixHgfdizz7UeZp/Pp
D89auvbFgDiyLhnolEl7HjsYX3zyaHsbGKFt4DPUdG25qtUEZHfJZ10oxBA++EkA
D6CRF1LbxLxKSvQveTVu+nqvEseY+h4vW9ByPtggMseWLCIP+cUf9Iz3MOolac4y
9DUONj3CBR7EEIkxM67gwISYGlnmYb1TYdQtQ7kG7lSX03JawRcciYE+7AfBB+1i
0G8qMdt/zrera9VfCnD66scQ4eSN6sUfOODFhpqhSMeZqfGrALbQiq26Fff5SDVQ
p6N8wTCzokYIliWrLXdxfkdNdieKFQagSb3JjmE175XuqZROwq1bJ7XiSyOs5teI
7mzWwT2u6hSjPhrd6dlXTZKFErWAWj3l6gbLENPvBdtJKpUZzmb1i+wcQFeiBG66
bxi2yK3JdSXChKvplz+ADKkE+MvCNxLg7LO8SYDxjc0RUd4aVS6wLVCZpPA+k5fN
y7lh7p7WrG6HxbVzOwrifKCr/rnZWsrkxBPA93cHsRYNXt0STHKZ0Qr2l/L7WFYp
AK5y8ee2qQHpHeYYthSd6Ydh9UscYgkUBQP3qbj8/D7jUsXkIKY2HG4jardVdKhk
yaTyVADgT8eZLpXz8UNkwoVatkK1ncPdVni5Z4xs71klRSd6g79ThnD1ohuApAgW
SXZmmMw2p5DRxm6iMhGQjMHXh5k30DWZ8YppfrbLtAtCeqqpkWbGyC5CprRoInlg
gOqD4aUQEY6/60gwJ/TfLaC0XOam2xciOn+oc0Yi2nCjnDmAmgmBP1ru00ws45ed
Z0dwC9LDV5h1cQ/FwbiZgk4X7XqXJpPHJATLiHdxpmgbaxlyEacEma/eTaNX2NJx
Zc8BOlCXfDgGCN7AUVLXt1AIQHLJecP6/j+Fw6mDH90GPCWojfEbYeJ9e7uP5/Qn
e5URPdbIJ6BwFczygn6jrXQswi/Q290Yps1x79W/ny/kwBBi1BGkm1BeZuzYn1VD
x3f+ksrHm5eYWS0XyGLVs2+xY1bp6CsF5diK2tE+VgAu+ToytXCjtXP9voDZYGhT
gmYHMcKqRlUKEONbiqqopqdap/gCgfk66e1VXEWvdnU0g9FWmmqv7/V7yILH2Ye8
U5vlipJD54l/3Cib5KQoCyd9FoTKTuPiVK8mCjmVAd5Q4RiFNu/dX3Ktsa3LBlBc
rkNVQ0iyFhuBWSI5N+I7iaJcUEh60oUvhSAXWyRih9XVQ9vBFbIJEIZSEw0cI+SL
9XXc4N8Zt76lNPI5RnQ4HFN4F4ctM2ZhXd044AxnpJpPhzLPMFEf2XbwexkixJG1
OGmOyzfRkiKgBVIKewiwEQdj/eXt3Ee+m/QNkOknX9DdfeJZWYGDZychM/2crovi
5C01WXrY55GXrJgBgTRZbWWaFTf6Bn4rdJnJ6pTnNoERl+CHr40iqoOy0qZgP8X1
3jjFpA1d/8Zz1JMAG72waCoXqw9psMw/AAT/9qOdg9+4RmDA5ngwBlOkghTbMH0/
1lmugt9HBq56o5IP+W1TndmsK/wc5A8gGRoGKo3iQzuUJR+4JuHw3NCgKB45NB2U
oTm/Rk2YDyehJDOaCIMGG2cgUN3Ec0USSb/MGZdmqJXeQh6toYizqn81dwiu37hL
5zb/nAanjXLzpxqhKz+B6tIKlCtaFd+SAaXn1aCRpXt+5zCs1VRdxFM/rgJR9QMY
7tm9ZV1a7pbSd0Ad6F+RerTb5MBvyQfAtI3c47RHUrkg/5+EiA55BZ+C3Lx6vQlh
cRnXmIc8C/1KwKNFmMPM//6B0xK0H1M4DxtCFC/429uoBPQPo6f8EodqrHv6Ztv4
0FMd/Du02jsi0+nW2g9mOmzqvkJcA5pnXK/O9rI3Xgb2SsLB0XgDIQQj3kl6yd2Z
S8OElgiRj8rMZiNglyEJz7U4KTmYfyo2wbMRQ+eVb+Em7IqseDEoxaB/iVdVwLA4
DdTWfS8SF3dNS9WxlWTpja2uDWRsPn+2fsIw9JJtUHhV89n+Xd8Z4krc85tOLXq/
9ESnJyx4SEd71WSZJoF6rG4r534S2vIhkW34xn4sVFUnQjV17ZP2yFQCbxv71jiv
QJ20rZ7NRViDH9xrInQV06Y88nFnuQbMj1K27h+4cU2PgSPsPwiQqEKSdLV2dqFV
OciW2KaHrC0T56SqxmbcvalpV5Ffvuafo7ev2VZg7NUT00nJSrMi63C3LrU0j3Re
6bf5yUu91QoczShm4yEMWxdBwObP/mEm+l84qxflJq7mHo+IcU/FGnMNwmTkUT+h
YllFjHV2RiSG+VRvStqqbJKM7ngmrY1DTh2dGP7g8sade2wGzB7Sad4kciJdip/Q
K9Msmv0o+AFj1bHHFsNyJRgbfmy7DDOXpsqGwTBvSX5jq1RiyTmmn2QZTfAw69oU
Dv4eFwxeeoRQYiX2Aa5/vGzysXXMUnm3XCpibwdmBh3lOykiVDSb02uAaZvoc2ku
/FhDI5NbN4J1Ln+escy/uy41wOQVrG50mcFv3743lZ6JDVfcJiUuk0JtrahZht3f
efzlao0npjupZPigcH/+K9LEYRh9nRiCxx/tgj7XSgMOJcimVFmS75AL+GP0EK+v
G96XBRUYAaMb16Mm9wht5SfKzCPdFFG9ySB9wDbmug50rmDGFVZPj8aAndk+RGUj
vCU3UiOs54E+V6S+iIwZqL4eXnM8fgd8ywEH6irG/Ti84CvtOqU6oP3ohouB5wWR
oTotMSriAYv1EfKgH3ZBuhtfog2qetYxjkFNecpRnuF5zEXvNFQXuDLd+QT9pCTo
s6Pc2yunqvSyn3SmYQzVCzzShwpo49Q0q9IauFSp4Nb0GC1vvlUuA2HDd5H9AHY8
mVfLrQ5yOfGc8FeFtmKl/NOqIGb1F3SRSrQ+YMyIh4xItt/4b9tpJLPxxDbv65WS
wW/jM0HZVvzmxwBNrZ2F5o+PPOIdsfVjslgq6W7Psbwi6p2o3umeGc4EsbQOiNB0
6YsiGA31PXjJZz5l8vtvJ8w+OSQKE1h6vtsdNiPm7O6nf7KHUW6q+geg86lG8HBO
k+WLiM66/zjCCHtGBKeNeADlajpXZ+eDVi4HOVS6U2oUC3hzZsPOXLdKPLluLFvf
a6RgujXZjILGbZhd7ztqOyu7oFPsNvAYs6+p7ugq7MuPurB5iLI3/9acEcSsMnM5
aLtGbPjzHk3wQdAJe3RRaa/XJ0SQjwqObTaAAszl0fWr3fsA/tmO6jKi0AD1He/c
yQ/BI5vkz4TdziYrszPicpiTC/GrqB01RP7Eo7axqbQpvUzvi4wivogtUJ2O4S9L
H7a7unUdlBpA3de85Y6ChO8wTxaFirfX7YbiqmVkhgdM3T82JLfkbFgn4D7RotGJ
pkUYDrgy/U3v8cMgeNlfUXJIEsnqEOBU4WL4CZl0kCZ8S3aYedO6zI5/oJ5QzHmn
BDZXsvkhgmuwyBbqawcmej7rfG146LWon2Nfk6B8w/nMLNZCYcZWbqyFnrK011EK
Ccv8JBfKOAxk/r0EU5K4LD+PaoDIWLaZlw2Yq6jQbY2GCcHEsKLYR7K88eqrJgKr
bgzJHcnO9IdxzeTfgjSPvFtcFlU+KAQCkN1xTWwYolxHyxIE7wpjk1Yov//cub3z
BqhCQ+V6w/GQMTxdYJPlyITrilXEG9MTOXwY1g4vMRhBnIt1Mh6jYbT+eyISCFNP
2s4bmJCBIw/h7Wwwmv3vJxR4J/pAesC8EfxfF054RqMlN6fStz72LL7iJPiyF3Gj
tBgfLcdJk1zby4gbneluLqNyKeYgxEQCGuF12OOoWASw7A7fYJD9GFW1t5+pF3BU
GvO/VJdx8Jjt9gc+g2su7Q40FOKSEb0tUzrzo5vK4AUL581qLoJryGhzvJtcv5U9
5OhyMMDmg9Lfvz0A8756AoXQZsfo2VyNSjgaCTbaPTno7IckzfWfzFCTSksP5QUL
Ym7lNaDupXRgNFjY/6dv5h6gIXjISujLn4t8JaxrogWHCEGgco5J1B4B3wvMc3LB
T1qOph6MyPAEch/IjN8CvsqFA2AVFTubomdxvHzS4HhVxHMDT9R144sUOgCpD3rs
TThOFjmMliwI0t37uiig+KWTN+SD2qpP42qiZWqfBfzZKQ+AgZEdwCttQkzOuz3s
P3vTxk/ca6gm/IUKYJgIm9ZTwERpj9N3tp78ppZC59LDzJ0JyG5NcMPEgufQea/I
2NaijayvFAoNYdV0VAx9UMkRQ5D5vDj3lFTWnCusLoDfe+FhHrGt9UTJsW5wj1YG
yJIF7aKuJ9sY1tlOGVInIMXgSdgHbPgY8UcDlpMl/On8W+M0rAhmdRvIM+CvGCzh
0MQlfjqAdFt8lluZInLVa9ZVwvx9XUFy0Gzf6O6ZDPsSr0CH+StayeGxQrl71DnF
OZYwfh11zadbFoNqZnGGNOgAZUm+99N6ZjknnJUGEBDiyHhxK5rDZt0b7IV3NiXw
Ddzo/Ajif/pzIo8/ONa37zcoW/R0bJY/Xjm1Cdu4U6GjEupl11Ahu9PHZ0SHXrRW
C8vRbNA84mjqo+8ekwdD7ftG2RVAY6KK2DrB1XzNA/DdmI3zpyPEwGb7cQ18sxws
ZIoxWE9X7Lup9A536naFDp7scNHhwnxfo160h34hi5egLQDn+NL06Mz0dgoF7kVF
GG8pwqltXkGbMmf6eIAP2wbObhOjx2+2ux22IqlVfkClHZSq1OBumo0qmt5haZOc
ZSs/IZ+RVM4GpkhpfVhHQYmwmVzr0/gj0vKUjD9dtJ8hYN6UNEVOlUFs+mr/2Fux
UP8HyoWhrtP9Tv8XmKHMsp/XOkP5vJFK0Yx79YmAaXRfB1v5Tfb+dS6DnWhhbM0V
n7yzLT+CpGstK/mx5e+uaENKq8htJlWEquZ9xyP6y1Dzzg+NrzkEDRvYjVd7+TGG
SPrUQRLdbNcRanEYhqCb+uoGVBBOtnExc4uTbxlZnkUrFJKBlqZAEo5UnyJakgdq
5X287mV/0ZwoeHP4cpZ+uKiyEdkE2FF2nfs95DoCVX1wG2CXdpru1fkCnTH4PPYt
GSeJw5c2xtTqRfZtbr3PgD88K02ErFCfQvCRE6fDe3dhq9mlYfNIOERgiioFY/x8
TOjyhjFCSMlLHbSl1D2mNI90GtIvAw4joGp+WBEag9nm7roOZ3qYEUm9ASRyeYZV
B4z2bJHxMqMsoWnXi/WY0FA1lLzXBDeqtBGj0JJodnRm2/jsxfR92a9Vn9rMXp0V
SQ7pqebIilpW8XUCuD87ugCesy9+mziTxGprRITtO/tBiTjfoGESb1lFny7HmenW
/oYrPFSMvuga/LGTfB1siIWDLoFa5ORtgQFDGetV0MGgd2+JPG4qMQKYUFUXG9FB
BczhfiEHPPKojHzHof7rPjpKdfKMheibsNKAYW/eUEaemz5bdCU1Q8v9CeEC8S1l
+LVh8g4Cdt5lAH3Ixw0OdgGl0de/4mH+DdEiXoNFbu20obFYEsYSC39nsE3L3eSU
PCvFQiV/YLYemcJp183Kg2KaZcKT0F27sUIjm0603fWN2Yo5z6GspKsDuWQ01vjA
DnG+SOhNpQqLybFI/zFcsGmS8/szZW0EZtGdvtWkYWsL1me3Z3lX8Yc0PialpX7q
iH2H32qsGp7LE40d1l8b8Z1R/QZs98YY0fcOjRWLV1SfnViR79qyMpA+d9Sq4s/T
+ICKa+1QpzjOhN1+oF4F4jqCj92Qs2Vg40iPODOXdmlhWjcSZn+R69DOaIi7Z69C
zlYWjlnl5qLq7M96kFcPgtuSUIT1zbj2vyeN45gvg7wgOBVVW9u7ScmCjujDQQcN
ikU+vbr51p/PHsRKQccAvoxFgSFqT7IqRKzLekTzvRPlhsfIF/6v3vmt+9b2z6Xz
w9fGNozSaQ8N17m6uGNItHlzMv2nSZGo/wPPZX1Z7+ipRlkGoxFw32v1mZtxZff3
ypY30heXyV5Ns5yRTgDG6i/ucHXnYH49cIGGOgbVp2MLMmX57V/374z8KC3OL3Iy
b4yyhmAOG/pxbarRWkBTKDfac2Qj1d+Ob04+uU8yW1N31p53lI2QXAB8KrAtKNke
gy1UcqRzxL16A5VICBOaiDDnjtEou/bfn8tyJSwlzGGfbykh4OKJNeMycsLmxtjN
5ZDPvN/AsaaIocGwU9nzTB2z2gGeQGH8rrVer5lhsCkzaGP8y5Rym9zyMY9JYxXb
H+T8/38Ai2MJOyb925dsHX9Bc0MkptOje+WZFwcI62Q6gSx5/gfU5IogD9BaE20V
saWu8GAcMwkWOeROfPNqdyITYQp6RroP2+Bjsw5vOLLmSlUKtUba3th5eKiEOLJH
gSf3llAx8JASoA095JMDdqwM6OE4iWGaZFltH1kcPeAj8tntoLncxfE1mPo7LjRq
Yc6H+1fxlr3MHWygvc5O/lGIHRQJX8CpTdFv1URVxO0Y1R8r9BPesVR72DG/uKrP
aKiugs14uLPzYUwDFB/+k5820g2N/yx+MP0tGvJ5GM5/KaSaWN8vG904MGGa2x4f
dQSJGHp51/xZQVHeQh4Wzk+t2dCBuMwJVfs85ROjBun9q6ZWgXC45qsL/fwLHdt/
HhJc/TMkIGZwezTIYOhdyLW3cP8qXQ+RuCXpRdfeY/sHbYSiknV714tQoifSOn4k
nuQg2VX/JCqMY4sRIjMpFq3sRxuLk8zaOYa+wmG52PSE8edMLzGYtN8OO+Y3AFkP
qyfPcfrLZluT7MoMFFvJtFP/5Vu6ih9kzUtQ3B8Bilswt0Oiq/mvLS5Xv2jJg6Hh
hqbQLIm9W0Az9J4wdyhPgmr00Y4yvGANotnltoLmKBm9KZEgst8dc7pH5Vk+knXJ
d1lMG3GBxYAEV3s6DQiK0asoemvzOetZQjWsmsnwXpuIiFh3RykJKla/DpuiMw7w
m9k8kgxHmv6B7ALWK0DbuCecLuFW/8b5QKPt18O22g/bAA6QM4IFc9CWCKSPFjCm
GIp380e30XLVkX6cbiyETMaoq2sAoVkrpXX5KhQiPrw0DylPErG7tDD8fdIpvr+b
cRSTSr+64E9Jck7tDO9Jc1LyU/F4/unofQrLeJe9kLvf69a5Fc5RjmxakUC9hDCZ
/sEVPQvfLrMLsZM7t0Xd87QlkMlORW7xdlizvzS0stUQUUqSjRTGevxnTLVSvDMa
pn5zKYOYKTd40kjp3HZScyL1m0lPEUCuLbICiIiupD6kfabLm54hSnIdVyw296ux
qcW7+x+69jgSiJmCD8PzEvHJ57e+s7rFstV4jXq6R/NGCIWyXkR2Nif558ox/lBD
ENEDkOEZpzbb0lyp4iLvY2fEDQRpm/yzl6xILHvC9iccT3qoGR1ocYAI5W+Auf2B
GD1Pg/lUlD5tPWHfbTK5El/rVTEfR2DvO89eFuK11lUWDlN9U9PW1vxGnoh57qix
mmpyG1ic56YF14zo8idQRJi6xiE1Ok4ltOIcGb80nCNVM/RG10MmSxuK1Isiw4gS
CDQajhgHULNe9xYrBP9HWInfCayzzQFL4T+62guNVSY+pk16Dapt/jNBOuYf+SZZ
rJi5+AEp/J6ZMurxKCs82PVFM3ll79u61NFI02SVS1TcflY5WgFchikNl6RMJmTE
Vfh4/haOPvcUtKNjP2OCCq4Ux1vmrjHJyqbaK08Antpx55Qpp6UzFIdKtJpre1t3
pEo5hQURnACARIzDlRH+N7nK36CdmOkr7K0YPEatWF2uXqVRS6GCI0oL64bfEQnQ
DLSXMyQwtdnUU8RTnikeS1LJw9mGpF1qO6KUx2hE2vdR34ODm+J0OyTt/d4r5kk8
I7AOs8OQoWBzLLX0Jk61pfPsW6JPMgAfmRT67t/g0oWke2aLyClykWNtrtyX8ppq
Fv7b1y3Rp0UgehOP8aBGjOGiINrygFjRazxFh4//ghhwoClQbzPArMlMwJJ63bhk
wUPfQ6ubxzFOUImMQBDPTfaOYE3/sxlcZY/zhmsuOWuwalBfA3iLUz4K2i/U5gGU
Nsu+D/ApsHEStq/Z1dxJDyALxTkaF33haPkUoFRPRBk4VPHFrbFN75YdeyoP4aIO
xA7bLHDpRdupygzH5vsf50tSrsfDkilnLUrO7n80kk1qtAj0RshCP2awGPnHHb2h
rHCRJZ5hJvdEHM0HpDYHiKdh3GqY5y8yqUziQnFHut9a2EBC1lBT+am3kMWkps5P
+2topRmRsO+/AUVLX05/0Ox+c/nXXCL7C3lKtK9FuL4IjHVHx/Fe3PpDget5pk0k
+xQxz9t7kLd4Uzn+5M7HjCsGh5qu2xLPiXhw5ZCGk1fhtAINtasH8BSPShifSZ8a
Z11L1VNltS3Qfkodvt+8F9Pp96odzdmoxc/2aY6G88OuO1rujav/AXlCytH7SEQh
8axSKRo13co3wgVcBIFzSzQ02/UuVebDP3H2nZ0zfO7gm1a5F/R3tyyqrAR3Ib+J
68u0i+1qzamHNYsf4oz6thMhhP2e5CzYUnn8A3AJ5PMri7VNKEcIA5F46HTaZkTd
MnGEtZFgx3QvQCNHxLiWf60KJ4lExSwnjBW0I/Vq1p6Go1cpP9r6c7eSrxVK+WdV
C7BrqbXFjrGUNvMpP/re1yN8IYiAnzqmZv2AxnoqEBaxeqvKlybPgrKCOBwulC0W
cuUvQdPugKHjzjrYj1QPqyQXtfz8QTvtScRDrvOY3wUcaFkRi/JdgNHCHk02HR38
HB/tE6AELOb5zlhLEN9vxNyWvxhlJN8MhsnlTI2e1aac24/xohx++W4ZvImVFVFS
arq7ekCWT7J0LUHCR7YPyu+13Gwg+9uJ/IunNjjhbAacdQLVEBWFk8aAZAw7bKKZ
rfG67o5arpspNYVz6AEN9c4sH9Stam3yvgcWMk0ETKVFd4TN3/BXP6NjHW5on/mv
P6rBHXg1+ONgpcGPPERTShv0Igs9Sa8VDnrv9uNQF5umP3cq5wJl6OeWVAo3uCE3
Hj5VexCuni0cHIcPaEvEA3Epd/p1hx332/pCdF5L6dW9i/Qlx0Y14vcRUUdDjS22
6mLED3lWICrjLixSTpGNrU953LXoBOZP7yHCSol/gLRtYaP4pxgFkt0Hg5U1iP6U
cFsJHJZ4ClFMkTb97HFcmqG/5v7cG5wi2ayqbyuvX/axxEYb7SZYU7wp6lkj1HSW
Xb1d5yzY5oghFfOP3XZp3D86L4tiwrRFAl4HNZvdaVnwA2uhcKxi5UszCQK3+WrL
erFBlMHPE5F3SjYbFmbYTic7pWhn0k2OjGd0v9YhengRm8xE8eqmeNsk5kEZ8djI
tTgTQSfCS7chjrHBX4Rgm9DL+jSOL2L76fSuLQuOXUkLP5tzaSgiD83O16Pw8cL0
WKYn9CY6u0MlJnbdHCqys5GX/wVrU3uCelS2C+txQVybcKA7ucXGMcrEFxetImIK
Z/YIq2Ibr8rXpK5wJhKw4StmhVN4iXZPjtnJnoloMF07t+LelLfYmCcYe1SlYJDF
lkiAwSyZ0cBWz85apDhIZ8s0b0BStNvRO6HY/N/4TH9+lT9lgjjRgEj4SFZtXP3K
rfmdqY0QLTqe0Vw3BXy4wsgy+MJTJsgPb/jnisCZCEWwjeocSIoYmqPE6YwW6tC5
KIRAG2Ly3TkPu33mdFJSHVxGeIqv/Gx8SQ9oNwwIPeHSo9xI8R25updsxtBkOWJV
SQ3SL9H0BOhJcyuGe+FLsnaEeNCHqjqGcZ24GczwrnlXDCX3Q7ev9IqWJh4hphqI
JzxR3d8ULaUrsarL8OWTg9pEInZmItzL1mg8mJ1vuncw5gfRkq/XYKnQt8SkR/cO
O/tk8Pq0Uib8iNkmVSVL2u0jjo7KAEgzHdvPdwm918B8i6NUy/X2nn8ZttkhH/Ei
WQlKarhLR1MxzvBl4XM4tWF6TltYswTe5V1bDS6ehRibT7tb/he/LA0+PShamuZW
QqzmVXxS20mxS9YNZKOINFM/48+/E6Jn2Ai+aXgIyP+0xTurkzXZVEDEGWJyzGWj
2E4pyNTeOEHk1OY9qjT8fCXh8jKiTluj3rd6Dm8qkdHzgKbnaBbtHBE5VMAiwVb8
CcsqsE/w+c1gHEwz7BirLV2WhgZLRPSa1tM/iT4hsSHwQt8SIZZXJC30uSnon45b
fVNIzv9FsWqSaPa/nOtYH3vazvX+BeyP885ETtxlPbg5VEJoG1SJiklBzoMYDovs
mTld/N1D1dEwukjVW5FQGrImc6FGmkFVVMKimW84Er/pNobf6ctqvaAnV0/lTG5n
7t+r77y5QT/sRIYeBTlKNBQIBaGI5olu+Ar9l0WZK9KppVMxcOz38/nSucgOZb3g
eg4kYLQMwbOAVPIno/oFYa2rwE1JT1p3QUtRQe8+zVnZ76YduTDmY+eBQkWjZPqr
l12Zw1Dz251CaVBUkj2luWgm+3GJSJvwsXUJtA76jxOspouNub6Q3RLNOpOs7S78
W+nXzBqfJjjv4Hage97hssGh4Eeh52tZtUzrftNrfLI6N4WAFnX8QASTzqoyBTMd
OecntmNkPSuxxEDKATvt5xmBxZDpamK0UDD+SWr0QmWaNlVq/5TwcPRyFSWiypxa
XHh2XDZyt0KST0CMcaRXbLZhrJ4aE2OzbDb+Kpnli3OcQS2n1ae5xjNNJiZufKyk
iRovVKUZNtzTvXUkhbeQoLNTZ0j4UI6eS5bBdKsiOCW3k1tITvlmT9YiQeXgjEK6
GOQWu5tYQrkyA9Za4nVmtTlA/P4gMhCHcyJM2VUjkW0+mM9BhDaKZfn092eNzCHl
Knc4JsWjlk/Yy3VdOpfu5V7fyjjN8gn3V25PjqrAqmUgqEezRsoGwTYdth6DEmWB
i3N6jOnexyaxAz2mJiYXoyO0WRfQBl6NqYdW8DN+NcUWcjL573XexoDiE+hmkEB+
+acGEhj2oz0AOnZTH7NtigmUTL/2HO+rVpnicIAJZDIAACrp0GKUet9jDHpi/H0M
Tgn96/y/4KAOjlz1zbc/7JFmtxh25Po+C1O9tbTx+j23Y7hfyxYsRUckA7QgmLQd
FOWXLmksN3QmSBj+S/ry92WVV06XHKNB7jmc8ckqCp8AO6La72Gbkdn2mpAGvbEl
wGkpN3Emm+dBxvhqG8Ps66aWfXRnm/EQK+z23KkzYjBF1kUKgVvld9hqWPbI4qUG
yX7aaPvWsovK3jH+EVF1yorbLXPH9oyE7f+E46fWBrZQ2jhzCLq5RNZMnkJMAHi0
wuNXBU1CHKxhlxyXsys9E7g4kosWsWcex8/1PryE2Ar39P1Kx+ls0ble+VCN0nHg
EVPENmLdqv/i26xdpLI8Jky1+xhwXL+ZKWDjA3XrPTTCG9lLQFGAJoe6G40I+QPB
Bii1HxMeCNQV41MYcYcJMax67nJ5Dt5zBuGLFfJpzUkxYa5HX6P1BF4kHjG63NYW
T5DpzNAaxyPnpGN8NYx7B8ksII1wedjrHFNZoBy50OzUZNkT1XJ2ua3UEgw7pdOB
RMdppXrWCmr0EzMCHbb6yHNd3iRdGgKc7gMQyl4P6XNUl76IRIF3RNzYFNxhEO6h
7iamh5T79RgwZaKbVVfWANCrX3Jv6gFDGjDNbUe0P2kO5/BosM07uOfNOVqsfYtM
qmcmWpoqRDqvNXhtSQo0598W/doLQqwv+bLERbkKeDXmoj8G3/Q1T3oCNQRbUMd7
Esk8cwmqJOFsw1nNw/gZ9M7zZi5EuW/xZCYS5iJaeBS3EWqd5brewnf4Ue+vDK53
rmz84dRgWHED8q2SsBhlGLCcrci8BqR1Ip9iT4YpNvnLqJWPCt8nZc12hYWBqLfJ
udl8QG4e6EAciZ1Oj09cXVKl/FhlwkobEVFO45GDlVKwXbJEUH4KoRcZi7V//1OK
aV34L2lHiMe5mUX7f5YD88AegQ9jDqOe11RjmJPfKhYxygtUHuzWGfjzXNJyrUuh
vu1wgzsk6O0oV+/azfquQ+e6ReS7vN0rM1f64QQYeWJejsRHBiwJVvKimveBNu9H
O6JWDWzla69ZXWibE8P1WdLnwj86gEFe8AtkRXT7QByDT09eESpGu9go+zFaDEXR
PH4iT7Uj/RGrPyk3atZUz5l8lsOyxWpsNbXE7laGepoLbCeqP5LR5vRldkh39Yhm
UOB22bwp4HHR2O0pPPyNBkgnMj97r2gUMzSfrqt3DmBJof45U0Hk2/rZeJMSj9sQ
HkqMu3tWDqh3C6+MWB8mkbkJKAyyCNEH6VZsW1RTDqzuIZ7sY3/FeBVAv0XMZwdQ
ujLpZsmM0HittLF/E1R0rMKCwtIIaATEWtziEqwMpUoN/2gu9OPz4DKbJdRoHwRz
e/4pbvOYpI8iqy2MYTyRMlSFTQ3Fi4mR0o+kRKjq684NwhlXqlXtalYqsvRhOyo/
nPUGxngalvvZrdigm1tTet3aTjw74G3fY3dQ23/ULkCLocqbc98+Vj1V3BnS64yc
ic7lOT6Jjk6iMU7SfPW14XuQME+rmZKX7H35/KXJYfC+hh225o30V+gvlkFI6SYP
AW4R4YOpzoK+orSjQh4/38Rz9xG0uH0rxBC39Rm3IakjYY+cDge2INsU7+/pQ4sK
PlxPLneinGmRBXlhc51lTTCcgoDWWHT7/jtX6MAzhZCZML0BVwY1RFqJv/WeVcS/
qqfmQU/7Tdkl7BSARj+FFO2j2zWIlJfu2w+Ezl2rx7GoaB1/P32wAN1126EdxF+Z
+vmE44gHIqQy03cLcRhhiow0gfQvorHysHnntiYBKI1VtYgOqqIs/5REN0xG26Qs
LZUIxbb4sryUh0fbrjRXa5PGl29OC8KGgeE9jBiSqVn2csUDBvxpWRU8h2EAqVgA
13p7XgjUiNok5s2KpGrfDRU0HeF2RFnijpsxPerw0ckuQDumXzPbo06PzUvir4N0
lVrC6nh8M/U735u2JQTURAlf0I1YzdE6+5w3V4zOzMt3CBCEONVbIqV84uHbdyzB
5mt+emVIX3JT6gu1N3FQV3UvVtPZM3WSANLCKAUafjsDVqR22xZ1ZiOBM7p9eUIs
8fjnQ2/JudBAdicYN5HzgVtycXBRwlUjqq91s4l/cO2ZxQ6+QeCWfyUceBH9UeTg
I1Tq4WU5JQQomUUH5DaVW4MbrMYZJYKu93iuQNLJ+mOPVwzs+GDTukdkOC4p0kkk
aFYwDVVqMyeLOPPDk1SXiyeIQc2iDgDAFN21+1d7OZS1IJv8u9UomMWLR6Euptlt
U++IdrMZrGT78JcuXd7AEzJcm2RNqYMTZ+y8/Gvgl13h7sV+HdykH/p17h2osxG4
keJuMfhES2jC0zD66hG3jhTeXELWMDM1ut/452mmUiY6i9J4/e8teFhHKXVdmifq
h4nR1UN/+6AcP8rxgezMGq4++yRuY2p2BUVDn7fzTPgBTDPWAPBsNJ8F7Qhaofv0
NaZ6ahSTXZSHvRDawcWGsOrN6ALHdmd6SexqOpeVjubipevxHaXDY40lwpTgxWRG
5qT+gv1Whx+eToHoQJnP2hU5xJMKllKV+ucZYZVcyAhHPGc3Er42CD3YKtm7NRph
5c5PRuFZaT52Jsg7VU8DKsvIneFO6BVY5U1iP0CV0aRNupL6fYFo3zde9vhFrvkI
Pxs9QZgZDaRjtLo83ZFzP8lDd8ojyxTDCnnMr0o4vG3dFliDWqcT7SO56br4QktB
6wPIUH1IQpYiYVVEsXTW28BwAQWqgJijAEE6q36zXtvvs5xyKA1J/9dvsTK7eFGW
Vps//JKMO1WQjkMlO4rI2JXWUJSDW5nn4+DhJQn2gts1Z5IanVZipFhjLfEUez+G
WFfRCZo2A52qUbPyyk/SSjcSlNx7DiFz7JXXL/tjuIgDi3qQ4v0D6ZGPaRdC+JIe
Pe9geVpLVep+T3URDt09Naw1vH9m8RD9ZzkM1aqdb/AUIJUx8c+ahd9SHUjmT4/a
Upr6FMfvmKLcycf4mg1V6irPEqSlL3BbqhJqe+/RP0vnO3VAG0oYl794I/OGNZr5
LLsYpqAWsLMzMDyWqYGGK805FK1jZZmsfxv9TVwer1G4KRfRwjRPtRNCIjTmcM5p
bh/YSSgIa34ZkDXBGBNooIGGHsvNTh2DWnMAIPwV1PRgwkoTh6/SPKyzA3ymEIhW
n9BHBvt267yLXjMoUE+jBBcdESAQu/joqxyGlWzuZSj58yjGcqV+VsXvNB2eCwcY
gu5QLkk0Nf/yhXqjFbosdTjwPGJ4YzNPqtiZnSfbeqeIfd5XXQXDDfAsAL0Um1at
va2nkGvo0WYU9ybB2+MwNMcbjdTOiPNtuFv2X93xFKLbEQy955BJrFA+DKMKS4tU
3rK2ylVAzZIizjICvr2kI9l2q9uBWJ61cm/x0CYHUcDlU5nfOSCGZ5HUNiLJCCxH
Re5kNKySfI2i1Dic9jpP8Uin56hs+U59PqUSDlpcB3XXbNeh5SX4Wkiv0PEuPiJn
rxphS2zShAh8Cm7Imz6XwGNdNksL47VXxx1vrRrt9joDHVNNE326GIpfuwlNWDQv
bBC/WTGpmaww9lkmSNZFlPyM99Du1N/I8iqbN7oZxXA1L4wglOYqL096gyPsieL+
FCohSni4TAUa19cJQGEwkbXL3cRSILcjV/Zcjqoe4Um0jWf9AkiBJs4TpphFmGEM
ePp7DtiMRkjNJ0kvhRzKopjRzx32P/MHhchxbHnfBCc+Ws3sDHAW375pxAtNmfdt
i5NtCKRFvg3f4fFtsgxZ3ksr6cZb4sH/VgO/ZNPTE+RmI67dHbAepfekhMZqj7gv
VNxpZpXGKFkkV3y7FZysnPQnXBZEWBdsiCEXFRpFxPbPkPeibpZlNctFtg0zXXhA
ZiLn4hSQLcFRmkgaO7aa1GPTAIMcBIv9eBefOJMnIhzH0fNUt2SAM1a8fZks0kQT
zW+gNrNLoD+2Vt44wysIoyTWXWqWhsF0LIvWvz7MxWeTKXm8JcAIEeyFfTA0kar/
OLaUo7qI7IfIk+4EcjR1D8OHlLxjxQO7Fa+fZTkBMc/mrnfU2qJuFO4B8RiLgeAJ
vLu/G5DOholT23md0uhlPrlsNqL5wvIWKi2ZtQSGuHdWZ/3ur8CsTNWXjfA6ITJH
oqHNjFH+z8N1zp7wtoG0/V/xwuW0Jz5sTsy1rwIA8zFWJzy+aAC3LNft9S6yrdqq
ADZHtFhrcgA0wvDgmr4POdcuLeAVdPhGO21gcG7GGRv9mZyi1KUTW8tOq0Iw30W4
Ca3axnKDAvmAxdq7daKoBxn9FP2TpaBFwBdU+t9vtQzBrAJIZNQV3V0/TdSqFgje
mP71qqT7jTL2zJJrtoG3iQdhfc0ejZsGMtoL3fokSL9tvlzfNb654to0kNiiAldv
8Nf8CowFlmxJNK4DHtZTqsaMEswW1Y3XNikgP4aFhtSGxdf5YdEt6u4RowVI9FKV
3fbSe46yWIj73GwBbGlunwmQKMHXbO+8iXNXB+QWDKLy+SJIqX/oDl5xEzbsRIyz
FR8g/RB5uxusGP0gJaj3710Nxc7o+wF5vtwKFPHXSE/QMtbkTPY1dPLlzFj2rc77
pc114v+IGlgBzzu6G0n0wB6gd3FrvR2LfEb2sO9Ijw/vKuIxoHF0RBSFW2QqS5bS
fWRUtP7YQxAsC6l6xtuwM61NZ7wHIn2bn0ZGeIzE4wC4vLFfDt2gsTS7ZTdWNs4y
HjyoFSX2ojtUM41K0RRkRPaTD31nhhUv2y9UrIiIYJXsGE2wt50pJupdZnyYUfYE
dsU3U2jzTAJ7csBgj9FZIntI2strrNOYXbEtld3HKGPKzw4GXFf59JRR2K/Q4Cv7
wUcFCw1E/v0xgmrbE5o/sueazhUDrTAv/fjFEZ9DVqsPlkXgjbleP9mN4BfPvkps
mv6C1fLxF1jDawaNkLLjcdNUZ/47H8IUsPmR4EV7ZmnYf1nDpFOREo+s6R22lOHI
HtfbLbGVl4oTf7VeNZz7/NOrH2hFkmLH9dFG13x6CWp++hs8SwdRC1OEmoVmRi99
yUyMqFPQSMdmNpqRqgbtHztTl3bidnCBQirHBRZZ/c+0+zcsgwLsniSjoIvE6t9n
DGK5pZepz4nUzGsNtIixIWNW9oH8qKR37NXJElM+kv8t5/Kr74Op0/+PYfdjWL2A
0uwkrnD4SNcxdlqsCHQOrz36rA5jE0J0NVYRBaESOMBofchjZMb/oqL79I/U1Vxr
joOoXsJUJbNllh/+EEXocdkisNpuqGqZ5peB/19vqbArX4+rTZnQO0mOvN1Z3c2S
FsNutMlVn4aIKQ05z29oTXAEapAoTeeB38nzG/rNoFfC5h28j7EALpfQhpbRuxgz
JQlSbBN29+na6kmguA5R6PxYMPI+QzQ91i6H9x00kYeD4gQ4J3KGSXLfeGxPDybf
6lcOM2Bj7IMRFCIQAjQSAqeoJiEb5nEyJgWpW3RvC6TLLuuJwOJiXyonxUYRlDbS
a/zSfw57TefDbK9p7K2OF77P4HTxKG42Auq84TImRplGQjMJtTC+USw0V+OWbQRC
M11zC2o012NxG0pY8JmfLDGepYTrnnT0IQj++CICDWwj5VFTdGZkvjTHdZuzeehO
rNlJ++TiQ+7ctBLji8M6nDwW1Uwk5ETzi0QFqQnvimcWocycqZFRZO0tV45Syshz
j7Z1fAB1NeonOisP+gVRgJ5ENcCiqpC3wkp/vz2QPSfYHS2ejDVxznMKdfYc8YY2
BoyN7k6ng8bRdCzipCjT3opVrff1ME+ajxfkPQpVAqxbDrmGvBJ8VfV+Oo46GO9a
euRilm6SVAXCe3/62UmUnrz2KAVFCTYO1BB8W59aVyKHZ0FqtBpx5FG93gtr27sG
Utb1Z/pPCKnDo0A/lGlGrRBvy8GsxyoXCLnuQ0oDyURWG/l6fE9BT0ZPJVv2Xken
/OfpB2JvdBgmWPnAGrG62OsC9Rmf2B7R/lOch8MtonjkPOygWcu29oWyLFRxd74j
2W64eJ0lrG+GFxFOmd8gZSFo8ffAkxMvXhTUucg48uWfBL4PzVRsz1qXYkI3JNA/
5KEuum+cYwYG1OqkkH6az4NH8QN+vNhPy/PgHLV5qaNI0s7FLYVjt+vVO4k2cfd9
Ocr4ufMlRJVhzPbGxpx0YraSNpfvmf0WB64GnM1U+AhWhgP/Jfbt2JtCUa0lw6v8
3lp/icZXgY/E0CwQnwiMwKLLNXFR02Tc1tagiQZLxelq3yktMp6EymRfvelcz3kz
1YxcvMjyo0iIGTTIWDktuP2F+H0r2MHP9Vasbqa9qXdUHAqqJWDyGuyw89kfq6fW
+LVgo4s++5hwOJQ5BjBkyJAbrI9DM9Xz8ATYEkzYwTSVU5Ytk0u+/rUIojC8mSCc
3hlTW05tqXP0MH8r6hKl7N7EHQ9e6BUKptPNVk3TisukKaPG99aT11QvGozx9LUd
Jg+16D5TscteSEeuiipfkSwjcoGccXstc78FzamedBnRK82wvWkjfLjku+Om/ZsT
5zy/WcIXOHu1MdoPocSmgmXc468bbpFsP2x0bcYB7FWTpg87fGm9JBo8bq9iwv+L
jOY17y/OxW/hNxukDn099rDD8d23hVMVpf8TvU2Ac+two5/DUnv2YBrsqzA7cl1t
LvlVwCr1MFb4+Bvgngb5Gdw9HMbTZEVVQwZ9ILknHWom167bewjkYqArJH/odnUS
Rq1hHiHw7O5JTMpZnHP5VLydcOaHJvidL1HpNPoIwL86VWDIS9bTq0STZpxPQAu0
7amZ4kTHUCI30UH2oqw1U+4a2bN8x3nJ2GjjbQOPQkt6zGvo1/bRm5EZV99H09ma
SpIYG/qbokAY+qMUhLgTvX+T/I+UT3xyiEY6C2bysWywX7oobCvzT0Sztemahe5h
E595Nr69iqx93D9DetPH/VOyUNWScGwIaCxVMKYUqB+wQjqfeTm0hg19dSC7bspj
YQqUWd/0QtdW4aMeVanqET61aL1+woei1H27LYn+EsmFxObEwvo3Bl4I9Dgpg7aF
DqpMqTvw5d0ifEv6IUELdg7WcaXQ6w6NVKUjptK5QL52JTtbCnz7W//fWIf5PJEb
kCR9260+sCR/2RxJAvnfimO3VH/FXX3VG0XjMvD9ioVDfiRUR7CL8NmJxpceiqU9
iTe5Ya098x5k0H2wFDwkE9UWMAJU09BBb1igT9LKifow+eCZjMgfz6Ko9Cuym+Dd
WAyZnl9SxKntq4pTKClp5FTF6pKjoxSEnCNtMKWGKyaQhS70MzJvhqnxqwxKxE1x
unvsaDUigvBCcZyOEYOg6RhJHbXQu3RT7AcxrQyBtXjQXwOMJ9fP3O3rRfYfqOGw
MvKBkzoNhQPAnkPr71NDdiMXYFCilW5piqifIkPHB0GYdHbyu4iSz5GD3o/DmCvu
Rb13V+6p/q6pssd/TUysryaDyON49Ipg4llmQKGfdWvY0LXpRuQn0d5/sgeSm9UJ
tFytPPJNtYHnAcwuzIk1dXh3Hk9cPlxJnnWK6b53KnU0d5T4ocNEu7T8J6jy6Bz3
aCB3u5PRJqO7mgAftxd3mCGPl+kQ0Ff1fDTYh8Wh78wC5onqkr2UMRmHn4CcB89O
34OUN+KDCFKtQIfWQEAkfQPCeqZHovSpedlIc5qQ8aUZErr1HAcYwRiuwMdxZ9yi
sWCQpxLzOcISN4R7BzYIEJYDeC6QamLfzGIyRhD3FO74CkmBAm72KohFjQpwsr9S
gfxZxgWCZx+mEgVLb+9q86fAJ7CoygFGbSATEWEsqFyiZblq0HiR10g4c/fVuGPM
eVFjBAU3bARLc5PM35u6oO1HkAiQDiKCUu51/kC1GPCwIM4arc7Hf4Bc2C2LkKwF
BMoUkkkvLsSizK45Oj4m9RYLn1LW1QcXhLCDfrRZBMPb41nsI9Q53N3WnTGksm0p
YNV2Kim3w5ShbH+qbsb5YAY6DdM0IDvf+/Sz/9jOVhb5XRygRmFVQvN+5228lb0R
XUzVX9RevKzODevKMWj9m6JkOcplNlfyq5takT3Uio/RmbQbEsEeyuopNWlVYKFm
pDHjRPB3bjb8QLc/JOWl4s/Bdmqv+O/oPEtK81dazrKuBH/yM4X0x2VSbNtNLsDw
vCsFiiYS0pgsblVI3GFWbfjIAtP37hE5aq1IxTnnTxDk5JatV+mRqQcq71D26131
w3LAXl4m/NS1lIIg759TZo2CxOlya/2vxP1j64MUny/GuiuVZfKRtS5ahyjDSKbG
BH31MumZnXtDfGtR1sq5arJsjm4v8FZDfjnZVfCoXCNbRx+U3OupAhWn1MUsUR4N
fr9sb8Ev8vCQlnxmp3ygAVzM15XT8H5MtIC2D63UBO6KLR77LmU8P+7d9LbeXhzo
wRcTe8lKRRLpTv20kiOvwYk0yAlPMDZCQjb17QGZFh5nXPo/aCvkTzmpW8LgZJxV
oPW91bydyC0Q48M4HWeruh6oc1Duz2uVM1WlCBvvPDPqA1HOgEJwVGQBSQQL40Jc
i5pcG0JoBbYrxvJxx/+CjNlA9tKwe4nkAZeZDPdhBoOg6zo51AxRtnCk9epU+GJL
jGk6HG14x4A++P/Ht8eeqxtDwhRJszuvl6/mMBBUevoGgHytj6EoTujsnZxUKKH2
ULv5jnigt+S4hgcKfjSfqu/LFBS+YDB3XsUbznd9UADVGBha0y6zIhlNyTAlcffT
UoHh4KonAXVl8NOuc8jMGEyDkdbQBpYdM4b2pyunz9TT7D5Nrya+Q5BdEyNk2lNs
LBV4QwC+gVh/s8V70sc467qNje+dvTx5RcMEdLaZwpk9yCEVokm6E0mrb/tTLrwG
SZwk4FSn3rkaJQVaHwltj/odyTRGWAnK+f/Tsgp+Ve4VjbN+8uPFSWPI4a9RxjYv
uT1P4NgwBnYwgvY20NE0hpWEn9+/kLHfaHMjA7JRN4rsJWnEP3c4WJryz9QirsgL
8RV0iD6KNKUiKZS2ZfFQIbKS1tNksXZx959X984DMDdbPuiF/xpeZa6J0tkMNy6F
O9wvezz2fRuVEjLf0F2sVCA1m6jQSsV5bzdDA3sglaE8hKCOIyndv5l4ON8ZKi2S
X34kz5mbbHXxe8gUb1PGEb/2ruf+E2UXOobNc1qRxPZBA68IQlGN1y/iCdMz7JPQ
67rz8lE+foJb72pkmSlZjE0N1++ZH7mlVTq2uXGdjoT47+7kOJUAI/LL+s0R7Fls
+/rqeCdsAFWPPEtRA8A3FuzXBoYKojpTeJEWdtmysMiK0ipQ4mFerSALA+vAjMSV
+t0pBi7RlSay339zra5Zgf3Lfu7WqFYRABtkrenzEag2TAy1w1+zIqWn7liPI3dh
CyvLC4CvR4xXE81p6b/6iPQr47cEvwSyZEtFOLym4/40k+RevVe8gEk5t84z4YpG
PgUltcP1ieF0ddohHw//WrQiCS9PsYJEpNEnUb3bosMPk2j6VUDo8O8GUPEREEKf
X5IVo4QNSWZr1Z5KhsbkGQ4t/zzejlcayPlk+GIuuUWP2pLt8UWHhZOj73mpDtjr
sC+pg8tsco5K7mcAnHctwV1YDg3E2MNhovZvFKM7aFzUQC8lwqLp88S0xQWPMAes
arhijT4dWFrYEXt8FL0d+wSNMedVrnIdposx0BRXdtyUpx4OIsz8I+n+g0Dpic3I
bXd/4DG4k3th6KGH0GdiuRp69KnMn5Bq7zOtrga/IIU7ePRptStZhG35RHNbiVZ1
nSRgyEFUA3ej+mszWlUp9zQ7bp9pVJs9I7v15NcI+Eq7HXSea/7hDGQAajTpcFnN
vkae++WZhg5U7eV2MN7cTSi6Hw3Bpap0zUKSHq81oN23PgB9RkkrKM0QcLUa7AHS
DDz+y+o4jLxEsACncwtTjUSMGnTc4+nW61u75s4VPabvrACjVcUGtgjM6niPGhTF
08M0GTDsafODm1hpJbvbTaRXnY1JCY2bZKhLGXZkh2E0e8u6iGhnqM16RwQtjh91
/dTlukeLGleOo1YzG6a+5sgD6THqviPEMR3bNTx58hfIzff1SO2VzomdL0IHXkn7
nD/y+gY1bzgRT/Pfz2MlhlAjpcoV8J6Rqdnsd3d65DEPtaIVjDvq6SJk8czeLS2B
yq7DgfUYpajl8W4aWQ8nfraFGvzdWDPF7ucwR06G9w+WzrkVoWupdjZmTtFSUdJZ
ic8yn1ekbCG57lpwSVj7QFVvXAIiluUU+7iUOOst3HJEG2dx5C+ejOigsv1XOgpp
uRC+avi/uDnGA3ePzKwd3jg+JHyIPPjDCZ9Fz8JeZ4ZahPYUD5Fv/bCthy+r7wqS
1ogf0ZzkSIFiz9lYdtN+NY5GzMXk3huubfrXiFaYaClZec8I176lm9a5UdZQFt/U
mfd5koqkmNn9ZH/p2Yg+xYEpvnu7ORBWldxA4wNtg1TH774SpmXyKeZEaOyFdjg6
m9cmCqxY65FOI8k/oWi8i40YHurcoJw/ZCNkRCr2mQHV2x91dxsBWAfQXS4GhDpT
zQlyFAJJKNgrJrE07fLuazocYwotEyhoNx6hep0QD2XmZHN18jAB6rwJdbG23W3t
jgCk8PsbzJRJZu+gsce9ZlaeeXLLdNZk/s4jCN1GhG5GYF3gQ614+I6lZU0bVLeH
RzMmMxuPvSmtmb463ITWZG/6wRy0PlJ85rg2cJUljwxvywe5tjrpKMFikF5zdcxa
AzJGRHT2fCgWgEzbDwcnPquc67M6Kvl6nWqcyQ2xRRWUL7bbvNP4dSQYqV6AYDpP
kcd8xn6DKU1nAhPIvp1pGOhEU4w0/4oXE9WYgTU+ZSX+mwG0CCyo+qcnb7GyI8ef
qpKneoWxV75SFakBJMFzqL+04Bh1tKEAwshT1GlZz41cdl71YKY6y5TrITVJCXB3
MmTAV64ln5qShA5ehyqR8Vcj8tiC+PIMDvhzJbw5PZuphXVJkRf908WZTDUgOsT0
yuoSY06UevSrt5I/X7ACHeTrjPsfKw+UltQ04YadDRyL6PMqlfH1VC0skoDCYEkq
gVBV7kisaQWjBQos+WhrnprZf6D+aaYYUQzUEkfFwO81eEznc/wN10os+UEbeFNb
Fnm0vYCm02xd2FnfMiQlOeH0bdyAN7wB1DijzkdbH+LY0fl4zr2kduU5FjkOKX2m
oJQOGvz/yLlALoAp68GynFqOJbS/BMKWuhsNoal6qBTEqkbMsPhFqWAH1U+5IHUM
tSE+yl2jVKjK5x5f/OYTteVTH1Y5zuYs7erbhNqkWGLZA82D6c4eNfjHtJNaLNy+
CoR7zWd9wP6qvQ+4J5DgDzz2FuNyUUFqsQthuShctsSdGCK7yOaczruVxmAxGMdk
K/eShYgSspHQrD5c4cwHs65CTP3diJPtOvHmdylHjuvZPB0BaqWWHWovhiZ4syKu
auFUxn3zcPvSqVBqmow9RFp/0b229NJoJPGov52Qx0CsNbHexmJI8wF6f4O25evu
LXzHYQ+O9Pehsh1cSxvOAp8OMFyiNCzvQE3EIW6ED53iOAT8gTA76frRMWdEqEx6
JLbEf0d4FZU1fUgdMz+NjIgWbEiMHht5azFfuadhzJhu1bHKxhEn4eo0SQdMWhiC
fAQeZXOvWF0eLQ30hOcip6V5X7TnCK2o5PIC0qxySHITrLkPqM7R96T8iR+2lfMT
zAGWzjtU9vcG/wVVT1buZbPXXdaqiMMp1nSkNNH7TVejWn2pYAeo7AFbPB74hSSx
nEFRUzFaoz1StgtPwgrMgSCUfV2g3icgAqDKHn9RoTxMUrE8FrH9NqvUeY8Rf7k+
/7xq1Yl4umcWjX8AncHCzaNU7XouemneJH5bSfILFODFmGSHHQ1pM1NgnjcYnU1u
LndiR6mmQh5WE/u6TDkRIsSFNQ7/YncdF8zBQpkTkzus01x42ReMNMCdFftZ+ihi
AVQ7FQ1DnI9WkcAQQPWSzWLBZhpMrFv+RoWV4lLurHev86YJfMZKchUzbn6rI6OV
V6h7Mlc0DMv8i2X/YuIrS9zcBpywrFHPMf7a6uNPiIuxXc6Sthtnb8YgUnJeiJDV
aAE2sbOWcIFmtaROIK25mwlrDoDsOBUoTqEcooip9dK1bTcGWXciA6LKkgNftG6T
J86PuJdAbhDXuAnnpszkypUmU6qwEc/lQHB7oyQ7mR/vJ7SgbVKBJXhZF91Y0QYw
RWJE3oHBmzDt3GDvMQ6dj5GxCrN28NICqS0O5Sxd2KziQVeHgGmCOvV+8QTrox/2
0+Y0Yh8AoTtldsohETQQPjUru3fd0KdzPYmv8IJfI5znp6u4wyY0m1x0+bqrksW7
HdyFwLQGR54K1nVV+psvBFvPoJwQRKyTHX51AbD3vTKNYau7RIecimm5rbeWjHNu
/EXwKCcbtAytcMR9gbywchpliSTVB8cm0P8IEymboMz9RL8VKaTsdE6pUDGPYJOX
UdlXjyTJdZX9yPUCF/tybwaqXz3F+HQIa5WFvmbiW0VPPieSmNdrPVgA/HRzXAQy
9amAUJSF5Pi5iAvnMZVQtXCCcMJp3rMazd2A0m/qXkxNFSW+jmQSQCb3cQFXEJWT
vaLhpBcPU8c3e588r5v+6NZUpkwgUXjfYY+stJtGSqVCD86jRL2VA5VetsdE/UIb
9ajH4hESzu5qYpvKHq3rbKATaY+SQ7DclW4JHAXiyRW5yWjuyM3va6BMz9R3KKN3
TdvHyCTew9l75XuVXZpourbtpxcjaiGIplaQzlFrVMyyJdz3+yD5D+5VvsUwaJQk
eHNVKyYIueGPwH/kiJAEAHQxMMGutVmZT72+tAmwF81R64cmPsWOpHD/OMKASXzA
j+hYBheaM6jwZSk4/z2AlVsYbPSKXiqd00cbBgAKC1wLWDi7Fl3icLZ1EO6n7P3M
QlrkkqHfYJUlrOufAq87AxPkgqAGrMZx5QtWRAmiHJWXVR9HkRxnZAHgIFsuURyC
8hWyvhQFE5B3yfz66pijRWr1SrmiT3H2oSefnc8KpaN0Kyqg/lxgFmEyMeLVKRjE
TZKXb3Fv94DCjwkLw3EahMXphlfCqo74fE2gtpnuQxex/m5poxIkVoNY67ygkiXS
XeqrpHRQyluI7P8SW243o6LBqKbHd2gUfAsFGxrK1h40zIk+z07De600dciz0vve
3NX2viVMATkwKG2yMuEiTDtK7Su6J1NdOyDh3OhGBnB6VsZ8NKXrqhmhh+S6VBt7
zNpCFqC5Zs5vP7RvJSndU77vPkPSjZcOaRoWFwaILDC1MLckFCFy/+ONZty+1/rk
EwohVPI1+9P0sd2tnuZi2f8eVIj3J+gEg36XivTDn8AuiVYv9u+D9IsNC4kvQKp7
gTeeNbjMHgyohve3oaaMV1u8LZtxtGGPGyLYh78BIwVFzqBD7kQtMRamTiXqCrTV
7FqZXoAdQK4nad0TPT8AOnqE3+9s8wXdlokkivM3hajafT0TeRaRLrtN5mb1RITW
VSi3ZRlHvLd0H3H8tJiXSoogE/+vIfN+mdIqHpdwQsd5+O8gPl4L6pYwVc4Um1dC
VcbPvgUexUXxK81dp4/t6E9HmJVSgjL3Uo2P5E91tiYw+n0PQwGeDqKfg/VafQw1
U7sYZJXB/L4AjNqB9RQ8BYMj+XNJ0Q2+tYGTsHzIjZq753/fyya+lD35nxcRgFNc
wdmU4eYsmOeaV2/PkSNy9b0zI57CxE0APAMtMqyoysnV6ObCzUyoJsRFtyUt3DdR
i4Ryy8VLux1uhNmdqd5N8IBu583k+r3qZlsL9O2QFOh/PiexZfeIKoVTgg+fJgUX
ZSuidUF1DNVEvwBrSykTc9HLIAPT7rarynLcF6q9PspT9MCDLW90OD2gHMkFLJso
602BrYpuLkKB5N0hf1XgZbGkqb3G4XXuaHiALVplhsqF+B9rbQtKx3zgES1yN8CU
ZBaYXOckioMJBpDz/vZWipG7i5Jl8L5wYwliBpGi/iAY6c9BzqqPelP40wvZYWEU
PnhMKx233ugNPrQPk0U4xve6ZA9WoRgGp3SRomGycZCCmRu0uPHLht9LnHKl0AsS
Uf7MfiOkE+pB8fRjYEWLo5GP/0jw2Po7iUQLmFh11x0158PBDkoB4GiAKBeKwPaZ
rv+gEZXqQCQgo6lxZkVuzUeoCmgir1UaZ6FSdOoGPs8Ep+dOVeiRJTvtNECi2RwO
x8/zH63jJA2cLWrcHQTPs4nX25Rr9CpjfMDPxMqmiuZtDUBotRvI4mosAbO++Hck
JNSuiM+d+LmUxjdVCdZbjNLpETIcrfx0z/iOIp+7bpXc3oJFLLnWviCRhQ/GHhna
q4mPruXq+MEFDxRaY+BF1Az/Z/H+n0aUBwHjQi55lKFQSszlNd6vCA5XhBL77hdr
iSlywY3BYUhkAX0ch+LFDSunxg6R9XLQCI1zdAqwBzU+y9F4nxKIms/97xcxU1iR
2HvIkuWFvGfEJFnHqjYv4ueeU/t5WVplFR8lbtOFTRqq4Nl5FuORMwu91tatdbsW
7w9e+KKZ7m+rStPdXLVMAh0/Ff/Zc11yVbTcLVGa+cBjRYrmDaEEmcj4wj+64Csr
na0BQkpBzerafawsZqjz7O56svvCPPtrNOCqav87nQmDq0inKskdR1VeThdsa6VY
Zzl0QEgY2JuZmsg7wzP+ZPPly/tCoUKaSbacurkKqtwjGNzeg7hO8zG82WtVhtgJ
VA+WGFBFuoKL5RB1hNpZHGhAPq+2maafA4gWJk3Zsp42VI+2mSF0QJ0hkJKiM4Mo
Tc0V1Z+MiaNvgc2uTB9/LovULKl8ZxW1KgElZtQ3POOrO0deO4fPbMuy6wgJCIIS
RgU4VXNaUMPJW52cXCjymlg8zXa8elEaq2/2KMh1dQhobEVJubl7gXNnYowjiRpF
sefr/HNXyNU9hOLGzR8UMlhgpz9VgfLDUsxLW2vOPestAUw0QnlETEyvK5xMkIFd
rZpe0SJ0j8IU/FuBgYUbjGyFI2awZQjEIcV4lh/otKI3JQ9rwBj9qpCW16RK0jXG
K2yZU+xxUzhkeWIjlsLcDAls49t8Qq99mPjArj1yaG77uWKkXgLcWIrDeNxCeQ+0
HlzkGpF8kMjeZmRx46kSuHFfyHVfLFGARn+GMUizOE8Q6twalYQbWEcETR14IgSL
vFFDyGqvrEwNCQ2rxbeFO5Gaw1S3Q0G0WNC4BpVaHOural45AaP6eUKO4ksQvnr2
JxDG8IS6FHWzkHU9S4taeS82KefE3i8DLCCTyN4Nl2vjdv4XNVFajyPzLFedOxxP
6Tbm1XKevahCoZqCVVX8G5ybBWoWTGy+KJHaCGfa9LfMsA/a6RfYror/7jv6eyE5
/0ytrJ1Obw7OVOtt7BTxKEGd8iRf4DsoF20dAbNeYc3Oiy+s1PZ52/Pz6ie6Pimo
PZ9bNThBRfYnbt6DQuxfIcPUayzgK2ni9a21idnnxxcpCb8RdgEQ7IxhbUZF+CNv
5MpsW1LuHD9cyPRc+KcOwnJnpe0b8oEvkb7jmHOsMSM5aNZTpTmKY5VOQymBNB/m
gCwv9J68AHdBdimi0bmO+9jDH7OPNTbuniudrcZjV/qpx4xmgRfbut6+Nl/wm+5n
UH2OAT3KHnwSZgEqTiRGX3y2nxYFbjGUp9+OEgoxvb+UY06j7n+BWzxjDRpNMEYO
W5+VLVKXbY99hFjvzh6/kpMCZFH/v7b0+pdjRZk12sqzRc+Tjqws2k+rsm+DRi+Y
igfALNcwP7FPdyBUF8w6JKuR99iUVL2UOZr3Y3tk8JUN2w1k3RZSTDHEjYz8dbQD
isg5y/YrRBd3+vbyEq8vLmtbQhnjJPCM2CioX2bAfnr4So0Ug76+wfSWfa+1OiF1
rFvQ2RUZV+wi0bD110T0sh2js1Qg1DQR7RZKOqh5lzpSrPVOytOGL9moNf/CXdJB
DHKyeM/v8xmJQcqq8q9dzcGEoJhD3vxNjfBUy8MzQA1TEZ85zkK2bACbv1gCH46F
xXmv7VuCLMcivF0kPi0mXsc9JNUZN7uxRr3scclrwC+kYLdZFr5F/MaIQRNqXW3d
WeNP29Ie/qg2DFXNQzsAyibYocLYZkJ1DV7uUi1loI1NfVaoU99HhbcxmWUDIN/j
1v1POoK8g+Dqgn8weYt86tyUDe9SwVwp8lhUSQMoZ9Y8jMBrX2EgI7dcNiznjroS
6AAOc5EaDiM/KK1pPnsl5F7l/KJI6DdrDTP0NfPT6vbXGuJcqFT+WGJxHMKCvSvm
tbzycrab6O6PrPV3uBNcwx+t+sEVnvdYNQoFCYXQ2Egy1vE/AkIJjoZ8hiMr5tr1
v5PsNiivl9JX0fA1OsRwxE1OrdPIrZvTdE5ebHzzERHXWQsKSzExM/5UFiIGOY+u
jNU6sDxVwqSW0LnqSPkockt7Zx457Ck9YtxoL0AeeGIHI20Uxoo0dm+WPGuklmu0
XjLBz5SuCrey+8Dj41LYbV3UrUZQSR/Rnn3vkbR4etVKkxL5bOueMLVbo5CEXWTf
v0C1dqPQse/Ix6IqkANbSqkguakybQia3B68+z9fpz0GAYc1bkrc4fTviUer4P3v
7KMaTdOzXfq5HV1+6YSDOx4p/+dVfJmPU4nSusKuQ7Ci6GxqbmitVh4P5Xb5C4ha
XbLCK8KWGLdQJJ5waaUjshHwXuQE3Zc7WbPpAunVbI9sscbdzXhORSZmnRk80lIl
dfAA/QH0n5lJwhcEc7h5LY8f4hbqVBfsq3/URvK9wnSuJShBQU3UoEaCr8NRZ5vd
XdwTkLBm3nXDlxSo4JG8fZ6UhkRZshO6+9HNCB1rNqGnIgvb2xzPiMUupqPhEJ3K
EByxmYOX8Vk/qrUUkqjSpFmPKTHo5YCtCRwNSuMpDEswAWOzKjdCNeIzI5+QsoP7
OUIPxzWU40prKr8VUio0UuukDLVau/KlRQA6UJDqjnjW4WMj7rk7HsU4n2MwGDbF
qwimbgNq8AKdiTV8QtM//9R/17IRTkqYM3BL3v6x5NsyiqMm+UEekG3tN1OLwFwQ
NWk6se2n7iq0kdpI4viia9cfFIDO/XvsafoauBcBK+gxj7LziHNW1lpUR/9xeYvA
dQkBK0tkDZW3TNPqV4Q55wVLBXxNhJEiG6ymVP8Nxrar/Rs54tmPpli6jE/hMCq9
oMA0IMdcGS2TK7W94vj09I9kBxvA3qrYWyOrKYQZ0LkR6w9PuJzSih1/DxQkdDfW
04joO0vu71pSVaI2NKzj7gJaxxemDN/AZYgtmdKuSLoDZfZzh0/GgPnzeFnkGLHB
NwG0hogSjHAwVKCsnQdd83ZeheLRsJ2d9kGA2A8Sg/IULLtyXFLw44NLeTaNUKdK
bYjaWXKQV3dhfGKfwMUyXUBGPjko7Viy3/gkViPU7zx8atO3C0nZvQacYwBHtVDN
evye6N3a90Rlyd0mmC4thKjgYc245dljhdJJ6fVh1kUkUddmtBn5IHyXrfocn0hE
2mPrqZOJOopD4wZG2MglK6nnE4Id2uu+6TxpdJkdtRpM0tyhKRyiZwNGVEg/AeAh
qtbpyb+T6nWyVoofq3D641zB0M4oYFg5/fcQloCDTvbobmyQFUKb3i2/aA5XSeDc
NzqbfBOauCJbViOwwuqnTNjJN4V8IFafLy2bGLKPxPLC3F9rEHvtYYxSj0fwGviS
qdtH+sTD9aOSOwysNCvUjycu3nUT78C7ON7yoK3HF/I+PY4za+X5QP/zIf+snP/F
r1rOjaImDPLt6hZqOhivjbBDMveSiQoJ/WYDYY6DL37z8kO7qK5ceDCro6TNJ/5F
oFIuuiHNdF1xl9H4bHlyPf0BP7fh9pVinYFnffLKBZjLcVokiRq3KEVKQy/6hSCY
yX9Noy/KvZfQHtCDUttjq0PP19Iu8WUXjuvRdckO6DybvtE7YMQJ8FfmeJkIpGNq
c3WW7vwnWCbu5FqgWipebaIszidVV37cOyvCvNxr44xqTjDwf+eHAkfvLR6UEddo
LlB23jTufhB/VVnEeqlTMas/kPgXRfTOtXHUW2ABQQBfhz2k/6qqUS2l7OU+JUd/
ZITJmrut/bP0cLDdAguCcpasAUMvJhzMP5ny2adNJ6O97Ats/S+uIUEnZDFcYhXc
6Wu81bBDX6COuPVNpL59Z2LeK36RkN997BosRGaF4d/QX6TN+EJanCJvs9gLX+wM
ZTyshH6WZgXkHLhEKNaLjHzCN8bfWLgMeEb3fEVEhpJZ/J8o52kVtpQts9vwan3H
zdnEPnwACLgJtOXME6nNj5leVSclHhXYkMrvKmBLAY297ifdGRkE6dK6Dj3j68tY
XU2W7UtYbehLyXQw5YOYbeNrL9Ys1Mc4CUwPAs6NJCjc5SlgTrZE+UINSvNiXiHT
SmgA6kVGjP85h1J4i1+F4wqFoEkmZK/81+REu7VIAE/mg45VtoHtk+BRFpDnEVlL
qItc1XT80K7fZWlcdzsmszmn3O8Qxuq10sUXP+zdz/+Ff1mx6iRrccwH9n/XG5HD
xaYriLVpjqD0gUjKIOEha3Yicjd5ew17vUsIjokBom0URWc3lvSh185opuV/757W
ERxES/dUeAqj5QYVUAVbT7U2hinLnjDMxzH6AcXXaplKFL3yKHwZxAEKRhnY0N6L
dFyOvyqcYTkzFSIGiGBZBTTnnsf9MpW2i7QX48cJM2XGL1s3A8c9FLzUX8WBFkjm
2VQqaxqrl0U2ewtA8A3C6bFHjG+2AIXs6Uj9ebqTn5Uh1ULTe+/f6EIaSzPnmB6i
dqrHUPr+qqF9UCQ1ahVTpV+U5jKZx4aiR2ME0tkrmVsOV7YTtPaS9vckxRYS+UcO
/NXlG42deA0usTMXBLVDXJvas4kThlUsmSKURwAd8rN7saahS4+OWyN7u30k27Vu
DpNk2GPNUwFQ3xm7mab1wzdF+Q1OYU/0eB/8ENWHJ9Ek0j0kyLJGiN0HaRUUnccd
dJ65VM9LWv/KgqjqRkbDy0lOZYEcuqALM4+Al/epX2wz/htXfoxZiIhwjLPr+VB2
JAyEm98NJ/ssuya2tqReYWjYXcM/0HH423eYMjWOBwol/KNuomOyDaGAgy3CXF/F
n7O7aijk88OlBzioiO9NwSwg2cw7+wGZMK+NbQfAWhWyx7aHjeoo5sMCVpKrJizy
qMnWCyk0qIz8cM7od82iuLTMspc7DHrOO5Kee5tOBa+GftV6zt3U09g7HMx6YpTj
FdvWou5BLCQtrp1Deh+XKJnruyQoiwnBB7MusgAiWSJzR1IGO3x+9h4sn1gIzOdX
1k+EFvYEgmI425TR97hm9Yx21HYLM/r+G4NbmocLRX6y+zp1yaPb825ASiUB6SQS
jfeXlFjz+Td33cjLktBqCQ7Oo6U1gcgbShma7eZ5TX0SNIYkSJbKs51ys+CKzqc0
mLkr8/Nu5dVd1V/DiDorn6+vROpuYXfYo3DlOW1caOceuvkePugJtgcuNFn0FyVX
7J+wq6WjmMy/t/15PhB5vOUFenM1hmtIeSYU5y+fMAXVga7rhaz0JSMwB1PwUP7C
9Fr/bSO0izUUqqnVyPrBBB3ehbZuo1JSsOkljeXyP7Sfnfso40b7TdTpgJlyDpr0
l6TjrumnCkzOONXhYLqKYwVWhPFmb7sAa+HwMxoVi9EbeklYOZzVVRyImRUOqivi
Y3j1Kl1ykQvhUn6X2SXh6SQeHPMli6L3PVF96D05BUNrPhTZYBC1KKZ/8wKa8Iz5
Pgs0JDisl/yGkB3etFZyUK8OFHzuX8jxA5AzEHFjGXiP9GzBUeoakD29Jj7GyzUZ
6OF935pzUtNBp17vwkOqna2l9nnoGjIKkmm4/TKM/NoQSQH4IAEHHnKjhx27+IEv
uKbwfOY0s/M0ixUQOUnGnTbFb/LXu+lXSCMb2kfg8D2Sth5MbMI+AeY32kfxRzHl
0YNz43qQoPrtKoTAte8msuYwORTlogVRUvBPLxqDwClBQIoQvtk9adCtiJT2FIYB
nLBJgyLm6kU5VHsQ6g2MzKCbtqKOCYg7phYU4uHyHqS6DGa8odat/uvyLawWEnhV
uVw78E+peruyR/o7v6NIq4nhZ/ThAQ5ndVJat59kGg+bB4e0L4mXZ3FLBFMO8tYD
dX/QxCTOLbazij7dq1bwpcCjZhZMGaaw3cndxl7BaJ/nMzTn1l+En9oaC1JQlh2w
aiiHlFRfhfF4v/3LKDPU6l9iETmbMxI5FeR2q0WctMZ3BTu57BYKn6SIIzRpSd9i
VwgzyUK/mWxPPCDj+l/HMVKznL7szjQ8zLngX802VD71rkl1ezSTwVtATDFrPhYs
PjGEGcQ760kj4P7zl5orMPrx/PbotgYYXU6iQU9tqumCpgbiaBqsTg9Y0FM/bQYu
1YGUshYhNr0GTglYGaC5lNTO9P1i7oiPCRaB6DKw2RZqRnP0eeoY+xebPmg63ISR
tzkD7cpSRZXG8gelZKE1bCmxRdv1VXtCcE2abx0MXmBOOvBUb2KYWNZNAI/7NFFw
l727ORCxP3KwKx8VziXlJhLRTfol0lApQI7Akkz406i4W5fnLnMONWuY8oJPTSST
3MjoO3jXuL8jE4BExmzpQ+Sbs+NBE/O+IgPOdOg0mrBbfrEgw33x04PyHWg+ALq3
veQy4HtURbT7EQaegC+Iy6XnUjcY3L82tLw9aFUHlsjg7lBQjBypgJR252ay6AK9
KVuWadJuTt5Vpye7CbfIfYy/EncaiWfkEz0H9gpq+VHkoKtFxO5GRoVCu3RhC+1O
QwpdhhfwqwoXIuAZxISoSwjCkEATpQ2dVSy59vbhDCKVm/Y1ZoCXPBXUU422R7Yb
Ku6R0jcsXZZ0O4S0paNxWwqj7hICaiAqTPSflPBWYADYAYc7DdcbGKOzicXCtBnb
EEIvgkaYW64VZjaJhSSzx9H4JFHKmuTsimivdMDZ0XvKF1omIhGVW3lA8KdYJtSw
x0HNzKp5IJhIwRzE2pTK+AAouHNF7xPx+nfOok9IwanFJ7beIz/Iy3ZHi8e0x1Kl
QxchEAAEDe0iYgQgR0TA5rVTfj9in1SsnGU9KMSGJwdzjEUkzYSi4UErx6au2jLe
wuqOZTk8mDNl6p6+mZN3FtQ1EYcn8Ix7sW1NadAju8KfsdNS944mOXlpNtPWmDOC
RjG45BlMN2YMpOhoOLRnE/UabO2As0GkF6cFu/Kv0BCc9p4/9SrYN3qw/h0+LTw7
vP7x6i0HtUEEnkIsyxVLbRi1ha4bembORTknikDNGuVLdxnTuGFJYijNAjSxPub1
mwE55uAHPNcKf8oumVoRvQMnyQWm0V+SZFOAJ1uRUgZZQYdsfnen52M4YSuTcSlT
WceQoYcZ4sLnFeh9Zt/pCfKA60Ywrs5T95pMirmwVUTuRuwGpGgaApK29pYpTmME
39C8OBwCUrhaELIxY92OYHasBC68wt07UyrKjmkzQ52vXDzMfSWJps2NpUQUFthF
9Lg3hWgJ4oMPOtyCd+WkegrKfmClQGvV5xLkt3tY8WMWqkkUGNcXJ8kzO+kE/bgO
v4tYcyLVBVbe2SHCp6j9mxaMZxoAnw0L70qR9If/B7g14F9czgHdKCefFF5ehVlM
uQiNBYybhUXKFYD3GxcWu8q6/+wXlKruIpkbaM3nwAMZOqiWeAb2B9ByTSy6PfEz
9BovdkcxP4skkv4zHMaICBn8TyyMwz5fnkT9rcbnPbPUuOQV6sPhwQz3Ncm9e3+R
FIuX0ZaW0GCZ9tX5u2v/yC45qcQLv4WtUJ5bQm3eIHbxtx97vx4Mq21YlfqKjNxm
1jbePXkqjgDJ24jDUJzfMAbWuibFkcW+k7MUHV7G/DrjThxSC+zohY8qIII3ICup
RsH5bWWgNd/JA2jpjO38lGqfsYniSmY0q2lARQJGKg5uRsczFvzMcbt1LMFHBnWM
8SlAxiughZoy81J+4Iq5C32EKfItROoAbqwKP2+F1VshAjlnAkWgygs+vC46mxu8
AU+jigwyjIYhC/xumVSH4lwT8C13vepqDw5AnoUIVPcyqhJCxfLLgmy3M/WI65UN
DNofMV71cPuPSN5+KOJTK4M1JySJej3uSzPQifZIM0+cIk4vLXLb3FMC8g6YmgwM
G1N9qCM34ToqIBubU1dvczjRmbH1VdOOjNLSkQdHVck9NsWCFITGRzDRNWd4Q4XS
EhdhIjUXT32mCiz9U0wMMLm8KZl5ncaAEYZ5IZn34suGyyJfwemlrengjyYiFTut
5BH7jrcqfmOGTzP6sVe/HDa6Tm5FqUs0N0kBI94VZCPdK723l1EL9jdj1UOIcnGZ
GYtANMG5WX7Mk35OuITyOFa2FJAukHC4vQXDvVcNMq14W7JjCf+EDJsAZYcQGqZD
dXQHbCaaH7eOdluXhn2EIlIakAKWWGe6HuJGLgMuRmNbe2BrtU+suqYxTRvcHxaU
ZT3DBp/XvD/QPIGfxga/Emx2CjJh26kzHK8e2lih1hmo9LeQWG0vKaL/1IrS+jim
YTH4437uhmkJX9tmbsxLEn/n660TCnhCXanaC60vP0B0Dw60iREfOTcfiE+cH+7e
A3oROh/HGl51a4w0wzkTe5g93v3zVuvlgndbrWpqOBEKeqPgOWq5rRWxWn9hrIHg
gLKUG4H8h1vSNthXnV+fVJ1CHiWkgdJU3Mug8OXWw4wl57IcUBL64KYJbpY/f1/k
SaJyF94Yawlqy+V2CmqX/ih4nbBNoCIlOgFwZwdgVYCFg6czGjx94PagbjMPiDv+
tPCUYMD+XGwEad3m7C2JPfwaqBwrTI6f30vpw3r4rCasBqmgGHeaepzNDVIeSzXC
TGxBHMYziEGYg9bQBNwmUHJYQxPTEG+I5iPbR88u/qAIdy+HNtnw3Mx8rsAQS5Xg
L5fcOb5sm/z6Ak76/mimVADlHcQ+IIZAPQlvsCfBSWI0H2NnkeLvCQbd9Yek1k8W
CAhkdXB0UgxDEgyW4xjyQ5elC4yAGBq9tjTZW5tM58932PqAN5oUJgcju5RZRlrW
TPFAZSIqD+fPEdVGT4kmN8ngS3IygRGMyOCZZPjYNUkYzPER9lXAQ9GIU4aBR/1D
feSbrAP0SJmKSYvRS9fyXKr+Ri3YTFZCFLfcS9c95bNa/7Ys8PVk2/cFmJKFGOZI
Ki4/3UGBJqNrvkKq+zswX2VA/SS5RbE/YnY6sIGIec2bS26tzrWI/NpBwBL3fiLf
dl8hRZzXEewdC2UB/FaPFuZiv53RntcqJxz4rnvALcvDI0ZnVYOt9lNVhOi+YJiu
KurVlPMNdrGuUu9MbDOR50lmsd2UFgHgFjUvQZGcqBxFU1FSwef4qbtrefVZ2G+1
PrBch/9zStq2zjcjoOjkzMBuCrkRE7JwHgr5przCsOtM8jbMQstlLW6FBWWYvOwi
BjR3oGI1mtkgraJij056zRuF7oWXxXgvQGgvmV9dASDMDTTxAEOiIePmh9y3K7v1
Z37RtkNF2oRdR9lBo8PY/E/SPSw7g4zJaI4McBAiMQtf79HK2gYe4TWrYOg390qX
2/cI22UINSFn2R3Qfa1mmAu5TOGrLeFT/4S2tmG4kGxx+holHhfUrAhOeGuEHwuG
4syvaF5On/+FRpToaY5oeEcxqCnMIu0P7U9P8SFXXL44zng/fGK/9ndXLSTCxBHX
akWRz7tS6BHLo06hvav5HSnL7EKPFujQTgtKHuGV2PKcye8h6WcHINBPK9RIzAr1
Bx/whSBHAGmGugFPDi9BBYu64Fj/uN7Nldypmc2BimscRsyINXJ+fr1epM42RCec
BKO6WUiJYFiQdWtit3UTL/zIME6wREA21O5EQCzFJCfxM3BFZoNYiwJL9cLR4q89
OVyTs5Dckar3EbYW426s2icN8JbrXno7wfZ1AjxmYqU+tBaOc01BULsfWJpcSDDb
IuXp84vlFSwkVsCezciyPQ8qVBBBWqYOwJQ7rAqu581QLQ+KVI1vL2jbNNOTGpqM
r5eSb6sTdC+g+dz1BVrRa2M8ftWe2HmTWwn7acZ8fFq+IjMaWZtfVeqKUfujrL+w
iHwFQcdjZJUjWjVBBfvYaxuvcCFat23UfUjB3dk4X3yCnBYzExYhCfFrM33YxyrG
kx6R9tamCx7np7r+5F2UhWwTXqazt2i4h0sADmtFOHSAUDuPST8J9OzTBDPW/iZ3
Cd3Z9nfcleQzv0sy8MFF4EVmCQcdjExJH2NEhSt2E6/VjA8X/JqNm6s6NLh3DqTf
MnahuPcdCvi83Pf0FnFaduz7gXaAKf0nEF2YSzmWz89Wsfl4BjCuntJ1BdjL6/at
rtl/vbvcQHUeih7oQ7uUdMnrLMpe+IvL17bYs8N67tAmisfmfQsJSpUCdNI6Shrz
XsP29A9l03+0Irchz6s0IrDtxamFRtMMWqND2ozhpeLrTMzDN3N4dqvpR40yL7Ig
Bn9pNUGz27WJ/Ei9AIL89wn0Rgjiotuk75z9jz0Cs7cz0MAxFfGIVTczyM0sCCdQ
QZ07daE+bWXGhi4I/q0Jcw+vmzRUA2HktAmXBP9U0kgKq3EuHDc4Qn0AA/3ES7d1
f3YnaidfoyqzyBn0NJloGcc4m6cb8r0jKhRdiIgN6F5Rg/dyJcYz/+qSbyZevQwJ
VbDXIIO9tafmSMN2xCQNh1Mt+eX3CXhXNScTtDhgowXFSJpAoXg4ija79r0OHuxT
ly7kKhxKr/TrtVaArrBbjTsA5Xy0RBfopaO2iGzUtMkAPLdV9u2N0I/bagVjFptX
5ALQFh9DcBEaKfXeTfGX9ICnzz10yfGJfRwoKLOm8G9WesLuUuckT41O6s4X3mEC
J6XGQ7bk4hvvk7m4S8OpSmNY1EbWg4mNP6O//iOdghg6HEoDGOhoLEqjnJ9fvXYs
N7MXRukFtfk+LRkX0dKoNIcJHV7MVXMDRM+wmPHqxe3Aktq0O1+X7kJaxOK2hXDk
+ApEYTwkvbWWaXyWhW0GbnGhH+Egs3eQEVy7kG0TaxsTqrNXmwKjb+bStc668Z4W
c+DGfp9qaCGpZZCe/3UyNOfFdrHtv3ZQjnVWZ7JU4B5KWcNgePnXNuE4jSwEfmXQ
THdbPo0iiTIq8QiLibfqvT9Ae8ZTcQ2vzV9D1IS9LEiRjCrSp7P8jP6+QNcBfDIO
rPPiYI6gYfXza0LA6KghvKRPndXKlrPk2/DZRy0DYeNRWbcYPnGfHfslcqWC36Qs
nWYdjzDJScaWiVDfKz/1fC9a5tkrBjPGX6I6UZjIPK+Ho2GwU3Egr35NEN9D2cQn
xfECdjwhOAMFQi2O4FieNm7YKu2yPy9oSpX/9XLLjoE0ubz2sFbtyAuP09y0F/3M
DvKpxavYVWGWy38sDShj3FI5SYKC8VFXWZsUk1KJvrcgMB6dvYuokIT0NIgAVV2I
mehww9+YyPi4mb5+lSDJh3FpkvtaEaqt435we/kV4C54vUXLvwSHF7BOtEgtI94l
lC8c6uI8yyQt/aJXT3rTBnhfOp952lNzj1Vnxk49fv0F6BWGpxwnsvwN5caWv+CG
cMozExVSXJbyMxT50pRRpxrizSlosDJyz+zP4wAvHyGy8AYKqJoTOSQg6NKl+wSR
jPMZ03iInS014ysU02ncStJldsCdVvNJIneon1YHYFgGouGKhzu8K1d5rGRN2Pu+
frg6OzeF6LKJOZgEQmH7Bmksl98bW4Q+E8GVRzeQAnPb4oy7MXwSycShkbOtDRb9
tqOHR3r7ee8K9BGp6cMX4uxe768bPg0jwkeP179fg15dSFUdVvC41qx2e7hPqcSI
lZtBkcsSDD+HT4129IKeB4++pn/d0NXguA8ofSytRHM55Y3sEMb3yjUzpkZK57LE
WtfIOoL41+UTNYnFlLwB1mNd0BsottyprjP2AN/ctI0W/w6XjgalIcWX9TropMD+
i7rgE1C1CRXTfUNGILpEOoptprh3zaxGAWyxFxCBYuS5Dj2jB5JPDTHyC6mQNXnJ
RiEBxiQhy2YAJH0ExITLP0E4aK44o13OuLWum2k605+8Ob92ydvVCVIA68lxBYM+
rTNrh5hJkLOdR0qAtWiyp4+bEPHL9foyfEZvnGh7d1X3vwvRTY+PFCbKIT2c379U
rlh7simhR3u+RSxVFydXDczQ5xY52eQEz1LgiPsgM8qT6yVa7nEKH9gVm5/EliLL
I4xxzw6qClJ0fH7Wtk61Im2YbFUlp1tm7UIhJ4hDRWUB0MH60v/PmaE5pkFmKKmM
3cbqvZnXPyfRYK80yH+TSqJGbx2UM/qElGXRhsGxXv9e73zEHOI7xkwFzjUe8PB+
GYMIsmbs+XwMuu6buoxZ+Pz0nf37I8qMxJBPD9L0nv2C2Zn29TMCrWw6QsoacoO/
Fr2FLoEhofxjszs8rHzNepxmxpTclV9UgO71n1Rx+sUmVQ/1oDS+ZBgmDmBssYFg
0pSHZmUz5YEuyQH2J37ha91WIdj12xMzucBs5LUpqEYorXr1ua0wrUd18xzYMoUS
ZsvuI6HM2/k/DrDGlrlHPb/uKntOxG2988ieW3qbHLSc8uLFK8SvT5TIskv4qVbt
WIxP71QVuEUXy0co5HsJQrliv9DzmiX2e5YgaLWxb9kCEzECPuUVpUZycR+NCieS
VEM/TaK8aDfrUqI06jNi3rm4Eoh7K/twQpmzBkDY1MrVLpkjcC9I1XSbKOI0IGDc
uTjpE+cHo87JNWDh3lPyKtcHGl6pvCHhRuaNR5Oumw0ZOMKug9Mf+f3qA3sCndgs
ooFjQ6HCSjD3lRjVvDiyrtwooN6rr8RhSiGSutqTRKBG7gGMV9utDEDY3UdsacUr
w0F18z7JM4Gs3fb2q9aMzCQ5HdqX1rc122/MhbKo3flUlzVFQktagjlSh3W7tGB+
s6+zazVl3Jlix/fLQWtK8wCVKP3yXtvGKSn6BZdKud50R3HFK2TuCpWTWZxbLaQN
foO1isg+b/ebqKl9aksay+ZCaAAXmhYERX7RRj7/7pXEXX5wi04zON1W7bK+dWf1
lEMf21HccWumhQ9VrMUaP9K4xbqHyLpASSpg+J10zvIWPF3GBuV6xCvJaEWQVfEw
rgopswovyrVoQm3RUjQUA1QCn2bx49QeB5Hx57TumpQZHOp9RihB8cN+VQPEddU4
DFd+NqtFeS4NuLsZ7JDcIcTnqx9NrX9EojL7GLdm0/00lS1rSRLjwqbMjGD301dc
94X2qaTUqZdJrhot8h5IpUx89pt6k1ZyQgvJxJ584exmsOSOiyoPjwCwRZqNBiB8
u6k5SIklCmAX39GM6Mh8+8CjpWZqXmh07/L/9+l36KDCfZ+NMCSzLHUjoPSRWXPE
q3ukvj9IxnbA/1E5yJfLQtTDCEVMM/XXD1pGjZfl7NBwsofmPMrXO19E1gzzJVOp
dinQUIpGp0URtliMlKdyTHhcmnzobF60Nl+LqZMDAH5ZSBHePik9ANsGSo2Smul6
IXE/cfp6B1UjJ+ZkIOrBbgO21ggIiSwvHQzHlmKxh7dkxYkkQxrf3AOl16JIwW5C
cBsehWYZoiVcg9d/EIf2DjAeTiZcPiV3jv2Q5KNvW+wL6be9WtCyCb46D+tBFEq7
Rk2rLfQo/y6jyAwo0QLoeaT2JWCF57xzmYD3F+hLEubp36y4+lMktxSKNPWi1Xne
5s2T1+4yf5rPpZqZH2cdF6pgKwxsBs/Pd2H8R3X8RazmuJIMGAlt6mnoqb9U+QRv
8+rwxfFT75UaIWb6GmyUuHpSsvxmTukELtRhZQ2JBx764iGAyaQbLQj1f7iXY9Va
qRTq4uUvppolnmQyVCC9FGZbD7ZATCHZADLrAA0W0DsFqK9wqDLdSTbXmvQOIO2s
YC8gol92YJCN2Qggv0LbTqCRRB18PCT4VRLZ5p/L75WUZhHtJDweBexoNiy30g5X
W0BtNIVe0H5Am1yfBucwC9EVlWwILcn0s3RQRgEkjqZ/szEzbAKaY9bjJPPyN4BA
r/motwrb+HX4qidUiHtTy1TdYomAsG0UEokL9H71j3yBLM2g0Xlel5A4LURshHKz
0Yx4F+bSSisN5wYcHWH3bxoVVSKR249fc9ff1fKIIqyDLX2n4NHDF7y4aSCndSWb
l7jlHk1vRUQYdfwNJI7JimGqaKshyU3GTZpxILw7zqroT/I+5VrBlWnFJFXE6Ceq
xcyi7R9blKPgqHgI+lZMpgcR+sGrclsscWk3us/Z2QtUV/FbLrHh4TIm6l1vmVuq
y2e8sn8sioE+rtBaGDPG3KopPekWo7Bo/KrHCluOTzN3dz56hsW+CGC3ME5ohp22
MpyM4sGUhJUCnEeT+TqjfCzDOEft9afVtrC8f8m4aQ28mQoCWCUwvKLoA6IMM4/6
7aySG3U1AZUJ1n2Xob+/lp1dnHDvwgp6an4Kx+McyX+B+rmLuZxBB9FLqilAyVlp
YaHDQlEfBWi99ReqFFu8GTGuTrB+ZeNrne/m+uFCWQKra34eiVV86k3T8GWziFhE
q8+Al6M9bMccF6oNZH1Cg9Sm6D5RtfNKKcKnWtLhUBlIc3G4Ce8B7bbr3faoyTKo
swQN/8bkmJN5OWCy6EH3aV+xUQ76Sq8hoeWTglsPjj4PljnqmWEhMQoewVm98JUS
/Sup3voDi/1RcJf6CvqOpSvai5IedZ31B7wTQCuGmHhEoBMuLFXUsW8aiMa/tLIW
xLZ6ZPYgShnOdnlRX/trJq/hgRvqdoxKMjfbLo27z70eKT5cAgaqzXk470wQLB0S
tGMzlGrh1DlxYkBTjObFH7uVclLdwLIbd5UR3UiAP0Et/Nuv56esceTYWKZtCEkE
360hp/7qLbW/ydjKkyqXU7Jq7wsvbSh+4ZWJWi4euksPK6sZmGINh9izAD671nF7
+ngV5Ijym5vit05w9XlkiDYQvujXC2rDjisscvOp0IrO9bNl5bsyk4jo/yKCn4V8
Sdtx6R32oWL063UaCihujbIXeZaJ2MDPbTbEh25YI2lP5qwMtWHwh1VuuXxEf8Y7
T0jc6e6f8uTalqY4E4DgMoxXNsAuqJA+qua5851QxZuBuKy0uZJShdF7suo6OQBN
PWHjPEoQbpFKbeMzZnPJgPv7NLswWsouVlomU2I3ti4m0drBp9LOh2OzpWx1QLKe
ZZblYKB2HlktEovYude8e6B0avkbdJ2Q0Mp+uWQGMoWxu770319oYj6z6gbz1ekB
+ClUJKrbGvzENCI7hupFTsNzPPZtHgyzeU6+hIl6RdKSTHX5VE4djB3Rniy94ORq
5zNW4cmbx8+1vFjx6CbSYjWQ+Rv2/Tacopngs2nbWFwsWymlKD3sYu/PZc4BDGlq
lrv10I84BCnHmRe3GMwDxstotujP5vxlyXgeL6VMy/c/RzQyFWqwVIqtiNU9Ibo3
j7qI1aSk7FwcUJqNBeHVw5C4yGnPk3rn9JEj7nOdqt6ssDT4QZwsperzGe1rxF9Y
kkTHltv3zHSxPwH4z55B3PSA7CiduEUH9HkcNHaOp7Y/dcBNKMTxDZWdUN2HzkwU
TSJmLGMZUs0D387C3nz4fNzWYZz4OjrMWZfnCWL3ziaX7gPPcYm438UJRuuSsERD
t+NnOT6fUIph4ok8vFHU8IuGQYPgURDuPplQj+Akp9WTyOLOhHziJIsNJGUChClG
50sbxKQH6pTE9bvBJui9iZERhsKWgNWXdZs+tvvtVQAr4Zsy2icoEjOqjfpm73M+
LSzfiXJYSxohB/y12OYHxMfRJr+Ax0o9uHUUueIKKYzX4Hh/yd/95fr6o1nEGBNd
ZnNkJxo/eE/eGf67O4KF0EKDeLcsaLZvqNKZyBJC6EktBpMw5kdSQswGqJMam3CT
814G4817xPvQM8yTECJeQda+36UIIvwEZfJPZ5uydWDBM8k9LqRZ4T0RSCOei69t
dfv08/+DHOmpi92AaaUlk7aBMduicqPD3uZKS8O699tMUR/1KN2EV/GoSe1vM0Mx
Jtxj/ts/9GsoWo/05XBJJ/LPNvTmkrohKhfsXclve7tuIJTP/frmHawu7LndjWMS
rCdzbg+T9NVqagC68a8QoAJO7lgQjbTOyshPicdJPLCBgzy/5j4fwZJkSgETRDod
SZRhIF+9fvmQBPFd6Zddd8qfiR7Cr8LZB9S6eTKodwSJAROeDIXTkhYJ8i5GNBBS
8H4BzT669pLJMArQ237Cg7lX7ipyqgnV5fI+6jAgFtq84vtUnTZGq28kP9RxqGfN
bi1WR/yjC/S6BC1fYkaJc1Je+TD7AoNnUIi9PdetLMct+W8tqVU/9Gg8L1w7g2mQ
/i+AyrL9kyp8LODsjO7dnELb0CYP8QdAarfnj6bwHPIbXQJ9aEkIimqk5aJ5WHKo
uwXzL1iJIIEFfKj+NPin26fogv42eIb7oBiYh1Uzz9GPuw4nT88PGGpZ0Ay+oxLO
f8o9j7+2AkbeHrAZuyHfyOVDzl7Llb1/mMt2TFJlrBsItLWDkOSKxaM3wPc9Hkh/
PYQ0G7UI/ZSHJxNRjz39bMmH+uXFiqNlr/DZCQCWPo5HkM6i1jgnVNe9LnzLGf6T
eX7DFNCyiW3d/g3HoBK3i1iZzo3Dh5MJve6LaKBj+lwQiOpmf5egQyNpI0moBBNf
Fvm0WbKLonuJRDTLW9MLSDMmFrFR7oEn6DVCopFSlYPHbYR2L9eedcK3+mHOxr53
HtHno67Irv172QeG6TA3uR2C8LBwoJpyi1l7AOi96lyLkfWw9JkacZ3QdvC2nh2H
SHl/4un1uVz4eP4GRM/3k9eUfNq/FqZXi+DUAggr4DAbAm0hOoVGGODkf4Kas6BI
NSVNj445jnnSVLCOmPZvZas0sVbP+dw1X91sk27wOCJChE3ujbA63TTXwiIbaNTP
kFnPC4bhyUnqY33CgAHfXE1VFf5fRfYJvCb5zyGQ7FG/6gK6FlxVlBTSDNNuzF64
YZD5pNL7uNOoua9v82I8MF3vxQbD7+Y5le2nmrGJihlu+a38Qyo+VRN2Pn9bSNWZ
29Qk1yS4uNxbrj9pSBNioZ6jP/M9hwbTMPyO0YyTqH20f/X5ueL6O+jruhjdzwmO
ZTvSGfHSo22wVghMji+9ewOLAPqtANetRWjyxu/AUEE1TTGkqA1eArLfTmuNbwpB
5r3euKMjBoMJgNFoR73Y+V+m7Ur7mvxxXLq8cRAlnVAIJnTTiCIvg+CcYXnP3psF
c+wNBD69MVv7Gw1OPZLxB15UQ9nR3U9UUVE4yYkHiYHBazmnlT90MvEZBjh825NV
H67wGoxPv76BA265RhSZ08D0qZVXzP7wS3F1zKtxXRBj6QGlMWOrxx0XodfgrDgP
y6Tc1uSmgqpWMw1GhD4WZmH0uBtPneBghzathBKGr6rVVNOxvxYGdFkTmhLcR/1Q
/hYVtGZxsh4mPSyk6wv/JK6zT7c+6PsUdfw5CT7JZzFmOtLge6kXz7K/aS4kXhwn
MyutBJMx1HavbHIs+xjNUBrqcX6tIXklVqh2Ek9ZwGP2Zd7MkKcHXpYrpaSUw+mM
I2RDZ9CHZupec4KCdNGyScub6eVhJlv1Cz1+cDNOSWBwUXTxinh6hUNr5Z48IVwZ
P8tK4cXf7QZcS+pl5A+hKgRxWXhSQ5VQ1RRSISnZRA6PkXUCPj5Sz84LqT7ZNbly
lx/on8qPiLIjZDloGZZlkNEUMDuNemH7PXFi6NcLs0DB4eVT4XCg6pD0MI1Txh4u
mXWspOdSq7u4a3Aa29P756uq3HA+LM9A2eKSCtE40tHysBwAp4bzU4y4qNy4zIVi
vr0gYz0HflelFaSbrKaor4lBC8C3ZAiA92SVFFjtbXiZiGvKKMu52f/LOc0HF+en
RrTcz1Tjz0p6rPM/apqRaeIDLJbI5QmwLLT52AOpyFMu1z397/jC4mE6V115a7BJ
La5k/+ONvxGR5hIxoJOm0mNzxJaZ+ZGpj6sl6ypybVcNUttcjUjFhn8LkhblAzA9
AoAVgUuiSY3BArxUN68JjhqscMSRoFITA8/kmU+qluXIPy5Ud24jhHViozcZSqbM
xhdc+TWYHu3MB/+j6ns2Bd26D5S0ZCf+7B/Y43nWpO/h3D8wRS4JYb1+y5sfO9kl
HN0GRPQWLdS4k2qobhJoHccy8W13pnAoXRCz8tKn561zIqCC4Sh1WVp2i9fvX5RR
B82QVkV/3tNCd6sP46P/a7weBjIwueQaqtJindeXerKql0hcc27AcoamFtty1c8A
/G4GyfbAPAGxDlW9uh+F7LRd1LHWd7WL341Z7nMulVBT+gC1X0fTEIjYBgKXDZa6
xZGHUDgEr7sgfCZZ3mMaW4YF03/TBHD6bxnZ8ngoBZBlV5/dtxEHaGXNotfBNl1g
WfHpt8le+XhrpmQ7xhG3RPIQUsjpObJNOW53+J+4PMNQu5lVlIt3fi1dz0zvInyp
i1TPL6dSgaBErEergZROhY75jz6dxGGoujTFvxrtyhtEYzx4uLVsM+0zvD4ij4w8
qSr1kfvSXXaLVJ3wb9s8m7v/vJ2l43S4uYJ5OhS8X13nNy69aY5hoc023SNdaR3y
rkyaUdYKNh6OgrXkukPh8mrj41ovb1Th/874qJ5OTRuvJhkntEpow9HhYKemyRB5
nzuyCxqSF96tnmkN9UMmi/vnTqIIUihiiAW93/CyJDq18juXPyMigkbVHjShqlHo
cpd574p2o3Xu92FEiHhP+PDMofi7qZZBk8YcxlCXBhTIc2BhebUjlgPMeUxnq2hu
zeDjyM4HQzIxhaVPLIUdclbNk/MxaMVtElIKBPn9iPje1MKrUs/PyaVswDEWvBJl
QCgyUqdekthzIb9sEIEoIq7nv8HOIjK3QixfeRRcjv3QUESPwlgA1FxKahK50H83
wvQCow/bCZ5+Wxxjg/coUJWAvB67XFedYwFrhtwuOtKCznU5Q0mucWKkDdagEfxK
apsZw1YQUwORKlaML3hmseWhvk7E0YhTP1fw9tAgUJMqbKE8PXOpvIkwotEZsTh0
4hMYny9tpspgGDqe6Dnb1PaM1ytofT3ByRHEByiPMP+Dyex/LDWhCsRjUAVOD6f+
s8YnqsdzeBeqtyeaA69NKKT0/P0Fzs9dwChktI2gQvmmxv/g1XAaHuKJFdM81AIo
X+cKM3OGymkMuaQpOSIoDKCrZX6S59GiOh+GNrfNeuo8hTNF7eE2Mi1Ng4xKW1Cz
qk282osnEXwkW9eoIQmgqJBh2ik0Kl/Qs7/tgJSNu+Myb4MQADo6hFZ/U7XM0hZm
aL03BGKUzaMl1fqvYVBDOIjBAJRLuc3Qe+hIZ9Lb2mAG82PUq/7ckv3T9Ssl1g0D
qGeXTcKuVABcWGnM9Oa/HG06SBKDRv5m8lHE1hR4p+CEpxDyQ82t8uxZW76cPrWN
lx5dLagAf5z5iUXVkDFl3IhM4diQFTIzJs0++UwcSTtUz3Af6GMf2uNbbkt2eySY
NWfiTZQdQQ6MJoivv3pNvkuaOJLRkoH7NC/UkPnUUFue+t/40AKNAPyC/rL7WemK
NHCGAchDqBpcnkRDjMK1eXZT+Esfz0zIp9EidXaPdBcRgLfZyQMOQchQ6H9LzqsV
C5GSK0cBm5ymyeEyp5mi44VN0n5aSBnpSxPYE67D4Dh57ab6GoZU1NK/XVEz3UyN
yxTSl0q5pVCfRnzLCvyt2cj9IA8T5LrRI6rb7JGKSMW2vEPaBjvOtxUZGWBpigdS
Xqlg1zyCqmbsw6Qf+dofTZlGDXx2KqJzvmnAqad61G4CKqd7hTgMGzaIPAYtfx6z
Db8/pSunVErqk9iyG5yNoCGe4wjzdOV6hKzHerNSijgjwtfzNYsGyrmQPNf4cM+m
J45BnPdcOtDPP71g4TJtvs9xEmHN0/JqjLRP6lfnBchz+1XhCi/d9dPCgAGfUsku
DfZEXAZYNyC3fxiIRm27AoJZIg5gZrnP4mbarAJILKVd/LD8wGUFh6L1ep4s4s93
MmZXSZYhTcbQmlFHWhAY5jo48PO4YMtg0aXT3wHf185sDTGH910oKNo+xz64h4JR
C1bWBgy6IN+zjqd3I7chkQngwHTK4bXEMvTs3JcFFd8TzOdvKHwWsuMwAOLJnM68
6+iAqjgavz1NZCxsLyuLH0CUoazCcEH1fDs823LjmAqtO2rj6Cky8Vm103EMo6wt
PpeVUzizJjdpM88QkaX6QdzNs0+IOCFdZfndSaoTyiG0Ts5nNlzrr6gfSzMJH/jn
4s8h3ODqUNb9Emoo91BzZZ9y1RtdHCCo3UlZQMnHhF0zBrAWwT1m6NVW6LFW4g5Z
zcrEUHb6EUmaeFV8EdQuq7jQA+URCI0Zfxcn5ZSxIU7XP6XUdHhhMQMSKkuIylV7
gCI12iJ44YuXv6f+X7BNv0MqT4eYWI4LROrTepLL1PmGXofUD3v+xhGxRamFp5AE
vkvhOJyyWGy/H25VUl3dApVB0LSYDW6bG9iTW8VQZClJ6iK/qrcCs2YuVl0yhet/
Ts0pX26nCdfwdjAj3Nieqws+GjJAenLlCxeoTMwHxw4oVYWi0yFP9pIAAVjiSFi3
1Tw+OaoPpn1gsEJ0sRJSwevsVVH27nmAmYS9s8OiDZwoILxPeOOdIHDTbRWQAaCg
eTGQ9+7HkJNf6wosk0ulGpdszgsedJUo9EMDbWgZnHEKbi5hJ9lLrqbnUcuQoPG/
IpUZYe2NkaeFtUlWuPzxw9ixOeKUOII50DfgFL/bBYEcLRKWiHxp6Ag85THEwzEi
l9Ztp4tMk5snEVQryblNpnxOO2v2DMiZRvCyTzLL7v+ZU5fp70o0vZ540nIUBwez
dMCvkMpEbh/P7xx143nYnFm1+Xr2kp/nUtOMV/L2mo3NG0+QZbyrjepZXPb14bNj
kAkDMnd54RvfXXN5DJ4G6WL1KWXyAI7LAQVZeScbnSQqga36aG+X6U/+FvfZpv4d
4YAlEdOg4jdj7WdwGS2jxrEhwHzVmnaqj6xkmQSmzVrjRTDdvZo6f1qkDzNv6w3F
pWK4sjeeUBNi+wKbS5UkbQuhfrrEfh6zrqxYoOya5thhDVMBe5TrGTmci3xBEAL4
D435Er+8P/rcq4g93qYoD39atzDuQnARznu0+IU9FdFK6gZliDBLEioqgD4zQ3ei
7+UoGaH9YIj7W3vwjEJ/nhElCm8HpLpIXHp+3qCIOTjtr7baR/FfVCWZyL+JBkiZ
EXQSEi/v6uMaom1F6lq0Dpis+T9VHQY0diaKldTo3aUoxLgsjUWRm2tLiswX0hvv
Ut0fl5J7ev4mw8wwnnReVMd0lcsjO8LJt9xPezXB1I24AaSTI3U4Tg9DE93RQCaP
JCfjQIeT6qD5cqhi4KIab2RaaY8H7SqxlrZ0BA7kQ5pkfZHWUY5MAZdRaz9mZgfJ
homK3EHQ/cR0efVHblPT0Lq1Z/aZHzwpUBN0s6oV6CRBGoxF2i5vBo0cpIL8bkqi
Jzc8BP3P/mvxb/Ec17ZB9zRBugZbHss+YLqYeRNlieNGvGcy4J49scbQB7XRyYLl
dxnIxTjkgUdEbI1NTu0UdZ/ZkWSxRI0fOGOfFhZQTxzE5PLnPWMiYWYXJNlrOqhK
Cpc6NFJDrXTK90KoeRUP9++yMjjgNXo0jF8S6U6l8Q3LrANnmpj/PSnUyUPyTYUi
qP+TOEPOxqPrRGLa9HDb3w2Dvig+4FSuUFaFwqxMIfSygpy+XS5nujmwgkkKrfUd
ilE8958KxHv4AczZmyCXqq8e0RvuT9FyuynUukdK4x8Gl2P1j/g64ozHFfFU4r8g
0dd+i2WnOzSz0kV/SMd6TuZIIloJCKZr4SC2HKAv3YEiq1lkolkn6Awde0GKxg87
DVh87drmC1+LIwy737LmrghWOX7ySqm7OVaZ8Xb9TgbgwwTYkoFASvKaw+kBoCyO
S93jec2l4tDKqstwksoyrD39el/5CkWxfSy8wmmimZ9n5JNKGS3tEEsp+4h5LyGk
Q+mTJCqAHkJ01mOs+7uQsAtBuSYLGJtwk1wuuGKuDxDr1Fl7mUUaKfFtE2fQt5F3
KU6pDIcVzrsI4YppogjWInHunOWt0chupf5gvyrmgz4aM6F0tZ6Dz88MjYwyUVsc
aq0tNBp3p5PDUTnV8PEy/n6F7sNtCoouDvGWo7Z/kVWdGN2C3sR/qqxQzbllFegs
1zcCQJclw7AF45qYQOcQYsXLIt3s2cyMZi0cHRhqt15vE38UZ+sacorbFRiOSWN2
P0SI5+RKPjOc5qHw/x/pOZoDBSGs0XgbTBx/vfU9K5a8gEJH/CAjSJek7ORIxPjt
cl724i/ojHLQ3qOwgitXfKxpxQsXrWgqJdWa5qIWiKaTOSiwnLAMwzt2HDiOBPRB
/z5jCQ/AzFL4onyxS3CGdkwwpNF1yKmxuxx7RH1/zBWzrZH05qga96vA/DeasAY/
CKwVc3QW30ccoNDq+oK9khAgyoYoajWWVrx19ybH9C4RY4eClwH4T4E86ubry0R5
LEvGyU8uIWg5ngjw8IIWojmDJvto23G1eevY5ACG+3czi86TcW9lAeCTuqIFT6Oq
BPb2UiULobOZePIRBmXDXaGWEtZVsbri0GZ9+ttNf6oW2gejkHG6UG4M0+x4ArYw
J/OA3andlbI5x0y0TA3jg655wDpSh6MhORHP3Lup5Qn4szGOF4Nw9gY6AuV0ZfdV
xrOkyGsnu6PPOVUBeTt2PA8GnSdXFAO+9i4v1A4sOEBAxcHo8JduDxXCIDleVJ5+
w77V0qG0JMmc5LxDs1cg8gQdO0WHkGoGMuFEUZZL8sG82bl1Ex6qXhnRfjOVQyNc
goQVxxlFhhDXgY4bAs3vuOdxaLACEpoobPEvvEQJW4ersrO/tYRvrnvJI3MOa2eO
3AEbQyU+jE2d/BW5H9fHb2/JJhHNO2iegpQoL6AjKkBK2VU24sZeWO6iZYigHTMX
A9NZ/D6szuq/nBAcy7OzsPQYTMqwzbOhsvHzp9ydh/CvAnpDxFMAl8UY3sBOXS5F
vv+KXv+LHB3JVN+LBXUruQzQjsFlGFqvVRWE2Ai4k4k6g3bigsDH1S1P/IwluS/l
odPrHHjDqZjSb1yhyVE7SGugXVCZxGOwRaySW0L/+Z6k1NQVCiyIfR4CyovLhDne
5QufnusmMobLq8LcUkT/GnrZFriiexyVi0EwUodAfgWx9mO7P1oLijf1ohpqwt/x
ZZjprGAv3QW6lpY4xrc/XmDVrQr2Z96s0JjIH5tERhVL1ziGG3QE64EUg8jaVl2g
YRmYEcIKQ/Jd2huzNsKONUahMeUvWukKASsP54yoRSOk5LEcnogrFy5f1Ov4iUsb
qFfGVOkcp1CnekjkyLh1QmDxrR03uKFisuGiLb0yANoVA0TZqbm6slKgvtkiQEyD
tnM4Kg5aOIZnK4NKADzP1fwPOy2gnRNnnuR+BrpU9vLma54jnnB0qj/aLaPaCLtt
y5mvps/KoXgCeKpyucBG6f7oVzNoviEAm0qXWgvTYKQwN8d7CL8rXbKIsCuFfQW+
MyagMkxDZB7ADxHnsEYxoec+MN+izGZ2bOBfHJFpAvWOnqTSyXD3N5c8WNCZJxVR
DS/SoeKaSqXa+Kv8ugeteT5e4X4QRkrCpPcqGINKlXHDpbDtVjj4lUcC8OR0X08y
Ct72vpof+pl+Slwsc3TCtBWQ88VMWIQufBLWN02aChMgVTEih1oBfs/yuGTIuDl+
rJA6FCGLVWGsDFMc0T5bp552YAgc7QyMxrOssqTZlmylCtsi6dvnsB8V2pGfCQFD
RiaApxY7ieP6OQbdSBqZrNtAb4rI0sFPZlaSvEgQwBQ77cjFPHZTGPne27f2kSsB
rIWTiViQ9vA/zVNquKReEh8o3FwIencbnG5Cbw8UhpAgzm46Jde0C7wmKOeHL0uc
TIBIrGIHxnsKRw/R0MDP9YS4fL2a13rPMpbclP9Z1mOz82FR35t9qVd8Ich6CJ4V
UYDwa176rhN/RQboAPc17sZQhzE6Asbvlkq8PVErffDrIcP5d4863jfs0I+z2fg9
uFTluUf+yMh66J/GzWV5awd3oZpK9bO699jiOEEOrjCnREuWW2PQ+7jEj/hgDOzL
xX8tmnzRH9UxHsnRawXN3LMCY2Qw6/GVFHm4MqiovhKQwC4LSHWZVLVhHFhCs2qH
kjDsJg6+4y7uGS8mX1yNuNdqu8LofRzsUlssdmCAzUZ1oeNGbzpZwbWlOXmvuHBE
QOV75PQG7MgZ1APmtO6exhzGMLPkXo3ZxPjsm8h1jJMRXMkjwWcPPcIcoCK/Wss5
Iyb+OVs2pfNyr1j/iMXrQiFNWFOvHcXFUKRJrdzZukSVkfGcO7jmvCtqe+kQgJn7
+NchAbiGxy4xzyGEItgXKddR9KQoysVueYObSeyeDAW9TWz3x8M/r7kS0Qm1J4Db
681zManbWmVetbbI0o3rJuQRg3gnUXhgZcZUI4ccPXgt6VMe1wgIPGI6QACXPNZk
VbcSHeFXCMK2iWIF148vE3Fv2vtIJ35NEfF2L3hT0llxuCErmcisqqF6XyplZ1dd
9nzP29O4M5s39LF2de+3MS3RMlvwHIEsVJPbim8eyfoU9xizhE1fRC0WwMlxNWKi
n8Q2cqDUI0ApXtmnPb/Gni+JGlQaz4XLzPrFuIM2z6VX1k4ys7Jqz7OoqhA6O28E
/GDSPVWsQ4eoHYfitv5Fo4dV7b9D80IHn9ZmDq+8Rpybq9enlFNAtmmA/SCKfqsp
ImjgnTC3hRZK9gEKnavDxQlOKabMjrqw4l7SPj8ThR3KH0+rZ90v0QAO139OO5Pe
xUlcaNW2f55k7lQP/JzyzMySuiqiwROuUt/+cvx/n8TGUlo6SBT4bbby1dA3W5wP
Y2WxyF61PSNQqoVoeXEhBs4UdcGulodKo2yK3xMYbVAwEIubxihoC31uc3kjB8mY
riR9X6Ut/1/bnh9BfZds2hMSCdf86+KMSKq8ofojxWFKld4Mco8fU9OvTDkExFun
Y/QsNTRDCzF2xwdA75zYY3W2bszP97ap/O0F4QaRsaVdX2Iy2AEWP3OS4dzlFG7N
EO6cGcevxZxOOn4GtbbklbeIeY5ivFJoJv/C9H9B3Uws3TkAfuYj02HJxZwww8rW
rlJxteABamnhmPrew6D1IrmpOjSRTgpQ17MoqguPILyQqnxPkmaIEu3JyyNULZJ8
crQElwwDWeTCtuMS5dKOL4hujoUTncerri8eEfu23MuceK2skAZoVtpvF6bq4XRJ
9kBs82Bh72QU9xXDJMwl41A6LfdQyFc9RzaxRuYPcVbTIDYQUROV4CHQQyjkvugY
FuYWFVLJPHoX6fiqt3xArUWoHE07W5OaNr5iufyP8iAoxfS6vI2bIGZ+aKVhGRnk
7DgEOVTraDQJbjwOxBVY7IX6X+dIA5N407UuGoJ7luPGXpqimDjWAu/pcQLK1Y8F
BLiA5Hg9oilefau64OaCFOgPFlNjD7P1nB6lGga696NaE/FTk0td9oVtFK88wxu0
QG7JwfDu8hkXE5BvSIbmweigNbyM96ZfQeYujxDn7CAD3ClmmqrAoEABoOEGPAGr
8GKSUcYRYZZPLgZwWRic5W/2+sPAJB4oMa06xA690cosZlptKtjop0z32EA7I+7S
Q14Y690PAAhg3yD21wVLxyb6KqQWvUr/9JYHGnl4OcdYroRZ3UR3Xbmyx/jYDKkF
Kp7QYb6Avj/50dEUAtPS28ZG7VbQbw+kMqS5Z6240cDRiU46qHscxX5uznRRnSXM
umzdGk2J+iDq+0KFGt6dncE4DoRzBIT4QI0tx89U9/kRsSWHKDpjWoF+wobEYH2q
MqFn10jimYx7fV9HUT51qVUWloeiaa8HPzMMPHICYh1QqK7ZXb4ubE+9j3eSa7YR
3nmY1IJBF/3rqFW6XxpJWWeSFA8qHtN4ohEkOJVKsNJmyRI6ZisMXK45szsKbi6s
DAaTgcJxfQZSMYiRfwaUrAH1oaBfIna34buiSF6L71BUAqd9po6kvoeIOHA7Oe88
RhgiIJ8cK7miIHr97FIFSE984DEvdMIhrb0PbY7fGq3AXBAetIjqeSi+IKT6QwtI
ZFwBOSOaNfO9kjryPw0E+PlrU/guHcni53YuwNJ7PKuokcZZ6mGVgNkQDKnlDV+v
gzzIHpyjEBXq6S1JQsSGeuSKW02czPul7A45VwDzrqITwNXJ0qxiIMw8lxBvS4J6
jUKgEACUjHeqWR/HsyvrJXFxnD7PPZb/9TLiUWmfRqtT8zsqdx88y4g7mXZW9Ej5
6RavqoY5qILxCpnsf0qEVAXdAImk4gNZbIR3E/7DYHrbQCqj81tub7HJBCbvPVu1
vfLkcnNS3DP8Sq8Sk2C2MO1d2Sf1ZvFP2/WGAPIImFaCNofVdgXpQ63vwJMRmgi7
CZTBxq/YLqxFJbj/1ORrZBT+ZV3K1hm7G3q8IgdXwJ88Tpn1/M1N/OXNFrJ2ygmi
ovOd5yUHhyVg1bQL78yNnX+Axi0llRNd9gl+WmUdMYxkMr2njJ3mm/fxrMyMxwNh
2925eqgL6pUt/BEB/I4ONFGRVRH4ci725b8qAOPrabnr9AUvrq0KcayazhU+J2bS
brmJUYN+RZQoLzJexbVec9GErDQsATUMg22Ypmqc5I/sh7A3jdT+LWK8Bn6GTeue
Ce1hvAqpUoK6ZMkyy0Wy6DHDvOftgTHYOCLrKmP9dDpCW1f1XueOSAapku4zSIYJ
yqZNemn/LsA+Ot5cR+OojCAUZcOh4TW0GSL1Op/ELaFo5bKQJBTcauLWkw3EqfHP
a0Zpt3Hl12OCM7lr6Q0MZawP5CuOtk6fdQQIZx26CmuBULwsfwXbh4Zv9s+kVH69
SNLhcLCz1eYCgREHvRUg/Jf79Jia5bswXT169nIEnaV5wMh15RXVgh01cwW0BfCk
I/7XH/8c7eBwJ2aLQf8SNYPaf3Q8KCNGIOj7ELB8S1L5o8GafHNBY3CuOt8LNBrv
dECD6PktpIQxAgkd+34azaXGfXSe586y0bXdstBTiaN92my/ExKHrg9yQLp4k+oo
g6US7HQ7I4kYP729ZLqrT7WlBdntEXuIJnko58apZnjw7nXaZ1BNySoebp3KULVt
x0vU3NTeGyqqAZmAq0salNow8g/jJRa36S+vt1L4KXIFz2EoIuuXs+V1OJXRGmFD
Y3wEtqyeBEVrLX6mLLMHG0OewHhf8pXEw3HZ/q/rogylrD7OOQjOAUaX5o3q3Jck
Vz+EoADn2NOlfBwcRMFIjcCJtC/60tsIxvGYPGmypKUQqf/zPc6f/C5Jl//B2Ecf
Roo+N3ePYo4atijSwNDAsE0wlgeESMF/7KCTtz/u5Hey/J2zpTPPG8/mYFl0y0ST
y5MIa5LAYu8YXeeyLDTE++JZIMFR6vSs1k3+VauxpFxFi3rL8fZLPLm4aqzJeVtm
/DzoDUmu+7ezKqlPL8RMoYc9DCfIUuIge2PARD5ZKw5mMutm4lmnHt9qdwVIUJ5M
qMdUZle8QD8bhaJvGkcvE0BJjVTdJmEbYk1nFU2rf0OK3s2FUSiAthNUNYfBV8IO
AcJDNIXKxCIKI3m37ukRm7gTD3qGrHfW9qsMJroqlZTkqQw5q50XuJ0z329XPbtR
0OYpaJZu23Jvjv2dUNRNmB5co75eT1va92TvrsvlZPm+neLXnu4jMZQeVfMxNmNZ
wz9ze3LGH2OdJLhJaHXaQXgJLwnfSZ5vPUEMNeGcxDBkYuX6KxDlfb2oVPKIIOat
WLkWhPzBmIYJhaoHgjXYTEqiAOwHCBNq++8MhwAGNUdbMExssYgqqpYLG6OoCwAD
VrkjVU4xxYVwiFKxLIeSO6gb1NvtU4NBJSQIIBNKTrkNG026mvv775ygbliihsJA
u1pNpkTHDPbjuuyEpa8GMZdJTWB3vz1BkRP9z5WI8dPp8+5NpdAFF7GMLYCNpgjl
7czuFfTuqYQxYPp32k9qeW15ZUM2GeKyZ9wQ3CBVDAp1L6l+iZ4lO6IrxilOIKuV
7rA+SQF3nf0/ekUK1YbLVtugfBvgvxmN5orEEOfxARG9qVj8npajR/Cy2/0G5Zzs
3dQQLhKBLhTds07lR8VjvG3OpX/drJqwSHQIYF51ty6WFm9pv9VYk328M8ujDkmr
bFJkRf4aM0LURWmO0UDsSYMdaUYnM1eCY/EeSB77MM/5Fh6fngBbO1WVCo7uMuEJ
i51vbaZTGMpFpxyvceI4pMNkw+3x3Qb1Yqj7xfBiDrnCQFdVIASAqni5xJXWHUqd
FOHH22MJndWU4SfrBgC16+QZlWJDTLDFx+yMm1XouI/KqwWang5tLwV1/5Q97ymF
1e+caSWzgPGmFiC8liSvETSvkGsCV6ZBXIvo1i/y5l3Wf0OMWVqO69ed6gxNIjZL
sFpD2rpaP4/1qVzZN4cigV14SweSED7EoyseHrUM4km4JRCHyHqQyuXl8hTaNxuX
rPe9qbGe8ezx+K56n7KIg3nekPvCbJUiFtU56r7nzJNs8pXv8puep0IXn1P4DR1s
3MUz0N+U9DJ43mgLTIR/aOOaypzRsXyxdX7mbyv5th42V7iY4hgueWowmVeSgY+B
64+hVqJxyRpI5zwcqqqUv8xudFuLgQxHhMBbQSfyWMC+nEs7LdgQhQRF1HJ466Pp
B8O5QqT660xzmDfhncYrXVM0XylU631AqBRz2Gc9mm6bg9Gc5f5STJUtiBhgmDKd
eKWTsZfx6Yie4AYyawm8nbLN92tvnwR/AK9NCvBp7G1/dly0NbYPsiaIvr6rhklz
8riWJHKWrgDVja2i8pSd/84DbaWUTdv8xB/Et6V9DRG6spu6+ffkkF3OPlNlWrMk
dQuX+/Mvy4a9ISR9IdnVeN3WBFotyPbl9mlOOisUOSPKF20R+4W4+WLBQEb7O6n6
qs/3Q6cYK88noRT0KvA6WcikNE/D6ojE3A5uQyBViGV+dO2//hhrgMWyOuK2ATxV
DSVejdgG+r4A+h8jX3IJCSO/tiv7cGFiU44JQLJ0AxXJtKkzhMBbFgqvvZGtQSNW
gva+m0Li/G1PcoPkWUrQr3Qwjw90t65n17BTVVLlKGZmH6KkEXO1YvzF1rxFRb5e
esxaAJrpRHpVD7/2RJ9LFasexpi/o+rPHeoLjpVXpB6NgdS6CmCNio9ri9YzCyTZ
4shnmmsI4gOkWQCQvkHR0itqzRz1WBfW2tI44HXpHrqxNkk1XmR+u0Zyazh/FkIg
p9ZVntZuoiv90fu0fgmep09MOHB6T6d7XxE09SADrnVtmBqkYOgEZgxyKy71XXrh
0drXwf6Obkb+BhWAIXVKPENl2SBxT9Vd08da0ufMJ6Kyf/iWraTf48NXAbKLAO6J
vzgy4yfJHztx+iQ87Xgl4ch7KlnSv6IZuC19Bx30u+/BsYl/abiV2PjSTCAHx4HK
+nbTQVGIUQHWOd2EURCuRsMHjIY8f8T9gIIv2SnPL610AGv1GTNAhYseCpvXGMIl
wcXyd/uPW7St93MASnJSJQHz1Zrf/vyDn616C34aCFTdKUoh+kuOy07rAk4vkAS3
CXdC8V55HkpvjrYMLJDW/pPDaUBL47HEVmEQn+IjyPeEVh7MSpkdcLN++NQ6jOqf
BTrkAijyLDZCIHupZqE3LXOOJ8osa84kkzOScL2xFmrDRzQEc6MNvZjKulsUlukx
wCn85RA24HYF2eNpgAph4GdPhciZyOylehHQFPlTrcagLNzLKOkFgEWd7GoXFvqJ
WV9SIcuy7iBhkI/LGI44ReWFKfUAHskXoJeqQ2Fj5qbPqtgbAGxdVfuWMfjDfhLM
JfP+WF795y7ffMPU/wfue2cTn7+z8MFnwFK6cQbMTx6WPJte5afPkmt1R4AOZAU0
774S47C3bICIfeM3zBbYdyPrrEPcVu8nhRSfRImrRC801WeFHh5z4BEL265WggAf
4Xe5gcoVq3sC3PMIQWmNOja4harGyEVgBHkipZOfNVo0YkPyff4KOjZHO8DaZqVh
/IPJbxgtGaLTIeWC+aRxVMlIJS607O42sdeIh9Ruq/hU+fErU6JEVXzatCti8UUT
tA6RyabHSOruXEhb24CbhdcEWAqoQg3dytIITX84ogOxwPgMCu89z0H0UW+4JUCQ
Cd45AnW3lcoufl54zCdtSK/H57micvpecl7qZgt7aKkTphCrcQ4zBBMKxaiOgivZ
iwfv0AMhMIqmPC1E1UactGwuigPQRglEWPz95KKil5JYXAoJSSKfzKhz9h+H/gYd
Y3lgwwYfhJ5MvRaNwxyk9fQxyB5KyKPBZn6emRK1lJ6wqxfqqVST8sgkKA6JG9a0
3zmMAbbeo+dCYT4crRSPgDM/6XHFT+3FF6vaPBXKZUjgksXEoHaEJpdOO22/3pp+
RiBGZ/WwjOghkmg8qcBcqY64h6bHL8gpIaoU4ZH1tx5/9GQd6zXtnMa26WVcbkdr
KV6/yKvsmHsMw0z1ZexYApRhOyReIJzV3A/+w8RyFfRFqDx3mYLcw9y2DAV4lvLz
vHGE5U2AlCZ0++eIkOmBra7JMCS5pWfzZMsNXZH6YBiUXcxBFzlzpWHwgw1npelL
u4WrKqGct7eIwkc3htO6YzgtT1YiYV9KGawm2msriW3tzmOoEEMAHHaCWJKDQJFv
Dm1L2LgTuKzWPhHFgQ4SyJN+50TLe7Rqbibs3ZaQugHHMNlH2mUwbaefyAAPtoOL
P9zRlqzrKyQ9gndlSUWajPc2vY64sokUAHrMpm6fk/2Y/XWLDGqv7+ob0GL0wdEr
DS3aDHBUykhVn10PvIHwwb9pSRrsZjRYIEM3faJFOcuTBTwj/g9X9uVftXjUsg13
reyFhRORMmmDendFYer4ZqYd4PnbGvzE9eg8h2/BiE0ubufh7RxOvigm2zuhKx8s
HQuqzcy1p6VHsE7fHCdyfpKUTVlalkJVLObdoh+dPBXY5UXLy0Qu6ZdkyYs/feuX
DSXqENdtsrvZB3zQjYy0ul65O9ROUSXhIGSf8UyNsLICgIToE6R27WW8jufTxU3W
7lHu34yARfPO6k+bLjfhyg4vtxB3Ue91DYq+a4Xf3cbyHjK1B1O4AlAQCCOL9P6Y
YpLqiBAlwceYgUP3HmJvKiGvrmAbYoLFJLoi+FCzfwwikpNZvaq5IXazxXYJAJa5
wCZiLcDYPO9/qVBObBwFyOLmxfL+5WIeBs95N9koJfkKouHghpNy+OBW4cfD1AS0
TbWhcuFDbTjLnQ4SX6y/UcKZPWRjBkk5OQcRtay1SN6XT4VQEa3sOjEgl9CqEDjF
yJvR4r80IeTDLQ0B9RimNLtY+QvhoTr/+QEu2QcTTpPZ35hjanCxYWexm6yobxMC
9n/ufxHlLMaCNulz8PxYaJe7ERr4SONp1nJNs2skN+q8sa9v8wnQ+QBZ/chfTccJ
TFGV6rWdae9xvHQrnycRzExa7rWCdMkhGxS8JO6JljAuo1+vyhtnlD1V47OFcnE+
+geBlVo7XdhDZlQrbUdP3tYKK0Bqq58frZOTWpKMUFSjiy+b9zrD9vXiWvPAKjfC
UMnTYCJ7leTTCE8GtT/uL8eMvHIqMhcgVwoh7dyUhGQ4jpULqeTN4JekgUEOic9d
2p93uHD/zY+iNVDWgUv19YDOMYsWnqXDoxemQXVU+Fz+GiKn1ooEmYzA3KmhfEyU
DdPSLIpagYXPT4Z2Zynj7jyUak2siysEqlpeffUkdBGRGBa07RZP6I9+DSZf3gwE
dNKDdE+VBTdiWl4Qe8kmpHx8O6keaEbli5Vijl7s17g1ZWkvq+4nfGJNAtLHkM4W
4PC7l9qOCryAA726ah1m/4fLia2NzY60Qr2s4z7Z9MsMQnlLFJa2q+VUZI9d7bfJ
QI8OhsN+v2aq0VgTV9apbadyiQifZejqgeju4HWFxZWQHG4m1HPuLv2d45mAv172
YL0u7ldua46JXL0eNzwVznzJsdT/ToN5DtIqDeDzTz+XE6cdEMwxz67rFGkCC8PK
2+3rLwZ2ilsU7UEA9GiIbfccycps1pE8KE8eLsdt5sPj9Jnpgiu6fOKl7NrkgajS
rNJNEmB26aRL5X9XdMxEKgURC9X5PYym4KHDNfMXHe6rb74qKNyXnmW85YCukd2B
x9SKRPCljtmOHn6DPiRhzyjiWnj9OxeBzCmuGdMRoBVX4cOI2PD+KWKRXAXMidGQ
lE2a3ew0OcCNKXfA6HDDI2OGL5bP9T3XHaEWSaY0NLw6rG4NNgxMPu4inzL3KiBi
Vf02vNXhx4bWSbyaNN+kQCN5M6Up2YLGOFWi5fWPJeS8l7VDNVkOeEFdi33MU/LP
A5dHiu5GBio/tFh6sds4k9mDSsu5wN2QRYiUkVSsscrHfu/ozivW4fvIFg89V15J
q7RhUCnHp06vcnSTB0VjCMs1JGoJBPfjBxOUwWmhiX+Lr/2LLQw2+xc2oB5FB7je
qz77ZMo1vX+3dUcnSYLn1LXd6wyOD3r54oTGp3ULfJKvF1xpxZe63w3PWmK5vYKj
itprY058vn/QRAVoxm13UvBRGWRxEG3d7ilDOYjK6IbGtnC+mDap+R/wjH1lKBjx
v/UCkdQiQTjhaQUccUtU/0RBagyqNRrdNuupcFbU3sMySsfDiyiLrSL7yaT4XMfc
1uZxoIrgtdCvEdoSuc2008ECJPrZ+RhDH0QwPXgyf530imCHXP6OfkWP0pAm87XS
RRMISKNkinCgvbceCOHTEP+GpgpHkt22qzVJErFSdMrZU5zitR8JFqv6tf0gNfes
UXBHOdjSA0SHM0CcEabOswK6jcBkg7zgLa8rmJktAGNh8mQXsg9KB5VxaKUqlwZm
EFdccYv3hZc4wQKGVoByA68/KL+m/x5lNYmNiHkNQpuoQsD41KyTntoTzcB2uRhG
utizyFixx/RsXNNghne3/LWXj93pvaV62pK8YiHglhhacXUTdrKFJ+jp/CuQ+EGh
PgN4hUrYkyLlPt0T9BmuMTQ6BrwvpED4NHSN3vicXYkFOS+phCwy0UJVknk16CEa
9v2ovpvx7uM+hcww+PfK3rgTcbzEWFOQVUa9B6oyISkKj5+SB+WG0cPiBSicAEAA
gW6w7MwYv5U5bZMDyUEHXXA7PRixKAGeNPijBG9TCeOVu57SP7D5EEvEj7tilkAf
vct6F04zTp4NXnRkn4wRr0vM27Iv5y15k+EtIWP9qb1OmU5uclFoiQTelsVRcHzG
NNAvX3BysoDlKk+P/+7/ev8L4WC2mQuVHPBY3ek8LU11OXm5ApCrllGbO8aMvYek
JG+/sSxrou4ifD1n1gIHWirmyzpohH1StgQ6Ik9wmU39AmkbWxGBu8G5ZF4vHXK8
mLpqcIxgn/h9Up56wg4rOhkDDtQzu7HdeC/SONjX5JA79Jjtx/A4h9hI28MgjUwH
ptzIKZN8vxS6FUuY7NznXHZi51UOXKd633RhUTJ4d44mioDaV+u5AXmJtLQa18ys
GObFzghif1N06s7TFX4bzSZCZvqHyq82IxapccO4F723NTknGyAi0cKdFgQPKLsu
A35Lah6XHT0VFriVNGu6lWDvPPoOg8o3ymjkrRtBhMgkkktoo4m6hs7OZZ32DdQ6
LArNffQ62uTEhkmp4/ozjoBFmCWvLNdFK5QKf7S4g63C/pCxoAg0865lVMqp+YxM
L6PoVQF7e+26ALzfBZIeWbb/OCyVoilMyz8qrEchH0zDmOD6oPqVjigLwD0oSxkj
b8oZRbQmyd9d9EK5Tuw4VwHF7vHmKBc01iSeXWZ4JYIi/Glw9Z2uVOpUTUpWRiYd
fd6vRH7mznvxmGYnGKHDqes/zVvnh+7VKCH1e/M+PxLC9rmjgZB+qahYnMaGFQ9C
UUEzhDHewCvvBD5AQ2gnwXAT90sGGlJ3IGTHmqn/M9iB0BmENoFOIObCtoFHBzoa
KwoohwBy2OJhvvJg+XBHPLfSo3YjaCybb62/DbISrxeBHk7aVzN8AFza2j8zgunl
+DVnRO8p5WgoahHMHDFO5LpDGo+fia8kCrzaPHNBFsoQRjBdBLOt0R9EjEFuS2ca
eUscmzb19ipBP1kcaya+nw2o6XfNsxeFBVV4gi+jdw+zZR+Wix3fnOhdtxOGQVZP
AWGHf2tlAfqdylbbJYZQtCb2iTmKMJPexLoVUBINhAiky72idaxdcERCTD//70bp
MvKUiGvq7lvvAbCuvVEZv02o2YEeJqVI0v0RjbsWq7nOsYed7WHx7p5vcxRtG80R
VhxCvYOZyCMVoFiMuy++MT34uCUsnnGDjbro0WdZ2PCavMmquc3FgO/tnYksb4tP
ds6CyzNzj8ZvLT7qaE9oncO68HsBYO0VhwjcblztvbQzgi011DwfQvukbbSH/lBP
DRGJhxDT5+S85D5EwCKOypydqqz50mpTeHWXbpcclhmMqiSDITDrRUes9fENt1q0
pH4GHaJksEBitfyGW73jYMu4YhhajYVxC3JfqcUSQitqCFEZLuqnFXCLsOXb0jAM
uQBYeHLbQAhiYX3oT3p2zlsTS1XAzetOWqLUar8Txi+WMbkzjur/nR7C9DzanTXc
haOdpd1z2v+T7siwmqSXbj44ZpzD0yIMyRrX+GmIk1XVaVcWnuSfxf/CZqOVf66e
zqQdByx7GOikdRZEqAYiRcU11qle+hcp1aDhumrIWmcWROy8s4SBkt5LXSXFWZek
NrJeJkaxmuCiTiQQzGlNLILBI6tf0R7jmBt/saY8zekwpIF8OWWSDVRmu3xaUQub
pHuNo9rRsyfv41FFZ47BLlHzTWRarqw3AU6kGIcR8vHdk/3cVjpVlKWkcZ2drHZw
K1NKNeiWzxP1tJQzkBV4shvk1cQJlvw9/OLSW7jKvGK/qUeLDVNwoVKdTwGUFMHP
nGvdCoPNajg59hiAgNv8eA9+h3toWNK8wKKeb2P4hrySwVydmUrVW4/7SlFzQgaM
Zlh3YjEevxwFK3Yza5JdqzSlLxfG8tK6oLpPqPqjAeXQFUGE/Sp+N0cp8KxpJEHn
OY7r+tJuGThbfGBhOFM69pO34PJ5CafrPIJPkNtze/0T8zsuIWcIi3Jc+M2o/Tgc
5sJLzY3BWhmXgLPvF1T/fzshEa+1Z4hurlMmoaGzW4UDMiCXHyAf5q86DCMluDxx
TRHyBjbrwYWLC8qNt3JrohjWy3tju1oablRx/IA2EGJP9rWQUEV4sNNO+5ywI8Je
p0GATTcQaWY0qbf6my06xMtBNAXoUa4leMPivT94oZ/o+9OqpO0JeUtO7rem+hCq
/HjSMaoZILkX3qhMVqG7Odb00Zck3B/dIwcdzD5LhIwc7KSPz4LnLwl9UWG9YbhK
O80Yul33+MYF2kKRGt9JqEVyeJzihhsWjiOJmFKXN2KVtvhJMAORh9ARmdcEgC/4
/C13nD7TSrYb9ULqmPf/h1ecPIvYRlCs9gmdsUwYGZ5P9CitJT9nySPtJS2YkWqw
4zh6E/WILXnIQ6rMm9/pO+gmIxbzQxNqadJRQnTBfl/jIHvX90y9Rej8aVtVUYI7
BSzpnU+nHqyI4jwbQPojvM4dnYaYjjugZI7SA+VbtcLA22HiIiHCKfzfU0aPhE5w
JNS5I8rEoMbJfFZqjrpjf6eV7iaU/Pcdi6iE4Er3J2Tee47EQQYFjRgNt3XqcEp9
IJgYn1Jn/ImHPUbw0GsjPQaF+YUlEW9OeuUaYdGx8th0sK4knggca8sj2CqUFDFi
JQCKJnvhDc81XeO5pmICJOlMeGGSFL1IEZuxVAoNCIhmg3D8wpFfoPtDD3OKSpWk
DyoAF6kK3umj0KK0FYYzgkvTSgckAma+bE/ryOa3Cp+uK82a8PUWzSdHVZstPz/y
7i966qv/WKGa9ZE+s/cItZ2pq2Ji3qCavmtNe9cPHrzJ446/mrEXhxX1peJRlcUP
mGp98QT5ztDnupVyo7JlgbikSWQiq//z/BIAzHMZmzNPFg3bx2wHFU0XMd6Q+L+3
HBxbB6RpoRkztuR2o+LeqEG/ll4m+8g9oGaGyZvqBDyee7UAp5iCTnogXO+nlEAz
eu8MpZkrlsmbJOm5DmQOcixj8a0ocaBFRQaKoabwJHQbTb2r51gSlaZfC23/wIEY
LY2GXvUAt6Gf6La13+UooF+7X0gt/zea+JkFY0HbX1dZ0wPPZkngAdiRF6MBt/2j
lb460+eTYYriU753mxsyUrWrl9d52CUaCOJ4MDNl1tL01moZ4usy8DDYp9qgZKA3
AJ2i1WSqB5YId6ZdCnEYVXk4CXamzsfAwWxP5YwJ4t3ZYogh+nBxfpUd8Q2b1Iq9
/RjUWm+ZUE44xF/E7VT9BMyW1BcMOutv80ItJr6K8z9u1osxUpBZ85oQalvBDDKm
O44jwo8Acf1UVp4GVsgOCiZ4LPgVN7Sf00D3HysDG4ZPMLt7sge4xTocYbK6iuLF
3/d0fB/uHmBvGTiafhSDXhLckuu8Cck2Ci5hpmgjpFygl9leEZg46NRRkSjq8FuG
DkcRTVDAc7ZqW6lIUXnkoD3c3asg7O17DrxUNIFDeGdyAbraDS6J/OrlakTSyuTu
Hk/9xC1JV8rf2BIUgEJ1b0kyL4qKeKTWxngmgW59kiGkNF5V+Eg4KyP9thJ4TMJR
5nh+ORUkZ3KQEqvRkZxoTM9009OHkj/IXCjHF9px89ZCU0TtoqpdBge5BJ1rc/BH
2vDsHVLPBJ2t5W8rCXWAZKH438DNEDt4i5P00DEObyszKpxNQibUrxP7hx7dIPOK
PrWMWb0PYDy2+xajghCY4EpHFpOD3F3cRKTN6sZxazP3zwRM4EeAdRqb8beYFDqZ
E/VlvE6b/mFdsNwxtSfkvATHbNQsZAqeXLDIxCYKd1ZAWO9QMHTxPl9bo68pUQq2
BYqr0zJwQQP/k2HH8UHKLxi5lLVJDthNOEpesluchLlnZ7IwM5Ej19icwOL61R3c
i5V84zOupQ0e2r96LCQa4utIcO5tR25vyYyk6ZRNoKMcpv2jahQXhMcjNnF98qEr
Rfh6Sd9QsRMi88O1j148II50RlGxLx5bJWwF6+Txm6ZVaPtcfS4R3QGKvyZJP7xb
PJp+igbNbm+s7y66tfAZfqAr5muiEmYXBGub9aWQb5o3KPeLbNPkycQAXGDAmnZh
2CSPf9HYWUlcl2ZJpv6I9ONFfY1kQE74I9ivCE7bV0HZnZ/rOTQ8uEBmD4pFqynX
UWWSXZhmqhXzf+GDeSRO69yxJgi0GlPYG/bqNYSxpAaZOn/yIABug/+zBQjiGEHT
rV83v91QY1vAWN8AabQGnci3ufw2788BZi0713N0dA8qwGLG7NB/36IbOnci0gZI
FGYXKUewdmhHU2rF1xrenrl31Cgz4y4VKzo+fiEkU1hUU0DpUXRJJ1xeRWDDnQWq
hOzcPey1WdJVJbIO6t6sbPqCjk/j0ZfJSvMvzKzFjhQGH7Xa/rZHE8Cb4KnObrcq
pLIG2Qq1hJQjR7AGYtkNM8a2y6dBpi7F1kujPmT+CgCzvmLQEDpIhZuXz4a9EUXZ
lRMhq7lwvcQdsVpMc83cOc2lf1pJ0Gq9X7wOW5U+cWEKCGbg+Tgy9vlbZuDACwJK
ZoUM4wlCmVnbCCcDOl8vm4LCwBiDBK95BdIx8Qj3DXT5U6noiiX/75gIIGJ5OTBz
VQwdfMkQjdZ6v4n4cOO08Q+JmutMQchMW68u3BCtg6DSxs3swF7cZLo38XZzyxNO
/k1Fx0zAnT9Po8VcVSPGcySvaKl0FJRXaABVoBYMo9b2QXBv/JTYUBJriD5hgfwu
Jsr+HsBwcyCdZI7deeZyRsH5dfxscUhIk9MVlNn90+JsJwsIJm8W9qxWjb2gyhSd
SSQyQQGNxj9flIjJva4N2RzL0kjTdaWJbZuYySDJC732MJjm5Ap+X5ct1ueotLr0
TvrdsaUzMX71QfvQPEijJNezTvp7KlBX9yvo82JU0/fAyoZWaPwIqP74Pi0P1BLo
Y5pb74rgflHrKMQn32uhwjF6JjdLiD0P4MjyfpqWESjK9IyPwTfEE6r1aULCJHVu
eQw8XROlowFufP2iZbzQ4GAa6OcF3k8JVqmpONdqmGuyAZjAFIhs2Dk6MDz1sdt3
rjCoCpzT6s2LFi7dHrZ/+JfwwkKFFDYfSUWw2Trkq0S8xDuXn/L9EkNxpi2qwZNl
+EmW2gaxseSh2ifavNo1BotpoyyyTEI6rQ8PZZ0rJJFYZnfa0QY8ubJ+O4jZA4Pk
ROTO/syl8/PkXj8CZh8iQUQvcT2i3/jv5QEajSqPKWQmgT2vvE9WNDzG94RLa9OW
l2EwSWd7Yd5EWZuCRpPIQLqI4V1rcP91MIl3aK9aFeL5W4kQ3K0HOJN7NtPgod8H
bLAmKti2rrDbJF0Pk4+iggFFoKOcmXgr89rqUvqB1jKcqxat0Zapce6pHxsGdDsW
4PdKMXanRx+weSud5GI7RwGVKM1SA54JrGdiaHlYfO6Zzu3CXAzIbUuukpGdBRZU
yMeSQYX/2+ZH0g4//OeKVaOT/FZcUz/47LwP9H2k+6HrJoW50/f/yKU6ZeZl7w3h
dK/snVzlB/1jhIb9izzzMlcS6LwySr3T3NPcCaTA7sjG2nl7AOogwgfK1Ar7wujf
uxdAozl++vuxN0eR1/ZWGLSfX9mAxtt8KllCtyvC+3m+QXnA0RVLvBzTaDrkdrKZ
rSLgiBqc69hU8TNnWPxqhK8K5GCJDGPClayqzc8+70TcAoGXasjUj1CltcT1wj73
RCxpqsP1GmPZT+4PVva7vO9Yi2zumpdjqGpJGAUK1NnXKb1HEYgXGuVY2nJ3t+x+
yvPmNzaiOMiBK/Ouc7snGUrTcOTiU9/a3zOpUr1+LooHqvf0jba/g1sGtDOQpgh6
Lwed9uhkSKVQl7Y+CNkK1QPhewnneHWvMBReMt9qOz0nfzRkfdsbT7jJUV7YJcqr
jH6osgle9Kf/2V5jXZM4fZVULsjL2NkoHKHtxnMNoCvekh1ADjlFWGmOAbfw57od
rQQ9bUaFGi+Uy8+hH04yR28JKgEmMSQaltAaxWc5N1ih2YTUTc9eMaulWTjdEmMh
jBNyKonHKPHcsasoHV4FG35k9CzUsJgR6xWD4PnFqHWK1dB/l11tV8fXoJeN4pGg
rPR5+jCLIVLW3vNloqwqV9K0GJV2Pdfk3sgmJe0eQpMBMsVtMDsRgKmUkbK5KOcU
UOBq/8CWCQ88NTlGf8cKfCYo4Y5p0KDOm9wpY3leA9hr19P6AdMf8Bxls424cR2T
uwXfMOFPA1Xr7tLmaqPiQOjhKlJY8mkgJF6g9FVc+jSWkHzhofVlaxtnIc1TSEq/
v9/JVfo6oX/m+ZNIOUHH5E3A7PkhoPKqggA9Y+I0Srux0ARTIXKlJyIe6vklGLaq
RkSTIRmKQNgysoFChENsPHA/Zt2E0FgALYrpyijw6M8qA5ee+sYWD3z/5n6AG6PX
zN5SRcsyzQtVXoz2MNUvtQko08hVV4VBRxTezS+rST+MNG4xzcEiryQMWVXVdNiJ
olIpdhxUSz/0+gEQGV7kdzaPiv4ydTV/q1mXsEpNtQB70AZDHW1Usdl6jlc44d9+
kPs8h/XLilyayHnCXk10sAzKHIRJPvYnfZWDw65nhKOrIf4b94giZVK+DjkvYCBn
Wsp7wUcGMQ0L3uJWd/5Q4q68j1IetrLAJ9aW0Y+JerDTCWQN4lma2klBKsjJN8G5
0tODOzfYNO8VcIMkK7W5ZrsAmCRVFqBDqsDqZM111hbRyA/kNGgfuRVW/ZRjCK6v
HaHRw+ZUXO07gEaZ+B+37Mn0t21ZhyQpHhzOw1l5Ndqwo4F0KLVUrSM5BwNaWCXP
LfmhkZXNl0uzpyIgm+hLH4BIvxhx8Kn+y3OSNM7nkl+bEyFMZCHVAW300357JwEA
7L+cRjMa32ANj7KkKjfVQ3Mk+sazicj+GvU1l2qBkpIfKv7Tmchffz+JDt7Zscxy
DZwWByc9mUfq11JbG7iGwV2yqMFQtFBndKXcDTfZeenoc5DmfNKzeaSbPvm9oDOi
zFHsaP3Do7EC7SuLDkH3e/XD6r/3rrU6I4eimUGso3RK5b7SoMmG4zvmAt1ueMJq
E2ltx5Gq/XN+tIaTpslp/mUpqFIa+QeX3Z5Wymrmk9d9Tc+QIvDDsxdwHlQKi+9w
I862GnIJ4NY8IWX1A7Vvnj4zGzzNsSLJ2dtT44I2Vk+cVPu7Uq/+/z1YNSGCIoF+
pilYrg6H8m9IgUb8KldJrt+Sdy3WzDtE3si+o+i7UUUPBIb8BsQuaIkAzTYf4flM
dxRO3HtMvUANFkgiraX+l/hhRMfIJCCpKXGpFktqp/bVOs2RDEk/2cnpxszoQVle
OR0qJYUSOhwhiFu0mEcPngDwQnAkTVeowG4mGvcpk1AQ8OHhax6d/T2FUmTXwEJ2
5KYeHBhMNQXnPApQVeiuA49MYcvgCsiE14h8Dz256A5otpaMOZfaqHXhuvGR5nUF
6lhLxM1kKqS5W3Y5fBtce7DjvVshR+4LuXPU6SsFbgzNOS2oto65/gq1TlIZP+n4
gXXugaILr62OSjmwEemGiNMT0JEvHYmLn5NczGO0s/+D02CBt4jQDz+N21adKEtS
23WfhHpygSjzg9PI3L9JsD6+z/UeT3FpMfjkS+g04XGNMatgUlfqRDNlhJdftBeP
UJMnGyAjjUWVR3WMQf379UzfwlRT3gFHMgzrVsdNQfr97DIKHHC34l7KyerlOswF
LHsXdEJcREgyiIOrfT/fPRbP5mjz6Tcwh+2cxsYOQI83o5Z1boqdYpGhdWWpal32
31LJSbUQJAENUH5fISBDPNIRj8OO2csF4Rxbq+jYiysfeAygL3yMgP4NgOK+wEgP
jIbxklYrAhxHZ15h5nHZIQKBVOY9wpEwFWs8cjFIgbLksHPAe9/Bz1dkyyhcsCqD
rVkDcFN/spZe2Cuv9Dwam4KW/p3ZugzwZxOs8pGDBOMufit6QNkNQZbfN5iEAFev
YxNUz2E7DuhMDbB7EwtpcV4zNCEATmQd3/Rdxs61o0niqqiSeZOxpTOabq2XgdnI
YNsNyUpvP1Bcu8nTDXa3iwKXaNNV/2uk8dgr12TfRi84oGtMSqeMeS9MhVrxag9V
e5WQVXc8x73q6XQLS6ExaIz4jxhQl9+y4Ad+qgbC0qatc5A39RP7lCSUFeF1sqst
KHLxXPsjv1VyTx3rIygWdraSw4L8SrbvnDUkmI9MpVqYEwZ0yJ7KCPXC0txdPwGJ
UfO6yeeNIooqcInwIRpdtVDB+IofHUFlKD0c8rS9S03zu4Phra7JDpJhimC9UmFP
DuPPheQCg3fRelgToVX6FuVHKVjy4dJ4FKm/voKA0WkR8QCRSGy9lJMe8kW1jPbx
IBz9dT6k1JS/AiazgYsfOmoLefnnMsir6O5HETSlqGwmTUPGAwXYUv/irf2DCCdU
IvkTA0TotnoEP6nw3jUNPm5lAdqCqp2KiP6qVG5Ur4pGuI74eGgSBZm8wncGmJXU
Yat8OInyQR+NyBskBpsxsvM3iqU1Kx3O42gEKp/H1pixOXIq8jFzjxKBPnOSzdRd
oM9/GHBIqas6mGYsoyjC75Vmd8S93H4aTCVYPvigQS4LCOQlAQRDoDfZXbM/ciTy
lHe1GANM9KFrhm3IwtJ67txEwzv+HVe1arngVepjuKmcEYTvd7EMHd3jmXcqBlcL
UnchfRQX+PCa4U5NrMcVftpM6QIcKkmo+qup1H2SElJ3lcBJtqpcvs3FnDZcRnCN
NB37KywB76+wnuAQPOxl7a2PKemXzMSr2LCmg6AVYJMFqg34iGLfM7YSgtGP5sLh
mFd8NK9mfyQa549+Sz5PdIXf/Y0iVBec7yGs8MP53UbtfV3zt0wmWgVtLfC577XX
GfdwfJb6dsN/SjF/4eMLylo0BOLnyqmTPK36nM2YQ+YMyO9B7ocy6pgNxF5taZPf
e9w20vk7ZbVXtHBr3ncervvgWchNT3HfDiJiAf/mdjHpXi8WWMdot/WJABBfi11v
lFGK+AaGbl+s1uEmvDcLUOnVAZAH4IhllB6l7rG/sIbN/Gdk/kWuNCVyjJ10vL3J
KO6KwxSJ9tyeNRbaEF9yprC8B1LrpYFOXibanQKobhqAf804s3cYqXYO/MXmVA0e
JOZ3RjEfaWPYoppAAmAi9K+nNGnvSUvGEdAK1+8/FJFZ2cMsTsjfA8sArJJSPSFg
4xdt7VSw1fN50hsTG9XpdbpAxJzQrxcMnHkkAVWUmqzfOAvBqaqZHPJ6UPhrkb/T
3GowgKNEuUE8+GPNfHpoyV+12mbw1jRI19+LNCcSY8BXrntsUtY01ZQ/sxp5Si7f
Y8pw6ykenMPI1yFC0/GHTsr8nlmCFeaJSvJH9Yy8RHMK8aM+XR5MYyHB/L8ef5kw
TJAWEIqdQhooTFH5TF/0QoQeZguK923NUPnLBWGpTYZRPrAB5pMu7zvwS0MGXXib
fufsnCaZJv+LChvddzY80iqORUpzbYBk6QFrO+Q6rEU1AVZurcSS2M+nHNceDKLJ
X6yBDQoDjcZAOWruS/tj4rLc2+KtR8PqQWbdwZecQsrfL20A3VIip3ZYgrdlMSOq
nvtYGz7008bVBgQaZtj9MnmkC/Z2MPuSwclHE+YYYwABiVBoaffE7u9iB8gHogVF
KMrNhgYSMgJU8AMpn9VG9Z47fKxns/gGKw22t5aqyTtPJgSE0SVelz02l7tJe0Y6
yvTw/2a+ZE8Ddjl79B41AnGujcO2PLAPyfPqAry6IEefXUhtTE4qXYL+8OF2C/xP
C7h7EuI2M5zA43cRQOiokUpXDdL3ajbyCRVTeMG1nAPk1QjdKCOS8Lp7wTajz2+X
bBR+wd7CbXA9NPKWpePkECdleIsNuIDvNskEXVFPuGYVz6L7JRqKXX85+ZUN7ApT
hGhSjjzDX9UjfOT9/KP86l6qYURK0Nz+0vdrAlUrh1rtrl0uks1bAQFTrbKJaLtf
dL+IFcmsy8rZNRJvzbM7i74Gz2Pgiyz4ce3zqW0RwLEC56rNOe/ypKdiJfBsA1NH
+c+DKSjEhfopwZ7iw5PyCI0juVGEEzpUc9uF5z/eeArltt0SeQW/DgbEJhxMqSLu
xy1QiavSrMMDe1uQynEi/T0jANKy+9vKYTvjfD2JSJfQuSd9wwgQt6CWiGrJ2qU+
j+AV90sx51YuMJPqOYCDQuo75c1+PB+S/ZrlIo1mcOKw/+nfG9Ci7f9t1bQbMMCC
CFRVkC/+OSmPV/y6oPVsUBKxielUd2OIHQOo5RE23/jeiuH3koLQNHAoLkqEJ3/3
O9mRQ3GSe0zjuFziYTIpL/mX0mCkUTaDTAhVhw8NKu7m0uyOQpXeWMH63kM3K16d
notDg9IsGi9t3sKJIwmhrl6rQEYxqfq1qDBaha8qkQ+/OG5eFEYzV2jrCO7O7/Lj
NYIkwl3uxCFDrodL4AYNhgd8CJal0+yGDFLV2X69iXCBLb0sHH2MNaLsaWwPVC7F
uH5eutC1J5bWt2qPKtFM9+OUmTsgqIZE9OPs9RupZELO0iSJwp3Dgg513s8GYzTZ
AaL2hyBsbek9Dtp3/JIWZDuTILXzZ4sLfp13uT9R5Klgjeh6LSXjI3TAd3e+nPca
MPenQ6f2GrMz9UvnOWiXWxEcLjPcayP1oaCKj/rlcERZTp1JjA4LE+tDKyOi9fEq
DtKIMnSTPdEFO5UNIGK52tMSKJu21AMaReT1ptyIrDzq1/4Ci0eyub6xi0aD+v3c
aN6UXCIf9EhS3Ldu4/KBTUxhZ5JeEZCth0J0ejoJsH4SY2rTNhaG54h5WeKX2yFV
CW1ofMJe2aPp7XsHpQ5jQhDoD5nncndvq4JBxHDYBdLHphg2I275UR1WttcmNrNw
1n6IAaZ8w5JHDb98bSqIN1s8iqLEnNEZ+drDIaKunaRiT+Q0l77sPwCl37kIRCD5
I7qC81d52le3PnHyO2DQyHGn5eh+FSs/UUVGTh/k8G9RNkhLl8cIBCgILZej9SHT
JPUpbqfr4pcUR5NNNicx73Azaa3Ls/4mEVrot4rQQwZ5/PdwfOo5V3jCEuZSNT/o
bQIJSRiBNdLfqMgXmczTnVX2jaf2/sAXFtinYnB61uFns43l/mMXAzoLeSs+B0Jr
HASqJh9JfKMayMyuiPgp+4CuxAZm+9nM4343nDtgTp9XCG2T11KhJ0Zwnp6Ngiju
6uc+YhIjvR6BhnayDoCAEQ1rApwwadl2Yy2du1+YfeNoLXKYoxsKpCuGqYNCTT3/
5933eqd2mbpSVGDZ/tUCDdgIGJLXG9OgOcKw7jrSotPyNlCiGCo1LeAMXcckgDFA
jOwpQyU7aL6TdwZBPNAnJGj1L2sdqbY+39X/sZ9vzn9keK6oscqPBAXcWSDCo9m6
8Qt91erNK9W7x+b5ULmY5WPzzYVZe8K3zAomKWQdezxzGDtDscyCMw6Bq0ahTik5
zD8q/Ep8tB75Ltprx/ZaEoOBaEy2phosKJsEKRvoKtF8IvUpNbKDFx5LrJUvMqdF
awJG77ealcs60UjQ5sxrRTbahkJyewgIXrvTZ9Rt5AJnbYxKdmvdyCen3i6o0A6E
rOZjYL5tuj75du71YIYVfUCB9ul8mkqFsRvupJUFq2uAca0Ou4tula6VjJPfhbWq
tEwA+0VH1iDRPybcF46/Hne6i906y9gMTRVYmc0bBz3W5lSBj3uKUBQG9MWQo2re
S85Y9vGBnqMGQaRt3pyKPz/fKxn3pdTQKqoSZudKK0NGDbHr2RZmIYkrJCC4ORVM
foi17q6Z/Aika4yWTL+9LbRA+qlTLRiGPVvb9Td9xiarrlsFr9CGnyCe+0DUwzH+
L28VgsUHpMPWScbr3p+K4RbrD7ThVtDtArGm3bKlABlKI3by6BsFF4y0POeEolzi
zmSLkT2ZqFJWduUzbVK1BiIS01qfz54rOK3/VwjOADet3iHbU7+fOm3uufDL7R/x
Wp3varfAK09vzaFWza59uIr5+HOZZKYAnqsZveA6d1ZfJhYjEnOn3ee78OC8MdmL
xazXiQ4P789fbBuzRife94+o0xKZfCRoGXuYMpUDBdxAzbRl5vd48T2E9TklzGVq
iJd40bC/v5RWtqtTv8L6XJKiPAO/JfS+nEkqEDZELt9jQLDPO/IDhJbgR0B3JXt5
pRkEU8lDykP8k3uINYKUftFqKzbkheVnOZ4i/LHRDh68WmrVKZxFzphrp0TaoXgh
pczQUw5TqktRbZZITreNNlGZrDbZwfdtuPIcWC8EZqCl72hRQGtpCbLbDt13FiQK
DIi9xEeS1SyoRdlJ09+01TFLnslX2svB1pYA1su2S4RecS6+wRI2YQHtPgdchVCk
6iJr82bX0DNTrWM6ALzvLd3UApb/sX3qXCz+gpfzxvJTPs62HvXVP6FJ08LYRvSb
eMWW7bVNp+KCPhwb//TvE0VG2B9yt7o8ni6CcVqxhoBH5nm0C3B6OuppM5gzlHJo
LmIy4mA08ge8SIxtzoCb7rd/KDuVmcaHvrDygcSrWYqMGc/ZaNjs4xv9SZoTpWNN
qE3Z+yDTiYOK5ZizEVVfii9fwb5VHhJRtE107cmbzoREBQs27/HT6VU1x23xH+JW
FtDC00KrQJn+sh6ydLu88Xv9i7OrZj1yb8i26InHMvun91DcJh5SUAYlq2jfWYLq
4v3vewwVsq72+wxAkgjdvai8pgsj+K4YDbPf1vGmnU3d0bHmqgtxaOPdM8XdA3Rh
h26XK3YDhDnTjti6jk9/rK6w6uuKD4rs+XfTjp5slM5Uo1Z/4AAIRXbbCo+mxaye
d2IUGMjV4RFDFLo2PtOnPd+N2l6Tbo7oKo14bXEg0H2LNuy3mQ9wGJn1NTxBpuyk
+q41HGRtK/78jOMVyO7zfI2wU3zAD608aGf2w1RG4tM1C6WlDU1vFK8aYzv0ofSH
XwGyUHkaP3BJCwNKw8WxYnHTR66mneR11D8Y/ofouUfgd6v3YIBHFXY3HnjV1r1G
PFqlHWW9FcNguLe5mFKri9kdpc7Dsn/nq/si3Alnb8TbX0zxCOwsLu1aCsFREhAW
1wbFfU+NFnFOLNgVovPoqlf4Bp1piYgWucCOTWicdmCBrF4OA3z0M7k6Kq1DwfFS
bM5qBv8MbxI2UOTFt1R/WbWvgVYTAY+LGiCGluXt2yMJppes/eMXYp7KpuUCQP/n
6KZUyKuTq/SenJEOmm/UosNHvbIHTix4Bs7Or0rUg5Hlk0LKX5pZT1MqVeUN2M3y
VwYeZPMXBkAPDQ9x3q7Y6nxMnZFtoh1tHGzpcUUEaw/T3Y4sdS75JjQl1iHBcs7/
JIHC3r9ra6h5rsUYFgXjvw1Dlqq8E1J9Qmtd4P1sAuXzQ8h27Fpb4RVWSCCFNYdp
gZRewmB7h53IT//H4ovUNABHsE5wnnSxfhmM5yVtrJFZjYm0xULR/LfHRvB7UVuJ
2Pn/Kp5xAAmBecvqksR7bId4FBigTZcyTXpUxjRCpqBErx8mMpOmDe2U+RDkw4V9
A9pY49TNgtBmo+g3Q3QB3ib6RO2ZMggCCDIYp2SD/+TkencFlawAhu8ru1Y9feUm
gJebR+cS2bTdCb0A8BCHTRefxSzY3pBcTPxaKHMnLTvlRvUkVWjDlHuH5Yz5JSrj
oW5dCVtHyueAF/diAx0cAs2/df3GJVXmhkG9a6A9OcITO+y/a/EmOTn95+ivLN9H
gLwcqD7HCPnqYvdi715M+z4rzHC/JEv0Vrb3HKUh2QSWcM6NiaEEdxcwn5OcMcht
26SrHcp5uD3b6s5uCMszabqwg7uVdBcziRku0DN9YyJnWqNDZPyawR9LnISp8QK6
bRPwBfCCq5tGirL/zZ+lhj/T6k26umrRemkdjFnuVk1yAdzh4e4UurCr8MMPUNgM
ySWkx4yf5i8nydIVfTXw/NuAjZ/vDCqfdtqkthn+ku9K4RqcCdC8rJcAumo8Loh0
jpKFYjXwXtRfDj6KQhsWinZo+qa2GWTcq3zwkGMlD7nIRXfaKXUx6NvaUMDVVjYf
9Ij8ecVEHSjmPefxfMIvqmRkQ2MfFtKJl1TERFBcfNAje0tNZbAI4pzbpnjZN6Fw
F4EhPuQYEpEz6w100iAO+M6yics5s3tc9io5jDZ5pKNGpsn9vpvc49O5YyklULoo
VE7L4qLAHXcP/IWhd9lPzA4AlgQbdrr0xkaNiofyDuflOMyG8dAsqAiMSGB3yIqb
6VWIPTsVkITmeIiLZPFt5mN3oN+eeeH2iEIc7wuNWbLtHivNOSHKzUJTwRCxtX53
BtwwMb9+GMbzyxgOiPrgS9mTGpeIqAEtbPPXdB1Kbft8p4tC8H2Hc+wTfS836nRB
793GIKTfzpvrRNslLPtAuH8ks+4HYDGotC8NoMPGXoR89w+YasIVw1Bs2SuW++my
NWJaaHNuyCmxfU2KqsbtiCoaZ0pO6DcYArXGUgnHhHjLeddVJHv808X3zGjAI6oU
oadOkESFZnQuZJt6BeYtPBtdcL4nuEIzsvOBE6z4pM5wdYChQ3SeDHWYGwKfjM1Q
3RzfT/WDpVwpnFCznWXY7kVW0YevEwSlaD2y0DXcVVwrr5hCSjexpMltaESiK4TX
oA8U36cPiZwffwdzUsLEI+zw8wBTTU7nO+usOTr7zpsqFB+7l3HOkHk/v12oIauv
pSFC2/dz68mX86gpowqtMgPKfPUrQSwK2Q+PiVccsbxEL+ykRYs3yF/bjNH8xPdn
8CkOIVvjrfuZQnVALOcYQi01v1yCSoGsnqib4Ly1KN2WGMdh1ix/FACk5xOGl8Ab
kuyYxKFgSgXoayxLWSm4fwp6pJ3PddvC6PVmX/NQK7LjCIznhjgNDW8yE7yiCBBU
4UWsggCmPKVZSCBhItPYrEbOvf53uh+CxSk8fYqaFFUCa6eUeWqw+ObKwur4O3eb
xqw6Ng9/9Amnvc3NedVstik3o1xclPnQomLxotIrBUwOCLS1wZiHZyBHkgT1r40+
Vl6zxQW9z6MoZ66JLfx1yRLGWg/ok4f0G5SAQQDw164Ti1LJHav/QpcsC0Sk+csT
XwuP3xscA4Bn2qkOxRS49fx8gv7VyVYslAsa0G/vVHw+e81OIrUu5AuBFe1n/7ju
QaJtSJW7KbzojuvMtP9aCBJxUBlJ4RXHU0sb6fJVWyIA7cwx3oLG6kPWv6SRFJm7
h4oUcH677x2wFNgXha3s/x9VrYBaJfmBQTTNElyXzj36OYCk8xN6TfLgCk3Prgww
Lu9SBmi7rkTWAe4KeXtqjeFW5QYWzWiIQi/IX54Om1fVxHLw8Yy0dK72VoxGZrPr
n7ZUcDNboOSOVqQFdFVnRB9+gdo/CNucDPBF3f95rZQLB3Z/QgR7FsN5qPk8FpEU
K+dcsm5kG/6V/5cC3GAR0TJKMzK1figKXgwBeYSRX1PN5bAZ/9tobLhYSZYLb8nM
2tbnkEAZ+nWZogope+CoFVdS0J7WJhnNbg8cm8D68w4moCP8aNk50OtdQWrVGwyI
OeKAXYnSw2kWmUYIpJmB6UkXTWVZawCB0PEyJMXWZiT2MrnW5wJTJz2DZ2BpNwkr
7xKf7ZtU6OC7G4huuPT5XP4rzKBmZzhCuZANUcwogl2OlDH6Y4UmecDiIuGkDMCj
BSBF5sqFG/BRXB7HNcyNnsKhaST0qOIniLX1GOjUetfV/F4ZsHntF3M1GzI6tDnr
JGfx+PE8eoutjkM29TpSEgqNAVk4cBbBbEpmrDAn5Hn8MqoYMrTrNw3P/8h6dxsA
9NvUZAiykPc6P00D81nzALRdHjupCZ1r2A1lA/nD5l/OzTr/pAUiZbdOTYLa24vW
D72AFRKjLBJSIWHhbEpQ7G+a/qv3wcHhFeaDiaoRf5l6VwryocRkyQ0t+R+PTTmh
9XLOKxC93rrgnLuaSNfgYNFJmrRFx4Z3uXN9cfHZ9BX4RTEA/gX33ce91pO4BrvP
NRDNuZNzgYPWrtfRNTIFrDKizcir+4YHtigfd7hpM6tkd5le4T0xrjaKlBYOfH2E
ad55CPpBtNwnxi+piUAUD6CzbQ1smtOXLJCK0CIcwq1Y2apXpgDO5NAHFs54Fizd
a7wqVhz5do+hX/jxoyTpX7vPMamb6FQpaElLQvfjTI7/xFqO/qo43qYqPJcd3aEl
j4UobPktnCAR4raPL/L5Ptn1NsQ4mrzOaf1AIOhQW+yUZ1pDej/ZPPHKvUR9Vmwa
kl4IwvkMRwrqe9alQcDgReJ/lg9Sj45WKwnZSV+3ry4Y1Y0Io3DM3qx+et50ex4n
8p612BQLCqwjNLThxAyhOgI848nmC9MowRv+zlOrI0L8jdZNe9HEF8IihSPCT7TK
RZPbyERtDw7dpEt2LABUVMqIn9gDR4heeRp8P/nXHOcZe4sCHxxUlQGVRYHpqxf2
9Z+gOP+iKfDkIiMbOrZKJZxNxt/tISZVkaQZMsooC+TOvh5W+iGeOPA4WggY9pWs
yow6GIjeBLYIRJLiY6MCONG4+9DzUGQVx9/tG3jV4x31w6EBcCE4fzMFLMHwaOXW
M88GwtgtQ5T5W9TXxCbNJ2CB+29rX/kBPzor0jlPvaFuJWqCHpHGFGppKGG5421e
jMUjkVT9oNCaedaOOv9UBrdB9ZsTD/7PgROD/qf4OD6bEs9QkBzY7USzJllIUaOl
W0lQqgNpqtRYwLGEPk8UuSb7L+upiA+ieVf/dho7xa2ORlE/wiq6LYBMF1+C8RB5
JmwYSCqKtndW4Guec73WRumJt5vNzKsZ0FzuBEsoLhm+OYwWONY4Q9XrsZNoqOuA
Dv25QuJirJbbH+WRiqaw9B0hIUVb4pd4A/w1yITsgbMXXmySleYHaWu6sPYmBLzf
l7omwIlP0A9egE08ZRDJtrrQFN8sSubrd143nfs57hPlXlra6KxRjCuoYdor6gSl
V/SGLJf5Ya2aZR5wLve5fIpZzDIQpRRJWztmPWCE/nyk3dMwnzTj2Q5G3el9P4kP
jsQ8NSui0XnI3UjLj3IQTS6uIefql//uYtmvZRYFmxxfzX4/vFEdq4NXROyHYafa
OEWlkCqhRZq4Y9zKFxRwKVgTw1zLLVAsEqvdPzwDBJSp4+ACTVwRpIza4Ty8T4Qz
23A1kfFWBt7alUbeVUYClZPMF67wFuELl9o6XlI/G/DYLv2zo+rrW7Oh8Gr6MvnC
ZFAT687cfCCnUit0l1OmMux7nLGVy45hGCAKrHQ7xt9NnR8OuWRvOD7BKui12IyX
z0BWLJHsteztoWjcfgRR02ZpqqJOesCoWMvQRQHSRthRRtY9KZ9iQDtDLdjuF51d
XE+oqCMl2XR0VjwPecFVCCIqNyEmCzWuD87f7yeu/dNWyF/zXs4lKAGcIOF0zDVz
F0LWGv5ectyLEd6AjPAQEdpV8hYjLX19v995MWP+QNpgGk1EBCwhgxZKgDj27vQ4
cqWkPoMRFbxyU4dWnzc1z+djScJQhpA0B4HfGcD7Ze1h7qaPLGB4T8GwczEAs5RD
21d0OhP9yBbzYu2bEH6XCrTGnofcQOQZR2zBduulH9wFG5fHqPmEdLBdCjNBvv/O
eDjgCPfKMLQyuVpnp+RVvRy/Yq5RwD3Hrow/mFn55De2E0hvaAjH0qHozOOM1ARD
xyoI6m+lcLIMn2UNQywlpRozW/VHNXlrsKrU1bsaOJKDGmxIrDInXNLjN14Epfa5
O+3xcKrU4IhYCLrmoEVYY/pPsl56sX3aGN5Xoz/UNv5sHG8bEuARo7IP6oa89OZx
SWER4rBHdBd2SB4TjCqM4nfyShl1YIBvoD/ZINvddxqG7sWiA87WtjyY+l6WFS2t
TAMMm4Orn5JA/Cf1f6rp0mKzY1qWJxHQ7m96SCRLoiSA5ipXDGQPO4Wzf7Dbc39x
/ONZyGkN7KpQAU7jpavJdxDfcP6HJnPZ3WCN9Zq5bfBr2BYyO05XpUw07BUhPuJZ
EEkOfEKmNvXkgKUnK8/OxgbHzFHkfuoGNXkTFBwAU2/H0nH6bxeEqhAP+J9q7zoG
2oaGedufSM8F8qG8H/QNWDBAZr4EFSWyBo/6K1Jtt2lvg718xVC4B4twPrdI7VhB
1LBr63XvIqtAkVzUVslc+aRHl+1ogKHQBKtwM2MnRiYnbrf+92rmAgXNCTpskjQo
75a0OVpOal9NlC8Zfx0zypXmh+G+xaO5jymFeTNoJ4v1gYfXWqPEa5vpdLRJr3xm
JtxFK9rd9++athwyc57naAJkj6ci/Wd9qbrhSVGQQMGJo5yVwcbR4l46BEHPIbpe
xPXrpe7LnRZikQZGfhkEpwsyBjWoPicbJRAFK0e86JA/4o6eV6OdvOlel2LXXAn1
p3Th6iU0ptAMeMxOms8qv/MILm/N4NJ30Xda7CwqsqSGLS453y/iX555ng9gMQ0v
W+ACbwZQlIyjkhvAP8ySaCbRgoU98oX50h7TGn6+cBEkNlIBbBDytR7J5I8N5yCI
8aPKK6iZEwkI8Pi44CvOivkIwIJ4ksXy7R0UHV+m6dslvy+4XgLRjACf8z8Z2eTP
AhsfaA+B97n5HaUinahIZIsZGsp/v12IAI69W7Iop2NgWMrm2T8hbO5CvY69vERu
lvZIPhIOGG8MGkMmEH65f6osGc69PdsCB2Znz50/hERwV8ENDlcV6/d0K/pntXFf
BcdJNekJ3FvwWMLX3uSmYZpQ0qCOFuoSXLqjfSFmMVGgOReLQAyG+G8MLqVo9LLn
suMv8mO/AXSUxzrxFMhcX52xG8mGSDjYYuVQF/ueT6jpq7cdRM30HEKHK+9SvYjS
BWeWsIA2JZfTGJu3ykjQm8kYgOdUziGq+upNx6vvpYbaswCKdvvCFge7su9LvK+f
BfPUKuyzR/WArlEKggWPJRYvWE1bzWV82odeKK52aocPCUUl706ZThgJlFglx9eZ
2B12RwrQucqN85RbYNNo7G6NMd7H15grFlm6y3O7I9w9Qn/hoT6fp0SljN5wcAoj
U2nD1cF8bnE88LqWohoNwZPpuwG0wPLCwdvvCeV2Dk4y/NSyD7LDd1CwODsyqDec
s06bq1kFYkjdEPKa1cXqHHINCkc8BpIil+h57YRtRWn14txArvauNVuk7n1iuF4G
Mki7HdzZ8Vy99/uYz7VG+UB/TaFlz6C/esFAtF7487hY77Tr9m5dFeE6lh2lxJLj
H9uIQweb/U6tAIzaZCZI2Uh5k5TQmfL3RVPXJ0B90dUErFi6iQSLuJdD6ZcNVJsD
AIIhp3u3uNfXEb4OOIZpMGQo1B/6yFkoiJfAS38jwPoAPjdr0sq9tlE9yLqYgQNI
sIKZpjk8IjMjEDNOS97AN1Gy0lDs0wvqsgTpULI7Pd7OrIO67eYerLQUF4MSH6wy
MCKDnS+TT/TljR4mnMiwEsBRqKcaK7wLAHwg5VBXmjH0/ISoZZB4SfJ15m1CkWyW
9/UqPlr31bm3dukm0edGxUsniqqaXdDx6QJ3LT4h+f2IygNaAzCxh8QfR2iZ6/XN
2tIdkaHbQEoj/pUgWUuEKqh6+6NIZzDBYKlU3jdGRnDErs4vlMsgoXBazIFkDWuP
vYeXz/5XKwbnm86nXea5jMjicbCXdrK/V2MEzwjSXXzjx/4azBbAvHOqWOzZUQSt
FQLjDi0riOwiQwwvh4PE9PO7i+66ghzc/hJb7CI4oD0qGMQjVgVedfsVtqB7byPq
OpjFFXh0oS3sQbrEchfI9EejQUan3em48zBs8QhVa5Mo4nkacL31/QpNKK4nT4Ps
Cm40coZiThpUCrHOwi72kCI4+hbqIrbH1cTysPnJLAOAF3iWrvV7Wnfs+WDDRbNL
CBa6wHGZR4Xb19AzfMY34faWCUt+H3/x7tbtVyg9TNKsC2G7GkNJvgMw7ew1E+RX
vvLRppWYVwqL3TfnxlmaC3wD2v0dvrzlb74I/mqGDIETq7aZSooEWHhkIU2UgrOE
s/bI3/3nc1ZYmyfUTVoq1Q6vBUcEuAz/z2o/ufWmgY1NR6JKbkXZq49wBnTXBMWV
FZojPZKa4NqE6Rzja5Vy92bz1efYI653uNF2VF461Zwlw/YFF7KHQ+5a97CITPKS
+pAxynh3/bKZEx/2ErPFdBRHBV2byrJt/5ZmSit0ld7Tbfic3u3ImpYTtg5sigtq
3FBMnnXzodEBNBdcot7saVdtYVxwMJLG9iXAkndCHEJ3gETsex61QAaNkdmAMGck
Sx1DjRJwHSXAtS04wocU0s5zPlYjKGrVWHOw8p4yPrFt6+poIin+JpjQk7N3XXk4
nnK4JVSJV1oKpuiVMbkl3Tz+Jdt3egAz2ymDaMGJuKkCiQefFHjhMUrG/h62NX+B
WsXBMy034/JIeMGVAeRdrYmwPoutzL1H15umc2g0APbz93V512tA6fAESsFauHfG
V8dYpzuHaSnN5/DbxsDfWkGePidp1L3Fe/1zgfOfVPDwEYA90PVOCYwulV5Sah+l
4PjHY3teoe28EFZDn2kht7Ek3Gx/At7RY62AFvELw9dWLFW346sN++WMcRrtrQGI
X3Esx5agRKrgGdPiJ/76D9mOWkkmuVXaRpXs1Z2SdkiWHvvVQPB65B/UCBzj0lPs
FZQ4I+Nv/XID1aJiEl/hlf6eDpeE5gn/dryV/TWGkvGFxrUFaEXqVFSKY23L+aoD
Ssco9Hbt/yh5+IQQ6jXVxdSMSXbuPZ5XZvmmO9yBgaPSFOczOyMLPEfefIF5ivVr
BNiAGfyzsAe9mvbJZIMzAsTnlnqYcS6mSmE/ZaPXrhykvPCnb7Zkse23EQakuFpA
yuNtq+aZNphu846O00sAL/MDe0gyshTLqXS9RUA1k6iFY82zMIMa3jJn6sIbTYhU
+TQYFm1p+TydKW7QdgWeDiR/sfbvA34dOXEvJ48O1xtxRhzhn8HPq9cpcM8YsPIG
jieacMz6xmLE+7Kt+RZmjva6yTsSKHMfU5MBQPv5xgbfS4KyoVoUJsaJZzwVqpYS
v1NvdL8yfsP1za7HiAFds9xvxPlXAQAZHIDL6VhVVT8nvpu7a4BHNCB9kt9AQ+Vg
JBgquDbvSdTbnXAdLxduihLWNKT885zvmWoHGDkY4cCh02o2xmq7KMfCiR9t4XWc
N5flGxJrxzfGF1WzKI0ZgRmrzX+jHDNC0LRRHhs5CecTJQOGRaT/A+mW3q6Svl9j
3qrO+qbrwjBAps2OE1S47FDuerNsZO7pralaY3X5dYmqaYfUjajbjXKGA+/lYF5a
bRiE0zNFe7B4nE3UpUcjE9FG4oa24Jcq5p+Nx5KL34wq5y4rx2VDnin2xRgoMl+9
oDPgJYzzF7irNV/RagwOa6Up0VvHUthdUa40wxPW7kKcojqqRrnLpWkQmEAcP7dv
nzJm99IOhHCRW+3AiPt+qUHN6DbtWVZUiVQVfOq88VsGczvDCzp8Rlv+A9wlu1A9
qsX1g7EViR4OEroagBVYnH7+L/ANweO9SRtM6uFA1XLk6b3GKA9f3JDeiHEKa2FL
sCIdgXerSqsXwQiZm+fBMgq//a3DO8vPEi5fmJqEd6vyUtDrI0OU+uh2keeR8Vry
DJ1HkkmsuvqnVJ7WqBWZ30gqTKIw9m+7tZrwRbntmlGTedcPD09ia5rrj7hYnMO1
YMB+eCuQ+9gS2ruNob8T3JMIX99MGeAkI2/aAd/XPv0TL4TVXkbD2rG3bcpPRp7T
bEqDnumMid7R+hYrgA9Hh5m+7ISbAOwT9ZAVgf1dg9p0ZD4F2hcdidwNO8T7KF46
Ep1ZDxvfZnwJyoez/CHcWz99P6lDYuMwSuRkTP4H19L89ZEJOLUlcFTYVlM54Lyh
pZgn7zxRznfWjs/5Z7wRsWqo4cYTqwZOVYZYiNkEOhoX2xhyaO7cn3js5PaWTMs1
+kSb94yv445+fqpCzds0rniQrNqHjs+jHSZ1aXKFFRaksOGmmlnthT2vRNZta6H/
uh/CaD8ZKalUQy4CstxrajVIy+7CPq53VEJPEV29R9Y7o3986PCv9su+EkD8d6NH
wv63i6ewilIjukRFsjhgvgZjs8M3EkKTvzze8xRexg2xSvzjqSrKxI8USQq/ibf9
ovZJO6x3mfEH/ErhyuqAAmsdwzQPLiW6SE8zASws2ucO9Bu4+/wFm32VB5hdGob3
NnhSXDeZJoomyvNc7+yEvxEi59/Ie6ipjTVsuT15Sx9WY2kHASIEYwYhf59piZXy
N8D9indY93ALIpPvXO7hlE1mepAaAsDtIXKVxmG1b9bHeHTMHQ6Aucq0NBL6l0/h
EhYkPV4RxMNpe3nPcHbFdCt2LSMCOS69dBLL5vYfLALO23h+ZJgcNrPkBga9w90J
JAzY70fdK+lY0Ds9EkETLLZnn0jD/n3JmuO9ygM3jpNtNw4q021+vvc1MI/qooQV
YT1w32huv2e+S+QeHeixW66ZR5cAWBGpDp6nK33VQN9ZqZJvlG/BG4wKctbRZwQ4
bYSt6Ovzxsz6RRbJjkpdDh5Leybq9idLieeUmYdOIdwjvmmt5tksvyGHzQFnLSR5
756rs8d7pbVDPnO+qmV1bjm9DHM518zs+JAqPJElfhyxlyoMA8yLzqBuHUOU3ZpM
lUFD6eVkiZeDl0donBIbgSoD9sw7g2zOm9nY/wzpDIJWAeWfGXfx/oySdP8SgBSu
zp9JYzg0+S6b9ZlAV6nXEs8rXctlV+Ga2Fms69MR7/OBxWOnTKp7x2B9uxoy9UGq
sFtDffegO+GSBxvDpryJ39r1saPjCtt2gNyRrNEXPl261UAoY3ztgn/YwKcMPapl
p0N98zW4U4HV1Tj7AD0XVXDdcyyWnWNWdODBthQ+2obdT52gYMeoLzrLAjUkb59E
zE3pJk11seKWDqZAY29DE2stLasNz/VMSodho2lQqONPhfBfiWstb70MCHJjdGG1
kSCwQf1MVY5hGg0tCL1eeavc5ZGZR9quBggBhUP9joP8YJf7jTpohegrusOY6zgF
7oTZHLiuR1rSObyxliljF1aO25S3s8M9m2Cl464PY6R4GtjILg+fFpJUTH1y8Zkp
MGU6kV0bKDfkXv64Ups+mP98C9aj4Jgbzl+tew0yK97pqP6fwPEIa/A7sSMf7vfo
upUDCE4EqTXuJ6BYpTfKCK/ElK4oGZbhYnltAz6xJhwbcgyMHYoZzXBYchLpd1o+
MsoXJn0qgX47fPMeQrvSYDnV9JIKAX8kf52Rv1hAE3TcXeN7QEj+DqH51deDt9lT
c6J2Q8iGN4AHj5oUHnRldV9jEzQxCOUAy9BlmJFOIpOPGksQjL21R332xeZGSIf7
zWkrqB/gUraOI4tQDdsMHo4sLLdhCE82rQA9IgZg1ntIY5Ep5VF8L0fbz9MOYrri
W2WSXguQxQfq1qbgWSj60V7vqh3+rerLgtYWcByEFh3yGbe7WVaWrvBxd9gH4xM6
v0mFKP2QlL6grpUEIEBDif1UpLmMGn3IWbHr7K3LHjfgE1S0wHwTQwb5zYZ74o/N
++5D9YA6iNqWfEhgzLJhx3ig+h6KMWY1fPUJliqL2xpNJVRs/r/pAaQ1tKanmDNQ
qi4HsAbiNh6SDMzA2Dh4Hk4dF1bPr47/y3ofEXoZKLT1n7AyjxPmEp3LfN3ImnwA
e6VfQX+zJl8EvcizFEDRxG6UFiSAcIrJUKVYdFMNaDuUM0XIgVeo6LMwslpbebHj
tsvRRGmu0gIjVjuANuQDZGCI+kkwZ5sbUuLQN/ySCeznQoGHDj5PkNWdBLUavs+0
090sdD7ku/J0HM5wYImGGq7Wf58cAo3Ts04qQKfl0wVC6HCkFYNySfTJWJ7cnnyl
nwrPNGKf9YqDe+ORadkFQgVhYWtOwEni5f5RqhseQBFPQ31nYiC/3ycUHZLBNOM7
tdkWUXeFlpB8eimAACuir6NC8iul+HdiaLhsrvZ8MqrusoZObiXbRhQEDKw0jxdK
PcV0sh4zEol5r/cwPGZ6DrI4tubI9a0/zp34Nb6r5KhhQyQaj+TKMn8oZOEbHKU2
emSvOdp9gR+RXTP/CJsNfIDS1CI97ZpDwaBz/QOgByFZhkTa+HAPdxvbwwiPPrWr
I5c+Ug2XplVWD7ayjbiDTP9f9xSoeWtCPNV3tNBqE6KPQtx7LqVGG6D094Ll0pJY
F73DE6jQOSEJbtIpyRHeryr6fjelPtdFT54QXEa3bXT7XzRYKvwWd7hzLLt7k2Eg
pcYqwrpvX7KlTr5n5hevxyGMfqgbzcHGvguJV3fyOLZi5EffwD2Lpt53n3yXIlTm
U67Y6y2w5jAnIXMmHL/dPd7trwohUo+N82/2xmY308VjCf1fyM9JRoDaRS9TIO4P
a12+RG1PZZUdqlMntGVJqFZhP7oG3k7LCRXQQ4X6HQu8IafjK/5uIh9mKp0Qs1aD
3gGWxJZxQEnoa6YG1kBCEJFerCjy/MOsThsA6VKeNfisDUfMLFhr8W9CynLiyBrB
1TzsU7g+sxOF+i7uwJVOuqthz/t/w95GqXGMeC5qXbrlNddiqPwYZlBGkP6n8Dil
y+hc9lTLisb1EEtE3bLdlFYq2H5poCwAYB4P1kCErl7D3gFCz0v+KUh08T7b1VoX
LK9W9kRecl+BtrmV46UfL5QkE4lg9moSshbkMlOq9JE1aLB11pQqXO1LBcA3kpVN
4qldljYUc8RX6pAjxm4H9oKpPpzNu/qjf/W4GfwGWQ5MowOtTHnfC/icI/6O1JKV
Qs7QY06RVOEzodXlZwcgV9bZ4ElVPdz/WO+/1o+B4BV77cAjepSGWXpw259CDiWy
470E+87Z8Gd/s46XKWgxyOoBUKUUNONh3ADNfRGp4Mtmq1ZKZSRrloWU5w3ieUpL
yB4O8NEqlLsMHioa0udnrg6e+a0rJ0CGfu8R8KSnLWAd0ql8T32L41EmJYHUanhv
n6NbuhotyWryq9jjPKSzRFdVH5jRYRYFdbHL05gsyCD3LmGZgPIsGzgwiPyTnKi4
CjclwH7LGqstXEPENUlo73Z9Y/agrXJ2j2kQJsPuFPjwztk+Zz79P7RTHlWkRm+L
fJVsyWM3oL27w34u7MYtNL3/CbtjVszUx45mJ6e7vhjAalLXHoWGQPl4yPZvRFeS
R7Gl51APrw2rnp9W3Ar6e36WNiODR1OCCRUnCYqnyiXGWfySrI8XrPBRnlhm4AlU
784OPt89KgqbKU4NGtk06SaYzvIfrPNkizOpaZDZ7dfDfhC2wYNYxqUCv6ddWgdd
iyztQeP+qpHnfnMketOB0k/o6SrT6JjeFlrEltn8S+VZWUH6s5adv57R1wakXRc0
3aiOx5yOUrzY6w0hbKJtxvm8y8HR9O5zlkEdZb65N6AU/13AIzO/exyMgXUZ8+C9
OP1HgKqpcD7C8RW8Y0lFldCeDKschbmcRXaI+D89e7uFTEvWI58Eu/QZxZY1I2DV
JcPd0uq11Yq8DzcyJvky3b34e4HHwQ5L5N3104LmXEUkFVH1UOmK9K926xIlpl1Z
7CT6sN+QViscUPElbDp8pQCJetgXJzNEKhuSKI5PpgAHnznmkdCNwXFIjmtjKxDk
b1fnzErCTLkQPudnXNQpVPokanrS6yN3JaFvrs31lLvpH9imfPxFsl5PWlGWmYHV
230ollLWRZpVsplb5d1oAwetZZ2UMwG8QgiXAzr2KfwtQZR0/KkqjZHNmzCqEfdb
rxzPMQFdPE+RDZKk/Nad5lP+/tuadtxaCHAoF8Fl4SSRl0yz7zrdaXi16MZyCuDp
kguWu0Go1WQFoibAh9s/raeMpgvY8Zfsn0o0quosyTV0Yr8wOhOftdrzv3TF5QH/
lcjkygvYPZb8WEyGm06DAUR8GHsxDgrx2V6rF5Xa783gq/tvQoSK7SzVic9UO/7f
dgaboIJqTPi43VnQ1B890vZia0Q8IaoLIadKuYgU33ivzMi8i/YRDpt+Sju2C9uz
0zniDBRGAxewgVkLnlXNDyDuhuBbGzmhoenYdsBgovgXM5zpBdN1t/GGNjmrMw2h
h0b3oJ+SSa0A4/FvuMeleIt2y/LcajS4P/eWb7O0Hgbhee3FtPg9rX/0fNkaE3kU
fsUT0ERBTUXEZ2ejW6RujGkFcOPoDcY63SBwQZ3J/ffqV0srVclnPm2q/hQspQG3
tQn9dwszc+K+0YhNRLiZw64rwzFPIA8xK6MIJoXB81WdZP7PZHP7GMGRPiPMkdyj
VAfwqGJJxSASXt/+/zG9hGAQlLsHZXNAkdxkH1mmML/7xLtycUPXgpjmypavRJGJ
SUibx1072vIPP6A9XrbqtiAObXR9DsUTXUFTini0YsBc38m9JpK6D1OVAh6iJp7Z
1XOIyv4iHk9W7KF/AkD4QUevtDSrCZ6fWDIvNbEf4+80xBwiPKovDOWbJyMxmiOs
2u8HUdD8SLzIpu/3FSfKC6MMb6CYHnL0eNRNuMlRt76Co60A+cijXbiB5uKktnQG
yqCB3tjlqzM1mQrx5AdVjcRGV582zfP1WKWEyuCuwSaw9gP+gMtAIFImDijVhaIr
HOvW5vKSab2GE2nqhncZxQNhaYiXSzGNt5A6vV+ygXV15yl0XS38/bCGTJ3yV0NT
SKwamHIlyuRkzlTGe2k4K+IY7hVjvnmDCihu77wK6DYEZt3ekfoPjFCQluXw6Pcg
C3SuWlzRh0DGva8B5tp78u4XMrGEXS/xlY5vAbTkL8k1Dhe37zHTCQL40jOP4vA3
FF+mk0MQVKe80l6wjn0RGmuRX8WnWFLYjQX4MnqrYZNykAhy/a1TIn5wWvi5oN+E
QKkPZ6zxGw/KT/EkHHohvyiIFUMJVhCdHq7PQ+loAcLYxjOACmtZjimPyh7AjuEW
dZ+ySRacfMVZD0jnDSf7wh2/EDHd65P5A5w9kcU51rxrXTCs3bPNwMWCKjRwqUMN
XU0VfaBfGKyzsPybZy92upCltp8EhiOAPqbQmbAAZ3EUZUfTvr9zcOplbkhWT+j6
hKIJ//MFFdQeQ5apMf9YG4+p2tX5FfAxeCQzxORdrMowkrnG1GYddwC3b+yyPDXw
wCGS9s6cVQbZAGPkVY6DuO7gwM66jZGjUqtfL7HKEHIyXuncBaBZlyUrI7L99h+t
Moeah5Axr6irVFFTA98NFd0cTXVHZFJtdmpUQVT3VUErcU2x5etVkFc745TFR62L
oajFrJyUNCLEcHREULGYo1Ewk5oU3Qfz9+JsKVpXocSr97fijudkW33/HXuCQFSo
Bh3CUVyp6ONmPoWg9aYz6L1RJgSwmn1pD+2hYG0CSuYdOzj1ZZ7f/gpfvrCk5Wpw
OJXci9ebzYddI0orjHW2rch/cxHn6bfERhfpBrvMAyC3QhKATsypIRiMaFtNt22V
8GsqRhH46+ks0sSe58cCuNuMxJL0cB7ViwodM4JFrwmu/+B9vVllSF6q49QrTwp5
sj+OH+4TDu/YRWEhSl1XpZY82uXjtH6z/wxHzwRfO6AA5rca2SEPqF7kn2fMmbgF
zrOwyQ1FaCw8u7oH0GoX01xvDq15ZZ2PgAcwnfLwhAVxzFINKoJ2xVCjyOGwIMoG
uz0ZXapIUx4QGyt76CWZvJ/G3LIJLp1/xbt6QxCs+pRTfkKxNlK+ydUFrRjtwp6z
cVb7JY9gRLhrUzn4sOBPTbUq1psccO8KKNXgSc4XHYxobzY+bxWTRVgXAyHWAuup
c/mvNViNOLBo2RtDMsvcu/RaWmqEWHsuVDK7plauESMXBEBMbjM/bYrmXM7TJXDk
jXj7Cz4mYf5Tea6kE3ZtokhnHxxEIQQElku+iH8d3PaTIexRPaSqpBt1MGfPo3PS
IZctQ3GsHT078wxks49YNNg+tivUxawirMg3KYq7DGrKdDVXXiBBChBKAK3Iy86E
o5GcUVx5B61D5vagvtVwZP4B+NR/cifJ0O5nsYdj6osX04caVZ+Loqm+Q+QmjsB4
po7wuiCI8cOsca0eF7z+QVCSR3ulkjTroTiwthZmIQcdVdvN5Hi+DLS/D2a7q+/t
BORTd/VhFz7KQY3OPM5J7LmGFMwn2AQCujsD8HlJxGqmLDMX/6Jg2vRg7aMERbj/
2Pzh+F1q+aopUjHJAeVou5bUeIaCwW7P7x5LiRrf2AF05M1Yh9PgE6bdDHpI0+ZG
IVJuU2/zIb4GKWoCSaw2UxpVbMrSCR9Z2hLlhxBcgFRPsk6SpEMwRqoZDz/MuUKA
q/UfxAVwV1VeHl3NEn9Ba0mVCgZrEVGWT6tWUpUDJLPQtDWG179qgiQQA5MJQR/j
u/Zj1tIYqTfFMYT8q5zC3xOG2H2MhgpZVp59dXwAMXpHiaPP2yvyPZooXnanQ5qC
UzNxIe7ChIDUhEkDxmmDPk+sIiKXK8ayM2YaAqyVBr63NuORadg6NyLHHm2KMbFe
nNoiwXhrCYW5+VLZsa+r2Y+IL4yOtvsQbTHIfTUMpw9x5bh1tisEB0NlIxWF8G7M
N9xty47lSaND0cjaJTCnpItXtZhRX9K0ydMmTdLcn5L4MxJz+pNVr75nzZHu7fYL
K6EEbMc3sHjk/HEaw1NgMANSwHT+vJgygiw4XVKajizbMkqZ6eIAcyYvtgvuWNWn
CTzZ1YFCF5fOBZJT6Xuyk7J8YxsitYA5mjS3pkDkmkMfJViBtXXFr8sXsi6BEncx
sxDPFiDHQ8VLKqVV6A2XupNzZPXL00LvMMSd6B3vsHkAlSqrpC2PcaOLgpyvALhz
OSL++gbhDHsJ0dLDeUrgJfRcDJ1HO2GQiOvr4+Ruu0upM9eCXLzxzDnnZlfmodBQ
Ls9ZUY/gkZFJn5fz7uFW/EOYGzCac6Tqj5zP5Knd+yswWuGBRF2tNkSdrfghYjnX
lduyjh2Wj//FaWP78WE9PE2XnQ8WNYikySSHieOxIW+JsqxIvelgvCYnmLSqV+oB
CkkfHMm4uDydm1yaXBiV/J6Umm6d8yaxw0pUMb/N6z6SsZDbuPREekXhmOHUIIs3
W4MF0+lp4U4KyzTvE7eYflUiG2MwXLRxindZ7dphsd/i7VQ5eMKxmRyFytYrKF+V
3wGTCWWPKz136MvJIgBTSt4PH9g1imnSeif3w66VJgEFHlcNWUJ3HaEgyZcdG+Su
8ncUW2v/oS/xNoq73VvUrB4SFctjcWDQvbQLb9Bjs/Tk3BfAt3vsABFV1JdX5QRg
M9UMzTrMjTzjUiPOLyqpAOO3sTPcTArrU3TQoVZviR6yxNU2Nk3lfefGz43Pqqir
+/+/wpNhiLw5/LnMTenr/vMJ2odu/p9F4qy50fFE1vaTliiMZi4aYlhOTN6jrzYT
lGHqIlnTMbkdLSw6ECbHKkLtHxb59uOEcYwy94ajM/LzWDFCwInPfXmrsyM+CT/r
IXcAqnSAj/B/DeETOAo9vLwhbe3vPHw/yKR61pecaaMrw3qLrGg/mdwUCNwo/Sfi
NgOUl4UqGqkEUEp22wrEzkULjdusYNFacBlKxOH/lgtfGSbcwJxUflQ03/6jjF4F
9h8k8agZVDPVxNKu+kJDhcMM3gCaS15xq82bzixavKgF1Q864C8KbJHn0Qa9kc4K
tfhDOAY/hTjNIs5DGOLESwj3k3zvDdRtT362k73ulWDIA7RwXy55lcrkavFBUWb7
d5qTEYG4DAJHeNpR95uUVAUGU9JMOazml1Ol10q+BA7O+dwWmyrUNn/1JcdFKa4f
hjyxFeatggGcsT+dA6Hw6vIgW4msdCpyWy9kgY4wBgTOV+pDNqEnG11KYE55vK9H
t4niKylJQQxJK54C5rNJcB1GYvl1hmnje60cYuznoHnhC0nbPQfuPWbPWvelbFax
AZ0x/vYCsesFJgFWJm0KGpt+Fie/xn719iIc1txsd89ekX2s7YLY4QfvVBoS6L68
m2zteAA7FkXFWrvdYDJ8KlT99VHdnAlE9UQpcjqGn85VtZadUBK1dvH44O8BM56p
VabW8yXleDNlNtF3ePFkXBOVX1ymaBNZ9TKvSFZbxah0CWKfS51K6WgGGdt1xDhR
0M2eRKSjHJCMurerQkR79vHUk25kevB2m1y5hyfzLeJX5aLPEFnKZh5GpD/BT4pc
uYyf1xj3uOdojezRaWDE3h7qqV5IRr6xdHaxAWKHnKEbDwW2p/vwhJPUERtKlNS4
LNaSeoRZuqk40Atqu+m35M7VtdX5fxBpNjPWCzUbX9Rtrg2Pi1XLMieLHKv/+lGO
GPKzT3GLO1NLjHYkZ29hnUdV4nBebhf6hVnmspZfZZ/hmbgV+wir6LxPqahRw8up
Eer+ggcfnTPZSSnF1LJGoHIp9Z/cumlt/Cm0pTCxWw5Wzk7iXq1TUAKiyVFjLSdL
jQvJRN8+T4u3EmwiAe9B71EwjrZ1iRN4xfUZchs9c1Fxt2Ov1nNYTSdLKcuAYnnS
zbCP0RSYku+1ksoInuQyTy01F0F3vDS+DQqBMtaoMd6iX4BhWkiyvGRIxSTuOegK
2P6FVzfFjCB0lZMga7Da4djZam3VYrhpqEP7i3+pNqCtLOPnQ+eHkD3EsincN6vD
veCD431/jrLN3bZdw6zUdpOjaK3iwbMqBH8Fgt+NbrcgdkESk7RmEZS5aLhwnbku
zyaMmhKUwbRCh3HsGNAucCODp/HBB88aJ6K/WH0rmq8ZSyf4/bgwQqrSofzxNfoA
NFAzciQ9rWTFjMiHGPAG6LpXc3S/RydbagN7yrAm3EIOMy0NzsYyyX8FNoCEKvE5
0D8qLDa3kL+xjmnty8vjQU35vDJAkKmkmnrRub5UljfBoPMnADxQe8jO/SS+ab5g
Y/W/FYZyT2LlIeht+DhaDHWivlAHUDVrmfQaEe/e1APfSpcSeKQHNabiAXk0TqMN
4ekEukXNZiNJfOgjVhxdlmecvmGEBB50wPZhiNyyFJoX26JUalPmsryc0bvFfI2+
IAfwuuUk6BFOQ/crC3kiFwueb+F8gUh1T5dM8Gs2Aw+tW4h+1nWTrDfH4XrI8ExH
G8Yw7wqmB7/Vd5RU9E1NdJPBAuw4TFEurlZFuS1fuP8nWfEOKOvs28+t+AMN0SlE
RYLOEcZ9TwUvJFMMa1KuB6iQ4ITHyr7/uJGAmY1OypY2EKIo3Pi/cIEkVyYTUZ+y
mMkuK+N8o3gp5vMRWsINg/sCXAemdaM5qzPwwCONLp4ByYm4EGJrq9dLugI9XZOD
+W3qvypvsPoufE41n5K++TzXmusBWMCPdTRJ9+r9y7JlBAwKPKqIcJmY7j7/vvQQ
8WufQPLJoyfiIfIQW8W1F4JV8DQPuuoqYHpfJ/btdX2mrYrwvLtU4TXtn05jPldq
XCE3ULWTqBx58KtDKTigolFnbn4wmZL8FPP8MU3Fbw8dXfeEmobMX04vBerm5Iyi
r1ujO1NcV3NxMnRp35gh9Ld2hojMSbGsRPriqbGG5fdyyFjOUso2QZ68gUcmFQt4
Q4YBLEdmzlAk0QcnH8nsKxjgz/fN3IrJX33pYc2o1XqxgCFqICf7uJp5QQ2ZtOCI
8vyGwYaCkAy4MVJ4+x2hIFbQnCiTARitmsLFBTe8vLchzN6QqyVx8NpEAQ0yhU26
ood4sEaFfGWs4P+ochSZgZqsNF7mZKkiYRCodmtQ9uT7WuNOIy/fD88XYMiFJIPD
cuAN/qN6rQQP7RuYtOG3gvbzjVX007KSS4wJgz524UiNDqbtw/XIn3dya5lClNXG
q9iha46lQJzXybecUPt9+Q0TC/BqrHG8brYOiaQ4t/Zc22+dK7aV3NuXtFGrEfBk
JlhqruZz019Oz8Fi0BDpbPHHkaahF2TG6zPWvqx7WfybBW8R57CpVCzN34wLF54m
phIpmC8tSita8zjuaPrF46G0TSzyyHKcfZuB7yBerN4YP9iDuwk1oe8J+fhf0yej
GZ0LoeY5g3AnXemDg7MfRnFTZM3hciHWrqbr0KpoUU1651J/Z6JreOFzEka6e2pl
xkR9fkdDaUDJYHPLN2Ki4yQUHAnzTV9QNqpzpwEMIoQVsu8Cj2jtrPoYT5IQicYj
cMs7eGaPjjqmA037HDoh/RhIyIRHffC4sEQy4akqpnxnUacTnPKUJOqgcBoVZUp6
zZ7BvUsrnU46FbwTMhT+nc9VBMxZILQOGyIqGXW9LuNF13DTUShW908qUQDxgi71
IyKn63q7lkhJx7qmZ3oDAdwe9tMRRgaDEuRof/f+uis3WTwiXJasx4R51jZxuYJi
p3ynb8KSH0lzucGGTRvbBF0FiJkL/b0n7ENsk5SsqCzCWZU70+33XURFyeBC7YLz
YuJwqrGEZ4wkXiMjOZIoHW4gGfn2oDMYAXBHMUSU8BfqB1XcSxx+ZBRjGh05+VUz
sKdMs6jh5lnvSAImnSXDx5IyGNWWu4feQLy/gnBUn73K4pht0N82/DRSdQ+tjyL0
fdoDm0atFj4z8Gt2n8br60Oh1ELaMVmTWjuipWmveRqdp3xuwhcibiYA8byme4Dh
8DAn0ACUfKxzYvhcq6cEkbUlEfz1YQoDSAXO6gIv1O2TpboAFesFmCjbVNK35CXY
++ds+k89NL2N4EhqO8D8OZQQ57+s69u5FaFDLVUiLS0jjjQ4e06IXS9nhLPmXo3K
zdZmDbJJIwDTPEyy8C0pRXvuEIqvO0qvwBd9uv9Oz3wNB1uLgeUPyxZkrLiYhimT
ONv4qNuT1lfmWGlurii2vyLYpvP+1vjLTAJ00ubpCFLdV3slNYiMz3yBZ5VLd1t0
HCAC808FbLzWrtbCaRP2mmjTQyHpPgOXxO3y9z9S+/Llu18Vj6TTpfhtp9xCN9nC
ySxF8uQtLIJQjugDJPncKW2Fh4F/DSLt0FhMMJIdqLHNZKBC4FJRIzxYpaGozUf4
5Kj/Vq7ypGomAnUI2uhkuLN3fWtf3RqaQGwmFprtahTBhasqBLZ9iB99HjyLNl8O
4fX+DSesZXsQICE86KJSguA4z4pOPRsVubXTyobcZxQsmZ+UuKv268c3VQiEyeqS
iDxEzsHkgR38R0EnACfLw/f3nkglUuIHYXj5uN7Z6YPOlNY2kBZ0AbkzjQUbGMTy
tgDCyCTaeIn+2W5GD/8nrwvRySdeLpp48RDHzKRUvNuuyAIvEIRY6DSCLz3Am0e+
nyOakdh1P5DXNNLouNBhhuSvSNMLWoUbgrg2NyUtlzquxY7DJ6OScbAU7nqdSjAg
0zccTwxaC6LzmpCeCxL+8GaSmGAz10ttHDUcdia95qDaMcT1M6p7JjWhXbQm9694
FcueAsN+MiojIxo8CIAzG3ZtNHvUVzFznKEYGJlGI33QQTEHgp4H85W6xL0reBW3
IlrYqmFTZyA4PfHcVe7jqRdwQg9MhKNwFrgCpaJsrIkEK92+JwqzgIHa1C+RrYlU
3xfLldIITXjF6EnIGd6Pwwf1AFe5Nmipn3U8mEtkR/27RCqTU+dHtXnQB1A84S/w
QONXx6Zcj7sPx8urO9zFvsXSiFqX7olPB/Z72pREC5OJWU4esDW0wF0cq3JHpQad
iyB6T4kCjS8x5X+zQsV6235liwo1eX4bQ/BiVGuiMazJZxRqy3DOjVb8ZPB7ww5R
HjdYeKTIPQNCPRfdy2hXS5uJOz9A7ous1c/q/53Q8chUVcEt5qhD4ZWPHaHWaMwk
5LiYQ3ohXphdNYW0yHGfnBHHHAsSgBNfd1oQwfyt80ANFPjqimgh0NZ4jB3su7eZ
YQFxMVZ768HAzw9bIHjrVJj4EW3eOtNt0uafPhWdtymCKp2T6xU0iXMC/fa8izVE
VVs0n69h7ks6iLL7HrgamcmKhBVv7kGov+GsoUiL0/sYm/Hwa4j2F52NhBRJLpvr
bD5Rfnxsg4PaEIyA8qSqAhpcJ7kZvsmNJoU6nKJ29qGoUHygM63Fu8W61idtioqP
6RJfvMu1phm4TAc36ufFh2FiLnt68py5b8cFF3G8CDsSh4JYwW9UObiHd2Ev1lbU
L6rZCE3hpWolpkK+xjJg8dbAiHG+4p+wtUOy1BBoijUCW0z4+g+ltpBvL1nx66Kg
vO1Sw8P2GW4uj5iG7lphdJLxECxkJeNkSDuXmuRpJA0J8Cje7DtnIos3IOwG32Bp
idD5J3vZQ1UsWFXFKr0GWNnhLvI2Ip4Be1LFDkUNVIjbcDBcJYhyq8OL1WC33xhB
Cfn6nk7/7k94GEqJQGOWgTTUf44rEWZx4mP2euMsuU3sk4FmyxK7qB+S2j93iYQ5
D15b8ze8OE1CEOSt0nzSB9WjIcAqaLorm1GLs+V7Gox90vfhpz+G6lmVYlspaEtp
PxkEJfowdzKj2XOK1ShqyzvHEe2X5hAbhnVLGeeDC/fWIfI5pL/qog1OIYuTIywO
z7BXZdlZC6xnHzWhPKtrh7vfu3nqZTUvnZiTJx42EdLF+ZWOO4G5bpA81nFPxjQA
7bFl80wb3Oxyl5Vqqq0n3q3O56nH9xf0wR1A0KktgMHQwEIAp4hHqNBvD3IrDQ7U
eifMg2X1glQzVTogiR43VOPEjI7Pv6/dCrRhMFERLYjGJQvYfIGHWFIPutKDl7sP
+Z9Gpr3FcWcF6Avl3hSxr1LoqiUbCMMtIokXXEw90XvocPnm6NF73Ttyfw4b4M1m
NHPY/fmvZ8h5/B73Y/ie+2zboh6q/s89AFjisZ/FjI90hJzIxr5rP5IKGQ8BZ+8p
NTZ5gMDyhRrgwh0GnWgVtd+GBNF4X2Fb4B+lPFf57O7lCzMWVTHAjvRTyW+DsVdb
YFElBboH8F58l9vaQyfiMuOf5JT1jufIlz4O1BSX48+gS8VdkPAfbgRLlUHWdHkq
g1nEMSR6VyQenJfZ2Tu7n90GpFAUbCSOzfuZlL9bLG+RCGok2wgV6seMIQMYCDug
dF3l4eIVfTmrwFFF0VZLrQWkp+rp/npL2W8RiLoKt4RJrnJU/Ofc0PkQXhJ7ytlw
gtZSGgaIIOa2jOODU8N07vy58lQTmCjcyaNI60JejZ2ZDlq1keQ5fnisLwwUckww
/10Q6ojzoXjVP8OtvKHNaE+wIBw5SCs6yq5mXCOZiV1Aw9lYDzMqyptSdP2i5gKt
yWyQqmrpL3nJVSW2zmE8Qgi09fI+quFSmwOHpIEufV0S4iWkv4H6SWS/doysU6IT
fSF6ucpPEORvIDPONgqd3qYAJau6nD0hUsbypYrnT73Kg2uCYFMMkkJkCmD0aPuE
BrA1L4cqYkeSq2LXJvFOvVoiKVpU506hRR4P1ux3VdPt0mBiFRdSL4wxqkJPBuxH
54I3m44mKHmXNaX5EoA3n1rWbix/6kgcM+iaBkJKoriU6zUNfiQALtKP8uhBWqxV
u8gC0yxilco8Ff8UbD96kCx9w8irV+JbWcZyvVfb/s/Az1yK8Y9rguztgxH97iFZ
eUCIpG5QTzqVDK04booB5SUg0AXkwttpHHoXERIZXPu5+37e/rndGafVrYmEBXz0
O+OoA6xIziPdegSuAyAU93jAjGjtsWlsz0q2/8+J7hD5ucPn1OsLTof+QR9PNIps
Xn/Gyub1A29aD2lyySiBn85qPprgdK3qbVUhJl+YoXaOJnu14ORUYEvOcCVp8633
iBowmwyukmeeGS4Vy2w4wgM/Ifs5UywfXknQdtsHNGCWT4vFdXiQMkbu/pBKr5z8
B/SP38hr3VG7+X8zd3b3nqIP0WUrXGf6j94HHwEdsW9t34BJdaCi8DirZ9hEg+17
yrnang6za26QfFC95vkTBsHwc2cFmTMCk83HnZEahEvLSqnX/jdqDuD35akFjXz/
QOnpiAPXBWGF254Qz9l90EHkeywRlsjNK0a5PDI/HggbvLu33SPRmigX0KokrX5U
Sh7n77v2KB6M/2JVCg9TB9fUu5mCWU4sH9DUgZDRUIFyIPQE3azvQHp2c+vX6LUi
ht11si5yfYBkyIEfahepzAkzG1+xgiDHSH6eFluY/80ELePic5bvpFiXMoRsxVG4
84oFlIEv5Sr7k5dKMfaOBGOu/pwLwfxgciWNDP6asz/L21tLRGNJVBxuiQYVhw0N
H/C53gKpgeqYAATRhDqjY+N8v7q0KhkPZ6Gs1DFrWjX7kxv9Dn4YqvKix3fp0V4V
RBoOVgiUc3hZXMTTA5cRkcPdjRKQXgP9j6m82rWJTUVIxbDeOpwkmE5Z1ZoTegfx
TGPIcGlp7wqZQRM/7amLZJ6xCUFQLMl/IhcspYsT9PN6RrZ2bnPorR8VDh5KC9X4
RIBIsIEx2hnHmw/lrhEmNGSa+WjJbYNUN56eSnYhLpjiEs1l/RfLs9lkHiK8eRKt
r6CoNOats/DA/NZxuPoI1ogFBJUmsHr9PE4htAkugxAeljVgarpKFhUMGD5Acvkj
pP7qxhVvuEDMoUgHT6J016qom2fJIVHCo1OJftYzYUDpRyTUzv+EEnrSx5HOyai0
0Vzx6qpbT9jXCP1vtLvyvFLdK8aIZ9InPZM+MQaaX973yFqddBoULsbxcojSuo9M
n940+3+y62OGHOxVPuY30ti8a1BqI/FPVNhiZb+1vomiS2O6YedcsQKXv3VWC1FE
8U1/fM3r+sQh2KcyJ17NbE7ydyfiQE0w01nLtTc83mOTWRMMgIUnm/88pLejWjGP
XaZKryvRVrCrBrzcJ+uCffL+Q3cHD8QhypbKWxZ+/nVLeaw5NaTgPjEeOg44cJZl
VkVP8iOnS7DVQmfAl+QdPSRy9TumFQx4+Bu7cGo1RbhF5cH2XLChmlk9Z5Qn0qg4
NGsqDjLDqbXySD/AWdXnMTDtbX8PV6ARo/ZzhNUA5lzF9PI2PU2ECOXWnCoUv9px
0boBXsgR+PTxqJzx71TrLxHREw1KIF7hBVofCqE+sPeqYciCuXrweh0J4ly8ZkpR
A0C7bKyscgZ2cgzdXdkboj995FjzzKt5S0ytUfyJWjdkxf7WuIB9pmd9NwgcLpy8
SznmscuwSt4ODLqyucS/MOdbxM3303/aB+LGwt7FXtOB+JJMKCFgKo0uoVZUwNmk
TxdTg1Cmam+126iP5cnBUwXVDWJDr7DBZ0U/ymcFx9BxyR0A38zsXgto3uN1LIlB
P+WMF8ft4A19/Kewk6bCGPm7O9WJq29+UDVrn1GCj7fGNBOjk7nx9h11/kKYmqnt
jfgt618glKUQ0tgPUm57MJ5P+xuoR8Xji4+h6ByQFB582P6fOSi7mAcqPR1Vc7b5
IaM7S9Q4ETysDnd6fT6YPOcXhgmMvFjotgLEfnZZfT3nfIY3h4mfTa7PZvMbTDBU
XZht6MYlbEM+JK9hJ9E/uUObb/pgZDwnEk7EUNrXds6N2c9sQEBneOaNQEFwmD0+
sOmwmrZ2r+iD4LHYRiXWfurzvAhyilme6cdlEeVJH5p7nkHgSWm52iNeWu7i6XTO
/vPAxLw5dTnxVDn5gH5ag+ZN/Crf/ByE36yfR7DMLbBnU9MFa39g+JnUuwd+ogJp
RJfndSqXxOe/dg6+lnUokm+NXDm8dieOqc9ln1o6hehEmx+XtSiOncG3eJpoLcVx
t+4cVI5j+zIMCEemk5fNPpr/N71k2ZGzU4+Xg030+LRCqVWOWmWdc+J6nfDlAWaU
Cfj8bkGtA3DADjjC3h5TS6WMO4xKRSUgn0ohNSvrLAmHzQMBgZfCe5V+gIDcyWx1
ayAujztx0GqAyLkADb2Af13K59+nKlzCJV5F69z9+gjZBY9jiQYz4gzAKCbK9Awc
6tIbaJXen3xiuOCNF+ftd5fIRpXNBydC1rgn1wu1bV6IUWPcTdwVGGHvPZY0RPJ0
7aMLDLVG4IlnIlmnvarm/qaBmJGN5ushcpew5ETrFZm37Vz2pE2jAIbkmLcrk83J
Zv0VcDmmHPsE0SPbH2NGKctXc2PyJrKBJz+ayfDBZbkvBb6sf1U1KtlRi0eQlk/M
m+sCMVtc+O+VmLjYp2ceZdoJmEblZ47DBr5n886aQXd1n393Cq7NWf2WV9A+999c
cnBhonxSRor7lLSRon5ypYutbFdJxtvK0XAlDgVsTbus9XiTHfN0E1leUh5RbC5Q
xphtgJfRC92ctG2NRF9ECcZc2rGjsx4RYjlYFgzKhVqVWFVt8LC0d2dS9BdYuuQ6
rCEyIfFe8VDDOmRLrEVNbjzsoskKxu8E2xYSUwIb77bmGHOfHhR6CHB2v97CLUaU
7YeTzfj6K0av2FOBrypT5Co0NSIx6NvleI/+h6o2UNmaAdX5HzUDNMB2Tf2AZQ6M
6Xo8imhqSOFBKiWJcbvdA+rGJiPuCqSnfgZnaYbNmEZ6ZePDTsewzDOhhvEGfoDh
PRIqUJd/tpe0M6LX0KpcAlUqRE9ImT4x7wZMPxXVGv8+5gG0zNlH95H5yL+k+RNv
ngcu5im4CybVXyTJ9ijzhpOXJYJMvO7uvM5meNXyixrEgr1mNeNw/DSSW91W36Nm
6yDg8UM4z+NwDSh2ezhKrstiR4o2fM0VRq7FEwTvjKw/PePQDhIiu92ihzsWF+FN
2b8WDudSeoQgKhhvNoQrjA/zH7p6Becn4ZSHqBoghKrbWBKwFR5WsZkebJONuDzG
f2ckb3DAXTiijd5AlGU5gbPsBFPKDFYKkMQ5gYFUNmD4nVRwS/GT8uoxjtBx7NH+
Ik7lfelhR4f+KseG6MIo248FW1ZxgTohGzkosHbVTa6IC1RAKmgAAVrwEvU4ejkK
QGz7suhGAUURXipws9nDrWzPqI3PPLBmllsDCAZkCabEx+JGBqUK8tjm9rvEDrBO
o7A2hGcodS91pMazTYoxUmShzAnlvouqDiv0Duk+lrgmSk33QOx+YLEyM8l4lSAl
FDdnPrRyGPmPM7WdHXejWLgbU3pR929COsVTfZjZCHZxQA3a3p+lUO6/248e+9vd
H5mD1bUp42/7VC93TnrKR+x/RkjvGqwr14U1R0COVczFRA/2T6aXRue4wj+PsHZi
2Tg4a+jt0zEYrdbOd3f8eI+TpIbYz1vhMSSh6J24UVxu3vDIItb2LfEa0wSASK+d
oqZVEJ+OBUm2tNriZuq50gFEtxj3ZjaNY77yRV84IEMyYhyDd0ibkiRtQSjKO1h9
EaJ970xCpJmaT8jhNSJ8aDWT8B1+2rYS5w1lI4GjniT5d90AcAZddNYB4bQKIYtS
HNhUvaCuE2ehWBPUQb89td981IwZ+8wHkPrmPmzjeNU4DF090bClDCtx5GvEGzbX
hiKjuqkdjz9eHKrNor39+LGqgfIWK58bhlQNgwCjNHdsiskOmkDLjDW1xHCHrpTV
CyKNgvUinuYHxx6JMgNRk7ql/JFITEvbyZRN7p6ztDaS+NxTVymxkcU6Y6KRVXma
0JjWYyox7RuEvIoKdu+vnWs85V6YD5TnESB83gCLxdiZOVvg6vjgTIgbrWPAvFZ9
/dwJXsrxxRy1MdwMmNyhT3yU6L+j7sdg3NEbbROk/o2qWh/pOqRwszrisDltlgsk
BoISyuhP+gVOAI8FXWpNk7CDTg8LbrXWGQKiLiJXqB3WnSrVupN7xkJnbpuzVVAm
r+p1JA8HvDy+E/k3IDxlKqdmsmmNs9Xy1RxaFs3sSip28K8GnncAJZKTA2ovu+Or
IpX4PjgsoursIJqm9WgJ9lZ1HuPDxMfhtA3xY4HE1G02aICTVkAX+gC+wrt8SgFH
SdlP9ndQAwfMgIQ98kDZtlxNk9VqMRaXACBVzEVwhk+Z6WjZkxZhPTAoDqAaoCXr
MB0DpzElzfNbOyTDEMW9iHXdXYDfVRF3hALlKHqSoVGBIjgxVcUlimEjZ808wr06
+WJiLyUEIj2cUcObgwbKx8s47nLzzlH5FLS3Oni61sjz3oTcCmaVJGUPYuq7bj4d
w1G91zEnI39wGpZ+ONUmbLAEm/+nStuldJNt4IZ9+RpDLSvDoXF8MvTYa016Oopt
nhRimDHg3wqIa4KWOYXGLdwzBfc7efnBhU7XgnbEhx4Kc9yiLE4eecDH494Oxw7/
E8PN5VMQ6kXrg3NNz6HyWsZy8LuYm5EKbd6oRs4MDKCWmV9eVdp9Fjhz+/e1aoa3
5RAoVX0X9A9Ta4h2lOyc7PWwa+6NlL6Ww2Mq5Vzj4snYUNSNFYyBupCsU4JbuHDd
m/0S/n156sRnZPrQAecuvlobhvRhWQm/QkWqjuitELeLFsohpx6o39xnVRAMvFCx
Hg5vdngzcHzZ4jisPyGlq2aNPK6DSN4g4Tr7+GhNggNydgqf+HgN0TBgIuF8ogM0
kS6/aP9R1YUul+YxVZHSfmoP49zJCCAFqPTCrlLxUsbYwjtw5WnvK1xsH5NMQpWy
KdFnFvC/EfpNRarEpAhjeKfDiaQ0ipIxXF0TYv1z+fTRe99H9fHKGemX56vmRMfb
6kYfViVTD7u96xonJChm+DY9FIVd06l4RiTKAa36BASe6zI7cTdaQEDquFiOYOnt
IYWy/uJd6jdoqDpuYzhFAg7n21YBs1KqA88AeBvXuLdTy7kBXJxaJqP6eKM74c/f
b2bnrmvlhWkCCBzKo3yqqb0g2p9CQttnLQJQr6TofE8mMFkgKks0SwQgTqOkRM7u
brMBAK+r+m0wFPakHMrU1tMtr4ELNGJov6uDzXYZRsujtuVRO+mmwlJvZV9Z/Z4O
8p4itkN8691NMCttIO+0T7dNGvBAXgtAuty8WiD/VfTJuDfwk5CAVKBKkojzfhD1
BB1aJWhwFRVF4UOCl8dG+ZRfjZaCmUKkE4oiaBxGTkQrIk4MFw9v/HMPcyl+3Wqa
l97PmaG2ddxrZWQFt1hjEPGYXbJMzVlwZD0J2ZMuSOa3NqtGw/tLamE7/DP/CVXQ
zbmaZ11WZDcqhuv++FIKXnNrnIIMU7DPxDXnxKN+qdrKIgJk/TTUyCgBrVtjPby1
fk9M6megkicY6GuZFvRnmE589JOS7Pmm01AXY7OLBTjQg6mBhMXGkFVsGg3g5B+o
h5VKfYu1kMpuZmnVe+S0bG4davS9Hs+36CMprcbimukrOaFVogAw6k4s37QLHr2B
c5oOIvn1tjgzu2mMRPeb9ANP+ybSQrpWDt4BnRlrXDMA0IMmsfAcmhIvyy+5fOIe
RV6l37HwqAog5XDi0G5bHPJgoz2AO+Iw8DjAvWHvmaiI++PoXXI3AQZSc7qOS+Y7
0m9takzIjYHWgySP2ywiQyOkGVt8RMgllYADFbnFydqJ+RBUeCyU2DcfLVxrUFjg
wMQ8DrhxxmvO1IvlPA2ew0k0SKe/xQUlEcGu/Cac7jAHZG6ZgxazVN5x5UsQuBb/
x4ezfw53sNq+2AL1sGv0hlrdKA9hNO5craM/p/jdxgdCEz+6Df13al7KLEAA5WYv
mYg1XPIs5ia+M7E2Pf3Hk7jEf1qY2JKQPvI8v/qneosEN7pbI85doz1W6mXxaPtF
ym44skPUq8Uvu9Cq7NStTXqtLMYv62HtMZkhE3mmG7e27iIVLXf6/tGecLNbP+FI
bYCb8b/Jig/WnRCCs2PER9fgKqltFI1qaVfTknkc3xDoXDwU0WGlQ53VmAaWOLq1
gU8ndLM0/bb+u+RjcTh4AUEZMd+Xb74WPLF9RRTQFh0ozY+SmU5YTEip7Ml0wHc3
/NWJn0l67uubqUJdNPJcMJVnAKc9UrmwB7xwOunAiHAKg/pR+NwA0onOilCCMGvH
P3RoqiC8PEZgM/fJIyTaUQ40ieks1C0AjJvQULF/3aP8ACr1wxUDg0HFBoIk+X9a
buTDRjn5209Q0+/gl271jR0UrYSWYHYOMI+4bLQhRyxqK/k6EodySW7ScjbM+VRE
3dP+CZq8BZPRI4Vj3435oTTGCvu9+CRinF+v9RPrVPdfr9zj1zGxgX0khIRmVW36
zz6A1vVF3bDQOmsz5tOyU0qanhDSLOXZDIsB2oSGukTQkiIAGNmRYFpuoqvDltOX
JSDxnVkE/LoiBb0kKbTGXrTlm8zz6bwviva8J0fEshqDcp7D9Xoi6oFkbUF/obUd
UatDwH0W6p9TjHrSPu7xvdc3YwWT+jt8rcHnpoBuM0s0XxG189KTDHzwJjHODQEx
gqig5ORlKfv3f1YQrNHdGzsWc2YWvTrG97Xn79nQvj0oHxHBgoUq89csa0XH+xKT
vat3irzgWabHZjl5fhApAiqVHMdLmkEtNqv5EyOkT4VjpMCRPycYlDvHBkdLisiA
V/YgKInKmyaQ4ncUll2r2yZhrjfj1WlGcot+iBMoXeqjL4jM+VL1NeCKfH0P7iXH
7d0JIaNb1A6nJ6gVHEohV6jSdhqrrKzS4ga1SdrCAnVopJh2t3rmEP9eFgrIUYBB
6UrgwBeMI81d9E192XnZZo6PkynuB0z4J0xtRsCXQRmBs/UylxMhV7Bh75yg7NXy
Sa8fQDu3120F4nZM3n3FbwAXvjTkHjuZq8qkVICh5PLdTdOknEtr5MyE6nmtrblP
wwsIWkBOglGfGDFxsY/GrrjeyzEyRGdbcDuLDQUgDjB8J+vlpeM8edS6kWLCumoG
TcWbXylbbRWbNmQY/ChJpSk47OhQfD46L6VlMJYmHCJIOS3RhvfxGYWKE+q+GbF8
tTlU8pBFdLp0J+VnbDovYkQbyT8Q7udnFL0jBE5vmG4uExiYBJJnUGBEMbop0068
r8nwjSykpfiPvhq1DZzzw4Y29NCOeWku/8xjylZmxQATVJY2y+Om81g9iuHnH2nL
LIqDJ2YFjXKZGywNyfZEXukK/qV+bldxZgzk2At23gW0dCTpt/WnQxV9FHSeTgrA
NuM9V+OwpbiSLQto8HHuGBBkJXVOHpOABElDzJaFdysvyJ86OUwF9HJ0ntrc1sdm
EHhuDFTzrhLZfcLtZZfQmCe4U4DxlQz+FcVh88Ro+xTopS8qvGzbObpPfARcAgHj
WE4wjOLMZa/3cnO0hG5gQjOCMpnaCFq5y3qyEqvJANNnJbQwcfhVi7QJebkws4yK
+R+aOKNqJTK0QQax3vl7J5KAEsVSO1EBSidc14fvbgVPzzZUr8l0K8Kr6nEUMYFH
qIJgN2hhUelhGy3R4xhKlw1DbbsbMpHeey6x4UwSJ/kkbaCCHf9zOmQUter56k3o
iWd6kTnqedAyhr2wGKxJtlrbb4wy87SqnO0rTg88+ijwwHcXP1pEvXnszIPOM130
M/zOKm1aY7DValL0KK6WnD+bT4y6GfTlRjJ6CWeM6UT1poKy3yn1F07R70aCJq3h
KS3cHh/bMKgD0VGUCjwMDZypXphWkzgW2IeIHSqSboEyhIcwcBVZ0hwmkSfnpQco
Hc+NZMCblbXJYEJxDDpQTI6PLYAXlu99Ghbuy2CclnZNB2ScWMp3k7C7MWaVfU40
el8s52eu2uM+i/Vc4Z/pEb2nIYUkVSrYjlL9VzHtwli4b3MIs+joPAhfgKucI8Pz
RzFcYL8rjldmZbScgAqj3XBbdlQQWhoDUm6TYv0gBiwjRODT8FAsxxb0gd2Iwq/K
+ZImWcUVCgC6TOG8yCB8ffILptEjS1aj1Du31Y0IpxHkJ+GZ5Fnh4zcmJoOhCThU
ERPUfzxaDgTa8m8Xd9+vlgbhyVfFwBiUIey4AO/9IjFy4IfD/wPJMsZIUxP4YEK2
vfa513iAz0+qM31ZZhHemCChWomQ0VJrQfFXnxqIPZyZ0am1b+R37CjBsjAbGV8Q
jZoVao+/P+L4SmiuoI9HHnwWMNBvFc4WJ66+LBGuAPt1IFLCBHbVc5Y7CpD+NbAu
o2GLMycjKQsYn9bcLK86NGyKynXi/eLjd4U9n6aDruZuGnDf/3/kuZkTSaKKBY24
90qDy9YPP33VnvRIA4uTCOIA61r6t0NuEKvBvgXSIKbhKrcBfEPaXoMgx2Cn1TRR
c9iDG0+G2BDGIGmxY9czaKjsqSgmiTZLgENo07IHm4DxOJK6lsrBckcqxROwX8TX
eT1bnMLD7g/llK7V4LsYt+4eyMOMtxRDZfdiFa+PncMBlr1AWBW7ctrjbQLo79Ef
OUJH7uKTiBERip4fYWp2j/0lxoMKCJPNZNKMbJ+QrDhO8fhmJk2LjVpzA+kh/jXW
XNdIvgcnnNiqx0+ilt1s/bGdRcencf32+V8yFYkRu6uUbswf3F4m823TyuQYzUGe
khqvDEKUXS83UhXOVnFg47ax1dDp5LYSa0zX77VgW62yOHFrsgEAJF+jyECP1FWg
WKcpYyiPM051tY6Y3jyfpe+Xzs6UcDKs5c7TauoGYO65+T9mf1d4CHXmw6Nk6yzF
ORdGvFBK8ZZWaaNeumiEF2sCdKbn9DMb2Xw0iiHZdBjzCBgdqrBuTYDfoKGtRNZm
DJMOkgP6ApBDp0P6bDUS/NFwjYO5CdzPcsKogvVdPR14eEcUTAJ/rLrvJHtrqFDf
HXyIfXpAbvoAzfRHrUwHr/NE7h9ymkgqhdau0jLlZz+Azd9em4Leys2uni+ZdIOh
1wOO0J70I/ZJNg/UWKne1vPL2sgWzyZ8lfMWN4ieMn85cLFhaZQpcGWQCp6dQkRA
HqyteGj8XEGnWm4OwfJzVJ2YQdQuW4SZKKKKgV/psLsH0QCIDn9KSK8XzilYP1In
zdhN+ku+3Q2dIJJ1QimhEQQ1B2ytoa4xgMVU9Opwx+G5neCRXwA9jIwngzNxEyGx
rqucg1W9Qy88SrOw1c3xRdk8XS5nZ8zU6h8uiz00vEB4i/TOjVSqohz2Cm44Zy5J
PztmhT1H2e+gJn0ogdm+z26IIZLLO8nIZ4q7fzBNZludqR9g6Ahze5KYzEzbhxJM
2VQaim56muhhB0+CYFhs4K3axjTITNwgiN29PQ2Iy4+7116oz1NXNB5yAmDbY758
uy9+sFgRvpXKollcEYtpwbm3bDUmujWG5Wmbr8GahechBbk5iY68FNKQHkYcWZHW
aDHdFqMG3KsrRonWcaGmeb1wH/f2eh+figggHdCnMMf5B7qOsP8gcxnRT6SJHpwe
XU/jBpCieQ6lQ29SVX2FpAys/hI196c8r3XPs5R/XMe2XHc19P1vdWcJ9RyzuJzT
4rLul9jWds31ew2AkJtXWvJf/wYCjd8rDW7C/gsqf4fi2OKIrD1v14f81+5BsVh6
nFmQT7G73pNKVOEX20yqPScPtPde7HP15pUF6JQNDLocdky2XYgftmLttiQCyywI
qh8Suj4lM1qe5mUG53toD0G1ZWw5kb1NQJRJjAaKG7Yy9lKjZLj9ThsseWc6XY/5
Y3l/M/N/gGN5HcheAvbHeLkkfMmzvUtXcbk4m/i/dFv03cFhCpuwJVVclZ54lakt
ghOLXu201GYIy8wrD33U+yu2oZN5QKWEhDeNAt4ZRYxMcPwzrWQtJaKv7/Mo3KR2
dRcPQF1MFM0BBUImWGmn+DTzyO1GnVPkrXtu+G6gURsRsc8nk09a40Y07OpLUS+9
uzxcdScwWGWrnL/UEnjhaWe6TWWizTEhHPcFsPuKceGuZBjFMlRWA9m2sovimlWu
VcIOOBEWlfASmzZiCyxfY+ZibJG33V3dJoxM+1XpRtUzGCiFQ8yrw3y7GrYFfIk0
WoQumNF8V6DM13J7gJ561b/Em0JR4Hmu6boCzkTsdo54BRYzRTxc3P4czTeijmTD
/k2tDca+v4XbdnuJueqIwEtNQwJ6sgb+H3BZso+xKPylGscF7E/J5k5ikRy54riQ
TNNY3DwWWoAJZKosApj/akYuMo9mWunEoFsr/DOye08ypO3x8HnM++LFZaYFxUDi
I/EPsVmreFGDhH8dg+lbNY5w9HsxCIH79hx+lOu/Ny6176zdzCDcIKHhaNipwBp2
hOct9TKCBrb1PTJw3hGgWE4NxKrdAyRPkb/L0yeXWlpJGrYi4Xg5siirRhALtroi
vq5QEeTfa0anphgcFx0kpH5NrZky4M0BUr7KhGZLr44bvdxfvuDgBr2UVygZrogq
GL2T14wTvHvE+5CXlHC1/OfpBHcKtRWXshi9GGVRW0UaA2XLdiudPuRlUp4IIDNj
k807FW//+iwAZm3Ax+H6cknxSashrlFtex5rxTDilNapZMTJMLIMWKvBjFFZ4n+z
/AQ37NFKkzoIi/s4+mhoXAuDeKIfnzPcxPUCzueXxqMHp7AacrcgswZo3lywg066
IFWrVpcf4Xiel7SNxt6fThx8zS4J/reFK2+KhnBmDKirceEraj8N5tYc17GVNEjA
XUT/VqwXuWBQ9c3DRcZiPa77rK1EyXldzzNvb80BAO/Y6hpulSRpzRuRfje2/g0/
hePkWxwiILLeU0hUmNCfG8tcd1QPYLer7K0ZPw9uru1rNxktRXdc5CMxjUkS89Wc
7r/P7vjDkM04v72sDM4Za4V1HJ2vnelz0gtalmM0BLTU9KEGVssFVZoh/Xanigm8
fQ4pziu/CMMaTEZuMcCnQMliiCqAVbYKI9729w7QFAG3RhjboOoMVlT7RZgCVTxq
RwVUf+TW+zBy3XaFKFEqQYMu3LCm2lsu73QOvFQmGpgfWYzjXgGlfXX0N06Je5uT
/2I5Cxi19ntyLrQjWWTqDbd7+PKgLeSJooaZWsffmEYbQj0QhxcjuKtN7Ohym1Vw
TqKrAIaVf6XUe7rzkOdqHIugQM/LEiKhM4MpM8n8vAq+FO3KFyUUtpLPHXyCueKY
oSUwC5v9SZH0RBlinhoMZJIL0mTu0CD0bJwAPlLe1Gjmi+/ThmZugYLW5LeS/U4f
uHjLwizUVTK5m/YpFWVvhOEHg1DC+wg/GNqAzF9ms8jXIlytM/MyUIkbv17NdNaq
4fD7i3aWNiynn7R46TZFnp+lxh1octnBjWLpY/JaqAv+KWyS6A8/qXKlN1v9E/H+
dRHmBd0aMpHvIdnGbO4A6q4y59aOI4jzc8RiR4sfUB3Otghh6JuqF7wLd/LO/9Bn
wodwTWGfTg0a3v+lrywtc47drscDO2UUo3jLQ0exqQk4Rmq1EtaXTHMKpDqI7kca
bDp+HauAJUrdVmjD0PjLfQTgp6Mwzn+938ZbljiyTa06ypFEv8U3lwT1hMyELNjM
Ey9PEOFG6FyoD7XSEy7yC1Az7Jb4nRdaOv5EYfrLWqT9beeWkL9Ztn28ryqXw4EN
87Ymych+850//yCT0ZpBjWIIqiBrmuEFYhhY6nULNZo43Grvfuf7DOcskZ1rYJVT
jU7/7JHQBjPwqGNkIYDtvvjnbVKNm9+D1jFsxnip58JDZiYkT6GbvM0AlW0V908q
/JcUV20932laKrTen0yev8+bptwp6WjNCoDnQn4BofVbedICyMjaTHSCI0m7Q6yY
xlZqaJVy68xSSu+FEAXBaUOubtE8FMXcV8NgI5KmvlB/vSlseWGtVtZq22jNmKAW
HymHHnufdeqxVxdeCTBoGQpJMDGoQYpmIf6pHe/zI207M9kgF4fxZnS/cJWxcaB3
/YJCczaMHa/cDe2oVNpKH80F88qRQSvkii1aWvx0eVhMO87GFSkzKqCyYOYRyQsN
BZ1pfJj2IWU3tbShKQYC+qGjQx4dG12HMgpHbS9yk6hlUakpb6eTKmp5x/JHmCJ6
AiKXORfijN5gohwf9JJCkokjCpUXASzNuDP+XRTUWLFTYc/tQr+8Eu5JDdCfzaRK
Wd4oRIuATQS0/ocl7SZFSkFgSWxTedlieprkD/qcbrc7MjnoddkLpQH3jooM/bqe
Oj9AWrpVCo74KWoVhEJgjBO3l02pa+Chks37ELlMrLBJnQw02Igh/TdfFqC3tJ8Q
G0xAIPbDXi+kujYQWywleUMDZ9FhHWJWTi9m2yY+6G9hGvZYKC9TyFyrnmbeFujL
3kwarmJZayPRA9sv2bAn5cXuwkG/9hm12uYgpYT9HHO4ZVkTgFs4NJ5e+8t8tMFV
jX+KofSQs/aitChr3ySoeUS29V7JQBggzjXVIjpiFZ4ZB0gsagC+UtzhF9UVOQRZ
PBZoKQBJexd70vTAUWS40s037teZQ/bmxv15XYaSFxLNZdIV7zGUJkuu/Dhs1jzN
of1TkFvYASUtYAIpO88hieTwKZbQUvEZ3ycEFYMh2MRTr8oFbNKqVe0O9dRN3w4t
OpUR5oKfviD/uDZjtjkMo0X/y2GaNLfINzbFJ+7+HVRC0prxfM1FYfTMHoNwiVjA
oBqo0bvRx9tBMcqhfXytvWYGFqRL7DfEScXOq4BxqMjS+xKDn7Z42jc3Jm6VoeZN
bjsASwBFyVSOPNwW5tnREWCm6/ytTAa5BzNuxh1dGgR8Ni3m7AxVWksTaASY2im+
6eN2MfjyXb2UQLw+yuD+InJqyNy7LvlzWpEZEUocr5Mza70Rj5nCQQfqk+LDKkLZ
kZTy5twZxawMP/sRck37G+Q5k6maVS7hymrV6Tms1e+g+5WC1dwoLttnArJIOg2V
2S4ZnEdGR4pYCnyS3jKmengPes5kUoHNTjAV4l+XTOLFwl5JfKuobWsQVsl8jgSd
ZCKA/RM+28m+wEGRmZ3++6h2NfjjNmCSW9p6f6XXcCDCnC+kKb62BadqbZyHKkqn
jAHjx4myuCl4p4Rg8I/dZkMQafEzDU0qBZKp/mfdBtKx3bE3N3I8cUuBFz4kIoAw
Vo3DlZcf/FnW3VzAOpxxbuHHNfQ9MmQA6ykjdsDj1YV4eaAmbpOlzsdgZl5gq+UD
r/Zrfc+NClifPsxDkDaJWHfLXV+L7mCBn2YB9FsPZ4Rvw9kw60SUhiBaJoJFA00b
WsVGmT0REJ9H5FapXAmrFFbbYZokbNtvSbAnbYdgw6dky38kRAs7dvAz4egb+sQp
6qLbvZMdni9+dkxUrbkItnw8gWI6evYUULREUzFGTzUJvsgLFdhl6+p5thAmrZM4
f/hhz1ZmhT4VwK4q0ua3QfdeNBzNkcXrlRjNUu3EGSTx3ThAmoUby7FpD3I6RMau
8zreu/CO6Psx2CSM5fJZkmWBeNfFI2GLVrxti2TZp6+ZqzoQrP0+xrGphFOrbKlB
B3GEFgf6W43ftfKVjlYYBcCp+ksQ0sClrgXrDLEmJ7Vg0QN/i2JVVymQAaVfObFl
WgaxnGAv+wJEmgIAq9aAfVALkg73CAQZi13dtR1R7HnqodDbCtSVOal3I1TlU8Co
oJYE9x9GXajO36eddeUb3CPUyRWVy5M4Pb/mTDtoStdFo3Yao6TJDuyj9gtHlwR0
o7OwAehp2XSg69pO/AQNuz5Sxf8ADTqHue8dVkUPb/zHk1vpi8ENqj/k4qYfU/xt
bILpBqbmOZo4Kcbmwxap21gIp5Eep3Wb8nSIbNa8d7iOw+mabOSI6f30sOdehLf/
O3jsczlcx9Dg8V0yZ/e3MOvEa8GZD2DFACrHc1Jy3LNOCbnUhud7e0XCH7N9dtwC
S9ZShK0HUEvuqcS8m0eEuF3WJ5xDUtBmEtAviveTOL+wiWObqWIVx3sSifFbDwJK
GQUwAxE3u8SS5eAsJjK3Lpba/+54HdZOhGh7iRewFAwR4cJO1oLohXbZIZRVKGmx
NiDxzLB01wr++DOnqIWsk3mWCca/FytPAZRjY76aVUpGC5KLPtfn6AGc0wi+mnqw
g/qwRrofoN8qNfQD1eKcD1JzPX+65Y4eChvAmh6PmphZEFtmsXrCMi93fRX4pTns
FwA99k3mfA1ZftPZ3sYcByxHbixyrFwsBFJ+PyYgFqPmbBkwin1DAeKHSnkss7cm
CQeiJlpCSIfiw4auHOE23Te/OF4I0izHpBn3Hc3E7R/7sFprgu0Cs+AeBbMD+kh7
I7s/+je2ijxgeuFEsflA8LXqAoKHfYC9wQ43V6o9rVXi0WsDzy2t02eRx3lXowIP
R84nKtK+GXuZ4A+e+wLbDpAsVPqF1gRy0/dUUEN3XT3sD5WVqrRxV+MlADo8uHU3
Nhgx4tN7LUK9M+yJTuPqiMvBs0ZBhu3Mlbj+QHRKjWOmFiAOrWZ96TAM9zGnMwxN
rqXUtwVl3ZG6Y4vMdE54AO/jMxgRQfKxL4WbrrJkvOpspiIKigGFdl4vGrtJPJDZ
ttFkTeDSYegkKZS7YzheTN7qj77166CfXFWaXfJ+4rBfgs9Yr7voPFkL71zNs/X8
sXH/dLi6BDHoNmX25YJ8VWVM58IqxMfp6MC6z4/lLkwTXbWlRuVlgt7T9SRJ1uiu
kN00ST7Ki16feykpR5fVY7ZIHZ17QftcLmT3Eun6lePGLEQGT9uMwIjtp75HJN5w
tI/EFAvvCZfn5Uoo4RIYQZxl+BaCsX73os9qfkBFGyLrjtq39xMNQaZEnKuhmJqX
d8kcWLAvz4Z4nVto6x+far1STV+nZkt9nHG8hqrVeXWDfSZR053xQTUJbnRrZHf0
FnoiX8JnuqSizk2Puv8hsv9DeWPGvJeVvhv9SrmsBMEEjbdtV7RuUBzCj7lM+G7n
boOMqrJ+yHnoo0Ihzd/LFMHCVSO9EHFYZkuDHIZrGcQrA/mcQprTCb44tDCYmlJQ
n1T0BH2m1ta9DsdfTSXaeTd/qCYAsDRRvraBIBDBVws1p6jawPdwYrbrGTo0mjSc
bCXpssIS5/LmTFPt7auiDxgq8bTXAr6crEDNyhVK+GNnSmBfGlbcPfq9Iyon1UVc
bjZ/4SR075rdYiWsYDNwpP/CrJvsoyz/Qjv6vBH8JvVoANV+KyLqC5iCeh2MBjwT
UPcCAh2J+WJ13LaXot/rogMyrnsZhAfGVk+rFp8EwEKAZdZu+oBJEJH+dVJOw9VH
QT2QsE8H8Mw4f80r9qMKmUW2+Ns0uKbhorJrpdQs0XbabINi6jeNVKiCKlXmVvJN
HUAfNglrdI0NflntuYaGM4MKtzI+ODqMmv0QwbJ60n188C3HKpCwRmxTILG9BMZR
MmDPmPEBisDoGbM1l8II054l9y1L/fvJTVOxShHt3HnbAPpSvdnsbvsA1BJaEZ6C
fMAo2MIPEneZzVn6MhdqBCqezQhb5qNGwWb9Zn9fcL1S7gBwslBGipufSpZ8xMAS
9+5r980xi8ZgCPqdaV+M+5TQl2cq6lO40qd2664sWPSFoDlZV6mk3LO4wyETGaIu
sozSnYLP4d/SEnRfn47qIOnci51Bq894gCeRBakqf8033bpmLBrZv2Lv5CmI6q/8
SiXhuZmj2276upG3ZS1FTUzAumoy8y1rAlj7YnJaf7PTE4v8ZhNuTdjoAIfb5nhW
r8ZpPzZKDw7pKc64cIHzdf3gwfBmhpWu8SJpcSfoSJvtwMSGIgAteGkanh5ngdpd
lWAZ7iUDEKp9V+RzsG2vwHzG3+6KOLHzTLFYP0NNd0FsTqYzgs7WEYIH0cj0Yy+9
eduCVujy0NCNi6Q/JI13XgDFg2zMWq2cCgoNLoS6Om+jii0+3x0N3uHbyIUa81rs
8NVOg3Yj7Wj56k+7vDt/4GxYsaSsIyNdlC8NJ84GgaCSwBgANI0u9hf1PpL8YKJR
u/j6u/mBlum9U/G0xRp/4rt4Of/9DCcKjUKtR5VYRO64+USeNLMmLmThUvowu2Je
nweWzSpb2RNG1yXcrBJ2abfNvcR1eSdGeQjb9eYlNuSOtsr1FsErOvgVa/d2Jztr
2Z2B7kI9VwbWN3TxZ+p8AOodTgP0IVmaMF0qILqE2BZz0+8HlBHt+29rBztAnoUG
2VdLczZX8/abNSPHARJqrD/fB/4B4tQHtuycyJfvzCg+kJkjAAoylcdXu0g7gNfZ
ZfaADZJfToSUT+fXUCKboMAcEPGB/Fs9z8iltnacbCH7fjnFBz/bTZg3pz4KY0O3
4HD3SBLW7Lf9NJprJWxLBF3W8DDACpvnHUiN/sBnnaHBps8y1TSLpuzt4bwMxZBx
FOheNXqizbYr8a8oy5u/C5iyleuQHc9aqkok0tB0TYruu1RaLA9JQM0/zfjmiaSK
7kCL+z8O410cgzeTAdPCqbHdBSudmZSgbLBF37VkbFRdETsblRWjH1ZRDPXrKWKU
nX+jhHXKRBT1XfVX+YSIrqIdoP6/UJKtXOcEXLenMsoV4oXGxK4i0r2ZyqHyn+C5
o5ofdEgJe7rrOdPDx7v6HRcoYm5LH94FQqa4Lj3+hRmAq661HUmNEBGqEHqxgOoh
v35YpNbCVX9MScmrHCGuTidXo2Gh13KRtjNQDp6TEqZ/ImPfa9Zt1e5qp17Z3Snq
JJdIP3KGTzk+LmdMarESajuEUuj2ClxM6HGz6KdOVzlxWnGNbECDJSC9FMnCFdYf
q9qVBb+5+Wnmtm56KYJ74Ghtl+ZFvREzjb4bq2MXrQJDS2QqTc8Gj30mxAxCK1l/
pETLar8G3JNuFB05lHPVYxU33g7GAelyEiEJVqFsv+u/aU4najIFfKZluNcmBJij
HOaPKb+J7GdBRAOXnKdN1LVZa/t0aTWqZIpXYBdIzsu4YEcxw0NNZsc/RaVpIalN
sKHE7TXRSFWHYsnvBXGBxrY2kq09tcmTGbujbGKx/pvfZCOsSnbYsNoK3dEqsfgm
u0jXSbFXiohB1w0Xmxd5AmoOgf7zAGiOIxBljf14G8RWJun3BxBbaz7GRB5Vey3Y
UEMbHMreQQWQETtJLaaOODANzhmJ3sBtSC8xtHk/AckfvZ9S5a8l/oqGYIsmyJBv
TZeMAvr8LX/HHQx4VoY8jcJmJDSmjpNLgt9Gh1AdGQwLQy8rWFo5qdjrF73iig5v
eCME+UggV0sHxsIOB8zy7/nPKeFpEO0YlsmHZ1gHGAuF0Iu/GPcwQs0AeRESuoxC
3MvvFIfLrJXL5i0AX7mqh4QN8DfvG0CCRmUww3jutSFEVvjr5gdrueNLmTxF4up7
3xgdgUwwkbctaqK5OiK3Ren0WVriIK9B6ujLspiLSimKh29xfN7lXWMioVVvazLy
ll6/0XPDusi9Chg0W+m/33v2ryav+uNAJuWH1UYTVEhGU/pfND7ashXUf9g37wxp
IHPUXtu4Vn1w4hdwhg1yw+uGIvUsQ+dKw0g6joi4f0aPKlRNQCof6QLuwdHv08fR
5TQpI7iDtJ2VL3mTpTwrwzcOoJ6YsZoduv201hBxLAhYgujVO5a7R4o/LWR8Lz1V
09WpnG63dzwTlb/sh0TWgmxlh0lZWt66z3AnKLeonV+fZnV9OJ+5Okfg5j7txkxV
pfU4lEKOJ9OFZUhjpalEJVNhWT3yTP7L2S3Unrta+Tbo0ztyipV1I66Gld35ieqV
OzlQtBB6ilHcxFkEZSoHhUp+LHXaj/nI748nNKp5LNKPujPl4zSSBH+V46Zr6YnS
r0DO7+NHrwPCDqFmzE9/VeyubrL8zsnps1inVIM0d0JRbQhfhs6K8zsB3F5LA3Rt
HPjyQPfOfS3FsIYUvQM5X69obKG4uYD7T1+pAgyAd8IBuz28cz6ba7SBI3vLJCrI
XkmoxeGT93EsCE6gAzuRYkmc57E9Jz+MFlHXDzTt4yNl0Ru6+pl0lkjnA3H2XCyr
nZOJjD4wUJOfs5rqtCC+336NavHm6tztB7O9NqWQYK0mGdA18uawG+gg9/2W9OI2
ws5U1xTYai6PM+QoYfSwGvDfhOlvL4mUObUWuvAH8aibEGX4E0sTUCNKlokdKjq9
NbAQLHA74UJS+in+5j1feEFnRWi9qP3vB4ovkjCpCp5SARomPM98ccWraVP4J58d
yLnO/npwuYkqOdD/pBn0GEObVEBKH7t8JX2xrR3RZa04pJcsx/7u9xh3urxVR0Qb
TU4TTbswSbJSlFXTJZkuiG1HAcfYYrsPmOEzYOgIAs8y66jh87FIGp2SOosTRyDD
3WBqwfTSj4HQDCwvdRGRf/PGgmIaAgl+RQEEdYBTFisBgZRbL8AWnKKJ5Ymn8hn+
pCiaonnOpelnC6idmsP2ZffzcItYTgjGqObLa6Q5iCYC/mRvL/NO5SHHcXXGtxf0
J/ayol1KRPb6xMU7JdcixkhGdXQTtyNqOtmMDPO0kk+1HJjvE2yiQEA5dj6k2L1x
AdXwim9qRVZupFHVZFHonJDY2oRP9r6zu5Ma+UNis4Ffg1nDZlErsZV/ImfjfmZ+
ckBxXL6O3qmjsAiJ0LRW7wCvRRtXc0TCNSU6uy8Taypt7/HVn1MJZeu1zG9Wojax
GQs0sgQFYJgCX1gIWxmtED9F3j9oI4x/eSTHBxEvu4c64LXzIxHgC6Ew6ynIrU7f
uA2S6bfrQUsmz4cZsijpPIXAAc80g4emgZ+3IP8gHPdfAvT4iOiT2+bWAkKVQlej
+lQfDk8iIcFSS+hgZLB6yUn8TxFM7XTvCLSt0sLzq9NiQmFmEVPejLqo6gHesmzg
3mnctTDZg5UkpZW5KJr47MiQqTVEObtInzRs6+f6OYve5Qsy04wGl8wZNOGBv34T
0wGRzdvWiCrCOMHkLvfBAACJq6RUAJyeMzatXbYyMNoej9n+S/E0MM1JPes+zt+m
1aFb9zy4d/iwQO+Pu0vF7aAhvZqDNeDxbI9tOUoMDX9+ULi5ZpGwlbd5aTubUAns
8ko8dvHyAe9j3mHv0UHSd6dLTpE6rzY2HohSG0Gm8DUlErghw/SMAUq1Ugi5p5/j
nDkphZIpMqDAi8PLTZDJH5RpcQ433ujGi78yWW5E4OGUB2IOMzpqCn7QPBAsx0yq
jIdbNEKRcr43u/4j3iDPamZKsFrU7NXGCkPCxEJLJC5nxYvAmYLEscQxUV6SMThK
37gKjCaGL51tsTv3h7rXCKzWnprn5zkrkYimaB0o9pkqHcAlx17Z+UHxclXS7N/+
N+FFK666WmkJ6RQkhh0exR5sg6LBxNx3UqOgqu68aXu56gy9cEQ4SlbZ/mm+pthA
3zra8DzrxppR7doz401VmbWw1ysfv038aa+XLMoDz8Ztf0E4SLkD5lI1zZ+fnRr2
RsxovpgFuv+lFvZfGJO5mZ3wLKw9D70fdV55QPbhwhC8F6sQNqz3jd6HLzIobIk+
QwoaQ3rQt8qV/WvF92Oc0iYlcZXlRNW4da8hw8hkpWOO5oPk5wKXcxuAF5qMDtJV
C5kw7cW5/rDBrU1L7OX1l2tps3Uld4WPEWFfjwfrq7Z2/hw+tenT2QWpLeVt3T2Z
xau+SIDifIXR3VcY+sEJIFCTaoi9uEZnJUSYwWMspFcRJYhFuuK6KlH2KAjNTXAE
PpitE2lNQb5XfnH/cGx8COBRo5RcUvlVH+HrWDeF/r50QPnBwmLrXZlfHPiWv9gR
YzKbeB/Sa+xrfcbMOL6vvm/SXTl8qqGcExyD5EQeLyoIU2iDT7s5oiPzCbT1oxA3
fP7oi+5tIA2zLjlN9/M9/fVgE2QCEe9xdNCYHs1/lAX9jONKRhBbaMmLSLHz5Wg8
5KBr9kmzPhE800c9U5rJnJxu0LG+qYi1BU1lwkmCLi5nZWZAI4jEwZCEKtnzPT4I
138IdU2uWv1jLwxfrUeQbAF4cgrXDIV3xFP4y6HyCL4HncKI2GRPDzHaYQ9lksun
nkSCd6p/+aC2B6bI4Ir+hLgj4HwGjl53eT9MMcxTXQkrajCFoXx6sfJb/7qSipQu
8xKkADl71bNqd2aFbeMJZ/xFT94dgRRcQ68ODxnZuJMDZjto4OgMg29ZAhveKGFP
GfUMCbcXoCvVIbwFeRrZXS6ePWMN4+TkNn+2rac5vwLvWTr1RpyBdskbnKllgVeb
sE6Ty7wHYmm/iJc8AImHyxLkabqXsVJpaM7Gg59DqlXKkatwQ1d3f2urFe9od8T8
I4zmC5YhrSbw94Y3OhA3i3V6NZx/S9/NLIchlCsxmlJzRfz4tSORRXpl6EAlnKIt
4I8f1XrV6TE1gen0giOjkowDis5b+gG6Iz/d5kYYxNCS/4/wGhOpJhM1BWIapNyT
PRByB/Z8cdikKTKZYCr+unkDv31mWYQwEpcONG0jVVGtM8OoDHAAL/kyExy066Wd
wo/k/h93n/NIBA4CXQ+EbXU/JyrZKFcH9fTRV+2mTVlKh8hApLJlrCQTbzHZtmGA
iiL9D6OpImmxta3ClvTJtk5P+H15CRRGGoV4LakxwqLLjPwHWBMhMgP/EalB0J1D
WyjEB9DStCGeI/w1RoT1dXnGuPRjWnsarY+7BZwD75598d+TWR0impkUyR/q1SML
HBHmeLkC/m8uG3vI2mdpo8iMeD6oHlacnK4bVnuv+YD48je/oyF77JjosYj8Fbm/
ay6nnzDB6XlO2FczdmXlwRRfCYzBH6TNCHLyf9gkachdeB55nVHbdPy6mI+N5scX
9T0Rw0FRadaXS9zsNnk5nef1CWNizlOlNFr8l1/MuSWZVWEbeEzDmOKWsjxN7jVT
B4zA1y8fqAP+QZY7tYrbYela1uz4bhdxO6SCUwVZDpZNqdX4aC1Hfjb32OL5D9uN
ERrNXXxZLIbvRCSzRo6gtYTO2K/vrYOZfZzS6pmSxUoismyRRzuB7uwkZbY+YANa
C8A9998yUVp62xBKY5QkOv3+cRHIQkjdxFcqtLFYNghbjAISdpFnAHvyRoKIyav4
V/TCw1BXiqhw09fMn2HgtHgVaT/mUoTgq0Fq5a75Eu7BPtJvJ3Eou0C67oDl75Pz
9sk02NZbYfldNGhD31sWe47icHoXTDrH74sglTbWSZBXHLiPbwir5o4Umz5b3iBv
JDrynHHEJz+Un2TxmmtZQxFlXCBqwYg4ZYnfHsiwLa0KIuW1MJRQGZEIj1tsZQAk
eR48vXTE17CuUzKmYWlcVahpLOJN8jpU/6ZWeKoiq5IRVpUInZrTH+cD6VMaq1J5
0XzlkJmbpdKyOjmkO53R5vQ4cLHwZlWrC4/tmZA8UAixdlDqXYOXWpMOa1EhW37l
UtjewE6rGzeVen5qGjGwKPCotmcd/vrV3nLkzeZSQGwpvFSjteVgTvuETptUc338
xxDMXzU9AvJgwkF62aIajuFx0h5o0EKg3C3ZQ8NXo2U6OhPi5XhFRIAjVLe8Pkik
N3ot7OSAdd6Fp24tKIqamsO+95xuG0aey36w1lfPYWoEJMnYZEES1oFJFyq+pEYh
/88v5XhvJ2qqXNu8YPI/1lOTR0uHFlqVwfaGzRyGByu5CCe8Vmm/wvdMqefADg94
Vq08HB/XCZgFmofDrjiHEgE+NPsPfXDr8F/Lb8e7vAiqsK4+TyXna7o4jAjX0iuj
O5nWzyX0MHG4o+fXFMPInBp9Zo9qj+p4+9NqXU4AFBAwhOn3chP7To4wIDzWmRZW
b4k9Cu7F7e2xEa5jTovd7bghHObwUVOZfo1IsOu5g+UCATWyN8ikw+VTCjdvyhxW
AJo430ZuINbU0GH7BA5tyr6KXnBktsG7R6Clcn8cIymH16JgqK8cuzTAdz2KetqQ
LuWwndLO5MW9WwE5K9XSwuv26+SFT3pCdzJGvjoUsiX6h3Hip0zdmk0qmkPq7KkM
RwNiY/WwbjkFcPNb1OypX62aGGpZuCKtECWbhba3x2HZRQjt5nu6jjIGtJldNypU
xgif9FOqujEKYb2D3ZpzSYQ37QQNtYs8mcn7aoNE3UIRiqajTnLC0a7ri21gKG16
evL8aMBuVHmOGJzgDZcFVdlKTeXSdvggH+09cCCGPb8Adl8sDheWczCynkMHLzq8
7xeZzCBuUTEOgUuvl+wsHp3Ixxv+dlIvYiG60Bi7g/BSrODU9LLTQYGqvq59H4d3
rn28Hr2VO8GWZD42whik4NFTgy8dGLKK808NQTLbRRe4eC8cE3YEB6wsfv/BBIrL
ss+yfEVBGa18Bm3XPpYlkASeL+7prmDAmoE4WkZ+4+/GLLXb9PyAKgl+m+gpT3Ay
4I+kPdJkUK0fX2/1QkFfcqy9kBokYK0N0hXsBtD4z/1/6LQ71JqNi6txzMUrSL+Q
b01C87i6KPEp0rAHO0KFIK0sZiQK4TxvXlecWLB2UhbtBIU03JfUJYwS1gO/oIxT
3wj0OiTWbe0Rqpp4vz9EBR8YkOHWW0Rg1tZ0cx01s9O919rbfbVjdS+UVniodwaF
tia7kZKhJAkGmNLtOoFBteXat3zvbHxQEHZrhBZ89LbFeXnUaruqhs67znA7Pzmw
KAwZanY29JaN/1x1VbUoV177vPvEEgBfcZmnT3m5V4lwJmu9uOW1T/HE3eexrXoD
cF86h2bgwIrBA/6xKVAJp3OR3RRac8Yl5EFx9PKxxMHhcWEk08984YU7chw5N0l+
9szDKQLlLioKPYNDa8qekO7fKTSrjQIn9Z5eGPufkM5AcRoWej4KxygG96htTMDN
EecS1Hm3bCt4lvXDm+l+VgJUAk1QtDIkfgZXJCChH9QfLQndOr8jDib1SCvzK1+7
DSjcGxniui0bVVoD1g4geSTj50hSGINEKKWB7wHEm/jc92RBd4o9rWbtjCQUrzh7
Ke08B73dFNdmA4ZL6SSVWnXrmPk7euJX60x6zds5FfXrRJrB5gJZe2PmpG+0o3VP
WsUiUoA2J7A2aO1ojS6w+PTtMHlRF31pCaJLyryuHLxhWY8mfp1k/TE9lT6sXL5U
tAIqiddyDyEzviB/jAs1mdQiczKNkIdoaF0kGBKGTuw4Bp8+Ju5AzIkCK1VJJbD6
/gcVPatDZfN/KIXAYg5C49VpTBk6FmNaVXeIRYgDlqLIFpiEsW9a3qrpD43jNdR8
wKcFkk6sdXypWVsBzP+RPZ/H2ZVT5SYCJF+W54YLV63g6IGJS8333CaNT3K8JAEl
6DRVeOIYZcSc/iAOeJvRwSzFV7edX5P+f0eXl8fxYCVXVIArnqWLO/mVjUmiWKtX
wM/J8jj/k+0/CMhsE8c9U6eLFJFl2oZjClU/mBx9MznDIFDePwzIhKLU8FaiBbtL
U+KqhNTDg/aqDPlRjmA7AFuVxgavNeZLk6T+gNLoaanSCcjIIaQFoXCOwhnKOTZ/
UcnG9oVM+A+EYRqgsCDsfMbUNgdRdXyys9E+Fv9hN9HNSUZz0wuAXtW9IobjN3qv
5iEO8ZDYrML5Ctfze8qpWCMztvrupJEuBiWETCvTToVURRcl7+jspfEfJaXcvZbh
v2c3pYGAdBfCk4Gp/ESv4Is0TnwxTKRveAf7EMQ2I/oVN6Oxx2/MxG21n7mW2q5q
PuQxXqaw5rNhz2U60Cfsk9WqKHWlVgzPejpJJByau+c9nt6JcIr1m/Ue7Yyjwn+x
NIahM1E1Ar+cBiTg8WF9ZtHEUG8z9fS2logiCEHg9QqA3A9L4S7REyZ3EYb1TTcF
okbH7eRrD/L/1WSYuK2cvoheoHZkF9SF3/J4rWK+mEF3lC9i5HNx6ZxuXhg9ozHS
5yJePjlD1tjB+h1HzIIX3ui6MAhGEOhu4Wy/eRQsfmdGb9IvHS/xMqzKjECJEGOd
BqwgLNIZPA5JU4FBsra/bi317FQcKTXLDaMDYkDbNVw3mhHWajrKK1G88FUhbVw+
MxJjTClcPGvznTKV4oAAOUKr4RxvEPvYU75hnsez48g1YsI7/L0wX1v34pioQZyv
fqe8bJXibWK5DUQ1/iS8kcpgS7Rc/hjyg9022N4a1L0k7JrdbfQ7rrk2xDPW3dvm
DpVWNfNDbvuYKPmp00AqqW19/c04HNI7NlvvSdNDXvp3CxQimqLNSzHaH9kduqDY
VFi75rNXrGNdPayimJI2nyjWui8zZNSlG+42xdz9BCQfFCeLhDlXqghEH8m67q5A
+FJOJD/ihsm0mbco1+FgJjnJpXgsBQoAIgj7BOND6XOpl1O8HZRF4EEm07wuV6Rq
EMGbQtheVN/XuyNIgEOpjxTPuoFEQcQsXU81M0HJxgXYe8DZ6T9t3xnyEnqBzs/P
NvsImyMDSgUrODxZteeIt9BZWX+IOnIMySneS5qTWaiJrZ5dwcolub14hGt17i+L
Cufd0Tuzz0lFkBfYBN9bcaZiZSBMkfCDWW/Ak6ZARptIU1g0tMhCnuwr/cSpQBe6
CK31Ah2vKp9OyCbCkGxyMAhwr+mATG7xK5G89Vdu4343YbZ7zgM/88HyS9sFH0W0
4U5YqiuSYgJsJrZOGlHsT0lDeYvc/q6+JyjNXKstwd/0OsEI+eX5KYwOrHmL9I5V
4ZYdln1BaEx+Re94NoeOcI3fdFTX1jPTlMUwdXsOlPI/W0ej1WmVZiRoiu/vkoQ0
Jkpmf2T8wwZlVSG1ztisxlK4Ww25wpv+vObr4sL61anKhOr2TVD661vGEPKf3r6V
FPXAHjTyIMBAU0MuFQ1ytGVg7fkgoHpzS0V+FB4TNrT5QwESl0c6cYRziMbA5Yub
QpbGC+NO9+olnTIxGaG7osM+JomXgqvcyxcPGMbXJoJUsVpct/da7a8eVfvNnRVR
PTexgUce5wktLeWzzzou6DzqKwFlbLH3z8k6c/8/5ZGi2scQbW0UP69c9GkSQXFH
v2AfHmVwNNw+g175UbXzeioXpILco7yqIPUYlzA/ez8eXm/oqOlYjEJUuQdLmVmk
2kEN38uEZHL0ZPtfQQ+m0RnPJ6NdgKk4ZMMSbJL95KKGqtLAULB8/KDerRAXyRif
edCj/a3BP4wlm6w8KiUQdhgkeBMYk6WwIiYFlaz88X3LSZowh6ZebTg0U39Y3fZn
icPZhApjofNnlTOHBdHF46imNasgxfT4SbDCJRC/4r8lr5MNv7BkjofhzFkYeKWU
g8+RLP0J2UD0s8cG4RdkEQzYgvUlXddItTSM23Xkrk3OtZPAjzEj9YyhyGFvPdip
/S7LHwibeGzO0XUcM8KcNWzBJknJvTfyTBnBjgg2LFU1VFzZWStZDU8uQXsAvAYm
kISCCQ8ZxdTxLlzgND+noC4V+2rHc2s4xAwNj31lKS2g58z/G/UTfhl2Q3t1bMe3
M4jbGY9F+2iCx+aLeqs9wVT1eMwOYTIHq9wLvBWB0gQttIH6o5aHAZ+sUs5FVhn7
biK7HuX/Z3NTNACuAtN4jl0l1hHtyn8kWG+cSPvSWlsHJaE18bYaNKhr1yQCDL5x
gX3g/8q2dekClsfLHkItcPnnYR1i9EBc5GK2NjzM7d3DY1zvw61hQs1sAJkmsRmO
3XHEDzX3JUqCfnUgqcRh6ADvKhBVcrgVhkoDM/9UwHmmTOJHclGLipdjFz2tBhdg
TzyIwVuYXuJZN87JaSpS0ZC3zwwkH4k0AWOYgL/WDOrCUGrEsIbbdfuNpbk8FfKl
rkLO+eq8qmWdzHTgd4dpaZBHnNKhOfYcatglHavzE53J9hLKWDx5hxbaWwCdyZnb
F9WUhrmjZ+yvSWhLzCC9iHRfn6RTsuHs8R2cv1ckhP0Eeo4NNkXLwkkn/33msgFf
govTdJAQJl3X877vRwwn/LErQy/lIPvK4lCkKLoTqO1f7PDiJDyW69gk7U5WEGmf
6r85Cbve36QXfw4KkwF2mBgDzwd69Rk7boSkD1QnkfuBSm4vTUtajXQj7Otl+ObR
cb7LNfgv+kHTgkm4FvkdHfVOU03kqk7jARllNRn28lr/lGSsbGFAzqmLu8IDxiZd
+1VsTOcKNVMFdFaqVYM5zwKd2G4JKPFOaToJ5kbigZgwFxum0Tx/2fvQetAEK9Ao
H2Y2CH0jk+vHLgo4B5P5lMICbGo//18CUggS4JSBuXz4BHHb9RN2qXTfpB0q+zvd
Q03lEb/cHWYLET8bHa8udY2tsJU2QurVdNWl7hKmLgYTGmbfAmG1MJxfUbDcIJtR
xRHFa5fK70IED2tC9QL6ilLPNpdrdmA2m/UwX8oYtvT+yf+4t/Fr0lVUYhux1MXO
v6oy4t6rpkynG+vhDEOdj4sfXWUY7T18oBSE+f3QD3/JXxwqYw8/0WqSfq4VC5cn
2WVtIvqDujQONkmiuuU4VC4FE4EsjRa60TnNempqeuMGiOK1SaBjGcXJxeoM3kms
4tLJdQ5AKigWkiYKgUXo5ZBbYAJaKEgrMsQ9HfP7GuwfBisRLyLXb0HEeyYbiRNB
ElAxidu8IuhDFCVzAp+1AA8EhtlG/Sw3ClT6wgacf+EgUuW8EFh7464dKUsmVoON
scy4hReU4rK695MpqrBZmV7QJXDci0GDkOGhh3o273wqRCM37OkVUGwm/BtROV9L
Jgi/YgIdeOKzwAq5WKPWXdviz19sZxHSGTJ9d1ivep6TFt5c2gkX+a71daoDQK89
Jx/Uvycs98yDp/sARoEejuO3KpCKMihx1nj2SmhSL4u1c7yHrwZ9sbL2pSt6u7SN
6KIsUZrsYw9ViJ3Sac5Aem5XFdVi5dVLa9K1Cqh6quRI3OeWJgw7haPIbMZRgWhI
TrQkuGWbyaj1b9qsN/m7Ql54lmqsynzkj1RQrtLngzq+IKJdCeNvxKTPhXjN6r2r
dB57GrOiTprfVTfF0AWqHXIdsTuwa8StdKfXiOdc17B+LqHMLqddYofG/CaRheRS
p6/EflU1JwEf0RR4zsYjVEfNktc6mUwUSvzpnWErbLxt1b4Encn5VJVlr/XuljmU
5+hmoP38YE/hW3vvO3GpdWClZrkLuBcXs4qm0wGZ0LXGzIyXsE5US0ABHuXZSclQ
p12NP+qSkYTlqcOcCSouJ36Yhc2NP3ybXFnK5F/5APfNr6HH8kiMfq+yLrbhshMb
oPgHNF8HKu6ZOsXXrSy4Eh6/BGGPgkvxexHToDKCXDm59bt2cW3PkkDuRUrsqtmT
3wwqoYuB1gFxmB9XBx7A2sJWu0sVc9ZalP4kegVYU2Cf70ZBjscYUA9+GwUMCdA3
csbMzFhF11RKrXzrE8/ngvHtfxwZ50viKeWHUrtGSkE1kurJJ4PLSaIQtbUo5dYt
++Jw99D4aH4EkXKjBmeOvOthsPgSHH51QqlrM4/dEiAC9f+4lQVr4MaFT76OpU1W
1pF+b3nhgE/3+QjRNajiQyWfK+mBgcPuXcG37VPL8x89dNuSVB2llwE8QtHM6U7+
5uKsfztZ1z05r+m73giNznbvp1nfNY9y+guiDnx2vep18P4RnYVpSzWI4G/o8Pjz
PTseWOsZCIiGmfyR1gxgsS/YyF+pJGmMmpD2oAqj4hoieFNqm/85HU8n/IX+JUlJ
BTHPltzHhaA22B3wqnzgZwZe37W1/uATyy+lc2YiSBatA2kcuGG5yfuQDZUxFv2n
OhQLHi06yAKaAhkfZ60mLrQXAD6HtaOzF2wW1RYUUsD/rpT2RCuXn05DxDuL4deD
mWZeZ2nnvM6y/39XxBTVrabe8Mx3cIpT5OFVYjr5E1C3IrTfWZFi1Nsb2PcqLOjM
icRM9DVE+bEmZ46FI6mti4l67WOonThoSHcGpeQ7CL9rDliD7GLF1gEV4fD5VO9S
GJVXGvvOC/KK5jZ+Po3VfTJ7Nb+xGPKpmD0HMTYx8J2eVQvPvSYa/F8QX8E2QQXs
pC2ybxlH/IbsTeH3sv/qf7eoSjBh0ItAgp6r7okMIwO9bLH6rset+wyWOyvBgthJ
o5uSNz0YV5LuCXRxfhQyP7Br91HWlttpSPgJ19AfU3ehGBbmz6cfY7RlMCc0EqX2
hlJ6EseN4NKKjWnCaWwsV8U2KuNMuArGO25V9lS4ojFKLCG2NQXpeKG1ts7louKI
zJfLXvnILJvUzz02AJWa4dXQnOsfwVEu+R6YlthZV7RquaM9DwhWd4PGDRxPBszr
uwcNFq9FQcoyx/HSUy2vIg4nus1R4K3XVGNrwAD4+xJTWH7zmrt0ot/gQdso07UJ
7XNr2XRlfs0tkyX6GqxLCynbyHJpAApUoXO+30rjuIe/remiH7XXpr8bpNQW/OiI
TaHcoabCiNPsWLmk79bgmne2Y4OsVVQBfP0M5t2VSvZAQM0ncXdXmY7dHFYBgmtD
ikuSrePsi4u6swGk0GEH6NmB//S50u42hxgQSgWF4okLWuOgpwP+omD9naHl4QaE
WROYDmw4nAANO0ivzyStsITUdNAljslZAl6vfTr7zzMAu/ks/pgQr9wekUPPMHUa
UT7xis+3krF/SKIHac4m19oyAis4wSHutfxcChPGVOsenLOpJFa18YjvAuTzO29i
8loJEf+0JDULJKvR3fMVCGvu6siJHiCOnQrN3BOdgF64DmbPKiy2KIk+cThrEwL7
kacd9ckbI1vMF7r/qbmheAHrSp5a46ELPzree22wVdpKiy4ooiNe1iqyTwdEgc3r
6Auyi0FwDhUODMECM+LmUeoa6yesFso24VlKVRhW1UJYpsF+IFetAc+/hGMaUhIJ
3zJ2CJxrm5l9FKYGTUEWQE71S5yZg/9vWj7sdj+1zaeB5gZ57+tYo6sHZxb2UDsF
gVm8E+9M4otgvl0A2j8WGNK1UjWlq9FIXkWxewGBrDKfvZjsjKmW+0VRnljY1BEp
22Ac61nCOHFn7RCTKBbLF1WH6EFdOlhrjRsuxGJFUf5Gfc6Fg+ZcKZWax2lmFo2T
UTls9KrLPtRayZkbL4/os+mtbvSiW5AOQamymuIK8NbMVzjm62qWIBgYuED037JA
//XwlNp30OskD9Dw6ZpPp54flGiTzOW2+i1y5avRCGrv0xP/zveCLgv0Nd3TuiHW
WpXeXZIWyvUXAxqWHgjXfrisZRVZ7Gxgv2WRG/lSs5bnOs5scSHgKKLGCjXsWUMW
gy0yV8921bIRP/h2h5NvVfcGzgMPBjK6zlk3cjwYEGyJ9Iknlnpqg+/bIHlp+Ihc
p9P3z3qSPFPmnWPuWom1H6PLCUXrRAFQjXLz9ZlhWjsyA7ReLz7mVN+TpQ6o+n+b
uoDcle5IXUKAaHqINF4vTCHB8pU6+2glbwWfNGSb3f0YFtMZ+JyYSINLlRXg16JI
bGjuQ39UfENJXlu5bboLN15kvo3pmF/2MGF2biAak68Spv0Y1vR0+a3EO+kzAzB7
9MAKMxPAuGWjgW9+e9tgABqP88N21Nocx01dvnRnT7Ghzb/dCtIVbvhR0Jme+sxT
2nL7eI0+2qUOfzqNqa7R5LuXZw5Qbf8sPnOPBoxdttR7LkhVN1Km4UiUDM64jRI+
0LmNYYpbLSL6c44KOOyF29QvkMQHM2+ip3latV2qvA/1vUDi2LKbGbIZD7ns+M/m
czZbEg5XTwMZWhYJd2wQ1ft9UPLKA645F4i9cK02KQsJX9DQcBSneh+WO9zTgSKB
iq7x+v+ODId0I/vfiMssPtg4bHkvRn1wfS3R6ut2G5AmzEy7V7p1ZSEQjAADRncF
GNgTeAK2UoStfw6HMmcihGIylR+B8gc4LpGJIXcuV+sn/NLwiYFdxpMY2RISpHem
fi7ClmQjn3EV2vrrYJ3prwsgq5bt94PMcLpouEWD7OSniaH7VgFK89o9i9+K2/d3
f93LGIqFQ0JlS3Mc+xtUo/70FycwAUcNP4lYGX7vQn+66WMpvJkltQ7pHzZ5foRA
UNzUvXJCQPGRFS+1t9DLdHIwFB8Y6qwL7gn7wzK3sN+dtMr4XRVE4ThZ0m3O75Oi
Uvjp2SeDJ56z+uGwgS2M3lc4+H6mCuJ8+BjSE6uemMUd2F0SWNxROVa2vxl7DE4V
xmgCKXZXETkT3SLjo8xW2tbTqFb9PFBob3pJbOw2IyQ0yuRNpXnVjr6x9xRx/xXr
OVgEn+WZbhynbBxk3YB7IM2y7H8t8s7MMEYzCeqLST/mfbe9LRuz7doeAOR12AZT
ocLbsisgK+y3DRSmpyqh3vzyjOUpUaJkkWE5jLuycssXZJz86ZWgT/vW9riADJYV
bY2CeTcRD0VqW9NFjBlqfnsCFdHrtLXyNphl22mWwVXTBvaUT5aOAYm2X2rfHr8p
aGcbQHS9f9jKrHZR9lvFEQWZZ/8kaXr1YExG+giXjpuVjc3llay6K82UDa1ss6LS
o20hJVrO9w/tLZyie4dlFjkUQrEQvA/BFwO/UtApej5dDdjJSKDnODitgF6xRS3B
V78CPuf/oKx535X6QKNPN078qTxEAIuXUdPn/5hKUiQ14N+7t2HyR9s7NgbYF5xy
FF3zb45uUYFWxqjPl3WAuGjqCzhoUn74n6mbB9EDFZ3G94mxiECkVypxfKggeSRA
6SaIOqe2l3nTKXq/4RKnPre429k2Owi+AQ+RLDZv2OLHSkvvgMeGWONClPA77251
uEFLBnwgBO5593A7RyvN+0Uvy19RJ5WnK8rlR47W+1ei6zHFP+8t22x3N93HFz8w
qHNF/U1r7wtGiGJBkYOou/cHrIb+V4pfGASfeNiO0am/V1nCybf6TXLcdF5BBgvC
i8FBKnpjMZOOzUmrV9eGdTrgUCqBDK8zOfwFdWKzdbnIS6sLCzzQ64TZs2He4CtD
CcpIrxvp1OYbUDXjNpAgAVA8sL9NRoQ4lJs4Rywht8zOk1iRV6L/1v2ZFBlzPSuE
XqLmFjz/WtjGO7hkJ3OLz/Eo6beL/DL8BHlwQ9Lau7mrape64j1cq8KKMrgC17uL
8kxdbsUxV2Bk/iE0BLlvqc2QBQaNIT54xMYRZN1cBIsG/wvN9e+kZPkf1zXEe6Cx
25WSxL504YDiRPLxCdS9J2CjupWubLQcu1eGDOogXLwitUdY9UN63P1Vrb8PSOQl
nGP0ehUkmOqN1OBxBz0boy1y7c8UW5WNY9Sr3wxqRxFTNtBWRfEzhEv8R58LI+U0
5eWVrKdCHJDSVKM3eO8PyTNBfRB+LX2N+9/p8BmJO7Jp69CgrBnTI7noac8xOcI8
6PDD6FdsoW+d57YXqCnE6/xmzw7VClHEy73isKvF+vuToHyuEIYO9RJOjodIVK84
dCv0R6mHl6clsuA96zr4tUXMSYAJ6ca6osAChZPeC2TwK89/pSjyKU3ru/qi5Ctm
gcuGrZmCLE/regSq5pJQ07jIcopQ6s4ba+f1GKJcK01TOwsYDOQRSYvRwFc9dY3K
KTz7N50rkSX0D+MmAM6RxQDQtOKKUXTdhmsd4aZ7EBV1L9FuDjxhpoqjB2BnspZ0
wX+t3tHH27ZxPjfInyW7WzgnAPclGrjW+BxAJEA195zVb/uK+UPXesYzoow4DECt
Hzfa1BK6eX2cgZtkNxMrreRbr3HVCRpXYqlHjhbOcFjENE68Zn5Pakf1lGtvU1DH
3nXcpZXlGvrlnO1LiSe30wmZv2io3lW8GZ/Fl2UGcTyRfVc2NGvAF7YWNC82ZvG7
JkZleS0IeuzUNflO0Kb46kH3ZtQ4oc8uOv6S/JtReGKoyhTBYEDOSf0ZubBie3wG
tor7U5ttXCotvtVRwGXggKaXjLbAzGGmPARDligYp3q9fQwqDUTWTQvwHjcKnQ/v
WufvBYViMQwpyHqoyNobBK/oijqeuQBG89iBuC5QlrxGUbgTguxnsiungGanrnSS
ABUYC2ARbkFP/qDEo4YOpcMEXmWP8K/L24bB37ZAz7S1uh/sd9heItwhy02ifz3T
UKYY3RvzvQuhSCbMDtJF+PiKU92/Y2i/Ufs2wQE6WZ1trd4AIHQvq9eLq1yXpXIP
y7FRv2rY/81KlquYhHPHtIsGOEKbQlwRPSWl3QH9vdfjunxm+3x1okvWNxEi9J4s
Ho8lytj/GFTgQIsGEw131DQSoKAWWhIIXw8QVl3Gy3KSkutx34xrwm0v6VgOf4Tm
ZU6V5Zk5xY3NWqID/7/Ff1I/P9JoHSA3XXwFOTWfBJpRTuIt/0Y3DcDMd1CSSuii
R/9wc4iJGwAoM0+9aL5u3hqE32Z8RVQCq+tllm1ofDjcCY2Fx60+MqP9sfoL3vp0
qlXGDoLRh8iw+CT14nexomu219nW3Og4JsX5Q84SpZCO2QNxXbG+boJokoYhWVSQ
2Vwru2eKkXogt3F6FEos9mIf+ZyW56zliuv3IzsgbDXB57+OTPxv1+gQPYId0+VX
46Vqf4etYVnp8qDDWy8520NrFH8gR8CeiwIaI9R/nY0AepcoW1rSBJs5J7DZUCaO
Eyb00I8uxVVRbfGfg3+mI51WQ/LMIWzMFTFYSXj1dNZ1NSnjCB7uxZeB0qJj7bQx
KuqEp9E2SRnFh7unYgCGCqaZyBNUICZT4yofTZrqmKdDhZgfKENKSLmleciiMS6b
UmHOGKqgtOKo89Q7xFfJ5jR33goLqsvyG3zVb0o6Xx6GiBJuYsm0qHA+iSyZVn/k
vyk498YKjZZa8aSKh1YdWhn8lWOD9QV1TAWGOfsRGT2UsYMMT2xsE7X1qKfWm22N
3va/lbCGzXyFc4vDSxEGMoY/360RtF9I2GLh1kEu41FsnNviVaZ0GkB0NJnA4rCF
10mR2zkT3fSJ6ID5ATl+P2Fuw1XW5SEfCPbCEsY453TXYgDAIPWu76B1gelx9Xl3
yfJtbONLkhHBUleegrLgHZk2iiPBArsD7jgsoQCioqlZFTx/ryJ7jFzwGQpSKtoh
T5XIazCu9OVDO928diWE0ZJxIopnzRWv567a6Pq0/gN5m2ZpG00ZtnRlgn/eyp4z
RhLhRFiHvosZSeUoKb1lxZGbVZgL2X/Wih4ZEvzFctkYdxkX1FGaGv7BbSFg1bWv
lz1xfxsFKSmKeQZ19MAwvdxDpjLFWkRP2MgNrfJ+Vng1GPT1nuk/UpIMZDWNOGDx
0R9srA0OzfV+uUcjP/pWwtEznoM4BxzlelGoeSnPoh/ub6+xZWbeNbWa+AXQDh3q
ABNziLqdTYFoyqJQPOpjuchOLFrRLakobe3UoHeX94ekxiiaMYIdxsvqo5Ml/3ow
r/swSfiyxs++/y3DuGSPHQa4LFpScNrNadEDcy8BDojx+oecn2lr0Ro/wxDCLddY
lR4kCKVZL85LPyoJ30D+3Zx/JmPOTRrA1BoCyFYREhJWezmEv1kK3/mE2kdqdPcr
HZmBif16vClqigvswfmCKlYqUyUVIfM7mWzXjOpHiblJvpZnxEZGRNqw/S1JWio2
j85Hso5eS8gZrpsbLhIQKjrppoIefYqKrRLRddQaCJoOIb9qQMUn1xV1TGZG8ZsN
CcG9dEG6I80GSRxIscEcj8mPx+xtt16kFU0C1ecKbBTQw3vtHmvvVQU8lF0Nr/GA
AHH7jrbPgDZkvfaLQWPgTN9P8L5T/wcu9dLN9B+PclrmVCtJkOHUv4SQR2MDs1X4
KKWpmqZetMukqQwccjo5OZGNFQuSG1KYHd/YZIbP+uYC3MFwX4KMAu2Ma9ODxIih
7SeiO72MVavbTafUJmy1o5HlYfjPsaYaBB9z7wdtjRL+xXvyMD9go4ccv2eUlHhD
6ngwOAGImoJUSj5C4RvhdHS6eKntvioet/JeTYkJ00H3QcEWSUfWAuvI4Arqpkou
d84zLuYPiGhpp8ZjUt7B/02MANAGssunFMngRcWgFxgUua4viP6QVbyP+JwWyBJo
XSQuRzfZrP/pToOpNeC4U2z0OL8sSZ7U5B9h3eEVyor2ow9qulwUJO4BsA2drKUw
goCkqhPZA0Mk1mgiIeY8yN6Cat3byibUUqE9EovCrTptNlvU8DwMAD4LY34JYo2w
MqORWzq7VxLyT7kynHm8PwtWLn0P5h92IlyzZs4sKVeWy3jW70E26kRK6bgUghu/
4xtUmX6SzuqFYi3AC4iI3C3CT17B9z0GqHnfsUDdHYFFTZbv5/tAzclK52kKtjmA
HMklhIaz/XYEKeiNPe9xOEuNeP1cZWZo9PPe1mphtHVi2NGarlqXE0BUrx1YEQdS
G/NObaYDgw3rbq4pBleleGEtCzK34kAkF5ytSczemJh3KDaF7VATp92striLYFVe
uEopd7IvAgAs7BKsSlFYll7e0IPG8v4RYl4jZIUHxtwRr3hLNhJgCv6a8CoaPlnc
SiialOGSVDjbpQ3SFRmbYXHc9NJZnyqHhDqOMUapFQRZ7TlBTVC8ZVbgKPbipPSE
Ev81gGqRAA4bPvBnkYDFRA0qykK5DfPabjxJF8L5IOfMKkywtIp6W47tNjybyDn2
9VPsgq4orqRa/QTtuAMlLv8biHdL3ubMFKCZFkiNx/tRU3DMepyu8vAly4AcTqQD
mS9MOzte7nLecDxpj/4y2IaekLgB+xPB+0a5YmTgJsejVl6HrCgfwJH/NRHL8EbU
264DFP/uWRNGyrNrx5/X4c9p9+yOfny4tDxZZC30HZMHLTGdZKgaNOv5Q504pA6A
kRbO+mwvscMsg3Cs2PjqPrD8Z1Wv3QP+zLwhsx6yuWFld7RAzYnwx31SlmHWkPex
KZ/Fl7xryMScCzIFR75NsmxsSU13AJmAJX6Z2MNha2dcuqkGcpuw/Il2qCazjxFE
Onlp0zx+LSYcEZ14sFmTp72B8cxrdDetTCub7Z55rnxwDiELC59FofuSVKExBY5O
Nt4eOHKz5/dbfAWXOxXCVxGeACZx7IJt1YQI0qpcpspYC7qD/MQj72IRLkSKf0ZL
wG6iJjPF/Db5U7+S8fj4N+wyaUTGZCo175wbsqPfzsPGPLkeFBpdd2iUyGEM3dKo
rUaCWuG+0QXsS+0nSkf+zLzVPV9efahDSmeS7cbJ5biCbctk/jlPQbxf55N37zU8
ZfnA7jwAH18+NxGUqkm2lTYmUTp2wATowiGjG42F5n0hlW6zgyuVi62eAALWayQ0
90asFVG+9cLe88KVMlhXL/vfNlE44N8RrMgPCRjMeR8x/fbqPHpfqjq8UzIZqa7B
dAyyjQZvwx4TL17yWrhockpOVGmutBGCX8UV0nO2C/1lxI7pJnsAZna18U5s5gm7
TvBxYoCCioYrH0l5gYhFg6IR8bpuEDcxtMBEXizLiaIAmvffyk9KXitcHHDkMIkw
TPRyLniuEQ8Ea/75LBD1zFLNp2YshJ7+UZrTt4qUeUpn/hkVAACkKW1ozTMPrp/M
HGdhnDn93+BOJB1tweQiUuQ2qZ9emuU7TB3559BLADJHgzc6i7IrMz51dPpAFPWb
Ubwri9VSh3YCYiBbumOU3EkrxUxz7BEOGz3WvKHexUSwchiGwiPFVcRY6/kzZ/DW
vKaicbVHv5jyDSApVvAe12YUMFKzrXqJ1VwUBOP64Bt00sxe7uGBX9I7WkGhLswl
VlgGbCLavXDcIx+PdkUre+baGfvHly3PybTvNvG9W9yiNwu9lUgj1EL2Ej/BKsQq
NcOuGKr+1V7UxW+wJmaJ1+eu3qcwTNZgfWR8wi9k7s5vJZQ9AOOqpaJpD7RqYzwN
z4tVmCrb1pzGJwzkHJ8gkX6526QOfLMkoHsksW8BmRfSkPYs1fwiq2bUABAT4wvJ
3bzKPr8XElgS/+s46Saf2ILc1iYrPze7NlC/3nHHBQvlb6Ngja+U4R4wseeyQuXw
tSG825/HQOzM9a1qsyU9oYz4GNLI9g4Vy5A18uLzv0ne4vGo0n7Q2XjK5dz7gCxp
aeUxQyFKcJQyoP6jBsdiCceSdHhDsh6oKyThdVoIF4lF+9bQ3lj27Zz1pQVts4hX
jEBmzh2YK0Ql9kncXJ8B9XIXhsPwU6fSm9DnoTKE7pGqSHBZbIIinV3gS3Xs/q6M
ax8pGAKVW4VoqTOq45v8u9G6YnsL/QFsru/AzVPheQDzORlZTOs8fAvCeBc7RGTi
DM6zZ6IUZwrTjgpb2nWeLudIYje2hvUuzSqh0KckGF2Omv+gUNbiPNVda6/S8zsJ
ymZeLQLmlmpgGj6VeLKCHqp23VpmhEYznxWeaGMwCqZ4jtnODI9hm61spVDG3jEx
RylcR6gE//+yzScwCboRMZsn2W0G4AYvw3iZdk99cpix+gUGS/RL+Z0YH0zuH5Mp
CLinXkFY+1rFngEu+KWyFnpeJD1pkJLptb+vvw0a4XwC2l4vEPVUnxzefTKMo9kZ
0sMZ0uQUVWixZCbBYtXikoP34GVWV7cEQQI+U24p+KWXv4RLT3DKHLYBo4WdARgZ
ynsccZaRfiQPyYjPBAF1P8lwlM+ERfDHoWZV5gDVBhoNvde3j0onw2OVDt6TUI7z
NXNe/VB1LchqvAekbQs/013S2xurIUa+n0ekEoWeuxxLG2sNJcpk2CQnDjWjD1Wm
w4pG9N1985z5kolxSD33J0qqjN/8nilenCp6Qa9kwLy0NQ8RyW3eaRul8HEnLSKU
un+bVZx60ys4adSkfzyqz0pSLRxMJER2oW/jOOpBo56QaTlueo1zOcnuWK5MW7Qc
femc1SEgznnvy4NhP0IybgYUtEIBHDbYJExUiI1A+FVqhuNojNdo40raCYSARp19
30yVZ5u1IgDmXh5Tb2ZuOmoexeGEpCEHIhJ22tEEPTydqHz+XKuK7LEvgumF8qXh
65zhXrA3MPcUplJXbsViSZ3gOzs1eoYI6hUzeaUICD+0Tl0goOoNvOytpufwV7P8
3R4PI9RobaO/3wHqGX2NomSgbJFZvk+KSyRogLHnYczogyt+6zGxBSkcY/d50vev
gMh6rzbv6cJRcX0PzTqVt09Q0mYVxl6ikMtn5ydwBcHBFn3ySs4Ie9OINT8Jshnj
ru+nRHBVmypfkscQV/onK3QCSot7Gb/RWns+IPD6aNYVBkoQh9BkyNIU2At0v0Ml
K2DjHTZ7unI01mzVDzJ/Ml80Lxd2AXKXRNJ7IXkvzLBUZAZ8F7g/uGtRszPHG+ZG
2T4XnoO8MgQiW3at0xcgsmVPSzcnql78jpIsBdBourKWOJs2ikXxQf5gp70qtCwH
RSI3n2viHqQG7kpqoBgteqcHDJf7cQjrImX8iBu5xl16BxFcQ0PwrM1pV/e2OJfX
ZVzZVIz7cqzn+fwCnDPfAYQJentBQB6r7t9X2R2QaPufNFzxnKQOApbhR9xwkgQR
flte9jMo2l8IDCjDZhvReE56mmYA7Z+uxq501OdoGBWtCNBGRmOU5HiDRbg7CoUw
KsD9r4KtnjbzOC9IJdDrMpE4cGHUtBgxlKqboW3VE+qv29eiH+oayCefI0mPbUm0
zb/fp3QIGBS8e6P/bRQ2uoLAHDWQmlMChTWSJ+A7SO4zHCMN3PPwNECNe1+3oJ+c
zv6Dg+rZYgTJ7ZQwKZ+b5FTM3qsW42wxjtkzQFH0oQlnFSstNclNGKVtEj9k2FGz
lqzRFhajbR+df2lysK3HgwRClwW+TpwV9OR7JgzbPJG61/2T7e8/ffmvwr/Kpa6E
ISrnECXK8gR7A8HpLVhf3NiU+ua7WtDCabmaJrEzmpngdOjhC8pxGoTBgaeV77xw
tE/EzR+ARiKJWKOb67wZ2TAOm3HmY9t29LoANwDiJNc151h9iptBMd0bb6fPW1+h
e9lawN8psQ4e3sFWPOqvlfr06T00HcBTNZ2Z8b6rMd8ebvva9jrk+X58O6HjTpdf
Wjimwft46+IP9jH3wHnpaQZIY57SizGWigO8z7DvFY+6EZ/QmLIclYyDBtxRiVzF
dkO2zfufj+fvBGahBf223TMknvnXyeDkvXOO8rRRiGMs+xOQRdUvuLgk9n0wAYzC
FWRTgiBEoGX1CV2YFqPMSWzgcCT7coRtSGGGLAPOHSqKY0I0OsxO/BNhig/YEYaP
B1oF9ijzx7uX4VskOKg/fZv5cHfIPWhD1Up42VRvRCC/ZgmfynQBRIkV4MVDMtMH
UFheJzih48jJ45sgaYCveDloMu9Zf8E+u8Yxv6gQLxkK5u9HMp9Hvg2f9hfxq/UA
n4iQozncU7nKV+Fz2dvY5I33n+zoNb8ExXBNhGqe92K+WwN/k8Gsp3pv0yuF8RY8
WJ8/zhbCAP3AjqvFblK6a7QQfDBCnZeM3d9JZWYIkOP92qcAhaZiAJXlw3CzY5JO
UzMqTcPXa+h+Gg2mqCgbZ6Wjm8RiZhkdMHQyasYIi38glD7eV231iOBc9c4uwK5P
11sLM2Ad5+6j7n19mqI2+kLvk7qsIijFJr0ZKu0Hc94FnZmIs1RACcLoXnga4Kfw
94dxBYUm8FL6YFb99JkQ4ucB259lg7zkD/f4/O3B/MtybBGt9Rq6W3AVx4Uoi6Zy
cVE7GjJTDsOsQsO+DREbIFnLCSPV55hZn/fsGkG6v+fKa1PfvwojW/DY5RQ6dnQk
r3KGdWQAzoXrR6svciG7SH9zK0mPXep3yqqAuWTt1N6GV9QA9uDfLZ/TyIAdS70x
DKVfeL7aWImGQ/uhiUJ5RJdTgmBtLX0v7zRS8KDDllqRQCMSRaxMF3yP49U1SttW
jaSXuk2K8byWGosFme2n/57mxaTWexMw7+DDuIvG8CTBIyirnqyrYyMdCRF3q9DB
xY4PuTvHgnaKQFICIpIhUt37VdkR3vUcD1H6Ks/fvEaE2/6CJcq0CIQiU3btGs3h
fJhMeqe6f5aOiVO0ib3x4w5jE4I7SjiZ4csg4UobCVAi0CeEmHAu58TU6aR82Pqn
WjKltz3txCNZayJI8azwcPPtyiLY0CezCNRkM8XZuSmC5Ya/OQ8oEiGwjznOXX6X
a8nyP2cPvg/FhOLNy/YD0dmH3mwU2Ry+aiDzl+G+HilwERF+qW37BANr0+GqulDu
ISaJDz2euQagJ/EH5+2/QtIyJhcUzB6jadiapFYyn6YYlSD7HOpVyPnt8dgf6nXd
D2tSlfUb0fUGvBwrzkP/S0kDXuIULlJRuA8rsF6GLSmAUzOkktYwtJRXVrwSaAoh
St13ghzsrhFfen4gshognTjQGgG5hN3gKgdVndIjBX2kjiEa+1kpTXk0O1f3+qSX
pG3sUaFl3apfHx0rgE7OaHR/DVGtwsYhuao1EhQmWHp/Y8tBJ7o9mLRyGij1UYWo
CjGWQBU1AtX4fBihtfrRMg6Yrw3bE5iR6L5cLsXIv5Im1bUYAJ7n1WgyXva940o+
VzFZmZqPjUy07aB+LFW6KQgmCZqavzj5afIlGuM2Tr8TPyXn4p95fxrMSDESd4jt
BwORKzJVU19kDCJgwc7lp8NV/WXkiAME6m0C6vjvZmIwGU4LqfM2vvQgxezEeZJ6
MoxRLjU7MDug9LuGQoicUic+nX8H+AmbZ6RlhemVV9FIKmjcSKjxhLqvwAG2XimY
HvqYHgfD2P6Z88mZOG5pkrlllipJS253fMFL2Ch5GbUAN1IXsab8DcnGF7XeoaKz
Keyb3I72JOHU0ahDiAHKMQQZg1ztR6T0qqvuaWBOEPhOvUGlLBUL0Iu/aodGUa/u
QabIvFqSqeHb+ah5oXbDNhQK4nMGKBoHBguOun2l0hg54IVcl0GPZhCUFaOjSS45
I9nRQJj2Z1YCbF/9MfJeQiiZ9DFLCfZ4PDCufqvGaoPz+PuTNGxX4c3Y+gv1A8vd
oN8N79FEqKel46mWxXBM8foP2wW8yhlLv96W0wte/WlaakNyjTFUGPXGV0uqIC1Z
nEX/oLVD+hpfdJrHVwX8tSxGgV6jwFmGxa5Aq9kfPK1tPw+9TT/Ewc9vptadZtUP
zZDXCHXEEBI+iZorOMbiwBy9gJ9HdwlkDvwAw/hbY1FcJmvjncozpVBk2Juvzk4v
f0aRaphh4WRYawEd1OffAszZQTr7dMYcSDUkj488m0Rt4hWKjS6DlgKBkfh4eIvx
fe/t/rFcYr3fv7gNWFJn8P0wrJtSkNV4a5TNTzOPseuCsdHkjqC7y5ngC2TvXBCT
JlXwQ+F4CuAB6qgGJyn/bvP+fe24nZCJiJ3V2y1Qo8P+MRGj4r7qa5YgqoVc2Rqa
0HuPMz44NXRdbfqVNnWgNzyEKSfXYKd0U1XE9pgogYizOdKpTJpduCAL4FhcbX6Z
DQZPQ21U6kzdMXRPEItZPFH6xOKde9D+iWf0q4cy4vHJVg+/gsq1zXprHTH6KLO7
8MjQqTGr8DWBML7Npm36WnhU5ozE0hVpxPOAkmaKJ1bcW25gY54o5Ubqu4vl14SA
LEHVfYuIUegLZIigjp8vID9Rn4bMar4BJN0X/OofxveyiY2d3m4wq+J3oJMBMjXo
dLMySW5AvnXPl2qnzTMSFZCy0RBxUHjAJHKFRRMp789COp2b4d70NrNf/0UKVAJt
B2NDNfLTBLM1eI2E1jba7J0j84IZnuBqGGHX0GK59LS6Wot/LEBw2F6xEaX4c0JW
Io6rgY81mBqRcgCQBuhwfRePPhAKPL3NS7Afi3RO0K/gWS0+x/ryV39r0Om/7/T3
FOxZyTmBr+N0nGWGhbhI3EhCd6ohC0UdBHjyj50ICJD/espj8/XqLrieXbzLM/mL
/5nT6TIytIqbbLM0uDzevUhNZ9PSx7bmqlQCIOWz5asMwa2jidccD0oCbVm1wHWU
0nqY/QJQheIsYRrOIj0GRiGLOeYXI1jZEQas6pD/5/3pfnePw9/+GrY1/q2RMc8o
Arf0rrIHjS47C/fM95MUagBkT90wX2HejAThZM0NoljUfZp9AfA5Y9w4Qd64/u1L
YWYNhrbrDqq24kKHvL5q+aVH2v+cR0DtfE71cB479vGo+JLWIOiaa2lTKZD/RJre
RLJbr9k6wARG8nISDk5b6nqpm1LJVLuuUCBpMB4SiqvvmLwLf/ezK68vZRi+fHRc
8AJkDvPfoIEjrMIEVV5kwY9io8XQDG2uPMAEdSXX/5kXHAKS6aJXeJ5ByKKzeQk6
yehYEJE4jKpZ+G8aQ6EXqC5/+BLP2NcUHTlGuc8sU6XtylcAGIQyLwlmXQtqbLtQ
Nt2zWqX+SbSaXB9LhMnIhwxUgJTnXwVKG0tP2ar98OX88BCAqjWM13Gtvdk5IRpE
HCSYw9Ak+SwnCz4Ze+mvbQu8/IuQpCywWHVuFTcRn6VOZIBAW+WCwe/s/M+DzrMX
RhE2jnY0Fs9HM1O01SaSvsv67YgxA3jmT/pF/tXkJWOVnJRNRRQRJrypM9hTfaha
fqPHEsitATHRYGGlKynHXM2cSO8qySoyZ5zgOW6XQzZJqlAwh06vbCwg0Aq03aNi
04eZpZEAODCQwBZC60tjtSVwthcuWVGv22rzrvAjg/Gqdjvk7e7rfUQsxURFCLBR
cWSW4YNA/N+8OQoWF7jPMv2CmQ2MDinElvc8nhVWk+pnQtXKOVWlYaQER+OaLsBo
gir//pFP7F66UzF0t/nG5vAflhvhD5R6XsuEZQ75lYSD0pKQuLIQxLzY2OqQTI3M
+25Xd0t5plqHa2mF4XmyrETKlV9qN+7VdHPEnvFlkIHcCEgbhwfQfROAeI5VFlIK
yDEIRZfp5SGHsj+5FQm0wY+2S0FOEOynQuyt2NCE79hNPM8p+NnhKs/gKESinXXG
pp9MqNG+tJV9kcY5E+ZxfO/jXT7Imux/9/n/iykYpJD0eV1KnT3IcJRmNX+rYwmH
Kthb5bQWiPCtR3Tcyh+SshTvzTavJtLdUA6z/KBmitp+Btk01C5skXKAoNwXqqqJ
EU1pydKP7nqyhjEwIhyk+p9Xj77Ly9S7THzy3BgXwFTViE3g6b970X1F20ss8nGK
ao3hv0GiOtdJurcpw5QYXglaiFHjaYDI9ryz8Fp/d7+TmYrmy2t43VvI7HQxnGkJ
VmMlxCZ80HsWaRMx35LeEw0sT9MiX2nXA3VSe79EI3pnPPaZKRqf0XDSoNCz/V76
lFVfZWL4qSJwrbgAHBz3TnlObIzFrfAk36A2pth1W43lsH3Fte0pjsQ6g1YVB3Cy
qQV0z4zdVNROuSc71Est8vXZZQRCEpKckFr1KBKb8LiX/BqrTmJhOYjkxxvbd6KT
GhTTGqWgEJOnkXpLL7G5lrKoDb16DPtubh6wM4vv1c7+pu0SyGg60zyWwE+KGQnx
3EdYHK8pG1mbjQ616kwJ0CfKm6YW/C/ln1U8bKPGMRick+WFfEkJhWmT0+nEtju5
k0rbCvhouPFwxXkax3aOiE/T+qRuTub6WbrslopYYzWyylw+6O1sqzbLO7puikK7
h2AagtZiXCr/0/f9+LNLJK8b3jHIKje8uYNc38mspnRoYmF7IKZq7tTcbNF1NgYK
LOTWMGdNavWe6Nrzn6HsyyRj9K7yM841yOiWUg7HRRSCTXWNgNoDxcHtBvVbnNIV
Nw9/pYMdegARbYi7DNLamGfH62DqH93/HGXX7QvhOPkFm68BI5WjVMv8hae+VU+b
f+JYTyPpPgwEUIhqudpjq2PCzb6SepGhcq8vOA3xL5DErR+172u2QBWwW+bsxVRZ
LsNB0sg0SeC7Xuv9bxATiUe2Yq7EIv/ssBXHadqO/pSeYet04aInsAgSGlMFDbBU
TyxiczPkSjradLg7q1LncTWya4tQ1HoLuiAFuHtkuXt7Ioqc8LOu+ZJMkPajxVCD
jWhNpGaJFzdpoYpzRK6RF0AENTM4uaJIFFyECvMvDjoUivunNkilvd83nFPVNc6P
V4xsyHdJFoWqPrPeCy1p58EaN4R6QRiwC/RqDCEJg2c/CQdp/P2+xiA0UVlWyCXM
CYv6cpads9hdGexMGEyKUziLcdZvzAkfNIpt/2gesaxh/y+p44tnSB0uQY/aPIW6
YBtzlNWqyWy6Jch1/rsabc5P+QWaWZH2CyQcMtou9hKMdaVfm3O1aGx99FybKx4G
9//WS30km1CtRpGoy2kNGicKYDl4AjEIS6JqXqlH8znDpIGF/Hyz/qDuV7WS1dqm
V0MNsquet48rWXkWbDYYsoGwnl5JDr3zI0uPezeFEaKB8F/0DAejlJAuMFo9787o
irW6Cp/e9tlxd8BQxv75hgGvRq3F7adOl7L7H/q+M0P9UhWJJC9ibKAC78Jsqb5h
kZrsVYqIVocuBhmOsg+7cSOQ7RVNrTRaV7QM9MWJ1qqM9Y92VWsa5AK5zPMU0Wit
JGXJb+Y72wFsQOiiC2vzan6S5jmcm3ubsQcKrRbg8EgRyW5SY3r1hCt8b1aCa0n5
WjFw1KH6xg6EVBcP3fb9J4h2hbJsMgimgbnYrHernfpLvV8TdWezm+rlKLPZeFel
eqruSYzxSW8xNSHqNDRyvimpYbtvaSaAAoKRy/ckcLKAoqfCXe98kFQwymmmekB5
P1u29vnboY0ZemhaRHuX+1emkyNHKzhl331QZe9hBOg0U6agoTunWFZys3y3kj3Z
+6o/3QJc1iMgxO31Ax2heDYUiNZ+YMfoRbcPpobE0RIyqEXsF26dxlQ7082V2HQL
evkGWNWvrJMM0Zc7+IbOU8MfbX6QKQh5y4Imu5cvWy9apMqmirpyap+Zuq9Sw8ko
QGn8/STbV6u1VyiM7M9JDy9YpoE/fHhpvL+XetGgTt2s71YR9yOk+Sf5ks+fQ3GK
nzUEpydFUYkFEDI2KauVu2Pg7ZgHGxO3yNY3hX7cwHDEeMLrvGEJMvQ3m3H6zxIe
rdyLZxFIpAEC+lHBY8J2XxZAxE6h4rDI31A1ip7mUuNX45RGKNHMZ158Q7+njWvX
MoNvrgzqOzvwitoxl4ZR2pXnv3XK6i8gCl606yzkAk/eM4RH0RY3ntO+oqT+cC9u
YCMQEJcgzokRtKAcSDYkmku+MnOXCrvvYXEADUI6stJQpm1ES9MzarXkLdf3JRh4
NBCkctHDOaO6qzVv3uk927bvInOfTz+XNt72hoqD03OqdU7fPH6rMpGItx8FgkZp
tdg46ytGCqAa6iYNCSfYIZ3hHtxEPmk9ZHKqn3Y4HMpkgpH+cLnu/L61KhaETu4j
3XY6H13Xgqws4ihdKs9lqbPxAoBvUOcU4cPqpxaAUJLo75WtmzvsUMUdJq0XQVgS
elWfdQRaZUiCPGEbX6YUl6uV+iTWPAwmGVkyBHxIbO1WwU3vl+fVaBqmjDzILoa7
veMUbTyfLfJmejy9TiXxO4Yr3XF2bJSkkRfmJoAoBLX11sFgL+/TaiSzyrkWu89H
jH5dqcsOzMCPXXiBgkINa9VdBfzP4yNnGX5h60okmQgniDP7AzqcNXoc9FznIydw
gY8/GngF/yANzLN9Tni71v+kfKxOzCG8srcd9o8B0aXtyYK+lAA18VzAfjhOb/Tp
5PH9GoY1eVQ0/La8cUxXWEE5Xpa64W9qDfR3LQMkGq8nuXqFAF+SsbZhoIdxft14
2iMBAylMrRhLWM/XxDVy9bm9zoXqrRp0xcl7+Wi7p2AD+PUX30+KS6+kc4I1EH/t
eEm76piqDVlMR/CDEHmFsPR5GJiC5fUc8rOh3Y7pbyqMx8Oo/1MU5DK5U8zFTI3u
y7A8b1M9RjUbY0Rh60os2sZrsouTx8pG89+ZQuAwuGj/2d6r6TK+M72/HvHpR+bB
igjF0rfdpqttxE92/GGClqiGgp+oZCQ3AYWA0h08NqHaoT9QPw0i0k0cG2viKTjK
I0uAj/KCMhgGTXX6+FkXp7bKbx7WANtMHB/pdByw/qDssqxiVZpy1t0nSSbKYOSN
YAYBIU7K/rsJz+EE+E8r6NErHkE7RJqXLWjf18tmFPdBHK8MyfrAuSQMJPtZ9JHu
6N08V/ymjCWNiKwlmplf4veFc2UYR3IOyT+qrKJWEqeZyJRSK4Hix6cgIXutjZL8
jsUkC77KyB2S6E2SL/zt5Al3G9meVF00bpoollMRoY7SpwwrGLwudtNrAQCGqY3j
a0R5WWNOaRVXlCCRMVftslyB7GbOMAzqwMA5DioAgpWXGwKwaYta0Eu4QnQiyCxJ
wbUELEUtQin4yfkOUBAdWVKecN38q6KgxBwnk5fu6cFHJ2NYQ50xGIqGrvuD+i4w
oRWVVEZmlYZnJVFFSCJoVrFmjKMXjHgd9k2x5vf6brjbB4xxZ5E7hazcWYTdTiM3
IcUI0feK4QCQK3YyUqrrnmwT1/zO+KdgjIUNiFySQcqpkSTNLb9u2D5ZZtsP3ecP
gUbLBqOnM3ynbDw4EpdJ1chgfpQJV8FiRe2z5rnUVz/dDJZesFu6OVBxygik86xJ
mLDFqDgc/Gt5hj/bUndyMdHDAaM4eFlSM1IdgveiUzPFOFoudsraERoeKOrHOxOu
KaEDT9E54yGGqhsEYh6CfPPmkRwScJgd/IK/7QYnpNigWrFHmsiI83WRYlZjs6Md
K13Zy6h9zlETZ66C7pcFWVLwe9XfV3ii0omeOTDFBqgnjqiXmMfPOKWCzJ1h/ktQ
s9/v9V9LLdu/mCBrDCm3j75Y+dw1UMBuDsYSSmUFfZ3dwtxocA+FhwczMG7bvpsh
8q39Z9JWB5QAiBkvzVnt2YjYVQDcelDcH6UlfXscZ/fNkUuZZu0wNVBy9eVF9sGL
uzipPKsyaUpzgugkN5TaxqpZDZYHUQz9LhxtvVRPkHOn+bO/DrLmsudfnx59FkgC
Al8dVOqZHLMx8JfG+FWzEuXoXM3up28qo6wJ4hXnkGeDzccdgqDEOWBMo6ehL75n
NIvFdXv/1QqZTtyiubZQqFl8nbWnGVS9LDZNWQdb5CxqSY8cJ/iDaYcD03HXfc40
vPVBVRUbPylEIzX2dMLsWiTkpDKETo/FzNqJTt6EjyasMlpyzRW3t6jL4l7rtegz
cgdLr+qUgJV39HEJsPaICaZmN+dzLLOa4140L2YJ0cnqxH/Rl79Jocc8zIQgbsO8
dso57LUS5CNOSkCiUHrihQPLgdryny8B1qg6Q3RUbYunDkteH8UhdhmeMQHvKpTy
wEqhTe806O9krfrtedy7x9yVCKyw6mDXqpZkc/NdGJgAT5Upie21NJKO3sTmin9m
vT3n8wlFfv8TYQk4eae5M2XOay25ywQQ8OVmh/Ic1RykvBnZ92NOmh6LT9aXN3HD
GXl/Jn6pZS6PS/rypDITFOnivfCHpaKrJXR3BRDkvqcnLzlp2wB3WGoZ8IITGsXg
wAreUUwZDW18pvqcHvedTj1tbtav1Ak10JJoMk/SwF2ptbA1w/kfrIbOUHVGzWDo
nnD8AhmJEFQ2JxpR8+cgVquj4RTNaHimjz/Y7+FPg7RQx6LE+Hff5VbLSxlS/1k1
EkgS1Evs5iPH7Vy+97LwGu3C5cYMQNr/Q/N72OnsB6mZrgWys0LUeuaolSjb5Si/
WXhrYQp+6paTbGZDm/1WqCnx6X/z5nAJsxBZ6ogjVco0E3EV50uQeENUjqHIHu6y
3NCaxJJl2nRAp7+puSqwy+zR4MA2aTKfvd8n4n5ZO+zctohER9hSDC7FwUKmyXtt
uwoliuwqrjXJvR8tAgzM5tea3KW9G/zn1+Y9nWJTS0eJ/V0p3yCRhPbLO4J+lI5i
XnQYskE6DrLaZESLGsxcdsFK3KkC0dzTUiM/bJrsy5+A1wpednMU+NNhR9//yGTZ
tiKQXXfoNvjt1MU/Td+C0ixnpwO6TjH8fkZVvwqmSF/MZP9Ddav0/zhCg290DMbS
UpngP+aijTMiRlDAh/QqvITEnnmdk4jgBLS0JkcfEJle/aPRJ87AxgsnHn4XgvNY
l7W7lCZv2zpr+SYbyycD/qTIeJd0Nzn+3ieQbM8PYLcV7TWxuc/6/kiVh5SUSsm8
3A+OSXq7TanKNuCTCizPJKU5R8edU7j38dpFFRin8EAIpMCE+Cz33xNUgQiI24AT
rFNwLZOQ+WekedK9l2Ebwp+ynNvg9ciHBjPxN6UBp+mhekda085aLovtPnTuKCX+
mlAGudLAw/b7gp1sv8ZOvvZAkFVdJJuuJ/mOyDlo8Aa+49+FQ+i0yxvgDLphltoP
+V0S2dfPaWhpLmUv3C7gfGfO9yFWjGhjiRQfJ/6AMKUw1zVd50Bj7Y60PUlMYTxC
gz5eQj3zsJbqPEsCS6mrMmqeEE5dlc/FnO2e14fNW3yklCTzsMl+pfQzCKWYVRo/
cghi0kZ38I5xHZpsC9K7T7I7m2wxCBi4Qv1voOgqb+1TNhrtdFKIuL9GYS7jnPl5
4Z3RTWLPkY/Wv++3gJ8whaMkGNb1Q4uCjF+pl7wR2GO8Lva1enQVH3jGYj7ZBLdw
da9KeLMC9ZhazyXeWyfNeuZw6awsJ6BLz7NkPnd7zPn3egmve8ZktEQb902P5jqJ
HXUVnakjWD3Fg8PtcFyVk1pQd4tbigZgrFEq/RMBJFY6hLF5z00UkX1japUQRHNR
D0knbbG+SZ2Zy16YsBRDkw7n/Voyswgt3m8fTs/cLJfzxS5Fne/MsA6oIbVZMV4f
NvUBfviDNsvmgRNqUdzUG90ei//G2ZPtjPDArMrtPvArIfKQSkyIW4RPpLaVVokT
epR36c+R1zUKqVGeanTi8Ves0lAxnB8U6T9/pvOuP1SbI7cBf1ooBwB97UgPdesj
sqm4NIG8haElORsd9/mHPYnXCKS1vUKBUReI7PFedbzhMX3ZiUwKGZPXZQy6VEgT
ZdiNU1pe5GkYRem3UzPCuqVoPtfsVJDxsG4iKpAoyo6M6qjairkGkgvURgbEhLGH
raCKHih93xUE3bBeGxS3zD2AVFc95WifNDSE01aDspNWAfsA6kTGn7TuhlFaYOpb
9WYMdbyW8keXUnOC18VDXGKu/EDnQNQ5/7MV0x2NcXu7jb3vKpeRxnUnXY45e0LW
AXJCd8xj5jwv1URfIyYOWV12IEM8fWzQKAB6HPZYR/WJUcpGPiOwItDDPu2o0myk
e/1WR8qA9XUwyGwV4xAEpjkYGn+ULKK2jB+ezjHdxdrx/LOzbnEq1qfFhXWyg3O9
ceke3yQlZAu0VHe+35wXBxVe9yZfGFQ1dFKTnlpGwf+/4JCt/J3gvFHDpOh4Jrjd
aYknN5wkNVyUiveFvN2ufCxXNP6SI//n7qn2FHfwYfxjPxMtD8ScAb91zANgWtJE
9Bv+G7twlsDHvbZeHZW+aLD22p7RiIfMilRwh2FQ5j4wPa50shL8YEfbbQ6Fef1n
VriBTOgW8XO3sFPBQwGaMpGYU0OkWYFM4/jvowDtlpwJFxCUFKMwRP4RGMI2Svbk
VqcKi4xr3i3hKyNKUI4+s/AS6HCpxSpoX3+p4/9A+ywM+XebRl2UxdbmBHc4UQv+
huKfK063pgXD5viv8z6ZCgdWBAEY8pyoIuaYP55Oij7CpnwrCzOPTSsRq4t9wBLJ
XvOWTLk4QjPBtb4YJaCSfNgA/4fJW+L52AKirL5OIOW4hnelVTgHSMU+6nd0cVgD
Yx1KKWOzF7KvoON7pSIP1O8Ri815fLY3k8U+3Kri1txom3FSzat9Cf5oTDXGh2q+
Hi9EYPNiaP2HStZPjndR+w4b7m8mUA5NSYvdu3NKGEPH+dMS9PkwROkA4rg8O2GW
xHcda532dyQHCK3fJJC8e9mHF/5/B1oxxhCpqLfj082fPYFAFWCGkCoRFsbazJF+
mkf3W/lOPcGTgAQHnRBAmNdrxnfcl1iKcDupbV86C4jovVKR35UIwUt1DN/SscK5
8DfE2j0TN3BcawrBsA/ZqDkuE6s3eftDC8W25lORRPazJKsqStpokncdVZKsXDEM
Ck2s3W7MNhy0l+iL13W/6+V4hIP2bdQabVVgxsAo+aGXp1AgpBmTBC1lKpccmuOG
aMK9qRpN7MpJjOES45uc2FUqkQQezVZAqTx+x+taHwMot/o4mSV/RwZgkaIKQCaK
hQdcMPFzXtJn3CbPgxL7NoSG4HvI3J4fPcEc4KEsXM9whcoiMPfcZqqMYcyTmBEc
6Aap8Jx49yIhdQTsjCIC0ihTSKxPRACy4j75e8gWFGFxwSPh5b8hS0VZUb7rtCDs
JrxOSOMZcbx87LBtZ87zbED44xxuUOH5lBMB+4ngaKosEo1PJUNAzV3sPsFHzfUd
WImaS9kJv6PZieNVaXL5QSk7XLocDSOrkB667Nv9AcZ4zuVMnCzXfSVm/jbjPpG4
oKASF+Rbi/xMzFTDtY1T1+NCSMMy74md22mLIg6hTCcx2Yk+LufSbamXA6GOhmN7
2gIng8HafH+XZ6pTj4PiFZxWeppdHriqP6cGrBAcAhqt49YvW+7MSH54JI+FfZYB
WvWer/b23nGRYZBiYuag4tBF4iH7T7sH4E3r1vzdsUXiq6QdgN6VNDNkrzwnD3/C
K12GSvXmeDDblz5V00ZYXGcHPcuP9k0HvV+kMzWo5ncKRPpEAtUjLQcuN15a25Kd
HD1ADALtvRkdNfq8djyYcKCqk5ov+6f5JCqH0QYS8ebv4qXsnPnj+WNsaR/ylut8
12vPBQj7GrVClF7CQiUqerj+aHA6NDGcVLIydlIrGcdKxjR2X4HSVdr2q2UUK80y
pl1e2cgbHqx7uujxxn2FSE+ci/Uc1s2mLwYZhNobyIrtmxCBSWo3fOCUriwVoUkm
mZ7DXnij+ufV6lbgRclGqEJf+Y24K+QJc+cwy+Jm/N2pwnCc+nPod/uKM5sQ7SLD
jqeuXJK9RU6wUOZbUe7n8HwhBCnIcNTNuqxxCuq053hBDvEkWOrXpW23cH5SC0eH
5beNEM+MBjYV3XykCMuryOno8VoJz6NRYDGjF2XDOp3Eu/DPz64JzLRK6FSNg8d5
xX63jawjwZ2Sq24XPZ5hSM/1wCf3l92pjJG4FMxKlZoUfVLy9oc+eHMsIaCuoyKp
Uc7Biok2/VFHo8Ic9AAid554VmCudRiEcN8VnPubQLyzEO/eNtuTGVZfOl8CN8rR
2GWTbV7kJJF+ZUvQe//kf2wvghv0UvUJP6Sj+mQOvXMJrowcsAwhAGBZJpzWYETv
FUoSN3KYxAZpVP3BOPNhYbxA87hDGfDwAN9qmiNFYlY0ptkqtlyWH6h7N2PnYg1d
MY3nVsSOtwf9yvwyxVaXdyTHWlcZXWA33VrR+cby2d4nfMibjbNx92yVwMi/7qdz
bDe9WeKbenVBSIrK0n7z1RjWtJqwSSbh4LUuYUrbW9PLJpn4kCeKMr/kErlGuKVx
cehjI9fHUKHqwMX1W18m564Wh2QWBh7LnoGuCS9ReptOd7flRkayIHU2kJR9m7rK
vVqHUPwS1JxOlUQ56QjZEQ7desOiwgE9RYOHrizcyfbbWKHMLYy7Nhmnlum+coW+
2XzSlRIVWBPTmK2OWqOBpHCdhLeLDWSuXV6QG/Mgk90XxNhKLyX3y+ivLXtvoLar
tds4eVsDz4+AZ0BXTHHY7Y5+xZmxL/SBsdsbXoNAFDZMforLn/eT9+6LbPw21HVw
x3DTAPurQMuzjszEKyBHGbEqNCO6N9t7V5vyok6lnZe9ELYz7zgcsETkWPTuWmhR
Nre7CBQwAPDClgJt5DX+wNkgfUavuPIS0uCvyNfHFMSqWLCWFoeOsiXaPLHn/npB
Y7cAcKolcWddS4AP6KcLTTDy6jq+9SjMVwuvKT5LibhyagfwxlingyrqG0lGAruQ
FESqAKF6lmevl3uqDxJJbS/3AxocxSMvj1I8gUoEFo7XXMXAbXARa1OHXT/djcNL
EC2NJWg02A3oyv4WSN8PCifknkceQdHzEMufMaxwHy9F8Uuuq3OsP2leIuELcvBw
nidgNovYJl/qmOga69FAH+vh6YPSRNIMTN1NJElbek/4z6GJwndEXK4eB8j1rFj7
hYQwrKmGj0V93cjaPYmfh3bJddzRYG4QNa+DmQczm6yip6i3DI6YPdM6yjDCbz3a
+7rz4kRDy80vDMZNtK0fbIVb5VoA1LxUs9RqVxOfygx9xlNiD+mf/TyRTMTF9Rsa
GqbFDofkC+JKqBLgBhOBOSs7qYkT3c5nHmSgv2CA2yoNdUX/Jk1IimnNt9Qxrb1w
PeGJZBMlk39kRAwEGjtQlhYgjOAyZq0omOJ8ogCNVHIzrqCrS8Y6eQT+Y1ti7Q2g
WYCSigwQdtfhMLX+BfVYTQhoChpOAwPJ3wly3ypePz9/QLkawaTOqtxbBDP3/TRG
opKsQDjbvy3kVsJ60plR6L/nSPcMdRWWvzeEE+KkVML7ASNudBnDvx2DQj4ENAke
t/rkkPMX49GVxaICraEchPDh/diV944PIHGGkGCvgRpNVaD93mHkxUhow6gybRj3
3SG9VsfSXFG6rXdLRnX6OWqgjx7iIM5jinBvYyB4jFUv2/9NopVvNeA35EIqyH9b
RlI5zZuHAb7exeuHzMeSM+eFnwbprI/1ZKgRM4E/pczOiQRFabtSjZH83krXJtOh
AjVN12Z0xbEF3a8DrCNGPkyjkdNM1jeX1HtN4d2XJmLxlCFbKe2lG4NOocKknqkk
CUjv8W84mZyL4OQ1HvcWlaI+9N6z3RM0y4JpX150oLwBXBqsrV5ksQiR3J3WEiX4
6fwcJKlUT5WAzS2D5PU3z9U4W47GhA5IfyPXc3I490EKMsOOB9gy6A4spB76GYS9
AE7luQfl/n7raF64kKcexIxfO8kNfXXGaM6GSXFjrZUhRcrJoO89lKeMA87wfa28
HhFfUKzz4pgJ8M6FznP/Dkmn6lYL3R0KMbuhN3q/8gngdvtiOWuNeBHOrqxBH3n5
VuW6telDBnDWqAVHRrOp56Ri21i8omoHuGSnIYt1IExf3rloR69t0MVOWhhDLav/
ztqCRXVn+kR0SWGF5/Au548RUFGr3fF/nCnCTv1znNTPqRk6ca7XPkNzOc79OPZn
VE/HZSlhw/vDpyuDlbLsn0qfcn1fdpCv8mDE+kPRxTZeGMxjqv6uNziLeI+6rnZP
v74CAMrRqU1GbVDWvP8ogmrnokQmlO0OeoYQXz1A6CM1kKA46/8XBEG0W1SALLUS
ULrC1GIh4nHWmWPZcWDITGw/Bm5FCIOMFp46nrjbXz2w99X6NCGABaQH8kXSy4El
aU+cQCpzSHor0pt91jeRtBJkqqUYncSfgldJgM4THVg8xvK1gCaF0z45Nd9mv5Is
rINktg97jocEl4SrXP9JVT+nZQnJGE678OQKfQ+T3mfx9og55RXI+kMhJ4SBwkmY
6JHW8A8niioAWwzFcpFSK5j7m1V29SjZl5MqaKXv+n0U++l5uXw0QmdU90KGs+OD
MBaqUSsqJMtUn17uvTfBkaWhv2oPviFeuJLxs4JQDNO0HFYm1u7bXpzlyt0MXOoj
y1SU/0ECIkIuI8d2r9TsmEecG4yqB/np4QUc049K4SSdNUhDtQ0ipSdg76ZKFle/
DDynNcZ/K7kAJDHNrAJGMb53FCpOpf4+vBKIb1carUmz16QzcsFrgIi5NZFqFfD2
PpnrdQpivJVA1QKeRKv1cOTM1bHpwsSd3xo3xGChoQK0+exRuigd2v55YUX5tg0U
zAk6TifWOHr2n9NEDjQyA3WnRmL1/1AFYuCI8fn+nIQ+4f708T6weUrK6bNV9EPv
n6PgOyGWJDZDJLZlO9YNy2747in2AN1Kc8VWRZKaWru7YIsMsOXAbmargQ0lCo+U
4lFN/0Nft8lG/GPU4HIFCoUJ/hUQcFwx0pkcJXP2eZOUjJuDH4LzHtDItdKDrt3G
pUL/ucmNdtVgkZB9rhIDoSCNGwn8TJ/figoIy0dQJuhEDN1TW66crf4rONw+z7vf
DzzNOgXMa6kEYdrlDvtmhxbVlSd9qWv2CQgHGdhtZSnN0fv68SfE8bLuqFFbfvMS
Cel/3QnH2ytusEsLryHL8M8eE4QZK8A5OB2G+VGnFY02Aesjzdhi0c5WqnM7Mw+L
3Iw4rXEsEnE5wcko985EpU81QkH8FszB/kgVmf8cili6nw6aB7uLlvPvJdnvkhtn
lwpQ4/WHusDUnGnNPx2Wh5TGv5zpfVp3WCTJYvCHfh+qlWVixSB/sDTgxt9l4HzY
U0lCURvtM+NUs8vr46D13544OVQCU7xsN7Z8A5sYbGyH4eg1SHuJpDGvlv6Fdet7
1ZbpJe4jCopI/tb9OVhGP58jgTZkvikAxdt92i7lw6qMW8MfgPf9NVA/JptKgkDV
SMoAb4XwGm9nQzpuGzPiFY7s97faRAgr3qOZ2KwDFb3TTcDmf39wtGON2mqmfIrQ
Y50UfOPkHlr1xNb0PoQpRjRJRaQqoBTeUo08PcmKgIDNEf3HawytRgTCL6vvXToq
AlmzQUG5pjqdxobTiVUTjiNbEtwXjTmu0i6pVYGN14jkNZ6TMm/PQ21BHfPHybwZ
EZ0sQPDcz4+QI+y1Y48ldija4EgIy8hrBMX8TeE7YIWfFw9pLvwiJ2JNUdafCfN/
c8Z8oEcAM+Gx9RvUEGOIhrvwSJm2OA3m7esp5DxSbnE11RZmPbsTJpYPfQl+E5FR
ICNMHgtvQBwO5WnHpv7nLrwZxcF72tdL0smIXJqrub7Joukxk4deB0qdpgOfKq3g
OmT30ChmTeJAWOLumLk6THug8o5Tq5ULd9KHl7TnUWcfttEbAYLpXXOvjmTwxKXq
CGWcQnJ3EcFj8ExY3efkeEbEVfar6X6Klv3NmKDJehyicB9iTEBYONwCneJEqdTu
xj/Dlgggfa52yHUVJeOsIioXIYxdpusZ6K5eX2Okl9/w7d8hX5+tDy2GkOr2NIUQ
KCaIP5rs63fBF7m6LqPju4547qBShARtsV+ZPPBZQRtLZojyFuXiB/NcQgGoF880
dDp70nfglLnNxbz3T45GngYByO04SJQCEBwrc5zbgJUnFMyW92LBAf0+j8yWNUdX
bkDyGoQYPQ/okMNqFBK7MCbzp6lR66yveLHX+u0VN4V1lDQroHLZAw78dbazPpbw
COpDxNxxrz5R85JdUAOcSx1GHAb94zEfS7v7MbrzvN3qr1TCM1jjwpCdWKnJfHmq
O00SR8iC7m1CWZ+YE3ZILpni2A0rpac3ywueF5ZkyqiaCL7JG/q443whWcyAgOk9
eJFk6vQpHgJ0KA7bdlU+I57PdjJZ0BAqlNlLDaB4vlxY9lZM7EJKLE26BJS5Vf/K
M9fWeU+v8nRnXE6GnEmchNps/tnsjyNj3JyIktTrft6hq8qpq6cpPVqHkQ1fRQ5I
heA8v3zjJN2n8qmWp16LFRvO6UHh6Hmg2s3wfteLylKR/2vfnYhYa4uYduCFCyy1
ZrW5UDGy+eUu5kkZDDd77Kh5hqSei0ypIfKLHf4bnsjIqtVrbsyq/CwHJRnC+9mF
xurBapyG2HiTYOCyTX8WystoS7RwrvYxHI6MzWXCSClKaI+5/mJ0KRB2USQzn9Qr
0ycXgzBEBnCqd7nqlQoMOXyAd3hvJLAf+c2b/qOTv1LT1fMUP7/S2bj4OLa6zOHh
1KBICkzSsZO+E8j50GEU89l3vP+pL3DO+NCmGroLlkcOgbVBROsE/3eOwcdRuCHL
Qgnd9ECN0A1wRSw8VlcNBPcaeTLJZlgYKTAEmdMn1tUy2+KUO/l8MyTUG7CINvrd
0dcJeot6WEWRYPuq5Y5UBYQ/Usu5FgbpMLBSW+gyovV3oZuAyKkJqsqhCcVIlSx2
jLSBoPKL+So7tvt5tuVeLXCTHH+0arQ3gGjA2OKBcq4q2+LFjAE1HOLdJ1zN3MEW
hTq+9Bisa6/fS+MaXKO9HFBLI0X4ToeVoeG1tCx+JoTZhL/sK6mZQE3f0VHQ+vb6
d0aBU1ElAN0MNusv+fwPx9PpshKCGvHYU6f8Pb3+9Nsf93+C4fcfFug6QMGE+Xda
5kMoYPX6F1g0LMMewae/QCfB33Dqcdq/pl8Y6lZZkRy2d3W9lhALK7GduTY9YFuS
+gRlkGzguOp/azyZPLCcAyzfsQ3Na4CbqFkzh5EUufNgkfNQbFBHxym1+6+2yauJ
qLzFl9DZJfvG4kVHqpYJICUraMvzTkxy20Sjd/HmEPp0RC4lfJ5hyL4nJJOojVuR
xDeKxmHVHcwfD/JquCIv4WdcEaN6HL3dM3CM0dBK69kvPA19fWV5tGPQ1x6QDrsT
rdRXquwuksvAC0V7NimpYVvCeuaDL00kP5f0cytA/QWbDQRoNEEJL/J1KY038apc
+2znszpSN69Ko285AHCSI97CmRD/JD1C/zOTbji0u9p9CdGYooAQ2gazv4trAIsC
7z00nuE9maw0k3NEtIKO6jr50dzOj1qjUUk32sASBW6TZOpv1wtvUedjw0EfUZ1u
ea/v3VIzsFP925yO/Qb8Bc3cy6UgxN415hHUmRfH383Vk0Ae9/hMneullBvQjBp6
b0RUaRR2BFZ62IHeMWiA7GDGjJcGzOJt4Yikpjuh6z/lhwrZmcNyptqbSlgKMqku
DvHHFTGNfRHaL+kN0i15fp6GdzJm4PgJWxWOoJtEnPFkdV1niUs1TdgFALGyScKa
bd5KfnzMXSn3iQXewWxM+uuZS/u5/k7sbPjDoMpixwWG96a8RcM67NOdhZ21P/Vr
WBkeXIDAhzos+0Ktm7i0cBnddxgZUEODTdXpzPxnfZyHt6II3ribI70m60dAh9nu
Vf1IeRfvodXqo9pGJuNygQeYLvyi2KFiE/LR8J6RKNL2Lfnz9Mp3JK5UEOzTgffe
FqdYJaboE1uMPObGG2XvrS0di1q4JkTCwxhcl1EnDNFneEi4VKafvL0eVp+2G3QH
YLALaODhcLXCR0PvpiI8XOsyIPcEeAfdk/NvgSkuQ1I8upIcrzdVYdgl6sWKArQc
0RKht5dKEqs14zhcaWRGc6VMKTGBVZsYuOYqiqp/+o0T3nCoSXifJYIfUKJVpcXq
wGByYJn7eJSRKhtVx65PlXcumtIGz1p6+PvqHTosVFvXb7uutGG+Q6/JVS02x3wk
OMP6+QKYoZUvCxQ5Cvtt/4V7nQSA+Le7/Gcv0izHRPvuq3fNILJ3ESzotGKxnEHM
+HXl/WI4Ste5L4MLfy9L3Gmb0gDqO1dmAK5O2oPK6sUBlqx8EJEHNnqQjiXM0s2B
NFut0MMgAdEGKORTWz4lPUgqU+94fjEBx1xJcro1ZKEYzGvE2UX5B7ctrT10cq6y
YZEbJipuHD8yPovmqk2jJTStS0rYB1WRC9VJBpgrQXNVilGdVbL8VcMD7JiKa1Yz
oeqS2SDUyJYuBHLXJG+UQb3d2A/OOVsVgVnNq4zRPd8zGwhALp7d5LFKlFQMc+8+
qoC2H1fB0LAFyzXItEW4ByiNRFJoRuIpFNSTGBFXQqfZaGYeU3GycSlCYVqQtW5z
Q5Ru4jQxvG4Un1bmOuwx1BLSm9ucyCHUQqTvLX13u/U/Q3U37lHbtltbqN5nFp64
sEV2Rr4KAVkxkPPjyw6hMNGcVHZv9iXnrRjaBmtwonz7oewqXaBYefMYp7h83xpk
TSOjN/M5mm6W+C3VIgjtMZ2Dy2d28yvuhNxGYo5G7m0EXsoNmNUfuEizykxc1GFB
Jl4FjlZjK7Higpmz3fXyYmGNeZ32tZFA1isk7eUDK+oN76gwYMpah07WlbCrQ6IB
UTb4Lp3rBIHDT1EF8uyqTreZTyEBA1TZVpnCmZYbq6SJfFCxYGy84O4ZfnpnkmPj
GXEILgI9z7ONA0NzwqJu0xSVmfdJxxujBiHJOdBS+kzH0vR9vIMXSK151CafjzTq
D6LiSjde4A8VE3IHMS1j/fQhuSGDrgbiohJ/f5QXdMwlVNLuOAEROLdNKuFcU5i0
2kLlPq2PXVv0VGE8773Xj9d/vwvi89ewmsVJ2biWs/GAV5VbL/N/B2NYRCRPDQSP
dsfT76c6XegM8AjjZqv87FW6H/8WmmJHDE1OfbnsBXBgHZNDxSPpvwReILhqV6Ao
QnZm2eHJFoKCpnu3MKfd5LB0WOyCGFiI0UmMEqnemRK9i446z7j8PPRV3oiAxJXF
3fvv3wFap4im4/xWc33ihRS9jhUxzN+HbEIo+ZD4YzOhRB688gIvPEm4Lnn495zb
VcbGecW2PbIcUayYTAwRqlkLFMtdwTg/gtZ7EZmOkYeZKyhtVTPEhoLcywuxTYbV
8Y4CLdouGx6bJ/dTxIDbVLvSr313pnOeQ2rmFrnfzjF8dg69fx+1mW5X1gpOdD2D
N9HXWV3rVUKFOcvlchSKjhTNwOyEugwnKG0lRxZ4ftKyEqn1ZLO0uEJ4O7gOCcz6
GfltnbHV6grvN42tFkJKoyyoVQSz+8GSxrjLHsN5oFpseH11HpT+a4AhnyQOY2T9
NeVt+b3fUFnVEmaiXRTkJw76vh3n/RHzZp/P/Lv9EkZa8rS1njBJKvc45Oqxu7Rn
BTVCBgzQ6hhHwkqiu2Y9vW9jAf7BJmgaswPy1LC6wzgfej5uTRqUdvsn87y8e/Ib
7FRZ37ud35j4cyqrFfainZtmuxCBaat4kzosdR0r0+cw8JSsHf5expAKJX6mqCoU
my0pXebace6+itmSVkDHkWhGTRpeotGP3lM2cq68hmzHswIBf1nozuhwqxsFJ9nI
P6AhVN+9GZOhyU/TWhFfSlmqae8PPyQH9e2KOUHIf1O+4uWnaXNwOisfjOkfQwyH
J/x+UyvSTLNt/k/esyoZWHwzvRRFG2BVvFln1h/ZkffZwVfwmi+rwdXZLx7dEzhG
sK47IjLHK85yEH93QpIWVM/R+3MvYXYu9mdkD0Ein+uQ0ukgGqGjhOko40OYvp/1
8usneeTQGr5RYPBxr+bv55162reNVqnwIbr1v1jfOp6NWW5/GXukuOSTOW1xtf9F
q8c6yicuu6qNqOFqZK/80kcwXmj/kf/2Efw/LpGBC7NebBy6s+FUKOLTgE4phqfd
55kqOfu0rIn4uHbgjOnCKTjrloA0MrBzEZxcjju+yYr05FNvfFKrFCIQEpPAgQM0
l7iVNQqt4ha/CIe4271gaDcDyhSTgUGjDTbXlei5dmYhHHKFlI0TPw17Ufvr0giO
BWeFoESwrdCzxr6fB7VV66+YNoRcz01uRN29lvl3yzDzQUndA0T8zmA1bvXam8qu
AnWbCeHT1BqJ2I+0z8yXOryQUyQ1IRzNLWYua5hfQPw/cA4o7n4FCuM7b2ar4her
Tkm+W9C2GgSRDo3Cc6Gm85Eh7CnJ9j0krInrzXseKxzMWIB08LFnTFf77ocmtR8x
fFyN87rruHURpUyY1hlbw9aRZ1t7NPCi2Li2xgNhsUm9RMnJzw+ks4HwBvRYCvCV
nLOT++tBG5nGkUpWOFw8VyU7c0h5pcTDjNo9aFcaNlKz49GFBspXVCMtISVhnwub
hds8gvW8Dip30t359Y4pVMsOj5kQ0kM3TsrejcxIsTF9MONCB7hugGsWvOGrNogn
xkfW2ZZ9qc1ufp6vaP/7JZO/Tn+dFqP+ltoRL4yyQ0uvoytME44Z2c4q3q4N8HrZ
AFAhsZCaB8RZLvkOUeiHnlFFukk9WQ4uDzlFexvl+/7M+g0hsL4A3LrApJZZ9N3t
udg7ypjmkY6ZHk+tfCSltVyZJvnUAqYs/qw0/L+q6ZmcaIbi6t39QZPikgu+63HF
uQ/K6p1baMRl/XYvsI0vURm5jLuzGlMMrxEgMfphdRLu/uSHwe6CVDph1fKg2UZq
++/3wR5yrVAxTXPhQhVp8nJU9Hn1FsG8qA5wgriJjMV4eLZr8KmtlBMtoANuuAYS
CSr9TAHGKu7MWfu6Q2WOD07F+nZt+AYWuEEX4MNdSP5BsZELi911S2rsl6dbm23x
nesrU1Lj0BWkr5UvgoctnB4V4xXJKc8XeB7UJdZfns7PWi2PW03Wvw420rLk8Dmo
9/3I/h8ND4l/6PdPvn/Miw6XsxxOIjZWUF3QnJL711j0UrukIAjRpAU1NTEhHiEk
Y+i9zOj4k2tNkgL9cXzG0b25QV92hBVlOqlxO5drPNeu0GLkZRna2BReE8xxvVzM
ye3ALj7ulcvTGmRYj4xj4mF3nywGWLBqJwnaS4RbBrHY03Q1M9VfyPOqyjF7cDgN
990oSNestZxffqePJQ8ZeiHSYD8GyCRjGhBuBlw+gELvxDu61LW7J4RdM5KdUlO8
4rcnacFCyxfoSVgiJebrgBDaj1sUGmFvfETg69cvBdwK095+uKeOjiCTWQLPDxcu
3zJ22qDVe6qsxEKLdI6YYA4xHKu6PAI50hcrlZNDtIR1fsOEf88unfXezijFDSnQ
n2kt1NKTAUo97nlsT1lc1ZpxA3sEHX7kldtvL2iY2lvHl/xvfYJpis9PxIFqNKbJ
T48kypy7iDgnBpM5/3pYjpUhtByRKbC+IJCCURDNZjcmDCza2xE4ULXd20yu4tFV
WETYI9yxxMa1GmLKOrlkBI34GpiF31hPctjSeBiPrrhs03DQSow9hWAmpabInHhq
+ThpZsEuuHoN/+PsB+FnJoEucwLsirDHVyM7xUPdL94br0gwOMuNOQiQjashwFkO
VxaCHvAl7kicQYvYcpAT5kLuB0posamSaGVkljsshZ7j8CrzgRqTNvllSiOkaGJT
PODdwC6iHwJ3ycpTGrsFY+P+bkIMRFfI81BskhtLCRYFSLySmtrOAAYClBjFvcTW
j+6IlG8eJSv3GGL4WauDr79fAGILtZQ+mnhDh7TN/emkMCnw1EyG2hzAGJ4FbB46
uxBHUcNpXQSWOVZJSXzialR4APu7931Lar6+XgI2SohE8nx82cr3lxwxl7zzVJen
TXI94UN1Y8XMHDmePg+hBJhZXVXA9VExKmBjqCU93wc2p+dU/0QWv4RzWNTYh6gD
c6L0CF0zynY4RTkZK+69U/Su6x9Bu8av93wLWciuiz9Y5S1/Wrg5u0+FQHQh8jPB
ePJKDRhSPg2iBPJc2INYI9Fr1OMaO4OobGqseo3EPBYRkQ61uUC7AqfR762TRDMc
5a8Js56GOv3uj1sVcBsymlfrYMWm14VYC+O/l2ias8ICljzCsJ6CzBo1OgiO3WU/
Mfya6/m6zNsnP19d0J7dlo7BQU4NsPKxG4t24+tyqZQZ8hwUedx+tNQVnYHY45BF
x2QK9A9+cl9UmUilnNwf7WIgdemUqA1X8QTcEBUkLAeyppMCOJ+OcqG8xDJgsjDN
u546h+0rVV5zPuvWKVHzVgBl03MAyGmAr5/DTND3stEQWv9adiGOLpkTUM9YJ0Ny
mAS3cdBt9RcbhiKhSqP9lCqevIIYdOGN1CNp3e2BvedN3BY/p6dXhr0no2mG/pam
UFLBNu+URzUuDCz4yVkX6kA0N9WZDpD/6CCvzAm0SNZmA3ssN4V7jta3bE0dkFQJ
dPSos4XhRPGLjTFpUyZH8/UO+QCZstZuLcPBPRl9vrI70ppMkAQGT4Bi3KdBLQ57
zD7j9WDIANMbnSwKzuCiS0VvG3KWWVy7diPeeaoZrIFP/QL0cGM6aEzeFZ6XPjur
mILpfVrcbtFT5xM/SajRWrev8HwTHynFrZkW871bM87pLEHWNLNSWcmQHsDtR2+3
txySml65pcXCwP8D+aFgBzUDhdwfItpHyJUEiNYa9cAs0W95AjdqGioybuXiwrTc
Ua8x74yeykAmGVfoWGKL8BElR3wg/EdyiH/6aPoj/x1+p6kSXb1aFtCKBQTcoKir
xR1wGDkZwtEgXBetUHyjcwQjy/J6Dk1TR0mbBYhGFXVgZfuX3idSkfk4H5kho39G
tjhZv6FEgFlYswc/wL16nWxnF8AW2DdMO5vcYOsw4wO0CScrZ6PFsWuOuYdiVi4S
cU0ySRB+t16N4Ppq+n21B1oAp7b01fWGVXSsVMP1K79cOteAcDnsRrxd0SmEeAIS
ub2/QdITtVh03q9zfNTy1TxiQ4hpJC61/JbmQdgWZskMikSFeiDU8K/YyVnLvHTw
thgVgPb+L/A8d8Nf31E/vD2yO2P54UxdD/Vv3E6zVobQjdsz3y7dztx3IHjQzubn
lZx0KaPqrTCm8/KnVQkGP6k8Z91+DsyyWdLHvMfmv+UjgD20FPVhjuw4JWbZ1+Dh
8232kbJL8JZdroOPbetK+gynbe2PCM72CHZD7RfIYe1pi69PeD380IxJ433xcDYU
AVppsYwZdaqLuRaYfl/i+wVBNLACtvqaIV6bzMjvjF6f8ALn1Xey0nn8/oc7lCqR
bxjzFstMbvHbF1Bl08elcI4EALLdq6zOPfEPLhMwUwSE01XDUuPT6G8yxdoJYroL
TehNSumbtkwrnHMx6a0jUbrQ/+yYDC+MRIVeGHrfFNFpHp08SmTepZRl1wpt0pEB
KmC54KsE8F9OFkzGfI2sNwuANx3vZeE3dHpu/szqebCShEmH8psa6V91i1UI/4XW
9Ji77AexCeWki3SukQi3i7uooCbGdHkYiHtgenCWexolhTGwvrZ52GP6tzne/FXt
LpTzxPB6n1hch1QvjPBYWO2R01bfUA2HWJei5R9h3JFqslxICS574ZJT+G52uwqR
J79ZEM4209gAcxtE9WXUCyRWAUo+5qfNaAPXrrbnhvSLhxrk7xbusFPJdeQ8xCPO
VLTVbF2YgQMDIBAYpqkrjAFNFUBSsCIQkJFItbnbPZ+BYKEqh2l0SPwd0KX/OzAX
2pBb2CcZZmuCnr6LY2rBS6CzBUnPE58tpDQvdu8uINzUrO+gdqjxCEyETfRO90gV
cyAWBKF3KAQHwYCr3K5qA63koGU+4OIqy6V3luEOBbud+pAaKIg7M4gXEljWVVRK
oHkfxmWSSddhwTCRgRzyT4vI70cIvrzlZotxozQ22jiVFB6oeo+N6zYuoF30YZdF
eK/gRgfY4TwdmIt/tV0z0dys7GZ6UGB8c3dbowPqK5Ezi4bhgdhjiQ0fc3rUygb/
+aS1un+Hxw085i/WX+XgrAgq1lu2zbdBiJG/QCT7wawpS+dS0iSnEGH1bq37MD5Y
d2R/8Nvr5gFFaoDvG+HTp+Q0uL1GLtApURdN0N4VkfNjhxGSl56nVFDgqKfwP7R7
JieLIYaRdUHc9zSlrX7agN5236yrCsOYjYSbBYD5k7QbBN7t675E+MsZaXokXsIR
ivt21/Wjm6Xb/pGfjeEFjmcRjP8M+NoWsqRXJ68pM2tuk6VzqQLw8v5b5AzxwvKD
wCgHcUZ/hGTqaApJkNRMwb2DIa6weIbxgJGuAft1uzEECG4yKNGMdd9jU3+ipETV
5pqlUyRc4SsjrbWF6Zyk39RroqGIW3GH6LuTEEuSxCt/LwLz+IsBrRbSb1FFRBqU
aoBmGsyXVw2Q6rgEAtCC3Arc59WD3bX8oxfdzT0dlL9rJzBOdXWOwPnDgMEcknHP
cJPyfV2d3OGMcjsADR+x+4VmnlWsobNODW5Zqp0L5urqCQwKR1PF3xFb4D8SZleG
btnzamAWmcR1O9/v6HqAn0SVLXg81OolG78tK/Gcr2bnCl4vrcb987Z81XBYouKk
D6tM06mzifM21OVTV/BstJqdQP31EawEWFmJmo/fYm080NZWtfWx/v/UUb6EdmLY
KT76bGS/Bp52LTz3GB3wj+qTVnTPIHdmXBZHkhOQm7EQclke6RfESvivnSnEZ1HH
C3W42BBSkLANjiakv0n7boT2tLOVgTyITuYmlodG3m80kyhGPvkqfHD23xMifX9Q
YjI0H46WF0jVrwB05jz3IZj61zNASVyp6MAc+VIUhUNiTGUPdKm3JCzZT2y5sziN
71fwpFx/JFAN0TjsZL2tf+sMDrIAyEGt7ngN74ZReOVxTq3wHM81EoaFksROjwlY
mBNHTZyZkshJ5dgwbkGUTm4umFC7mZCBt5Uat1U6lsaRru/2R2mwwDw8p2av75kO
0oz3+E08UUWH+a+F6iEtrn9jGrBcx4Qu6axoN0eIhCbMoYeMJjxYtxtCxzMSA+IW
cV7EWpVa4OnQ9dqW8HRFgh3Wb22bqZGPnqKh9MNfJZI5EnXw9nFrZqocCimbHaWp
FSqLnWTrE2hF2f9g/1cuY6L7K0zENcGndutNtIIh0YlW9pslAIcravIGfs1dEXgh
g4WJXUCW4uJElUfv0VDuUwv6366QNQh6P6wdeqxqcVbWuMC0x81VzrkmjHuMAW69
9ERV3QWGd+rxhKAu8yXJy78IgdZQi88xpn8/uO111KZaM1tom2DMhmiE+keF9Mz1
Y0YA1tIQ2XXHwStaTpI4oPKzq6x8RUlyngneFn0M49XEJJxxsvk9mEljIsj4W8e3
Wx6JLPcK5aJ8WP2hcw2WSXnYF3ueNwj2by8uE4enQyRbsTlQsIYRZZF7peebclsm
N4Pz3Gdaoxs8SxtcgopAqJWK4VKY5XxuATj8jz6ak5dRoka2Y/u7baJCm8UgFrLN
GpGHodSUOzvukoR8sM/5hgQigy1gU6LkdfpO3VFlC4zwoC4Yt+UsAZgjrISYFyqE
OcKJAybxBsM6zEpQwncFstrP3c9GotRhpGzT0dDuboR+KK03IViNmrh+tMGfRb9D
8412Hr7o+YkcsZgwACoSZo9WzBl+zoLc/Ec5tWwOiejQaztfGFYaaCk1Sr7Cr1Xn
gT6s2BpUNZd34QEcwk90Fnqfsltp4Q9kQYqcjKXA2TIb7vPpEdtRLE31S5sSI3Ry
BTy8CnlgSg/vpxTLfRAPAiSSt8eEMzX9F7NfC780qFkLW0OCXQ1joQwfBXW5rkQV
Y+zSb+MG3TyiT5ex4W5a98Cta/pIsji2Ah3RmThouLa8jn7ZDNg+8odyvH08X4yh
TQhcjpKWXKbMoSf9nqLTfN2K0IejX/rVA0wmiYdF5+ozWTzYgmfUqMfyCJxjHBE/
f56pqy5lkQAHZEowC66aQGCHJk7LQJJyY65dMfbTdoP8zm3YPVt6w8Xuc/p/sILV
/RuXbCBL3SlGj3yDrvJZM/8l5/3WSCjgycucnh/2xHWkly0JzKNpYl026Jf3vGWj
AI6wUI9MXC0dVVaHeRqJs5TR0oJPSkoTLCQRk43nRzrrgtllJpS15Sse9m6WFsyt
KNJr+DL3i3xlEtNzIkUezuVUlMrQwBjZmt/QImTvUDejT7YE+fO9VxWlaPrIkrwC
QHf1N0K7yKm0Odf7B1OH+N0jJvx8oCSu8ZujH5HbThZQPgyfVSUTS60asS3+fCjc
DRK8LI1qFCrlBWPFobT940LoJGPPvRL6QwlrGT8F8u8OkBC62HLc5wj9xt8oKHft
zJeFsj79d5ILOASGibgrINbzZAccCRJE4ThH5ZquTFYzSFzDSSnZ6OpUOaDmh+VI
G76rfE16KDbKTqLgXrbhPD5MHGfCPodeonAxkMEYK3HhU6/Khhwa4k4p3XROgYH1
Y1mWiiu/d1wTsuyqLrP0hHfNIMK5pjJxpImKtbn+Ggv+yKRZT8KOfOpLvyfCY5Cj
hJT/hAQw8L5B0YfB/6FQpejPD2g/tyfM3Nd8b0KvN4ZUPc4KrFDi9dLtu7qXAoun
Vbb2D7GQplp7AiRQeenVUyLTWFahUiI8bOyCA32oxdeEuAoZjvko1Nr6sQq0upes
EfDVgZmPQbphe2zpWEYLYxRz6o8uDO8AcS0/yY1W9ykSkRXmAkFrItWQ40Bx4hSC
MfbR+h9h3RdRHTalBb38PpyFn2ac6l9o05dFsjWDoybH0WAdcEIGvJC65V9owUys
cf5oRubL/etWnpftF+N3RmnIdzlapn+JjM0PPsCCaNXUMAzQaM46HhQ0UvHlT2Z8
xa/j+R+gp4+gCFXSPgVlU4+KrL6VqlJI17o4oowHbsWmh4UPZdDiLyLlxptkeTV4
oADgqw64FqeFvPHpdc3c0SWAajE9BTy7GPaQ0gy5X48ZrI2Z5BaoNbg+Er4Ogcjz
OCzbHzmrcB1YKEzxfoguqHhe5fAxpxbMsxMafeUxNrrpiD5TSvYqypYrfQOKR7by
uVwNwPwkbx/E6qs+wprk3hc6YPmEQtb1xT6aj/XrTBT0pnqHqL8jv802fTUzfbRK
4oiLhrtrYw+QOowA8b8lDqj/tnWAamp2asEFWsNX7cuDsIYbWqp9LWqSMXA9uo2I
Sh0HwlN1VjlIPS9JWi5jC354HTkewpcH4Kv+0EDq/qRM2Csgrg2J3PrIaA3/nziJ
ua2XOJyFZU+ti6e3f0J4/A0Lc0M5JAniVSY18pDm6ID2n+7eALz/VVMcfGJWxWBR
EX2V4K+YUgsJVTJMnsqJYEJ2lLir2gJNviSQUc6BSWCveA9iRAZlEsITTIcTPuxp
tEWj7Y8s6h8DYnFe3MCQDzAJ/y5vOu+sP7Tuu0x+pjbCWuN2RW/QQAwoqbpQyeIb
6bdSQUMm2FqwfGajdA6A+VVY9j1TJKZpkdcJwXVi/J3RGqBtCTwYXVKO6QP9kkWT
cZzsjammILvDsW+zAoJyszy58sd6KzeUtfLS9WJ9zH7nkfycMtoi1Xuc5tasZjC6
flOmHmS1sz+ZnMXdBMkrXAIGDD9GqnVFn6V9u/hpQaAGnYdgUZHho/tbHct+61Qo
1KqTt1h53YfXIEjEzIEw23dmjfZgc8zcoGWaIqmdG7xtHxmdG280B5svxSEtZre9
6qr9qjvgHMgDaaveMElAsMmF7FR5VXRbikDGCmgVMCasSX5qLhhc7sK8hfzrJLMc
ouIZTQJxGybH5tWn1yaDQy13p6Zy1hkZteUY8/HyiYnN0p4nqKqOo3sot2T86hgj
TVIZtzPAONyv2DJxPc0P1QbnzmrG+BmuJUo5zJuJAMBeLk/yugpGqbtzZIUsJsTI
RzfD23GvfUsKAx2oaUOPgQNUdsT4ZH9UXaF2GhBWlKo6wcbHXIb3KcuGCXmZFnLd
pLBh0U22iGwpGYFpFaawvKxsUyttMnm8k6KCgX51So49toaexUCLeAxcHG3xlNyv
LEpxqzx/XJ/u6uAZ17pBlgKkXpMGgcLp3s0d/aosn350zj+lFkDCMHnKRekE/GXs
8bOs9oVpxxRExhwb2p1+IffSKPa9e711AU1H/qQFDkRzgj6mWIeApekTLrJi4eE7
/Aipljr2qbCbKXcd+ura4vplapYHtSc4eGFpVpxWTrRbvPYU5voed9TYxkmlCMAI
aXm0bXx+Z9VmAmzbzYRnXjxiCwGwcyD/8tK/ehG2RDpNU+Qc4NhUHojrVjh7/whv
L4KMbyy/NeNKCXFEWRvldPs+M3j5qtjPOga6AtORYCYJpzK2WkRH0TGCiFC6Sw3t
6BkLe9pI+WEpMlVXVOKtTFPJbyP8QhGmzvKOMYJpFGvo1XPSnOccHoyCg/q3h8SN
rN/e8DU0TwFUfxppFWq+JrVKTNNht+pH2bmV4wMcioaKoysmCRfBYbFRkTZ2AKI0
C4kpdvf8Sse5MVyYFXFioxmJCPB/tW3BBVyDiW0tdXXmQi0mmbICxx39fd2Qkn/Y
t3nT/0PxtVQyJFX9p79blJqLeMpe8g2mT1aGInz3bxW3344hFb6CbbSmEWX0QbJg
ZXb5eDs+W6hG27Alw/K9MNAQ1nTnOawZZXnhkuIRHDpT4LsfVwXPlVjPumncsMU5
x7l842Eo21wQ/W08bqrZHJwfyGVmckQJUpo88GsD7QNdYg6Ab224IFcnCZH0oTmY
0Q2+W5+IS+ybi5ngl3L3dSVdNbi8kav338LJ3ouZW+dByrSOfrpid4yXlrxfjx6r
P+btJTXCFO7PzWuwDrz5w6ERg2Igd5Mdqrew23OVlJo6kPK+VUirJck2JEzkmRWe
AzDTMSA0FnbTlP1r5odMC+cFWq3qp801smvp/qfcC2ohwUdelwlW+g6VPvMTwPTr
xEyD6Hdzx0Y1jfN//Ep6OmP77aTx9EXHOLM/hDs2gRdICFg7tBdJ6eupk+VbZxRR
5WxeKHPXkhlL6La6wysMh4S3BmDaOuEwbm/GvhEXDSOjeemttsgSEGRUAJoTGqeD
gWEYrw0nK99dhfN7FlHZk6XTHsooIU5h45KnhjGqVm/+P2//0I0YghtujAsbBeAP
sdxuWrlx3Uz3zL07QvVrxPmCtDQtMuhgvMT0IYHO0n5iHI7JI/ynhvF5qRlZ+Odu
w+wnda6hfMVQuYEDFaK2klQwzWtogYnsuEZAFQR1akD9g94ICaJ1AU6qyV7jnm92
VoKzk9D0AMPB/k/8RMhkLB25ItNWJ7NKn+MqNTU2aqWS0ziztjlY768wlOWAsxB8
br5Ldd25ohe9UZ1kXjpuLbo0pAX+IHpELCxOBlSUaShX1RL4jOXROKALE4IDfOVN
dtGfC0ujrEWzViEpnaI21I5t9nsxPnWJ6IMCjlxjSQfoZdpmJeaImw8j3Cpb1nf1
ZGoD/JfAIjY8XdRII49HX4zgAFC5iKoYYc3L7fV8d0CXLgU7y4x52nvs7TRH7trS
+ndYuCUq3ONN91BscXWAfhY1LJXVgNYGj2xBZIo8iai7PulX3yl0VpspZs4PBlTS
STMQX2LCQwRcrEfFbmgn/GDfDPqvVgnPzWBq6S4JQGwnfZ0z8z1JPZGRM643/99r
CeYW3+n5v/Q4QTVQz2MijnAcAUx016UZTTO4a2k+8zok0OuaXRkYielBYiJ4WbfD
7/SVyRXx0UJMOgsTelB0eJzWHd/1gQDT5Wc0o9X1GmhrS8tRpKQoOlu6PZU8iT1a
RX9ZnV63W+3P1XziLhtPvVhrllHycLxGB//aca2fpm18bEyk9TH5iEBcLpgWSMu7
jhUYn+PbcxhCMT1OhnbvXxrtQ0Ejue2IPcdE8lHibJfUdYwBA3mtjQpsza2uOLav
+SSfZkrrkzTP+EJQWUpsSsl4AQtHdw79VzxyPi9tUALajkZbLQRJJVSfR3oELZlT
osCjZPcXHs8P808djBcajvlV55JKoHBEIoNk+eA0PusMia6Hp6qFYXJsHszxuHf8
WyKiijTqwdJc5JUnJHcXhl37PYjOebc/lVhEoIdGRKoTec07L2yQDAAG9rxp0JIX
/hDDsF8b5WKx4SZkY0CvgIIc56iVt5cixKIHkmj7RO7mUzmqJom49B6p7KHD4jc9
5p32cleGJim7rVD+lkzhZ7kaeHITOaqCyYovVIdTUdf/BPbl6tP1o+dcFXHRD8Gj
Mo7INDOhqrZ7DhSw0vsAbOlhrPs7pYR8cTuQ0VAKPPyRyIlrjlB+3z44k3b82/JB
JsIYVHfm/tKJ3JTi1pdL7eFNV5iDhFJSZ5tjKcGHR1Q5FeMIdLTMw+na/9yjZ/Ia
S7LgAhjOPztgccFizYXWJO4t651NOJn0iLTvsjdsfV2ssRVM6nAeqqlyCw2KcHZ/
SOraZaG16FUochp5KF9B6EWtwiWx3XYeFDdHCn5NNG9/dzJAHvOJymo0jT6Hj6Zc
B66HkAPa/8S0zQlw++LNoUE506D7dzWNabHM9wcCeGmjCVzJweUuytKOOp/hIbMs
ES7z1ZIsXe30XTnB08Qm3Ygqbgmt6fzjfsc+nBVwyugBkkbm+wKtN/R3Dpf4CRy6
Aauitc0CXii5s8pbu1yHOUa0PiW8DUr+RU5+5TjZ+5btTUM8GfJKszxH74v2N2cx
56OLAjn3kxiU31QuOUMKvHYJA/17Kk2Cni2bhPYjHACRqeSsCkUPDJCgNRohSOdR
IX3T2XAOjbRlBVsWdvmNuB82umWAhBslrCttJ+iwcRh3lTP+xfsVNB/uD33hMUXf
vEgLRuU5bzzKaXdQCCTijRw3jZdf1oTv1yAiQD3+b4UiSUs0BrEkkq9J4Afems47
OxaQmRgyO13rX3HaO+tVzygSMwDKj7DlkTSCRWjcn8nK/l1/4zNkWb7wKyNdSRJ2
v8ryjWIqk40EVXhgSf6hY2os/Lzkw6kqzoA3XH/jKWSOwUAAe7PO2ZbPPZxhgwMg
dEEG8ublE4AA0mycuUERLs5hxuyB2SlLuU9fSzi+ynRmmDZHv007YYZ5L25flE7s
Tc2EePcWSC42mqYUOPitKusgnF1F0/W69B9pzu2fP1GyYE/PdZbdXWAbofO0htki
pVsg0dzal14GpLmL/2SJUpMj7r/wlsAC5EfJMhP5xWm7RwO36hA8KC4Oz4AB2cqr
Xsi6usBwEf0pxiTElCYiG6ZUC/HaK9HDlYIo6NQmwZweiZ202h0Yu7uLAZFPov5d
1GwtYbFUIQsmbbWkIfIZ4ttVJ3+T5SXvRpfy7x48nU5F7pML6iSplurX9ZL4fGHX
MuzZBma2DR260H/60UlsN+UHd4A4Gd2Zon7oeWo3U/4Tnd4CtQNMYpV6YSYKB+gw
th2ONgiL9w4UkV6RLiHrWLy9Hoxa9PH3wFMcqcNcEjckEw9uGgqU4uff2+sS5yn/
sQzCNAbTu6Sm1hk6qJ4lS4Cu5VS9k3C1HFw8naOkvJOIr6PWl/2ia/fNhIa20/lr
n1pj1GaU6K4W0cxM3WED+3Ztf12TbSPzrvDGzrfmxW2Sxr97hw6AMqZ9Tct/aN4g
bFzJKI55RKd0OtxdpHDe8e5c2lLFoj+q2LegBUMkcKMawaHPhuTCl74ylEuln2dM
O9hZQBy5GWM+8oubetg/c2ZPGONGdeWVkPcbAIq36kd/IrgnauNEAkmsjA+DtDxS
TnxyuiK/9EDyBlJTVcpJM5rJUva97CVGS/JrVP8WAsQ0nkwRDKvGb6VkPZ41Nh1F
hYPNVPT3xut1aO6nQFnRjJCcIm10h3b9NNSw+vrGwysr94pxlkW5bD3A+R1uMMVa
0AMrN+HCyFC3WRI9a4P3bLh7A90qdcRJp4ilZGiVnvFhcZEPwV7qW9Jbxik+AHGl
wFjHDqCroyASVudpKn0o7QJabOtlKn0wZbvwAJ3YrKb/NpA5AyuT90jumzJYUlBP
Ppd9kxwX/7znNZLKQZ73moPJgkqf58rzNpKhciUL4nHxc9LNgnuicgshuIYTKRcq
SEPdzgfC+KErQMHH0vleD3sBpYFqFyodSmoHYt1sF6bNhZmQluJWO9Us3MI5aHm1
ExeXaeaOu890H3It1dsWJnphc2Ego3r/Qbt0G3SU/Dehu+AGPjlhEEl6NizBh89s
atV4wkxAY0Fw5LKxLf20b8ZYCXQPDs7GEKPOmc0VWfzYTtnMevddMOFOJgGhUXtf
e5tluXuqLY04v5rFe1q0DRDpkMReRPElZglzknh/4WgcWXg0DTO7va3oO2F7QIe4
Z5L5BYF05y0LYO6fzf4Iqc9n24V8f+YUO+m0bkn1FBgA5SPDgnf3cSkMZ9NtfJNT
jE8n5pelNI126Y3meDkcLFarPTxVV8r4Tq37AYMRy7ugGLJmajAl+fRH2VoOjvM3
wLmutTxCt5JR7zoTpLjKB+VJpTyEjfhTqZkxAltlhOtMV08ak/+7EsCAyJCClt02
NFYHBrKC0Not9SDVDCMKkKjv9G0uTxaSSBlw58X2Z3iMNHJRFwimsDoPUpJ3I3Wq
9glyEl/Aex79KxbHUmUzq4DI/LODIPNzggWbPYJqvmPf7rlQCR0Ya6Coad8wTRV/
bvj6zPu/Xl0skzmjQSHuKwLSCWUGXMZ/Sw8oxR9LP8vXetxAR8DsCCaLHmDQf+6T
ODP1vSSLS1O3ZgQRUYHmWuXAhQ1SFWzqu69u66y6oQmEHqGdvj9qIsLzP6jA1hm7
kTtoBMPF9IqSrOBJsbfKCnXlRGGkXNFQghICGGCgeJvatvGL69OR6q9Ycg4UPUwe
5FrKt46XTwPnFekKCRODprkDAvZJGxQz6nxeY7pM5DQvzYEz91LhDJ5k+kcm7dtX
EVRoa0RqbEjXXpP8Sn3jCOU91kp0T8LZFvi3CWV6Fc2hxVbdSeEFKKG6z2RPDTFI
EkjQ9EoQtAjwkNK6XsZw/HN/MoGAFFwxU0aumzx9YkP9IzZ6+2xjhylUgk8SvUYq
84Ct1mEKAYmHm60BlW0HHAm0qVgBH3JS585Rce4klCdMHI77NmyvXeErK+KbhOj2
m0x9f/rvgI3+LTffBW/7VvnGlM1oVv6pz+mGNk2/j5Vp5OtofDIiNl35ktRkgpkn
o1qM+FYxMk+0joeQsSMemKV7n7opiphaPrteXcp3jB4nHkngucW4XP8Sa12TqCtb
vLEBiXxgb/xKhGfKiTsXc7AuU3bNfpl3MwiOoh3cPhaOwZKbRgI9cEVVUVpN+ib+
yEnlHAIRi94cmInxtabMd+uWuZIz9RNyEmiVU9LHNTK9NCAAmBgbRqWX/iFs3Z7E
V8KWPL3U0ZVMvlkhxJ/PyszFAVTwsm9bLYwKe2yI5QO50qtoKcGMq46099/82sI5
lNvAPkizrmVVA3Vkfr3r1FegBEaUbPK6bWxBa5xMokxDCxRibcuAhaD32dy8iujh
8y9GFVaZIiUh0AcpzT4EpfuIso4CFvYBG8ARceiR6GHyB4WN5i8Ueq9TMm1L6lL2
0BOSGw8yspKOha8aS7esm2kaRy7lUMBgwVUW9Z6an+3Hn0aOwqYFeZSO2f4/rr+9
+ISnwrdtSvUhDNi9kpvYBrTosFYJ+h0rZGYPb38umAtScGhV9i4IkU9M/scAkUXq
SWIfFQCXRXg/27RK2Or7aj02zq7IIKV5D0W1Y79Wp+Pdh8ikFqhHeOEVM+cLLnFZ
gwtqNSrfKtxIMveo26dvXp2hwIYKKl60fqjuaKjK8GfIXXBxFOZQglSG3FETNF/b
gm+1i9jGx36WpCHR20KlrwlQjV0TSnl9ZqZ3M60rS109Tvn+Nc9dxGCSpG+LxLhp
EWapPwV6SFLqs8mznBVLLif4r12In9QeDmOx/SG1R2GUh1kBsaOc2F6Coy1XQJKo
QLW7JTnES3Yq92oUGmktJZA7NO9dvQR2Z3FMJ0NxJLuXiOEqyHstBrNy3IOyou8x
5L1Bj7M9Yp7HTXlbQ7xdC2CO70Dordyp/eySEF/60JXOlXjX57J8Q74gFJLHWe4D
W9SEVrGW0v4rpIFOOsUt4C6dTA0+tu0Kb59Tt/0mpD1qwX2uGv50YFNRs3NNqEEh
ruU8s4aEDbzghIgYa0gO+G1A4slhKI3/2Oy1M/aScTLaa/c9ICKlf08MIaMYgepV
7O+BJib/kfTx7tqz2NIKNkwJMojDGOViXkLy1w38tPHHbR/3jZyILXW8zu8kKAQP
edC8cnJlxRguySrFJxODvqseaJOUc0G2QaaNZchPkqHivdEGjhybixmxk8opdzRL
sUM1ILzOB9LV2Lmf4viUaWpNaY7i2QSOlSF+nh+tjVNvSrPqv9QQLwRQDUj4dyd7
4HN3sokwjVDQzidKVnKOca9ChRsocJTXACbmnaH01pMjVxo3tG8uhOQ92qWqY8Qv
VXiO06y3/OuyyDSNeOxse0wiW1GaAspll6XhDo7KqxrT2oUpgLH0ahwdf3Yn5VIi
kxwcmP/1n8AjRjahyzenRJpH0vWImRkfuG8lxi0Y7F1IXwhewv5vtkupztRY9ITF
SWhsjxCoY7/yzVmwNqDv9Z6lW94YBB+HPYGOJMFEDIwooI/sy9yKEKuMLx2ijGdE
KZe61u76jb7I9jvCo+tBSExGCF4Klbm3bJbY+9AIqoW0Wdw67QdX/fXz2qCVCSnd
7fDi3UJQXbqpEIRM6nTITyRN1u2aqIpvHiR3WXGteGbQ56zg5mpRhRI0AMpkKJkb
Nc5LA1PXugx1V2ddGP4dH690KDOd2DTGhIAmbjucVAQeDaMvV/4VRpP5XUX0nWcj
VDXTLj90VWiVs5mLnfgoFxTOKxt4/cSrpMeq6bZ/ZfXU9Z9XQbPAoX4iqz/pXsWG
E0mOPfxbLZX8GWGGf4NI0rABEKGfFQn6AvnBuCk8SurZLzQLdZL/ufr7p30sNR03
KbjcVWDnrdaopZ05zK/93md74fGQwtkiMeoJDYqL3VlhCDqMatwMsvSoFDGUf8Hh
T7J3IrJeQbRtgaOcV2fs6YillNJb/6T9w7HkJ2urEGQsOl/h9ZVjuGPs3UXcAUwW
nBMfFBFIZYRPuLBpHgVAXYGDtm9L/cbIL6McFfUsW3TUjND3IYjUg7m7IQhaUfxH
Zqlv5GTxazuTtUB0Mfag7zGestfLiQIKGhfliXfvRt13X+NwBT+gfVFzDMIiYlWT
RyejW576mbV334XZoUpFAOAfbUtFChTB2s+k4tXgU5P7IAtkqznS0vwCAV+u1Dzn
awWe7YvflKKB+JNx847iK/VWHWgoSGbjV/LA3sih+4VMmSuU+55JRQRiXGWlBpOr
C3LtFC6IBYCt2b7ENg1Ghb08iT8onCvXbagQfN8uS1g4LmYu2M06hGtAcdqk6ahr
pQmZmPypAz0YrU0bWfHk8uk4l8acRqzHr0JbhTKhk4Qobb8E3P5XPva5Q5XavveJ
LbehnRjbuILCn9xudpc5jFuzux11+pjo7A/vO2Rl9SZVvbxr01zmJ8Pmq7zstkLo
YH1oSvCR+j9Nmq3tdLMNphVQ90mBHxnmxc0xXmNQmkJBbfdZRkBfUVlwGlKQ3Iai
2YQ3oVTKMDWWZ4YKVeJz0c2ZEXXF0LMomz9+4/fCuJzwMO5P9lzAiOq2Kxfnbf/t
GdJPg5tJ0UT/dK/isBYLmb2MW8qh3bJmttk++NYLhp99ZzofKbNSb7HTaiTkJ8g/
6DNhuf2+ea4QXI/qYa778Zve6dRXNvc45+RMTE/Spr5SZzYe2dCACTEbkwK0SC/Y
IpYb516y29k5WaMH2mwxd2sSuNu5K7LAo8APEFtmEv3Yd6wtdCjHE6ug78P2xJ/J
MAmksPshOOO6LOukp7NGAbnCTQkSdq6F0bMW3/QK2602IO9aUfGdNL/U5CwNOMEc
wkN7gyGrJUWhlpC8OynOacQdoCT8v/yXTHtoeoS4GGIV4RHFj+oGqA0gAB6y6vQN
qOyEtbzEqlbX4BSQ3VoKL6XvgncBwhcrLHkorVZxPTvcjuGVbOPWrhfBd5ngapct
aJPf5t9ugkyUyQ+/ipwmsdTl/XqMQAyZjBEDVAG7/N7rYIuJpelg1ydVKT+uETKY
j7tTxDsIfgt0i241iSkS4xwMS/f2k+FyebmiBfqCjFEu4+NvvxhQTCYHCxjbBdwI
COGvmzmoEfqM/B1GtxttluqYz67eWhKOGGMG8LlQPsGaMMFYvPqHIIMa/7czV8fH
q3CtgzyJeLbI0+fNs6P2Vj/NgMi1p2EvuUM+g517SsJFpM9x4adOAg4PpAZMybCd
e9aAvI/XY4pE+3i2nkv87m1vjRcmhMwGtdFP+QGWUH1ZlT+yj/NxwaAXkjISz5iJ
NoCsFOBAm2ZlDri7LiJnyCHy9PpgLvmm8eWIaSqvNdx02wyFy7ptNwkzFiAfrtfT
jzTL+BYRNJLe/ukDzyPCmjjaOwaDYje9ByD+IyZgWAS7yMHd/f9bNHhzy6NDyMOl
yJjBgHET+IQIAyWXnDbATy9pYsZN5OP7+V3jpbmECBX8HDTZe7NR4qNFIug1e8nF
ryb+aM4WUsumVc6vvJblP+OoCn9lePGpoGLVMhDqc3hcrhWzWq1yV9E7/UmtRei/
UkRou2CkFfFQ/VW9na3uGOYMbvOnyjoGRdzq+hms994P95e6JiCLDTYRSplsC5AZ
TzLKnJSBGOobkta82+AAH5tAaykNFagv2N7dzg/lqTSUIzDlQHUbtO9UkB5GroVk
SloY7fFnFo6aRLijExkBvJhwuKq+On+4c/U6qY1NwL/RkFUOWX6C3YbmecjQIDeI
1UID4DyW2DaAcdn9MJ4zZlac2+zBNDLKzk78Jfl0L/ls+t59/OmzL0b2U4kL69U6
INUNZiU5wuIG7a2FsbEiRANK4VUGENme9pW5YvFa9YFbrlqahSsGaKFga7cerjFF
NLRrEC/QHjDChDDhnpL7xTkgbhWvLKGlXxUNf7YK9fNkIMhs8WlHGO+BWKQaPsHd
hdFkcIZo8r81LgZpIcrtijqiW6wdWkQKe/lM0mBJoeZLSctIF4J1k8XVjGQjcR+U
KxwU3JKbW+9ypRiaK8DfcFECL+GnUTEAU5S0veo8a3ND/GAdcTN0iXkBNN0ePD0O
Yp53RACp/+0TKFI7W/rji4s22oOPJmOC/1jOAjreHSGlXf8m4a+LSSIJd80yZ8sw
fCkcuftODDCqEnlvSEEdtr+F85lukfFRMj//oTTUO8e56Ee0fyd4JgKx8hD2HDE7
CrKf7QBL7xPOoVsliNTR8v9AGWunzcxtkkYR8teNQjQYLXZ8pkJRRpUMvbNdxXxd
UJfkV0+0UR8GpHIeGkXq6uVam/t15SeaSP3/mqgGEZwBhjZHxgCGohtf0PfHHgSC
xCOceVcv/CSKMJKMXUBhs3wQ/Auub0McIB6XZYie5o6Ep9e+u1NhdF+/ZirneuTe
oa7bviObGGAXXe9fNZuDdJWJ2uQNTgjAggrMTZZ6EVpkqbqv2iBhYsg3S8k1C+un
8cCcE805bD9yJjVKyaV/xYNiZ5cCZVe0Fbc17Y6OUBSBfwB61xuoV2D31ooWl05J
7bwPTGdsXqHeAtupZcfyUGvdVjULS7xRrlNPS+FEIq36eo/Q1Dyg2i0IzyCrRfD9
+Px7dc/XllgMMO/0A9W4C8QGUXSvlC0Aq2u0yilY1Tgu2kR5X+7I0mb3h0VBuIDA
o22gX+ppscNvYD3BprsSPVx46fez83mv/Q8V0JzseJP9t6J7U0lGFPJmVOZvOT15
D+yNjNJhPGtg08r4b9LiMdd6QTQSzmwie1jFE3Gb5ZeVj7oEXFUqXkHyMKHfGlab
X2d9RDnSJkYSB3AV/zJMm4THb3CjA9yELskS/hw+QRyYE64avzQWrUtdrfggIWjW
vtqgwwnxpt7nvxYyV26Zj3r7yDRCFrX9PodKTcI0zYnLnIbhpcaJEsMbpWI44mPa
VsKPeLAKU5gQLegqlGm8Pmu53uO0AyYt+5IRVPn15Q9AmAkXXENMe+vIp8vDjJWW
nQSoh/TeHy9t5kFOeMvTAJPaFcp0fBxAxTxtmAzNzP4D9FQ+Lk9Xj+cQ4SiqAAsG
mbbHZHy7SzER1LG3KVhXZr+QY66koPRWQavNiSLDD5WMSWhPJUQO9oDBuLbbH23R
GQciQ0zrZwqZwoit1v6E8Zt+/TWUxGrrUoHg6mNJp2u9oz6R6H4sB5KO/HDTQ1pL
/ElpFDj7AJbt3It8eShlzCYbjWm9ycjgf7J5aBdOioY2o9HN9J88AU4REVpjuXnn
e14xNyMaMhBNtYcG1naif8zYeXu9Fyj3vPb7knM1gRzVviIUZB/y0T2h8VArqZci
p6xvXsP4JGs33OhiGwHF68nLmJwfYbHgzLrcrRC+sCDN4rqND0FG7LD2Gp2NGV75
NL1DOQq/vFQm2NVp10YV8GwuC70vbo3tR/yEyOrm922C4Z6j2NdEEx9Z0AuTyM39
d4cN5VRMAioJRQiqDQI8DvZHlrXMp9spIlRQLH7BLYeRxem8hAS257iHlg2R95zb
cvG5V1QLzqY9NrSIdiQqmtPmurEaNMfQJEjxJVCDORMHE0yd/Uo/Jds6j3ehsayy
ThAdr+7/7xnTHPJ0pmlVFABivQYkF/hegntQ+RA9j5RYaDFBE/zjy0K80tQ89ZJe
rmoJ3QiqPCyaZ09IGsoJYfy+Q6Oc90iBhMHcTZ+yyIdQkrdcXVl9JCfTrJTmzJ99
+mgOEqzyqG0mP65xeFNyatW4Trc9y2DUv1kIyjdg4cz9qAZr7Zk8m45wcN1SeqLK
/Uuxumo1w1flAVuQvfMZipZWId28cmp9N1WizR7MuTdUXalJc2vzXATCDU+LxEUm
Fxn/pfOpKm+l7exOqVW14V+4CbgqjkxUuLDqoRg4N7fDZsLXqJjzRKKU0EiDDqqz
DDpZGtz0t1ZwSgBoaK1GS0T6UN88FDKEUL6bc8NfEq7pwD2qtr6Dlq6zPd5lknWQ
rBDQyo90Rinq8ktheRNr3kOk9SkoNv8HggxsKi7evz9y1Jo4pWoKXefv0IIn/mE6
0Fz6PklJKkkMqk0h/a50/UwQFROY0qFFBITvyRiVQLJcouXh4eaxxP2qa9NR/Pl5
0SzCmj1Vq9TzRukeByyJH+sre8N9aLBHUvvU1RW+UlFulFdVWfdLiqdRATb1BV5Q
sleO7UcnB77SQN90gBX2LSDwJciCmjMSYvfnLkrpXniFAAjP9fQHFPeqthrLedhl
yQqNzsGIbOv8oNz/5TzWv7koKv9i1rFVIwmDk8WV2KuhnROjA8J+PWwwCBcCL+FG
Ev75EfVy4XOIvOCqU8nl2LjM5qebBmGHdRn215U2Zdjrwwi83bo3wLXtQpKa9iMv
khizJLViePYZK78QLd8qvD0XStESQl0/a9FjSEP8p810h58pEb4OdBl8RrH1J9S0
6h+3fpiP60JuT31m4v8KmK9gTePhxPkYAUBDRfjiVuqmJdAANsUr/EX5YpDx7JHl
iGzNzpnow1G+kMjtWaX1lPnZlK9t3SCkTlhF06V4pl61hCry4CZOQgPCpchQlnbg
2Q0EZY2RXurLQ4yedHyVS0FTq+bXOZO0IHkVMPJ7m/R3e54JvIMQlWOe4dO+ArHK
F9pypjIVIKTzUVOsX8DEzXPVGYOHw8dgC9zgIeKp7+xSKDZEk16sDIGnvgzGzemc
RKwAlbSXqS8eZBesGtEevXsBWDZ+IyFpjhiVYRkEPfid+D98AKuhf7TV+gWSl0xg
8RtbKp24LRry1w6SUDkT2m68LUZvJASfLOa9Vc44pFqGjd1JKZKr5CslVdJRD8iu
QrsVtphWTULZqF7f9rW2nAMPM3bX/dejbBCtKJYcmJ1H44waNiGlD864c5vGdc2k
1l4kUbnKlhSipszfKeKkkXCShNi67FK5mUGGY2QgeBK0JsWGrGUAnNpwSCxVXWa6
o7jAvSd/OA3ge5Pe/6VsU+kwYZKhunSD32ENTrq+Fj7rCTNYAyxLMoswOM2lcPRN
DM40+IjVUyi2QhQaE4/UJrMqGQe7GzRnnRoDWzbdJjfV8Y3CTxrs8xhaOfmMkA8e
eppunkkXJXbLXIA0HEDVSJ3lkKnENuwX9IYmOEUbH7/XH42oK0lT4hgaNZltsHdV
r1XSm/z3Y03iB/HVGMl70UbyPOOc/NitwZFm6LUT8JSS3tsSxsYxyJ8ELwrmsv1Q
sO+Z9dNi+MCb+kpjkMCGYrju6zpaVY6yurGzDBuv+rnaLb1Ah34U3hQZ8NuggFbN
rjmGYEAGg92qC/B6HbfmYE32NsM6C/XtdQhz5K2uMS2vQd4CTCaKaq2Hs9R0oCSb
lT097mFmTPVYAX8RatU7IEBZ9szLKXr4QECeVR5GC/kmT4SRNgHZ3CtbzQzDlzCw
rEcMD9kKR/T7tfyCk6Qei9tyWgtulVmIt0LF74fAg7+MTVJEreUhkmzf/UCVo/SX
Atj0JYsT4h2/JuxTU9QgzXBwvrAWHzHPeeOouTtbnHL9+b40r69enOzVhXJESE+o
TN94cVe0XgjW67/BYwywS+nr/3l2wWn4ZxtYnBCUkQBGfxzrhmkhhRY44ywssDMq
OlkhYBtgfpFrdlWaP40oBmms8a07a3+bK4QvZ8qsWT5hp3yo3uYLJl1aQ6/mQ6cX
p44KzkIxvpKY44DIeJUBjIlbsFGOfTlZSWNaTYraC7/3kI0z16Xol81sekYSjaCd
BHtPGVAIKfP7xftdaQGhcIlguw5X+HO1DY/0rxT7SYH9MevGsMFSrAcBgJLW1vnr
DWmzzunqTLplemg7Y/9rdelKaqr35mig5B0157swuWB3l+tDAPFZNz0yC+npSItn
txmslpOZD8iGUJ3QataiCj2VuP3/7MuCrx2SPECVyc6jvN5Wr2GtOSlrYFAOSlaM
3sWm1Bc320iWMAQxzIkLOlg1gaahBla/l+bbzY5n7WuBXn7/43j3PjujT6jbdAgs
enmG9CnHQLw+rf5hUQR7hI+rIfOc9M/s3m1JuWgnoqoj2dBcfUIRHNKjO3vADDJt
TCojYuC9I/6zzV0WfLd8MnB7HWN9V+JWMc/PYLmPN97rZbTLjBu1hLzlqNrkYYkf
tIMbCdXwA62zp126/JAa/SYkWrJZ0TT3DCe+cnn6mJ7GyeRl7NS/XR4jH8NNhevq
3ggk5stWf33IBMniGzzMnC7H8tIfCDmhwcNsOh3MZmlVO4c2J7HX3vMbep1pWetD
lFEdrb3O/uGIDgVYxpUdS3CiQx/nBDHisR5Iudet1vUMFlYfnRioi6BmVmH9dWp+
eIwJzXNq4RHjVz7NRoeoC0jHGCSw77FsROYyOfFNMFQg1IuEI9Nr+99NyPEIaiNb
RsnRUVGzK1H7kbmnKUJ4uoABwvCS3Kzq2tEAc+BhjVpuiKb+h5c3jESvJbvNtuJ1
aRhVW8/zk4qDKXs4kV/TZrczwqZxx+ir7gnDDZf9hzi42Iucvs7VUyjVlSOFg1V1
qqxDDHaWbdIvGpOzUgyq5Dq/su7KktjBHUMlMneGuQVIvavEgWL+rbDESQWYbsGB
ac09hLI2GIyI1egWdSIHopfL2UpXVz4BBDhszm7MELP8cO7BBtzdMqYfAdujozDJ
oCIqz1MeIpj7iuijzI2F2x0ABjgrfQ2itxcjhK6Bodr56agC1xYbz58vEAM9cAfN
GumtX2uAHmu/hfVROnuP6N1KxuXXeUQ+LQ0HdTrkcaj5ajV/7NRF/1aCPlB1Wbmy
ipnUPwvgLJQ8Jk+/VtNDznAYEnrJzCT92+JbbTBWrzPvc/aWi0w/yWSjXLYNNAzd
WdgGWGTihuU8QEz0y+ZfA//20uT+UibrZQBYqhbKx51jM5qsRGS4PXWbVBs4sqCC
db5okCSrH8/oXrsg0X3kiq+F6eTvkLXyMrdurNvxzRYpOw7dIUUjZqev0eoUj+UB
moG1NL3BJuNLc6gb0IMWldVdg9b+vct+Tm7Q85HE5MiYNP9X0WGgxmLtva954lCv
Jtw4x9niuSG8jNdubqdb36o4aZo5xmCNCXESqfpMdvf+DdRDALC5JJXt6FYAc81h
xgOIiJFKNUC7t2WFAMLlGHQVXPhrN+co8DrlDyFBbWxa8UCzVarSU78blvHSmzih
Sn82vvmZCRHgXv6tj3aX962Td6VkEaePLI4g8b4fvARqR7LmyprWtgK0Eeh2Pze2
S4rs9eRjCuxSV5IrifYge1bC7P+k44TICr7+YKqVBV1clIkJkX8dDDMD09w2YqGr
vEHg21G7+xNiQ7f7EfJ0Ot5Yz7HCgUkBPQq/jVvJFtBIZVuaywvDU/3tbJawxPMl
onzC7JEHv+H9VrqNd3nqaEb8xYBuZIMECt2Rk8Z+yleEWdwzypXj43aU0abltHIP
58W6PiD49ZLr68BEtw+231+J+5EIama6icNuWVeIx6kpvid6MBsJiqL3obX1OUhE
RFdDPL0iD6QIWTSjfkvwVMXHsKVFPJXgN4fdPupYD3PPfakPSiScNagraeoMCzpu
Dd4zbzlJXwOYTinZi8KcVw54owNZ3//YSx3Xq4KyeqfzjZNnAmFeGzo3s8XGyvou
ztWltWyP3Lqf8KGpRwltxZemqG0fQ9JfGFZOvcBLCnEvBIoYXKkP6UIcc3TYrPqG
RDDF3ECEwz5R6zMAqcIiUKt48//SPis3ifPTFKqEPz6NqkC+FDkZeiA7TRwYfhEd
xd8pFEwCwFF9wYoNZgdfGWQeCtKPxEoE7E52H06/RsGzp4qOk5ef3HSnmmXt66zO
Xcr8lsEux9zO+sljoBWxXS5yyONgsUNbmy4rR5gY+T25UKh3PzxygPvpN2hqm7wX
quTVeQy8B6MARFAU+iNLQAJw43GwXoJb8UGhUIRxtXXKctcIkOpx2/eQm8qWDI8n
qr5BF/xBgzN54vsHP+mclPsrwxwLOLplbwEak0KQ4QtKKsWml+0+PEj5vaDBSFhK
ThAGTQ6yZeLW/Y/JeJKZ087wLM5TQsccyvR93tWbbMVcPTfsGOssqx8BGHl+idio
8Z+Ungc4cbRL8jG1ilV6FDRb9bhsUmNF5Ofpd6h5WmA3D1ItVcdcLfHL8+vyIdZy
2LVntz08ZCfeRo//YlmqFZak3BpBAnUewW8gPadhLQCGqkcaDbC37jmrVdGlATlX
qf/MRxelM5e+NcWNiFvzCj30fkyI2/8ciclAk53talxDtVGOJ5ZBdc4KnSbdkYv/
TJsjkpF9jfynZGuQoYKXQphlfEwC6HlIDlHv9x+xJkiQLML/U9uQg5oRmqfI5jAB
wyiXylAYX49cwYUJbH22R6MjkY7JJeUoA3wrgpkQBkrx9CleTZzk3P3sOVdDBUvT
/RKx50ART6D/BZfG1S00d6PK7AJA/dBK8nxUmIzHSN5lF2Dajm6n15tby9yqXySW
ipRNJhXp79uMFl3nWaD9hFZ3sRKbCV2piB/j/06ZPVZqRmUdNZC5KO2YgLnr245S
Z3I+A9OywJrMn1Uo9aI76PAVGMSJCfkV7uVKwUrL7txw51aoXyMOiD0XVQBnxU0g
UjXKW/m/Tl8nSNcRY70fBr1Yge6tTnD5RJuXvIDJfrIT/sEvXketPcgbNcX0YXGo
Zms81qJ5L4TOdPVKyd8b5rQU0tnuO16QP4bP7vm9pzxWPiwVUkpMsLrCQHsykVm7
RqMeFx09YmEDn+PO2al4kAAn1PnIUkKSgpVbA0iEJs2D3VSkNOR1jTLhsnIMKWFA
jnbJ2b4PvX0s9qp5I1gVe4w636oyY9a4MgWIO07k0v17gJFu6/o0MxY2MHmeI5p/
tRdh/gc2Gr82BqKDXsgtccgGZll69KsFMfJhSBwMkjlEuqjCDI4tWAlUPqUTClxk
zkm/q+5QHdmjwYXp/U2x8PoVpR5j4k5XI/volaOlZ3Sp6GNvCHfJdFIAloKPyv0q
Jjd+T0Fo2s4FhbsueXR+5rCQNjlXND4r0hPeLVxHzzNlMECIKt27g3cr5lMjickb
tPOLGhesyVg5e1MpuIafLa0WK142sn+Z8s+95nlXBYdFQOgoiKgFK1sT47pBsG+8
3r0YbrwtYzCy1EAyd1CxyL+u+bbJTFzucmAIDc7IV8OQ1NB+/XWUWPO8GrXFGiip
6jZ0VAFksZ8i+GY+BrXibTQUxke6PsQ/5v9c53fOnOCpHoOP6Oq6jEFfuGGw5pzG
jct6ZoMnAzD5cDomwCYzk6CIm3kWDGgJ/FTSR9Nl4tMouEGdfHKTsaSEhw6u8jze
KqvZJToqeEuyctmEcfYOSgJscd563K+6PxWZjl4Y4ZTrbOGC0ils3NmBUo2wgRhq
8j3JcRe6bnaVoan9vGVKjjG+m5PZjQlsMnMa0SspCyaGfDZ/7MHpm6E5tJFIqTT7
LQqS/XfHnPbuVz+wjC7dPCbPD/Q9m7FTh9K2leR2j+h/oWPCbM0jYJVsl9UBvZQN
tbRzt+hC7NSjwO3tR0fvb5PQMsbfw1acRWbaPnvGzXrnsNlcoM3w8yXJ9rETrSEc
JP5XN2LuESkHKkxUaBwGTEKTtDPlJbZvV8IK/PyFFdH7TBIDn+VYZ2VQP1eIEkGW
NkRN+2C0dDJdLhtle6u1Ed1k54SP5dBLzuK7bLhjEp+idTeuILsrp6TJBOV9Ubkc
T0ZBiz+4PWVo7DvaR8FkTCaE1TmU7akVNAOOn1kwlOMOJY87l4iPC24eF/zAodCH
dOMSBKltOyc1LVUIA+SvJytq4V1GfEl3gd6XSAn+sS3Sh2HXZaH3pz4WR6P2i9s7
aky1me8CBXsfv2V+veoM9sagJnrAjdIDoKrlH3mMvtGat7gFwP6rRgBy0ZQUUzEV
sRMQhd+fjpOGR1vltr2vvgtrgGPY0wEwlEhcov0tjYTwqDRCll8wkZD1zqlSTyLj
OSBIQdsAvl/sUYeGjbirbVBcATw6Stlh+/gQYtNlYlMZf+eu5STNSdAArFYbJhX5
rlxOrNydzeTHFoGRuDURjJITHReEybKW4koUhiQ4rxZVQENq//O97bZ4R517N+Rm
xpJV1tXMc9pAWp8nhMJ7O5GTEJjMzaQiNxowKGAoea3OUNjCE63gfoUyUeWmmOIc
xwqS1Fltm7Aa0L42iFMrsJZTTO7LdNNjwWzv/Yer8CZBE38s6RRPzIzJmxqvWVNj
yJyoq/lQ2dV45UfbyukJdLvP2H91D8FnBWZhLhNBe7qgbesQCRDKEGMH8TSKqf7j
kLalGlGOnKLOafs/OkEr0E8g/2ZYvYsMAQNvcGhdoEeYeq57I8AJsJRu80/ZczAY
DLXWkCVgEVaYyFzNnwuht5fWPMtUh7wQ+H/U9mCOfHcacachg0AuXUKhwbAtG8xk
PV+2I6amtcuNPl9IjWCJUQqAlIwnep1O4T9VdzjltdNqLjyIDSrhaYq97svS4ZP9
v8ZMC0o92ZietlOFv0t/5v7bOaui8b6qlIBVRCdNY2QzZ2BZo507ttaK2yJPjBKO
nK63jjkk4ZSpiB4ybHltXyIIcXfa3DtQ1EqgdkZFT860fkoZ2QshM0BA6oyLS5Zb
ZNZZdiHu2ZQ1Hw4p1AyRtxKpA4J2a1o3UcVeoUBPh1bzxyaDW7AUqIT06tH7U0Xo
xOEX1yF0ZVFg6s6G4zkXbKC4dPHPGJzMX4D93GPEtuc8INSWWimRTaRcyIc1FJAQ
Wj6QhQgAp4eq1WZQctxkCP1s4yMJeVba/QMPaPrdIpy5UrMtgH8VUqEJ6e3KmJjz
oBMh4W6tH7RkHuiXRj0uB4eSq7ggnONZ0GhqEsdO480RmOpJkU4nTcNFvcbbjyx4
X1/IU9vKZDypcm5z7hHP+wGymt38AeStR/bI7wzq6RAkY9Oaeo7f8VXzyZeT1C9s
U2VDD+R2lUY99hN0QxYcdFb2kqyZ9WPf2kgmEjeenU75brwLXKwysHZ1pDtuBTnT
Ltl11MUNbrSJjySkxCEuxBUyLaMHoogS2ARKwnMQFcqiMvFrkMMSiuZMB3ZrwNXb
x6Gkua/lZ6Z1axoOQVLYeUhGPf+5dramgYll783TPpiapJUg80Ea0XwqqtkP4pPw
3AV2weDQEfCribHTaoxkLJMdYhL73C7Nx5pgws7KxnY5Fm43IPXklx2EzV4qcWlE
/QPCAMPLg4Cy9n6vRS3bgb8T3t9yv+mdg/R17KqUUZTIPXg1e/e4F8mKR4vxUy2Y
o3qMba89srRNKsxGgZIwXJw0TbvWX1JzAjWF7vkZeCSHHM1LhH1Kcc627box6Srj
0GZOIqRTSwecQQ4Lluw/LShL7V8xTHjBtPEjcIYmaYwTZUmd9m45ezQ07BdkHl8m
bKUoaUvwtXeryT44dCsR96rIbieLztctRCZh1e8BDQTz+ZVI1ZlOvnI+8nBV+Q1A
xCYmJrH1EbUvmvRtfUN4fG1MuC6sjZOwITXJj1xuhPMGb+G5uAefdk/R+Xkjh8L6
dklyKRGP9N9sZ1df6jCphkcp/LE9yX5g7X5oxjZEEKEPqUrSrbcihQPYO3hDQazt
2BRx6k6rWNgBdDVdbZ+jjj272d4/zq3eXk5L2t2STgzv67moL45Z/76tYFiqSiTe
xUhYw7J5LF/JL8BJIXJSD3i/dhaMDgjvhMfviADsZa0/k1e1nyaohM4/tKTfm6Ff
43xM5FNmHm/Fnb/RX4DY57vkhvtZqQVnawRTxu6+t2Dw09rKzsjwm2sknI4nO/Un
3sS3MTeNcCeKIWRMc+1HrTXabaSEx3pTzQjTv6qEYkx5fZGaFE6JPqu7jiRcFCtK
ByVKVXbr4wvwSWdQM2Yp2ZkXE8x0NiSx9GaythkSgEltJvZdVogw5VGmxQ2aDmqR
iOXpyUNq4jZJYJR+9Y2Ujj711TnDVL9Hrzb2JAeMttKQ3SununCpakUTkawL6z9s
Vm9kYa5REuH9kLxkuQgZMIxIe+Ztte5YVpRXkjxN3PPm+uMpGaGj1Sgwz6aeKMSh
plqVuHhxRXmfaWsQygaY2Lsyy6mwNC1ARpydU+w1P8UsZb/F/TBQefdNQ+GaS/P/
zmCI4wrcwK3xGDkKoEdi7/ilbPll8BsZCBColBiraci2mBFwwjo9hUAhg7XlnyQd
0EhQtX4l6meL/JXywXl+Z2XbCqN/a9RBihmiCwhFQQ7Do3zS43l4MCDRzMg/uZTn
WC5T8xrH5rrMgAWJG+Dk3xBkYaK6g27w4aKoPaI+8LUbH0v0n08+fqeaCCpmSNJQ
Gg2rVA9l3R1iZX+JKbfJbLLUnnPvkg4KDc5srZ4ZN7zwb1+7/C1T33JeEMk2mhgB
mD+QCNUxrrMqjiyKSPSKaE7/tDnJ3hTz5gFDXDW3DkkJIOL5GScNgzDbsN0V2TzS
6cA48Mn0BTkalqHCvdSgB4tfhekqRxo/F2gw3MvHIHbMRF+/DRHMaAPPdl5dJ5kw
mROkazIQx2SofEkR+8VisdmlEnwT2yoVCHuNbKbE80powIuzPxOuALlcYQGvxE5n
cxhb8A6XYoBhSUsHvGmC77d5YFVJodSz1cK/iaaPAahTUKNtesFMGk0loLAuJuPi
vkcldBGeun9w5cYE29fbI9TYh0ySxs1byCtrzCnaekOEdsCIXXjOrb4dsKCsYHZJ
2M+BRw6dvXXn9eNpyol+5n87jmCwWS0vowap6xA+iTyz86RigrL/yctV4dgKR6ex
EqZ5VVh8kysQXVGAbv36qRsI2++nbQOcJFyaSSxT3nRrPDTonYpOtK+Jt6sbbo/6
Wi2i5lqKlLvkvrFDc8MpiD5fn+c9ykTU2ZJhxJZoLtqPJhTOz5TbXFp/Idsexmuo
E4ZEfYzcAmeucRicx1drldSauVvAn3hLDz+A+0GUDI9uNl5A9bxVL1byFNO69iKT
ZSpeViLumIbY9c+W+PsNkeikVFKfdPyIClPtIdqrDWpdJwWv9JXDnafJlGbEUXP4
Ifz9C6RunhA8ypUa5zwJ3FsKttvuEO4TlOq7jn1mUsXUnfTWgWHkYedHnIsJ4vXT
u8svG7JkFNZWTj9zH/CRbmRTUt72U9NeUW0uSliJva7dsDn1iXPpE8iWKauVWFgk
DvwhOWGeI/n6GeRTwvYaCkU5pCrpUXpCGDrgSUgXax1KJe5cNArtT69c6/RygSh9
JE1Vue2jJXu7yWaXOGLWoWOmfI/jwr4PD1KvNEv49y8ZYmhyKm6+JpsOtrSRSLoo
yqXHpER+VC9wAQUVAU1ENFp7NUlrDb56bez4PpvMz430OiYr1vqzPQ/3/L6bH48f
1dW0Gz03uF9VQlhOeZpA8ay/D/gNJlpP13VAwMZ2qiUXnRgsEEb7WyGo7MmG/I/c
Kb1tg17nGrj21uz53wPHQoIJziV/DagGoqL1VhuB3EM8Ag4tfvvq9BZhFc46Rt51
OMYkjcLOFxmQLW/bg6q6fpldzZMaAG7Tcj4oaBqEDLaoI5z5VVTRL6nSzbBcagel
uGB5AmRO+6fD0su6ntt6JGGaLMNVQitPwz+jA32V2bL9oMBjgi8annhKRfKBh4dr
u3KEbMjrOL6Z735SawwtvnST5UKj7ElGsVmCu7x1v2ri7Z3J9xZ8deTWxZAbN8Ph
uW4ef+UIEQZmcO+bPA0PwcB+ekFuc9IzLCFItNzSpZezcOvQq7zfEw5p/Iikwn69
2P7PXMoHZQ8X76jlBx++Plx2I0dKLfd0I1VnhXJu24DuRKJEMJMlbW/zian7RNTz
OBJu2sAH4zkPfuOQixHCPCzWKBwntFuFqPEKOY2a2K8ji6RHmfo7adowonWYXs+s
wuSKzS0Q0OmdcxlL+Yqdaw99hdBzj2b41ME3zHbGD32S64oVqq8rRiVYumBFUpBQ
ux1pDJfQs1Y9V3mmmHbiOTMtFR9Nk91jkDLcfBwqW3iNqyCwC21V0+AoCo8oE85N
iRlDS8K9mWTAr6HIgs3Ihbrse1b3gMY9vdIG7wZrnucWwl/S+U3PKWZFa0mXXUbl
GzpHVJzX7qiVeMdj+mnJy/jrywl7UplTzVmf3mdygIgCN2L2l1OxEu45hRLZZVxF
s+eWo+71gX7zPgWKpabYSafqNbPysOpzK7gZ4MIbT2h0G9e5QSYu2vnUPwA4+VnC
OIRMKMh78wi3jKCJxy+I3W2zfZXNcrmWQyh/17pA1tlBGS5p5uSe/XPHc37ondsR
vI25j1NVQACJZY3Gwjo+ME/YgtrzN3aMHpSHKwCOO5hdqTxJbhgHP32ciWTXyDnN
kXhDHdQe3l70sjgkyOZojMBZKjN4FWBeHz/6zPkpjZ2utK4wWSJHfYiwJVhuIP/p
iDSFdmr4Q7EqrIGE5cwm1BYoWLwhTQOZ8oNGBJoeQCmelqEsCQRYTalYaEgdVKhI
ZqVJsjMvSSa2zCI8UZzoaSYv6/HVLZii8DRbd8jUsJWygBzAQyY9E2ruSzE6frIs
vUEiKue+lnbcfvyPMwBjUzAhnV/hCGzFz8Dt/MoUqGHa0ZmLqNUfn1QvC/1hocGU
rPwE2K5EHySq+W7x/DnegXf/TEn9kH/dD6YSyiYlWbRr8eFEWnU9JoIMvguuH0nA
5txi7cMh/oaNoHveDdZFBxK0K4ikzUPXwH9hrUltQPFYcwYGWesvkdpKcj18djeg
fiubpTurzLtGy89As7HF31DOQwFGK5RcZ/JlFvTIVVa1O5TB5+0BS8Wf/TbtT5AP
bsy2hXxStizUlMgrQstM/P34JoFar79ywPPumb7oG8IDLRzoblYVP/9o+KqcHAHH
Jpm4KCqC/qs1dlcVJSqfeNWk9RjEX2bzRP7knf62W8USi29wTKUCF4hgL3gFSHLU
6NtulHeIwFuC7Qij6rI444uwYhK0rrz24/s0KMmWcFC0v7DcRzBGyZTocrDFE2Qg
4jl1xYW9Bk+5Z1yuzp3fj4gIkLX7eaGR5cqETZmObAK7KZOOcj1uIkgwUrhgYuVC
dnkbvKUhu3sHqEErsUGu+e6NTZXDfdjcaGk4NOWRPsF4J++dq5K80y6ssJ1TnKpV
gMZcgFgwxY4BXcbIU+Vv9xY9cYVWf04pTvmnAjnP/eLjV0zNnCsVkKaYFL/r0yLi
cUftQkLcQ5v/MhQ9KkIsZhTSFsLlzX1/7BCWgnA4A3roiC3WXQ3bDtNCT/caPdhG
EmqGaKeLX3QejSoD0JCwuvqJ63FRpTUrNAbatWgtbZ56MVEmoS8UuCLmDo01nqkl
EJVbzIeL0TBThPYTtUSQ3z+UJdZBLhDhB0BU40q5jc8SsGsIip7tYyPYEMpAHPyT
GHhxMcV9/8DYbD/x7tMi9OOggj89iBM1XgHF8KqKG1WxPm52Dv+ePHW+olrB9wk1
DsoibTTRVQnq+jZ+6aGwx9hJ+mCrhTt1Bp61ERkpZ+M0Ct1Jk69jSGLASHq+sbq6
vwz4kHdLS0Xbb1ESSoXib80wI92uz1PddAoWtrhevfoGjsKY2qKd4sbWkvjbPUpC
2qJb6vEQ0AtL8w5sqRVAjuyJBlsw1tq/yP1fUGGHgfKaFHG4+vS1e6OF7c100cO1
5p5jmv8E+u1kHuUIfzEysLA9xA8gsyVce+OqkZXeL4dXuFXLg6AVN53bD58mURQi
wV2Nywe4OAqo6nVNNrpQJl3kXRCRkuCLflETDaUJLBHaY/JytfAKaE8AATjv1482
/JTar4NmsuacMv/iDZzNpPaivwB3BEH0p0WRrfPBTl8+yUFh1+ZfmbttLkUSF6wF
01KQMQYEDG6hKAgL/ySNibnSokoUGglDs/8XJErPs0VOTY0crHmCVfvc484VGuMg
lS6G1Yvb7bzWnIEdMs2MWvjaYqvNdR3Re6j92F+JWH79k61D2EZPUlAr3GZ3jS6I
elKjOEPXxYSQOlmjQhtF7Jw6Sx2B2soVQIelQiBmMRrRYYXx5xJmayDY4m+loWHf
u7K80MC1BVSX7Qzz5SYzjBi2a7GRgtEb2VjU79eSKATi8pnc+Oa6s79NvZMfUgkG
NQPQN3bJDvOnxpClDTsnarl94owW1MPKUx2UznLx3CJapSwCxVkpgQjGV9z8sPOT
AP8WJHQ5brfMIljYIBeeJCMT6PTX9DvY387oi+FSAfoSfBBhLdtdJATvDtRDacGm
Y/w9x4k9wBoDwBBgQnKgc/66Kqz0eNmPx9Jcua9V2t5xp5PI+p/S11qoT2oYx847
terwmxeFqilQKyMAbF1dvwr8LikTJ66HGCH8c/zBl3M0wyPsHd/90n01vSuPWDjA
vgLwKosyhWMwqfNE2/r5C15X7zr3hTQhuOvOuJpBpXvXIKZZrF3ndQtf6WLE8WzE
XcEB2CqmI8lbJ3UQuKuzKodOt9ZZ/kkVFVEFE1atliSuxKF1e6IxKsBjeSX9YDpF
4/IHih7ir7ZmmqxABp7waEqRLYalmoHjqk8o/whO5Ri0JRQCM/f3lOHfFkyKZkrx
dsEpUdawN9s9G1rmCNe6O0P3ax6u/rYvTQhtpIV9BBCEaYJR9Sifb6HGPsg7Xh6S
yYG4Togk23vE1ilpwWKUXEQ9VbpTc5ylGrtXR1voxNFZpmsxTHTrfRKsloNeoZSK
AqBqQumtDFkUOrsJ5T6TeC23rvpyv7x1aXSB/YccPejItld9nBheB9nBUo5to+D/
uocqMwEsxK4IrDIDU57omIkD5fBkosJhggks5P4SlAlVRrVPVHluTk21+R9xutEY
+7RZE9BGeGdxlMFAVc2o4/c/EzCZ9W+MfXj8tpvyviHUh7WFEHBmFZHV6OESW/K5
mwK9J7LI05xMvL1N31djSbrQeB2bAYcES3L3FZLCQo/ZD1FCtTB0GXkpMo8ZUm5X
bD+rIZ/63M8RySbiRqVCIuoLCYnaF17t3pA/W0r1kLk1bNym+Oh9ncINimzAiYsi
mX50J/Fz+jsXJ6TLwERCUTEenelGNSdL5hGhZuXcU/WrVOMoc/VhV50qDwq9+a6x
m0OWNlFCJTS/b+RNCS4t2PpIpo6U8U5mhMNaLR1czogU2DAC8KlUsbP00PFXyhT3
XUM6uKJLImvBhVxdQkV/OVl3vZ8J2aYniITX/T8HQiteIdT9/cueAfIKu1DCbaF1
t2gxvH4bIST8kWCTQL6We2etJ0KRi+3OF5pIeS4zwPzBoRlkFMKYXxh90kByLAVy
Co5QutX30lkhNF/s9T5JOjbq31CJ7zuTKJr53yO2Qo9Z0eaRaEaH4JtLwWmlDq8W
6kHVwSry37XZC4pFedgz6ccr+9wH8HTpSUGZHVF1yIN/9q36inBo+2qgbS98BFjg
i7aS5Yik7h5q9HqUtWxsmkPJ5Znaflr6zZ/dqWBog6MN8iy/Qj05xoAE1kZndt83
fAksspMtEk2s1lbjZvBivC/WzfPZlAaPxhhsepUTu56nYghs9yOpjng8EYv0bqC3
0DY8hbHxq+b7hDrG0McQl9Wna7TPbh7u23iXVptHV0Jjr+dN5SDEDYfZP7A8RY7Q
yWUxmhqpr9P+uhYvIYjMoHRwnMuC6MldZoQlfdXU4y5nWNLQ3XQmkH32nKnE+bOR
AO9p1wWYmivr8GFIkzL1CDsUTjoknaGWVdfvIQ0CfzUbt/S/6US/ZEm2QUCHcTTV
apw/NLBzP8OP//X29meUTmJKbPyL/WWj0GDxzFvCHirdMj/F15n1UZLG6IBFP1et
jGxmdXrtPP8N/qm4C0YT77LQM4Hf82BJgNaub2GXlfCRowPuvEzjTJzBaKejvtbW
kaueKmyjdkEBGtEX+cDRoBken+6HjEsNw2L40kHrWqUqIH1s/sP3NhPlJUIX0To/
0d7LBuRH3yy6NQ/RYvX2XOyY0BXtIqq25aMtAL2YVvCaS6X6qoMeFMVQedsXxALo
sQnMevqxZ/IkmJQnZSLk8e+Xb3MKjAJq8W48zGQpHi0xL1EhejGxns4FX5OhpwuY
2C3bIc/kaHt8CzUIqogTVSFHIhpbpHnr3MB+/dndUbBN7HadK7pLe1g1LapNpIzm
raeBPgKziXEIy+aE/EK9HRe3Cy0FGS8f9XBR9HnWsdiBsUG3DFSFBYbIDOfdazfk
bZ63kNhmSP/fNNklFuM2rdeyawfd0wVVtu6fHmBtbBWKcdGn50uDyBo2igSz4te/
+3XA39C/ZWgE+E4r8or4vx6BGmgmV5YKPTvyhJFBuXo6p4KolQ9jOKkfUlXvF8YY
RIzFa9vHXmmXPou9sqaqW7yd2BrmCeqAMiEwWRRYilpjNX+MJQxIwvDDgjZ+2I91
t8Wnv/PVAa+iJQBpOfIPzSRacxyjr0vpMhXpChipP74N8nidUEvv9zixFWNMXE4D
0OpAtGL7f+0btyfuz+jmEhJO9ndaw/FnoFhRoIWzdsR3tnXXVwwvhndcXz6nXklr
os07eWOrakQMGB+5lAFlQZLEBMMhXSCy/SVAh3lY0ikfYZb0TjbEw1lZMGBNHOhi
lzOkogd53ZyS0fGu4ueUpw68x2u+uttNMl82ql0+Sh/XP4XekQ3i/4/L/XBdPljD
LXb6bbQAU4Jy5GSEkcDXHyJ1lBubi7M/jYnL/asTFLN5+UOxCrF4E6CUynVd5qiE
4MtqfPA8kNFhIx8LU17oJkpwjGtVCJX8Wm64WW/LXahmqDjOvkn4KEFCLKdtqOch
eD+ia07k8kFjwCybRq/08ozDqR4E5/+iaNSHgL+ea3aieWCGotFddy4QwZcEiVDn
FORXCkOfRrkji9jVLs4Rev8o1p3K+dsrPWUJaDXV/Nh+kdjnbeQMP8A/5J9z5gLD
hMDluyPZ/9ShlfhGs9PjKzYDJO0H5E+RqeICa9TrSvAV4EY8CEY4qDoJNKyWgGHP
FO/Acx0577DmAIP5lAVeqLkBvG+KW/BWwx4ofudITwrG3gRud7dcI2rKkRcBUC/U
PfB9FPanlyXOfgEse5w419Ctsry0aJASb4jDVS7M/qZQ1pGHA++MS8uFBjYC1KhI
ipTh5hl1pc3eCB8E4gkiN1YtYj9V8twf6e63naYqb+4tUy3qbFmMjf3EOGA0Tnvp
XPR3kDKiizo22X6m7y7qFyf4JGxZGvQNDssipImeJERd+yuxLGedfXbwlpZdm99t
ACv83fVAMOKTLww7qw7gcPwSKqlYSwQhfIIFto00mRV/STUReXCckmeqNc5fqEn4
Pkcc9BcdL0qeGWAlHjHPV0zKp6E2ji8TsBuapUAEuMv2qyq8+Ps/MemTCbkQfXyz
D44mymS+gLmCxk8aFdk50QzUsqDl0Sa8RV4KxanuQ+YsSryOTDvPA5qtojknY4fk
bXthfeMmTUqGV0rHUHypOQlNFYETmCdcbuRjHYt+eJ2kmUqPx80ARwjvzq/cbcWE
492uWMUe++6tCgNZ1MyZ9XoNbdq7aQaXHnPNbGXAdVug/KtsMeDFdUCodBku3yMq
M2HpnqgO4VLh9shydvPSCAVpCUSTmXv5Z73hzRYucnyEHa8LhXXoK9C29coy2tAl
+YfYYN8iONf7KpPRVE9Q26kEKSCxWy7iYPmTxkxcJok9juXlf1TnS8E146+Lmu7e
CxlQsI6lIYUg0xEUanEZ078VvLPH89anfwZ67d2hVRA2FSmti9x7awXnWTDjswhj
UjzOJ9ZLjAyOurYymDcpkSAaA/tjm++cn+WA+tIlsX0/nSufdwpyqEqvfrERkfDw
nYWEcDRAuWKaVw4Jk5VgAZr7Ah3jO/2mlv9cpy9BiCdoOuQYt1UC3LXl+wcVhCus
VrvHT5am3+EFrc/Es5A9vmjwvaNT//Vlo8k64cjMfBtkYB41YFlDUoUx14mFvum8
+HwAGLbLRZyoseFMkBDEBgiYqfsguHdTXLCbl30MmmF1Ju8jCjK7A8JnbzegUbxK
njFzvJIGBSxpnnJIBpwCxFF0kWzPZCl0WKP1om1uFppTnB7mOSQboYUuj3yzA5kh
gQ5Xi/KJgk+zibe3HcRs+ELtgY/zfT96ij9OV52fORNFX/L9aZrIlG0RGS35JhYO
mPiZ9rnYsNHzsZBvqXR2XbW3oIOqwNwHOvpZDj4VHupHVX4Caq87nFVKTPY8eA9M
3P021b0T6yWMogYDbOPs5zCJia/RacNkq2LSGJlxT+Bg1WTPEZepC5fyMGyjthm7
fLLgH+zitfMOR2B/vc2XAiyqqLUEkyVFmGQw402EZkllToCI2BjJ60cOnymrLNLL
hV8Ig8es+E3Hb/pK8J0KDDFIZadF5wP5+70tMEnqoiimlAQcodmBtodqVHeO9fzW
OcgxChJFRQGgjV5iKsqaQshoGgzQxODDhNiTRmCj4K2zr8xAHuqM2/spSs06hfhm
Sewj3oDCu4nFJYx1KuiZ5bFisj7NwglK/03X2lzhT5rE1OEqORzcRCX/OQ0R7A0/
dwdErprAmdoX4RG0e4W7gw+N9WN51I+fKcGhplExX4G6A7pj/Z/h9j6WvmWFuCrl
6W2gskWdtAdYGcoYgAwNbdKz0YnyDdBpK2uC0a82ZDVe4FQwzbKvEH5Ugz4NHVZ0
VIfz134V6mv5NryldFJF2AmbhvtWKFBOTShNmNLRVub0NBYWwq65Gu9VLzBN+Asp
gfWiRlm8pCCS7y62V/fyTazSWRaktSWkMTGvlihrBMMDxR2SuDsPhaDmNPtV+xWO
3R5UE/u0QCOVTHJ+e8w7YZ75LI9gKXRTcF+dnDoS8DNW9I9kkYxw8pRs8l/+CmM3
7Kifpm/xxP+P1QXe4CAlhz0n+kvjQ3Zm1SW19bYTid9MBsj52WkVkZ/ZOEhfq9GW
MoYF/9lQx2EiJoyRaYrPSaeMc5cQ0vB6tNSZSwygRI82TMTblT9D8DemjdtevBIU
5tj6vw5asncVhyQG0PB9FpUajY+ZzBS2D5/PhukBK8RTZO5bQn3hPdd9G0E2FEQ2
bnnS7PdC/ktlB/BIjE8rPeNMUVFKTVPwC/zy4rbA51jEz8uMIZ5ee6HuYghrD0s+
cziKjrudXSGwB6NnFIyakLpWJsL0Ja5IJVfYUs28DmqVGiyCJJsoLji73UQy1f9d
IFJMd1YYksJlkohL4HhbZgL0FklRsbeC/HLgdZCZhlEgO15y7nWK1Eg/EjNNw5Rd
fBUGnMK2QwycElsG8R/Icx4/NxOs59rBLvSdG8sdQosxN4tfO138Nt/8TJKnPsr0
WH6gVlvfhukQNMFjiDVmYB9svU9N304JmvyeZ5HzlOyjNqoLwgUteDxJbbYhR6Cw
RT9f6K8mjRqWrMNPBzqaTkbX+1aHfDzkc+lmBWEQA1euj03sVwZsm3y8USIggvE7
5x/nIWZlvtNysHYumpO+D8lzSGUELALkPoRB39xWCG92gzsOa0EPk6HZlj4rJ20P
m5UD0UR4WymdE1sXoi+vamAs90SzyJzphxayptqrSJDObf5rP8rGzlzFHThvnpPO
WMXEHm8e2AeZ3pmNK6O/ZRl/tQWmnlHTW/2gY97Wgl/S/iszO/wT8fkzncEAmtoj
OFavpquRq6ZDbGT8YyPyVRXiEt9N/JPmMCPYSGBcylyVuGstAy9rvQqwN9OLAYCC
O46nBW29HfuyoPx1RvyL2tM95l8MJVFqrV2SYr5k2H+ostnf21KjbCxxXJLTMvZr
lo+rl1jHebZ2UhCpI3BtvM0X92jv3zELAAsp4M4GRsdFGPkU6GsLl8TzFTvnFl+Y
gVPwQi1MTmb5Zpi5lmFPsTKTsW955u4Vb+2LzlkWfrKlgx4YB/CtEgCAMeIcietV
AYuKZ6dEVyRnF3TAXZoIJQs1VBxgNRe3E7g8VJBnY7kLYcrPWUBPxRSN5e/vWMVW
WUCUFWAtIthYEQzgF5qJkOEQQ3Ybpf44b8+HloN1uTJgaJK+kucaThvWRPmW2O8s
3GMH5JKFdKnqQ2hOVjZtSxWZty+8LdLy7QDA3Ziwm6qH6aVTwDbjMc1cmD0Hg46R
iFIqxYXEqC/twYT5ByHwcI+mCqIWAKFF8X2SsDPnByMUi4IL3eC0G+Fwsk4J0ch1
FG34pn/R0TQYqIVa0TSU3dS6895Ldsjn9BYMJ/8bEZLpRbAvaEWbsEK0ZJPwHJJ8
kHW50OGc0yhoLW/eQMNi4s+USKf8F7KpMHWIDlj5znqUs/UOvGL+XQ1zTL+wyXxc
VIT+Rsb8Q6MLUxxnHBJkNcCuwcy6MBPhg2OoHopp3OnlHeh3g9O7awn7Kx+6OjDJ
AQeVMFEzfOsbzQMcuOlBUV8yMuusXKTemdDvdrc14oKdd+04uoxAuKFb+f7Kv8pR
7AzRY/52JpNB1WRMhUY1XAdfhZcAyMgiLj3py8rvrOfk5t4nbDx2X2ofcPXBI7I0
MZecv2kYyZSbh+770u/INOhnx4b6Cqf46Bas0BEGg71Xzy/Jo7TMavgZ94X9cj8b
yOTSREH32fWMIhjPNc0wDjBofUStlqsrdN8obLPn9UVEaMk9TCM7lGmHjq9FVpOx
TlC2OMjb6bJqYn+1/HtBObJ4F3R2EJDMG/11r8VhRpr3dGE458FvfWkF88vZS4ZE
cv6X/onhb0lJaXcvtdgGPPW7pVX7ahi17aasAr5ete/U4pUwfAs0sYYELjzpEUp0
nNyGNNrZlZ5iGd1NZmnKLy6iwtwTG6VEmbqUWBJX+rRmWY/Igh/H/u//WqC2JAIP
VMVh7C2nEeXXb5pcbLkAymjti8Zm8W3M9EtI+RlFW6j8s/4F16BE8jsO+VVFPV4A
MXD/tsNkzLOw2PZwrnft3TRwKETBa01FWEJLjRLGAIjp7QScBcjoMjN14aCOp3r/
dv2zvSixP8ejPpY8cWz42/YXTq9+XNUGZm8//jT3xbujyHKDAlOm5aejqn0tnvLW
O1lVL9eMRHZISrsNfPnx9UVlPc9iHRhIW0n9DSwR3X9DslCoKdds+34/Rwhpaai9
TBjxem0cHQEWjIH/BwiBVi9bosKiUs10hZ1JkomXf4UQoh9j2hv+/top1jvHewoF
71I7Ps8sOznhTHIIha/VLnatD3HyA1QYxRo0E5DAp5wRx6rJYBTmZHNnxPmjUkxl
FOVzvA0RoUTpRdTt8Eo10TKpVO3OqRcpAMfCYKqJh6xzqz9Z20TT79dmLGjxqdbF
9xXNsXGHT8JiqpXkpeBcUUkPv3i47Y6EAaGGZpNJoXWsqumPy9C46xvn5g64M76s
VC2fUWCL7vuInvRfzSTjWWweIz3Dg9dfTLcgKR3gl/m4W8G3xCZsntlK76KPpovk
buPYQOY62fK6rgA9smhJkLiaBZqDbsqFDrZuuYVvy4S8UW7xhpjDcDYkXeX53I1V
TtfnY4pIsiwwMrgNPsZ6LT29uhMc7L+Ihb9UZqVFGZwM8SB/QLdaJFfacjhYoDPQ
5l57dGVVJVbLh9T3E4oquy08RS6glZkAJrZJBMu7eg79sfRlKvkKvnE1SAk8p1gO
dNv0pUG2c9Xm3PsfbvZIZubxqRSbOhQRzJEg5M8Kx8cryxL7hDh8x0ER+0VBOGqS
GFUVvgxGoyknzj7vaD8HrQlqZL+ZKIl2od5ACeqj9eZYLP/QyQi0zClrIWylHU8L
uma/1AQr6fLtQwKzBj0P8V/CK2G/w81iGXwLaA3Tf++FB5sTSlS+9unV724VTWZN
YvVSDURoVwQmKNYliVqcvHgVnQVFkd/IbVMvfQ0Jszp1MBAdFIbTAGqdqXEHPCKa
F/PjrZQsmIiBZsGuZk7MeLRyLHpjkNW3Bu/u/OfnldddUw4fM0KTw4251a1PsdFj
cWAMvJeTn/jxqKBpUJUR8JQQUCmZduAMOBQa4nVeiOdW3kmgG54NnUXJ6euk4Fm+
n2dp/mt8XbZ5i2+zWtI8COP1SbQnswDHIoq2hCgQjuGDUbZZ1IOUMhEotBuogyYL
p/yxYHgFUiEZPBQM6bVusxNrYPaFz9GovsbH4TboO9MDScNtXdI7oXIfYyARLj7X
4kpL+5MaqSPjPeM5LLmaf15IGm+Fpam+bf1bNdmstgN64zk7bBNdVuS2fknU8Zdv
mMYUWUiQNK+CJG8C8d6jIrDoITsf7Kpglrvh9RFwxzW//GE/NjEOudvemcM/NxBJ
yA3z7KnHp3PMd4IWeqfvwk42tjq6yIOLOex8x1MSt3/oVvj+jICaU9nsz4okDTwH
1cT7baSkwaUFyFuGsv9QpAUNjYU67zREU7jm+7/f6C9rOe82kU9uBK+wYKJDtTCU
9Yw/XbARwmC1UiQ/E2GQVhDjGM0gdWmojwBSqtfhh8KdxFd9ZoazZwtzwWRcJYtx
kLlcjplAdSWg40ucfuG0c3+cRfxFeVCWQ3ABqmKptVHf/2ATETLPO8FCbXnvOmUz
oygIm54M19Iiphn9Jpspa3KAibA71whGO1byuYxqhq6qf629arTvKVzVCRFx6nJZ
qdF8sO/R30ov8F1XYn7fnCMIY/vtd8/AHugpyJNNal3kzshv++wex3skrp4cE1E1
51ybtWaDdABWMFQjxpYWT/pRwzQ3aSYZqBPS4WHLtUusXJJEz4NKahWFy+Sy7Iik
vmHw8x38PQkAGqIIbxKI9dZXxYUnxuQgUVaI4DELn/h15ke9zYvoOJT728wPU61u
Hy97UB2SB7KpORhp0e5gciGWvXaH+Np8hbt1AQzLSzO4jIgGUufWJFvD+GgxLJp+
jBrK+XFzWwC7KZCCPAgxR+VchJrVV37y9QlUYa6GxT7bLRVt+P4anjp4jApyL4fU
Qp9V/CCkM1aux3hqTOsLv9DrYg3C/vZSaWQslX98AAwPWY0hUtr57VtP5wE6RSTF
OeWyemhfaSdJP99XGsHJYq/lRnlg55A31Z4wkvnlN1yiRVgByW6vkUQWOPZHnt3Y
SXLmfNxfPPKHYI+5jPFt7YkVXSy26JzwZeFWARX7uJMkT9so/WOSUvAKjLrx+Uuo
0p67ScaBrOd5POjZT+F4C9mjXa1dw/GZCQDHjS1BhbGIVFYxzu8PADuMK39qtfZO
+DttR8v4Zo/SW1GE5sIp6YpyIZdHlC8SPxqg86o1B671EdRFRRCYlbWg2BcwvrYH
QqaRIGTYI+QOWnjilAr/aow3TIvVfWoU/swQdWfl9poxM/OP6hNOPdc1UnaDXKRO
0Yg+Wya8KzwJrbGC+18kXEpyj7ekOZigNOLPDhtCpsCvdRbRFopC4aFYYjEH/gKY
jp8hk6FAVQkpo34N7xAFeqTrwwaZyTZebywvCKvbohMdWdGXra4wcqh8A/Q5bAd+
xMNXEuZ4fPmEjYMLPQQtkZk0oVszuF4sm81qRKsfgSPXfDu1XBA9VL2KSDoesT/H
sppoaId49yJN/RiW6R6v1S8EsVxbHIRUmnMO4NmoRVN9fpN39cDH9nHxwzlICLig
Oe4ot/Z4gmWK40L4pHO5OMgCx5jnR9w/r0c81/2s3RZ5DoIRviSY97Fyx6uWTGy8
FGW4pUjKfwLdNGXkYJ52RLFQdGBOSg3owX0zdAk7NDPRwNPp1Bm73JaCcCvY+sqw
mYfw9EONbccv1MaSUEwSrpA9nQiEhVZhtlU7W+lEmO8dTZ6jrc1M+d/alSGDLydN
dl/FBDURSQxp0M7GfF91GyAblRoiatUG+Bq2e8fbxVSO25A35VdoYprmR9ovkSzN
tWn+fc1m4cxwCAyAMP1+edG1XXO+PymvfL/b1BGigrEttelsddAnqErKjyboFNrB
svv9CrBQYeHF+8Xmod/SEOOMXi4/P//Jj4JkA3pHArYeAJWMBgIXE9dhUD1F3Woe
Svn8GLKf68TTbOnV8+ITnbXoa4ygYjtTFZy85rBJUV4Ha0GgoVMajDsIpPKEFMmR
PCck1dZSrLcJxA7kTa0B8o1RLRfkJ7+0YmvPtuXFVzj7dWtCRcDSZhLvqBq11UXT
mYMG1WLuut1/GOV5j/Rc5ge4bhOXBzGvM5TJh1oMkoVx9yz5Na4wKF7u0CZzILQW
/P6cDLW35r9AHHAvej02rWrMVVa/F90bIauoaUMTi49GulLM2R9p2bmzDhH+YbXX
3RdzxMDiONUhQZULmMpIgWBefi0ok44PJisySPHjkNKKSIxjaiQtQjPIQ+u5+ZLY
yhpeLp6zbMug5qRi+hJOEou75UejNNn+pvyBYOyBtYoJcJWoF++SPVze3nYdauNe
/Gn94k/+51Tzxoag7YGvu8CnAlzOrsyo9TmSBGUuQT60a966IogHjdSkYVRVlPbD
pbOzUlquFstFDdhakUXoY0APpvDcWj1athKaygS7ru2ftfhAJdjBkTUuU7vfW0BX
CE95HioLkc74hJ47Z8QeR2ocJTlNcmTPc65BtdpQaoiXXKS0jRIfFmVW7fydoUUg
OeVjhPG989lIGCL7L5+0jQgXLYYwIJAEOG++SHNAu8g0OezHndc8sSEu3uIfM6MC
2yVvVqVBdqmo6h030Q1CT7zRochdVxdrs5FW8122eIgfCnrgd0+jsFnYS0pmg/i8
W1c5G0MLcMI447YBWoWZzlEYkgnEu7NfPRJ4tNqTxKzFEyXyiUJAkfqmOOM/T/YD
RQSFtLvgoPmbVUVdNkfZ/f3SXWw6rH8EC8OZsyUIblvSllqukeJ0xiI6K4PFKRjr
/ArA7Dq1SzLg6d/lE6KezS7IiTBFE4kecrKzHeMpGb6q3JSaH4NkcXl2FNVVbZKt
Ue9iB5kHfLlXObKGcjE5LCcqtaXOc9LtYHkamXtPWNyrQYLy8yh9WjAxxc6s7kQ3
cZFT+bpe+a6Vc3rwMv/cU8lm1LcT34AAQzPgoGJNudv3Df0sB7XYc4hoCYaJjl50
8ZoIph+H6AEwHJmHmceRceslBrspQEXkD4PkKak6MYbRJPR0UBlkIBmX8tggTHVa
/eSWnD2nrqLu4k59ZnRUOup9iwT+lnznPCFHwwoAGrBKaDticdxkYs1EehMOD6q+
OAn7vfdUuhwvnbiAR3GOYz/0HORb8gtiKfLUQaFJaOktaYqtjCFZEoeDtiTvUuF3
Y/mRTd3tbDJ77jjzXU7jy9b5ufY3MLyu8iPHboJS36YAnhpMs2lWWFB/3P/oWkFd
dOibRzCmic+MQOtLcDQ5EWRlWDqS6x9byeG5opnqKedRAJAsBbKVGSpgbaB//aEa
3KYZw4omHHp+Vm5sFbPS78KGCqE41SANPRR8iQIjy/jEerhvDZMlCQdFEy0M3T5J
lDRGcigc1creIPD+RsCPvo/kKATF2yQs4pbRSCCl+f/ZBl488fuBYQn2q3seb7m+
tSDLpuRkORaCv76gQuXHuCMb/TQ6FiMmVRsYpkHlBGgE4uZa87yRCbcYY6vLeNft
LtD1yCnWZsTalx/lrhGV6ckbBxjLL50MiPIqoWimQnW0iXZnWjn3zHZrjyXoGeDq
P/8wNAr6PZM7RuRUYBSbLAR3VMHuyYgogA3rZ3TjHKkNp9Tf9XrmJiUPn+lbHXFF
MfBASfU0QaNBBcoNWWjl/64c5odoWLw8ItWz5MNb3Hug43srhl5poWJs01+EDxP8
0s1zWsQOi7MHTLkZ0EhYn/CbLNMdQAMyqztCCRB8CAB0vFmTd2DEKOGkevScCY2o
rMXnrmVlXh5uQL+WQ2Uc4nJqdtxWqHkR5aHJz259obVkOm2r2N607w1V8yPtWDz/
sNXXRs9wDVp6aduJqah9j/i14kEINx7dHGj6J+zmyv6BfMdwB/pIIIxLzRwVcf7a
ZXEsLOoDtGBGNd/LG1X4yaVt3jeqzawqAuEoWeqBoDdmchZhYeud9NSCQYo6IeUk
Q2PJuYX/6BRvmObyOZVur5wvbX42S1kUkVEJ+ZnDvyobRR10aFRfGj/bXHBQ28+4
hM8ErTiONQaXVYZcKrx2pBSfEirDDV1q5XFM6J2e+y7c7cWAu3YmLqLNHu5iyb2t
DNegtZhMJwjGyEO98FW9zeviTIPIQ6lbeidhN3nH4lhv6jw1LZDqu7Uh+yeDL2v8
u1tQHpofdaBiLgi82NGBKg7BXjxdzAbdF8tL3yc/2j7gHaYQEocdM03DcO4GQsV3
6u6RT+bJZCejfP4RNfCgAtOOHrPEbuZBZe9fg9bZ1pU6T4opH0g0NPxgKZjagAxJ
o31dL8GEFzZsDeKjlgOwUD3pKPEpy+BGpH139s3/REoAm8+Z/3e15kziAWGrAXZd
RYxwrx3vwltvD81+hVYSw7aeGDIwP6f8CHPIGKPQZcOXZZNkfDJ/rDvuTzogiYe3
g2tvZXkJZpQ1TOB2YqQsbeqH0md/4BbxoyHCMaz7hQ5nj3jIZ6dmJOltPER7YTLb
OyqBTydxe058gbCISWCYo+ZHxHp5Y8yFCY/XEyQTlFjPhSxvgp+WjHccrDLvIBeT
agypo4VLDbJIoGnNpTv1jls/u+ZjFnGAbeXkc0gKacNmYY2MMWf0ylRh0obQkNud
npNFw+wu4vl8Xc1QiU1U0e3K4/g3mIN+IS0iRvdB7OlcA46Y9gch+/gLLd1ywigK
QvMaTwdbBv5f+Y+cdBFIykNbUg15auF/W5o+Y/OpNLQ2y3n4gCZn1OZeqMCPVA8m
Nvexd3FIe3R/OFpj+v4J6+srwHrX/cQf3krMIzZTNkpuCinLMSXOnfaDtQX/+iqK
ltqRqw/4Ii515WFXVTGTziLzrvdfiEsc0uh/T/4Q9mW2E4J6yx9N/sdMd5tPok6X
XYHukWaScbT+hYqNIyDIW4/nXbyypgu9HKzCPCAS8BUP0SNPzM5z872AYgbMyGyt
ZhC/Pl+6al3uux/1rSCfkLfKNFsO0jW8NcGm3RgBtGLEHPpZIv73P7/wNkw1hdbs
yR+v0nSA2PkuY+13MnZSx/8VEcRm1AbSe+7JZ6bma9gHMf0Yh4Q1CLs+CmAtgOrc
9OzIjwZNNXd9ysW+tF0gUg9LGSheSST9JnVLWpn6ff7BQ1eo+Ux2nzsZZiiMmXGS
fObKcQ7muMNu7LoFINVvF2fByX2bo7TtHCwSEs/RM5BYb9PEXBFwfaj2xOK+WyUU
RmSxxbZWQKosnOs9nxNQjrMHbOliPIHER7IyfZsiJmPLajdKFCx7kCSqyXsuOcxJ
TMdnHToVpQyadlWnLKveO/QtTRhxNBrgwUYJ+5/3NgqN1D7fBqWg405Nbq5t3j1y
5drSSoitJxQiSKFlj6e7EWSSnbGhaxR9obew7Hp1/SzwsHPphv/1gSs9x3yn+KfG
G6hhUtSfcXOOnbDJ/qKrjV+awZG/FM1VgthQgrGtJd87yVng4l74IPVa8G2FmAnn
G63F4C9l9cpVXJ/fgXl43TtYKnOp4M6o7NfRHhoa3yvb2snvC5sW6eMBenvNUSk5
PR/kS57kUNPu7SdBe/pnwOac+xqx149pDJ2kHc3ipydG/LTEpzYmQu4euZQ2yQbC
ASQG4juU1TqwyvSbtoC7pQjPjbqeTqLZhSSHNrjucXlMAKhi7cJh3pJTTsQo/exI
qEb+a/Yy9XzWm3a76cx9jyPylulF8mr2AIvb+vMHvV+LiCc2nco6x0zZr8DxnCAC
/FAJ1Amv+tcGqYJbW4rbbcRK8QIrHQ3HFobvJg8QkqGWP4nlnLVA+SIbcBchxI/w
GXeukTQIwL87C/jk1dLMr9KI0bV4jHwyrO+OHxj90f2vIO7ckvTaSwg7t+sg3qt5
gAuZJxJ5Jr0XtmuhKdmTBfCjmEwQ96QX9ncH1lNQyL8LpQ0n58EI0575VX6fzBXA
I65qo7oasPdLUEfcxHn5MEb9Hje/977AURwBjZaHxUK41tytQ8+t2qG2ziAqvMoD
sbY00QZOCSaWDJ6jX9X3SpiFW24GszSjRfbVQ7g7qbWcEPJMd+s1dJljRyxSonKS
LP+TaaJOWL6YKFXJ2u78356DMo/K/Qkuicj5/hA7XV+sbUlUQG/EsC5AoDuB116B
/SUx+4fFZh/qTr/GUDG6S9h6A9uw/FQ49wvbAdeyjno+SO4I7ZRsJRO0xsWOHDt9
W+D5FpJiljfilm6wsU9qXPRAOh++KgSSo/v4BzBDZR/IoSaEkI+Eo7umjo2XI2mj
caYfprJX6SsXPBBA0z3gQymASUy2SvKEAkpGvXcFeKOCb7bh8kCiB1kHgrBbiZ/A
ZVBwEum++pvd6xQWnYjjOjfkoDDxqWLRmxarZcKAfF+uO94PzOkS7jebDiAFdOQ9
eQ6YH0c4uqLPHSj0rihWsglBrWnMiz9dFsBxZkTLNJ5tnHOF6eY3z3bFOGdXxQyC
inQDcvtz/txDxDTcj7up8FSWMOCJ7O+WvPe1J58tNIBItWn5h2j99VDABQPLFO+M
HxubhKIVgkcVKMp3zGGY0LOOS/f6W+/y7J/SwZMnqZvW+e8BN+fwcjEaq9A5NIFA
4aBCTJFXq/89vYF3wyYgzNSqDqLHm7fvcQ3Pd8pR7yc5718B6U0Urf+IIFnHIW8l
w35s9XfaE5LwKW4cFrQGgWSK+7e/jUtD62CcOwTRh6df0Env8z51NBuuSJ4soS0V
wQu3EYQcjD4k0p+/YeYKTGIj9IcL+clnE875rNL8JMVcRKxrVYxTZGdi3MlEgEoh
kEB72UPO+6MkctsVk308sn0tk4NMXLZ9vQNOerqSlTiuCh+6q/gI3YCSYPIOnxDX
5mjNe9v8MvHv3Pb9THwi9fEdpArr6TJyXsUfVNAkOv+UpCrE3pBklJkmkcbrMm6q
LBlRqsQsHbIVo1p7QyjqYdFzf5RKSpjxUkgeq75qs+ITaPcAmyOl8cBkMwFq+v4E
YFIXgBeYa/dE1jjrtDMlUtntozWG3Y2G1Kx8rZt0sjEVLwojGN1a+o8BF+MRpz9I
e9781Ppsd0IIMpagz5MUck9BWqHFzR4zuNe8gcqfsNVodXOtLqtEm6GfLNhmW3vM
eJ6EKFHnOrlhNY8h2bjst+18POperzWY5US7j39iX4rwnNZZ5odYEKNNSd2REKVB
R/x3rdMSNz83kWmFKhNuMkbtkcSclgukmgSdEK2/kqjxGsmwaNfvJOJcE2myQxRA
QL0cpzF//mftre0Y+DnpgomkMAP0e4PNcKhI1BqdcC4QWXpDhrCgwKcFG7gNEpxm
LJai8BN6m39Ol74QYKrNgL1v09wEa336qs+Q3RmU8f8UzziwyFsrtISkxvfLZDhr
Mpwroa42ajNSutz4O0ruIiQUD5DliADtKNYn0w8PXbQC+JfTI5UcdMcMxfJsnEwb
ollUPcSqPl20DagQ73WB5njArwdcx+WfFi339vsTObC3GWFrnmGIjLE1I9W5NqFC
hmh7Bpypg4pVxwXfx+JDKexTvbzhQzKhtokVKrPdr+7tHrAUgUJHm6iV0fIxT9j0
GdITHHfN5i/+/eLXEBEtZPfgHulDyOn1pAaYSUj20BD+za5v0zdCTrqn9Sj30Th0
x/EovwsG+XANoKnCgvEbDQ9JsaDfxTFAOAhmVltUuz1fs5UU9nuALPVJQX3bbqWl
z4vPZCPPKbGCgWZJn+y2/qDvM90P/Wr/plkSXQJGHdC1YzfSzmFl9Vy14hasmq8O
TJYyQTexGNXVhoH75LxTHA5CwJdEZeaC6vRiEbvY7oMd4Xla9MvjO7d3rKEDWqKw
lZRwwd5IDUbrwHNgn8gChKJgYmyZBKjB5VBDbc4Bu+XY7bKOIBipSKZ3Pab8jWHC
0IuwU32mEMzVCk9LgbDpKM7GMQ89MQBFE/NNU8ilBb7pjR05cA+XcZ+vYsh1uUl6
zhjq13Vw+581Fv8Z/hbf+Av9/LP/hEozcIj8vOTyTmcvgJVJk5sig5M4soeBywjg
AJAAlkz2myYqGl3y7Yn67LT8GO0GYYuqq1QFbDH5htM7rwlRQ2+KpIGVsqQc67J8
/nqjpe2NqY1u+95mm/7+EEbPM81vgGaAXAeO801V1poeNdcK3YMvnPhxob+MwNsI
jFp4mYA4lHbN88SH/rthy+ZUvbbpWGr1EhcEryI5NF2FUaLZLtyC8trUGm18wLT/
RWjw/IxhB2CENCEStnFnJ0HclKK+xNtWbxpQsRxdVu7jOMwF4eaTQrvQbiQLCMPA
/rAcQRZFvMdi4WtbUAWD2JmxgYeRjnlCwUjMeJjNllf+fKoyXuFHqGHuw35qoChs
1SzZY+qtE5F2UEgaE3T4Mk7Yaeyni74kaZcuIc68VmT5tG8FVh0sd86xURwGLJe8
0woqShEksng013IsdhpIwthqyczRcGCcsKQehVmi87/wcc7sIkh/bic7UORl4Oa+
B98n+/a/UwtI2sKs6qMIdgOIGEaSFKTNrRoxBk1yUWAbKjcnqneIDfjbabN++Qh3
iYvCojcOCdwJEqUerP4BBLjr+dyfXs+ksoyL7tPifG/B10wH5AUeGF+WOygq1pSk
09bqmhOjMtz7VMe0BD+RhJhj/kbe1m5e9Ry2IRwjgj4Oh0em4pXZTNqtxp3tnU4z
gaTL0etZlHCATXR3ZG8rEAsCKMZsUKH+Y5ClAFFxgqtZfvmZ85dWw5Xrjxo0/4O6
By31MHGx6fn//v2R9cKIAzk7HvPI+W0XwwR+qVA8uTEvRswV1gDhtCYHY+tUPK7O
qyDOOBwb0/3nhlMkkizIcXIhe1GQA2+BycOkQ4zl5mUhckw2T1gTdedl9W/Mue2I
gbWJsyNDQbO64lZ8I+bciV1bllFjCO4kHtxVRnBRFbz7nOXZxiZdPwbCudQqg+EF
5NbweKR9e9gVHmF6I4eIlK0xOjiOKY+QAHdqC6gXb6l69yLt44LCBVivMEzPAZDd
xHGTkmEK/8mwVjhv3qzSEbH7xt1/9dVEqk8vwE/qFN9VEeqCbHhU84EeK9g/8ff1
mOmSsIO8oked3Qt9DSL+KZFanLj94hUcVPDTTnA1LM2oplhXFeLgrqZH1mIN7oo7
r0FwagbP7UJL/UinmeCvgOXZk5LHOldOs1lc+ouCBuagy0JkTH3cTxMFommsLpEH
pbBjTo1R4BTwqSpkQtkNGkkSC5RNCdbwmp16N/75sAdoHP+xlA2KbRfStS8C+fHa
92RWNY8dRakw5NCccpJTv6az15h5rLbtuN8klzbjc/OD7cb7dHqC30IA+0dbKSm/
74PW9V6ubPsw0jSKDW75mmL8iQzRrrus4ur4/OqwbhMkYTzdnJqSGx5BGCrYnCVd
xx96RNDsE80AzZAW+NcuUUDJ6xdgTARNYWBR1g/lrCV9Y3lknjoZTOt2dcRYjuY0
suWtdPHaWMNDWe49R1EBIbzF/tehxTTUiyzlhWAOy338yjD+GEwO1sCQlN5WqCS9
0p924za3aw7cfOKsFAnRSsbvIlwA91MtSUrRW/evT2IVk+mUfBzR66g5lcN7IJcY
0FBp+RgUX/Z57ytTzVghV4Tie5Vg4RckCz+0VLqKC/cT02j2d6CuiG5QNmYVynsV
oupdlaXT0x6l2kErY3VsAknSc2p8kLYp4jEblpv/DmWEbKnN4xy51Y6BDPJH1zTQ
CCh1NyYKNk7OOakaMTuNdHrUoQ02H+ZWRJzfT7QwVQ8cHJOI2VMYJbl9cjQI0aUR
LK7hCDLPAequM6aiY3e9bAYAEdOGRGK2EEEW7inRKbO+CBhJZMcKNJs0TwzbddVf
tHqMuPZcwmWqxLviZaAc5Z82F09jXpPLKh5iUhvJ2tf3OLuMwOkbxor5nZMiR+cT
WcOl4m7uzj9e7s+2J0GdcZCR+XmtVAETDgjPBi5EKMurlvcvYwIuAks73c8I52r7
vIaZPwcQqQzgI3eu4NVx6ozf7Smu3Q+LMgaPAwhvkVpLD6DKyMyAtt0BOMt9n0wC
DRXfY0dQqrcNrOlNlhOjMzSzi/QRsirmWvyYi6IYqWb5ss4S532+86eZ6A6+cpUI
9eQZIYci8KwOo0BJ4f/LT6nxYUQf3HnZLUp9h6ob2cTBbr5yVYS3wS9hrcv112KY
KkNhoc37tYqtj3bEGu6WFzupd9FLBtOWj7xUcZO+BRbut/RL8jjJULJdzgUOgibL
nWvfkAN+3wDOV7lW3/aqMTz3pkWA2LONONfo2ed7Drf6b2qWCFJqH6tAz0lbhU6x
I0fuRnVxaYOqO0pKL3g7iq/V4R/lF2SuidTPlyPfIu9wYUWkBWxb2zJ2sGuyGJdu
XuzawIKz3XJ+8o89sZYXvkqBTYCZmV2PEeALHRoz8t/g8DF9AKoUEViDp2MNeXRI
8erVxN7zL2Nwx2bx85GQLlc1WWqhwY3SG9NqdMmTxlc/YsNBYpGITvXytkvwzmrO
3TKu2Zveyip4miH3490gzXuXccv7jege9lv0NXn6itxCihM9iKh7UuUcyemX18uS
8sJW4BpGc/T5DR3c4WGmwVCFE2fLUjdxEoGbtY9QEC8sMg3Tz/rtBstWNOvwS+Jo
A4TzREeai1d8rV/hl2eF4MTYKkgTyNCHtPp2tlrN7ff3x61zTnSPN2DQ3I1otXDF
G1UWWduewhyf/Z79jKvtNyzsEDrFdDbL8D0W4rmEpRlwHM7PFPpK5hEwPtqpNEod
bP8RD9lHVcaYQPgel51VRu/SNxhaAZz30/MEqaE0eLDN5rwC++kKpcmeesmwdNi/
aUzNXZkba1ONLASdfCya4a+Ody4QiMMN3sgKOxSxgihsyYO1h7ZeHYuA22NEWBst
wq7XGDUzHQ3nNvIZGQy4+29TCHCRclWAMPfvjq37pxkGO9K2veo4v05Z8+vfN0fL
6EQko84jZ3+vdP/S3L58H5UX84stTEPJI4DxRDEUkY7aazoxThlVPrdXvVqlsOZw
2I8AnOhun9YPcmbPseNo38E5h1z7qr+wPCgfETv0YffSmyUuSyUQSEIl8/zV5Bn1
IgM5lQsJogpIG4rNEuofBXetm8ohLujteGobqSFNsnBqXZ3AMz0qFFy/0fA1B9qK
3bd6rHvnEXPOadfsJN/1lmju9wcWqT+BLNgsR0fKAx4xRHO7Z+dePkN4Uh8TvEsX
JefwUiBVr65jyocUm25OD48ksuma1x6QJ4iRV7mEosO45T0441hkeTdFZVQL6shk
r7Fjey1lUX9IQCknW9zLq4qppFEg6DcI1Oqkxyh2mH0UqdRxZjpM3LXQI5VNQ+Pq
pUktVHui/RWrA5URJeBKql1cDdBTst1oIsjlbeIB4j7L4JhhiNzoHa3rDDCVe/4s
zZQtuLBPFPZPpFKyoAXwDLAu/1m+Ako9QNNwi5kYMonbxAxtEaZuD2AY5/+LXiYN
CBebDWtawtN9NhGkgoq8oJo8O/aQARmZO0Iol63CAqBpxkn1Sr6wktA0yo0PYcZG
aiAMSwexVnRRVOpeKS4EmbGcFocR/lx/AUKoy6r07WiI3D+6W8HWB30EgMXI+hmq
YYY5eofui8qa+vjk2GT5j8AiqpXgNlXdhGrAbznRT9TLmKtuxGoVv/80R2BIazAN
Ye3t6BQ3yJY5YBITA8bM5ardh7g2wSU723+DH2jDtRtQKZMlCds0HRiMgpvkl+oB
E9SBpwkURB41+Y6tFjXlqQ0hRiHkJUN6RAHv7n1aH15TL3uni0W6+Vmn7a6cdBoo
DLCIM4H7WynrQctdwCHKWIxscypjBJCTiJUK09F/f8Y7ejeizPsbiPAI5dNwbHrO
RVJ+Of6swlfYfaJGbi1lXb8r71b+PNgR/Azt/7RovRGBGENmBB3p+tJZF0yyng1M
pkSMCjQ6oq4YrdOEW3Y0qt50+/iVHxPeedEx1UFcg6LMt4TdXtA6qWdbhr7rARDK
EzYHZLDTX/08Lnyb2B3q6+BU704y0DlZT/N8/Q8uSRPtxwDFzrcnjdfWpA6BAmAd
yJU8kHN8E2RKGgQsjMYjaIEdRDdTO1Au4eerm7FeGRvvD6hXfxDrQzoaMNbJzjxh
udjjfBOmjnwXJ6ItwZHBn6kywgGBrzBcnB3M+aSc+XSAKTXTvAjSt8CWmKpzpw4X
qkkvFmzOgEtKIMKsW8VLsr4XJd36qTz/1vCAWoIC+NiN+TMexo0b1Nz9CuwM+HtO
i+Sm+ik5c7EUmg0X2edQINMZjnCCtDRpF/cEEaTUI/Lgnkw1uXjCEB+TLxwzRNiU
sLV8dTOEWssEtm3HcubZU1MIDvf0N78fDBAds6f8Bmajly7E1bEzSG1ZW1KVJNju
Vlsu+5qabcJ7+Ld1Hc++zCPPtWJzR4gGCx2QOPl1U0NA0M7d/3KcmwkOWUkUS/BU
sul2/E1jt4YaMxkKDCjszp5POgUJg3k4sl08WgjQvb626LvhlqUab5t0Q0Ok55PG
wI0VzOlCDMk9m7KwwC8JxQV4H7+jSMGsWPgCmGn6fqd587Hc8L6dcmax55se7zfQ
n9G3oVpgvC+pXUAxPRRQifjAcE0jmlA382K+Lh4tJLP+p6o/XRSQ68pZKkI4REZc
FbneveGeMG11D84wRrivwxAzEqRwmekIEx/nyR78CD9776xA1vdqZThgmOjX5i1B
+gCKBJZKcmWJbQk1SWeWcf+MhWuhAUzxiMceJZjBZnqwAncX5YyIJrTirHWxZpf3
Xd2fxAzvDig3E2LIf9UaJZs5eBrlvmPHgzNah3OmvNwPGKxw61cf5ZMs3ANwzeFf
SPFItrOl3N0sJcnX4PezZ3NmY7eEy/wUGt6hCwiMHLurraYy4SY7pNu/62d/EFE/
Wlr6WVsJx/Tnb3NdlwLzvsIUCV5/5B2Y//PmgiNVAgp214dR0RzP9HT5KBEP+2dG
VO+a3hXbYgUU5hBvqEKzs3rTHIp4qsnbYKlytG1Yb6LSibL0MErGRqRSe6hjwHl+
9s+J6OVZEBkJYimXRY271MYJonD4MS46cKC/a3oX/3Q2iUbPrlLOJJLNgNioDDYW
NopPV9rucwW8+B72vyE0MHldo1McR5gdrw6noT3ywRvqfhZ1VEHootTfTBEY5ccu
B+nYSThW4GtVSektjCWTx5EzI2hbHwYNKGYLRvLynisNTb1DW8M4d6X4YI2yVl/2
fEQPMJ/+pdDn3Mz5FwFJ2lNA2jrafyFAlmLPiavJ5A1JZ7nXb5a4mKs3VzqIG0On
otecnQMRxldqH+6vte7L1QnwGFFG0XrTZgjMAkdqCRVDnSCVTXl/mOQrtPq1xtBh
Mclojg3mFGvhseBlQkHLEKqSAukC4Deu7Ip/TUxP+3fp1tPoh+f9z2ZRCB8zkBX5
9CBL9M7Dme6goQ4LhLe90AMG8PoHjK6vJRHvJv+gWxOfsllN/cRh2KzphWd9NAGr
bzO/497lIzZKUS+YxPjiD2fYbzlKFBb0yMusfEH95OYVd+/ENJ4Sgw0WfhmEv7zs
zPRqHMA3Cexx0qpIZGqHqOrLZ//aPIRoZKSvaZn8ExEA4nFZCLlQF6M7dF2GL8sp
JQtlYG9hkZvFBmxaWlZ1IP8+GL3ds78hVdbKjMzoZlXGX3mcJAEOA4ooRrLMINAm
RRdwBm8lnbROKXROWhD2qvQ7p6UKZHMq4WMlyTqeo7UOLezS46KVD89jV62bEaJ8
XcmBg5y709S4yBXe18Z6GLU9Mv0wgrG7rCAR7I0UYprBgtZUaWPRueypPZrpJ7UE
D5HKkv6EOjd0X2dWQuke+qAWBXSyZ/b568PCdH4P1k143HUIYgLDXOSG9zLlBXrf
p0WHx57pnEifSvMkyYPMooTvrzICEK5pqQHG6kD9TGm4sJkqchghFn7FGqP3IMKE
ThOzBOOY7lWbg/HSNjARfN6aKQjSjab+rLkCGHVy+ON5rEMZRN1Y4cOfFCBDp64C
pIKmwQAtFMmnt2zRDA3JiAtPSVVZQtScG1pwBqMvkiViagQ7lo+Qh0xEHd10seAY
VytQ2Xdnx5QFgyC9z9OUuGId4G+e6gS6BiVff1zX551laGKsmmPUWiAH6eLkSjf/
64djO/TbKdVhi/6bMRecYOvnRhfLg8K45TNPkDPlB2kqKCH97I9Q1Q0Cqv3QdQX1
WoZPeawq8efGTWlHWNbvtZTa9NeVzI5aQ1UIo2iBGp/FVRnWJB+TvKp37DL+qeAo
h8qzGpA0fK4MwV03MjkA9WBXL+5a6mgXGcg8c93Q6HGWl8lCh/pnin4IiApn0lTe
8mLa8eJMtt63mVxjzTMpt72jDZgGFytyijdOAYM/P1bINxOQvhEapr40e/f8krwa
0BDfrXovEEVFq68f9qnPBVsEuzPFyAv94V8TEEs7culLBFLLnuqQjCFson1ILo0d
bwalQR8nJkN8bZV5uyalhEezyGtJ9lqmt9Moy6TmQMUUet/VBY0tYZNs1aI5Yd0j
PXDY68RM9g4d1i1fNPDUsO+vplh99/nlr19lUnS1vyV9Ycb5SJv06oUMUfAXbs1z
YbuvTdM72x3C43rdO1ph7QF44ZPUx6Okludnwb+NyIo11uqua5EhASy5ldRuUMNw
NKNWeGL7vUowIK2q1QiFiEcUeQroqMSwVg/tVN2/Yr3cNO+Yo+HyKTJos6TVhplH
atLkz4e364SAQT3j81rccbUBzRlwzHFlPcJrez3okDiFsW+A/GwYQ1zXVjL3iB3k
kLY37hLYmx6qUmnPm2BTkRDHyJPMlG1wkYLK1mk4fGhM0+PKWWpfosvgQm/aAZGX
Rwdepzwlf3IVNvftfzH1AvMampi40KS+WpgxxaZJgCZGZHEzbbj5NS3La8wKkRz0
myCDd2wwNtnqc321IQ/TDaMUAPClogMMQv/ub7c5k1T0ChbG3mkVdgKNxRBihQnM
A5Q0X4J3j9yUkHm+x7RW8m9KtTMw2ESILqKPwkYPIVYCJ98OfS9tW7wFEXcr33Nr
WaWjDp/JR+gArwLvBjsUFXwEN50dpvA1+b7ANud9vxeOWAQqx2C+hIQ3QvwR0o0G
4SAJ/rop34Hkq/2RnJQ3AKYxZBwNMETR/g3byrVO5kPYMo8k72BSmBYdLCe6Uqd1
FNAz6VX2UAy8ncn221OmlM6cQ+xCegG4WMB5CaU0mP/rcCQEr0LU9Zz0GwVH3Ynr
71FlDaNFEQbPGyXa077+rB8ZPMhz5H7ISPlK4Pz1cCwaLrvtbVtq4wZHVjhQlm1t
13shjN8BL4mGk1c8Xjg0APr2fr3P7HrNPPjcmdhOE3KEvyZDcsOmFL4RWUdmI5cI
DGH0ITn51CWhKijm9Y64/Q5qZdrJoJKy1ZKMf7DhMKMo2lHntDefPNSFZsvtRTjW
pEOuHNw2IhddJBF7226yUlKip4YGmw7+aL+yABsLAUtEXToxoU+4gyhNX0RZrPst
NR7AGea2HqFCZQTuliM5MnS72z+ngJ1HR1n+3iCC7Z3zSPiIBsiXfTJTDKw2Rim5
sLfwBryyOBFXY/2OtkMHMr2+8eYW4IlSuluCryDy55rGG9HSOe91llSdL5YxX4Oa
xBdrB42D9xfmp9Dz1JZY19402pod7+DbnXp7V6zFpe75CH3Hacbv0gucZTP981VQ
jGUhurpnzsc89PMaitPY5/9VUB2sImhd4VXRkPd47qQa+0nR3WX4wLRztI60OgWH
CzHWWNxQHBoBdze52crHKiL/mH9P9SoWgWHWBBcqU7CCSYfxJ76K7wLBcMhGjjDP
1QjhUuYwd1FIg5D3p3BEgM0eLdhHRNk0l4d3I7li1ZVEiDumnNt77w3EGeiEPjGT
DyMau8c2eBFgkFCEtgohMtfuMA6VQ3mp1BmOPQxiFSeFTUJ377Bqi72xFUnoGp5S
HJ6HocwZIUtgyIU7GmkjnE0NMDTELfXlQqvMYA/p1eeX57SwQqcHV1knsbZ80VMt
W44CbdMKIlcek3twolMt0BDAX5r0m9nRBN+8PemJqcerlE411021QiOKLKYyWhcU
F18jRBpJQ3SuQYs3qS1JfntwjKvfnaELeaSBpoYZ80gSGI8cXHVR3ZVEpIg7QYNB
jd7VlxIoeC8K6QlSCuXRA7VFrHUps8cJrfOlhV1CoDGE8QwZNEiP4ntlzeES73cv
WtohZ/1+YwtsBtfDHJIcLJ2U/mz72vXz82JkhVhkvA5tf9l6AxK93PVKTe0VBmTx
uJcHdgULKmuTs7vEICaV5yXRttS4qcGZG6GmqPTAmOTr/4YE2cRMq4ZmTPZDGPV1
h96esl29KO/1mYpppSA99pOAkmap5JwzqEa82QJeEvBj0dUeQL5iwXZPuAN9WOTP
VCG9sUuvXOE/Ef+ZMBeFBHZRZSBujfFsHgNSnvm/SNbW5D77S6qwobbplzUB56IM
dMOem7xz/9rUNyDz4xC9tCOEmRaTJABPpeSjw9ABCVU1R1EikFTWCszc6BeX8L9z
Ggq4KX6kFUpwksmR99hRXThcCguQw9P9EBEPGp5EPzlB2NNoebxTWay1atBbyW/I
sjVyIu8XdBC2AWa3VxPutNlSricjydJ61mpv59sQVYMinE+nNPTlwimeQOaW2+n/
dJ1bUyd3VyWUtlPtjGjC3BuET7jPJCAxWLchqZWSj3iQVNe5OVQAXgZR95fK7VJ5
j1gBDhb+3uqJn4RDPacwGdjzA3GOULGKhLloUNXuHqbpEGzANe+aQYtq2kXD2NfO
oIQhV+tYqnoDNlF2Z7vQ4egbrz+ykhyhutibYoDHJovKLPCusfIwfFQdMH+x+aJ8
8LGKmtpeOYwcXVzSnkirmeqjw+XXemwpZxVc1sOiLTr5Xrwkf408H+4A2fcCByLY
xsfwnA4oHJlfQ9QCor6cBiykbPgaQ625najEXCVXO4eZB7kJjbpHUNAPZoW7nF06
xXSCx2eKYvhAocY/z+jsD2F2JKFkFblfYBIfELYZO65mU6KFfSMxoLMiYq8mCthU
1ngFVdLYFWGo96gOgzDBlggl/seS5znF/wK7TSVpX3kRFOC6sda2T92dhkflYHM2
uwtg7PeUn6NTtaNtmlnFUJ15eeeLS2UbcRcsAkwW1HbJG8DjtvX3t5sv4Zc2ss8/
D5PFvAlmU9t4hLWkfq1QgoyHA5DXktqcX/QmOcw4NAICWtUhKwlN8kmQv0iF0T2b
W7B2Eduaydi2GBtBDAMPCrwtuI2Hqp68sqxVnpI9+d7b3Pk8oRdMhvERAJVTR7KC
krb5cb4a13MHKGsW76/xIILZiuHDsO+25+mfCyujyLHsS5+5JDrF2LB6AneoA3wH
lS+ZCX/5Iy94HvCiY27Y/gMM1ZrHZl1LquQe11PhnlrGXJJWum2bmTWRaC3iErgw
w6LtVlDbXtgUYCkXPEb/6UKCpX6TfwJjYBj4WJSNO575D2clSRM6VD4rpXplVg5X
Nm6nQ0FUBai42EAZ6QplCDnJ413LTUAzlSNuy9wCUZqs3PMi4rV/p1fEQMgAs/6B
WiUtBEL5KS+TdObaeUBvVuHg0WgkYKzFluMqP2ABHjcfQMiuBPe/PBXA55BwQgSx
STAICzIz7otrtUI84xCaLE06FD49GgMiPbPbFHBfQnfHarHQAzhnHJ5bawCDLf5D
pMuWDtGEBsT3sDKIxyQ8rrKAvfLw7/hfto9ZHUVSBdxMFufcbpXmETys1obOikBe
SA+vCvxnKiSCUKBdTdUoDYbqvUt5fhsH36PjWf4oT8ELJE27a5r4dHi0poCw2npA
Az0OUz9U4KBPbLh1h0O5SzaPy/rGgz1TdCfeJK7k7IUyBNF1vwdjoC9lG3S1qFJo
ZcuxmywxTUvJ4yiSlw9x7lSO0ikI8+Qg6jW7+NX2N4Or4KCTjcGWs+8naL7ZUkHq
IKIIPSAZLpya+3WuzIv08MqzbTIMlNP7GRpk0jpgk8mIrEgzhTFEuLQfFvSOAQ8M
V5DVDmhUgJNKRfYUBMYgHuZmxB+PccKQM4Q3/0y56M21/OEB/oEsoauKcvd6CeAm
Xb98QF/LslCOJ1mVn4XGQ8n5pp+8yyqIAbzcxkUp4eLXPmW2u8kseGVLKW6M+Kb6
KiusDTWYT3bUh4EfoLvcA01sxOedfBgkuvKLiVs88Vu6143LNTYgkQ1iyflYTz9+
gyYdRtQMpuQdTzWR9aXbe4rA+gkZ4JwRT0427a9qwdh7zbMEyverQX6RA7Hurjox
9RfB2c67MD3uGz7oGIQnvXgzKh4cUZKh3COymXeZk8NVFlx0bvv5ulOPBQJyhcUZ
hxFyCTyqUNriS1SUH6XVw8KJnKnbTKpT3WlqVZYxPRDqKNRbW3gT1r9GPUJRdIJ+
Obt82e3cH4vvAaJFV8ZGHZVUe4RRUVIuXrv6KWUGjDb4yGLi6uHqjThMw7D5GNE3
EBZCJHIchLhU9dikP2ILw2P5zZm9ypqYrw/XX1Jf+S6GBOL1F5L7p0Z08hZc54Hq
syUT70M0oUOoO5LeAxQIBkGORwchgToNBQgaTG3+NJckxaC6y1kgZZQ3u1JrZ4zv
KntdQ3GhPY5UeASlS/3M1ngJO8oe7FcZV6XefMSGpT+uZFQfLeynkTyAPaPyS02c
9o6NsIQcHPIzaQ4ZmI5pK6XZYEDuMIE/VGOLtwjRgwJ/91DTjceExP3MYS52ovFq
/evm9ylN7O1Zgx40BRAVAFz5KLTTEOLT3HbC4Vorv1XH6nTQLu6PFIC1LZ8lXOU7
w8dF1d5GqeubY8Sk0pwRofq2B0GAXcBnmOGSTrvSGjaYEXkMzukLiQKWbgpv7DKq
EnOYztCzO+49sTzKkStLw+Px/LbIQ7VHfaB97HCqkiKM8AsFVG2i2eDPgVE8wQfP
zurcDyWPp5KUx1q7U/VUd9Fzibow+9/FmbwzxPW/rm2Y7gyBceMGxTq7I6CqkGXi
MRl8hn8QxGfhTwsvVGOe6ok7umJVyEPy6E5TTH7+yMQTWIiwxSw3CWSpz4Q+Y18U
FycTlgdiTe/t3wkXULhMCc44O0hX+35XoQF+PEwFjPtb7FE3Y/ZEEYuVse3gtwIs
23e7Qd++ca3+UDXhhiOVHKC4d373agIymTt+MVAFHy1SOPU4pUu5EwZ3ON0S6e39
m4bhF2Qmn0172mkqgsUe/7YwnsLhzK6rpQgGaB0HaU15gHkSUXcyd3G9fRG8axtv
+FjHOZivE4RBidKu0PMMPvCunLg1i/bPm8mrkoEEjKBcleNWf3A756cmZ8fF9IPz
M3sWBF+4fvdJJOrCRaBMoNSU3+pqbegiuVCFff08wOKseaMA4nHrQ/fsiPSOvuk/
9t1aKhfOT6WZt84NK17jkQtH5kZ2IQeGXSI5oN+BCKo6CrXA3MjJ3wK2mBUmobfK
JRj1bgLLX1BJbTcnC1f5q4moOCypjtqnTaznVLZ/vOQ1+Npmvecy4voJhsMD4X7l
Sb5SwUgxLwZb+UTOZKFc58cQjeKDR+sK4/oxXyCw834drblQ9tfyw8nPQ0uULm2f
X/yHWDeOkV/nCx1NsMJGW+2zNGb9XFxwR+RGQ+pMldwSyv824e47sKzlQ8+PY4DM
HmV3OdlFY4qZrMm6wRapRAGyK0kUcWhwe7gF1sL8s03r9nF0bI2Io954/Qvf2Bee
QQIMxj5bXh/pRDtMph6ccLDDlptVtaT5jQT5UfG58UJPos6G36YfTfVDEMMWIxOM
cI4s8m1buzznfRaqVpL8Z6AAt2Zs9zx7rpXLHvvblzBgpdjwEZz4HAMuioiag1ZH
pdKIe/amTdg8uVuxRaDrQlhU5G2lMVoJ7V6ELmkIqzlxspHDjaDxU411D9ya4Ujf
FbVma1x5KlZoFdMHswoAJ+fFIy5+Hn/QgU60TFbZr045XVr9jYy8daVGAdIXa3QQ
1Q8Gu05ee0kcR8bn3blnbavdA4Bj67IM/V5BLKQPFB3tWxe8nVSivrSW+QEk2mMc
6KrwwxlKk8zaEJcgrUF26msIadnU2cu1FjTa6xj+8fyhF7fEZ1k/qg9RJLYS6cRM
lH+CYGHaaOMjI3lakYL53CuqXDMvdSYDZ9AcgVD6PYJnpX+tOy9YoC99S1xQcKAv
wmGnqLTjctNAWM5ovOtJLBzo8FtyRNlD4vpmSKwankp9tmAaqPcLDV8IsFszURAU
ZYXGNNHnNH4OnwA6GqACc4u5F48ymDEP4SGym7fYOwTQbt0S35wbOuIqBj3yi110
i8gmpPORzvQAcLxGjiUF25foMR6EyLmG1TMOKhPaXug/hHB0dOAYpCjhONVF+pxx
Y8K31iJcB5H6ahDn3YbfhUTiwOuIAFTJWzxh4DWJPeOReQsh4YgTh3vXURCoLxPW
esvBVy1/rtCtTl5jRvF1vsc+oaepm5Q5cMvatUKqBfE5Syk1wSqbOE/0PEww92Ac
/RMeNDVXRZzES+CstykiKk9OnC9DyCkk6sLOuwsUmolqUOQm6LVkT03HsAlNtgZC
bGZTIQNXdM5izDk2B+yt5uIrWhaQMhSNb3bKrJ8UJ1keka6BNGyRisFvtevQkq7c
SkJeP44RmV+VEkfTxdLayZpGI9c4YuetkP1hPtDvaSArGMbjZgVw/uxvnUfY7k/g
RQs6NraEj7oVsYD5vMrc0TKUid8CFQGAAojndCO4bz4q4ERkbCzaLDf6EYba/nEm
VLOwC3N6JFss/9xIhVSxjn2MSibtpzI1AsS8su9zwbA4dje6sG3QtHB1RImYCWd0
+ktBJ/efycbyMOIdOlsw67hIU8ICTTbZhGsVlYUBjq/M6xPJhBP7vYe+4w0XHTvD
YDu7LV719Y3tx/YLJKBuJYZjO17dzUAA/yE3RE/HHxF8VpVrtVi6Fq9aJapjFpzr
bIOVAQ1dnriesTMEq55vSXHSPK+V9t/rgfC0T4uTbk04kXD97axXUfwV1a6oExWE
pEsiK7JYbnoXag5XyXEMMfV9tXzNwpMj7yn716REpdDIffkSPSFJign6Dk21TGPU
XzxQFQv8Ih2bRe8A4hSIOe5ilNw6/KIPBnk4CuTvGqavUbjzweOOFtGPT2PavSsw
WVeWwk7w6BZuSh3WzGtgtaAAlwVETmdH6xqrJaM8HCfwYtduF0/hOvfyN0tEkwD6
Npnl7JZjE26ghchnNG9e4+FAiQgckOjRbimRtT9kaLtUmUQHYhpAXL5flByqQ2Bg
oZr0LJiqzcxYYuBh/LQmfbCmhCP4tITuz+ukcc/CIgnNuIVIRdaJVWzhL6MlBFEr
6oD8cU+alsMR1upz893c0q+SiwHKJqu9pAMENCIrBtiN5VE0erurE8mEyykMw/0Q
a6dwt6OkewT4uL5wVfVp4B0iFRk2NfUIDG7uihX51V8KtPYpW6KssZkiIkGFij7K
+fnmHd3Y2ZkNSAjkC7jU4jpatLnskFr2DW60sZs/vtOrPL8nux37R9MQT+yGvY9p
7zn0ZbGIalgFOPF9rPUmqOSO8C86G5Q2uG/K7JL6Up6tDwOfdksHUgOdcFfxXlBt
x9fiIPPXOih8DF1WVHx2RdFyaX7odWoNPhQh/Id3BBIt2BIoffq5SY0Sam1QVOY7
GuspFXPfmqkWCH/DgclRaHFXvrlMJIhck/zHH1aUHz2Q8+FQGwJPREcl8t7p/ngn
vDWWw1SX1MfjKifalln2I166rh1inuB1Uj618LAuwUQW7DYzneE3HStkmTZ1eLq4
iQX3fV1p9GOeD+0zgutLzAETVt48jX8W0z4UniyMIxLoqTrJdPFX790Rlr+ed/3w
EZWfI9wh2t+77hD58fi1eWdQwUylNTIkAAPQRMIiCJlq/3RW9TcE97w+j0p7W1Uy
CzsaerK6NSfsP+wv1J2DHpUOAJi7rO/L2QCkPPaPPKHpdFoPxbeOnvk8tI8u2w1T
0K7dOtKKmMDiVQxk62tpfl5JH6V3FJk++6gtFNz+WIY1y19K/CQmPdp2mrGMeDvk
77ZMkzNvkeprd2GzdvyMq8t5MjSqqF7UXS8FvcIKHi5Nfh4lwo74Se67rlKbXDG5
8TaG7ALFiaxud9bLK75Jm6io/A9nSsjQYzJ2KdMzw5IwdlgipcWg0Z7NXiWQ7WHG
d/N0T4L9JX6ibYovotW8kkw0ETuZ+vLbyfu5oo53AjTpNelhmP+ohPAoXQ34FOSL
sbViMsEMlFqdu45H0zE8QqW8X3WSzD8Wupj/I/unfrrSbKtZbJ1nlo4bmy2rpSiS
UvEDeYx6/NSDDw4RK1NT7pBU0h/yuGaz7Ts3DzPUmUh8CBucLo6LQjEbjNw4/K5r
7y4hAqiyiu+Jt9b3LG5ujoYVoibQlVpcj1fLqoGgns1EGyVWpH/17qbVlcduvoFw
AUuxAWso41xcZvxx8+dlLAXSiSQfGavQp8rG/3YtTBDqan6fGseScr4nAKs+gEoL
k+gTNQFuB5XYiYpZM5KKWk5IwVvLCfv2xmPOsrTu/BLDQ9RIFSwMDwwJrdgaOS4k
XvtIej7hvmWa48MfpmI18LWwGV+J7wpkE8ykY6ey/bPttIKlzdZtkp0MM3Wbojtx
Uj6UeBIIlyL0KGCstXxU+fP82EQ6jhUgSP2ok4M17GS4awtp9MjHuD46wZ2wWTx6
DHi/0clbLcHHQVuEoxaMH25kR0F4hcIAHYxtzWZGgUhRHTN+q+V5VlvmO74RJdnb
ljjDkB2J567Yz3W/dpFXuQERqGtqd3kSBCtJVtENW4Wl4oYQasTJMpCYe0/9cPlL
Mun/fjPN36pzpQGteFGemEubBA1n3FbWOSVM3LE0P/728Dg9Um89NjdN3i9t+Td5
y7moL9k0UJPtdh36fAgRwb6UJ89TpQsgWQpfugEhEow55p95qyjuIXpRqaKGqno2
p7bD+JRG4BshIV/tQUtFM6F8CD06MOgRRHrRd7rpTySVrb8bkRL2NJao+WGJTI7H
Fv+7M+5Nxf08qnD9j/ULtUX9I/X5LrUgXNblkO2aqiczUlkLX6Ma63lJ8koRcbiA
+lw4y5PlHVwwtY8tEexOy6BLuiUzm29DrKlVqTPGHD9tlpLWK/02hqTf7cNWayQy
jP50lwN4sSrirgvE2HrWwWpzQYtQYwRMlwqrP7FV1KzF8Wc+2pVU2/5K06q44jvM
sXtfvKLygWgFGEQdOhhq3AU8J8KfF//N6DH0uPM2G3F9mkZzEVkms29cZ2RraMtO
BNyZL0QlDjw95TwjDVHDAy46C8QKU1GsJfYhbmDTmuOf3iGdR67DrngmqxOjWFDM
m7gvT7/7foS3rNnp3rZvni45FjCZ7Hb3w+XbBy20Ozb8xebKc6+fLyO6TS72LzIt
YGCA2s1FwsTEl32vX+gWyZC6M4EIjosXawUXhMJVowXG+at/FVVOSquLis/l2I/E
zK0vIoZytXo8dTh2ceMYlC/IkqHD3+mTcKVtf+S19TTdIYSny/nsD7Rej9skrf7D
fPQaHR5hFXOZ308MCj+dnlKxQEuAz/xu+LrGu1mFfMdqHiz4Y/hhQEATGxKcT75n
z8rt4nrPMmC8b0fErQSsDE5X2f92I4fmFJM4hruQYlGtI77zgoHA8ugYWwyU+lLg
PDL//HrDhC8dFeCYy4aVKu3A3Vxu/AvjfWoIdK9HbeBFQ8NRmJlwq+nxc/OJRY87
/78qTmAI4OuaFN/zCx+nAfO9nolG/XhCoKqC9g3ZIo5nBQ8VA/4vwHo9CoPZq8jl
dBdeQrh06vQEhvo94Eo4ZnCCBhDblqDYjcnGW9G2lyX+b2OEe8QQ6+/DgJkDqmw2
cLjovEAPJvXBhpcbr3IYXuoHnpL/uoI8AigL8lGImsAgQ/bCXM7VJB6zPxklbHvF
DjRw8Hv3xIgkgemA2PvwpHj32/HPiqSO448K1S1h6gcYMPOjBP0vkUXswkAkGEKd
j0rcYBNh/La1LODpeXPA42hMpkqjJe/3rRzLZ/HKMrS0ABTNDPiSgxtzlxXlw7N6
MEsJT1nyru12VMZw3Jb4pWV/wlMboeT6rAqxbv+ImEPEp0L1Zhz7jxlfl2aLN/Bz
BDSRHFzA+rBFJXW8K3LoHA5YiaIaYpACbYcV8/kaDBM4eHIcBeNa8sOVthhWgvSy
JyEqNfZ85d0pKCxCTwSPwvR4WGS/5EAaL8b16E/bwucPI+XF++4JdlYHq41DVW78
7j5fVuyEUESzDJS8TYug2QNyLqlHXvKzt9N7CN2VO5mfQFsJjTH0ZdrnC3t4tJ76
eIbFyS7PPqmXXM+1DdTz+YUcuaIZvA5ANLh+OKl4m6h1/v1D2LkL5pSE6NinulyU
v6YA4xJyRwb6yaYl5gmR/FKQkEj4m8xMlUmEmn1Njqg0COmK8TluSCCUxMOdAIZ1
2oBbMKYZ9sXvvAZ/OA8gAfSCZCxauPHcbREHlRVBFWompJfFyT5Z9+L0a0xqur1p
iiyZsjrTwoUI8mHiUTKMpMgedLKc2PflI9qpwM8/zPKrW7BYFwgd77OcU/ydLKl6
dN+AGrpDQUJ+gkrFLenMAGq3C8onvBYfLchShYpWhkQjxwKDE0jgFFwUj8E9HCAr
+o3xvMwqXltnjD0mvn05/DFPdfrphMDqB7mtGFaQ/P04mRAGKziBKeZzszBVfeWw
xXysViq4ZIdLkjTMklTo8G+bHtGSXEKi6ImQ175BZW9mZ35AD7UKuuqjHpM75YjW
95kr+TlJeL9G4pWVteYHTIp8n8/QJyGaarY9WAI9S0rhGQCD3UFQbVHg0YakRxih
9k2XtIPUXidTwQiGPo7ZKePU7oNdgGbCAhwaVc1iq5pYM1k91xcokCb4Jue7IoVl
uxpK/UfcztsubaykoL3a4IHOmB53OYuSjxO42KNpnQlLMaoXj+iD7nR66Zyf46Kq
/xFI2dfRrbq6UWXqCVhQINCYpyryI3TmGBXICok6iS3UfUBhoWv8Okm9OAZCl+Ac
KSiUdAwj0abKgwSfRew0rADkB1cG2T16eHkaOO2LXCqIDFVY6hvhfbXdD8/8uzDg
RevrSv9pYcq4DaZRdK5My6TFURqHzJq/k6zps1jx9QFc3cYeO+MXH4nlZY/R7Gva
BJHhCP6pPIoo2o8ETGi/VZHE9ksXNjMnrNiUmTW4sGbwIk7dgitR7tKhki8cDwqf
8Tv2jUmmmS32Om93T9Us3KDhh25wPP0tDfka7H8w5oH1QsyQhUlMlK0FgdCVi6E/
uU/NAMpmLR79AtkQFu0q/xpHAM9Wlw1o+Bp3AmklJoO4zbEEAkXhYCRL5joTBJZw
b+mDlvQ5NqwcDUJ/a7JybEQgSZDEMrlkrlxJyGT8QoCjZnHTjl2htbDOUp6W4s45
W2gwd52mdx0DZbEPhAvJF0Lp+OVP1+v3AGy2LyNuFM/tGwCJ7ctdgoYkQoup2Jq5
sqYP9cDQX2jg+5cbJgyo+j6QYqNft2l1+Ujqm98lOJ3tVYyGbAahGc4Yad7scU2H
+XNmvvUqggEB2eFAFfyWAtM3mu1UVGwoKz3AXps5njoVYpAlVXPq0CUmhHCBit3W
khKK57E4ReFxRsyacQeY6SBTRxuoqXqNSSuzh0xSa283Z12pNMb2HLDqKN8kZNju
rHV/u78LaJqQOYW8C9Xb2ZmtaAlei6hHJgYnhR4NjEkGqdTX6xIJLMLaJNfwaQkX
Wc2zTDH7OJgtsZhJe7M+lupiQ2k9A9teQKEBRBe17a9g57Ti3HrALeLM9OkKrw8o
2CDAvrIh8nzDmr0rUxHXObQY7mVPgmVgkXlSjjwONxWK5/47L7xsUjv+mHRKSPHT
0bi68hW6OXH0qnPSxJdfwLR9oCQkc6LhNYuIlS2+fWDOJxvZvGTN56moGOfqcO9x
DMdB+orNCJsHylfMp/pOGSyt8/bATnmiYcswnoAH0vtclX4D/RMUc6cYYP89yp52
69C15aGTc4WnIiXAX52MXRWL14sYiUBtHVl7YcLPt4lTh83gsUslOKGrwEHZq0og
Ezrzo010LKsMDYymN428cUCgW//BIKaUmdHfR3Z6zLQ0j1kljGxoKOEooxbX2rss
ooF9DgSVLVNHkA3YhtimcFjrnFgbpx6zAc4p+CdejuNnNY0reUFGmhPlrTsHFT2A
I62IsY/f5YDUmHTmk/1JqrITr8HNI/mJv90OJm+Ir1v9N3ENc9apcwbdUK9fbfPb
dmSZJah5Vdp6iT8gfjqax8xiS9bfaVsKyAoF8iYinXH2lG3/B/x6rkZjqQn1ewLQ
huBi1152gf7r1zlrqgQSDzw7d5NmC3qPXqOX2zO1LnMZoBrKcqzRbKAig39GD4ic
akxi7y+NSTGim7qt8nWT8+nT0j1xNQ0dihpl+2wRCtKQSeJS0kDViyxRkykNR/DZ
ot5HjuMz1+QLgXiOh4e3LHbF8iYH2rH9AevlfkAmOAQAs0uq6ieB2U98/DKhAOBP
xm5MhziXb5fWTawZJav0nk7CPdPAYZPXTHdwxl1Kz6LKBxJcfQARyi21LwLjqHdA
ln8EVrA4gh/lCP685pgrKAybScVrX4cGAZ22dDCxH+8o+m4gnme3qkXSn2XAluWE
X56IeCJfDHbLJ8yZkrBzjpfQWC5gO8DihOC9P31wjymFtxUtVkveXSbLaHB9ETee
vFV9J7X28Dq1rmGWOFElEwR5C8ig1CWSeHEaKEj69OQQVzDPNa1C8vrnnk4NTceU
M851VrCPhA9Wn+2FxIL86LBOeqcQnClOkHcOuOLAg1VwkcLsYtZYTzU2mBMZHlsu
nnzFKiYFvkvOgKX6o1q/Wwx9QvnTFWsN3+yjxNQft2jChIbKTggg4MH5p+5+YBDQ
OnFavKYAgemxnVbV3zJPXrRGZjjS7vNxJC7n3FmM6Oi+EEEIL1LSoNrhZEKEYxvT
cO3Caavm0Tt0xn/Dg+myYl6rBpgDNPbyr6NNVwB1mCmMTv+d08Ua2wJmKFwTuysb
FxmuNVPeznyPvExohbaeY7dgHdIZiqJjfG/4OBrZXKG5d1AGJ/k87qI+jmIYDoVP
pvKwqVPCnfFe0Fx8DgdGbgqn1YdwrHp6vFk5tY9SwwmJG1Wx+IC8zkeRe3o1ttIi
MSY6QCx9JbqyJTARY6XKBuWf7/hwQPi74aYj2OO/wLfr58V+LAV/gAnpVST99+IR
YVBHW+XvmEkH8sYICg/G6P/TbtUZQHBUm7Dmp5PJdipWxQ3mGHSR3iHEfwxzgT1n
Wz2VtaYJSPryJfTmeQk6oFz6jluO/YrQhghKTuyuuCfzjS/kgfas+rRcp3XsafiO
uCAd68wkfKpZsfFQfIgcL78xeMKU36rsat47uzmP8fQfuodVkqytscedBZS9jH6M
rTP2Xb71FTRc29UuL4+uERznBnCvgJT8u+buy0pX0hkFGzSNEgt9lqkS9Hsuuf3U
4+XfzdYU0ZAMK7Ko9sF/whs+hDC7g9KKlsoADD92hv1BAd/zlcK9bcE2+p92CtyL
o78w8ONHD5ESQ/3lrC2mZ2AlWHOSGxiPDEy6QfxRdwzEQSodDZ0SMramHnwul6NJ
5jF6ZgAfuvU5PwU7EtzyhjWUgLz6E+5z6dY2haIE8CI0UwndJ1NHRYJ5orPj3Ry+
JcGsRq8RyjZupchIF4TbuxAnXICmz9OmTrm6M3FDINoSimF076MXDkAa8MZ0DLt3
NwjmeRg5WsX8SnoypV2n5Vdd3LByE7bdxpIiaj6UQm3UKEZyGvYT9dNiVy3qE87l
E5whL6i79fW1Gptedm5qz7dT5Zehalxvfa9kdSllKsS3mWgpP2xG5qnNLiou9JS2
q4l2DbifUqFbgIdN7BHtQprdunDu7AFDV2iy+gpqXJ+usw53r2ZY4R6eaom+9ov5
sjusCRf6uu3BYVOiOPF31lVxWGH0Wf56hifEcq5FDzYn5QEN8W/XxoyxTl5MzL4c
rMITftKDeTtFy19Atr78PWNX6wVykMF11pCvFpJaVpW+J0hTTrF8KUPT6kNLeaLU
bivPh/+nrPQkole+AgN2xIWgysBiLU3vMvKJFaEQIjnrnfr5mmKExx0gmJfseTcT
K27GBS4ufy3G72gjxQPuP6fwgJ7vXqH5Ko4jwbbeRm9opmRJGJWt144IzKLcjjqN
V4USsLVPiHEvqGTGcXB16UseB045EnlKjZmQQ2AEMC/gH0XDoIzwCzLmUpTONnAf
JarxTOKw6jVY/a/CH2l+qf3LHDdpHwVtCRu1cQPbTGGc9S4aUypYsSnLJQZyWA+J
gUno+YZ9RDeAlVJVScaSVMspygTGkIBv7WqLNCnZNU1L78hmJOzkyqPm/Yaad7pJ
af5ZzateDOzrZI5Oe4NPaqEFx7VL40mWCiSuaZNxXrzjIJE8C0xtAPCG1TmkaVNz
SZ305tqH984kzugtEry2IGMMPSVHJVIa/iZMAtULaTveUFLqWMfIz6JMdSXkjPZh
YG9lU/AQxTKQBJDEjJ7zHZ8nBeThu5BAsT+xIM9coNUSN44b4bmF4oaiWD8DOoaR
BP5n59DTvT9FlwajmY6Xy+JZY6psIwVdXUBYQmrsmrsg9SxSSyK7opBTyqsQGOu2
bRmuhnwcEHdt4bOxkvrPTv8d1b+okMKB4Bs4g/b9vWoGBofqGrDGkhh+8eR56VGR
92pRk4G4HbsufLcvj/jCFmU17rxjtVdJHZdBzPTiaa1GSX5UowH2+jgw6gQwkvbG
D92AJkKotH463RSxL46ZfkBvVX2Vx29ElqZo+dTfPW/nKZpm3Bygp/YFGUQiW1Gp
0PSvDKkFJoBCiwuIQXxzItAmhWg3yU7lpoxDZFwQw3BcyLGTHWW22uy+qmQyakOw
Fa871qgw/0Qv/VBGMS20GQkjqvq8kfFFx4j250r7oDMIrXYz/H+/79b8HnVvsjD6
u2RrqUySz5x+8TQT+FYUCtK0XLglCqwRPans9V8vTvIH6xKvJ0ccksu2kMdAgE9d
fIg4yvQp5a5NGmN1b6HZ/XRlMliyZLsfSsTWATkQW9W1dOqLhn9Lj7TmfunPVErB
o2v0fz9NieqLnfE+ugaOAM5YWaHzQOZ8p1jXv90TsONdkhpUUa9+UTgGpZAKtZgb
dpZjZAHlmz+VDMMvh0QDQ/ROE6F0Nzz+R2Y/yuY9oeMrYWG+oHLvurG53PsCVGWQ
tilF0wBuNZbxwSyjJIyxIgHp3V6Yy0Pg+r2G/cNGS46280KI5fgYhEkyAj9+GV6H
rs2+YZw4TxmINdIjBJNUbkn/2oiCoZ/eKKdbbJIiuLuIvGv9jHN4V77Xxgyqlzy1
yYyOty1Sp1Ih48EZbf3KURiL7Irk3TIH118HhiVAPr/f/pKcfguryqe2S08miT/i
HJNju4RM1cV1771VRT2FOhM1CrdzCWZ/yIDnCJavv8KwcUkKSM6aMMO59jfD+5Vq
ua1AdTgYEggni3qeovI4bwGmed7hZHLU0wg00wHkmwjqlZOWX3eJP9ZJsEqNwIK6
P2WyphoxPvtAzP5zCkY0NVHInYOveN08E8itiycms2Og9iCanQCCFt8c5noheBWN
FOI94097rsLP2mRLmt+q0McK/MDJBwH9fXVjM8GIy94B2BNyrni7nKyfduKsLHUZ
963k4gjFSgFPXRMbDlf0WIF5N87MNS93AGphR10lRJS5Vfq8IFvJ3l7ap6vvpdcE
nAco86yLzQ/SJ48mA4Klc2UXTWeP3sW/X6LA367lfLKG04bnp4BP+STdNPrdzBbw
F4+o9dkBJsr/Gx+TAZTShMK5Il0xqgSoY5y63V1qjLHMMHAtOECWK9mCiRosnGyi
Ov8Ff+D3LBGOtZhr/8t4bIrQ6zUbLRaa/vl9eGx/z4bi9XhohALzSuEmcXkf0l2N
VtyY5LjOMFMCcffYkNVERVwH6M0RyRhg/BNu3pbcSXmgMnN+uj1To99R3pSZh1+u
VbDF9s/A6wnFA47cahjv8yjVZ3nRg5JR0er+zpSg5eHDZ1iO9T+wQILpeXU5l11w
2diR8CLZARBa3H68W6h8qu8cr2X1jWyMcQlsrhtK9XIguJT9seuPsRKXFENJ/rig
7MxNmPSw6bLe4MThnuf0AC6i4EqZqPj4itUvdffAzd5nmt6QDeUj9wa8uCJoVCB4
mAwrpZsDEzxJpt/p+R8mIzjYSeZLh1Ha/gzDx+Fgu1wZ17GBmrATToPnxvOKS4WV
w0KKro/R0SWhz01sBNfQ/ESBephyqkZVFlPrScRsxzpA2RAPHQcZ6vQSEb+OMlqH
ymCHZGwKxGeyJM1/QKFOcJNkQ8lybcln43xBkN3xAkOt3IwUxVTqVwDjDUxvGkrh
TyUyF1KVjFpkxx+wL/YTJqQb4Y4YFRqOvQD5JlmdHbZTh0UMJfNGT5bKAIBMOry5
qELkBY8ALHlhQ+kVw/c0dzChqZx/tu/7+yj1jz1JqWuOGjO1+fbVMKxwT3vv3ZX7
0cCCjQZWZmDcxY5gGsfu4rv2GJFog0oo82jg/zmSdr7N2Dhsl8Lp7+q/wyzjyCGx
A+1kK2hE4SvKJ6Mmf/Y2Ki/SHyfICSiLqfFaz7T8iTUd5bRhd6IBHL+Ta6Btp6ai
qYyl8RtHm+t+AY/Y6yHVJ+xoyDdY+IQiPGzk+qD35KVGq5BlfMjZ/Z4e46Uw3TYz
dqLVhAYWlII2PAvj50kC9DiBDuim52XlKXIvYseTRi/k9oeKgAjE6lzZaxfD0LEZ
RxUIQe3VHGPX/XJdNEALJ6RGUmBQLXzwei9V9MdInyHWVyaZcbb37t4vgoW1DW10
y+BDhgUvZV7ED9Cdbz6tlbjO493/2+daPM+4HyPQtqcdyXhzT3uVPwXNIf6GZOpc
eQOau4UNFNJUNd1WDNweOXSxg/Gz26SJy8wYdjcNSVvicaTPyLpJfKhp8CtDUmeF
g9IkpbrOqNkK96zHI+CukUCB1RGfMx0HAa5rbuQ/rTjrV2oWgez0Gn4nJeNXKAbu
enLWqr67DlEo6zEgNNo/QMwNSuQ3mGvHEUeJHVV9QXC+1githSPqG8sWCSauaCzm
uOuejzND2L5zW3cER9qDS0nKLS5hT35AiG8yiiOgN/GLptCNIaHfkfPQSwB4gOa7
tbgwaD3+HtLwMQ994CAPTcUcB7Q6cCzNo4CuP4R3I/YUs0jkQwhb5/h1EuP9dm/z
BcTGzbmmRa2dhz+6tuoR7oVGO22IVm/J5Znw5ZgJjtGbtQFLgET4h/h1q3tis5oP
My19cvFQ9pc85641o2FY3ko8TYGvjsG3mbrnt67qzv347sM5KMU39zVlW2BDKd9L
DyTQxvQZyDnQjPipUhAR7/Pu95oWLPHs11G9Hp5MV4za9lhoeWrb+mmKMNJQg2lW
mhS598zV8bsWvnfj5HPtNg8jxtwahCH2K8NV+nDe5TFoUocGPNstJM+7HTwq4ljh
XbGzgEdrXUaYKVqtN23ZFBa5hXK+++t6HzS9ZJyOJ3UZEMxEkrWzxDmF2U9af5lO
+UeTdQR4Ytx+kZsrahtpEOOYkLRpmofUE3mqLskzjO/Oig2PPcH2BQQ5Io2NxLqZ
FASK9BRiercEQvESyk+fhR8gb83CBlFpcLVvQe6vHaYRYqkNK/aelpZGNJCzSXma
XX+qx7Cw4XDqjxginzX35CxSy5gP397uxr5oiA7TCfQWsCnWm0vmTTTDbaHHoGas
ZbPHVyE0T+EVzSZcCu/RHDQUAXCB1LMvY/gVQrSq609uQfvIp9e622l9cHAYZWhO
6DWnV1btgeB051wOOeUCJUef9lIHLH2BdXdBOIwUEi7zMNPn8VhuHVnkBP3lznes
z0NPh/j/yuFJ3nLQQee6OwgUgBWv2uWRL87N51bYGz/elvTCLhP5ekhyvPD2rCVU
zsIOYGd3DLN2jXTekocQV0PuTTu0Dim5yCYhkN+wRcpKDF+MnNOqEYO+QQ/51Kfb
jzrFF7B6gNMESkS+Kr53TaEQiSocV1uBmcLb4zaP4T41l1eoFFuUXDuV5ghRzYID
YG4iUx0ugqgvIfflwRTYA1zGY1Jk9q8O9EmUwqLsg3YgvWG4oLJxztyWNvH3rpzl
PZr69fGf4SyYME0SUNxQ99if46XdXEgN/Qv4XxXpLPqN2ygKjybRKXUFrYkP54hu
SGbPetb2xWwSxlceBFMFKbx1ZK4X3Sz2JEmtXPOY40OoVzx0wIsg8ixgOS5p8khu
qYL+mYnoVYmZRsf5fY+rXoSWTxOoAqJYfYIt2zKiCr+BCa3GKz7gSRuChR5CEsRA
ATRGT0wf6DFCUcHLbvAHynL3H8JJS1PYE6JYn3tfnLEGb4eXTSu5O8WmUpNKkvhh
U48ws5P2Yml7OuG1Ndz+q08cUD1UE6/kkSVSOQ84VUJr1AFN3ruCSYD1n6R8NKoY
lSuwf8CKmXMsDl6cBUh/eRjYGwhXz8Y23/wq6xjOKRkrN+OZdSO4WGbCU4hGorL1
57I9xtxZqwLoSvFuTOewddMgM9iusnjFl/Wt+SxfS1S9iR96cPw14Yof20KfD/hz
3tTFfgxm3eUSLlm2ZzyF6GFTCjaCxEGqgJpKDrzOmXt7LKAF+hpIXNCBw4gjt5tM
ElZUnM5HdTRC5Dgbm30H7k7MI4Ka5eTV3zvcgka/w4aP2r+UXr3GpewUezdBp45P
gdzsTCIaWbZTBlB5JTlUZc/+cFshkpw21K9KqZyTSW8mLWgcNXTnBalpCyyC97to
TaL9HVl5OqO0+UDgCxXkv0sICPUVLOEU8gOx9exCuL6dtuMaEAzGA3VD5fwed2tj
KFkfYLdyXkmyC55mKtIxmWtMOFtHtKPju9LielRkjnFhCxK+RqaZsxMh21XUbwg6
30yoFf279q2bciHHcMixezxCBxlH/H/1mUASsE0zIpvBQ0u+z3zhoYUk3PKAW1So
BspQI2KFFtdpDJrY1rHtLbBNPPuUzQp9WlY17b/0MvFmPBv7wzwPuPXMOahlCPhl
200AI+miEPLuJIR5DDoHQxG7vlEYgerc0LDDFIXyynWaWKFL8TQ3Zf2BXq9v+/Dv
zUUldmLIjQ/Waa4SZVZUZNbi/MWbB09WdswLJc2i2POvus4cXnTK5GC79W5IL8L9
kQaEESvOwfaL0SKHYqBp4ODhuSjGhwWzGWnBjPJnDFpzJQJS880+RtoZMU5KoJvd
GV0/eVUyiyLJS0vT902BvImIjB6WA4JYAV45s7sxXubI5yF8nNYCn+M8gyjb/7Tn
OzJ0T6x+IA691weyFxqW8HV6r5n6aPL6pY1cAgYESqsGxv6NokWNuq//Nsqj5fDD
kFGLh5R5IhxBOJW1QcscvoStupOi8qbGcAjXr6cvch7EdZ1+5q7UOQ+RTLK8lNxD
DVwj5T2MZrIL5SJA8lyRUuNIa72/lTxOMuo1RT9du7XMGxRvMB8b2eYGI01EQLoz
Wrn23EjouxGy3/Y8yWTyobUKcZt/EOf6gDmm/XfPdiv5ycHydgA1rCzsnGpPlNtp
8BG8/zO68BqOph1+yLh34GU3E+BWExk/HIiV3VtrSyCXRmZrpte+04IVpTizY5vS
VEhanZ6NhD2zC82qVBGdY1R+pJGp/nCj2UFtLxcyRKzC5UZA/Z3HPvLmSqXq3nEZ
ftj7T4hXsN2natcEty1ESrqX2LGwtEvQG66w3ORkCYLdYMq+xDloafOt8ACiFZAn
ksJrcdGCUmvESyeLWutGr/JIFwtBjvtLWH/fkuYFCXpR1nlitldmwNeBa42j6fTi
TtzJ/ygkmBfxQ9hz6dPrinj6MZc6c0q8/V7Me5ehbMFFiP4r99u7Inud5lM7HF+9
mC7MDi4wmomQ78LhyM+8Pn2kK+V9RhAjx4mI4qqzcNfA3ceJd0PYdtQYypRwmcmf
jsytWYxCmc0QNfas0jRnStBv6YZY7CxXDK7rRiAPHUgLmKlc4YYPYr/2oW4YMzdi
mI/SRg8hQB42tIm/6bmB6/Cs5pyMSmN7fT9hdIa55Hn+dQqEoug7e90RQPh1ZAx6
1YMUAaJbQoP9UCGA3wSLFYP8ip4POvQ8l2esvx8/jhddoUkzmgNsJcoesZ6w6qcg
lj3MZ0ZZXcFftHSBP5ipbwXqLq32iEoi5JSv0rIcaaWcdRRLNxTQ/P/pj7TpbhZ2
ZIodxTh+DBDujlDZKJueiBeDgPIr9FRmq1UhgUsdwln20RxnnWxv+DtKv7qFn8Ui
n4armqmrQ7nXaBtqcbcwfCSr0ODWgaDK4LV5jWUy7KNYgOWNTE1KjpdtP18EEzNK
UyVD3xr4nJsinbJUluoKJCahvlZOuVjfwg37lSuzEaqGcsUCMF9++P3gmWAdRs8d
BR+1cJFkICRymX9ShrlSGgdppkUSDUT61O7FNF6WClPowcLv472U4Hobl4Rxo4MB
U/qJtnIF8xyvfpL0I3jptG8CTS2iVmeMv4wjIc/yOHzxaJ4JPVF7AD55Id0RUYWi
gPhYwQZkmOHbP7r7RdG2A4r75mb2zKC2KDokW/nF0TaxJXNgAv2YZConB3A1xDwz
8QV5xCZakzfzDps51okFoxGFfsnTHojMiYpyi6mwsOi6uHpUdAmiDWk1FtKOzhSn
/zvRqau8QlSO6qxfhmcjP5Ju+nlpTCDrVdQM8mF6TinrtPG3crN7LgTEOMiEDI0p
5F+6JnyjAvqsaFa71z4sVvxOshbEoWAO+ieC3M6iyzho1O2LdexADEmP55EfacIR
bPyoeYDlBudNBhsCJ1bOogZ8kBVngJT10T1hLHvINCKYDj0RXiCKELxv4Uv/vEtW
Wo2UDr5zTnHpGbR+urj5jJe4zCU1hZvJwhaxOc0MOGYIojowAuKkbtWlMA/DplLV
rF6sHt0hwDIZbJz5iOOgGUT3oo+3R4u7p3ltDVpacufuOjduxduWfeXPWHYg/pg+
JqeA/48cqATn6kkwDyJAjLHSdmoavGEXExZ6rq41fRoiDTpptS0ZrLHEqMa5lqq6
RCHv0jf09WHbEW1O7o08ks0e5YsKPi5JO4zRFWVjynAwUEtXEyilWpUU9klUGj3a
rkj1LZ3VlbwQxCPfaKAqT5bDHb19zwdDKyZ1+1Gr9Hd3aptSkOMyWGZ5FkhShB0l
p2ygt9LBNiWdcqhBBWMzR+1pRObPNLB5LuJbY+qveyh+/XUDNE6vzGa5T5dN25cr
JIQbGIlmQu744x/jiGcdeyl4+I45ZJeT2j1IpPgsNO/92TfcBXGQ4yXMpTTLJ2Rt
CuT48c6cUF9EaELzzpcmwfnwhrx/tf+VeJNECD4K+tP0aqER+h7sOndUSFWEb44t
kI3w9e38/iiiJTEQblYgfxsLJQKyC8scx52oOm9kpU4yWlcPV+FQabuM32lEQlhz
b4z3I2l49kB7LIrtFI8Agsq87biQEgn2EncooAA2Hf511TAOMcWqsLCmiZjHiZn1
Nc7BXEjBmslNOYDawepeQtUzkHFHvzZtlouEYx/rtnaAPFd+64V1/RyLt/PkF5ir
hsoNj2iFTI/kuSm+RxTgzcyFwywwHdK22/SyshcALFwii1Cbxntla4Tyq++i3/yx
6GNqwKWXs8o35ylKk/g5CzO7koN36U1UVkX+0hsWaX2DoKr4ElW4TBhbhmxVwq0q
fey9sjQQshwrRt+7oKNstyHRz/10wIO0lh4W8a51U4kX/uXTi6XBNqO0pzJxZqax
kc6O9x8NToKspM0IBbA8L5EFzd5mQgaCmG8+Zi3O0QbAp6KWvRvZLRyQtmaQZwLs
rDCnrgeIdP4Y6S+efPPbNQ7nSnj9pDwjunwqrdH6TD4NBtEtzR9K3eEsWxSCXrDm
c35m4b4dgcqYNTqMQA/udcEncjtpLt83oFTL3zVt5/D7SiYrHu+DjoWyZom5FcRn
R/DplsxL+05lTJezuWCgnUeVNXNNYIdhfg+e4jr2F6albzHu1qeJtFxTBHbStd4w
7+vasceK/IXqLJtXBtof8Mhsqz/G9M2NiJtjCJ0GexuPgYFxFdVg1AVVHUuM2F1z
KhOP1ho+esT2pWDE0/fvRrfZTljVmz2kAemFuc7BYwXneyjhIvR6JhKOk+8driy2
auRFX+m3br3ueBuRueHUK8ocn87ufncIA35LBjGNPysJnzzrSxqh7raWuKPhTX8w
seMHKTfGhJ/5G3B4mPJn6QYJjC5taQN3hRtwR/L5Wnne31fOWVhz2W9C7O+NHNWG
BDHaqqgJ0EPTb1HonsMkYt8HM3tnuovyBa8C2Daoc0YIlCQnnJPjjbQI1cSNmCTs
A6Acfwe8QreW/qUGXeQs7ycgKfuVUsiADAaLfjtV5gVhxeopxjzoIAO/VZGE05cH
3a94EOCf6wx0qWXQh4L/YZwMplrJpSMnfmTINQJKhl722QNglJXkKWLWtF0adISJ
kxXmXrEcXxpcyJ3cVf8FOLIceYqoiZ93OBD4qqnVKm4WK32ZpJ0aZeSfBhUOX1bJ
HpHWsHaXM1vkERhAY0crkvRlASwKvNltcaQmkfhQCQFEtQWxIA5/vQIJfqCIBU9a
lh8cPgy9AJs2ZNNkSOwUQvKcwGFOrvntu0qhKTJtgkX0Sin9PXwMMoIEC7obfD9o
YNlQUpip0njaP+JAB7wk+E16fpbPVOWeIfLF5rd98z9YJ3M6aNE8v5e+0lYm3XzE
FMZN3bwhoK4PtCdtwwW7/fKLOhNa4NA+YclZ8v0/IP78gncgZ9FZ2DTOW82EYpcn
3sNC05jG6HSJJ/6ABDBlX0aiiPnvT3ulc3f63LFANHVx9KAp0KaVw0FuqUvVdnUk
uuW1XVveQue0ghJUx9TESnA4trfhNQ5bggO6RG/cDD/iAKjo+0V0ESB+PZfo76z0
Yw9EoFYiMX6XltnCi5kQW1M6d2sm1jLVVOLFVuF4n7xvt10ytP2vxacJ/C7RbNoY
EFUzSsDZoWKRqsgRWTjnYwa0VDeE2PGYje2tNuzRK63VHmt9ViLwVRLFPYLK+DK3
wHVOiwtnYDJWKkIASBRRDIZHwAup7UZIqTWy+31UIr+58MJ/E0iMMx7LqJWDrH5W
LZ0nPs9HvryKIRnsRdJQSfwiOt63CiyExIBxm8mv/gQqK+4rZdmMGyl6tOoAlvZA
46I4P6UZp/+VDxTZn7ioMfZCbllYRUHqrHb3HZzTwc1DOqZFzov0sxUpwpwSQ0V2
8Dq5I9EXqFJfkHvejWM/6OaCQwKPuLwhN5cqKaSQEShGznKgoYwuAxbzoL/S2CQ6
fvb8jULLY3IavZAMeZjlHzd0/Y0WeHNXoVB7K+MwFRmWecGK9aE/sOpF7jrjNK7Y
X3379gT0xeMbw2e/HKSjUpLelZmzE/1630y+XIxWtyfvCuaEtslf9Dpqn9NElsVp
pnm47wdVlgebcdSAAYxSLCs0Mj5rmc+D4iapoM36nPV+yIIFss1R71gE34DlJ2xR
vsUG+B2L2we6vYfKyG+PvPMM73wC5mITvX++nX59uohyCZzsC7AEzbamiwuWNfoN
eZI7LVwTHAeaLwbNiXa5fW8t+hznAXG+w2uobWw/Us50Jo8w0/Jx9eODOqqCN+G0
m6MJMLsTUx/wGZI6p+NTzWLolSJLtXV3U+FJIWaJJWO2gQ/sp4YWeUiBEq9S2crH
3QDS3RV+tSExqvo+S71XdiyM2AoYQ9rIEtoP4qh5l0hJwfN+SAM5ypgYbpJnMTrA
rIEYfMi564MGESaSkHtJ39ZSp3ze+6yU7FjFHLXR917QuzDOYiNFGVDO1Zi/YaQJ
rP27krPR0x2ndINLxFW1WwUuTh89Emm+kxm/e4cwWzJzdWyvmKy3RvcknyN1weFH
k50irWqWT/5Iux0ra6iI4GtCkB009+hRhJpQb/R9wBCESk6JTwuWmmEiP7NXh/aL
YO3QPohUkUhVNrQjaJph7s4LvlDM8anD3HuQzMD6/kn4XSpTYBU2SsQki6Oc/oui
578M3To1TXfIiMVHOXl9MH56UAA8/9nQ32OPHkqJT55qdmhVX/Cd+X+ME8G2GKMd
k3VokA+P/l9DtyJr6QCC+o9zYS+cDjpk4QCnkBahbjrdLbnA8V9QX62zqvciND1G
ddwP2x5xK/EolhzTHhkXCWjGO0G9r5F7RFElOeBYNkDwdRi0wRDUs8MYcabZuipv
xJeYEre7pa+ZUTCganlB6H5A+pSlTbdopcEenNpmYNxH3j9GuY0fx/NUx0UrZ5Th
0Ao9d+UZ3jPe/s+MexVKF/f2PxH0jA28QoT9YkFntD6sYh8SzMdbzeP5+/me+UV8
wJlZ+/LCv/+g19o6qg1bh2cTv7hiELkh1QYMkYtx3h/6gIFZJ2LKKvOq1sBdZj8o
dQRBe7Yo5WjQMjMxfOL/VGNYmGb2APuMHHxr0oRX+UrPOaeZOkf9DyBTOjGigCXb
3M1JUZxgPDLwP6/jx0Y/zjOfaQFjouEIlgmPB2CBWSvAV65kxf3S4SZWk69hD3nm
wLwJnur5Bx8Gw7aMDdIn5rhX2JmCXXzy632VST7OZgkiI7fIKntuHLsyIvSvZ1bp
ZOu+gHdP2jIEsIl+fqJbBAx4pBE3EI+atImMVwKRyQyhT/FJp7XGMI/UFR924Q18
NGfI0/GeXzpj5L6g1xtGJDLtbI1EkSFJtMOMRAurM/eC9FOMGcvYrXqgh6GZ9TaZ
TvRf94GW8cOJDJW9H3wcpcYSglfUhbbvXIed12u/hc4gN0xmmlCVpAfYyZ771Uph
2P65lrEC7FFiJ1mARszYVl3oCctovT/RKV7hWMKQ1E7Nu1PH5I9Jnp/ISptRfOUf
ubJFFbIP7H2WGGEz7X6VNUaPC/rU1wzSyuMW+MOk5meTfGVpTjSz8hZN88ilV1qE
Hhd3bK5xCJD7dZkbgA7RPEAukeuhHkzOV7PefNoPs/JHKMA1uD8rPMk2Zd7yc67F
XQoWKT4qyWePf4iyS0p7JJc+3ZunYx9d2F9zF4LEEZTnITYVuUEYPbNwlani7VRg
cme9PCBBQlyWNYLDO9+UfUzg/VvPpHf2WHwsACGfZFhwJjihYunuL98zFsv2DAdg
zGivNGTNftQgmgq8qOjY5XLDPoIncjJnDJvWlySROXCcfShf7Ng4T0sdjEx6vhho
I+vhxWlET6ljEbWyK34SLlWkRRbW3v1EVi+RJST0DuFT/xFZyQhzpJNMq4fr8HC3
JZv1ydXoB/6sNO2h6BJGF5fzTYlBAx1foPbzpBebfG80wkmqvt/MmH5uJEiFnMui
aZHMtltD4RGhhpLXFe8OKvpMEsycEFEqQweSDbE8HwsztgNjw9wSIfd2ItPAYY66
kgHUp62NjSU7gvOpwttO0tRCINFzxCqsmgsNEiiFsadypfatClFK0ddJI4v5GyfR
RdN405nHYbMNJ3NJ1JvjjF6/M1v3dSxHHaF8MBefq3XTB34v7NeDS8YsGSUw7g6b
2IQt+6LwBk5VXar/Pep1m48V049GcIM44MyPzXDsAseGkt7OnIcyxhSGMJK5evSP
G8LAdobt7hPRjVHJ2cmcxcO4+aF+kximaejQVLmJsaJhGA9kUcqikaRdw0Y7NqHS
5qp9DjFM73HDNze3cXUBHj97z6WzBkKLYIHgjeXyZmv5EP7DS6x9Uj0n32vH1co/
Md2j44j5mOEzm20z/t3C6SorI0zh7SkupEKoELcObK+3SHdxIPGONdS/ldz9m75V
WSfswHHM+z6tuYLpfFp1VAOAaad4sWOKWB4XMqNZzyAFHRpH786TdVvJ7gbdQnbi
EkvTiNooOMG+sBXOsp3mOLc2EAV1uXfZqvLFExdBBjxnx8iQvOJzYeIWjIMQ+ZP8
/zmQU20P8mcC6Nrb0NLF/wCAZejxMxFYYPsDmPrMwWuKMStHQrfJRUYSp6RFJmE/
YHsn4Tstt53eOegQDVTwMZiv062vWn2Gp6t7SK4GCF/E4BvvGFGKLi59oTDgCwXY
GVabYUky+++7V4EoVLZI/NLLp5QuGhJzGVTNEIH1YyrRhXZMyONOmhKhS7NXBdjD
SiyBoKj+Zeeh3sw1AVnu11JMFwYglF8k7A0+KreCDowoSmrSnqhY583iSglCR0y2
psvVX9OjlSITOwguTZEaC60Z39LSslyA9lrzERlabb4gMudwKrY0lAuSCOWbAEFC
a/nHxyxhAsoGijWPYENTMhkQ8OPgqQ1WnQW8tNv8O0hdHh0RhlG5y99ST1EFLi/X
UDSK9dhPO+q1FaZFX3fqlEP6yfWgslitLUWHEMlvht9vx6OJrzg7XhGFQpyN20A9
we6YlLd7ZUXOGyKSW2haldujKDBCa0iZZE9g22HH5hUGXrAxCuesHnitk3ieR9er
AI60h1OolVI4Rs2SXdXbMFFjBNjpW8HNT/FRlEiyck2eXnrQH/ToCvuBHU+5oH0y
3sEaCsLxfQqcUXhumvS7Th51bTm4eh4/3S0NEMa3tT9mBW5J8JUpqxf2WhTpzT1C
kqc0rYafJfh6Oc8SjcoJBbLkTs3HMCKGX+xaa8WhlUBzUsvm/cdRif3SHr1cF2Kt
6yk3WxWT5++LYEzteQKTRMoci5JzPkVtean4X8sBLw1QxMvRwNZy7ynCXfYI/+b2
EWObK2yc6r0MrX5c2MS/rl3wrpR+ygDMY0Jydw2z3ySfRxmGqTFbJzcX9pbLpkA/
UqBY5tUTplaJwEEnb8K9s6vj/NtaIIVI9VcrJfD+ajmqIlWa4YQxaJgkqoEihkh3
/eUQMkBKwgALtCpY/msvohWVqdD8Kh7zhGz/QgZF17YeLlTQK63hiLcJJ37ESfgl
zcw0Ez087u5bRSTBxAoZm+aIiPXc4GTXwJLviNTWsTNKMfwhi9+fmiqvwii+fgx0
N6Zx/0o0taWBQG2+BFzWw8FzsmtTIlNbu6+bQWXV1AK4iI6Pre2zCtoxVVLwV1++
rfzX99QKM66AvL3K/Wst41xqiuGr66jsgjp6NnKCSaVQIW/WqrZcBmKupiC5ubVR
4nvuXVpEQsdWhhWj1DI9s1rbNrmwToCt6OI/EWJNrTDV0BN66n4Cm+xd+TkVKCHX
LUOXGYyg/QExPLr5XwL7vBVodlZ83zLJXrrGXdSKwgMgiIvL+BJLwZ+tz4qlhHqB
s3/L2N2Z6ftrCKWpXc8NNYu9BZdwmWYl6Qh8QONEXKyG7FSJCIyq3qt7ZQXyT7pq
Qp4llVVn3AlXRHXPdYxBdtezYq4Vu5vUp5Ial6LUMSOcjj0/wWjRS+h+u2VBrN19
NEV/LbFH9dtkB6C1Lpdt30GJO3H0e3j72plkJNBO+EHOnWsFs98jpNIeNSEUsceI
FNhleluC+1VBucRz1VtO11F9vOtvkHHPL3uy8TT7AdYhfki2uZTIF3Ef2lRaiDGV
/yojKLtPAFyUApDUP7bfCJzFIbvSMomihIXJ7lfIecsjGXpXefT+DgWvtdm2LdLS
tnKWLIYnerDpkOhEFuUyN2WSbES1Dbry+twCn/rHQa2y58vswcHh1/QGx5nCPAnN
wmlvNizMEcWX5PYfKkp+1uruPXy5n86S9g6IovMal+2wXWSju4rxxB0PZ9KMpM//
vbEKxmbUic/2kKc56MoLZb6K2+S/FQeSqyVaXGf7RNTfe22LcGCrorM1nFYN0HM9
QHA3Xz2uEu0W6rLp9/0qA6UxqUKEkmgP/+CpHAuN0y8RXfJho+q9M61LffqK5LQW
am3go3CVfaIkJRwZsdDnHhvqSWnQlcem8af/d9VWJ/v9q6HLBqVgAPwb84lrNORi
NJNuPXFWvr5/K1rS5GLwgjnIK+FT81bQfBy4fiTc2Dua47uZB9ku28OZ/MY7D4yv
dlDb57i5IyrhJPVLMnPbEghZMfbeg2r0JI7wLpz+63YagXy37VgOjp8Ofin3zrhD
0q0joC+5vvqxYS2a/zACycsoHgqPXOHiwM3qDjXOMSJ4mWFIBMmVcwShWFofhmyZ
mSnC4HwSOIrjEKQjf6AlhnBLlOT/BQOGv3DulGEPUdxydux1gI/d59aewWis1pFe
HWM+zxz+HE8c4mZUoKYv/HCc1INexA+xS9Zhs52HVyH+cE3s1fCX31lkVQhKNjNR
8Nq/EU5xDAwQpdETHoVd1sf9J+OFAZCau3rb4uoxDla6uSoGCR2wCvTYVJf6+O6g
f/4r2sVpxeFAvKXu2MQIFShdlxia81lnvSRWWTXTSm23XXYrWiLJy8Ue0j9JV+Sf
mHlFEh92ZXPIxzZuKW7H5T0qjTb2JsB6izBgbco6lbogWtAAn+VOuj3rToKSF440
Q1iBjhXkceP1FE6keG4IRbN1RMAZfokHc1gkao+lolRQoIPh+9Pqu71S1TbnZA4Y
kBduGnP4lVlvQK9XLO+FgUGXUWo25opvZRPK9W/cPZ02IsNqHpBmAhM6FpsjtF3x
4mSkXyriVtQ3F/jBF4HNr1tRr9AY9Xo9xNO4igCWATdOLx4WYxvwljuwsQ5Deqw6
0Hu2PcJXF8HBl/XMWNwpDoNwxrOzkms6/7aAUHCEWHZJW12RofzFvu6MGw9eKhql
vDvMsbrFkdPvMNMmFTe/hRVZrQnSIBNY3ihGV9yN4qTzlbWDcYB32SvmPhOg6J0z
rYMADkWq/q0V7+SiubyBC80g3fLi8JGF7ZJ16DCYzHv4VQJMONAyTlaS6zGEBMAl
rNHoSaxW1tJVqXuphiHIWYEmHjCqBEOzRDDh7zL/tJJNWWTUxljWj9iMXpkppiQb
gD9LY25XUdoCqAMu8f3wFrx2uGfFhbzxUbvUFM1IUUB9mvgil8McOA75Z2meB4+W
TUJTBXiDc8VoTL4dGBdrm750arFSJ3WU4GlWtlQfxtQRJR7vrpmwT+pTMS37eBfL
kcE4WfKuh5DiElG1aa8P7MKZlpvzTelOB1El6R62kk5Kf1Vh5F8bKfee5J6CQJbc
2qSAyPDOq91KGeS5X8Z+cn3w56G0CainWKB2XNXSRp0Ctw6BJBOJOb0gIjdXcY8D
MOcMWhZtV3Amf2X0bzzHMF/qx75bdQf8LC1BFyQFHEw6DOylLBL3qYTXfNYAPR83
OT2QymbAYvBh+phImxib+cLNdcqXLpXCSotKga7Mk6mSrW5qwCOacBMCPEdEl9s5
VMMnBUkcxIUPuqEnk1I2qwnjfkrCbI+754CIk6LcygeJwTdb8QG268PTKhh8jAIP
ujlmk+LjVo9ILfAN5FUvX8K7JyfInzcpcHV1XAhYQUENkxO34Q24rxcsbEpeFVP2
p9dTuC/5O+te9ljgNaqob+OoOACY/6id7I9PYrzoB3+zl+w5/ODcEzARS+toc/Hb
XB7qNTH9BB7p/hjTbfLpLH9bAAPqK9ZCHLF5Sbv4uHOwClisF+3gGdP1fN3Hpa4O
WnX89AMdHKEdfs4LosiTBmVPuPVxOvoavtk5Xck3TEX2FDTDBZLXaosY6JVvuhha
0rdfV94Gt6igX6GWdj6xe3IhBrHEb+cl2d+RbXr71NGJJIFJVsthTZjdlrbZg3X0
bG8HCVIjk03dY12QtQSA9Y7eWm8WrTr8V55gt0+BAmP1vYKzOxND3pEyA/HKh05l
iizd7uYjnGf/7gqYN/83dkyB9B5zIy4bjmPRxvbj+4FBTG9mVQPxOlvVjhrVB4mO
A8YoZRUOp9EvqulhRFnOEcR030ts6OfhXym1sm+ceOsNS/O57AmIgMqDcH+4tEoC
tzNjQPRrVivfbqezGYo/bsJg5EqyXdVfBnhTrLiePzaG9hwFkrXBsKfVnleBJ7bt
HD0G+Dn84QA2AtOi+70BA1calVTNFZOjQJp3cjXPYois7bKX3bB+a5jKzyn+Fkcu
rih8koqRGLufnYQy1+8gxAKuVyOm5TPYAVqNma9GlUu+g7L/XCP6k4Ou5aaShWEq
xPP+vbb9eIJqgVsXpJgk/92yz+ErkcQf+LXQNLKUrQZVtBPkVpUvPSxvyaYLu4cm
Q0FMGkuzfQwsktJ1wFm3BmCEaoQj52nITbU/wtmNaztVLb2DO/YTrOKnPGFIzScJ
v3TFWLCUZy/KfMp71IFt+7Fs1xxv6S9gwqal/t8Q84cB71f81v+8fmwin8z9E+cX
JzCxeotBIG+/lnwA5VNXUA0YOx2yDzX/TB4nD5O6/VlqzRRcG+s4pOzh6DkZ4W6i
utsubzIAn0JYZAA/M/iBAa0jSsV1SbSvgVS3hAsUai76kfpAuBzU9jVsmTY1P7bs
pP3a2ryi28wZOYbDDGNcjP7sdCTfPV7HEdmrDDbE4cxDwtfYVyJdzGDGWbrOU58Q
DXTM/8+PDOCKuxgyECrp/AXfq6nVzFfrctaBvPPx0Z5teMa+QoYTv3u51sMKGqHA
8DTUYHSS/Yhq8dntvm4HEMDLORNuLNYUiNpxLE9tIWPEzh8JH3qMsttJzhBBHM73
lAMSn3dfCyQK/BGyI46+9rThGJYgVvABWQ6j717Q58f9XraG7bZsBI58boSFltKB
5QlbVFMRD1p6D1jqG1ku6wGm5eOAhA5sppSNKFLDfqbXWc2WKUti6Mw04KMGiYed
cYvdyCfMbLcX/VSxNXz/hpW5x0hJ7EOs8Zg+7eeKJmUzgYJ076+D1gHNJgbKpdAG
3m28KJM4PyXoh0sEepRqa+7isrLNN/FVHiTOErZx70/yZ1hPDL21AjIhxLLIXhaB
C1NJQUkg0+kwsgaDTXMLzVZUjlPxemHZh6eOp7zHddrlCTP0WeeBD2n3kAkbmqvf
Pu7amb4kWN13H+6SoDWga4/45Cfr5Ke0FZkr56RSvVvK7ftu3zeoVF34oK+5RC9N
p3LVJWNd8tHkkT89/cAA/s4xZ8qieqz9NEepaoej+ApvL+2faJlNgTYcdltP+ZHK
Ytth9rACfcjAi0qwUk+AcJXHWksiz7NNNYL8XvDWha9mI381FZG7KCwG/EODktFL
OIm3F4wNUD10Bg4uw4itpOvdfB7xXbSJBKUhHNY5ro6gb9UuBI3GdWR7j9Usv/0I
M9lr6kXhHBDqXyKD0uiffIXe6vOokumvYNWGgf9kArT4eondcBBUouFvL4+CtYSq
44ZMld/uSs5WSAF6gBN+LWdg9c9VUcGCy829voqVCW6IVhgJsh9uvivFICrg9gXr
ERFDY9AMmOkzmdo6/hUF5FZCTiEtGf+QwDCgPYJJ1/u2S/g0qHZ9LMIepF3Uyix8
k9QsXUpQ38QsJkjxhXs707LfU8szjG1CmnHEpB/TwAccAcvq5yEdbIdaAvchMvKg
UCMenC8AFPX/Pow0f+WT+ZhiyweekDjjVTX8f16DiIaczsDWDbVZFnPHyWy1KcHY
r30a2mAZJX3D9PU2DQAYuhdY/2J4DMEejXezxQHnyiCAhOJrR6VhXIvaj3vcp9Zu
M+wXevHVkUb2BwHYMFkFXkf8NSwiLY6XD5SZdL+EqTEOfyzM3IZy8j0l46LYhBu5
+JirU6tqF1xByBhLbWSb36uiL8igLrkI5j32vh78fpQVwGnlKZfm8le/3Y8TwFrn
g6ofxgTocCt8CptRI9ZGQ6AkwrZAZ74lk6kas8CttCpA5dWxGFnY75Dcr1gwev2D
oWn50ATNFYlZPT0BnqtSfQfDwUvSnXBvJkqs3hXGdjRUxJJl7IZn1sHJGaNJaecp
Q1YB7XPEUs9+vV8sN4z3BPSsI+NNY9fFgG8Oi9tJkaCB9KNwz6UYqkUtiIer9YJP
Zy49lN2D5U6dDiIZEAMzr7UO3T/GtdHUtw1x5KXw+iy0k/zPCSNfuJ8JMNTivMht
zOB63cty9eSm7GhiKdJBufvFGkdZuUEwBeJJaIpoOqxSSQMEzzrdQGKnlETJ9y2g
YVXUr9Tp9LKKK5qnPiaxjizMn+ONP0coBK3FF04U+xEdpjLr7EFquv/asB3KrV30
IAYcFaMieqXy1bEYpzfebIg4e/RR+8tBtB3SK+OC38PjXxztPzksZWuNY8FDwRAH
BHfMTlsK0NPTnbGDDHhZxBZD0zP4MWPYVDvXka5MGCcxVVJ17U7F2r7O/R2TrxOt
KMoi0Hepw5SH0qOdnEgHxv9y4wy+iAfpy63fQNdw0wjTnrwByS0rQeXoCebrV683
vjewK5RpQhn+DGP6OHmO8HXM0tQ6q0SPa7hDmhVE3Rb4OxtqGn+AFB1OtDAFDQLM
eI17Ts4xOfgUIfHCnnGEjB2OcTH1/MAoSUGtYPvccz0RDl+OpwR0kis7PzvZQYUT
rkhGTlCDY3HaLXSbPIGp+DVXfZvQ3FgImxYIs/0/2Gd+d6mWLmnz1W4ZAh9670kP
xm7DL7gSpAaD1upDBTdDVvLzMxSVLSmNif6EoWatK2WpXP+NvcZtWCH+eUcb45cL
zB62xTHK+O1JvGbCz6M3ou3stgWodb0y5VORFFG7/bRkuJirRsoPZ5eA3SoKTFNw
NKG2fSosxl5/pYL9imObMf418ez+E7bmZ0NQBhC1B/PAdkE/wBU9pWSVzYCD7DnW
JLGc3qP13CnoOYpxNIs89CGpqSARS2EVkwA4Svur242iL8JFozxDGjTf1p0dmXsN
vMInQe3WV/kprThGOByWaeIsagNl8HT5j8XU5PzgXGsUqS31MG59DVXeq0RkbLxU
Wf2/OOa30riqf/uXq/HMe5ccfKSKVOL1Qm40uTZhMs802+X51OdIqeqrgLAAeYiy
qqL3UMZw/H0AruE7VPpK/BXMqSXUc3L2wFzDZoKmsnEwcS7lkefK6sW+YwT0yLjY
Cn+r+iQYKksuOG6tJ3Q+OfQhrGwwDmPJQzdFBhPDWCq5b5zFLeUDk+hQTwtV+ZfT
P2ebu8AEi8zXxsxs4ExHS3iSsHZ0gLRaDEv/aMRZC40tEA10em3JcVJm7eOOyn9V
QmMtgTFOMhv4kUw/4LE28efz5pTJxFs6H7hnrC2mSCpoKBrGMGHYLKeTL1cUDtsB
oqCGC0RLGq43Q3RR0ajZgrQ0YikvKZFpmV75LWuB4dOjrPbyInZGgpNKHMKlX3tR
tyYd9tvdH2vlit3dq8sgj+PjgZTJWJ1ERQG7n9qNj/EhbT59czDr5EX6alrESpxG
BwrnoRzU8J1sLgOF8e/eJ4DL0klh1PpDUl2UMw5k26p6JyDrHf0YPKKgvY8calzX
jZjraeTyLnoteMZpC6bVvbqOQ3Bn+HPtujvR/+9ZZm4leGIcnNJ7Z9VTXxTNhFuX
NkD23Aw1gA3d7teNmv4IEgJt4lDkDO3zN/8Kddpw0zSkvo1uAwrGCSnghETcU1ey
YsC68M8Mn7NerPAFoFLQl6jMZtr/Cv02Y6Nyrakwo9OA4Eb7hTPoVQfmJkvwCDp2
I+Gc3LlcCiEKVxR1eN+0rpPA4IYZj/qqKprtQCz6LtNGsZZXDwVOt7yWD3iuJyez
IBnOu5a0b11zv5wNbfh2QKde+OIg50S9MoZZZI54H7/5kTSAMDMQiTXIHTkCD+Oh
RnlGxAAdK8C1VDBg+TTDDLisN+MzHI7Gv40JCrilBfJINUQMf/1/j0IxIbpB9Mhw
2ghy/NJ2vzwTkgNmUKxPb04NA9Jaq17OxM8ao8PozBuXVXJBzWme/2yiaFLR6mft
YgBXgfJhett20Fcm+JZU5/7NZSX6EK10PwTk2rmFcnlo6z/f8w8XhQfQSXZgQy5F
2Ta1aIHjPX8xkKpDgcLbOwKHUymycFCpbwLVXubut7MNXJoZG4pEIKciq9n9mctT
zqu20G2grqlonbyJO9pcAIveARa4cyW6JJ/6PnGNMf2pcJxfR3xH9CEi1o73ni4w
fWYWdK3FmoUY/QYJLtaBJWqeuv/g7dRVSlcl8KJMRoifHIikIThHlZJeaouXp117
B6P1z1UTmCoQsDJJk/O3ucdIYQMSpcsELQ+K4zrAFeuLsk9gfAz3ogRLGuuNjrGH
ud90c6nYq10RkYdnuT6GCYdS6KD36qlbV+kpPTMgcEDhlsuHo55D5we4pYoTeeL8
JDbvVN2UfvePsFnLio3MZTiAzH7Z2KLEb8ZRCGv8c6ZmXySZnFFlN8qBvjdxkAeV
v9lvTkAgqjA3J4zEnfq/0mWhRIv52UQl/hABUgnlLaUVNfFshvpPXg98WCCYCFZs
vaC0MCKm3wfKJBkwN2VhDp0qBaKtaE0zybGIllpRXz4HTx1ym3C8nH/l2sf4z8yi
iihFSNfy37SG+Kpxzjq+VVS2WNUVtQUJip8Y/LR2jPtp6qOx+Lh5HEgihyki/fZm
0j/Wb6myLX0/t9vSZOGWD5R0IFguLuGG+6nwKxbBHq3IPVvihTfngD1vU/E3HlZ2
YhbxazI6RkqcLMTV9dARKhRQHa88FK1cmxeJ4W0DWwJhyA6jViyiiZhIwj1gAECu
Bm01s6/ZUgUjBTl33otry7kCsED8lAh+3WZDRtboNMv/6sjtGwkhngp+ApGapOoE
6KL35wil7Nvby2dQDe1+Zwk0cl3ZtJyjeXIf5b6yY+9CklCUWcmNgRc+HMDJI3d2
yXCgSSoba3mzMnuQlSk3e3pTudVO31wHF85+p8LHXsL6jGBTETTuUBq2eUrua8qG
0FhibtXEtBJFYLrDIJi5TL9I4DEaH3CMLAs8rA0zTvZjFvZ/vL+pKySIeZ1+CccU
a4RJm8/Tf75FS+kbXnan8CXFiV+hG1ugqgjNrm5kBssKOZxZT8uPo1V7q/n+wNDz
ELdHbk0yiOQSDlHF7ZmjWI0hik6jzGoUiOtBfiCof2dvN65AwtDF/pOS0KXqVuPI
x2BKnQpUw+ojs2RiaQmXeWwFzIUuKoIFtsvdLIid49uhW4ghTQdmifPIYt4BcLU4
q/u6gJFkRHRu7C89MHJZRAxq/uEI8tpqBpbPSEdrzfiKf3Htv+w6wzQc+dDim+dE
RIOUj9VfPWvmM2CCu4bkkQ3bpJUOFZ2/Scr/QjfteexrEiFlsnKBhpV01kPM0Gav
pw1innIjsKxdTrZCsnIph9FQLQeYgrUJZdWE8kvmxfwrfMmQyEnwkFKWppSRY/t6
8qhfovgUkspYclOW1L3LpHLFwu+D/Wu79skHKB0ljgm5e5a0LAkvhMt5uKiCQWqv
COv+SOfDJXoOalgFbz1evqJv45fXUTENqNJyrMh5oiJGtDBtS5Ex8qbIEuRdhxeC
8GLKY/XJKTPAihhhpSzlR2yd9U30/n4BNz6hXIPFcJH3qB5sIaVDE/0oFPoAPzfn
lrOR19HtW75xip+rfCDhDK2M0QoZXIIX1gfZbnQsyoOzk3ZSG/4hTwfnkfdfriPC
zV/JmJc7uNAHdZ1Zvpi1KpPVZe1kXoHzX2eJFW0en0uOupoALcssphck8DLTcWen
3Bi2g2JC7tpwX+YpIbxUiL+Qt+NdzhsmUxIJU8GC13na4deFB3uVYC7zSgV21UBw
RA/Ioq0zQiY1tNFLd2jf1bmajsLc1DndsKHFN4W/iLx+3alqRsfcr0tVklznGApE
aEP7gvxTQO5CfvKE9Wh6fA/AYt+HenkutjwhliYtAHK1ljJPE2r066c/jIQQ2Hbo
ALm3XqOp9qJ6cG7t2WbEtKJUqOxAuelKkI0Je9gcSHpkud2gDOsqGy2vuGv338ht
S3/8COj5nq69ml0eYw1FTs41hhdlLgXZFYClKsuMvY2S1zXTB6fQkJ/vAFwLPaLv
l+lwCY27M5jQG+zcO5u0daDAS+jlUv6VKp5pJg4JufxfudkO6x9uLWE16HRIqAKp
dtTXIinwhenccjz4yDgrkU06my+ArsNjzf8Letrq4khsQg127SXsAiAtA3Kxyx9c
8Nurx2quvc5ZETMpPe1A4Qe/1wwue5JW3bq3dlONSXwZ90sw/O0neqVSgRljvYd+
hdQfcgETqeVnhp5xGPAjVQYRSwYOQYUv/KJh23vykSUb60ZSnRoCMKy5S4RzmqkU
cfuYatuZDI5CpoWZzp5B3z6CU8e/jwz2prwMhTP0ErrsenQeE9l5wgtvIiNOcdNa
tcSDwkmMM1rJDe/FrruRt8y1suYtn9EM/+ikEaKsZ8qFiIgKX4w2vmwecPiG4zGR
tALGpKJNwVJqDDxU2avSwNXtFSkJEG4mYnkYAsLT4wFNUoswFJB2KcIHn8EROB87
yOUBJB4MThmJ1aCZZiPXokpr9GS2S3SJOcmiMexurq9qEg21hdEKOUCjyAKwUgf7
RPvELbrPPUdQ47Z+DpzUup+wQnrx8IcxtnFRiVjtPWwwF08+SJWzTt3k5sBEWjnX
DeYA3nVu8ZBNNqBNsXS3oLWzONo558ISHh6qA2neda/K8LQEl5e0R41Bbk0PZqTe
VorLe6+xZN07Nc5gex08OpCrivhDxpJeaO8a5smG3GklH4C71p5PtUzBebsO5CfH
cPPW4YIGUxUC+9e+4XegR2yqkbCFh/w7+No6N+ph+UIv+9pn008xcY7j4f3pttN9
eWQblerxkIAo1UN1FYZIvT9ZjhEckvq2RjS/OpFpvj4CRJ5AuFl0/duYoYIqY6gt
0ZfL98K1cEflG+VfnyM81YI990PV95RjVCutmNz+L5WCOdjHpUV/2pFedRIJrEd1
8Wl2c4xfoEMi4VbR0dozc+RnQZqA5GvLqpFVudgxVpAso/pLUL1VWWiHTBr9XNuF
pWavr4Ba0emxgSL2d3xSbp2uP7DXg53PUXsW5Qd1ay9920TNQfl3lH76fjSRq0o1
x+qtKdKsr6t/+oY78dnDCKbxKgcDZZIvEv6m3ZF9CkYzsHSYSQt4SGzhuLiwKNcD
miFgmIS5kkucmuEWKN3L1EdKoepfbdagXvXrO9YgrbwlzqDp9vU14CY5u/uM+klC
A+++Gbxv9I5CQ+uCwN81ee/vXe4zuq9i3K21bxAF6162jcAJp3epAIbrnCL8qL5s
m7ZeSnXxQPvl9dtuf7YOFZa06napf2D3c+YbD7AvuCR68Sw0axGSN14AA/n7yRnD
unW9qyirAsLOfzELkcfWKt6SPl0Y4fxlDLKtce3pBK1qd/Chjd1f3V9zMIm0Uday
vCzE1Wgg3gpxb/C50AWoOD0TZH1OMLdZdlAiE3H3Y5c+k2TiyX6cAi21RjSEmKnI
UvYxV6Xsq5KAU6d6oiGhsjGAkrDD8IhxiDSOdpt4+8BaAsTlNgAfRRgCrOnr6J1B
0uGghB0H6q1cO3z6IZedCdxMzWxoLU/DvzEs2yi9iifxITRU28C0nMZL1n5YpSSB
qe96OvXV+6bzqjEKchY6HReI4TOwngaU4M3HEqSJVObuDlGb5uFskYHfB7Bjhj7h
p20SGK3bGofzKymzXk5y71PGkepBes/R/CrwoPtohfNlHbBuHBILKgG78OouQrdz
bYodMqD4iH23NrRp9tKL7NHWVHJ4Mpm6DA4kX5HHWh9GSWSBP0jU+UM6UCktNxN1
0nQj5C4iR+35KGdNW9tZA1pJ/cacRTuovH2h+jTb3a+P/XDPcZm2D4B9ViMR1SbD
FLxD5AIeJRTwLQ7BEC8L0U7v7wHPlbaixfP/Ipok12Ss/xJbrUiOd6RgD8PoksfF
WuomswToiJCAN78OgiY6r5eL90jt89hQ4wTKK1egDLwgD2EfktdnjXmaW/gA4h/Q
Kb9zvfZ8Hkqo5TPipjMDUqtL1CQVSPUR3sEsuMPuZ1/v/KdArrYCAd0sL5YZEvxb
rng4lpzDe/ETqgKeHJf3JEoeV2SFid8+p3D0JD1d3IMzduAWwXcS7PCnr8Ax4hqy
xFbaBhisJ6aYuSK0bINd7wYgAKk/vPUrsbb5oV5QXuHSwfJ4Lmm8045Ld/C0mnTe
28atVTv5/BrwVTmSKMhik8BWFGMqvyg2Dv3I6wbM6pwIAXTBSThglcRrEw2rs8th
/aC1eghfwLkslsWvvuRyXPgu8BFeCUG+LYxzzuM3RYF00XLsItO/AtkUHTIbuO6W
S3Qaaga7xb6bZDRiQIP3yt3mSz5LyRY9Tkvn1FH8G8PnCndSyZJTixsGrE2FRUCv
td9zncm7x/dWbDw+w5n0KoTONT7Prgkq9GdC+cSbHKN9z7/wtUCnO5Guk+eawK0I
lr88KMMJWHigJVo68HI1tZGX1kRPyHBaRyEhC8qKDEA1mcHCGOcowmswk9IpMwNB
C8ZNDpR9/rqXKHh5PgneN/zPrCWW/RTpu+Of4TCJ/RZ0+v7DYRUgv8vl3/zmba3K
uBgZKNOU9LHu7PAQU68dXvDXyRDV1WBW/KsIRF73D5vcT9nyZNRSr5U5U5H1LHen
BbU5s+iQV/yFT5Wh4tMXC4xwIX1BVsNjZCNY/HAbhc5U6/cT/pqFk5rkALadGtvL
4yf5GLpC5OhlLKze8gQAclUq6Xfjp9AocpG34xmwD5z/cdWNPEhNuldqbQyKIOzO
36Ofq64X7q+z1EjLNrbdGdOwcq62FhxqYHsuM2sRknUybHIBqMenSJa6jN0JQpHO
HIYd8ipTtGfbc5i3zxXxmPUUqDWNR4GyljOsyy214B3w4B49P2GJRyMfUQ4YgymD
4T89gevyrOgCgIf441bTj2Yg59sCWkznjjYsKi+cJrVcEUhsI8YqcUC8+B55N+3G
u/lms5tewLxNbMv/OGZNJ5FXk8neZE4NgBZl1MyqRup0nIMrnkm2CJTklIh2myhE
UFfS6Q8Kxtd3hDFxitzVRbnD4UBEo85p1cejfeZpvrW60HSRVpic07ukxO2Al//2
t/o+plgwx97URs+9721dhkpLX0Ay7cit1fINr8yV9xLAe5+MLNGHSxw0W0ygViwe
PTbEjyhBJoaEcY0vRD+p/eHVAM47N3ZMlKZfA59/0Jx3rp/gbfNIJsd6bjSlDlmJ
ia5p99ENxc89jgv8+rj9mFn9k1Kj2Jl6uid21rBlXfvksJ3o6n9YyFZo87uIfv/O
FP8sskwwR4TPAwQW0ir/tWEZoLRVLONhYpBMUuougtZUJnOrdrw+XuXpaAUHyMJy
pkthYi9TYZxIM+4/gaMF2VNDzXyMU0zJJ0wazhLz/0NWbV9U+gfCRxZBrQlq15OW
2aiUKUaguOdnjaf/LLP4EatJMziiZNGetOWQqZIuDYSyWi5KsftbtJ4RZ/6wcJny
HI+MnWHdBYqp/Z7pJzZ6SCcJhEIphXpzfDQ86REFIrFdJ+5lpqvHbH9HqCoF2QbG
TM/o1Wk45YgR85vlXyj+aUmasvNV5Bc9nt4InfiLpvoZcMXH3vWLnpQpa1Lo5QgA
Bkn84+I2qTFlfW9RfOROccAuSDHmYQ9Qz7DHEpzdNBDRUCMbO7Dkx0JYP+MM8uYY
wNDysw2tvfULd/0yYUVrYGfTHpP5nKf2EYUc4fZy9cVwn2vWC50OspYvpRIP8S+T
AF3cE8A1CfnSE+v1htexo9l77ArhVaGK5j4ztibfzoryYpt5AnuBWCYayC2BatDw
GdLoLbpeS3PqHrcdQjF6Tb0/3Ce+8GA8Ax5itK0AbBWMxeBBk+hH804tKmiLUwPh
5jREM8YTMwkg4ao5X/26VWdfqfzeYhY1cl+V8rR5akyt3hab7IzyjQRhN0l6TN6s
StN2lmutzhsYk2W52jDtfkD4rJhNl2jP685NDlxVO36xzc5xLso7knlqT3vS1Cw4
45A8RF2OTv/dl/pYKMR4wMPNj531sC3NB6TN3D7eEHEyiH7DkScfBod+ZJFlzyYE
MtWmbEaWH3FM/oYp3So9nRIgYbeP4tw7z9BwC054g4TRbB6nJxm8hmOrE38jF9Y4
gxwNTru9W5FSW0uYphwywmDRkola4jaLfxxlzo+LZL2KSDqA1TkuHvbpPgSiZWqH
+LTBiwWEPvBO5E7b1APhr8HF3CFmjN/rOlAzFPuRfu3Vcpzi6302YRxWTeKUcmeW
RIi+gmLy/Q8kzO5aCShlKNmfDFIX1b1TB/F+O+zrskFcm0nFXFPzEJ3UtmRVCfVb
BtB1QkFHqh4Qlgmt1nLXN4mHfwk0TVtMfuIobxvwlKom78VL+Ji3jBzIsNjwPrPm
nnkBVXTnqvu4NjwBJdpq95m7hkk7ey1G1kC15Xq9PkrmA0lQdCV6nyExEMqwxfLY
OR40elR48lYR3eaw+jagMvVX86lOhJsH7gV5K+UgRpcuilAsVhFTYjA2/Mp/+oaK
UNAnjLu5QsQ+I5uWKmM43qAhnLe25D8IoxtkN+AazBQI+CzDdbR12QUlYvLcDUzd
pvglvOy2vpKGD5Mej94Ge9dRiTnmnG1Fk/vSYkWmIrEjy67ENn7FEflDntZn8sYC
WjmK/ZBjtavYRtbEV9kL3UM46Qvqrzk8nlG/jC3SRKunTHB2sEPKhT/kaPnH8a7Q
P1Yo1MUOcH2NkiM8KjGl1HxVtbsyt7u7PW+Y+YE5mpAyl38eOt1ziHoolCve+nq/
eEj1iwv0s0Ov8FWS5xs1myXJEuof5K/CGSZCzTN6pX3urJzDlGBd4zsmzE3iUoHo
OcXRLR3YatGPAKlUFY+5AyoCXkVAwMml4ixiWQvCcnOJhNCNfosnHDXBfmv656qT
Wxb+VjTDZgKIkmlrjhDItVRWDKhfM6cltNwA+I+Gd8/j4nenkX0jif6VxqV+2H+4
X10KBzECWTrAB9r5KtuBWzOIh4+GqkHdgTXzy9MqWWY01DrnahrcG2McSM5jTOFf
0IGhe+XRrGxGlQ/awQgBbdBDaam4z8VeRBFWZ4HprfafTeteS3UL2IdnN1fa55gO
iDiiV5Dy0gGSvzvfQCGKdQZI+nrOOIlDQwwEv7cYqBv9Q04vaSoluX6NK1bAkrM2
222wrSs1DKcyTfthnlk9VkWgFofh2de1jiA0ciMeKhPUrI6NPIGDHElG5XkRogzx
X5n9E6EHpC9nd4TS3W2Z7xTo1GQ/B+aArv+Eu+ij8EYjJ/g2QF58jPRmSMePma4s
c1/mraZSumTUTFIGuPm54449xHGOvR3QZ9YfJ25e0Tfz6v5atQsAtsti/NCg6h8/
sL8NDvIuiEV7Y4T1mP1hRVhgCBb738xM7DkHEGRjiq3T5UndG1J7MMCofuD8QZFO
WheN1CDL9wuG3ZiT3WN8RkoKjZ6ex7Fz9Jl/8MfFW0l8GqNiX5I9ByUXogOy/xra
khnmoI3UZEndZOGmjvu38Godf8cUAQofy0N3rDs97DTvvdMr/ew5v79TERmXYe2f
a8EcUoh4NKSaQhnfmEMYAsuspWZjyLNNWTjB3d5kMkkRQmb6O9zBP+HQh1lwTVDk
NelIrGAH1Lepwa4l/9msnOI70kauwLYN7kuQrH9qm8WmnxlSeYQA8b2WiV77e4Le
zrQjLjhhKecbgrUYySGOmhymZoPYwFHaEWikwYqBVK8KcIpaeMo0VgIbuufT5L++
GKZGAIW3a3o28QnwaCDh90Ox4/Wa5jEW9SL3M+8/tVBVGaGO5UTaxFq1sd6zA5QP
rl/Ejr15aetDW1pJLVOB6j4DHrd8DwnrhllUQIOgjfHzNnupxP2kXdxLHeTJQdWn
r+yP0iRqh7N/rs4wnmP643twg/Ej8V/lkJJ4u2IPYgwgBglkPazdDIOm90tfIj5f
juO7xvqt2f+A1lQXA48/CK+lSYM1gChCFaE4aOQVM6hlxGT36sNUFjKL6kzA3uhc
tSfIDZnW9TEnxUHWC3S9wuloe+wmQE++bV7Doz45Rn9pQ8K1p83ovhAfc07iWw9A
ie1vBVPoyoFSXTQQrMlTrjXx+cBUgo0Z4hcQBak241c1Sj6aZbV1/EoaJBtgPVe9
7bSXib0iIw43AniGqByNfTLUKjmLpQmo7Okpt3NMIazYTteim8jP+QhN9BLQMomp
HxG5J0BnSlEMhwPFaFim6Wv1k62oIPIc1ISzm+7Nn3RkAjfq6xP+Kc039aZCV3R+
sctaZirsRL705A6W3QXUq0Bv3DQL/jsAvqfKcFTKF3gmeNSNjk2dOR37CLmWK8uk
MmcrQj2PdJcxYUQGgZTlvRnvCUJpSZYSWAKGm/zy7KYqsYkGQuh1iwO/ZGQBuU0p
YgCrvbgKl2kFPmZ/rX+FWFJ4Qgq6D6nsa7WCSPpRFhQo6YWMZGW0X8Ub46AUs2zr
Le40eLkcNy2rjiO+1Y/Z2cv56fulFDBTvzDOXZzJeWZWqdAZrLmKfiRLoJK9BmjW
rK2reKr0owSr0lutfL0SB03YQSs+/CpIsDpObPClcof1PPPP6rMudpNUuylv306I
ZGMAKfZMK7+MKtbVhNvLPcBBVeY50/HoKKcnoWbbYb7gDBoA6Azzy87Dys6JxQGv
tZYyOMyi5/6Rl5U6BWWs7KQDuoOfND7lAtMxbiWr8TjiR6mWp7ijf+ml5+JUjitG
OXL42buV9qYGd31X13jrzbvxazlyWiAKn026W8yo+SGeSXmx2nvXWRy0+0Uky5bW
e35QkDhGmF0gKy1s4mjG2UdODbD8llZtI+NUE2kECSQOGGU6XgkqoJ3/W4WSiDA+
CAeBN6q8gbH9ErwMW2pBrwA15ejIqIGgKIUMArZLCdZ4F+hJEmSX4SV8xr8Fmuo1
/P6APO3BSswTeypdQ7SII4zDrM7/M7nnGPlTAwqTjkGsfjWntsVefr9pucnYkdSf
RRhwg6tBYBVrPw38O+K5ve3FHH3DcYcq9qCDfjARwZIz7vRfN/MmlX8sMd5cfOy9
QrkYt31HcTNgvZ/DoAtaH7PQ1BTn2YmNdCStZZQ+k3yOGbj/35zWPt9cafaNmB1w
fKD56VBL8INouZXwQWbdiViiYZamDtZScjr47TsvEyr6Ua+zv94zTgy/z7ddzqge
jBiBs2eRfMp34Pe1zoteeg5EMlKaUkzmQSYgso3ImQBJBHR8StsGlBBWbR5BP7JS
dV2B1qosec4CRiLqzBJOow6Dlrny0pY3fj66lnzAKof9Ouc+mrIfRQxmBgxdpWyY
34wScMkAR/d6Ooze9/ULFColgZZjMcMcAbPuw8bem/1Uu75/xe5iASGr6XRBZTs4
WBydGsoNlKIu0+gCEVg/octDA2vnsKVdEzkxXpBqv6rB4GUe9iNa5uoD2xp3H+ny
GiekCkC/AlHgwYi5aFq7Vm9X75vZdiYGehp9jtA4TBu4l+UVgocPnvs7zfXwFUkY
rax5w8f1ZnPPjqi1h5QDzOukR08YBjyCgF7tk1SuOQrdpUGI2Y1FBrUdVXU1JDEx
GJX+dAiAZ6l2T3SKI5fxUJaeYMaGVPdg5SrkhMS1bzUGeY+y7W1QSXJ4jjUy9Ent
/JMEv63pRA80FgUPue9jZjjYWmJkcQ6KF2Drooa7nSTPeoXD05pb0nsk9vT1ikfl
TE3bh0DUHUdvfa8boRcmQPl6eipmPGvNhydLyQXZmmnOnBGJYmopHEL6gJu8MRAZ
FDX87gz8RDypBU9z879GeSCoTsrRp4mBbsvCgsfNGNMInZcgpO+jDp0FKC2VX3Qd
fJKl+jiy2naRsrJH8BJOMcde1hXIOA9t45NQqKbzRACv+c7Wupt0Gv9Hkc1qlQxp
SsK+9S4ckKSdDZhEwDJEBnzninLOg3JHeD3fJAEQKpCbdJoib/W1tmn0HRUCTddz
ThUTpmQmn/V++xr+A8jVqRPGzfnZz4GOlRmEx2EB4ZtZYYO/ulpV6+HqWykHYbmz
hqNHheyutL+utQt0HoctbutLrDNxzGJCqknzSnJZXelWqm2xC5DS5UGQSU+3fpl8
KiXJSu0PHba9/ea8XsNSl8uh2hn9Ws+Fi1pI7wiXgspJ9/EZr4S76BpXMR/BO13o
zKIanGRvPcS7TDzR0u1DrJVrK7+mPLSgWfFXQ3LK44N7rJVpK/lMq2nNghAt5BHt
Tw91VF5wjB0x5t/s+FPb/aslBz6bc+R5syzZetRDWHkcyXKSQRi8emNvU8obuODq
Bp+fyfkrtCtPvEWTYc0qNEgS6ey6n8otqGr4vSWL1fHtcDtQOl7YBRlqIItkNV7E
NCkBS26AlaZpau43iPjQ7exZlwafm+JKDhAiIHsK/yYVAT1rPk4/HXgo2md1J03n
nmFPCOMMiybu2tN9Sycd/m/yHLf3Ztcfbbg2+J3lMvrRYaVlErJ30HtAdh9+9Gwu
qbFIdyrubh5Dg7b9w6iWSRD1Qf3MMzmd1Sn+d8+f2AY0T4YrtRnJo3enheuYRWnK
m02Sb+tD9l9MsGZogUTU44WT1/bnKjB5T3ENm2SpJrN95+LXB6VhFKpBA061iKQY
xTi1053EyTVfSBWuA8sYL9AhDv1RewlGRYjdYDuFeVlA621TrCV8FIMsJVQ5cO++
MghZV9RUCDEHuP3ZxdsaeS98nG3guGTxH47kqmc7fJVZsp/irjF1mAVij6eec9rU
yZPog2D85VTzDz7ustfGzCUqUfW3z6TOMRh38KEzTaMmhETCRManGlSNk3fnLdQx
r2Lp8Z2DhX2iCKBLDFm40hnecMtkMMEvmWeQjQejsNoqiTxa2Obm2qzJIoJG77j9
u9Dd9tnUsGz/tfWl3+O6/i3PLNj6zptsxMbiw2BVCISvhMUg5orLEybDjVQyj/+r
YXS60x7E8zFOXAtPwiml1Gy4BlTRaDkjtaeEsAkFRsXjXfxpy5SPs/dSEPrW5P2Q
52Huqo3D9OCwodJsZ3KZLxNikrJRvkYSehY/u2/8zo0P6IcakyRchnRCFeaeHx7J
oJrijoaOaB1QxeI1eSKMXL6RSZmTCDGGa7TI3YtI1/oQlyQ8DPVcZO7fVeUAuncD
/wvxAJJIf5GsJXjh/+nAj1go0VAg8I+X85cxu/tU9G7tjTmmFeIVTXo1ijo+3O8L
uLWL62vPZCQJMU+kHddHDGclJbVhOjvQu3707FfcuoaOweWPDw90BuNAQ4KMn4fN
gewO/NLnrH4VpwXNZKPO9rU6Zf8FLzSM6XZL3wK0q63WV2wMC/En6MjstPyoJK1Y
H5lRdcBhMGU2U6BzQxbhJc/sK3doBS+fkzKtjYWIBRlXFE5nfeA8j+NipSTwL3jD
oVQJ5g0UBW9S10yU58y+Fa0fRBIGJJuSGjKq5ibuCoCTs3D5MTsKfPNB4Ix+xJKx
jP/fV6YDQ/9rxKQISzmXgoScAefkoFMGZOureJHug5521cAPHsFRwdp8eWEseG7E
wr4eNY0klaEqrRsmTPvx6tnFCi7xZb4TEeiVBxbopeiacOl0YNtP3XnURmjHSNTs
9dc9q/KqeQVvBErmC0ImZ+Z1l+MtD0XTQZK+FSXWrblBpIN4t6nqqJJ+2vw8+OlW
wvzZSUW6yumMGVQ5RGje9Hd4w56GqDhmiboF1HLdn9Qf392YALKTlAweEvSYBYAp
Z/lRjTQkfgd4h34G78xyjQg22xex3NZM3HxCT378xfCwoFBccM9uwg3S1HKQv2s0
iKFWP4HGUd32iTRaj1zc0MMidY+0+k5HBKkXiu+e2X1IOpl0db7Vm6qmNP2okXdF
dC82rJfwlDVr8hYe5khK8IDrJjFr39WWcURgHahl8L6KGI63OMJVM4xxx/a+nNeO
2fq0QeYS5zZ3Ok8XtzNZeG3G3woq/qUR3KKndUbt7iBp2kkyX8xYyq5t8mvrjNjK
I/Dd34qShSNyvLtY/ASddsPgsaqNM4lYbWfhNkvMzA/aTYfZIZ1gCN/hGwKNepZ8
IQAvlQWYZiTxDAehgeQTQIV311Vr9VWYf0QucT1Zc8LLtaEFzlO3+jHUm9wk8DII
ieyhl+6GRXWdA0x3p6NOqZNi0TzvXvQZaSueZr1ctKUbGeiS1Svi3NQ9kFrTiF5V
jH2y65LFOjgyRkJ2s7zuyPHQPU66Y6LEbD9M0gKBdhDVmOSzsTyDC1UJITY6vuJf
z6FxEawx1m984i+Rx1Qhf3TFscaMj/UJIBf0mWn02JzQeXzyUwXMAfKk01Odf4yR
beEIvlD2mT3xl5V5aVy8xutopKYQgT476nDbBKfo6sDsgRKPW3pYQzGOZuPGwaKZ
a+Fc4nY9b47CxNtLJ//luNUY9Jya/ukaDKUdhWtoaZF3ojF/YahPOL+/JZ9asijD
PatgHkWQEZI+sGLPnJ966KQ/MAe16PaX/IIQQLNfgJoJljbQf0PpxNEJHgw8LdI1
0lkChk1ml97PkpQ4zDylWkSkf5pkuXjDdkhqLkmh8hnoSNyYeuR/fDKdubZ+NOg7
Bn/IjeQy9jslwPIRYRF+rnSZw8m75jUhkmmAY1b73yqfY17yhaL+b5JUQ8bd7nPl
/E5Om9pNTIazH08aV/DbECBBjkorgoUHLfuhURXSw+PrGQu+PkjdNB+2da971pKQ
E+2uMdLp8dzeMtnMSrcYt9IFLBWQYbt0Q/mLK35Rb0Nl313c746r/DkIvXHuPgBB
HaGI/EQjP0QfnNl7hZzKXwpfzv7xLNylYELov75BLa12iUh2DMcFlq4Im/A2BONX
IiOZqM3uvqIs0vkBW3Ts6vEDOiWX70YiTv+pazLR7PaPAI/PMZDDYDz/xKiB+CsB
vCFhNBJ1hK6doHofngwNQfrY0vMYguDDUx60eG53JtVcTkikDXhpfKxUBKIBd5yE
cPKV7b3+DkkbZ5O60ZWLL8aIAX3epmTG+b1N54MsJD5HZHM86FPq65S3upL0aWPh
GA8TNeIkEv2JctbVDl+/qq6JIGxbcXcJoNeXWlI8761GdLIT0k39Ev7tS/gTuTMq
17j4tP4IfXDyu2U2ZLckIKKPdgcm+CUeQLLOtUiQo1Qu9LiFZD1Ub0DxhOWRtSiS
Z5H+L+oWMjjopa50vpB1WMXh802jFHLC0XtDsIm/Knfhl/FKlLdCFpTktj19pp9U
73nv1ZjL/QVg48hIYP2Ygk1bw4FRmn2JNw0hsmIJzYGkpROJxoZnwL3qZ8D2ZaBe
dd/3UQK88NGQ2p/n1lN1vpOUAmdC9nKzN5K4oxqrgSqfsfJNmucJKVUQqYPHUFrA
xylDJOQoPkv9rHys8ekF4cicRGxO6T5h5J436w7SAghyYIlT284F8fXJ0fyNKwvV
ST/iLRFkszMZ8AJLWoAt0eiji5SAc3oDfellZvZCAsbNBciH9ks64yB6As9fMCyl
LkS7m8I91rmMhgPpjDJ5t87z1Aop3NFe7BdWoBADM9bS1O6jRAJ8pX/mJkF/Xol1
JqkLlP3TPQ/Rfv6Xmr+eUhSXRO9nQqjBddXiml65NBoPBh/8cuLNbsraRfVLh7Xw
VDl9OOpHfMP42//tJOCBqDNhJrKte5CgF4LCROet3CEPrBJQ14IN24nHCuhPLOPl
CBkdAaSc9xKACpeAfQV/aJQ0WjZa/okZrctv5Wea3Fgp6eFPQXWA9PpNtOafdQLw
5SGvK+5UXZPU48D4Y88CkqAYefEQXjk4++IXKS6viFVSBP5h7pkIFH+VYPGlyNeu
UuFx9MMGnKd11huB4Sh59Sg/u+0b3/PufqruWKzwd3pNWh9upZBS2cnpfg2jyEiB
GxpuanHyT7kdwqjbYTRU3cOMZ2nF9+8UwhZPw1FVUWz9HDVIygytaggfutCJiPcs
B2B2CXVmY0r0KGqSom8oqga+yuxTNxVX6ZhxZLOTp/aPMStNjs7hB+JaUYfIrtP2
dV6e0n3rnVeylxYDXaO64Ps5MBi3aQDt3Fgr2MWv7X4QYhZqM/7SwzT9dXXEXZHE
9v2NvuzjpPk28LK4zGCdzE51AtxK606PLr3OG0Vrp17YiU8wf/XyMKo3u2DMFCBc
X5/GKXXnO74/AUgiwqSUw6Gd1n/FnuZo2HtxfmKYpWvjK+k3x3dLxqIPbmwhOlLP
naRG98DGWgPUj/9AsvVObyr6F4NyPGN/peyxc0wV7EnJM/8JkWAir2MnE73JyQ6Y
rlAHpnSPud1KG9CE5F5+hUXH+W+eRA7P9Yzq1ypR/bbjL3Gwzps5gZko2TH9Gbce
AEhN7m7vRngFvZ40WbqcqFOOTKU26F9k6ni0zuEK9HIsRD3+tiOdg48pQU4tE2iY
nU3AptGuV7L7iIdW+6G4rfoBdLx3mLZlwSOyf7Ma/rlXgG6J3snob8oPDVCsRRnK
Cl3gVtkOOK62GB9fIZEVaae/Yx3389nsLS2f084TfSEEJPNdAnnn6HnZ7yDX+keT
ffCgvUUu+I9KomBwCMjTO7E8L/Wmpji5JfHlyRPgRHutmrrkFpuxn7i07rPQxnEk
Ufoqc/k7HhJhlPIiYic7M1OEf5wAC6x60Bh3S8OMmUJcFZtbxLRdIosNV7rbgk+7
Qz2Y9TzH6S9f91edBs7ZB6kk5lDG9nWbhWQ2pl0GIEHC4OPDC71GZyXSPNwWLUao
tVRfnTdMN/bZa6CqTfXdSYNIxwKgp3g4wbei2bCk3R2pw9oDLPXpB3jwFuzl0z3L
A4dtzHPsDOlRbdWyYsUk3+/Rysy+qD7IDHTsDydBSzMGg0KpjNvf2fQ9xHMIEsUX
ZOgBfR3z9ITYEvEbce2z2PmDVKEyIWQIS/HrEZw5f9huCEqk4UZQp3zi2D8GpCh9
+hvTH6HczV4HZxkZ/OJNx/eEaj/X9AJUyF2bWlP5LzsXG5vq/9zEyXFJ2anew0DD
KW6IE1EX/DziT/mruSAprsezi75u2Y1+8jZ/m38bcBr7Ijfm171WvsiNY6wvVjWe
iq7w4R4RgGRvEgd2qZCv51V9CTf3vO3umNFPcRxGuPmzzORdpWH7RYg+C5wZqMvF
+BKKLVm2Wu+aJ6q3a+PqcADtITMK6g3ACM1pdA0zmNn85zyF7+AU/C6yHdFJmuT5
R+/rw3vOfsYfn9QlAAN0h5fEF0oiAceHzuM+yN0CeEmC5vV76IeSMXPtGf/XEDYj
8WURfqW2SL1TYc1o/QWXRgRf+2TQ1/vxkKoEcV2o4M8+flKNCOiqVOpKUe4aZGyT
IXuTmG4YdumS8dPaUp2Q1DEiRdn437i1aLVNQbn3i170Q+UmauLONqEqBkvc9L0K
VNiN1hFeW23jeL/mvpczYqjVOZ9UoKx1aMfjaw1UvWXHY2nt7s3K3TinCiENIIho
qnHw6hzCdvZRuby1ga+eZgc69oDVkY1rXYqZpt2J31MxXdf2nRk8zF7F72pAjVhT
i8ykpXWTwpqdQ3VqFJeBnEqGnpywiN/iE22vasySVddkMbWsrm4eegkN1ly5LD0B
TMlY1WYhXSiqwDAeZzZldeyhG86vq5OIMZZb/uZrSqnrBKuDfMEt2itkHDm3WVQ6
TO508eyy9auJZM7OW36+VS15X/bN1+Ae9XQGjzfM6TdKcypBqrnLWOGMnzOdeut3
VRveGkNpIcnNOorlXi0Rv677abL7MRM0J5ipTpg8Od9bt3dmJTs+p3LbTrNhk6tj
GopV9mrTKAXSbwcrh3oekRFxi6SnC5jFU8eDH4BH6C8kmIAtXIPxnjtKkJx0+++i
hWWeKIhKBgwHXzV2VneSmTDUNbQ7KtwVx/60nl7+RMsq6Q1/2Y/Ofir9EVJLz/VX
RBX9JKTjJMMm/NjhKiKum/lJQo3411tWy3pdPOpIcnsZ75jswUUPn8pq5cfEo6PN
mXGCDIcHLH7x4gxhzAOHT0MVcVFbXTgadpoTTbcIDjmlvHSqw7oMUl/YObvag744
OKkpBm8cwQTPa0xNw0ilgvb6PwUuYM5LnWZ8OrjXHNwaq+x6tM1y5hTY9s0GVLHv
K6fioEcVFB9XVsbe53UKKCaC4gKLpL1JkcPf3AgIEQoYsePj+w58O8WwyJbFamyW
cMhhxKT7V3M5c2PT8Xn7o73WaYvk5X/NM1FCXEqaKzPlk02/6+7llEcxNaKVEOZ4
3AcC/I64QTuDfoM2ev3TQKpyrG7lCGMBulbweLQWgLWqcCHQkaXZS+jS84q6AT51
TFEuuXvn1mmbRbmn7boLxygevVbaQlkPJv8ya4BATwRzowP/gcIjF6Rg8VmFzYB9
ubBASUkdyAGkhEQvsqHruHkwGTjWiNBIITJOin2Nn6zZcP+3Mr8XDRhZ4QYR29gx
+6vyB5rHs50ryNP5RmZYEXdO8R7H/2MWK6XTVuOpK2b+Vo2OT0v4GCeX0UzqtAla
N+PzBv2xs9cjTLlvJ+ofdh9+v+Rbwjy6z4mc9fCAEVw2Eg+7L6tuVwXjtvfkRlE6
f4GVdrtcTaOHw7Bayi1n5cBcPNOUl/+vwAdZz1MoOof02UU2eSF0FcdQ4ko9OFRO
vjVrXE9vWE+xrpzwjszeHlbkPNrRtNmZXzS3aU8IFAMHGo8865/WDWqNMfSzhWny
QD5SsrkF7t8EZxCmkjKY6VqmC9lLGAeIT90GxqrPsz47o2xGtCZHtPxNqVX44oNi
tNXK8sxgOseCNkG59yqLLE4b1Do7bbchJMO0u4bXdZhpYHfPHqRGsjaKGlI6yuC4
Ka57Sm5SU5t/q6wqAr0W6LUvxBnIp+luil6E8KAblmEwA4rJiqQsJNs7jNZP1l0A
dLHOI/DRNgG+/r9Oh9FfBbqJ+7+5HiqnPpqji+183HG0ub5NZqmT5oZ4XVTwqSSr
VG8OqXgTwNlxNp7X9rU6lSgiMb6wG3KR1ltPnobeJ1vQWmhpP0guux1wd/As4spy
6YP3R44WP8a2Qoj8lxAZDo28E9QCHYNIgM+sCNNPkOGds44OX/dmfvNWpJ18S3Hy
jNk8MbPeT9G759+VEZMFM2hO9QDL6+EH6x40880+RZIpkpHOjmsAxdSH0Fg9716w
gCU06xmDG5S0iN2jNt45fZwENGklsYGmoOh95M6FOCrUBC8Hxf4aQ6wjpxf5+qXv
5biaEt8SzHahrfsEaJMjt+X3ji4kO+W5+l0O7c7sA5HeS24vO/z+zZWUHMFE+mbl
hoPS1SS21mGNelGzIuOGO7MM0eqVEcAr0fp3DK+0XyAOhfnd8cGCAzTAtddONxBG
xRoDIGbDoKDxcI5H4zykXmWTP2ZB+K3VkSTA76xmeH4d4/lfMJzPjY+XY6vddiPA
IdKh8S1n4ihzWbAs5yJw329SsAlI0sE0H61RzMpSvoiI4+QZlvdjf02DzeIp6ylJ
zTGpcfWABt0gfg3h21CTVUq/p2GuxuELQRe81Kr3jJ6HmsfhKKW8K7RnvOvl2sqj
5ka9Pz3+1bscZ5MbXO+WACknGBOTeCIujhivhxmZcoQES8eEJrKDx3h1lKryfh7N
9rj641taOYH2PNiQDh1+tvvZ1mSNwZYVRme2lOT52IOANAHzOb+maVMfTKGWKILk
eDnnN04dOy+1m7wh/KO1VenXT//WYY5Avp8kkt3USdsYB4XRmYPl3xIr3RuQH6q0
iLgNL223YD3sED2A/TjB8ARc4Sj1spTm2AG8b8ZH/TYT+d6PDINMTGL53aj/6lpc
mFdLZB62IIKytiS8YYjr3Adf+/VYAP9CUogWwYm10yy59ouX2NyQFc9VAOITFFVg
pR1KZETmIoUHFJk/xtYEz14pS0OsO5SvAOO2y6OExYDrxSZWPQ55MiPZ+hnlC5Cl
ueEBFi5DkNuXU78u+U00uWmZJXFDPg6FSoTf5tVJ3fUZNxs5jyYi7Kgmhm5ipk1w
SCmKqhxZIwJjyZVK9hIbT5LkwnQcRQM1lE6TfOC+j5lI/MhOGjXT+V19/wyAZ4B0
eZ45gB4vJDC+0reOZnUY29pANxTgmQHUxYBHFp+cSPiwzQ20iGACLvl8J1Hskm4k
K5xUAorp7Vx3012xm17Eor6VYf2UzgyJ952Qryefth/UZiCdEtWlHl8G2GozQnNF
dnxBsepmfi9UgpMqHnFuWzOwWP2DbmHjsf+0V8i6vetVKEbpryquPXNhkbkte9cu
GVj1gcE4xFtuYViYBOjy/C1v540YUUSOHHvAZMBNB39v/TK6pmAWAhV4FExOBufb
wF9q6or40009dkzuhHqCo2TghvY80xfJbuy2eZGccWxp4+V5Z362OVg7efaKp0DK
ZWcFP/LeE5KmZ+LKiCnG7HJDDIwEgfnf/MPG4T5HX0cafGQVs06VEOvrj9iBdOAw
2XPtrtpsosgLM2Mc89DK2ixtwV1Hib+LkLKI1ZqABbB/0srsEs0ffxe29el0jAW0
Eay2U9CrDeGyXJW1mGeqvGsHphcBIMlaeQZCI/hN9SG8tVHjRSwiYq671LB+LMbj
U87QTE2idU75xsxFGoDNk/OQWkbF4gc8kYX20pvuVywcdj2iu96vkvI2fK4PSiio
VvIoNEsln+hjp5qfOT9uE+JnTduGogXn1gMcCz3l/QMlcaB6Od8CxzVZpiK9tzuy
4rqZFQ+VIyc8aECwkwvRQJaBKUxnfP3DGWeen4rlRSWfRFCOV/72OR8XQ40aXrt0
5uyYCQIJS8lj/8t+Ir5EY/RIeWK3k3gS0wVWATfR7lbwfQmLyz6GcFZjcQLsimK2
Ia7KtANF/lKk0ROpodcP6bfZdq5wnmXiVSEzQFa1/BVX/lKI3pQOBWAXyFGDxOJg
hyieaFzB8reuY88nvwnDMp2n3orU/1b8Gw+XXVQubD4m9vapi5wYyh0JBcWTV3j4
Q0PocWflgXnzZNJPvNE7MBk0pGAiC6owE6T3YDCBu9hi2zBmZHY9aaJw7isVXPJR
YTya3ixKNdZRZ84GE2A4k/tk/fG2g3bQH+lQdhcnUwHWNYBT4dPL4qWWcMgwGpAh
2RmTSWcuXAolo6VH7qVJ6la/sqtjwnbsBVBCXSbTTL6HUMLIx5bdHZTAz3o11M9j
hNLvA06VpXqyRI/McOcKorT9pwsEs6+BvbNtszoqAaD9fvV/TQWi04VZOHOzVv/3
8VHbDH9hVyg2sQfm9LlU1Jtm84eBGqHKQr2zNTQ40KQU7u/f5sVLUlr66XT1FmRN
SR4XIxYzGgvxSBbsqi5J6DVUkYKa2aV8VLBV5DJFYcHgmgSAXSCwGF57ArnUu0bC
6hLFDMY8Oeggpz0IQtvwaYigB6Z6KVjI3dyZ/mwvEfClClwiH7N8dbq8iiBh8TcA
141Wq7ZKFl+VDGu/NZ8NbxoQkG2Pwe7wjVvkJUE4bbMOESWworVajgjiWCikJWc1
CLVpL6xvxOq04/q8CNDU3MRWpBQprJfpkiLu+cfXwnAOmD1/DyWxY6ZEfwuNluQ+
LWhUFimJnFjsR/gXQ2xpmNDUEVjw4D8kT6jrcefJjGtpWaUVUGDY3NxKy1Bu44Jn
0dMk14USCfL6c2AuQQfefIQ+5j+ZzikgjDdDqbEaHL28i34wsavhCWooNyDPK5OC
NPLTq/D/YhTl8yFErpfZoOuAxV/KiWryzK8vwk6NGtIwWKWZ1uaLwyFU4FOAN60U
VijEg67KLpu2AtozTMngAf/UN4YxMBVtOc2smVui4jkORcSfjA9hphqIKxtnxDgn
ER3ONdSNHstoDVrzjcIuD9puwTOgS2VUK3L+ImjPVVUJ3R5XXNxBCQEDftfguRJI
RHdT5TwB1Uvv7TxTPr7RfhWT3QvbV8/G2Ux5V8XzoyYJj+wF2X8N1lIxTGJ5r9yf
m3sGGoxNCkML7whOvjc24HmA5DMt0zN/t4MJ9U3yHb5FREvsz/0BKtypmUMGC/XU
QhY597vsuMzDoW9+ph9HiHbJJC9d7zamL4frBjpoCdSYG+IGOr3EEE5VpWCfFgdg
qvrNrwYO42Kbkc/o158hX1sNKyBEOzEp8HM0xhcSSMo8RofT9zecVYRl1ZzzIqDe
FZvJjOskOpL0F+JT4W6v+IM9XMMbpzCmxvspBBG+/iK05c7JSUTIyb5r3saBdupd
xgWImFPkmGsFPx+gsU/6cJTIfVRIGOVDPLeK4g7Ag+4BuyNJbvMTH5rXpKtGoHPV
SDSCElQNzJcQqNqlG0vpBX/3Oh/D2zjxNt+GN9xcz1PK08HvwuG5q0d0MoeIOvGz
izMDtVaAb7rksSCXPbPTYX/Sur3KYv7TPbKC6mQ/aM4kM6Zokh38OeXMryGsg6vp
0rqNzuBhMOj03KnYyWuNunTS6a5LpsIY4OTxxxiNBr4nDZnLPLU8IQj1gT/nQUCu
QHgMHJMzIgkpG9B57EuovUWYMaJR4eKkTCNF+uHFnVdZl2+bHOdnTCc+eOGB2voZ
4lHqLRyU1IZBw0LDhyBx/o0bGpFmasdAAzD6fXuGsWW/XKPsrH0b30/e+Gy0YyP+
47/6Dk1oPuSpYqNj4gr68fpwHfPbtfzLeDiLIz62ZS5P/DYDkVsTL1GBnrduYWMB
sI/miLCnTK9kUxERHOQg1ugZdXChhmjpdvj47nXUv1brXRaV3CIPtOhQtPYMcaVZ
uCG7nmex80QjOKieFEnMexz1NOyyC6b2AhQQAILG0UOpPJEavYtw+lpBU2AwX9Mx
FwOLLghbXCby8XcfjPR2UEoPZU7cq/WLgoCgOXeSDSfIHKeqsbjMyPpcSvrvm+3z
c1JFawtn6yiPi8IViuhSS521uNTEQZcuXkQV9g9U/jgpBwmKf2hjiyHXA2qSNLJw
I7x1x7Hr+SwSnLSaW7oNlVFugFAMirTBVOaIWZxtcqCMdpLirkjqoVJg99LqtD3s
1QokId6WF3cqNZ+eukiwMrQ42yQ+gejo7RsQr5GXxbQ00JT/MWPxCj4e9H7uco5a
6nWqzVydzR+Umbhb1Ev5lnU+EzIPsWkGrH9xSK8D14LKYDOkpVWVL1JIvi6PVG9Y
GtCq7R1eYevv1sEk5T4CcKzcJmTT7NSpi6Hwus/FwpozgXnzEWxR3EYfPX0/z/LF
EH8Woboq/TSxhoWTknne0ZIX24s6neb9f13ySv9kqvXre3jqGvteHDXVLme7ddMw
qWQmbtgF0MuXkLY7OMxeDoPzriM91nL9JWGX6lJSLBf0XZ+4ryhfnrCxn8Cu+bMa
rf1D488wWpvfIKwPZ9s4yOcSqMp/HwU9sMwn2F7I4xdsq0FuKo94LD2tAslbdh+k
ZC9ox27JkmO2JRqMb1X+MXpJj1lGJ/MuhbuBlOimxVvU9lNtDjauBJAOfmQ+xm69
Q67CEL0qqQ1CNB/evd94CZyYZckulZt+Fw0DieLXqM1I1uIR4EeFP+6nNO0qud5T
Rj+9YXHisT7iKZ/ouLGIq8NyMVYznbDXDxVhZGNY+9kx8N8fQdezLSvE6bbF5Za1
CIsWpBExOdflA3qmES4Px2nP7zF9yoyOK6VngcXwsS5G2bZX4ekFzooi+YRAnPPU
Bbd7SnMWDqWttv+gQFdZK0ktBJDnpAoCKKEqYAQiytOPy5FV3d1VGvguZM2LMwKO
/30H51TztYAqM/2QD+37TSWCWdkcjxIpDC0ZGYzMgvPgA0ww2lij4ovoDbGcyAOd
1DnlOkzWTjxL/pTNJDSr2G51z95hmAZxqXS7w6ogf7f6OwaIl72mcC30W+4dhY1+
sjyLJrkLjOd65z4LaSKSTRvNtkkDA/bhgojy3Pj6gS6oIOhfxBamRVjv+UyzrrIo
2rqX0wAu5hFC78LoKHUM8GWK10P7lU5pghiTQZnnZSbBF6VIDHzhwm45vjpdcMoT
pKsivo170LBbM3O6215VkdAKgb1INFuya+VUqhUdE1uCX3uFLp+Jp32iF7DlquxF
PCrCwMXMGSRUWHrWUIKs8u5aqDi2e1qnJYvvwzc9cTQq0OCYM11gRsaBUpO+aRKn
3qA3twH4AUAL0tCgW86FrCjfBu2XBGE1XZ/RHp1aq8FKQqmzJD0PP9sw+K3aOfF+
ZQZfQxJ7DPPYqxJOD2kFzHr6kjb3r51tzcWaCAyThmtR9dtCRbhW6m58+e1HwSNd
aNGlNn27IVIsRgm2EdnkIhBmiYPYzXSzoWddL5SQs2gV+T6AvcslIiLYWe+r5o6h
7UUYQKg3zraKhdt/ACy+gtzrWi/4a8THZXu8fUwNkNoEovrF4I35f0bcu6h6r3lu
8bXf2QNA03h1DNGulZ1QG05o3VUTJQcPicf3XXSRQvmJepzQQ/QEyWqgXfn73x6A
rfhad8+EIAAKt0sKFdbp2TeJNsbrStXDFeF+5r8M3tmZT2AI5EfYvSGvua3rsbxs
fjf1SHj3t1vB3hrvXkt6ZuXegvRRtFrhOXSHu5F4Xr90QIbLmLC6HK250HSNVi9d
2WF/QZsOxkkPAvv7Utqo58j0/pkBMtNJ/7pNdCO1Tl4Y1Hf/SheXJKJsjzFvIf1o
T6vV0G4VMymYLcDG5IvIEbX0+cGfL88/RzXJxt3SixqNIaEzH2UOMqIE7evxCQzs
R7/CglBUtvscy0ced4q/BqSgQnKZqJVJtvb8APWknse486C1G06O87sr3s6kBz4D
Xnhmna+cbS0dV5gziUxCg0T9GybQgaeQ/q1c3UQS/YncaFnzFb7IQnTBNOqfXhif
m5x/oFAg7qGUau54t0aaDa0+lpS1zzatOLIaPAcRrToVIZSj+K9OI366joh4RJXb
jSxsUoFVbQqBdYf/QCBDfIe/bun1+4XVWcN+e/51fazCVv8nBWiwAv9DnzDWNqI8
QZeB9SwSkCETJPGxU5yqjaooHAaMae2nTfXcnCa8zQei7Os1hdLXMdQsk6q+VW68
jY/YboDCK7vc71jf/tjLaw2bKmJBc+MPrGgVahDjsE2INI/Ps8bUfx60QyaoiKuO
jtUBs6TKz5oRBDhr3+8d2L90Birx0xExdwoZaLt+f0kyPRQHVd43TxQ54eUsJ+0p
iwNroXnHOXYiLujswU+oQspLNBI7MPMP5WvWqjoa6pdhomCk8e++J+9qmBgrKaeF
AflPyFzHsYQgol3ci2n/fcl8hwesA5lxKRwwcBOb8xGd8OB98++M8PeJKvoV21nH
5zEfv1IqK6kfZ4ja9hYz1/QQbsK+w3hHl37PqqZMXcq/e/FAp4OJV7Kh+De+oXao
SrougdsKVxA/eOTTJzBVU7oUSEBTq1L0kceJ5sFA3Ph4l3NlRb3P5LzzBZ1QuxcI
e1GI68srfKfti8MLP0q9C3ALzopO0KmeAB9Am+oNjoNvuXa1dMQMnWRAGTt0GInz
bmfJvuzTXRz9H7dq9q9hapyks4WbmmXkfAdqJh+1ShdAPebWWDyBdJK+le51/xrp
DuYDxLC6GowKXDW/ibNH1tCf8JMfSO3fqLdFLr4C1dovP2MrU4A/WxKtHmQdmRaw
Q1D2bvkaQSXVFg0bfRno+h2gtWJISpA5WA2IMyTbWISqqLvkD2kn570IU+y8OsCO
ZfQNKzK8Z/AfWqwj5xj7pkJAioKeKC5ZvJBTJNuQxzPwO7Mk9LVk0vwJWsOUULU0
m2TdlgRYTen7xkXqDYLsL282WPpalrLuRJfIBZSFt8NneJrl6qLheit9F1/EnlPf
pQyiC1/OmZgZySYe3Ize3oi3OcpzmVCmxkOc+axGEGKw3j7H/jRjJR92JrI+L0G9
+aVBMXWYu9rsLrwoVHUApJLJfYadTCgdiZBzCGXiMs/y5jf0m3NhzmEL7mmuv0Vl
Bo+PmcRi0K6G8DCfB3yG48v2QyEdMw4H6ioHeNknoWJz2giNANmeHviwvt3OCpyu
qfev4puPCOazQCG8HkhScevvox9yVFLodhM9pLAnIlAFFPR+KB7zU66Q7Z9k1YsG
8fxeNsIo+XazI0gsApBhr6XTcvmPL3yCgQmuOjRu+WbYU9EKx8wqaQf37pFopQbE
RvQLI3Wppi5AMRaJjzyAVvzdtD1r8OazGFIeXnJb4kTX9RGpOss5BgYj8lzWDLpB
2syA7n8/miDQpHfNKOCMaEwJmtWTSdBeyxChwGoAuUEbHVzwsC1bmAM/Pa5ODOf4
JSAewb4iGx5NGccoXqiYCU00+lshrSjJLshKnE3q2oGRJMknnWyashtHVsG9wvj0
L8N8PQHng3cetVqmiOfTmqE4yzNfJkNMtCROgoah1H2xz6pj0LIgbBgYAl+AbYVJ
3g+gPcSmd9XyS2+IG5ApONpN1d5lQa3C1jfSKi6uOCf5Onc7hDItCPJgB1BkzR8R
4g6vyvjNPEwMz9wwX6hi4sEGmV+SdoSeH8ZJfwW32B4AfUhvZPZXwh8W3sCrSJPy
5/6A1zRYITsXX6ZSJabS/B8cbuOR4J7Rfv6M0oylJu1tFYFjithvNqhIikoK5s2w
8XPakzNlq9SpjVpYhidGaSPNlCYxANfeTRhxdV3iUPkTRq6HNseHQT3p9Xeu5PjM
JxxvD7yvzQnNr11HbZbBeZqbfBwhYDDlvJmnyuNewFGg7UV03Q9BEW0MkF4/Qf1K
7K1dqxdiaO4zVAPCgP24BkoZNzhZsSKvIJkDBFuyzodFbcP1YoYsqxNmmN1cHs3i
BTLPEGnaz8phq0pGcR70LM5HLG9NQaRLqjuaOglOZ7faLhD8z8qyOZ82ti31+j9W
2qj2UlapD7+HiSPJjgajp5kGss3aUUoiRS+KeQopC4pNEjeP2VZKiMXFpP26VeqF
4XnQ8j0OoD1Q5JebU8gVWVlRWNTqbi6fkBZiY1GEX/is5wKt0u6xMbo30lmWMYRc
5q0A77tnYwkc3AVRXNud0wwKPwZONTeXrck3xcw+YzfHsupt+oz5VwBo1qWtyhJV
h5BMWK8PGmer7zN0GMuTRs3ReKWWscpovNYt5ijOlKHRX5uSd7y2W26anNrkmn77
lTa7IulEFIKGz3G5PS2DErhbRVDUgBbfTvBz4bRwoEuSIGPFNx40SzqpErNYdO0P
TBA5S7dykAgQleY+EIVIEzcPR8X7bWjv35Uz5qrt2vNAAyTDylzucoJ5JYIaOKn/
Z1NcoCD4JRINsVJqHH+/VvWyObJwJfUrXq+YgOXXGGvZmha/U7Xum7SlCxqfxN62
njT51BuBmS9bzwNMyFJjOHpf3kg88RzWr6mD9HYq8Okvj3NVK9Odf5Q/Lx7aRK9d
6G0DtOPiVJuNLPxxMV7L0UKHibS0mniwfthZjrACWBa4AcZRm+JphXm2yoKbX8GV
kOyyHOxZSnbfwuqzt1qqIdsCjLXbGgZJVbE6f1GmBCLnfzI7S0ecw634UUhNmHZF
W+SjPsMlWoEalge3qLlEqMLb1w77JXNe7XrktmZYBT44m5o8SXHA4JI5R+EoyedM
AE1kgqooTMm1spjaiCmt5OG4sKW8z0j9NFUCTCUS/b//QQA+bWARNrFIu+ySLwa1
su6GQyRWxuvpnf+Q7Qv+OtVynyAeUQwjON1sTroOJDuDACALLEBnJCobR2RtlsNb
huHrlpk2OnP2X8Me4cTyol7W7kNlmbKqej4hVP0VHe0sDw4sDSPIvAjck2I0b/Hq
vdw37L2ozal9jWQkoUnbRd00o5KYrqTueikn7S7m3Als1EhM7d+3S2Oc3Or4nnOP
NWN3ikFG8mKlq2uq6SnO64/b6rd+VwnpFovUHYvGSl6bazN0vBSlZemTchwU3Cz6
WKsWZ63JkM0ARswL+J8fu2DHhd5egp+yRiTVYsF678DMAeQ4mpXKwC2cnUdFvX9o
WUzBZNtqLXR9V/2miYM5iOKys5NLdCt2V2m1bBX33Sn3A2FcAhzB1f+pwymjdxQI
ifMoQbp3EGATBOQiHAun0Oc4cYdP1xNJICgyM4WCFi9emckTj4lTKAaHS27AvUip
FkYZQqOHaAstHHFCHUH6FrhYN5UEFsf3otS1WzyMM/5h1NIMzUcaXN+5NMboS4Zk
+XkxQPLjFCFhyDK0GerzTJgp3QPmBlAiVS+pdiF89eV98fFDGTBwq41fub2qwQJ2
Z4cMpoS6Vc1svXT8hcrUhzxCEIN50j1cUX6eZFjwG4B1vvlG48s9DPk80q9i1JBW
MUeEMQacZ0jm4yXjHHXkTH8HmbuUmkhqs6zEd0a1g+lk66FyRw8SaBgaGx69+fEB
Mc6mF2USsCC5WPduzbN4bCvs++2P0GVde2CuGj/URzMyC1Y7TMh3GxbdaTfeIb73
NGIkhWtQNjN9IerUCYWck281DOziRie9Y8RW42qXp1xm1RMv+1wJJqyRdeaynCmX
AoYqm8RJE+gKgykYlju/ZHBIwMlVWsnvpm/VIoCIm7r5kpbZ9FcvAXi4Vk59sKiD
SAGVOSxwS+Zdh0nxVwS7tG1ZBh5XMtWDqVzTr9gl8Gv48aLsdoW5vSmumi7X13qr
XhO5dh6KM042JFXyciVHBqIx6ErWYblsJ2QgwhakHwDn1SYwW8aQrdqXJ0807TVd
7Waj9TNq/RguuUs1UCTS3WNSbLoUsBLwAH54Gg60+bRmQWlqY8QDvbAGQw5XI8V3
GITBzCjZhpfRNBANw/xXiRhMWQT3W1K0dWDBt8oNuLCRX9lawwXQ/dXBimQUczWF
viQ+L+Fse/xJ+gF8v977ZLjf4AUw/2Kv13L+hqpqzU3UL8K82i49lfjhQc+1gdCT
ESC88hyJuoGmFnxQISkpW6k1U3Ov3nHunmauXPL5lEpXhpGFCk2k0UU3+kAtLt+y
bNVrj7TOXu+x3CCP1PRjOzGOUobpjyhpOQZi6czrtkA8doQmi/2MuH7sAOOVy7US
vljHf/NZ0NnYAn4iXNbegsqKXt6pU9mSJlhX0/eVUBsGgDMItj0/lHFL7nbcm37g
IBCMauR6lwtIxIkbnRtERFu3QhVprJOcb2PmX76Wn2tQCtk28quD9KRGxXoVx69T
KOhKVPY8c+BYdZWmB7T7skXW6Slajqi4XifQeYi9/5WCb4Gfs7vXONqL8FqXDkK2
2UAhV/5DBAgiRaDqky9yFkckVad5ELhLAysg8JjF6it4pElqtj58158y3zTuuFev
edYa1kmaW0l3vAcgiFauCw0hZoeDj2KadihR/jqAIyBouz+vw5GKX2UhryguQjKx
BJhXy/tx4IV478f2sNwoBvfnxixpk4LQye5tSG2ShUCuFkjJ2nfBWp/4cLnmEm9I
rm4tWqUFYHgDlE+LPvz23vc+ZIzsVg06q+ePGPFC3kneT8j2AsYwJW+d3Cd+lfJn
lJHTzf/4zHOM/ONOGOE/jCrJJp6CSmUIsWBEJEDLsX0rkwWnu8xlJG3feFa5F+0M
zhTE4goG0/KKWq10gYAsRfzKb6Y6x+1qGQw5I+CBgUOuc6Gea8NaBKvNFCAap1pe
1TSK/+lObGI4MjxlL72m9udegEYdP9OMnoWXOV+cduF8xeUNNlYnGwBYC3L9NJS8
dfB1oYMjPJh968uA4X0FMv/ocezpCraw28/rRbiC2PNGRt1NQG7U+NY7Fo7cNce1
u0XC8pte4KhHadCHnSbqbikCI8jup99//x7QQ7WW+UJkwEUYYMZJuBa7d479dpAa
LCVMpRzGwAxKupYIKRUKuYgser6+fvRi4G8sxVshvyv3uX5dc8XNEQ+/Cxy/Qykh
VKE+Fc9830imyiyr4RybRe6t8MyB+gb/D6IrcntrKCwQkGspxKhHmut8SumqkWJ+
Uopyr3R3RYV4ORjL0heKmMPfeh6hBCEJFW5bYxNCTtHH4V6V/dqGt8c5p6Dez8t1
QceUf1aZ7VRNuLTG7frzBfgnFSrcOM5Xx09Jsr9dJxR5rmvY1OgHDMLNaCBeI2jM
wB9nu46QOtDZfmuZjmHWe69B+wm9SIamvLNeoDLxcE++8GX/Hodt7VaMaTM4yfXK
KSe9nf8w9WFvezARykIvaW8Sk/zrzf8X2UMHJGGtpN17KD0BD5AyQIJ2rFcT+ovk
sXmR90hwjFG3gMrOTDx6RJ8b7qQwmJhWOLxYgI1d4gVlQxJsNVc4vrh1ACEkGqGT
H1ZebXLuhcWtiKZGDasaIHzWfhrKXvrjVDD/tTG9J8NlpjY2ny3hplFGDKvJu8ib
xbJIG6c6dWpw3lFKYJYRCz11AOSewnmWrfY7KUg7ygc1C8ZSp0wb5dhtyzpgsEWp
RJSQvLYTdxzsM30I4AoCNFDa5OOssKMVwNctwAbju3xijfDd4FwsCdl0aRebTueh
vWmn47hQ+HA28DjywBfObH829sRSneTHgEqCR2uVb2xmVCX1oehYUbjVOg/xTEvq
HQIDk/djHGm//1FKnOjVjWRid3XSNJeonFt38bXxOj0z1LcD4sK2jgH5eafTxwUR
QOWu8StsT/NZ4iKOpBsMM5dWHwFj2lxNuuFjKg9L1ZHhCFp9iQy0UJCpN7THYJ/U
QxXX1ZKH0/NwsruWxXlwbPHWlccmVus857oZthUP9tm9+iygDmd3CYIDqrhJg8k1
p1JlNELbdQX7GPC5UUffRyvhk1u747eQb/SpcuxM9DYRugoQgeTe+NW2D/IF3/df
cnTzBDIVOSNDb9BkUVPtgMoEB7T01vjjXd2JbfrIcbv9IL0wsNkYd4IRiZG8KA2U
tZOo0uqDwVwNJ1dCZOFi3nEkNs3NfxluhxFdyANhoQ5xQgaERQPLqYWuKI0myaxr
QaA+Pqtw4ysryAo5kTOtTcJvUGmQsLHH2rDkTORcAXoTXN1SwC2sTtaijpxCSAHb
daD9YkSwOuL3Vv9n2zlGmYRNUU5HOBeKBhrR/AoiLNjU/x+G2UgR4boo2+DE6H5f
6Mm9BSMYce9AgPxKOvfOBplGHdrk1ICrJPLeZ86oA6OhjSCrAz41E8oNO0XTmvSI
XTE/WpN/F2CZO63G+1hxlZXbJo5AYpg7k/ypEF307ipTsqVHP8+fZGIr0nZ2zF05
JiLZ0yumqMyu96aYYNJnMKc36Vbkg8ijw08IZfDFxm1BVUhEMTM7jAwBxG2uN516
2+YzzSuZP3Y+W10LNvPzaofIgDXSr6PwSkl1qWMNRQM+kffZtLeWEzDgcUP9dLXw
jRSGWW6+MtK0MMGSpJzsjFDiXcJ6evUUUUVtCXuqGSajOB43X/wpY0kX6/mcgbh7
w/NBPFYgrMpsKpt+Xp6kquZ+dg8WgJ4FN3GqrR2+Av38gtqNgZ5PmG+NIQ1whzeI
3j05FjgFTSjYVY6jy9SB27ciEcykfT0BbaSKoWodbNRubs6GgcuJf/MK8glprZfa
CCc0IgDEmMfcanvkGbUcXm5ZxTOPszmO8Ad3MABtuJbvylLAy51ZmnAvL27sKXZY
qqWrQhCSPMww4ANGuaAGlj1L8kXHagJmjwUaxjtILxx4Qr6oezvIDR7fVhflFp6A
leUySkqV8q9DAVGz5OuVhGOFcagYuUYtgLJj1doXQA8YOrfZIpmH0Vmvr/6Wguqm
LOfpIOtPcA8mm2AOj11J4uyE10B7e4m9v42QwV/kQy6fbNvrio3haNjIKOPJEr5N
6ezh0ENBdbU7PxjgiQU8mnMgy6fvkI4crFmDyuXvMtvC0S7HjVTUYStUzbzcUDU7
V/7oZ+oW/5Ong1TDEUsehRQn2sxpIl3cSIW72BrumvkQNDqitJ1D7LQoL548PCKb
nFiPUzY7xxtKEVy00818G1FP5s8mkgxoBJLvVR3S+pNlVhskd++Bh6fowS/dyqpD
e68bkG2j6CVuEhm0nRr7I3qhCeJ5q0qHsR5SM+WaHHdUM790TDZujfgqzihM3/jU
Sv5/JeK/SqBvvjE145d2HzoEC3EUTyiiMdjTPVZ1dr27LndH699R2uJUQmAubcJF
BtHzUCrKHAFhsPi7OlSqQeDbIISL9i5tugt17w20MZdVKlZ+g0L341+qyOzjX2A6
zlK+tu1CFVP+W+0PDEoZVwTbsNO1HnajnTumdeB/nT1FMa3ujC5gyqEQd+hTcuoc
VmbsLHZS3tRs2TanLrFmKA/hbJnK+JE72E49zr2by91s2qP5kwJJ5iOS1+/uAwGE
p1Uld7kU93D10FP98ixOdbPik4c4EZk4ShHL4wQOHFHmTpP5bH0npm+1TknrYsBA
SBc0BtsHhw79ibyf8zWX6h0DdWZ3zebtNjeP5Fc/G1eaXXFhusWzpNkH0Xxw0uYe
4xQx4/CJsvyVma1KKKwCa2RoJzBHzqDgtD/XkWHDZ0IWxAPzPuAjCeaazDDt+pPt
tlCbsRYMCnRIjxlSrApJJd8hcgeANKZSKjS6EPlkvm08btCAbSbZu7VnLkQbn9oc
nO4jBJUzG5fQXi+uYttSgj3yp/wLNh51W/xmbeOfTBN4BcV+jkg7Rvz/ORin2Ukv
ds2KZw9/pQj8uv7m4Bee9U0CTWZDfpzL8DBgn6h840FyEjtXp8nMrCdDajiB5rw2
WTJRfTrUDAMRIsgXl6MBsAStU+9qPVqC3JuL0fheHeV4hHIYDv8foqXE4X26gOl+
OoQOOAntUeRlfGBpagpFekSnLtPzA89IA9ofYya+hDpvalXPQnZdzsLNSlM2iiBs
NMjQ7T6q444nQrfAJbKxYzGY005aA/sviG6bOrBpzvkYotILiNHCvBaPKqFJfgvp
XgpdoVWjiX4DLu+G2gGV3HZcTRemIQjVkM1jaRPjVVgVvwoCg39jdVRbrtbcn1S3
1xILUTV+mm0YsR85crx8+/SnOJeoZXMh0RkSHcq5iFAn0Au2i3iGB9mBDbiFvYtB
ILAMj3SV08SDxcoZ5XuinOtMfIML2ftfa1eBrAfKam5ZgVNoydEb4pesE4gFQCAh
Czxet8RUhYnpQLF7qrR3cbTEyO3X+qUaFGK9ZkWjwpLqClD0ngqBiURVhFkNu5xA
cr16601qVMP0pZA4kT95j+0NwfaARJnkZuomGZv6u27Rr0YAOOh3bWaloJsfUFlu
59QX2U1phs2b27azEDifrFYsgL2oTfLtgJ0gMexVOnxCMJDpfXQwN2KxWYXNopA6
neeFHCLptDNHjnhGliCuDr6hS03yviNz4manm1pf9W0T0JPKYkVtbBXsvc6034QQ
vho3HYndvoWtqeYTHdtOtRSHSap6luLV+ybrJLHeCfFxIie76Kkg8dzwVqw4tV6h
+f0sp6Y9BdmAwtSUdoPWyc+rkzU+L6PUjx7/+KwY6IoHL19INyMvOlKyGyeoLVXi
3aao4eDA+EgWGNzUwH70tDZHXoz+MTevm9PgiwjBEvwGFvx9g4PTNrf8y30kHbbv
cN0jGOBCNVwn6k86HA5mEu3WXx4KCIhN7jvjc938O/YOF09CaG3H0gsSdhHSSS25
bqa7PtJvW50SY9BsCS97fUHMVAeewejFI4C7wcdrLzB7r6ht+U9c43zpQtmULL7h
WSu2NBObcwvv5w1CCgsRQFFeZSgxln7wT9vytZtIoeyfWJ11+wGWuXg3Gw2/EqDG
cQG0vSY20LLeolI7mfhu19U7uPx63hGUC/1YtJIj2cjsx+bKwCuIqrNBI+B1TpLv
AnUkfrHkCFYHgBUcvdoCpiOjt40f+0qhDokoAmShAWWgzcyVEUlczOg0q7Hrkg6S
lIFI1sV/FWikescG7UNqJHffVtLmAjzS7Y9kgwfTiC6XCZmqxUJ2NYDOzqTb7M7r
k6QZavhStlFrpGzjmPNW41qzkp5OGa7EHqCQXWm4VFMco+tk5c+MZwn3I6N7fVWM
m9qpN5WCYJ7W7l32l135hIsAzLU0+bvD5ot9uG5O073LjSbOmV5c7lqrgFgCz99/
G6kR4Su1kPWvSAMujc8tGMJzuy+OmvFFH/kNqTKw1z9/5ZJrZ4dPS5HO5fa+e8xA
b1Yhn51zEf4+eKlggaiJW3NX2SNv40pVExuc/g9ckqoJTCA6/n7TyjU+inn+ICzP
iYHNgOoRBDl8enH71e4nOhfqlOJNk/ZcDUr0vwivDVgG1sGQIcCMaik/n3Mf4sHI
XGcCZYtP32dds8OM/sGZcn8BPHI0k+R5X9EThgYwHUzBUwAGSlpDRqCQvW9ZYr9G
Th+9zoqhEd1X730oZeQ2tcvnJkqYVeVXUZgmb5of+pDtl+1xWaG3bv5VRkhGXuGJ
6b/D2viWZlCx8mxuCgQePCDfDePZ+UkISRhwX5HzrTeOGzw1oUKQsWhqFFqIettf
M1bal3Fs/Q6yZU2ATAjdK8qGxwdkU//dVQvFdNPRatHVDpePqAKMY1GdQzVaL7ot
qM28bwBqod8EkpQ/maQbYqPuXjlzXRSGL9p5OjeSHrkbFiVqY8heuRYMO4kuIOoe
uCjbKu/Dy15hFOkr3btpFiv0RjWyv7RgGI0FuB7IzGesoedTTGw5Xp1eSCkEsgnw
7NnCcYTnnOnyg4/7Pg0FQE56pLR2gPUu28BM8IslhbrSvmhnZm+PbwtYKh+ZDdYA
XuCb/LpTwlv/zjv3cvkxLLr/DNaRzPdOCGM4AIWVdWXvDySrpgmyRMdLdo2GPSCO
lHdt41PqGZltT2Hp/H0CiLaelW24+wak4pkuh4NR7FZwd2qvsfI08XevUGn68ucc
8B7e8iVGAtikZ/iupSWYzcgCmVik4AikMqySH5+paryQPRUzo2WkT3WyNoeL87rF
b6zBhPuPzkH3IGV/FMJa/0wmDTvXIdyxIVYPcAP7fXgbE6aIvyQcKiiH+X2Ij8e2
nLhQDQfwDkiD0zNLc8tOPVWmm7kXRIxFSbogH4jmiHT3HR/hWKIyH/BpB/1k+D/M
CkktQGAlRhB+eNNEDsu4Slr2aD6XVTOrzesDL9bkWGCXuO/uuMmEOB53O4iVKlf5
mbMVH7cosKmY6v/RN0bW3FYvdCVQ8+lt+b8AKcNjLT4bjfv9XKdey0tIGOm9OCGy
Hw2TPhCI55Egnwsdtau/u8IAVrWaP2oM/7mJU3LvreyQZbTO4yry+WZfVJnQ7P48
STase8evDXPCsYVOiRYy7vwcTOvMYvbYe3E8bInnYA7eF32LmivYx8nxk1EK+Wp8
DDOJf3uIGXq36M+rsBDZIyEgbpLc/6uTvD5hBn4lOwS2rHmP4sr+VbzSm4g8MyaP
0lRbiQl12ZUbGc0cVuXigwcJ+aFNgxZcjpXJgo5ceT9N5Ie5mfnJrj03gcLHTrk2
ikMYZR6nu5ufkHxrDWAdiFTgYpYpngKAzmez4vU6WLCNEKjz1gbpq8V3RFrOrxhl
ETmKI9mTwpkC9rVoSQdrw5v8u8JLVC5r2XswkMAhXcqT+BYBWXwIZn61MT86j5Lj
awWne0n7UktXfAVShmTgukzaJjLTFvItnSyCtnD/n70ucCLOQTHBfnPDIb2wjlD8
mrbMBRXIxk3htj6+2jKj7S9c2N2UfNo5WwUyQEqjQhLR6fw5y7UG0AaAKyoiaQda
42edF4dO3gzlATOP9HEecpNwahCN7V8wUn/VAoaGdYuZypESzMALs+gfCh+6I9bo
m2JTlN9opUmhUm3rHBRa8AauZWZcSX3eTVozS+0PmkFUfEUit5btSQ5sO36nc86Z
mt9EeHCb3hohzV7LKZTVqIsAvctoQJbk2DYFhR+3wQ3WQ1i/X/pVLDuPuL37UBeD
DLmCBH4p53RLitsZXeozUWceILq4aoeRS/PpHwlmDHl8BIjrDDjJVhOkyeeRTJWy
NFwALgKjEzViMuipCJnoT3IQonljjlX71eaXWQZhy2njaUNp3+ok2jL+yAPkbtXW
w7Ptc8wAJZ8vbrMEvBlbRb1SrH0hnhM32UIUi9TbMQPV6I7hxuUah401z4OlI7d7
KQkZhAVN12tQ9jBBUbcUiGZDFlr2IAoc2l8CXg2/pjVc9We8f0Qp0YHtl/n/CicK
Ml1AIWh/UHjLhVmlnETR4wA4Iwa5Oltgdd+dIngel6Hhd63iP5ccEyGwqb/KxD8t
429XBVvjTj51nR7oGj8PlFv77cbUkW6teQvhCE2htk5N0FdLcFG9goujjv5PvLFI
bl5Ui8BKvPEdcnTe2ybiAOSxbijpL2v0p8oAVF2sWPeFqLmC2XczsyIfHrfp10B7
+J+JNODmmvrdxKWiHwHR9TJaseKclDZPhpwRd3LfTvjbP/rhXLr6d/p20HGx1ptQ
Ho9gAx+eDP/son60vYD7ndSh6fDTVy3fGUBhDxqeOjq9bkSPdbtM8VrjbNRrPjFi
hSpvvow2IZ1nhrV8paQTtVE4EcI7FIesaYlic2LYBkVsGP29xLbJP4rVjQBOqc8N
SouUIzKfk7TVURrQEk1A95I+vYFft9Gao9tWv7eLwtEwKViMRWokGG5tnqdPkc45
9xEf7jFnMoplYa0YTEWk4619YgwVflI39D85c3tJivnWsu9n+MiVR4TRAN2iRgPT
uT0yC3o99cx+9cvhAwT0akyY41MjzOm28k0OQc4Q6yGsLtnxmE1IF1Vql+FG5ZeW
POnmNn8pDOeH6+a7N48KgHIGvccCRPFBTrGrCdbuH50/Xv3ICPE/aTBeFJSJt9NM
OANyJhXnMJBJxx0Na4fjAwq73t/b7O6OvEZw3+a7u8lJGDd+L6FkXfQJ75J9rccy
ZgkxiDG890NVCt0xlOPr49A5Nyw/bun99fKEqiaUsJl8KlVx8zt7Erw1soVxIRtE
19jRRJ/Dnw8aXX9P4DiJeZLiGuUt2ZZqOKl9W19lq7rPqrqzJJv0fDnqZjukEtBW
aHaFoL65+KHQr1TfLOuSvO7jNxjCMXNsNEWDli8UwJW03Z/fE9zRUrlJYmKeBohP
hG+od3f3YMwviRHlJDpdD5ixRzATwwc6n5I7hAfiM3ks0JI92PybsXqY2gpddVnE
vEWyvt4aEJKQUgA1GaFmUoTz7zQNdI8hMJnHNLZJJtzjULln4a7mZG/9RTAiPPYU
0ZuOI7/wJFECn/m0cXEBizHhVdmTslEN4YdNp6bKIs7fa83GAYxxyupx3UoINMgz
3F/MG3/w+s7BOJCTo902/ay5J3KGdKTgi6xV62oj4gv8PCne5Y3bkWEnAvBWn5Bt
6sWlKjcTQXTMj3p9lgumnB124Sw6Dkmtk1Xzc720Mhhv3HUbc0RRx2QiI761CMh+
6PJfxfhrmeL8oCHpDJ5QId34QJCBCY9qH+YyONN3TTiYOvfHCHii0MD1bywJCzxA
f3+w/b/34b5rua8SiGkW0FTmHjjL+lJ7pYEC9BdSnY3CtXZuZuFMb6UL+ZSpIptY
vtC/acoT5Su6uTl9PE4BtH9z2NRY9sLn3tBC6ca3tDwu0r0h0dc+URkMebQGAgKI
ZvX9Y+NcCS9RXyrsJyMRm7nh//b6n68DEwmf1nzivnjNGL41hPkiwZWcZArM0n2y
glTIBwwifQCAUa2jHTgeHGyYn97QiteARTISBVReCkT8gIyZwySTp5/XIXQCXQEx
7PLtaFQw1gQKpTeTzVRO8TIid1EO/aDvzloRLW9gKaQ5D0rZfY5WP/zXy5fjAgL7
hdfPjA6+/mShte1CpxnjRHos8hZ2THSfaoOsJWmbaAQlE9Cj6VSOvclaJlA4gSlM
F3Ab/LjAPL1j7H9cuTQL1+52rdiOrq8sZfazjc8cCmJvQd+/0GDqt+qvC7cnpizf
YxBcT7L/jtJ5fPFewrZxQXeBzt3Ez1FunnoXYEXHDEMKKIyXPdDl+Mn8qdp8cdVP
KdOe/TPdKmHKwUV7vieRhlEu/tT7JSc3NWryFOc+g13X2Q0V/6oLuPkRD9Dn27D9
DjKgxdUmO2AtJgu0Wf4pc+V7k5DUzq5TxRCzK9Ts+V7J8qMP8pqL76VYOm0ZHW7a
fRfKAy4LVf3GXBiIeApQsGtCWv20ppybG4+PXMFa3m+JOwGzQE0hGvXVJ4zlA1xl
c8+21wAy2xJqJmR+HmO7nOyNxynog6PsZns0hgNHqq0kiwoGFFnLWrNBr2oAugUK
9CwlzosiRmgcWiSmQF0TgWmqMSo8kz1zjWamqeUaDz+qXRkyS55EzzRjfNsACswH
M1cMXhvhcoRVqS9RsGv3XzyROQBynByuzc/a18LNG9QzgcTtgUk0bRUpAD/rok3L
m4PxISsrr/LT9stjEeQnNFPWDhO5b9B9k1TeOq4nV3OCMmzuWaCs56EM8i2jvggN
SK/g0joeJkB+j/uuwUnJYcO17oDrywR/2Ltl4xJizDpBiaYxDRU98Bv0k9rmkeqg
DwsNlKdqJKqkHZUf36N9murrJrr1OFYVSbWqtEfGhoz7x3G2gcZdKd2yRzKnjl5G
X9thUSDMVaPxgR5SARLaQx4TE9Lm4gEHnM+TWEupgViq3j3p8hiXIVUa2W6TZnwR
EuJZdUlncmii+ztgt6yyaCKYJxvECf2kGP5qwGOuYNDR2WDJGXXgxmVN4rtEVVDh
COBoFXarOAqpCRI6y4N75TOY9V7VUpOA6a1Ac4S1eKNj9TXHD0vHhAAngQEUMa7t
xTYz9v0Rps7nac87Y3gIsvQePk5tqmCC6h9Memje8LH082rTQ8ApdADQDwqCX5lG
vo7GflYVQEKux705cc7NHRI2ele/E4pBnrm0FO+/WdQaUJglO/LSGV9meu7iJRnh
9jTkUrPQ0o22GRl2GqTe8rjBCtD6dkCE0q0JO+PkoOrAQMgSkGSGJ+JzrSIRYOZp
MP3HkYJrCtAH7Eto/itJIXQOIRZl2odk79z2wmHfmbdxnrsI3k4c10CrRJujg0to
ZTceQKrXempq/SBGAY28NY9w7kDEHy4sAd1/qGH0cMK6RoLTwUqYG7FhPDeRpRrV
P9mYjLA+YYmKk0txKNNN/SvNSNHqDJ/HJmdZy0qqLEeEXinsqFgRmWdwH+rEErlx
8kgbrUbO+WHM5+q7lkn6y+YL7pcZ4OZVkNy4MdZX04Rhicc0CIclgAaXX//gXz1A
wl7Kxb0xCb7l6E34shiOQJn9gfpPTA955g4snl6ieUTVjUoCU7Vrb1lVM0lqL9cL
PtyBW4XfKlbv1kRuEw3Q+0OI5hS0/CKnR4cfNTqpUPuHJpirOMMqgCfuNGExFUg+
plcisuM9ba9LgBnTs5q1fFc3zdUBrDqibJZiRyivoSfrX+1AjvPJDj5Jvg8PBfcz
8/QAAwuNyYbV2NRy9YaFsc68Y8R66m44sla1YOcgJgCuVvlOKppUaEAKLA9oyboU
DG24vpXpcIajDB+tiPkPniqWUiI3iVLVcoxV31YF/mj3qjyD9hxkB3z8TnOwHhhr
OJFOn9YlnEhBit6MfS06CS8AaPHMXJJ4qtwNUZ8pzEncYCv813ikVcnMPgj4oYP6
prVWWan35ARfea0aKpjWI2o/FoEWf9TIZMTlSpV2IJP1A7QeHjmbj2FTptbg2QVy
uhNMq3iA2QOHAiCZeC0Zr/GWfZQK7W2PHa0EgQQrRjwMcf9yp65Lxe1ubVDaM1K+
4eLG5E0O61h772bRg9zKgGHLzyJ5cZ1hLH/EJstBIfmtmwboX8XBY9tPjokZQfVz
ufjO/QIZem93vWXBmkKxs0qKegzpngyjipfQcsMPcnRbXx+7e5Ew4EtZ7YO9VVWm
vqP+e8rM3YvMuKpOkEGGHWWkYCp/Magb8F4pyFxxwE+K1I8J8nPBFEyfPSf7V/a8
nSPwTtJ2a1DqkitSRD6OBWKbrkvByZCPYj/ixvjBHbqBETRUeKg7AY+9BUsvpaf0
PV6JPuUZs/U1e5n+XY4I/Xp4RmD4CX62fO2fyhJF+Wv9oiK9ixhjPmAaAC4d2jAH
KAT0opXrjWnjJ/teL/x23cZG3iyvm8Z9aTcfhp3loemG5iBWVXUpm8pw1YBBXYAy
KSeU3w3QBweoQwfeRTO8QJJLEMJCpaImXpZSBHWKzndHaAFx+QWHh/UqDG9xLnD7
OMHlYHnlE148bydpE+v4mEbpqlBU20smE4X7BFh8LjhG1pN58Duk5lsRQi60lqa8
gwM2LjDGHsrkwId5bnV8zOxmf/B5mifVhzCfR3I3k52hF1XgBvtsTOvC2CD41PJy
75qH9Ty3NVPzNuy5nXSkeSRQEP5p2hjeSBDXL/xHOgISvXxscgYNA4yCrIMN+Meu
+CBiVJNMqadiZb6zNZbVRY4nB4lQbehZNd0cBvFSS14H07Xg05o/MVzLdrZHjqrD
Ij5hUTFqdLJS0IE528NTdcCTgHMXnRPsgT1opw9Q1lEzBkMq6qfSxp0Lzh9MUHyH
7i/IzyMIrEvVSz4XzP+eRur/eA4YZseZyYxZ0xBiDtNUPsEK6xIxCQHSz4IATYmD
SEsRbRsCs6WvCLfqLq4IzrzcNfibs6zaQbu3ChlzF3oK+RTFNZ7FnbrjWUlszc6+
eCxupqm7/lhWJ2MRoy+QZil4mxOxUBb6q9C7iyGuNLbTGlvdUoL/GRdq4Lgw5+No
1N2A7QFE4mgTnqLDMJvUcF0Dr/kznGX8bSiL73pGkvjAMosEGKkSSjSqKN5Q+5gC
gsgxVcy3jvJi1l0+4ogpudwOKtGs2UEiAFPXqwDCsCkoH43fGqUi5CpiEfnJymWD
NcLLRoh1jOtd+RDtKfx1et4MqRT4hf3yd9eCnok+sGcZmGH5Bx4svqjlyetddJRX
1N59lmn35RcnH8dVAobnKEP5dljKzKX20KllMrvkGWLE50SBm4j5vamsNioz+4B3
FmAsPeZG6jjSuCbjdNqkCNdb3ig/Ls/SJkekehfHg8qNbAi57Vs3p3e0z03wttER
WieCMxaiXLjkDKr88urvjkBPy6UY9WdNfdGFyl9Kh2QypMsiJ5y0EuSnwf8Ss7vA
bujPeEYLCJ5NPKaOrUFj7I4+ZtPoNhkCOZ/6SpSoymDWSLWB+6Co1iWIgsXHzE3Q
6cS5Io2OUr87XuluDeS8KuFXr+CnRpN3beeIvx4PGNIAGMdiYV+YeGyFb5ZZSq+T
mS+S1kXPTLGyl1SrmVwORnZg76Xq9XNeqxBjbuaBgiNP6Qc+kkbHAu76PCAKirzy
Ddg/TSxOrmFMJZ8VWMc4NlAvy3qvSCEmaH46wkTikmY4NNQrzWfxFijjvixI1Uiu
Z3jDpMPAdVr6RQuqNGHTtuAdb4gQ4hPyYgHS9AVVHVrByrX057JwTeVGxy7crYZy
9L8YSiifg7ht7OHkCxIMrCN5BXokh8P02cfEKBpDGb4rgZAVhpurrmueFglx4A8L
JKPz00vBS/FHTJoWZFaVaKM/g+mo6n7onSdOxWVshHGY/xno8I9KtuzN6tnPRMH6
kqReBcEn1C52Av0ecpVmT1b8J7zvOa/GaxCyLBYAFiZQyodqAAgPMy12YFBSFHXm
A8vQB1eNFRvMu+uOMi9TTDs+YuT4ARZxYxfM9I+tX5HPPm2Q1LsXs8xsGRVrci3C
viVz3csMa9tFSXzbCsWBD+TuzV2XFgS/eHGma9hybBvw5NJFu6MEeDvoMIWQgD8S
34EbrAfvLeizJVxxWKxGLaF9UZ/MFOtfR6PUpwr18erbGvYryK+YyDzAKtLdIX2K
BbLm4sKi3KrUu/0qIY5TW6vG5CBo58EYO3sUcixBCxpBaAtIrd764pH7O4xxQEoV
lApn3afOokOAJgJjUai91+onWNKX2zluROuX24dtN+OBIQXiVeQpu05zWcWXQ72P
9R979plLV7Pzw2VeMb+z3N/yMdzZL8TThywCgJhw00OEGOaGMT2M+aMcCwQsAMOZ
8UMVfHgwd0NE6ZZmdzfilQDnJBcKyWU/s0huddmQBzm8PMVmgRtPQP8CJzNr5on4
SpxBee2504/k/pZb4+i1RSFv3MhvE63Cu2FzS+27BYscnXxvwaiQXkK4Tt9g5Nhl
nscbW/AvX6DzldhfOGOB9Q6dyCMwYApeOvmz7fxMDy0Sg2+jssaKHel5PrpLP6O8
7/uWspuPdk9qxXDvH+melKzqYpSH2FauIGgvWAEpJ5SVOEpylQ1Z36qLqeTpynHu
/YJyPzOHBGUsYLPwj3J9zVi6t6vfvd14Ll8++M7r5ZmFTOEIMNydM0ynbwuJ5Onf
rW7v6C+kaHx27l9AyFYtMm0H3Xwjm0q80GuZpXJgmJIczuzDPZjieaZpUkZ5KsD5
fj2RY3ETaA3spyWO9vRb1Xg7CIMKlPLP4iQEGYWLAC9AduE+r73vYo2jQjxXax3Z
tfgXll7rs3JNFMgHRPFZG4Ceca+DBhg3tfAbqj17K3x0Yn8Pjb6jfafl4URRrTry
696Njjq9RUKSugsKJ9WuIfY2gQokdFhWSXPLGPh9VgxKt4wbDgX2tqpxZFhWwWZy
uESU012eGKamQJoL7mKKPqlA4819kNnWuu4DzGLgn5zBFUtLEArTdyoHdvj3ZPl0
RZ7/JM8Y+IGi6Mk2Wx28ndATOuIn+ZJOaeTgHfyp/jla7IaJIIWoH1WzSEq2tox9
NJUjhKUY07COTvMkwCWhQnmKzE4nO+eMKqvbC6SiqZv2Q6532AOoA/W9l74lUeoP
a7Xumj1OU6tcnFCpSvbm52ZUR9fRKUa4cyOdHt34zmhoVv8sJFrRCbwCPPzd+8+R
HZYnltkstH9xJr2gu9fQKvRj081OwGJE+5OOUB2o3D38/aKUUPkewONte37jKSeX
yEPnqpH9pt/agf5LyA+ntwvyVA+U+R2rFedMphwrrTIzOQ2w1Mtxa1mYmJxRUFdy
Gq/N6aAKNwrdA5tjP8vrED6+DPAtE9lBwJkaovvbbRC1g7s407w7H0s3wJNiX9V7
tEFUhMxOvswpm5QoFuLR9VcZrDRfXB4VVwC0YMTzttnoqWTRn3H/UHQsRyIcWX3F
3J2k2IdiIOpPMDLOagpvllALu4Pgsh/ai7F6m0VeumpfNSM78x2FZ0cG+jdeUBvP
vZh/bd38I1sK0zgJRCbcq0tV/ccq4CMfbmj/LwAbxS0o9Fqjjo6aRJ3SL29G87Ze
LV1a1TYl7Xl+j+OeSCdHkhgWIHfNXEvH9DnuZhucO/G4Ohyrn7AFY6tnq86Bsov1
zC63TlpVeLQrzph1rnNy/+Zwh0QXMzQYvouwzYkIpEWLU0cTnkmZ1YYNBzxVHE8f
kSdq78E0tZ4mwBDb2WOHOFapmWnkFlQNfhW8VxFeLLni2sntzlx4POWc8Rwcf8qf
/TptlrZJUDaG4aWisJcPlRkGFjlxO6fAMXnoySg23tIYLz7idSPa4FMJWnHzciTx
kUtSOCWJOje8gMduFqeuBGtDH7dxuTkOw1DgwjPwzKFvb2i0Zbr8D5HxowPdq6X+
VOK6n5BBSQderykllYJC4njXn+qvj36fq1I0dZxdUd94BSmfhB9PcQKi4Br0NqFS
GTjAythQ4qbQ7G2B+bp3k2cY0gMkcBgYswjiLJYS9D0CiHkXHFoGx3BzJJswMHlD
4aIWCdajePQqTa+KdVgyGVlc3dQwGSH/Rafl6PZLvrxrqcNfNxIsjKhrfYXxL4aj
HJe49LQ3n+84SIjdL19xDZ2Dq4px87TUET2dEqf/82eYDsO+9iDhMdu5eEZ09H7I
BYlbsrYWsvtl/N3Mq/nsQAVc3M9dKMH60cRV+Np98hT0SSuK3psw/nFkn40hFHMQ
4OO1KxNwhiAsIt8jOy7IIYunyZvCrC47MdfRFVIEMuqIVNZiLcS4wFIDBSVBSTOl
gSsVW8ljiAFILCMHomBOcZW4FmVjM1xVuEhzI37FC4DZ8t/Otwyqm0d55eR2Aqxd
XU/GYSnRgP691sUpj4QhGeQzfuooBmo7NIIcO+7UADz6NPiICO0Ywi7A/OYn3vSi
fd12oj+hZz5rvH+QJpkAkYD1efbvrz87gtliSK35XM+5UF+KzzGNZGnWq4ZnSOwt
Gjb0SrIFUdBATjAbdv+HN4vtCCYLJS0HTp64UhZllRTWKrtiG1dsRpzTj8kjMkyb
ycfGFY6BicgkzuBAoz60JtZCipHHVIYcd6huPVrQgNGpZFgVXfkVfb/7ZYagCulJ
QAAVak6/77LEP4y/4COxmzzF54x0uE0FghQgp4kDVmGvLM8mzCFtubPZGoTIucAF
05RRbbm/QjZQ2kOmPaXbKBIHW6dIpaiPmE19hgHj2enBO+OQs79ow1ZyRRGQIZlu
/dKU1nEJz/zXoxi9hMdK4cokN3yj+Gp48Ur0xEmKjbU0E6E1VUsYoSLuDcnZu5bR
fh5nCKrlFNk2oiPq5mOHUvEMDZ6f9DZKbARK0n53xSshI4cETzTAUNYDPXx9Ate8
CkFUgQxQ3ovFjgRDxsFCrpltAM1F2aeTvFygzInsHetdgvt2ZdZ7kbEvg1fdWQNV
l8dR3SMNn2kiIVTCXNdsL0wmhCX6TilWE/CiwSfL6mVIz71TR9idGpv6/nrQ7iCC
zGQq6hiHndUFgk2f2warHK4KqdtGtV1KUW5er/TawILDFFRfQjrx4TD5JsMCyRhT
pPsTduU7JRWyqv361vmJcn6nKyUTyaUOUPBgM95ZoDwU9j/pIhXCAvPS4ewuHpmB
qEKsH+irjs+sU6tWBoYY32O1MBozgmb3NCXtTIF8oi5iDWweuCt+zykIh7yUJ6sA
0PwyZinBBt0CVfwcC2qKFiowbYXysD0hlna4PGNR5B7GiBsttHgdtNv4uFo62+6T
SlPv/gIYfB2dKCeY6qkgQ6QBGYpUPaTW2nCBRVk+gjgbjCkf464jU2wMqNxiGMU3
oGr/EmXBB/A8zenz+38W+LReBf4jmlkR2swZif9+M78sRnR3OXZEajRG8FgSb3Ns
jjKGKUIvaUtnNN125NSsZGf8woSQmtOdhaoXN24GCDt+fxwFSwzB2Ppa91in0kLm
eLArO/bk0ab5Nr2kRzDBXaeD+8g8gSt2CnLoNGLPgAB9CjgMFcdPDJs/FpKbbvnF
wW0FGLiYp9l7czYijpB2sA/Ut9RUwX5OWEoRTGdrqOjU2lQ0TKHXwxvvj1O3OD7h
AjDYay5GlPXXoldjqQSjV9zfs/DXEdTFp0DcsGXIPM0VtGpBO1aIv5TYWJtrrvL5
HFGFUO/VSEyYAD8k5+SKZ0Gr6NAHxmiTkUePGhlQa2BvfvQQrKeYc8qHnFQHTO4s
nPptvpjSusrFLhCGbIo/D+xN7AayKRwALD675BK//sg/ih1AK5ssXST88lwsTs2g
ySo9CeFV1H+m7npEiZe5SyQ3fXUlB0BXmwZR4qqTgLYxVBRiSbAKL9X1ZTOEv+zs
unehz75dkV5YJH+CBz8VpS0GPOnnxXjpvAVebLssVmaa5BEJNaOYoTNUIlr/ujFu
tJc9QjWmw/YA1UDfFmvGq7UJEqu3dDoiwcSKJzv3Sb1jaDktD9auMVpQ45Xv85II
p0vVpzot0iRRbxI1z488XJyi7SqIlM/qZ9zyQwO/CJLcOrEvW1rJG4Ba+spvJvQ7
d8NJ3+E+AQgxyzCaetFxO9/79EwLqjobsUgEUuGlH4FFD0WkPKWUk2IOivyrPZkY
SKlSF3/s3AX7D1G7pUct1gG8gpCZePfmedDWp6zuCsEIFFwz7rARNCMd0qt2KMOH
aF+EuSUwrd/4FoIhrYHnqDleg2Rju0hyElG/pY4TNr/StGiKRSE8DEclTcPIG55r
RHnX+Pwb5M3PJ5T1W1EQ/jI3UJJoErtaPkraXMkN8l3I00X5hZ0LgdDu/V8x1oaa
Nfo7gKb3+my6Z+PWGDE90+RdQRA3/keM+7dN5GHF6B3Z/aEc0qa8s05e/k1MSAri
V4uoIWNGLoGbMDlJVDQwZEz90oWVJUfzoFywC7Vv06G82NQkILVG/UeOueNLVkhv
mz3BoIbKNWZV3ikD2S9WujJ6pTbdEJ/5mn218fvYUbETpnieYhe/QjdJYjkLss4e
iQpvAHFNlN6NQYvCjlCsu8lpZ9V9w06T677581Icg36b3ntLfWpqbKKPm/YRNSmG
liSM3G+++9IZjadOBlsTpAcKK+0RYAw0dxiqUg790Rs9PDu97KnqK0Hxf7WwY6vv
+9paO4I2FwSwes57sZW9nq67YMr7xu+GmFscsQiiTFtHFWPpcaYBE7IXR4BdkNr2
6J59eIH/78QNmBMjWb0f0PjckyNh8TiJjJ3dNbMR7Sh5477qZq5zZnsE2Gus0d64
EnT4DZ5sZdDBbXhPV6lQ6mZRV+7Jy6084fwD7FCeB6+45qtX2/U0Of6bRhwwTDz2
VG74gL8DJcK9peViyaVcrgtNzG9kIu2yLujclv7BaoXxlwBCh5DnFIpSIhk+VLG4
hjSxYP6+ntW8IYChZMxhmEUvk/Wm4fG6XGf3iwUk7lQNy1UP3CeUtyXzx6Z509/E
biWH5gcpJeNmtcMHV8ZqtLEK99g3AfmVjPO5WEmmbZjDttH4KKEJ+DawnO+I6Xa5
3a9ZKDf7kH9a+yct34Xyr2q+Ew9YziBosXtCxLMlZ+sBQvsjojMnaXTRVgs2LiM6
vVw2pNQhG0EXe/ATuEcf/RGITMLOIsfyBhBpRVf0Azo0ZLVVCPwJBFNIRxxbLMvc
RYRJIz1I5nry4PfwGEOr0sh1wMRMEDM2oiEw1yhKYIeesisgC7RES5Lp/lOI1fBb
/cUzCfUaerIyJUQfokeOYz64WWjhacVO6fjk/33DPfobT0pGod/5zLTv5dbB45ow
EoPPZRIVE006ZsiJ6m6yaAMe8WgXy7bsvI3oOM55Md1imFepw45Jlt7VE2DcFHuw
8/vbrb8QC7TPjhTRZU+4Vuc0ei0yiR+fnDNbi6l/PYWwfWEtLLPYAGLmRTyVfJg8
mWYsFBm0RSh+1zybXowOiu+RXSgNkPue9Vq32ZuFSaVEx3xaCURXVGqPq8ozIn9f
fUnF9pUJq1KE6lByjk/2BbmeLwrqjIPypQAx/Asrs/qodO7oMgspECAg5D511YPX
m/3IaCIHawApWXhDnkIkyWm+oaFrnBlEoV7u5ZXn6KhjiHKscd75AVps0xBRxjqK
It2pmdh3dCodErgLdBOatW05gcMQ7drGpWcTFv3nceIP/UW0oFJiz7m9/nYl/Fcl
bRQTzP7Fq7pIpQFlmrLzDeeq5E3NdWnvwbS79StXr/vC3hwgveg6w0lRpcFAUyfe
Ky9VFzB/ZnPHLWHZHS9cXVR7eUcX7vd5iMdSexga7NsCQuMiduO1wQkVbqJyiq2A
q45TYupLz4LczCoa3/RmvpqLO/Hl/gyEUs0RY+LVxi7rSI4gMi4MbnBKFfvSI8Ec
a7ff1RV/g8mHTOCz/qfA6bxIov4zMitXGjKiDCBrlrxN6BrvqZ+ky9rzqvCWz8o9
eAIo+ANTaRBDRzvBMHlam+WGLk5BwIhyve1/fC5O/8uQDrhivzBn2jBew64cKMgm
hDNBjeil0WCir8NtJdrgEEjY0ebyywSj7XpSak8oZ3lvtiTBi1wlKT7P9/fvuspp
LHkGP8/Ei6LxIa56g10FkPCjR0FPhyjQkQQiLH0TL2DJYx2jhQB+rmj2XPAeGhsc
FtIiT3EhLvzMQqHX9fO8/Yv/5c9g+GW81P5dXYm4XZ0cx2CHTmCTXJR32pRJGsi/
f1bPKnwnDj6T0AlNfAtkTErpUrhei7E2tteoSResYiY0f4NsWyS10wibu3Z8ORLI
EVoaxi+vBwXOdZEyidw/fX40Rfm41YkU7dGU+YXbeM7D0kXKXPGv8wdg1eL3xr3K
qHS14UzFWXbcDVp9aBVEt/UNPULF4KoU5ZC78G5OYrhRAdPrH9sis0wNC9JHrHKC
vDrrPHgMHUXOp3CV+dtGGiHJU9+2otIMNU1z5DCGOX9+/FxI3oemcZtPu01xOYwl
/7gYcKKshbQoMKT9Ph2Yc3c1vYtJMtno37lRTo4fgbArH1KzK4Rqf3IPOujp7511
PJi8X9Y64rPkdBgHxXEZIv/jrpzJvGnpm2L8h1D1c/ozvax7iZi5DDGzKUHY1k/P
1tc/r4xg8BsCy43Vphtco+0M515A1v1d+BakIF7qJ4tvxLXQIPv4KvoM9QHtXX5F
SMa67xU7JeTG44iW4pU2/K9/1JtMjTcIArQdST2b4GUbox+x/0nErBuEGGD38a6Q
vFuYIThcmivPZpun9WtbPAYuwalp9dH1Bg21naedbNPtk/BcIeXEPrzpF1Bwayzk
/FF205l+5/1m1VMUmkSLXW1ldq2EhstH2LeYDbuP03tvBYQ0GerRih4buFMs79eW
E1sGZUeFtXnYX8gLLMgs0aTuPm2l5pYmV559sHenJu0kC0xuBQ2vOOc/vPHt1Vvg
6ePD4PCb5pEvrXLsv9dxb1Z/98c0GO9JaanhO+4pOTxqoo87S2QvvUPTK7qkG4vk
7kr/ek+ojisYs0D1dP4be9G2amcP+z+CiNbx4TfOyszDVhrs1nxg2kLQh1qjAgav
v2CJCeHpXYFo7zQ1a8AgeOsaEI20dXdmt74gPzflvNB2T87hUR0rHFlPTKe1hF1e
jhCBFAvlD9QDuNsELz0Yo8AlwQm9mL+/qNBdftqMej6OuCZUVA6cBifu/McKKjz/
qaSpXpzKSkh93emUirR3G7h48Lh9lH1c2c1BA+BCmHGvRuld3YChdSLx30rHNtpB
CSdkvdVjd9BtBaLfJuo2lpY2aBOKGvrLf6oNklguSmPa6CPIEjunrdQ+hRH+5O91
EhALjzZ6+CtNBFkJl1eYlroPlObZq6cNaiZy/FnSqrVlfMoipHOD8LocX8650EDh
gA9W8PQzo082BrwKCBW94ez4S1nS1Ie8jkXOBeg+MSwRJugV9bgrTvEjXSYdp24b
SmyrnWxUXNvaqSNZIodJCo6YrNXhp4f0iSD13vtQL0xQ9BNpk4ZynoVijjIyWBIV
JgsWOjYz/AGgEbZeqrCl8nUTlaEZWxI5rIoJPAbi1nd4AC1d0V2tT5JbjDxuJBau
ehVSAw2fNuOMFv8wRAtQ+66cq8rkJ3EkS+i/31fU/kWPAT1XATYpJEV+srHuTq/d
1EEWwFKPcSl8Xadr5nUmhMb/6UyCmP7Rn2R2psS9vMeWY4p7UY30ITFn29Yxw34C
dYWymV0DzlrvZKm7rDbBnkefAKTGEtqXowxRx3MKTn4yTsVFz6mf9C+YMdojiVwL
O2SxqYy/r///IVrJiOOTgbtAlf2ZVLq5rUUQuvtXeDmQmrn1Ar+/aJKAtWu7+1/H
kt09QAHmfMzLeOdWUwBnPrG5mOR8k0tq1QpNqfQM2+ADxJDLBB+j3xs0iOWq1BA9
tqxJKVyRhn/GgSptONhiGJSaHcJDETU3zcpGsW7dURzc/a9pglmhSmz/ngtbduq0
amrsypGW5RddXzSTwMGnu1tMLLlS4wxKzgAXnGN7Bre5NgEKTnveDbAYRGqJrVCz
pg0+eQ5e6S+CZQZMnOfY4DEcZ6RqtwOD5U5JCdNfN0Ct4Hodz9LozqjUJaB/+zMV
pmI217Gmye8Rb1otvQjLrjzRygyi6EGIql/D++uACuhLVAJ9CbOFvqhB/uUHz3BU
+Al1qa5Cvc3FQLOP//+Kcxvm/rOsfj5iCU+93CFOmdCGgQemnSoa5zNZjgq71DA7
ykBd8JnpA0EhUsl6KrIkLPvoe5EVVi6yIHvtLH281jqtSD94CNri3r6n3uDIfQEW
8GE/o1InCh23813VuoQ2xi0Bncz7GS9agn4fohJQ66EGJUbFFZ/47P7GjknhJy1L
tfIVKSX+I4jTuK578C642TpQcw+6Lh4fd7tdC3RLT6V+iCkHv6Tz5ThvbSIFPKBc
baT3qg0oYrnKMNUs7zgGGQzzNuphxetZYPSk3tJc54MwWu2s9nmpwza5a4on7FQ4
OfAgAAT7DZ0QyDDySuBRKyYryMq04jCAfOCak36MqNryhvq8wRMlYtIbcj6RoBgB
MZoZPHgmOBjt6pGGcaIJr/zMuoYRXuqRjUAnlHYfjCzCLC81aR583WrLM4HCOFY6
kR4vITWJ0HhunQGzbkkPpssv1+A0DIwdd4ZOmE/asYPZHFet5hmHGjHKW7kgMcpr
Fx5p0fQjSJJdv8XYOiW3OlxxfpJ44FBibhIdWacUOMaiuVgCdf0O/VHcr9o7s4Xd
YwtVUujz2YD8m0VkQbtFmjypBbVllKdHQoT0mJbUILKIiDKSc4+m59gmEmSUDF2E
jJWCnD0E4+HYT29PPDrzVNPuchwKdvvg/As87tamxFXUixVnsMO+oEnfF2o4S1nc
J0xtguEGbF/RRG/jTIso/HGqTIXPi4u5JVH8jFTTwDWNYSiQ9mw9z4D96IU5GyQf
lnvcn1+/gPIEY4dq+c4rPlih/y2oYZQGF/ZhcM0PIfBu9JvjAyx2ZBKIsnB4PxTP
sViEEiZvrr6i5JbU2TGMv6k6fwSgvm5ggnRIFOgMVGmDpmF/+4oKNs9/s9VDyg/B
FNFuxkLsmKIs2ZFnczhVYHtaRhvC+TfVuXfyChtinNlbPIlq8937PVB3nVdqrvjd
OieMpihtiy+gC3chIpNgTudur7qRdtVoZyWXgV1qGjkjy4zat+Jzwk+28A4GdwX1
N+0ipd4srShdtdIBUqXG6OHwsvulaBSL8JDbzycYU+n0+oLNJymrEyWiiv4I8n4+
NybxU7CMG5GyeigmXNU1weO4uXhRBK7IsTwPmyBMD/zIHeRTaHBoWobSIIv53eK+
8HOEQD50XVOs9pb2SGd0y+RkZT2XPxaLM81yzgu+tWMBnfvwikF4ldVQ8zb1xcGW
CEuPnvvdOfPbpEZZfyk5c6i1YO0gy5V2wZhp/ybx+cVwp2EM7Vz8zsKahrhLOp+N
joUXXF8s604vEbBC7zBJtX05D3p3m+l7BnT//kYTCt7t8Iru8qPrsA9YFRnQyWp0
JQvF1BJgA22xIL93KmJP4SKwyMpFsrBmCKoS9g+P5CiuD8tHhMUGu49rXPr56Hdk
AhFoT9E0TKyXelW8+qATrXBNvwkzOGq/jDjUvMPtvmuRrN8RW6SKVUEhvlJTQOCB
nCXeztWZM4YvmnePEAZSLg90tz6F8b8yXGQigOXhXqEmrP4XRZzH54bNGp5SHJVq
Ww/FdfBOks69rAoqhKoE5Ne+nY0giBEZbCoxOcVoM0agA6Z9XqgKs3zPkDsINjEL
m89x+5d06K8VBcQsyY4tAAQxf1EARDm8ba1TWr9oksGfYJJce7g0iuv/vQHdFQr/
I2lEDX+SAawFpA7IykzVFR3RwN4ywP/FuFYrTs2o7IHqClwMFbOv9d6tdbTGdR/G
cJ5rqw2UJpPYWwsG2cxdM93DiDaYEQYfw9gl0HDvsj4a7Nb2IWKSbgwhp+G7LDEl
6hsoY1jKurTvhwTSjUbVodI9W7xxCcMqedeJNTIWJvr9lhA9okXRIwsw+NRWd/7c
isitwH2x/9bfsdsu6pCtEAyjhe9AKdmpICe5Zu0Jex5L6gwouuuO932l7HJhI6F/
eQZJZRCFMRQwBo/DxRsiIgqvrYowVhJ0oWfUfR3RyyUekIOq2gGK4VW/SyuSPIPR
wtp+x2MNikC/9wXhgbv55KQ5wce+AoFcw31tlZBya5q61/nQu0W3DJwtifiYaWbb
uw5CWoeDLoyegMNzmW1n5GZ6fuP19M3lV3xf1m9TbnDxjMKEasbmZLh8rz5FOIfV
fELYQfVOD9QGYwoMZ8fBq+G+wjC8COoFvhXnxo4L4NGFHlFc6wXxLsuPy7o2jETl
s03VVlS6Un1xQxp6xvmUtzq46/ZEsYKcF7mc3zkfqMWIyfENjaKLzrVMY3WBkC5V
ecMJoggXbXsLiUnFUUEpr10yc6cb01kCdqo6El+wPIGQ4HdSwULDK5VT7YMMT+c3
bfQBHqToDym7CmjLbpGWKqaiwjwGy/VSRlssbDNBK5yY7txaX+7yHcq7a/DBf50p
6FONxsUotv6Ouq5obwTL/tYvFDZSl3jLDYEd6g3Ia2eOgR/6l/TeCo3QY7VNr5Ht
c03Y2gO5TV51n1WOPoIFoZ6cY1zH+FfrNON2MGnWRb9RYtY8eidU78RqyPcABRBo
gk62XqJ1DeYnwNW3hMsTB8aQcsM43nkBNOw3k4Cm/FS9n7sjdFTslwhBj+7MzNAM
Sk2S3tBsQ6OnMncz25q+BZfAJg/w4EqDbJMQILGoeBbHI2/ysLglU+xljklcpcjh
C5fxEab9RxiPygjqXuXlI7qvC1L6UxCbOUHQWRgz8LTXs9HH2bWR+saGihIbbPiL
iAoXuRXaVrbM/k/jYusxoIUKYPiz/6QQ4ItbZpPSuJSBbYojYr8sNDvqGDU4jROX
4Dgku1NAEtw16YHoVT1hEkv1GtjEq0tNWYNjtpp9921FjopAxHABU7vRUIOL3LE9
7/tTv5g1g2Zcl0rkcl69WH9yTHw5KEYf/LD+bs1U6ojOMFsVZPvMuN9x2buE6cjX
X+5wnwVNzXEy50LVNwcr9HMj/hCKMM84E5Mfz3ZdO/VKynKFdiI1vQoXLzGucRlV
B7sL7c8Jejfsu+8WP2QP21x3YtIV7t3dzuC6sgT/VFDWYBqNt8pBU2lRuMqVZJCL
f4AV+o8/VJr2kMdgaRBZhY7k5T5kKIqZk16KPVaz3CtF7Y7O8ZD2hz7Fluc0nwpG
HVQhZ6zOw2VHfy7B1PFl/dIwKO7X0lOnHwj66utXMa1Vasx+jHCGOuMMbYgRKV7V
vHjsNU8K4wdzMYuQtTUjqZn9VcQvOG0t8tOYXr6abOW3sdtpUtknl+X2nXiTM2hA
tJxS1Bd5bkz8AzlpNV7gSSdcV4dMvbvyyrjiaPx4xINx9n5JCYX0APYjNkmELGt+
vhBfml6ib53o/siaC6+EpldmoTBKY8MduEnmrXjzZsJ+0l4t6EhjnXkaDlqQw6UH
9Cy0KWERMICcyGlRR7zTrDeAZNEK636zfbjtu5cQXg6aAEFs/dvey7Me8CU48QDI
73q/3Nzs1iCDcPX091SgLbRpGa0ShkqB+zHoExXhuGlnE7EWahkAWcmkVfrdoTzK
CE5lDRDTEpzUD4HzjG1Pe0B85Tf+6iAfOFkySnw/g7XPA2Hy6BkW2VM48AAV2B0Z
RcaJaaeWfE0tEDTBvIggmNRXMqtxfb0fF2/DaeLKpIEC1lJY3spC8n+E/fBQIuVq
4abaOIpDrtTI94StPaTRaYl5/rO3QoOYDMwpH8foiPslPf40uAHaOzjeBOgcKZs8
Yz5yF45V2i5AEoPWuV5J0JPLEGshI7vAklbuvPiRcp2GgmG1uU/ZGGSJyGyzeGFY
qfXg7N0sTWgWxa/YTkbEENHnwwdrmvrQYAxXxinePRNG3sOCcC8FkhokeDoYfOik
bFv16V9V3GZCc6tZI8A5oigzDFAkzGQYv+ilVbk+z8ZcIAN78TGrzb8SpFelkL0N
mhBO/RySAFVUbIqRq2S7Rx4WXPoPRbVitI6XVuhu8FQuWRdRufztVPXB4rimrjO7
GdIWN/er1n7W92zHieyMYrd67PHgn6oFbAiMlj6th887x9YozV49vcQLls2fCc4P
uI+Y2nneev4c5wmbg+Xs2zSQ5mYxmr/C9mWb2r4Ve4Wp0JmVNhsWaBG0qwjEi7l4
+d0q5aIom+a/4eU2h2OyzBLEiLjd1zNd4S2xyMY/APepvejP3TaJOIPgZxfzdWel
ItQJCtREZQsos60JH1PaSbZZ9AvXjwJ39iPL8S9B2A9IbnQMPMS8ff001Ub5err0
ZyAxFjbnY7W7vjpjzlqC2cUUt+BQycqjjR6fyScJLjnXRQkkm1DWUZ9YG729Hfma
ElHc7KxrGK4mZxlbJhaGGmfBxnKJmC7hnxqJpCuttLlYEF9jdfDPTZwm/8EJR1oV
+BRAF7BSiGA0qTdxvE0XuJcz6lMOgt9J2mEeEHljGxfA6n3EhuNxrErz8FfeFbov
wHSUKtlC/A58RXD5gEWECy1uZ/fqqPPixqoV+ycgn7GnVoWyxbsRMYF6l3J81LNk
lIgpRt75k3hsJK6uFJ4hhmk96LapE/ImOJw5GY82p0GYQqFcq7Xq/BPNq/uxMWmH
SXfGIILGs6FeadvuruuOPM0xdK411jl7MwkGDnvpRwDu5ivv5FwovOqkXBF9oz0U
FsCSwipT9mVTIwijQa9MowBZusuzT5KISA0A+2Klr8tG7RRd27eM9bRqPtAxJgE0
EbqnV23EerKAb3vCxec0rngIhrrmI0+8nwAt/SWhE71KUFBC4LFf7uFKrrHsKrUU
1O1t0sBGMr+AWo8qYyDSqT8gU97pr96vgfUVqs/AF5m48hPP+sXVghij82H65OEe
GcbU8sJZrCvSEAiSrpnDWzewmmi6W4u6q06uNvPmR0oKZ93HtMOHSTRiJT3Zay1u
BOK/SEpjQrsXrL9/MccaXKWngvJHPKkkuWppp5SbZ2ZyGHRmfK2YtfsAZFqWZn70
pWgUfpkjNFH/g/gJ/d/h58b3+uQYk+3s+GOiCniW7q63KKP9LiGUyQbi7YV8RQm/
gDzkb0UsFKCBP8EJ/+bT8j4pFUXhBhWDfhkly9Dx5IywbGh67lsK+cO5t6Ljy2iL
BPAJC3nKRH7bD4C0NMKcgwOK28Yiu0RpWBJebDNL1vLWLac47YxYmWZvf9al3B5g
TpH56l4+tflqOlLJBZ4+6sR5UyVnMeIk9Rw+Bk5IvlA++2jxTLLzxvaLVyXLAQ+G
eAVK+p/M3SXPezqz4Uz4i5PDSr26tDoU5zrxtXYtYP2Q0KNFv6s7dB4m/2FHQ8N5
lr7UjpRTroYhUiE9FhuNHyQAc2LFQsISuNJzvn718tFmEoc4XKENbX+XORB1+C3E
o/bldZv6nYzSoi/W5xlqgegC5LdPsp+65OgKl7lIsJ6i98FL2/zJM1XzUVmIiJDV
qayXPL8M2KsLY/k8ItxdtI+Zm7bSdls7/b1Y5fczd+CEKiO4qQcVZdvYPN39k+xc
IqEgNVkmHTyb1igdsE8AkdtWBFzJT8GBQala3pw5kdJdTl/aoVbqO0z5VsTTgnSD
ItqyRA+nFZ8pY5KN+ENKPda4wQ0ZqENH3y2o6Q9bZgcy1OezGqWl0iQWBFJD0TQc
jn83/oRtoY/NCmI4CH3yV0xY3Dn5uz0brQNY0yOsaj+h2ZXBgA3mYo0jN42Xtkb+
wHqRlJaJ41SPicaB/GK681vzjKhyu884T7UWPq0bBlmNClht8+f3JRNAs9s2NYik
F09ECcuF0Xdkszb5MuL8W5Gq9AqAdL1Lru4cKe1pcbHCHAJvc5i+JTDBkhHAKgXo
2CfA1r1jU6dTMop7dqYWt8z7ze7sMZmlJv6LBystn1gtFLqf0cEe+iJ2RCRsi1fJ
jEIYSZtEpvqTq8r7vPt1wYeLkn5idaLU7c01qKXMQOy10Nr08hJ4fAajMsgglBc3
qoEYUK5KmaqprwNEDuGfCHLbdvd7oLfNGi2NXfqkw0j28f/hA94F03iu4jNLmmip
3RWzYHEHBgt6+Sje4+UJ6KtPkj+UL5AuEdyqwgrWpsEakLvfhd3Nv8yZUUCzGMEy
93FI8ffL8Y7I2gzTvWM/7rRvm+GQIaxJ/ZLQ5Xkek9eHIs4bnKhHKxcSN9mtMc2v
n0PFi/d8afxIq0VJZLQnvBhUQxIT5nZWrXYVL6/1PpFiot0Di/alJ3PhUCnIz6fC
qsr+rUez6oGIEhUvWZfl9xkXFZGCBd3hXX2ubHrfWhZlW1JKPno0jAPJj7e3zaUc
Xwm6oBfApJbEdXEei/9vPZCnuZCf0lqmLFAea9AvJrtKwWqEcQXETk1LEc4dA4YP
eDyIHcS2ftsmF/4vrya6pgt9z8+oCsMobHIgh9Sd+UnpcXvtWH0eNGDbIRo9SN+S
SUEH4dw8AN/oEFRupgyMDEiboa7T79JOGbSMXspUW7qJGs5NstkUGB6ppzgUaIRZ
5LUEX7UELgf8tib03vESql0VsoP5K41Io4dGTNlcfb715+Tc8/N6dfAWcPGAs6sY
9U36lAY+o2dKDWCGRsqVWBHkGu639khSOw1bsigM+IZs28aaavRQaR/aGKg1NldF
D8rP4X1aI8otLJubrxs9sN73HT2RY44CLB1SKzDchkjpynVEzYzk4lQPjYGiMJp3
PQTWJE9Jm9a6tO2gRHYGfhk+bWJqYmTSwax07/gjB+Xltl4zKQooa4sz/1Cnf6dm
fsexNidJuoVMYnrhcFmHXXdNgTRLSIDzk3KNtpVm5YWKMNLEmPXmMGaHDI2NSdSZ
AkuSUmuoi+uAtjflC76NmIHUN1bbfpfs8esucGEIa4QvhkumrRfKGIIxpV32im5n
YtqTMj8hTJ8jxp3tia/M2HMBxPYi1OrgGajq5gUH993psX0ZnzU4PyCAgAvsu9xu
QOvL2meq7I90F1BOremYy5p3cgOCOG3pCpA+wYHuZotcZCwHzkdOJSQeI2t5jDds
Gy5gzX8Xz9Bdwv0mz0KQPQuxN7jIlW/e5kdnOl06+VU5K6ZglZXARr5wbSBibpjD
8E3BuhvAdMUyot6oxrZJRZStL04ZNFABbKEd+zsjzIlqaWEjSY0ZT7eTWVcV51D0
d4Q2P+IK2KYJhAmIXtnqAxX19W7B314KzZxksnBJIeSQ5gJjaHTyBtPw1/Io5Uz9
05HeNUS0xhqwN1Kj3+QooO6UXwxA+pa0UaOaQci9wPxwItCckcKIX/YFAeojcKXQ
ZwUTsok5bVqnnIH39aiPyfLsAz8kSadAQakj+ee9cYErpDRqE9io0jvaxUTClKQw
Uk6hVOYDx94nKvHlVcL9T4TkCtChsh4+I1SrrUV0VmuSozm1sTe1XZT+oRsiE6cR
yVltkRBgcsh8codUThu78Nu3DpDrfkxqPSWxMVn7gXS3p3Po3lpmJFNHbyVcqSaD
Y5SoZSC+HZd9DPTuh1HFllEsKMOZpLa9ZhFFqE8SmQUOOvv31rzRZUyVCHq3UxQ/
FLpKmYfnH8vFSGeg5cYl6Xj6hpMikKX/GhA26qx/K1Z9hqoI2RTy0pf58nafWcKU
Y+euCc0GQLZUi7kjUIpLADTiF9MqOi4FGntc+bJAa11ctfQNby4268YFppriucS9
zfjj1kF2CPl2Be1NHtVKiB3K890RlWPpjynQ69eenXDmRUWuywLhdcsS3nriO99v
VF/bgCIVeJxA8wn0/elB8Y4U+SEiwHJTUWndWYBNaKhOG+yWINB252pOlSE3iQNl
muS9DWS7fy5zINI7IndHnWbHPtnpxQxKOR9JaI1hYiQlsO04XhY7t9ozhQmAOnLY
NPaEIWvKU33UJdBOxo8kU7y1H9t4o/8uDiTZojYSMW745pc9Lu0wDL/Z86gyh9lq
HbEDSXYc3hI0gD+/F3N7VH1ICIsVjUy7zI6I3Cuce2mdykmIxfkWLH3GXidlGgtq
mYE9UowrLHkwaJ/ha/5XQgneDI+kQnN6oZ3bfn2ijvIadU6F6PIJylnn7uicXWzz
DwGAKRVFpUs8tQ0Kmegh9OB0s59WPgnUDXBLT7IL+CnFXVl1lTlPZwp+O2mXLTwR
+3+ZvVceKHYE+q9H6vURimQCboyPeEVNPxGRxAiqYWWg32YwfUE23RHw+j4iAF3s
ZXIb+hTXLe1z5VpFWv8ChMYEjp63g0PbA8yraFADi036Hb2nCgNd/IqWAgHRLe8b
ac/xksv+UvD6utA3pK6MPxV6PQgrfifUhINXSF1aSiJ1CJTahrkDmoizgv5mJX27
bqB+r93MMfUvEalbwGZ7ry9KSHDFif7eUC8tjMN+qHs1+4UNep4mi3ZXGZGrNerA
IBIdiwx3Gsd4X1aBoh0pMvbbNaMMotZQjsE1C0J9DfRpfOSFMqBt8iNLEnXP+Mcj
bMvXB6HYgIXdXw+8IIqIvBDUeYGq4M6E5CgEewOWjupzzXZ1acZ6jS5QWm1foUkv
LSmcJbiZLtnCsIsN5FIU05n7Pox0yR2LQGqtNFvSEVzeFg9CLvsA2LeWO/DAMedP
u7C56ydTq+7mj0M6GSsLdxGXZCZl5R/P81aeZgEA7BGxHnSt1exzQC3FaH2drLvg
QlQo46Mho3IUdXH2ZeAVEh1mG3MR55+w1KY3OsVXRA0Hbt/7SQa6JQR7cE6e14lz
poRPbGY9D9MLtuiadlJ4oioNSORE1nWGbQIiGTqKsybZe8YdF1ML3M8aFE+KjROm
vjENLAVvHyrj4JVfKENyXbWGls1LWVwg+OoxX/ZACiClY/hLX+Ho5y5FoHeua19m
c4wsXlL5+4MRF9L4PAjM/X2M8CQA+qnpdpU/6B0JBDSn0fz8cfg2OaEczFdNF3Rn
E/cUkFm74MBVcg9HBWTgNxOHNot9rw+1mOWGlPrIiaCR1BMJ4JLE7h0E0tEn3O1J
/o9ZVzr+pgHYCwt1SvtIUTXA3+UGOcwXC9HE3ZibtwjKDkGlRzcKVR89ZJjM45YA
BUUDUaeExdhNb/520jIZUhj1a/aaurBO9GO3c8OP7TIGn8CDmVwSusilVQuueluA
d7E5U4zDp9aXqv4uureiTXrEl/zOXEN4gDTd5a+XWt+5r/6Hu6/4Cq/+5dLu+EVm
jXtojDeCL2qeT41Z8JK6mTp8ori9lqbL0fofa3tOlhpdlyGEXzlg+bdMJu3H5WSb
7rJK4o5UwgN9niycxj8sTpRHwCGZkesYgTdT5+trtiYz/5D/S2NDQ8l1xNYbwza4
SSlFtESqyM84Z8730oa6HtaO0vZkqavRjmO1XXCAs3swxZu5KNWfmdlU+7x4qs3w
166tLqJ2vRt3DG+ZXna+Jh2GUjUODh8pTUpiIzcX/nXCkYDEcsXlzK2KiP+Etc65
XOLJel5T0mkL64ZlBdFZ+BEtK9CY/9lk+0BO7T5GmRp6C1ce3FxO17jLO3TuN2fD
x+Lp/IcJfmRhpEqfOqw4r6c041+gFdK5pHnAUHcCfE3ANroShvLcMs5eAx3BE6Rv
9i5rj3UiazN1Hs2bsT1p0sbRHczWeadv8z+hUXCXi/3qN/3VTxctwjqBHnjAqThh
3XVCyHALrkwY8kp94FY+3/cPA2MZyRbV0txqJNNr6VtMMo5+eAZx+XRkw/DU4OAR
TYzHFZ7JGAJrLYn1NA14apnNstFQuiKgyyfpGyhH4/fzBI5TqR+MN2wAhUDTYHNX
CgAerGESvnj1Wsfstz+Zl2NhgRr3D32Fst6BZL5/HaKQ/tibnuBwqtm6p4pb6DDn
5sD+rVtVrknIrIJc/BZHQgGUCoeFXRhvm9/70vPit+Oy3Ah0sEr6JNPKml3xZLym
URO1MLdbaUJ6xSCIEx7dWFQRIc+yYLQwhLnPEjLeRy60kcA12BBwRwWxYISyQt+Q
19touqVUFJnjxKTJoBnbLdbOGhJmHkF6gCWK/JtUizAJLYJoPDHtg3Xk2X+At5O0
G5Mbl5x0PA8h0Qj6bUV8zsYsmHu6ZOChs5TDuuIw4srSqpOvCnBZbikB1SfToki7
Ukm8dqapaAJe+9pUfndwLxPk22EvHexjZ5yEuLFmipZQQGPqo/nR+yOMVH8ZcW4z
qNGy/yMmc4VhwgbzCZ0hWai+JaBQb4IsVeaU1EeSyNjal2jHILklDxl/lTjrsz3b
NeDA8TLokDa2V4tPqZ/qZ/LSzNUqgctmnUXTTyXCQMGZiuRSIVIcl3v/BGK96dFE
7yfMJXu1YfluOqJ1/QyOfPIYJxv19FokWXAV2ZL6c4t+4TuIP3tTZRVnXnMg6sTZ
ZbcGNfbO/g3RnlsgquneSI9HOAM3FhRwZoJv/de2eaxtu0O4nNtFOhrg9038yRMT
7QZ9v9chYrNGRYIP8KvSd/Sk6/W3IVcOH7ch/vJjStXgwsvk6Vz0YpPjxSuNC850
kds8uWAvDaZ5KoH40hVTXNUmYefqYjH0iWY7YvvI4e9LdPF4e/QTK2hWKEGgJLsa
c4jA6ZU/e55H9lKLAVm2FexDtEt9kJVUBqkImbFOpqekeVvSPMiLN7IETHTaxKOE
Lt+L2soq3AR8/fytJ734ieOsVzuxh2+RTh0UcNjq3VAf+RrOHw+DLonp8vXqiJd0
7FlDBa1eSdrA5xvmisyFI1Hw0KRaA3I1wK1Yi+xqUhk8njhnmCWUukrVyhMrxmox
OUClcpSNS4xcmjd6fE+git0bzbHVe8f1rc0oYd83B844TZEk4whXBImN5bhifYT8
OkaUzQzFnqZXX0+OSuW8XQ0XIgXvJRJRnQSfxdtYZjzwkAU/p4KVbZIdrYbHos44
dQkDQG96fv3n1H/qQY6k+KDTwD77qFOgoDyOdPFuHt0QTq3YY0EzBNUcBM0LtkH2
Bray9TxG5oR+AzIyxiGJpEzpnm+M5P3/LqNP5gf+nZnPTKiVMsHmAh4Lgs7dztp2
MwecpBL0z7y/B1yIIW7kc7v30yzThK/kKUyOrY2tM0eHisJ1j/CC7/2zHCb9cIDd
ir7xW91MX2RFuzy6HKR4vIVYi0aLxvgf0aAmUVpfBmfDwp7+LSEKCEa7ojdqBXoT
0ldxP7KDUOzjvZhTZ7Vr+DZ1AaICSV30HVXcInJRKHs71jQvK0DoE/vPM51GvPnu
rigowF/++QLWIwB1waKuZCrJCaXJISTrgwg4mEmNV0sAJdpQv9V1J7CkJF3WDb0w
ZV5+fJHWC1gQOfMJW5kbQeZ9dA0ZhNFrXZCTDy5mPZMNwyipZlyhsylqBmLcC1xS
idNNnM1rCZLA8IofYmjwTMzPhGD5bFAepInzE1lH35+aZRZDosix+qSX++4UvCJG
KUEZHNqRVynBfPGkFw+AnXwuJu42GDraZ1HbIeRUg9tI97JyfXtqT1TG8oQfY611
CYRh5+yDgXzvKYjjrwK468Uo+X3re6AU+eXjEr+0FD3Kyqm+Si1hXe5f5O/jQIMB
0tJ/TfT0HiLwDgOl4DG4+ml8mCM1taqE2nU55qHVjCxbcU7Fz1t3MjGJl+T7nT+t
tI0nAuFYJG0t2otpIZGG5cZYIDP0V+75A0gYclguJofXgi2or6pFY04LZGY5fs++
UqgcevEF4q+w8pnOU3u/hUNqsweRbeN88MT9ljl9q/0TNQvehw57rU94rUO9S+He
PjQGF8fM6zS5iuuM/TGxUMgVM3NI3ZkSTlNn5U/jLetsDmOd0apkJew5qJG7FSZQ
lUn4BMD0Kw9qVAU5cWnqzxQkJ2yYpxKZHSPBZa59vuX2fSi54TdWufywF2/90PiB
ziQiq/dm8Kvg2MqEwL7Jgn/p4UUNRh9vzdkl4Nh3rXNMw9qVpfkTX/xrC9Mj/Nwx
9qKzjslc0XYyP5oX3+OtZxDpp9ItgMiJmwo0cPeS0ywfg5Hwq+Xb3gKlhHa4F7vt
5LtskGc9iz/i7uNuSPV5YrCKZg7v0M/6/n16ep1s5uHJtmbj/kE+k7+qs2/1qCZP
ILOmpf3+qDfR2XlJNjzvR+IyL+t/koxnnLLlZWempZhSWtmhHc9I1yan3Oxe72KG
GZ1lTGwX0DgZ5ILo80ARUj+xYZT8yXn5J3eRkrPdIHIlkn4iW9F1knAdypVn58o6
vJzCtlSdQlXbG68tFUktO9jcPuQppUFIJZVzAc1APrPYMRdWoiaEcG6DSxWSUkqJ
6SS6e2FEPrFCedEk9FxcOGaVWXaAHir0+TOwk+hAZ1s+C9S8101brRJeFZoYuVLc
5a8ItlVVpVc5StflewHZcdKRizuQVCCinQvZfEOF4O7gD+rQrSKZXjKSQXaggtax
2HpnAK1ReTgkxlAZ4geLa9yCDyUHbvWyQNA/u9Sd+AKu4/sInUIiU04Caq60Ipg7
zx5wc4BF3qMG0W7UD8nrl+q5LQfQ/u8MgVSikXhoNQo701Tn/LRJ+cenv4J4yT57
pEhFaNU/9eYvNGMXgxYG9PAwNLjFjOJx7geNO4iv6wsTBnvNKg7/6Dmday4LCaXu
OBYFUdLtzuAs++KhvvCJJbRileSaCLRuLp6A46n5qeKodNECe0/9vGgQ3pxFAVRA
BkIMRFDXZHsQFNf6AXTNBIvWlOUDH65MEA87wUoEWsuo2hqbVGkQtVwxPbRUqVT4
SL+ttdKCgaYWByrzQYAs6B/qkIxIHSlo2S6PFiakAv/8QdztVu6tjg5oAhri6mra
U5D6owRFNb9jXFkCcgUQSuKi0Y5fdYw2mXebNzN5jSanQMu8YCe6cm5X9fE9Q8Ey
mlobpjnvpZ4m0yTJQjN0Bm18ij/+WviJsts/ZeXXgNzUJHvvAcn2U1NKLyOcD9QZ
gRQPaGNyhamilZiTymwLVlH5rydt+Gt8Hc3MvLrN/ena9sibxXMi4XX9lFzeFCp3
7ecIb5rE2bnpZjUSSyMaoprl8yQ4u/CDx5prjp0bGule/G1pmsI2dpnnWML9qLyo
36M+ROALfcg+ali7sU6LYD+Eh7EH/Zyt7GrPhS+eewkXCPMc//gBzbg+8/NFeAsJ
1RkaAJjtQPuLy1AsTdACzQWQ2Zki+7VCcYSwufTTuJSqF2ofYKMD5rECBwH25FWB
dFCRcWCnJEKaoPi0I7i83XP4El0zHYolG315xKDDlqKoC2MTD6+VMvRDO2dsAazu
v2PCJ/hWGGWfrwY1EobDvHV6qoNarleSg49ox1/7Oykp311Jb01WTG7A6fX4Hle7
AHY3mq3rusTEH7BznT5mXbELReWPrBYmDuPhvJtetzLC0v9tJQLPOVf3iS48QK/o
lISrNIcgJZrKJTttZpdNOf9KNt7WVKS4e+BmGtaSRMst0waFxw5NXWJDeDHQTS0X
WIj669Cuw27+b6XwXNHg6XdMjCy4DunjJjDXHTP0b5FlWkdXp+I9lH83VqRC456l
tC/LemDfZzxGAGSsayuUyppUlFKH/Ohx7vnX3JK4Sk8vuTh4Cy93G4MXlONTNYaD
1EWkNkHhpX8fnFOPvBYpITTI6SrucmKzcDO0xI9/L88zELAZQHLi0rcGQbMFf6UY
QZ4Fwsg2J36NWWIhxRMtSZLJ/oTdkNEB6Zfyiwml4Dk3QgBnpIgD4ctPW14oXPFu
yxrQoqfb46RNWk5QKMgRiVF60MC1rlLsTGuctIuXLvMhnpEs5OC53ZXlV2saQPze
iqeiq5FlHquRh0oDa+IJWQ0cKi55xSRwVzoznuepNwas9nnWLjxoxdYDqDiwCfCx
0+HNZ+FAWOBLGOeGkdBQ+y3Qwose6Gj5jQ8ou/PV71chyBJ6GaG4jQU6HbbfaDRN
2iOI3caYh+YCiEOeFaAERp5GusOfY2ZYf272hmbYMEDkJzEOaD8Y7PIzYu3IcHIj
23BMqG7bLFptpJugc8GyAKqt2wBJzsDpOunP49CD/FfTeSsTJYVWeH2i/jgI27ZW
jR5nVha5SkrhF1kKHBNHhVuveaacf78GPDcKnknfzAK/EM8+4X8UT+E35stvZrct
n442N3joEYCK25vFbTTPBagr8S3GtIzb+4NB+oAAd7qpSTL55U3LndclNxknplPh
Gn9xuXIQt75iMh6Zpo3rrge7PbnOIdKB9eKv5YMP6zaB9WLBJNll9n7qoGeshkgM
4NykIcpG//X1PcmtFnRj5EvT/tC9g5etmrvPiDlnYNf8opxL8NdGytogcwacmjlj
iNyZQTWpMwtc/jmadkU1eePTjqIRzBFnzkwvPupeQwqYmK0FIo8w5w3emkxZa2vj
vCj5Y11ECKydysSnoY2n39B2kYypWMVoQ116fsdzHloqlTRAgfrDm/ITAhjAxUcq
naI1WhPYkSOCntglrmAQCzzgF+wn5N53OrvovG6BQzdrrq7uz2wv2NMH+RXdXpgB
AHXRKl0vrzXOfOxNYNQhy1Ms1D5yF5Uhv8ZTcMS2uU94/3ASv9z+hcxqHKI8vTFb
Gq+BVt7giHR9gE8RDOYRccxsEjxNoEQkJRVABFqGVJU0BM1WYZDXVfbQ9hfWctsO
GTB5cN5eZZloVITagbNoV+nviVt3iDjCSGpVh7w19XwxTCf3mt80igidau9RIwqR
OanDu6x+0w08iiYAa7JM4rCI3b2o1HKxZ4p4+BFKsvqRD4NlvBt/1TJE6NY+BXhq
3b3GIHdLxBFnaUh8lQssTX6um2vcdkAe2G0zZR4BdKmiHJAx7i4uw1Uxv50ueaB5
NtI2pTqaWTB9v9Ry/2iy4QjYy5UmVs4wHp3bvDJ4tDDRF2XI8SfluZmWc+n+85Z+
Hu8ePkiKg5YPSTfzDaGvuspl4p0KUYw2cAY8l9w/D8O+9m/z9zM4UAowIIKc6eyu
kchLsoaFgCMLOpZQvdO31hoCCrXtoXZKbVWD2QfIV9PFoV1wfhmt5xPnwBVbSaPH
haXJDRpjA2jLqPfws+zCrJ7Au6PI4smtYbGaFdZTi1UzBvqxyQjiYLV4PusSBOGn
t3dEVeBIH/WGA7x+LXwFLHtyQJIj2AbDAh32NQVuZm1hYOLShT1OOBZm0YQ/9ouN
sxYY/LdXTMJljweeoyZQ4t8fPmxby00bFovvgqPwXq1+hoqdVF0tfmQcuFw/AA+8
CvTshPDhZhxGrfEsWn39QJZwIKmN8x9Ft1gyNLkamZrBpLUbQ5tFuujPm8viaZxb
zB1gfZzkLiqet3Q7nwAw0wbnY5ea9EORwV8+9QEzkHZIB6sqJp+OkMv0z6HmNViJ
3QHKVL9CqcZLIsfbQt/vnoHebToxHt4uhByI2KQ2x9+iMCZv1WvoDMud4xpTKaXK
rwirPHtGqlrLJWqGpzWMPuqB8Imx+4Isc6mANygbH+qOmKf+e6KrxVzsClNExLbN
WzlAvB3hP2Gw4bc1Qplug3P6myk9yOcnNwdWkdyQX7aquadMBz2JnUnL0hdkLWU9
4i6jiFwykjfh8pASDwUM/wmvB/yRnamLKIz0QiowSN9vDuqYlUset+3UK3lqprrS
NA5XHP1qw0wSOAQGrGBtJdxCCjZ0kw27HrJN/c2U1Pf807tWhJRsQIaVlTvzxDEB
0mtysHTXT4+KgH+Y9SpL1fds+FOHHQ4ahZ5p0WdlNCi6nQFISFiZrKj0gCo0eBNi
CNFbtf8jy20D8k8BEWMBwgB+IVnEsHWrwk/lFWIEhf2ONQS9tuTbfEXOGgxLtdXG
rKrPf5/9oQLDLOcfv2iCRfcIHqbJC7FdGknAqmIpfLDIWf2CFhq/G3mt1hV25hPf
btO6LZnOg8VW/b/VkirmLLGgDM0N9jh3HdfigPZ10hDntVof/Js7+d80NfmdeS7P
xx/0jqRhD3jW/UeH7wEMxXe+Q9BQHW/ng40b3GTkm8jE35bcAU9NCOryYnvGbHRL
jQ5zBF/00ijilpXnFo45zQv3BSNiedFTB5zrWD7Ib6C2X91vgNxai+bUEajuqhLf
y91U+UXKWYEotXiepAsdbYIkowZCMw7251HU5+7o7cG09c2d0usvizVlnkJOR5QF
qIhia2xlcAqfhKBBb4mRlwDfSzE1CpIlCkDzvO4OZ3wsL6GX9h0+QCLSaT+wqnll
M0DiDSxLWzRRm9bicOWwr8uQIYIB4PtXIfzFfx2LRnzaLYcrdmgl4+wmRNtsol6U
sNjKATSj2c6HbjLE0WAClTMZS4opI57ZS/I1V5Mm535jObNMyzSX+BpfGsDXiGLj
Sn180Pmc///C/v93DqCI8lKP0/5qkFKYygCjVoX3UzXrjBs7h2b7Etg/6f16y7/v
XUw6nSUDXAZPvbwgQ9Fi2W6z0g55ZvCa8i5+tYyfA//QML+1C2gM/Tmt6sZjNqmi
mQMd8c2eLerBRmR+M+158cSmVlR1fOzU5b56sve3n4weYtoZsVD6bP4P4DLRUp0+
pOFPdRAgLQNcWVW86yxxVvW8xf/INz7dCCkCb84XkNj2Iq7EHqclLWiN2cvZ8S9a
r+3SBvW1+snRhvGooORmKDWvDfA3n3m1V29yH7faXT2lLCCEikbjNLxOd/gmxOdg
5uV/Q2XwPenL3I2N8+jRDLCxhQaUIYhgtCSw+lzRYUa0hr+DSYkfaFZJ2SWPMmLC
YvUq0tsqrHEnRkAMjO+zBE6CJpOj7tEqVyfFlSc74xhrpUZVRFeBCdkRoFBeZwok
gogPwimS1ehrt32J1Z6ou38Z08p224bS7mHNfntLOCoQcATwj1QG+B6pF/MhsXpf
Z+lqRJRtYyEdloHUvvny3fA37AKZPBrLKbCFL+RNIA/94pNBC4985jkMzXCyR69f
kfyjnOaPKQ8jb40sZadqdU5TcPM5xlUUBWGmJqRe/Ht4O3YHvPHlRPyOy7PCMcDG
L0KOze/dcmQMobjZdI2B5a7pckyDqYBjM59WTD/JmXFa8vFns3Cw4HtgEnxLmq7o
weHQr1otzftVOH/mQIR0beYJ2i8IB2PsNisPfz9oDvKFo2NPFc75r1rBU5u6hYH1
pMRzLbDd0Vj5qQ0R8bxxJvXV1BpSnMoUYuiYB3MOlMLCNMsBYfkWybOYZhKqPbEa
grEy8zuUQDeCUelZPd0WAaWR11SEnKER7JNcTVTGz4vcuv66N4Zf7NnakP9L/cC8
+pc6udRllEMobTHBAXTx1YIGDFJrU/z1Cn3vuCqMOxdVFIuKJbGQp9o6esfWQZPu
T6SvdY3I4XHzLLLB16uuJFMHWnNhHf+UcqND7i4/4i/86RZ7dB/9TEVB5EvvFN5D
XzkL1sJiGUEYLa5arHAYQkf1QmYBx1mPJhJk4IYX1LxEYD7aCfLBYwg2Cp8jUnIT
Uphq2AFqiWKQw4G8Y6I/GiVfuttufqfdlpnvlST+Q/gPVtkn+i59mLKYBA+ywqgG
eq/Jnp9nzsNRQwPU94I6pFbXZisBmR0Ljj0FNrShjTRkScxVmVVT0A+oU/N1JWLN
cqtVlye/u14ssEKbjDkaQEvtS0G/WpHqFctwFMxB3iNjZNn/awqgInAuXjv8Dmut
w2hG8ZOrptWilWxOxEUwFvRJEV63DTWLJXldVylFAYDr+peFmEYCUXw610TTrT5W
iu5PevnEIxanDz5iaw/17np+Ls8qLoH7NhDmaGZIBTE2faGJND23dmvunTwWacrn
b5iA42xgwNa7HjhN9aBenmDYeDrl4/ZIJ7AZD4HTO9rKlwB57f62O87lcf7tQN1n
F8ydpkUvll/nSZdcZ9zJIIz0dDPqfrArbX3gj65+zwi9+TWKvAzbtGOKT4+frcOV
4SJMALXsrfywk7cyWrB+DcKV1z3g+XBekLQLdIySjtvh7Xsu0W3Yo8b5lDLfzZQ2
xTvNJOaqNodMbdji40kVwjJxedW3B6e6J+7PA0jRPGRO5wzLYQMvocfz1cmGSspX
npYFgdrwjZ3nInWiPNlv2tIdDbfXP2u3wDDi6VLZU0crZFzzVHDaNXV3dumWXTAW
64jcJ4n5a7+AsZnF9AiOhIY0Ixp7rrA7z48tbaM+HBIgcilaMWAMrzMmRpQTxHNo
TEC82ZSAOZPI6j/3Xy93ad3Fj4oNL85QHaNjRSYCF/S8lDY/MT7TjB0jQhFULcDL
jbV9vlOa0eQazWJVKYOxNo1KtzAay1qkd04Othydmmwsu3YniUFx5JL2UkwKUJov
EZPOH2AlCssig5IgahWDI76VVOZcq6AgpLxarBi9zP4c/1k3pN2g/14CAHgUEsac
u2vZ671nh1P9oGyKTdu6gKOg/GHwOFNIkeFf/FenMuGLWSRpHYtTzSO/aUBfFUWN
yPseYH/XHdI4SoxvIICTPv71VONe9A/3B5yJdufZXR1aPhqhARIdb2cGJPZbN4dL
rGtxgKTEDsna2xHBP9SNIcY3D1z+NZzY4rc8ReDAJfywqBPLiwtucmuhoKSdIMlI
SuuOXFqN0cM1fTwm4onAiOIttAisr1xBO20ihPVSqBz8ULNtKwrOrUfEXbORXhbb
SSd1Zyggx2NOMUEpOAJhaLzT5Th0LJ4SZvcOrQV6fYZ9qE2COMctX/G7a069iHkd
WcunS47QAlu0/VfSNeUwAQ+vrv3KEEEwl41/RcG8YK6eZpu91GF+0Tuu20pS4K5S
B45wTNm9S7IZ721risjYj+6CjjourTMs1nfgeeWfBupfd6cV3wx+FlThiynzFwEk
rl60tuhB3Zd13uLjB3LAkMGKTkptUV3A7hvo223JfnBkVuvsayJiYHmkNJHPvCwP
S3ry2U8FDyDBrg29OmjuokJHHjaK6qkPgeZjMeFISEk9XsDOUgPrs5yIXTYM9fJp
PYbIbhJltIjEvL6qi9Q0EXIN+D/st+1TDqFvRLMUpo+n90GrDORQG1TvjSQ4Jupg
Pn9a+Uc/ADN6RcfP7WHm/5Yx/3ERUmrxyphC6zyQoRpZcmkwuuOfGZn2gAuH3Poz
rd5Uq4MuwSazbtuM1lz5ouSaIy/T2AeCVSqKGJv5Qnj9c8TIMgLMU3IDmUb3nrxt
yUy4YdG4o39QwsNrf+FjwxKmgwiU3BFXIjWuGsK6p7N4cASBMM6L3k9kpquBl7rs
UIV8QkVq9cENx+HMT0TiyxaxZZjjVg5gXH+l1Wq5NKunSpRAVISMyu/3uodY3mxS
mulbLAmJxIe3O3o4pmsKmQ9by0ulduxRGjl7G9oGnasL6i+QrcquQygREdl0BUCt
vFZ2jy5cK6/D4t1piEmqgesUfonUYBGV5LWBkJmRZw/fbkdJ57+pLHyWKHVel+NX
mIZz2y5swM74gnYRF3BOx+PUqB37xLccI0AG2/NjiLl6Lm2CR+/ByamiIVaHo88n
E0Fi20fhgjKqT8L2QimLFEc/5z4z7ZKROsDsC5/UNXnZFB2yzKj2V74ZHrKXiC0X
pcdOF5JbuaQU6uXK7gySg4hOhNs3Z6c/6m5v7pd9HKvc4Lu2a4xg1APi2Y2uVLuO
CoZHmznq21FHCJPIdbPUyu8pA5q12PmS+IsyovohlwLa6Ej7ifvxZ2SUEFI4fNLq
E1Rkqd+I53JTqVsl8XLmVpZYvR6WCxhdoohW/fpanc/1jYY3Y9imO73krfT8T6+Z
NAOFyT+ryaDK0eA7VKPvUHEc6m1iY1Yjg6u8ExckRCIZhp4SeenBP2K2UsPfhCL8
uRA0HJTMeiupT9ove3N9g1W6Q64BYpB9i25o80RStg1mFVPTbbIJD9UGEuiT+QPy
/Q4Xfkihv7WORFAn10lnUeWmGszdDY9SIZgHbEgsF2Qp91NvbIWTvwUdBoJkCxBD
v1sC6C6PMOnp/Oed6oPTwX7t86LHbtKO8kyWkqBra+PGnvJuYt5PXF8pou395vyg
EtGK7sbKvU039QCdKA+ZjnDlMh+tjN1RRUCNUWXjpiQHRgd9ty4uw+gwSNQQZ2gW
enaBTZolUAAPn0vKV/N2LAIlzOQqnY+ASIuUjUyYGoOxCbfXqf+Ae3tdnTlrj21U
93DLN3bWHfnvR+wmjiwB1prezX2T+uIbGUH+Q2nfw6pdttY8T2FZgYudSy4yjoFP
3DrGWjEFRRkZk04nLc8JzhChDqZXSpZ2ff1K1RnsdPlBIEkkuxlTsDQKyB8XToIV
Oa+UUo8hf2P1oEm4G3sedsThSysdF2hhARe0etHbiQ5/O7N8D9XIc4bkST44Vhvh
YbQ5dvAJAHMDZjqSXbQh576EEED4SFn2NihDMa1B3h2/jLzYRXsP2ldqF/HOPOeg
vbIvHL/nOpDIv21qVXNnjzX+JeimDOwr8BLSwYxG0534halupM+GvQvuI2aKFp7F
J71RXuLIRU++j9GJrC54Zocs5IhBBstzjWbjSsF6f2K9wyXOuA7k6q6rnrrqvokI
/K0vwGWtj8Gi4VMYTSQw6pmzF+afuX+WezfOQrTMMo2sEA4fYJc1YpXMFsC5Vd6k
I/CTUcuUnwsIjdaagmrEBDpPeenI1QPi/tzJvYrFe2PdK2dL3ohDMDfD7G0qTGmZ
bKaVrnZno7YVjO+QPVSAFLmt9vAYuAZXoXd3T9w+jknmuc0TqblWFGe4iG+90moF
dqKBfUNhv65CBDxHGMDrERqIMMxvC/oxD1/AOxM1+o3nOig8QFhCF00SsmsxrJ4T
v/D1/cEZ71yfeh1lEJ60RvQxtWy7PYg6G2Knqb7HHKit1p8vXnJVhJY0aSRCWwM3
Gk39MoKh/nEsueARXGguhRPQOz2x0HGf1bO4wgdhF1v5NgnuStFOKGqWtCkZK3M5
vF9mnx479Ip/gUqJ+SX/IA5+WS5zn6vNuLoBZe3ZqtkfNR46quWdOdS/9wUPsD/B
vBB2E/+atYZ9fzPaxS5zRLgUe0R8RGXbBEq3wBYA66F9I8Q4G8/yTak3XKme3pOK
dlqb45vrPo54J87sqyJGQHDjWELRnzVoPssPR/T8enewfhFlqa+HFrQW786wMXe2
wXbw8NEJVb9lMB3fjhpDJFXIp9uqoqGvALFTcDcttmVbscRiv45alGSOeOSRxWKT
WsyY8Xw6j7AYL8FzGbW4FHgVFSxpwUvXpJtB6BsQxSol+NjIzQssVpa9QxY5nZOz
JRWZEmdiIoSu7WgcGqbQsKC3W7kmuuwfNG3cdnGiNPkGVJWfkb2jJYtzRxw8wzRz
XkyApfAILD5s2qu07YKtrTprkvqNhiBy1frnx1x0eBlBiSqPgiChUpJe2sqyXTUl
vsaYc1D1faLWKJuvJx6Ski2u8ssQ25XY9gML14vPO9N78yBkeHiyuq1FJGCL8QBW
sLDZJFdo2ZIIRiTr1ugxeymlLTtX38wYml6Agag6c6HUQFiHXgqSt15RSAg1voTa
rgPjqA/GX88ZPKb/nzc4YDKxyofa9/SqCZbjIC5+v9UfIkjVX3nNy+OpY79ojS1f
B1o+tUEKnOZVH4ZKPejdyUjT7dkW+wbfsud7a2p5h0KhcZt5TeMjRQIXUPiimPIE
vMqZM0N2kwqdSbxHKX533umyT2s+GaJ3dpZFshbG4Y1iAAr5EP1zHEcfriK9ntdh
hHv+t/W1oNGgc5FMdGT9luPRkmo9RR2yOm7oO1+1Lwlu/wXytY7SxDg08LUJXpHH
VZH4+J85ioHOzD2vvOG0KeP55595mX/9EcNrhdB+VYe770CixHu4CHG/DOcMIyOg
AQgmJgCA4XB23mH5ACBrsvxChENZJiwfHaKvczLczJIjT21hYr0y/rhOuz4wkhXY
xJcnObZbCH8mM60Hsuoy/vcz8D/bPmWfBVR/SupU847hQ5/o1k0IyR+TWA/Z6yrx
4MeK7bPCPo7fws8+CWzd3SIh2p2oI49d7wizcuxA+FUZZiNlkeeDCLPRKActlbQP
7LfVm5J9igzRxaK8MSqdDzG9AStN4JDcstiwzLQPEg7WrxZWdT7LGivJMA80qrh3
3zWlnnrl8KDcmzSJ4qW//4BN4iXPhWQ7Y7l3EBJtmn81fcmhWbPJ2W9PECHpntXS
/832YZjFe2RWNzJWJzCz69fFYBgrBDdXbNPyQJzXHhzvuRb57dRVo4Bd4swLN99N
YgUVUYKe+iXkY3EIURFQOaI3Ou0e6bqSgQAPvziS45KdgwzyM9tVSVCF8y6v/Pl+
lx28xT6zHpuMU1XbulIRuHj+h3TagtOa9rJCeKR8IVC2f25VCbN0cNqqNliT751a
39vDLabfBkvtlj966iMtwRVDCJxmGLW77331S8pkYE+lnYiTLjYSxdKUww46WLSY
8a//yxYR0rW8yIwuK/w6Vap15LKNJcUa5AcyPmNXJ/LtevnSSJYE8Pvn1WtSFNRS
2sCy1RUmWzARS8YusfAq9M/PnDb+/iR3G/lvE//VaSUSrKEoOgISzOI2KWxq9XBD
o/RkahGbga/MGUaTZHzPw1smWOnbx8XU/57TlYemrWpxazgmEfdrR2eAVKzYfS2o
fdKHjOMBIN1xtAZneWibi9fAS8UIWM73fUFAuGZ44cq4wFJta1gkxij3fl+bOA9a
mv8S1BI/l41gk3+pLq7FDVn1bzCxKWL2ZAL9O8d32ou7XsXeSSVr4yrkatbEt2CN
A+rOCRa3YQwM4E8s5il9RqPPhyUsU4s5KbF+HS+tN/34MDgEb2g+neKKiI+XYWS0
veHSnhNV/0rugJYH0k7kj3noh5DLLN7YHg8f7fzHiJ/aeF9r5BNcQyTj2/rxxi00
NK5vtXCJRZTBmcTCKQ6YIALMsnGRqIlucVN7FL4zLWmTbKDwW6WprBpJllamNHlS
eje1V6KKTtOQNNc2gNC4c28icBn221v0Rxm/7rjUcMLoWG53p+5eP6+yHGFgGnOn
M8S0lUr1sLLPt7Z1FsYcP7UkZtOu/2HhRX1x5USNCrc16pnU8anxksLxEK0YixcL
f9gq4Q8nfsgOjSSuTA8Mgoym0WuxadNOJI58b/M6v42Y1YYUfk4O0ouRpt/QzcdZ
VIVOph5ag88x62BCvVzaJtvkst6un+yCakDJGVAXcZCds4/UKHWUvvXRsKbAOI9D
4ke21dNuuxTo3Ks8C11OdbNncdijH+uiLJwJtKmwOyzbP+jM4zm1q1HTeUD/fVJ+
ckg+9lOE3YOr1gj4Se4NiuMi6i9JM8LtBd6lWhv+yFimDO3hexgX+Jm+5lxvtpgS
kx+dJ+yk96BQvaNlSSk4JLSPgtQLx1MVZEMiGWwKS4oU6JhTK838WWLTxclyU/4/
V1DghU8JYEcduT52GxRqI8aiavf+sJiZWn3bktaeGuMct6MV80BTDFHpQ0kVEM7N
oTPP+pAH7pPfM1JYzfPvjmNG7jeHBFuqdl/SqcWDYSET3N+VsVnyZLLB2jH1uQN4
MoIsF30AFSOeM/8IwbogUJBlY9LKJHP5/RFyD1gLG1iT+cGB/C3/Xoeck5h/q7YB
106MmXxzy4rRb/YM0qmddiUQECpXqJ0btW0CTh1cWzL37ngv7alntU2tiiddS7p+
fLbb4eSHTXTdga/jEkxw6KZDQ+ojuO2xBsj3hqwCTZLxO8mLhXxDvn743xzGJj1o
/E7NpSWXk9KYC+e9cfGS6ly8VwSg/HCNVAZ5ToKelHgj0b0wl5/Z5i1pxPef0a9p
/LAyX9oN0xWWp4Jbc6zEsFoUKh7kuvZ7o0aCn4Gi9xUfpOfN7K7VVI3gaLajpsGv
p1oqpFEINv0Lfcd7y81UtpO+DWEbcmntOjVMbONJmYkX6PWbK2/ChYhIXDgoMMAv
mSKDdkWdwmBCedOlwLChny+UWZKYUiuiUsSztGodH5RtRet0JjALrx937aKC86cl
Dw6EqDfNRnQYqfz9n9WE+MRANXM4GI5ZtJdppi8eoUkxV7TYCAcav7qVINc2BDQg
o/zuBun3n85pQ5lLcqVrlN6gcdTIUqnvo+H+/vk4fh0jQIeprXNKKmHZFXxU5T76
1A5hvUObEBJ4sJ3QU5mClQqnMtQjG8RP7Eb3Yv43X0RzA6e1fBYq71F1ZMs8N0Y/
SMF7PJq3Gsk6oKFHxt1u8IoVlKM6OSxmz8Kal0Q+I2Kz9YAcELqR1vNGCODKrGMT
tPzrAweOrf6x0xq7N/8RAm7jDRj/Wb4P4uf5o5RmE1Mjzb3w2K/bXpGu9UFtGrww
InvfgkH/DL2bf6Nag0XkQs+bQLRQIxsnig5JnbM79RE3AWAKqtxAx+Zx4TmdEM4G
9P+6QwiS51hZJNHIqL56hR3fhbdNzWGWMVPK6+nJThLddGgSeNvIuvuDfzGMamG3
H//aCQtC7wT5oehuqGzMydyvsOxQKbA1Zf6LI99+sll9nxVG8Qw5/QHumNie0n/B
dBUwJd4pO2D7kzmIwa6xD4WHakoB2NS6B6ipKG5tynWaiHiy6WAfiFdgpxNgQ6+l
k/T0IL55vM5nUbbkh1x0SYbt31yHFIN8sqy7BzQ1MSYF37XDDFqLjYOun40Qf1eF
DRc1Ma4BOp5r8hqhdn+ylFctHEXGF5SNa9yjOU4pBwCFKBgWLksOHPFQhKtDQ6GP
2pMhTlg0IWXMydpDB982cPYB6h582FiEY91THQ0T4yycyrmlQdMmbheLNYE/FUnR
ngy3DlJj1Q/Edf8oDbuL3yqYo4LsvaQ6JFLRxQ/RTTiKTAEc1PdP7K4W1Ma4xVAv
LozUbLWQ9vxii8OEa4LDU7E0jFuURfkcnNEeZQlstsPt00Z3Ugz3fr7v4vLMo92G
8lNwd+vHQWgixEJ5P1EhPwO3Xbw8hX4klQr3so/5nmEelI2nSSq9qxldp4nR93vN
INs8/JeDhDDPaB7J8ahrL9L3EpwsGrP+kc/bmyTyY9JrmUc/TcJAvcNzzNq5Ywjg
dGDJLyBI29Xcsb34wS2lLCbBW73QXhHO8Ag31EUssf5+Qw+0+IWsjPRBYBtldfpQ
uR1woyPXMVB9RTCn3MaR6ADa+dXMsrZ9v6siGnkPr5VDLhitI767VqO38VkdwUAc
BnKtHzcEe5iktip7L2G7UeNcadurn2d9mEx4tROSIV6T3Ri0fs+2mLL+/VTI1QUO
hMpNArttoL4eLquauw798E6eobGbZt1L1dHg9DC+Ey6xK4YiLfUxzPMU4UeBHSHj
MuLiN0l3J7DPdL0MEvSJRm6UZFZidg0ifhzO98vSu9axvnM5/diZE8Ux9BMRkJ7x
7Wd2cd57/7X+JMJwPOMDmyOWLfSkuSPrR4rrxaMrZlfksY4uUwBb6l2+5eVBGswb
90hkvM2XRp4HIso5E0KnxRpSvQz5tspX98e9Wp0Y1bs9sthY2y2v+s+q+0jdqtqQ
qH904VFDB8lC37/H0NID8EMKnHcaNTXQUzMkPTJ4RU184NvG/o01fqEv1y80sQ+J
TAQfC4kTsVEgiZymFCc/PoPA4SIP1hGMXwWM6sJNd1cPKdnozp3iWaxvwrVmbZRZ
8VhS2KBYqAbzEkCEd6KMtEBGQWbQYoSqx42C250fyJOxgVfQe0TDDG6cqvgMXvbz
d2Uj0vPM4aWV4/8+Fmwh1Nyp4LoSvfKamMW7PmWlqW51QqPuqDjbXDtTITMkhOUn
FF3NQY3XiZSDe+h1ziixs1JyC2u8xHJqO81qVBYia2QLQPu9NBPDXSxNhjLf3M5t
Ku/Q3cBNaf5QKTw9dZ9+g0dNdXHUBunl46UALJIo/4pxfS485ZdKRNqRplDppnac
4ncq7Y9gZrgviW5UASN4tl58zEB03lgXrSWswPj0kD+4b/zBQ32XsRVyQcXo7CZ2
7hy/2ThZXGJ5UT6tjcopmVqKm1cSy/IKjzbWtB58kv12Ig6RPIiD0w3CiiEuNg+y
/PW7gtzijFs8Hcm7oSHhi2WDHdkjbHfY1QopY4LOaL3SHS3vhR8lx8NsJRcS0QxD
xB77HotAzJ7Q8iA1OwZdxVeaTUdDwhHEtDAret8nkkGWeWCT+0inZUx+mHOG5mfA
vFlv3jf+lfnR325y7s77yEjvKkM7dOVZp5m5Io4mnVhIvq6YgE2FLmxEgRdqLeXI
0lvI40/qiD0H3ywBGZSZ6YzM5hKtqWJ6vUI54L+3U0TNyb47i+5rPpVXlEWk6+xK
7JvK20lCBlDidPBWotbNxfmVHdSL9VtehDbU21MZZFq34A28L+SHx41R1hr93y+N
sKrxpKTf0rHBAoZDdGggBM76UvkoXl+sD+YC5fqBLGVnRfV5/2a1or4Li9Tk0pFF
HPfsZPxPVt7TvayOrcV5GbU85T76zUguWISITYQvIEUgrlgWqHQqoqto14cNu2h0
iAG3NhR0LpT5t1ISmdIPayq9QzTBYEB3GpsPENdSuDerugwagZwwAAPiEfC4+fgL
nZn8mWQ2trQnfEJoCWUO3uMmRHTqfaLa4fOdJWEmUDxmaOgcMAe4VesL7nomHYdf
wjePu2gcd524PRfP3eA+Liynj4X+TgRlo9zjKxOjrRDo/pyInwuHflsLyNZtghgu
RIkhEglrr2KAMoQCVBX4NzLxjR0APHihSiX4B6Q4mE1wOPlV3jZGDePS9iZVwtbj
p1Vk18J5a0Rq2JJ1Fi59SHlUbqSLqFS0v4UV8PzM1rXDvDVYh09qm3X7UxqvysCh
IpidqIPDlZrSB4KOERA2DB0qY51zebZwn8Mt/NGgcKRUgXGxQ0OeB7fNFIJE6Fcp
Zuhgxnv0eREc3ttE4ZjrQza+q09YMVXhtb2Kj7Li125bT6T4TiiYW9d49DnJKovg
JFr7m5nKjRAUFSVJQ9tlTnXsQmOfQBP6QERzjFT+JyB6Ev3G0ezGVrhVTNwHK5PB
PsMQ2S51FP4dqUKDGkPFJ1HfRxE9bdWW767B3WUlUq0TVMVOMMYqt7Dn4oIorGtb
lF69hy9xwbLHmKLMk3imLA5+uah1K2ITHcnXsW45X+m5pJwhskLALek8lNAI0KgJ
Th48ddoQj91DTrnG5YDti009bvqEDgpXJJyAQYtTQpzThucnNVvjGJyJIcXNTDR1
eIu/LPn6t8JUpY+7mK/Kt5gdvN9TaShnmmB3rwq2IcnrdfaT5xuOwSYEkf22wFte
puyd8zOIPOQhNtMMQCT/ziK4lxFUmYZCDnGquGiBfdE0FinH/1rbkqcvtkYY6kzZ
QnEMkZXrwNYVgcMdr9YavqvdPtDFpB0/5P6NKrx9PAIP0sTIP6XX6dziKz+QIezY
iLsB24Zo1m5Oj8qgUMP98hzG9LiuJ2FnQMqPHoKiV414uapt7QOb4FW5JD6MOSPe
kUHNHHPwITWlt0cSxOK19cE3Zjm3BxzYzc882wS/qkuO39dV5fzncclZRwOPw7WS
4XZPqSKsPLsQUj9mhZAmGd2V5SVhwLUXAKS+CvpuOfcBazQyTGOd4FQUgta4i3zO
qiOgWWcYr8XRvnnR1zTxm+bCa9zSOUorsHrfCu+dPvaT5UkSyozOt+eh4VwBg1w/
ZMwvwk5hunXfbEFZ65YjKhkHSwcA2O8IEkk2lDUJv2oSj09SR/xm7I45FkMsMy/O
mSxFfzRCDq7hL8YOiJf0sinSkqwA6ELPlxpL7yp2HC/fLNYIXyxHo2kJImqvuVpk
tCHb46Q9f8tqmwOPCC0/niVjkWsIAExM120fORl4ZfyY7Pueq4n/ZVPhZOHWq75i
MNRWtBP4FX1sxnIdPrit5rAfmBIrF3fTbVsDgb2zB/Y5qVLDEAhqnu+SsEa3kijd
8goQmlcqGpZoK2meFTox/XTxvJbAZBc/flm7XmoJ5FSb9IeG7cFxqQLA74kq7Clc
uQ6QZTsKlUXH280pejb0SG/WVGgZTpY2Zw0jWdVU5W+IOigbQtcYWYZ+NMmgASY7
NAlSSEgIJY2HFvFngKAXXQudNU9VN36W3oi4s/jbTmzdPk+DCFATI7jwF1hBvscA
Fn2Z7OCPecSkE9+p6oVNJq7nattAcQwGWF3iZC3butupIRye5pfV+rtdEIkYqiVO
malXcDfjiMN/U64nEvW0QQzDOEHXud4gsaIwaw3E+iR46v/7by4zpuOrGrsXSYm8
XVtHXtYJS9FQdPhPTN9spX/bO/inDnpDLzHYdnbL5JCWgskzktrZ8ABiLZNJuB4G
fKNrcz4osaSCYsaBkexJK4p2tQbvVmnZ/2E5xQwVClH0OxrZkHDEkTG4+aZw8Qt7
FNzSbLJbOmtGC2EZGH3/FqMm3vnj8xIebeb6nMZ9f1dVu78M9KVMadisN/6nusxh
psqq3h1Ahj97T9+n1zyHkJ6FgWS9GJ5QwRoS3DZsLSC55GqhFSqnl5h1PDMLhrUR
2Ln/yp21qul3AeXEHWj77EEsd1dZPmVQQOvF/uoW2c5ituZkjmbYW+fAqz1npxC1
o6W/shiK27sEHXVgvviIKUjzO8iZ8yz295/RIekl6yPe7boDnS2V2rcA6QfwJiTT
xR+hA8sNjpBrFixoEKepa0ngLAV7nSfgtx2HnaxfYi+tGoHRJwvhfmvsNTnW1j2f
k2meW99uYfIEXzFfyjslrZ4d1n/tMvZpGpeAVVczomDB2ElDc3iCmjSUx6YVohXY
AKzAvjwBQGBe4o0OpMDKM4fkBrbN8waIcNnIWL0icNonTeaAJ3R/eb0Q7NID9PZa
rsW64DHNaUX5cCnehoGom3fJXIDyp41iyQJD14gPL1mjSQYz128N74mZ4KXBU7oc
UYircPeqwgvdsWYjXYf6UOv+9jaV410I1uImJvQoAJNtXmOemv9i826voq2bNeoE
0UensL0E2fMOuN5ncHPaywImW3WoCNJbI3jyyfVmD3qBC/AwGYdf09+hqqLduSlr
TL7elLplt7sNvzqmq87Emv2H3X5ekWkFIp9XX++beJS1bB68Qj7Nf5pYr2bX1I+B
6NDM4VYs7/eYlisnZwdyzSgiqSE14jvVsJ6DzMSC2oZTZh7w7235ImDnDgTjWH46
CuQpVyytCYcRDkk9iYS5G62wyPWVW9ER0NPqBzect/O8u7azmOzyLny+JDm9kCy/
n0IoyryHPwYVmbxtU2TOjgRzvWuteMMmfPt6jQZBz3n7kv0UuZUhScxYMsn6p6nh
euTCGrTANEDRpJq4Q602dX4Oyzo1LKhSuiH1Pl93VAhDVo9kfoeLSgrmVtsjPDLQ
+AtltFKb3K4n+s7T710vczJf7gGnmyEt/29ND0p83YLjywMEbZfj1Pq5invVb2mh
/duAgEPPqLr0jSzGJI9lhqHmzay7SgNcOeU3aSJbKNBjYgJJUzRna8GgUREJmAFi
DgkZscqgEb7XrG927F9PovPxBJRvtzrwNBPxb+XcwggXni72Ay7BXeVtmvEqQx/Q
LxhOF91ECOU+4bKSpvsSe55ebZM494q52d0yPQPP52xhfdTj62rOUNG5voiu6Op9
MiE5t9wuYVs/aTHDwl1TFbJkIal/zC8CdNuSishDuENpcX6C+MjGVZ06El3/toJq
IB/Yhp33Io/5oTjf2TqrxvqaT52+S8inFAbYuqKfn8IvifNJZB7cBW9o6AkEynq/
Jnm0DA2bLseYX6JMldKA+YhvfCsy+cVyN02v1AO/ySWV1rwmpvfMHCc3qo+zX22l
/qjwrRhBcQulEfIjWnfhZdiVU6tmt5NkYfhdEXfoJeOUVZ+L4zgg84i1lYKva2EQ
rYrBTJQJb92AomV81DelFp8dY5aNWYXAGMJ0v7l/2jvpb/g0p7zmIwsWLP2T16xd
fXm6ffPyiU8BMOql9ZnESUaHD//LCbwmw8a5pyhL5vuENyQ2qAcvozSSNLUtBc5X
UKanA6PQuMeJLLEyASmuLNu3E9fVNKEoAs6c3r5EOC47CmIVMHrGA0dc/8L62MlJ
aJgqcfx7XUZvK4AJRFPDDwMFBismIueM4bNfHWe06pW6wDs4+ucFVdt5QeNun5Rv
CQtaRat6jlcDu/6fWni1aCEcsaIpiilklBRSYdsZdqlP2q5OOuBDnbkR3+dbssqd
8oJBQJSdswnbk5bWekAIK6AEyW/b361i59Ct56UKWAElRku4j1PSfbPANMuNe3cS
UKMNGpOy+fDCz58uCbpUytB/+jsOhYwTGlVbob3B7k0VpC3ezH/S4sE/DNFtojQo
XW7Kb6kN9XOQ8+AsYuD/PJyzYFTdqaDuW8gwD2bdu1cMUI8nyIgNyvrwbc4YYqhm
UV8uHKD9FNCsCqzdqYkBNUTS1vFwo6i3nL6WetQDc15wBo1y6UoYfC5IfGmeyoM6
amc/0oNRSm0RAJ8UZwe4QS6kYEH6C+o+7qKmN7nRpCWuH0YdK9hr1b2eyFvHP8GN
sJDe6ExlOnGNUG+46aIHisPEmCFZs3XPyKhDQYQqTgPXC1h3Mjnw/IIIEahtBvJb
GfkvdD5Hkz8ClYd4KHAa/MXokbY897ixK9+2hochTeh6Ko0uOYTZsipHZdasa6zq
Y7mASmCVN7JnP/uuQbXWUxB/Hhwy8hYcYduId0RvxfNL8jny8bJ3QOhS4T7PXObY
Yyy8FMCXbSvNDij729imsa79ipT6EgV/KAI3zox81qTCHZ+QQS7SJmIfMhMVOCBu
baqMJChjfY9sOPw7x1owMRSwc3m3r/2GGFxIoC1oWruI5hX5pKHK1z3mzz/ZylEC
yoeXdshGuQUPS4icRmIaW5NlBpM2jJwuK+E7WuiBSlRwHPA5IzbrBEXDFlJXSTTK
EvA00+IJLVjJRRwHqfSdjtJ7w8HNFfg5mNmQv/fgp/dSbyQLyr2Zo+nnguC0Hfqh
HQfXMhQ18glEELITkcep8FsYu6gPcc/3Z1OEAxU8ctTHGoPM2fYWOzXA0r9SqGYB
ZptOJTlCoR9g4xhRRbIZj/4rAXRzKERQZ9qXnds6McqlfunlJ/NVeZEr5l2EVRfi
/WCyZEQem9H3dX3cX2INL9ETuuw+JoM2kf3YtNUrvl3bx85/uywdo5h4fNGCO6Dm
JGn3G6zyaVJo0Ma2Nn+7ga88r9XUAFPjUQdjzJ0Ia8W4m7tm91f9LhbtBiLIMWI+
HrnEbCORyfRSlhxcTeJdT1363sqYsg/oFbHBHEitQO+0sSZZ2QEVKTW1E/cgySEb
OqXO1WmkwF+Eec5FOJpREQwkIVpc7h4ju0+iTFUz5UjqvFvC8FgA6t+xNUMb2ZQp
8xDT985ObIwb5R8lklVqzqNarSVy5cuJPG0pswqUn6k9jFlACEjCJmcCLtC1/L4W
PPYC2VtRJTT+DylpcyiioS+RXysmRUYDF1yYaByYc6EzSGYVkcvg5A9OxaqikAc4
HQ1fx9z8bIBLMx9YGiLMyYIp548CjkJPyAkigWy8ErevqMuL8YPd9I7X7Fi2VRKq
bvo8Fmgr/T1OsInHbMfl3qdQhe9W7dkcuPJXpK8uC6eTwe9T3vIupicFPFzd3XjA
y2NXQl8FblvdAgx23JCbT2NqcgmU7I0ltp7UNrX2PtPtTF488sZtKnZ0so+vX+7o
tbdQ5T+QKEk+WvIs3aRvNoib8qbBVHq2z8oaSeK/aUVwZJoOXP42hcMJ/V9cS6ki
tZtUOjoHjgOTqLMtGsMZGndJmQdfbsrNN9TodjTxlqAUqGfFlVPbXW7abTPbmy1f
mcDTXPAZSF0jf3CXAJed4BAT0ZRwr0nJCBID4WZf0Egp+1FVGU/EzPrDUtk5yorC
/of9/v0meJ0M5WDxErEUsDlAMGJtPauEOEn+nvI+0y3zU72fcjMnITUFpLy8w9nU
0oUXLwqsFpmc1mPbNxIlWnQhuuiBFLQ8TbxnlpwjR3pye2wgazIFeZbABMiIQ38A
H+23p1wXixA668N603HIRUtQayXerdPgBEkrOJmaVwM9gIBSIY28A+uvAK8kQhaP
bYEJUdAhPi5lRuE12ltXOd9Bx1+O3nlDplff8WJKLDxyC6sE55mU5nLC26JmLIuD
pwBuFV7+RVS6UICEpVTfLInko4t3TJP+RdVJn+tWlIJ5R0KKMcmThnd4trJdGAMT
twmddPDFoJ7dZD4V9XSMhnW7fxszT5e539BptPYEInfuJ4c4NY+LD7s87wxaQFd7
ojbeMD2pUvQu0+K9mqknyj07FthIb0NynJVzkH7uAHOn4AEolcTw+8QFtH2VIm5u
iOb9AdAYJLmFEEevaxIA8Pfxm+YdB29dRTt59tpn+VUO9YL1vtEeyDwgnZ5xvrJm
w9apyHPAI3YW2h5AvAVE0pLaR2aqwiJq4fzS0AtFygFoTSgoJj5+E3/D34k08PW8
HI0QZwE4Ge3GkCkFEpDPv7vqV9DwJeKXgLSWF6iCapM5YcuRzrtYADaBchvgH+m5
/DhVFseaIlzOAgEoS8tU4XXY71ldQbrbAyr/3RESiMmS98oNNGCXNO9ZnXTo6Brh
tkauzs8rJyXKpfiJqkC8nbEZpveNh/V++eZppMEQlzPyS0y6NEzphBGTQiOdnX4j
iU8nJpAOelF0U3w+xKxKCXDqLaCyXMoRDVT7am9+n26tB0046T3y+RC7lbtRuPKA
Jv2KnUoDSzZvpfEEio9j08pxvOQm/XDnznQjPWOfsvq1v3Ba9Iuz3FHmgOEf0ffW
XTyvUBmaJzrmQHWcfnRdTYO5eUPCj2aAeFdigWKqAMwNPmJDabCVBMJPqAcl0aId
snfC7/Drsn719uWKU9KH2zEkI4VrcMZsDCUCJfRZ7Urpzdrokl7mzHoLOZUKd9xT
4cASyy4LNauinW4pREWW5FocZP2GHuGvMjcXIWY10DU/NZEHOQlOlz339ljSpXRH
b0py/k2MQ1hB0vGl1DfaJmqO1aFbi6N2E4mWqVsM/lzmY9e0ViWmXtttJ3QRrpu3
2DylAM/xXjne6K1O/APpbvtXoCitkAPRRakFCoVRTqyLLJKu01Q6/GP76oLvrWbO
lWU0nQ2rs+lhlJL+7BMkyiGCsaNiqGh6fGLEGxYpsTVaePS8f7321E32AJIswrNC
GvcM7UwkdLKUFgrcKEiaw9u7nL6TFkIbwpE8xvOiCoBUFZ6AXBp+CwxGQcjb241W
mzgt1CEaZPAlxsfk52K6pRZr6NczSSZlZ/oZquSJQKJX5DdWICvtyROgIxhykj5R
DEcwXS7kfQ3L7Ya9r4pENv8iujVLAANpXfdDpPB3d/E7ERPvtH8EpGAEvW1091GP
MH39Wsb5GvgnAOVC1Ju0t91urd+ilHi5FtnV1xcSdgNBZDt+KQC2y+pHVEGZKf9b
c108icyWUMIdHzF8wsylSgB9hIEzcxlnY6+pIO5ONiwu2Ff8mvchsFOaja/lol3B
27dClwEk6sptmI7jT3vWfM7sP1XrjnjJWDc+4/8D9SilC5fa4aeL5hWyAdMzdN0R
iOEB0RKKBtz8uL9tGqT4tkThYabtbTDm9Sh3yTQLj/JskgMRw0z0+aHZu+Tlav/r
UUipy0UD7VJ6J8rC5KOSaJBI4/+yxFftrER5fcLve0Dkw8LuIrsuBIZs2FXfr1O4
muWWqjmZjNLLvn4h1somldyxSLIQLDtEoCjxv8EA8o3o1cCAj+KPJKBEj+ZuBCeE
i6tJOs++t6S9y5AGp+ZhE+LAd7C+7IO+J+UnhtHoxvrB829d8AVV9BrPx6IkFZ+h
QtSS+RaYPEyW+C2ULxJbZAqLXZx+cJoSfjKv2j+3oZfFvt6//8u9DqImMxPF3AOk
2csCkErZdVV0723f7jbzOEvgJGdA+3MwxiYwr7qMtCCNfMhZdd8E2bkcnPhK5fT2
qP2U9Q7PCu/YYojc+vzeq4oLQWGGNqaScOCHZHXt3HEkMMrFvJbLKuhV70xOrRmC
Q2IJJLN9nflPkMWF7Q793u6zA33gkXmxOh5UVyNtmQFDM83zzROkbePwqvocsk3x
SlSLnwo6lcL11KjqbrEbdFuH4GjQheIolMKVekefoUXACP1AHH3WExNqfxsN5byB
nYiGOkjWdpPeIAkERzHliLHn87ZONQ3V3fQ0/dpXSfpfm2Xerk55ezvmwxOri14q
RYRq2HbaSybtrhOYaaXzuNl+45tuXfy3D8WdGbN+WeYNOsgP63Ri6eFtGI4V1sCT
yPjnZ+AFFQgbI55/RN0+F+496Gzee3B2gic63vjRi57U+xbEKjBtk+m/nT/GH9Ls
znaRGKQMPNxABqgmLDdY9X5QK0HdZK7y8mJ1dUm3n/BGNZ8LAnCoQaMP4IThYUn8
NYPkoZvwhrHudlfSPTYsqFElQL+oTSj2Zut+drCZiF9CnZEaLLnM6YAb42y0+MlT
DQm5dwwk5nKF9V/XR+o4O4SICGFNTg1cYsi4usNPQcKinuigGQpBAMk+sLjt9bhC
uBoqo2Mjm41cyOkbTmOjTbwV0YN0vRt7+Tpwr+dLRIMH1pjDj7Ycw/8csiYCrO1z
yXDzmITzkBGKPEw+84V+K/rl0LFNAPMM4/RrP+0EcfDWpFK93z3CCNWdzCz5qNvU
Pc3yb5P4rD2sPzh1ljhm3MZIeEPwrHO6cjXpkQZwzGsefAIJBgw05xH6a1dzvGH9
8jaaK1td2D6zRFX5pX4YQmJc3wEiuKoobWwmXw13aKqsPmwaS3Uko3fhrFW8Uvpt
RfhpCjuv96KeX4wPfLAikcjQD3oxunxH/TOiFoKMe5yqVlWLfNuP8NAqRJG+a5M7
Zy9mqJjDUDvtU5mc+QsqbOba/PwBOl/D7aKa9R+ytAZzP0+oD6AkYljVAT75ds8r
/eYkkIrn6KF1Fc+g7b1sbTqsocRvZIJ32fuxkL3omjj1Gw9VnySAFHbVEb5Yg7vI
2oS//9k7fw/Fcu5y6opab+7ia4A3KP4ITvAyLL16xsAVZEYlk6HQYQQCc25jnjtO
DXwuwiCkV0Cg5onz/qB78oeBeDGTdd7wZbs6Z3xa+51GBm5ytseWObo7UjjHpCBX
3gKeavLrUaoRAP1WguypTJE7cKLmEG0xeVS6wlQHJgLCgUmhbOCMUQEHruDH65wq
fQ0FSrLptkxuhgOGVXR9NjAv+QwHh//gyyKVUcmY6WWix1VXMleR93OLDxV70Smj
85gWilY24M+yIxPKFMGdeOrJRm6QVEjFtbDySkqvWWquVeY5LrAIfw/Y/Ta2EH7s
PpvzayCxXR9pLqK2AzIp3mcrgUrYzjEj4ISjHdMLjgjyEl2CvSzAEP0MQp8RRUQo
x6lmwjI+fnSS4O5IJ0BqUuoWn1wKR7p5uD/NNngk8Gw7o5nJIxqcPHETOi7BxHSd
9wYvPRHkR6izsqDXWBBxHLNcJYLrr5hcMvQOd0xC71Ff+lW5X1mFGP86oF96OP8n
n6gmZZWNFy1UzY/I8m0sU/o/MVgSNN7Ttat3YWRP0A4kQjsTEthHahzZW4UDf3Em
ZNqkXF/S059xsoYTDwqpMuzFagattXsluoRx+mxJtwpi9yBcyPQ8swcNYpvoikS6
s5UbrTHRDlB3hyiDBvHMvDhWLuRFR1G011QsYqEEVhN6Le8lWCIKH961Fqa+DHPx
f3lOB9d1Xz/dqRgGb9xe9xwS/LdJWsMX1WKn+Isv5qXa/xJYfPrp2Mkv/MdyZALJ
FsX2Z6tK4rmgRtP06xzl2HKka8uDI+9BYMXpTjHqeZlbZslLNF4uMyTPxZRfogx5
dTQpLsLpDJ/bSVeWRBgjhglLMQzbx26f/q3bWRkFtjT4UpUfq3bsZAiPIVYKFhv1
0AlNqwb9J7E4fO6L0pMoZM1qWkyQ5W8mOGBJVOcw8utmSawq3PX17zl/01h/YpkA
oQ/OB1pImZpAb7m+yDNsE7xzjdGbxkz8DmWIqPmZpEi6+vWR9D+qkaHSFiIwu1gw
oq71Cn1rZO6+1bTYI49NHVyaZH0tU2v2OfwGIzgM83Zgo2tuftDWziJpoOPx4hAw
vErW0BJ/kkIR3g7c0ndhMrOV3y9/w2Gcc+7Ptc70BGD31KPXaOc27ecH8ccAjwuD
ooDpXLMc6W+XgxeJMl/QvMK4uSb/4tf1mYYdgVEKfROn8TyikYrk3Vwk2Xa1sFRY
86f2wZ2aKESEwc2alzWSv0zl1BDxp5aoTiu75xdXsyFgz3Bhm11Q0Y8cWKmhqfk8
csqnQCF9UUzc+MXVVHsIYuLfeDGIKR8PVnAPZ562EvRTtRLFS2duxDsudTLBdoY7
lUw1tNXxQr4xQ9t+bR2F7HDTazv6eH7XxwokCsVQUU/cE5esBlm5jtIo9gTwxJtX
6qgpdEYJ2vP6ZVbEGd9U3jmCiXZB0WjIiVOsIwxpMswPbU+9Lk7FB9mqfISYEhrI
61cyucCtxCST8UbCx2jcz00Lx95xxUlsm6ogNsOCdqLAjh5KGk8+lUX9QMQopDem
cEK1CAqxZhgnXNh8sJrPtXhWmqbzg5U6Nst2AMO5PpLGzUIJM4m2rdId9GcOjW6M
WvCGLq7R66t7I/DtSuPUksBfjrgFPMUGcjG7aJsgRaHlp4s+z/hUrHwsCpGv/3Ie
d/mvBQ8mkgDx7VKMxPjzdaS+z/1j7caXw4o6SyTM//dFCRCPbHfyhGq9GnHfVK3Q
+RXF8Y822t4/DhtbOpfqU1uev7ZeB6dhL52ZkWWkx3cBz8KjUtOMhX6+x7lMpT+a
ikJB8cIaX3C85Ebo7wqYj12bfR+UxjWeuM353Jz3vCPS45lWThh4zfeWNbQOB3pK
W27UkX4tF/cbaYUr0GIi8Y/2G1tRkHB+8eL+jbicbpkPp57wb3t6BfoLUBO6c7bc
/l6XxQNjTfGXL61VH8+9gAUpLKzCddr67B2nUHtcbyVVM3UF8aXh857lJYm+bpg2
dUCEszpnMTZL/yZILtrrxw/zADG42USduDAw+6X0Edb2OjqZEQv5+gpNP4GsFaJ1
3qFSC3ApigudSQk0tmYaO497OMt4JDMKMr7c5E0jHSDu1x+jMehQX377ENuqPb0p
Azs0N7T5dEOZXh9cXEIyPeYYK9pvpZy6gXHNMKkxcPEIIhZZGQfl7GLfmALG5Dhh
D54oiKyletwvCF3JMPjj8JdoeF+u3xlbROdz1eo5xP7W/0MkXPTzxte+Tp/VQLTw
ks4qVEY8q7PWieeJ9IXw9CwmHYuek0LFhj0Ld1ZC0ZFDaSY9AyhFrPLWczSb5Gvm
q6+KwWBV2+MkL+VmlIpEExmofHg9nLhpEgFkbgTlN1S5o377J97aghp8qQTVVSeA
2qCa/vmcoqSEzfyehvyFpA9MZpPDFcotNpD8iK0DbjjtzuT1hgJlH9KGX6xjI/aK
fP82TTxfY9sX9vmzPDd3MM1uS3pS426D8fSLQ1fLVQD88WAZO/am5xsF0Yr/OUYG
zcq8eeUp4dXBqYReihXkv/XaAYNdLXuYKEnhst/kzgfwmJ+ZNjqXKszLp8k8VYyF
fc7fU2irAvAkMdEDugsSVZh8FuHL8sPNJ2VkuQ/IsU6DyQ8Gy9rABV/bC9XGO32g
QzI+YlMXRCufuSaOTtdzxPYb9sLsVQhoJJCq15THgiFtMO0qSRaLtDlMdtH0/hYj
oY1s38o4etLkEaUKvbL85ePvY1eZXcZIkx+aX8yRbr9U8gUphhZh56Srunh7wsQz
cAxohwfz40HB2sCgtuJDHUcgoQFj5KIiPjvcD8A/FGrpc4FecysQGh1cxAgvziwS
4QiPJpDS2c3uy/uWOYk51kCinE444WlDk6NJlrirXo250lpOfgSVUy8gfP+A/6UI
kqdyl243Fjm2Ztx1iqUmOxGLkDlqEkRD5+7NvTdzFVn6tlQ1lpaWOAexHvNJxdVI
0NS5IIIDsVerZ085uQX74nrckW9eG29YK54Ipr3fHx/JGcB+WL7Z90D1mPUYOuMF
eJk1TnPPRdSLORVd6OCRInFQ/C72Sm19l3fdJ2WM37Flq2OrJiv3ACypTjwN2cy5
O0Bxw4CsDu/DGnNfhYA2E09t97HwVelkwiCTVkBs4PCPOZ9fBqGqEbBLF0G1rhuO
19x0YPzrvRDoeCESMJmn06dowf4nNbXztKCRGIh3jL0qk/1CW8y5eJ6S3zc5fOoL
e898Z4pVttAMuD9++P9p5ZWjaHUX4AYLerXfuZimDr8LkiZaxia1Gjmpqf8EE8dw
GZF61MtJPf+iC4YpYHJQlo0Tso+OumsIy2RvXs0NYraD7XfTX67kxWQDeHMYXQRu
WFxhtNIk1CkSgVUgnEhUgFoELhFBhLpzI67g7MuldeRtfi3H037i++hCfuahu11p
ceF2jexvVJtg3Rap9sFumpGBBPzcN3JOUH5mN2TMbQ6cSUMZAzokDZHER3B1eXJd
o49c4XITP8jJTaKVlskMfZUUYffnd/TmX3cJtqO66g+WtOLz1+K0HDhd/8XrrKmh
qIAWPzPMpJLvUDx8w2Mfcxf0Qy7Vr40ipgTfkbhiFJqiHz3ALBzJRpA95KsLJdG0
iEbh0rKT+NCx/a6yhriwBc8iBzluvZmHWqtEUgU/gNOQnbdTM70dHw9r9wqtyYz4
X4U5/5crNbWuePQSyDG9JmVyUfeWvrAIxNCeSSn/gaduywwe9urO2DGJWT0p3FkR
DnU6l+O93lK3cyVdb0ircd6rJIlqetKTnQoFObI6XkUgVof/QCEjA0Vx3WA3XWCV
5AJPer47WBCgo8LNrDQ24YnAKfojeL9zcRA6wJeBwsTJxo9gev0ONu+DWXj/78VW
vA2/TvYhq9MePhIzvTV4nLeNQUe6RdA8LAw7NU4Lavb3vU13lZyquMX7utyVa1eV
W9O/n3wWNN5Exzu53rGpHKB4B5no+dMailHSTdJvKegtaEx5OgagOEbMfw9ucSIf
hv9KnV6uEC1BEDUch0r78ywIsYuRtSx5/FJ2kh8WwI7xqtssgsoJ47giHqdcp75S
K3CWk7e6qR5bvoirFstXxw6iNNYIDKRMzTaAq6odcEgAGxiTjCEFahG0JhdyrtGn
pMZlpOIV0js68La3bKWOMKJ9AWxJ8bzN84umkxBdDcVTux2s+zKof0X+tCJ1rHvn
mAXjaBS8Qomxi6ZXkIFv3hElNdmWx2N25DzJLqkx4MziTJKdYXzdcHpIGqCu/pJw
NWczrRDtnYRLug29s4iUN2jhG8pNwfVHU/SdqN6acfrn4xFTBJ9BbOYcNCf8Gao4
Mm5g2GRga58UatEJ9EB51pCAnvOnEJy02Pb2Y+BqfVg1iIWP+mr8gzW1MLuWQP7l
F3sNXe2gicUHJVj3lx1kkKFI+GeBh1soNmloruRzx1fyaDrbGk2GXPb4nLsxZqIx
ndKpOFS2sJYxevusLjU9go19dg716aYKO0/p7Izn0yC5+bPdkhtCHZIdDexi90QI
Czrde9jBRxoL/cm81ThSKYcnk+gkUONr+/ISua/wQfp1AHMS5nK+ZJ0xdqHGwqRM
CIqNel//eAKmYd7DdRoT+DRCZz8LLf02XDaeljuw1k2QT9S7BjiZlBUYMnrZRjDH
1cTzHxXac50yJlwGAsrE4+AUvxWZUKfs520UIFxcZLMI7T0peMYBtgv3qd0rVNQY
O+QetmNAmwEc1Z9H+YW6eguOdhwNHPh4Bqq64dLuQ38EHxOdPTAoz03VCytkGh0R
MFqM6/paf8vhgTBp+T19NpiDW9PJqgMIPXog22K+fcxJBgUrMffqhxuePjgZNvdh
uGl6WIDLG1d701AmBhr1Aqa1kZ5tHLkBveL7ROOC6XhfqYT/ldmH7rtGjxsMU8Yy
NteMI95rAj7pkoJpIsOHijT2Q+VeiI+SNWOhrQlrdyppx5QU3McPdB0O7DxyLaGK
OhEsVc8L6jQ7ZXecAgyxWiB6S5nWR2Whlh74TZV9JClox9XKX4oDBI3eurFh0zc+
WTiUMj306YDfs7Wa39jpMUypZvURoq47nkFMw+ZtiQ7WiDzSKrjkkATB0vPkK5Cj
EBJ0AI9hZOdqzniGSvMaqG17nI6mSvQ/dwp18yFbVCzuPPIw7Z/M8IUjXmCVLLfG
jGycQAc/YeB8yQWX2JEhnnxufPg688YsT9HnruFDb/+HDNU9r6lQxg3O41FbMyyV
lWvWZHmBBi/z5hHTNSWlEG5dsKEMKvJuBMDP50vcizvuCnwKNxQJd54NAa2tDPP3
eeTzjP6T24wYIndc+AoCrELGwNAnKo2ZG8j6/8hUGzHhyJt8W8ZRenhjA5oielRl
YRan3k7paODyRLXQpaVRyrBPmii/kCOWaDPwIASpKH4jyUi1a1mTvY2FDzGUbT9Z
7KRfs8WBV4duTvSpUaCN5QG+2iE3SMDnR29PhN1OPSBXJiUuvPC+5+S/AV47smKw
JnZVI5135Uudxzqam8tCiUutE2jThDSPYOIpsoa6yI/2BEwXompWEfwH193J2NIw
MrSe524TAhpi2FWtwxGl+TC8wkSa5ILGEV6yq/LDyoCGd4IILqo0Y4Wx/4Y54jFV
0C+Ix7mwdtQn9fW8UKJr99aQbw85x1MrcEoJ7Ebh3QlyJGdgMp3eiXGG1s0ot9ge
IRwHANzTjmj6NJsMPikNmnW/fg4a65kmOYlsycnvfgN1TZF9IOCrz3UFhJNP752y
tHTkzUVIHe8sTGi39hB4O+CWfH1lazm9sFhfyqAI6W81C9/P7BAWB9jSwFCk4sh+
k/WbbvfnhsomZH0kQkD5Np9Y1nQv4n2W+iHQ9WTFVfQcn7P8z7qRhRoMkfcSb0VP
TIotjT1tTN1MkSODUKY02hCQ4R1jfPO8KrS+mlJy+vfHbykoTKwPebxPRSkUO2OM
p+XY0H1H6OoYlO/Dpw5tguSod1otFEJW+56S/y56IGfxyyMkII2XNKm9VLdlk0V4
gSTdBSmd3alYOMoLaIi/k0r1QkqOm/8VCW3qTFJ+I5QH9Wq5ILybb1+smN4wLCaw
olZGl5MPgKsRoZacS5l6GKm7DRXl1rJnpU9b5SHYU0eHcAIZzcl/2jXLZhqVa/Sj
glC6iCD77dOwQQYrX3knVoia7reX606La1r8ymKhmo6sRmCWV6O0+WoYlzei5nvY
Sh3Rxz/3B3lsyIVrteCXr7Wxa98GiOES+FyIJD2MeG9Bb6sv+53ktCYk7VaHmnoj
ipHw0y8Jxsxbq2n62Ac0WaVspqz6jCQK5H91SV1tpGd2KzO1AvSlHAxnvgvlUQcX
1bJUpANbiDtQPtjpb4AGbSIaIUlxO1BXLrtA2Ixsmmyes0kuv2HrZ0ClaP1gqTgg
1zAtbJ1zXIOjQyig8fqAyHnI0KeB3Rpj2yeIrKWHsnNXpQZd5uBY2RMqGv4ESUbi
PoBMxZw4vWaVpwQHARjvsXJO1M4lKs4BkCvqY3zKbQ2sGzvOZbsfFbYBfQMfIZqd
FN/0brGuD2X5SDd9OEQJHY/vQt2LD7xjPLj0AiE7dLLwzcfsih/FDSa0q8YLEkDW
bMYF8v7Je/xx/st8NTcpaQnC1Y+BdlwOdD86Uu9jSMKONGQdt22DGaBI/dlcQqZu
qL6Gt3Ww+oxol3+5ezWjj/P+VFOAk5VyZNmTil+X3r+Wi6TtO003NvTABxNoRdd6
VNNh1UgWqJ4qadFZdc8FQUdcsCJjCf+PuK86zd73f76vpQt80EsRKFGn19VBpn3Q
6senJuqCin02XWF1vPMytg0wSIkHGrEdfxn3tDeWp3lnJ4ogtS3FPOdgAHlp9BSu
S5G40E1O4/4ZFR/KJBhvfLMVag2bbV9EzOXtHt6roC9Z6YGT8x2rRcBAh+6VIvet
EDkpq1YsBv6sJLl+JkXraRb2ESLDiMLkKPKY/iJEmQt90KOruz0MoF9hc0FVduzE
5ra70wT7SjSSL+Bf3ZpcempSFd84j8fhwKzfXRA1XJ6TUHzZIMepW3mmGJgawPAq
A7xBOMaZs3eITxdiYf2PEa6Gj6EijuYabFXq4bWJqqCWDMa3l3+icCVXn7vVXzjC
QKPlCvb+/o/NIIjtusfyzymrxXjuKBIWmeBgctDYrqgYLJBiH0h8yc7FhFtHklM4
bJKhs7nvnd8SQYzl4MbYzjQh/gxnqLBay6Yev9cO7XlQYNGDHJ5VI44FL+xSYhRm
JoN5hmmtbVXaG1Icl7AGSqGgnWnGnNwdLNWNbUN7N+wWIzHGODUUzf4PlWGoiQnY
LmcwuLtQXOSPBodgn6hfU1k1s0HG13fTlLVUM1qhqDebbdECBkRZFj6HzFdFPAV1
ztakoF2Rr8bCjUTl4CoNdYgO9DAbM7oibuKaifHqyCidXYw++OkNHIvLhUG+mybk
Qd/NGbD8ovwC9OMxKial2v9rNeFt8u8/57GkrPzWWaxWc4A4wLutPm2HOkt7PDat
SROfWEDxv66uN31Q6kZXveHWgRISEndYTJPAO5I5et1+yN3OPNeqi7nWLCqR8qG8
gUewZYUYhpoKOuzhPkfkREXa2mUxp+9nOQyYp4amHgUN2tBeRwKp8D6SgSPH+7Lk
IaezOyk9EfvmqePR35hrXGuyn1rQV6nJapx7KkzImI4513lk12fm1q5pZq/U/3a0
xZ0G9t87VYx2/KQC4UBsVJVvG/U1eHYulrKrQwUwIyihLW+YqZ/Ez5FmO9XPDiSM
UXOwrX2mNe4ryFvNtOUrZco+yj4DRAZQ2+BD0A0tFyvs9olP+NkVMCwuTh3YyClZ
Fg3qOZokiUJy+RcWwNNtvKm3a9TDvvmf6uxoVV7cnS3tyPt7fsjfG0ewMh+XSy5n
VFFy8NvqofPQat2GlDFSCH4OJbkFppTipp3in7ZTkr3ztrTcVBDnKUojgod8cHEb
oO+OtSE4wHmVtAwMQRzrLrIrjCzZHvcl9B4HGvRgn8zrRKxlTrLXqL8wzaQ9zB/7
IC6ikv9ybd+a/MoHsGhiyMY1Owvq9QsZ19uGvK+MRBnUBW4ifdx2q7nAh8gzCD94
MS6Ol+upH2MU2kDinMNeoerTZGTPjvmBMNqPFOADo4i7SQmH/MBT1NblE1RFTuUb
IUZk3pC96IB0th4K7kOwNaCujcYX1ejElCP/v6z7udFgTJPSVLtD4GxkBpu6wzdM
h53JIwL3Nx6N0sD34gJhdZBOqLiG9rJRKBEBdg6xCKYzZNLwVJ6xAxjRLmPrRtbz
bvO5xHR4QOxltfkEbpUiMeTxX/0k7gDiKwojP0Hg9F4a4jx8w0Ecu0CMH9OreoDe
RxJhKyc6nnNOfsO0gsgGUIhJttFvraDnLfgZy7eLj4vjFHrVFOxrVrafLRf+KHLo
t6tfLMreyPYBqsI4ZKD2h0pZjp0xbF2RAiI15drz3774RmQDkGFR1EPxKaUO0TBG
luTZyeTaUaliPQ6rpBqTwheQf+Y4EqMYdONfuTzlTdYvsvAmOogS9sUdLGms6JiV
WU43xE0bVtencL4To65e6AD9LgNmZmj9b8OwlS0vgl60CfCoc5gnVaDfbKJ5LfuU
tP+TVZVw1OkLZjpCxJ24YtaOy9Y4gdg9+PMdG9SfwHXgCpB1myG3+OFpo2E9YL56
IILNEIlNxD1NgySiT254R2T+wt5k/VOKVT+MGdG9VEfgmCDvMv4UYb7xC9GooF5M
SMEsm9AwomZpZ2mL8Y9CzyJ9XOVIQ3HSbKU7OLdbFjPISqUMNdjlQKI8pKxg661m
/4hnc7Gqv/xzi/6WphUHUI29EsbFstwJyeR0O0nHXXgtWTmLuzZ9Zy1AAh0pIROC
u+9yJZj8zlvv8PtDkFJk2arJb/Z6e6jRy/Y34ISNoYTAFK0NOnHbodnfpMzzzDte
xMMT99KXnkHGBdVSGDvXk8L0PxeycttNvUys5PZMXCvaUchG4465YF9jbgQcmyHc
lGC8RMNzBiuX9w2BK6WawdJ+Y2ZRYLwXC427yts+BBSb9i9F9Lx94xX87AWi7Iav
kgCAaUu2g6PTz+FyoM/xWtXVJ6bEb4XlJt9eosH12p8HnxasQETZ5e0yVod7xZjD
9QGdQpfGJ5ofsB51PWWTmeARFpnjCJ2xtAEl2/nSG1bZ81yIMosxIoHJCnTm5E2s
MWpRens93eLswLY8OOPhAbM6IQAhUMvhFrlXuN+GQt9FNjmIVQgh08j6rPfvRfTj
Bq0itUPTG3roQEbDrXsZMcImmocJNGtFwoda1WMZTETXIxGmt5wLYNy+ystj7hqi
Z41xu2qs1pOYi9vfFuTdbV49bdUvoWrgAiWH437RML59ubfa+PttAJ2mzWHKX53b
ewlu1jjF2y15HynFGfJbKKVpDzwXUh+j9SsSBzGbDq55TDhv0l1ipCOma6LiVNL4
xKEYh8tMuxN+IoV0WR6J7/j/c4i4NHdYk3J3QryTFlU5JOD1unAY3Nq7+4OUvaq/
5Mh7GM4qInzhXUK31acHprPKVi6WOcHzn1rUF+/3CMudegjTBS3IPpXObcPU11Sz
p7R6t8kpDbcezD29l773Xx16JHFejaqDyPb1/96x91n7IFURH5yYycVD2MFipq78
uUl/bOoa5nmXZj5HPSwtrTDrbrE1UwgyVDGtXxZIgYNy9JGRNFgch8FH8W4//SIa
WLMfmmWDNhccrZwIcmsYRZ8aDTcSotMq704hwtoBW6NF+v8SxDV8vl253paRrdh6
hKcTW+QvL8a7vMd0g1Z13sLESfItcBe8l10pwxMtfm1k8r4n/BiZ27nh/OfEZhyB
NPIIwrRwCqpSPY9LzFclBbBIqQX0tNmO1qtyY2+7JqL9m45e3CHeKF7U9aRQO2AT
ZdLDHm6gj3Z0xde3OXByVjLtbCIT3c9HC/4iUl+mCgdRPg+ZKkyTjvZUtMcx9Qh4
t1Mrrvo9X5pTbh7lXgKa8lF5U/BnYongCOOR73gy5oSx+q3BCuSk8kBTXvQ6f15q
gZps1bNGRKvfRmotYFLNgOdhtPcpyXxfS63/jUFEGi4CDFOf/ggC/aD0FSzV1TCt
XE+zC0Yl35xz3hjjUzNNFoJ9FzSBeJds3kesyr/rOh8Nv/1p8ofFsnn5LpAnkylU
5I2LWDwcSFSQ4sEZlpQaLV25NZnMzE+0MX7+ofXA1Qj9/zYk4ShIqrOWE8CYKtAX
F9/NOXieCFBAU4byaTXH8O4rLhDmvRJzWqXRlCMndt6lgSyUoy7Qc4qixZwi5nfl
rkxvAO9j06iV2xqFY83N/dw3LKuZeLWNrjZLwNPgm8HKmzWDad4r+PZQC4RkgKRW
drXAfkqwd2/n50BuUVBEGv0ddJjyJ4+/ivvigIb16RG0NChG/bZtEVYDLbKNpkj4
atmJwIrf6fGiaeyZmx5oLUDwyZoe9uGuHP6Jg/lrbhtXxKdgj9QUtbM0Ydq2Gxy8
Nq13Q75BP/CzRXOKHPs9QnNdUu3RSG2bxP5Tj9S1fKRljU1+Yts4mN/3byV0x7+/
QFHInHRfm8ipA28w9mM1UWz+0S355P+nzRUqGI2UJcaOz8RtQYSPP752PzjzwQFM
bAW+jSl7jgmfxpkuV/dcHqGGKmjaoyKj01wEO0l2dsbaBNJo9KSvQaPLRDfoFBIr
J0rGr9JRQTZqnm53z8W6TzfdkZB83ltguKvHsXC+wFbMB1HjS882pX/XfCjfmXSA
sxIy1Vp4Gg1IbLq78MSYZIVtzJtv9hwO9VMBsnJBOsKhNDRp+vJGTz12r1zh7HdC
/1yOYwajJjdTx8GYCjRA344roY1GkTqqG/sqD5cbQiwwVIzsQJcSxYLsYVD/SEJK
P0Gca2Tkk+hsDk9VPJqTn/8zM5NFnHW5CSClQO75iuVNQ2OqxWG81hv2KpBryYce
tllmLTjFbO49+wL8sHOPmjksxQM3pqwyJrL/ayoF8Bv7k9EMknMGPJpYX/Sn4g9l
sUNG0s5/GBSEJ5KAemUj6t2hGu1/NYMQPuwm9HSwGIiM/pK6DqpLI4goTrtwe5Jq
vqw5uEuKU1o438Xvw6VDB8vs8xIMSZf6SxEJgof/fnlbXKPiYIz0UcgUS2b6BdzE
zBK+14FBKzHaeFGSvx0q5mou9NXjGFxEv02rERNIX4rYx4unDlZVGOgpjDNjvFgQ
CjoJZx5iyCCHckpJhw5wcIpy//QEPcLZGkWxrXpL3AkrxiPkwyOVtNVmiGTn8Asx
FsQRQ9IBX4ZCDweRLMKQkAZgSrnzH/EhoB/BIjpIdV0DS9VzW1mpETkbyBO4yBkJ
zvBQXldtUey97Ju82gY41NRSavNdDXNDxjzL8Kwn3Q+b7GcRCL9HOWSPEATegTBE
7aFGuDDNfQJI6CYmKnH3WISwkqbsqlqC/2Rp5HFXh+G3pY94T1qg+r6X99Iw9x7k
PJjaXTs28HZQAZBaFNWuOqDH7iXyEMfTqYc557LaE7p1HWnBtdSHPYM7v4dcoD92
5H7Ux82qfKbUvKx2c0+V6Thyqj/bPYDJV+NecOjFn+cYELqWqiNiqw8alPwgJ4Qk
byZeixqpKHQYa8eaxwljZxS2RlOjFJ3pzblFYS2BUIBmPrBjgHKMIWARWK9FlRb3
6FF+EpgNamnZxoZElM6IVGI29uIppSrLnV8QkRXX4ztGz0UR6fAaEOURbeaEqKpN
AF1ag/urpixSXp8hHRHtF4G+meLc4h6XfKIIt7ZSqL99wY03Qn50pf9gd/utCEKJ
TV4CoPrtFCTN3owiiGwO7fxa0J5ZzByt1+lWPe1+mxJOrQuvED+W01Dkf7zg9Fxp
GA0+1RS5DjyIbLT9YdAB6XPTOy8ECcifpECuDl91Sw6PvvkWmxiw6+2EEAh2/fhG
qDgf8uX6shgxDx20MsgvxcXlcs9wnTCrC38cClAocofUJd+tFT3MekzWs5iVOn8B
xJDU7ai/tJKhHOOPrBe8GnfQoaxFWMZR2lx3esiQ1qEnNUlW3ufoF4OMJ632uDAO
4gu5k/rxML5wALbrMxFZH6mZ0INvqSgEf8oc8uB9w1bWCP8YcjqwymiNAkxm+h4z
uIrQxToCSu5sFHwMWQeN9oJEEWXiNwYb8Mzn1VUqSPvZVbfVH8n9g3tF+F+YBYih
bfm0jco76cOYXxo52aJha9Wd1sk6H35hBwuc9XvY1DtTCpaX/KfmgehGXEzaH9/H
bcMVOdJa7MlJHsjRT65dcNeTjGYMGUvpWRUfDYp/1n5ZX4zU8kcNs6d7MIQOzfUh
0GnZci0guiplmaUXSf8IYwdeOUoei9rCoiiYtinKU+TBJuMIELrjeI4z/nOpfBPv
Nn/h/O7MJq4XiHsqmv5+gUVSSp2UbQMM3nKWk6TvEwpGYH5YVIe4KrrJSyRhZ57N
t4CuVnVTf6WlzEe7I4HiohtWckK6jCelOEt/EdY9I6D83pcUy+eRFeraRvWQmCJq
y6OuzxUPkXHOIvzUAb79QIagnOVZXEw1iu8EBFVa3SK3s8ToegiceQSY1ol6/ne9
nKox8OPrOCNntWETzktdIQcvGlrOm+zyRxBlDcx/AFBEAtbvS2iHOivxkXv98TC/
jDgCshizEJqfCvqCf0/FcMVbFhZUomTRqu9L7vYSevLT+XD6XM6BJppXSq8qBTMB
iKFYUCX23u09naLAv8wm6wB7e56kZgR1AmSi3NV5Ycg75PHh6hyepi+HK24qIyWv
xtHxuDHBozcYA9YwOY0A8CpdDdRZPIdS0qxfbWUvfb1EHef2/krodKF7YWX9zynE
gN0bgSd24xyj1VC96fGKlVAerFX0ufIDFDiKiPPVq9iqFwdZbJM0ijtMAWRiY6UO
9gyofdMWl89dTe9lMQymsUUMlCiJpjulRXJ2zkUh/akMj9KWKwiubmVcDECynYd/
uOguNdlv5WZrlgzvk0ep+iU4VTX+CUv1BlXQ1u9IYrTuzZ0O7cNLJ66HxowmmehK
l7Y6ImOZOHG+/cqIx1DmaiEGzIWPXFkr3aGCmlgWYCHHsiL6eYhgbtx53qhlrNPg
sMxdax6tACQdZkbJTP2caihBXp9TpBk6R9vTM5UdnNrg9PZNLKwRHvS7C2fRYrdV
29/e1xMaxOHx7R4LIumr0eeEvsuc+GfJ3ux6rsYNjsxC8n3jbj/EmSkvTEtVrkfN
/LbgiMHQNzgAklJufs3cAE0N8nmsBmohATJuE9dGZnwFFwPENNEqfR66dsJrv+N+
szM5I64MVwrEqxDQ5ruUM7RxCdIO8VnQ47OuIy9GO7z33twmSk8GonnDV1ZVHpVw
wWtitsk+9l31o5EMtZr9/H6VtPDZqrJmTEZR746NN7d/cqXS7VZQ18o7txnq+ZVB
0EzaAe6mF/gIkvfAG87ahp9zUqLhD3OW1vRkBTA6mL45Y5peDDzFKeLv9u2B/xHj
w7FUU6IMHkTgsywYKIppPPWepcYRLADNEf2wQePGFSzybjwjrJM9xOlZ5SXae4Rx
Vnt/crl0OO0Li8fDFeyYUkcwjq5NGlqqf+z5cGm/V7g6cv3j3sb+95iWO+r1pJ7q
UsOtxET0lqgtS01vxdTALn3TLpCgJGioD8Qr5Bfc+ny8ybVNeFUvh1iM6Yhjo8zy
jP/22SH7BTFGYUvvdYJGMgzCZZav69/6mOHEl+iYL+KdYdVZqloOO+0+p2zbBDoV
hrJat9mgrF1ZDxXXgnGPRQOgd1kDl1+qS0zZ4buav8a8a4vglPNxzQwCS/kUPB3P
Uai/fdmfNCfUHYSfpCbo5o9XZACgNlFcxgTkbVlywDIXgTlX6MdP31+1N74SHlS1
/EE38cVVR53/8yygFckpDRQ9Eeqwfda8m9wZYpeo2/nC7epl9yEzhrgghMiUWjRW
GFqB02t/EFgFZxT+CHOGHZa7LvrfXNNS/NVkq5cduq77K9vsxid9LNxQI98j9g7t
bmP0fEXHgF5ytVccpiuhNidnJCoJWkffK6cy9be3+vxGvXHLxq3njjudYHMy52WA
OC993R4wVFGpAvKEND9CdUn8v6XJHuSAstrWeglRLt3WUcJIS+/7zAcL4VcDRp2C
QDRoLJ+eq5HSXhF6rx+2BBQM7b0NubzjWh9+1q2fk0lmtTTWWwHixMIvmnz+mzss
OZLxWd3WX5ixdLB3HfQ3WVezZjjYDihjU79fkfBkLKBvGjTrNsaGcl+Y/JkhrtPs
VamXhJ+pxHVX8VtpN3VzjbP37xUKCCCkGcDWabQbSRIrnPkNbyQKAP4Uhm1UjQ2O
eltS+DN1zloDXz+6dZ3uxWQ+ghAaUBSZS5r4ixJ3sfm+o4ELxW0FGGflYXHmRh3N
ux8JZbvkUjye2EK0pNRf0y7KueWV8Id/rn3YsdfLNPurZLGJvjOoDoMMT+CLNX1m
uHmu3JsTlgmqHkR4NBJ5EBEj3P0CrKRIyjxaUYz5J9vMObtbHKlkmADUXxW3zfKL
79OL/7fGCRi9akgJeASY8mdOXeC4t8m2G/Ly5ovZuIGs/D8VENNeFxu98jj/CePj
AJP2QHHe7EDVzVZdP6Jqv3MwpDwQdnrJOB3fynRL23I9RESeUOYzVtDPkMfaA36+
JT42RBHBKUGpl1ImX7psnXpqzHXVxxSrWdER0TKBQRUq1pCUl9y5adypdE1F90Tq
29OSYaRqVLsEps+VfqHAP6+MPWYE4gNzhqdbfud98y3xRvwBroFbQ43BB1ualsfb
WwnHNBBTNgNVhOBR4uz304Nl/WwVJqXFQl4y7L4SjqGJilHzNQIpJGBx+yXifC5E
rCHhp3CLr2yTif9PtOwqlbeTEnbPY1NRC9Odakuw/BzogR6/vAsIVBYuAat4Aask
QH0/XSZgtjUzpgHl8xNPlRBjK1w8ZNQoVUPaOO+7WRHUyadZNn9irN8Zw59BD2G+
cK0+0J2zsLuoFSfc3dc33vzgCeaSiSkSp94dj8dJ10ly1+ivH7kar4e8QDvPY4Nz
vGw+zViFCmf2U/sTrOTpPLTXzFMb0qdAlvk2i8HUxiYfwE1yZNuXrLfufBDNDK2H
+qyG4Fc6n1ZQiPTPoM4DX+KD5Th/YQmacYESrubV3c6qxnK1Z1LNcVzsgGwH+qk1
n7P+C8oVmj6zaHDYajPYt25cHr/pNa+R0wxiwj1mj+WEs0BHMhxOXfjW4dM7UhUN
FOIoqTNruiHt5wpYE1oQIXDEV1QMCU9Mr14qngJiNoBTA1wkRZdL05AAvx20NkV5
PoGNv/qYsO/xpHI76h9gceACzWQJkkgpzH3WTkwdx7nf1nUuTY4aqT04hvs5HEG9
lsrqGTXKubd27WNxcjqyUJGLrVqwlIstaXHOwRX4AMkRU7HuifbCsg37Quy3z8jC
XYJhhjuxY6aH+dE/OxSlZvzabh16MkNLaHVxCyVsOAtdmuZAaRA222OsKBMlgEma
socSTCPA46+usfDnxaZ+py6JVZI4GnnJ4fuQqcc/pAia2geOxKMVJOPS/Z+c0DeQ
109xIYWgv3wpSn8MOc6wyZE/4WI9631QEq5VUWOKuAqHho9ieV8FwC2gd4mo82eI
6pEGj1iuMyA2jmiM7OIxwEy56/v/ADE3KQnzT1N9f3vtRg7AnyJPRYJFcOSqqGF7
mokG8lApNRc4NQL2KhOi0QxrCDo6GQ1GPoHEVvGRdQl5tC4tA8Gy5gnClwb6dCdf
V8dapWx210KMzf6d+Sk0wxGyW5xIzPtCnbl8VxppbKneYvmAi/7BZnBBmlgVHiP9
eQyWKRFHs846/hq11CTiR327qRsuzCrnRs/NxjWwxcDRN0K2UDXW67xt0wqZKgok
5j4zTX/JQjfB+wsNHPxhq7jtBm8S58CSGbc/FZfm8axzZUKtDjRrsXSM1NG3iPRo
R5r3+ICveVABaTn+6yAcVdWlw6B97XZo+xygtb38lA1ZynS/XjwwjoSMwg7NlMpN
sxQEPkHXPmenbaUK8LlUPZ5ds2jzslanRwPOP2nzhiWFZ9uyYnsnnHxJ5ItQgNdy
cSUQwtFz0JBMpWT5pdiGOTkhNYy5KAxOgbSbsXVOrIxw+rFe3TYvDS0AZOxYqXIz
Fupji3PWrSnaUJS1Fsyh6vfoj0DLwiroZg2RxkuMFriyPZicrDPMM/IiLvVnw1B/
vVSTCZmjMnCrDYjUIpmN9snh3W00E0hoDs4IBy3otk2rBgPIsUxqzvpO3XhIkhBt
58RX9RdOJxMUM/CY1+f9fa9TvM6aFviuQcEZCrnVkT8jM4Ym395akFbY5CnzLjNI
jfKZOqR5+OPUnPZFh7vFBXx6XiySTEN+keXDVe7Uoivv1G5+ChgTwX+/CSMAfXiS
6t0O26+xwnpi9kazNSmE3Vv6+SSA9T0bPNRs4SlNcIy9Mg4rotLhJwwh8RfB5Ejl
fqCzQXRCo0dIMGpEh35nUymcHqKy87QqnquvTfvgmaIM4RcnaXo/1gXtHvdoUju3
KoR1617vUcVaa1L4vsul56W6KhF/iw+KC/PDBLf6kqrxXVaXUL4pk+fwEKnrFhCu
12CI+QUMuuoC46tAk9E9EcgKgpYciLKaw2HwRIfCAO+w0GOA93Pmd39GjS5R4UTz
qXKCUs83fPYfu7X/lHxEFlFRpGxdgQhDx+kq0EsDafbQd2Nihbo0R3rte33Aq9FA
JAeCPRu8qbBdC/Cdz05efewSfhUmzDtcJoFYjS4Ze64F8NGjZmGSjZFlcK0Ww5Bg
c94wzg4giOjH2pSd6DJkxZjP/SpmlqXr5lzG47SVohnkFqzHMWgtNjFf0mTWyZMg
YDRy0opRFiB9F1Y9IM42kd7sAzLy9Cv2U2VoK4ULjW+b7WrPvLJNl2qe+1vBD/d4
5QOtORSz2wQsd7HhSOO/HlIZjxUqc8UXLxkPXdaHPqMe8c/p/7mAmORKmpCimRVa
Al4cbpI4G70mOA+3vbBMb0w+ws3nkLF2rbZEt44MEOGNoaCOuJ5yjBYXRSqy0uOZ
6biIIhPe3wvaC7ddgIXiELT6g8kSh8skQEMv5Wy4/w6I7otfGFebO+dz0kPwMJn/
EWPIqTpKq7eWCrlgodnTFrwK1DSmMvOpgMoIHH/oOjaNPFA8AHW2QRGlEF4xtvty
iXVcPYVNnK8qqz1rluLRhyJIfaNkgr+m6DwVLnF7UenHfSasuVbUERdrm/o2XNG6
FQAh5crzhzr+byzuLZbNECC96VheDAbjC65PbSK+iktFKl+MFyaYId9adVQwvG2y
jUT5zxPQoC4n4ThVENyWD0kHUfNKdm0VVpSZaVpXn5wYK+Om/CSx0NZBTVbDX09l
15xQHWGu8kgJBkS7eSBoHnBK5BynGocdVtNJSNeGAtKyrAeEl1cfiUU1Yzjtk/Fl
bxXd8k+svc+L9MbcbTl77rJ1+Y1WteQEzvfctnvfyJUi4WdD/oO5d/We9gmmwkOM
hnTJUGA6izhMTTVWeufLZmioi/0TE0yUflJ5fqGzrJ4hab+n6PZYAs53y8AbLUWc
c9Z+zE043mNaQuhbP9DsqSUOGYzIi04tIi5/xb8AMd5le7Fbdi1svpmLp56cjwAM
zjFOjzZSeP9Kr3FsasbVlQdVT3U3icF2NJoXNbtKtfn9Vjs8yBoG+i18N54wTwBM
EVY+nRSz97NSWYlr3l4wzVzusR9GdZ6ALQYl61AwGuOl9FMP+cTtxKtnGAAKW8cM
lpv7sM3U5+TdEJJP4TADl0YNKnLbNWpEwvvgyPTjCQ9HsdEYreMQiM54B552z1cV
oPsUZ0PIRGUcvLV4eTd8rtlAi7t2SexPrafgmfrGWWuRDLQ7O1iRPXCmsQnHgIh0
/CCRVR2OVnc1u1DLnjerAE1Nyv0NN+CHBlMLCi4RcEb7p0gLnVpXhaTE8DZxMsDv
ZEGPRn4KhcuKjb90GexTzcgVMCGxxlurmm1jLyjt8PYCE2kl4NnhHq+wIJsHV4H2
mUcWxIzn1z+e+ZBlIZZ7p9Zhw6iVUeL34p3LkT8uwoxJ7EaMpyy/TjWzDLqlMxo8
B6v3FjQCON+DTy0uqSncwcbu6tD+j5SdgiIywNMd1LIjtMMxJ5teARNUi6wipuvg
7PiDt6Og1pwM6Ix6yZQTEl94pGMntUkBLOvH+VAHA4gaqyDVoAfHdHC6QxNwrXZn
kg5PjuXUTZfRlZVpSzx+eP9qUoNNcQwoVRPfnu3mUEVhi8dRW5gBvhKrGeY9Mwiy
/VoDnw48+sOVtyls+d764Q1jdW66vbqL/JQaEFh9xn0gy0rBMJ/UpeWL2r6AnMjA
jdtQvg6PUkv5gMdGRMbIzDQ/JrykRuSbzKzzL7JaT5i8fPxHTp2a8AMHKR+D/FxP
qODY3yeXRNHrgfHeK7c+JD7z4/ooA3z2j0N7kFK5GJlIYrIL29dLXV87Nc6Y4Lvi
jGcyOdJSb+MKqKXx2lGavyZi3l55U1APYD5u07BSHoVxoHHRQ/EQQZBjt0Eu3I2+
rJkRFAXhCovvhsFgG0rLiEN2GNRIVPQVUbSURGWg59IhGRaFFLEZqaqX3temMNra
htTLS0J1BdodmT8TsDCEzobMNImTb87cuuew8ShuM3+8L1Nrr+6+HIJeyBY4mbe3
laz1cwUB42YbXG3h+p0ZHuf8QQAJkmXXNpK4Y5u6qPIi1L+ZlDXv+3ZTvNTD/yiT
qQU4sWkhEHcTuZGS0XExrbd1z/mt/9cUR7a5/iujpBk8nvudDM84LkvEPCA9lwDB
T8bIgERkenHCuRO1CC3vukdEZ9Vc3tG1kf4fykryUgVQFg8jpqUbhNX7uE+Zs9iH
46RYSAP0u3uhYzp3BzxKKUJryhym5hRgK6bHrj484iitulMSogIOWyHK01WFdt4B
S63w7FvqBhm2hAsxGfe6fPgP7RLNycnApVxwux0Q8Sq4FO6/Bj6+XgQEmtcRFryW
6Ta9iJ3QB7mNDyJqsgWX9CAGeI0KL3Ea5UwZsXx8ovGIdfyCLqfv7uTUwX9ARm3V
AblmgEJIAV6CagFsjyy3+rJTdDKuyGtyNm1memd5RB+0WJha4pGwXBwHM+2sFtxJ
MMXmZbXbJpI8xPYt1yAHMn2tfrLGvhwuqkNVUO2maOyS56iIU4bJZT5VGUWBXtoF
vdtJ6evcRRDOf7s2PWo1P2i2Dyns5HWM72B1o4nCQJQKbcrt2p+HBcGIK5SkuD1J
k0t7HB0/bcUBOHqiOGbu2VsC9g+SWvg8f7wbpl/hQjWHf709PrVuW8zzEZkM5ryV
GW63s2wtgiGR5jgAygnmoj5SRkr4vzhz5bECKuSZ+tCWyDA6apzLZEuducBFh1aK
kFGjMVws36RCXbDIi7fNmhuiCOSqFQt8bkNXVQDc7CckKrfQGmt7IBFXwz6l10eg
Eg2sY+AUX1ormXzlVkyMI5pLHwL1bndd6+xkxIRDsfJ7YsJBEz8qDld+vfrKSk0g
RFaAumvrn4WEmjAB67Ec85GLticquNkWDlBTRKo7HEZlsrp9bG8k2orG6wNisY7T
DKS6m9LaVvCX4DcXTGiNgYZSq2geSjUz2mUkF3DQKX3TBwjzU2h52PuBTuBYwQLI
HEJkuzsub8fU0xt6kJKukiWvJ5wbH+NVWSzgaSdlD2FhbRRntnVCsC/tAKwpR15l
VoLkQgUIhEKgPGy468pIxkRguzvd2kSWVbNe+jBDUicN7xz14P1ynLfxzI2FR1B3
0Sp6cKmBVuLeH9Bv9f8PYmH3jb5UVt7fr3akI3+ScUys/MDaO16mbQafwCZU8LfA
RoAwkzlGA8fBUlaHGmqYpxNKAhkSasQO8a+W1THqUANBIfP05Ki7Mz8Qa8YN43yC
A4rP0t22sqCO72zAI5pQizJDuRvGjqQwmkvSOykvMs9htb6+nJnBfjyjx8+A5/xu
CbeiZZP/KIKiXOz+S4Jn2yAoj9a1vMVAJL7NgPsZwPEaDStdhy2UiwNDyVqqSk/5
S9yPtXAlICjFWTJ1AECnP5FfBrEmZRdl2K4Kj2vMoBoWp1IiUXE00R7URVuQ4CnE
hzJMEuWXIvZfKkPLoyrYV2t+ZFXYD8zOL4YvQ48scQwVW8K0adlRADdSuq9y4vB2
A3+VY8ljvz9buyOLajy4BbOsbDLK0NaLbimdxvXkAmiKwtCm6LpbkfODEIOPm+od
G+Tuf59cO8HX2HCWr9dbxzgU3QrAPMrSwZ4Cz7VUjLmdLuIYJ4sSPjyXflk72GjV
H+RCUtCeer6j35xbGyiin0hqiR9EZ1xLvWKq2vCJ7g6zNltb1pmAwl2CSYhqEdSo
ae2nRt0buTj24o7gO6MpbcVjdk5ZDvO3OB2YvekKmRg/CtEdnrxnPx/Cm7oWI3oc
zl++lqFHcbORajMQLFjr8/QE8nEi8LYHMcSoxp6M/GaJI639EFcxeOr13d+KssW8
c05cUYkm3OjQvwhX2U1xDPp0luEe/fB4kZ2dG1yeIEsKa8DioU5McyzHbpVREaW2
DnnACGYmPXiGESIMZg9VAd/GRdVFryqKr94XoAKB+wPGW+blusmaugsuCAouA/zL
5BTDFG4B1r87S5wgxD9aKyPEOZaHKTB0x6z9OF9OeQq7qibtpACPX9cd3WgSwXbe
K53VBxa/5awA/Y57u0Y2MEk7qkdAcVOZGtMQtUSLcpzytVPHApgAW7tAoRusmcXW
cU+ce2MOL5MoUhrjvI5mrm5kNX/nHZvONRIeHja+OV+meLMVAYHWV5eovT3uCFC0
+xhXeY6mdxaN3L0OjuidnhaWakl3JAwOi9N/vKoiBdKGvr14hS/suhMD7O285ESl
2BnfOvlhT1vfHO0WJLEbUWNZlqW2PQ8E2vNUNnkftFnDCHKtGJ4nXDljtPSgmWYu
ltETtdtzR9vypTrdtB6BHxkgyDtW7Kispr18YWoXnmehGJFYRKPfEhug7SGRPDI2
AjpL7/qJd6yzgmdVLj9XmcfTTIPxdO4U04tcoBxYibIsBclP9w/ZDrneyKSX12iX
Zv2563QusiUDIk+e9K7FWMClelSlWp4d5P346ujVkx+z+RgCtaLYx+KHD+cRw8Ic
wzn55UqJ25+2ZvkhRN4ThTXkPHZhAtH3x26oyv8+8+6+QbberXvJAw4Ys1J6bp4U
5b5gmI1kM2CLEQSBpTxv5S0akTR3yb4gw5ZOUigMOo8PykBQRaPyqaWzm10kNEzb
U0GAjsbHPnJWjH23MzU0clZMmAAbq3gKsqJnTUz8kos0xuwMV/Mtt424z6gwaFKV
4ER3txH/W5fRiBQyayPf1GPLwRu4bD/N9X8e0QqBQS19Ln1KmjrfQ82BQy+FBe95
8sQQp0G0vdKYXd1DyaqxyqONK5gHVpHJZawY9z+kJTqsMg2bA+ceRSolt6f+iDeP
dwOZhKjzbvQ4hulm4WuuY7Tgfb+rlkQJPzDlFiEdrH3re02M9pc6TJpPJCWAETPl
BUwvdB/rEj2fvHyDK4ec59XsaH4Uh6SPdl33tAQOxj0tA75vfpQtuBJRwu02kIal
c6MyW1jCfeDmduWvAJQ5mE64aFTjUpzXT8jkCBZRFQ9GDxpFhShxz4kmLZEuEyht
z769hmFxSTyeWOKNuGLpMh3fIELCmVtbaW0PDmNcgh7CG75SNccyXXFOSEXRpudx
C0acRQ1KFKmG/zhWgsT2fw+q+e5VcPCtpmydcSOiOMzvV0K4b8OgICY2C7EWufo7
T/0CAGQQIVJu+J81sagjkd4P+nIdMjQBAmCkw9erHYfF6ublRNOjW0dFdToU6OJo
hChb+n/vO21XXru66/tlz1BoaQIOlSnhx4ONHBOU+TsNeLRfN+3C6kE0STmp/WMD
4HMjj4WQ+Va2J9UvJM6hMrlOlBexjQ1e40Mj1FDSfRZ6g8N4iUHqOjH1vqkw8A8b
mnGZsxpGUqJ5GMTtro1CQLSdh6Stk7E4o+JVJLHYJ4Hcpovee1ktDoWvftYk3vwS
v4mw1zZGVTqqVNYLkrqxgOGJt8lbBWpamEvFUohptp+puZdVDkboPxnEDnzQN/g1
DsqoKsh+AvR6BRnK6fPNyqy7woBrIX0V9QzgXwrkw4OBYniuppfhifCKCUCC2ziC
dqfdbk0AffvBIaYNj8a5tcIp5wlF29TBkR+wNN18fIZ4jxOBOWwUqV6QAn9fANv6
yf4rnCVBRoOtmRRi1KXX13GJb8NfzQuJzyTWrA3opnA7OqzsdHQVushW+t9UNFdD
gGAhe3GLLilrnb2xJXhYHadExW9m86pY/4/pYe6R7gUGdawJbpI4kbC6ycMQPT+L
tGyejkkKYSqGVkila5iTAXxDcdDSRfVd45RS6Os1worVdeUK15/ErwT7IRhlBJSM
5aBcZd1+dwzax1ZdX3PF2IwP71A2U7nQFeVE7BicYZlWIyllRFudR3xNxefhVjGG
dY5XMOZCFC9Sx2Ew5xpxGGmBclg+E8ToObiY04YIjzdAlHy5DhhA4XuHidYX5FKx
eJ+TtBvBcY0OTJ8dHaHCJ54h0ZT8BnqaTUR4pUF9t21EYQAjZbEbQSK97QaIf3Zw
+/CEmNU0LN3LzvVOHzvKS9unSzC258YlYBRVEqpvpwMsx5lOJzVcxW7KC3L+M5ve
74OOTY821AzffDHyf+c4O2VJpOhsm6KNoVb5tOMJJuHJlnS3RGGpBhbw99h4DoOM
x5bMlZGaUrkW00OuxAey1aAjTjn15t3qh9j22hq54hvShiUP0yNWPg5DbvmooKen
G6dTLOgt0haj6F9Z8G5Idl9vSnffHtQOplKYPOJQ1yubDRKOMm6ycNK2yrDG8Dt+
S/9yJTZUjG5+0rQCU65/IR5ms8zH7YZal/k2PBLM+QDJpENsMUTt2q288/yQbuFu
MNFpoI0EUw9Sn/28zu6lQMLKqibhP7GTMTLDpuPMoYi4a6Vqw9NHTO8xrjJFL5Cz
XoxQFi1RlSfNvZngrV5VtDSvQymysWIKQlzhQdM5/NpSuU0+G9Wx/aK8copMbmS6
IdW2TmwFD/ne31QXdOcnMq8bfDMizDTW2EWrTOTbuA2LThsDgUjdl0M5d2/h8bvz
YmgDGjCbTs6GepVfCuqipUd8YpBTMFBf1oJduNVqvaT4x6Q11Zp1IQRithMCdBKX
yT/wqtwtEaCFWk7kqMy51eJN8ek8TtETQJiBU6ce4s56KjyY98LusXKUZXZIJIC6
cxsDU1VnPKgWL6lvpoP4Ai9S9+IImkIrNRMsBnXYSAd+TwtA9vtjsQVhR+9we9Wo
qkdqDI1lZvxwra4TFR/sYDlN9F2ojVEkBLCIhOY5ORw5DE6LuMmIOIv7XMBKaRDd
AAMpgizRVjax6y3kiWU12z4wJzmzGkcNfUgSU4tKHUhrA0mzqn4gkIC9rjTAd/Kk
+KJKxUy+xG2clgAmtn0sCok2XmEzcGY9Is/0Kv+puRnXX0IZSdHURoAzXw27QdBw
+yPFxQq5D95kfKWhCfAIWsmnMjxswweHbbK3GsRA7r8hW4AA+hYjE+Psla5C2h3s
7s7prCMNV0j7524BTSj9rncQzUxrcYomOlniZcZWpfueH3m3iRq4PGpsvmC1UzEH
7JYbRkbtrXp470g3P+SWEnaHPcMSf6U/FJhXkzduV6Vy4iCQbGOS2/PvJAzfmh1j
NB5VyVvHfmOwvzknnCiCdpPGcclSlSwnxsq/8yxp5vkiVPvY3VYD6ouPRVIpye9v
QzZAdZPCQ+T2cIIxg7vgFuoyPsrR5dyBhGblb9kjSQ8Xt4FL/PxuDO20QFIQHh+f
rPjrRGV6ciygw30u0UakESkCo6LfIu2HD0d/gCrvdYRcupTY7K4UUmXuYAzsGoPA
Ms5WnZ3F8FfIkeyx2bAU0QP2sfYqIX35daFpSZigdkqK6aJ7k3QXiCmrAbeS9gdU
PPcg/OXJZmnBOxSsQkzVj+oQH/E2EHsBPo8lq45FiMnIvjzQqEzrEcBPxifESDhG
Xe/+RSbVNlhhYZaXY+lHdUVqCzuhBj7PaQaPw/HmHK9N7TG1+aqd7mhUJ0FIfIyd
7+k0G/lLR2Oar3Ve8MqAr5SlPxXHscscyS9sg2uMNDIdhqcWVQAB9ivQb3j4nH9N
g0MPopO/yHOB3sCEYQG0CDiAG8zu6BJzcAZ4JvAjoz7T9deU2yPYGlyCckUTc70o
wXrJRt/XoLrBNJkjV8bYSqOUGdAoLOMeTYKf6KrWoHoOip2WZ/bVgznjrtntSx1X
68SonsdsbKR6e6LQT41mZlOaiXZ8jVQnui5l/LGCB87NdEAV9rj978LSRrVIsk9g
7aMiTKgVG0c/65paJ130ma9Z9iFy8xBv65RRKLAVGI8T8Regn7nSSUoUqImM2Rm4
BoRfgTClp22HmKv9NWenwiGFNc5F83uRSJgLbGsnZCuXYkZ4X/z9jZSbN88hLL6g
jj9VCfcG8H+q7s5Bjro/GBxHsb9A+/SlGB5+dOmEn4ZSYQDnob2AUbIxMAiTzO7N
k3elpwfCjMVeDwmT7DCoigafpOdn7HEnLJHGjIwNrnIz+MsnZbogdpqw69NZZEPc
JVGvtq52nf7u1XD2tcyCWB9rp8toMfCx/G++HHEx8YWJ/3z71/1+38909yFzQOSF
GuCAc9ui0oz/TtVA/hpf0DHYI5kELBj3kqvoXP3UB1yFHCRduPuBuQYT5ZCGv3+p
WGD0i6zIK09cD0msmOpi6NZ5eBDdhflV7C5wFKNF7RzoNtxhJHQZdKnzjYetSAn3
UlgF+q+xwyIB8z2872hmu7PR5drwwFPUzXfbzOr0eRv+vBP8Ceydq4df0qE45/HF
LKsDis0MFNwQJHlRjqzPEa7uPyVsCxGRaQD54rZG+uIYMMrquVlX0mJiMRHbuby4
Ss/ZId+ssZcmeKFGRxE94+EVdqlni6d9qLnjBExFj0IQ/OWpFxbTjkkpqnpKiOtq
0cDsPFsFAZ10WB6UxVh1U/NwJkW3kqpzbQUmhU7z9brWXfmjqy2zINnFb0gyFS6B
CeJVxnCJIf6uaYOtqOeo/MCak7/NmW9MXEb7YMp57+YD1qOJgdE9lGhcVheCJdjQ
H94wi4k3hdV15JkqnYNZReWEM15d1AFDlMSZQDkCiFx7ekyXeCp2bS5jgWJM2skm
pUoTso7ftny3laLjDsSO21hsqRz7XbJ35qi4d6/zlRyflApn3/O2aguEVU/maDoO
2dd9CHejOprtazByb5Iis0DVIHibnTsjMqGtdzcjer8qDybP4exB1h9WcvRzMCje
htRkS7J7ZaI4f/RlaZhS8jXdVPMKSt3j+RPdEZCJoov4g0F+xBFFqs3NRf9OiAn7
64jdejVI0jx1PmG5pisDIuOE1iO/a8Nx//dThnkC13W4DIjeNhwuqPbVtkYlA0f8
DLD6GyXfDSh7Cg+cEwkzQJS6AGi9aHQgi65NXa4QxJGYUV7WnKq+nVGdftJtRy/6
CcXt48ePujX04Xcx1m/OOsM/W9nRBKAk2D1gUhpkJhxQQZDsb+4FHRvKKMC6ZjTT
CfWQxTf+YxCt6Ub0P44tjuwctnBc2aeD7e1sdNQvtAo8b5pg8//3uamDeReo+AJ/
YdPKBFToknTBfz8C8vRDXhf/O1IFAUey0SA4Q0SVnM+jgBKu8X/JETw5bodZ1oBe
GBSAul4jPDMCL8LYu++1G27wIG0Hsj3ekgybmz7lAumgaXBB2niN8mEYg7XlsXvl
EaGOm9PeBODCB34xbNY3TFKVkQtCHPryYY/LyY/VN4p7aZjMMILySqz5Z0Ragt8J
6hhDvtomvArGuc3X4gVQdxtSNTi1EJu92W5XEuR0C5ZNcUIdpzwO6Ser2bbQzQ3k
8rUT94tvxC/Bxvd8YkeRBQbB74gMj2MCWY/RXZ7IhHpYzaYHI7PaDh/t3rbheUPt
z5m68GMcbxiiDqrDbWJU7RQSRmlwyI5r/UfBCevdaSGriMJgF5tk6ZzIPr4TUmLl
s8RJ1XPGJfT2m7npWQKymvnNOTEeeTF5tfhyJX5ji3rB6DZiKFSOJQhha7FDsUeB
VbVeHrzT9eEJTTzzzYEcZ5hFOy+wiU+aF64Mc19vtYd+lWXjDHLlce/d7tyDOvpU
9YE7ZQp6mDS5SOWGhReB7kaxNQFqNV+3P2yJqjSSONVCLANp/t46yMzPbmpaEdet
Y9MRUYbWSLnneGFOVrLfWjhBR79orDiCjHsdn74J3kfi7SrotXLT1T4Tcxl8wneU
7/dmtM+tEWxwud+ffp7TIJYQ+a/WFJC++R1/328yM5TXsJW9+n1z0AqIenWDEkKz
Ws51hEWY9y+9loh9N7+dNWFuZV39fvwO3hxgN83dLoG750SVU2z9cRCBVKY38z9T
7PfFeRxXS7434KkksomIemstEuo7tf8btOHx52tTJvXj82BWwjxaBstoLq8pMph6
kgzSsIb6asc9dATD+iy4Ii5qQerdJsmqUSjvPoWPkqZr5JCrP30EKN7ehgM1tEw3
gWRswWk2M8ndqWEx74h8ClFgJIIHk2b7PMuttti+6oUPSdlXWMl/kfRVNw3v1fqC
vpYf/Xd+FZV+xbPofqKIPWjeloy3s7Uvvy+wmQhFaxXTKqKxGMHsft0E30BrhhcH
kruVbM0ho3QaRK0yiMwDKo2neRRZp057jNLOsmj6GRJqIycGrt9mEBmcXrVYNB2y
0J1pfXAmYJwISzlcG3H64jCr9+lSDVN6tOKY4zYhobKpUKbJhGSy7pWgEZgwF83t
ccr+BfMIOA5KotAe3xmttuZT/nq3XcaHHEoZHmr4NMWCF9rRPa6INN78BrahuTWZ
ge0WjafI/CHlC3fb3N3Ee6iZzaJ5KIwq2vwOQpd4h2UiHcjnXa4c/Gh2zl3gDV3N
nLIlFKqLMu5wKUuvdX86nEDTtQQnp+z7XBEaUmfMwuW4Gj6zynDA8OKQHsCewrDU
tcJTm5M/Do12btWPZtn+wYg5PHaFrKzSqXPb3bsHhZbHnUduOEVeZR8ot0GZnQD6
G+2WMIpxhEFQX4VBSmnmcHvWIbjNMAjvrnetivxg8s0texG+hrDfJv+/CiYjdANM
6xE/erGzwnEvIzohfmHylE2DBoQ8b6uGQbnR3x04G1/4q3Ih3V2Pliq1f+wPm3F5
U/ErUcIXXGE+0c0iOhh1fcqlinAM4GoYby1dN1yceQhEgeLIz5zAdErLLJZaXe2+
iA+PaepVqPM663zPSslDSWvLvlrTi40zA8/wXVK7OwKxMExC08Z/Vxp7BwW07KzG
ONlaNWujqRQfQpBVS1WbyxyJFadMmRh/iBcd+J5WAOFpI505w7AcH5Od3xYolgdQ
oay6lSPlu8RshiknhN81EWM+XyRLu45QYK31IY8W9uQ72yLb4TbUo2aZNPiBUfFX
CDC0cwlhQ+QPm8gVZCAfzQM2ULLi9R1b14Yvp+PUBmQA8tvd+jZI2KYQUOYj7/7l
mKHO7r0uCppVVNKeOQd3joDdVa/Bp9Jv4GD0MiplFWI8uGkAHq2miB7tIPaP1drx
BqJMbvIuYTf+H+LbW/Ocau9DMbnWxCqQwDFqupNOvm+2YP+RPvlhOx6nMBYZqd8s
+c55wiFPUdK4EkphNDr7nFbXyqPAJvWtVSKTBQnu9c0DZHRrmBYq6rlsU8o0PiL5
hgYF/gRZg3qeSQN5q3zHB/F6JsClLaryCwOKV0eo9GYXZvuCJE6a7Tm4e2lmfKlZ
EqYzH74llSIwcWLwU6g9xQ4RJ36xk54reNoXHaH3d7HTtMb19iYlQ69Hd77abPoz
Fs3j+hYxHWCauEYwvlDdEtjnsAYKIt4sowrrjGstGjd6PRGYc6PLjzZjyTUp/l3b
dpyCaWiWAwYuYkBa+pABvYr77/36PVEqGt4jFsvF9XKdY/9Wcb2WIEd6v8NGl1sS
4LFmUqaTQ89yKBc0vN0nWrtXWwuiSXBNs9PHltup6S+VPHkkgmBFGbquOGBtMf3R
tctoWIbGKOsaSNGtpQ//bfukRfbePruMTS1BlVvP04PwV0ahy/4NJkTckZSBtCdT
09DPsOnnGaugBvaYfCIX9e+eYeu3fVNeOLME04RKG/Z9gfAkiqU2T0XUUEMeSMe5
lbfFi5M0l4VKlcuSazEMr3xFSxUH4DzHPq/XTJVhdSbx26ioKIaB6cmzfR6I44e2
Igqc5ZKbOvKesQn7fqdMXEClfAA35IROnKC19fIcyIuSdz7YmB3Pz48vibN+Iw5G
Tlm7TlFp6xh7KACUWAlimjOkrzyKXiFnaP2av265Vpr22Q1WvyqFQYhcj0ysVnaM
WT5Qiviov1iLlxpsvxq+6o7Vf/zhtwEFtYqZoYkFKWYbxzAXu0d1FxehY2MSYpP2
nF8KAInL627zh/4Ky1g4rp8juneoWEWuRwnwJcj+EXAK5gSaeA/GEqvPTwlJ7mIz
sNjC3k+hR/YWQHqhFF/XF6++N9DEwiYwEKfU5Xpq55sHwTsHA1uQI9o1J15PjcLF
ftBvwFmt77vnnRr2P+a2puWRQknBTARUN/SxbWVOpKkVv2or5drqFxWi4DbPTzwK
ZpsO6fJqJzglJ2pRQN79ek4uhJkqx6MAjUFmwOnFSUYjXzI3iyN2zp8nDyGCFuG9
FZWxzvcc2m6HOeA4oWAHemNw6Lw6JPOe0hrGRvaJETcrlAWVHFqTMxtYUMm5ahPJ
PgeC2yBLrOIMAKJ6fMzyKFbG5mdeC5XtViJzEX97ZeHe/yEVtH5tOv7VBl5LEmz6
lUlLW9Xk0Vlk4FJIpz37WvocalPLy52okTyKPeYD9mhOoVtaiLMCT0TIhTMsS62o
twtWcKuE7lKR2HsthOPPeVDlA1pOVIERYB80d/XCsq+x+gJ+XladCdjs3IjtDyXj
VV2i7E3A2K2SGUgBXq9KnVyv85NRjpjoNgtLbLWJq0JU2sZsS3MHIrl13M/0PQvc
oJ3g+fCYU/4/S63SkVpIJBpR1GcNzDiuk6oaEjRAlaznBQX7PSs4AmIXX+TlChLw
G228VFWUJyQ7OfF5r5L49PlRHET76VSOOGupPaOBUp2BKvHVO3Dp+ninD05d8kEb
aKeSY6FIU1a8+D2FUbAvi2Z3d9VzOAtp+Gexm2ZI6bdItUPAsfb1QPu3M4rUhhTc
QLMV5VduEIHVEzZ1ECALP0XjB4NfpU/CYaIphgtlf7Q4yNrQdO6vYCVXVUJWmEAc
htNfRCJk9SWi41P0lQ1tveH9x1N2Oh/yW/wmTZFZhQRfnPka2oOo/gsWueQ/X0lu
160GXX2xhic1cRTB5Ocfj3f2ciZfslvi1ixzT5rxwa2ny0/JUNfRlEAF8+sD9dzP
iRx8wVHIMokToo5K2AiyqV09dTxEyQAd4T+nUFnD4QZPkx/ot1v/5c6OmDJjHhqq
4V7seCberimd5tygOJXh1Ly0EfG55YtMIFv41g4buoygAMxHOainIrBaDyjsiuac
gses1OQYEhH/FJgh1tddH0LJ4akt45/aRt8UDDOGHDeMjmsrNJEdkI1GY5WgO5WE
4IgrI62EDrsHbM4Vzav+myqyCbagx3QMLqbKOqeYI3HR9rn4mgi1TbDdsi0Pmrz/
I3sQpgmJOfI5lOLdkjkueipxH9tvG3nucHbU6V5UwMr+BJ0X2jM5V7MpoifMuBNZ
EKcGUJhVTUDzP3SLe99v/QYYSNkCxuJlpF7yft0t2NX8wez9LCU01zNIGHPhy2cA
R04BoC1973el7OzQ/cPAiR9A+EfaHp971iyXVW/JWoCiHVN6k3IfWjyYgrjDOKkh
NMCjcP6UALPl9Fsc6qrTQm6VDDhXj758ORRyFzZFTdmLdjk0hrRgm3NmK70Hhu8U
+z/imkNAmqhPbMcCNTaEGBUOreqqA3u//IHEIPKgqR4f6tx5iYLZvLQj72wj1rml
NVf41yZ8lOMG3mKIx0+kcaTPFpWlakjKagwHhViifZ2Cr6naUkrT1O6q6i/h9nek
QtelxdIl03DxBH3Kcm/2sLIzsLjz7Ij4AtV5J/Rr7RAeA9eJYSJ2n9jJXaYVR8WI
UmWXI6M7Js4+44w/mEgkZuSgNL/wUszHBObMRsPVJen1IGu3aX42qDsgXOs66Dwa
TFs2AObaMKvd7XAmdVD7quBEWEyCmChB2g6J1cjbYyvkT6YO4S2vizNZ5N6cpi4+
c9RquF+BROYMK+1Drln78D72pt6b4DlPJljGH/F/8tm++d+EgWiJ0GyEnXA5oWkw
lRzfopcGC4LO/fICuXCX4wyfVrrRB7gBoJqIKNJfn8RK1jaQzx3i0pgHN4qWNkuj
olOluN+1UI9/ko0try6hv6bp9Yp2KXprXgyZVGUI5ADosVmFTEfUtK4qUFwB9QTF
F2lFr4lTznkqX3NRHszl8awpmCn5yMcovIgdbnwxfE5I0Y5E/8o4Cd8IHntno0hF
DbfGOmrOc8SwQJ19T4MNQY8Dm5EwsmfsKMlOLuAOgfOC7YXWKZvVGDL/UMcpuFKB
juFWjJypnMDKFmcnzhG/OTUakkWZm+AxaDsZMuhM52jzMFydtUr66FKObjsGJJ/3
IRml9VoFa25yvgDij909rQ19+FDS1/Uk1jqpU54CTQfnpZ1z+ifxUQ2Q2DUVkX7N
42HjVkZ3BmZob7Wu3kh72lNaMpYSJelmyhSGWycu0XhS1DkfGCtXCGX8NfG7Zp6k
VjParB16g8pdvZ3DA12XGwCHBzLwh+s/1DTK1NMIDjZ0eNt6kd3rVjfh/vkMR0U/
eQt6rYoDY7YFXjlPdgLXvf59iTiVe5yo4gdcFr9bcCGNPo8lHKqo5pDBbhd21R3O
X3M29RgbVdhEqykPIModTkgH9g2sqj6omf9GCMxZ9up/V7cbzQuzIWDxOjPqxTLD
21cCAvzojWKadT1K3/WTt38RZnqYKagWVenoDpPOgKFHnlAYdcTBLw4MAzC8eSYg
eeK/DR5SzF7Ju2tgiDF1XEd9JP3JiyPfqbkx0sloBQWh8TLHkq5smoB0453JEMRT
HEW4RntcibwnoOaA22zjrjVn2oEG6I/SboUTvzd5h1BZFRKR8TQ+GngqDn/L60Ob
g1KgYvDjbCamJrscSuP+hXoUeXzkAKh1xRSB4rWxUmrHEhGl8Imd3ELSmbbsYLJy
qKIm8jQh/oRyo2FNbmFhaOanBRBWZewe4k4FQwOLwaL4bUrlofHrPOMrdPPj6Hrf
wrrm2Ym+/z/ygcfv23iAwzcIvAkbzER/Zfq9pRMgzaFmcWncAVu9GH8JGs460PtD
D/mVsImv9c7AHPXxWhtIw8kdhB+W8X7zgdNREAcgziHyfmTwU4zaZtIIUCQGIXQk
UyHvJJEi/urVbB6bEJ6j+s98Fij/sIQCsFjklLuXU4L43ac3NE9afo7OYKNANhoS
GfuTR6NW9jH39DByGvy8Z2pBuXDCwwpVTn9HrjIz5kl/DDX+EDT0hANdto0q/hTa
z7C1P07bbaO8rRMV+pBI2Mx6M4pUINSsPuTvKbAL5Lv9Z4sMznKnQ4E9tFInZDMb
O2cyKiSEKPFkx679K7f/ZT/R4xyuX4AYWWaiSwZlkymFxssOUPXFGS59ynbIQ02F
bLnedbNytMDJud6I2Ba4CE6fXw+EQErGLICEoX2M6ZNDJoOfYXfOuChKDFVWN854
aT1VZwgYTWc/HSypH01szEoD3D0/RWjuHRVrujP3N4kgAw/Axkp3DAPFGX9VzHj7
WgmuT5bsq0Db6MrBeAWxNSHBhH7Re0NHjjDKX/0SXiDY+hhIQzsRxyMJiOKeDY8x
hswoNkuMfZcO6VCwhGRst/VS32R+s7GXubp5Q+Ivo6Pemw3oqVTbGOyiUs24eypJ
F/nke8EKnU3mf2f/MuNvUAIL4w/DZRd9/rynC71qkQ24j2h8RFkfFQkUQMFfwPfK
0iJafpdV/Rss77iO4toRQkjuhyYUiwEwmYAbQOsu7euxVE4Jc4QkfOU8fl91jvSH
yJRQFaSX1ikRv55EgADM2CoPsNdO4Dr9sWQx4P/TFmWGSiCnGiuVVcNzmT4DcoMB
fhSqcMG9VBvcnBntYfJ1MY2N/HpvidE1xCLboOtEicoE6qv0fy+mMWZmMFgSmJrF
Pn4vKzEaiIPEU1+oVs62YGwxfwAw879GTb4m5jrEpdKFyIMZgy+ukGcudxLbOZDo
/nyBU7seYOpOCzKrTCxUpAyJn/wzPvjKMFnN3XWIOtLKuClxx/J9izqvC+mvZAJR
d8wuHnd6OaO1+OdSuLaRlMeAstEGQVuE428AS0PXCYzHnqaJyvZnzftfibfx6Fbm
4kxPgrUPXTXYPTCrhy8q6eGE/ZqncDQPEELPTeP1kFEB7PyQh6GJgLY02PahE7C4
TP2Uiluyj3gYOJhAOmPG2HC2EDdzGOHnki+hMvYQVO4V+WzOBo1pgEmrop5YSM4U
5uznbftD5dIs4IG46SS7iZh1+LkunGBGkzAX5D8qyw/Ft/bMc+1PowYeDKsIhX3H
dTJFY80FfKISGibyojK+nB8wTXhGpPaC4pI00s8TcOcWjNsOFZo6YThJSbL9Y0Pl
RXfwLTKidbflO5C0q7Pwa0NCxnlZI6/U/ljV+WYo3o1xWqGDtvMIiidxYYRPe3mG
5zPb7JYgA5AZgBPA52RElXCjDKk29ZPnJs8MtV5ydP7YXxXn3tQustzTCC3oS9ma
vLfFYp/0Ba94mBLVZWTXBiSpJs6YJpM6dB0mezrpBXqSEmoqe1JSlQ9dFi13P3Ze
vXKipL5/FWB5JvckpUHUg5Xkhd6Vni5jcqVg0buPq2cEXPEweQjLMnhU3tAzyJgJ
H1AxdrhjmBqQchthUSS4/ZsiUduZWIdO9NCZd8duxTW9CiwbsGBHBAG5h9HtdJAA
HJU/CmiTSG3vSK2JnPnTXLLvHgEuteFGlOz/i66K16VYXC3UabW+0X7n4s/5SDX6
qjyO0T7FiCQf96iKJTgHOM3+8fZgQIxD3gc3ziB6HtaEajfUzOtSV/0MtvvzIPxr
mhzgt91JAiDCx0gIPqkmU2RxvL3D/4DxbCRF/GLkq/8kJ/21RHjtwlbR0G1EmuxH
QQcKSNnJTKuB8ATvutVwqjZ9DuGKGUVH0ohq225e75lWjCJEHT9kF++y6ZB31sl3
NQI3KadDJivDyYO2737+RsCT4VzeNuUeilmXG4mxOmB60XEkKFjIL5PNxsA6ZE3f
VhLrpW9IqJl2z9uax7lhk4VckhDeEGboGEP76x2vNA3veZiQfkjxykfp33CCQ0Ji
Mpxf8Lu8rJtmQKHsZJQXC6lmRMBzNlXsSErEIxiCk8n9HnLWMOe0ATH1v050XO8Z
2iXES65J+vyE/uxwHW2YGn2vlHtgD69hmDlc9Ul+BD6NW0ZgkidAn9tgwsp/KtF/
gPXm5u5wOHt0V/xo0bg+hGg7ReSDqUA5z/OHStkS7HXVzJRGo9wdNTyd29weqITp
AYiIEO92cr9tHXtCuONDVC7RyZFCZzPVW3bI4ZqnQCmguitnVj/mKQ5cjjtmIZMU
qdLL/gxJ7N+YzBAMqbBU5RabdY3H2AsozmuOsPu/2jUW7RYd2TqnzVTIkdnrEU8I
OynhFzoMLxEXc5Iufgzlq6P7KRcrh0mStKk0RN8e4CQNArAmWtW+sBNo06rXdCnM
opljYM7n1OeC5jywKlanEP+vZdaO8nLjd/jOqQwVLWH64t8mG/l5xr/Nm9ydQHmY
vukkQwaHemA1VXaXWaicRxHQY/BBvxhR1t6DWOMXaNp0dkqR5f9h4HJ28vasDJ7d
oWo6io/cV2zqVRv9cYzB9VX1EkG0sqsDzpIwvitZDGRvc8nAKvQixNWBoeIrGi2I
L1TVuiaMS8Sdf1JT1o2ZqHKTN69w/mdBZWy95DIsSQSLeWHnvb8tRW1otjFZlV9k
JGooxhlg+n79GtoxbK/qcLNNxfmJCL6rRRLDOZI6k8mt7GiITcnfs4AC37XJdoR0
Eb+Jnmv95SQqzC3PCg8Qim122TwX9RM9ZsJJL7Ul2K7m1T1hSHt4Pr0heuM9CLmW
CxIRv3Cna5RokFoRP1s03pUBqJ4l2U7YVWFuSFi0IxRxaSRZPs8bJmzz0DHesRp0
bgO0l/MaB3e5YiAWA4aFw5Ki9zRAZXGnMVcfuvHSRtQPKvOKd1mv1dA9LFNPn7nI
fmjBHzDDZ6+li4LdFhQfl5c32f/fj+WWftHkh5n2vk/0kGgV4zajuva5vlZxcBmf
lBs+/x/qY+Hz8iRsDvQG7FtFfDbwAfQmpcnI75vVXQUEuQotplXv8I/PxCoiaVsi
0cwCkOCt/yg92dWfwglYRGn3O/fLPxm6PF01RrXGgoSyfKkUWbzBtVEXazlLvdGi
oKwb96/lDc71rv36ErBg3ykb/x8UEWJUWKlroIa+hiQ6NSwK9FFkrGutwd32WyXV
AspZEGtNKza8hYYu/sbslKZt0RPrxgzruFLGib6JajPWLM4AxRjfeIpcDwSZdjOy
CvpBcVfBinVD0C35un3Kmi/Lu2QAL1BPEh7eSaAWgw3D6fL5HdY5dKuE7YE/0GVI
r4iOiuf+tFR0mVsjW/KvvYi3omGEp0drqXJMnGErN5bTjIzGEEYuFJKDkVFXSEiD
DSRhKXcAFdtdXKDm53Nl8+EZJGbtCNRxnBBdqDPV6So1LHqBqb29wt0P2eF4Je0g
JvgfndnR9hIoHInC5qvowZjAbR5K/nx22RM78MuP183+5hn+FnFYd+TdR4IoKRuo
Tn0ExEOCGv9r3jdlaQ/UvgDu7uXxrWzBzpSe4Ne6NPDsqwW+sqcLn42Lw9PGGR8p
2mFkFtfkdwoWZA0A7QgR1g8TOr8jdfyR0POtNjpsQfpeKCL+af/044+7uLgEXhn8
ahHcfIhrK/YecxgYCgyt3+sNxFj30jwsUssO2WACagC5rkfV1Ee7N6ZBBSPYLf4b
s2YtFC350YfvVWhKWQS+kdIXPjrmHvNZlLxQzC5uKwaNkJ5IXmrozX6NE3AGGTQY
DOEGGn7KGeL/UXuKUeZR8RbDDt7ELOwBBzQ0N88tcWOe8qf72carhc72qa7cS7pX
DInZ4obXWtnHrTndx7kgxRU/sILR727v6j2xluZIoLmMa1ApszlFtYMPddhNqIru
+o1xGzvCiN1EVOi2zzlM4JIvG2FY0FqXvK8shwmalLjpcYzHwa8dr6wEX8elRV2J
jSpFjaGSUWKLcc5wWw9+ANt3InujMjlatudqJtqMnuqGwUSWJpSnHkLQGaapb218
h3d2M2cn1iIyetqu3+dSoi6f1mQT4N5d2t9QrqElhY9m8YIkNGGKq4JhC/UVKtHJ
fKQeKYCqRqjQ7wv9G+a+iMGauJOTfILYZb9q33J6s0uPI8LkRDWji1NfPv9kbySv
zHelD/ofLQV8yNgtv2apZ2EUiwjfqxx4UsOBVL0upcs8UFKuqLzyGnEci1HTGOR8
M7lRHFcXUAJKibBqDxiD0xAOQBhhgzU1kGNs0vhnvwWMi85cnKVGpwd3iUHWgYO4
T+3fvZBS6nTttLiHFkJ+iCYKuKoSrXQiq/8W00oLOofCv5uPTwcSusZuc59z9ytd
irvhMHIenHoa55oQC/cz4ctOX5BfoAR0WOq6WDsgI9Z4PKE8q6pN5xJSczlXHaug
UuRc7BYtOKzCt+hAC2x6rab3ZHVipMlKRRwRebGHxW0wLWGALsi6B7KWxrXshJu1
nSeiiQYcoiL8MCKo2q7pE+tem/XxPmm7ojMyLELzHzdF2xyl8RiN2/ShY2RoiGnm
FmhXMQnFSb6eTd4KAuQ5FNKdoTrHvJeXCrBzv9YlMXthYQDHh2ckv2bz61jXqsg7
SAEtNOSquLyxxhZlhWDO6nTzkRFk4dMToTkNfZOjIQduOvyFIypDPOFVBTpZXSfA
IEtdLUFVHsJovlHDPOFAJgiaK7hcmXbc0Gk13fPHyGMUvX7rtTtyimsmVwmhbn/c
9oazgaQHIOHLouerDpE+wUTtGfPP0GiJu7+H51xX23vBn5vr4SSKrg1SRe4bJrMZ
gtEPVAvNM3zIWUOHgjfX6AYjAe/x8MQrHLAU+dBDNFpsJXNs6KLJF/caSXtMrFh1
wNBWr6iZ44zwPYaCqtqnS2/HJMr6R30W6O110D9FUAnPrxLLMlu9jgHzXalWS/tB
6tkxcs3Q5w/lVOyFPwT0Ev/BlRJacBy9sI0WMvMKZ9l+9O67kAhcRtdpIxjKglep
YEAAz6+mmkdhi3fBxsIJrO6F7HpSu+IqleTxPaesQkKuiex2QIYYha6dltRCJ+X/
mfxSqpYgxA75WkV5I/hO5/cHsaPYqSC/GohG3ZfJesdmgMXWBzlCsxai3iSv9R+C
pbjdJQc526k8AwbqfCpkqlTFcXDHeDVmoSn9BkoHJ/ZeXGvKzNgQ7nSNfav+FO/9
3tCp953DbRKvhQ75V5Ci2y795KR38ynSfRgmkd3VLygxKTFzqwNM0sqTzc+AAYsf
/V/Ln7sDLWUyLGznB0wS3M/WYdECfJ1IEk5/LQN+t9iNWLCoqhU1Qdpq5N465RNr
YhcCjJ2Ey7XDlR2l+cTK5PBRfkbkQ0haSKWWLQ4GUkIXoek3arso0AvRDJmTxoke
AJtZ4fcRP6hlL7RApxkYm8DrPxkxzGOAtjS7a7vOteyQF6fngznMQ+4N+ksdk5Uw
FY+VJYuR9ujyC8NpWHWzQrFiqNjFsBEzD//uFr2L9bucRAZ/VHZG/gtMA6va+wPk
w+oblsKhEEsG/7TTwJAUGrzuRS2Ult5gD9VJfFvkvB2s8r+Rt5B1UBRHlrE4PEpo
UbTgRP9eTrdvNnpRXdh+9fQFYoVUY/m8EkIzZGjJlQ4Ej/LCx2P2HnU5K+3l0qJ4
v+snA7UTCuWZkmp2hOHbafZzHIC+PCUtmh2jk+KFKkN0VTtLp2anEUXeuqR1fR7C
uqHav2jFPVtbEZZegUzxdzJ4UU57Y0pe4ufubnZbCtnfVvAz6FrRBbanllc1RoIO
9l3nZGvkJBRfHaS4MGs+5FOsaO9MzWTRlshLcJMgTEE66bmt903YX72h++OGSXAQ
854BOYjH6iBDXTLb1MMC5nLHjHuGjfroY0Zz2rfu5JXaTHCDJItr2VSTUtnfkvcn
V3SZPZum2FcjxVsoz53FKHAl5rV5/1cXwkNGBZRPDpG2cB/NT1N3otA9Ltw0TPXy
FnR9VM0Uxpzkdyedk89XQT20KOocuaczvgIjQ8QzdLvYLVnT6uOeWErp1LJk4Hs2
s2ntj+9QmDtkRaLK3V3ssEU+ZJyzstNvZWlnTvbXIAXBiyAYC3mD6zLJDaVniH5B
IJnShin4d+FSvq4Bo8Ywo3AlLrXrYaIuyUzKdwru/TH/Fvb5OD2Q+3cLGMAWQOTs
5WWKfPCSU2rN2FU8LaD//Fyo+KNz2inmSCsGChNNiV3zq9C7rdZXn81oqzb5s9fn
LGoWkDsynL28HU/ej5xcWKD1zxq5LqtWYQbU1LfuLNureiKVEi/4GM+1ws2YL0VQ
OJ84pLRXn4muSGY1E3bzFeC8V1yzBz2TCsZ3BxN+EmamMNJ4qi1CcenSC0wRYlV3
shXiUHz5aaYBc72C8fRhSKr61lyUZEyAfwM18fViJVE62ameO5tLddQgjpHftOJh
TCeS6lq99il9L8xFODp2PxO2gUGRixHbToIYM71PZ3MpSP9H28ZfDTaghAJoriuL
32xDBysE5FgVEMsBiIUCVvN+Vg5cy8GD21RHaT3I5beoJZqTD+OQ0wpB/M6rYw5i
sODg1IduG9AvPs1PUIXQM4aKSYPfEKL1kwP1i0vgyLKKsLol1elyRHmOTd0uEp5y
Fa+uY+6qaXU4rFW6NlTteZ4lB9jusgl0j8W3/SiwWOs/Z1XXdmK0zFtFZ8boh9T3
1fWI3M9qp3WXFss8afEsHGRx7wiATuY3hSXu3usmv16t4F6N/S/KfuhPDgcC5cZ4
s6gkXrHalXlY6XlGijbXHg3cvs0t9LVBp9ynFmtV+7R/wvPhQJ8Rb22wRvfRpcMp
bGL4CSuzFXzq6YV50LGurd2TNEfYuQI6lc4RVtDxCepmlnz0XH70i572s/c4StB4
PPgBt1nHztzWEDoQRC48E9YIcEfcMRSRKJVIiH6cQjg00baMkfGy38bz+ElDTT9B
TE/y0zrydLT3jsYje2MJnNXKpj8Yd2V+QIXNE5aoR8li4BLvS3CIhIjDSQ3JH4+8
eSvCZFpE1kB3+hYj+FrgCuaStABr1aV7xzUymm/CWukqJDZeVtkLyVR7TTyP07w/
8pcBm7VxenEBjSkD+JZalX34B+VnTn6qIJsudWdDZPtheNQlrbHqZKWhVQ3EH3qs
HO3gjHqv7DbYKpKWULH8IbTcG3tmESfMZ0hUTOCjO9TZklwZ/gW317fpBrCSHC5t
TBjSYZavHc2Xaeue4oIJ4BqpKfNss6UNmR7X8wpq0k33EdZNyj/hiK1IcTV8QUjC
tpuMbDU8gP8k5E7CgQhXJQTAHnT9BEAbaLlMzZtSqqgBBmoTR7C5d8PNR2oHSzDt
5vfS3q/eRRPBcBi3Fq3zV4faap1y+LhJW6OGPobv9RFvRZ+PQ6z7yfsukDkHHeZP
NRmuqxLzIkfH83X7PEep0SSZCoo/eBoR4ZRexEHoHYSvyCtnQlMQxZS5KQZgUt6F
n2QY2iGBCHtozrgqiYwupH9u5th5wCBwxopDYsNUF7FSwoKm3g4SRBzM6azzRE6F
4UFSluCxIl3T7jrJrr7fKNxA/u7FY0SNl2S7h86ncRY6CwkuXDK43q+PIPnftUu3
gtxQGU9VnUnQb1LlZODJg3IGuOuHlX2FsIFZDBWP4C4xWenJ1NwXZBL8Ai7pV1A+
/a6ccwj+RgYwFYRbs5mLJnoq+lfFZErLhJaKnDcgPBLzE89VtvzRy1HcHYQza/bA
sV/h/P71aw6lUAraY6qgGLkpj+V56nSs3QmdhhVGw7HQtZbAQLEKp72vuq+wQ92E
p3Fh4wOja74kJ7HyOTKA5nv5TdKhrWQRrfA9JGdiMorDeH0hH/BBTZi+Z7X7pG9w
fjLFR263F1tb7R93C5AlNW7a4vYsxiHMMDu/da+yEQnMyhEsK6WWOdQnxjbRVux9
82pr9+nTndJtIrn+aUxqZWcMgM2D+yNnAVhh0Qqo5C3UFXSefZze84KfPGeKCfnd
qF9bH7Eioo5ECe8c8CUMac5VRIigaLzmqdWtK+zkmaLDefjIjfQaFeVcfqJWE4Rv
sJOBfTcHTQH6OIL0Fg0AUHOw7GFkoiN8QH05G3tGjjKy3/DAL5k9Ak0mM2GP4N8T
UKLU0XYX8ZBCPwp0py8tK3cAFWDD35mCFP28ZXCS700/AzZJu3iO9GbNvICR4xCp
to0HROJMCfDSSa4Ja8w1hjkIwLOyBqBoHBJ9ak2fRD7UsxH2Y3foM4a+EiEBXjg8
FKHDtxlcD39gAS6XkvyoMi7FMBu2de+/KgwxiA5wVxZ2jveN638ZYl9IwiQVpg3Y
jVLwGfrNUeuc8rp7A9JMm6nymQc/BPFshcMirdjvjxOQU5lIoQCx51QtOqy3gLmi
I8m3eme6gpynewWHdHFLR9gUnP+AioVoObEqPpiq284vFLrel1P5Odlu5bmnYkDM
qXgxXb5PCJM3wOktfRlb0Efbm9+f18Yz9TJQWj0j2eo7wmNiiWuAcPu6rFWv2m0i
0wk7LdsBIXaLV9dizdL4TQqrW839ZpZCcCaO2Yxt6t8SkdLUh2eoX8iQYtDZXPiG
TkspZLt8alpf9C2mtrCUVU8PFJ/ImzBPKm812k6uOgfTKsOCju9YToSF1Ey9S5xN
cejrxOd1BpIu1S5leXwUpTpNTCy9s3LHoR95OuDnShONu8wiL15j/4laJUfgSWn7
Sg6aewIv44fV5J1kMcphGqJ/cVwJsax/M5n7E9y63yYSOC300Fe2y04x/cWHRdKf
va/Q3PQ0gHDRHSAVKPo8bJNhilMm0/QBwFQyiCSQ0OdOmN80fc0+2ao+o75Px5mZ
GQXONiTH3iR78YwEky4yNwH4PkD/CQOeRBp8Dx7tiPUZGXlH11qiCYKh/wpqemiR
hkMnVPijeCd5y8rRo5IXua4G9MsC2bfK32XmPV0UrEtI88ZKmMI6lec3v8IV9Qzb
Y+r7A3g00SZ20pScFphe6C0aBQ8880UZgzEFuYnakZ+75qXg9L8IE4aWNAItLpYN
XFqrVplfCBtifSmc4GnIqm95nOsFbewcaxZMK21bxgVmUVhH31lx5pBZb3rLudOu
9SGDfadQr6fd6b6Nc0BfVJAGoSLJIow9Y4ddD5iWRrlfT6EaGrq8+Cw+A2SHHmS2
iorR6ReThKcHii4k0jtwh7T7JEAUE976IvNo/SP9s6N/22YogcLx+EbfuBRsSqut
dAqcwl7C7Z7PtJPID5pRJi9jGzUH4Skqy5PFomHymtOfd4QctNgFD/aSRtBdO4dh
1WcOvXm2nlSfPt5AmWEaa+8tUUI6bKMhgPENT12N/51FOZAdA1C4NyMdB798ssMi
Ok27ZWuwCHeBFRiDk/TrOQ7xEUJCroKnyCKrvBZ4Q2+wSLvXFhCj8ztCLAhWICVQ
UHhBtHI8FvNocHiYjmJa3sNoQnj/mNQJ9pOgEEHsKJFgKsz129B3D/R62Z3VQy+4
Bdh6XSiJH16eli/NhgNgID6h3cKEVeJbJQcVbGB13lmDTtnK0CTLA5Rp9PH7aAgm
+UcA6WTINtc5B+y8vGoW6mRYc12yjtQTJPuOd0wDev9szZdW6I8MwDIjPNNgxmRD
kbde3Wm2qI/9QANH5KEf0v3axuTJ8b0AHEHoV3ob9+jnOCj0/s2EzixferFwbQ+5
/p0F/xkDU5RbCSVI4VkMM+Q9uD9zinKnz/jEu6MPsjO/qedj3NvnGpSmUggBCdaG
OUiTmAx1kZWrKp0roKRRE3CaeJTfqHu/MDhXhLiB/7ftkvqdo4NBvP/Hb4uT6I71
sKk+hNRNwy57oaA6o3NJqZKGD7gUNGyF+YWIIrCgPMUU7ek59bpwkQ1jZjNI+lCN
YV75/Dq5wstUZ8ba9eS+R5mOks2sBslyIqA/G6GBJhiBdi0URdPgGpzlMfggZVJ9
YhfwtCYvZJnSMRy/eNnVAfKfuGTQU1Q8TZW2Ev6lzMY1AqsFiLQEI/hF71y35VHC
7Ts/HbVY2QdTK8NRJdAX+B8oPXOoGXqA0J8ZyQsWxqrx2d0SaLWuP7Szy7uD1NlC
wrXUqSQECAo4JXE3zjT63qaGIyXaaTT5U7+lZlEPJRj7mdYGbW631Fo1/cvzUlse
N6b64v+cgs/EmuwRieFeEXEus/89QiQemLLKO3lt3tKBzg3EeqwO3Z3hKtGA/gVK
oxgUf165A2kxMflZsbdzN3KdmYnq5/9xQm78ylj2uI/rmvTwy1yn5yheRv5rzwkU
xtCA+GWe27dxTs+BXzaYoOxNuv7emT0a1MmBdavvFUnI7nVcKggVQR7dtMOpR84M
nwJRcrXGR7srx24c7ktNUb+jBcYqwe1EVgtZHXnXS9bdk5358NImTRXJ7bDvK+UJ
YVTQphp8QLNPTCiSMZo26Vlay1Aejk6oncvkIyvk9SkbPH/5ekp23E6wWiQee85a
V7xE5oGoNxfokSIiPatCghM+zI07HGub2fooxHRXc4hOQhQWc62gmhveR09kPrWh
4kqBtHhZKoII9BbKHi7st+c/3efEXEr8hWPwKp+6JojNDPubmtaPwOoIC3KHkxig
PV78p9Zttp0PudADvqbQnV/xQxpSB9gLRYpe8/gwpyHJES+FPT2gZ1dPAyWwtNTe
vfsGtcip5ZF+0BGz8/G9WLlttRwKPsrGrrOWZt0dZsRC1zgeMWR4pX+b5NejYtaD
PavGohwPlUf87HgbyQcmrGmnBhg11eYI5/qertxYOuFPviJ7ZcpPJqdYdWxF1zTn
cvJxnHfXsyLzKwwSNY1tuMFg3SK2E+iIfLrq3QF+8H8aCrGLwBsh1CJCDa6XmQy/
XPibB5o0scVzSEVS87aMUgeqFoQqGKb54t23qnxCulCnsp6V1D8j9myP1qX9lCqu
RaOFgclsDYe70NPTSaRRAz5xg9ZtxqnOFyCWWmfwSiDFkjv6ORcAomJKHEOH8uPY
iU4drCgQ1uWbqMs+mTHwgrCcrx7ejFobai4VYLGDNyvzmIrNBz4uM0sts/t6Cm1y
3DqMhEzRArQFs9gONNL/JIPUP6f9sQ+OlZnaEe3u4wbobXNmb6IhjmYf9jgHCKiE
lO7ql1dGTGSkIiBSVh57tQwoVZBfwwV+5jAiRSUrFMK6HmRr3z5tDZv3gDMnuiU7
itmtXPOTEkYFKKGuP8X/nG3l+MzlhiN6zyDWkKKHKyn3fkyzST6aXAJRaWuZ4/iS
2y2gPAx+AAJvigfzVc/zNwtWsUCIeU+uUb47IbKaJZvWeRCZVHMtSt2fXvhLWS/W
t6XZg0aEHr5UKIfXOe4jl3NP4FFcr8YBQlqovWArKWOcT/M3PmFGBgMBVCrED2Xk
oD4xba/NOIOr1Lc2HIVYI2iTG9QhCBnWG4HCCc6OYvcUPw7MOtySHIypwJ27lCXT
j2bT8ASCegQ2OyaxvoG7KB4Qkz4VfdkNRJreVZqVHP5bHU1kUX2q4DccRomD+G5k
z1RbPeC8K6eElgcq6nVGBO6PvlnSKA1CP+hdELXybXWVQKKjN7s5XleFm2+6vG2x
2VaG7HIl0WnvcsICPHn80daErKsa5qpBU5W4d4yyWRH8KDzpUiKGD7j37F6A9ZHn
fs2z660JjwQOhznfgYbontNWDIrUEvzVwz091mIEJouzozeQiAnxmMPzxEC83frt
bUQchqDBytotG6KOXb2vgGUkMT2PtAjo1SPQmO/M7XO8pTCKQF0Dx4s6/Qnb0UNX
sOfCba9DDIhazCF1wqcLTd0Webcoi9R8SkGTPZ0kUruafbxN6/DpS0HpXkOQjFhP
XdU2/5hMDrZBB+2yM+o0/H0aDwxLItCbOXfRUAX2HiwEu9vJEtlKdQlxA8DZP+cD
mNy0tVVlUg1Y7BvhW2IRuxl/lYKafKPFrQM0x7lk0qEPm/qP6xGVIPiZUHHmwHIk
pV97WfnmHkeaaSEQHEnf1V2xHJmLFHRMJkbXkcy3nQQbq4op95pCMbb9lEje/800
OAQHDzCsmsJs7VbX/lWyYGoZW/HGUIDot4UBo9WN/4iZGep5RdAUoQ0H19GDTWC8
85saOBqWiaR/xC4Mvh4DdBoOQiIMwdtwCTOlSaP6OWsTe4AONzYVZzqg/Pc6gIo6
upSM/tyjEMDmFt2KIkMVhEEvi92XYCFIL42YmeOB1l+tZaHj/5pwwmEC8NuqWFHv
WSrXOGVapBosZEqrnixVq6TsFfTIOogGeUn7i3z1VEmmJVWKEb2s96rkjJGZjQGC
sQ8y6ZLmEsSDW22U77nwuMrH/+l3ebDVYzsNXXDP+grQy7ViCsSQFKisaMYRJjn0
2X6wmBS6Jqd9EmBNKXYTjX7vuw/i3k3pKUv9dQKbckduLTA1NoC/T5USX81tNSqj
WUqsCn8qGGxcx2/tZFA/MMkUO8iUiesvdjmdF9UQPuCLEjK2f2J5Ch0qKwOXAsMJ
c27CvUFuAMSVkemU3W8/QueV1NwxtE4exe0S5YVN4/oq+oGMsDMrcs1DursSMBkM
lCsVjOtXGF5bYTqcNkTcjMh6+2OGpflgZnzwOk/bt9AjjRvyaBVgAVIFsjP+zvcE
p79OOm4MGmpcSXbfrmGveffT/gnPduhJ8e5QpIzLJy5FuiW+zMV9YmmiDEcoZYOG
0HQPku6fmBmEEyRPS2CB1ZkLcRoSV2vSKXU1qTJ9aygJzAKTDxwjkXz5K/qaqLXh
h/kCJOoXuud9hMCBZEd3eGY/xf7MTOoyU0KxHVwilMveYt4XttbHN5YK0VRT23Qh
hYie7hjoUppyOEkspIzsxx0kAfyyO8LGoGDMrGjBJfSngPDoD3UlL3MVlLNkl68p
as9imLG5rMdBTituC8AfP5jstKbZMx/Uib4gdG785rfapct04ZUh8o7xoMDas9mH
vBN5Fpa8BM5d4DtQvxasNsEAFh3HUJ/k6RCmq7/+670uJIH5ZsFL/vRWXt8bntl/
wnO4ZXXDIjYe3q8xtezsrJJkYyc6DpPUKibbEpTtlsiLAig7eJLsvxAiKgdhyFxr
7unmJ2s5CSWCUJspuNRSsJqTws2zh6Gi4YFneT+5NOSJDynxTyWLk3VYP60jhJpW
LfpURT6KgClRA2v6sgu8EFf8/bDtLnyqrKqm/A9phTjiHdqYLlTUQoqk55vuwxzM
Xtg6kEoqnrZWdK0Gd82Zpo1/eP7t9ihL2zuDG8PS0W5J08tZtZl4LOAbsnpXVPzG
0/IQRst+RCG9iGfLtHCA5wk5tiga4wJeXDxgt95e3qhhBRhQjhhboSe6UD9Ailg9
MVH4j3Uuwvl7/HoQfHWp+5E7NT/rAEPe7pC9NE7+ZG77hsbmhyoH2Ijfhv28JwyA
0agMEu6+aJSUX0KNhFJGL3fkZieZCXXQpXgSlqzOkhQDg4yKxHiSUuT+bNqimedQ
hLftWVYIzjXyTric5d6Jt8uu0nst9U8NgsDocy64UU0ZLQUgL0wIBqaLeUxhjTNi
/c3wSImyI4KijUvC5QpI52122CTgJ71rCHntD4VHzsnMA5qIEVsLOxYA/K7Hmqke
eHo1TMcMSnTNXYwztQ09N0itfXgPONQYqC2oEy1vkAS1lAh7GhkvmqCSwTfigAhN
9YhQwrDFwQjadX6nuej8MHyYHVHFguvEidhPj938d4dFTsXg1IA8il1Wx9cE1SLd
o9tOd+xz/XForkSsXiXVzTz7DjTLkbpThg2O7FJ12b6FgUU45reWkyU7S1DU0/pW
is4N7NVb6w+e2mc0wJev2hueKe3aOS70yVUnRa8eCQN0v52WfryLp5cGUqRlwrJt
mRKYp7R9W6ra5EpwfKxtPYtmutasFMqephc7c1dEV50tXA19+8fFLHpngMUNUEB8
TMEr1Gae4Tut3bNCDK3aHsbacGGMmdgWMpuzKjVTyOkEpPsqeY5vS+7vp1hqYvv2
WoLzLgkHJ4Ez1hFbkx9KqxWHKVsWx6sh6k5kFsfS+W8nyDehkfTmWO5NnkwvVWqu
38Lk5z/NpGwiAU6xm+Gh746AM6hawXqlWbTCXzWwrSdMVYZ6fXee4QV51i21OiEj
PN7Ag2wckn1cLGtFA6VFTBl+dNDanzvCeJKSp9SRhX1Rok7e2luI7pCilCbBAPhb
7cYTPHnZ06vOG0m8hR1fwqJPpFKmxO+WSICLRUXCe+jkR2tsYK7aAejUSwb/mxzj
V6dRoSxWxv2ysKUhuKT1hZU5Z5onKmDBDogGEBnzznCAOSYbsB0LFRwWPcSgVH5/
OtIGkwI0E88H0v82RH1vDJGdGMvC4wjCPNcMa6CL+NHyvNvaxyljPWJzIWsDphn/
1MY2tvHs7lztPZFiyoBMAMhpPkJx4BLKp+zRpF4/QTMGtgZkaJojrnVk8G5/xMKB
eRBBuH43P8y7i9iPJOzGcBEgGlDbWI4LS7nWRTMoE+zFGrvDocyVArCds4DACKzE
trbBbwpq2/U1Ohtrm/V7EYedmFReJMBV1DLZZ1IFEP7nlG2sqypDovFBessEMRSL
AReggFYQFeXAFK4fqHobsiJ3H3dD0GsawytCLj9v7XW7/lP4oIMexjGSz6Z/hrOt
avsO5wSxLfmt3oz4qboHBVsgeaRM3XLFy0H93AFuNG501Db5pJgLL+7T5uipIGny
LiBaVq2uoAny0DOwBJIMONXe2aoxcwvmSccxQ6LyY6Xr9unO4LGGqHTlYzz939Ji
wm+kw8weyR5CDMqCWp+v7b+weptdg884XAoXx6VPSd0C0Ld5w6tahSy4pX0/oZhE
0XNrpxu32JKTL7mv7HZii9Yqd99N3n8Opmjv4lYUABUcJ2BW7jqtO0CX2FyerUpx
B518fx9wdgbQvtoYz3yOiwpiyE57Qp10Qj+/FJV4Tm33IJxw4sBhOHGWOOFrejjC
rfhkw+++1Be1L7ctFqvMeb4R9VKFLXrCPzf7g+saj+YYrZm29IxKlfeiKpsnnEED
OZvZAex019ID5UgrVvml/WguZ+R5v4JTRDSS7SuzNk9dZP8sizBYg9kTjjAd3guc
w5UUoCx45tesFQgz3L0h+QNwiH1c2IFaBbcDv5nilpGaaE3ptoqepog/2igtrPiV
2WPlKc1r4sUdcvTkS07otB4o/bqDK1yPHCxHc1mnlHPTK09KdV6TL2thsrHDPstX
nra1SXITFFqdSZJcK590Vg3eoecRH7tuN4dsd5hjNXZTabbEoUMK7ARcoZbAn03d
ifMNKzNqrVwj2JutgYNZk/qJD48WrmYiMjEVh2NrJG4tbr+onJfB96qgFyDXEbCg
xX756P3eg2ynGw9jhw6xDGztiqE4Vx6MaIvWPe51YJ+OWrmNt8mHcVhiMGJI/tve
AkOORnicI9sPypYOLCzM+S3EubEqK0Z6+62s3wfqIxpNhvEnHEHz+blyPKpBpQlc
NGx4MnPjPt+LMxFPkVdh0NFakkJrRZNrfTK7dbud87dG/mXkYESSVG3nB3c9vozH
5zBEYc2d+Hq//fuvLWhD8aVU801KUkWiEmjahLydQpgCaL7l8JrAM5q8CKN4ZXm4
a6MLPIxIz9Co4tF9LcUrz2RhejZw2tdTk+hUUXOZ1/KSfvYV1nRmFjsxX1H7g3Fd
xA2xoXVbhsS+R8QyCkbEdYnW+cZQsD6KBnVe8haJtjVOh72uys0T6WBWnBz4nlrY
IYI38XSBq+VFqKWBvSji44326i5Rfzb6vxXpH7+H1wAzggKw3lOaOqJKmgp6ofey
EXQiqcEy420WhKhOMbvNvai7UoXxn5PPM6XNcSX8x/PFxMUiTeB8l3DPhZJ+sMmL
nddHLpDO7SKLJggvxmTZ1Nnldy9isYBAX45qmFQ1vjuj6EM9SW9EdoqLQCp7roGf
CpcTEUlItHK1yxDMq2Nsrmg8WIMQCCKnxTZIVMjj/0C9J06xLP5bvClC4oT1t0I7
9hmgx8YLEWY2e7S9uZkCWamWzonF+uHnxL0YlOCZROanD4elb9N+AWYW+xplSS1R
zlgQd100sLwhc6mtjEFMulHx9NYZcsGNCoQ5cpsDwFXEEQ7DYH9LGfGer14Ag3Lq
OwbbrtJnhZlI+oWrVnNWn2kq+FuHKtumBVqlP51y8uXzl/xUAho2cX+Gx2x0WXSL
S9Yza/m3ed4c+8igSMH12fVg0RwXWyTsjd4QKqBsxQqgXVrEHbHe/E5iDoNs+Nvu
VF3u6KPSdLqCX7BtuJOH9p1FmD4nU7vGFYaVriRic6uNJJEl9xuyz/b8/C8VydQ1
LPGMWDEaeJFTdT0YvnOnide4Mv/GivINTpWewErDGy5HPfITJrwJBoYCcGm8rB7S
BUJbmsggthkM3ZZl4+msqcjhTjS9LxhGoUAt28Npocr72J485cDLDLRidshtnBbz
qVB64s2aWkL1i4nObgQnGDvIXO+becyBfvAG6WGuuqb7W4aWkyvoaqeXmGfbx5AK
2jnpuxAwZfuwGBYCAhOpHqmAofYyyvsE55QUC/7gGQrZN3+lZCV6BX8YYeh+/PyP
uBTN7gOoFKRhd3vJfTLO8tIDUm6a3d7A5eYsvjoFIhy6lE/hPxyBodrNzgJ8xlH+
vgpETU7siGs6rBoFL8okL1kHS0YT813IexDpUpLYiSdd7USWe/4OjbaeaFZjcxEQ
pjrWTwtNPHJdf7O2lO4x+U+kQv7naxeMFjGuNwdIKBWY9dw4uCSnZHgEzrhB7qHC
sDmEiPgA+REA9FqlLTKNShvFaAy7Yu2/l0Uj4OIHRJT1NQbJwNXHqdZIyASoci34
rEKYvpE8EUjZQV0dkarpl5mPwR77fuZz2EGvxieFHvKxzEuwKLBQ3P4YyDyRRWQP
/tB2pALqoaQuxJH/FR1le5u9XRKMvGMmnifKPc20RPbjzdZJ6/SfDr5/OerdqkFS
/QCylHeLpjKesrwUcLNncm2n/KtDQVyw8zBzvAGTs/K6s3puVVuLRI4ge1ILCuke
zyNktafIast7gYnCALr/BogPV0jcKDsrX9+yq8MAUJbBkPdDDcqz5YMczfgbs9zF
P7y2bWUT/lX7VTa2gRBos4SUaJXnwPdQIMHOQqplpeNS+lfteb/c8Q12Vo4MKs0j
Cb3n16H5MWiSkFCuVgnvEmDTeTJanJj5MA7hMTzT8/J9OYIIpUgo8l3BirgZistu
QCH3C/MJHuGl4k9SxMWlf1ab7B2/zo3dFvKkFggLEDMrgar1lS/JavB1oIqblQYX
5H4z8S5z0vIhPTtaxD/K8Bpjlp8pSoo8C5MEGi67USos+P4E9biSO73cGrrdJRyN
Dc/0KJ6mFpQcH83H3uzOc297Rjp2LsPBoHjJhqMa+2IWjqqaqq7wx/B3seFS28bD
KYDoQr7HTS5bILByBGa8R40yokfWPI5CYGcppstF5Ywb7vwA1RdLwgUBqkIt6eYC
eAgVE5/lA4a8OPfIC4PgPPes9GlTGC6ATBztiH/28Smi0b2GcRRiAFDuu0HVWw92
nt5sDoKC8lJONr9ssiFtQnN0wDX9+dmF2jtOjmJJFJC44b0xNPb4qJCmhwBJkCBd
showTwlHyuonESDxKeqUk5sNf34dKxMcjJaKVwcILRmRtUcqT/fk3CISaon64dCR
R+csXy/YxeWx/gEYLGO8AsP7crfxc9bleNEY4DSyOfQvPssT4Ucf4MT4VOYVxQ76
v3WxC12doSY0WoXGYBN6sLtpjkRw5PJOor4Ri8dhL+D9zDeReXKOiTnTkLeR18PM
VoQWeDd4T9jS/GJe407zdbSyeZUE4GvqVZs1uSMJqxWEox3PzTVluthmMH1BD9uz
pXvhAvaNFg82YTZqR5mp/kgYxetmeZbY1qNWceeHM3lPHAA/MbKhBL+7DERNX4rT
1q2ZihiiiWCq65mGIkeagbEmd4B83BZhl2qr+i+O3vUR6g0jXVujF1NFawSVodds
SUbXfeJouvkkqsrjOr0gH/Joqr/CBsr/H/ekajdISwezZ8UUiwfG1TeWjTi7kkLG
AzT1sUDTaZGUvC94NNAOO0rDsW8LVF33XTSP+cCUYvW9k4IKBNGUvrC+WgFe/rm1
2C5N6Jd8mpVhzFVrRaaLZOhljkphVGp5sKOmSWY43KYWfltwdykEwdIkuL7tCAIN
iLiuOZNVIDy6vQPCQhVPeJkN3potih1ZupuqVH3+U72Tww7pIw+gxWaFjXBwBLls
o6q9BVG4mCkmXqlApsmHN4kT71CDAUUaXdlqw3NHUJgHZQZ6IfHXGYcUZsvoSnlF
z4P/XZhlI56ythhfYI9XIpMkoQw6rYQZZY4xt6xXxx4rGfskQR8mw2DELAnNHXTJ
5Hra9pyaH/MqR4rWibwbjEhfeD9NYiTNIlUVajBYRmQfQZNEhNPvAKF9tKqntFPD
hfQo4MTU6+5iObao5j1h87IGhjVA4Bz+Q5i+bheaQqhJ1ZxHIGfzJ5Mt92zyTniJ
we2KL+TgDsd34qXlgPD6jlG6AWZBUG/qg/a0DFSy/NEPAQjrLhlPrJV09+rqX+dm
YV8SF+abqInKgmEDVVPrroSMZm6WQ8/YX8A7TtAKvbAA+cOfZh8NF+Ng1VQHmF9g
hX7TAZSCN13pt+/OQgpFiOCR+1cNEmLWRtG8G9hIQ6CLPuQc93nMtOHUEa4+X7HB
BX0eNj4ajaTIRDxuRDXwtMELEjqKdDNZL9wUlttzF4FmO7Uo7XF02OgeqO2pIJ7n
2YiTQW1VXB+9WvHmeOnA1a9ZXQyEKfy+cG4SZoRgSKGW0RMP7KGCRfAhdz1VRZC5
LZX5kSxzrlkDLEmQKIPsD5Nh8w6NFxCD7TjNXJjlZY7Lf36hQn6vAlK8e0qtwsSC
XKg2Fd6D8XTb9wQdNqiGwIhWMiXNfY+PKegz2M2eCYw6c72u6WVm16JovF6xX/Ii
B2iNf9YXSkZOfFggcN0i6zM8Pl3M01T27eh2EUkUzEiPo/ui7IcFXrc4UCKgFQXj
SK3cU6mT4T0+I2JhUhLXfFjaapJepfXaThHFVpXI+sn19ky2zXsQtrVLZceKuOW/
xBQghTjLHtTZdjuwTxuPK/OIH/m0OT2Ps1UWnXBjCEh9iCDzr+qNpZ6gs1q9TTPt
u+MaAG0ffeAk4VBnuh6g6u0/UHsMxsFL7K2EjGhq/3G9lT+Nk6VV5Zyu7Ln8iXji
M1Wp36I3FYoptWhI6/pOH5niBNC0TNd78dxiW4U/oPIEQftaRtuZYn+X97PWqkBp
UxpeoyDlsRWAYI1ZENVNNSvcCfpDH2bUJI2BPq7f9+3Ht9w/II/URXxl2aFkOxb+
BfWXwySXObO5Dbgyrq6AqwlIq0fP7X47M3VVohRzb/nq8JLFNHSSbPzM7iUYhtGR
6r3wiTWJY/dQQEYokY3BC9xEZxXl02UzMJiZKX3VUW2wygK7OEd1PTfAOgA1Pdsd
cwAEEKO6MunumgivhK0HSyJqU3OTS/mcIlg6XDKHdYJaMgi0aRojmjgC2s4XnqFs
wJzF6TKCrvKU++1hoR/Bpbv+BgKcn/e14n3H/x9WeXAX2kW1e9hYoLA840hWBtPV
yRWSwCzmovwTCyUnR7wVDoK2ugvwOs2UXRg9rx2GR3Gg4os/wuWeHKXnYrzA66lB
4b+lqxtb3LHAAd35Wdioi7Rhut0ofKWSJ7F4x5FyfgkPseNruajl5e4IrgjU6o+l
SZWeP157uV2KwVu5VkY+UEwkfSqQ1XrANHEI8XCetlhG5tbj9NWmgnrCcLHWLlCY
LppO1qo7p+07dL04FBGG/O+7mpxvFWoESMJV14LA0ybIGjbi9AtRAkAUtPWFwWR/
TTAl4YJX5AFnq4xix6TYQreMaZM3Eo8uUtcOhZIKBZmB0e4kyLb6nVTVkkEiWUSE
3UZiqLa731vl8k727IYXgHxR84ptZlXfSs7rlZLCKSFTApM8JwZVcqvthtYa77QV
wapQsNQQ3Do6GgPTMKnnFQrO17Z/nSOZQbrPosGyXfT1BfqLi/TtQ3Cj644p1Nly
fxyQRAPXYxd1/hP9uU0xOY711iwjEqprRKoeWvfnlks9pibyqzDUcU+ETEJCWKLO
6LP9yBsaerREVMwua+Uf26jS9s+VJRCJisx+XiOWBshglr5hXEMahzboZ051Nh4H
bG03bNe0hzImY0odhR3yan52kRGQCNLdtwBhGwxnzRoGtEVJkcYn/+Pl3oPwyK6U
s2NRmESUlfr5QKH089j2ha4TfdSCiTpk/fJopo9S7dqbvbBaVnj84z8mhDDzoJtC
NoRZOK03pLSNTY53hbNpFOg16JlXbZFD/EcavqJlml0iwYX52Yx3Auybg0G2SE7v
jop2FaDqBTb6Apu7R51K9ar6QQ8x6755on9qmAW0rHGYMRtb7Ln8F02iLTQ0Sodg
ndZ5/wmqRHzy8nuzDS8RVlK+Xc4JALxjua6TX3D84WnQAh1k900hkCF6c8J/x9W7
SJ0mZgVpPV40tc1DFgNz6v2n3uXd53zWoAMgEHkkYQ3bBQ8MD9hUh895jOlyDXtt
Z8KxCFGlw5MoH6PTg738onXh1lwc05KWkMq/qnMc1+qGn+++FQDLvv8ARkzArmER
XS5T5+QPcYXHu5rfbWfuho9Oe5jtRrH0xAXdUvoD9W56Qhj28x8vlC+hdfrbDtiG
XBlPTWETLSfewxU7Q2KRkxreOSJGGmPlzb5p3XqRggBFGSLbVWM7Cpc4sr4TImyB
dkstL7XYbSvd4sYred6XV6uZE0UWMIh8Rq2AmtH7dOemsAYZV3y/FyuciGSoJsCA
tgYGSQffz9h9J4rqDn1PmlJrsNvgQxzMuPcf2SiVx5jEFbxmWZlAdwHDIrb1nkAA
mBpxF11P7V32qqtZriKCmFE4EJ2m0h/b3Qatqw0IUqGSs14HPqAn/kI7Jl08nqLu
x8e8En0Wq8XW6w3nsXEg8hf2Y2NkPsvB7qsUFCwNnvY4oAtJppuPdLkAmUhtLhWN
/MPyUxyRognxrrRn9095lxP08Q5KjhZQSjWQppdKivFXf7lfzvgq+vDb1ofkh4KV
p0VSVB7lyVfMC1wLzz8/+ElgkqOw/peL6Xz31mG8e/rW2ysxuLsdbZK15i9NcG/y
FoC1534rARGNJM6bB4MptnW22pwq1SFQiAY/8mx+wz/TaeiaxLPPplTLyfxXix0Z
SmtgKl9/4BnO5fOviq1gsJTjqK5WoUcy0JXQIEM2xs4rYS0gP92+KhNd0VXATCa9
SR9KP1ITJ/zlqvJ1YbJbrN2yy/9Af5HzmsuawKGpnYeVRckHw72mmrS6JULmhKZX
V9SFbl+bH+Ftnc2g1QdkZ0O1YOz2hthmX6Dww6k2SHRsu9G4oUpPezPxrFxy5WjZ
p13hioAmvGx9KXrLAI+/ErDZ//JJmI0AMGR0u9BSSLsLQQZ6mVi4h7kkNxvkeHw2
XnAMbQYYYqsNHoY2fxfTcFgkJVkAWEbPDpH/7AAi9MFrswm8WRzFGGdKkRNecLgA
wkX6QIoZRHCCDDyR0QMXzpGY+aJ9bRqqMtlRIfYFbWzVOnacWyd2OS4D5pWUopwT
S5SZ88HiwtVOBKWOsVkxdxTHlVG7+GQECpsg/JL6TQcr5TYKiwPfgOLsLPcZd+3u
QxkLSmViDLpk3xmI6xV6Kha3kXAkr6eFGgYM9Cv0olTz6d2QmeSItFRFKRUgKfEZ
Ws23EDaIvd2YDq5dr7EiiJG6OiB08AuV84Z3RT05dQY3YT+lFQeabtH4nNm2vAKT
IapCU9Vhe5m0146IaJklZKN3AL/kt8eXynTYiIlBVC1CknjLT6OR7NdsUTVwrY5h
s01Gsyx3yoHwzOT6Umk7t2BY5EeNPpiiyHJRX4TiL4Nug2Lr/fcWL8WAtm+aTfPB
/m+wo41ZZR5djNCgx6dW0bAqxWSLoVS5sTTUWXgxR1iqjqnVzRppnifcM9s4BmNd
I08IktB53CeOYuxe/dfq9jdzlprw74BlZlogTQKnSRW6pb0cwr+32TZm53VCq0Da
XQDnRqFDkAFu+quE75pCOwhlAcTjVlhS0vNE/k8E0SrPNKnyX3nSc1QK+nfHyQLP
3P5LrxDHxxTV79LKHswUHGqUPya+j7vqOnKbqNghu158+ks7Z1UE/I6OGwdKs9rw
vnczZiyAGNQIl0L8yVYz4y9lcSdTunOTCiOTawtrkEYi5DsuAww/RZZL/gyrEzmT
UapQ37MiW4Q04RaKAAsxn88xflY2WJU4pKHiSOGrGLT7Ct9Q7FMeIvX8caFP5hCK
cEBKZFcor3bdGMcvBDLc5sFTnkF+8ep1D2AMn2Z4KCRxa0GkX0s8+dKuKu3IX91N
tYWSwe9ai7iz1PZJX3aE6gb9CIuZ5GeBZ9ZVNw9xcw2v/gebJ/csbCnz3f2IAC7h
XlW1yuYtoaukbYcn7YjwWGkjd/i68y0mY46xffXNEubZil8cAtxlJ2z5pFBHjmf3
6n3hiJIF5UoGwGT5ZrXFKoDvJBwwnsur8ERvvl6S++o2JFZVDL141CIhSC/oPVQ6
gfSkA5kVlHtkQbUCv/K1YeT+t2JYVsjhU1g815xdHi7SkJ4HJjXboMdeZU5IITFh
n/W27tiDZsgqck2kVhZI1lMFmoh7ZYIw41OftUje1xllY7b83gNOD6i2a33P7pjP
trm8LrWJgmv1iJy59XD+aZiJdYZSY0gWt6DzWFkg2Wl47J7L+K2NLIEIgd2pZk3A
NBXe0LXu78V7sR6XLVLn2Mq4TWAkL3dwhGR9Dw87yUtKm3tjhls1JRHVJLw+ire0
oGX/k6iw+C3r9UoN8QM5f0YKTuLRsRjfZqn4Iu8xqTSwyv9ehokd857kqV1GSfBC
bJSV7zhfsdB6cDkafAvqkKZ5bjM0nHblkfRB/2Qv85Byz0yLnagonbbqQlc+nY2I
myxIA/mz3Iawgfjwnbp1UE0jWBsXYSkUFOHp51KiNklGSw1vO3AGs/P4hwElnciI
j5qrXfXLQk49RqdUlqw0L2xNKz4/DmM99wJ+9cmsUfHelhkrop8TbEVLGmJUD9XY
TshWzvbzxP0C5EvYtbMVlODML/XKfh5yxkgD4HWGUM6KkrZjlY6yDZ+uLwKafvHd
YIMyx8Jk5ROl+CWB6VS2+9HPueQ/DJxYuNUk8l1Kvg0y/2l7BOeTpjw9ULotEylo
BQmmgo3sI2dqaTJIthqS4z3owYPXG3VmhH4H/cagJxAFyxis39UnJGIA567t6Z+B
0N1eYqVKb7eu+zIYtAllU6rx4ui7FgLGlm3JvHa7N8mE6uPEu1m8ZfqKW1dwnSip
HB+HZvlZ4wQ1K41l8riglWUBWmjYzWqNfjYBu75xQd9QN0n1lcvdCC/OOLtA8VtY
v6MLxOUnqAM71ehYVANIVtOXSUGGicdfTyq+VRoEuKXX2mz3aM7/yV3Nt4PoWbi0
SbWYO46/+zujF6ulwM15uGX1Gg8MLpYwms4IvJAvUPC0CS6rDZkk9C8Tvn6KfLJP
BCXuCozDwKUXlwkOEBRWxzRD93ZcTseDr8QwODTpnv6lo91l1zUnLHAtu68e0ydD
C1O0nonFns2F4WkEeZPvBjw2DccXgzyLSV5ThiLGLHxgsu87aCbhWNnQ3t3bUBEo
NCv+l6SUrttQGv93K0je6TLyWztlTikR4jCpRh6mHQZ5uouJd46CVWHnV1xBlj9m
kleeKqgHTTJVWpMZgIk+mW14GnSZb7nlp6Sswk5+XvQCS2e5y9NRcONYoL/9ywEN
f7MqwW6CMpnwun7uHIN5MbIWVKDx7KOqzffxaDXRB+fapLYrznfI9aSr4OpOgN6i
wvd0pSQl7MVdYPQmC1HPWv4u6fWqNxS93ORJXNL3zk2WTk2TLwIvUzTBnOOcdhy6
mnMiKW5yG+RnAYjPQa0SDcESi0+hfifr5ujgzL7m7MJanIGlVplNyU9+yJS1FJZ5
gLb/Be4gkVHcy1YMP3hQLSFetXf+6WqG5B14bIzQg9ZNY49C4kI56kyGWM828lR/
Az36iqf8sIQgSnEjz58JTgj8SEwHqTfYlhuTRs/VPPadBiY316j4w4KcO5Sg5T/s
DyQJv4dVT3K1292JPBYhTb1G9uC1InFH/hOfxCBaLlzUq4jO+4iEI9sQXT/76zme
Ne6+iIr5bLeT67u49fwefS9ok6qYtDISgYfcFg33YcXM1dSrRHbOA/jo5CsbqY63
L1WHJBRXmPSftl9Gs9s4flYBjJrE+puPv+eBILJY2oklG6vhqWkX8MK2ewk7WcMk
yBT8CMtC7FQWv53Kfqd4705kZz/V6HujuIewapSuwO8Mloz+xXSAtkbbHfrFjK5v
5+OtwO092oYS+QQ7ie0ESdi4S5wACe8VtFuOlm1t3Jgm0oSnKKG6DRuIDFFo8PLu
q2uN6LEJJZrSHBVgpJTAsnoRprIH0AA8haSTsnjaPGz5gU02GsMzGHHwuA/V9Npu
SI7XMK5KiLQ2A2lXbbIsM//ijs7wlA7uiz3Wnw/YTkp/5Kcsgk6pOKOahpbewtyG
EvOWf9yZIms/GxUgyRiSJFupz+DV2N7ZqDZWLFnPS2hTk7xmz6xgnZ+X9ojA016s
vhrxI+tD9hgRpYKNpnM9dnJiDBS8GqaQuiUkwQkSfR5zsOsN02IgRC0SyTCbyKu7
7r8Iy+0YiKQiye9BZw5axO6CAvyuKhsl7JxuIRju8Qdl0c7eFBghGlhuUb/dSK8r
96+PwSxWJWftTK7CR4D2HDLEqjR6yWTWEr0Y8MX96hAuZGpVChyzngW27NLQFzOs
GNgwG59f2EznuJYJoLiJ3wPlPy2K+oMe+7IRPWuT092MYXge1hnTfMZrKVHWriLm
UsLHIzALNlP78kwBZmxikUoU395laZmK/0t+r//w3nUnfEh5C1akcQCbV2Slvtdw
Aez0UQrukPnkKclYbomww41JztBiqUFsJ2euHzbmfLcteetxYkCmbS++d7eUZhft
OI6jXwRckZGlId7a+o7wrsmpBn3wTmVge5BrtUALLrX5+eKh64SrJWm5wlgeExmj
Ah+zIst4kdOgPDa0rcNb6/vwP//+XUcoStylF50bRxXtMKwVXZd/o+hxa1gBwIgg
RreWXUftLOwJmVcSZ2QcBS7nQ6HW2y9ApMQX0S3t1N4cuOv8MpyOm7/LBX9pzZjH
PW29KgVoNd5gdL5HJcXUjrstmOmcfelKxPUBbhCvb/cQY7MT5PlaVHiSZ9kWE/89
IZDHLC8GRdiG2Tx2v7cPCgFARb/HuByVwaFFba+UWYDiMp4FRjsBJY9Sv2JQ6wyc
thQIhM5ydXAEZVMOYjehIyE1iJRqeYGy07RaC3DJOvAZSUSSS/ny3JMwA/HPzX3B
TzOaXYAWNkz6CB5Y4bDU6COc6RAkgg4YrxkIAzWPS7h2JHvNDXHV4hK5w042vTB5
WabzoYTe7GeSdyYJWLlq9G/Q9Gryv9wLvhqL7N9VCEeuAySwwNZ4cYl8ZNMj4niI
qsqx2nqKhkfpAdK3CNwCP945LMUgVWz446Em0fZ1F6z3ta930VQfgVSHrrusxvvM
09ZOjetlwbxMeqXKL1+3znKtGjTL3u78bfu7zZLGfK8Ekjpu7KqJtwD03mpOUov7
VY4aIppZa2ZKq3iBzCCzkavApFUsAcT5/wcdqDGE2Kddomm0ueiKxgglVCgFTcuS
+SIJSMDyAeg4dks91J3IRj8OzFXhvshQVbLRBHXAoKYcEJEFLolvLnnim9891rXb
NMw5cxCITEoEiG/BhN6iEpz0dvZWxME502S4nrvQLVEarDesh9mAuYV4D8FDlcg9
VoQeGead+ld0mAasokQI637V7wIQgNaA2WbBtua7YBbPenrjjIUIPRGS+GR750kQ
Y2W2KNJAeHaLBO6ymRJMT4gf6RN2dkusyQR3uirbd64K/Uf7w0dXavd24azRWU77
DhXmQZEi+VIyYtjjniDpej0Xolb5FKsD3JWwrXGNWvG3g4mG9Owj6sdxBfeicIp5
8OkBJieix9bHAeulzYTnGNTutcxtwnSUaKDz/7JytOSwLkRNqS6ehUco2R5Gjz+H
Xupm7bsKBM2a2URiQgR7SKlFJWO4y80tAWZ5j31cE4ZNB3v7QYxt8TqG2ejqVF/X
Itfsxc6XfN2Qk3bwuPCG2ggpx4FSdLz9iDBR4R73AcqvO0JUMlW6XLiLNak5NEMo
e3Iu9fXFeXCm4RgcCXF0AQbDKlFBiBvJEPepxRGNG+Rk6tO2A2TLGPFU3ym7UCUX
D7O7jP1VpbDaywTQN1Zqt5omm48Sul6gKBv1msyTwcOJrC/aBPsJf0KnUGUw6Z96
FMkvRBlQwZD8z0tC2ZiyzowRdksC5A1B4sc2xOR3V6B/tQ3xqIFhctI8QUM25Euw
C15T2CaXNgl7D8NmperMDlDk+cO8my/N0uzOuXq0DkuyFV0EiuAr18F0eXmTW3h7
9Xl6MRnH5PkPo7K+JyU5WwV8XiTXNHeQWp6V3tDi102wCiPoDWnmanCBpBrkJCRf
sVfrL/585jiBHFsWDejlNpimawbjIR01wCoTjuktTbdKibxXy82YrbeVCo2cg9N9
iNXnERdkzhDshZuCSj3oRlfVXUCPYVMqs571ieyJjJvwKYWrIUjV8Pb0OUpLZ+VM
sXJc/iVc17KM+xfDHGLrQSv8nFjHoKFEPbYR8YygBsnHMHvJ40jCoSuRg6gI7SfE
jEhHvChA7CBbA2LA0vkwXthtwAFgnRvuYxWPzhij7vacsU9OhEG1/3x51XA7+PCI
3R+YA+vif6afIgrcmXy5UC0x9zDWAwNokMeanyH5M79/ABp/62Vdm8t7096p3iGO
7rNCtHYGcCCX51cHfcuNBCCJ5dSkPeYfr/wxftpe73jlJR0s0b63Dg7Zka1nS35n
ujlmFyklsAhePsoNU5IcGuqf6Vy4RA+fzr6cFTqBtDecAt0aJWcHXBglzFdVqxjs
RlvCVzPj9RXsXtMd11IIjl+gOx+khRIW4i9ZBU8AqtuM3PX+yIDDDofmU6GlIWSC
9sAg6YEA4VR5SmbGk+782nSzKN2UPlL58zrOYt95wz3HGYNcGyWVkUmyjdb+UEmH
gGIt0ugp0ClPU5fK/UMS/hNDaCfpdNFcnmNcVLODaYZUjaZNykjBIQ9Kf1wTnIvj
3ObTnIGEQBTNi0zTqu4AH3bSQLx4H4+dIWLi/JOGZ0XKruN05uHLyxdTnMxpdgoE
npEW/T5ba8qYcEqdfsEo1aOwzF8YyX5YrK58SykcW3AoM/KjECbfwfaqFBM2u0ti
dYDnK1ovENjmJnQfvsbcnkr09vCeynXiXZE9BVUxZ5uPMavvuq2q+V/NS+hnC2OS
mN04VM+STlKupf0wUCRRHf/2malsBvr6xYtLxqFY04pV3A14hTmi4YavpXjjJxdH
vSAdZVNypRMpWWcmeL1xw/ibjJYr1Ppnx4NXgqrgEr/MetD0b6Dv57jTL4Wbk+EI
zb5U+5PLyF39VJKRaIQhfS/6LmO90twoopsYfS9MtSUuOHESNXJR4ar2PXBcyvQL
mj0Weo4ZtpbjEtBNu5O57jTO+Hhyp9D1xpHB2dZJJAmM8w9JR//0VaMOXqwXgEOp
VScLDVesaROvgDH5A3JBZuW/wDnfNvFwVOopqV6eSe16tRioLf9wSpzpd+7wUgWW
L1au1i/U/qKS9NOb3n6+vnzEnw5EootSkzpfUl97xgiflpaEzdPalTdcbLFZAqd6
eMqxthPtYsugFIIFBv31UPSCfgXTc+khkD/zlgDeCp9PL9DQ2Z+OoxN7t5YekyNk
T+6BOBGo9LZunc3aQq8Pkk1vXdz4GCSFQIX0vWI5MPvBs2g0lg25t9UprfeaXeGg
X11Ud/Vuxma7Er+e+BZxewF6RKntu/Twkjv1l8PnDAeo6QIpF7vVUuOdwlOimsK8
JS+qt0q5JMGu1Y1sFCqkxDtyYOx+QVw6yioysWZ136DhKguerqEWJ206Sk0dRah9
zox6qFZbeJ1oAujAjslY0pH5etBGnz0XW8j9d4qciOsdZgcNP75QuvzCqqY8FYTB
E2ZKqAdQfsqRhn9qq3HyGg3CfB9MjhjWNjCfrRvXqJGGokQyJt/kmlavU8qqgQpu
6U4L3kPt6BI0TFDEFFQFjwnPJRGsqC5RsReYvJh44T2xH0yOFFmuBQXu1dcDGgRa
xUQhkwlSJnSnTS8TmJ82AcLoM/QXV89IR7DLWaCO9LTdFXy9F3v4b1L4a8DgFYzQ
bnZss7ErTDeuypme2bp4EJXN/oo3IeYmJekT2mPjbScYYA6+2aBKnnIgMuCg/0XT
9yECi2sLHzzpUJSs487XKzffCAemH7cNH25wXgD2yofLiC4iEEJ1ew3FjtVpnRRc
LPXFZuvGVMgilzfKNFxlEUmC8gCj4sH0U5HUD9SmoKZq0hFyY4jwozKy9PGvuRXQ
z38HWse4SvzPFvob3Wv6iq7hTfH1H4aBBtncH9cM/2jXe/3d7JS8/rrwDHxODUdH
rwlS4DloMrA5e2FPPPjlKcKcYYCbhhyiSHjXi3UzBdbQm3iL8M6kE9LaG/IVwfIM
I7SzNgeEgAVdXiEdtNuXJPslD3hVLMu7bzILBt6/ZdTFBQJLVLMzxX5SPgeuhd6u
hOO1rSRNSKES8rl/fuBdcINzgyn0rVL8a3QgfwDsrvwJvLqjX58x8Cvu4U57UJLR
aFLqI3zNZyT91d1YAdkgx4+jiOja1juhhJkUAwN/4/ls09lEANcaGaLtAGk4gTok
oMv8hJ96oXcFGUKxCgtT3lbcwZZFMBKsomCpE5X8w5pvlgLDgONjrd1HPkf6QW4n
LhEiyzXCc4/4P1JZ8rgL6bLn4x8ppobaTMKg5fyOBIX4yzpJEpOLibrmp49kUan5
kvBQEwFZNb72SUUnKFUUttpsCCEyaofEbL6TuAwkYbhBnlGJEpC50JNOqX1T9Ajc
lvEw2rCCO3w49ShyIpuPf2CcjR6jfxIt9nSaXGJkvxOPpt7AxuSf6qglbn2XYLXC
xBX4hepRS79Y2FBucFCVrHga+tpxDL6mc9/oAz0yrdnvCJHZq2aiqpaSdgpEuinY
2h3ylnev0Zl9hp/ybBMMUeDmTHr4GzMhFO6bwGrHjH6g0pymbfm2asDVzTy8kWDy
qcApnjKT9oYJszfJ0Vr8FsMehcEiDlplepZIx4GeNpDNDb9L5DRWkzVUpcSnby+p
8N6ERwbLUsTVDksx7bwp5FmMx1Uum0Xj2M6Va522KTCJcmFOXmwh8X/VxhRYBcUX
6kFh2tvdiyTXe8nWszuGE1uyCbAnSLdQ02U+REjSH/gLBTkTrb0mdLtf8kCUA3VF
WF8LdhNhaD2rEa9syYab8kx+QW58VilwCAiwRF3oAj6gkb/RRmUaJ0EYr899nU0g
JDyJFyi2ZFN9fmTnqUJlS2CGbRdyWrRQhQoH6mzB7fmf7Hb09UdyM7Nq6AiJ10Wu
1QZmzTCPbcrf4GJwsU93O0ivvDApL3ECjfBiElQf3Ttev+ReidAE7L0havyFUToy
hLhucGUZu0lS/pPIsqFizKkZPmX+XCmRG3aO1WqdwNn3woP/YUtI8O1pJtFpONrU
Xw+j+NJ164txxX38fIGxmnJOrEo8mRUBLz1zkBZxjxwfJ0zkVBuxyllpe3Wadxgd
aVdOD1MinADqbIEUmjAA1yVqTobq/C/mfZ4u20YzLuS8Csa38Za0oWbgIQaxF1Bv
lJniMpqFAIQogjDZV5RRJCeJ8kG6PDbs6micrI+dfQ9Slvy/eEazDLJ60pI16fnF
7mwEjTxsrSDKOz3k5YkMgyMopNjmN+6qexJJH1eG55uNSPveT2zQuthAyBkkxuOO
s4jZrFBK16IQggVjGAkN8ya30DbToXLPeMXAf1kZBaaY6yi7PG6t5QL+BElnkNfh
oig2fm1G6msgtUIVOW/GlYbVB4h0Hcfvg6JpxKSwryf2Jnj1PtxH1/uqx4FsEl7V
BCCLgF1s7L4UDLPWFfyagUmoMAbWvp7nAbHmPh4i5BqQoKRAYgjwohkjuJ/oyTqF
F1uV73wHp+0cEiIVtDWFiAiKv8R8YFNBzP4Fk4LafrOCN3BfjPQS5r5v5c9M/sSv
XF76ZioP1BZwoHwrglMQ7MCbP+TzHivjAIDu8zdJ+tOlzmefiTY21loh1Km++KH+
Ykr5m3CB1/oQJWHBuVPUvaYylRXV6+GMJIWcLtzDv/uBvWQbu7istd0gblC/BSZO
V9B0RaVp6mPyx9vdmzUCd1OpVkCjqInudfxvpLOLjMvuLQ/QZR25a4JaMW/pU4Pg
+Frl9kVOMXdom4NFqOZAB+jCW0eWV4zEnaQmB9Bp9acXXf54EJyVa1tOnaHru2AP
dk8x1MyvoDGzMT14OIV5fqBSGpBrGojAsZxhH/2xOR4yQq1bbFnr3eh5Twe3Lhzv
0nvBrDRi8VdO8IaGfPTzW6Biknlz8TM40bmfy/cY84oL0z1zf2QykNZRuE4zOX4S
P6eQCVlsr7uBNrPOyMzzS0pdIm534hznGVqhYkbcmugOt32u5YRGe2QUyw0GQv13
87H0cpII/TjMCx4ln93moDmOe69xaX4VFWzqP6ShxXWcmkiqfqWcQbdpHXnK2mVZ
zdjtUFvMT/TX59IVBNecXqWNF6hJlRvIHW3Gt07ahZIz8uK4IAmQefshaqMHjmIF
1EvJWJWQWGTp6vocmNcTPiKxyjZnp/OvRqR1pVxXQFXQDdEsgRIXzDgi/LJ8uqBC
bRXmNw6UuVVUIYSPDANqCTWupfAuy4mx53pUxYxXDL8UE/LMibKYjFJHZFFbfkCz
5tyRXBzvaDvxKk0hisl1xySGcv/za3mbfwVsPwMeD87Ue8gHGV5WrDiRl+A4v52C
IurvNDwzr5NiKyNlrnoy96qYS8eQYtqTXNpHisOdUyelPbDnQpslwhrKc1ptzuLY
JfPRjEhGRzUS8+2ydhnNVlHJjX/Cm2EsA6EZ3soduaPr7DF+X6iCKyelRI9c1Ft2
/0KtRBX2+uNCeYrdxfa/Gk+FuVc5Len01e4kBIhnWDNQ8Qf+YooGlWw6NDMZwXoG
UMfV0yqNQ7Teeu2WuG2FXSJDih39R3xvg8SY42Ov0VS2uJAnru++CtSuxmUx22cv
ArJ8VRZMpNzCaTwPmsK/txHUcD9of+oKpOyLvHcZMfMz2OE2VFIqAjbpZa8RsLfA
uGHJCkskftZbs6h5/BRKQG7VJXlTEmOjhpmGJcRSyssENESdHJgWdlUOrD3+tzQ7
OM2t3s7V6JO1LVnepLziHQaoNeExomdGvQvdRvAtW7VaNGxzo8qI6fQ7LCfX/OEZ
lTrWHYby4tHbM6/vLvRJbZM6zKImv7oR7ihzteqHAfaj1hvDKO6NLu7rGZ8blK1w
ooYZDOsWXIyVl/SAIG0lJzVxoatdkA47ijhXun001EEIRMhGoU+Zonv9dyU1bxgu
494cGkarBLGiLB+Hk5hRpnjucfpQ8wsYkJQNkYPQilrrP2uBTLjDBgUvcGbcm0TN
D1G5YFpLO9l+zUSGej2mvxzgRtzJz1tB0hBU44wKa+jPJUy5pDyCbJFhL2a5CwHy
hpiKpkAX4UdNVzZQGgsNM1L2/iGwHluLpMEgWCa2kPjFhCF5w/fONQcjtgYRiUmz
GjBpzb2Fp+NP8F6IqE5QorO0wGf5R9Y1IMcLNDgtBkHvqDK7/0EIuZuPpAiMiPLk
whSRoIajLoX1sWkC36Vvd10naELv5VFXNjXD3Wliw0qJUcUoyxxmCYcZ+WVeImvj
70mO8L5gO5W0faZn4XMXBLx5AajHycQy+OEBD32YA+lu+V+uD52rlqzK87UimhuD
yT+UjdIoM5wC+qlwZfzzS9OjqCv0v2R9KNNjg85VYGepY4dGVK3zFdYrE3/AkhNh
QlL76inECVV0x3b3aOLvyLYx0HJDv6LOXGMTwiPwmbI62ZHX5g/jF2yZNukAHk33
i3go1FodXPtkCjpOIekjkT0Uyol422tCeOnp+gDU33++WH+0AdD2GAxaOyG/jZpf
5xtptT+xDQGU07iVJwRe0VRjf0a29nQl08qx++mylG+Xhlv+iXBWV1fNSe/GWRMK
x0C3sKCidAx8/4gC+6gRkQUq/MxvrHndKrXatuO/bSLAFdWc/OgJ3QvNjYiq8pYG
HrydgY37+XZKdof+EhGcowoZ3BYYVMDXVoFDRuanKy/ihSZa+u1q7ZNykuRaH3XX
RFPFC4nNJTS6DwvbM0hviYFFZWlnlF5MbBGYpOvi3k9xwcQOdMll8gxitRnokePW
j8uaLI9g3YvXPFq4x3zTqf15JbT8TsTYbWpC8KEaKTBvOI39/euHEC/lvyJjheZv
nWKu55gaetcX1Y8sr7iAdqPPqQTjYaECGJIw9a/TqLjxGa3mkqQuI7ghPiFlrYsF
f/FUHfklYbLqkHqNv1YGZU5kX9fJFYW3C5RCetU2ygmcaTmqGGIE/MRQ+Wixqnv/
/nP1W0mm4CUonD/kuLCq2IZabaIChG3J6EMokWojLYtD2u0RzRE/giVYzJcL/i9y
XSNQA+NSVloas0Wy6gbKhzz7cAKMMbhbaW0LuPOVYOx4XN+empYw2FQdU/QDjJNC
8C4X4/p2lM7jtDzWOwA5MkVEy4ha8TwEmLtncn1qKtFnCcGZuZI/bXy8cMa8HOOV
2yhQn6Gm/VrcCbnqQaWEOvw/k6e7WytDfqN3B/0ltVnohcNoLwAwcJM/JDscUTGA
ADiSz3IFARfkzC4B0qOLqLl3fq1quTPzSfg+RH/mJ23yZg4a2d0a1avaJZNY6TaE
pwcBKNQq3NZr1OuW/uNSrLA3ULEFemeIOtmh1LwctNk9f5TI4w+UMeywcb042yBQ
MagKQWDnkJ374jInUln2KhGY4eGmlphYiKPgNjiYrFkjh+SDaOKn/fs9zxcmUmtX
RxFOMnCxM6rmN3V51U+Tte28xzVgQtVDN5ArM5p9AfEgx+QMX3F84XonMXE5/2nM
CmD9vd5jl4qRxYMH0EuxfBsYPxkGvkXWIj8mjg0oq9ph+S844uk8PncLlLE71aP4
Mv5O/sZ0pgO0aRCGRV/RzeGe+Lmr5YC04ACaPDm9Z5OUjhf1AyAsP75Z3vcUHOqG
3FsoJVrnxqKcZUMvivqQtbwYaYkiovlb3ttyY8tPGe6BZErzDO45dg68dOWOzMls
QojPvL8S9tyXfInxOtztQ2d34y1KE9GYVz0zERMnJgBfxJ3hnHSt6IizuP7SjJhz
P02ZFhQs1kBRqBoO7u4+uPld1TMj3O8/sWdRic/k8zRjjywPcn5Xd62Rq4diXOq+
98T3wJcupHxr854gki54wmXdepJOgd+ycC4ZRhJRbWrPVNfl6enyI6Pm/wXzmdsI
NVPDHuzGOGFcrYPkcc1kszi2ZcuKbSCqYbvtRJiNKeHXSx2VUgaAd2bx8qtkUeb0
+fwdi14nvUERDB5qOnT8mvulmklGYOEAVSl7BUB5s1Ob+IXcYNfiTLwslxBtMiH3
5n2cEpz7NAWlBH1lrb3RmQYqjOFm0PLSQf5raw7BI9qDzujF4INvFVWwPQ4OVkHB
rRfMv1oKDsXv+U/E4Idzh1HaczgVVxbXqiljiLbNR3RO8tdkddm4GyoAd/i0/ia9
JSKBnmiHvYR48rmb68RYLIERTBrJA+ICbuIgZmkf+xZAXJLmW0ZoBj7A4lYgwwUl
o0VvvfqFFM2IGMq0KiW4pxK1AkuuJt0vmvI3LEPfpzXwfjHx+pn83+KxsoBVzY/3
WDepAH70U++tkjHyNZlq2zwtwvbuwV1KUVkgAWf8RDNMSvh/9vPum2oo/jeLjWql
jpv67PW/C5X1VhGpkdD58bfQxyNyaP5pPodyolJ1ziBciHG6LXpFcfssNKCLQHww
Tv3Cjbm9Nm0utdYULomTbDW+enE3S1KdKjk3wM9Dvs7QufD3jN/HlpEDDnex0BeW
phfK5q6dXteFoUhooN8rQ1JKgmir4zsOCwkt1101JavdtenDpxddqOMQV3bQg/kc
Q+K0h7LFvwI2agWHisF7e7aMVEsgiSwAnQtsgc8RI7EHPq05AkPsOy8sP3JYwL4m
mo1Uxvc75Chcb47VX2gNR9ZXYGqSz1vgX0yiJtwXkL5TwQI+DbKwbEKmZ5+wEbC9
O0gE9hiIYGwdalvL9JtSC6vLgg3FW5d7rGyIT23sSsja3R5wwatgzrPXg0AtUkFs
VmHpwhCDwQXNG7vLL0izfYZATk4bolXFkIT2Ub9m/DhyfgL5aSUBo5YvZAV6VkBD
PzK0aK0iYD/5oI4lIWsVAQE6wwXMvourLAnbfZL5JyPtAvYaJwmNY7Rw79NiK36H
6tCt3oFeltM9cUcVOoC37paU1qreo+C7K0am/XQBIBrqiddU4F20KYve/MplyBgr
37X2j8iC3R+y5KcuAcfvnFvYGCsiEUAbVkSBOoYqsa/j4RvU4tdASARmA0q1Ijyh
F4B9ZjRjh/rqnq0swNm0sPYDpHJ5jSuUFy8VV34jepK9lJ/Hxggv7Wra4LllDfVk
ZP1o4gvxDHNbLzUCjVSpq/BtW5pP3HWo9/RMd5pH0p83oRZwAu9y4cZZURqwANZF
4SjrEt0H2rjRza/tgt+j/mmJ42VwY9hiFfjG9YTS8uz/RtmY80OAJbMCbJbKfzWs
UZvNcxGxj8a1PFy/M8I9sluCdFCPcZc1uIGOuEReEfiZwU3t0DjBkNaBHNMQBkE9
oNZbAmbk7N8ZzPvOeBqkVRI1lQIjqe3NlB9hyT5julNRI1aP2CY5QY6+gJ4sl1on
ZnGHckXlPUGQipZA6KSolGSeBMQer4kz2VCDrO1zdhDiG5LEiD5Rip+vtz20wZds
Z2mkSNbJk9GbMgy08VrzTsCrz6xqF48Ve62Tvx/LxXwWsutZhi4h0uqWAbzZBsfK
GHJUNKKVwyAQoyY8SXnTOsVwM+wjlorV++Xpll+g/kqlFVIgnOhGO3I45NJMP3a3
80FaH5Wzo56DFkP2DMFHok+GfykPR4oV5apSLpbqSI7w89kY+A71ESY+7gpjy9iY
ivn88y0AvSiedR1/1IV39CpmCqsK24mNm/KsLiTiJ1oL9bLEvYXLR/uhmnpxom3X
oZj0lxVzvpMvGvICP0WnHh7qMI3db7Bawi87KD568VYD8kGLGlNcsBoab+vbG64m
pt+6w9FR9wpF4O94/zyjrH4ixH5AOJGIIfqL6AYHuS8QwvXf21DthL2rhcl5te80
uyz8n40C0HalCOkUAamBlWfRLKUaEXUvmSjEeNp0IpJaxcTRDThG/MLB227DBEc+
Bxn5o4NZ6FNy53Yqsu52RYWeloBhldmXC7hOWgSSnQ9DWff+73Oxqj+zK/wJRjHg
35uPEc0zxTru/uWYcnhYI9Vh6YBGPQHmHqR19SbSzJKzCYhgAq0Wrt5CDuvL8DqH
3TWgxRJ04WllOP4FnuiDqxnvNhhT2QIeF0lC2UoCGjmGPZNj2mxjAVCZ1srallrm
loqW2bSOsgCpz0Jptgo1c2RI4OwuXB53z3nbDakx78HubKdANgRDlQVXVU+Kw6RY
VGHmXbOqF0Q7eFuKAOmOLKLtOzB+wP80WxebSBhbLSbVFQo35Gq4J8xA15zTp6fQ
xSkzmxDKVJk3ss4RlLwTo9ZDX94BzOi7l4n0x9/ECZ8KqG3si9ztxaYdSzjfLRXw
lqhLFvOx34Sih5wZJ5nCZge0KrdD7HUTIvJ9lC2N+Ye4/ryjFWU8XYj0RdcsM0CU
IwtSXoAfKx1JF/V/jRQMc8ZekT/EJCk4KUD9LFGrnmN1niTovyf7dTrD8u1PXqxM
husfCgJ9hfd3G57+dboiGcVvOF9oFBfjBF9b3e4IrcQ4ebBGwYbasWmS8EbFo1A2
3GFaKDunEr7DiaO22tc3rDEojrMzz/MMEg6srycrvVUJCmZjBubTvY2Bn2qsU2/6
WGMxQnYKWRixHzjbYDZszN8MTPeKTeA0Yfs6Hk1WGFFILGxvjP4S8pCsM5YKZ1UI
hRCkJ+mkBNK7sE6YugwQifUG6TboVxybJsIqZ+d8QknfoL8n2bunwG4LvRfU2us5
EdhTl/eK5Kqf/pFe4iN6pQxiBBqEmCmRg4eOlvLJw3RcrRODFrHsh4aeVGyApisR
kk6FMo5icK1M7G0sDeKhXn46M7wmZhsTjJ6V/dH3SxEsoh0VV8WnBIC9oonJbknR
11GmQzPA7qIvquhSCWvAuKXiMouJRFmOAmz4ONV8ulFGqBi+3/HteoXi/JO4h0yx
IrtkdyvrpsUWt6GOz7coQ7OgoRWb2vNkQDiHx6zmSz0Vxn6iDQs7Z/wH2OigwZPZ
IDn4su/BsAUbrwhlM2Nyg0rGcmInAP/W0qLnPLhpYVDpNkP/AWPE7G1TEKCBL6f7
7vcNp0JEWeOLdHzaLwbjR971FCSZAY+IJza+LJpKPpV6Rx5vKxW55AXcAm4eOnh6
8V0ZQXtqFAfcnmtChLeWWl92TDqkpkYEqQBz29EnVxLHxI8YB4d1FSWOjCX4UiVC
GpNzgyzFouFvnQUJTuPkb5PLalLz8AzlVVB7R9zIF5Ajr/BkCXlLAb+UyHYuOvNS
jUM4viVEGtyvuHLwvTEeMuTcR9t2bWDVbewklGeZkUwRN6W1U35vI1v7Z6CRTZrk
Y/OdQ3IA3XhQ88tKaJBNzp/sNJ9MV86uM/9Y3ZA1iPJccVv5mXZFdrqIQM1lTitt
soMvSeS7UA32nJMgi+FnXKStGAUja03yIAO4e5YwiG7Qbe6LQI+ufzIvNx3RDGSH
L0IP3hba+subyMsj/JXDbLTMYc/VgrOTSCOkIwmsoCV6/BD8dil1qRzVgMlcG+zB
1JxpSjycV/6vofsutWbURjYhmaqhHItmut9sH5X/BcKpbOKAtQeD/DxzsBJHnNEj
cSLfl1yLhhx7SYRQKaxLiARMjbRu2hgqt4GtOTNg/mPxAycKX8ZxeAtNM8G010hS
SKMFtFg18uxARhu9ajDJM3Sba/e5u1wRzbg6xOKAL3eAH3Fso8IDiWiZdow2MLXN
jCKS70/GK/nEoJ/4nd1JhK51Pp1srhJBrZd5B4z1DVB60ILbEfRiQvNXFdF4huC4
3i/ibZlj0emFLLaWhuwwdEBLY9aGowJ0CzxPubuljnmch5mRE9MZuqgUfN/t67xb
XRrCmkxE2RAMXNqqMarIl738MAfrqEf5SZHA+1iGxw67hy0VYJTMPb7qxj5ea/6Z
9LlS9Ck3A2yoktliKlbHCZAt/aS0yCiElXBGovjyN7Etglhtr8iCW7MuDurZioHy
awUkYdxsn83qygV14fWWa6LGzIulfhioJfN0eH724Lr3wQtX2DMWayopZCzI8lgv
SgpUtRITbG0NPZKyLI7vAmFGcLTL/g2Rd3Qt5I79TKcapGIE4WQhemLaLkw8ryKp
OKEiUqtK6HaaFaiNFMWkN3e/wAR1sqV9LOi7f0LAkBxHFBsxvWOUp59qSKjM6/uS
E2jKFr6AWBkU3tXD8oC7ItVYTH+RC4uFKT2xiLiNQpl8OMZNk4/9jliqKrpCCfDG
/g9LyvyyLhejrhu8xxf3ROC8Y50q3AA7Kz8EqezLFFYA4qtABsYocJdcGlqYcbe6
TtrtGib0gQ4C/516WVJybokUK7I+0hZ+f4YAGDYxSCyklteaH31s65agYMqLjgqc
0z9oGg5b1mbocwYyI33Vb86CKyp0KKbVqHC9iUnXF4DRf6MlKmmoZCSSruVv4qAF
8RJXnCHuOBMir3w5c0acBL1od41JgzZdMAu7F0QX00hXUVj9gpSalxw5GIx423tW
uc2YzTo1UYdEekhFVegla4gq7MicoZ/unP6K9UjW018Ts/e/9vGFjjdrtSM7g+Dg
xpE4o13bfTc2lcKA9OiuHYlEP/q5bPk93++y0QKxpDf+u0oL6V9/mDMOiEUFSttb
n7TJ6KG/GWs4C4cuZH5hPoYq+c5qO0zVfBhhEE17qC2hz/2H2R32E+/k6tUOozBZ
hG/UPmqJdYBzH8SLyj6vILJXj2bZEXEKdCtpLAvSg9SL3fetQI3VHegBHmGOca6r
59NCxYxj6x4Ku6ux4A4sFWr17OA8liY5y7ICoDIEwhnXf9vayxBcO4te5fLXPLZw
iR5vIfMpDuugos651QKrUTnUl4mLOZxmHekRsesd/bvfF+YlcDMAKEaD59Nda6oy
wpDrfVulbuH89mF0vLlGK3/oYlshB57qAKU6/SkkwG6Gr2OMvLkkhCZvbabjZ8od
AxaRI3+1zzSvMh7lNW7jesYRjr0iOWmUAoUqa2HZ75cG0Ytnw9fZMIHkmu3PJ5Ej
g/dgBM6JQH0F+vOKJ4sW2GGC3Alkb7YiOVispKO3gJONiXf9FHVbUPrBelTzPZle
3R7Lgk4omY0pRZgjgVL9PSyrTXPAW+taMINK621XlWenQAaxVlb9+HnS94G5mbUZ
vL2xgDfFKugveD2m7BVQYkBda8+JEYsoY6qjwfcXA3YIYiA0F6bnk6IL49xO5ITm
BOeLn2BwexBy8ffKk+dvcUj3a7rZMDNCIfe0xxN27z6UGMb9YLiQg1HkAH+aA7wY
ZBrej4o9qmgjm+siWnCyAnQKxczZdDr6/psKOpEqiJKkXUA6CZGZQRQmEnhoOggr
/7KJC3O/DivC1t1lppLIdGpTWwQJ+o3qikbSKQp6B8sxBGzDx4EfO/3wAMlAYP5M
jDpvtzuIqIutNSnxHpiqotMbq/RsExItGzyLxB3x4IN4Xp03i7JlEwh45OiLy5DN
Ws2NlSUtI7/pdmk/hZnrcxuujl91SVJRmwRLKdmGEsUpQbOUqqnwlW9vPqDhD4Ma
wNvCmBVhKy2ZEKFck1ZQPgT6IYyq/ayGfzchVZUSM/APrUXO9/bV5jvVobo1WpV9
+/pgvgu8pBeS4fC3+ZcDwnWj9bylWOcg/+wwPw0lZf+I10LMd5Y29TE75tkCFxz8
z7at0qrXt5mh322gFYe9T/cm7mZy5MOhwltE6J8BbLzRJKgAsd+9k3+tzIalvGlp
7Lw8sWlsfQKPQe4IUFwGZRBQ4PoGoKrR22AnRq/CzReI5ILJKEYyaVD66i/JzXil
2Qh3oI7uHpucUaMdBnvMxJdQ1MGEElWs59ITUPkxv4j3twG2Xm4jVBDeMdt+onWs
MqqCRjlW1db96AK1jXTJ+PU1AV+rfu0uf/9L4zXJ3hYgnWtip+hXPtzpXpI4NtF+
IWHJzV5vYEoJlvDRpgjdJwgL51RwA25bayCp2LQaGPGqf7pOHyktnDWKf6/i7vdL
jhVmBl/jwEMuTYY470CSkduAD8TyJ6rkFZeqbQx1ThAS3P0amzQ23yeRN1uMVko8
ufmKWvKWwkJMy7j26eWBxbycwIbyslNolbmvnV3RJGm/relJM0SNzRbD7AkvYY6p
Wtw3XyUK74GLaHiHO7qpYKSoCUesYNnAVt76s5GJb13oUonC1mm+F06xPIcUR8qV
HgIn6/+z2yxm6rTT8Jc+HIERVKkHdUHoAAPdECZpJNkwhnf0OEaYWPNzBUOyQARg
6AQUnHkyQwIIcplo25YIOgjQ5FaO5QJ7FL76X8MOwBDdqe7VGHaL/pdBKmdT7BkP
+alH7Z+G+Oau/UXfAbuGf3i2budkD8Eq/5R5Eryt0duR3aD2mDJLhnIz47tto76z
3n8Nt5bqreELSnNiMae+MsCd2XWuFOgue8OB//P6os1xPI4nFzN3dIuz88EX4TrD
x6WUvlq6ZsvbKEQH7zGZq07/LV6OjR1ITU0YuB8P7RNegWIAykGOYYtJxmSdVa+Y
ens6wkdcGOOLaRrCi/gQBjk/qP8wYKGlx2xeu9MHz7UTe87WdXFQdVXyipqIVtJD
TOUjvOCHKiJljZlFC1CarkOztV8BX8hPkI9/Tyfbv0GHWMVD0MT2uezjPK/jUx3I
yNZxLG5+4/5Ymbww2ublTzQ1w+KATcuFInIVtdKZXwEYqusR4mLMdn8du9NwMi3M
hrwqrWiqvZL7vR0R//jqHOx0iAnnGcJhtJTF2jm45xIoXCGbO9g8pFFQlTygkN2b
Ci8l+t413ZahHzKc9vuI43wK7ovriF1RvAQJybQtx6CmaMUA8c/zSqKxSMzL2SCy
Iir1ABAFf1+PiBShX0rzRcMa6fYViED56NQrv7tFAL3uZ4/oqU0pTxMTn7CYY6o6
sZP0qzMcrXRRqtmXkB8tRZLvdcykxQe/uiQuTZ/GrMGCSbcUL/zhqpl9kDR+lfJk
+afjn2EkJyEHM2Mwc2McCIOUv3uMKHY/HvyNcguFusZXbDa5pI7eT5ZKhIDP1Bbx
d+nLLN/YH4+yDzTBV3ymMPJKixsYkZvbXAZ9H2uZDFDumtS4u+xBwAMsBWBZ6cxY
aOqZcEQaTwSbnyw3i9rRyuo0XX8HfGEiopWjZhsTjQFxa4opSeR4YfHau+ly7bNG
NODAVTqSHsMRbalKYL7pp2QPkrJqVi4YSXRYn9fWowYUIUR08MYHn+vhxvtiahuk
XHoTKFOVXl+St2PNDAlm0Zkk4629Fl4YkX6TJXxMpBRV2OaKtqfBeqihRZaySmm+
SPozdqF2O2lK+e5R+RAys39OBgVc0w+MfRdZ5Kd1bbDM+s8uLtIV/amLpZXxc1UF
tBLX5i9Ih6+p5uRrWcYLGcLLJ7VzrqtfLhEG4w1MhsdeY23PTeK3qUEvwyDK/WLt
D8auyfRXHnhYn3LIYMcGJNz0HvMPX2XrabRbZbJCjWj7jVxsawFZnTQVBs1gaElS
Q15/Qa8E9GCFv9X6COlcJqBDEqqXgpc+wX/74ny+6iyIgqZJy0Ci8WkXV1tUeVEo
w7RcNKLuM8k8xMeWhptyqzYYilgLxMwfgz6yfOKHY4JTp3GNlpapLAbO9ThnFsbn
i6wPKqwVagw7PkJe5jfeC2+YxsUq92RiY1pVMWgVwqeobvhGj2ex56U2/jwMWb8+
vTwnmESyQ4M6J+FX5J9woMz+jEDL5R6VmLBXAoJQdv2fsQixNJwypf0/ZyDH2Y2u
rM0QDr7cAwnHcp0C2q8qdDEy6B83RH9pIE20bxVt7yKS1ese9h5Lct3bAOHljJBf
DUu/lAOdtqVZNuryxJqtOxfbrDHkXoJlLrYipKcDUtudOE1Zrd2ORcAMC70HcNwH
CZh3ELb5yiU/1gPfy3lUqpVZ2/8H++DbRPlG8RQynbTHGS4/LTxyrWs7Obua00oE
WG0/und/4wrpRtdmpz3EawjVzdI+75n61BvxTxTIRZcdJdQKN5WewznSQT7Yuski
+G3aWxbdpECuhS/lDt+RESqaXJ/ldvSewAf+PrJiX+x/AXKFTzP55QQaMPdsK87/
salRDZS2WiBIylIWiRoZ2cY8jK2hR0FlPfDqGHP7BSlbJRxtTV5ifraC+TDichaR
kKB8sGG0aIooBj83j0ukcA357kHTpYngnOqGt0eZ7AlMkk0sKVWVdtRvjbOUnoQz
Xvx4/fE7KsWelnlO5yBsDcWpeskPNmJ84a7kqkI+Hi+icNSUpaAFJqmy6L/4Zppu
TwNTe6Uc1u6vtscc9JBP7idgHRVMfLLw2YUl43fT9kcBM9s+PsNMXFCIbatLAwKO
fEA7owsONbrcX8vLmaXjwswySSJclfwOQBINWZhsA5NdeM7JrJQYV3k5KHJE9O5x
SM1dp7S/EWKXYDCUKjMiZccnG3qfUjpYgEtDBnNnjHyv/TKgVbpGYuJE94/JuEa1
7bRhZsCGbkWAVlIAFJ9i1Fm3A9Z4c4YtWNr6ANZiLNGHtWjZUBWRxaXZfZaE1/r5
wsbrTUvdkIPHigJIP4pnnfRax9dzcDd0G/x/AO1r1TDf0C2Ypc91LLTuG9nKdQeh
F/6yQZl19ZmxjAG3i2ih9Wfe8T3Gffx/5bMPS1No1zF0GSpBPnjqwChJy5w0yvGw
GBRiaLXd36Jc4tFdSgXiXrhOk+92GpOc+Ge+G3QxRh24z+HPBWn24Y2PsCxwfNbS
UlvVVuT4UW9EKkYtevsMX266hM+TycSjW3QRJECFnE4krzm6e/4w0T50h2P4ZVzh
uWGBofkpNgm+vc25Gn+glwJbpHlxPWkAZOpynEfSK8jDteViJDRMd8oQ5xi/tdh7
rUrDei0MGZ5B8v9egN2HftjVmu4bOnYMrUJOnNJzeU9DXQQFkGPZMLWX3xQfT3Gr
SKr+QSXEfeCW4TW+N1CwvXWgMNeLZtKpVsCft7R51xQ8H+g6CAcyD86YKQmEksNX
nj5S74SH8xfXvmmXeQPBizyOd0p8awdeTdHOFGXMZbr++ktTdvZWqP3V4Dfa/UgI
610QFcFuPdcsrMuNhtP+a6Ggv7vhGeDkofAHTceK6h37J8bk0HvbKPi2lcSp1uRv
4/lfY17ryzBO/RrTMPjF5c7rE+xBNG+KLJhn6zhLA1O9XB7LckXdzfsmSoYm6ueD
PBqucp9EH4gS5hU4edmv3INbPD22Y+JuDihN4+rbu7GnKR8HKZutAmT4a6g+CR3/
pNvkdAeYkZk82pdsCnrride8SdGUy+xHoogRz3Y1PPf20fVJ94UG91WGoKE2U4RJ
pkGDEKo6PFNK0esug51+6YFuplpXWm/GCRRsTbr5z6qUCKRyv6KfE2HxpR0O/+Z1
HLx39XmHyLZ8KbI1EgqVGBKptRUIzX6WeHyeocmjvwFUoWtSMGg18AaagYaY6lvJ
ujAD0sRuYbK2PvPS9wBAik/VNOOgFqboaTOE6F+LjIRhXjFm9hGlh2pf4y3wasqb
TVeiY2pBjh9eXAp0j3kX1Mx1Jn4nf2xupE/4FvgZSdvDSyuILynENa/W+7ZhJO6Q
9Xoype3c6dRqknZk7icLhx9ng7654zg2B7Sc19BVd+78p2mMnxNUSbNvEjcUpwwZ
fZPlf0SR58XdUaeDyFR++ZQmpNh3TawklVKmSufkfWH3FFb4Ue2jIIMFUeRpydr1
8d5D3cqOmnUWr2jGXNqY/H5EprkR5tHtRGB/lKl3+1Frdd0MCvwirUXSVohalQvX
3jqytqkVMRDGYTHoYMX/sPfWsAlbJE1uKOls0mwl3HF8mFybKMQq2iIPIGI3WZIZ
Ekj59agZJghM6b+v6mc6b/H/obx1MNL0vgs9M9QxUMpPhzh/H5yO1h5eCXN50RDt
SQM1FG5AuWLuHM+gNIJjQbmF9Oynxer3yHB8R4HWbCgmWD2utbl76bkJoxJyGunR
FAyno9inUjQVUlIncgXlyxhMxa+3VsxKxKWGgFbQ/WrXX6z83vp2MOEwDo4NYwUQ
90E9YIM30qArXvRhwkTy91jVJfmlzU8PjsidYH5GTybznzwAFoiPhujDnz0sU1fU
8o66VXKHjBorfGH7muFlaYz3NUwZDaTeGt4HgTOk+sIcRC83Re0ubpDZSFq8C/sP
DIBPKYXmalGTksz9S+4/LA9BF/Dck1YaUNiLWFYhSwKctJnRkBc0dBZ9GiQaXCKw
RKktMaCQdFnUDuWi0G6qG/pDtyOVdRolM4W2Jyo6OehV7i0lTxkIopiHBejwnTeu
a3hwR8UwwelIiFpF2DG/s8bhEK/MPefuwTVKfgCxtCeXdRyfA6RwSCPFpEkzB5Os
+AWMIOJz4X6fxpDqddHw9WgMa9Rpbg/1q65eT+RaaB0DN0pgUe2w/KjghdwaFmym
36R1avh4MvTjYlKcpTaajYPFJv9L00GAbeWxvxM6ZPDcVfzwORhkveyiaKde0MNl
/n3R+CEjVSy6lfZbN5EBPuGTtBxaHngmfv0w9Ys8GTSARIPK0vzY6F58tdop3U2G
k8v7dSklsvcQU8URP5ZWaqppE/GHYYEWglvFDdIt75zzLACDgNcUdkVeiWqgwlxO
1+uznL6U9k3C0qz42I5lry/rhvdyo5D638Pw2xpAk6hjKW390xLv7hw1VCiQL5/2
qY4gqz+Z4wzdHMrJSLl7ABxfRtQ6VYhPG8oO4X3UN1NWW248/GA8gZl8HLLNiIJ7
GLfz3/gr5O6RodhtqJZtaDVeAghGdXaaEvOpd2lIlLaa8eB79QB8XvrKRCjq4kiF
42Hzv2upJfwWOBopSAC9kZsn5S45bWGDRZlIp2BClgo/Sc8DjWwdbcQcMObEJnak
kYsuYcMjslxecld0NHIVL9nOrUzUnMxRsqDcbhse4sArX9GrTiB+GBLyXijiJJvm
CI+pTpltmVU7qFRWLFH0nKerE/e/1B4hEVHcAW5bN0u6lvi4rRloDFIV+ekHKU+i
Nk23YmZKBmDpvQanF/7MVmkv8Rvk5wROcbFMIWN5OxACeIOuEgPEzls0U5DqkMyg
rpVySTUInBityZS/5rzwip9X8nfP8kSqqJbMvAjWFz2TgL3ycIZdopnq+HU4C5HB
DviQmXNCzAkD1oEy8tqoRzRN7s+wsMUuNa79IYxaSwCacEyGh3l9tAHecWrMDPCk
38F5UyWA6Q7TjXy0hFw50bfa6mV9BJOX6vtKHvR16uDRClvryDjO6kk26InNcOkV
dibNuBvBe/3FM54joCsuVfu6AVHoADavBTjNf4qqwwCGKF5ql4ig4acRjFuzjbrM
b8wLp3PK2VbvsMv3jy9OFTJtc99hro0br4jTK3DANd4Ak5Uitj5dS7/e2hqVJLr6
Upybm47oNw4KkdaOxmZjC6bF4BN6/uhG8sCNnb5pX+PzoeUhyOGWlBZLp5gugcgk
vY9qWzkfEcD7EvUWdSRehNs9vxHLocTzYasT2bsedSZycZ25YplhBWmccCUso3ad
dloJX2vsBFCV8bCDmVk/C+XcNFU7aXI3tqvGybObk5SQIm9ZpXwpilHZQ+/WrwIW
+WCrFj4Uw4FLtdZ/znadQ7FPk3dvsAg4p8pt+wlXQe9Ud9i/5OFsb6E+g0ZlN5n7
8en2InJ8+ycCCKlrpk2XHmixbcvmUOwgUtyOvJi6bkIgMzcRTJeN9tJl6YLfOtbL
4tKxpCbXVHixV2Tra8w8RWBxDVPghDhFAA5HBOaulc9dRpQW//7a2YlbmS4zAnU4
i921AbVfbkiOlNF+6FieXTNg7weDzQ2pDwHtvPoHEtOhGzjst5wGeGz1J8FIRTqW
So1Te7kxD8ARMci/kiSHBQlnmXoptHa1WmJWFGsbNQsaQXx73NGsln3iX6SzcdOF
p77sWKV08lvBVK5EQ543tSI8zYhwOyn6BVm1nYNgNvimPLiPdSpIWBLKr9k9/7wd
qkYTEXr2cBulPbFx2GBLLpWbASWSD0Bt6u0yjK7J10X3rEuuNmfqd03UdvnO2j3i
dyIoQjdEuphfXynbHbvjytCCmsND88XcPxDO95TKMLY8+jEHcxbFcNPkuswUugbN
CnHFtufjDMmxYksw5FDdLKRX4g80O2CDQV3EzEbRxDwW9fSBepSGK0Z8Fjq7xpim
aTGLpKN2QiWcbeKhPFSSrdpb5K/X05Ji9Jdi3FZ43vC9InIYCg1jWJow0hA8aG6N
F6DNcCwovRNUPhudK6AXlu0HGUggKRtZKU7MJO9xAWNRdvhoHwRcvXOwGb2FM1Xe
SFaw+PXLhm9e4eiFO2ICPnRNTikFD37I+FVuciRsZjUE8OA3MExp3srtW5fPx3am
qR9QPXp09b6m+iYXh1F2wM61FBT7cMpboN4LRfgZ55H7xvcTCC3qdhFDNELr6AMt
SBy7kbw3iBkRMmfDUcuSF7RHPju9t2O9ApGlazjl35hTTRt2TCB7ha4iJk8gY+qV
P+rsy7F3AdwXBBdZXwKyWTNKMQLDx8Gk8obu37VZjuJoXdv0dUaAO3W+D7/ZLY8q
b9hPfVU/58+ouiw23t5hOmHqrRQoTuQ9FCfzQQAHHWQcq5DAzKUxqSoCqgWZ5j4l
tQVLDgtoHigjRWSMWusKkRKtptyryIS0QUXW+MWZnol5vXvM+VjGVvOdrfOaQe7u
6LQlCEtI1/IE3bt8BZuvqXMQFmJbE/4w2dcp8JdI85FbLgrWrciK6wXUM4yC33kY
4T0tFWN2uNEZHfa3VgcLLTNaDhaHdBmrfX3TKa7HbI73W0FLL57I1CNY6mIiT6kJ
cwFFBPNGmfCVOsV7h0XUlX6ep6ZuBo+5yO3E1jzhubxKVTeIzEygby9mgbeBouTL
9z7VztmzHm8f4wvzeiK0b2qGICaTmICgL3ySL41zqoSfzlI0YLTU5b4bI/NJj79t
pmH79kW+fNNp2l8ghHaWUMJvCHPKqzwPjKqEhtL8aUfUI0h8n85nsFD5fnMztkIz
47USsRz0Kcf2YdRld4739t0OaYAqdqVuDbUn05RBM7Ab4Z6dqD08uSYBocLLJbHd
inTz0SMejVorIol14p3fxLPsrltoXjvt1iav+oBqLqESwj6b7wlz9/JcrW/yzOJV
16UsDj2Fnb/XiuNln0tq0Q2GvG97zkzG7LuAeSVWMW9omtYYWZf9kAo0Xy9Mv+mB
e4f4MzdBBnXreEWLUufG/rncnbVokzW/4BIds9PQ1wytXx/zaiOkk0XAVlWQ7BMh
/1Ms71tfOYi2xDYm6KgElZMFC53oHVTM7NewrTlmXrGGslq71JUPPG0BVgccnwGq
mdO2SmbvnQ8xHeh9uI0oW6F+MznDvicnFvFfCm32Lu8yZh7tzrBfmiFoHuW5H2jh
vqSXRHKJUGG1YEUDnPEmgFPB7QrqlBjqE/yke+0Z7R6pOIWYNpudoOD1P8CvPa8H
60ob0/wcvpOp3d7DHEcCX/jWZIFBSFAeEts1cJi+64/SnJOzNgtQMbvj/o+LNeFu
wgTnQb3iOP8GwbQmkry3zHHV99HmV6FVFvZa9q4iMy4p6NZ6klotkGS6oVGpHC2H
w1vF+MqSwK7g0XbOFkL3kxVuORvTh/6f/8a0D8qpotvlJt2XC4aLbPYKDTOQFn8Y
wQsl1/0GenuypsJdnEbn27MT3dFCk8WG2kImTNvgyV0Gfte7D/0Z38ZGHNhi3c4A
WPznmE73vOKmX2AT1q4Yq0AUB4dEJ9TmwkVMP08Fw0NBJ3hL0DWx9rWViu6lL28o
YkauBmXJN+2qyCI7IG2DQdr3pmrJYSMjwXueocBDSyMNnB93sOZMBV4q9DKlsthk
y0O2v3s84ogpITNM7TrXkYgEXsDppK0G2Zfy5n8VCSJXsUO73FKxys8CKOMqodKI
DadBUaXfaGB7cU3D8VIYlXIoVzOzIwjvolKsvR++mWuF5WCVAD76MnQEgNXsyXMV
uJwTBsLNG5+CgpDEffNOfDorH2mEjRHnV1R0m66hJmQa7b8lL+aqHvi0m3y0QIon
6wfYB4y6yU5jfcKZGoqbCbfo7SaXPWYt0YWa7F2ZRs3NGdTE8U+PYgJS+GkXWXw/
bZpcDIdGb9+GpCUNlO9OVYpL1ayC86KSZQe6Z8yMsFc0J1BiYuiDV4lz093DguxX
dHeGZCeku18qUejEosXps9fPmp6QyluJ/Wgmql4f1OYx2W6Qqw+PZajwc5UZkEMS
PR//+yr1/1DVPkgdpk3ccQfRkC6DTOepOSfIdMVYtPqc832hWyo/ja1ckqYeJGrc
GjzNZtCthZA2Q2P4DcIQ6lAaQwYQtLA6vX0BHAfVPMjHbWhbTV/BL8KLZpWYdEgA
/gnisg+8037XBH0LOsFDFmieDNcTdzG6sRe1rrMJQAUpWm9L+XVkplsyDPSh2NOQ
sKvgt3jnRC9oUMhSWVTd/psL1OzWjN/TxdpHMzeckPHvDGac+B2zy5mUU6b/3DuH
0ZiIrPYFNtIEy+8Dks4GT6ss7OeZUtmD6Ia5D9BVTso9teswqjW8EwCUiEItAB9Q
8RAr2ESLxCv8F1D//9LDK9iQb1N2zyemCBkUQKD3Ypq7SK+TjWpRsMaaCaOlqW/8
Vxk1vt1u1IC6U9Q1ZN9oQn99H5I4vPrADXN8XcgxXLhRHV//OlOtPgxZB5SovWqO
RLHDgj54K7deNa07U3CQpnIccJvJalGKdXX1Bkb6NF/88ZDlAyX09r/rx9vu05Va
UusnpGaYwbkGVG9EHkoI/8sahBV9k5mLvE3JVmQMA5rs8IWwXoVhDL/g9cVwrGVJ
rPuRJMsMkJYG/F1W01rcNliFzR9jgFdV3UsCDUkF3HYmndfBaBf5IxTYnatOwO1K
ep32SM6WuY2iL3m7kwQWOUAFos9bfIdcKDtWb3tJv30NGi3XkTugDgZNBAwTySCR
6rsl+ByDT/n+nWUPuPZHTow7KwNfnTCh9PJKsbNgQuEeTFpBwirheX9hDyGtWdkb
kJoNRMplOnjnmg8zXy3ZieOkL0SuQIELF1QHVUnzjalpccooW+Byuzq3FlDSQwD7
LNcQvVeojMmOK7hG0EPE8K3ThXfMASOvOpkJN00pBNX4ejLfoWhngguEDyyJpCwa
0frua+DPx/TpSabSLc7dGu44k+/wb8OO2FZgMSi8CMFWtn647WbiNKhbgBMzrD1W
0plbz3iUR+TtiaNKdsd3MqvMYcr8AFmUCVLeusZJORvI+8UmYt/VkTEk8Nes7bTJ
wBiFNgRFNq5Vb5IRS50zNz+m5nX4xczVbfwY8yOc+ZxHOQwjzET0AJyl4Ld/UCps
FB5gM0dzJir05vudCror45gIUPGDZWXdBs6HSLC5/CNLRu8a+QDwL5pK6vbWU9ib
Y3Z5m9IY28YA5n+yYRE6nFtQs2QtoOK0dsgX8nXts5WwnEUXZP9XqAqyNJaRBXGr
fEIAqq8NHLKkzkQ8laQQUWyQDtNP4Jsai537BSc1Rk2CSp8W0+KFEEBUiyMleP+G
sz12lwMJ21Ax8AoAxsoJw0nD+up3qn8dkoP1uqjqkqiJCL2Vm00rUAuHSmLk0oKm
st3IFv4akTR6aZSTJYmWecLFQRH1aVmYECWhcA/eSRzH0EBZxsjawnmXzERN5WXG
9usR6EEJcxdHL/gVbGlKWmKLZnY74CGhmdlAFc1QaB/P9I4lWLxqCo8tTwoBFEeH
hdxPYga67TgYgBzQiA8d2WYgCEVYIbAIYDUjjoddFKaI41f4uHrclvkAsNhHEKnI
8NbRlZ+3Nla0c04oYKj3twKFMJq4e8Iik1pwmEmxb531WPflmjSB41AsS2z0CFlJ
gANvZne4KTxzoU1bNuazL0kcedffA71NWEoX5t/1j0dUQWrPUixHfCHEKtHyOOrX
dVvPLlvquZrPhn6cuLHaMYNzCR6aCeahkYgSMMthfgNnR58dyLVhXWbllyja4wc+
hXUuvHALLy/xLichguEc2zv7aLzeeiGbMSA7u17sclYC/DreMLik11B5rTJY9XSJ
RxDRI8mQfRsB5722GEQxxA1cxJ27ERGP+YnEKtdj5sYyrqBtL08N/StkPTqSTagL
ebFfyEzk/Fi8NMzEd37qE6paDINBFgHsukgkpLCKOz8vwMvX9xUG63LjIMv7ojkb
SUXGloJgobNh863LGY3IX1Dsst3+bmXUdVWcEjT1ThtmJ4UmwTA1oh9/VkjuLOg0
P2Ik2vXNJjl+oATIyUagnn4HJwLonR2nRAuOluikUfuFFK2ADhpM07jrGqFNVivz
txopdYR2dZyFp12AIMVSChiHvAhvZSrVoCGknTSU3/K6e1o9hFxtSH3UMYOOA+8f
BfxIZVjYz98fsx1eECCJjhHOodkDlpzTOv9DUjzVHY87Op1Pzq4EZMfyPViKEVG5
yHKRsWx6Uexnez/FGRN9Dj9Cs3kQ/uCv0FwbbvxHa7l6/+4//vo2YU6Z72QkYI+z
KxRMxWDQyRfwZ99tTlcSv7ERCaqLY0AyOz0Rq7U4ifjshvQvYSny0IotqIpTvi4m
p2hayjmvwH4Hfry2ZhySDLiVBsVC3kblHr6L6lAdOoIjv+InnkujewbDU+DWJKRr
cEN+N+dUs5tJklINSIjgTEUh+M+2gJwwPJL3OTVN6hJ1udA4eyB/e5Mn0anFhgDV
mWuUTEQxqt0PBonqA9U06PmzFxBui3fbJXJ8LGCEEJZEF1Yz/g2IyfAo0JvGwYgI
sXwZFOits+uuvkl9e/HT3idw5x+UNeDfwPAogLWEF5xSshQy8ro3aUKl6VS8m5sS
YmlragPB8qZYMMSqwELdvsPE5jqhP6ivRyilX10Y5rz3JfC21tCfjVVOxpxS79T4
jFG7eX11vpnm9dcamCPENUgt9pUpxJv5uzq236elKIk+Chz7PBZ6fAJ22zdGA1qO
klHUKjH6msWvM1tH4HehExDLMdcSgAQi2S6WCbkWaMenZ+oRMfcIn6mUk5ABP9WK
gnskbJRzf94fYfHHKWYcjXwB5Oq8ZpGiw7iVDoWqTm2No6DVnXJfdMXj6a6HOngA
F50IcKbje62khP7k/bUSi9h0mIwujE7pzdT4HTh4wLhT6Pgjvq02ZOBPNo4Dd/VG
LHJjSsjBGgCpj2QP/JVqRX0wveXDnh8d5y/V1ChF8AxYm+6vBWoDmMPRW5WubKUj
AspXGsZSRN/DSsVIkowPftZgRPRjQFh5tMArqynwPtZ7Ax2drivnRe41YCtCfK58
7uCiVUOXuIA75hopIB/ezddlbTh8qF/39VdKeQx5Q3i5S7c003xRclhe/vxoM0ko
01rmTbhhVDGVKAXs9qytqVJO9mtTycSPeSR5IRA5hgGcWbg6ZYh3Iujqfp/PhgUr
aWUgpY51yCsuGJqdH+D5+GPRAcALC+FZP3Y9Dth2WHkMRZrr4ai1Vy/6/BnpE4JP
2gj8aNoZMJmx2qexL8/YCq2wfNcBRP74n3XK7+UTkDHPo9o8oTRlLADCA1lEEBn2
K+8PrA2DVnwy5c0FmCeGyCT8LbJO1lkw/cw5/xeP25nN/Q/oRY8KwvGb5isEJNmW
x6DNXZKvlrpWLGk73M2qfdR11oohCFcVNIl3fbvAhVwe5jrFPEfg4kThvePEbXbB
3v+Pp6I7XqJzXb+Pa6KY7E6Kgh9d2YrVgEArAfwQfuJ7cFIskhwKiAGENGMEhaVl
aKXpHQc7vPcYw7Ydjo/LHJl+JTB9bifXqzwoILE72GyMOLgeyuSGPZv1DaDiQMAf
P40BIJ77jxROt7tWoAX/MuLe99G1Qr5rz6UNh9dePlCEV2/zyrgbI5JXMeWvcv/L
V4LeD2SOuee5ahbh4Sd8Yww8o3kCAW4uyfp/LQ1iFk8RFupO9iEAA9Ya5jvfoB0j
ysKAsT5qX+oZJA1l8M4+o2eVzQokr85X0euO/WxtVHm6HfaXy3X/1ObaVv+YoY1p
zyLA1eYG7+xArD6bTouR187GeIkmE5yKrPlqxC+j5vGIKUOqb9M5r+5baCSmPpZa
0r4Fx4thOoQI3bmsYjRXtotjJO4KtlTz0asnm3ZWo5vCFAPinU3U/pOjIC5Pz+u2
LqZSFWwU/t7U24BlByTjzOINRnEWw2kavVr3o36LG/16+Z7zYrFPvmDivqFuzJ5H
TfS0EYwLiRhhBTvbQCz5ie4MF/iw9JCEMZvw5nhkQJp7nA9q0z68qsey5Z9WfDr+
JnqwoO78IJTcuRhyVrhQNQbIhraOYAejF6D0Iv+EmcMZTT/Ns+HL/493ba6agqT3
9ujDJDQAFMUngQvr/t9vNkEzHGnDxBtp/Nrl8RT1gHofKxTgwXa7hta0nThlWtkQ
/8M5o6vHP41GqIpjjf5lujp3j5OpQWfpSft8HV6Q0KXjZIX5t7axgfqEGXcnshBI
KqJyYIE3SiWORHdX2JrwVI/Buq158xQ8AuKjm8jq6ZVZ7DWxiNGyEOhiqJBQDslk
DWp4LGWSUx6ZcMQxuFX4IkWsT/oR+MSlrCWZ3J5r8tf6zszpQJIgEjVANOl8BxTE
NhBURaRWNvGHMtpG7z0Fr6zK44PZQAfMGTVRgNbndHKfrTLj56usSA35lY8vrRLC
zCIq0mRXQJXqgQSd0zGWB5o9MPt1EU4TSndsltPQyql8uqlNqY5xYGvnY1J172LC
LLATg/G+FFeyLwVKrIycnsHErXkdMhoG4t1/jSgHXnD0LxcIUCxflRCgCMaR6vrY
2Xf7etd0RnzlZaHw62MFWnbUALAAT3YaetuJ9RADI/5t5d7EJrXjKhcq8j1SOeUs
fsahYJ/bWYMpDZuyBVY14Go0M+khcKN6H+aDZVptqwkFxnTsjGo2CewEgn1ocarv
L7Cg6iZsYFRzo5GuRfzb89+e1duZ/LCPFxmTb4O9oJ13Ok4yhJzgcHfW8w5uMyym
xY4gKH/oFV7BR08fLl08nY37acl9juWREt21YZkdSa4kKjxuKqdodBnDHx98S/2r
MjmzowbgDSJHhOnUX+rbCnpssZtAFRivoiqwrA2BS5F7l0EzpEsJJ6RHlzYu+62z
9hUhKapDOVAl7gStiPjLbt0mYkAz1GeQF0O52wSUBVBLs7gNdS0GJemQYb0t3/Hn
3lclkiqAc6ovb38uYIyWtYKJSDMdySkB/NXpQF7rmZ/rKgjv02TFr9nXPU03Z+XA
Vq3mT6bTVRhBeO1hScobgmW87omBMaJW6SiVgrhIznb60KNLZkKNe5FIS3hQe42b
KD9gKApyVMpPz8T2ubRDqHqEuaroY9IcOejYgAvckC7s2vvu2EuL84LBuyR3Cgnl
KKQSoMXuvNI6eYzFpVDxroMnd514kj+PRd1ZIKcwBDnnFKrcEV9pQXWLyPuhs0tH
pvvY82wVluXh75ttb/qB4I+uR7/dHCKMTOkOjzzFN7nOo2jyNYOd3zK+c+EBJDy2
p4ztw/XPJjIeoJd2Lha3fGryrM+tIzplGUqWLcng9cNgMoQX/DxI+O5mRJ7Q1sRs
/oMc1xVFyhhx0Hzb5NjO+VNRA4FWqqRrx1wmN2quZFsW3dWB8zTijZPnJJ5hRpQM
TwJqUI8L4wVlZXt1HB18CdDXML/obt1mOKmPx5rfPdoR94M0sbCNbPiWwhvAvfH0
9+MEQCp8UUujyab5wLSo5oHWN2c/3voglliUHIs2Dgd8a+K4PBhjHlatKb8M1M1x
p5x96b3eyamOxecVbkhGRXCvCq4DNg1aN+PVRj5G24Z24CFLQBaVruBSZ/SStGSm
/NDO924rf8eN/JTSsL7nYtmnodtyjAuXOm+uAHC/EoWwuLN6HceXoY+FFGF0Qkuk
XT/jGWxxFcW8X7R4oPXEzcXWuzyXUC+Q+SA6M8Gq/Te9qFraWsWTZOXE4r0Wzk/L
xUZBHIBBRizfzd7ofpDvOntiqgMjz7vHxZTLxUNAmuHsitn0uNqv3ZPeCBI1aSuH
6qterprph4Va0yBnnX0pHdX1y1xys+FNG5KynjBHVjhJOn8u0t9U+BsUsrlqTVQm
FiNPvJjOuchZ0sg64S3jQ0p4XYTqjTIxZ8bExrQJbKJxFKcRAOnyf79Dth0jDvkM
gAssPKxE8MlB4XHXRPYVg5lVlFt1wOt99W4M1H2PYI3XKT8noKJSAxpDbuaKBBe+
V1+n1Qrk55vyfVU6nOYCIXt/K8AePd4zSgbHSBET/xiZyx8LRasycVWbYY2rOStw
NpxNJ+6ByNqG5jleHbsjqufzHClNSxaPVELEnHbGRvTa3yfibqNAB75k9lygP4QA
bnoUq4UW29bhLAdbc0M44CPDLoiJdJxsJ5WdEJxRgzrcH9ba8unqoop+7WEXIoDj
O7N8aIhc2Q18QJKyTancWGGTbAy6/yW/UzKeYWfJSPB4EHr7g9cK/37MfgQMviQ4
zDaKgeOiXNFJMSYyo6pYwzCiHrKBrPj6f9Jm4JNFRwz19kIgANYFMb3TIBgfGZvy
EMkpDf/c7ycOTu1iMgorxbxWAJlutuxjB5bx89tItjlp/0+yiN7So1qKUv26PkQu
gh5+4bF4f7Bl6sqcRC/hVnEZPtl/pY7rbCaT5+SreEOP0Zem6JPKHXOFgpi9gwjp
cPMXHWtMkEKE8rCzkREHLY5M7/wxxCi/TJl+nZ4BlhJAh6SMe+vlS0nKqdBSDGX2
kYHBx8HuRMjYwCwkeSlCKrchGY71SwUaF2bIDKMu42rVjiJtkLf7YEhZLO/WEGPI
hvSvBxtPtfzSn60cOrD+42Neaei9fWn8xte6p1oDDZKiNVmp3BXpkjGfBDTOcRSC
UsJrYBU081hIdT118SZZtaX89UPKBaIT1VojdOo6I+D9i/L0sEmQNxFo7UUqmJ8R
XRNzD1dAP5gu6jSH7+imX3wYiNksw89O5wXENyNOa7ge1KClLpjWNlO6p6L/OV6p
loxyj+lOCMjqRPapw0IvV5mat9k9V0spAey7fI9hHWOJZ7ZSnEoD7k46M4BTiHPb
MwM/CMTG9o8HecBOe1umE6b71bTlU7/bMxFI8LEpoa0Qhdkbusd8czpP4viYtuq2
3Ez3oGaX7bcovqWLqsHQ8SFh6Z/tfiMm5ZCwEo0lLe5TCgyV/3Av6RR3Kn4Po3UO
EUubUrKpKWjomuDrGBh0KzrN6ZjYIDLIJxXoCOnp2j3gaDx0vz9v9rLo73NmwjF6
4De3XlRl7fhsc+aM7F6U/2JQuHQHYlFgtum0cgqr0zb2HJDWZSWmj0nJtUnkQlXE
yK/OADTtzscsQ8iGauVcHKZDY/koiqZCypOpBFezfknHM36PtjK/T3pKNwVDrHJ7
Zx510jdZE1GVCneMxvkbSc6tMxnp2Czoxi0bNmSAFcxMt7zOY6j62BgHlRevF3AR
hxBmOdz933R9dmEDbmvJGPVH+wxlq17Y8mgrYetEq44ibQfkbVVX3OlmfTQ8eFUu
xYrnlVnmoZ48OgyFwY+aOvd1d8b1zpA75FqaU6/DBgu93BpEdLMi+UNZfIznvyU9
zRi4MmDYhEC8g9td31/EjSrG3KZLespRGzYUhU2FjOxbtrubYKqU2uJUcsGkriyF
WrQPVQf3krhKzR+f3QBXpvbj5/BxpsgVHm7W2DYbi3g0eRJBRqFrmFZBF8YJ9+Nk
pSa7hgjej+lhj5HqNZgwV4cQuvRhe90TdFFyOcD4GyK8G6qn2pny521/c1X19Ofi
EZiaSud7uvvNatlz+Y4qA+ERv02lATb2JkurNalQBF4vEx47hSTtGu0R7h+OuCcM
W+LF5gI/pvjR87+7niVW0FhqAQ2Az6ocKS9/5MuWAimQ7pG4OWXWDzButX5Pdwjr
oRy2uDo6+/yqU8PcRTE8u3BZhtPwof2c4UsMK6xNKt9sOsZPUMgzOTS0ADzUme/p
FbATVKpNjunObA83O4AsfNFpNm7p6XRssdkqoN3wWZdoCX8jRiFfGKyy8EtLH9WL
LMZ9/nW81HT1ycYBGtNedNZENUrtomSXFoIlpyk5nt6fFlfXoj70zYq2G7CDXA60
FUs3FYlMWgnL/Hay3s80AyvivrmtIKnNzabUb+PVcUX6sX0qgqEtLiG59wHfgFLe
uJ4C3uRvjNit0yFE3cfu8JcDrQRC8mlc10HBEZ6EEd1yqwGdvts+Vntc/a9fg4ah
rqVOoPdiU8p7DOsqavyiisAem7Cjg63DpGR/p9QolYBuf7dGuZ5vrFa7NLNoWakc
Gq7FNQNf951j9oz3lTjTExbxsnKi6kBShZIiQprMfXvPcK1nqtoQsgeob9As+MHL
PP7lhZAvzSMc8wEtWqGNXUTW/1T2qDmTYGzNdJNYwMFRKtj23z3bWo5zD+xRDPNZ
9qKF8XAOfuJNV5nK8slFfYpGzPMLivpSP6NvYivkY2Ig14VUwd+rlRIMUSdcIoqj
myJsBm0+X6X4HFZ/tfRDso+27cbWyMkzNW1x20EjKbdlSihH301RSpCdqwTfzFRu
p8J4wI+/fBNLwzn0bl/vqs86qVGi795GBoK+I+EKyabuYwdKMp7PXmN3VoTVHUOY
u5Gi+MJN87zQn17DvtL2xZwkxQrRmjCT7FhJvoZfGuauiV02Sl4HR+ouGXd9VGn3
XFq45dOY8CQYUa9Wt7lGohfDHJjdUM71WOqK2drgIbIB4hmUAzZxHvQtsH1T0F2G
pB30gH5BAWM3I3+8vulgStHCactft7vV2jaRlmYSwwVEah12vWw9qHjQ0IpUAW95
GdwKB5FRB8icaQyk+mqeIORvwH/rsUwyqdderraSQpPQQgTURkXiFVDhR3AtjyMC
yC+TAuBgmRkdf9zoq5UIV7WLelOZl7tU1TJQmhwFM0o6nKesMIO8n84r9atlasKP
C2SFy+VGy02S5DOq9v/aaqd7s93AgQZjW5pyJ0HCjMjp1SdsXcY7Oj5Bgk7GcYQC
BchJiVZYuuXZMmb+uqYpdIVI4bdsLZXlACGAINjbGdQ1M8eITjacDJr8bWj/uSt2
xtNSN4Rz+GFXH9qT6U+FuJrFGip9Bgwk9NWWPBG51XbIqNedfL0MYlzYZtxPqPOA
H63XRsQgBUajq9BoDpdvwtVcC8T9h4Gb+EQvnuxmtl5yJoRYeuKB2bT3A3icW+jC
hI0qKfxJsrrVHuvU3V4lRUoUotsxo7atfUzn/HAM8jxdqbmjisV9kaQyOkTvmsJD
iep9al1kIu9/2v/3tTUU+XEsgqrQkyKiSHS6sQ+u1WnWDQVYBvvDLtkLVqGgvP4U
MtNPxIh3XSLrWJPwaDsY2k7zh+Mel4wR3SiTuC75P8FX/zMkv8SzFO15YnSm5VVf
Fn253Fv81Y2jja9t27sa/Hu6uPae7Nxq8+x+7g9YssDAMdNECphr/dLE58RwOkOI
oISQXGOrga8Kloa2GwBzl/+ksXvvPXyaKRjSyw5PpfJRpZaMO+ZxhGXcs618Tte1
TqWmAsz9HIfQWm4Jx8Y+8CqyD4tBHky6CGUuBCjTTNG8CfsA66/Uvc4tMBZ+TQDj
eFC5z94RvbTF+h4vdMqxsHgPOgY1SKyzeHOPIpoCqBpWJ/K9HS6PYN7urr6m8NXv
f0y5LKRqESVWRk576thjVBoYoAHJpLAAfcSGW9nmP8iWHfhBNOMOu9lOoOFARr+A
iKQEvs7odpimC2WrwoO6f5yFGLXV7eAu5+eEPJxi4hOUqxB8NnYx8vk7qVpI/2CM
x63zQSUG4ZzTY4v58Moja8scEURorVE+dKbs2OGU87YEQbj5I67cim8DA9ySo94y
0seNR9vNCNrw8ecQC1Wo2QU121X59wlfXhldHZLtjWj1RZJdt0Nlstcjzmawzm8T
zhDSGweQzcj5KAUd8Le/489UzsfiGXJaDQuyqgcrtH9tuy+u+a63rWEdRHgMgjN9
RwOi4KJOaKl0JzxnoVABFqw0OcLPXW7NcmvF6YV/+Qoq0t1V2Zc0GzLZC+Itebml
4nPztLZrSmZCpmtOpLUdw/v0idRJ94hJcVLBS1v4aUhU63NOCcJXeFSNUtyj9RAb
9oC//wAsRMYsvGFLmlRjCubXJLVNZydLdziDy/mmTcxFDOlYzttU9Uc0ePRR/2Hf
0rVnFQg9l8wXblyUnKa0l4LxRdC/mXz7GNF88UgkTli3kagaDDdHgtZ2VtUlVnIH
X3+XLL2g4yi2nfCg48ObzZsJ0VsBC5K4Y/luLNkEGMQcO7XwAQIEAkaeHVtWaHdD
yeRDeIUU7T/SfzW/KeAa0SaqrCoB5uIoe8nhtrMR9Ex/xXD7gHydK/4PeOohUPLC
JadiFgQHMF76xi7j5n3TwfqeNE5Q3g1t4FUMuXCfMe5+8ndiNozWg+2X7nB5COFZ
jLvHtVhE6OGwLl2oSqK//6t36Oy0g4qaxyBh0O8HQWzAIn9agBi9jc1U3pnjkbDb
DBvYYQoPemKqhp48SpW2tyXz5ZJqMk60i8Qw0EVyaJGgHg85Sxxo3Sjk645aNxec
krPp4Vvi5uHewuP7S5YQQGXPM3U25mvIVlEkHqf4FW6M77V9fHWXUzepthQ35IPX
6CqRhgxB/yRfz4DiKhjJSpEX1Q09/AT6SgHmA2B+BlYXox3wFbwys9pfn8Qt7nZh
zQCgBonfSIhRHcvPbFovlgG1f4OXS3fEXkI544hiBzl275AESZ2O89kFgwhdPhmy
3YPawdRdmAGm8Kg53xEJrjeNd0y3kaiL0ruinq9tdADvolYt80VoLi5SmO7LYW8Y
VPUZ45qAxeI9wvZkys1E4kyGyTuwkzdIILP4h8AS4rUzHIXvn4gq7a/hK56LssvX
VabCFzHFg90cA4oJOLNgQ9btLGMd0PZraUZ5Z5Jm/+5ZHmLuNmYNuYUXQechlj4+
peuN0zyp4zBQ6eSql2uL+k+qQtWx7Lt1bODCi2Ynv5losHeLAKTCnYuFHEM3ZyH3
Su6DxXGp7z8xJfmheqMmRfWi2yFBVKIADsET6W3eB1RWicUxPn9d+c82tmsCS9xy
b7r74PqbFuWwYXcfOwGwcr0eqbvos1WxwBAsXiwoMkxgxMruD0qY4n6GhDe/ZQBx
nksEZDYcELPESc1mdDGT/pZkb8qiu6I3lj4q2wEbxvFtG0B5mUT56MrIBC97QzRu
XdajwMpi6r4vbdsLM4Uf3kt5K8wFq5Sm9UzlsoDtyLaK7nzcTV2tbWNxi/OKXTqB
tel81OIJAvyCU/3UL0GUFBxLNT+fzpcPIbSAJ/+pPvfu+ccwlRky5fV0bSo0wKQI
F1KCdstJp2e2/1/ZY8bIHKwF+M1uSl6F7tZQW5w7RCdNpiLPJ4DrRb43g8/Kb2zH
V2CdVb5FrnxZMyndJUrBH7jw3JXBI7gNiX2/AjOoqHyNHFgDICOtBvQ1Aw/egK1f
+DFeFR8nkIvsCETzxSV7xAD4VuoCQh9OiqEtOTepjLhmhOXlQwDGcGoXYcBrqlql
xQWsYfPlegYGDmt9MzUSIz0mRE5d7lOqMniXdrkN3GWrWpq4pbB43+BIKcavS9hN
NVSJDTvPujcprxa8AjHlIYxjtGw7O4GujZrh3KOSRB1rr9Ox5O2lSSS/Ueb77Q8W
e7DbaXMfqVRM7QBVqBkRWgHeACe/UoIBHQ0z61voZJU5RdTKHgh698TP03hhMZnR
cZL60e3UAxKGBKFq9dYSy4zNaZ/1qYgrQHiOUYJKsFz22rSVOUatNHkFbRN/zxCd
0ezzB2R3xWY2+c0Gm06nj1mybmxdxC7/HzRaPOEfQj9MHIwYr7otM8xYv+N1dPhG
tQSUPBUag2kwcXqGWN/qj33/qboyK3W8uw2j7/3XBNlOn9vzCWd3UjYHN8W5YB/k
xLwHOhq3nUsKCc7eEYzXmX3PllqYZw/x4wF47j+GAjVHPb8/EazK0FgAUrhvM1vH
Hoj0gDWEFdBin10A9YNyECn7SojvZTUPgg4gEcWKTgATsHWl8IkMeCb1YzHv5/RY
VW090UIndeU28kS+m/l2xyVgbdj7G7WB/gdzV8alov8NbBMLeLMaoIWXFYjbRx6f
TVNJmd9dDmwjN12SVBbL+BKQEoyUEiihl7NyM4bCQfCkPxNP2RBxWMg0N0v+ypk1
+JehS8+0s4UkOfUfmpv9fc9qIib3lVlbpxG2W08f0K+8v2LMv/CQjtqh+DzW+yc9
Vnq6Ab6I/j6VmD0aFSEszgKf1J1U5vB+7WzXgFegZwBhHJSWDshldkBxRq5g5SrL
NFwEOqR1crlyNkjcJu+jHwTBtt9pt9uxFbhm2yq/WGOP3Tx4KgrRrRnB5GvmdO5S
d2JUs8do+nkGYma3deegMYxxSV+Qo96Z85hFp8crA4V1dHi0ySlrN8zllZUIM9/Z
5MwrwHpBLPcQtJdeILux6pK7ux1D2HSB5ePLi8dPOL2OCJIFdHXSiEv4cqJCOIn4
QhsoK6KI38+7ejU+kWLTM0bHcPjU7CaJmblAI1LyAv9dmKLvt0RiEmh559vq24/2
9/JUBwofmp2tFyLRatNXDcQm5mVz8mmHChG7OiMgInwZUZAdbCYkZ6TBu9k4rJ/O
s6hKnBVk6fqpnDT0dpSWUz3FIwl3no8zVH3XHepIP3F/j9MjZoCrJqkW3cg6DM05
Ayzcof8BbgXD2hQxzSJEC/pGl0WeUq86tJRFGKRVm8wS6y8hrwWpcbSv35bnX3Wc
OglG/u0O0huSZXpVIAFht9ZZ1cAKXabB3kyyrfFs+mWKi+k/IEUaJFrVZi+kbL9k
bHoUhG1f58ls/pkMePHJ/ToKFX7JkGnvyxmmgiIDokNY7zIJ270PFfZtPeeiChGR
qZsshKkXCv3/ap9+4mZv9P9BtdPS0sYAddGJHUuIjKQhonUQfwNEBqZCvsaiJXZM
Z59spdI7cginqlYlw2gMDH1V5Dr2N+/J8Znhmrxs7iYJbujLs5KtLV4XBFt9/Wf8
6sfNhXCYTLGZnrAlv7o/oH1Qh8U7kG9eUAcXtzM1OB8BfH31qlR5zOJJ070gFhbn
ZzyiSRUO+fAK/yCB+SC0SBElNPVvhkG44Zfvg9Fj7JowHe+CrNqP46TjtdgWjHoF
qTGPSBPI4OTORnKp4iAC/itiraAs3XTDng9QBxjgmqli/uCnPro3Xqz9i6GwBfnV
JGJmW3DWHbRob0JWKwJIuVdykGmxlF2xs3GuNr/SZJkNIFx7/shbwaiRI2eUTRxs
3a7twbLtneefu99NYPrFR/9Cr2Evpz9+ScXw9klQ4YbHxhLEmDgPZPW+s7OpJiBd
BZSo62dzSrgwJnYwZzCqVI27vky84PoQzQl+NwSes6XVQ8EpO6r93objhFyHiyqz
gVNH5Wk0hjUnFqnSQ5dVV/K+XWOGSVKVkHSG9pYAPn2oANM/UtQ6E32miXGNEqWN
doiYTOwUz6wVju/SZ+OvU+oepf2czl0s7newd7yYh8Ak6zAK8GxzLVcCxq4T6DED
NoEb3PKiQ+f/rI2fMfJ2+8kh96ZunhvZLJ8k+Tuocjk++BygXL56QM5WEidcLgA5
ToUjua7tmSuUA++PHSpPwu2mtxHqpqyu26SOpG9GcX4P3O5IuBaq+Ile7SXIK7lz
csddACiPfHQcfs/65z7/t/Aivpb6maC0CvhtEzD9iTZGkRahCUAfQOCYB+ARnp6+
T6pAF8RlxBqZRnpnCjwsyCp+LBEUK4TP6/PCbHR6lDS781KaXIdL5ZeudZScaLeW
bjamxBnmX8YPDXNafBMNk00JLLtgIBQKfrhejgYc9ql0YaaY+vTl8uooCGwuSoGD
h+6gR2vdjVZ+WVHpxGOPrjXE+JAzVguUxurTzs3Urs+JHFe6Q8T24RBlUYGuzTqA
zNvBuzt7gJxnC+/v11Qchw5XV0dwRQU8ehoJeZWUvBNyP+rSwxfwjftd3JYEQ9Tk
ZRBt5/vz8VOkAKuVKpewZaptIKnXvl63P902MXVgUaeBOGiOEUnkmQFPKMtHNIIn
zq7faKzUeqJjGBlMX87UUztVlYXvNvidFZgMIU0E+ZrhPqJR7C0RaolLf6qqFx3V
ej9Bi7U+DHm2InOh1GW2wGwc7fHN5AwhOFTdNrNCUUhjj4VctBNDJGBKCgYwMLkG
A/A/RCQaB1PariWEMt4Vt4NW/8Fv4AwySxAMIPkLE7t5Llf+d2Gbvm/ak7LD31U3
6aGXviHCZJZPcsvZihy1KaFa7nUwlQErzmRRlxzxkWYpeWB9MpVdK8GTru9EpVO6
unLUzAG+tu6XePMbsweI0hFjNtnf3txsiaX/kb322mseitUxZpZvzePayJIFjas1
iQDKUDWOAdbgo/FELoHsF2eiCHpeGySUGirVclbJVNmJsQY6mxHMnuiyZD7MzZZI
lTCugbsO+m7I/ADhBMvFFbx7XBeBlVIdQGeqexq83neXcwkOaFE+zvoTR9jr6yY2
Ls4KGTEPAzpaK6KanoS+I1Nv1gykuLuM+rpq5aWaO5kQ1OABLYokKsRQ5aILF/KU
+Cdlm2wPK2xYgh3AJzrdYXlp8Sja5mA64Jfgp1Syyq383pst3RygDDTbnAi6gHdw
PYksR8ZqXL40LNBIOlgkVuJupqb00kp0nJoei9KhawfbCQLGPJXoUSKM0WUcBUrf
jhlmqwtvEV5q4JaT6SJV5pFhTPn0ZWjvPDUfJKDzeFDXkAo49hmSFAP/1Z4QN5bK
PX3NcVj4tSRl1YSGX+49LEI79JKM3s12GUQrS2zgkTS75yErIscqYzTQ3slVAGwa
t2vLq/mkWQ6bOixv/DPnxPhoghip2zPb/4oi9XYNSsJ/6CWOdj6H+J+rhOCRUPp3
sDybVgSlb2W1P0O73b9n5LI0/w7uaentcXk5NyOFKGIvZvV1hyQkYxR4Jidrrnjt
tnsUjujzfOnILnARCRBdhGK0dWsOzrH3DW2oHXbo1HbNvMiRcgjetP8YLtXaVzVU
sYYgU3WJ3Mic3k9vO/9UdnwHYvFHzQ3jwixIeMZZJCQSIJAgV5ii1oy8S03h0Ryg
a1kEgxol5tNpt2nfci2c6PVKtD92sFkeY8RL9w/D2KgYhdwtmfDBrieQ+WZzTtom
6gKv46jlcQr8CVg6jZ8Rm/LHSYNwTHk1+H73MMSp1OHRdZqBIT/ZPwd/PqAadiLT
O0/mHj3Z/Fsowdq+CjTwXCPkVhm0NcFV5Mj0JTFZYE+hBofHDBT3t+p2OaApnljR
Pq5F+uJ2Eb5cIv7Kgc4PGl3Jyz8o/bWZQU/AG2HJ2VcTpUEAMRfKvLOTc+90yL8J
JSTvZoNr2J8J7wDLP+VSC8hy1rK/muFjdFwtowrZrdcj0mDZjRluw64xC8HerzZK
yVlyzIiavTRbMoH/I3ZNS2NqK93gfZC/TKYRuo0PgPhxYXlunHQp8s9mPKVKy+m3
RD0rXJ7OFo6RF/MdQN/K8456/W2QVkmI7/kMfHN6E4IWrUIUX14fPs2fZlhlkuSx
rsMG0W1d6bkZXRYVY8wenFomdDZwTGdbT4GOVTJpG1jyrXgyyAakR4Zt4fWNfH2j
ItdMIS39tj5pFqP3rBQXz2QqprJcpkHlOkavfbNY3vexLrnfPQjv5LvNo7AVTWqc
OMDy8mQNQrNn4FlSrgi2TuDLVHPMVy9Jv/W4J2ASG2syCsFd/NJf2k35lyO3fmIJ
qtw7zQmiBlrwLv6ridNvPa6S6LkGQLuropfTW8R7CvRU4IK1NcVLKtaf/O7Yzz5n
cKeYVH+jsSOkha1N92C6NXthQ/XkrvomJxaZ/RGfGKbOZXCDYrVXlKvUSZQf1fMb
JQ3RKbNfLy1B13dElm2O3cHZWQbB1dDMxdgr6MKmvGpQUyFn0TopwEvaHqsn6IGb
HEyJgsHX1zQ2UNSUQLO+WrQwpSl32JRSuZs4Jf3Cio8Whzm4eOF2QzLma1lYWCdg
cg5n+55AxExBFhJ77Eupjz2DPqXiJkoPw7jl2G/9OFtkQ3ZaDF8F8uDL1LvZW7ZW
796TmRVhP9Kqt+26EGCcEKP5qZKyTIU1IKvnbFQDi9EDd8o0Ll5izItev823WcnI
jEjThkfU08z5Es+hNu51WO55DmvUz7jaVLR7usjU6EasA3wdoojHerINCUA2I7Ac
y5rSoa0mjyZOrJTEon0Jr8EWzwr4O6q7td6e/wEfCzZDJ+T64mL1x6gLFtOvIoYo
x6xaN06zpdFEjSkkgu+bS4pnVU8/TfM2kDlfePq/gyvHyNcJusDSmzYWEtNk1GH+
yHUaG/DRHrZLWGHg087N2h6HQ1UAg5m6C0HMfXGZAEwt7Xpc1jt1G11QjljvsgMY
lP+4nNPurRemRW+40mS6785oPcP2bVCONzKo5YVC46SYnfszRI3Ne5uH1VhaikuV
m+RrIfLdnb/7ERFTBzIsFgZMG2lUVaKzWr2+mjvkjTqpXhVwUPTicBrm0qitmefx
OXFx4HzI/TA68KjxvhqKLdd/BjfBLAEsV9SUa2Uy2pBkBGVtOaM6qhsgDS13oIcJ
SYV9/v1S4VTA3Ieo/exp0ov1gKmoVZrQH84TJsUPQpLO758+FXwUqquu7pj4Q5Sf
0Vn23Wusg1sYkglG2y021xz6QIAWX+HsrK1fYtrY4FV8CEfyDBQOb4q04iqGLQUn
38bWTMFo3kf1sOrE8ndU/5uQuJ7cH58KgpkdKSTbEfYKywqRAsevGf+2js9Pqwab
cEkh/9GpFZXkmLH43UovKGm6PAz2LVpqlz+DPM0G8Yvy3qZuAtveSM1pHVOB+a0f
dSceZPQ26XbszQGEqHcFGF3kyimWfPriNbou6jA9Fj41gnFNNvD8xdAYw7YHH1Yg
PAg4RH12Es5BgaHXIgg1m65lKvLDrJ8CXJi6FGlPeVPdTYht02VQVw7m/6EwtUGv
uvOcBVM94HwqMTt3SYZk2oMq+39TyK0PE/b5L+qSvuamxK0MJW3SmH3ZXBTMloey
X2a+7RBHafSuBg5lkRAQUvlNddCCVYqOzR8OTxiF3ITjlcxbHbn9WWgJolXwpsII
7e9ZiDCpQryOQY9WPmS/Fm3dNqMwKBDsnhgUl5p9FRfo8eRkTW+cnR3cjwDphUC5
hgcZuHrbFkGFtIooDoxIOu6WEhyIZm17sLLUbE4NjxR9RELysOEt0gNxSCksY+N9
tqTpaDF8d3TdSkDvg/86eQTeZOgRa8cDE8KIXZqbopo9TbDYweoxKwgA+3a+4m+7
FmbTUSbgYjNmfbDyVV4HrxhpmFffLc3MbV7tqGISYhzDr5QTdxmNQQ23R9R/akgp
gaA90k8sKKJdDphZNKVaXDFrcXA8vR8O7LC32gfcX4GhSnPBB5okEhfVy77ShJRe
hbymwBGvO2QPU9wXPZUv/ept6t4o/JKpFxifgttJskOQQugn+HvF1F5G4je9Az/Z
mGJ5edVqQsz+cJJWmLIvyUntFDbfZvZhG3+18wFY+HPfifLu1Hzo3wgEKKHH0zzp
vMs1RsdS8fcHQrSrmFHIOXS5AoCH65xwEgQiTioADga1VgcmtHhJ3qnt+FYHCgx/
x+uQhHfZJ/89xpxBcldB2+bmi7BD9u1w+UoS4/i8tE9VenE4PbnBEFhRRqq0AFuE
rBAaXnb6e4QSh1oI0OuFYycGKiBBUkmgNXfjat20lGAhCmGUTPXdFL7rsR5BVsPQ
8ukJH7gDW8d/uG7G4Gfp0QNpNnPa8le6DrNFCXQgg+lTPJUD53tx9VzB+2W80xdp
umMcQ3mpPaEFwTAFGTCBIl1lwDKdfGQG56ezK+N23ROFkv5w/mNMbNHZWvzrUsPg
s3Icnv11pZNV61sadMsqSKi7AQjt79oApoG2DFSCtKKNretYSor9/ZEQ4ix+WP/C
me6/DXMzE9OlnTj37RtRRluJy23SH6JQSZPshZBB4Hcr5IVix6VH7o3NyBIjuipR
sgddjwBDnHBgWvWTP5rrxzR7hBh1mVPbWAWemNtGvfkiu8mtz365TUFR5r2LjDDh
f4yu6tFEFUkTBs5iyAEloNJoisK5YnHzpDYF0pJxIphhaq8LOEor+4CXaICE6otv
kv4hfJb7OuAQovdNBxHuZ3/26W9sU0wzzly6izb/cq1LdWGL2kzyY8HTwn0/EJFy
BCvC4dyLU/4Lgz6C4maA1gkYfDiihyrbwrd2lOU3BQBvZNTywXCiUY5QLyw2Sg7N
/yuNOtOhvOZ8zfDzo3Q5o3b87qS/hI7kg5UtXX6dLoKf3M/cdDQlDH6cO1SfAhV5
BJncnKvuQUbeJjDKZc1y8XLkrMkrR1br1ZI6IZe1DW4Uya6qJePuzL4iyhJSmMSd
Y/vexPShFFDPj8jhwtMUDaskfKJ//Ys16jmtGNODrAkP+yumkL30LEIgY9GSBugW
5kZYI/Rl424OU4Q8Q6Yg/pJf700BSk4s8U/KXszUSMYrjiDYWJZmN5EqXCZtrLVK
UPyNLNt/rAjWSl8wPvHd4Pqt/b9g22OrVYHb5535LTBOl0UpvuxPVUcsMcyP9mrN
mhiE8jdLQEOzfJQJJKcs/fSk+ZHrIh6mWOR3hNmd8O+eueTlnm8H+vjYC69pQSH8
mAjp+jhALlL60JqnEvUsbmgQD7KozoKpzcTCX7BY0Ujm6PR3iZl7SmEg5/+MNXXe
I5zxVC75+GPr8xEbsH7Dy9VDGo4PnEYqOryeqpZp7fpK4yXRDC5bkmiaXz9ChFcE
ClXu6d6a+9RgnckL1uFXlHtAOdGD44XSv/vbStDB2gO0i8ByI+ZD6F1TQVn1Hb+X
gIuiIfwkba+75KEOORdJwArhMHFrqICH5S9ApdZvei6cO8AGzWlmcGVs6VKWWjpO
vaq57RUxt2qgjRnGXrsc9OU/VehKymTflUz9FkF6Wsass5V1gSXkPqFgfeVORzSn
de2Uj3fFwoxCEH63KkEeOjmYtOSvmLvwa8nWALl6VT/9MvVQl02HzZGsU6ntIYjk
ITbMnP6MNRn4ieYfW/7c3h/u+A/Ozw1LI2IMTV1A8hur6BNXo9ed4eTdt/9ntUcP
jqeQ/V/8Kg97qTL8eFD4ld9F0Xoag/2t0NxV2j4xEkZWwHrUySVKvEXGiITlQgHY
kylMDKcUul/Q04Ivw/dx16I3Wc5K85ohS+PzDMt30aqVzgxexIA2SBHBxfNHDsCX
22eyW1B/Dp16zGr0QdW4v7b23Ub+TsRPvHNtK/6Q0PhG72fA4JbiFvkywzP2YMC0
a1CS5tul3on2eJ55MhXvqnRkx8Hfps9IXsp2sUuvIs2Y83mW44AR8D86MnzM5DCy
iOvlCjR6ZGdh77sNeqdYcZBjT2iP/5nRgIOFbSHp3op4zlRIGQ7k+hO+vSqXn4Hb
P9gM6cnjEr789swXCwA4I2wdnrAOON4FxCykTwp5Vn800jw105wzPAQcGbk2Tb5M
PAgj3AxO16iCZzgGjf0L9LtdPhN0qEQu4LkXofIY+A/UcumoW21qgDMZKeMZZJFL
OsrSqD3qngnPRHfJGx+hDVvG+P6SQtu6eDeh2M8ZMmMWHxZrm7WQDAYtGU9D9aDT
WISFGu/w8+bB0smSVKsO0r6OQ8xrRZjMCHN2ks26sjaAWp7iiwO9H9WLxdzuAOWX
79QChMW0W7/qUNgAbL8Rm7ducVQvqT/hbrjNWSnyr2oXLPq5GVws0YBixTbKBw8P
xeyjn0lnaWMmaybfmd+KoM9cDvUztHDT5mXnxUG8IBJSeHrw4D2sLr7k4XfwmSCS
rNYytygSo3EhneGpmcskMZwiNbqve/Q6TT9bk7uX7NZmaDcVkdVEOyNJvIKnsp5W
Apxg8izc/Co5wnE4NdzkUGx8ci+X3nfmQMzoalggZw2I4+QoLuC3ar9TdGAEZmR7
s5Fo3C2jEwKPSESK+xyjCs/dNBdqWw3ePZiTp23CZNa2Jp7BH9J4ATMfCFT+H58g
rn7M41wH9SsVAI7xjPw7DNlzoA8REvaraDA+xeh+AZIEkQsGY68e//equfVHH4QE
STuVJeVp8mL3rDH/DUYTAR6SxAWwxxSjtYZgQH2rFTCK3ZmMqocxLLn9LcMg3y+N
GAWppGGVuwTdH67nsWcFMrntNtiUQ6znfNsWbtAIw2kpx5hfGcfMjGpl89kUz99H
JiPLZ1rzsgMhWYgG1i0lW3SY9W16FnurGlxqnOqn11Pbb7f31FtTOQG93nGhEL+m
FH96Kj2RUkqYueC95N5Nc67DWaiDrj4pMzg4OGeIfaWJgu8lhjRCH22R/Zzn3/gT
k0dc/Ux8vrjA3Q9pD0CUm8AaeQ1H3tHMjpNPg210LplYWU9r2Gb1iPm5/SEyoM/H
b797xbO49rjb+1M0/8km5Z4Hmcsdm2RdEKGXwlRbpFeTY9gJaYIeDEEa+O99W4sT
xSl1KaN7WZjLzjQ00gjKJmQHGEfmYVaNZXeNHzMQxwZ38YxTtzjpWDx98wjW4qaR
shwgGYMYl6aRMOBRQew4l430l6GoPid4mU1PEvACMGk+CHwxIyi7NZO4+MJ+qz4L
EP8ocb0dqV2IW5UhtOS+I4nUQl77Mrc+tdGv/L8heG8wLZgXMNUoVD9VKti8X0Oo
Np9ZSdq/PkwoNw+p31IWopu5u7KTaxqSiZ+OHDcB3qZ35Zsyyui9OBDZf8+UeraG
CYEv3vRSkG683uGuFIiNqp04Dsew9z34L8UZB5/igPcehk0mkI4LzicXj9z8EpJC
sbwvvFk43sQ9UYOKKWnTfSsL+mfEyX003fY5nmuH5dk8yGmldAoKmA0pfxRK4PEt
LyxH8bxZ1WVf/1NOZItHBHx1g2JVn1a1BHRZH0zac17RVvVg7M4lp6cEHNwDAbEC
IsDpJ0v2OnC0neW8wmMJ6m4sbfjXOIe+OnBJF+lm9xVScWl28eUHOLjgaC1brSIE
2njI7VXjCQ6PpXbAZWkbZfi8PM3zLxAt/kj+BkkHejr6D5tZYSBvl8DVVe+E2rjP
oq53vSRgOIdqMwO9XUkWG3ynA9SPX4glGO7NMymJ2UJaEyaZ7k1ZbLiXfafk59UD
u7xQ5H5aEE6HH0cCw9i0+g96CjxlQcEqDWuV9DFH+X1WnULkyMnx5hRs4+/i6X2d
5dvlghxyXmHbaZW6WnkuJEHAsLa3ClFirsfK5wKDO5//IWqj9OT/1gEt0x1he+KH
Xmfw1IZQM1KGT5It6J8LZonwH9wDStv4JyH3Zm+n/FyUuHw9oPuvSUKtTSxbkDFl
Fu0PR2VzU4/AX1F0qNHUO6eebx02LJ3VjF6CNQUNov/2dZ5JJzZUw4I3SpUWgbxp
4wr+IIjojGNXgGXkclJ6QfPRkGF6C/XIEm0HqYlKP/5b4/dybvGsak2LG2HSziMI
J3vVp1FZyWsN7abKujZrOYWbRhU6e5m1nb5EwU3a6nfAXkHiCuP2+EW+ZuE2bp4r
S6GwqlldgVxC+sKrEVobJitrFF6WOTLe7z6C1+HR8jMo2d8QyPakNbci2F0iKKzw
wozWPA8W+6mB81s6DOk4qUoAAQxJvWD/AYnPCqkW+GkNCB4ouvWbwUkeIAoEopvh
tg2263t6GotlrR/lm5pJL/YMbHG0ss49H95Nd4kVgsq7+1xhQL5BkF/+CPLJPPJY
ZOQ3mR0pP+bQev1+nLgKEjvfUFdItPVK3VMqhVkxNtGVFTfDaZ6c1SyzzaBxAGC2
LbvPaVh9DOwEOIYi2ErXwvtZckHOQtUdd0A3tORkDD7eRPgAI51l6GdsYEt5PU+5
wzSUv7h4Lp8KqJP1ueh8JzV1WDYWJDiMKkmGfVXbD3VKvBhU2c3K2CsEWFez1ZfX
nI/HYT47RHCpdHA3BqAXWVlZUsaVKLIM3XTzuiWB1tO8b09xhGpB/hFQYglS+1Hf
nc5/j2I/LfvVImE02liEH8LrCvnJ+at6QQIg+FYrZcX9KTdldRdE9lK7oI8zXyVO
ED5XrsB+833tB29aSggDQkdu/Qca8so3iOX5Hj5gS7z52FEL7IN2otX3sP5BF7bz
/+vUgfDpjcqcXbJVCLyAxa81/xg0hTE4yR0+GMIyvLXGuB5ouaMY0OiZLeMnf/Ez
+Ya+DgvDzYjBD7cWS4NeLiyxHdqejkSWOQqERe9qTjxmpVk8NTd3zHRrlUSCReHa
Wj0c0/9bzfUxwKWFu8G9ITdpD60tDJDCi25Fu71G4+jSCdQCYlL3RQ8Dj+zxeEGC
FcdNanG0Ttrz6EfesPRGIvC5C9OmK++tlo/WzqLF3g2uTUCHzoZkbGIXV65n0jUW
jDOZ6hDIrgRs9avj9pHVTHZ/r9EC41e4TqoRx4TJgXR4PGR42x5wYpsc40EjmnbF
GOqwiWpvH9aewrAVv9T0W6lsvyDCP1M7a3wv0ervOwc28gm8ccSUyY7l4Kedm08W
Mq/ps7MwRraFEmrc8OM6dVxy5UR/QImnHSjPerLuYI4iwjizEicHe8VM2BCljXr8
OUvfNMlLjCqYx2J4zf81Yl2ekm9W65hwdXbLlXep8ZMlLKx03cjI8wZUvfOsqt2p
sk0Jvk2u4AvygDASwvbYP09AgwfLZbnxvuwiMGUC5ijOhmW/iLoJIvuWMLUHmrWI
M8ckx60kQcqmsmQEjXbp3F0e2NGxDHS5nt3gJODWGqb9+/IwRmxFMTDEjx9BU/5s
3YYHUGO+cQ9eJ5U7SzN9ML4kDltmaxpFHgqRrULNFguHmNlovxEJ5gsl4F6eeWTc
qOwJPkXIkTHettgEp7O329XjyDOEh5DVr9wrpDzza/6csKviy5m36g5YfSQ3EHai
3rji9qlA313vcTDby1Suzcm5VLIu8pulcgFM7Q3mSOqhsXLetTCC6/3cr7oGO4GG
/hBLmFA4DehapShZnGR5GVvgeThKruf5KdkWDZjrccZnrJbMJvXvwL/roIF6HCqZ
8BiothEVvvh8kSMZNeKOr6klNrxlS4e7vNjClheFx2khzG1N5QfvWvHni+ZFuSga
F6tjTPr5Y7UqkBG2yPbOKc8rdMOkm5rjTvLHNQbAl0tFKvNdHMSE1KLCOheK5XsX
Pwkk6XBQVB0uNsW23NhdNVWmrpDs+uB3+OGWzJ4AbG5ir1O4kgpMWkHEBpOJkUU/
710QSOUfsb6eFNL3MeqjmzQOzBrSz93Sv+SIeEb5/z63mXNItPvULJ5i+/saNsdy
SSkrFgfy0ssmLbWyFCcdPBnjxjT71zJpYZ4rVGk+fgLf3R0bAP7euMk//A8/QMhH
zSnBJw1hYc228/FjeCafbQdtN/zU45WiW6VxJrGxkH4XXvcmPZ9cEk93XyKt1iKO
sI6Z2QdCKrK6XR4CynJbhbQ069KCOsLaXfnVg5ZKotBtlFfkXBv397oqiefAFRVz
wzQi+JWlEEC8hh6aLUXkTU7/c5yzBoQM0VzRud4kjMCfNzh2P5YA2cgeXUtCRW3a
wSSHVAw73X0TJke/Rq+/GlCxvhwrTYZwEGzTSSj0MWE5GYXTtHvyt53EAzlyWywC
WUNA6YDwJej2lCS+XlhsHBJ/X/QD9OJZKmIgx5nwRLYn6Apg0t5YPnq5on7yntfK
W3aSjPOhiAdHl75R2nvgmbHKLcOZYLjSSciKYU2RMUnceGieWEQkKvzAMopNr/QQ
deOJ7pezdubS3Ka35Z6fe3BV+Z+dcip+sakRMpMB0K8Hb+ijneuyApLTgt6XwWY4
kLONSXcQfc2XFx6hOH4GvuaNMqy5rSOKq5ILs/Wzz9cM3i1f+hfF9N2nP2QBqYx/
m+dN+oTzaaypWVIEQguMn0jbEsR3QdyHXsF7b+rQrASYY9OICvrpjo1h+F10AJ1m
fnz8xuR5c4740mstSMAV0E/0aHHBVZFyNUM++Gwb5ynO58bXGVqeiTE0bk/rRtHz
OGzcUofhzlVI/EFZXhMasslmRUkBxfE8HVUy0YDzOtrNdkh5gYjtPHHwYOt+YFjJ
+hQ16wJ6YUXazDRgQA8pXKG1Ke3DJb0F1hZm/EnGyEISTTdl4W4s8eBbMR9oHAdw
ICEuFxxgivxm23+gZhQR8ppTTmhnJb70jEGWB/dyXpVmGzMtpjnEYv+Yzifxie7g
CWSaQJ93xZvtI68NlciiEIgIwBuXT1P0x6iN7vD06mD6yk7iquC2UEf7Cv6uB92Q
JWYjGekCquI4BF54uqiP8ogVIOWuegrJP7nLS0q3Tij+4FIPi5YpRmBEFeNeI5DY
+Xsb4BgdqqcuJJye70Jjvf8c9O8c3RGMYtg7hi0GLWn6w8xkIh8sOzvtnXKUle8r
r6gzE7dZtZ3nmhqKTDrHYtm5GCIH3ryVFgKApoEX1PTT/8TNm92WZmEX9acsG+Q4
g4PRdQTsX3Y9Ur/9M0re3tLzUFVWeP8YSRNjYolTqCBbgjHG9Ns5dXZqSgMuy5bk
E6R1WA31hdTtovo56TG03bH9/AeUS0ZY0VdJ/Fi7GDAMR9aPZax0r4JzLCPCbYtY
/e32IP8yO0Put083Pt4HTsRXMFSAUrnPrsqfTL7+wADgzijUiUHSQnUze64Ur34J
zxrHOLdEVitdSWoxqdf0y9r/+ZQV8UFilDaH+/W81Yb5KuMsxEOdc5Ys8oh4jWbS
vInfTEDnePOYmqgZk/e4XkLG0wD+A4pcKTYRt2Jd/Udu4tUzrlAdul/5EmPt9vpb
hnPCogJehuhPKz5tyFNLy1w4iQyjSGcN9ot4Kfq4KhLsSsjsp7oBzXu+y3e1jxYl
p2ub8VbnI3Ykp9uJ/fMxFYGcJve+1Kmyh2Q2lJwc4ENGbBMtIRcOPqgomTV7T7I7
cFZQtsfbq1wUe7A1nL7/EkgEPKoFk5KaG1Vb+f18k9NX0n6jHEIA6wXBk7WbO0dc
1kbvh7G4zJv6pHqUqUvL/4nhH6tItLDsX9d0L/VJS21xdTlD0bpusF1ZvPYTsKaT
m5Kpi9fXHKupJDIllsUwCnVvpeIqjTxVu3hT/OwxB87S9aMHzbQWCuwhIpvlLgFq
RKKJwen8wD86GUN2MoJmPVJXmC4+Z8AonkgWARrMh0QIfTLpiAiZAt6XMN4sHi2f
Eh3iN/9ZxEdSOa0ac3MN8mCfs/fN76+MDCCBOx+gM/ynTjqWIcWzZ1wihGNKywch
GnpRDefb1kfZL0SMPp9zBk6WA9BqamGwV9fC2dRFPoRd5J3F+LBCSXf02fU0rv1J
J8l8MEf39/RmNb6FNPDwri/DyzdH/sAdSEhN5TJkwXuAX3PJfIEJJe/1XD2+eN26
7dwbOh4MtVu9e5oVAET1e1CtAypxjrYg90sD6Zb8yQvIJ/8pHQP8cRourBJOor3u
kfQpnPJpWrLW5DArCCIPn7T4hOjtD5Y3YZCKvQCTz5rTKhDXDCFXuoNPxFqNISh2
EP6Z/7tLvL+Tg3hZXZlgekIjXHO9+zs8a8opI7iGDzs/YGAXl2TcVuPRWkCIDdvb
EImAJOlVJPq+USxDllvLNTXHLNXum+sNdwp8PWremc+MMgOrZjJQXsaZxhJ86WmN
OkrGiNX/xaqG1g8IE2+CtHyhoAB0xEa1ckOaRsKM/5PPYeUEuCl4yKp06drSwq6u
mThlNNkNZW0x7xGntfYTCyBQttZBOBU4OGlhaWg1DI3djQUrVzHyOquaRg4iurDG
pNZgJUhP1FQ5miRckhxRNj+hwCrBMNzXPSE838JsBt12AYSIxpD2I7KtMhAacjd8
WF2cJq0yj6rzpqY/zeDms50DIGKdOLm6oLPBDjZ+CyLly0+XXNo65JAa45OZ90N1
60YReusfAHmZbSmOURHthFwfRogumZ/7AH96x5KnaqwrEoZRx0I9Ix2j/H/CUJSr
b7ohOh7x8K4ht9WCYcbMjZ+aox7cHL1me4YyZ7pOIUXo2Tkix20Mo6NPxIh2m/ng
MghnAtvFF4HAED1VGphuH53E77oXMeVSwPLcborfZokx0Om/ntpGBAeFx4kR8YI+
3JXcOCKd7Em8hxRxBRr8HWqJ3JUrWGlhLuxfRilYoInhSe6/foXhsCgF//HsrhSr
PpuWLG7ujWGPvqH0FIXRuwLF2K81u7WBJq7Kt4elfo/Wh+PQtUv/rwpjfTibo+6u
6DYLdGOmBTtz5Ga6zmeGox1nz27sIoLpcP15y6Grxj1a46f2DLhCfjG64gM3QXeQ
P0kWGuzxHolf3KuHJGbi6PCa3AE2gQVcmnETDfzH5Jt72FrBK31c1/hrh8MSPrk0
pw6fEi2CneWwzdyHHk7Nz+8zA0499uemkjRoWlXV/MAEHkD1Aq2nuljk0KS8UHke
2alEeILrTSz98cYRKvodRfAsSdIF+0zkeDjgiLvL58wdIaj0C/NY1CmrfgFispnU
rUE7R8EU3xaxKAxQd9ZjHvAMuQhZ0q57xzoJuxfhzlSo3lhSGYc9U9HOGtAj1PpD
A36/2yhwbbt7VJNz+2rq6cFvxU3bTVFeDh1HIAvix49voBk3dMhMY/MHPEVxlRHl
uPDNGgY8YcCYOPco09E0fZZWpQyj27NbpxcS+T/eC3K2jfVEWgE6UhIAn9Np59OU
v8uimSpY2dMrgzcdE1jj7zqxTHU9T49MkvOpSu1bcUZvIXfFShK4xcrWRRZb+QDO
2XRDs8W76SyaE+gjz7sWocRstvUd7HRc4awcaieSrFriGeHFTTwQ7SSWry+53d8M
hDIFg8uXQcsiYUwFx+Ez6evgmPmF5UIxwlqZUPK6xtldyl/FJede7I014cWEV30K
AyX38wZVzSU5voLBAcQIaQ6TyRm0eSbC8vUoGCXYSSTUmjKhkOCXJSBbS1jnn3Ht
5stu1xbjjb5PJ5udHcFQnjhdGMR8nYZF6nwmp08mzYNvu99NODN+nZFsEXf0IGpB
/VzgIcLe6eunGrb/LuoDbcjjGeNF4XGJ+eD6voULsb2tBsQCFDcSo9TSKFX+ZIB7
z071gReHhOh/MfTeUOjSDP2g7CD/JnLK+dLdvIv2w+Se3ouuIPn0joFNmiKnUNxh
WzZy9V52YiJwswikR0Zr6z7dy2k4mlTJvoUMJxjRDJnqo9onxTeekdET82xC8ydu
wSGEYHbaELwnw19VtI+3dVDq1ShGLLKByM/A/7OcSdZQ+bm3JesUk4oHkT0vvxse
+IuXWrh26/wKYaMZ/YM/RkCter5jCHRYeny8XAMK1fd5glre57ZfJUEgOl/4l5i9
fkYOuV74ZICbvQqcosHFPo+q4JjdvxfMnyyzNa1Jf/dV8jdHG29fUEMu9aTCIEAW
lK4g1/dsK09Jcf+plhGU/1WFKK7oatp+9o0xxF1auy6K8WJNT5B1KIiAh4MFcHf4
2lATEg3EdTkPoRyGZHbl3RI8ekhaShbBj414HSiLE6LEYz2f0BH5pcMy2ndksPl0
bP0di7aE9mgWTPM79KjAKtbseEqygg4b8xDnSjlpZJ6hYwS2H9hKO6Ezn+n74jfe
A7SxzAO6SwMQWILRzw+M4reIVJHJmqXbA0YG+un/rmVSQNX8Dfwl/CDxVNI69txb
E9JTkpsxlaQPkbvNqFGlHPLZygNvd+QY1l4SjsTJlRM71/o1iXALdFL10BNi0413
Gn40LSzN5DtH7c+ykr+gx00B61zu+Y30g17LFqCJyhb17d8tEy3+J2BcDmb3STQV
gjP/Pdx0wRRT8lis6pbSQotXZX6MCJKS/TdCE1xq8U1EQplAgQ8ADN+KPRKkvXUf
6UzOemk6sB6nk6lQNf6eokLvqwbwApRjHGf/ISZCd7GPjQEXqTehpOBewEYGKMs+
aQkg3V03UN21ESh20YV0FdN+Tsb5DOj3eam/XJuzIbpspc7sc9XGWgcYYUiVdVOg
BMg1oLBDDXfqkykINSjrCIjDfIpVUKlYzgquWocmLJdmls/+B+JCGUOyY9QoB+Wr
2M3eKnmDW7/+werAHvwXpbw+q6GuLcIR6wV4m63BvFMT8xV1yQlMjOFrE+odWr2j
XJaPuOGqjX6Y0EZfZZOcpQKiPC5v97ghePK9AKeFRspYkFQvr/RG1eQg9t5fEMJX
GOkRmavJnkOxzQsk9ucSQjz9qXnSaQ6ibDiO3mZKSUbtJRXXK1IpLJirwdchl2r6
dCQq+F+QSSMLn5Zc427NTSu+JZYdP3eraTmQHFtKnkp7MOXipn1dfTxjgZYUE9lt
2myH/ZK+R5bt6dCb8A0UJ1yk9KJ3dBXg9pMU6/Hy9HsZ3D0YU7S7OCJjbkfW/EVk
SqGqD63m2a1zxTV/a6nY1BjPi9XbwVoqvR5q7Tn+A66xFCfpRqoMQ/aOkhWK7Jpd
UeyysgyRSSHxLt8Z9XA0W9lxUIMWoi1hOq2512ykucjbO+jjYjsU98EwUu77yjUX
HE/ugTCcXaNUUQJzsORE8VcXYXFEIlk7l9mGhPjUfFWy7esgxbTmPlqYt3eazxfN
akolZoh3zelw/OAYhGXXjM+Jm00M2D9jBmN2SiLIqDF0BAlqnQnePe0o5p8sF5RO
lz4dFmScgtEfR8gh1KOhcxbkYahs+/nrmGIViBDbq/fSN0C99qClxlZ2ZwFZHqTY
fMqlmkh/KPE4Puxq1bv+dLr39A79rSV3Ru6qYliUV4pI1lWASDJ01kIe6wSSO/9J
At7N9H5WN4g6rhUnpJurhQ+V/s/9DHOl84461WtF5D2XqxxCIHyX/FdxkNp8Zjmt
PLiVi0c+hV6UGLlyTSl34SkGpU9weNhp3fGoyRGwRTY8Z3vSRyk+uU31XB93uUmU
NJeDUuC29BxcbMrgr90oSDsmxa1jqz8djrPwgODufOIdnXjj0ybCR8AsKIVcCTSk
YfyMYv+bgrZoPrJD4Wb7FNdeFF8pOqyRZGRWtzSjNHDIodq9nHO14bqE9zSXvfwG
NHWDtodxSd1nBYCsiBZ26z++KSpALBcYzyBwk5xrTshVVt8HBLjwgzxlZ/3GF1p8
PN89lhQGJ/7bRQwZfJ6YhLpmDfB79fJj+j86kPKuzwOGUjZjKo2+7tqqzCV9ZH+S
lu1zb9zD159DbosfzkknMM2gCgYUwau3TchxZTdOFdLJFYE0LLrYrsY6cR9XV5R8
fURJklTd/Wn1uP6IYOXDRC5iTeM+gJGjVjIcOoQLZL+9N57knCMI4+oaLktVjiTt
cULVcDIEQn3w3KpnCU/hdgVuVUd3W11tyKF0E6dv4T98wmNeYOJiG2lV9l4d5/GR
l3SaZXB1QlIo10OIj4Q6L23Ab3E3tRKW2VUmXM9KFF53lyzx10t5dKJKkJSHEvMp
Ne4LI5pycDtiq78pSM93VWJLu0npwTEKCSttJTXnf4v5K0hmYZBhN7dPe/7ftXUP
oW3IhmkmyxYDnAo8NcykNDCjuZ9VNMBbQruGdVmR5mlfjrmaRWtOO9CDI551IdXI
5bmWUVP2f8mZif2ArmNaifognfrj4ijZS9ySIkWOpDSsM28YiN6NyiQyDAfMaI2R
x76dTXz3Ng/ETqW8xE9WzEhKm5AXU45/CzBwzR2CvdZ3HXDSHQIcr2JvHG9/QQbl
zY72yJTdRVv/y9GGJrIVUXPyEMPtdTRNdVxYbls2AIjLbkesA2ysAcYOkq/Gb9YO
U4MjDIo5giTw+IJADmr9VbbnwhrQvhpj33jFJtIw4UiiK1ADqbIEiC503AIU4CpC
tm/1mWxYBGemxwvzXI4lqgXLeQXjqjT6zARaPLMdL80hNnPRyCrj0Qc4SWTQyfZq
A3XjNwC4+BDbCAUwhLuAcbegas3CFlshKIuKcwUjZSmesOB8BTKsHLYoaZXDXpxq
8o9rSwvU7ylhWNwqRg23Gr3K3/uVbO6TMJCVTZkJ04HnjJiGw2k4sVQB1SqlVJWp
AKdwtAHnIG/YBJ6u+pdJHTfneRN0bqBL7WiLswh9Yh8jlHgxnShTvJn3hOqgtUh4
+ME7WDBJJpsiGBq5l4xpwuYXV9i8TbjsPSSiMQHeYzIRNJhpT9+XYx63S9nMkssy
tfHu5YPeigrNAip86TSaoqehhfZMDb9Yq3nkSH5qxKsrzY/RX1UsV6168UYXs8zv
mjjZpQd41GUZJh8D5ACsfsBRurzlYFk0qfjiIueS+rsHQWetbKmDs6FymoBxo8oH
lh//sHjU9phxhJ9asRbEKYAmk4szrJ9oYr/hpu5F7EbxXBMcG+J4Jh+spnIdEu3G
DHXZW775pTiwL5yp1fh5NZ3PCdjtJ0dW40bbxhJSC9Flb9obSCJzFiGDzTEyg3WD
WXrebSYlmwiHD8wXyzaiCBqocDtOzJULdAofFIEaW/FiXZ3juXFGYeLmm/YeukBv
FwnT84u7C3jWkln/ZA72T7kGPGEnI966d9KWTQqBfvQYHxap5Tmdsp3evBqFX/bz
42mKqRjNZj2B2dhmGdxldKyY1Xlo+e0XbmDRoqn5yAmowIaLT+/MUjj3AIQyfDyL
dBfreucSjZfUcmgf8xCuL4GZpKQcvP61tZsNKAqzLaH9onqwfTjEaEUCaDBS0vIH
uPoSBlvZDSoAVMmzGR1czQv6VmK5Um36J3Y3cOBziBFoU42cQ1hos7Nz+u/ctAjw
E8ybNFWbV/dNvRCALAjKCT3U9frP5TCGr32tSI+ol45kISVxF5wl7bCUpQs3/o2j
5umxielilUzJV2T4A5T5Fm+qcR6g/4p8foEJRaivP+4b/1r+TLzlQ+spDXLb8mu2
DYLSi5mAD4lJ2jEuNQBPrUFVD7XtnbbyrTz68ZNtYF0WIluUYEkMGITBYeUcdvtw
dAGpsJIDg+9jiggCNtKCkMEROmQPez6t7wj41dQzWzQpRVaKFh4Fd1bI+HuuaRok
BAStoHX0bFy4053YyHW2nwnUKe3FK+oymesIQbK/Re9qG2SQ74xGSHwTQKK9QZVw
l/ggPtF+nl9qkwlj7dzqg++4VE1WsUHgeuLYapKwMUdiDyyV/9R8atYMlJV421xU
BQnUHBIRzy85iZ+uW1WBIILKVJcTrD1JgzxfGHFs/sbQ2gqOIekSJldANZyIjzFg
pMgTcAWb2XPUHie1x0gjTE5/IfRn43nmWQ37Sqs0HA3XFskyxf0Zqo4thTjoaKtg
/YBfAUrnllUelR7g9AzPuZ1LzxjfMgDD//Cg0sH02L0XAH3Jq+QsV9BGpCf3gksz
vaAtaTE7CqpjRj6xOCl+Rhq9DJiWpZCfWVUhDiEWZKXNym8UHOxNoThVkNG7bNOO
M6STrpfQ0aeoIzEHzTqGsSd6ylYvViCsM5dnP8ZF6g/Df3D91WwqQQMS8SngVPkk
7r1PyjGr4VrGgl5EDLxiKHFejd8a9vD4AkLvmuAwV+i7Mg7JhbMqN/M1i5upJig0
xpcGyaDQFtCW2S1rfeskJw/0ozW1MRYgIvj0SZosaKPIeAd6szSL43Q8msLiwjWL
jlIhWZnPNijXB5+THS4wVQ4p2vtkNprQ4suRQJHhcK3tFDbANSnXt62sGKr1a8x8
4NgfHf/X3EPprjwx3+ICXN+LI9PudyKT1MKys+dSpKgPo5evAFrFwqCA0PXeX+Ne
BxFmAz4RKeSv7W3lJ34rAIKwP1gOPfv9jCMMRViL/zM3MmZv2KEiI0ujp+jdR0er
NcJTXXjL5J1Bs/yQH511cnWN5ogpf2WwXykWLKf9Ug2xD+j2JwOllzjYkOf0/F9L
y/2XE/fJUQBofAITHgnAQJGtFNzWTRlmak3tu6cyCsfFeBjw5GtEmG1LAK6tXmbv
0uIQb6t6vZyPxG8Wgq7+aTqkiycyPLOd3AJvnc5Gc4rbt8B2+aBgvSfouxMSn12K
Nvb/WX08HBNwGdzwHzYj4eMNuS6tX+NGyN/bogJLqK4XUZfN6OO4JhU2XYprp2HA
eOhPNTR8n7xoSdkBgkCT+BFPlrp3A0nlT7QVonIUId+nq2KAks4i6NFWNrZ6UxOc
KcPB2ZkLVwiYfQy5mJOIDnp+bNk/vomi7b1YIk4g69PK8huaajYeD7XBOQ0MSMqE
op2rTD2XxFTx5OEFIF4F1T8a/KzrwkedGbrR3DrCHS1juwV5IRv/ykD9wKlSP++Q
HeD3LVF8QOHaWxP7TEdIoK/p6syguBLpYwN6JCnoyyGh0HvnAil1A62xASq6dTSb
hFd7g3AP/mgybpygFQqio6+35/rfr5rIVahO5SluV0OeIYrk56kdbezeJ1k3ijys
ouxzTWuBLzURWvOUvLUCll4g6nmYNRpg1fP0Es77JL5QuFEmhoEjMbBEqPwUu9vo
Z1+U8pdXQNkuMSpG0J56NjoGK+8gc8i4RNIxQ/FlqinhgvszXzWn6c3Il3FbL5RP
3N+emyhx4SIrHezKt9mgo/ebXQCajy/EMiw0Xc9lIhQJUpI5aHgKhjMdciZ9HmSW
2b+19upMr0f1VJ7NdNXAYtnXy5wUfRbiO5NB2iAy0LZW6C3ESeAGUKXLpI/0GHq8
fiKpYhl3T4Pn8qbDwuQXHoFnpleRi4cp7GQjsmLYCUI24AbCtGmUxFE2gloukZpt
lyz1yqbzbRZkcRR9xVLlDVt8HuP9Qem5X/AwgB/rqMVPLhlt4Alou41Jw9ZfbZ0X
fwM5T/hH23u/x6OEtuJEiBaRhfq8prtAueYxY0PcDkWpoxWC4RzBb6AorDnji9d9
3lekJRHwLFukMTpIkYnm/lGu8iQhvP02jgSsUfB4ZYy3tFJbYnW9iHInrj25FfSg
e293/CVnW500KJsb5hoaphLaHl8PpFbFydue4zv8jU1bNW+3in/TpYuKF7W/hRoE
L5g02nfxvOkRHPn5lQZHlZowBa3J/iDY17Gc57J9+QjWtwV9Lg7YJECfTK+SOnko
5esSOLihLDw3OrBNs9uh8wDY4GN2qU1/UFpx/X4qIb56rADST0EXgiBng+NmZOSN
WCYGAqii08QEBGcfzREwqSWx4tSJcflk4OQZ4TTQ5UX/H0muVjsbpAIztvrNx7uM
0fvjFp9DOk0+kWHTNcVTrRoQE4/DgnIOGL8KxdSQZCZPaK9c+BS2vrqiOPw6daqC
BgNgmmjaz0f4c+fqOjwqVsFlWUHjSgcBPE2cQwGbqrCI2EXWn0Y3q1qMqsEFIs1H
oJEKcTe+R0tIJjh0QO2RfmOLN+q9b7C/9+SXC9aSTySouRUoQV5Lx87fIMYC8HPy
x7XleAS1xbD1+NLfvD2/EFVUPuVZK1TvZbr1NlNKmjwqgwZhSCYDzJAvbMpDgt4J
q2xBoYClHYW1piQdYFPcAwJklVNv1F2Wo3JxUMquTOQDG1b8BuBEaj6V+QIBzdKC
TySGU6lVYxgGCTKKrSocz1qqLQMfpOJgOBwlTrchzecCL2NYdwARNes9q2q/IB18
Aku9fNvOB0UaK54zDficJQ4vTQ3zln4/+Zl7mhusH9P96kQWwp9niHtqoCbCdVTm
wuX5Cz2wfG6XDigg3a3vtUOWaX3UoEDyb6ESAbQXkLCAVIALg5RDHyh/u3qCE/ZY
Qar7oDxEzvN0p0FsHTYRVl8KvZBgUJR5g5bN7S5LOJElds3bqxZTsdqvYouJuE+X
wdpCKhbi1wYeFRqK8fPQM/kPyYJhSlOnjP8Em+NcC/oIOJ1EuouwkizI5Xc6StMQ
PK7CR9nHHZeiq8gt2s7ay4crkajimvYv9uWCMdDOuWVULsNfDg4nEUnWUwwxN5CJ
ZT08NTevnCKLxwo6So+xzDIAYLrWzGwtasgD0Iau1yala9VTdll7GwM/d9e4KBxr
ANtyWKSM479GU+3K6Yw7dXy9c+Ne0l6gPepkbjyO5JrF1ExkrZPU8ETQoYh3/FfC
Lu+zBpvTw9llZSIimkDuJ7uX5Tbb7W0e6UfQ1rGB/qtD4b74fgTpS8+HHnL/kPQi
M8/vtYFai4jl+NPxMQL1OZh6aerseuRH1Uc+eI1KcYnDooeneEpSYLhEEob56UHB
jwxQSo6z0N9GDeLe8f6Pfwpw9Ax5hd9mk/gOYwS5LxnH+CnKf7mwP/P5kS5jvZwC
sN6/oE1JEXpzLylmpum2J93RzbL8vN3TrUqPHaIu9Vbptn2IQOvrSKym20HjEChv
M1S5uHtmmOQhc4mtHKJII4usJm29DvNRcA9MR8Cwl4pfuYiCR79CPzDOVz2O6wsO
I9AUxcoLOi29iSo2m+//xXsEk07NjxwjGnGJWjQyjA8lrNUbCs0ZNkBi0/1GAJ4v
AKhRv238dO3KQG4y29dCscnECwyHEa4Uf+dTPnILUP4oQ1yfjX5Zztfy3BTYX5UJ
IIG8raj9ORNIeqw/GPbhliyYkHn/vtvc+2PFQPx+bTv/+8I4E1ToNGmawq04wWIn
LQGMvevB4YYHIrZiLt66H0+dJGk+gb8FQX/Pcp/bqXIyj75GI2fS8D9dvkOlC3mq
6l5QGBOgCHqp5eMIcSdkb3Kopduh+k1xB8ILN02azjdr7zhyEMDoUrTr2jcwiGl3
ks4atRvm+YZtvfOa+DEaaOcqhhfhR3vs37cE/SjlOS6Pd8GUx5fENw+aIh6bX+ef
3M8LfILhlmxrDNrQAhkqG/pp7aYLDmoZL5EhuWVS55IijQFmjafS5DWZKjhNJFJN
MdVLJKBfUsuKtKlodSvUjcXiWa9YQOvA/mp8QeU85CFon8m1yEt5ERo8dD4F52w0
92yVivIp2/r1YLBy7PmbfSvoLJTIEqeN33F7QAY4mTSCVxlFfy04Bt58TbXlFnM6
YdSlFqERmJX/dKmX+j/ZuwKPXJhYewvm5YNgfA40TtRL07PYLE8hMlhpLAMshsPS
JB5hT+jTKW+yPRC9QbMp3tKVrCWfAqLijThcC0sBHgoeI1SO1B7u+pP8Zfveungj
esp/4Ge0k1qRsMg6RYPERhgwJehw3RhsIV2PAfS1eTahEizfeKL3ZU3kPVw4X1ks
jp2ZQt3F57FloFHmKuw8P6JhwYp8CtXN2m1AmkkjocXllkoda6Y8YtKPeMu2FEY5
7efH88UjTfdLK1oCMv9ko8gLtUcW/3elZmq0fQmL96ZsOVw5zPlr8/QBmKHoEw9E
RQDXQ+q3gfN2qNW+tL4BizyRz0UMedMlXkjjRO69hkOVk2NlF4xKfH1OO2iv9DwD
O4NK4F7aorFXhcBF5DjFVevTe2p9x0tyRq50sXYvaYgIfipbivuDygiyO5xmOY/Y
KCH1D9eMbnjLC7gexlYuJgePotnmwFIXUNopGKaXZXgMDEuGVzHC/69qK63y4AjK
uNwHdc8rCEl9j99EXUt7b++/qlE4mnbPBsD1SacM9yTPPJ0NRYZWrf6Vy/BOgI4J
zkCP5vtz94hfdy8b56D2NEjHleuFC/yobHUo9LxOiVmwO034rA4TFnro4EWMSo8u
4Gf/tJ8lgTli6F8n8YbzvHLq7JV1BgvrL/3OBCsksKdACIS/xYIGQip+cxlka0aa
8b0+YaaKd/ZBg54surirutEkYKJrHDopKAyal57yjCskkNlQoNZ6WXQVDnDVgK/Z
Mf+fduZYnv8kte1L97h0xUSU4KtU3ionULIcexx0Pf5NZyDcwxs8hASKQIqXTlVo
23rL/SFrHcZEPDGqxgnhYgIwZNsygqv5lukiPwUydlZA38U8v0qr7ovkktIAtU5d
F6glNvc0jMfvXUHU914VEQ27s70h/cRmCVU2p/5/ycQMZ/UuqdGV1DpVk2UGsLDT
cocOvMGMRblC0tkL7mAU9c1LqIRiD9KhNs1j7RaCXmhjIXJO89+EWQBq6XeczumW
gVDy94rKpRDqaphvMlzzRhJGQnCKukEzfjLDvIXJMS/GUIPhj0S0uS+O08kM35He
s07bE0/HpSTNIDVj32Gmmyc25KPGZ0vkiaNG5kLvwjS8JMrFEKLbV2/oMGVl4CT/
QdK8cqb6Fg2As7tl95fdnRdNofs2qFP6PRXP3lKZWFFFFP8OdnmhFwKNk+lZo0XZ
4dv3Rm6b+Rn1EUm1FXB5kKPI5Xr27lAqP+51hXBgIA2gHYN3pqqoRb9vHDd45Gj6
YuJBF94jmyM9hk7mJwnh24aOW711tTBWAmIzvdt0i5U4VS/YrwyunUgU9MGZyjBW
IpURlFqlkhTf0OdU5vM0egtzco23k1z0WwK0DnimhFIskvwt0wTnPVv0F/SUh1u6
y3QEcGk+Q5KdEqVbKRCUIgFXu+p+RbHeSMJtNorkiDnqwluwrG8FGWB1c518uX5A
WhF+NrQTEYf1QFLBePPWq2GCQwo9Rbm2x5BJoH3WSyhsTK2CiE2h8gqeAnQ9StyU
dDPcJ2vhHScZ3GuSjqJ3wMX1A8uuPc7PXdn7hLPx8tVhiYmizhpbKF8D3cuWx8e6
p4+9M7WCRZM1HxuK+YauhnoEc3W9iAb4XvH8MdGlt8S5bXnU0V0hL9tHbohBEykB
phXQ63VTE40TG5uf/R6QQCntoscq26k0p9EL5FLtD3CLMtST3iCj/zHtXmJiw5Nu
Pb0oHaQwgZfsL8vkOU7cIBJwjBrDilHJ8Ex9GgxgXSTztkbjFrh++sylzGXydBWx
K4znPYFwHMXavFamRYHaSKuzCAWvbF8kTkYmrGAMlxiP2lbA/K/97/UwttT9fJl/
w70xwiQOiOtQAMNM1GWvinA3f99YYBJfpDT7Q0xo403HUszQY6e88K3ZmYIbivXz
kOQs28bbFzTu5LXN82rf1e4fS0Pjoad/aRcioZF8x1ibAFixb5IYq/DmbJkyXRcL
fDiDZB8SIsM9KFG60rBWIYGm49tqetjWfWokKQJ+8yifJl2jZB66N0+k5dulvibQ
N8/ZXGHHBtOlMfEOPjQRnwbOu6/zgLwKfic55Cd77RrmDuwXIUSNOj9BKJAchWNx
d48Ne04imMEGWcOAuHBGQzlNsfr6QsaQ1O5pV4Mpstpo0UILRAZYEyXc2Z2oSeTx
izv1GGdzZIlqNGNtvEjLWnKoDUuD5Q3l2v9aZGCcB0ygJHOTGrcNMPV4OiAFumMo
9C2lnjGdXzFNDRkMJ7kK7dSLhTU8eSCgextFOcpVdtiakav+/djoarZM293kVOC5
8ceDesr1SEWNKj3iUjf3zI9+jArnDIvRD7it63zV7A31KblZBMUWPg72o2TRbacB
F+bkXcaVFiEvc2p/mZg2a3sitxLlQ7EsAHBTZa5/47V1dzp+lRFiP0of0naMg//p
2kR2OIRhbeuyNPuXpxxTJuoxrADjq9DekdlOQfgqtKk19EkzbFCyjGRbjx9GQ5kx
qPm7FdM6pz61VAIht8eEkGdjDMviEMLM7uluELSQrLcmgqCOANInWGUexV8k9U8E
lqcLWAteCbHs+zKsGzU9s94Won0pEGGJJ3R2LAa7M7qLUW4lYXfws/I9pG+Z0nlm
aiznamdMKYxIx97rcwfsaegJurIM+pG5U49V/uvz35fkfIc6W4fMTqQxA7pbTHKa
8IW+9mHTUr3VAlOrhP5G/9u8XiYrSVUwx9hI2n7twTl7u7UR6m+jmKKvZDhW4IxY
iVysIzZ/Mrl3YgnnxZzcg0PlWj9CIAEr4RiY8GdjN8HBm/vnNTMNVoqPRVYU0bAs
MxiMzG8RyGrlAGzRO8dgmWdu6585QePgWlHit3YeD8f+ULoVp3lBP0AOfv0MchTu
lWdcoyVsomDzQ6Z1a32zVVpgiobaOE1oIdkbG1mFdrRw0uiek5n5XbbivcT0g0oi
2GIvIsVosLTR/H2Tx/JEp5vInuWd0sWGUNdyA+lRanE2PbNKSiSpyfaAwkMob0nw
eMmLP24hCaBTFv/y4H66Oh3AvYK3DZaygEC/9JM4ygb/pk9BDvBP2HgpuH8h6yXS
eoK8Equ5+xiFR8xcFTznYsQhfyjLmlsjRUjCUgZbGsQtBi4zUcBOXYjG1KL2MhFB
fSbPeKUM0RkNx7BQkL6nOGsAwn1apjLeny1dBaU4eVJKdOC2L6geEeYd9RdtLBDt
HnowdwbDMaO2xf76HgZDN+2xjkBo9bTiHu42UzGdPg6QphG+3qLT4u00GiDIIV+C
JPxhSjkvJLusn8oiaKvnzxsh2F+l+PoBehFGnhq+xTPqd/ar1uNx2GrW9IVXSq7z
/LzGLK+czRT7JBm4gAxcA2179tMucRIX4zj8tALXYCPyL4pia6xupp8C6nuU01Is
U6pwhzTD3Q4ZSM+4m6sy1Mpj1BAJZsoHijfZPZdD/MEmqCbB/1R4Qp7SdJyDYN7r
2o4Z6LzKD6j6Jzi7PNugyF22mWp8RlKJ8q5shUMBsHIvpCsQwzeb71ned4ccERon
keL7bxIWKxAjAIHvFwS8IBYKI/mo4bvsAXdd72v9B4GTTX7Sd/Tdy2EoS++njMkh
ZDMp07DS8FLWoO3rvqolxv27zBTYTFTEoGUMLCCWrCXCY7iXsI2lvySZCiteUzcS
5Zzzn/8O+cMuXYEPiei1sYkZTD2D02sxMRSvYHiVflIXbqrLfdhZeXNmZzyJFYew
skbhhONDbKCy/e3DHAsa7qURbCfORLZYKQnHCPXIt3d+RdVYyBLvjmR7vYlM+lod
vUGAL6P4ouUAZnxtYuXU3prC3akGyhXCw4JNpK70p6C0UJZyFXvN9uyXLb0a6nOM
aK41ZeeCV8TLjwf1q0DWakLoZKgGi8fsv4sHvJKB1fRNcu3L1GJGOfFY6dc8GF8S
XM8UwbTo4o/lwURXhtgWkbdIqZrJDj5L2FRZE/YVqKjtD9H7m0dQ962fWsUgwJj5
VhxWWUEPlFbOSu6yq0+WQBBdL/0QwCODDHaq4+3XqCCRqYcshOPFIgYi2YSn57jV
vkmX/TcDo8J+f2xSva3RPOd5z/OB+SzxzFfzuuw04z8tTWQLW1SsXBFEPP3h2fLc
T49SJEB14BRhlYsL3Q6ql7DNaka9jhbMW3GHJFNgBki9HvUKe7WlfyDTmb/nuaaM
Pg3fN1ofnTwbN4BqT4zINea1ECscQcSHvwJ4kFI0poLnrAlGNlyKPf85FM3ri9ea
SmhV9Iron7OM5H7cjx2+PxmnMeiFHLdTjlLyEIa3tqK5ugYNlfksWr6f09jSr63R
QxzkKs1gTxkS0sxddTazYb5IMvUQ2AU3W2KBrxEw9mGh8OWasniIMPPLmII46hHH
58mkgGfiEcqQ0vzUOMkE0fsGLa/3GZOjhCoG0o9YeazQVVWIuGI841SEmeQR11YX
GlkU2a/tIzlQp7vu6eQXS2gFxLs4f9jWV/MldbYJxMwW2ksr5Qrr63lyePSI+C9e
q5LYxdkJKhMNR3YqR3X7viY/0E9JyBjeH17IJBApZwd52nVzHr/1lD7h2lH9aLuq
8PXMZbi9DsGYd6nc1IgGLQv3WfLYnnEhYCxfs5NKGnje/HYVFLDIsf3p++TuVLyB
jrcCFwirFkDS08BjhO0UXeJw2PvCjXQ5NADvtavfX/Y8eEsiwTezxeTSLc4D7mi+
Pjl6cgDQ594fX8a9JraA0znU/xvZMbqfK47YxSpxZRsqEEcSiEPMZY3K0o9LQhvK
x4QEmqhdDRWQjXOmVuDcFzUaS4JWB/a4vb7KHvGlaqrm8Uye6mMUPqwgxcWGRprY
y2Q9AkkeRuxDAdKG0vi4rI6k2HLWnhM4H4jSFlI2ykzFhWr9ygyfI5W+vXfNl/YD
ErdhrIIwqkStTILLWRFBZorkdupxIxnKXgATra4ThqN6pbi89qdOSCtpm0Nsny2B
s64GCRVSUdndBz/S1hwYTlV3P6sIZ2C5MGs7kGxavE9z4T0FN8JhqHujfRNmo9qu
ZyIduHgJ89aiBiWlgu3XJZNsmLoo0Ht47FXjbvZB0PfzFYb2EZXbVUE4xyJLwYl3
LpJLt5CPt7pNmh3vhvQBpYPkiqjCTqR2BdL4iNL4nOLefK/5haE0ocY4r7h0dnjK
ktTDHQAITQ/okS/Q2QYzJaXgRYPfvcnUpI9F4Di4Rg0ed4Y8VEeqo1MI8CRQLBnv
/kJJemXYvDCuOUlnaxEk2ZyciaKnCzfe/Mf8hkRJp+CxjfUQ/0zSbZFRgfASMIll
yJ01yJt8V1BgwxJ48CV9Cu/9+6A0j0MAnTvuqg2HvVYZ2HHIW3AF+PM4PlEuPmmB
X3RSNw1DJLLZOWxvznhVxEGOKIlkkkfaj6meFr/QV0aW+zhS3nH34FEFym5PlruD
kWANIZmzvi5sb5TSd+StLOZ9JIsOADr/06DAxmEjLfsd11V4J0s7ap2zg4yCTb3W
hcucgnRmKn+Av1lAA4kAWdfbZuRTeVmV57nGIc75dt1ZMcyIztj0PNGrqrGY1WaD
VBcnvH85dNSOV3sURpKzTMPOTWf6y6wlZr0ffGnfaTfKa9/tRHFM+3qbCA0lsEuY
YJG67auDTMP6aI5bPE6qCdKW8xanNmsyDi19YYnzC73JatJVNdF34hXIJ8bpuhKZ
3VfWtIso/qtJD2wlYctnyR2vadaNXnjFfteoCM55B1adLDZ4vK7NjWr07edJwjA5
d2DUZ0cP1FUOzsRAP192TkrHdWOWGTFmAr8IOasCbO/ZBPfpbZKGqniDjdFMDYY5
0BBTWFWer5hIMuAqWXQID6EUFf/00aZIIc6FUShxEHktDKmrCZH1xHN8fm/s4xl0
kl66PBf+Q6mlt0QuiuH38mvy+riizxvwpBO9Fw+E53uG1pVOlHO5/x522+2cudNI
RVIlIOKXcghOJO2K2nAScch22ammwYwZAFCV570Uaw0B2VGjWc7Yr8sCWb0XvWaE
R2Tv3jARupBtj2mZv6TXwxCOhqXyqtvNSlEwKXJHJZYDXUeProoMC9o427EdJsXF
mpoC2ZfnpqLm0LPEEDegNqgKtr9GZqVh6Bx+7iwuKdKOijUYq+qpxyJM868sKPt1
VVtBWNp7N7wV2Hn6z/FblnLdqqsy6veQmrAg+2Srvj0gX9tWNRcQQkeUD8nBC5bP
mqbLJdVbKiAX1gSLawmkmlQNAhyU0ubR4jH+xWVbjMrm2WBHbVwVimOaLRkQRFMK
Fawnn8NaifZQzOdlsjeIbbaj1/cpePxOjo6LWxkZVc3937IJ3Gt797bCcpFjLjGe
hZk6AJLTgtjELEt8KWKwRlffV85a/TfJBY2kkMfgmq/wamNEHh5xWK56eVfcLQTk
X10pcQBfotPpPrtpAKBha5RE2qLnGzVVeXkHkdC5ke8CNm8456QrylQUm4+bGu1h
UCh4qqbj9YUMWTCz/emu6JcaU5lsRJ790zb2yZgJYbnl/FHaEL/oVLgjJ7e3XgyJ
HUzBkmMbDHClvXWgaE0+JV5BhTUUVC6Tjd9We444zD2vUQppXK/JqwUhXNIsH8U5
YQ7d5S+0eqoReeb7qwft2sBeWraz6seli7t1GfUZuY6Caax+Ro85J8+bkBNohcdT
xdZkkdyMoa5NgJZ5ZACGGyieCQGvCNik5ISk7lBvllC6Dln8+sWUts9pYoQmvzTe
N+U/x04jXhx54v17CRBr9V3rjB4ipnjtwDUVWqZmbEoOL1Kbz4b671FmWaaOfQT9
LEDnpzgIUujeSH7MB+eK/Szg4aL4BIwcLNtDNNKqBej5NXSjeKPOF82iNYa2Vv0o
oNAUWtnDLu++CuB1IVB7cUDocG8h2GyZzDfUX5e9+CCR3szb4GDSY2prskb07Oul
HndASHx5aTIXKZzGPfj5nGLlBVyapUV3p6ow/3zA2lOMxe/0axlUyT1dKMr62e3U
t8zjPSbGVVFHhoZYEvVFEHc3UyhWp1xh2F83tc1DjPgC1R1AC0ucetDmfsTWiouj
0CcF0vkWTI6yzf0AQwPy8lgVjDPfvGCqDL4xkAaJLMfEdwv3iGQn1OQCFlUHY+rG
9kEIGBe08KYfP7LF58Zf04QuI8NXkRGAkeODnQK12EU7zLu4NrYTuKWcnJIor7hV
BiIEbSDc73/RGGmZsUlzVupXDBBsaIwZConnPlnXMz9wMi3HwRE/juFv+Z28zq2I
VUAWHp2FpABIakQHsuT0kaYzHhATvyspSwr0+gkC3EATmwqb4x/Gg+uN/Cz2lCuR
WHrC2OBxvftSZ5Dg+WzZ8BTn/BH9czds5h1yG+8gTZOeR0V31uDgbPuIP/Lk6OtL
bF+/FKbgJf+sEu/sCcLsqVvxXMPX9j0pIIEV4+JxLmXRYmRDFIDMgAHrfLmYGOty
8pfk9Mdk4NVRDpz8243oXU2/Lw5KuCHAryWkShRUa0nLQH1hXyuk+Vc8OuyktXTQ
YrTa+KLCsxvSzAz2xB1Mm6Nl5uc7cw7mcLheDADKHLUgeXx2XJr2IN2jeZkYwmav
IZvokVRaTnCetCLXDE8KZSGwxxPMFmvE0sPCbzb96X92AIRkzVoU1TMAIj1GrIgY
jJUG/+4PFloq4R/PuKTdqMUAUPDa/6fGHqPnu29beVeWA57GN0+0wvQ/y4EE0N7/
ChIB6JapoBRa9UPSNBFNyNo3P4U7+fmcGu0rGL3HOwQjOKg+DTUFqpzzSkaqZ8ZM
I4voLhnVWjNi2GHMGmog1MjXKRVv27EPKlDMnFV+PKEUSHZ4f/iI2BS5zRDol5N4
hsaVohKK41IigsQPhnPv2oShX1MfnEWu7L6JeOrh7G4ohCx/NQp1UQwWmxsqCLcQ
HIMAWO2AxNXsR+TiEoOc8tU5T/pMtEsnfE4Xhuf1TOSCyjYK9Dp0unWgZYSYwLNl
oFZZTxm+7TMExpB8F7Ee+Rx5QTPYFaD5kWv7at2KfXH2Z10jio7oWyO2K0W3xqOZ
ZXxWRYOrjOVRAU5L84IKoKe1j84joAj2CyAIC86Cl2/BM+6EyFtv9FJzuxNCDhUi
42n96IIWL0nEog5ctbhQSC3Y1FXsyJaAhS1cXz1LhMhZIPVORLmjiPZaTE6v1+ZA
kriy3ZeUUJEDvSjvdVA7V9srw9PnU1QtYlpArKoA0mYqrW6o6/1NwYCXOmD9DH3Z
hw9ropF3sj57QGlxkwvAPANw8F7o7S5l9js+I+JVE7ru5tYsH7jXL+/eW+sqRWtw
BASIiUQjlmuVKwe5YXPGG6gTKw7wr/9wdnHPlPA34gkZcKDFaNOBOcpQ7tmIdU74
UHHKkuvhDyxJPza78R6uHk/tOMgs8AkkzI7oc05KQkg91M3WiitcmFpB18Q7ikhb
cCihNIn7UolYNUbs7tciddWceDUsNk+0tjDWs1YsT7g2WYTg/xRX9fTdZAOvHcOV
MsIUCNf+oZL27lqIGwNEdLvr/n6Ud1LtD6nbiIDQ1CT0vgZG2o0FVtALRwl6MP8g
Tj+KumMvj4w+o6zRe5tKW+o36C0KnIpSStzsoysWLExrSjR728GokG5rSZplW1Dd
D/afuGALcJ51op2cVAUWDVQusF4DYJJUcIQ4+EGRmNjfgbCYlhWkb78atjNahrr/
D/oBSITazLS2Jz1t8dvN/OHsWP+GcWfm6cSEtJDCq5+YAlkQ30u1cj28fBSJCvUH
wn53KJSGdtYx3pN45JaCpHYwO8iH6ZjgUDv891IqBciF7+4LWKfwT+un8v40BVyG
rXMhWfp+oJE/ryvNIIposfH5wDtASmLoUDKj70RESY8WJTyhBfSSn9C9UP6RbtZ+
Tlll7sm3+stsR9ktd4TjsH5EoQquIGzLsezSGlfRONblhKgu4nFMPXXhe2uYMf6x
usQawZaMvSgbzgXT7BpVR59uKVqkL3mgsKPTIds++hY5kwc2SfsGAWIjvlfImn7y
W/VkpYkT/SDXbznYwiCVXvjVtJm7CEdXnkwfTTj4Xj/2aTG7ErN7SkGDQD/D+7aT
daApOsDy/gvJMwF82LjZqMfJCai+IHcHe3z2psIcV3UcI2xiCAKBjS64RQOhUcWS
koG+6xPRQUMK3TK+mBpuywZV+TjA8PbERE2S23LoaBbWPecY8a/u+gcaPt38dHMZ
1mCFORjr7O53amO9lCAsCeKfrpg0Ptl2pQLbdxgxIJIva1LNY2ddTN9SV8oXb0kZ
I/WzDoOwiqLJrn4N4MeNUpVmF7AudqPRQETeIwBkoNV7iDgvHDMIqe6LXMtlFfwe
/G8+TgdAGF4WH4nGTmrxEqoeO/BD8T2us/zsQdMVyhee1PaAHu0TwQz3IK3MG7qQ
dL7ZwMpyXF8wtiFZjCxxqGrEJeZgwIhmUbclokgKFgQseuhwPy4HTZn1wKQslEgT
9iDyFx6ofxlnNtJ6Xw+q3viTl2+UOSv+s5hjskUM85eBu8FvGFuxQXjhB0XLg+KD
yR2N+3AQys2n/n+nl7ZQP3ZI04AIQxIAUKDuxHykSVQlcDy6jx0C07yZAgXrUsDc
xVUJFpjDsHlSqXwxpUHWHZAmd9KDlz6FpVatzhAp9IaUbsOaH9aPPHx3pYto/LHx
rJop40zjuuoL3X0yIOYB4Yvs6MHyKP8hJtLHag0lEPGc5qpB+6FHMF2L10bO7veY
Us1uyPQPXj/iaQ1UvwDpnwcFYH4B0oDQmYLMRsm7KWfSDo6W5LDFaNTmHGt3Xt5m
qTQBj8N2nLWTOrZ/RJBX3m7276gHj5nhWqXWmBBoW2vjcB4ru6C5FhqczLTOwqy+
dUUeKZSmET0ApMpFuS9zg61PlrtKvMqlzl8KFt5R94sZJdxuX76PRYNfwqjYkfgs
i52TfA1aMSL3Wa+Zy6aJLGT2BsdtJ7hYVxaC64tTGi3jAeqH0bJP+LFAvJ4PT9V5
tOwGtwemIKgP6+lVw197l+Ai7/vPDiNgrae7KF3BNBu1okOQuiBJ8yU2LIiD35+A
C5eUV8JjFJl6hjnq8vwkg9k+/FarQD5BtaBvTFaWmUfeGkzTJPBinZIDvbOSXq7J
nEJ9VT5mctfv+VsW3K1xxDs/iWwWDPzQD7OPYOk3Fm1SgFSjB7dv67DF4Lny5zRT
UnYAMfKaui7owBOF7AydqfknR4ZKBr/DnF+S6VypDtdG5Vm1q2R29UNNQ/u1pY+t
x9IUH/L6jx86i6P9WV1klXAFCBijK9cyF8FreSNCb3FxV8x5TtaqJbg9bMnyL2KW
gdUQCVtqu+Gh/0BGyWFxxOxnbPrQQBs1miKsqRQC1GxSJ7dAFLZpcZaagwsrhs7B
qxyy5dobAklNOQaGz1PExJkMdK4vumZVBQlZVma2j+I71snW5g7QiWYswPqzpO8i
IYlijFdMsWEaxYM3ctZ5LsCowWYS8I5rGUmXOQN8tbbfiNEGJLcL67J1FH9D9Jlz
2DzUYhVV6Ob+62OtM7DdE26Jj6gRX2lSeNhqKhRaiozQJb0vlx6sTiXLWgqSScCL
cYDu4EqYaISVzuy/lyFKF7iz56eZl9N42HrEk+k/cEOsoj4AVi8HxTnQoE9Gtg20
LjabYix5DjV0u4/FPyZ1P6usEikWyvyY8eQoY5/mcH5cCI5sJc/VFuWYJDZgVEJ9
vmc5QoxUTtycpTTC2lYTG824kkcpyvqM94MP3Cwe19PYF0Xaehjwf85h2plFtM3B
zsg3VhOAtFLUWwF3y2Z4WknnUwM2zvm5/V1Fo8vpk46NDsHEZdNjH/x1HWmflWE9
WgyNEML2eEKWoibPa1mlZG5NbOcfPqVT8muGc04sDEpmhP5yAypdDWvKdN78qFwM
GfyaCzGB+MNE9Pk7oEGFnZm1Nh+QDH5g+vZnh+QEXdUsc+6BUcaA1gipYQgwIV0R
9vEFp+r/TFRsT5HSnc/1MLkmq4qZNtIPihnhZ/zoa/z5nuItiruakULObGz7X6dE
RzNMw6hyAvtxrBHHPact3k6p5OY+v/SNg89lblMHRi+LxcUMdka2z//nxvAbMnd0
uFfBpdJbL7UolYTREt924pfIPdhwRYNBsZwpz88kiC43NOippm5Wwlb8ZxTs0WTN
WtRWfp1ioqxeQg9gprECUJYV4BmSsxbT9vvfzzOiLmdcESMnz0QC9yRC4HGpTvaq
VA4zhvAS1nFC2i/we1vRHRdPFd/p/292LuFheklULUllcF/WQOvKyK1z0VCwPt/G
lA793cVlRjA2OTJtCugJoA/A0gkXRfQhHRZA6Xshvbdt0e0ERUzxpUdEBIvZ3FkQ
V4+vxLcC0A4Fm8HgeCkLbldi3IPg2iu2Nh6N3Cq2QbzNkOXDO0Ge9C+hB97173Li
BFksEuTSQiUmh0ZSqHo6l2Yb5Sfxf7igQtArkrm0CY5b+N/YX4cpnRM3mKgvmvPj
fILrhMGFHF6SkyBPZKuMsws02AgxPWOKUXTUcK6VrzPFGWXDBvQ2pcnH/X3cBLU8
lKCE/d+uRYk2pWKXuqmS62GvnZeSB3EDhw5p79dE9pi6/PyZJcU3yFbBE5hvYV6L
2xE04EnVgKOHC9DYqHLYmH8R0TZZnpOUh5Ih8MApvHi4Jh3oMFn0t8Aun9ie27Ax
CW7joHnHHmYQXdhPOWs4hGfL8vA0ZX0C5/QmnO7+g/8LBM8pnUuTNc8cxL2+SCq1
lJ75S+k91TymFZXVwrOWo2IYyFBq8NrLSY/0k0IaGejmRNpBEknBTr7wqFAF1Irb
G5edRMrHHU3I8e2DTkFWDtifzRyDV+JVJL/Y4VIPt1OsSI+XLuNlc+gUiXeFv7/K
bxp3i33RFjdSv0TUBzppP0NBE9qIvXf2OhnMj8NW64u+psBlS+aRjlo+2lJaVp08
c34p+Box3f0Y/onaZcIGptxOC4kUuO9V6RqaORAkdFEA0WkMPjtp/ovep+8ZW4ex
sFr0Ae3brOP1lcxcZXNVPk5rru76UvBzBOn7Z/Mf6DPEJpbY6bLAOjyqeoxlU0Kd
4ihznb4tnsyaJUboRNkyMjXgClejA6mwdf57dsldxBMR/1c1zPc6YW1nP+Xl2kkw
tnqUEVhRyas3vKm9UNh3XqY+ZYLk0xbkXVJVj8oUEcTZJuCGfcgH4GWu3v0gSqEo
1br42Eycp9Ny66mwMBXX6FGb31RRQHl2MwQj6q+hRlmkt9xX0VsO9giUuNobPRl2
s+EEIwiaRp85NqCz9nwmlxpRi5AGjhfMNPQDlkeHHmytKPZwi2ecIcV4bqSCxI9U
qlu9AGIxI9AYoSs38yVM0pb9OConKfVmTta0HoPArpMfdfKufm+E+eZ8HIWqFnbW
5SJcOlmckPJqUdxbW7tb7OQkEPoqJOSfHVrYCdr+OIwGECZ2+Kt4/4DCzm8U2OAG
T55mIe+x2nG7SGTVk+cOMIYtj6oC1xgJLaxSVQEsvvmanZSdOso+9gMRg/gPvu13
5aInLgJHJIpJXtKCGJ1UIySUQ+OpYtl2Dj4Q2TgJq/ODn85f6oJPXu9CP8+0us4F
hT9X20X0y3qmjCUIkDtz1oeqGT9B0bEao5zkaraYma9IE+1K9+8Hhm/HpflePsEr
PpltzCXU14ss0CKWD/FhGG/5ATJlKPyBnx5s+vYDAiYI1wPZlYplciyWkyiWRZCi
XKR1Y7F8lnQPjd77zeF4DquA9bcMvBonKBmkywGEYE8A5RHdTu72Y9XA7FRB6FM8
2OJun/FkmgiUI3n/V9iq8yy6vXR2LVTj+2kHZd3/SSwjgGsCvyah7g30dAgmgYqI
YxBngKyYgnmOAb4rUhFzaB/78k/TGU90fOPPEmzPctzXT35rKkrx3qPavlvJDBgy
5J0VNrg06WCxyX0SQ/Jxge96p2q93H9Dmwv8f2FZ2l5UbFcPPUsAsMimwBlWoHxe
dkgbD0XsoEjuIrXrl3uhkbcXE15BCQk22E+AKIr1iRm+dS/LKTXL793H5hT6qTSE
PVuFs9ZTSq39ZuKkWlUCg0Bucs/hVZT0skR/4fsykMD5SGGocGh/lHMzR57S7mRb
L6wY6vrgHRY/drNOsSBJUl2jroOsqewn7++kiwYfSW6DzrGwSzE7lKKcxNpyNzEh
RoofF2DOyve199fCDK78DU6qD7NJwYYwA5caVc+u3BtSDc6EyvrrjtQrWNSG5ga5
PTC9DFJzOmlZhRrzPuRRFqYmg48R+J4zoGb7SvZwVHSR+RDb00WPQHf5qT4+fBzX
jg0izSybFWAa0bo6BLBQmuyrYXKXO6a56mJrMZGmBJ9FHKQduUERDMNEHgQArZdV
jvITPTGCBQjRRPqhhNbagr+WffV8wSXQ+SPdU8I24lxrsdm2ecPbKpmhtCgCJWMr
ZojvCcq7K2ksP8yHac76elxhcUdOHrek7n6+bu4pz4KSQY8dyU9051JRhifab8rs
bF2McZ0+qfif3meu/NusZq+uJOjY19gHJFMmR/maofQAuWwaw28v+coU5265s9R6
0VbO4wHtsP9LBY4uFqHKSwGPqJ8twssvesMf9eU9o9PIEEhRexqqKta8q9qIGt13
sAFcoQWnuu240iFRQEXSJPeGlunz3CbVPwDA6b8pbFyu2prLmn/MNqEJb4Bi7mgo
yOasOsTF8oN5Bt5zriVZQPvmxPKoI8iM0IdXtDCqfvEULMGsk2tir2APbXy6C54W
oDTLotKhP/eyX1ti278XNRmhPXgsHwqKT6yw/ua6zxoglBRbfWqSfFbktsAfkZMG
4kd3cuglAspFNQYv1lSeyUFEK0MvL9stXsgb+yBgVfkv/GFnSvzuVE9Nc3tF+P2t
rxDMlgX5I3xNSZCrL212kky5jJHoZMVUiXTu8jwL9BuYdW5B4TP/jR9nzv7OXdsy
qXgMEMm6Z3MG3DxCBgEEOauFbn5gsCSMc2zEnHd0NloGEBqq7WksgpmJcL2zQeb/
dxJkbFUAHmivmptevsmhgl7sKL+eqynP7/Gfe217CNeg+n93jgZxwxs84rXassEh
wKSkfXEyO9Vy0g6hMf56FzWPWebrL8IL/O8YHn2Q9TyHs98sk4CmxwQQm+158vt7
vHRHtOD/zXt+khEE3o639iUfjBiUVFSLT266qEpBBvuLMlMOFlhSs6YRJH2/i3P1
UchFmIP3by0yIjKP3PknKR+Mq7/+RwhlHiGOUScSgg3CLxPZXRy5EDkOqJ3Q+K4P
FTTlvKAwu53ta/b8QAjQVkI+bktYiK/Zc/RLBQrN7eVSUPWwqPxlUdvvgvairgZ6
foG7G8jJ5EYBhWe5nC0W6cDxKggewAzIv3eeeL0Ao/5/fQcCgDriGgz41UWpleBa
UylqNjtqM762WdDzJG3l9OlGmNm+6/nrsY6GPpB9HD6EsCwEYQ2AOcuRoxUscmZA
WL69a5kPXQAhvzT5bdAQFweuocUyIuExM6y9dasnlun/vMOVXI6SrQjUaL1WdSdk
q6Xq7onahqJdj08mbUwDiq10xwm80iIp8pdqmA+FShkzaJUBhQkPH02TLl/PCZTp
TNa3BZBV8Ex8YyO3jNX//nneVkdtJKtWltp/3jO1O7SeyXg6wDYaThrG1KDk9TBB
IqmbMwrkKu9vxWv5f7jMkT77/E0XC4tCrxuXpvmBW0mpjQ2LxppUU6tom1HsDm5C
flB91EHJd39F1paB7SsV0LJcqTlEMQm2WPu7b227TnpMGRgiL4tUbgRh7Gd7y7/r
6bSKT+Hg0X302C20HPzNsz3y7OFGU6J0pEiZH+98ya7ceZwBOLpNRfHCZvRkG/sN
vyiJ6uWGWwOxEHBeXSOH9p5nchfynE9uQ3ki0R3/tp010zSU1cuTyqsWelcu7syV
uWbl+6Fs8BlQEmLXGMl8K0cbn7c+NmacvjgiKzow3kPGxMfwm+nBZvrdLLppQkIw
nVQIZPDnrmxE7hfZ8bUuc7jfO3QqK8Gwf1bwNECExbj1Fs9KkK8CtkLZeqv0/dic
RZMAWoCJXC+3G9fQYOQav4VXyvGxQm/Gvki+DA52zuuwoofdV0iaDGXK7iO21IFq
nqUKAHI/aVfZBf4ZoOxv7GuXbFTYVhulwY6y3rZtIIKWBpjcnjKi07GvbI+W9LLI
QiInEcWOcRJ+ytOweQaZ1mPy/gC1VdOw2Flcj/JpM5iaGwLGwe6QgE4v4ebrZVjm
jWJUVPAuQAKzLofayLaK2oDHqTa/DeieMixnbZsjO1DkEx/I/3PTgwMSBXXCkf5U
bEjiaYSfDOYMbZV0xX1Z5q/4DkpVe1/es4MbmCHpNz5kjtfscTEhVTlXTadC4vNL
GqGvPPZPdTVYAMnkdK3v1LYtYRDX3LFY+SoeebYpxICcyaLjDTUGONcJTjk6+uBc
J57q7xGxvUDroccFzvlZcK/OuSIYWAdjqL1bNV0sMa/7IxIqT1z7MFuCzncuqaLV
eo/Js3pwJdhcSkKkDIgORplHe9N9FeNjehoszcRFPcPF3lX33Rq7j2Hkv8VCoFdB
D2c6TIN3UESygUUVBZdrJOT86H4MzfiSlYCv0EACLtYjypRBF+qfIE43LqP7on7Q
UEJbA72XrcFgmP4b+nDVBVB8pu1GXnnyBwZgRi0A1f/IoCTEwNQlV/6jOKFMWAkO
MS/0DlNgw5u07e1d/rJs7jcvr7BMdkXRm8m2F0aJgE94PjlpU7CKyBNVNRLMfRif
kgKtUhCPlhWYSQsE/mFOW78jsnSq0I7RAToURCurNNRNdcP1Iu1uXuq4vCnW5qlw
nuZGqA+BPCbQtlJT8ZTxrOi3rIuHJMXIjf04hGi/DKU+Zj4hh7gBo4JAxvKkKGAW
3aNU4nWMjmRH04UjcdgjaaQzvZ5GUmxTW/EOenoWjapP1C7O93L0qdG0M/aq81Vl
caIOH5KRM4whNwq/4pAPAZInqANppE7bMBKYxUwsYJeEhEgjZ3/a+p4gxTY8xCg7
Ba9iIGyQo9+OwbSnVMxmUq9NA7d9cQFW+bssSfdEVakijd+i9DwERqFk9xbeBc8J
ebsXl7pBYE1LQeE8f1ul6h8J9Tr1jNAhNRMW/ZtG9K/k77GJ4CsCQxcuOqZGXj2o
IabeLrl1V9s9t/fq38oN4zPLa7CcPdeFNLyjZxYVuq03IUgkJNAbpRIuk7dvKMUk
4ZvcyibfRx91jMGbWlT9DOUmL14SIz7tvjhmVYASXbi4d+9rRpIM8ktIyoIs9VQ2
Td2x4pmcl/pzzXMH0z3T7cjXylvvh7+B4YdjvtMFaP0drNX216TfYAyrvWeMvtFn
1WColaKGrduZjOWsOERY/qsX9uXMkgih1jv2cs4xh/6GudUZcrV+tNCVDFMbHNrH
ake07cPeLd7RzmFkDMIZRVgHzf5+QKt1tWfZjHXCl0rkCN7EMHz+YZBFGodpd+s9
J335kW9K4teaD1EYJanv428hd7OoC/v5xlNbL8xyRrG/MakfSMZ/pqLA5jVn5oI2
sg2J2mmujRiwUvuDGBjN6Ldxqxtg6bVEcBkcgSa6u3YkmejitJ1SNGf8jWPQcENf
7iodp3zyrRs4OAPcHrII54q4zD55P6f73ZUJopV3taUJepOVmLvECo++KWZe4s4e
rrIXJtVcQXP9jTs5fE8iWJbdY24Y3JaIsOHlsQAsEt+KtdFkVf6a+M6dPhW64k0I
YulDeELwl35wY2zc8hDzv113pmCDQVZcFgtZf2blVYXGLs+wLBYL088lNsf00F7m
pvCgxKuOSdFvAuaAuFYsC1AmBIzXGPkhNlzjL5xIauSxwbKPCjNx0OtO6B+zdxv9
rr3u5SKMbKj5HTMIcFNb3B6lkeUboDU5RZIGj5UIVEL/udtbYW5LBxt0ZlIpjumn
qD55CkYNzUq0M2nUzr9CgnXMfW1C2T5CJN3uI1nFlDbOj2dC30B5qSHbe984hkAg
5xw8U36867iFgl9V99HW9TEZoykHaP+CM16lbJzjp6lqExMh6SKo3Mezc/vMNo03
eOjLYmpAH9snpdqHAqJEDCxbY/HlTZ9ByejZ/NkSE8EJopSQQJ1JhSdOwSZxspPu
h87/OsgFM0y3j7yAFZfqa5MKGLjjxZfbyP+ml+0EjoWSWcIFxTOiUlWcYETicuS/
zr4cVv5Pg1nTjoD/gjL2rPVEu/uOdQOOlOYBMgYcE6vYg7untmT2cWOfcmGJJws/
s7A6VOV1SuaB5t5nEwTxBFbsL9D4fcQImkQz8D4p23tXULD10xbo3K1758n10+Rr
1242wXIsi1blPOTx4dqlq2/yl7+Sz4AvIwprAGrmkRRxrJfLLLZH+z7kfFcv1ChR
INumDSHseZ69Vf75wv6Nr3kGUQL0bcon4dB2+XbJLvH7ePfmBmLsoc4I5cyR/m01
V2VrgCgLHeSGepjFeaA6OAxih6clwG0joI22r/lahPAlnuACFAcA+MijmpQIckcM
xFUfCQH7Kj0g0H1pqxtLOoEGoDzEA2+UNg1SDKmGKjbsoF+ty9cqR3zyGe/5f9o7
Hm00nanphyj8Q9MMr2mtzgzIuFR0dWDIbkxJCK3YJue/t5wdjQVIkke5RMSsD3k/
rvEx3CJs6SkylPwvNeUTWYH71J0yNpZ4gtAfNoZYgrSVG29xzi3Ooex6GOla64Yq
Se2GDTH3Z38NrV7XhPXTWvp1DRGl9HbdixTozFR+p3w52kBrRGtiF9HPbS4ZLvhG
xg1TfkSiE1fy3rFPwoXpHyhMEZvmaSiPPPvUvcn6AwCInfxEQH5m2+5fdnubgchC
rN+O9Klzh2AgBKfHP2SWr5T7jmlyqakxBTAeUO5sQw+PgK3UR2nfe3HSnELEdEtl
GVShpRyQST34xOiQIqVmtpfY+IVgEu41eMS+8OIXIXYuyQE+HwNENgKOfgDDwXOp
FS122nOJx/a0Lh1J/+f5s2af5EMfPWh8qu9kGTRJRAwSWaC+hrJ3aVF0WzWQwWrV
hT0ksjCCKkk6z1zrZJkEB1UEWNWeDb8U2w1IXBh9uRcWAdYKQIdtT0YIk5CcMP85
Boqbsb+Lu4DG1+LtXnTYqXpbI5abB3DN018X+22/Zt4FGCv7+pXERHoOqzEJEVxU
uoCq3n1+GvfeyqO9aU78cTm6AKbPqM5ihXJP2sihyf58k4XxIpUmMVf+x1NhcWN3
JhOA52mh0VOAeXMeB9YOABg44DJXA3aRMlnNpAWc7N2TPySsMeeKI+BhZskQ5s5Y
1vj7AiHeNrFep8QsOxdMMIW5nyiHt0SvafWFZLsveCmUY7UWqHDna0tDW29UHZ+R
QOcHOp1p5ypBMVn3MbB8ZIaJYMpgX1JvySin9cH8DXOqyGFRfMHlrb5KyMf7elbM
cjR/KH2RQZZpvkGpKU5baRooXw9s7hq1mkBqz6DD//C/IKMkKtw/+r8pLpFeR1wW
S88FfnTs6iZg8hvwv/bg2bn5xwX/1kIoIcKrshhjU5dxrbHsp/2MwTnVQ0yQoKFp
MBpj5gPynBvvFCIis5Y226VjA2AxtazVOgygsSvWLVSQ60VjsrFi82zVZDCJtuDh
H5rPMHSECUf9OnICuteYOPcqAsp3eeKbxV71FxUaZWq3YNDRqfZNyzKiKzST406g
CzyFVXC/Txb2fkxI+vmWke/lP2FtxrvA7JH3uzYXhLVyjXn0Ds99bnOQHrDEaswv
rqeBG1FgoT00cNPPTpKOFXzapOLZmpvesJ1F9sO4dmgy97XBW+TmvdXHwABe+sIx
KLJflQ8XfdiDSofznfTJNsVcbX7QT+2R8dhREpTJcpn6uTfDGA8qywAp2DTWAMMD
S9uaYNA062SHf974NeK4X0r/VZLJMJPAxcsliJXjHwFUK8i/RB6xeM7P6kF1HH9N
F/HmrInONGm6vVjNSTdMtUkqXtndf74/aS92Sxq4L6BVIgAhzKEJFu1FoMFGeBs6
Fgo1E9fc5cgJUlrshYM5iYLze95kH/xPeFiHE0ttEjb5VZlINhYsNIku5MEPdJfd
/jjp89l/jQSiMqeFgYDY5NL317d2CpjvK+eePJv5gt4CtwK0x+C0ZB5K4AR2kZdC
hdu+M6ij2Zv0GlbBC7ORnreXSOZOxHj2nto4lkQG8/1329n4Xv6cpBxH2ekCnk9c
Je6ouHy6ly3c4eMUcaTlISeVt08Y946OiOstlezqXHbmKyVbbFptjooz7FahwMJ0
Y05XU8lIRoDE1rDubus3+Q/oOzL+q6pNTnCmpQR30a2DYHIUtw+zLmAfvOHNNKNx
4USJ1shP1J/VaTskeIt3i6V/hRhDhFsZY8SpatrLkX2uPT+c9mSnZluQrwl0uIx6
LAISFmCCj3jGX8e0WMbIyZErGpXSbEWrKms5VAIhash2rX83i6LC85cH4Jd9avqf
aFABccmgftvs+aTbl0W/r5iJvdxzZiREy0kBXzDSWm8/3giv6rwiT/vDmyYVVr25
4DJ4PLOB6pG4z06VfFudzKML/9Hwm0Jq57C0oLcJxi3u8KT4wlDmqZkdC3tyigSs
/2P7QfN/2/JeiSM2bs247WXT1G0Fi1lkeZYPqUELi8fuHCtsy+Zh6pbD+Gksym5r
m2CSQdR4FAmZybhvCeR9FTDr/SKdsps99bjh6I6JLFMy69OLdijlOI1yUZsSqjqv
B4r4LqfY71AtFfgY2PdaMjgNybsTfcKPjpfbL7Ophx2PB2ogg9rDOzEYEmzisHD2
VyVQ3gnZbgJL2HEpcWp4GUXXG7B28JzppYTrf+DQ/FLjbg71ehnjk55XAKEj7xeE
Z6xaQ108dz9gvATPwwFP0qb3X9wY7rrGyIlZ4YF3WHEmoucI8xWo5Ddfc8kMTA1Y
taa5FIGIhJjxVZb5ZykpczhcTkBQky9LPj16OAa7EyFRn+AFJZc5fvr50ygMaTss
Cz7mTipeDBIVxbwYQmXXHou/AgWgrat3GX8pqumnSOOPnlAW1krxrvRJeSeqCSkX
O0+u50p5XZITwKObcBGzf5ASomti7M8iiLnFIry0gwU/vOk32eyyfN5BfT0nkObp
LnQzGohD12e9Bz5dyM58DftosQsGZZqFoUbJxqPB6txB67mYje5GuYm9QJSoGcls
7xi2XK2hJipGDdPq2ME66mR0f6ROj2BKnRH7PuDbJ64xTgimd3yW9pnPHyF0ZKoO
Tr5v4r7+f66ts15kv40QBR+mT+KXAzAA7AIxyaXLaysmkEtcpYrUlrdPr/5koXop
ltNcGm/KvND1r4odi4bzEikVc+HoSp4o4udLdFj7VQvdgHScAEpvNs7A2HZ3xQcG
TVKpme5EVdkK0BVjb/6a7J2AHNL9xtPaxPp0JC9eGe6/qcogyWZq32KLZ5fhmvOH
H4CfkoB8ZisHMniHd9GhZQqjW1MX2jzbD/GdxQsV85og76b9vdn7iiHWsZGVPt+J
MiiSUHGxu4lqzFCf8UrQ4yeuF0r3JE4mnRjVFKXZ+l6QO7gppnU/d9aQT9ZRvp9B
KHfacuW6gGTJ4tn1L0gaO3c4ChiY7VyBa68rd+i6TaJFkNan0f+fCO03iZKC9qrg
aZD79gXZyEtEGQ/XvFcx1WswztCzF+RpHVYxS6J4XjasEsLBKDK4TrzPiBD78Gwc
HHshfeSyAFXV1MKInKdLXcp7V0/QAxBvF6HlErYvsU9LdiNNo+Ou7WuuJQgQl6ll
iG9KpkITCt5IU/MndTqN9fxN+lJ41nO21zpqHfRwvj3tThfbmLt+apFnmA1FROCO
ek+v8I3mUpBKx2AHaTmhroh7L1Ei3ltnr+jdsq6gGKjq8MPkfo0dbawYHWynkaDA
E0p0aS4OKHELHdt7DqnFMpo8OPcXrk2YxXae02heC3uMT8xNLh7RrBKWJZ726zA+
rUlbchk5BSe9HMQBKurvfXTkT+Vtl8CDgVwL+ee6Pxe46h4Zt8LbNek4hzPbtolK
A6kIe9Wtu5tp9Ic4xVUybknuaU6+lwvaLLT3EBMLbhGG2EOEHuLUxE7xnHUPDgJf
P0MLLALvK64LNIh0vttxIjBw5B6GEv4ovSzzAH7BYVgPQMKIVVSGtJGhrsGhEbC4
eo5a0U1nYKmYug7pAFyCyiIVvqxhn5+a83YcE7G6OGIp2F/FjsZeLEtgvTh00VFC
rbMwvLpUBVH7MXUF/EC+KVC/eccg5yPDkYyUb2rWxY7ILIkjKZQa3M7x92CeVb0i
RmtGyo/sMbL7VHb5EU9GYRwdxnZpUOViZ+ZXpzpypSMI+p1wPtfj5Xq3sjGvpeHB
lsrXxrzxDZK1geM6vAD9zrdgzy3p0Q6MkTHI98mEEjdHtJcU00UL1RLpfJMRUe8L
1A3E0J4Rebrz+FUZEQE3e+K2aJ+DbugpWjtXqtnoHb/sDKj7anlR1A0XUwqSrCGD
81XIA/3dT8/qKB6OkmcI0FiO3AimM9zV4h/EHgVXAGPPq1Lkoq5z+VN/swe6fpPD
yn60s5X0F89e3jfNGnfKcEs0EI9Xd2YkvEvVncR9+7Eao2MIPvwElifQnS1krrkz
s7EPNEnYRnZVbijkz3R7hezpzsueG/P/9FQ5y84Rin7pTCwD9sAf5us67ir2zlCh
8yZE0LLBkT1NZqY7DCzPcgBY0nDveX269h6RU+we5WtZipxhO+PRImARa/XuqMDq
IVv8I6mR3VsoO80ORzhLrKeiO/ccIPi1UwMK5/llv+YL9V8Vm8zUF3Fk84LDIdqo
nlf8kY+RLVoa28KGnRR4DG+KOWgcHDiA4r7Nj3jX5X6pRD9uYJtwsH0JrFGDt/mH
Cjlds+awCZ6zDgy4fv+6Wznc1zqi99ePfnj4yA7oFfgeEx3+uxiP/yMdEDCt3jkz
IQaM72RCLrbKR3AEGciSnHLAXk/PrBE0HqPi9TOXRV+J4uZZfNLcWcaSHYFJUJUB
7cI+qF1DVtS3AkKzFi89VaLOH1U8kxM7ZXWCHFmIMibsMam5xMVXlqoXiYR4XIcW
m0tEIG/46MoLCRUbLn6G8aZhAxngwfOMEjRXZW1NIxbpvM8VWHJ1v6CVOv3UU7xY
ETzctQTv6KJVdzXIlP5MFJBoQ7CzIkgs8L5d6d0ZDZ3CuNOODuXD9evTDGVlqTJp
bsXyEkjYg3IvMqN08zJyh9UFuRi38lGvbp9/IB2rwi/BlUeFPWUZeueI//cLQPCL
vb2/zaHaR5gn57QGdTz3zVw6jAy0bBjc3pvyWO/XBOe80B8H627oyeVKZKmf88uO
ZdzM2WTTGm6DQ0Fp8jSTwRY2fEltJs3KK8zZl+/VSawD1bciEIBcwV3HKhLZwIsU
r0I0YtbPMG+Y5BZ5gGc3a3OdTRJUXnqfBZj33Ia+b/K0Z6HnjLT6hhnt09rG6hoF
cw0nxIIIIt7OqZ+lEmnH9fwZKp/N4TvejIBpS/3GfnSH93X39gpm1kSznjKFuYsV
Yduu5SU/ve33toXSWMimZV4nxaqUVf6ZXaSepLs8WlEOjsG/tbEabhiYRqY1ormS
eExdhilNxeCi8YTJWgKR1q9ojnmWwv3mKyppqjP2Cz14zmmjRF4lva7/ZPQIQfAk
eX0ldBQ+6fWQ6nDCoQmX/zsC+5pAdskzAToc0f4nDGKdH8tdD+oIAxQVTe6CyE28
Gz8fUc47x9mlDVuYLd0OLpfgzZorPmbaAsZViLFaXYUIMdeGdsL3A9DPC/nuOGxs
hFy1hgWUSdLQlT64zX0z4sw8161Y6zqBjYcJInHVhDr2iutKZnp9HNn0K4kwyUZN
PRbTHPrUTMz1TEEtVETIqihkT8PKrjQ395s/NVAjbGBwtcAZJTJ7UoNstjY+RmEn
7vQR1grsXWLwP1D8qj8SB00ELkewE5CLnLf3XcxdO2ZGsYOQYwUBBdwZ7RJR1chW
alrNjKFKPO2azJJ/WEisxUxi1sDIbjgkfM/I7LpVhZGU5UGAm7GGC6auRQlkVaq3
BouNmCvxBt7nTNEjCHosXcSl1bU7DIA9IU9ehdEZa/HxJ2yVwsa8j0x1s/erHKOH
vu70VSQ6rX/Reh9YW4DZWubCT9YR6kUFWMVS2W2wLqcH5yfNO335G58F6cWMGW5o
b4jOMeuXGSAcVebBb6RzAUCHbynfJoOivnFQLKTZsMWeIuHbScoLvRRCRNHakceu
9CpHbwW2PsSkb+DRXA7CTMwYq1iueuSLBSPkonxU2oQKHS6TjixRyihZ0Fv9+vzF
hTWR9Ud9DqNlDAzoKAhsoDQ9Cjpak+qzvur2XSQvyCZx9rozQ0txh2BihD+UL6lu
2auY3TX4Z0mY91amRJARCpCwvFOhzURaRX+V31E8GNwO5CRPLXFu+9S3PucFosUh
u82kr+7XmO06wMOHet+U4XPflOARSrEFNr1TSxE1/mJdctNgm0g1uk4Y5iL4US5j
yjQMPQD40pY8ZSE594maYL68G1vBsVhDcE4Ear35XS3C9U7Bwxh+9vdCwXaNa2hi
OXEzRaswireCg7vPwfFqJFTp4k/Q/eDug7NLWbR/8ryKAq3OKvyUP1X/rrPmINbC
RQUyKikDPGMibCP0DBeKi+CVy5z6+Ee5Rqx7ui1TWrtY3nF33mA+fS7jdkfjMvTy
U15YNeKYr6Ul6F1KGtqmRn2QouMuJfEMSujHP+m9Nc4L7lC5GQB1cyasfkPZO7Hl
R8utu3Fi/YKbcyizBEAXWioCnQq9PTIMpBm2pWD3vDz5gyUIZM+XZTF84l1qDvIc
8L2wSmHV97yRtCNKJ1smaOCoVvvD9c3u0dkE479ep/CczQ1UZFTmtwTX6GgCIa9e
i9ItpJgBIsDdV3/nhb721RLhaiFgXviM11BCA6ZixVJR65gciMOHshNBhtNQo8yr
7vdLsUAF9wXuW9EIMQDv+Zk7pb+qy0yd1CnXXNFx7XjKrYY1sknhPb8KWGOMP0U7
+u3p7w+pThIoqM4D4TgyntAqTmNaqY80bwchZpurYg0z7HTFL+8RfT0HBuhDNTtD
3FD2qmn5Zc5VBWWdI9xJHZlTf2D+cSeSd1YggMKsH9WnB2bdjRdbJ9xU0YVolChL
3TEEyZykrOLLXVS3tpP5/ZFf1oxGzSIZVoD/9fZRe9lBLy6OPXj/MUoGGBWkRp6M
6Xh/5+LNkX8feGmmCoFcvBnREzictw9Ncr6vFwgD/VYov0v0gJRQ+fqRR+t8etHG
NOdYuIGc2C+DSlahYsc3gB59aUhyuGPtgltXtEwsM+gbuMG0mtM4/pvRRo4yJQq7
aArokeDqGxxRSD+taoOPW5Ey/L9Jdjd0TyWSys+xOGGt3GVooCdsvxHu0rbjOMiq
EtDgaHVREDka4vp00vFy3MFaJbXycxZBp05ZjutJDCSd/ECwTnzH0f4cWAETb+jM
/VF4hGlFQXsn3tM2KCQk74JId84NnCyCunJU/kzKkg7lck4qWjvLvDwqeVGKtJVu
/y139s842C+yAe0iAhlmcdFfSjyzgj5CwpmWOG0h/IXO7OOhJzMxrLuw/vYrqCou
Vv7sbWYLuVp1fpdjhvrBGHye1xdzPrRrwZLaT8Y0d7kLZolCBuERMTVG7KsBVEZH
eBxF1CN+weN3xfcdGv98wI6GBO1V+Nm3TwKD6570XjyU7BVQOGpQ5tkBX8tBbCU/
oaz3Kk1GzclIE3apejAkS7YlOwQIAwATIpgpHZFF7oDhe7qOZfYg+hIf/1KSqlnB
TtHYRP8k6SeJskYf7egcQ1cBT8uFXC7MX9Pk/K8Mz9wVR2srzRy8Maw7D8pxbd6x
oAdM5n5hcbwj6WGZKh4xhhsxxOcHboQUg8L4OXl3tY4cjh2Rvf3whJ2TEucy1o20
5UbSOkM9AwD7PRN5rkOR+qAieqbftlUMK1ir8EFEJd+aQUr3l24466W0wGd5Vw0i
PN0RYjvYHNsURERnpcGK9T5cHJQCZOXx9gmt5HaqhfpMU+2YUiyF2feN24nl++DQ
t2EcXhp3pzvxWFRo3ecYTSqb8F3s+rZRhCMF4tu2i+8cq8qkSwiBmWyujYlNNsMe
N7iQ1GVIzN+hTNQUaB3SBwFf2xWJoFRbqeZKTQb1F6s1+T24plyQyADH7whfalk8
vgdqCC09t9nbXHFcr5+u3ffIkZacSpNG+VEl0lxNQETuRrjtOWOU9jjTLRNaym+s
T0+otWlS99o4ehZ5stkEeSkJX57uyXqb6s194BdNYAhEed5s7JO4so+wicf+fP7A
Wlky/zxBnMYWo/VD+6Us0A9eX11yuRttkEo9IB2IU/upsidD66HTFqeWmsUiZMxh
lQj/KBj8jGDsEcZ/MOeX82iSv/zhAXUwM6+B5FnC+Ba/+F/t1JZNFT6F8pjKvgZn
LDqHSMqJ1X4NY+Inb+EWl2cUg/GQAIqyoM6DnvGmpfhIHNHQ1vac0sR9TSqTUMlF
fF/mRG8H3IuxQEoOX4sjddcUjv+pIBeAcDgGGfSbyY3Mud0V91s+Ef33yGKsla+5
sVh8C8ftqNxSkJe28dLI8T1+Yp6pmjRzOLRZcPUggycyyTPBwBUtcMjUVTmxNle5
vGN+E82GOKNbJYlGQgAMf90RSoLOsPJ/6SzrEjda+dSgzfShtx7Ltg2OW7qNgBoQ
6plJEKA53zzh/9aZTCsKdhio2FFIKsLDhnqBMaRdkJWvEU1w3X7RsM5ar2Q1f0yM
uVh9vTd3c9V9YZDqaKxMi+9WIHmLiaMSb/Nb+BgLeZoDPsIdQcmYnd/AcS8mMWmC
grM0qakze6J75s6eHAYBXYLeVINdu/I72v7q/Zzlj+5pIK+t7YZFN+r8fSL3rTda
AHfIGL/9hd9WR6PXG/mcvPgeKlG+3uyZAgAha1lm1m4PHbZv7jlbas62Qj1bhzdt
d/JOZFqq/byQR638/eg5g+XmZbdVrKhzuK9V7YloNa7xoZB+OKJXxugtUBvftha7
a8BrlPcWC8Vg83a2P6QKxtClJMVVvkoERK9mUTW6FMkV8oyDN4c4+i9WP1E7ifZT
E2OMV5HW09T4Xh+gpqzMZL6jg9ejDg6zgLZsO497mBIwgeQ0p1bSrJ5FrV7NR7IT
YTGDGMtTBVpkPxjcRno1v4FEw3ot9v4rohore9dtuBsDDmDwrOKKgCuHv10yjMxP
JfvE5rCqGCYLbAPyQhyK6kONC3xw5Y7ejXKAtGInty4dhJmx0kgVOSqJ7RiDApY0
8qhywasPPv7OR5/09dZuVUWeX4aopjiS6/iGyYqgfQMKviL+WP8778yQaanTnsxd
B9ZYALiaP4FmkczcOg4d/13Kz0T5zejqJ0k6Rl38TMNSaB08D7RQ/p+GFxLVobmu
nN1cXgfvtoqbruBNlc+f2vL4CVlQdYmhrMo1hCehxz5cZyapDr5Ct7ryImeq2on1
nJu6r47rzadiX4kBahkAIlEQXWmxIFfd94YssJ24kHTDtGM8o/dA90QO/CUGvULf
fMUpx8pGnif64GLF4sI5LwxglOvdJdgYdt+YMVDGPxbpvrCizg1ejy/PxjLRhWAK
UzsNX4hIfnyiCh1EtivqHlUSy0lvIWsDwkADtg52ncmoz34ycDQs8aSJXla/wBgf
/PKV45tYHcndACkcqrlfiE4u4pv2fZ7FTHLkkTEid73QmI197aAK688xzFZ3HoMY
S0fjHLPrZk0iaVIghoebyDIQ+Bn4FFC46McZ3Nsh0CVTl99A4nC+djfhrDS9mB9e
7qhoXiZHnJQ8xvb7GSIik39rjcbC49ngZOgw9LnH6VW87YZB6iZihkD/Gno6iOYP
9xCvd76QIy/u7SOXRl9ApfXWrvO8JkBnFeKnXytu+fifSQyQAdz3yhCwp+KL4zdf
RMOLGkU8Essi98xOlsdVvCy+qVe9+mlZJkLm0hFGEBspz7wu+AP5y4opdrhxG9ud
lWihjmswTWZsU1HeV/uFsVe/Mdk6pn4zyNEmrXAy4FVR2ICCzWTQrWj1iiLe5KOh
MKKIOu8RADBpK3oMVNx7ZB0r8cmw6FphyvK88Zn424T58rR27f+X1djoKTnmxWbl
yZUlqWUtY7OUCRB2hE9zLaHPOVHAqbxrY9Bio9LFVjsz5ac5BSgGf1JGSehMf72R
Wf4gBed6IN2iAb8XIoRK//UY7LuFNSv8SwKrz3YzDNfxZZ56CJgYvBqVg/Pmx+ZF
ud7lMAmV2luzSo4RXcmFP49qqchX73reC1ujb5E+OHawKAwRCtAJAMCsBKTzYknR
a6xpvBgSjc4+32kIPtITlOO9FCN0VGOXY4L8nEM29kP7O9b1zuyT4IeWJlN3Mc9z
u5rGY1Cu3w4/IFw1toMDVqI0SARduPW1VdeZJlLZKuLIiBg2L6r4PC7PGK3yAAyF
UntMQg+VcZ3Lyt8E4mgO8aagO16+mYG88z18jwHYzzRbY3jis5dqTq9FL8s+zLLI
AxbHs0Lm0UqmltvwFS0kZmijiGl6OrRCD9qwDjfUoUvIVGpWbT5MBbtmK6oq7zzx
6Rj3iPpYWCx1XZFZzfpNSS1j8le83+JAlF3mNS4pa2RXSRU53XtmZHZVqMsz0y/c
8tUNR84laiSnKxow/YeB3kDNnFoUsAP6LYweYV0kmCGH9AiDMRYNbyCM8P3zxZjG
NCv0U9tvl3rLUv+YvlWcPrt35iVeoiP1yFrp+DBGJDXRRN8sxjjh1hNNT5WWCDtN
EyQVsDAvG/bZAfU9rL7UPhI5AQ4yW+rKWx1FrLtMCqlMF79Id3WP69RDZDHmW/la
51ku9/Iy0MbnQk9TsqYXsiYHDnmODHhN9mUonHGjuXGaC5F2t3pYOrOeQnD61gWp
BORq9x0+odwfFo70i+tqT2Tm+aDOVuPsmE+fbV/IH3q80dBm6U14m8OO9ESMtSMr
54l/F7Kw3f15W94SxpVlGDIaqle8WG83RbZISPFgocSfnXawRDrMedpz/xCdJO/L
KTF0KhAXBMcl/Fgy999XjmnK0shnb6VaagTQC64h8/5yRxXGmnrwPC/BITCzHXbw
hGXF14DnTDdBf1ZrgL3JcHOygSpFhKADNqG9oJ732FxTUoArZ2pbOo7CMWV3ZRHR
vl652LI56TbQOp6y/o5rPLWXMfMh0Te/NQrqQ19AOP68ACdyKVFZFDDhAPgZumzM
wmPyMuZkIQViYZ3vesdWKVkM50b2pqBdTzYFyC0Ccp0b75+MdooE+x1L6krE2OyX
ZoblOz3KB6/DJw+X0ug1grKY9IVLcBQ+BeZfMkU8u60Vf6M0VBKrm64V9RqXxP8z
EogIWgwLdTdFZLPNlGXJdzf2jeZuwZ74WeHcaCaW5sIPWAD3QW6/uktKO0mordxI
mR7aMP+54i1COg966A8Un9OdlAy6I3cDVie1B+2FwiUc3sN9vGIohBeeiSIRgF5h
BY71eWm8G1aoFCki14s8F7HYUCjxvAqAwLhxaxyfqzHNBnYSHlCb+gWsE8C0B7P8
mxdNWWVRfjoyxnJuxS+WsjMI9U3GuIEDOsR4AIv/S+9Xdi188LxQ5WqkmJL/71YG
NZpKswb/RQG4abjwia1MzfpvT5VX5Uo1ZtDjdY2cVAdBgJxBRG0kAILvwlv4oZav
bO/wq3rArAwxfZzN/VcLUhxR+QRS8OVejj2Ma2pLD4EJ24otfHw1kE9dU7N9DdE7
rk8ZNgRGCpNFwHzayy3EnAyTKzQm3SyFcfaKpSvo1H/PEA/FvIbQEsPCgd2xjBAZ
ZXnIIVllhzCQyTMxVViOX2UBNmjFIiaoCif+kVzdjdCbyek3ZzBX4mJG/MLbDvM8
gR63zrmZEnCrMeqqOyjXbjL7o4vLIMjmdK0gigwwlzp1xar5KuREL9HA0f6tQDse
1ZzhSQqDYm2ho204XpsuTVHST1cKC6hVpU2Obu5nKVR32sWgQMTXLfsMZD+BRBo5
z06XvwAN8BMYFTeaNTq9UNupaHkyUcck2axOR91RQmSq6Qx2qpjJvd71J6YkoA/A
DAg070T7YSpRRmYUOWg7O/+aVgZeJridVo4qmNy2t+IwSvFI46n1onuLaOaLpomO
N1e4Kh1pbTQN1oB2CoFt4BrRw29TFjZgIP8tFxR5ONsVcVWEr0VAd0WtzPW4cn1O
4ZrzDRvCOqOCOct4XgxbSY7tnBW3anL9dmsSqy2xEKlDc2gnA79Igfigy6CxSIun
xzIYavnjMRysmnJiScqi9jhrRk87rorts4G/nhyybdqubfsdNIfAKkUBiJMnXTxM
NEtQYpoCECf3S/R0cGA9RPf9bqxeQnQ5/Pee6avC5VRSHWQU7WCji5ZnQuAZDuFJ
aVU4nZ6qfBflqeypVbjkysk7GFFP1fuEME9u0iG3k2neyJtO3dWUFkJxZVfM/Lsy
C1yadWPKtLeGLzZAqTYMT/8CjIxBQWfOPMvGQM/yI9NFKb5gpegP5nN64a46HCJL
48rtUWhxx5rW2809cxycJ+ZhXVp/Pnz1wQFagdGCrMr/udg2YCRIbQ3ITWJJL32E
0r1+0DrWT/fKvodxiFk7k2IRZ82PqtZXy4z8EHqQcyt1EQlIZtE0pJ0X++EoTvnP
4Y2OQcTnotqqHTwRIIhtLEHWtwfK3qbNWaOrhDQs7cq10Hm0jtqjPvalj2DFjvq2
gVwrv0lY4n2mT5uiVRARsdhlSpoHgV+MP0pl0HTm5strBWxq/wMJL637mRZwU+KP
kN+I4jaO4RABoy0wo+2TM1x4Av+G00uYhzcnMynnW5S+LdEwCkqVgtuwZGt13y+b
b3DSnrO74dc8pHhc3L+YrScltQkuzHZ35u2Stpg0cnR3yQxlIZ9bndMxG+gWXGdU
hLmFxyaE8oelzh9rM2ZTeXJNdHrL/nfhy4qmm97jVpBdlzfbirWUiN1JumW/JCYN
yzU2s5oLiHq0JO+ZlzPyEkAsJlzKg2VbbjmMp7evaLTWOkIHJsmtZFWobR0+N2JH
9q58OcQk6JRTILkxfnspiIlKLWM0idhgSMzAyiVvEltvxc6RT4wXPMKE9U0Pj5l/
8kcWsu0uq62/Fh4AY0InWOgVgnKHfhGt6lu5dTvXq6eOmjaVRIEYfc2mfoqpk617
NziIAt0bZLbwyS6EkLknR003gyF60WUALT5wdsJElV9ERwIRqrGHc3jI/CzFcd5Q
DDVb/TIjN1IJDtABtu8UN8It43T3afJu2grHamdb+rmvs4yFV8OFeqfHxgCtVNVs
LvfIGA4yd660O9C33gXPqYUut0UT5sNQxSDR3i34BP+Q6ASqD9WC1mLu6gC0ZlXP
DR8wLW9Y6KtIVKMAVa1YmloZyVOoh7okgQL6ifHDs4CfhiK0li2HqhgHbpIIa400
3Mq6Cb69eFDjCFPYSaC68JiWBSe3iQdU64lyarOK4DCy78t/qH3QTkgYpP6NW4hK
fD3E4iUBOF4/dOtPhV5nhBTlmC8+MQkQmfxu5z4em/auHRqjrZdneRoNDl5FgMOt
+w24rblZv4uMy8qrP/t2gBKhaPPls9MH4hJZa7w/oGUkubic8gF1llzo7elBMSIf
gKyHbea74rFiC4DgGpy4bMfJLFI60EAFn0iP9VKx0de8Wnzc/tmiV0Upr8I6GiEX
Wb0ZZn2wLUmP9knwoOv3QJ3K2ZZ2OexndxtVvPxGSxMShVYj5O7Q61TVLq//acj3
IIrlCyrVHzMATvuRo9SsGjLOiZZP9ozyH6noYaxNdvNpNhpwyuabddfYAIrsA6Zv
4SSbPu2FGHqZN4TPqoMtuVVUnGvg/m7bLqGK5a0P679TtgfQKXLZNUJCVGxWrSeH
bryvTuNCvJh/5ACsILn8Bs/L6RduEA6wSQTTaK4KiEANPQK2YfKaITV2qnyImA1u
ngmFe1Isl+YQGdkWQQyWoqU94lyinqDLBugw2xVKeTlJxrf8eiVtOfsM8sSHaBTH
fIF+4Lo7JF6w7TOX5Xgzk9c5TbqxUajuL4N3gvx+glBvZ3NXxf6b30PK6NUap0S1
SgbBB8vkNH29dDyUSj8GDik471nm++2d8X8wVsbrmjQk293R/Ve96R5SIsNLOCtG
PXKrKNLR3ch50/swLyVs9foJdg4hXgJxe2kXUDYaEZoWKu8ipvsmtgEu5U1aNO7I
4YbQqUHHeOPRPaUxQXQ2QMp297B8K6F2ujDmy18gef/MbEn2tOS6Qs8j+M5WMpkd
7+UaA/TJ+MwiTj7ZfOUDrzwuLXoNL/VCISQ+bpwXe+GqPvm4RcqRNmQUuR+KH6qZ
qnZHCqfGxTEIqUb5AFbyfHKE0JbgwYvERatEOaEtJifFXd1dbivs1V8dqTdaVIKZ
EvAJhfGDgRIOYxYVvzDucRn4vJQZRhPXh8ZGxE/Z1ubd/EDsKfB0gGcHWqG0Ybgm
e6OQvagLMEtI6BGgzFgQtpDG5mDiDLDMVTWxfBG39yBBmMsSCbcvu3WudwK+k/ex
/CqJOz6VWqT7+puw3XMXpU6+z/jDQ0/DIc343eBVqedcnEbhhoDKHDHFsQsiJTlU
LddqKdiQG+b2XwUtvz6PShTd5VLynnYyUizCsd9AZgHnrbPv4yHveD6Bxn3lbyKV
EGHWqI4HdbNahV9JeFVU9lf6rOO5kPIfYF0QMf8KC1eNmSt5vFBnDGSKe073TBsF
z4VO1UqFzqB0DvyA70apCNeEQBZ5tO40ULDiibhVhAWqSn1R3s1YU22Hi9pinrIs
KmRbsXABseNK6BkAvI6cGwPrn1fD/Vzu6GZEZ7P7VrF7iwDi9+rmYkL+qwrUDyxR
r8GekGQxiFMwaK3YNIAs6WCfLPlF3AFXq2rJiLbPGI0bnHypUw6Zf1mMenQOQDgw
PYlDkJY1uhNlxvR2alH9p4/0dXb6bnNk5NTeC7YKY0IeoqihtaMd+n3q7ohj9Zbg
oWnY8ii35JThBWkocoXRkY5LPYTMgGgmJBPVBq5tM5Mgg34nNafdmdMztX9Oy6GQ
xS+o/geECvrO/XobgcO3dg+8WfhBaOPgt3hIQ8jsMm/caIFzJ/CvoKaDDEnVpu08
QVn+i5CHCIm5NqhksnmiISG7GDGI7GO+t3EOZ3ViHXKzkxVKo8oqsr+//B+p0/8+
lkNhOWrvIlLLlOtdlfupMhECLpDXjze3xMEK/ifFsREwQzLO535UXd8tHhQs5yhu
3yfhWtQtWu73vAEvs1uiwNoKydX2zVs/SSC/ALPbQdSEEMZwSviaXct8lqvfPUab
tyaDkz6ATC5brTqrXZBBSc0b3mXciIJJh2VFZ563zl2LHY5w3P5JqvETMCj9zhXm
9rgw0qtzOXwS4Kt4XLocHZ2FjCpkqZAWpMdrblkebxKEsLMYEMDfpih1oEkiRi1+
rHofSavSvLwnl83BloKLqhY1X9LDhH9SOEPvZI0BkQH9+yE9YpJ9INbfmHsBtANi
R+cuIXkMc1h1pJDPEhDM0RPzKHDSUY1bFOEOFRS3HQCI+mxZ7bXZzb/vWk8KdEuz
yK480fCNAKEIaOnN/K+sJDujika+mXlqkV2LdAZinhGrGGGfLvX8OF9gcD04vHK2
puG+JzEQaS0h+rcIKvPG+zIb0gYmlRqisLB7hGwrvyCijllbzlpYqET009XwPm1l
3bg89OOQ67WuHA2UGEPmAW8sLuqp8dvv8JOosB6demUh8+4ff4RipH/mUaSY76Xg
qKEkjx3UC9Q2PHeh2ef8/RaYqw4Q9vfAceTnH7umjRzHhbLb94wjoBqoS0YfXFAo
PMeIfVWD7ra03RkHbD0iHZX3/zNdMBF16EEEmu8NXKhpVhBj+gHoYLafgS96G4dl
ajaI5ITVnlwmMwku7fOHRRt4Al1M7ZM/YhWlFYt1gBNs9jaOF68ZSYTm+P/zJEgj
FD7LcxPmT4XAkxtM2vq1FH70xmDX3j6mGXbV8OOJL5vJkGaTHEsr3HITLGw2tE2l
GmTqn5aXgeE4KEzpD4sY4WhvKfS2jlp/s9AIQVcyHfkKDuhL1KBJnimJTo6wiiJS
e8TrKCsNROJfJifkSrqNZtjLH8XDYpozdZAN7lrzaRhG9Fi5V+tBufylk2MUhfwz
Vt68C2i2a4ukHXdNz7tXMpu5sa1V84w0ssZnX3t5ydPWyuiF2LLzbw+0V33Vu9Ok
sRILHMue2bTPY0GVaw2KiwTHO4t8NP7GBWnJZ4Gg+iW6uWSOfrba4cExcUhywxNh
gaZiJ0i22XhovjBGr/IIX8LYqIyBHmBeHnaDUru4u4+6X4bi75Zt4AKIz12VJjza
18KpeBpq13m19GA6q4UunNh+svT1H4qq0WqI72rSCiOLROJOK+TKPpxS1XU8ogi3
177u+H2/hYmsssz3Mr3QD35AAyFDe6oyXMHUfrZQBwE9hFaMLaashq63rUoZElUq
KMY6qWYkOA1XnKjwZmUhbXUiy0nAfXg/om07SnQtx1BKyIIr90H6outp7QZp5vtD
nmzFp9pdAFYZ5yEP3RRwczvYmOpCuZlR59FJUOoLGi9PmhiO4ke/rzr4dPgDSBII
0IgiUgUaaCc1UrJhtzK4UU2Tkf5qilCrgwtSTqa7JRbomIGyMPwVrE6Z5ZbdUiNi
f8soPvSbjxQfkNp2HPX/3rCWGkbwQrqCedLFqX8aviNQgk9UeqELev+ZbNXa6aPk
heKcGQtPQlOzQy5O4htVoD+kIPfyV+FOh6nezQVjQnMjiWdxXpNM2s4w4k/zsk82
FEPa8ygJScfh73SniJJ90K14KpycsF0JhaoXXqIPK8sR82GhrcHuiPmsblR0IKeY
4jZOHU3UPoDizRsNGfxZjEk3ntvj5leKi5X+wISmPnvxnnBTBR86yDf0/SBcUknv
SBMSxvGfaDKGZ4tz8ahnxZr9YewXur5qcqfcOZhO3ja61IZg4GUGwRf1IxFxPfq0
q8zjDG+JNX9OfSfggCO5DXJWqrJqA5XEZN46IJ2a/+1bnh6WgK7ukWhBlKbi3QrY
p24IrCLzU1brGh5LoQRpq0DebeVsULlPEzv38w+s0S0LGVMPDCgH04D9gh0jgxVS
A30SQjXzY7Op1/BJBVKvRWULNoP7IkcuZsGN7Xi0S7g38F1t3TYkF04pVdIcBb7R
uxepf6ppByl4oXIlKDc+2d3WZY6+i6YdGKx2ERNEVyTSFjuU6CjfZ8qdy4tmZd0f
0jYB4VjAesQLlD4zYMVWcfvaj7G+pFlMXNhssxBMPFP/ZM5BUpqmjtzZwJDmJWr5
2mdzTs0+on4TxpR50ZFfhTFum7IGCXwnHSDriIngP24sRTn0cqrocTlUaOKx2cHz
FmE1OMxGrgu4VQPJNMZ48RfjL4+HzUL+zkZKSvbL+NG/lLc2iy5/qWwnuoQBFuMw
vlh6DHVzDSZlmR0+GRWa7+Pd4QG2MEA48ymeDcpEJfkeCUXcU9XJIBqgJ6C7sPdf
Ya3keGH5qhrxMpvD9DCkdPFSRIn9cUMRHYfYsKD7k93qXfKCNdwvdATBg8KO7CSN
P9qGLhFfIo1cBdNMLtzg8CYr8ZsIke1iCRABbH0PpdCBsbMKZyydpfVR7Lj8pxff
cD+nCUmPfn5PjUcsXIDxdm8QsvypI+t657C4UM0kD8yK+i/C/Q7tTjqLvD3MQ5rQ
TcdEqMcNjw+mdhaMsR+JCmrEH9vfItKfAfEG8dSKX6muXk9lGU2lLEGuK7TzeVjq
4JVSNP3oUx8pDkW3fH/opYQonFhgzvYRVUqIBYLlk2ym1XjqWzRPaO9ciKMWVL/m
s9eQpT/WbG4xESbPePqluoC/IUx49KJoogQ/FEmn2VY3iA4fEG0akUBKwXohzFXU
qcLnRwThrpMM5yjMNVUlQzWC2CpCOhBM1QvZligFTKmLmtnNJ9dhiPhn94tXe20C
tdIaD9T+wZEtdwE9exwqM+zvabDcKdPARvVt+aF34zhEhD0okg51MkRk2THU+obr
tp0ZPc4k/tI1PIRUSVsV8AAoFdSq0jRjlVECTWmr6EZj1p8UioGl5p9ygQasZTuf
7DTVixm7jPeBVnIepE/UrMo7GX4ZVab8/1V/3/W9AFde877gSnIhb/jbeLSnE+3n
abPc979DfBAfET52oLrCSLY/t0451DVSI4jaXTX2sJ+i9shWJART+fR3wYoKr4Qk
wPxv52nQd8w3Hy8YCIZeVrAYIYm7HR70Ukecxyiw5y8a15IUp226ojbXG1o7ZI0p
IZ5AUk4voA2je/YpalHco0WLEkBwylGeKu3oH3G15grAc3TFXBzI/ClC3SRKdoST
hKYLeLsjjBbq14eUp5h4E7ys5gJa6su6NBRtcRIoffM3tH1+uWxFEiDb4lhrh9Bs
2UFcU1wJ24Hrt1zqYkna+AU+QZy54L2yxc8BEnPJQWH+MVpbNbWmLbImUPiN1sjj
r49290nu4cC2xbmFiGSpSj/uMSWi3PyxNquhdYEskXvDQsf3HuU6XO5q5pYkQZs1
mbYj6ZVOz5N697uuj/jUSPXHWpRWEtMSg+GnOv68mdah3V2q34aNVHnhmBYkXpC6
SDZw2fWSjDwrtnZcYr82KZFaMNqBTBftOuLYSaUVgZ8BeHs3k+ro1tW/6ci5sx6i
IhL8uJ8vjJ3/NdEHxrLNaPN+dSvF3ojhQgLsowWNzbYEof4mrtVHRwhSrdE1zORO
pSTP2rBkdMtCovl+gtQoUn2P3kGxSC3Wn1M9EREkgnMd24FrBcvHSGUy83k4D/mN
eWrJkJsj9WsNtDtu81aqVVJkiqCw8A1YRsu+ow+PJauHB23NnaPmpQO4AFrsffVV
2O5Z5EtMn8K5IMCbEUoCUAeKX9F69vBaP9R0S9WMzh6iJIXLAV5xiPK3tsZB0np1
aFC/wbFdEaNzkTdVJLj2LRYFfb3iKPZiPbwiJHz7ib05Mps0/10TYucOiC1nI+BE
s6+tEzaSFNL9rUva4/LpvUoeZoZl3jLTDhnyl3xfBA5tm5iKwz3Y+WCeSuYWDsdj
F0eK7n/GUUqztSH6tFCxazOHTQKZ0RaoHgroit+mU0bJhN2NfebzmFsutSU+fWXK
xrd+JWdlmy7ryjl3R6WchbK3SNxVZRsjZ2cJwlAKSvzm3e9kpgyJ6h0MWrbrRulv
/GqKXjZ5uuii5pwFT9AnEf0LSz+hI4jvUdcLBbEvDnIzpdmI4GZVuT7cYTyulgYL
xSpMbtKKvlsyHQ+TZSiLF4LxV1Trrbitf48QMtewexP7bJ4GOeNyvljg6CAcxceB
opZ/30Bogbe6cbpHtYzWZLxmAxZOaWkYVwaS2QISOfKQ+9W+Dj/mWEvwA5diMZlB
5KDlC0/yxR85ndhzIOOuEsbwgggdvYYRvU78KyMqat9n+G23BfxAQMXdl2qN3850
GfEoTy8yjYEpyBfEVCgnqo8frG7MxMBsQPkIG5OG/XepCaJ/7kQULcXtBqj1M/4H
Jf6OvEiRqRLp4bERiFboY94PS+FR9xo85ku90EBFfClbkkdVZwi72a+o1bzpvYz9
QJ5vvehv/iAf53mnezzh/POGjUwuNA1GJZCeU2jXDe+5dObJMFBXji3NMFj8KBg0
Cqn3VQIeaXZbb7NhxmNQHjtpOw+NdFZsKxIdRBdRyZcxVJbD57F79+vDJbUP15l/
fDA868YpgJdKi9lFzKGH62/3jTIRMGuu0xM0XSgfaufevcheBAnwRC1IAP96M/Hv
VjAjnKpjssJIo2Wfe/CXuDTQox/yt4JHkvXKRkz1a9T5ERZv3ZLXa2WS1VocMO+j
2NLQxaxq19/0uCbcdV+csovlqTANtkc6Xso1V8xOjj61q8Aqsh5BS+JMRGyoJrhz
229nLthvB0CLGxInpJjcQxA7wJr2hNbWGyzxzi2RdAVGpQIvOXIWE9gqGNhzxmaE
DMhhWns5Z4bYRPGbWRigtcRxdfehwYJ+4tlhFTJiuzLMjCG6E6ccmUjtzBV5xOew
TddSKdeQNTslU/j6Y5whRaqoHeIwy9GcGc3jV3h9J2DIefthlmzozxGFzu/0HFGA
22r/hvNbYfN4KUMApEXRfRe87FQgyFk07adVafZubHa14V6Y0F3aDaMcYV/Rx1kd
+IZ6Pc4sjJLMAMGHoP8II3olPesObWFhgngTqZVnVc1ZVOZ7tT0AbZaFJh8jRMnY
1NjTv78tMwVNoYtIQpUwyxqO4UAwWumhYonLR0jhqQONL62xhtOguBmhxeNqR/42
sSHu3cojx+wX65qoNcQNyCQrHy+Xq1NfB0lefPAmYNAd08BDI6oFDceFY2g+moQH
xDda8wv7sObxFkHkMZpmznA7RjQ3B9Fa6Z6bKkIc7LDGjgQhNb9Lv9PoirhnekDg
O73LpZfQoAepYR6fdoEnXBu4y/NUlTWUbRdzabg6lNyqilXyZK77p+neb/ycrLmT
m6Xnpn9Mu9E4sL4O0AsAHPho/f1Jw3RMzVqzmFBeSJ/2BAkaB6c2uxm3ZF+D/YZR
GRjO3MLpRv8dBawpzzGH04lFsRZQ49KYVe6uT9TaMJHfSfm3FX9qbapX/Ms+cdQ9
RiI17alIttooYUjb27bkZ+yTXPE/DF037GafHHLmrK/cWVAH/MHDvBfL0UavHOFk
WC0QKF/GxkTYaVhGlN0lWX15AeyvzE57FW/a6SdBlLHh/a0PP7MrroMjK8AIU9YD
Ah/7WLqt/9959N4TQtwwyhwAqpxfwVCithKt4keY8re3SanepsB/VkPYfzRQ8eio
Yagqo0O75FMoFmYKiTTVWrW36HG8OmssLllAfQn7EQu6nPTmwlp8cuqIo6heJk0Z
oHR69ldrS7cgk7D93YX070dlH7zo55UP+qkfMnS1uUiolX4qTw2I/kFl+1h2iJNk
DOHQDkcv60Z6f+sHdLvx7GIuzOvajEhI5zUKlRG2of4ozOFTfwfB0fE9a9H47dkx
tNUfDHJAzaISl2HMfbxSIo2QRcBhdzHyNSoeQNvz+hAgtLWB5S1d/w83peLLKoZ8
BpzBzla8ixZBc+AzJnL3YrezF9UyRLHoNfTGJoA1fXv91sUDZHQ8uJia9Oft3AH5
UgzuHzXQeOFfysQoIY9EYBIoyJtBZ0C1+xf3lWfmrIUh/m1LTLflqnW4jbFw+Bf5
LpU76560S1ipzl2Q/d+/Ub5icXlww6SMOtMZtLd/DltpempvBEtYUvJTnUThYZ2d
Wt0ZH/6EbAG6KZizeZO/9+j8bMDW4tIfFXNRKhVti8vMR/gJPBFbIa2APtaNOP3h
VkH7Q7tSwA0O24g34xkNtosD3P9GPWwpeG2G0GbksMo1Fdx6796UMZN9d6oxhtq8
haqqdIw01DteGEKD+lEil+bTeLuXchoqCWntMPLAMhnGzxPcKvcDM8UYy4r5qSMw
V/shbooM6+Swo5zoOMer4No+M2HXK9VVhsHQFi/iW7yByi8ZZaCVz/eBpjACzTKx
38SiYUOIjFRebu5ipI6ZLrzssLLFzEoa9GdLQOjBXONBeIYby6N75A4uN+H7YGZ6
+3c1YaYZCkK/9EntpTCMgOpfozcSQcQT/qEKlhlUI3DA6mTpsp/W5ixI7okxq7Df
qkVd3A9j0kcoxm2ST0iTVuB0E3Eu2DMEqNeiH9l4U5HY4V1GEhIDVrfGdUaIKmhl
sqAda+7Dkz7iuWApFZIvrne3GY4qmDEICLiGy8DyHoqzEqXFwE/R/tEPSBok7kY8
nIGRu5zisiYTIAMojaKXC6Ys+vLdAjZ/uQZgCzXBtG/VWzz1hdlgpthj9Zh0nkcZ
bAOHGQCOm0iaTcCAUT0ZkkEJOlKv/EopmAf5D/2Wf8Yo05rruvMNrA07Hq8iIDog
kkk7br2JFsCeqV5mAl270PDKNXeJtSLwVpBzoMiY0FycnOWGg+hNuv9ceAN8iVEd
k6Co0XltJJgejTEQBGD36ERv9MAWCYZTNgNIk54J15eBPvbui0a0PeUaSrxNmDKE
DW72eE48ezGysx38MVBT6QBQ6YeR1V1V+VIGw8gmsEZaw6egZJmsCbFe7piESv+N
7fqkfsFxOArZmmi4fEqWjNiJc7wD5xHqqE/UGeWBKjhrZSr8rTD0fydTRiDoCTU2
kBDgiKz1PxDiNzGaFKufF3FDxWCzmFgSv9DSEiGPpVdYNzmGkzsmXzbWtCW3Ly8i
vvAJVWoWskQkxjcJpQU/0Mm+pdVWOM7Wj8D4fhvs/IeIY1cXmQIaZtDkGMX/3eSz
hsB9NSXGCqtYflSlyQ+ZwklrF/ttui8ejUb/zabAd9MWF5yMXz16OxjK3T/A42dU
Q7FFiuv4DeEUg4y6OueR0oYK+SyMbWq5I3n+eJbLmQJnSfUqK4f83sosfiLETN5R
CVgjvUa5MgDsUxT/UcaNWP8YMIz+dBL1mWrULhR+tAhLTU9VOgcFtH4w9AbqKuGV
uQkmEmCNMBvTfMcd9X0EyHAO1FoB1LUuc5VRXdijXcPKH+XgUnjAFKeRaoDMEf/G
caXWYuFGTLIgWPpZxKXxMMpFAcNQqWeGV9Z94k7gf8aqclFNleEUTVCQxm8lCfxY
EDxay+Kk0cUQK362szz7VSfvNmfGpFv0uWLpMbtV2oNZ7ju1rDyXiHcgISUBmoQu
F2v4MoDo2X8IO654jstrZ1XE89Tj56IuPMNm87TZpwMinIA1EGC+Zhq2/GjyAsne
wE8VUJGSrHyj0UGPssPX28Z+Y3jF2ZbEQfwkg4myifyRLdzotk5wxAQ0scz3jdvL
03tRi573x9qTXruxB61FdU9d/jD3YTkQKbUFZNyP+K2PkKlE4I3Fx0myKt1nP/vf
wL3wObC62gXQdJ2qzmrCYeH6jWfFZ/yRY02OBTJv3ZH3UN5bYRKy21/naXNi9mS3
GAlHdkOedGKj2a78JPLh5Q2t9bVkVsv9qWcSdbqmIbOyiACw8r1OkiomjEC7+shT
p34qO1HH1T4Ma80RTTWfg7RrKil7kqEGTC2EMLCMtqgLizLZ2AfLFT4jhIq7qnjA
ypQ1E+XQJR9+DYSFSQovwgkNo4P4r3JDpoa7tx59rVgzdZgy9nXnyKv83DBNTn3d
B+aLmfW0jBMFMOQSQGTlhr6r5+aesZYJLVntsafVo8i7WiENKdiq51HQ97X2UY8I
f6Zl50zZDYxdPW8024mHvpD8kWuR2NPt0WpGEA4+2zLecakWw5Onh1LJOZ+KiTw0
HsjphhDL8BRf+J73Opx5xi1h6YPlYJc9Pu8swzOdVhU9CW/B4sJUeDMGzyAh2U0P
d0GRlDEVny+U4MMyCYIOVJAqVBeZKbTbmz3pSrw3KX9YXDuhCR2sO5nVwPNWnENd
kKoUXBTt2GErauWVpEmHfWFht1uZcEKixbyilcSCvo5B2Mt6j8dh3DdN0SkHviSA
YcgleRtT3q76nN6cNUW8sx9PdnCQ4QIi8la7jBKplSallmGFlWymC83oEQ5ecTac
vw2vs+Wgk0Ldg8yEwA41xyP1wuodPAl6hx6he7+DENGl237AXPX5purNu7m1Sazp
yUvMdIBTxPCPGIVsWHqZrqdqU9bFA/tIDq6xf/o/xHTPcTwiQYKgvqvylQp4ujFq
KUid/pZ/XOJrT7j4CPVl6qY7Qdd6+jyrYnw9H5lmsvLZulhgqFupfVIDlcIVY9bH
wOObKH5hRRKtiTBxcowS+CnMRyeMdvAqboVZVTUDCkxJ5Wh0qJQFGc+f56T5lons
TJ6tFSZIQMn/y6EX/EHm4vmVgL9zsvylLMzxSbUaHwTNmbom4W/i8sqIZXb+G69L
HkQD0oTvcpTa/i9zg1lKcwZj2zhPe0QDFkPZpHnf/dbD5U7x2vkNZRXtbPQ+P1IQ
SzXSteE8kUBhAVkNOUQ9ua0hvOQWe9BsLb326r2wKJoWYKvoo6f0EaVKtKUfA+G/
B1tA9EbcsgECzrc2PbHlovxMij/CrfHhDITv1gQ1N8dW+WWAuBH119uGEIZoeIm0
o8Di+ky4m8YawIEPBaWnkznqyhGt7q/W1/EZMb8lden4hRbdLPzuocmLcwT//dZu
k5xHCTcI9XIKgeg+LB6yVL2HBgamm03a2o5gemJ+esP47wpe9GPlXmx7p4FARf2o
vMUOWTIJmDYkMP0NQ0ntHBy+2XvRydVThdH7Ptf0RCKxUHx818hnKAbWw1Ww1JqY
4eRewwk+fOajcoJasMFqpcxRLgHNqI6ucYA7A77cCxu9ttE9BDN+fTQaIM+VtL8O
D8B+dz/bSCBez0uPfVxd8eRV1shcqh6UUdXQQNtNe+fW4JdPWmvGdX14RfPA3MMh
7bWJwPsM4zUeJxnbKLDK0GgJsSAcWuUkNHXaHZfhCsz8/MkSPDH6u4yvvXFfysC7
R2mAt3YRMB7+Z5cQI6oXghCvTwRsBS272yfSk1sEAppv5NLLSpH7FgiG9P1jHOzT
JJK0S8c9UsEMTBR1z+Di6lX2VSON20OBccHOgXLt1f87E2NEkD+3LVit0hs+VQmp
jWAwy/k1ZmO5VegEy9XaktNvxJRqskBYnCmjVCU4fWU43YvF6KRgU6FT59l1PKjy
hUuaMmhauQeaTKc8VMyklJqzuA9Dt7tQoRZ5iHBcK9gkTXchUAs8BgEtaJn1a/yW
n0hyKQcWBJAo1S9HJOLVNghiQTkrH5JppLOsBjRsMj5Pjlz3XU91METdUErufIxR
TSr8D7KlTna971wQiOIJx18f4lbCGKyT/IbdGyRugTsubdrKdU4Sj6UZR7kZCdKE
VZ5QCQorllmklA+d1mUi0z4i1ZgQUbDxEjaSLq7bEWJy5F3uMsbfgLlIM7Ab5qH2
ZPMUeN6TFHaWlOnlr7AZKdV7+xKDgpwRR1NpItBWHd5z9x9G0SgBYVjocYOM9fH+
e/7kso7yX27FjHYqdojpnq2TuoUHxpaWW6uVtkAHga0gzzjc/gMYIj4V4awhRGE2
MU3RAaX/R41tbGcidQaKzzUNKetiI2CEbTyIZwzJxEvii4TtETTRu4096iKqAJGl
Yf893+zVG9Hpas8r3gPYGlhbmQ4CAIwOST73ESAJXMJbIl+2pBPLScstR+JV1sht
s9ONPqG6jitOa9Dj3tl43wZ5QBz8NVxzwfcbugQrfYq2npFJsfjmOc8aYeXv+8vj
H98WHvKUsAK2aMFwBx7OZs8ij0ZuXvt8aCzbNWICqKIHxYlIFOzKDfhLZm3MTimP
Usg5rSi2F60xuSFHC4oL7iyXn+Zbk7olXbqMSicX0AvRP6/rtvpXjB2IqoYQ955y
802LscT8xVfOH2mlFFeXmeEI+xheZhh6LreUIAKT3d8ihKJyHAAxDca2BzRW7UK1
bjBzo46UqxO+jjF6BkFXjlXQhq7qaN2ioIlMqD/yezK+RD1cNH6CLCPr3xqXsraQ
jXWYL+cwrZjw4vdHs/sXJ4cgHZo9hnZ1wNbvFLvJa5fbJ/Rq2/W/9ToGcC/xGuXk
NiUeEduq578NDrFokhNqJDE6ViTqlX9n7IjRSoYVa04l4nKKnkPaedmm42RPwoxc
eclx/ZARoEe3QBFb9R8yOUkf8hsmrrf0ojqyMsdGdBGCCneSPvdbEJ0xEngGr9UR
/Pe7K3sA2cxA9C6qPIoPjtBqWdDop6PXIk4eXT79tb3SLr214qSy3TLpj0G5r/m7
p0eQKcoCnXMt6LDBZvoay+Uu5uo3Se+yAtShA4Ld8aMJWzAYpFUofEisjBw+Pc3O
fb/lPh0dzq6lWOi4+0CHE3mxkpr/06DzFF3pcqEN6CILKFfIzpdNCFr4c9hYd7gq
WwT9RB+FaYDh45Z1i8k1M2SVUMNCKagPUZHvrE/KBT90+nzE16s34wESG+/z9aOQ
traeGKpfzYM1+pLVfW0v61T2oKZ4BlZ009eBJUcNwdfov4d56T26jCtjPKBTz20z
ZOvQZag7pKOXjsqJe1nxe6AAb/BDXC3kbreC3IhjQ+SAeUxzxqTSzY8JEBEoT8er
VNAX/ZzTooaf1yzcqAib/SaglQyI1jIp2bDtUimQY0fJ0f1mBnFCtJnG2qcKmwyR
tmY7Kjxti04zZj7VmEyLoYTb51tsgPQzl/RpGLlKFGbIj3dCGXUJxb4rVDwt+5Wo
va3C4VEqPl6tNZ8ee8pluUyz9JxG7oL4uF9WmCE+Zvc389NlfLmhMMhOHuQqZpxX
E7Ob5x2LiT1Gk6lSbqaiZuT1/gtIUN21do2r1hTKE7eTshaitPP3DCmsDlgyZLRF
sMwXZvjCCUQYiuxkhGf0rV2F6Eh97V153m4E0+TU7yW/KZAM5TzorJl5lNlAW/m/
O/QeyWNhkm4JtML9NdF5pc4ipNRdOJSAC1q2Fs+CgQm5o2tblLIoIgQRSIQ1AZou
EjFYWS/Hvis1VmnzScnE1OU9ayPREb3iIjsQl1CL2BB4RZNTn1jRlDSun7XwJsHi
SBQLxvjpW+0aDzjxYHeb/4Ed1QgaGzmoG09AvdZIO/lkZ91WBDYxtqeLbLcXtZyD
EQm+QypcHA14TLzIzv3R3zqyeDeM9M3A5ruzb6oQX8nMhxLxU5k3dYolcDVd1kxd
vOQejeZZiejE4uylbMiMSPcdRfAbWts78Uyk33N6AgrBAeaP9gqrFZcCANUrQNSd
TisCOLY2V/IPSnSCzyzvav612qgDBq3UFu20xg2sSKHKNjrBLEE/5EETgoBSUQEQ
jPS4M+jGc2qwdVy9zUCbYKPbLiQxYdt2k9ll1jQIdpIRPILy9JtHM7H+abps6fZa
TKi7Iae2aLbtb8N9usfMfYTH2/wTKkGufSfuLaSwkN3d+q8msA4xTjCJGyQtMe10
bK5DZVazh7Mtuuueav3F+fG11thKFUC43f7c26H36XR3TB4cWAuCXUQMImTGq0EJ
Y3f1JnS1ffgq4vWqExZGsIUq2xElnARwjpuVk6w+9dSn+DQemvRKgI8kShmIN+cA
CvO7pKdNM/tAQ1lq5QcWydsOSrgLc/KzzFrHmPY+t4VrJPYzFoJfByd/Sw3cYOK7
zAS2smsdESZgJ15Wddt0QrGhyX1hSXus3K7ynUFxWyc7BXTyMhsoOCJTXIXMWLzB
u7QckxyUkeM0bW27y/rPpUqWDmxLclW4Pee3f4V34ZiW2zpA3DKO22pdON3IutOQ
kCoIyKsOnd/kZ/nNQMXMpvhZqoebjT7Nz6TV+5OH1rmCBUT+NiEG7teiUsFNsol+
ZVzxijOJjeHgqR+mDLC9XUJ//7TU/1Mh7h/Wopn5fNLepH5uIDMv+Rzg06GNs6cr
BfrFQr0aQfZdpmLpKJb6H5K9oGwpRC//hlGg8s/rtNhqO/dbbHiSka7zrSz4OaEe
uN/8uyXZbBUd4vXXfQIsY5020KlMQuDBRpkxS7NjymKsUQq+MSw9+ru3N/3zD725
uB2SRUZHESDKASgt1c/TnAgOBbP0bpn34U4uB9Mn07j6inhcZ3hlDNti6pbIFRzf
x0MRm3NYF+nNEgGJv5AjZDTigFz4IakMGdpRXVKfT/RxsvS82s9FtnT9sXtg9C7h
55dtHpBFLU4S12/5DgFf0LvJHc6IVwJ2FtHqNhh9+UaftTveup2Iq3ovRlx09DDw
ZRIY6zRRz/vEvWmXxfVOF2gxL81N/N6PTUkroUKiOa0o6IFtz5zTpeixyFmMV3R6
LfrscJzfj33WxUiWZvZrVICIQXaRLNeM9EPaPLorRDMfZsHilcK+udEJVN1aFTV/
m/D4TYDUA0ILHW2R8zHM6KeShxsvUjrM4dDZ3Iac1b4e9gZxor/dVazunlOSuBja
b7XTyVI2xF+G2d1eot4/DnHUlLU4goSaSLMVKEV3lrNo4OpUcB/b+K5ZNHJzZcMG
310RMmLAk3Nn/ubnXL8mYdGnaWarec9IBviS74oGqpRdmuIrPRk4NZ/8HVG5F4EQ
JDwtW9n6lQB9US7rMuyJx/PZABUmNKx1Qfw/bd4JhLvNN+e/0v3qDAi/JRmxeBpD
6FovOI8kE9zywBq95yF+hIhBf0UbR4WVdg4VYn+eR8n8u8CUpWaPG8LB8MVygC2S
wfvMc5a+1hA1gduN47hW/agIihTTAnjHU0xOXKSmVJbpWYD9U9QwkVCC9+lesi8M
RwQ2H73VXUTgEgGWhR7nY8If6UMa9H7w74BPCMdKoPV1h0nbLvgtFrzepLwAk2FL
7dmEEEHRfY6CLHqwjwnd2AMHDoq8/FPebI87IjuN/C3436RXF/56htIWH+kFK33F
8FV5Z85SLjWsugGv5kqqi5hrdxHOYobnLexWBuYq6zMzSTQjzvNGeoGyzkhsaLvD
h8eMCc9dx1XRDxmzXa3rOsUZHHdqJKjFCshiVv+QNlouP73uNxj0KtFAERzlMddw
rpQeX0AYH3pyENxEkuMZTKz86z3CxEAHLHayfz9sAnFZPOta1mUVP8oooJSX/w0J
TiPhmlLaBFTPt+uYhQFONzfLAx9TZNwTdV3AmgLMHiPvSZl/gysjCeu+cbVc2eLw
2KYoGIVjuGNP20sUR9H3pcjFsOMMRhaiWlpRj8d3PMKcM35+jknh6vtkA6EKOSUQ
OvoTToUcTFzOvYw0okc6OgygWdDFfV7M2AVemPYqrRR+dNcp5pLsy5rgwJt3BNf7
AGr9TRqL5lZ0uEkaZ5Rbm9ASHfGGsUUbTLOPj8S/GZvGKjJzbZK8BaLdHbSxdhTg
sfSuIYT//YTAlUaRTu/JhT6vjpbOdEi3MNAwPSsLQ0u74dBsNnFkn8vsIXuxJxgw
egfYrLCmtg6qWCP2CWGAXc/koFeLI/5PCAQqFphKbxtpYQFQuZJUct1PK7ckzsWq
+zwzDKaqgQpLxQkMfRbTTip+zNlQurIwYJYUa9QLw2FRVYbekHD+g3Elcm6P9TVj
2EybuIqY4AbxEuhxBHOzAlh9mHgbQUor3S2uR7RSv87eCnm5p5+G4zawXzDaK+nq
ey0d/cqNu09t1XvhrI0XdxJ4L8Ff5fCJELTxPV3RhCOZBKumDrn20ddt4eYxUIrV
LA4uhx/qHwN+8LrXB7X7yv2ZVXQsQM99IgQjaYVvpY4H3YV5GckkLjSx9/0UiFCa
+LJZSInCu6S2wku8uZUqWkxa52cc7p1mgB162BIxTtSd0+YM8O2IjCITKoneVkDI
q+VJZNHjJ8bZ2sUyabD4fkuput9gZj0U0Mrz9E+PpzfBZ7PiVd09vA+4Qf6dETXJ
mpwONq5Rq9KjMIZTPBGWbvAG026m5YVqih/QUmd68AaRpNUF4mqOCFbmuLono+Fk
DZU3/EZlbX0p6x9c7KX/XAzl65JRuUU+P/b2g3ewmsKYLmYx7zx/2axdFfbHbH0z
iniDOKtYUVXNWwIFqzFcXAxQCwvabwQ17dOAm9LQWoioM/Pk1Ytz7owXD2zj/VLe
MkaFY/iec8vFSUhpbMo1XvEsVA3p9jbWmRvXqAhdK1m062KHpO7X55xHEzimUp5G
7zzsom9skxawxmz47uboJoqT52dfjMfdiGf9l+SMxZgJYe0f2dUeTkKZrneO75dD
+t19/Z2zyb0knKRCVtD9THcnoZmJD87AJ8TMa5Xa00EVk5hs6kvGqm1dc2dm34ty
SIlkwMgRp8weHbRwNGohlRYTCgyK00gbaHFJow9O76jUS0d9aOxwlkm8Sap1VJE6
Nt6pJ0+O1pLIdodZDAkVNf03yCRmBPy34K/yTqrWpG22/63Amu3HqkMrPLjYXl+r
zGkf4LGRionWIfbJgNH3TfyqVqI4D/Ck1iwbKedp8lPo+RcDUQqdr7MW0iXfPIC/
M8xdq4Jvgvit+nLjELANtnYdmQw4xHItkz9oCVH42XM7gZxBg88IeyS3JkosBWFJ
3Rmw/y2YV09hNwDAqxPNfl2FHAI//RS/9Jn2o1VG8Naf/gTeiv3HEsmPmh4DH0Yq
gzsYWdgr1NkGuaHGKI2ZK6+GtoK2La1q7utuYx7Uh/tLUoB36Md+t96KGvZaYJx2
wZi2cbv0FdZHQ8gFUuPbRGzpYXJba3B02QQzTd/6mhKoQ0iKZVBVKNMCwRWMZfdD
3pEcBxl1YeJuMN2FUe7nSxyqymb5YIoQEhah2z+Vk91++W4k9tUtyrNix3NRk/Xu
YHjVY7dfhgajKh2QTvOTtwYab1Gq1wajQM5HkL1kbNj/LXXjHx7VomkQSZBbvK2m
yAgCkyH3sgbCUrXX+hrSUp5fhfh1TYu5YeSPTLGDr8lzfysMXHOBAl8Ph2+8S8x/
wMnNo9OtsYU1eR17E54IJ8/354XlwJw8yXLgu2j4SfCQg9BH7FDv1tauNSwhLY59
dHGzCIetycGiXWUGWi+fgWn8l9SqasX6BFqGtyb0v9xNhNTkSfcESuANWPCBSuA1
mUH2d423AvXxofvPoCrysjlWEVyutZssgzCjJZq7gxadE280FJ2OAvyI5emX7FY6
56oaP12bXq0vpJeqli/Tg1gdIxJnltg42iqvzZh7g4nYXIqVPuZxjPMZiZ2JwlKU
aa2pkSMzzr+jxiqwEZdA/sI3tKA7oumBVS41JTf+NvyKzzSYc63QKMuZVgIcR9gS
m/5a7zByDDPF7QjgMZsI6cbLlcQknSYOp1zMMdbfoY8fBEqt0l8YNg8hAWTfYpt7
S8Z5qV/NVKPiROoHe1vGXWXVZbMhJXFDVF376bwNqu6g9NE+sqRESoW4wfTp2Y9A
FQHIESK2iuQmTpilfQF2WDaclkHI2Qgv5MMaaawgSXul+HlWzALcl4R0w5m1WNCf
wPbui/50xlOU23N3thQoWux/w66SGvTZRAvIjNj8UfhU7Zc+vXbG2YZKEzgEbioo
8sWCnIEWsFiznk4kvzIfjP4n6iDgxWLi28ouiFxMRwoFLrrY72J75HV3hBqTgAcV
gM9BblhRMNEk7lxXsqGuTKoPQpizx4xjA/yRGMvuWBIQNjObWeFY86YtLef4txlS
QvavG8aBxA2dm7zyt26ovtXR5f+cIjoUC9XXU3hfm8C93ry8vgT71lG9OZiQVG/n
nsXGGDz7JEvdvHYLjOXXcTox09MDxr8UZlQChpeNmp1D4HdpTTBPcaXizwEOlTtL
NQGwvmh8n/B1ORbKleytFRz0IZbUUY/zJqC7uZAubWJdbuvTDOYjTAJ+b1+aYOIV
o9KGmRsfSSKcZUixXsFy2W+UKvTsGssOBDFiUfms6EjjaZzFfebosH2CNYz5whoj
XD6snpjITn4jtXkOHsmmF+UZHOXlViKlDU5jfiKtzfhad0wqiwDy+PpukrUKrAx6
drdZSAznDXNojGbNG/9/SjLIL95uu+3kWICY1kzojSvvVVOZVgQ54vIQXzN1eUD1
FC+uItPoPxfhUzogmUcEir249+YR5pKeiAbWrX0/d5PLVAsStopXoa3UcdBFTEZg
90oLwYUbBnG2WDmPkIpReqjqUHQ7R5XlPsnge7Eif1DtymByRt9i93B0PYP00IiJ
TUSCnKac+ZD6ujOWsu33UtBIjzHlvtqTq1q2dvAsDqKDw6YduC5fNphGBqrSeVp8
fNue/VWf0vRrerW3Bwh3BnZbvfqRs3bsYlKUQO2OngF6YQMlTFspOBRmloALvM6J
BjKwALaS4PnfcEH18trNKE45F+X2Z/JoAfvNyH3SyVGpftZtgB95cNsLQN0B4Fmo
77Lbvzwt0dDM43sXoD/5o4kQ0zM551kuj3jE/ZYOCsY+pFulFnAoGMQG3WUP7KXP
dbzj/QZD1KVV6veCFPXtdpr/uYiY5GQxWiN+20DweSTXbN56R0VnFdXUK7IadipG
EgMnKO8sSW2AXRKE37LSj2/eegl8umS1zFtTwIYi2sNTvTqzx5YHS1rw/7e5Kblb
1a0bJpvCKEBMQh5k+UhzklxHSSTbq9cJOmBnyn0TQKck2OQghc1Tym7BR22T9E++
Tw72nu9ej7yBc7H9RilEcAnnyTzb1joheFCZ/mMxjERyqCZRyr5qjsVofmi/Ze0a
S21irRSh55eufnJ2JEuqTAZaMeuysUYX1s2x1HIPhvwsl/eGS8q7fYF3/jiwH5vJ
OoKMttqw+U7v48V731qeOYyhTr1+WToYNJohKybV98Pzp7yh8C3TvLgBN+DbrBFM
24/xdBOV62FuigsPrgyvxkFIUPAoJHWtrh9BVG7/ISYYQKvNE9up5pZic4apw678
i3hEI4gTkj7nLnmi1qHM9b/Z9fp4xaE4pZY4y/QX8BB5+N4afAkymP+M1bkY735p
fvTzNAlomdVw/YOMPjtWqttIn2eDPfWTXsrp/oMd6twyIwOi0oc2I+LgnYEfambX
lkWcKOCztxtdmqbXxvSwnfFddCora1WH9sj7tftG+ADnIb07zJpMHXtT2KsXEBt+
6hyG+HOjPrIkeJC01vtxINXZ1df3XevPa4rwdKW4rFOObE/5MtV3h4mXjrlCpcHN
vh/N2BSwvE1vlVQ+w2EA2bAXgUHw67NiMGlhFX1Bgf+q90t4LhU/rwOkRjAQSvq4
2CZB18xog8sVSmTKb3OQAYlvOSYc6yZx6bny/kVDFXsG24ysBiIPzuH6t0uKVpQW
8y3GJZn2yCYRvZf6zDO9+lIuah+A49lD5PWiek/e918ujYXxAZLLEvOgP0KagyMk
Duon9TuaxjO9+sXBaqu+bhSsFjXUzp+8eN7J8eVbZJiB59MRDBJtuOuC5nwt6gf/
1HzzJd9Oz3xOqrhjjJKRuzrvnvjQZqDXN/n55BWqi7mLcfsIoNyTDd62GUG4l/y5
8zhuIR1hxeJeUqw3ousfPe3Tp0urBxGYrpXUA8nKNZzfsr5hMOXnpROWs3ltLWYR
GU9BMj+1C24HP1BMa5lqbZUQ9YwoEg2JIE5klbaDz0jtMKwLTvYPXuN2hHADUyM5
ZKFsR32CQ5q4j0d0toWVbHy9CVWbmXrRlZOwx1ZZvU71nC1jGm2EESdDLM6uLyei
r0bYla8XvLfi4F+ZT24SOiLuZfMfQ+u9YKnR7j7iTC2BRlHACc5GmEuK7Cq6Zf5j
SCewVxbG8UM0RlImga0bTxHapZxx046fHAGx3xsx+pKr1Nx/dmzxFJBGL8izXIIF
Pz0L6d3PtDjmzIrWp1q+9NYn63bzlHpbzlmnVvwj9U5wxvkQojRRXSRyTjFcJa8/
jqT7siR9mFiMIe68GfQJ9luWznjYc1YrqGGYUli5ufNNsQZ8pUKwS9B3UiJ22wI7
990dT20jKK34O7Z7x5XLouok6sHyvvYlaiHG/154cxqdal3FWvNDYPfvkJNgsUQB
okWysyZ5aOTv2y2AY1Oq1q1kOczyAXmbl5eLo3TmYXWqIbfKFdT/Pz0x8Z0e1On6
ydg4guWv0/NIqmpwzKWSzUEyTsUovtxiAmblBtO8i1lD2cJux4AHiJGX+ytvQYo1
xqgAAIwT03iK6/760IzLfGRHgoShU57I1IMNqs0e+IR/s1C7e9sB3DfwaiFxpoLA
vYAd/40rSygh1EI16FnV6N+dA+4ZqjiKTTydSR6Usoe/sHZ2iW5XEwli6jGGP/gk
gL5ubiwtALCGmdT7lIVp+KxkkfpphOxasbSwx+UjfOzpibQLFVViRV5ARi9evN7j
rFZQC+COGFjigoSKbrRh/8BxU/JnhZWXLkDfun3aY01ZKQpwPCzCnW5iwumxhZR8
Ihz1jLEYCikEYE0zFgvCfDdrk7L6vg06ZdiLg6bN4MtiZyXjrUf5biVWgf3IWD+a
T3V6gzGFCitKdjufAEudtZNorL7nDSV6KKyf0AraOncaYDwAkQM/iYhZYDQy3sca
N9Qn6bx2+ECzqKdfK5Rnmn6z6cs3I9pqt2BDpcFW+RkyXT7teoBtxBL+QS2mPkoR
pvfsjD9LsqBHzkCKYBexnBGyRayL7Vt22w3vtzsQdN6H0YlsbGW7hOVLxgg2E/7Y
mancjWVYdlxrGakm8Dr39db9O0hg14Y1GFvj+EuV48rhn+te2n5JkaMGcJ7/5eBv
QyH2o/eaUBlBWF+yjd2tMy5TjYoY/pmPHoP1BvG3Hg4gutqyrhXiQmk/jk8lD34h
+kPMuacHzTBkX3l8l4d1RHsqITcS4Z7E1zqcJZclIA8DwCQUc/TWnP86tNFj2ZvR
ZYd/n1MOJtRcMFCrt19qe14jeLqgRQpgvbiN2HvEQo0eh8IlC1ohOjsOGaRwXKse
RYZGw91/zGuqbtnUVZEKyzypXMR1pvpRoMIkuqo6w9kAiPBurIhvzifWx2zEZAyy
cqak4kkUqgZkklTU06EwJU/uBgOB9at8KmgOIjwTxdB9jP5Y0MkCZBuxqGfZU0kL
bPmPc6BhkaYziEfMSm6RlTlRh0EbEwJsOBbB5yAoQy28wu15cHz+fxu3k/jBM3RM
lDn36ji9hmzz/qMlQcSI4kC1XUUYEGuJNikAdPaOhr+zSXCL+8VTt3zfrdkOZOlm
Tq9zLjzNtEE7p2gjmBgxJ8ZUwHPIBx8hOSsmJhamYBTReChmbwbgcV1dCtp8Og51
cO1wo24GxlC0DGshsg5tsmhI93jfTJdeXt18UcuPgr4qKk5WKIdMfJErGyuENyHm
qrh7d2nknC8SXhqT77TX31kN10FDfmVfJdofRz5o5ICPdH0nnvmztweht6PAk+g/
J2CICKsHaCVx8VbAU6Wfs+X6DdJJZjXFOSjxbSmgeXVnxmEDi+q8V3RlMacKSJe+
oyFUKv0RoJk+UXhHZkdIb/e6sOztvxm7iRLyglOaysMItwysgIU1AzqENwdyv2Mi
SAhDM8RZV0iq1cyVGlriYHuvaTSleuQOvwXBi0yHgc+1CuUKkz0VVzGr/+JsVe++
g2B0pV5w0QAIv5zrrn+MYhEAMbpOc1ssoNSSj5zJg/F09KCKSG34Mz3j75iqN3py
QX4WA+M6jzELPwSfA1QB0cWnosBteCc9M8mxUoiqId2+UqGHmgD+fWbgVq6oIs9K
Zs9m7nUKgnGT9F09FfYs9EHO7FiKVWWB16vfP+ZRq/+9tpqp8X4hTi8ADL4zzWBP
3reXKHPJsLsj4tIcaN0JjGYy/m7XOWKVGLa3OJ5Ub9FZVpbwSLCycD7MrqbhnbvU
oBt839av+GASDY1Jw6+jNRcuDBPsqtADogr/XVFKFYe3EShramSxGBpxivM/7e5W
uBruQkHqKXaXcsl3sfcq+x9pke+pldUW+NtfmFuW9LYeaAEjE3VWO8zl72cvUqbH
UZJLQ6f7x0CXEqJnD6oTnQnkgvdKDQoWrZEc0LSWw7vaR6G22YN9+PQd/YEpaRfY
5tqtLD6Ad0Nmb9QdubRGMRe2pIX45S8laL59qmWpFCKGZJDlDiWF0/UE9K4rvKXs
TV+KrZFgJHmsQeou5Bn+6DP5p83MGhs0i7ZH9raNyfiDYpVyWv895w4Qdaw7Axrz
0lczIhr8lCZ8YeIpkrD6teXaN7NUGZRUmyNoFatFqBB3Na1YorPG9l986SF7aeoU
JCUciM+EcSXegNQiMslq1Ch9dyf2jEm2phxDIBGSrOEi4AJztgm+LBk9gw9uGztk
NHhsTpPOU48eMQ3MFqqa2SKsej8wLabo/EYfoPMygaDXcm55XJbXajPiyO1PTxf9
S5/eCPTFEpW4HEwzQryfUci/D92WmyhjcMcm4JyxbBXSburr+YEmCVr3jvXm2UE2
+fAeaxxE/0CO4w74j77AIDMWwAdAL3WnYgNjAVe0KIWaHpmQULqQsCiNkxqfOiUq
pTNAdCPGJGWAPaCmVd8JcW0dnHYkgxYpOMNeS6GYwnelHU0zKjc00JBrfCdh44Fi
iZVE1lw9WbCqabqbgEYWaShn6Ev6P2B2HTo6qIA4v8+bZIv+fWzSme/yqMxCXtx7
Ig3zvOjimOx1df8L0y+/hisW5QqWyXa80X9gUyHEcja6cKb81xcid6WBG8s6Ou6g
g3W2Pb12CrPzW8c+HTZkIWhMF2kdVaX1ZjTYJ4ynq7rRhEEdRwfKIIOQ2kl+abem
m+bD6eXMMVFGzzxo3yE8oxh5HIciibCZYZ2YLKTQo2/dmcgYz/Xo5cQuGwHWAKDl
bXaExCJyy02yThbhQvgAP4AsRIR1nIxhd7AW/QByzjrNBE6WSCd59tbqyGz0VChJ
1Shto1SnCo/m4NEMoMwIPeTMbDh8xSzUuIdcMaGtYyiu9fh4AGAxkP7mUHsUvh3b
nJ9o2/u97AGHfYzsg1Fy+NQKgjm9+ThyzODpXDs4BDmRNjvc+yC5FnFqf9KMgN0p
Y5UhbJ+DNetZPqY67MicWleLzvm5v3M0Ij3GY91pniveMlwzGL8ICUn8reYGRqXF
i0i5WGr7fvaJOloTwcqZKZgqkjNMpxoH1Bxc+rpeGgifzALZQyTd5kYugZCSXJ5d
D7bfR0oknptaKVW46ETWNmuaM1vYUpek+8BbwIWAgWSgYyehavxTSr9JxzwuJLRk
uvf/KUvVRq/++XPkFeEn27xZsdPDqxbuJBkBi711fUe32hE255n0n+d4AVqZzD6+
KI3Z/tlVgml1xHs2dO7bO7Eva1TNO421CQD+2wjwZhYFyTRq0u4K+6Lo+2nZNZvD
cz+MrttBde59s/JtwsQIxzWfsJRC06mXW3ycoUK6S+Y8BIpYYDZZbr40wkJvqfB9
NhYHJI7o6jKUka7Wwmea1VG5KUbUNE1Q8FkzE3d5Wj97I36Y/jNcQ//LDSvU5lTU
7tXsUBhM+PGLJrQz6iOiPcykVeCbAfaIU3KVjN4+fef2ybHpQ74sgtLXSum4GBTa
x3i5GBMawzB389MeAMEJW9LmPR2BOpjFvCsWCWOCfAKoqSw/rXPjMh/aZkYg9Ra8
bNU5FeK4Gv0fN5S7eqrYoh3JPrrnj3in+OIpu05rn6wnTy1nUAtc4U12vbwkOlKD
09Y1Rr3EBwzpzXy0V8puoxw2lp78t4ZZcOopt/dESATrIn3MRURGnCvszFOnKvEZ
P42koVBAf/03t223XUm1nMgt5f7mirrS1QhoWpk8PJpoiqx5rn0kSWSP6pPkl2f9
M2/3G/SLpxFbl3Y59J7gyK9z50UiaY/1jWy6vgT8hEkuz+lGtlGLTs15d9qHzqdy
D0NGbIgjmfQbMTGB8Ee7e/6jwTaTQUGGd31ekGj3oYWNEj4cgU2JAOBWiQ3TOLV9
xLSvLqQX92jk5ZP0C+qRyuey3fjkFcWixOzztrcATr1qLcD9sWVdWvDZYNBU1eIl
5fq8LcqJNrNKymy82+bsCny/WpPdlqJYhniJKF28OS4bz7mIFUAKklQww5Qc0mxs
RC8GFsfYRz2QV3eYPAXGsBPAy2M0ch4CT1cfbrIMHeK2gWn3BHZGmv8/O5oj3oqE
PGVp2tXzYnyv8wkOSO2f5kw1UL+KP82s1vTqc7siygajpb4Tv6jSrQpfH4Ao/vud
PopTW3yexnuV+8eGRrgSv76s73B5RgCIZW9NUYIkKOTjQ12CWZuiV2yYZ1BF2HfO
WjMuMOWeL8CxodBVZQ6x9sy9b/AsvjWSWStJqR5+hqaAWei9c+7/30vXWVjY8qHz
9g3UUkw7oBMUB1tAnht8uzTRxhd9oOizW7yeobYcDA5EOC6brhVOysjlu5USkw42
QX9QAoXzWdm48PWNZG+r2CBBV1V8KTsHdSY+LDNo3olGbHJ3693/PK/7IGOWE8mp
WrwZ6JENciMAwg8j9xJdS2kTo0Tzomio68o8n/vR9R3T4DxiPUA+vYc/QITZlUJY
XVpEspxFDTZyEFiKW8sHRRvAjEnk2hHwl1QKOcw6/4uf3FfrnSyMd9jJMDv4XPjZ
IGgC13MnNCkG8Wy+HaqkxmFNXXbA6sYOjRCAuQvHnHoTfwZX7L7P7OLRql9NESpv
tXCNnSW1mJJNaBfSDpb6pJAb43Iy28U1xRKo/OgWddWoPibQnJeDyIv+Nu2He7gA
15oImfza0PlMhWYtqb81AmLP9yniVRDIyR1/ZDQpi9BFr8Vx3W6bCeTHTCwJ6yS2
B5nauYU3QOzLfwBy/eTjO0fU5PqLLH4cUZyaJa/ENa8t+fltEvx6C6O12P7OLq3K
6GhL3os0LFbmbIKDqRI2wCN4ipyIFg/XGF/zsZCVRcS+lPSL8oKWW6j9s1OBRP9A
GAdnOvO18BZrvFQs5mYYCjvLRRgcCYzOETNKvmw4ocIFRJHv673Cd0xMC9UKxB3c
YUZyJbXPinLMLUQGWXLBR1O5pAQnTSxomjzYUtcM80fwTS5vkGrUY00K9JVwjqT/
nlZ9HnPNI5XbawduemMzOoGVDx+iPTjHht7K2TqfgDWo8L64rbJ6DJqQ84Pkjknr
FfZVobnEIy02eX9owdWTsiiuuEoAIL5AmtKzley8BPa4sYB21piky8kOr+XHjPl6
AESecVuuzu8tC5kLUPiORdt1bHi8Bk8qJ8uvsjvS7dKVMvlXx8LnRAMeIwUwXJDv
hNJtfW0NZiLf40bi6UqjdNTjO+o0OtBGE7GUrRPGuxOyC5Qrhr4ci2s8awklLyqy
lo5byOFJ7C3vvcgZUynUNDQvheP6pWHtxCmjzpN7l8ZWihbH5Wwk0c+EZQIb5sN1
XfgMJxF6JjITqJG36K8+vJcGbWwXI36mAEbRsPmAm6r3V4Gb3ujK9R3ibneKP5YS
KdsWv95iSSRKOym2aWD7Q9BfvStCWy1DZJ/fwqkeJZ9svT5kgH3aP2mT91wtaTyL
tTlEu4A7YV3IBc3QTht2vcy00lbHjjcZ/eI76TpV4JEOnEiZ19dIAd665mT68SCm
MRbvrkoVgFZ9PvpKkMuFuGZ0Ac5eHi7vkbMol3DyLQxfSia+chUw6ujQK8EI+aCP
KOBt+uLYnarHHYA/XOatyGLSaSAD5RrGl2ecwg8lTzbmce8WWtGfS5V4vcch4bd8
uD8kyKMLSl6hg7Tzt65Upr5hyaA4n1ZEqU24Zh2TcG8XfsL0Tjizd8aoiTYAO70b
vQLHLW1BCNQy2wQIer5tpv5+rZuDOetqA9nfFJwS0aKytSE7fJMtMFbSK0eR0ZNT
kEFAEd+wkrfc6LuQLmlsS2vBW4rN2lLlgj9N6JHvgPE4N+Wf6K4la+zgqMjuGx8P
e11HwRT9qMWAqI6cq3SLJkN70r5G09NqKfQW7YuLoEU/GeMlXFi4SeqwlkBGP9eg
KSi2GgGCbkOlMojcjFXHNl7RXSdj0rD1ET/w/77V46WVDdvgVUg+kAPsUd8uUEXj
LaurNd7LnvJBtg8+CXuHr+w0BX28rjW+1m2CPUkX+FLFPPfPQRShLNXjXB1I6AXs
tUwayHn5rwTh1SxzJDjnR/7YanYfhB2m5SvWLhhVm+JlbC/loDI7Pq3OaXNoYSqV
rIfpSmN0DfnWETFrOI5LRqXHawuY+m6Fzbb6mbwzelyg0RJCfoHJSvjna2qWhRNF
fUsSI0ZhTlJ/mpNvJAoFvjkSQQtNzc2foZoGui95a1p/S2LsPbjGj8EfYXrTXgyt
RWg8V1FWyepNgaxBUtAIvCr7wPA4T4+8DTerdyGDCUcbzPY/PbB5XZrQsequ4MQS
CV8TRLfJjowNWIEj6EjCnLfqt4pu1090YUI+jtVO1+86Lvz//MA8Bp44Lc7OskfB
thh6PWgCFBktde8XttMBRDkW5y2NSOXKzpTo+LEO3IIleUwAzYL0/bATaNmfe/Ok
9HoVzHWIM4m0nvzMg3AL8jZHqMPsWwscONDV16T/taXvLzvFH5ji440JaSwi9J0y
LSKfnd3BSlBW0bvPVD1uXTlyV3QMaz7UM3joBPwCGvFWs+vs2qQPF3+bbnz2yEv6
xcXWKylucSKsiNkAYxYzyNIV8+EZldEULno2yx9yiWAmk9x9s3eUNKVPtMXEXnAh
vVIqhpTryjJbx/AYUuNdZ75bCe2elknFDKmFbEPe+RSDggShhA2gILr5bZnlmiTn
i3eZosXUoSG3w4Q65RtJGpvXW0ToHgT1Yh8MJ18dKTUYDoziMOga0xpP5/+EUwBQ
dd8DfKURejrAviQP0wJ/K5rUX027ApBvGNYWdFbVs1+Z2hrwxScYSDj+Xg/GmxKJ
smh6GYoE80V92bG+IfO2Pg6UvNElS/O+w6TqBt1FoqfPCkZBUEtqO6eb49ZLgGvS
U0MypfcaIHY88kpdops663gykzgLqo3u+Wz2dgXxD53+lZykJ2K5ioYK2+M1HsSr
6LoGQ67yy21l7pYqnJ2mjSX8vCXkEz2qPDPEaVkqzx7YTeNQNOx2gfCE4joZ6ZU1
HNG+x9S1iyuvPtgSIVi1GxJKrdI8mvod+ubHfnmDQPHQA8DmARE6TOKemID1pNfG
QV8aBcGGyPs6g8dggiB0HNFKHswj0Q19F1Q41OCM2Wtd+fhNLZR7D5qqkAhBM1hY
gG3NkptGG5RA1zJ79h0qXR+CdF3ksV2q2y2zouTcQw01z4cTpFfSLyr1564jNM5v
AYJJcl2qn+rplPSxYNFMXcoLfm91o+K3O6l8Y3KSNmXHThr1amwe2cxVNTsdJvIS
kPa/MV/GAku4blmgoSmAk6H6frOK9jgVN/bDb3/isp8i3mv/ceUBhi7MmVTc/yE0
sWHWdt9A9fORTw+3as/sHgD9zaMexh/L4kzj2Yuv0l6IFAJ2xYJS2u4ObURuqIVA
j+KijyXXGMW0x+WinFlTftq1apcOqZKLDEYSqPREuSGMaf1YmX6Ihrg7zZzM55X8
OHpFH1a1N3jcgBariOqZSemW0Q/+5oQmRN5Z7NuptKpqfDuL+i+HWXk1Jnj0QO+Z
ZD99nGE4ZCGyIFUhxJweHJLG5X+yRMdDDlPhJbddcss3Fq9/B4Q+lMeQXHzrdjaa
xTfEH5UQIclwnbwvytO3OVfVOa3sdkHA5sZx44Dknd2AUBi6PAOf5zLfXfghTzNM
kGw9A1jHUQG8AjHwBK/gpRagelIJCYGJMrfI2P4SMxz66GrmG7k9UC75BL9SrnqW
qkMPCwkfHu0DDw2KBCkFc0xaGw/crqFqzaf+GFaVu7rFWwqNTOlxg2EDvBJnzY5M
zT9g3yEsPIPgjQuvvyeOtSj7iXz99KkXX1oe0SmjNLjbpgD43BJxFBbfxP3gZ8sG
WKbVxIDLwYJwcrsFx1a+QZAbjCDB+PJtc0Ydd+09WRYWcVoLNMJCPVlNSBffj6s2
uiQbKh6m6ro5/isOAgcfZRH0kkotf22BRcxhMcmnnQQ2HQZYVxJvOGMpVtvkdnU2
LTJLNZKLbVAKIQPwlUURdGNH+lc5HGCjU8vNct6oImPPMbFsnxVF2wiPJ6HLVIgH
Vqh51qwJXq/juVRmxWTxOV4O3lNkzKffwQnvoSTvIrZM6gmWr3GUK0tF9p3gpWQ2
qmCxVrSwe9ifMaeosPTCF3V0LDpPCvB8xjfNOGlqT1C6XmlJjx6ARCW5Eooa+FNC
hn5uSiNLYRHHBqMZ5jjbd8EamTDNCcyP7sB8y1EeDPm+fY+wv67JIiYgyVB5+yxv
lRXuPaqgRWSvX/KhloTyrfbVIrooCoHMG1M8ah40jXX3d+EOZON6g+dKGA9CJCUw
75EbmTNxrWEzsOLPTGLSA3EXZ8eMgBUlGNLD5+RDLs+8ML8J1YHXTii8yYUJ7xtK
JKO0Gn9LW7ogjzgNxcpDFZsYzTB496OQh87pO9GtDFDBG6Jf9bdv0NFRcVeItxzr
1nInK0TUIcb7uoMK2Hen6OwC7CmrvI0fpw9yUTGawAufpgzA1EbXu1TWB+AZ0clL
Petih1SvhI0QDWL6XPk0Y2sLeBVdt5ihXrT4NbBMR4hDMR21xIauOYV40KAOtbGI
f9oK58UU91h2E29XSK41QfE4mjkaYPkHCZXAJMRh4C/Fv8Bz8tdV9cH+Fop+XH+3
bvVV7yrgeMZBgTHhfLfpRGRw3uS98nV/uNT6rDNZefzJjDp5LuvRtQoA0QiW6hN2
u6HFk0dTWbHU0VpFJyuUW99wGtFblhhjOnsCbHAvQE4PSfp773le2/qu/hLhMZRK
z2EhLPewdQt975Xurvu9fVgCIFOrwdWkpY1UO8iOZyVTun+FHzN2LzJ8fY3q9bHX
qiQ7KiIEIBTWV9gYlWD5cnypUlMktXlC7x0na+OpCLv2D9lUbOD+j4Ha9sEOzWHR
lxM2YbiYqFFYofzMguEG+gH3LyTeGYm1jLdJ452kk0CDxeJJkGHL58WEnRD/sJSg
HUwihRgqNFs0w+adtwvR9hsPLYy8XRsvzwHyqFecCaOdJqnvqiwWqhC6Rxbfe9L2
lwsqmG/qJK89FGOXg5/pQoKQm2ETSWH8ayAZyib1OuGY2qQ5PPx8mjTobHDQBFFY
VUrocNFYgZWLy8As2DCxNKcJZhpOn8vSUbEnufQmDaslVFvp3DXTSReCfL6tdF+k
qy+Ax+FmLLgGKf51NFbxknf56kAtu6K6Zsi1rVH7SlfuPFa+IsVIzSVWWaf2L1/9
TiUcw8N5PuLITW4Rq5j5cUJ6OufWWTLhfQ+lBOd9RN7jBNsMztWwpdw3si98fRSI
yg7v9NGNTL4TkmDVnULLBjKkoC37ckYPCS1evndXw6zR5TIC6UdEofeATiAr7Wff
OwRqLxanbdGBintJnR1R87IaUOv+PEZkOA0FDWsj3pJtsTDa2BQmXCe8qiR4jzKo
D1GzxJCCIYoI/+5NVSVCQdjEYux15y4KzqyrVCcBjf8G7q7lBYRulsY9cFMTub3w
KQ0EPHHijV9LihJZf3WkyYhSXOw+e4LZSU/gI/0CrbMTyVcE0EpFZxhGSerkHoVU
kZJAPpLtkahftj1Bf1XS0AYo1NZXoPBc5Eei35M9FZQJM1OvYpLNDHsjH5gVg+GY
/hG7wxSTrJqOU4I8dXXZMUu+We20GD2yPi0siAahSzn8/fZmyPil40novPU3pcjF
NeXDy+Hmh+pTE7QIaWEWUXX/4n6KSdBsXoJEhYX2JGCv04MKv/ypICn/UcYt8SVy
y5AYIkGKYw+GCbxLoeoIO35EYQ+V/raTEK3q5bo5p2vVv79nMYyzVGcP2sKeA1lP
NMxR2/ujhdY6apSnI3+aLJlNqEsmNckK5H7NzruEdDlC2erPm2XSyirdCBl1YTy4
MP5u4PhuJYHdVdmtirhoRpurAJp90GH0mwci6chcCXVFH2Me0qJmtjDP4CTVvlaa
cPmti9lL1rzUMiPsLz4CSqBo+CctdN9uWTDxD6io8tiQbyRCL2yENgFMB8VBOWO9
6mpjLD0XBOuLlEc5Vi3zTEF9RGiXX/NvbmwCOZNaqvp2guLJ4v9DRw3GU2L9alHd
3esCWll8RuNSnJndbO6LOdbO1HFE6BIA/TaI3gdXgeuH2c/UMs4AVzmNFK29YPz+
kCAfCpsXKmGpoYBDyMtsYJzfocgyL7ktZgrwtNyKJo0Cyn9auSuCQSCtZTMAE3AQ
9EKBsraSE0ixxlobZTttxJ4Wlo1sDYgLWr7i0Vlr+j3Al8bVGnEagkouF86hRYre
qAUmOc4/ifcmrVur8BeC9f/9kXW+V6R50ai0mGIxFFsOedbukbztR5rKqtZNlEP7
+gUQ2+o0DdC+0jtYA4SP6RTs6po2uewn13m+zLSDZsnpCm/cWFRiCFRyum0Cufxd
6/5BD6C+4xhONJLz/Xsp3iW/htnMtRRBAvpaEHNu2tYy1IrBtpX9wr2gSfHLDNsT
Y65CYSLN9Ej2qd7tO9ym0ZuL49UYaGGnIZVUk9u+bLvo6vg5QuXHeCl8KdoK+Nq6
asgJX2S0Djf0rxMi5PPEH18v1GppKwWehnrszWwIGDhToNcs3jreaNCFB52ty5Js
s+mnPRF/WvUF17SDaGBs3E8DNg5Nhmw1k7VWchHcLgeqfSUTD5wsV7ylscyZp3su
ks9t+ymciHa25zLwYO9PJK3Eum59zwW5wmk3NM2XTE6koWGm/g4bI6B9tKhFvXb3
+y6COP9JcwYngxZL3hsjgiGu5A6tIeJh5gvVqdavQ6hr4SmuhNad0YWt7opdQVjP
qfvD4V1QlQVLj1QikmEAAD0x9Y3GvR4aljdhztberqaR09b6xf9QJpIibdMTjFz5
sDYZDLPhGrBuOxynff0ZAcnqoF06JONSKeEYgoQw7vY9MOSAuccsTwSDK6pbfEEX
TZqNAZMzoUednyVAfe/VqXLXh/y+Z8yROXAXCt+3J1uOplZX6CgnAwfVtr8ax3rR
XcHhO1WiJyyvtNJKz7zmG0QYBbzKhskJHE08HDqPMV52AqnS6KgYFUuBVx7g5tfE
oKuW49+4YC3j159M5pbBzdFT6DNZsnmRkZK0iBYgH0nDx4LfXEKdkzDFeKgX05GW
KRzd4x5tA/SzfSnBoFgyezwuWuV7YC4z0fGqAuqno6qjtuRlE7GCpSD/1lRu8KCA
rghn9qTlPZzNKoTG8PQsTRVQawI2Ix5GdB8BhYk4nZB5ZGD70dYE8Us87xDGQK7w
rFkIpx4zgM7K+z0ELq18Rcp3aG3zDliW7TxRLDH9uL0tXmi+uI3OoWFopHK150Qp
RdKapKVG4yiu39q45AV0pYbSeB4++ISuDPBUrE5m9QU1k3Ig41R4uxIkv0sNNCFf
/HVZwzmAAPBRVaH3G9FnixAl4P8PD7dHjqc4WrQ1OdvdpW7d3w64be+FrqBZW9qq
e9QSGZKH9VGQJW3nxeUV1/kQEmQiyQSrhsIC7JIkMgPlxgnjO0xLucszaf1a4jaW
iZcK7aa8XMEpvLgbltOIgvpexuTA/a/MEhkZI8AaLLofHKPE2IA70V6S7yVZlmhc
Zyr6FFUMcZT8mepFHmilVaMP4hUa+acDNUZPqvyyXIyouLhGpUQIA/xKt7Lvydf+
uT4ZMPiH2yGlxYo7WdCCjHGeF9ZS/kyeQQV0m6B5GB7FFS8UeF10YFWTNjy6wAMw
fm1hapk/7lpCxbHZqHwui3CIySBlajRybdYSrEVp2KVjCZ/PYiQ6y8dwGTh0jWpM
5wLQUTbp6WvEIcC2ko03bNY1lUYBMVHIeTFNX3FEiX9W4ohQ0SfBw5NnnhNDGDvC
EISCclLgQgU0l84eQY1IauMXm3l0RvJm3S2SzSdbgIAcyNieIHymex30aii03CPn
4ik3EADp2HPYmb9ViyeykY0sQGbFoejcFvW0++C7jH6B0MH6VVtdtffYbahnx+a/
Oflm+25NOGfF81/LywCdYiA7KJwmUgrzu5DWndobGao2bRqehQjnSLOgDdHU8nPr
QeQmUBdI6GyGfLkUmhXIgCiQJQOc+WHxRcwd7+3IRLfwYIKQ65vEddafBY08plQv
pO1dXuHCh/SH3EDLkzS56J0gHAxvcP9rL2KESoQfkcnyhvxX09J6VbQW/U6aMUiW
tJkkOOP67wQZMgbU1wOPHFfGCz9b1ZPr9e9CxA+zdtOjwQowU5Mbyf9o4uTWom1e
hR3k4aB45E/c5kegmJ/F5QK4FX6aoJ2ugy6dymwR8m8bNG/RO/ZiG2WhFXIMxMMj
Zd9dQ0zIqMxln2ISwZpEn8ifbXoz1miQzdjdst+xnr5Za8hCyIantbsmo/0zDzRM
MllzUZmxttYfzS2l2Vz0a/z5SwS8hK8A9cw8yzLwJYqwOUwoMA5ZI1LSRAUh9ifq
iYd8XZx2OlWLGP05e27ecV/UmuZ61I2qeOxEcp/BV6YxIzrd9ca/ndZRHeXwF7NY
rr3gFRnQVbct1t/mzpmF9A99s2oKSqMLyBVn+rpSJAtKq07IhEccR9v8F76kEErj
FzkOTPvonnxK0FwM1ewx8TJHGQxrDu3DlERThh5G6pZPU5Di3YlFqxdGBOCy0Q7D
jTZ2atCGoWG++Pl1FypSZivXGS2K0yDU4kDcxIbBRKANVcgCR7DnFH6cQU8uo5Tl
HE1AJBDn1CpFrOxVqyhOgbb3HxDBIUIcWJPTJgTVkMhVHw7s/x1khmxExV4rMiuS
JhBdVnmsmYgS7PIsKZeDDBSpQ89/dgdHzGf9LRSoTkWv4hreNpA3gSPrKgOPwa+0
qJrL0qHb72WwS6tootmJct7uq1kc4rRn/NQbC3LYkjfuKWQNsCN3MTy9E6XMKDST
EJqO5yJjNAoX5U3BD5dvlZE6WHGCHXDxJOWzCa96mab/jyA3CD4SMJ4K5B1oUpD6
ddRYODtSlCbPLUpakpIA7ODPnxxCb4VXf0og1esn6sa9cxdx22MeM46DOeuKFi4i
xXifvYFG6UI7EFgbjPUBrgbvhNO3SUEXd4cxVc27f+e3mjdB8rEAg4GYubsSfU3R
zAvaStCxRSdB7gxIJL6oa63SbbRj33/tg+O8kva2AXuKFXhHaf6LWk/Hv3CjvCqG
q45TBPtYX6fh1V8+l5lMTWBAUZMS9hT1Jl+q4iaHWVDfd6JIGFrbAIuIVTkUcDgf
5FD90UyRmZ92pHPhmHawYwQvkbsfqGdMaMS5CMxLjbcNZ+jbA7psT/nCZH0DKd5y
2zOK1peQ3d/m9yYt8ChET9M2nOd/i81F1mIvZBQmgGffx0xSDRaC3ZhyUbh+Y+rJ
37QOKiDCTWtbAABw/dfx5rwEBXcLdON97eXEjc6pj/jn/L1B6vmogoIh/HISIB3+
CaySq8eVf3tdAPRVZrlbBzEdsykDuY3NEX02OA3KLXkovH1/pYEu7tbHicGF+7zW
xj89EWjig/kjF4qd3saJVStPFr87fXmyJnXR2A/Xc0x+/caNLJRca0sXYm+SfZZK
ksy6ho1vRQKs2tIys6ca7C6kDdtIfCMFreVTssCGhYwHIktXbTCbxoE7T1ZFW02F
YFwSI9Mt83cYi3ccTs372mO0wK5QavgYUmmP6E4Syc20x1VoQ6j0HKaYPB0QUlX2
1jUJoZFK9JbvD3A0PJ5ONobKGdqwHHCxaDI7kApNfMx0h/ztewabb5S2ssiHygOR
VIIt236vmnIRFbMaTJKsG9QcUUQ8I7S/9mSLZi0KBEXTwlgkRtWa0b6z/l0ePRnr
wfG79+3TQ9pBBJR382kFDbFfAYrU+p1NHtGRQu7JrOXg2pOJHh4srZkKowlDVNhv
bNfqBVT5zzk7N1UwNLxdWg0op6wpchcrgMd8yyXYcqzXzXcTXliOEwAbpg2KClev
MDwkfD01PD+VQjyyVWxj17ZjSPR5oqXf4g7NJuRHnTAJ1IuNDB40G4lE4oO9PNB8
nW/9GJdui5KnXX3HG0/xb8rZkFOiTWFFcw7siDF+bjDSkb1rAUHPpFBtWZioxWme
2Gz+opWbZj33yNf85MNE1gvyc4f1f4bg6+AjqezjgibUQbqiivom10ij7BGfLr2x
I94cBSra405ImIWR67ffmE+65izvvkqjrSZSUc2ebs4JIr7bB927uxCzrB9wUTFo
4sup046u0u7UD1iIUNTbdb9YyDTmdTm6DAvm4B0Y7Jkfb7pxwHLZHY89Kx1qzpFC
/6QoYdceTuRmLwlXuW3Se/yOUFPjXTZmN2GSyA7HDuyYyJ7Mqtr80LkGLea9RZH5
da01wh24EezKBgFwxBbBfVTfjBDBSoAdrmZZu/r+w/lyh3xr92C/nMaCC48PhrBw
EEZXVhTNEQXJR0PefGVVtbLVjAqRjLiMYT2nJYVmYtkVdcHvy8KRk+I4QNkkAIYY
iZ1vwa4EI/dAQonCFfghRcPPXizm3SA3fWNbnxVbOpTTQzPXbIm6+OukubGw/dyR
NIbKBziJzXzhtatC7g5LVMH1UjIbawRd7tW0amvkDt9+aPAihQGzmzvxL8eV6Sna
JJcFn9Xudq7g9w4PHuq5DpebX3CzYGlLqRdIkWEYoFHQBG2D5rqUpxAuIEtk7eTa
op6hr1xJXwA1ccJ30PpaeoB6ixlQWUKZB63Qr4lf0Q1Fpf2Z6Jw+vmEE9EgsfizF
919sry4mQIt1FJ/Zl6CCg/0pEPdmxQyq1f9na9Y5iJeyQIe99df7FeFBvBLp/2X4
6rFMWvhQ7O4X6F38ZV87SwtiqL0IzNCqVkB/Xj1jpU4ncU4u5QOGUKbbU2XbHpAK
oRdSzif0D3KHQmRG3uYCV2KNt3BC7P6/Kd/IpYI4H8yZPdkKkoE5kzNOESvkNA/N
bkbgqc7ojZItxg15TX00LtqzbDTx2tFgEpzurtf3OA7/BYjaAMmDynwaIztKJPYm
yo2Ff/CrSfYiLSa7KaPCXFLEyB4YKxgWDb6eUBDMxFhWrm7ex+F0Jbd41UFlxBoB
yVF7xQ+7mQUgTf13RDuzq5ynPxa/vYkXg5IhQm+iGdF21nSpY36vQDo8kVS3ApDe
qhSPYYrBTCrauJYTaT44BbBbJcdHtnDCMQG8aicRWb0qzFfT54R5nPgio1S02WXt
IXQUHxs5At5QSjHhqrgVD6rWOr0R0UZGBhXpWZ50mnlo0SP02FY6D8zqITAz9i33
2wd4KwUOg8xJnAwsJpb7HYMbCcRvMQmaU7ybcTFrbzWT3BYgEA2JaBnehCb5Vs13
s/PFecG4RMqee03aGs8Wd0bHQzF3UviOMgU43Hx5RM0GBmRsgJRxEpU1uYn69f0e
rTcbGOU8wDw5vCReBOE5VDoaVKAfG8azTmiuDK/wQzDgcDE8HenmvV1Z3Xs3aFxc
8fY3df7fY+I2avVpXXVdVRQnWd482jF+9kkzB8jVjAB7Xex6t5mdy9C9EVWyOoKW
1xMQgBVC9Q8p1fuc6G7qNqzayq8BGyGov257bSdi7Ow1s4Zlpe6jrn40hB0+C9/k
HLbUt0sPtfTekxifmSNYmjYnj3gAQ0bwQ5qeFSRMkk57nc4Cbq0FrDIVlxEY0ggU
MJgiuJ+3oEGS1eoDhKxWBU1/LBVnTezr2/UE2w9bea0MdGkrN+PXUz8Ob3/Z2cMB
WDFBpgepbmdjTaq0A+Zb/ugkU9tHUS2LfkSOHxp2OUic/VrliNBfok6HVhIM95tM
jCSu5NDybTr7NjGX4GiOCWckG8mqFfX0PblQw32ir7MkN+NbzyFierjqTHwjTv5n
OA0M8ooa5X/1dZlZKxGBmwgv2ELxVHucxYSJKWWeFry1cZXt78gOazolNS4eKoEb
3HywEU7/wwDXih8iN6uQ34HdpUDlfl48EsDrNQ7HRYuPCRHQYNnTI/UsyYaA1hdE
aQUPqsXntCCQrHZZKX2xjGGKreYuCSf42y56+vDUXjSgzZZkcYU6CL4m7qNXukig
F63XHZxIzu5MxUiOD7V2JHha42vbAWrCAICkH2ru98YWHEImDrmkGWzaou/n6U1l
mKNXRRYR3H8CaEIKktYYq+ZcKqq3blezSpHhE5epRD5sJ9uudmZK7E0JYH+Molrj
g2f0NuFjsiSNlgwPXhyy5Zu/uQkh9GW7Y+FDwxpk0I/VfGNdjB/5lzyPsZif8oV3
C4lbESTR8Bzp35krSXauNTXKoWXxqXkSNhLQylIWvM4JFAr7tmZSmENKTYUgEXvr
GYLzG7gwXqz6F2akC8Gjo1rLDC45Nr4yKUF0VlzQZtHbp+uGxf8RuixBUYa0TbJg
Ut6VInn00ZMCCmlS0fMTuYBOURbV1CAuGb5bFNewkfaoWQ/RI02KDDwn+S3gMBBU
abDGfHwJYPEBrBebm7d1m1EofXB8XVInEpkEDdkNEhut+11DRxUCOYt119GSb2r2
TkrXHcWlsBzpC00fOlAcUB9x97EbAvkxEMVTi/PPuuHr4HcJq8wRg1gXIV9HKpLw
lcjINeui344U41CIG+fQIvbFUPcczBtbayrKyLzwANnIZGw20prfdHVndsw2AMpD
abpHd6f/eqvziszFauQAvmm0gMVPF/5qO9Flrvwcc3tFBHDdMeEEVnWKdfYbpyfM
8P4xdee31/kK7EBxn9OuSmg5GJg4Y8Nx99ZGbRI8jQbvneea/qj8FsK2bK7grS1u
dG5aGC3ZgAuzVByjb8sDBjWUdRS+YhY0DMNFWKczXZ9bUYjC29jXaN8u4X6Yxq5w
3xqiyuxvBzGo8+3KJhsRaJwkWXleBavrSprG2EpU/Fg4bM++wh6hgAr2ZVkUbziv
+SwdfDI91fi+9eW7A6EIc0x8I1wl/bIK3ZFRuPI6krdHhqMVXAd7BcKMwv1Rg9MH
/EgwUHFXKunt/uuf2r216DCZbSZEMpPG75GEeoMj/YWasj8SdxhObRuWQu/mwIx0
DH2DNy22ZSaHxi6WilgPHRQSMpp03OZuzPtJbm8cgk30pC9iBDIHqZYeSQcb2ryJ
hyz6xxyJITeHphEUh4M3A5JsqOUTY7vFvpuZ43YIGz8p2MhRg8qyGwtqtN0Hcvqo
wPrKOTHrmvwIekgNz9+zis0UcNS3s5VeaaHBGbxsyafDFSr1r2X0vF9nas39cVWj
P2nwxWKuUqrXxb6gUKtGiLsItzJGXjzQhVmSBp19PygxuAaJv9aVUMT7fVHM+qKm
ZsMNAefQoYNexPICGovF0cAOo/wddb63cgpgDjkn9mlMVyFzcTLa3rNkCay8BIUf
1IMxSlhy/r2w4aKIS8h+jQKhtu+ubgJFRViRFgJhKp0DCTym0YNqxnFUASN5koXo
WG4ziFHrdrA7WCHvatUoltXISDAwRuAWz+Rpx2WEsqFladOhWwTuID7V2MXaBgaU
L0VIHVkwnWkXZu/MmLD6kasxkIRCp1UEranHuEWdvmEyeGB0YrC35vPCJVukdA5w
8/M9DekU4IK2UoFAxubXttCeGghqAPDSHzSED6CBiyrGQbMl0Tjce56GgIJXxpFY
G3wzRyjN8jcNtuCC1G0XGCW6TjqvSyUyIUprBiEHycYi9PnLcztf7k+RAKmPcU8r
1DWZVJcPfN+rocn39K2VmrIjwM59/IfP4SsoiA4/gYX2saWsoU2YNm3OT+fCnxLr
XM4tOL4KuTaiYo3T18LjMfoNlq6jWetpwQLtUBzuhst3CE6L6m1bn2noSTFQAC9R
7rMk0ED42wW7glR60x61AAY9AhofXS9ay2e9PBiHGCFE0ybj05eNB0oYmd6Lgqnj
rpzz5GGSEs+bxVFCJ8GS+rvvszqz/6GBLzY8cPJWkJ8c2Ltra0fx9viRYPSHsZmM
Pc+h/mtM6rl+xDTpPvd/Tx1cVpzr3gLsbv2LUxGeV64gyVExFimEdpD70qOTgOYO
aVB32rI1kNL96A+XPHvlNOkghyTSxkXlLSPX2Z49NEtzHqZq+VLDvEBTyAViBw+U
A7BdGlH2uZRG6G2sCz5eUvKdtn7WAk8dlm/h7ud8Cx8p2YswOSoRt/zReLYTJpOl
mTs9FJAc6uO1IWGl2d/GpPnL97A5kW36JCPUR14D8pmsUSfKcY9vWC3H5LaA7NRy
KrOMEXXIUaOw7csIViyYvJvVcGQVur+eD6hRiZtDUmxh2fk9AckQoVRLRhe6aUw7
zGIU1TOC1J1Kn3kUleJHhbyZtuTQms7654A2aVrD2MwRKuKEGXzcvcKnZ3nLjmJH
7N11mThYgtj1lvduu3UJ13a/kEudgiLVLen7Y+zpCAGR64rwcRKkaq0kqNrWvhHs
ua5PRbltvtsGuZvaPmDuhNAPegLJW01qP6SaZFNrs0J8LIwSqmYlWfX0IXGN1QGh
59xy49bDhO1ka9PnHGOIPuvaIOAPn8H6aj9l7RNxSeiPN6wpFG433O7+jT2NGgtd
ZyyBc0GjzovFxun0XynGF9cX7JoYDlz7lCI8sLd8A24ghhm8XzaN2Ms6o4UEA4HG
RogBtRi+Ph9M03JR1VC8MnwHqNRixvV93vI6Mb5rUZZxzV1ZQRLLPu7I2TTehtJS
8qvyfnx7WEN5hXQqR2+dHNbacpy/f+m7lXECBf5fir+5b8AMERIP/gCAZQoHa6qQ
0LdzkOTCIgOHmidmohEXJQP6YhA2Qv0JsRnd2ln9kg00dGn+jYMWKhF7otogF40h
NmJYhEhbv5z958VqD99iNMj/+e3A0X/oy6CauAKnV/guUWUjwdN6hoWodJ3mE2wx
GFUI6knF7iC0h5Q1mFUt0PYT30MMFttL25K/DDSJ7uDY76TAAwHDiVX9I8yPIlrF
JWjAjHx/6hsl95eqYRTkQ9l681XI3xfnNpfZHeg1w0XI9NnJnsLzh62hAtHCd8uZ
aa8vIXNs14mqfPlZoxs4vb0whfFbn0EACCnzbsPZQKquvgMBrpH52QYv9C5lixcl
HZSFxR8N7XgJPJYzL1idQxt8B9O6P5YOe84d+g/R0VcfhIFkedr6mxICe13OFxGP
zNIHqz6wY0yQHsu8FF92qVVOCnlIviGsO8RmZvDw43JI3YPppCAgxy9g+hRZmh0G
80bIEzXe68EkXCzK4YfTqxDJQrO0hroGDWLA98zKjpV9xYsJEvI603Fq79KtVtoR
f2T0TS5QKsKAt1AcuAyZ6oo5YSZou+2cr1+HajiQBwxXMCE2m349dew8oTDUZjaX
HvBm99SRG5mKdASz1wUUBd6A69f2CtSgf/cvPYL3JuGjFYItKgQ1y5y9XDABBFmq
rvdMvIuPXfqUhYaY3FTUWjwh2wOvtW8J4hitLPxpNu382N7SlWE2Q1kXPWHAZHF1
chh7vdGL8Sc170QZCtFAPxYfuLHv3Zd2gNyrNHPeh/ub5DkTtwC9DWS18+FDSZAZ
sd6H7g9bpoIDDoU47uMBRSKfYFAxfLMAbjNMjNOOWdSgUBfeSvqwxHn/lrTSieFI
lGxcx1Bw/HOM33sJWw0obBUm0kQxcIA6xNoznz1CBlfQWbnJ6vkDQaNj2vRYV5rE
uXsuJElFGWUoUuTUqP6b+dkuPC2Bzlq8uHWBQUtX2eTPYeyXOS/DzyaSIXnYfsZA
o+hSYFLz3i/ehRmfXc3cWhytgdedhg2zjshj4zxdHCvsGeeGvZQ8IErxv7iJSRMx
RCu878fBgGDUmUt3JAFsia0J9znaHDXTfxmNRbSENORo9NC3fbnRWQyIVHsGuRre
/ySY498+vqrMcyeXBADa2PurltF2eUKoR69308WU1UEkMu1j6/WnUZfrk3C1FWhg
ROlz6cMiyGkSyekgY51oOt3GJpwNZ1cA0ys5EO3ZyiVyfBfXOmjgBuC8ZSLYn3Fm
I4pFE0d13acK7TRQW1njZdjJ81Fyv0xThTDvCevt9AeRLEKmQOQbNL7F1pS14Fcb
UBAZpAsaIs2N+ShFPGZnHkvlVMMUADy/yIE45a2m4oUV3d2pbGQTNxQWHZu4gBLl
MrgyA9mUg7eITuYLqDe9rkElzaNbZtJIKzsgdN3n3m/gxgy7cwke5a7HSUDAbSg6
eHFy57TJCmFECiWlKAhjSolUo3Mlfdl3OnraqOqkAASJcRYYtsbQaKYP3PSM6c9j
h+fvWqMB7jk/LLKlkirdsSA4Ay8oLs8WdywyfHWh0aCXuBvEa1kjfNqWkp270Cac
HUSIgEtNaGPX6/euetLn6CScOykrPoqq61uN35AYO5c3x4kbUgpl4gJA7+DIjkIh
2SWa0s2tjyY9XkCiOacMQBMBGX6DKtTFMRgyL/0G2w07YGL19ggjFZ8C6L1UTQXu
JpSWVXDo2CVXm9gjgNf8QS12css7MVL2YJEjKmEu82x6zVmS+vVnZ2rffn3r2k/A
iWuC8Ph79UjxVT9Elr6p3cgp7asfQfD26gPOoVeotvSHj0+Wzelx5vrRJSxeupKO
kO8o1qnvClsEDD0SFxOYCDuaeDHcdyonGCQuuo6DdUu63J1S6eeEzTg+V0A/t7Bf
0TNZedJlj0r9GJE0KOhMP1eb2PljrK/YvAZ/n7+p3Vvno3AtryrBsmaxBUulGMtH
NJzv4Se4LVnuB6tfkOQGd5BaoByBZsudS8dHJXi8nwxsTUFI/FMGOK1mX5fYTqiz
wwpryRcPlQ2XfzYOEd62W0XMTMBGBAN7TvpoNdya5gLpJsjh1Kz5VHPPlPsOs6bw
27EMZhbXOgiRqeXqkpg5OZJRZsMRyB/bLORQL6+OcT+d2marvvhIv+6hFitKD/GP
oxHV1diIL5Vz8dmAigPYGbFekzhyK3PF1DeHG5UMXqVZ7LYUScBp2Yv7L4W3vWZu
5UAwf3pnXHYW2J9RYOND5W0QJCyngAhir1HO3vTTEZo+zHmLoUfw6tXR0CmO5i7d
uwlYEXj4iNMkGnT7gROKVMs79CQ+KSZTuqAOmR0Sfykjy8oZtHx7RXwL6eybuC0J
NoWpXmtnj6iZaRItkbwvDysjVmkZxc96gSF1y8EnKiS65rmvv3cUNUPLqYta5gTE
NxiFcMniQHoWUHLvAP2U2QHpOPVFFegUIZddWthvTD9bqXf732rPL2uJh8CgmR+k
yX/FEdZ7bzpecU2jM/anFUEdfjmVGY4HpP0ybV/u17JNln/i+42bxwE+PL8kxq6w
Osjept6pibczBYKXx0EqxS6DW7VfJR60BYC33ihrMiI2ucjyT2N1SUCDYuaimbq5
Aar8gY419CpgetWhxqq3vTzyPDL0ecJ1iQQqY4Zbyz8G7a4sg4PbkdzIBogiEOCX
g4rEY0SX0Ou2O/sR4AdBbMQ3JYd6nVmKVbkfitLKnJfpYhZy4ZFgGMeY+rcwGaZU
QyPy8Of5winhTm0dG+gPHn0Hsz7xfeD/j48jpkI827YdHMfoErS8PHLOUAErT4Bt
DaxQ9xKFyM7zGiCA5vQvCpQVlsKVKXhJf92FcHTrJxH5Ue7hEA5cLqCncbx/qjmK
CTDh8RCePmWxTqkc9vJUa7ekdkMuXiBIfN3tvowxXMLPorfz/NKW6qAfYpZsW8qB
FCRvpbGf3xBiEDSOicRib38Z6Ixar3YwOb6cfZp5Nt4C9xjSc7pzU/YvIl3JV+x7
SYSM9aortKkGazFLovJB3oThGH0rJMv/OA/zY+lqpNsMv5R91KV8NozMtZHsWp8Y
NCHmpVdqwpX89dyTWny93SXiXAayTAyZTy6WB2LGo78VKDRuOrlKeMQ3riMKQMbt
5nekTFoWhkv9l0GLv/L2XFR+ZxE9aJ0fSqDVgwdginb0u6yny3UtOlWEZ+SvR5rp
GunFe8iIplbgZAAMdNKpaBFSAJYMlF3+ezQTvR6UiCuyxZYCs1bWooq0tSEawztJ
pJvSmJ+bNWrw3fuPmjit0Do0tfGd+fK3nzl3AX7FDCdXOqVm90gVKZVmpDmPIgsI
jtrPfYJsMkU7GYREy+oEcFLXXgS1ONnmsLN7pLB79IgyQfaUw3GfZjxWaao5EyUF
iX8M79f81oU0hN91Kt8WctMPwFbeocNch6gOwNgRbB1Ufdgzwjwi6rDbMulHj6Yv
CvLN9uilQw8cu+C66SFacRYIF6lZRGutSsC6rGjVaYFwOceTmGyOzVOdeZqnRt4z
BXzvRyo/1UGBBE+lt8MqiX9tMEU+iK+R7L+JtkWHGORUMxR1vzQL6zwzlBWp+NB/
iF6M/gLBHcaAoaXteWrylu2SEBYlnrKdRhN63sz3HyiqHUvGfoTp5rlc7I2G93+T
Uaqex+VtiydH4fTfC8IwDU9S9EmVeX13mrbLOCyYwAiCfakFs2wrRy5sBheKelsq
WhgYX7QbnvQ8gaAsTwFat4bQa3BWKzucKi91wrMRsFyR4cYQFLOmlENpHMOS3Bm6
w9/+Z1uwgc5FsvEPfIy+wvhgyRtst7vSz8ex8kOGjItYfOw9vQa+ZOBLVGWT/Mn9
tIL3mbrF1N2SxthmwwFk0IdJsjo5yGLMpXqRtbnHkKBLacqXcfukNeomcvcJn1lU
KvdFwIYHPx+pU7U5Vjbh7GrIghnKEPjU7xSLdQ2bQ0vG9IPg79+chj0SanRLywGP
Zm6hQ64DzXWmXVP699WiJghiuY7u6yElBe/PQA9sZqEwevoqk4O0ktcpnTXmB8q3
qovq6H6fU9AIMIHV929EjhbMTeQ1CEzkCQR4lSkG8w2XCrckdx9pDIijVyBdffRo
lG4n2R8lhdBPNpDjUlNOMXiaY9C/qAmWdHyyQUT8fTcLISoqn7/7DHOTPXQWv4Ki
Anlr6SI/TrbTDpgg7WgpmsDrrmat6JSkjTSWf9Y6Vlpl2cW2EOK7NZpFvluuJ8Do
hi4lWkUbTuZflUZMlm6wmNNBGReaclapeuU/TIKaMmL8ZDjHtMMqR+SxsLjnPfqh
tEKoS3u1Egg1hUNxhjAGR7NsmOWG2szhbs2YSgUBSFOTLTO/P1/Y8uqZ+7BPhzxA
bjO0R7N16CvLo6zQkHCkmTk4yfAaQHIsgi/WH/mt6VINZ05y5d9vDvVGXqKKZFdr
0Ulkz7577ezhy7CzHxBzxHcq6GsY8rxL/HQ9vu6w/jOG6totNEJCE0pioiSp8mqx
vRNwBcOaZzMrOJd6Vz6B5sQ2kNybFD7ONiMuhZ4I5Gw2r6O3H1Qgnav/scgpf+mY
0JvzLZ+pBtAgY8sl/gXCqVmryR48WI4Ux3DawkpqwLSKG18viNPCkQKjOXVHS4Eq
ORuKA9g/46q1rfy75Kc5e5NPrLpLb+zIY3I5u3oWazBzZIwoZsJbpRIL8RiVnG9t
PqLAE6R0bDkAMChpNpgBo65vDtPgMDdGGyArVnpt45V+H7PAFnbzI8kR6r41wCiR
gVpYUF3RxK9bPjde8AsZ3T14NyMeP88DjNASwjVE6kkjP+gmFdiU4wWZ4nsT+e75
vC+CSI6Qf9zvAjU6yPcBctsDnfRVXhRcOYe3QY6G3bLXCchhmeYA49c7nU28qn34
XDyeHFM2o0JuUadvv6Bp/m2MVtFtSE1EMgnspGeYdj0KA3ZiZWZ5nPFZZ2Mk1fGk
5hQwxd5R+7IBHaYJBQxQENj6gfmFymItbZgvEgqlIXYQxSMK0Tm8INku7sK2NIfI
lQBtJal4+Qpz53c+z7rjzd/Buc5v5oVluTXcQa/NJeGd02xvlkJwVjdxeKQi1FKF
zF1SZzDB2mLzUpKedf9biug4qYz04XpBadIl7zXHPVvJh0Sv69Xh3fdU0zBvfhhw
5FENXNyggGyulemmbGZpLVGhgjrmfaKbwWnVaWvlsMrZPqvidS+2Oo0BQzlvit7B
M5gKkreYLEKho8jLT0VEbec26CRjzbQAINfknwpmbUJxHFfhN8CCzIzstpFRsjXE
+MbEkvQvM3bwAhyjK5SPItUYxhin+T7CrXhPQU6N0g31Zl+zWGrZZRujPopoF5qN
t6eo6zqRsgO1rtbJ+l0E71ZI+9xRXvtUVCSIiZ+RKWh0+PL+wSRiiwziygiu9gCS
wx3B3iVF9FQuZXt4j5Qz9OrvGzy7SePMnilasYOUyQq+ZUswNrsVJhi8f/Bursae
thn9ywi5UyZpjiOfsHVDAckbjOXhCLIy5iYLS7hAqlUY53WEmKU4aav2Y1ZleP65
Zeh/0o6DlCabOX2CpG3+TkBRspBewPaspkNatJpX+dDV++dEm0U8shoE8OKl4cYu
OREFGH4sC/pxlWF8nw507QgQAm7LPI3B5iKHWA8LrkBQpaT9juEBFWE3v4WSKmmC
+gTc52runUMGJsrlL4kl+SyvmYFPCld7VnrYHlxzK/otMNfIotC7U/p3MRNeLhU/
5PFi76pKqrOsHdSzzlULbaC2NPjp5SgszZpUV+ZzNopgrraT8emABxB4v28a7h+d
l+fcaqxU2cPTqBIjB2lO1PFfrnDSQrDrSRSU/WOqTuKDiDFngl58NQwRpGe7/Kr1
mk7HBxDOLlFiwMQ67nTKBf0Nc3stf7Znt+ah0KWhJV/Qgr+W1eM4Coq/fpMS2UBq
+Fv0zclk/y4zybAj2wMiyemAzGfYS8BUzjnPku/oLGdPtEPg/e5JsL+B9LPNXXs7
4KNzr/yYVlrY2KEs9pbOY6JEvoCf8rP3f2kRVOMGVJw9kOe5fh6KUdY6iLE4kcNl
8w86J9mgsGS0xX8GRLO7WGRhqUiZrNyC/B91bdAZfWUBXT4b4HaDVl+s0Cbl41L4
MWFiN7MrcQiRDmLg8iC9uiTmqTD/p0bz99g93TDLFOrT+Oe5gsLZ+Eedbu1jc5ub
xXsb30Snvv9EP4be1s3G/3YoIv5L9/5J1XAl593BA20l8HG1viGwoH/OSA3fZau5
2WRuua+4uNmCQvHQJrxVnw0Q7kcB1Fv2nnh3+LUuuBwcwpT2sYC0FVFpi6exSxSU
zsF5zsxXhg5Z7NVyeVS2ujXm/TnCSg1/S0D/GjSolmg+6GWEMfiXGHmt0is3Tq1t
ZYbhE9DvhunriVsVXjXqfZjSEstYDNy5rgRkwoojA+0z2k26LztIG+S+0aik5ab9
MTm3RQzyhYJs9AaQGFqqScN/a0qbNZnyoI6jRIVZKKc2LvUa7ieziXa1pLY+T8Hi
nmCAMT3zXRL+32AxC/t9TNYUusRnEAdklcQBlmrLNkgbCA8n8edalEeDlnx+QVi/
1bGNfWuc5fXaPUfzSBUIUqF6VUBQUxHeIauR5CSGfkdPiqiU33iO+JOQWkWnjfBo
XVSXr0oPlIOeWJoykCJbUMRqOlAdOMK5oA5V7+j1GF1z2Z8eQd6Waj/uBxeob2XT
tyhYuI4xbYnpTJpxjO6BXdcUjUaGlDXzxEVuq44t4fS8BR6IqikfmIjTkB+iJNNf
DPOfJmSnTvmDPQryuem8zDuRToDEdLS51WRldB+vuwkF5c6UlxkWHVV21TzT+NOs
+APjNW+U7AMvYqUAxf0P+kUYhwWFjmGS930OnR4CkpWtLHYxleuhFSkP6lZpRKem
l2gEZ4ARKMfqOTOzgCG/HMp64E1az+QDm2wdDqmzmOdqlhQpJ0DYQzk2ABDb4c7i
VjX4KcaACUzg+sbNESX+aVKo956fctRZ3e7do1fkVHPdbRSAHXEUUx+TrYwi/JU/
huJ5e0Lb4bqW5bmbp20GaJAfR07FVUd062vk5DhlT+QBI626LmhNIo0Qz1/cIDJz
iWauf+UolgsrJ6c2xhnEH6Jc2hmkT2ZQwERIcQR9l07Yw1rTLCM77ctbuzM3DiBj
6pOmRy/c3LPnfYGTUytaykiIFjylktcf0P5oebTJ7kDRg/SGG8MaNoA+M7cATPxN
mP0TP/r0xoubh8LXt/z5JLW7pNiUnYLfqJMnQ3wvP1U+bHGezC1/auYy8xVxxtoh
8dZ5lxgg6fhW+w4fPwd6UGRJavfsrJLajqDQMll1Ximwl10C8h2KBcLVH4r5o2rE
g46L3CMmmvyZDv95JKCDHiPf31RFIBFwzRhQz/sd0yJp/00V4Yitad13GNArhbr2
3sbNkkS8tCzEkxuTouv4LTITOPpBMgN3o1pbWg/zoTx5uzkxFLyAE0uIritijohf
hafdlgZUnZb4Bvp32TtVEnSAQPE0eGJTETlFe3UONBEo21qdH/l/hjFfG5WEfAwn
kBw4l1GujP4XSI95KV7ytLFNwIbNRG6ImxSw7nrGgKfFXMA/hbXhjN8O62lkhLbA
+pNLGI6V7/EpUUBpSAPJaPzczKGnJzf/clpiDyNoYMc0M1rFqeu4Jc+it5RVkRRP
Q3pHl+iLLy6bb8dLiaqUui1gt0K9S6N/6PH3f/jxWKm4NqJdg3+r0ytErbg4dbA9
Q8bMRa9v+9/U30j8OzrY2mnVtwc5WrUvjG5sDfSRxAwH/jVte+flO6qJ7aiWcaOi
2po3ztBhFRbMP6UYozIUFergOrDQYsnHx3mRjY8TZVU/fApIJoxtGZuI+k5Nwy0I
M5Va8V+JKLqE/ST0/PRWkqnjkoeOS7QUJEa7JNDNBsXLXHyaeBJNqbScNbbqclkh
b2yh4bIyRI+CJ5Kr98cU/cpPxWYuuzdO99Ec0r7cuBH8NdbmtsLFeW3DO9/JQUKw
Dr4C2Cflf/CMqRaHHgekiPRF2zpOGVnDwFx/XHDe/aHgJOq4hUnl/HpWTyR24jZ+
q3I8pWWYpbvlPOJnTwk5q0gNhg5/AfdHqdrOVBY9PBg000GyoZXJzspmjBjtedzk
jGk7U8jHwtslxJlbHaVmVsms1UiiaFMCICSYEm4ZnYZtXUt6+ICW7a4mL1uvHDPV
8j6JeCu5pIJCBPdpiuAHCyfCJITFBH54ik3Jx8f2n0IBnq274gi6zPuksra13eM0
y0ZgBng0SyYOaTWcb8t6AiMU6OLXqotgBdQg8EQn1lDNg4Qd63ayfV8ZRK2fO5/E
qTSJDObVQe0hz75EOeP6OXMMKSPaBGJ59xX2Hwi0resc+6KaBycnOzlps1pwPxH0
uQ9sFXbUK2/t+lZQe5kQY5B7q8rME2gBzP5rCzN+NTXBjZBCoreE5IL0sj9y0nMp
j/wyP3mb4ZLlIdgpTRlam8eYUvO/ULcOy0pjP0hBvSqh39EDmPI1bYQdTq/NlVOs
OlVJRTNS+fEbtpDJ+LTQTFlXrot2aDD3vGm4Gd5DY6wVs0OpS2cP4o5iHlK3EU9V
VuU8cmMD3BRupjBt8MDYgAnMpliHVO54hnxmBqUIW6/K3vIWRvEzCmv4Ta/TCQo6
KrW4vn7fxwoxfLld6lZGrCxwPrDqDeTdNpe+6hgbgJbuD/EsqdHPBsntUyyNdqzH
m2ap9GmkJ6i2APgXXh9yDO57+0iAQ7ewIwCZ7obCT2WlDhqBUxNvUhC3XHnXtNil
jxBkUF1i6nxWokR9UGGhGu/FP2fC9gC1PqfNmXAsL92zaj7NrR8XnBhBL3gHka/e
sjPvkyuwH5JPWSw+kshpBcx8D+PBFnjhKHJjcjDN5wVvk6AnyF1VWF+JyoL3iW6g
2ighI8toCDssWRotSug7PxnXrRgiPfWXG1anqrnp/5BHVxhbi+dzXb4xmjpCVaBq
PuftTHB6UVuT7cPFpIdklnAAdYgStlUOYFVIrlJa0ttvTB83eqx1xx30POSmFyDJ
WHfHHrmT5bKamM6uiVkrzazKCy8aM4OlhjF56cjKn4svS3FDh7FIiAKGcVinNg5M
L9r99Ea6yGMm8DT/yhvvCJJ46XY0Hu3Q2lLHpHZCMwXZudD3XyyPqYa+h01aCa9H
To6gJGPg8bZRMs24jE7xmfd3WtCw8kNrDOBTEZOPSyCmvTTiVc03dn3Uw57NnSME
4gwxnG9vOzgIO10o7M+CtKkuy4JBI4fm54/C2e3uCYGSvU3+zurs15QPTsex68eB
phuqFw776EWkonvh1hi3JtgUGniH5OXLtNvI7eseNuMZqbjiumbrn6Tteytgjmj9
3+54FpNs729/mB6dSSF7fQBXtKsbHR0DVVrhiosxEjVq3UxKP1jLxarHulEuS/R9
b+/vVdn8G9JDuk9RhPW1B0tc4hsyF/yUkh6Ofb/u4rJZrxsmwH/Yq9IX/eHNjmoo
9hxunIq/557iHgZYCIO+JtkkQrbi2PfSeZcb6eUjscqNDDdZ1rNUYJ34Bqr20X0c
jhgZhoMAzJrHr1MDrU2miIuiEcpgt2AQ3gSqRj7z6uHqJOlAdW3E4uIqCaOZiNr9
K4gMNwHfqdDl0lhaj2n+wfuLxlQPTwOdxh/I/RlbFA/apI5XnAIxz0wpEyOb0CpK
pVktkJqC4WOLyPNdacFhU4l8RmZaFzi6+in6ZevMlkLYo28Vt7hqcqyXRIN1z/Xd
uDf7EtBpXqgGjai+TGoB0SZ4A44uyTJZUioOMxQZpYIXElHqFkbdxk1zD0lqbWUU
vJGyFihxas1gawkWbGML8N8ZaluzyBkbWmJRMUCnSObyIo7Xbs7Eou7N0iLzNt8y
RrxxdggDHz/MlTbfjSz3KBvTDv2QjBt0pmfJ7mhqdCQaJQq434pkmX1y7Xxh3BLV
ZxXndX8WQNBt3UAxeEBXg2JutbNwE8WeGKOAENIgylfLfLuH1a/z99WFkLl0NMcA
pLJ4ou0y1pK1CqZC+cNWrAAGOzUpx0RslFAadhYAiSnqFwpjDD3XcDlhaJUN7Ioq
AoN5e1V2RIMcfq35uR5cceRc/7ZgrKr3yqpMW0xpu5yQbf8DC+nnO+Gu2m0yim+O
wj2iPYf9uBNuPCvSJJ9Avptf6WSueDBbawKtwBHRXRnwdSqV1C9NOUaF+AZ7W7oi
OWaL+IoK76h2egA5DBsOQxHrMhx2DilNX0fragYZqa/Kb/f7+JnpsU92V/mIyWbU
Tb6eXwrUBme4+FIrbkoEseAbamHqKRnNbyF3ioK3OwUf9opiJu9n/wITZLrghEep
wFIQMaeRqkFA4LMUnL0FOTW4Q/DeVAKTsT8b3YIxIrljcpx2wRsYd3sbNqomwsMe
sSUR0SZeX9w6wAQXxzOZb03Q4sBTgdXNFTR43kfbBLkVXOJG02loAUI3Eg+Ea/gp
VVjmpFsw7T9XxwP0hnGjNEyIlJc5X/Bdn/j6LaCGvLTjLJPp0rZ9bFykYabt0Thn
KNsVyHoFMojjAjiANY33YaucP1/KZ4eG2+fnq/ZNRg/5PI2Ksw0WefRDrj0Dqyo6
xcndsGp3pClIUn3H/U7DrLCUVoJAcxFWjXOf3AH6NwDyTtHpPU71tDbRKSG6dfPx
mj8c8B/envPf373PJOJahOtcv0u8rTJS2+hLxd6ReztDsq8NZ779Ubl0/Tgj2E7L
QwNSGRLJasz/uFBZ6QPnluTAQ6HG79FFCxt6lR+stXyuKwLwC+cOqJEQGhWiaVJC
1Dxg6U0hmyhNqYzMhMLR6grj143gCEas//J5WGo7ymGeDF5ybM/Hx2xZD2UXFlyn
TyJYMHc89OLAkNN2qjeCMS4QHJ7RpYdgW+culcPbDhFKAUXqGBwfOCwz3B/oJKlP
yzkPHI4wmp+L5ztGPJ/H9rebmiXMtdYLASLgHyPTWvcvvQmMInwBjBSr/E5y/+6c
TpFDtPzUhZ7PZkWvEduhxvxfA2DhtdEH9e1mMkr2WjfmDA3fLad8u0d0U/r9yTMG
C90wOQvShcX9ZCKS7eN3luTnCCU0UF+UcbyMNFcLdUNfvqPpMw1/A/fYEF0rS9zo
J5TeEJM37JbOI/I45An26+jeRpSbFnEIjXMfeGvkvw6wE8o0id39iLd8LBPXhOou
2/zAvN7PbgKI/Dm8/6whTqCmCHZfy+WkzouOvn3Mpy2FtsnXWGGZXlGWQpbhX5pB
0QRbRmCzWCYTuAWfw+nLkuzDN8wDdDkXjQYp7VAxpyd4oS7yGNKD3RuIliK7RxcA
sYpcnNVHZsyqldhM/VPFl1UsjL+6KKmBVWLg/EUnhL2memnqPClLDkM7uakx5Wmy
aZz0rrQ0FnjbqmilyTd0yPmZvpZwmZquaHi6HgDGULkZSjxFxn2gLKR/gPtatuwr
FHZKHWkIEULfhpZ7k9lTI+DRar+1dtO1tCGKt5RGXw0Sv+YwllfGq0k829PT6lNx
N2K6YdPfFcnipjCVJ8S+MoKJaJqjdzJRHy+HSWe/StZCUy3A078d38CgNNAkFC2X
5s4UNwGhDScWUyYfJvM/Do6zGc8L30cgEf4Jm/oqo0l7pJFR5vQ/xhP0tv25zXPE
Ph0ZjFiE9d80ZrBKUuIFlg1PKFW3nIkG7bRQO94/kNutDsG+lOTGKIvU8/es9PAx
9s8f0bYRtKsJ4w9im0SLyJmTmB9xrPAr3t3og0vPVK7QiYcMU08enZr1IsJ06t7X
ukVyZ3GrRM5IHPadbvlImdE/f1nbKzdNy9b2phNBRctqNKjixGpmZ+iPqEfJHprX
Y8rdr4KU85E5xWBwX1ttVZBLoTj07vfBPc8M6CL7kJeD61afdJ2ZwKBz2oYeiypa
iftgC4/jb5MboBQxlUPeid17BO2qIJvm6QfkinZ980vGX5FpErObJJtlhkqVZpI0
AyyGaIY+pPqPYT81z5MJuK6XfM/weK/LCV8d4PWlXDbOLQF32RrEmXYVc/sj+JfD
vqNfDce1oPU02s4PI6Vp5SWDkUM9sqY/OASgtkVinyD4/Tscx582kpf+biJmYEw7
TzbB65Vs1mqvYcV97wQOipPKFg0xChAWAO1wbDQuVasHxNzd6Om//Yf08272sv5M
7E2K2ReYwuMjBpjaX3n5sUSUAdDytg8JNHqn96tXtqluXqVCvwDd63TMUXAGoD9H
cLt8GoAQ1RnXXL3rOLFJRQHjszr5jaAoXb0GvF1I/mXxVfZMGphDge2l6w9HXXhy
41YjfRJ6qPine/oGIUMMvIFtc48YcY/3iGXFTFwLtfUnMlVDo+7s4viHz8GuerlJ
mPvlpSa1hvYnzx7EvgXj3sHBSqQKE2r68WzN7FVzBUJoUQiOiS+WzvYQn4Iry8Et
/xS+M5APaojSRbF2Q/3Qjl81HTPF171rRMY/RaG2hPKIscUGwfdLRIgWtUZetRYN
CQwhCHW55Y8YSUXzDyrrZZ9H7tPMLwqWkfxue2+0vrye765XKPmS/Jk4i+PXFL6A
9RNmifcWPhfCTumrmHwG5FvVru/kVLfw1jSxdeKAfDuHb0T54gFxlIh4ZljhDMKh
JxUq3Mlu7bejsZB5OkP21ENGdw4/RN8hw77di+pllr7WjVTyrPXNzLHNOuxElhog
O+sycMpiI9fi0replOJWrVovHqw1UJ2MfNjG3TT+fuDfEg00Ox+mtWnAnTk64Pg8
h1YcnVYbZ69VuVBMpk30ORDvIXMwFI3bgKV39DGTg8QeNlxvs5XFpx/p6lm40NaI
86ILpbrRQ1LWahDQj4K8sNdnfw1TkueNGPtvToeRP6gXwK9BhXowpWjqhli5BVmQ
u5CzYeaE/vQmxEyGL1XMHhO3uf3gnwoXA0ANChPR7UKP/lDBLFtjwyoply59bSKu
aePggXUDl/zZwFTFTn7/fCD/jEkwPPmPMj4LGhHqRb86m9xOGwdmER5LYg1j0ghy
FHCnkyhWxN4PHZ8mYYoaSIasrPPuHBcp5luHdlLLdpgT98qzZLE9cK8n0wf9T4Td
1mevqCkfjCHbBolW0YFhyrNRGP8iXTdEbVODZQ4lCdC7lnIcVqhlekcRM5adx1D+
77K+2XsM85s9WcxUknMvzTYhNuommtTdMP/RPX2jP6OCYsIRQdxoAnFlkBwx4baC
FaMrJpb6i9jy6FCJeYhBNZzAQ93vtL/h6cVeZPOSQb4jgh8U4Y0bGiHjCxH2Vpa2
tVib46eOfHgD013vsPZXQsYTgDklh9FfT5HVbvpMUiLWj58qKonCCtlNiOvsmrtp
sWaeUhZW8waFc5aGM4TCPMAAh7+z14PIRUIeggcU6LRlCXNOm/lB44DuyZBtZ+em
DC457jnRzI0WGMjA5EHoErijRRxGgLdOZXEtcFc3lMF44c78vPlRjRktWWWXZOll
Ivt+J2aW+YTNB9cKUGaqrNaizh5L48nOJQnErg94d2wdLDaKhvGPf4cwsHPHMEQs
F2YiqJvoCyugxgSI/bylsC4pK0s3AeSX4n7FFBSU3L+2kGdFd/YNSjXYzs/FNADq
UmcAPDD21ES6z1a7M7GWQx2QI4awBO8vqMmcSuxrRiWCdW9Es5KPOoU8LuUwdTnn
P4JmLU0NSXatQXjgSWFAsuYyCkfC6ZpZ7a9WE5sBm7g2Kk8s/DhsIYXc4zsu3Xvg
Ry6zC+FoOLau8l4cORgdfspE9hF3Vir9I9M3pV5aFKfHF9rSTEm3gfdw6pREZSXh
LWUIxc5SCtCResUvi/uHIV1tt5tIaWNJwoRazu0L4Lxl9/IE75jtg2x+jbxiq70e
FJjjxWvLo6l2HXHl8dhj1cpDYcbXYHk7EnKtvncKeqfsztlPaHKZIZOwVcXd/J/n
qGSnosX10iFIJca+tMcVAojjq5B/EyNUiBXpQPnekU/MTTagvCa4ZQKBCRoiecmD
m0Emvw84yMZAndATnO32YKUQAoDXuvBdXHVqXR5PWqVWb48KwJtx94dTs9Hag3SW
/ASoqBujPjawmsCh3ywzdp5+dZthNbQpCx2gmRBaG0iWfSZHTp6copu3pf1JFJzk
XV+RKprMF5GkSZmXaADCbReRTY4jT7TvVzB7a70D5YTxJ21Yv2bRR+oXK4dZQLrO
uGibparoQaFpTnTjZKqEes1fh51clDZEtCq1EDlJ27SE0yLZ5Lqe70FWhdtrmH7C
7Jv9eWvP566e66FFswAX3nu5J2NPmT6ev2tYXDU6MVQ9kQBb6o0CFtLDH6p4X4cK
wNK4emu5g+kgFNe2r1YGL62/hCBqz+wd2M+/Iwn4lsOvtDf4uuVjbkIDsDG0VuKJ
bMyxcFzS9XEeiDWw1Vu0fkjc5rJ83FVKH7ddJXckup4yaipRYKtHGv5x4iP/LrV8
5ZcxLaFl+B7t5Ly7SjSdtX130/Gk8LcV3jEVcZxsQTNpu29jNRemNT5R4r/JQP+y
lqHrZeAmLzxcfWw/SfJa7gUp5i6vUTIfyFKpTXVRigBu6e5cCXBxaj6Qs5Ee2siT
MnhUqh8RWjgZYp0FjIYGL/NpQAnMjSij1RD79Sr+9TAf07Eyloqygnvhn15EJpjk
jzJ4Ud0EazrK2OlcrPz1lqTUo59jRlWMzF8ILsR9cq7o3wj87ohAz2oqvXbGG9r9
h/MIdOfmqPz7du0zSLt5HbmsHtHrITj6qYqw9ZxhfFF+1I805RSqUyAaLdM05l83
I1/pHkS2drHFk3k/1wNP0a2Imcm4HgwiWGpmNTGKF8/MoFW783m+SQQbSi28+Js+
7BnhmkZw/Gp1PbbTAWU70kp4vfC4Q8ecY/4+PCrI100MW2E/CanZD4FKA1NVpzEj
YpFgxHBL3UMulgMk/N4kZ22zpkyLC+DqhCCGuIcJWzTzuYlOFOu/o/B74G/c1KV+
cAAzqRdXzRWgAjg9o3jGMCoioD1+da1790BwB8UBpm/tq235/AS1KgMZEvhpATX9
l+58XnLH2zk22Jrs/BJwU4dHFWU9q+No3GZhn5BXvHFRyNTV1iuz8jTcW4CFNwf1
JxbCpzanTiKmNdNHtQpPSJD0HL4lWHJEOobssagc8OxYILnTa/mHXLkOujzsqM4V
YnfBNeanjdizQYpFLwMrL12295bPyiNfdoBgxgSX+Lqpr+zm7JCuiTsFw2Zf++2j
D4uuDhMB54L8gv6p7qzgczNvlA3rFO+RZIV0ZDjSk307fCFN/3/FPvDoF2BfkM7k
Hl+SrUYiOUxC1yXtvqTHgE3BzUC04H8h3csBGX5D4paaWZnusTnqdMBzAk1htqpo
uWWQPlctm2LQ5Z3T8ZuL2CIyLRtx8rs5q+lhTHBkqLzh4tvgBIObCC6rX4J6TiG7
/A9Y4iy0qTDTSmY5qfD1gga6rKTtsWpvde5giJqHEztJy0l8yd1PHsY5xMxH3lv6
sjjrWXbkF0Adc49K5EcBB9iCdRRbLNf1Ek3p6fs9CAXfTIr6POTkydLOyrqXfaAj
/xiGLmkAn1gqeoWnhqUCIkkHo9QeZDS938oc9SYIBau8XO5EZ6cWV2HwLB/AlKue
z+rmeMtd6iZ0RY4hR5CDXd/uFdraMlMZRx1sg0LE63ht/mTrTzNLSAvw/VbzrR30
0BXb+59TDcKG8dpwUns6V/wptQJxle5jecCtGvACBGVhVc5mtKX2x0424VNjydhh
vbeLDAobAc11mRduxhNsr7+gCK6dkDFV/DTmGvmwgrON+7KhXAR2mCFW3MBk7D1s
PK6aKlfUBhqhI/qStGJtMGtdPv/22FVOQHlhyVkBTDnTaaNz0VPY6cBlIqKecuOv
XRklofYb0AfFldW3x2tYYbTrWaR1y2DhAHm6KewTKkek7jWqck/yaJcyCD5TvnpQ
yRgin2YwFvsM36KFIr75AJMbJ+PGX+5l3bOEK8UzgPGFtZPPhJbPniuymQXvHMfe
MZq0XvnTnR2YzQ2XniM0VaDoyB9/APCNaWsoz3vKk1ZDl7NjQ0pzbJ1YsNV+Ggvz
QYlhqwBsBOT3BxifLUU5N0lsGMVDOelwb9xRUzaHWb+QGXdkHnKfVlM3HGooix3h
YP5UagKoSK8V3yw7HMX3HFdfBbrTSllMAHTgIdmsOKGoSjSgQAwzdGV/KH5CmJIM
EouMZHjBtbcFPLRIQ1+pybr1CuL30o3iMzBFl5PUPpq0I2FlMFdMGSFUKx3l2CKS
lA9GsdqPOlEODbGu5dTgWWMuBOVI/TP7f8n4gI7jk+lyJNz+AEdxLCt7WrRY6I8l
iICpZX1KgxkcJCs3zC97DXe3t0pgk8pm0QR1iTkTs39xmnYDDQgmg4LA+eqKATQx
+5XKPm/O9YccxmmAsnKdYtoEjFVRu3QByYe+SNkisdTD2Al7Tvl106kgKFnJKG9o
UvmNvbfproQ7MXAKzyL39/amPwqGIayLDxgNDFQzQ674AWUK7DctmHgDtCCX+gN5
hf4LpphO/leSpLGdlAgAgNOFfkkly5lRzpGDU8DR9Ackp1Sl8KX/1gviZs9iYSkK
hwzIWDuCblRV/8WkR75aMBMXh++UaukFIXSEIxoqi47xFmY58qGsU8+X5vLkccPv
+ThY38t8gOpKUSm2W/DXVTB5Y8zlEc1LV0n537fO4EFH4NviE2nlLjtODNnf8eBC
9U/ujw+ZIjIRz5teTt856Y/+pwjM4TY/4SnSM/r6hdYpCI14KpWE8IyI+GRb/YQU
fAIhLKYh7QZUKv6Wq8NHY4t5luWdoNLobg+nuPfuflKjDZEP1W8pOxfuRV/RWrUQ
iOH5Gq4yp6mb45wMG/OKcOF8WH9etyCTHFjU67OJ2HotM/o6LhDoQlUdVyAV4OCc
I7WXczTVvkd+prUSIvjhri/LQ0o+dAg0CMMaXTogYSW0Zj4YfHr7Xhef0OQzxnoh
X6vxfpacmaazn6Kylf4CuFZ+3pRzC9AtLkoshnLhtyjEdrzqpnovQQPMUcZJNlvQ
WrPnax/Oevh/IQU37IzWBwGpUk2iyJPHTwrsuanyYrlNWyDrYm63FXg6UIA3pDPw
sF4mXjkKk74DKpo1nWhiTzwViqALD6gdFcVRUbtEIlarHJ3y3/Fa6CPlJI++musF
n4iWVFLyp0/M0DnfgfEZb+C5y3HdW1RRfxvUBJyusSpCarg2m7AQeubQ0QDzIA5a
M3LtRIwv/LzMw8FHR+i2c9KFQSgM+bkAGb5s1U3UPtbHfsWk1TU57EGBWfic4VO0
VPGBCSyXwaA17MpXIt5ne8Br9v0PNcsi4qdz18Zr/yGuCNvkN/dICUw6g5K+ddO2
qhQHH2BXy0CZnm+JMXcWilms/8H2Q85CTRy8zsGX0H3NMc4woaYPAQUP9+wMNtYs
Fe/igK8QGDl5h2uo26kvfNF1KeWOYavMFhQ3Lh9XXw1bFKwYOZf3hfFHUL17eDrR
ZIQvpINkxlQ1IukV/zfERMmlw3/v7BWk364bpiSWQAUUjRaQ+kLQeEvHMQY6KQ66
L+yz3h9eaJCAs1LayJYJe5r53yooyJjwyi4pbO0JNUSTRtYbarM9HW/cGIaLq5AJ
nDHSSJhZg9iy2k/qoQp+hOiURw6lwrh+/zO5nbQozbdejwKjB5bha0G3RtMSbRoX
Tij/yTEEnxe4GQo24HNsPN1ta2kUxJk2ahE54IgvYqyq/+1hVBJ3C0pAdfjgSqom
i04JGZFjCvU+qkIRNc3g993UEla/VMRWj+I3b0KBqtfQ0WKbbnJ2IYKIfqFe7YZ+
+YuSVxWuc54CWiqLTQLQKitJEuPAvNg/mYzH0RZDTHpaP84mM9uflmuawxzEUCmD
FA3TXlxQI3esxY1fjpaCGjJMue8Zc5Bbt1wNafLe98e94UB80Chg6SE2xtVPnNWr
1ckRD3TZE7O2VrO0hJ5nnJofYRUj64syIe/zQK05NgwxR5NQN6A4HOUUM+MuPNpC
PDsV2PaOiz+fVtjJaqE21JNHBgGGSn4uKw4nb6UYDvhlJYHdwvesGkFtTiQXuPik
/PaIAfosCRQmWiRK9mmdHCr4M2dMmDVC78vteXchK34jwkZijhQ37MhHu83y78vG
XVZ4KIABvLwaa8ivfXrXsPPHtciZ66gUfd49hXJAhWM28Luh04eLngZ9DcRQCQkX
iXYLJPRX55JUg39+7WLHQve3k1kpXJNBfxfkOELu49te7vBtdeZkfZJo8xQ02ijv
2hYYwhkqmJhIvIOqEtsn6otazUOUkrezDZ2+U0XduUHRGjVpsMkcptq8jWwGzA35
/rp11gYtzvsKaWAB5s6sf6TDwx8YCIRv+vDJ/Usv57vmCg9f2+5ciZYGqRB4gv61
uIUVrW2khCZe1oHNtVVLCsc5I0w2tz6N5idrI/yL41UfEQCI6YZjCP9eZxISUpGR
+E5iHvYvTulmf69M4Yu3U51QQfAjaj2Tkds+BLtWAqB3DdE6Ex1wKTQpsmj4I05m
n8UIHOFGbSa3dcol/DCmm3dqlfOj3fGtO0sUfPTpzN7A4Ae8+Qgl0JtyGbtgxHDe
BEdAzRrh+8GCKULI6hQ49rj7M8LZDNr61xOstv/TOMQWrebNsHMloq+jeAeSUpA5
PgP5UFrMQU2+XBhGkSpkHQWwwkc9ANP0Xmga4nPXT/cT1HCtt/hqqZTcFeKPQkDR
4GJuJIvs5Vvt4nuavCDvAvckK7b1WwU+7RurshipLq9kJw0B3vS6rrSYzOtEhJ2C
3Y/CwvFYOuAALidXEp6+NEId7bkaUPdlj6oM9/EIBUfSva/yDfImPJ2KavajzrxZ
VHFFLdXZDIymcuL+TeYuMiGTHqj2vE+iMUwX/fvu2U90Kqoe+spak3LxClrbSpgz
m4kHuCKJyk5yxOLVYjgOeXcVv+VmFfmBy7QyMBIRmoq9Khpl4wHxNG4Tu65k1id3
/3XGqnqOmsqbgZjGKbNaytkKFW7vcyeGa/dkBBiuURfIJwusVMm0+vT6kq4PGBhh
CgRjUzgkMNbD8r8aPuymdrwyNHnS+hvuqnIqIarF7CAFXpBwFXPFMQWfEBfe8j1g
FDvkmuaygJ9hmUTPt6y7CvFRQGh2HlDFG2gm/3VgvfxdRQTAha9JfbfZ57qCKA0n
AmnyT0yNaZPiTCwa5WTjFGhGmEZiYBL9UJ3yL0UMSu1NwEq4hUx1niMCfQkgC64Q
cdv9HReotWPvQGE0coPNRmSFsZ078uxzQhDjKWXhtKjlen1pTv/BplLU8seDTatT
BdL2N6wZ80r4FJwZDLSuvZGmv0TewqNFPAlCeci4zMe2IEKiexLKojj1mZfkTQwu
7StfukUJk7XqwMNVunXp9ZdBNb2l+BFCHti4Ion+YIJRLreJjTg+ZpABQmIEUFfj
fK2YmkyLsNVBi7GzumBUlAYwrEw7sdjQUM7AGdgcSRJJiW2EIH0sW9UDnDfXlpEe
idmgYetNLTr/NbthVbdrIV9voZercUMhB5KzwAubAqmSCq5wfyDcMYuWVLEwZ78L
v8fpy731x/S8s07EesYAogIjcIb8e0hEAI/uP6zu/b+hP4XdCX2ax0g77cW9HeeQ
IYKmkFb8+jLKr0/8zyWjE2D4e4B+UGiSL28qTe20kU5cZpvYNaZd3ZfxakwDtiWJ
ricTBPDwi5N9iUaB8sjg1QNV8WBRqfo+4uhxyYMiuYNKTqSWxGb42Ys/Qxb6/Vyl
XHNYhhrkIBwu3QxCRHB+ZRPQtFpU01Rk8K+gr/f1fVPoFFGPSYcf1X7bgo8QNeBJ
rh7bobN5vZe0tpNTYTCPc1hW/J7V/H1OVu7Rn9e8eDHQmHXoAKO2934dG4x78tDj
JJYoeqPOIyYadYLAThvMVo9bzvhC1ZBuC4Bts+nnQGW8r8+O2V0sS+RQP4c98dYi
OUQ+t2SYlGDMboa+uq4A6KWLSr+MhNso72llbXtvpKR1/852SqaTyVU/3vxsgese
mdWMIfd5SmWRfopthYU1GrNJls+l0294eNk1cXigEdT/6QOyf+iAAFiizRGC380M
16QtdI5T8zzuip8t0UZxwAdN9ssElJIYFATcwXykJADr42jNTrjgRAU4AddNzXjh
QcC5VRv3vZDixR4DpuxY7cDgWderxb6cJ4VB0PEuDnZY8mzmr8R1NY9S2MEUjgwS
TqDmk2PZcAE/Xi44GbOeF2Ph/v5XAizmiaVTemC9CxFf0G+08A2yD1wmZowkFkqB
AgrhsBQvxMyLU8YRloGcu2LoTyFUjXYYfwTZMMsVgWeFqighpLyTu5T/H/pEceSI
7jM5Wj7Aj1qB+B0gLMSMyWBRN61/9jwVQmqIryzDM4xLBDMPT/SHOjV/I0KDl8Ix
VMI2LUERIdDw9hL/A5n2kWhD7dCrMfDOZRg/teRT8WbxxNk8C6uyhOEIwVEFCR/x
Ppf8NpFOgFWdLA8yMOQjad6Ap5AO3i6HSAz198C/406Pw9obcgUYbcD4l7lvfvkz
PRGOw/GWnGirexRQYOxaYzlNlyzlDxpAP3UStJRseBj0pFI4e7lX/Zm1ULG9Faw/
tVOoHxInDyPJfXD2HzudNSra8M0eGhzZ3iH05hC1zI+dF8bYsQzAZWCtoqKqQ/hZ
D3vTAGgeGhmT2OPKVP9zf/uEqRfWKY6iVg9mtgwcZQEs5RyI85Y5jtdJfZxSFfHf
3HzUGlA1wbyLPoS0aSJdu0dnU6o+f+9mnP4hgf/mMYHWWcFrblEXtB+yat19CaET
WoFWDqtYCXoH6KKA7rUQoIgq5Q6CXYgF0Mp7XgqZrw/p40/+Pd6z0IBJRoTOTaoa
/pk8oMYMhUEYlnaCNcomnv/4sHsjD28lqXpbsGDKhkyVsnbeM9ypWbG0536ev+ds
eM2iGeb3fEXbWnrcntjZubjqpMGZLWl3EBtx9ExThN4SFqCzywXcTlUU1X7CB2/D
K4NWO5vfOUnaMei9/nFS3PBcJU8+bsRyVvL02WHxol8UxBnpY2AYusAb9uA3n9Jk
su0FLZQ6CcbhEGg1xxmWf1IylBEtK+Mtwe2RpoBOpt9PJTJJmjZKrWfM8aETJUdu
HJzX7ZdCEv2xVmI6fZDW8+tyz0tny9I1s4CwA2LvlLSXz6RgJVpoKOcIO9zUGCBQ
dRrC+vAmplCn3Me0HWL/Vp4qcHoSUBm1eEjl1aCiWdDSdfL30bXPhiPV+nRo537J
uJbQWZo13Ji7jqkobXBtvAc5oKB5rlaAQ4+L295PuGz8q6FqGSFN1BsH/BnNL8Qo
y4vQd/ZpbijMOARyGCgUVw2mhT9cI5LEUIRj6q/KToQxWZXKxM67OGKrBEvqQZnF
8iQn6CqV3HNsW85/B6ofvDYJjJqevQQ6r9/w/3ya54arV9ex/2Fdb+ce5UwjgbsB
w0Toqwi2LAWpWCtcSSZ+i35+hGncVXdjExk7zt6FRJeQr2QfJIWtHPWOBR6WTDf7
mCt+8TyCm/1ZF3Oo6oy/YYUdvxnUobSpbIIoUX1LabyWDUZ7fTs+lCrrFwvdfkTZ
sYmP1mvlJVfNZAVJoBw3joZU6UkrluxqINLUPmKpo5o9XAWFNW8h0aYSbvtZPzoQ
Uu2AiOOUT+WAejSzB2Hci5rH89ZX/P+ouPhINgDpnlTZXxkRjRldLEim9PPeZcrU
QAi481+5ZdfDCEbMHOuKXFE5LzGGGJ23ywizLlnGnramjxquthRUkoLqVkscLRUh
5IOi0xN/5WDl/4bpCZbKvi2j4eK4W+meqeOiIDIZA8QDNqxiku3dqQXnTtch3AGy
L6IbTYpH162XwjayKf4KpM21mwMaJHts6XibsGW/IhKl4XuBx5DYL7zpZucSL30Q
2WFgYQYCWk9+JchPDuLj/YG9bZ1xLo1nC79OA9c3iZ5vE7pS/J3bfPeO3xqSuTkp
PZ9ywQQ/9qcFQlHQQnmvOWKLo9YZGRz4Qc3BI8nKYPh5bwPdd0/w4PANSN5D6PSn
pqfwedBpBz2JoHe8aoeHwR8iRLOd/CrkRTvJx81LQ0WgPDDD0meFq93jisGXZtFG
paB4dk+XZbIW8XbEdrN6umktiaF6IcB1TbO9SlWAcHNSwnrJhDuX3dnNPvUV2mbd
4H5J+2wlEPJZGSa1v47vWUb04Eu3KZpqNRNShtBaKJL7OT73XabM7GGfqgAcwCr8
/fQcQKN+y/1tnVN5muH2TXSXZTNkdlM2gZtzXYrkbxLEd4lQSVfC5XxoaMG/kL9B
Jq2j4phfl/r9GKXFu4AgMEM+zuGocOjDvqcdb0cUaKCBzpp4riaD4mWmnhJch7ri
kTUf1kJX3gg23kGiRIgo81r+4mzt5u2Sl0lL4iJ2SQACKHObjbu5yX137p0OkD43
oIpT9wuc9E4GJy63dr3p2poJQ9sjl1GSIr1+XUN7drxuKb6ZaQYTYI11aQFJ01cH
j9vi2jETz2c8aFuTi/Quf3sHEclLhvgtFouTuzCusumZxjPhphiIafvmg9YdHuEc
ewiFr9KJ0/8N9Gkz9bHD9ah5XvVz/+5FbKc2oeYnzCqBqExw8lDnXN0ArasH7e7i
rAODPVyhfxKIUKCMMo/H0JB5uiVFUVuj1qOwUCc+2Wclu4UQZFQ4GhSB5RowVEK2
yey14R2zpyz0UBTBUV9DO3nWpYAZWijGXgJDrrw9kWCfNCYwY6RhjwhJi1gGliFQ
kOIxDNzmtl1BPt6Ejl9YzSgCmm28bgwWfkEhUsZIgzmOGxWcLB89p5iivyEY4kRE
BsjbizhZWnl7iqLMNvLxtl1Ibr40cbvbnorWgY6CqVUYh9I9Kj9fqz3d118YEy1q
3TnnSivLysG75eR5zm5asn/SUirM+03S7wAE5KZQ+wrCeVq6wGpVSrJY1gT0x1t8
L3GHkpkKwNxG8bSkFTASYI0YX6pcr+xV4blp5JQlrQQQUq7lEQ507x+mBNNSqJ8y
J9cfijwAx+mey7n9h/a7rsbkN4TFG8dD0giTdr1ecd9oB3aoPNq7bA3g9bJtDwOY
eA1558FG9TjrWvVhiIg1l7ODs2mNinnIL2mB0dO2xEftjnPuSMFLddhcST6LNOQo
1id6Umo339IjCA8GF1ZfXIv693cIje59hTzHJAAzILWZPwOFL2OtaBKtHuYSnfQG
8S8YFoxc4g6UCiP/zsuweb6ykq566FcAGsSVgRds40IpJxjeGH95Ek7SePTkOlDV
3lbpPfE90wyaD3owSc17XIQrmoQWTfrdpUultdoejZAUkB1RuFB45SbqMvnxf9Cv
l83QgmtUPu0V34xaRSUCSyc/2bf+DHn9AAwJeuku8DBENOA1HEUdtINwDUdRrA58
Sm7hza6IirbfCxs6moIyfym+ZLvkZv7mf0sDxJMW06MltnGr2EM4tm/+SX0wRm6S
3D0RSKZ6yqEivnSX+obiekxvJqnLmEhnDaMYFW6HWf6N8uDpFGeUmbqSt/YDaQIM
HoirHVwbt9sYK8AJlKqGWcqECA0vtVbW+RAkr3Kpr7Gem46Z/fuPB1Oe1/71QAzb
+SH9uTKQx0TlZTm02UdtDVjkAwYe3a8uZTPskgBjW9bHc43dKyOr0k2Mz4HQefPl
lJTxJmazjInwH8kJXzKGBicIbRp+8vDTQBffK4LFcGvt+VQggbQ0JAL65m3ugDfp
g6Oy5xT7tQRDAdKOvn8Ur6VRp1bMQ3vWZw7NX7Gfu8U1MxZhGgjFBTxYg0qj+vVJ
79Gdv1HKEs+Jk51OvY2a21d2zZULkrkHIQGETJJS8NfhS+wZSthQhwmximztqdIK
nCX5SrV+2Yug4k5c9w+jDpUyX4kFMQH3hiac5d1pza9B5nhNWpDDkMeC/kgmNlMM
4eci5mu9qpRynNBDf5vr8Vzie2FldGDODUmX0tDqCA4MU4PvIc/II08v11my+z7w
A06dOAWE0odhQgBp+i9qn8gSuY9yuCvENlsxRc7UQwBDdPtnrQ8wsIo9G+ZcePX/
hD+UwOrSR2ksMOxzBcZcsVI5ajeqXfXaWTf4v1O/HYkrn0jhjIn6gCw0Gs9I3NL8
J+5FhmHd3PZJ1rIRPdVje7lDbo009SpQoxuujH2hBZSSBopPY7l5ABrIjhujZJ+C
geU8h9qQ5CFQYIbzvurAS+qP3kNEggT4xiZRcmo1YmejedrFY1TTCYnOAwDeKuJM
nhJSf8tEhoIT2vqenZJfMZeDF8xPDaYlHAwGdnfpQzHekhesUVZFYOfHCV4FNocV
jgo4uCCWbFFgBosYo+YSKCb37gcgg/WxD6D/jkc7T3mHxTSUe958004MQp1t5RNM
yd+Z8MqrgOwdsGnp0igFB7+jG/2LTtSy2vPgWwaCQIkVS5043pUDJcqvIe7Qvd8t
2sj45F0ZashJ+KlwEcwGoi4+uBpzoaom86F/lOwPeM8TI6WaXVPXnhfzNToesDR8
PZYJev0gbgpauCvRhWABPN9JGnvfefDznCmFF6qOQCEUEKa0fNIEGsFch3tpVXUy
E23ClJlhuGjysDXmlhEX0MUXMsPwjLXGLpR+h6FexYJ27SpRwuW6fp1oQGzXw9P0
vtdNFm5XT/EHTkSQbmEruONEqUUizO5Seh46FiUj0ozjQX7kE/FKcbP1ktWQBsT4
hFveW2Py7VB7jBYGMs9f1ZAz3dp+lvQCAY9W65AGPvpRidzcudOc+rFSRnXxrG0C
iLadSe0bQdmIpyDL5B0NECGpja7EqXJxuYQetTmW5B1vbFL4DoCB6KnbXM33pQBg
uh6B02Ktk1ntDtmR0k4syPQKmBPbCuMY/FnYt42vt4GjQBsFyyn56twb+HD68F/9
YrOzP0qbKxBheG2TGjeuDruGMnzvj2O+0Sa7rlW6dHl5jgy+g0E9Oj+bbTzUEMoY
Rwy7A3wQDIAomDzJMjZXw4rXhLKn+Ch9luGlm7rPcBTX0UehTj/UTQbwu0yJlPC5
AT6gPkq637zuU6fKwmrERyBBFlCg6z7T0VEp+Z9YoUHxoMQ6Udp+LPeOtAIHgwY+
hEvQgaIgcLGKivnTvohTcEknqeCS+UyS+SNFrtEZlfWAXp7WTTifrM6D4Oo/483N
jLSXAExlMjcZVRQExLVbqmzyJ4YMzI7C5I9cpnNpHcXc9fw/stTo48Pls7PzKBPH
S6qyIwshozuM2FobXMHW9+M9/MkwOaSSUbZzYyq2r/6ebP0bHy2P6S4/49GT6gsJ
0q/LRXZSO40zkgpQZ6MJuL7LXdMpm+bw8qKRP4Vy+fKi7z41zmt15I5YDnpFpqDp
ou8BbS2hnrEoImU+bdTYX2Fiw7P+6wlOT+J/3QGzOMPoJGOtvznToGGhn4mP4AYi
H6kmZLoue32gWBtouM6GVG1bO8JMMMv2yswxFCe7QoXse7yLU5mFMgyae9UUNrzj
AAYweVRkaIIp3YWE7JhSqM0H2++Tk2GzFmGNuEwqJsqTq6J1sVqIsoCX9yBukvr6
s5OGnewq8FDo6kpCeGM9cxCqmyapfofZM5NbmNBYOeVPZ8/KjNW7SzRJEDaJNu2I
MyDkt0G6sQJ3KKZbei4HLFM2lVb76ZhJJVVqzpD9SRo+wO91DNZqfwa34KeWlE1b
PuyAtewGr9HaSroqfmtNxsk7irgQ/MHMY91C3TvOKRQN8Se9IY+pQcaLTkfp0YU6
ww0nGlSScvJeWVz9R2v0u0E+IOx9PBcDWrffCSdaLSWuW6GYcPgFgVbm4ZqM5D9f
o/06IPJizLXULsVLza7AuvIlV3SWN04iCAUUJcUtwTQKTTQ9hTvGteIi5cn93nK8
cOlpok7oPnYDJR/cTq/DJYbCJukGQW+HpHMFymvaen5RMMTt2ysVF5P5iKZWa+eE
vdl1FR3uT3dsXhGFQc/7fOUpXiIjYALZuv5gxzYz2VhqXaLM9Rrrn50H/7Zxok1G
x3n80usGOStdFAwbtU/CZI8AjbEQoENKCg6FeZLmCo1XZJzwWlExy24ajuiNMjZj
d6ZUecnNSmImLU3oGFTxwzVL2ofSRoOqHNVeA+E3YdNbOnT/IDTRPnR1o8NJrHvR
8cEmzi3Cfx0tc+h38CK3QL2V9zZo61kosigFXSazQRTcaMgsPCBZ16EU/PfkztAw
2twzCw0D1nO8CgcD+OKA7W6ky1r17oGsYOYRJojB/8cJc98N2RbHjTXwl2IC3r2W
b2W/EKWPM3FA0CofhLL1sGQJp3P2tPm88jeYAGCDS4YTlbIr+tVI1jhCRN7QATAp
kBLqAh9dLZKwC1/8KVTPv+d0Jv/P4HtIWGR/4n2LXKFOZPfkk0kvy37IY8F3Arxe
aOtmtdnzlvqKUNgBeu+c5/I08+stPAY9rQgttrvPLngyZT9wOL4I+up7Hj2L1LIX
tIZiK+UryvGB+auVnlL3di6deUGob1rDr0Pqc5pJtX8ZegSPbUIoRaMnX5jfkOTi
CB6X9BAEka2AY/7yOa2QPdcFhET8XCAVVdYAqOLsddDzy6LsLxz3CHfXfdtCVN/l
GLNqT3ZGDY7whfr98LKrKiVoQ59hvRsy4UZCr2flyJl3AemGdkBxR/d5TENGMfMO
uHIQK/fRzWFR6An+eAKeqZRYPQLLZ84B5P/izdC/yprfVQc1+aOmGF6viy94Lxyf
vv4M9DBNUWsjBVQKq+9LUg3BG7SGzYGpxN1qJMPsleujmgRTnhjIkvdnupLQRKNc
huLsFtVfuZPRZDV86fhfksusMKt5vZANJAyF719H6r/bEpsD69rhJa3qJMit7xHE
UMc9pjpsRamXIGtp4BR80M8dNzSzFByf198HhmvSpbGhykFgg/Dh6+7O/2Df7tQU
ULqDHQ7mxKkFygnKA/fXYv/1AOaQIEgOABoQEKzbxtgiCOnhNioAwKLjDCeEO0q4
8umbO7cuSM6tz2jZ8tAbd5jtBgE5Sif4428ks9x5Tliz0I6xwshLGIC5fnQvHU/s
zbflf70f4/fQVgw2FF8AU/uQAPXf1Qbf6GYkiPl5xOcJygwGWzC+JFfYDfFEP7Bx
InLNQxImCVMfaCxBTihyS8NToHXaaRk7V2XgofpdpSgpFAKEPtvu3/2lp2uVlfmu
Xqbkb8GY+n7uRUmCvdKLaoIrY67OFi8+ExU1yR0o9ePMEYfV2JWK2aat+6qKENn2
X9e1gRPS8bv2rEguuqBEdHGmi1HgYcDmA7mAYHXrM/Y7qqFC2YiAASySVsVQRPhL
aCKn1OhROl5HnzKt3xk7G/6PvyD3RPWlOupORwjz6JursehGaIAvKdgKzd2gp6we
GpPChEAPy1woGYhhVYwp2Wq4WCubaooNaLLX8jeb7P9zGBe9iwhTaTW2o/yfF7VH
5oULfhcPbSjol4rUihF8A6xAejm2qK71PArgOAP0PAKbjub2qFAJm1b6BB/rBOOl
Q3uqzhNYjG1NDgIgzJREKVTVnogPSYEtdcX5AM28OW3A2vbgFrzRcXROgjRu3o7A
YKjbVIsILW3LLQlKcLREAcPHjb5+WieOXkoqYL8uHtw8/JGPyLLJFo+Yvc42kubD
IzucjFo+67OikFbl3kx8TUsZxgI12o+ttITAGoSEcnJlUHLEom0PxCVk4/KoAqyK
kp6C8K+y+Y2pF65+90mGjzlxFnMPk3QbV1iVbPJ/ncn9VYwkPM6iJIxNa8MOAfp8
dm3JIgEQFgAr8DIrdWDy5mGOF2+MspCMC9nJ9ZPE51fZRYFU8t/bEMEMl3qkuBxJ
TXBXI3etESAe1Bdr57WSbw+YQPa+ipoPIrfbQgtNkyXRR9FfJBOa4jF7wFfFCLd6
BmlgwTl44cF5u3tjq6og5KWHyZ+GFsFhNPcybs5TDr3epmmH8ORscalJ9A6JWe3/
OFV2Jk96iMbwONCFzpCM5Cgk83PJ59NIrV3/6nQQt65CZcE611Rv02YhwyXGxVar
vTyBof7X93Jd5ULBHc+l6IZHWzCkhd/CRGJfkRurIS4Vij/4XBgKvDHw0hqkcjW7
6r8SY5MgcGAFM60/YdpRgN55SGdhOg6f/RfonUjl5TXDrhUcPYHYdKB5wTJGnSIT
iKci8+5eY11Yk0LMR1vcUItOMvcPOfIQZ/Vz0h4pzftjtQ7rseAUWaZH1oHTf25j
YGU/XMd14NvGSR2YyLLmAn/VrtEhnA7Y99WXLZYciTA7zbiYWvNL0ZM9UYYRJ5fJ
BIMQ3eww8TH9J+lzcMCvA0lyStz3fLKrV+jTJWedh8cbqO5dFfKVgP0lbOTZ3f7D
O1JqYI1CA4KMVI+YeC9TbCx6BmYn4c58Iy1V1kwG7x6NA5NXewwb2yEk63qx38nQ
Lh15qM4MlNtbDQ4CuZEUQkAR9SaA2JZp+DCtJu9h1vWSwnB/Ke8QaPeNLBYaJ5LT
5x95Ozw604UBlwUF3KZI7siBrkhsQmbOOzUc9pWHoVWHbe+UBNcfCsyHV2hsJT6w
jftiiqegUwsmrnCu+I3FRXC7qGELcVKJSBzlu01mPjLeH4CGRZ2NvG+c5jvRsSWc
JGQO6Ow6wsuYlpwYvV5inieadfTJOTRmY++N5DZn0hICaXpqazyNHhmGTtyq1dgn
GGW6lw1Exql5R59HyqIG8n803xHDREMjj3yREorHtRe4bBtvO23TbRJ/6MdE8A1y
ABKYdR2VFyQqH0nqu9EeNfrjV9UcYuAD3hAKqCj/iEwD9Gj/rWHXtPa++9/E8K3i
o3vK5SqBfeMq+RjYjPHozt4lgUyftUH+3TYDVi+GiS5GVLKkD3By7nbM3crl5gsH
KwTouFcWMLYS1XCvrTOV78VSvdIeDd5A+7kb+ASnnDZ9TvU1d0Clij74KjC7Fd1q
lkrrCtNaN8TMg5onw+/nh1LjrdNtO641RBZGEhztp7YEMIZ+5UghpyyuzRpZS0lY
7NYgU4tVT0RY+Jo+04nTIb11jV4IhK0FmgdujSQBJJlBV8ixOSQBYPKbFx8m+xj2
YewskN82CX32vmTRetidy5e4wY2YpYEFCY3XqwwuXD2RITJP9eA1zbLPVO33IC42
8P2HVAzCumYUyHCpsXOl6OkGYpKx5z46+2IdGheaoXri54+3XJoUv6+NEP1wyu0k
N/QGs7T5vvKE/gO5YM32Q6D0PxN2jp70FcUi3VgJG4HsWqBSz4QinX1sljfoRype
B3/raXJdYUCgtoeLlIxWMjRfynbziQzR9zusHKdBcs9J0dyCbmG3SNFccyaWAxmG
HAkSCHt+1/pev3H6dlpcyoxZuzYhx4lZKHQRipHUjM5a1KDXj15YOIvqTZDe4Hnx
VHmJHMdeZEQxvUIMzP4G2YOapgQ0tKVEKeFKnCxCgi5csTyUOK5/pG1EANxcNjEP
vYrGHCIrC+4vtdLcm0LGDUnNeBVp2D8wI5LgFtedo6rZUuRB6HlPYV99GtCsIXgS
Ri+41Zcunqt6dZCLJ2XzKbWDANTC2Zb0/gYKyIYKYhlCffNcHaJmHDRFezXoB3Sn
Anqg+yv0bpnPsbsDVPYltERdcyhOGkOJPr4jsx/7XA+xhK6rWmQKYz5HIIDvMy73
C0fEqwN8oNYPzHINf19bEPjW7BvKDBQc6TO3N087Zb+vDoVa9jlRiIzwc1NUjK9Z
WrgumyMN3okDTqt0GkGLaSI5V0/WVINewN/540eCbQ0mdq31TXA3QU2Ans+fWell
/k1oZHh9leVjVUxO56TlKh7uOBwlpsxfL+uE7RsfFUczYhoHTYerORwUOeKoscuz
cbkNkQ6lzdWqShR+BFoiYrlU5qFxBz2sJMeJWqBWh+TdW8ZfioWrqE6gpNPN00F9
BAFJagxbjp4hPBP7x4kpbZi20gnUadfN5zG+sJ4aexYXTOsL20z5qA337WEdajl8
StmMap4ZSdFNZ+eYBXQSF0KMzlHi3QheX6LVuTvk45XGqJ4a9z7M9R3RsGD9Ut8Z
KO4EMVGBOdsSnU45lKH4yFlWWackKsj1DKFYAGYAhj69ldNSV7TTg8Qjdt1Zvobl
pEMejutkWWzXh54oKx1DUrZplpCSQLkr7V9k42p9uUq1wKQpdzchCFWgYfdx3MO6
PG8jvXjJaRLRTevm0tLkFQ+cnz27mydcdUBfTYTuXyEDkEmULDIY3C+exvdnxndp
nDuhPzeSVqQTJbxBqZp6ZcV+Ev0fnT+WZPu/VDxr/xVV+yhbk3YpkwZrGCA+v+LS
WwtEjIMPg21EU7ll4GDa7JKJwfxejEgLpA4X2n2TQncL6RfVVnT/9IsPuxZgmpLX
9a2XBb+BB5AnxxCTTmTnXWGGa+BZAwBfivp1A3Xi8/DksuoN0Kxkv9Y9+JChMITj
6RzDSBkSIEmtOb9jHodbygUzrNv9KPLy8r9Z9uiUa/QIUizQsGn3WNe7W0oMOx+H
fZ4P1XJWbPc+UwydyI02bdWENhZygLgKyNDjLXAFK9GLCeleUVPb7XVHF/9/dbpm
iPbvIG/OSOZ75W1GfkHpsSMI7mzev2Fen95d/K6S4qYXSkR3UlogFg2F5DVT/nXL
xl3jFQ6LvbG8F1fI9Of+d5DcR1rwPow4VpBwuGQjGWe4E5T2PnKV1ukjsRpwZeab
qV2yQA6uw6QGfjXyglTUbUxOkLR4l+RoC95mRgiG4meLtJ+MihIUrnav6WHnf2ot
9yip3zsD4oDBDY+eq2GBnoKzgphK7XTkIioz80Iv5B7kt7oMihZiba+4C1ycxDxX
4ygKPO4HrRQnCt44z4R5wi4H9C9wCFkWr3K0Hfmtvn43VZHgr061OwPgJ3RpLoUG
WcaBXfE+o9H+cyvDVVFlAlsujvK3oq7BQ7KMhtH0HCN1ix2toRhCnwDweZfEzPtR
PvZPhYLjDByCBAGzVJMsimoHM4Dx2wt57N3plbhsuYnDDc4/Jx3dElcj6txW55Qm
u6LU3dPPdxp2jhmThqnes7zoWWn6lJ54JyZj0A4bdCDkRCWqovxwUwjpxiewX1uf
OafbkLhpHIkvCdSNl+Fj6N3eskyOMC8u6pxl9noUO1OqexVFLmkRJS0kftV9O8af
aYLChbM8V3872klLHjzpiNxgZsi4/w6d/K8su+VGhvZS6l+C6MOmA7XLR2u9mJ0t
mkA6QKcHfeum28t2lubPd2iZPhJpwmxCny0nTfytw2A14LIioCy5x9AT1Tr0bevr
l3ranRtixwa5jUJjRTRmJ4cIzfJHuwTS/CjojesGHc0t2pRAAXxL7YkU4oIqD9ov
gLfDP3vjlOWQpsdnE1eZ8Lnk14cei6EJJnB/4DmsLa+EnCugG9oF8TyZwnru8bhm
XwwAm0VvcyYQn8OslkicmQY5OuuMSi53b+jnA88ch7ACsnoDA4hcZ3M/WFybME/s
iTiMZ/3s2Ck9Tl+SOykfsdClVsSSxeoe0r9cOkVNOMqsm+WCQhxKxKBGBPoHIMAF
bXHrWK2AMXGC6Y2X7/iT0cYpY/SNWxRziDzaaR+SQ3q38H15r8rRWU1HWu+l8ktK
DEPwnzi987kwYkOTM4/61qRnIkq7icHV02s9U7gJmjIjWYWGAdULDI8yB1a1Ik5Y
cXaZiY0Dd0cVnfHC7ZC84cko3tzAJDYTQEwzpS5uIDaxXMNYb5nk7i5Ei+06Fz2n
CwbRh8+LWmTS2uVnotrG6R0E+rJdUj+okQFp9+iCb6u8FWVW2IxEXLf7k2FS0xA9
WmOVQLeyMDb8XmIZHtc60ynPZWYtb53boRPDzigxIiBKA8UiyEhkPqL6c4abnPUC
UeW8HrDCoKPV0qYOrq7MtLv6bYLEvEyeO3R/AHchocHF7A85tdYr6u+GKv9HYHkP
WS0iqXKaCoxF/NytVTfQhLBHU5lMIgAgkC1TxGFJLHmxslAS1SFdnFVrAFmTHgcP
4cs+bgbRW1iqVT80GleksNxUEuJ7AC5bOY7VD/PUag1Kzx6UeblYV4J6JWDqZakr
cJhsDFpKtCPjx2+3ie5fp/Y19W3uVwcTq2xlw3pYLTe8uUBJLZG9Vgvb9h8XC3EX
uDxU7NqCOi+O6jVYBQlTfYzJi0QmjOo6ljCiJOx4RLAkz/aAOHf5wBJ7tSR/JSvf
86C1fTC5zsUoSOKXQNsTi/jvcN+UmanbiybDL8lenYHaMZiK9Grw+WwAa5jRS6pb
leiFiPwND+D/LCmigajIeOqIxeT/mCJ0+ouPKTjWbLhXpBJ/xSolZfxDCOB7RXiq
eL/Mv1HZBnk9F/PRaCG0C3oLFw3S1CG6hDyIz8OYMwovvYX8foLSKu1BFckbfpeq
2Qa728Ylid6risX7ssM6NLvsrl9g3hitKbjq6FOmtI8Ll+1+cK+gJH43Wy+WRCd0
KR7R5YiRdTEbOr5dO/dL8AOv+ZEOU+COdviHKS2d0Ix6kPBRLwHD7plrD4U4+/mK
NI19FVdzbVgnSZtNIlTSqwP1F2NbjQpju6eO8BnG9L2WKm+hMl31ZhtqFOOaI9sB
ekNnhX3b7gBbWdAS0Staxn6t+0C0wPO8uI8yp31rwxqU2dPrJGSp5yqCbMwKQ+NV
44nw7EJ1/kPYpvZ0aNmwc0afYJSmDV0rPEsc7C0ONvT2BUZh8wOb4G11/y18ac4k
MvRE5/DBt0G2lmX8KMUMXVPkzhzM0wKjk+RvLxsv8sCAaxF07mHfZyDEUlrx5ZAO
7kDSJuxpwBn9uMlRMTosu4oNPN4QsG7gOE2G9juErfRBcSTBtvW+Chi2kIKlVhFS
tQNLKc86J74YY6L+YwxRjFAbXo0uvQosY5JlFn5DHWSvMIQa2YqSl6APMeN5Rpys
oQTzGadzr2MPkmKi4UKrcKsSTY5OJjNMZ8DQoVl2uNchofKH0CW2vgcJP0GhlT09
om8h8dJtUrfIyVigt+DaipG/H8cIe/zzkn0vO2TxnK7NhiChrr+lDL7fQiXX3yL/
zS26/qCVZGY13LSWaFK3zHWBitydl5oU0seUUbWRUk9KDWoL4GMa9DNr3eYEQxHc
K45Vf8wf4NkfIm3KkylcHwPnoU1X0KnUY42JWqiQuq9GY3XCp038cUUQqLBg3cZ1
a964DprZWjnL72d5ywQYOVMWGH+cXowmX9TgTBDcZTZu+//mWxtOyKZyIRJbErj9
iwgUvn6bEnBE5FkfdpCTXmg9J5s43pvpuIDzURtTaR0vkZeKusCK96B+g75fPwuX
/av9TPlNIBsP2cDy6fXoDwHY9yoZolDUoQbr5cuI+9QEgn5KEC4CSNazBTD15o5f
X1SezqghK9+irzSO2fFS75WaWRK/Es4zHqi7b/8i8Ww4kapkcNy2uCbwFSPAXWXk
JEDYjxQj8bTMXwb7VHOAbF38zgv0HzAG7M3np5KX7PHhI+HPBkOOPpTVD5JJ9DtY
mrzKCHVmhWSVjopJZO3QbdhYtIWG98U9C0VCND1kjzkzVhw87J4zM1WdfwtqNg/y
I/S+/Xl/NFwXF5sQLo+XCD23O2CPCuoUS5+BM3JxtqIO9qs5RuAX07pBxTMZbmX9
xQP/cN5tJ4YjW++WM0VRTBUoFTfYyFoCgUzHG7eakmlNKmpRRCQMLKzdsA6zxnyw
5eCOiVvtALdIo8sTlbDihvf+QXivk4LzcW4SlWgVIqKWlhwD7JJ+/xfbg5eguTlU
9rdZHe/soDcRYQ59xlUHakCTvwYmIWfzaOfKdMO8ZHL6/6UWaT2vl4ozg3vj7tyW
UMz9JJMib+m+SrYj+IixU0PMku590mfXZEofeKd7G6RP8/gBPbLBnbDSPtcwDqyv
JyFQQaTPnGSWjiPegrxGUDx033qlZjFU6QWPkgJGNBWm08ZueWAcOZRMJeg2eKrM
LQuUSgswmqrr7Cgo/YE78PFHG1Eu+4JKuWpIB4uppQx+9PrDFxIv2eLjtzRzJSBJ
+cSOJhtg5byLszOy3X/XjwhOtxD1nrI5atryRuglo0HYxEc0+jyT0BblFS73MArB
s1IlAaZPL0i1l6Exy6NKcPO/j+tP1Bfrl5j6VXnsVMCtevf1XXXkxk75e22/fmCy
+b9vAxzFpZ9smGuU1PmGQeylQ02h/puWdOkEDs7Pp7iykcaQG+RFJUdWfyGhwLsF
QNaMSFo+EALAJN4Z6wrSGr0sg74M126ugHLsYQjyy5bZ0XAPCLRxBWD/GXi7xgvy
nDiMmyo2xvqafflZ5GSa1ypai6sTr+ACHXvPFa4E2Kn/WY65z/EDvpBLp1pyEndO
u2aZtQ6Q5SxNcZ/oCaaqWiMncveI1i1Hvd6GA6QzVPONA7mkAnGIPe5pPdLiaZct
V/DaztMme0zstTWfV/9H2JUb+P8P5KX1t09J6YtvmiaOwQlhRzq1euliEyYP2GeN
44Euw+GeesZvu1WwXDAzVqnfmsdmQVMaKvoWJ5GTjQ2qWBmgXGzcIr/on82kTBdv
8RhmEkKl7kWfrNe634rBzjFB9+00M8g7DLr7H7FcOCLY9oqthIwe2kKxxmTnFBPf
/tRJAOddD/axHrrm3jVpccT1bNKuDSn+M7fUajesjl2m/44HRx0zvfEkdEzez+Th
as9YaTpnvbRORqjjv8s4R5rNRPQ9T/2H23J0v8YXGMhN26gGVjqVlA1gSSibQuhp
52IVK6Jwh/gUA4YH7WF1+SU2+yKJebfRXi2f8avDthw8C6FTj4/llNW8DvUDCsvD
kZTQjJkEvYF0GNGqPVizH1Mp7LglArrYXKIHWDuljHwgfQIgnjRvSPijrH4KI61I
px0HIpbuY1fsxm+sacVFZfwYYEi7NcD0+excs5hhdGQDAM20ilrOvDP+kPfkgXQW
PLa3cl1xi3gtvNFXeIovwPawBVh2uIoFY4f/xu3es7TKQVW+y95fG1RY9mu3jrLa
BPF4ULhBBmPtzhCTayfJ+iBfFUpAQLNVxn4KW7WOigMTTRdN2qxYfheNZrx1/HDB
18DctnGmCsnEUvxxleU3Ps8UTQRvGougOkQsKcOMRSc34fx+0uP2MMvt5FuAhL40
m6d872W1LXWqaC0sxgMp/S2UWC2gVbwC735HWMmDc2CHaKCsYdad8M46kv3fhXZc
WwFOkPK+eUH5asjgw46Y3iFsafepTPPlzNvTs2lK2gQhYaP1n4SfSLBjla0RiQQS
Kxw0zW1h+HheyHm6XrF0fQqs41c/JGFY+ZCAfKI7fbrcAxMWBDGFWhf1W96c9ZoO
m1tCxjC0Zb6KJqE9bVyIx1sf9KhHZ2JtXNI/cNCcEIq2ybxDreVa9lx6vlASdu4g
mlz2wk/tWDiCGfP46pKXpb8JbhT5hxoiOZJ2TeU9TZqhi5SUIg7f34FyODtoXh3W
DX7ldOD2ulhrcFOrUO1765J+XFBtdcYnF0Va9yXfewk4lYMCHSDwoEfxWSDU8lMS
YZptXRW6lYm1jqmvfE1obhJtP5R7gyyrg/GFq974tVo5LRUPOFuxk/upNhyKviMF
HaHLH1K/yoHPCytTgH7CcELFOxzZzvr/SpqE3EuHNHP0wA44GP92y//TTu7Ww8AS
bVRXu7hyb2829SYLRclIEaZ6QacaA1pA7WcZdUH8vkc2uK4xOwSe0nesgK2hmpV+
saik03WzKp3M5YqEgZ54WhbBxO6TkjCWMhsraGVP/76dU9Ev5qVArzRCjzMTCQrN
GWMjwH2De4IiJxZyqVFH/zXnaPMPWAkGgClbdENKIt/Zt/qaQQVOx72WnV0qBRgF
nRyu3uNEICYIz76mQPN7UUSK+GF62WvHyaBlLAcU3EefxCxdDeFwXukQeC/WUEIA
oFb/2CoFxi5kfH904Ogbw5g43DkQjM8Ejp6laUXRN9V/4iF1aZgZixQXt2KQxsWo
PvkAWs8gAI3o6oKVU8fbWfPq2WCDCG54d2vwrmY75F/u/IZqSHSJ1xYgm13P0Ims
EUO1EGYUFa/fZ11nWn85LPlnYiyKABAMJKI00NBNaS1Hfr/d4hN5U6iSriP47Xzr
/PEOqB+9BdEaYpTcUfNjQCbZvgPUekPoaEHNf0IH5yvBRGe2LqGr+3fD/vT0L9pg
pth8lPmw7qUX20zvSUglLEug/Gl6Sc/u222eKvTJ8WvYlFEfocwKUCBdVpfwpROH
N5AgNtUjV2PFPeVf/zYWjKIcKlnnDeWMn1I2oeXDMJS7u7p0ixfnYBd4/GiLS0qH
0knTL32XUGwKJ2qcjGQ9iPl5qbUtPuW6NBLGHPw6kRJlfsW61XsHc76E4e4WA4ho
8iWtVMNMmMlmbsX2VdbRYHI+kKmMVBJDuF2fOKamUwan+IHtMkBoDGnfqgt4QI2A
cwl7/tW7wo2u3WS+f1rj3ANePFo7p3OICyjW6N7wt7PR30F0Ukr5VfnEN/0qRtCG
JWE0L39UtCnQ9F8tIHAmrf2rImoMfGT1+s7aOClP45kV4VAa8ITEepMh7fASST9S
jL5O/8zu1oh3EcbeJSc5/3OIdpwhS/5/tgs2Y+D64WckjG5zCG4yvL34Ev9bUf3N
baWWXqIUu/bh+jtqdu8CBLDBAQ5/vy9OxQ4PenwhclvW7ZEOQrTmbsTtq9EuZbig
uHtBh0fQobUoIbRGcjfpDH52bFhdQsb0pt5yQrOSNsaXiNG98eWxdKbkMi7kt8TQ
tbS0Oka5QdbdslY0bR9WdweDqgFXZ5g3Or01F0tPRWd6wzo4io0eR6SPh0qAP/n+
W5HQuIcicF2bFTGWancnkI/6p8Zp6nDvunfHkNa3qRiITjAq3rjGG2tITtADz23E
HbnsvekZL1c+qA7ffdtVpPZ2oA3vSQv7tlk8VtI022c2r5m7TT64n2CHNQDiJG5M
4Yaj86olfEdzA2rxSWUB28N+avK2nNVZWijp3BLLeAa7hKYE/N+HEo3fYz3dMj+5
FIBHL5l68JV9QU9ifKvtHr24w8YGoEfNSRm8jgRrvgCNoniTftxGS8wUYPSV3PES
W+D1D8O0Jvz/4tLCoUGHE26CjFjQJYxZ5qw03Vp8lvb1ZpENN6hePgGUqvCFAgaU
YnR5vTNGu+4vurFGSM6ud/INjupFHNaCYa4ohBqZH34zEYJpVffsTbUT6B7ZObEb
ANeXd3+9u3SFQIm3KZkYJ9JuuJgf7Ak7+7xHPyWwt+dgDhF88dI20pH7dACVz8np
pNifWcMH0j679UseukdrBTl5nnv2Sr8UUdP/21hsSREb+eMlBS/O784xsp621GnQ
PUGMiEGusWbe9BBZmj4Vz1K5SPSZOL+ottAtRh2Jr1f54vzBO7x9RGfsPpu/1gB1
uxIN3tYEo/2K9Fvts+F4akC9jWMLIpCgH2bp5xpdEFKP1i9/fR5ZG+JtcrXyk5LK
bxez5VAJ/TJJzVJ2UzyyoCFhwngYQmGkayAm8LDwYQsR0ORMN1VUCDRrah5JGQ9Q
3k9BYRsZXZGXI85YrF7Ib6D40NGvqwRgZdzd4EQ+N2oz01aBAhWiofaXKASAPGXJ
zk6f/fM+32QSKYwKpffPAhU1N3JCl7hRfBabsVqhcdGrZpUwngxrTo7e4yu2F+Ew
M/ugpB0TlXq2b05BW8zF5J25QIQrro9oAucYdYiiNyke0ValBLjrW57Yypou+DOF
+ft7KH5NGo1yuSauWnDNmCS385i1Ui1ns6Tq1p7e0UfNNSMW8fqafZ5WtYD6Dxoy
/v20r8gRvGdgOdVAQ7ilrxl63wDxVf2hqXjq8zJAQQgYey52hCTkgKTUw/erRgho
w9AzIjdSMx/2QWvtkDvo9dscnV3P+fAgqzTBdAFyFLRUZbmqhGN4QUL67P2dppDk
gBt3iyvzdmES5yoRKtL27uZRxV5HBH3MpZ7asRv16phHTgXKJqxbgwcRp60P62Wj
cUAnxRihjlHGEr3pSpu4MNal4GFaQTZLKoPRgQassdEW50+85QlwGDLgtZFWkH3W
ilXMZEwR5lHiUif5h5uWL70og7l88dq7xFPh4E9dOOwSMA82bL2/lFz6PmlTPZNs
+eSu76tr2aNTQ5zuM/9vmzWb2nRb2LklM1kb2v0o32nh2Iz8KIL3hzejAbTzD6FF
7TR7rJzNR4LDQrkHprGqMr62qGzIGLUFVoCrYIWCmXKC6J9tidkM1SX50pMDZpMM
/CmUUMBUi8AE1sr25H2/41LETAfL8nyj+eGfp9Cfgl3B2MyFpCKHRp8N4eyhArQ2
wcnzXii7rOoqbiytkyvpZbXYcxJ8kNPg4DrGSjaCPy+xkALhzyCJYIxK2MVSMQ4E
4uRlIJ5ge8PpsrMmVheiUU0Y2qpenfkysZev3QCi4NrvwSSlBn26fVBAj6j3BEAL
EBtRIrYKcSZLqUQDa/wpFpaBB4peiRrV6JUXgg/8nywxSIMsJ/lIc7EMw/lks5AO
9YxUlebovhi8vF1aslZTdziMwkbr9lSX+xMh5Jg6MQUQqjizJZZa0wdo+bdO4RyR
oDYQ9Zpe5q9yYf5XJiWvU9qBvkj9HcbxYEdE197S+chnMllpSQ58hPDWfrfTkl6d
U1rfO3cCJkyS84ji6tdRd3gc9CPlrydpvMPjCoz13n/qP+S/ShMxFiG4BD7tkltT
3Y5ZJybQFn8QFTJTTJYQtrxbVDGb+lyaBBRzNd4jM0zXqT+Mt7RdJcpuHgvmeYJE
W2c8SvxSxkHRz9I09/0brE2tUA6g2Nw3Qz2JGB+8I7H7sy5qTiOjMPxxe82Z4FEm
7vv+U7wYwyBNEmZ26VxS6HYlTDuT8PzwRkJOMLh9/fTZHm0EyzDGVYKlK+nJbtun
Bt3WaCkcAHr3/dMYLLa6T8H56cRsqtW6IH3b0c07nrS2J6HauXAIvBJqbfbysUQd
gpx817m+MwOG2Ot9FSjziDsyE5tAsURq4OuFZ4k/4JRaWjtHTgpkdMLoZEL6HYOQ
AualOITaPl2n9o8/1zPJMqGHRiwOicFIGszBhcA9sY6CGXGrJ05dNbtj2C1yNimK
jWIHlVrkETjuHut6sHMpWNFzuHmSVgPagBZUhmdV8/NU81R75E4tzWS8eGEenVKj
MHsxYlwXEmNtJrrB2dQZgXv/z1/uTxYuJ9k5puboBlCN3cRxSuiSfmxGqeVxWDK2
ZgLQyffuWGho64LYHUeBp67daA2J40rrGq4qqhTe9CStS8OlVgPE1SVGba3MgDFL
vv1zAwbJMoljIBbICa8hGhiFI2IhIhSp5L6H0DaMKdvIvjC54Sptay1sLDuRk2JS
ZVnVGplALJMDhLWXrnrN5bLuzYbi4HWkcTQG66N6sci0sgfxJl/Tr/lSSz2Yis/L
k1ndPtLvjAu0yUVLNFc3rM69fo5E8b2+x8iv/pZcU0QZNk5bcEN67TpnR27gPTTz
gnFzuuLq0lK6w2hcjt1ldOcdK9qUtNBrDKSGaNc79IGg8vSW9btHgHvSnMDI6Dtw
KMzFQV4LvUVu15ObHRPyiXyDnVTp2SZ/9L3AiDcBHDZDKdoZgTTlh/3MYvPT3Z8i
p9Wk4AkzuPeSzeFyEd4FA9D26V8KvQBN55mmxnfOzIsaQ/vhZLBY1hWxeTqPF0EB
YsY0YER/gyN+dRUmlZsvFrcwchVhZKL1AQ+hwu7mZ0BaK+jJhoAEcNpS26BxUuxH
XAhgWwth7idMLPfmkoI3SPBXO3RrA7qz2DrRCUZ2mhSq+/Qgwf6OC1xDoXHfFFC5
azku+vZepmlSYWVl+aqk9uOJCyRoNay8ODeSds3nKwzZuiQTaSQ+aWgPz9hEtbXI
3hhl7wnBM8HdkuVjr3aDmZUB7P9xiYZ/mQ6cq6Hf4Jzp5P23DWx6qkdSNK82Ovpj
wP99+DgZ47GFOnAJOFRBvCSztVHYatX9abU+YCN9s4yZu9d/wwyNvfDSsvoJkLTj
j8FwO6+wR06l9m3Se5E5qcggsmka4MiQFKho+pNKY3QRBtTBzzfoZq4RIfV9bIoY
IvtRzbLg9IgJcuTDcMfOSJy5XfpwToKfppPDUSc5SfPZMGMq0ZJ8WyWBd8Kk2Aao
kNuE2o8C3ydcBacOEwk6L0SV+eLzpLwXlGC5t/ZJLa/5HsZofshSdFfMc2QaqS0W
qGJQc1tFnudLSgJVV1Ta9W9IFiLkFRj4vmbkjB4tqgKS3d2A66vE//OeiJlBOlx3
nG5ZEI0VhGbxM49tHT6IznpuGEZ8Axtcy8/TeeV9IbGp/dlkLAsBS5hxoK7qZzQP
jRTd6KJYlAIYHTS0qGMi79P0gWlRRpi8Bqpn2rAqaWGv/o66H5mBBovZPLZtY5ib
wyFYA3r51B00lBKY7wHSasE1/6B9KW1l8N879tCjlt1m60CH9xf1r76w3eXsfTIl
2X8fV79rpLanAK/WKD+UVruyhV8DZK57znp47243LGOGRvKi2Hm7MVh3vO/u6I18
IjYUOn0QfulfeSavtbIARIS0zXKFmEFpip9IHtnLH2EQkJLqOcSmAvvPam5XEkC9
HiOTdiTfxE/buXnodsAj2yn/Ptb1QhOZIhpvAZHHky5abBIMPy2GItYdkSJTRORk
Xm2nIj/SYy17yEcR8JrLiTTLhjpThydI2iDJJa15FBlnM4iHVOsvyi2sM5O50JVG
V94Ictnofsnxz3fDu5Ww8C2a9ovkvBGl79IYLU5icWUXVdtihffirQKl5Q46rq8X
zTsb38v2zVxCcQaXB85u7AKjcVlnkb2rIHL0/GFDNDwEyyAt883f2rwFKLokToG1
bkGlF3sUA9XJ7rWdZ7Xfs3OOoAyOEjjr9spz4EcEItgcAQAIwr8EqUY604ACDN//
OQZdGASBXt/Mgy9xAy1qGeWm/64a2gWfwvlQS2lvKRLjICl31afrlEk8XfcETq47
+crN47VhurIJcX1/g/twiciteIdQMd2qWnVrLSqP5r7y3ZfA36+53o99Nr2v/ixs
tKRlj092vcSMYDiLDw5JPieeJ66UnmDvAYBNxMXSB9WAisteMXPNGDFGYW2tHqtC
SBKhc+uUbkbnvQbxWGZ2SJKoL5q0Fr2ZbdCn1otf47mFR2wjD+x6sJZOPFL8HYlZ
yOsD1MAFgAAj0W7dSjQIfFmdajEfshUWDZpPTYCaxBgy9aNIIlx5N5vuaLURDQXf
/0yxA6LnDGjtcxIhv+JYYpcSGRK4jc4IXdLxvJ2SJLHt1weyofniNUXkx96CdZ8d
sUPQH54TAIYd3BPVdZXhXlGyzH0JE/tEJoQtG22eflDOk0f8vVq8LZI9P/LwaMHi
ODXH56vMF69BeumWqVwG1RN02ptiPKVHPEWSyg3IKTur/UOLtnBO3nJtGXKkDnJS
27SEroPspHVMOLCOsESPNoXyUjasN8RSHyoFHFWV2iZqXEj86yI1lEHbx0gWRII5
Jeik8/spj0s1X2kHX3DR3E54KWtlHTQB5QAoFP67t47ZmX5AJGE9vRmXil1CX+SW
63IvW2GA7kVoDQpgxy2Qi1FIfy9m8UGO01XEhQIZwTaKc10U2nLXr3Lsik+0T/Cb
IRAsTA9gV627XqPkgSgkjwthFSjUv52bU2nlTiNmAa7RQpUa8G3D+IISxYvmOr+r
/bVq2mKYPtkUfE8oF4hvPPuKfAeeIZFUPSZYOmSdRpd7Cu7wGZh8Bvq9NqPzpGJM
MLm9LSFWhK3e64AMGKXCDJbcogGnVW9S25wDaCLZVEJfaVPz7WQTN52s6ytyxDyV
iUOMzNZ8yNmKRY5EKsZatw4Lpi9keCVze8XxXHGIY2dmdzuxPB3bWx3trxOs/Off
aNdE7fInc2kva8ulZtjrdjggIVKFMAVA/IhPlA8KgV9j5pdRsDu22n1UXH9ch22o
GJPwK90rtTUVBcNm1/LJpl54BvL3VNpl7zj+LaeqlwvJLE1oFckD+9Z+gwz+jSNx
lkaKsSkPjwjwiTL9uOomdnpVSykOCb+ifVIzFPnujvJ07SSZrV92ILFueIc8ntOd
WZS5NrbDvLA2IsatgJwDlJfxUO0s60qyPqj6hAFvtpKbKSkgJzf+ju9C0kudJkPd
pVX2LIQahd6Mhg4iYxIKo7jlU9PVy3uTlFo5D9/DpBR2GmHR8cR0TxRqDthGVbDb
JmReSW5qWCcqqFMYwzItc24+u5yOcGfM7zlNDfukuX/VrhwqxqisplrR259sHm60
YYioNgVPsBUALn6Fr/sPcwfJKrijbe4YK49+DfrArpuygP/Z3PHuqPITyLcr6kDl
Z8krI6Xl8g1452AuNChygCXOjO4vtT4AvFY8HRnLbBP9KXQIqS6oiO2uogpUvcR9
DNg6KIqZW4gFK+WRDkVFO9nlZr/xHDetakGPrV8+K///TjF9i5XvohXwgQIYNMwK
7SsCK7BEaHVu2gPNwQ/Aawc94q92FfWOtiZ9Jwy8nhm4cbr65Y8SctZWytrOudEX
HKjIev7omvCFCWpeKWxakGUBV+mWikKYFvYPDeGHwonm0PMFTP03EmehQrBuy/q3
xC/qwxIvKhJMjlKnrfo6lW3mhlYP03fBxBa1SCzznm4jW3Bn/0sPDYSWYinAwWho
ToOcU9o4E/5QjlsjINFrXJoXUrQBNOeiCZBtkGxkBgOsET5bjW5QZsktR0JQodPH
I5O0g/Y6jZ70KPtUsqubrM0Ps3G8JmOX75dDVpFK0ODTUVk+XqMiCuyaAn/Nv6fU
etVie1CHo4yhkHRJLvQGtc+0FOT93gYtv/tWI554vy5I6w3heNBapjW8PgZb6jj4
UlG4TJjcIJiKLSF6XvPZyw68PEeuGMtlMJY361DV/S6Cf2oDWuoFrzGRAL0gMZAY
BcuRmHXrNKk674uBwh4Tkpokrg49yEBEU83UZ2iurl12uSqy6ovTjOU5DCLjC6QX
mAygXFPk4h3HUDFFjCrW/sCpWU0QyrqxCyLho3kYnyS2bPy/f5rhN1W/WuXTb+p4
m/TZxh2dejY4xRfF5PM19vzpQruEqXnHgxbfInSsaXPPlLNfjFqtuPJ7KvS2OW+p
4BbHMCc32xBW3Jurzj1bTPrcvXVC9PPg6im5sRZUvJh3cixLgInPb1a+hcGxi08N
N0XeojHyTIBy9BoLNw6RSBiP7KfA0GxGMGzB3Gp4QXDxwpSHtH75Cn5NJFA+GwoY
TUBhhJY8necmpuiiT6/0pth207I3r/CFlknyzi/SavaVvEQhDWtH7ibCAdMZURKa
KnY8nkdvwW4a8szsXlcccRfedV9eWpmWEJKKRfabsgekZcx60FJF9PfowIxNrKVZ
UcWqgXm37uItc70ZGOZq0oIRj/JFFkzp+7l2V2w2NBd8xL+GWecyhvE5chl77Oxs
tHcpaOfu0BM4S7HencMOz6J8DaYNMauRtsI9C0Eh8xPW6eBC/iPaeNG8IUJmAAep
ck5Ok+wwLOZGNE5f57moNbLbn4L/gZ8DcdK4iqV5DjhD7uHRY6Zb+j33TFWfVgn1
g0gzPatyCXBr1Q6vTaVLW3yyjfajucva3xnu5uCb0FSV07X7eoITdxtZvNBOSoFg
HCDL9+xKAXzm0ow9JHWwm/x0zjuPASGe289zpRpEPGX5j0JfhgUGs0LOZzX8mKR7
YzLKKXBbi9SRku9+U+dCf4nMxEnc1/HpfBFLBlynKbaM+BuPWtjICUiTAm11jqaR
f7bum8ZFppoM9yC10iaicFpFrrZJgoUrLwldozBnx0uFaEgYJJRBpJFcWvsYsomL
XurC4vWrhDBBisJmZaAiQ6bs3+07mHrG0ZRfrTdQIwUlURqKU9VhvXXNGROErX6O
uglaaP+KYy40c2qCR7UvWOk7NtQFa3XQUs6C7Mqtbc0TPEZlUC6py5K9rxmaFrI4
rXiTNew9OtqV2zVnu18RWs7bqbO4BHcNLMnSha5NzbRqsv9W/68tQq28yXJTe6tW
MaKGQlbFZinNrR8zEqfIDsXosu7ekNfT18Brbak4u7GusJkc8UfiYcPmyT9XX9+k
NWoBgkR6Jr3/38b8oZxeuzGmMXiB7DluXf4G8q/HUnVKxLTKOF3vhR9XRt7lkenT
VJhDSZznDGydtpUUh6IXyDLhLQkT2/zvZZd9EGYNfKuNwSEFIR+NknHSOupLKXZZ
Xt4fovpfhluxsys/liLNnmOT4PDCf0KzNRLW/61JKvw0G4k3aijAWJ0q377az3Mk
mxwDWnQ5F5CK+SI6kpEyjrEcwT40jW31f0yqQbNh3D4KRkT+Q+eyUOWOk8IrVFen
GeP3xqpLtiX5cIJacUXVQgwfNRLHC/9Qgu1MnQHn6FnWVd4DG2Cjo6PV2HFgSIBk
yty8ETB9O6E7LVhqMhE0ZNiC7XoXqn/XH2dyagWmvbefM0TAUZdCbd/HSjG5BqGP
0oMrW7OgIOMHXGRQiKTLc+6HysS4YmPelHQruQMQN/HbKnwKka1QDr0z3jeUIy0u
NRVI+/Vx2Z/8J2+5dbRH/OwGt2Ywkw+0kvUf1TPKqQJMMXh+djPwI6QaFsOex7T5
g5/FDsYqnAJxNfynzHzXckKcHyW0mO8QcTFO8oOLyoyxOAxgyeZfGFZXHEDPmJjv
f9iHfqeQ6arlvssJ7GGy1hZ2U1r0Z25afqH1WBMWS+mZErg5rS7AaU7gOyID8hem
4sOlO9eneK0CqCLE4KgkyoTfRJ7jlU/S6z6RootHnfixVAloFw9paWx+TU7Oqqde
P4kOVocyylrsNnySuugdgM7lKpCzCqDBLxv5bHb7c0DqxYSwBDrQSnL5gIeo5dYX
3UqtzIbZdJFXX3kqLlJBVKZ4E5zwL95wNkqBLzUCQQxZ347x/j95jO2ZuJN2347G
MiC4Mn6RxS58LIjBJ93bKR8iPUZ9Oszq+Klr6VMIL1UrJMF08EEFilz49xZRU5JF
34aWWgzQTg+bF8zFAe0LaUUVYlXJV4Csy8VBPL82rdWJl2+nj5V27x0A4e8rET4u
kiv/A2XvH/bjXy/YdA1bKNRIc7jNWDMQyvjK9c+SEtQpS8RFTSU7q5+xVaT+HZe1
0RzRvEl5aL/X6suYDrsS0LC44iu+HM4NJ5G3Ir4qli1coOXgFHqylH0ujD70tFB/
wlBAeR8kXP82OpZqt08cPwN8SkQA+dfETf31o16mLZmE6LdeetbVe5ElxoOJ8BBV
0cckarvSDQLKv26YITw6iIOi7PhVBRSwtRxi5dmZqfnzv9Bt3bcoG1kmEW46Lh2e
WlCmlBNoJN5t+oLJrxs462zFk0ZQA2cz0PWXArfIYvG8ZK7snmxosEaOqJpamgFN
hNVp1mnte7fJtagGmj7YzOyz1gZWcSfOvBVJ1ZgVuksrti659icmaht4T8IKPTPf
zhble2PeseRizW0sor3gqpw5F3nBjt5lo1FUrXoNyc+nR17B23YP8M8LHoTlRyEe
t6nG/4/s69pDVDFkZnsM61dJYUoTCP9j95Xo7YqJ2OiqnJx9ZDJ2KDSDC8sPdUVR
uhF5143sq/vppZSCa7Ly6kJjPb5YSlF7F5jKejWGLkL4eLSnd3f98TCpQGuprIOw
J1Ix9HCyJVT/TEQVqe/3BbYsAxg+TTeYH5M/+mn9cV6sCL1UDJ2k1Ug8u3MiFfUB
ZKvZaZd9But4bNVQdty1yPEC3TuTwC88L7Ysz+NOf/ynB1WqlklKwEirOmveXv4t
wxiDZqdHGnD7CqX//nRFI2akH7i9cIgkH4RN07YDLp/JpKytM8hLEVUWS9KntAMo
yglI6uq2N3Aq9BMXc0eOXnGxegkN4vMS7qSjlEBnMmnOcYTrWaFSag8xWQSkl0Vq
wQaOyBdAf3kS8JXeVrdda4h0yTkHnXkePM4JV7YqHLx/2ShHWypUw66pu/HrHHZZ
GTLC5LUbesbUxjHRnOCCsMh1J5WOwx4vpnFtwwGBs6kP9R0nMaGyuYAA30UGzwyo
g5bpB6go9Fc2cZy6HlxpmUy7LNsEYRMasxwUXT2ulNoS3wSq3wPOsOIjhQeh9c10
633pU/5s1GazIna89uuYxVwCgGpvEmlfap0k/G1S2xWSQDA/huWTkxkUPFfzpmL2
5au5NXYLmn41PqxrXbF0siNdyUX3p2L9cir/NKOL+AvpPTQyoc4YU1c2HYLSSzsw
iLhQ2W7MXjxuQibd3didNP5x66F1+9lq7Y1E+Yzk9FtYXglc02eCuW0Nwl1526k2
IoCV6eOmvbc5P6vpfjqJkDTiJwFSLUWjVM4ASm8q9cVaZ37IYkD5NxxWbLel+8GK
KRoHlxnmJkcO4/CcfF3Pt1sfSGiBjFeFRFlYwL1DFHWOGq3vkJHCO0uW+UzcvxLa
P1UjM68ivg5gdNqgTxPwNGlHI/PRB9cibSs8ThRlvpBpDv7s6UzMaKhSZEPEsWJ2
kNii3LAb8VQ3l9v9STZ2oUV64kei+vvc4nUjd0bRi5tpSD4zb0RpTwzugq7vHXI6
Tc6pcGeq9piKtjlewR2W+JH8mPboVwSGLxFDw8YZRTrieVARB1iM9GbTCQS1O15D
BxBzM0vAXTmz1rDkLAu4BE0x/OakP80quhW6oSPBwWIVk3yjV6Ft7dRU3B6hTA5u
/PYx5qlnSEMaXv4AJRK50BmbyytOO0lWNvLDW+Qn79tgeLEFAIf4IIexy7Km36/Q
qFNk6eIXEfrNP3WxV1g01r19tA6UISwz/Exn9cdpEeRFmY4yEZEs9KipkmDlVlY9
6GGa4Sljka9S2rbap8RbGC1qM5qY91guN0mx41UlLunLZnOPvhlY6rvOlYGCHrev
L1k29b2pe95Vr4NTxvtgClNrjdNQ4ghiIrHbeI6dpNdSVdQMFAaLcA3Flipm/Pt0
xHtN7Ig5KqtMGtXDxVv/AMNBRRAl4MNe0JxZAgxiYYD1pyJox/+vS0tGCQEONUfM
Z9MO0GVW4yA99/NEr1z/F/54X/xCm7F02WisDtMCKdsBl7ByCmGznb1g4r5ZbeSX
01Ubl1PNp+pCkywzrobrunbq0zreAfoqZGLAwq6lYB+bv8WOi5C0o2jHY2vwjWNJ
chWfBtAH78Wh42fk9vc4DaLHjauTXg+XaeB7zbjIOIWswfirK7XzScmj0wz4e9/q
psn++KqDD88AIhlF/xEQ3XT3A4h3sH2IdXoCUGokfVepDde5Ll1km1crVfB41Xr9
zg1lDgStzULEyPOp6MWZjhyS8FuRDK+gfD6bmMcxfo7PpDEdAzQVER89AOvHuL+c
7OwcXYkObjwFruz2niHzRYJ4gF3i/YZ2BfBRpu67WjRFdLt3BI/lGcBDUfMH2ywb
1GwYoHb/t+HT7OlCrkUwspwYin4bsMAU3Gxb47fcob26Y4B9asWBgPKIT+Z2yUJp
/RafS9N0h6ENDhJFs/gZMcKZz9fc41UcTOaXebeTObaxn+BTxitvhKJxgg46cM5y
ak2Y6VAJkmJu1T+JhsGK7y2Nl/vT9MTZywArCyPPQF3R3Lsjbe3tK9xpmvUNDWwH
tr+Qa6pasXaVfeAM9hySF1zIMr3aS7o7ICo7qrA+nP6pPf81dxojs8OjarZxpKr1
DwUGLIxsqG6KucjFkTXg7B6KficzSrw35opM3gcgMuxZSy33LDJdQ/IS4o0Zb9+6
6M9ZOtCKvVNtIMdRoGPImrxZIqAm9ZRqVw38YFaZXPxPeYquVYsvlK1UeP6T2hEW
xCL9heOyhmzaDlCv3xHYRjndbMVPoroqyT9hZsCH4QPcmmg/y21rNlHxojkihqH3
hoNfC2CYSmPkwr/jDZOYkBKVGvdRDDkAhB2qv6AyYxFty+HdvJaI7PtkNpkkSuFJ
jrZS9zgxrxf8uIoduczogO4cHHC2B6soX236kPt2uMhveyqoojSmF6airpcRBZNO
AbYgQ9ed52OwDQHWzP4RTDyA+Tz1VsDEqwwZH5BMG5kfhVmPsJTp8rZkMZiKcfdV
EDr0dDJ8nlYA7wLU2ILhtgQyzqqlwbMTaCCMygBlpwUYzu1c0CVGmvYxmyzA9med
+QCq4xgnyWbK5CIZRnZPfM/ZPg7geRMfukuxEOeMEz76pTRLligDWH3xeS3rFAIj
cRuXbveN7eKOOTKLI+vkafQ7V6Ddpai7TRt4ikxm+7g73LRsJoOKLyhqApPpk/Vb
sdAFqvVBUQ25HZCUbjbu+Cs0a39P+a7Y+eq+B7fMVE31gCSFi7KARC63eI4cPKjW
Bb6qgCcpMaSybvgNF2PFQgwkp0/hFLzgvNFLCmQp+rZqtYgle2KBgGoo4B6rzcoG
+gfnAqtkupZB3W6+S/bQSrUDCescGEO9pvd/9H0IE9osyUqFl5J+/c7I5zM2AHBN
H10OV6m4u56Bh0yzDk/laVDauw7npLZo75GBBp/p/z7JiPjxFwuNemkYxBGHjP1U
QXL1dlHPiKxbxUiSME5P59GwU5vo3ZM/yU3XpzRC0steN5T42owdbFwK8bsY7KiC
nHfO+lH6EcF6hplyHW03MKq0X0wlbaGGTJxugEsOE+x12gMaXuWLMj+0wVFD7MkO
dhBKYWFOGz+wBqHKO/9/BOYwanV5UJ91Z/h1EfnQAGq6sN1rWDbejo3M4uwxRQo4
hId9Bc7i6c/VkDc3Tg5jXlZakTvNW1g+hiIIunEnTPno2/urg7OB3Gj+TfFgHove
fOkjyDTd2tZhmw9SuZRrfcoYgrd42Embi3CoJj9XSxdr0x7i4om7ZT/sjVqNtyze
/85bP5bNxfsQU0vyaMiWWIYMKO1e8orrBf/IxcRaBiG49snGc3nJchl0qwa+qmWY
JWOjlt45YXaFwndLZw1EWx4DVYuNMXvxTLmKvzMRMIWzOjrFYSDx2A8ZPpxTLXbO
HLkdl3d1wtr8v8EOQV19hfg8cL+Yc4vRPTO2lq4sTFESAeFIT2n66piMEFVbSWgs
XVaZSg/QKA+z6BQbj6TIMKjmriRGPrvY0KTbNgsQjtMndEBFo7j4BaDh+ot5kpbp
HBqLOH9HDrST9UQ7Ndv2TrENS7micunouw8q7miLSC31t4dptbikZjFNYM3//Yxp
UT3bIvMNhFGPKP238m8YoFLhya/8NJxPTFkZ0XK2Y62mOb0lFvmu/pHegJVQpHpD
tMNSAXI7HxyLP2kehs7mYiKnJgCK2yk/i7z9UB+aepGdIOecpyX/avHHVoMAUnhe
uaO3zW8eO3cAd0duKoRZF6jWTGiTMdWdFpjeAtF7lesJNIBKFx9NMg6dJ8KtfoOq
kY8016gVNNopSLpnwLx22VHr0DCoSxPCHCNMYdxtbg0Rp1qsyr36zH/ANu9fQtPy
PJlrmqn4iAQ8+rU5KE/uianq3l3EZfwcR3MRXEFliITCl3f6N6ahfHRCkabMeID+
rvAFqcCcDZ4iRCdQmm2cJmjJaY99JwwEq9aAOTISEv0MF4HCe7IqdornHDPQCeVx
yaR8Sxbg/rjhZSJqWlIL88TbO7DMBko1uzpPSUInnvPO97zrNnYu80l2TLgd94Jl
xz4p5TYK7XL0CQLeNoKson5EQSAWKShC8b9Pqkf/61JqPDU7nhdZ4rh7qtmPk6wU
FRvFtXms7u6auibly3Hx86AtF8YOH5XkcuLgqgLDdJ/luItbpwqQuQZrjmiZllsJ
2pZGZ3sAwQtvEL3PEZgxF1lOE96uFnpPVGjMPjGCvMwku84hpfh2pVIYZabExCrT
VS6Bx2H/bbaS/CdGJY+0pj6yOrivfLizZFZMPNpDBEv4I69OWYrQon00cD10G3fg
taNApjVYHtSZ+xWWBi/UR3hhbwfs6LFwVVBnWuDLo5LIEC2kFYX6Le7w2M3fIp8u
jTHRaqdRpnpn7whrqWPpj3ipaMXjUlZXqCc8boJZ0zdUgSoAcrYWR4jzCs+u4A4S
kurd3LGdqHf8ra4i5w4MeFWIGXyaa7/HXmGECKm3X6t5uhv9UGPtLjPLYYBcnztl
3mbB4uKaC4iW+52aCH2pnckk3eHNePIbxNuR405EJ73Shh7ikpVkJvC9Kz/JsFq3
bB0JbkKL5LwZ3cyMBls/GpDc9Id1Z7LKZXvxlbxvUGyBKlYma2h+78k+3/OOI5qG
9fo5G6NEpwY5KlHBkQDuNpPNtgT18pulplwqvhdc+cYm8ksgk4O3wK90l7pa6Oam
q1NO1f1hhaLsBFixRV4i0N1ubzbQ2zktjF8CwyV7BbJ44/oBTzAUmCfgXsekf7on
PxiHCuD37iAokNXFwewwDdF0Gcpvp8HFYLFF6PbtKEoIAUq19rKmfPHZ0CpsqGej
Cbvt0LB8vpPv5sVjhXv10Ktn+6AoaIqiYnwdqUm9Uw8eH4REZyn4zqloKBjXMAtG
PQegbYGSbkM5gEcusSoFO9Eyf6ruhMWl7WFVLDaqnM3bL/md6c8XIRejNIhbzgg4
sUbirtLX/QSUYVU1YWhHiRWwHz5pxOcVmh2dEG2oPuwAjmOx9V+eI53ABJM8JzBk
Yys7olimrnQjOzuyv4BLlZxAs20V+4OMMxUqq9LwHiLqCW1y50TyUdF0IXVgjqSm
WOuA8tRWC50EzZ6iMBNKaWWsOyCfY7y/6tzaxaRVWu6jLZ3wxjw/72u/fie02Twi
kDlTCGEQ1aMXJpYo2vC00/KjMlGcTr17M4WNdmyqmUZnlZgTs7/G003pAF6UdEQ7
OuokBPrtivaccqgGnlNs1KxZ8mFIQP5A8Y7HZ3tDOo7Bzn9/Jl94YfXw+08fwNul
9VOK9sYSpa59eHxsxDfTcQBvj3cIvuQlPlevsOSzVhq0opUtvSBwZ2XUjjcIqNuD
BVRoYkYKOvvmE6Wzp+owG4w0SJwPbVDD+/4sWal7ZGGMj56fiur1dcLL4emzKWnC
qkIgrvVLVBSmy9HYaXuL3yseE1M1KgVlKjmWtOhcTXpRQK8T872V3R26jrplzweK
Eo0FPQIt0dOAfFziJkdVt3CaaZP8vuWVAqbcHWQnMim7FAXBccVwStLKzCRTy2v8
fU5yhQpRCr+9m4MRq7HKWvsGzaizp5ILVxmJCGGQ+zzuveTkgf02ICfxMFg1iNyd
NqGZqJwekIuq4bn5dv1faK6qQ1x9DyvW3K592w5I9t2SoHlAf4Gk/+UbaQdlQcm/
N/MoRfExcKlKsPP/sKSkiPwQ5qosccBpHD5stRF+WDi9zBDWllm5Zc1ZfWsttVSY
3TzmWIsuy4YqN6Th/+o+jtd3jbWZTK6nAEi34IdFSf0wfwipXTREzrTMXFlD1zla
uFPi23/JwTehO0HCe8cJvpZ8j726TsxU9xxXI9cmP4VCD77IlxSoQB70adta3o21
YyPovnAHpZqgDfHMPtNC8t0wz1eYY/SeS/o2Q/+GkDsGL/UcxAmsNYDkYE1kEsnt
t6agbaFczeRthqG3IWUGR3JhoI6Q61EGcenL0O6A+SWgmNJHVbdaX+Il8ChdTXZL
PjCaOxkGpCrRkMN3r+hEDUHYmLQNXpvu8sz7QEjUioqJRNDIt4h9faCKurnw7lv7
LcrZMzzYEtRcxxf2HmWXMJdrSyw6SaJNmJzz1BXplLJZg+Mm5pLUQZPbbL4AMjKD
YWGT/N4gu7nBYZfwA3wfWGltXBUSwMasBydN43/a7u2pNePbbQz3JKTZ7cstFITR
v28TiGyjJXQzkZD5CLNj90WbH+WCQDn6juE7F484mp3lsB4AJ88XrXRyBKTSELp7
pNwoypjm5vaR65g8o3z26RuFMHRn8gpMmxe7KTX10SMFKBvy8j06vmqhvnS/2pTC
gq+b00DAz8ZHnooaV8H+Av5L+TNL6h3hiZqO9Ri8Rh78nM0ommTzVtpgPPspwzwr
jIqvi7ISJwdHpUV9IMD2Gj6aMrWEFqbLpOoseocaMjPf9Ntz5EoNioD0BaapW72r
3UGNXWLnm9ORbof1zQmsH4QzZ3/JDL+LYzHgcdMMQXGanqhBbI7QlQn1Smtzfoa0
8OzoZD+Oex4605xxbKpnUL4fCLhhAQzp6uavqrFZgWSEhTVUB0JfPIN0vAjWh0oY
+TzkRAG5Z3MMM9Pd/11Lq5iaNug76QskrTf+gcAhNOzzAMAi9TO933MDMcCpoyos
gfqVrSGQdjtR9SZ/OTdzWa+xbe6cg60JCI1OX4INeKeY9WhlrGqWiEKIeYEOdWaa
+76dGZYObe0jTaBYSdb3jSsTCt84NdrUlqfZ430Dg8amJLqiDheTlPhsb/tL9+eP
3oCHsaj4qzrU80f/JHQxIPge26LtoUzDU6kyaO+1tgNH2UxN7/lESMZvt0Tbghr+
ry4vKRN39OSsel5ZYTbTY26s3JhuBT0vQIoizBsrxEtnnJinBikRacR7fpyOKwJK
EY6QD8S422WDLvSwvt0k6p5bmcEAzEEkb+hnbDK+nPTKg6fztg/zVjgsAxCA9Ppb
bhSmYDZhYg7U1oLdxxcvO+iJbLSfpK5PWZS8MDzZZ/EwaAdEjPJ+X5fZNRFQ6uKk
PYkkFb6ltBPvjA+xuT49RnNstnurNIMIDsRucXomx/VM5X6FHvQiFL6cUGso/IjH
RoBH0oYzc1gbE0IACyLZ9/vyKk5SN17jwu3Vi9Mc1WAm7f0CFoUDkMAvg42j9YCU
SMHJwfJUTPuJPXj2E+NadnF2bGDOlBxI1NhFfZ0/cQNF0yOmVHSaGLWNDdIkE3A/
iTC/U1icINxTB6Wo2CvwtYVgqkgapTLkbchlOqMcOvStwaf19Zx7q2/D5G/nXxH+
N5Y2SPN5JhgSEN6IJslufUWGXu/FzKnIq+KyjqG2u1ph069vZqjSyNkyX/cku5wQ
fE53uE/TBCmMfubyA8/ioJkXCO6x9psy5bC9ThbDbMAExeCyqlwaA1AjFOr9JtR3
aoYjrHhbeRqi3kmEkbCWnrrJOUKToHXq1V0DRF5pCdhHC8ZduXOTQlwg8RruWzcP
YOfuzpha+uKkKtbTjngj8UIWH0IlW+0UZHVpZji2U3c6dYD7P5MNJzYKXA9yf4WV
2tMWVBcFl1M7SU+8u7USHvqmGyC/pkN7byBZ6OCvrMJwi2QO00gItBkmQdMsNqco
nC8XrfngChZY1Lhm7gtcwEaR5aaMwWTyzPd76yJjgKzEbMLmT2HLn7vDf1tRFDCj
zudXkJ9KxzzcbCYtX2SwO93d0PBfjGmPGJbfuxRs9XGRViseM+AY8nFW/sQRZsPI
/DyTnifdy3zrTFN5Zx8o0XeM2jC/NPQR/qUQFDnUVC5WUb4x8nTf36YY+8Gftpbp
pTJ2PJ3waqRQdpYVz321puVLln0idgynS6gnxdQHtxb8iHPyDGwY5AkyEMWbUSYh
S2RrxCrcOAe1B+HNm5sqU8mWcCbL8WhPBvSyuZOERi9MD06HHYzwG4OF7kgylEwk
ganFc8WBDtBkAiAJbU6ZNEoq6UbqgKOpVLpaorxhi4C6P7lsJxOrMCO2M97ZvV6y
etSVqNyiKw2fsyaEDTu/S1FKlk75Co8JltXkMj0B4KAk6FUqQvjzq1RFvrmKXyGu
XVgEi0GF1QonKW8wOp9SwUWK5iC3A7HwQGpCHgctDBY323qsrSB1wlhzqkek3AM5
aE7PFkL7HyOJUhTeaRS7/w34W0T4CeqKni2DxxraBrhAHin7ay1e+vv96NF+D/sw
GvxlBWQ8pnKXWR89QovF3U+/VJ14MObYpBNOw+VSVL0zBaKC89OKVINKjPEMfGgR
eOg8IP2kSBBnm2LrSG0HXSDsc/g6cWQ1qj35cZ8Km7eGEJ7czU+OuTW5497YMUu6
ZYDkjJNBohj1H2hskIUnxwr+zrCe3SU7AOP52kUzj+B1ZkPfDw+IKLbLqiqdiUu6
QJJW2/ZNmWBDFw7skNGkDGsa9lY3k/jwk1Uk6E1lJk2LK6CGCxjYSH21/BhUeqhZ
P+INqrK2siczlV8sMzOLxfiTWkfAEq3Sl4PBr9VNSBzWuPEUhHj/wYLoEya2pHtC
l9Y5DiAYt7oU1zSIOKqolj6wfTxgy8EANFA8beqTl8xuOsnfE8TgaQ0k/Sj6j0Dz
3KbyAnrBTFNREC1u6FL7MhhVoLOGYAvHvw8QfxP+uOF1FkSifCAq+Em7j+DYvYHp
m3P47ZqssyvjUgTqOW9MtvfKGuWMGorVILsmsXgqxfkQkTWRZx5wH68HGrf1GP5y
KUUeoImn9ydoTRkCEO+qVyr2MKPo9InYc20gAavcwOgkg0stk+XO4fc3AwuXBOUp
9jLXvZt7ebj6GYMic97kT/VJB9BGxTkkifC/E3nw5ChEbdeWIIDf5DDgTrp6JpQt
YTmgXKAEm6DgPReIuUQghUN6T0knZpPRFJLDnFQQBqivFx7DkDn2004MPgWoqOJn
JAuVtx+jxlZyv0kX8u8efWoq23iKlffgG9sJkaeiqZWcC3T9cImZPKqVOt2+LcAt
FosjdeC6X7s5D3OttyiQBW9KK3XFC0eF5q7oxDW+W1az7uq7IvQrv3ClEmrc9pFa
OD3ao4CkXM94CxvpO2BiTtgtXkXiCHWN/tqCkxyb+vvc284UMNcIW6f3Rv2+iBCR
lzUga30Fl7rJedocRHresWgz1insr86MdxUB0Fuf5/A/F5Gh7GLloYYrrX5j5Zyo
o9QIpeRqedjf2KBVHp3W+mQbYU5kVVPrAbC3Hmad+/knYwZVmi7YmI6NSUZgkXXr
Wcv9gBOizv7CtG6XzHJkgdX8sfu4KNtZW9wTG9p4SmJVlrq4wxi5cIsEmc8nR5Fn
4ISR+/cIdTQpUGmjfCAcxt8p8fH40D4i4BK167sqWzRleUL2dq68q/q61YLyEtxK
ErlQi3VoSiYJ4CN2tstpk7csprQF0KclhdBM4FE02zQo3fYyY6gZ/1XcKF8cgkZF
MNiEIpcPPAdY50vKXPYfHlH6S3GmuQOjyzdGiqc6UZM2DTZw4W+J1EIcbOuK6lAu
7bmuBAeLdvnVO5t92pbW1uE7Zqccp1Z7TFXtInrltQqDjsOgX8Z85t3baT6QMwOL
rdatGd1XVKQ+iUaMiSmxDJwFkKVpdShyG8MQ1QzI7BzTvrJDgQx2J7PL+mLyXzq+
EyjKYDhQumGi2aKWzwgI/aX8C7w8DT+qjv8qlcfQpS/9N4qh5UsxtLWcBMQP0rkC
GY2M/gNmW1CkGQQqAv1zXdRcT+iVGwKWR/vt+ZmeFNY6evk0ur5Q5iu/n0cIOxVr
xMZtGRba4tlRy9hGLIK9cI0bQ3YAKSAE0aeLK5YWBWH/AbleovquiXH+yTyj/Sm3
ff1Rp1TVk1S4wRiiH99DPid6TgJjXH6JmzAIeyn2fowdEucFJcognUGP/AjkoVMm
Fut5v2pPMvj9dgVPs+fr6QFK/2Ulu4IJ0S6aR+m5ALvWmyEf0XeKbrTFV9nmBGdk
sA0uvwyNu07eakKVroSsCW1dFgRYsIzszzKkFi6wBzAhocbpDaQaOsoZO4RhD8is
4iiNTn+cCoAthuPyvX0aDK9Dg3upFX6icda783cIRNJ92sEv0dBzBFoPjNGJlsK+
nvz4EKAzD4JF5zXnAAbiNIZckp7wsHQ0RaoK/jRJaADTD1B0Q28bX4zfwQBFck8K
TVEty26X7uSXpqqa7xswvB4zqx0N4kqKpgEhZVDJkC37vAvLP/bE+3riw3SW0nr3
lo4A/eXNiH1/DrTq7BgpoOrBEvV1xPbtxHf9oPLbMcPzeM5DChAE23H5GxggQxEp
z7pu29hTNQYdvlIfPJkWyakgA1ne7jDd70sVwZ3wbSEnZ+/UE27Uk2cs4FNHx29E
Nf7VQQthZeYSY+PKtaTKw/gl0CgER1e9SnDCqorzCr2s2C2SR8jsWkPfyLe9EvwP
hL1aXu7PcZau1qABMn/q0n0ge/B917GlwnAXaSRdj14Ar6JRfbb6j50A6FRUPIiI
CPKNwocS3d8j5kCbQEswwcb5V6GLYKAVcEYkpmwrkiMwR9POCAra8TX4oDb0de3k
PonKBCgFGeTkT+vNI4wd2rE7wflrpV47G7Xj9918pUkRfcQc0OT0EuYAxOjpQUwa
lBXItgeii3OMZYRNUf8R8RU+0toN2XN/WioL6aroWpZluMRkkM1DW8Uz/aBAf08l
mg1vFbD+VNbrjEfKEpTZfeUWVfoqqSv90rQNIP+wHuQu+kIBq+W22Nz2casEWiw6
5rJQIaemqsmOC68rbXeOenFaxDnpqWwoV1+iXSQMbYw1//vHFGhOl6qgbFX8U7F/
9oE64kNprmDe975tEBe7Gu+jrH7+32yvGkiLc9JiCLXzzK7bIeU1Pns//GrG71cx
1x6t/I7rEH8gW0GUUYQtrq3PCGdvnOQ9iLh5aI/oVQzr1WzBOdkOMysKow5d/KNp
aViHaQBSgpTzazFZx3oE0SvnoH2ORrx+icRTxNId8Fn7Nlznis9EvL+v/z0VCbxQ
OCI0tzlaM8HKMm7inOeNo8vEkGsaQasPZzC+9WPLDr50SbWR4NuT9YlARus+eJwl
kbAfvHZt3eamDn+VkYqObPfzqsl+4oadgU3JI8Fdf66JQl6AOujHPP97FJScrvIJ
r1y7Edzfnryx19S1jSMDABEwgCpPGdswMFAQ2Xh5AsprEjm6x3sjD2O4yC6VZ0RS
vfIYN1gdQwf0vUuls+pIuRoAmrkUv7f71EljwiryTFFYA4ejwVxzSq9F2bUJaueg
9BvRZu+Dl/uLWNk9L3bLGhvEY34MAIXnZEfTR3WUtyGnCbg4PazH4c3Z3iM73t4z
wZboh2MFyLPQ/m1roP+naTQWZHj5XMW35/ghx/JPFZ0Rz8UgtO04aiRaOzxoNVwU
/0EClyVGtOHwo1goS0oW4vkGZLuO29HG4tW88j/WkPU7hvv2BpSr8+odqDQDHug3
ohI9uKR6bPh1TyLvMqJ+XdQhM+KkGQuwDOWFu2WNwZY9F2sEoZahM48wFaCIAJlP
HFxZZiKrHDyMY6VngB1cczAFQ7C3BSjBjkGOhWfu+Y3c356naGte770kzRul/XON
X5SZBxeyEIr1ZGchyLAz4ufPtaSDQqi2N7PjhrcIOBGjchPvjUukFio9kE/2nCCL
oKIO+iGxVOYg7Zk2w+Lz40V+o4rEgWoPn5+3nOXQnOY90NuvcpltjhtBY+mHLFXv
/h4HFbop4R9pzH7CrzzbkbQ/uPbasOVB7scbrRBg4rVNbZBOZ/mTmcF8XmV5zXGZ
2cTDyrVOIRb2ewI44SczKPojaDX6b+FVKbn32lVFF/ywouhQd8W2GEGsLNcMHXGj
VP7f1k9op8hm/kqOnxLFlDyzAKLK9UaeQhllNgojpD4LpIOVMZo5NIpztn80DI0T
6JGwjuVB0tvvdEWkR6bHPeQjQ9Ih3gZmY8SGurpGBqojutLhN3o0fMPPEtaovPos
GtXftrhn1kZYRc42xMnj0xzXGjg9dJlF+H5D8YF6X2T2fFu7GzjPLIqPHL1mW9z2
ShwK1XnsQd9+SilwaajJ2btaJQeLPnRtKYd5ria2nSsNjRX3SnKA2VnBc9oyDitp
UGlYMQnZp3vF2W++IrI31rUF8/C2hiKe5qyyIhYLs63ZObIR1kZ2Eon95UCkvaA7
ez7pCIxFiFkjx16LQ0bA5xL+pKecxgn9AVwXx+OTxSRL7dtG51LG8LZTPeYdmEX6
LGRBu/QwYC6zVduBg13dx5+6cjWULVOQ4NcEs/MSpZzgcSG0IE9+Z1QMA27IZ83Q
WZGkR0PzfVS8O0owOC4otGCo8hp4HbwqtZiAaT4GxH4rK7jTkt/sxAYi0srjLyV6
FIq9XEFSVYg/CuyBAYcPnx2A4ZUI4xvogKDvQ/OmEpoWQfDad88uNXBPt/FD0Rro
ZmvJ+aDPnFVRjmSExoloUzSyguirK4k8Thq9uNsfqxQhdmLwdjRokqx2TE1slTgO
xgPJR4yhogx+M5K421HHDiAhVD4YT8d5svCxv6Bom4EeyUW9yGuc9SeoHrTi5M6G
gHIKXJ0y+oC4943j/3sh4Fc3afp4Ot2YpEZwBCDTFKJs1r81nmXAojg2arcvCGtN
H9yEEKiz86GPIE5sJNLCdxzB8IwCRADHjjL4NIygSldNIJq1bf/V1XL6NUQ3rv2d
ZCc8mQtrsw/TSLIfvO2E5OYFGWhxdFsKiYPfc0rLFLUckfVjRVcZXYHXRg/4SiAC
Z9JB0qZQgRmSQNYZh8omPAslJC31VI/gMD41HL17AxQ8EQGIKm5T/FXuoXF8afEf
YL2jy3uHn0emkXiPAxXF/VlY8ZmDrJxel75g0/a6oa86h8SnKEu+OL/DD3G1q5c2
QOML7cfplNIUmWrXRu8R2as1Dvmb4X/dgZQ+7eZdsiMJ75q7+KNeUlIgYwRVJXRW
iz+2sz/uSO05GBm4oSL+/hW5OHKM0vVomAfzxLFL9LoTZN6cdiVYsZWqub5xmn1p
kObaLJ29s5JXi0hnUroZft25KXXYEoTVy5q9bPxXXsWgi/9QfBWsSdhI5Pj+tFf8
10cAH7lD25CbxpgR9m3yl6+k4sD+eicUt48KSl2CsmZvA0SHiowOniURr3+6N3rz
IiG7fA8FQYrFG4e66gUwLp9DdkKEIX8kG9yEefHFE5XM7XelWfdHN7zA9z78LoOf
ZVC/tLRZf8FpMO/TczH8Ic8AhUYqeyrZFSD7cbCQUShtZXoSIBHlYluK+5qnkjf2
4e5edqT3yCoVJ1V99rc78cTjraiiISiYcOGeCGYLPRuIYp/pZGvM4Jky3URgEcJj
RA8ANcrTaFVxX/6DSyB86w7RMZ09+BP6ZnK22vITJSkYe3PIP1zYqzoPtDIZOdLl
w97orkADu1dZNvCnTbW2jfaNX1o7s0CWQgCXa8hT3gB3oReuBAvLzXccFiS+kuWE
OW/lI2Q+9mDIfbJ3fKeWSij6ONlNbQ9g9tCxxtEHiHdOYnmkPOk0ATAtrqVIQOmn
RrzrQRRagWUENB7+8alOBcCXkjglxaHYILXCWnW7hJEEUyTiOmGu9B0ow9+ATip3
Ii2VQF6dE1DzUezu6g7aM3BIrPje/xD3qr1ztJBVlP4MCJRHEA1Fm4mzEeO3Jpyu
mbtf1NsSalRORLnBpYO5tJ692P39abZboMQgciizftxix7FxGyrcUFwC6oYlmb0I
Vr69qYkTCfD0NRqCipaWSRKyvOGdJMOIg+PwRcew5aktCihjO8fNcUSi1AbskSKc
xcTs3DZ6vAdiYYkhDLvdVB3U8QkLgPP5yXB7K5U6rdoR0pHytUaYOCdUxAEti8Zq
2jq2msnIV1HbuxbnzzYH7J8ZxcF0s0k4SNc93IlCuy4v9T33sGEPzivW72c2wLx/
CJ+xnZx/m/YJsYNmN8b5Ldw/tR3SnRnRFKsdEQ/hr2PhdqfLOShRa8f3l1/Op/ZM
xiOyHAAwqXQkbzbtxJBCd/zwGQt9qpA7uFXRtV0QailHu6ulc2vFVZ17vIuVkz3x
12U4eR0Am7GCwJXQT9lxOcxFKAIKjezP3jMWPb3S/zcymoW1kVehzbdGToxC5hqk
6xy5fXvaCLcpVphD6biiUEldKY+XrgZzbJ3sy5CvpbTdfHBBCcf66Gq9BhEDQPzc
2FiJOQ5efMTlC4kfVfNEqbBwqvMYliaSNfRCgE2T2eSQ7q/tFhnB0GtN318y631J
zjoZY2JN6sKA0C+BPfWjSXGPDPDI1uEG5BdOCBUrjYwqWrIwwOo8KzyLibj5iHU4
yKFmgxXo6QWBvropAUj6koO9IoHI7Qmb+xhuXCcJyeYpCPg0gWnqvhsLibGdgEvQ
70EMPyZQTVzarC36a8i6pnFo7JlpJlxBIwOOIshBI65Kq3lL906EX52vR8lgAkru
ZRv91ljEbykKngewj+lGqPeLIQ04hfcH2BhYthH4k+57bclzwWGTQ0P1XUn+Ge3F
bfxRhurmQ3nvC9J+s2378LlCcMU/zThE0Lp36rgndQ6RjrC8HFwXBIVyd2pQwKt0
/lmbQ/kHhXuT1giHz0iPQnDON+PbFluyNmhVQBsloD1qNm6pE7SP8ivyGRyPjEk9
YzmmbMVh0vyCa3tojnbMEaZpK8n32vQQ2Zx2FM1zU3emIhkT1oP1ZFky9XMKlMcG
IGR35OY3m9zRLI04DkUl8BwC3/qJ5w8lWDK5Q5X7gDlw6KRn9IW2jkyaieWHNScp
ZbIljjY1+FBpedjrB22oHWR6H4podQSFzIqCsFMSnQl4gM0fxiEGLoV77T7HhNKa
UIo093LTUxPusCoMUNSzsWdKMfjSNOFNMtU7wsDQzXMHAvttApXkrovNPRxiCtQt
R5zrK+jhNIK/nsqMZkhdhinMOqXSYaG6Ms3tE9H/DbqW9eHbhdJUtp/I1IB7qXaO
exiIef6gM/Z6MEyayDZSYV/PbLZCnxHThBkzbwq7gPlPJSMhmTfnNe2yPLq3ZqAW
kXreuIvGIfXip65jC0OIUXuSwLeHr+etOlws027l0c+FVukpetRLVnhiHmZuIKId
GhaHWGyNJbC5uyhjx3xf/IxCXfFn5hFVCLtneftUBscSztyYL90X2a848FzVtROb
bzmfrom8X4UDx5cUxE3CW3gVPGyAkbYW3phWd7CZ0P/wLhuqaYkmtz4v5CkAij9q
D2KBFUuqooFTpexYnPjchu4hLsqUaxykJPvsaiduDChkZn1/dYAHApl8MDtvfktH
KaUAKOxamtq6+UCrVK7aq0TGx67ht4KuGAuqAQlejSVGTsjTtOVCr8mI7MVMp2zV
918KdVa9qmLWqGwAXRumJWBFxGhn0yPgig8KHNzZeozJ4r29F2ygBJA5ZxNvakyl
pXbOnMzGKby9dG0g0B3NO3v3KSomXqM+oooRv6FIOvRuqDIBp3qyZwpxhX2UmH8U
23S1i24/3CbNHAUORlSUPvI3w/sZFByOWQWtpSLTc7ljydk4/6zSCsJpf0PMZV9G
c+sMDzd2YgSvOOl08rpt6Zvauve1bgprQPK9MX0YdsTdsJW4TuQNGxjlVNqzYWm/
4Omm9IWrM8HxySbSOHFwZzFomZrCXzGDCx+noxpe93pCoPvbHbtfUkrMpsPf6O2p
v4dokZ+ZePOsdFt8ghCai9/q1vOQKIfD3u5a84Dgg1REEbaKjWmZ/OQWhS8+rxA0
qzHi59UC7BQ0ReSE8AEFKNGnRIUuvTrTxKkSnjIUmiR8x8vhHBY+8lw0VRxSDfvI
I5pyfP0O5iZCKPKEED1od3JMo7FUQNUz7ki+gUTHWakTUHycPT8hOAWqCAuy85FF
vD68/2iXMRemIKOE/kebW0iFJXb62k8W5Ezn5nl2Ld4peqaTJ8+rMes+5IXZY7aU
froY5SqCPxjRdBfKIkCJhcqxs2K9LW4qiykXHRfgt3zMGxYe1TFHvmpTdGuzQxx5
/dW8uASRXM4mR/yGKb/0RHJpTvr/SZVUII5p/K9r39XsqlOf7jyM/SIMl78TtZWV
2tsU920/ynfBj7Rp3jPonz+0lKpvfcHNBZpbO3QwoBrGW3+czprTPPxXu/ZeJRrN
tXhOUj/vizovTECoDzY+RpxBQbLFz/ipQBmJU6slD17cC6AoSL0ttkdhVks9SHPN
r5Nt+UhhNIYWVHngwf07HP+Op/hp8KvpsFNihDWKtD3JF6vbGtXPB74JWVVvFqes
ll4bTyFbS0isSE3RyYv/7r85l0p2azVluCQd/mJlLIalHvYf7tzKIv8S6AOJndCA
MWv5ecll+Fj9SKtrL8Zh3rQhmPUhLqSLcb1Z/1PwlW8cvMD72vhn8E+aXK/PbBNF
zq1GeyItya4jrnKhjRyTm3DYl7GFI2chAVuEDPUWmgJB25NH7G3UdCJiEeneP6ew
ZQbr6MMKTWh7gHYU7NU9KRebshb1SLDhrKin6Xz+H/ZpP/uMFKUWPmLxmmkGtpjH
gSJ5dl4EDIOObQc/+OCGIemol/ZkPDmqV3jpjESU3hjW8hHTC9OxyxKTisXGBw15
uDNdVd1QN4rYOQxyzY7n/3A5/zVkhFWpDWMCaoflx8SfGSUMvHrGfu7dKXNwcF1O
0BHYrKq/Ac3yDxapsm9J6hfar8BNju9jJSXcxvqV6hPBa2zstYn0xN3iUqC8Mm2l
HmJs/wVsQKgxO97j4d/ync8kwyOIlPxkFJAVEbMZ4UQmR2N4parExO/7Tucxhq3Z
ovySZdGJ5TufL0IewQ5vsG93dG7FqTf5NsiPg5MS86BOUa2JQ2SGXWJ2QctK1wog
jEZImy8EXxjA+iiRq2ICADmDW/UKNhHBX9b0fjJLWmEqKrHAIXEskd4g+dqr7/TG
eHJJ7+3Bik67PXaciloV7SwltLhHyh1qWcOmyK/2AObcbRc0/s0Wh8yiRXMYz9zB
aQu+u6Ts3rHXYJrF/KoSAD3rq8iLYWcNaSaTo929PKn9PvTBH7Nd9Tbrj/HtLHBG
WiLqiqEi17XicmGKocLsAJqMT+CAxljn4yj+wLev6HHbkPuKzKemnGKMdiIzQZfq
t5J2bYH6CCpZ/lrzTCeopRkAERyVsJu3cUd6rTDk8Bo1PnqrLniafomiFvZTmj6F
ZBl6mk4AeHyOa9vdCUziCxj6dF8RWbHHNAzStJk3DYxiTTZ3RzUEnRV2Fo1FQxqG
qkf5XzGJMJ5GjLWeaGRr/ZX92S2QSksnKRO1fAOhL57Lf273uxAA2QKWH4q867QR
UZCNp33G1Y+isJ/Z3oyZ1UzkwdYVnoomsDsYn1oXD5IkDn8sLQbtizBul9J8crNl
pTu3yZM3NOmz6ueDvPNst+Ao0vaUD2uVTVanj7PthAMgTPhSSq5fM4CAZ3WQpUTD
l9HtyHUscxJsZYgbzYD5o3p1sTq1OGXiMKSl2zcjZJ3IZZxxYGeeTUXJKtsAF+6S
KN1VrsJngIhqfGipp7dkMgOB2qYq9FYGoJKDdzHlT+x6e5FxPLrK0bdpAcpcm1D9
qemxm9dN+lCha5rYcP4R4TfEaTsxVepTZLebMpSvnPP7OWA48hYy6Q2XhywZU6pt
EqzJSCvbPbl6Cw9WzgbsourZ6WGFCWO33x3LtyAF1BLxQ7Hv6h3L+aC9vKg4xarA
GXkddKE4XNIQu6J4CEio/PHuq8F3uBk3iL40plQOxZeyppvuQX2Pg7cR1dLb0FPb
2ruqDdUJvP+4YpALLJ3xepxfb9fwoV2NOJfWKMoIiLjDj514KV7fQrDJG1IQ2IH3
+/0DvoHYQLTDrbaU8TYd3pCLqWNEUkN8uCiwT+aPuuvWTuHbaDJLP34VgB4mhtyF
36WFSkS1Rre20CemDrN1lL21MRPY2ZutTrkCR+S5xuJMsadBgFoQlql9RAxOuIi0
kbJDOPkEoKrY8V6CF4qyelAR6oPM3dJHJrm8KuFu1eOzLeiVadNkvF9WXaPdV5FQ
UrCywyCPXSgUPGEM9rx2BHjBJirDo6kto3OYc4l3ewKLCt7sVtJqi0HCUtMj+HXU
rZAKIdV307nrc0Sdw/fONSXnVmK+mSvHh0BNqLsBN2SIOez1SF5jA+dzuiYJIZYb
67K4K3VXzS3MJtlx7NPgeIHnGITDfolBCuiBpXaGLkIEaBm0OKN9GPjwAa4GgPAa
MxYZEJBLbABnC+zreK5uRvoRA2DycK398p70DWAa/Z7peRsOvUQC6N//agnmxG89
YLtyELUDAuvY3+3xdw+25rSoPzfnH8JTc8+eOxaWMgYrpdlB2Py3an+da7DPlLlM
PS4hd25JrRe5ksyDBst9OHOIKE9vREtIFSQExg8mv7fb7IHf4PbVq90K81gUzJIl
fXzoVTSrhXu/5Z8Seilqr5kObSVuXUmRrE2Zv1xO8BjB/BsEd8zuVo9eKBi9Wa37
NQOuLB9flFq7O0PwOsnhliK1QSSkuByNkgv1F4hLkVISaIVbhTfhO6+2LEikxkwO
eQXqnuVxd9vrHwW/8MpAQCobqm5WtBUKJ11e1YjjO7EKVOm8B2+WCta1IyUduVgh
EY0aNZKnKvQAU5LNXvwW8yUGZ1L8S34xIM/4l45xsQexY/nsqE6ZIb5mviGzq1Cb
OnC1fBkHC9pW0W0fBsOPSSvFLlthfp7SRiroG6auMk6+vGE1ATFBZH1YFllQ2XSs
eZlF2KWe1YhKLwVykn0MUK25gLVuzwDvhOwGdERi3lhYxK33hQxXVcQVRwqfD6+C
BoMIvl7NuxO5vkHb/4dckaIheblA+xmHsaVYv+vFsIlw9Qatf1tHUtyUEr9dkhuf
PQlPKca9yzGxXa4IEbwnckEOWlLSsFdRUpWWP0Qd97jiubHy/R5dip8GnLDddQ0/
ROHaX1zFerf5Ld9/m2IL6pvvEyn4ORBaHFJJtKdKA4u8JVdCx80rzb+LAu5kKoW5
+kVP7h/mlLRiI+7rPaKWCjB2bua3VjOkheqHXiIP5WctEXke0obH6ew/UpEwvJ8b
1sE0lK4EibGSrN8V4CKAp+F4eEGcfC1mAptAUqU5cw+CjOmvVLZtDayTZs6hntog
eDoo5sJjjompf4ubGMe/SYdqwKzRtO7/jlRFkTVgogZ1ABPb01LNUz4b33Qmodg7
/ZTW0aB4F0wKEFWZGfDonAKsc7sm9f0PPXcFfUSkv8fMGx7RbkANHkRtQYf4Keh+
SEaNk96CYzaNfXm+DUMT+TZc517nLIIlQpXd0ha0HPdoLnkxweq933r1fwKJynBL
GvJra9Vln/p5kfLTmA0Uk2jYD9WEhfkdE9vcMcPC1ZKv8CjzW5Y/3ZMifcQ+Pdyv
UG1qSuQS4j0nXYm7KGMOe8zAX6eTjBvD9wc8bydUYegNzOx+RiElYSyVDV0TFxt9
DoAqRoro4UcCMT24RFk029Vc8iAN01CzneMHCkulBd3eS6X6s+35/douzsxEtwH9
vm4t9YLWbdE7Nxdyybew63QdfgchyPUbQQFrDMcdzs0BGhwo2d8qZJh99V7ngusc
/J8DW53xE+xXrOKJ5gyln+ebf5opm1u1x7ZunDBqo5gSojYrCzLao+AtZJhGCObK
pP7mhmRVJ7cobeACJsCMEJbDqDfh5r2cPuber6LAUqb8wT2cb2HHOX0UqZSa1D+Z
XW5vbXavStlHxdPVY5zP3C7RqK2Snc+5xHXvzmupYqBe+exWCrWWaySOFxWyqrPz
snjju2uB+9YCBDQGWNHbGgwc+Y25/P5ASIvE4xC7XKiA6F9YbZIPs8nWQtjU/Op8
aq8mXyeXd7c0tM35ene6/w7CzlH1cfutSzCPGNE5n4uGKuAalbocn32lXP01LQwL
W63WvhosRaMq6LSv/+gQPK2ImmegfFPGHWuT7DoG9Y/z/5Q+NzDHSDj9xl4lHrs4
1rQWEL3DU+m+ckfuTzDsiGbN3EMicveeV8CDgRf/ouvufIfvFKY/0yXWF+ZAiP2Y
/WANEBgoWnP+V2qLUysGGJPiw3Arbg2xZNw639G27BMfBc35i7irMmZiDWXSij9S
GV16NrjL9Upbk6CoepGRsUCrGXbbI3UTLWaVq8GUO1Eg6m7idXSLpl8op/5KQZJ2
MNF1xaYBmQ/hhB/VKomlQlTdPNm9eehn8F/YZd3ewkBIrcxmDi6qsX0V5JuzADzf
oAtiCHvwfw/i3YBVOmT2JkPckRbS4XthIPf1kTKH/ILTn8HSCzyA6iai/xG7u32n
r8TNGJIhbZkQH+7ZgOXRvkCntOcV5v3YAN2kYToQgJckkxH1zrUyKU0ZKMyzKsD1
aSaP7+NE9XEAGi+KvRVaIg3W6hpq+MUZKGHbs9dmsqCAzDBkacmwdTvHu9g/p5HW
+Zt290U6fyxnYmeJZmtuPsd7ch7GwCrCP2wgKprjlX8ThBe9McsbSlBNsBVA1OHV
2e64He7UBEhKYleB8V5XyAHPWwvAIlzQp6R69PwxNIuIQmWDAPlWiurI2iZ1g015
VO8pBfGrLKQ+qMlgIG5ZYAkikhyIHnOfatycre50j/yAV3V9gxRCHj6IRmzk3pRb
+Piq5JDYOIGU6CZLKaOLOHyf2gmnS3X7evp1gikl9ksnd/y9rLlIu1AxsXKb4xOv
/dYbcVDTz4U1JGYf9M0Q1RrirjJZs3e8d07ykPKCnbDbe079R7DthjVB5llGRm4U
yI48DPuIqDQNHyaWgqwcQvVGWBauzNbEQgaPu5MvKtFVVg6/cdU8P9p6q6HIHxKd
60D+TplJj8+mh8TC0KCi98AyUUorBWonxAv75DfT6K5lEAs8BxgYidPNf5/il0cV
zEHyDiHRCQ/gdWD0ZvevWyD8+qMlYPH1tWMlhPTkYyhlBFVR5YIjbod0/BDTrtxK
Ck3ier9/WtTsBQHSwaOL/fa3byeZwvWgrKyHt9ir+SC4ymLJv5E0+DLwGJ/nES+2
tZpP5/m8jwQmLKZb+EZvJ001TCOHWT61pb/BNj44v0n1ZuaXi5MIiGDQBf/9n2DO
J28ESZbU7R4mx7oc19Iv61biBq+adA0jHtwQkY13GxIUdGeaFQ/2MoX/j6L+YGPf
RRmPxNvv7W925syOzbnHAIgIC4MRN+4gnRop/NKqkOUfnK6k/g0UE86OqIMj8NmU
+zltGGmfS4XMRHRTQcbiBB/advnoCYYaDY7L4AVbMKeNaRreWDP8uRrXuNyheZ4c
2T1qimaNMR1cV1VlKwegxrMejQ8jAS+8JruYnhHI/VUJbBeOeNF7y489E4RHEczP
3CVz9qmUPgIdaBKwo39Y7EzKjZNJKpi9alYfihTTfnorMXCOA8JZh/e0I7KxZ9Wg
j1DUBTvH59ynVDNVwdfWm/597t1U/8y+fdFJkVxHfhKj91dCSGY1+xmuOtcrdaTZ
E5xYD1GoyrslIwiPNg/9QQYEGt4NLY51ep9Vc/dfAnQYPxjfaEGaB2Ia2d4fz2PJ
2GouEnDMmsLkjw0GHc56gUlL+TsZ3WPLV3cm1knBdG9xacjF5OV0NUj6/l0qpsFO
FL19z5aEXuIz+rSK8A6Gdx67DyCsdyyul0osH6sIN4kgueOTLSpgRn6VL1aH9tov
fmXrzb72+sbHIiCtjME6lroif5qsxrABkWMvKM24JRjBMOMrokWRiph8A66H/wZA
ILri7eDHSN0m2tYstq+oHqAJMjdMlBS79+oH/TgeJLExaufM9JA1Gtm+XxlcRKJO
dTKMySHpYajsTKGk/JvjeeCPc1K4/ER/afzImS8y6JZrIyQmUlKkMwLOeAArOhvK
qrdt1GSQgqj1ABg9lVvsVL/fADTb1EllvL/KmdBJnffl0i0p4ySnAiN/24Ztfkzf
jJ+YgMnCdpNlUkFdA5YgoRsDwh10L9skdUpxs6g2iZF/O/avaePNbWze3SMFfQfZ
narLtd7vn4LyPjdRQ0+jEr5C09E+WioZsokHz+qLD8ErQ4r+xFtLYXj45KuF2ObU
A5f6ZBB3e69Zq3sXt5fD0Uf+SNrFYNx1A/NiKcOeV04ZPUw0cvobA9nDG1WQ6jpn
cAdjuTDAU70j52ClWosICKqjeLPzQarZPdf0JH5oUgVJQseOQAfuPUrSWmQsKrdl
zDOcwkvbNXcu01j4xiVQvErH90uLEL7fy2AC4ILvcGWFwxcEpusNbVEKm+pFBVfA
Qtjy1TkXtutOP8/PbBBsosACgn0365pGzu/Lu/gRFF/t1RaS60hZ7VcSvFFfkqfL
l8lrXX8cTicd2XrhRocaN2qLLI6PQ7K419STllOhHqla0WcYMG5rfdIoEUuipVgf
nLXDGF2rBcKvOEfqAg8stUR1lxjMWA+KXFBrEsaxwgWam3CTklfjX25NkkuBwElU
dJBeAifLdlwt1W8uwxJBssRhCsG+M9ds0QnF/UyTisw3nUAKwT9DoxpxLvAIzi3A
eEQdWk0N+ezYqopo5lwjcsVXS7fNNVAAX6hijz44nLGeNY9f5KE7n8zqBcKzG++J
PIeY5QJFa1CMFL/FXi7LXwc5OZN9sygCGbnODvHHzMs39V2SHw4IkZamKuMgpdEN
oaq2Ysxo2JwWHsaOLi4nIUaEhjK5Dsd/9sRYJNuRxUL/WJXpkMC2WbYY8scRD8CL
NCZNkcRnryVZk+fj6354bY8pxU4uPcvxZmrP7YyTQHcy6aPS1u46MjyeSLEkcoko
3WGMzXnpYxVxhLyVUCpcGtUOKmH+NNPPi5U4uOKHIM0EHaiipW/RHC1KNmlvbUov
hpS1LAmxaghD9EBlNGyfOmjap9FmkmmObEl7ESF3ye5fuxTOiPUM7Ipn9O4o8UaB
qalD195Oq+D7Il8RKOHFiheko/uAKx3Hp2HEEn1z8vJo2dzpfTlPFlXMqSCGDBBu
9B7fYclq6I+Rb9ZVcC2q5s+Og7QHz9wTRIH7AyqHx1TWPUUzknV/Yg3anCh99g32
M5eEJf5qLk7yLGF+DPF0z7Noi0EYpTjbVLSXWVxYlMcUF8USVxYhS+DMRGLkgAyz
ESd+dtabyzAhn2jYDw0ZDNuAuOshUBPtYpYBppNaI6m35Jouq6cHdgiRwhwTi+O3
K8lSnx/+3NIIqBf50nqDHl69ckeWWN6IbtoCW2Ms+b2SE7cgjE48SoVQpfXKgWg3
KQUPBJUufxRSXLL71P44aF6ndjxEQFukZqUuJ6wvOgyPaj4muRQG5nqd2OY8EROM
onUGWdYgR+TkH5NP1FX8bTiE/U6BHY41c8133VzBkHwjH7tREEBb/HF4/8o4XrVd
9w+BCUz39JrDgF7Y7hG7TNBmtJYwBsMIAeD7RuFYLq1NpYqiTWvHnJZgadfB78Fl
2xIdEjAQaI5IGEpEZklxOJwSpDG17sUTfcyWLwu6D6oT6Km/WGPD/QcQO3mcCmrg
UFMe54np0E4T6Aij8dwvX842ka62B53KXHGnUZMbgZYGy/F7mVSRI+EJq6AUefcE
PATGQCRv2AT8GNBKy4gPLp1TB2aTE3khW8oZhF3DeZ0ldpwuokB+NNPB8mjSl/9H
ZX5iaAWvw7dr03a+uslOOZTUQ9OwD6O91Af9E1+fI3Z3Pslr6CgQfkbirgEi2cZo
E8crNvB53BTRac6Gj+m5lFrMS0bNHoJ8frlrvDg0GbxKQqO1MkeH29dSPPmsuXyR
Jt1IDHVeElLR9ImPJ1AjTjS3q4pwvlMH9aTOQNFFWtsNIlVQJ9JMJT80GkH5AXQ1
tjDc51mGgBX6D9izMXFNzmi3br0oDc4OccRQwU4yOLO6VLnB573EXctoc3eHrid8
9mwCqDHJz4njz9ktilCUQelCJNZ/NBxDUKcbwbtXLFvu3rDIBtSMrQu1pbGVzYn2
ZQsi0ATu9DWD4phnsJBG7XtIarGXfFnurgeL0LwsVo2eNjMb9wfrBrBXs/bdfAXv
0jnACCtUAA1MChjeamo8y5qZlXH680M4qror5nWI7U9ePsDTnmLqWEM6uM9xODWM
4VN5IGpH/7tMi90cZAHzsKjgQCGTXqv9WjJOMuhQLjsbeD5Ka/TKLVeLPE0P9HIH
npjf8Az07BWnnN5oMD72eVj1PKzbN9fleO5aUQWnHTK8xoTIKydU0YEdMdjYlH/W
Vgjac1gdlqdSbLCiGZHhCunexyRaKrxO+nO7mEh78WPoKtwb4AS8+6MsBT0okw6n
Clh29uksrLEdrEkxYR5I7MUNn5+pMFOLJlyNZeyYW/VuMGso/KCgB8j+sWoq1A5q
K4KjN1BCyMVcYZsU81W48baRLGaBlyj8+XJ2OQPlkxppifkGttz8tlGmkX6GMry+
nfL3n4dSsXro7WMxIw2uaFtYU3Rdr/bWD0BJZ56oqs0IsIHiQ/ntJ410k4WAgKO3
zzvBQQBPlE01hNYF0e0+f/qwZ3KvcDoT3XMRtuOa1cKO1eAdqgiE7HncP0En1OMA
x5hLp0vkFlQUFS9NIYDqM1IFWLbV9rPKmzOsna4M+QXr1blCCsC6GXKOJG7TEHv4
yzAuhWhhULydiC+jJfJUDLO67l3ar/EZfsajuKVCcJQWfptUkzeTh0WRT+ucE+W/
T6nb+rJKwm83o69hYqkLIyBJ9kcTPOvUgFbnLF/Pd2Ryu50CBL6ZTyDjgn00OfQq
Ku4ZDhqdIWXRXl3DeSfv1lVnV7nLuUc/8I8+93LkbMfu//jsDuTJgD/+3UEDAv/S
stx0Jx/NXvL71GDbUQcH/DSTQNBXcjKll1bFtEAH2h56VmRZ3k9BtR8su4a2JxZe
9Qk+hdT7W1AvbLXMvpk/brnyHL87DB0y7KCn0TcOgdh0xTP5GxFPn6DgAjqV1L12
NTs0VgqOGtl5wvVxJY9IU2TE6ilSQ1N/fGXs4szPlrFnUHAvUSX/Q6A53UWH1tnQ
ounYWar504awo9cxuIhlyPC7ZvJ4VNGMfAKJxspvaJTsOG0oTYAvrNKsmLfCp8/G
Pb4t6RgZ3bZeIRVy8SHj1XvyCU3b7n+NrsQmXCLaEqo28h+FBAbfXzQ5WOkL/g5Z
LbYBOAjyRT1anshmM1mh/sm2tI1+Bwc1iTVuxjQGB591WA0W+NrrWTzXcH4I7rhD
2beTAA4zcH9rHELxA3uMjtPi5SjwyF3PLJtnzT688bYqmifVEPTLjScJF85gQ8cw
yKf0y/qCJlrJ2sz7gbEkDVeAO377befiqsyI1NialJf6aPtEtM3DaZ0VVvr1Rs01
6vUlRxI+jqMa8XuW3CS9x152LB4ge0CRLrnbAZpyfunXJtlbQ5r6hIOgeoCoabVi
4MqDFrjpk6iHNjMSQdjsZFFxvrPolhMyM6IKraDZZPL1UDsAMZVs5XiclvAa70N0
HTsvq51TgEHy7Hn5hE3tAvfbTAIc85RdwbVMbx3c44MPuWE1XYaz1i2l+iSuNoKB
nKrXoom4VGsqxKSYsBTc0bOGYvyXzdATV/sa5GONskfeM5ZdjinE5SLO1tBX5zjx
gCf9JlllHsY9khzmGjbNUmY0a+MbP7XRt380qOpp7DmhpI7w4JPEvhnsX6WGimC6
L3DeEP71CrXf3fzHOqzm7M4AmfG1u04E1o+V3Sd/1GAhodf12YCKRY9qvgvY5/OB
NOOl9D7s4qnw1o0utNONnIYZ44YayOfXP3b9pEUe9eL+mcr3vlGN97XL4V2FXSid
yltdqoAXbwVCPo5PzA0V6GT6RUwxldsKjGtLz7YHvnFihdX6oQS+vY9/wPpc6bHE
kJHAE0ncdC4edr9+e7uq3mQPjT2t7LGMBeO7PYRsQmUQQZuTLRnrC5TQCdpRfvcH
aQ45HrAN9/PSTF4lzV2LGUHVa5Fu2GXksjuyZ50X+4UWKsc9QBh/KeTG5du7rVoW
u8JE6JuvK6yQuhxcc1pNKi3SfNUhSZNyrs2PZ3fUg4DiHzq/6ZaMDZPGozLVlPTM
xfpi/QwFnKR3uBAqTiwBnSx+z8kjvyFWSXjTbuOsFLDUsOt6z22O/AUlNlkqzf6h
SRYKmgc73vNwyiYCOJdbbM4lPLdl7zI3AxM7fIQJNaJpTBfchqvOk9vjxBZbRCSD
H1KCybi9CTlO1PvyO6EBEQe1mKthjAo6j5g+/R76uJY/A4+eLmevwYW745Cox/ek
Mz1Cr8zTWAsRHJi2QjuK9MZAQfjc7a/KVp1U6wmfIwyedSyg+fMqCGOSYRFI3sW7
4f16jMVR72Wzbc8gY/5qrYjOgo2IK8pvEpl/ojaskn/7+4a3c+6t7N7V2v83WVJk
0+A7kRjWhpQscH0ROLIcWmXWG1gzX8vY28yOxt5VO0vk3SrGX40ADFZ/xPopwSwJ
seuFXpuoo/EDR/kGLZnYxnZ9bQ7DTH60AHRe/QuBoimRRUc+wSdcpnbulh1dvJH/
cpY5DLPJOAxoZzPzf3D8D8sGsJCDiO2oUsefC7aZxcGrgt1mYItsnyws1yGpeBny
W/8wmHVRA/qbjQ4Y8ibEuhvCswfRo+oDmUKnp3XFtKUfhBLk926U5kq0/thVv41d
EZloGpS7TgXCeViVktI31KQybRRFnbyQo7t5+3YJNqCRgjTtAlkUa8M08vk0Nud/
eCt4bghPTEljUMeiD/49brpQijrPGDo7sYpoM8yUUzNcY9IX0rgygUb4c6S980Jn
hudatcpl4r+T3QGiQWISz5A9Okgce7ODsuJ6ctq+Gr1dsXZJHpeb0yEXSyybkWjl
xVUobKRlfDnKMz1SyTUCvoI3YGK5DF4rFe//Tn5Es8IQzH+eobdh0Y/J68iKE9Mi
jRIYYGo5ELiR0dkoibT0DgAXC0hRSpr8wS+yrTm7R2uRHd3p/pGwmx48vYcCpXbD
w2ySxPfVu8CiIj4FZ5ViwtGuTmSJV3afRqGsE0bz5bFGWi934x/fdUdux7yBBmKI
uI5WtX9mQNWtzD3RF06m93j7zJyBmf0nX6qSKxqjCStKh2Q5X3GuVAG+kti0BgxM
mk3OXpIigOIiFdH1+gqqHnY2kUA3gF5CMLAQehVaGmQdAMK0AbxRN0DuBa2F8G67
IdQ/bCJXt+ICSsMcDVxc/a57b14fQ6zgPPRWdcqBU1NZScSwVxFb0h1zc4ke6vCc
SWDQWOoSXaR+agtAec7xMNqK3ne6OQ72eJISnPQO1zfucRe4xTmpgnr/cWoVkUHg
cy37W1UNrCu8GZlRL5RVOTrcy8kr6EJXrCXIOabNLCoR/z3xJNybk2JGW8xiJfO/
mxcSs6XrfSiQIEoLAnmbv7Q6z9aDFD7alLNvRQ7DuFbKoidd5l1OSUcYdgc5YgVZ
RS+vuuU0gFdRjRzzsa9bXL5dKjs1TYR7eMnv/00u3GpHp5LKGKxS+P2v1OLSjXwG
NA5i7PMSZ8gk83n6178xQ4WdA9qW8Fpipb+SU4pSP5zXyqp4IXFXmxsA6fYk+/7/
tBOG4QC7zNZqu4hN35ciuQkW+S+iBiTliLst1EVZHE8iAShprx9o3LUB17Np0+9K
l3baDbXS1JPcqWJo1WAE843dS9cBVIKsmD2IU5Jl/g0+b+jNtg9jaVvkp0TcRiJw
Ubgt/qnPmOSbTEvTAGRuNKZ6wc0rSfY5lzoR4NiKpNfY6TuzjN5X1eLDRZ0CoHHj
91f4aR8nMcanY0Cqlcn61YU+RBMdNOyMErJtOedddpYOriQd9ue7Wv12oBVcxaNF
F/pa584ZfLV6lRp75QY12h7LKGl3LB09scB7hzRdsplpD1s3vD+5aoILFs+YKOiq
B1HDDldc4Ik2CYhV0A+tEAzBAmBGN8xqD4xIkNLonzOgxSprE8sTRI9jNBi5POA5
vpFCr2paQSl78JLBRF3pTHUgHo+qIEzBuD0TEdYZlkom0CKmcsUT7yed1DS5x3XN
UO7TuC3O461saEzf3FKbM6+eqNFBkWrVSWQ30mOMuoUohtgr1BBTTL9mZ0+Tzjng
NoeqcOn4DbZfNHrlLcsw/j/LU9LCM40sxxTgC03c8DEcVOcUzLm5UTzMUgAhaabK
ZIIjVt4vPKCtlsY/H2BSFrxMFPEK1BCKoAA0nYTnNhX39wvQ7hK102MwnGDIxT6S
mFvUtd+OQEyBqUgseWQV1Xnvmdh5l6uoZTT+7/OklAZR3/1nIWbXnAsrxGg9HtNN
oZzwUxKxz4oHosyEHqpJ1s+oiAYMRT95tSdbNWB142xzz0vN3FvhsX9mylA1dNq6
/h269BtoL+wh2ohNugXX0dLO5qX8OVmvvH4UhsXVp1LZ/8XDQz18Vj+MGQ7sJwQb
gSMH9WMpSVggxg5cVPAW0vpWtN2kmMWdOimZqZ/0J7aiwC/93pjAwiNJMuhN5PG6
Jnug65rkzkeHwp1NOXh76l2pzxS1xW6BkfKdmyoCrO82xxT2IOcuG1+xp6VHRsVZ
mfMNS5Fxn1kslHkiV9nKWX+vV30GMFLVtSvX5Xkhp/2EOY1coNzh1ddBvBqpt5SU
QgrytcSuM9FGhCjeOx8BeF+1xTV495fZk8DtJWFcLd+mKz3nqa8erOnTSCQ2bgNN
LUyCSywxOikLp/d6DTObBvpibj3lI/8Dg1MorOODD1PfePQwJelWw7WPI3bLciIu
dAfs3YG7HrAHM6EIK50L157Fvyn4S8QLRUvkxyUcBfD2w1XmltcqisTMXW67Z4Wq
BHRj6uOc8nm2oOfG1o3jGd4gex2G+9GWobtTMxwEQ3avRsDiXDVdYUJwRXffrTo6
uJuP3bUEF6eI90+ENIGqBdHKhtzcJU9KVkE28mAQsEaLl3K7CjA4bDCHzQFsIrOx
HMO3+v54Mcc8Oi6rPEXS2NhVlh3cuXlVqncpbxcOYb6kXU5igdB0EdKO/GDq0P84
doqDOVxX9QW2VocTudynWCn2Wb55pSx06I1O6UOVonmKu5s5U4PlRPkuNII3LIgY
aDpqH4H98YbD9seWDTbtn+vWowxJRUrH2JSowpaGrpr27/vW9yOrWUrm2xqI1uT8
9MCc/H/FfQd0Iz8sHWMDbcWcRKvbk6uIT7QW+xzWX+fEQye9lD4Ne7aH4EzeIu8E
MzqEJSJaAuUpfiFsU+HoRszNSJrJGyrCnD1yEfkrCWDr63dk75GBvEvt28ujbEAI
PEXuXj2KzHMc0Rr4/XIkxRLF6eeBeYuNN582Q0WTanlWaW5yjiQp5fW54NJUsSUn
26sgwqBdcMxOWe8Z/HmM9Uo7oyutFfkHYkN41VUTnECxFAdhZHLZ0+IPBmS+nQn0
DYDHa1C4QnqzwRKaeqfz+2HhnAuxMwOny40zfrX0a4ViQFhu06eVIBpGUQC8czuo
Z/sd7qWWFq9tRNjovCOYxCfjDZPJysVqxQuBSBmfL6mlNm9/FDwbuIeBe1D4m3Lq
95XxLTkRfAgDZkEMxZjHh4tlmEKUL2YKPQApeiybpjMfyIHqa/DjN231yzjZiLGL
OROI7+EObdMYmj3flFNN2uHGnHvIDQ5bY6jL+To0jQfIpOoKS8LlbKCxlDR4PnsT
AHSx+N1v1gHUgbSjpGwmEY2skT+dJx19+YQB3ghpk9UpTozgs2JsXuw/AkyxS7G4
J2/vtnomGD45Ch25PIhbOs4nu4e+1uHJwYE/0avWlIrD6/EVVZIMxfAq7HWhY789
MjemwVpIiJjrA7Tvf2RM/Hv3feSTukPCi7TMZTkh2jwnTaKTXY9HcpeAUm9BwCre
M44oMcF1JtEcUsTppzvEc3/RU8YQZJ5BZbfdYehQ8sm3wWWqLrh+FLuJKLFaYGzB
Nu8j/vXnc6voHMgSf/ERtaXUet7wPWcH1YmTQKBvGa4ZS3NdP55fKGy6DAl9thID
DisJkBK/GSZIi1jvhYNBH9QLItYy8hgHEZCK2+437Njt9IyKgmuV6yGYtruRghl8
og6r9od8ymQau4LSOCr7lguUQZEBjS+bWfbygHQ6L54ImbbNeZ65mlR+w/fFhqUl
jq3SQJ82qGsDnCz3CYKgAaySMmAwXJWNeH8XNUS+oKKKDCiMTzO8tzi/7swhVhFJ
CZR7+rOLZPPoevLI+rXUQ12DOP8YQ8moys72CuIewMEydtidjz++MDRQs8fBD3/2
LGnRvXmf7oBe+QZk7UArM2oC487M2nK119NgcucN/9zPTFzQORjp3LI5sh77kff+
aFH+qe4jTT5np5lli/QWcOKmEeGHfOb5RZqu8xkLvRlDPas0pk71jI2iqdbRLmG2
vKeRk7VBe/bs5eU7AB+tJUapzTKvNvQX1+r68/CX1OZSbvtvo+1Kh56wypWJYTGi
4J6vQNOmgWr3ZlFYZnVixGldmc7H3UiRqOwTzj2fs5Ynviq7y1zWMN5CeRhW5SyP
QDUzx/D24CKtTTM9zrutfdM8HlZgubcKHt/xkEFn/XrO83tNrsN6gBzOZG54UGFC
DrsS0coGxVAIxGoT/XvCGIScGfSb2V2YQQ5yykgM3dU7bCGcXfWlDXbEE3wHABSu
bAudSXzYjrRXKYhuZumshR/Yh0w2UuRuwzHj5vZB3BdPt6Fx/ln1amjM8a1mpHoS
CRv1PwciK1XWIVga9tPc0RcGuyrWh8oM/0kduAz1RuTI2Boubf7P9lD+TL/uhNcW
WSep+zpd1353sQPYu28TotlA4TBds7ulitvC4Wsx4sQI6tjFu1QrnRoz86m6ObJw
YR5Nanq6XMIucCLRqlWi1G2q2Ys7kAZYeOVWOA/Guz2Q75QLzLUWZMmoVya418r8
+Ap1FF8S1IDogifk1catK7sqB9a+3RTS62f0BJd4XPlLd1jQjukC7EsuSNtjVswZ
iezq95H3xj4XVsmtrQHh94Xdvww6m6Sc358bEJmdbf+OekfELnqRrNa/DVrO5R/K
/GFg2o1PBspxmBBDd2j/1D/H5ku2ACUEW/deHol9UxbZ1YFpPIhnNHzUyAJ9Ul33
SowXjXiVFp1fTvxr7Vhu6gSYwLZWwyd6CcenN3XkcQwEAtPxUxqAdKVFDIz6jqH+
+mKvZAWcqjUWmF7QGPFCtJ9tqBGeJVI1Fn/B63B769kh4O1+WwRTJmmEZxf50UEG
SboReuZWWnFNPd2R4hFQu/v/kaAtiLTgfue0oBK1WVsmBB6MVE5UN5oFjP+KT7JH
LMsM3gPTsAjThtyKveFRmvpR68CyBaD3oro/glk+W5mB4swySNj9zvJwAIRag5kc
Z2qw4UycdvD8U/FyaSS8kE3QibaeTLdHWef+jCTQGHJ41dpNpPobhMwHVdtiI9cr
T3oRPnuKNbLfSaUVSzAD8X5bwoJynISLG4Y04yJNzECK3FcknAPNXkZNY7TPTLNn
2CC1qyOoo1J3mQBLb/SW63TnzHwaNEK2OdRJC9Rh45C6daxQYnck0DhhyaWNEMwp
dATI9RMDrF7rCk+9AKpe6bVRDMO3VOxCYR2ipT1PLOMuECv6IGnTp/VBzqF+seHP
dSZFbZSsg/QBU2KDma7ihIi9SVTRwPW6JJXxqS6ElW1yKrkg+HgyIkn5cjOgbfEs
Qi3q3R1lAF4AYCQp8UT8hI19ac8zBZ9xXew083JUsz0JFE8FbRQo/M7lMj5Fh9rv
IYJS1tCjTrm6a9YXnQr/JJr99xr0IGS/l/UBR1y9VKTQ0Z/i5njEbnbFKSgvvP66
jCAaBTppEAfOMAxIHRlxXLfHN61hv885wo3avEg6dmJcHPT5U45smegrs6SD+JgZ
dKyZCYG1IkF/jgUyrqw+fL2mttJJyszdis0FGDJp64YD2+F4y59ZvXLlEryzAPgS
StDG5/h8qb7mAAlCYLp51WTI/A4uhvXRCkADjo7PrmBRAhSysAHceqVJ5XVYTSIg
OtDTSMyeJBSrfOGqLiWf65eoJi/l+81J+GjmwhbnT1BG6d+ONb4diP+VIOKi5f9O
s7gn2x0YY0mMju8SynId3IWnUhnKQZ4xBFQFTNucuLO55EDDUCMtAlnsqIJWuLt2
vvvjATvBrStrfiZxGvPZn9zHc5LX0oEZnAhmnJa8HkaR4AbA6pRvEsJxeqgVUQZ3
Rmxp8ACVgjB+zMhc42GaGZYeDhPipHG5V9QmSXl8/K/BOxb+p68AxBZq/YE12vOn
saIpm/UKyV08H04WfFULQcQvimoVNmSKv1Vo46oNfMtzhQU6avdYmqJJaw9E2msn
C6wC7DU3XkNCdYXeH3X1/W60Ua8soMgPPOXqEs495ScpiFimgdr/PvQ1xHB/NbX+
T3iXP+XRbyyGchRv9y38TLSc95VWfEB8NCyzm7JHVLhVeXq8oZpkku7bBOxXVK4e
9+kFFLf5F1cPb85IAzCBTxhMDqVo8kuQm53KVGelyeE021y+cStzNdqcKscZRCWF
UfAS25d7347PThOPzxxqJH1GuDe4j8SkolscC8Vl6UMRcPpcoeWAyax3UsdItdY+
OkZjrK499NrJNfbTzcSr7EKBHxLGl5li6sdADj75r0aKNARH2Fi2Kw3gKL+blcBj
zrZ2oiOXNBWkDZaDS92Q+SpP4TabmIwVlG0Hda5j63dOnaXMZLfEGoV4fQ+Dkn7W
sTmhbtQxNsH8OEMAJ94l1c1ni/+mkfgmZPHH49G/+x5BFmGmAkgDGO/2D+C6BVlq
l7CgeQQ3qNZjkNdLLYiFSX2rU+FqDaGodtidgl1VzOU4sv0y4lxwcHZvbjUoAFy5
GfZ9kmyuxB6xpe8PeltBOm0hswILHoGnIKTPzYjTiAhBCtSGfmq/lqRBB6BAtWUd
+boHDsjwKcM8YujA1t6yx0d9cNNQwEdxOlMtLjIytkClnV2cEQjf7LSncuu8WoEP
do8aW97aTCbUMJP1wPbYZN4SS7NE2y2rCFMvrRubyNQZIoyEthS7EGCY7vKR3lLa
xWm9f8n1cGzpccLHt4ZMTbaG/yoErt5BxIwD+2EjyIP60FY7dEOTXU8dZbeAfIiN
u7fl/SY2aim1FEdpWrGi8nt1T9mAONIcqapjNo8sDmKezoqKJNkFZA1inhiJ2pnD
tKicNDIoLJN7kf9O8tCQLuYEo2qVhNewDDw57zWyAh3ik8hYryc0ZF/mShaHvh4J
5zY0u11EHI+M/a2tQ8H9nR4Xs6HSbHXtC/dYMHTTT6veIMZ+338iVQthrG8Dl++J
RWj/2JSwg560kGBXsk4bjsAKbAJMfKUyh8l+9mCOFHwcJy35hsvY2lsX095Q0/yQ
HrlceC/z7kNW5A0ruRYX/U/Gp7AtX+Wy2vtfnH03UxFq47vdaIg3AyRqFpxgwTMS
f7Ea6t1z7h3aBB51dXPRzZqJeZ2yoLOoS3bAoPtywVTLKWWQ21FJsAgixTynvuzn
MvRW2tQRq8/W2VqNS0H27tI9gaXIg4P7SUCQCaLn9oI4+LpeNoHo4h1t+/XlhjB+
YgKJDmtWSEl3ImSaTC76b30K0NagvNbOqENZu+Hv9XorY7H22IhMUnLNGYmKj2ZT
hG5BBu/AviNTaQVUhQ3Z3F3I8o1ho/vgjykAVEOKMI++769XD+f+vudWTYTbWvrT
NkrcmqNwWmNSB5OhCswZAZKayiYY3K84bsBKo3V8ckEJ9J1AJ1ytb9l/eEl6B8zD
y0ar9CwY3vHcC+c82ajKdqKsfg+SN3LsTbwVSneCh4a03bAn40Aatlyq3YQB6b9a
lv+MBCyfn2dzETkCfbnsxX7Drl9msgbPIBotmWEZUwDX9qMbYsb/d0QqQtp/9dvy
yLlNYYPd/OvUIeuS/1eIdjbOhTA39mSFqB68o9W4IjERwOTZvzhVxA0yOXs5qEnr
fh0hguj7280EH3WcUdy1H3NXks+VNPbb7GPUsLeeGR0HoqTjDYlzLcJI/GJCaxVG
WJAx4d7qMEM4EB4bxlM6kSXhAi7J7Ev0Gk2hMqQUm1jwAOtNwz++j/zqkZKJhcGB
eW6s+nTBZWo0HUD5aIDWmNu8F/NXfQs7MPA5nsL6eaC1m3qmObYsrqjwli6i2RNh
LgiqMululXf2CHbbhXTBRsCC0ubIuvpO/vYK+jYB4E5E+rMqNh61LA2jr42SXlHi
5cNFpge5vEV8JrOYkyeFcuGAnn25194rJIIclk4m+gc+aLAMiPnBcKsXY2YihrOY
S6LomqgnTzKIr7vG34QfxOL/vdfXX7u1PkPnzxyAGL/2Ul5dj7Cvz8bbe0qJIMIz
L3U6ODNWHgXu3ap4vBrkQreGJK/GD9eo3k8EOZ9PJMKWrky46LXkfiiogvs7fHi2
5JkbyRHjxb8ua43yxPWGeKHbSWAS5nMm7PnLFELVZB2bsNygSQ8wzZa0B30cajv7
DOcP5xus4j+/w+ohWB9Nz1aHSjICf4E1DM+kpKiWJ7qt4vTW9f0vZyfLHcE09edm
Mq9MCDIG2cYZ2iiSd3Kv0GaUNVn7h3z9W90rtJZBYUgs4jUY97nFcMn4H8/n24+g
Q2bWh+X9N3uKZZuFrQAYTExA1w3ue0hZbG2J9uWYyIa8HxXDcW22/0b+zgD3hUbh
MYUB0iS6+kcYWoaB+zCx7Iaz8T86DsxaqVErryo/TTD3JmgPE4QO4rc8lTJoTGEz
i3GoPtcwQxGxOoejPCrktKG40tAoEVrBAOlFSZ/0VM20Q4z7Uw1nGrX/wPm8/0rj
6EM2Nai+tWNF2xWSdJa2SrkE0MNchay6ZDm14FWk7AWSSbwLXLqAN081knmIdrc8
wKihZFLbMlnNi7uYjKbNE04eRZvqFGNkN3NUrTlpES5YabGupvgzeoZQ6c7y0btx
4573lHq1mtCyuXNNDULbkghZkKlSNvYffpE+ZDBmZDE54+H3SwCO3/CifXxjb+F6
8RDHO+a/5HXyemxgScHTrdcoq97fFW0WC4M9PfvOpuS7uv24xULxFGKUv8Lh/UNE
0973bshaJViuglD/Dp3gEcGItfSiw+j71tyq+R0tnJLA4vamOtjrZtyFBYNV0lM9
5I0fCKWTx3IMRzl9W2n46r6SOfGYHzqtwHsmv9k4AFvtAOGFSp9Iy+tPxp6zJQyL
wuGQ2mgWjPsrfFVqWjFkorhuNFDmmCrJkjc06nSrnaB0R1f1yJr07PwlEN7Mff2I
PcnzL35W5wVWHpGQ2qAN+MLc8oZPyrxAeYXK+Q2jf7YzJAFxywormQ3SFtgXZk7l
StJcKlqc3obQczEdG5SZw576EG/6HQ103u8APnkzEArRqeYUgy+8M7ysqpOEXueV
upkz9iuwt1pbdZk12t0ss6xsLlwoOxK9+CtHJ9wFWMDEz+ydgX4BK6M9bcJrkbDg
NiM3FaW10mMou9m+5AFU8pt9I5rbtniGYMNBwA2HE5xvgHaqHwmu5GomHwQsKMO3
kEZOseQ71UQo7Z7VI/qg2IJgC0H9km2K/Pa0MW+aAS+hl07Sx86T7OPyarD15nLh
TK+BHr5l9gUToJOB2azHIIO69XgcGuKSIddhv8h0y5efzUXbqlVhvYxGfqQvosiz
thjwOk3DOjtT4m9vpZm1h3TIXLLrxi3jkNEhPjqtFVAHirErjDhq/K7GcHm1JTHn
vMaRVSSHYP+T37GWHDdD4Rj9/13ZHRNmJ7uMhqjxkHRSZRTEx8WndHYQNlyc4inS
WbQMlKLhuYUAwI/U+KFUwarQqovHLkPETq6qFiJpGXtCoWXxXKnBnMiAt2lK5638
7DY34b1VDA6DScxRb595aazPrPRPIDe6euRbBpdkbCa3PXU2i3kO0HamQD37B1X3
mjxr9UmEfk5NQQNuFQBXg3dYaoIwsOk+gt+Hru1KtPqTMhbwePZlK8bAlkFH/lLl
2oBsV31hKt5U/39EvrRTcUBkoGSXwNKMwr0goMOM5XJBgWB+rfMH55DkwfcYNGYu
lyhDQt00E5o55Uip7mwwzb4K99ppOxC/mVK0RMXuf25oYOFla3y05wt63M3aIEwm
nD3hZCurrHBa4i5uLOYtJkV1bui7RrvDkh5h+qLbbu8LVBJ6bKA9ACWXR0lnZ5G4
A0nXqjcXCB5hZOISLUXv1VnV9AiyrvSzwUJ6PSvSeYAjV4MBbv6J68PDtulkv9YI
cU2f4g6PHI1ibCHO0X4Xr3qm33d+XwiCSdNUYD87qx8W/K/Vez8E+BtOdQzh3NB9
E6ZK/5uDRVbjFDcAZIJOYLwx8vGOC4yq7IcEBYCPuTtzmXE7C3wQFLdHSfkBIQ81
XhFjwSVBGJOyGc5oZy4S6FLrxRDQh5wORfPYvcFIKmgoq8VQTq9gLe1JxFlWKBop
BVmjUUUN87AxTn6CfrnGinJO30Ivat4DsUOUVI3ltdCaaehoxG1tV0NY031JuFO5
iCRHQT3hGvZrPADBEew1SB/uuC/3+JDCBm5Edz2Y8OMXKrbmkSUeMzhAUNvj5AHx
w88+Yg2jCoCX9dU9L7eg3dntemZrsptSz741SZd1purytda+XPjU0/IFnfWfNETS
lHuAioCEbySDvvrR7kvIJF0/KwQ5zNrID8iKXBQo+cNmcj4Th3eMTxL89CCiS9rw
xMoXPVe7oK/OR5c4qRBVpgIEyAvg0ZTyLodZQTw88Esy6fpLpGGRnphvsCRlruUR
uK9bn7DdXH0TWetpZwSKDC//7tJvdKTD9dlk28qrdRBzPttiD6vukEtmHPsXxQEt
NAaSx1X+7/MBaWfzp/NtHkcpREblmi1DsgIoM34kVeo+JMmJkqLJ/g/we6V0mV7u
XPZxYoLQIoUOMHkxigGBf/eMfIeBNiuC8ilhV2aCXU2gMVhCO1rNAwq+a2M1JJoP
RcQaSvVkDatq2jM1u7xkvEDZes+rq+Y60mf29kWiemiN9cRjE64G05bRUq/4pXET
fpAG5ZSbYKu2GpNegeB+iBoSU4fMkK/fh+uW0jQ+jidXZR9t5l/bfLj00D/E2wR5
efFaCIaeGGW4lgekeXlBSXHAd2k01V5ZdYg3DqAvIim2bXSyYUl2M871m6K3VDNy
izTWS5WMmRRQOUWK82qER4Mp5fvUniMkHRoQ5ErMnrSjMVgjyMAjc2CMB2uUIfMb
TyiF1ci92J2S5JymyuCs3WKP83HenVgetWlReE7vM7wcOX6/MmQGP4XZs8onzOkQ
BKrEperrwh0YsE4nZFJUNQyT+0Muz8nPEOR6LIl3PtnZUQZNX89EXjViOvIi/60s
eCJSFU2m/GbldWxrhIwJ7HJf4ywfmH7enNotGfVseXlqtpPWTH95TV0rZ9GarvsV
ndkz3nG2dBYMvnQznJRruXWWz8JoILTTsB1xDuIThqaoNOmu7sFX9RnJIgIuCaiW
V/n8UAT9RBVAkHMUNNt1cV+eQHKovNVTecpHCaEzXyzWVTS1JmT+0zT6jUCmyNOb
gZkkTMGYW6sl/NJ3CBICOGMLy9zbc9pEVKhSj5P7QxOgyMOdosT52pjMqy16rvbf
4if2YbKNkTpIQ1A+TyIg5jDIKhegfqGljKJKUMw/ninpEnden8WU36KQ/201YWea
sMUPBy1y2ioYOfnOtCWD0IaaY26kwO8ScoxUpMRcJVY63EYK0UGFHGFGjd6gEJZf
G3K+Deg5fm39IigTlmS7OCZSoibsLBhvNEZ1v6pXNPI0D4bWqo6aVHpjmRdpTURr
B4soQyl4E/2Ynwq1p93YvU1R7Ct3iS4KcE+vCWfm0u+t9uZAen66eqo3vwMlUWDh
lhnyCCd+cPvFSXVENicfevfLCic7n3RjWK5W2Cok0XYC6KtB4HuIf0Bpf6XH/Hjn
3DqIdjrR/dJidnQFeEyN+OY4upW2VCsTyoa8ALZmxfdD2SxTH1kt7S1up4+tBp9N
oe3JNDsCvUcfqD0Vbx5P2HIJ4zk1LNR5WricXH9Oz9DeTjsrfEd94RxCzykjM2Ty
zC78e3NKIvRuWdeOkbqmT7Z4DHTcdbKRlOw3nDUmI7bmeTr4kJTKsreMy+Hy/oPu
/yf6zMApcB0lv0a7HTs2O3hO4rZ0iI1CMo2gWfyjlhE7YeZ9iIgMAUsLKp+gP15C
qkujpWazFzL2wXYrxJ/pIn6uXUtY1QA6boiqQOq7WMjGV8NV3RmNi7UhStt9jwb2
xfas2FqXMhhTUcZ6NleJIDzx85W870+9JWbUFegIhntdxKrodbj9uRbPt9RGN1qO
Rr7dBDCyTmHlrQmUrGlAzdxh+0JIUI7XxV0RPEBUDOS8qyN0HZ0Jb2Zy50gHm4b/
BLNqHqCwFtoYBN+XmeKveDTheeMsrDpzS1iDIy+n2hr2r+mZm557qrMAsXElKu56
677XMWXvW/A1lNgmc8GlI3vQ6Q0wkgxCM4LQ5gZ37M/eYSg+/OIKgbmcRKpt9bJR
jDhR61UrqUG5uzVQod1j+4VfA5Eho6DNAfD0SaMqGIY39E1fM68QSDwsW8jv2W/y
GM+n1Irx8QGQv9J/WpbCx5ImyAJ4pSf4pcPBWJ/3TeA9guBz0d8OtW4rafj13t58
3m0tEAQAvGtTXvN2xbM69SvMlYOJd2tNv+AQ49TQox3RY+VczLvz3Ol/7BTsrahd
SCj7UojsjBUHVIK5ZwKSIsNU8ozv+ouDwrQUaror3bE+1u0wXzaEOO3ab/zWdwVr
LxUKmI0Gv9c7Emri+mOsFojsEKiZM3C+eLpzjPM2BfuPhl2H9QNlD/jfViAAd+UE
31sRC/NkLi1jZF1M+ZxfIdTvZ3djKXPk7QDEAOqxAPQz9M6YAymkigY/YmWa3pcu
KJnJLfb9f85VQBckokLR4XtyQ1lSvn6/uSS2+EXYKhqZzHwM2Br4qTs7KwqkM/Eg
AM6K5b6P1PiFWJKF5Qd+3hCPUyRbGV54HziAXaEgL+SKCjv/YG27Zo5f4VFu9PDl
xlFvFHH3YqXsSP4a8XRsARoGZ8H1aLgV6XEUOyWAACbegh9VJA3m+3oSCRItbgad
tP4HQUWUENy4GF4cmci7TNYMFxjnvKNo06zHdmWUDxt59QiyzXX9tkGK5j48FR68
YrpYc0kxneHC7V+SFvOIAjluldSVnazmfgm52ZMLksQWjQYmfjHCUrWTq+0UhCPT
WpY3yHi4+DkWwhKfgR/BRdhsiwSlN3BX46rNppsC4X9eKGOO1giVPmazbad3WI1N
Ww7nd/JWupYMkB+dJbPM5j1ZHzIhHk3UZIE7WHnHX4a0M696U1Rp2balJFJptJ/9
izaNdKWd9zAVRBQk/QUUam5LNjfiubwql1Cc8uxc5lyXY9oQCtT9M7UgQcukkLQs
xb207057xWz5jKUZ5Y7I66PA2EnjOdBV4EzuuBWvR10qaynKDdT/gV4OxhK14yki
cOXyX8bIdePI3Iy1e5D/XQLRCfUhDhaw5uSP69mPmYAfQilc4i/w+GA9cs7OlCBI
7oHilMVEGpaLOo4Xrw7W2Pth5d2wrh5IYnHoPaTsioeUA+Z/TE7Qa3sMXxbXqVKu
t0GhejH77PU66adUDvPlqbZZF5FO6yt2a4E74ezBWbVI5C0Epoy5B7izlcvUGJFQ
J5lxjdlfsS/FrMOtA9oJgP+vfXus5UCbnIfa7O4U/dW29YRsNrdqUXKPYwJNNsT7
O4bCoTP56lXLla1PVdVYQiOXmUmLuhDsYimSMQkt5EEK7Qv9fTE3pUd7nlhSbtaK
udByv+hIWq07PrHWtDtQcAXuICsb3mfseY9KSSjRYykcaGa6FnQJ13WlQ3KGW8Qw
mZGF9gz/DxtPv5L51nwnnECGIZeJitfVF5JkuzuGNeMJodAmi6tZ0MVfYD7jH97d
9vybOp4FCed4cuGfPQtOKznwPXhwBgU+K97oZWTmgA4gM2CUYFFfVkfF4OnR2LcF
1ITdFHLj968DJ+40syT8URUqmeNBrIkK6w/5ORHYNFcTaCx5NgZoNoU0UMNAGJ5v
K5UzrKkyJSvpGOeBn1esIYRzCAApsbLLlUnhPsyl0zsI0g6al5BqXeYyZLPiZYAj
jkFFz2ZyBFhxuD9VoEzXLwPlHx/yTtm/u5QPheGUxfqQkqQ5MahxgScY5RdLy91E
FWF8OWblZTVOSoQ83AsEt/R4iiYB7WrAT/3pZ4ONiqnbRaqo3qRnonTw0cvw+0zC
4EHQghTHpeqAWRl+kBSp75BHQbBkoYW1tjPUpi2E3bU9ZnTMatq6VUgFEcrXJMKz
lO27aB8Brc57XuKZErDZj4mCIUOAVCfRfPkBMQsxpoTzMn3S/GoQmIOr6QmuC1yV
ZJ40NfdVy5fIgmXlVC0+0NWzo1fJAJ1v1oBBTtsPTsaLAJ1auAqQZ85cjqTsyWak
ZiQIKx1m2JYXEDHrmtq3w3hfYYAv7wNlbEhb+QGvXShqbSUHcuhAwfI9R7a+A8s8
s6e2eMDwiClk2jHJ+b6CKTctlg0piZGrJhhQ8g8QhcLVBUnBkAFHz9mZvSik5o4i
YQv4M+GJaoyyyytcxu2lG545GEpT+FY7isA2/lbWsoNw3c/C6pDKU9FUU4pWLmtz
32KSjjxNatFKw2wcxSviMaA481JgECFUNrb4fYux6NygeGEMx7v2ENH8krqmFGjK
4l6muiPYwrx5/k0y/PDvkBf4cYVzJSghaGfd/D+6wslElUdpIjavo7LV3LJQgnrH
PtJ3GHJOctlguInHeN/h0I5dXNGXyYh0UzKviuAx8q3wOxEWeTMRwB0cOvtGuIlP
aPUrCurVvPmRH79ZZy/PhueKBSV4YMKCY2J5R3P3EDW1w7Lrv7DO6N8qgADZkg1T
SXQk6A3ZyElxA1d5zpvSH6XNG6X40xrKN6pzXlXQ1UMNcIRU82B+W1t9/Ra/Gees
jQYZSoRRnKHIi88uSW+BfUJ0p5rsojCVL9wlgSpkwGFX8CDOdsqbyR/lZVqRTB7B
F3UkzWFZ9+K7tsXBqjfMkGZEmW1ZbyN2ui0rNufQyqaLsnEb01I+CIR8N/Qm0jiy
xfJkudLKNt2kVGM0VxLpx/fL8m4i7wShaxBr21nRYSOekcMZQG3HCDtRENCm0Il7
WxO0TnDaNkqr5R3cFH7yiESQcix4hEvqW3Tl+QaA/zVWx+MXSxeDnTK7S5hdwSuA
sPpO6K7+wCVqaVOf+zSDdj3cdzM0vpF8I3VZgr+XziAiiMKWrCJJF+djXURBa0kz
6zMBna5EVcEScTG1fNU0CggZnXN+lw6KxGxBrJkvr1J3pBC0LW5HPdBTHZwtiwFv
R9MaJh7Abya5rUfL4P7PqcCOmh+AvnJI9TClhq/x43AsDpVA1gJx9vWKVEC3CrUH
/ZBmde3jo0JqI5KgFFA2OxSnRpRcxaLGxE09Lg6f5fqYI45VrCjgNGam9NTglXXk
MumNQmGmGslTGJxIdl1bqNyEhkpB/3dZ8YhGEuY9exR1Y1nEkNU0en2wnN5I2PIV
z6EH/Pf4FLMdlOuuaey4StZ0sJcniydI5WBbbnN2o6LcTKvKcjiXuuygjnJGB/rY
lxCllyWq4TmiwXNh2GxTLQ+yROycduL8GX8Bdm9cOtMBbdUNK9U+/4R+dlvlAfiM
kyBQjqCokOp4RShXSc60jb1p/Wn9X6FQX4NbHJqVQTyYtLRSnCBpK3RgKa5W5/wZ
0x5R5mMPReSMTZ6DFeRRje0WzZfF9VgXA0XmtzXLN7s+kkBqDAoHw7lrDTB6AUaV
qNUsU1AR0BH0XNgtLGf4GVABsI7c0zdxpNBNe93AT4RTL1z7F3TFoMy5LOAJJsCb
Sv309Za29MWIoXfLlo/15Fb31wc0uDB2OOEDwj/nPehruYUDlfM7hkkIglKJeaYm
jK9tvfrQV1xnbQdBJktwQYvT4kH/3CSniojnoE4rCYp3hL5Md9ijMjFLXTWDtl3J
UFQUiLGHJtJkW0XB8fOLs9tTxW3XjNJfYfTjoomTB4NGGhfTW6R1VsRnryIpSrp9
3Xpr/KAqTgvjNEnZHqqaMdYMlJzyc0DR91sOLfafKVixqRpnTVy649kwdNStTcmz
dS0PqStavK7d/kxktMtQ97FYE+CZmHZVMi627wn7gACl55dP/Gcccm0g0KJ02MRt
0lApvkLNRDP8azCSQS1a/47JhbAhQdc+ZQ3Av7nlYgjsEqOxO8D+PXGsLZqCfjC2
Dd1BBohYLThwV6Kj7EmPi6HVTE+RwSdJwzESCO0/Dq9nMOQDgExgfcV6mDCEQ29b
NVRx85Ce4djxTgVGPgEzDyDg7FKTlkxWpa2990UlsGXnJzweXahXgFvbArOwzxSl
d8B8DHF2GM53OhX2gK+weJp1Zx0PBMk8bMSFj50C9FS0btssmbYXSaOc4FTHqv2P
rnlcXBM8qnqrqO0IhRd/ewB29eR4MTACweVxqGZ50xYG+U9l01RRbZ5BW6NGaUvI
hxyXNnLbKZ14kMcGJzprhEsFQouVvfawj6uIZ0Y0alsyxkJFAmrjy2NQWDggOUVa
wyrutVk5hmo+oV7+tsN0i6gRPMqNgK8ZkNyIMNH5B2cdNLhH6H0GOiAfTsmKp8pX
tSafpcYkdhD7zw+8GBAAPGAixPaRff1cvMBwBULy1whzzCACjvhhac023s8+/iu3
HFyEZAYvqaFQ7uHFdGbytJZuX3fH1LJYCCrQ64ieWPRchS9fQwf0J/O3VNpJdWop
X0dghaEBW+Bs85earHP3wrPRNu29RCwtbaGAsPvs9ydX+v6K+V1GzlIVT/tgFQNw
JIOGknE915+v8C5ovXFeSKSo7ONQutaJmt/mCKBhSvJW0s7jIEEelyVQ4tmjmb5J
kfsUz/NKDXpZ7WI4Y7A7yoBWFLgxZm5ScAy/DTJDw433pQv5vqDzrlTTKdkZVfA7
BhQb6lm88k6KgxxIa7StmyY545c2AXH9ExSAd9DyREEL0wCz9RL26TbW+7WJvzUi
bA77qCZ+UDlnoLU8lDUCTWLgaAnvYgxlmcjOTgdf91yiP3YLG/0xPJy/DJ4LgRRg
gVGN9aCAEfPRHw/lBEFl5nzyWpzDqpFKx1/Io2OZeGGYhHBUA9p2bcC8hlNwlT67
3y6vDuGu0FqTJV4xGohzM+BMkD4nEZaQz+jFe+OVN0mbtqKyFbAQMgaLzhrpD+tQ
zI25D39K6Yd8ieqPt7UWXwIdYbFZxdhCmQb1sowX1pqBvxLT4QjmZDdTAq6dpcQk
I9b+WMaur0qfhCyERRbR5tFZI3xJjeTzve8rShbh0tfmQbLANyqTVV/CuLyG5DNz
/rjCs3fOGaOknPRdqD/9D00swzo6vvtA/wbyDinqNRbroRFTz4ZqJEiHTxIvXz1l
VlaAPY3llyHdXOoGFycqgz7tw8cHmOd4/PITU8O4wkvUGRaIqXWwtoj50atm/6Bl
m0/j/1QCZ5vlgFfhtXjJqSXaG6pB3FlUlSAUy9PoFwpR7+i5hSPVhAbdS7nWL2gT
nbLPMiJIM/9Kw31aaeYdcngVIUWSoYg17zFttJEwHRYVlEbF+ooqfmcqcUf2gDJR
yLFAqmk8Ii56W71/LmvfhhnxXeQzppVJuu9A6ttcc826N6s8Hc55FtfOhabZ0KPL
Xg6CktUrzoP2xxCF+Ch0fmUTntIkD39Re5tlXckOLwagsrRvVAMHI8WHcD6UOxPg
a/i24k4s7A2yRZBzNmsVc+NnqHiEJyJHX5XTx1wgg5YIpLj3RbYptaYwp+3VRChW
ohaE6o8wpovA7mE1gkq5ErbH1D825zy50JsjgI1D2uSBBnGoqHR21I9pw0TeA/PI
OVG9ZyX8UUihpXQTABEXSX97VsTycSJs5wB5q5PiDfMSPdBYGLJPJP21zyy9Eh6h
kGIp9DY8+RPrpzIFq63K9MhEmRjhky4brnpR2wpet/er0Q3EKrNM+sgZnPU5focy
lYXQHuqQUYbk/NnNOsNAeRkWR6A/YpAksNMpdiEq0n3+5gzf08CsFOPKZ8I70mMl
tDfRrxkFpJQ4CdLyOO4Mdel8DLBzqBXJx5GcK4xOmKNYRnA/j+HDUGp9WL+SjezE
4l5pBmCols8a2K5OXFApFYH3dGJm7fGqypsoodxWrxKr1PgnVvAm+U+knGyAK2t6
w04pMj76vC5XFkAegYUco0ctvj1TKYtLcX+z88yup4r2SJEs3ytnXxzNXhr1xp9Z
ihrYVRK9g3LwDzOkB4JwgrmLIrtP4dUXH0k5by8zZWHa/Ip4SwCPoNCw7uHQ99aN
0ZVjOWuu8h+GyPoZp+7Qm7MgHYnpQRY/VKR4S8LUZyvH/W0Jv8aZpHmclXBxRpcb
l68I16lAufarojHWkZ6HZiFOapf5KlJ1inHaxFK4A88/3JqgEcefcnAABLL9n6X6
kzMWojKWGvGKtv9eKI/yf5cLm2L5MkZNS9xXGnmdhX9ihrlrahZ1eHiKXSKs3Y1a
kic/ajb91XCRTBnt2JFw5I9PYlPbzkiJdhfi+XqpI5TWlix8J5lj6U4RulUFUJ1X
stNw/jgXYHYhp2F1ErrAmm+O4WHXnmL5NUF7+TDgbt4YvOU8QyaB3hhHAXZNrptL
AquK5VMTUydjg4PlBHJIlAzvyW/rLd46D8vTUb6BgPuLVXrcS3PKpw27oBQRztg3
nXXbdcRurY9HIivTKqayx8x3jmnSVHWoK7vRDxhRFcTKK79eKc7lureJJxcH4+JS
fvQRd5CvU/KD76bNAMCdJgNpsdth+BjVdZLXOiux1QYC6qnMUg8vLcFfqcsimf7E
cBTihEaIB5gBl/dlj8A7INUC/CzCrp3Sl3siRkyjziYce8Z5M7W1EghoX09XGS69
gVOb49gJ+tpvjtyYX8yctuE7RvwR7CRXU/rzpp5luYqrqQxtZoSlMF7HQSetbF4O
zt/T7YX/N1M9cMCjf+RqIONkeig9E4o3J9XwLNjJv7NN8dWkw/jL9VeFLsXj+lI0
MHtGBGwBUWk/jQGaWv+5Em/cB0YcnFckgiQoO9mS56+XT2Si5kJPtWv8sFB36lt3
gsLS6os8oMjnULbm5T5l6ZPfsLekF96XsuQDpZgo6/qfRB58jLYFpD5tOPj3c+wM
+hGa4Ywq86Fw+0IzwLHswRgmxB3nqXczYjEreY+wKOklRcbEYvLo4tB3C3SBlfE8
XbI2W3pxnOjQJ7vGjjV7Fq0Hp6GRi9A4KesFzrIQDUUDO8QCI4gR82AD4ucEfwkU
kACcbfR4u+hOaD+u4k+esfIb09TkUXc1p2Qipao3zzxVUfDQy0ki3HcZ6wfPzAPR
EZJy1pU8vNQGcfzCIR9xxTlbg4spK/rkkN7+WHwG09kCARFyUE5WBiIfg1Q9tU6E
eleL/32obGKBW+V4o6H3i2o0jXW1ePxtoBxv6b2dPw3CJ+LRPW9g+IhdMsDgCJHS
b6An2584IQvfvYGIz5g5+oHe97H2CtL9imIoT5LWVeXD3HD81VHJ45PD6LJ8Cs2B
JFU4gsc2WFWLEW98R09DIwFihh1ZYaCUDGIcbfaQ1WNAdx39ojWCwEkFVIjCZ/cM
SRQAfQQrECewyOUsPB4blHM32ArGu2pDKhXVPTWFWy0xdvQyWt2mMHKZ9KuROv7K
FN95HC1mHHR6gWeb27aWzTSwvLmH3TvLE7OzYxDCbJMmFmLaEoqGESzMLhN9ZqnB
WRyBWk7oKDLMnMAjfSwNcyOYLBFp+z5kH4Cm63n1SaB6S+r4V1fGcqBxEXgKIOKA
ljWvYRj3rUVHCLSfmUvUW5pbOe1HNs0f2s1cUfrovqARZlmDSRTSutFQw2NwGwX3
Z1oAcYGipVYXON1b7qm67ZVOOANAnNJZLLCWJewRfl1VoB5R9Hdxi42ncYp5A/Vy
2nntaP5H/4yksmPpi/ZXXxMp2O1n4q9DQjhcU35iDLZGj5m7zEnvEeVHvTctPeNI
P0tiUzGHVxsrldyWkycJNL9NxWswC4KU5QGW+1lHLpE15bZspd7vqNjjkdN3MJxh
apxeIA/lWNYS1i5yLCiSg4Sj6kT+Iz9CXKGkg4D9dZcVDotfswsK3PoSM1xrSeDU
rFmf9ZVChy8/k/W1ISLSDr3IqbEXwwNnstCLNle+iG1rWnb00qppGFwEPDDOazZv
bFFCfZ0NSIkuqTUT5RcizbmhNTgKnp/UWrdQqd9OD6x7iMVGEsPHIVMTHkhlCcRU
pF37Ua9QBNaH0dO3hObuzzKFw11tttz/tBQ340pNtrV08ENF/Yxy6Gk5uYzRj11+
flQBvhmm0pjU8n5XcXmymiap4sH4Ow2f6Vpdbk09Hx3kALpQ4xyrjdV8VYZ/UZsl
d6RW2QzeXn/+C0NaYRi5mqXkpjfDl9LFT26yfUmDJldBFjuvG2W7N3d03n7qgQVF
yF4mj+q3z/7T1kJZXKEGZr5JKOIXwFaaa/NPyu1uf/jFsFSzRoe86Qldwlti3QVA
HgZmTt7LuRQiBcLfIH2oUU2aqvqmUO4OalKCE4uTpH6v1VGgvCgBYhTHGia7PNP9
eNcWiT1W1/t+i9L/spbXxFJZ0r34yWONu4foMjlFKfowHwBBhdOjWhGN7Jb6I2nj
tjXmZkLmAnCc31RyuJL3sNjmnPFUUbNJjdnexp9ovkjPyUW61+Er40HQ8g0I+PKH
B4ZMHfNxJEOUVl+1S3t5U/dVFJUsOvlPK5W2Fzy79mfPSSGU7yUllftHlhoDvd+2
UcpcLtuYVQVbalIYk6+WoRL2dsSebnLLxe/ubwYH0mIuGhQ+d98II99KCFFRq/ab
XLF3YdPt38yzSme+HE8PJn2Iek4QDC/Cpq9vJFibpypvfZ/pREE4tZw5cafHwVpx
kb7AMSp4F4le1fqdx6rmV5bYmsAVjrIC5MZkmSlzLcITXAzSjFZy5yPI5a7ADKcy
n88RT91Oc4aOpsEBBvxdwVLKu6esXkWCxwldZxFxi6Zl1yCfxwVG3t3Lqn1yH3RM
MHRcty+Zm28BNPUIKGZHRXXhKc0SC266y+I/quLdIoK5u9QMsvpEIXP2XpMgLPCQ
E9vDj8Ca2KyNIl0vEEtJlmbbmMyZGeDgtWSJr1YkOZX3g7eu+WinvsdIKRLw2/bb
mw1zfejO8TVNSrx23CY8jWl2AydBM4WNmVcSL+kuN5xMx9u2CVSaJvfg1f31SfBc
RD9suWRwnKSjVg4cnIurVFMbW8H57SEZ9RWafiw+1jJoAp3zdy97xpILh1dDYb2K
r0IIPP49S3D84CyOpfZ5wu3AR3c5SyQw8JEPtl7JEeA53K1USWiedJBlUpwnYZjF
c6ETVpylufJqtjUi457NlhAq/sMRQ3Ysmw4AzpGRMKWQWcu8Hl6WBubT4242Ygl5
iSkjl4l8lapd55CKnm6u1lFEAh6h3NCBFRdXOdM6L/A6FMNvfIkwMjlfAldQkr6f
LX2ZblUY8UHSX2TvSVV3JYugKYB9j2zugzNaqAOg2Sgfflu7F4jM9u8bwjJdD779
EkZiYnqdiqpeA2Up/TARjNdX96wFetreJbBnLhfcHud6x+7hRCcIML/5Pp+YGhtq
FtoS7/9QhKgoFhkh1eacjIsKgGv+mbj/LugG5L3F+YIdjZoFcWX70IOJC8Pe0psz
vezYezpE1njsoyzq19m2WCMMlXYkKRt0/LltVR0rqOTMbOIl1dd1tErZpjRpGOOm
s0SH7ivgwt80F+dRQRwr1lrKFnPFb+XxAryIYWNbeUtE0ZGDqarGeRbFD9AMTRoy
FuEkqLhHRN00CVAlOeemmkxsgauYEn+5m6viiQgbaQzQSzZxp495eO7h8N/oaIBG
XXTHexrIC13LVKL1lf7zD02pthtDvc+Ac5z9+w812HDfaL2wNw9kdIXZlfmt6ZNE
GzwZGn4FPXXyV1dcUOeCr+2pXR3q2nUxUvIVv8+rH193zTLM06I0S6XmBQObRtka
rCFQ5wCHKE9mZdoq1tiwByOndJGoPdvkpTPFWBEUA5guXJnEJx0it+NpNKoAn29C
EzLey9XX5+A4OkCzTD7iY5lCzdx+JvCo7WpK67LeLkrWPNfgPKhsBd0tVmZFUYVb
7u94/6xEj0CnFSSAh9nK4AEoumpg6Wjv+y5nVrXRdRsx7ezYF/kfFWLm8JsS46oX
wVU/niVsEhHKqmyrLdlIOFBpNdPZyixPMWF6V++ngS+/VAYnvpW4rjWq6DKCSqfG
+YfHeaGo+4wL6R8d11sW2XKESHreSwot3Gh7xwkrBDew3wxeW7eKZoI/++lUtsx8
AfFfldZaZuf8gs+mkSCprpLjMQK3ATCUa6CRgRZXFcOBiB1VXX/h3nU5o7fF80ae
s8QqYNwurh3D7pL+ZANtVMUTdH2+hcQWSl9Hw6aELfTEOqXzdhj8eHgtGY6abuuR
ZsJPtrsfUTUAOAU21LF9yPVKnfJ9aGarjXaFo98gpKcxr/PzO3oKtuLeb+dX5xF0
64672vX+74ULypRISyxPhJrzWOBIV2yDithdztXYelplULotJ9r0Mlj8ZuWEM6C/
mak8KyyLuLyZVKRKfdcaMvjXqCwO2LjgdPPDXc8mQo/hV/CPy7g0MbP/D7NS6gu9
v/mQQcdTbW1tOVVyIa7bHQNuijpZy/yIJH4dI8hTKDAIUyB3Gd9KSRHnlnkq0jKJ
aZ0o6AfKGcKReDPMNvHMpMmWi9Q/8g84zHSJ17jYBx77P2F4aoXb7zey7CCFOWzk
dTQtLklCLsIfwaV5ViCt53v+sqcddMPsZmOVy7gQpxPJfPJzvWtOsDkWS074XZyB
GMzbtOVjmz946slEJs5+sPIZIuZvPdr5AkyHkf5arx28uN7x0qwqh+e3Q495SIAo
IfQ/aG1zwDZeubRCHxUs+J5Qvo5MrgVrdydLrAEu5oDVqSILycg0u+FXRaLbBKbv
l5LIQIPvjo70osdvb5oyLJUVTarVzj/1kGgvGjO5Nuw8tj82la/3169rnjcqcls4
4wcKVN4SfkJfDuakoLYp05GjGtm0t6rICY3if9Afax29r47M92NuT5z024K+t+G6
w3ixqA9pWetMCnJgI3VCI8GzB6hyqww9seOPSDGPk8GsHsYpF0+MxFEAQzZK0xUu
+vtYj9b+usQrL5gU+Am5ip+suUd9UXbWNdIQRnL+LGPwlMVJqH0x/ECwG01EDRrr
H1f85W/rJT5KjJ1vDAj+PDVdYJdz0fShqy9tqVuXrC6qn7vhJ4fHbp14l39Se5Uu
Bz1L9/Iv88sAHzUm+bE2lq0aNGlIvP94P6Y8hfosK1si+aX8jeuWYMsNBTyMGY4w
FsysrJEz+gMsSnxoA1bOxHciumslUf1hjmnQC2Vq8spj+M+/4/E0auZrP4DhgtUT
EKWLDnsdhpwnxDlJEZ3qKid2g4UsEaqksnn0q0BeLTK/O3nbnryabvFM0gxh3LE4
iLCrlZaVzw0KwppE5wjC46z11o56B06b8UZ4wF5hKN8ZfisrD0EcPaUIST7TpEPp
O+TX5I6onlU8RQKzrFDXAFFKpsG/jhlJujOeqC36EfX0HYRiJSSE3veauq0qYtR6
wStUT36HQoBuGKeJtzU+aBVFDobppQ0HTkN3FzMG5gpsimdx0a0QR5vBMfphoL1I
a+FDn0pWaR9VQ2nemz0GnMnTSgLPtCccwwH6fZGl6RJTuzkV0ahxyQYTK9DsxZSE
GuM7n3ZLTTUjZGKaWew/W8pqp4XzMMas3uRBQO8PKAN97x/Bh9H46xKiJV4Dako2
FCYU62Baduy0WFmBocZKZbrSR/1frLs9rKPmknb8liuIHdlhB2q2jG9yIIk1G6qh
uSGzVUcDYQiiJY55cjgaKk8bTupaQsNb8FKBNqhfyygC2u3VbmfORijqxr4xzuce
PrD8wOMz7g8FW/d1ZSUQYQwQtjfYzAFKDNs2O4b7Vo2dGWVy4VL22kucuBruQQgJ
tQEGs2FbpYFt8vORKSw40zPnyaEEoOclqRmo8oDAoZRbP39U+rIAsLpHF4WHzWGX
A2X/rQJSeNNfbtIBuNSuzpSEfw7c5OobrcQpcodqXhukYHi+LiHYSx/4Fvuw2GPc
C72ltpfb2OU/5yXfaONZv/TzhzCFrc8LaJKZgP9SgcNFFHE7CUCyAny29h5Sx8rj
ulQIR8OXH2t8Yx5m2t/80SPeXFh9QLkEsa0Jb6lqGVn8T1XtDoqjIoYQwYjqer0Q
Y+I/Lr5vTcm6B0JwhWaLCvhRYpyhOKijM/kgiht5m44UzR22J5TLKOQRsQgBGOYq
mLXxHNOWXshgZcjUfi4kL1RTUi2/Blx0hMkJuuv/oTeMNgYikU8ZGjEk4a6G8ZBn
bFDgnx5iMKMMXJrtd66i+TsWIbdt7VpOd3NvgxyE0wI0f3Hm9tXg6HkRTqg2kHaG
fYTj3XJ/zWPkD9ay+t6P50f1Uwg1Xz0g0nRdiphPGukZA/pqsQuEIJURjD/u1EMt
fpBccy4MjvgosU5LjtePKvatQXTHSdHhylvLPWlny6iSjMejqTR8URgQOVPSUFVZ
8+obanN3r+DuylP9I5VwGsyk9Y0ev+kNpHc7C4wxvuUqn2Or+ioMfLt+x7gLst7R
IE9H68VBcMkKeDhLecNwqouNk1SZSaKrVeJc61E0CULNnlXyWXH3HhWFo3zQHKfa
2dBTJqWFZazy486vQGPYSrIjWWGsOuQICvJpuBRI2I+SZWc+ztgCsJt5ix4rjlWM
EG14jKfDbcHTduS0ovRdfnA/CqEvKoSV3vDU2Aba8k6wZP4pRIYUMO6NbF2GlY/P
cmr+ssJkP0gFIxOOuQqudSrCFwtEJNQgFVKgoiQh3zOXcRuicKXZrtAxEyvaGDPv
LT9lpFZv3CVNF/OmKEJytp2Q52d/CmpuymmW272yQVC6+9hO2oNc5Z+JAi2nex9d
uRqERcRn2dWZX3kIka8PbdSBcjG8MA253LeUk8vyM4FJdbEND/vOD9Qhz/DV2X1z
t/Vtlqcre5rCEEAXg+qewvXY9gyIfBfN0YKYoiHcQhr2IGFiutQp/j4h+qT7dPV/
3hJU1meVrSesDmw4dFCJvEKaLWklfuY5fx9xefmjoC3kMjZdeyMEFa3OQm1NyqJj
sbQbUcXeE+G4r0vxtBC1zxzYJ0bgff1EHyVNHWvIjWXy5KbC9+htDeVLwKLZ9LDd
dstkfa0mSr8ksm7fIFvQwtmo1XnsrnBcH8Vj1ux+mhFOUMYoZpyHMaREJwHqBADH
/0OUpq4FXexUFhCwN8KUAe/MgGdT5qkD7hH3BA5228TbeuGs1s0eKqDW1q7qxsW6
dOlXsUrTKvKPnPyqXjNw/i7XNYCNPo6w6YfAeyAYJIh4pfT5P6vHTZs27qusCUxn
KL3uz7rmk+L5wmLZ6iemZVzRH/TibfbPMDKaLGsRSIa5t/HU/JnreHOJZ7o4dyON
lG/CQ27UDmqN25+zWqvEiM8fjFVXzR4U1lSnKbJAPXSDIygRb4Syfq0inoWGeYk6
2RH2N0ulV9cPS7zULH5ppzg0qiZM7NcFebZhtZttmPNPJ0J3fxs6ZDX2pd0vGJN0
SC7K5nPeG+2Ygnw9DT79CXLR9BN4pY8QS8lWu8qFFu1bm994UCt+MauYmlWHECNR
1jG3Lx56U7/GBxshvakoSy8sNUAxXMFeKMHpr3Z+4wMYgbfOz3MDa8nwaRgOzu6y
9Rg74Uvb2JT0XPXW5zl6Qo8a93SqkijFu63txsHSkEYvkNiX5y2nkQ77GFvo6Idk
3Ha9iEVmb6SeJUq0B3bSNWbHuJL1/HdM95fjIIuOmdXFrjzwpj2+s9EQYwLV4dW4
HiaBuluBIkppz0PJT8YVMrB8QraPlf1EXhrfPCDszTdAL/BOM2oqqL3hBRtSySFg
TlNHw+lrVFNkPwjtGPDZNaUa6f03Wodz0CDoI9pgNfowc5ZTlqW1j33VnJ1NirCl
8TYrrVVrnYpQVQ3dD4hzi8irIGjT9mWUp3Kg8TRVuFQnCrBIaxIltRIZvO366X9O
Dv9uYfq4Jz/6jf9bFMikaV2SrUiCqyTRuOM4Y6ohjS0hyYsYbl3XwxMCPq+1WLsH
GobwSdNmWEJv4L28f4Xo0bIdO3Dw7F98jWUsnQX0DhLPws6OBpl76SkQkWal/f3e
okKV8lB9DcBpJnk8z23t0TzK7YYw9jf5ank7MjCd23zuQV+pO32mQ/xUCZ1oo+hN
yBYTvbR6/v51qqirhoe8n5/jBP/O2FNTMVLUJdoOva9qdwJopNJKzpvliqq8OMr/
DqFftEBaq/SkARo85/UCApvEFopJqD2Wel8FDT0h92jW1ly6ji025ipJc/BAB4/t
lSG/YTq+KflcnwFWIaJ+H/QOWwNVlENAVOpkcGntTLPhTwXQR7RRx6wrjP3DSt+1
i97536lbgXw35QPEHz5sDdiWrk/9newQ4O8TSzWYz7HVjt72R7v/cKkUD87Ngogb
8TCGe5WLj1Y1UmhNxr9Grs1ih32HDJ41mQg541sgOSMdBFnQxgzPJxn9FQHW0vkZ
jBzQCdBaNQvzpLQ7kTtI9BEVYF7aE44GnWN9klb61Kt9BslxZywtjmeceKEHj8Py
KxDUK4uB9H+BW9bvU749qXvUYy3D46axKM2ngstpoV9fWJ0+0LxhRKxTIl85/Pbg
aVHSc+7HwOefNV7yGOKQ3RV0wMUFaVjlxHkRix52Szl7ax0ea7AZ4oy8Be8E8Xa0
nYNjeFaa7QRI0b4D5txoTLB588RzJk+eVe552OlgJLttxpnjP2WszYwga3obr6IO
sJoReh2vV4zhMcrWsoIJymsLWpd4t6aMmdXWl3FHpaEjTNuz9D0MawRu1EjeNL5C
YhLyJTTelS90azS9xVv7oR4ifhwDo9Obx+VoOx/5/Vp7W+YWjC0bP6CXmkZeQVFL
t/oJfQweTRh4CaAdUtMX25GM1B/XQJa3+swqB7DUkOudRpgmPXxJ8zvIRvVSB+vc
7rGJm/0i77gC8lgANbirlzBLZAKXOpwobgdlHhoKXChZeFFzXoJPp1VcN3WC0tbV
6QW4xmTJ4ScENCeM24BXkWhq9RyXhADgMxlY5cLmaEBaaVsvs5JeqSe59p1yHVbh
2OLC0/bylbGI8ej4J61n/i3dsOE4aOCzZFAqbU7I0mdBl/xS8xY2UAJUd7MqWjc0
clIpeJZUYerBQ5HQlWWujeIRBeCa+8xoSCDAOX7v8FJAZM/RxifSM4lDQhHwDhQn
9TF6R26Sb+OnrixRnWeI28E/ZESa5Cvdn+CeKgPx6Jza6t6JW82sPTD63ATYu5/K
QcoYyeAx+CuPzXn8PqEjcC9J32ZtcUyEagt86RC/0F9FIoG2Swvj2n5cTPdc8EMM
eL5jl5x0HoDlyWXizt4l0dNFb9hch+NB7JmvdDcYpd2W0l9IdQNe8GaalboX0/3o
0+MsiZX5Rcm9txd5PoReywrjFfSSPm2QNd8E0LqoPDeYX3IY5r5ZBgJCzQfQrLan
PvnOVn0cJ2gMa/HDdxYEwDAVgCBlxBaWzVaxREIGcby0UnQ2Hwaw36IhEvzbr4wQ
MCCIuzt0Tsczd77JQ3QpwgRhrhkkWaEcS/gq2BmZOwcS1W5gISGEHdMsL3Aui70b
e+wHgk7Vj/WB5HvU/0jQGPCPDfJuaUSl/YLn626oKfpFdfvxb1QYm6vj99cHnJjG
+r6lO+RWB5dEST9h8+RO9SW07p6kAZrlLb62HFu5igR8b7GXlgNT9E3ue9zb72/O
pFN8VQ2UPLnIHUkcguFW/N6sHJEcXntxOdGRy8XRYsZtmJS/UHxwmz2U/6R2JWF+
5boI4Hx+HxiPx/U1qLlOLO5py29MjzEQ7pIVWhIC+o+FaBmU4GLOfB5q6Ls8u6iZ
5+r/jEc5gQXXRe325eUwntFDEGq7JWCGamGmpvvjR4DRqkJo9++RhbBuRP6TZ1aY
Xpx2Mr1I4852DMXj4YIAs66adfyL35bvBHK3epCac5Dr9CxD3/ks6CtK5v9U5nrD
csJ0q59EeqfesPyugD3yxFGdMDvM5mlDsuNPlmo1VB/WNf9uF5mXjDXbq6zkecyp
s9AJp0w5agUV/98Cw8KB7nL5KjGyS/3P81e2j/Dii1zZdvanvOLe8QIIy9CQ9ZP8
O7C3+tj8hJK9km3C5aqg2VbRBh5U8RJdhVBsWHy/xr1aOVN4Tmk7ieOvVGcva2yF
VPR3Vv9TVgXlR33K92B7D2D6Ej0QkRWQQGrlJ3Pe/DdpoCx5U4vBvR9g7HWNn6tF
W26whnzySwDDsP8aIxXG7Y6964+mhsQ/P+qM8fLAjFjTJ5YKwggq/sCSrOx//uTJ
3Ud+G5jPY5r6+m3HcEQXf6bpVuxnxoEdkATfpj2Ny7WbWzridCRZVsCacLbdIkWo
uJM+zcMzec0jGtHtchAyn2aFu74/TNoWDyLqF3nzi8x1gK0oPPVUNjEoSWqxO38F
2HiMPSW1otrAV7MxR9WVGFeKWhichmnSZA0+npD/qOPLJmQCg5F3/393G7EG+qyZ
RubtwixtWBmAN/9hqNutwH5tsLcE03mzto1sCgiRA4W2KGPeJvUDBWPi1QmR9YBc
aWglwlqj/NRGu+QgRnOIf8K1jsLQdFhfVpL2xa4bN0NJhPVC8ZgDrMdGkKUnfsYl
GSMzDsosHjxOCOA2mrKhvakgNG25Xacw+NELYxOe0c9iUNNDleYEZyZSzUp23Xzc
8aEiSCRihFAbqR9K222X0jZgIWbgLFuc8RPo7u6AekixNKZBdX9l0YH8jLzEt4z3
biRHvPOZvsFOYQWsvgv313FSsDFRS58PsV0lPCsB45XXdb3eIo3DW8HFPpIMixE1
X4Vg6d9UNNyzrkCa+oyXcVp6IAPGnh/27ky4LqXvxetOBoCTKw5tmWBJZjkdjg4S
qX95ykLWapgjQ98Pn2umEv0m6u7MJHcZWT91WRNwQPFigwiu+BsONSmxcoDSu/jd
7e1tiJXzIh/2PZDxSEfuvU1iNluWly++3t+v3EOZvvxbs4WAZUHPB23CXud1/wrW
DxEooEZh76yEAk92thpZYjPRqFKyvX1xlkHWaqSJsukGrtOWZLg0mRTxyOhODjbq
sjN7M8qK7vrRc5mVkW+hNbk0S5ViLvwEE83AcoQwCctvu5hh5LJiJT8yDu2x53LQ
uwsgW0vOjyV9KjzOJR7dcRZm5IaOVsK94hU7GUZJ5DVKjKKxBKnXveJ2h8kfVF3e
idPIZkErX0fp50twuyErhyUTU9ETtEN1OltzBZRIYfbttbzTVQwAeqJoNymP3V2D
y1/GupTJnEDRabGdHdyij64GUGhEIGuwUxGtrcJ3Mt9eWlSvKR+pM4+apNhomGIR
Ca3XQzDZa+ACEoA9hBpBoiK2C9irvy1TVLVdMDl6TFoF44VgsJmy4oxG96L18Twp
6IvX0uKoo06Q9lizEeJ5k8AWcAPBLSDr971Or4I3Mdn2WW2YGlUQTllkHBtqAX2Z
Xxcvng3V4pQyvR70/XRS98ZjVCteaM9Y98pPQbzFdvVxvPl7lz5J8pDzo9pJrftI
1CyZIK5piFiUJQTomPcJdw/TAJV8ALCwE+qOYuZZ6eAb/c9H9b2W0pUUTcubivXK
KXTrAnETt46umOALTVlM4KrGp67OoOauPoiR+0yEo1dT9NmEu0tndwhzyoT8CQCn
N2tiE0Hxu5WIVsytWOT/4j3ABYORPfCYqPy4M6gLxVpdQYn+1ZUN+rtC197dc8z4
T040LHE5Gwkt/cR7i4xRtO0Jr3/GMnsbSZyrxus+d48GD+q/hj+y9fn0LjC+swZo
8zZfLepfw2IzhC8Fm9PTj+v81B7QiAtsD2dZYSGz9mGAJ3icK7YIJRRt6xBxDqXF
UpvO1k3ZX3xfhJr+/9c86CF5rHRD6YEQTOwp+tI5Qrtd1kyFwmk9WSjTBoSB8Ppv
9wK88C2cQ/eJpY+Qj2QEx9/+ndMyWyBeIpbUw5sCB+L2/KIlx7xGqvU61UO42xpO
OKrZpfU9DmCus1r3zObgVzemVQ+atwR/4W+vyS7SSiQKbyKe2TrQT++u81kGnPsu
jBYjOgd1BNBKRdsxN2HT3N3U1pe3VuutWxssHVm+RsDBF/fa6JXlUxOPzSefVJHu
Oq1zmMIkMssDrDmTR033bW2ZRPCzqEs9EwUOZ5cjj8hnk8PiPPjDibOuOjeEQC7f
Kr4JfFdJzLCqBJsnJskUJGV4AWKmYQiAhcAfJwjUOttA+SVjjnrPD5sMu2kq1vk4
yiZCs7vN55p01jA50agzzsto381h0MA0t0323+EX+1KzVtYQ0xGKJRb7F70EEKfl
SOwsKe2tT99UwOWtklG/PMDcLLZbhpE/uNVgIgM/wmEKDfNnxD9A9G+x1my57/pA
T+xqTWOcJ62sWHRci6GyBe7xBcvVnE8tf6a372JXnFY7sdbN7JPf1Pk9h1ZZWYW8
Vgu2bHXBGhS6Nbf3M3B7qVL8LM0BZdgDqtieRJvUhGIchA5JLkjKmAsl+ebFOOYJ
mWKeXwKaF3uXTPnayKrmCGH827GDchiD/IvWRlgQagsYNg1jBdMOVifv260pbAks
9Ap0pNN7CzWpkkWZnrsWJ8tkms6xH1DlZKq4KErqv/lVGbyiNpWRTTy/QT5wwkJ/
pcUu+O9eUBtP58UKnozuMjmOI6YXy97mhmXsVcj9M4TaYkEgMuMFW99Bfu8XU9pX
7rdBvoJrLJK1GIxoGqqukB3rwwpYW2+GS2aTHyjlJrYM3OoAIspB9MfvNgC6AA7U
sp33MwmjXYmbjhGIheJYh7Qw3vOQx80YGwHQ+dKoEupOySIMVS7/RkUcyMvbFall
gA5hQhpmKMcZTMEWSUD93yigUr16XUE7Nanhcr66wFTdgTr0bVW36fc2gWmliJ5i
NIVPr0z4ggtmC5HO8tBxuU0aofbLIMZyeJYVfD0z954kz8egfuEKKfPgRqXsY5E4
qODX24kDYtZGvCPTt6c3w8ykqMeIgiigYxJ/lQ8CSX4IM3diGUVYzAkxl/HsEX47
ug/1OgkYGlPjVKM4nfI6SiYn3syo35vgersWaKiC/swlcwlp6whfeFOPT+tBoDrW
MkQ8dV8LXYOHywDL/hFGrM70mOdzXUYdtgtRIBQeG7DiHyL7W9hjo4KvV+wlHMjr
MPlnUndqf8eZOUd8GiWZkhsMITolJ2eXvYcLk1mLzqw7bBB7V0c+CbSxiqNnZAm8
1tNzx2h0wXYf+Q7hwmPakeNS+C1nn9oHfFtbnunhj4bnenDfk9dvqhQvzUgEzx5i
WQQzWpwki1wkPRU5+4OCw5Sx2qF2ZWi8yI2KOq0Md3jlb59SnEFHozRQqGwJpHjF
Dc4K5p01zzuHbLguVEYBp969Raz4DKSk7XztfLbbVSU8+a+SHGcCL28kCFLeuDmh
zSfXpPgWZ8zdXXkXiQGuCwuY652u1P9CwD7YNRkhXcWeAnFuhWYLUpQSFWm6f+V9
1w3BTz0elK2VW9eoBnr3c2gvkvz28/YT6PAGB5CKb6t/AIA5J2doTpIyl6iMRlIZ
BKQ20P5uR2s9cHLBXddY3zWawrNli+wei3UYKBsaAX2xR4SSDPDonzgCCb0gHrqh
2rEI+Iid1VFT3mCeXEi7HOf0Aeyi6AgVvRWCGOVhhKcoSRZeVq+YTXRYRVz7CB8B
0H7gW+lDXB/3wqC8zqiaCOdXfsWL/3Y9bnlargCq0Qe2fOnn522sdv5Uqcm1jpi1
zZ4d1/Wzznvmd84rq8JTk9XBN30QINfoLyiWMZCk2b1MhsjySpuHfQjarKxjEOZM
Jv5Ur7TObUHuC+sk/aCj2MgpTZVOSKgy/xjqlXz/hvO1052kHZOh0ct8WxjiQ8Ii
qxgBiSQj1hW9ovpgqZnikv09aJH6td90qZh7lP9TOwh7USdEftZPbGX53NHyjlzU
XKZhC2yZvzP9WXbcw8AuM758QhGHkPB2cOwxo+3Wj1odYLN0TM2pZOIY26yeKV3E
V/ekQ/dKE/gMRmSLfZaGt5YRTLYLEex4DxVfB7CV9NGu+CgySC0ew2NxPuelgdEF
PYTexTVjK7D1QR9y5O61xBViZK0i4mSG2lLCI2Ybi5hc80Dw+N1Q45IkciBtBcNO
nM1iXel3LzgWJUMy/qBhDJz17Z7fyfq/P4U1NmFm95gyN+RkBLYMS4XwM7BXCkK7
XM+ffqpSSOoJ3sUJdsh75e4QbjpDkSVADJ97cQ/8t1Ly7FW7mM48bJ9szt2rQdck
1me/T4cYMX1vpDcvYjif3MStPYKZoqvWTBiz0qz8YV0zeFVEyk0MFmkypCfqAl9n
ew8jCOKVLrEzCv9kRSYi22AV1UaVHNkt7BmxaYSCyieMNWR1BJA1giaVv2cFsCNn
pLXNXFCDDPSOnpNWY99QJM0wlmznvzONf+jiL9U2MH4kj0Ecva5v/MPlG0W0PG3+
CJetcyO5xW1C+vTCIucb+gGLS5Mbyw3buOJ7Da+lFXSd8HBbiNTY4ze8JOrMiTje
jSNPFoq0deOqEYjHF4Bmwz4HDDO1RcxrakTA84GI1vj+5pkqem3iy37INnYZV/fA
u4vTF+wa6Pv5BBFhzB451xTEiTQbuSteCszLC0LF2Dc/q+AOAZQp1EHwLJdboJFd
y1UnIC/jKe/Ckv3mmiH5aqE6XSZx6h6yeBVABP0Hf/BYKol2NmdEVlYINXb+0n96
Z5vZ2nRbJz0IAEHO2MS/vQtKWjBP1uQqcFa4+Tmollc6MTd8Gh9HPSUlz0jNaxtz
8bERfGskirKh6xu0VYb8NiUlwjRLaQUwuUGLgYjJXGyrAwWcbA2uHkqz1ToFnno+
cZDxPrgqzcf8YGQQGd+j0DHmHIb8+jpAtDt7dmU1daQ+lufAzt6PQil7CZrMo6U3
gJHp9t9ct40BR3UOm2VarMv+vIMXjnNOhcO0gWk8boQQP7bVmWJ48UXVci4ss08L
hBraeEFugEllvOUj0/RJh1uv7NmjuAJZLtboQjjvlRMMDFEFG3YfsICy8RoXAuog
VM1iKDUCqiRqnxcTPeUR6oHWOPcOPUN+3rKagxwx+xLgPen9FElF3mh+xDtTV+Ov
XVShAfxtESeMnXuqW6bp+UGNMYJjDi5bum6lw63Q9DkT17hrTqMi6L/we6qDPMUi
BhiqOEQI6aHUcebmIeI+azce9aRDr/f4wE+4fO0OBTeXCkqHLXVBhMl5adLKJLxa
NUCXe8d2i+xyzddzxOtMSkzl4jzHPSvBs3kz0fKYFCYXWdp66FipwsAxaN0V+XHE
VowjBTf0XbGAfx3JLZia45BgRoCQgioBhuhJFOPHcISGs+26RLD5ZFqHG06iZf/n
JetNtryIjo9w2VH1pzoJjwWDOKIDIYLtOHlGORjVotrVm9hnA+42RpoZqioCa0Jt
6sgBExjPaJmdCxGXn3abxJ2+Um+VINSNoi68gD9e793HUz+ZFl/Jjij9Xl9oeUPH
YPKclfAD88DESuUPpUzyCfwiCDh5BtCTZLRinUDH/hHc9aAtdu4B0nwECD92mmd8
dRCW8oH5D62SYnLL+rS6tEVqyZ6RARhVl4rFcr6k0onDGwHir+/tcFvpIBa2jXzp
uwUeu6ojawOE4J/P6EcAudhQym577tTGjIcIB9IgmDupkFVFIWVuHJXOzhF/bzQ5
N9X0azcrC7U7F0zj5UIbVfE6UufbeNKokJxcBqcK8WbUKQWKlMAme9W1EdPAfyjU
jOpU7GwkLamSKiQXYn7K99TA/ShQkdxltarjppDjEwRtAAuJcPKBdZ7EVOzBVZ4u
0HOWVAD/N7+5Xj37jxOPKMFh5KG1g/vkfgG7Ll+yFeGQKNN1hsPqmRqHUBpHhZ39
MSDHFAzRkXYIqE8wCwIvYQKVjjzsVig+QYTImuOdziX11KrGQ0/AXmvfjeQFFcUd
pDkOIG1ZAx9bL7yihyCj4W2kOqAQZamURcyfPx9f4cekZENtLDk5JqgHQi+DrTiY
OMfLR2KuKfjGpTeh9eYiEBhGeLWDhHAL/JnW7403LyYjyjiusTBEQ+ptbU+NtdJO
7yZoKX3NoTVFJGa4mGAEFBHLEoS0KKfHPK58fHtB6+9U60MUQ+0Ho82pj5Vul2RR
cEUFHluAVBQrMk8q+jMafCbnAe0E6LiHEU9yWG2ak3HZBv42vaYaA/bseVpPvA+s
RKcaCDyUB/vG9dD6Q2NRc9zaCvibup/VQjyYblk9AvwkUcquMYid0W9J8W6Co80p
dk9qzZi0CHaJNv0WwK+m76Yjh4HkNgyUJlFYCbZt9K6Vx5EzQHS8eQ7/nOUPLubG
Pka7P5J1z0N0bTJPBJnlF1mxZe2M9rh4XLxujYC1qcWd9iWTME9du+slRaKFNCZR
atAqQzgswXanmCUF/Q/Fs0T9vTokW11TUJQYWjnNqqPwFBDR2BfPwQ+UcIME2Iet
8jYYVLopG1ya1PTBLNkWuPcoUbZUwDgt+MDuMhZ/dDfpaUUuOiIsDqKwbH4z5G5M
i6HAFO9LFJi7RvfoSg/bwzM4ZyQOUVqn27TvKehKEREJxyRbzC39xOcDS+cGPDyj
JfbBgieDcFu/0G2/AVjN/0WiyYXHCrRgntuWolto7DtDbAZcajhW2OnS8S2AQgmk
f2GyFxXlutVxazlC3bnUVlBdkPZlDKpdgP8FotnfQaNCtHP4Y6zSHQT/sJRLwibp
Xb8AVmjCMV2PMz9tmWaBKq23BtMY2c6d9G+Z5kJKAxyOsWjFSrbot03pU2VI3jGN
1KRLMVZXCGy3DzvjeXbK95HrSkQ2ywJYcXPBFcSdFS2rcInkzFfHqm/oq7L0jerh
2Hf6CBNE5m3cBft2u7NOdTvOwebYGMXMxXVPYvX5c3/0ESyfTzcKj81a2f9DnJK2
gmOMbZ6cVZJuJMz4j67opyJgyGh5CLf/tHuOM2jLjPtAmcIOMmr13XMc1eKUvDB7
oeMzCbrkfdKvXENcCjENXWZbGLOctNcHGDLGwReRGa1W5BVUaQIyC1FaZ2eFBsnn
UiE6m4gmmQdEjOtgONX1wLoymS4ZuYBnC+QCx+XherPjJG0oQCwuMNSJfEOExdp5
AMCrNN5QWGpmgO8anADctftsM/RgvfIt1YRZAX/kh3xhd8F6oBqCeR75bjC62y8I
2/vEMwmsjAorj8jthzDC7EzlynT0RXoeonQwVhLzDc3sFxtAB85DZBXegak+5SUJ
BgEi3cmOi+ZyIbAKmfHrEAdfmyCwfrOqeyv5rZliLfj+0rStMR/MusjLxYLFVB3B
XABGkueXVK6B2YsSY81JvPGsjUqO5Rt7eaxKLWy4OYC6S9j39rKesPrpPe3svNoC
6+U2qtExqvp1u5KL5wWFTI/Aai4lXYp0ej++m+Kc1iBVyt6S2q0IbEmf6VtxCBT0
Oh2GYvDrFRCI5aIMLCqFPMjGs4kd7g0w/zuCrFKtm4lQzStUvSG2uI2FJ0CWGkcX
D2jDnJ+W4Zja0RNNYuv75uAoPfgRIjCnv3LW9k9+ZTUbIFOJK461cO0W3cbNwsMS
ZS4FPna23t5hSeOyRTeRG2gvKZSq3XWTJeG3SP4d4L3GiDPS1htjoJAiIUHseDnc
VfQEMGddjJTMk3oyAMPNl3vcJKc7PSYE8jGo7YyCt2dR/uU2IWXy8PaZp+LuKTHo
PdQRH4Ewe78ioS/82zA0uDRaqE9JiXF2JSFuQA1M1GF63kUDeTWVygofZFbO3TKA
UvQr3xjIgJSl9PAOmtG2ofIraQeY6yqU0/GaZsC2erb9ESGu+bxIYyBTrpy3Yfjk
oU8Vn6s9JkcEtYo/QbOcBQQ7O0tXWCTh27WLJc9OdLTTOEMedI5cJdzbSlg4HbRE
2PqvRopvb4vpWRz0tlkvlL7RxJvZngPNS6ApnBJzIs9vUrJpxrzzkgHrHigPHg3o
yx7Crl3oVnw+BPOgQFUeWg43tRTs1nOHiIwQeYAvPtv+70MT/+ac6eXEVRnhRKuC
ptgymIx9gUaMaZwwlFRjIuiyK3IaWmUqyavL7QiJuLvSskxAqaNzh5xt0BiKdUXu
o27MiHoeqk1XkTaLY+akLT/Vmi3jCTljJm8eED8PlJk7nb56dBnN26141XY/88Hn
J4EfToThPpo5XQ+Q2B7CetJh+NFYPPmlsyMZ7QvpoVEBQ6A1A6RzLxZElFkyNknC
22SnjoDd1g8wDgWkwriOg9sZy4wNw+3eOSO8FssyDLWSvJLASmwAASIFJ2vk5pfM
dVcSc4dE5srNYobMM1SosHZ7JIPu6K1DAYyJRBlu6YdzJv4IBfLhqq0NFN487bvr
jhCxgNZ2LFk9X+mud3u0ieMmo3xxv9PmAnpPr9vNFjOUbtr232slcO/38qiCuZnh
tsY6/81k2whkugCb5LP6q4CO9GDplUQX89MTVZVvKYGnCHu9wuthqHYSN/xVSRq1
n60/ZGvIb0PVQushVTIRRECub4hbogrJmbhl11hsU+sWNWuE01Ae7Bu0DmfdHLrD
f1E3muGtSt7nDadmqdSiwyIcNHIC70FOcFRgYc4JIDA3NgzeKdKPXcALRbW2AkKA
Z7IIAcwQfgf2llC62mc/K5y5sTyysMe6/MQ6EjNf3OhYT2pwVLirWCWyx1aN7IG0
w+x/Hpy+yI9l5yjJW58tXLei6sG30WnR1PDFFKK21VAUz4NNzzfWBGU/CzFYhEdu
S0h18rHjhjIeMj6mohOKDmoU+EkXM5ekQ4VrU+U2tgqwpKproUWNSckHUr9emP/h
2fYWqyOgmmuwisEjLpv4rf3hKSqjyDtpy95Y7r6fjrSnssAbf6LCZmlnzDxiKif0
JEsF3vI3cqpiLgZlu2cp6oEZAr7FJQkIgB9X1fP9sbal6uyo1M5MgjfIRLyXcY1e
tRGRuJeFbU4bk6DYGKkRQEgguS5wsx+dYObqxZfgN8obeqeV/8ru0tyO1ounR9E1
vziuYrOHcAJpLB8q03M/MgnbK65Nja3gCC1yOtA8duyfcN3wtm7QEFNmYiNJUvp/
Rt3yaKZ4Dov3Xw2vB6JnS2WAs9IxO2R0rJQHtYV8EZwgFUN2BFqs22nQ4BlqKKnt
QGDm0yU9EjG2d0FEk9J7qe2/eDouxaHD4/6u8X0lOx5riTKHTo5eac7nCMSjV794
EzzjTvPqG9ntn4L9Z0UKV5SvIIkeQtyGe8qlNlAMuXaPmZgdCR1RfawueCg0Wxss
MP8ZRQimyGaSZXJVqO4+rJSHOb6Rs9Ho8JHnzmN0Bhqkbph12q+zs3KrPJy73vz1
ZGy23I7ixvNSfmHaenpA4IxOGgfaeqUo9twlmurPzASNe3x8+GbzdVnpiNk7dUFK
8IwKiEHmfM0sQJLTayZ0nd+4A6LpCgvFupeUOLgigo6C7oT0a/D9/raPkASl32W4
s45WiebqKEWuX5wXEIBY2znNhJcey97pj0WtFHTccOCH7QzaCLxhEaneNwOEFrbd
nd04sycRjSjPQZr4m2GHHdQxm59+tHU25iGPBYABjfVj5r6yrpM9p0CdY8voXal+
eVoCXBPpO5sH9DAKHO/8mhLUOSHAnYs9nbgfMoK3W1LTFLRnkqRpgZ+ozbjQB8v5
4q0KdqD+v74tCGWgXBjRn2oC2KFQVulCh7tDq0tW1T6UIOIWclzkmYqHpYBp81b0
O0UC6Xgwdf+rL7sE7WDDiFiSV4l6w049bQ7G5shrjlX2IZxM9IkoIt0dqka1IhAE
kXLD1D5bseuZASREMQIFMBp1b1utX+uy3CDqRFKCqd2YnVKyLzZQe3Q4zjVUVIa1
VMj0ijRB98uU/Iwp8UD4AjcxJ1uXyuaKgHqxTufct5DsJzU9g+pErLFTis51KikM
uA2Y+pnat2jX/xpzrFBBGQVVSfgvia0KBFF433NffBhQNEqQqCkEzcJuiGjtGJ6c
OFsHHp70vJK62zJC98G0K4OrOtKaSaFqUq+6mX8+wE9e6beuBP6IITwwGhXd1J+8
jptzYEE4aCQqgW11DKOkVjvOyL888ynmodoEiiEBU1i9F/Sv8sBkZGOz43biRqvb
hE6LlBIr6CnKjRW2Gj5sbjENX6jspZwE//Dl9qvbXWUG1QSiG9kyC/3G1OhKLGxu
RszuZBBtNlXQUS8wiZhVM2MaMToLVPrQjcJVl74FRYBHR2GJtAzL0N517FKTkCuY
p8GPN2tMn1HgubK1b2KeOmsulcrpn+q1k6EVgtW1AGkO8fLEgvMa81f7YdfHMz+5
q4wEwRCYOHj07qOsE3OfKFC3JuCRnc3aTliX9SaDr2ML7ZgN2rZaF/RmI0ChBLJ2
7wmfWsLgUX5ejuFc4xVq7BtpxoF5kwhqjHQhYX4pbEdOwQ7gjOH0sMr0UFGPHpMa
P20+fIIqG6UhncDjB36l2iyoqhHMnYciJlas6shhB9g+jJS3mhCbPPboSdNpA04q
GmGy2VtkGwAeeDiNFBMcB7EyjmbJfs3T4QVJ8SDSLvO0xwhQt78TAy55uTe6dKHe
holGaJeYtEYm835dY4e5yHLH9dXo9TxvbawaNpNUUkYtBxMlyRBOyJdUeHgF2ESb
IiqRNonf4sS8eBeMQ1arrJBFZPikjgymeOIuolRHmcZMhPTWVFi/380cGIDfwcVd
qglWeZDPpFFFpYd8zBg6bQs68A8Ab4rt1BUM3XC8lRkKm5UZFXRomQd9QY+IMv3i
EqSXTzFHCHMSUtNWzmgfPOdsXPoKEZAmD9hx8cLmDPQiic/VXqgrP90gnLkJc5Nf
+dy/yCDV1QTLLWLWKf2A85qd4ELI2eGjYGpVipa7b0OaDHe32tSJEzD6otx8TSPP
tXE6nATrAzjbX/ugokaWeMReJyVsjyeis436MpIiFYH5l1hXE9Zk+VeWQrqCVBRX
BmwMP0K70eV/Pgcy4EaxghuwJRADTFdz3lae/UOlwwFVSf7ufbZ8iOlYA2AjN7qs
AwHuWGWkSs7f/R4PGb1+ZKOgepZJbHxDZSNOneuZGN2YPP8y4sme8fYeKVJXyz01
nKJ/anPNu5xVJpXGhPwKIoQZsH18mGmH9mD4+uBnekpGIN3Cur5NTvPxmkxv90ol
IJHub0hJG/tOdbS27ZGSp4toHFucLnGN82QlqbHegbmmHemWus6WmQViiivPtdZ4
bK2V3nzo5G8USEW2kLJ4Jkihclv9w6hV0GqB3WsEu2vm7j9R9XS39rmirDJYb6JQ
IXi2f0e7+L5+j2IHN04RM8Ka2exQ6p5Mfcb9XDZPBjcZo0xFov7P9N1UxEy1OvY1
XfGzDe5HN1X7L1pyt3muwCP+nGwTqU8gkd1O5KVoopHPd0Fl/QVx1b1IwA2Ga/hM
NdFyLH9v4XA5EJiM2BpgUU2Xcy+wwRnvKtpEVAqTGfTFM3Vp/1oLqO9D2ANseT5f
nazIadzo29QI1xMeQPqEuEJwXwHwtVwtrPHfv8Onxy15Ax30/NiAE8XVhkVPonBU
ivEnjMyv7T55NTwaJ747JoIp7dMQ/7foa/Jnpy6J1Nip4+KdIHt25OavmoxFFjKU
BPpGtbjULwe4tumraTBjvntvMqaXmIWkXA/wxGTtWKX2E6tsG8LeYqLABNLiMLgN
4nT3xa6rmfBEgmu2r6L8TexPT/P4ZNtTHKVUUd3Bw+ldbhl5p0IVojRZGhS2eu+Z
zQ2W/WwE6BoMMr7yQhZV2gAsk9HRV7jDiula2J0npIa9n4KOm35vxzpinYCLnYmI
RBi2EyeV4cFYMkBtsNhgEpT6FIE+Km87X8vl62bfnET94F0EnK4qdPYAkvRmibCv
gdSvgLPFWpRHxSHTx1aIxHQoXV2BvK6udU6guLMS25+2XXpUz6jMiCJ6DTrSaHZW
sNbaVDmDMJmWn0XpVoBLIxwcPVftMKLLYvQAIG/qR+CLrLBillRLG5epuFnzteU3
tUd4MMWZ11lXZx5Zo3Mi0ylnEQy+JxxE8aRwR4rYJfR6op63IfiT2JjXL3ZK290m
aEM09+hqUvhVMXwMb62hkD0OV+YfB4J0WlDITPXF0jw6TPtyuETuL5XPf0AhphoX
05UYsnEVWcXljB3CJx5zLRGE/A/vR8Z/hK95QqrC1nWXXLiro4QVvLRelztk3dP5
QzLAakAQketL7bSeRfnavRHem5HMvUSFItgqZFUYYDB4L4mf88RRUBrhPgu9SF6p
GsKhtUG4HkB2GV+EbxD1KOTbx7QVghsQLdkQWENlQ7P9RoixmlxneZ4ao/O2ikWb
v26Hk+20COMp6B8HdfeA7y5KwC/W+fFGDT2lh2BTpFAPEgNZ0HwXUpN9Qr/YRO1b
kItspMbxkV9lZqsX6k9Ps2tY8f0dsUf81vJ5XnNOsVwbn7JyCSC78+wsvqGMB0EC
wFjoPGLuq+7GSKXXYsWkWjd7nHThQFhryXK/6yqhh6zB8fWO910lqKHYXwOUnROA
WACzwu9/Hrr0xfE5CTLFPKWbrQrZW5ArCmRrv473DdDfvSV110h1JbuqkwGCaIMu
knISIAjTiXshe0R2FE/7RVzyS4RaPlEE4gKK49lGp9scqZS2880G9/bE3+r1yv1o
xo+J3YCVYGg+vuz36COKQ/5B07DvYou6bpmEERVeqpRbDtZVzZegIzpyJTzd75D8
a/4D9n9RcKvK2PmWr1MRYLwsggSTbpKLr6c7ckHSIxaqWgJJ3htleWLgX6r3Ytpa
gWZb89dGBK6iwau7qeCUOM0d4VvPZOFx2uDBRuLQzHcVG6YKRQn9vzRss4pW35tS
jRsicZ6JWDj1y3iSKZljrP8GrUU0OmvLms5jRO3wCA4sfPmGAod2cuDxNueby1RS
ttgAzGNZkARBoOPBUhduGgVzDLn8zKQwYK8G2vCtgok0DE6o6NFNuwnz+mz5HCew
2KnpmHAKwu1QVfhZREMCkBub3p+omDYIJX7I5wY0CzpsBqVeIelsep3xmbF1OSqU
ns42h8nS0sar5rxJiI6/jiQB2uArNHEJOs4AhayG7q2zzaja55ZL1BzwwlIrsLWR
WhfJayIhxXGrU1oyL2zyuAzidsVOv/BQNOrjA5d1z7P0eG3C4A+ixJLe5mlumI4e
oQlDhD4EujowpHM2HyJ8aU7pt3MmONZBI35ukdb4TAsAFFYTXdpZX7wxh7vI5WCt
gB1zl+TQywtaaO+sR0K/xafZ2XzIYxVJLfhz51DYwHm+9L+A+Jbr/mKD1CqYszhL
uWI2TqDsndKiOS/Hl3G7W+Od/Hf1Rnx5yF3q7lUyHOizdHiK9L/Ltl5YETd8zsZR
uWzbHklkVZwCoFCAjfYALrhs71wzeJ2Ytez9WwTh9TBnREPRKbQh00zc4nueCbwM
KJ4WGSryaHOf2IdkOml+i1tQotvvXI4XvwELsCRQ/KpSwX1tKQqtWNTjjcbziLhx
4oX2uBAchlmfylD2pw455CnP9YLcQJ8WhP2o/z6dcAKGRrLQysO6ArRKlnpF6kvA
MQseyVKLaJDzBaw+pSISULyuT6ql6QV3Fg5OD/LsHgDFt0eodz6bOplSCpWAtmqu
ve4deFQiv79GvcIQ1uc/MuWi+g0QgGGJswzWjt02HBwBqaSJRd+8puKO8OuJGy+x
o165Sd0x3XBLUK4To/+vtJLIzamGvvuvARiU6ARAjNo4L8tBJ5InxBvN5RXvhAJq
ywdU9AxIwNYtcnF8caDfiCS5qLZvsIPiBbu+9o98n4EfhTMBfBNEXsFqTMKreUUp
HqWWXV1TeCKgr6SfdjxRiOOy7fDk+jRCQfwAVB4g1ZYu2ycF764cDyZfOUVdZ5KA
GAqBMbqbFCB6aEEBqT/Rs6dYK85Uj1/WbAZSfdnHQTUQVGM3a5OZEcI3KoWb9EyM
pk4Dnnz2N9eBPj96WpfEk9Vq4tvdg1iQ6RLCUwpNDK9uRp+Q95/CReWXbuRrudVx
de+DLvsJ5na37ohkCatdc5MdNAckZxoywJIDbvNTLd5T04ITWjeC0oqcppgFCGek
prUiBS94QTsscRNU+1+W1fPT7f+YFiBClPDC3qI+fMZ5HroLsc1m2yQSbhWZPitQ
EsHvLDnLqm0+rjCO/fCgcBlf7gOmNsb87h3aod+1eZcY0IMolR1gm5OO3P0LcZO8
/QD/GG39B4quOMHIILj1yiZ6+gRPkorzDdEv/1sVF+R50WU054rBnzITSjNlzceS
p0yc0gCo8hXZoHCM1jhsAKYxrZKCFYEk63lsXpVU11PWXFZdAq4PesFh1cmMAE48
dal7VE30ed73kcYbCye88tZt1gRvIN7PEyc79HT7j/+vPVcIlOCU/94HkyyJPlQ1
5zmzDf8lRu5ck3Z48XSMONqLMW81jj0QEhzV6owSufVpffZpRkTYO4Aa6R0JkdeQ
skRgHMFoDySMvyO3t8ty97ysGt/G/qn8qJvOHp93VXpTvRRuMPyrwS2ot3wrv5lr
2XB+cbiQLeLKyx7TNIKvp9HNsL51vbJ8NRm4FFl4McKXUv7H9wdtxywjbi7WlvNB
EnmYbQiIRr4boeDK0dHa98PPvEJVgp0qPSh39vmLEChal3H+9RRuPV1A0TFiwgKa
A0mkbhXRlCj5o5jDZDoihxmtroRhKhpQ7WOt6ZNo2A7g9zUaNTskdzI4PMvbntcH
crgh0CAC9aPolV8Kg2HLbnO5wX5oz9Cxi/osIMvIO7UEmad5vnpFXjo6xC3mmarv
PIZ9AYJjp2PRG+WsIi0BN/OcyumEk1kF9Cg2BsH+gm+IvJjCLyhLPgqjFHiUhzly
KhippWt6DRtinK7FaTtHWzHs219+6N5U2e/T7HRnT3QN/AjKNQJuLPTZnLLxWd6d
97DSVq/j5/DFUhDX7cvaf6Zi7un06+BanuxduYsK0GOs6wBcbfnOibrPbAdvZ48t
M90YJpOg9ILXeLQbcliGY2MyE/frF5zHSEUQ0PaApkB/p95QSjxatAUJxx7oVlu+
lYHXxVyx3UDcd/Q4lmvzFL3q+4NJhuTNZF1so8mldhymVFPtRW4OQjs5YQTDPtFE
KxLFI4S/JwiknhvUrF45tL/mWN6Olh9Bp0GruCWy57zT977KwWv8hdJSivtxYQvt
2JFRI7FUjvCsdOt+RIDBRiTUh4F6/2MCiopNl7hvvfQItNbuyK5ooh2vHNpWloRA
H2baF6jexsYPzIEwS6DVBpDvJGkoDjccKaX8yUQiLfBnSld5QUShGKWYRdxq65Ja
f+JMP1Dwqdzq6tWkn2IerQb0KSfi9QYt5nVwdMDwaoqo3eJWsCyOQQEAKCS8ChX+
3NMXRjEeyZJHmKj2rewxDVqkFMkWYDDI4w96BOQtwV+h8CXa1KiT8XLoFVr2mIrX
1t+/f9mfdCdWJe2FH332I1+NAfCEN+nDWnRp5ibU2UvxsKI1tjOVoysX7n2Sw82q
X7RPJ/6MtzFKqEZHnhNjwP+2IPGAwL8zTftbmZb2I0no/OaE4CH318SjXLC6vt5F
qRFshyjE0xwh7oHUPwUhozd6s0fVatMrBSkx6eXM9AmmSrnqfXYWEWtsDJwlalUD
M1S/jM7RiU06XOO16TCy8L7jHf7UxF3U5N4CPwYePgITu6/2RS6fKb+Hq+OCk4UB
EnhapC5lSNpQqAo+f6MKxIY31Vidtjb6s9sOR/ZVQhSnUl8ttBg+WdAlnitHgBXn
oYhx7a2E5/3gBsuqm8ViSwc25t+ZrN+FeZxWmQJDzFSknJPuq35tP4rn77bsJ/Wv
Xuu5bL1NVHmm75pqs6fJiI6cUFPnu4ye4fdxliueEAjOtWDceRTv6fv5ZCj6DnC8
IR00p3WqkGG5D0ONp4MuTCWFRp3O5/FEeE6NqAwO3O6wZvLE+pHYotdbzImw9mDQ
LG92LEiVyIMee8tERrJwFFKXhbmvF0LjrGET24VXcI/zJ40QzpK+4XTdk5QjOfOu
q95X43BO3eGWTohnUMVlxL3HwYIErOalmBuf5FpqBDeZ9OvdPYKjxmrztRxDZzBH
C7O3xaCLt2tomAaZC60qyz2NhC3jj4ZWYt7ncwOgBDwJSLwyl7qlLWYmcsq7nzP/
sU9XT/ackxYE4ReMR2aYR8Uej9/rcib8SQ87ZGUsy/c7DjtZ/CXFj96zvKUVOHQh
gJUan7hI88EYD19p8+S/QLBS2GGWA3CXnDRnS45AIOOEjc0tXaYZ+j+ZOcUvVTzT
iH0Kf1okO5DOc3CTqQNR5xnuwdQQmXUDs+i/NOgSvOl18Z9El2BcWxty9zj9gNjD
Hmzd08O7iTJzHK/HEDoC3tIxsnvam/yuHkYR1onFoaMrtT9KGHwVlzSOvoBEXmOa
n0FNfDmAMyH2R6WMpqPJQI7ofqihJ+yk7iLtyT6oAjDX0sC2aleU58Y3doxGb0fC
skXBm9j9W5XY8WuzsCoubrwOK75ksnkehC3TVlMg3HuqkLPFY/1dP/NzUKuExH/D
AQRz7Drdma7zkzcz1PTEwqXUy2gcUUh+SQeVqXP9XbXg5t9wGMcl0YsO7o78+BeN
J1agn+lAknvwDubwyrsrAF9dO+AIz9N55rl9ziQ7MyozT1SWlxMbH4nLItvD4XRT
1nmY7sPBfw97oazN2Wt003CTOxRS5Zf2UVmBGK3JOd+Ik642z2dhgQp2G9t/gAuA
z3lVuqRkAGNXCQUfA6/vx97fBAQ3E9KHRGCFQtM4vrIgbqQIyijsX2GLt6/7m194
RoGpi7iS1ujSmvUXVLO+jsiSNHfBKsAEvcrZKAGpljS4Sk0VLhZZqUAmuaG+9Epo
SDB3SOhuTpT055ywlMutrrqvuVedjNmwzO0r5fHZpyjft8v8Md+0XYSsk4bOGMsY
795mu+HLJzcxrDzGU697VZ0QxK5VQahKXZwOeNT8TtBJIi6VvZh2HupxRNJp2kmZ
tGo3uhurI1PUKaLauAXiNUkkUYx1laedQEuePClA63Vn9lfRoWRsVPyo4HC6Z8bf
ccMVTxeqeoNGhrMToKnlt/ys0b5TgJK26ITidsQj6t3sc3M9Kuty6V46RRQvNjJ7
yAInNsfoCG4EmkH5+mqZrZrkuuklEA5MpiTzRhWoFiIbC6qfyFQmaYMSQgRzejK7
nLSUQaDanxWdK/Qy5RQejjRqs/p4e29eWb+JRdLeT0h1SiQHE6C4UHg7IAhPHACI
rrvyVGyBNIuGcWgk3MtixcrEC92qNJTbD32+TlcDOevttxfxMzD6VoT1GP55fDkI
3UiaftTJ2ABfgXO8m54lMyaFIUPHj0xAegxoBGoz9iVdRkHuhUNqOxMsHlcU3iz7
9CH2CrHbl2ue4X/uzwGqT2fRRkGP230/oBuObsgOcAEEM2OhKlrvjriJbieufbHN
0+n7q5mqR3vYwUmHk6n20R0pnfapz8jI0kUYeJRD76aet+Qu5A52gIbhNYoeG70k
J8B7IpF3tUUEgUm8qmcO7kRqf4vcWZ289llDUJjKImq2EwdcFZjhVGbbo6byM6Nb
wPB5Fk5U2moY63+E/6Gffu+IcuCMdnrx9A9ViIQVYxU+eHoW50dF3By5Yz9J1q2Q
UGdlKLZuoweOP2pQkstVKEkVXIBuyuFYtw57jDtoU//MvpmWdmCF+mq4avlHgQv3
uErcmZlPx/S1No2aRBbLnyFlct2wZ0UdAwJwA6uROVEMmHKb7qG0atcAjrQ0M6h+
fLQ6TqRC9O5mpIeHWW2UcYiAF93BOjB16w+DWrcKdRjVabRgmnjNdPyXZZ/nF3E5
Avl81goaPHiUNjbxP9FrEZQSl4kNpydLmUv2Id3pcLiKdZVaw7rP+gKCMBF33NVC
jNMlX/ASkDDqnKrIjWFKOd636dxTqumJ3FjlxRwPxdQ6RuH3gFJIPS/pXO9AYQ1h
WXjNSjYge5JqjFYy+KRAGsWQ5dl32rZyKYg1wBYOQKd7zQVZHFUa1jUFY5iLBsyr
ZeiqJ+Knze3VLKB6kM9hR7qB80Q5F6LcBW4InAaIl2GAx+EozmrnfyiG9/UUNATO
PPBdS8G33ivuhT5DzchUtMs/cVdh4CqAJzGJrxIPpPTEXgwciVVFM8fDEKSFvDlu
Q/OZG189evYROIe5hanaJ98i69LAPNWXFJnZE7BsIV5k01X7A9bCRDvzgd5hExHZ
v4okz1S0izoEZKf2fthH3lbufc0KUYG8zI645ho7mmOEJcaCPwwp/Mtq/cMe4Xf4
0l7hiemX5LDLOZuIeHhnbOQmnZlP7G9Lm1/fyVZxUihZX5oq8hkWEDrcouHLk4Eh
h3L0//T2rDwwWVl+QmARneJ0qens/p9YzZnwNM6Dn1bejdIdAZeZtP2dX8mT1xoP
+bBgR3I9XmLhD0mBmvoi9F0VIz7V8IhUpEDBnGrJAp+KJXpp803dEtBXNdDrWINi
zhmJjUHRB6TXesGPtB2MSmk/acpqFdCmwtRI6Te4vvyJs+WZZ+V5NRNEMD7Iu3qB
56jDocklsXiLzuKHbm1PTFMz3kvSvR/6CuAQncy3udR+Ca+XD4Rv54XSNARwFafb
yJoLpB2dvVRXru3j80PBaSom81OCGJkunlCtP3XvMQROGCJgav8K1/0lncmE4p9o
c9MP6kSK0YX6jBvQ3aMqUdfdZfPtIF5KVZ14gbj/8FDtD3Pv9qOc0krPw5LiSBh9
0XKBVt113C3Zx4SH5D0hNwg1HVcusAUNBmjRMSmgA4E+NqOPQaj5OCINCe+yJ8eM
Kq+rzi002IuqzPEPWkEFmaWKmwEAaJ0KGoZOhA+sqIOszC4p+TCUQNqG10WzWOGZ
9avlSA+BRY4TkRkRtgdAtPHTAlC55oX+vhrWYoUCJLxxT/mBXQ7F8SNbBFq5S9YS
1UnIa+NJiw8wehsMEd32IIaMmo8ZCwD2HEwLF5EV+Wj5Pl6uX/DnOYJZcJEdCOnr
QLsxM/dmUMDe1l068Ur+ApJGFWHnVm/dk6ehuaBMnM37h9Gl1RPOFwfDI1LpuKiw
KiL+UanPs6JjgHO7vRQVV2PCM+dh6wq7grFnUEsWHmJaz83den8qTy0LFD6SDh4v
K+xaWq5Cuc+cZKKJC8JDsKpcxdy6QewB7bFYdH95zM1l7unNtkMMluNoBKWBTfDF
CalmMjmxqhikvSkSiBnOu5FrNSS6z0sClMyoNOUOeTxA48VvRLFIV+SSWn4xUs+P
TczzbS5OWhiz4uu9hlpJX88eY0/GlBuC8n2I8b0hNlsNZ7sKMzhE+JOjBi9YgQyL
Omor2GjhKmfgerO1tyi7aPiA2wNU8ygaMkVQv9+FSVa5bVCJUCjHMGjWrjxx0yV5
xtgPWVaaLqVug1a+bqFSEFp9qoybK9ebkINuqph8KKz1eOmtXaXa+ozO7Vn9bY/j
dgXrtCw+HoTg0CuD0ZA6FXad1FCjJnyZPvRA2Crz2OuiXnFuwOQT5hxlBPeIcYVs
F5Stp0zeLsQlzOr4GwFsPXpjmAWlpysKLox3ZuI7rYtMPrWLakHn9NbbXLDZqMce
IX7ZSbqBrDV1pDNb+mABzMgqoLWv7wcOoF/8aQ86OE3wSJOI0bmVgTsRCH+ZwrS5
joMfnUkmxjCh6biSZv/zSD/otC25rafV2gai3mJXqOnGuOk9PtGiG8hOv9C++4aB
C/OZGWbpwnRS3SI03fNbt6I2+GjasKszZCrf3Z4UtS26MgJjx17sEbk/83Q5D9KM
lcZz1nqhZq2IrXOPFGMAw9TTzeXDkhut/zut5fbVifIUz3owH9Godmw+MK7UdGXq
zca4CPzApXGQsj/E+Dyy4MU9Zly05bmyr+9ZbtdF4ZIvvNTl4sfFjcBBlhGK/E5+
5w9Tmk1z5vUop22di0SjBdewBbIDgcBnsFospDrqirUlZV6GIFp+/fT0DN7O8Tvc
/6fPCcrH4aWXBkl8KsZiOZ3gzmSMOtHVYgRNeNjJApXKUojPG6vt3PWV88N80H42
OZeEpvy2FcULxkn9cXF8fzQEpVmnjfnbg7rh39Ef788KkFO4sYcuPU63miPV7gEH
2HaNOoRanKaBygRgOu1WNJHHuWSRYZN9yVOBEwH8OfW+u7LDeBiiDHTI1zNkeoae
nSSZSavRDapvKsCFdVPBIfK+3d6qtQaLTXvjea//mYZGst8E8aokGj5DdwRNFnuY
N+FPiB8R+Oz/HZ4dCcp+MLHD0oJNriBuzQzfy8ahJAU7MTF2YHZ5sCkv1+3KLzNp
vW4J5ZGjs4XC7fqW6t4aJMK3OoL6sg5JUzG4/RkmfoopmM+Kv5G2yA/zlMt3yeop
X8GnstmRunPEd1eFwhkN4prpCgWwvipzVZEAay1aXaQrMvwtPzLxfpfmUTgmX7+B
92yVTKXUBv750REL72uyQuX+Soo3lXTS6LjfVbxr9YySgHHJtM9meEseCwipywPR
NTVE2mXA6GDlJvOSAA4KenpAxhqVJ4FUXaDtW6GqirFGxDncAJZyLQjRipAquxjR
jyakTZJQKVgINKUQnpKbMXgvWoa3QrkBlrewf7dbAb0V2wUVXkamEwDRpKoMvmtT
IBRCYRPoCdeVZ1wJRCRaM/GC3gnIbLfXDKzE0PQ8Vdb1HgWbbHDQ6pPUTuVnhL6Y
0OB7szooS8g7liL0wsXH1ffRw6z7j+1gJXj6wjSOXEClTbB+TDEV8dypw8bfLLwx
vuUZ8r8bwDd2QQ+W9EgvFK7CaMRvI3VQTjNR/6Mkb4izOkrpZd5eHVYlo7F9fpJB
dg430drhG0n0pfw0VFaTxet8XBaAZDgtwGSfEGHel8WoVF44tolr0du/CdJL7+n3
BD/CcN/CnXDUc1PjpqmGLvyzFPRr1oud5jnREMBCznvEf1EaY5p5KpSPl2dzUmiE
3DoW9tWsI3F2iARc0RxOnquW62pkkqQdWqy2YWOnclwj56HvJiSjXHXR/MgnNNON
je6xf2u5+UGKSy7zG3/wJrWlieK1H8NNBe+ybeMpG14Aw29FB1SvHBFRdqUL8Vyu
/aSWqbQgQAcxK3wWyeiltXe9IlJaBqDAIq5HHJdoCE+7XNcIa06pa8arjilArQ5y
l4Sowc37NyQVbfB+Ooy0OhqQR2IqLLD8MxH4oi2r8rafCsLDInMHf9FBOWmTK5+y
UjHKVA+uDOmBVgJw3mS8scZ/wOFhBy/X6/xeM0x9JlfMoUcAEPGayn7PlULC0cqY
ntzc8I1JGximevvXt+8/p8eR58erpsCo0CviUFsffe/IqHJdXQwCocJ+rejkZ4aa
IDH3Z/U10FDNWDzIkUxLH0djaiE0+wwLtANfyNjfk98MzKl8VncV+fk1psn/IRQU
Y60k6rq/KxAO3B0mOKpHlPeWnWA7GeOvJMx1iI074JyfmzdS0e57cQ2jy/ArimRY
AuBgWoLSgvLtL5Ctrh4wM0eaZeiCOCmMndCo6llYJ2Xpt3og6lmYkCOOOCZgBFju
ACKKhmAPpIekpebuLneI8r9mKFfAjLKCq+sQpRjTsb71TTKDmBpjQmUgrVhKmkHf
ZXFykap8fH69l58USDAThR03FtO1Glhy7UV7LWT7gUoPOF1rHFJobqHzcJ0JluaM
pPMJNqWD7qTLsT06zQfUJTK7/6slticJE6dJIBPRieV0+tS59KPRduVdGnqvvxHX
7JZVDnw5wfPfe8kmXhaIVcXqtMQ9RjBHd23FEbzzMAZ50Pg6VVyz96M6nlawdUWB
wBUnKnW8v5WBWnwSYqi1aMjIrSM2BzQSrf3Eh5THGxsOZJ5aiSaPADejfLM8xDz7
WJ6UTsirDTDZbUgy3OJ3Pa8BJVXBWeCKvgKdeFzjuBfRfjx2KlSCq4OdLFj3TFII
ifxfUZC/UCyzuCxDpoCNo4r1nw1Q2dQhOXMdX9m9/+8vpIaYnTGFT7s7rJNnvjb6
7mjUbIIY5mMMzLNwPWsNtBI8D0Ze7gTSKo7h4f6uYm0TtsgLLkNkAeTkbiYuSGrQ
V2muN3EXlBx/txHqEo98jRwz7G5o3Tw4bspJyDrlp1Rn8nNE95+cw/Qjsy5xCi+5
p4dC1QEyOIOoCkqKv7zEoun9n9d4p6GHIQiawxn9vDfjKWTvBT3UEq5tmy62EJPH
8zjYS8t7qiU3U2ybhnN++ZQbDSYeZ4tdo1ORSoOlj15AnSooTRAxATa53lHnbc1i
XTKBDQ3PjWXc30Le1nd3vQZtwtRpEHu15zC6Q5njOY4XD/1PG8+bcffSszm0IK3w
5M3LLdP6IvhCp5+wzR4bDEJrtw/65pri86eYlhxLXjLbgkn/o4easOJSTDw9G+Qe
EWzwdbTA4HvihxbpJaVv9uvKW2Lrs49EpuVzKUTmonQb9GNeRygj5thUCFmj2Nk2
oBMsPpxZMc0O4M3f/7awlTMPzWu1woAYe7kAMVMwScQt3kndAsb54skO5gOKPxBC
U7Rzdp4w/O7Ek/Tv9PXi56mxTWkY5ven8dEbZwqKGLyH16SqPM3r7QH3ZbfZuy7b
f1t2yr4FvTle8w4VNxtJhSX3kNQoCReV9LnFLy01Kyc57LFZAGuP/vn4erF7b+tN
xSk8122BOERjhHfKvqa1gspZ6vOqJ8ynsFlpHrhDiQX4b7PpdIIOS607u19UO3qv
lae3S1M/wgqgU/6MIbzWtPLJRSr1ZWJlMdiBUbPUVLxkk8z+qa1IkA6VToSdZaBU
MxhIqtQ9EfOQKV6XhPj6ffu8T9X5m809Auq7Hi3g5ay2YxeTmb2kf9nlnAqU6b20
1hYIzAT6/Mq2++C/YtAQMeutjn0Evf0T5fONzrldOZPs6Dgb7pB73Wq7G4uqd/3W
XnvuXYcC4c1mcuJtW9prnTG83oq39N2kxnUPBACKURZGjjMRsSuL5OELoqRiMY0J
RI/gQoCtPBWRZogLBNBEuzOxP+ropbw2Es9mQMEwxAGoRgzNKP9tNOriwODIOgcR
Fpz08s8BjXMGmtpUn9Eh6TSMkjWqprjKhZ+8D09ws6vn4nRCicR36IShMmsv9X3b
/kgECDpP+tsiqEnM93JKrP7gCSxBnTcNEktymBrALiNfWKZgiEVdLAHozpmRUbfE
4IqEyUpL3IG8tRnZDL7cRx/dg9E6fq5naeSWhlCocllm2WWsTQndvVGxXtQkix2J
wLQ7chzIwD7rDiBH0GA6Ks3mSL3oKm+oXlVDt+ysbrWG/7+BEk4LlbnDSQ+DPO3s
UqGyzq/l9rQBQBP2NuCrtmPquvVKt5EM0BkioP3Zf6TAxkGRD66hjpXzy8dhQ5FA
mnPbdLVntiUctCffuds8R4Pmr/PcRmlQvkM9bEO7yFdYJI21l0W+oFOGi62h/14S
whZxLEMT0vmMM56KGRZG3QT1UZpoDSeZK1MBDx0LKCsGOvIWc4Pltxeab4ut5Opr
zt9SGxME2vuxhWuHoe4Kwzd4v4EvqWxq8630qBys4QbSyrK2RoGfrlweiqknSa3u
suMzouZWbtztykoYN+S3eEGEueZ579S1C2sp78bZbjkfmsU3a7aD4SSJ90ymwtMW
X/T5bRkfk8wn9QctXfytbsJoJ/KlRr46I+z88HEfJ7n+9Gi8I/Cfa7UWTBmUGrFK
u7tJd3lhgOW0NNoJHd7cKgsukYLGta0YBs/LxIOQEGydvYqQrtaTNWvg5joz4LIe
fjTcsSQmoITD+k7ZTgFR+3TcCVbkLIH2yp/L9vhdC95Yy3PixUYHccPiYM096iM/
cn68tiSWMfwghrFIZtCw6BvKVfRly8UjlOvLKZt2MtAnkpnPrac9Hr3zFRpn+Z9J
VSxCq2U/mfCCAB1ryPJkP3Ii0r7EgtW3kXOy9QDuQ/Rw4OLy0/F+Kfy7At4u2L6C
SbdDtHeqiohgmE8WXakhDSdMlLKYTPIbGEvu7X0KH6AECe3K1tE1JKswormvug3r
FPfNC5M2w3b3QhRh8sZxXTGxhEvMQPCsTD28CtSxHT31r9P/3K0BN5fxkiKFkXSe
yC9KvNhTjO3kwLoqy74eCIx4ZRl5lKxeaAoC8dXtZyEWR5D9CSAGEkx2l6Pwe1Aj
13rPh3PI7xMnonGaIQUvu+rO5WCn3/MQOUBTijbF6Qm+CgcNVuiIoRkHk0l848ln
SvKpqw2cYZ1+Jngscx4i9vC/P6viOBiaw72QfPveVXlwuuQxwjUZS63X+C0tyrZd
OpOIFFt/h0GCPPw0+CdunxkxSYAcVQ9PV7Id5QYtN/DNwtUgC4Kwl7X7MCcXycLZ
0eHwWgBrZLyOs7w+gDEQeHYnQiBAUdsE23//ynPWLZq8OlrugVbQskFBv1UnkTjx
NqORFe6nGjJqUgTZVBHH5buzqaaqwZo2QLggRHSv8i6Ojmof4CN3HTpSySTMCS4N
8kWou+1IrPa6zQw8jRh86IWM9Jl8x8tu+VsYBcGuak0gNx8nXrN/LGijDYFiYHQn
y/0GEmweb2JLj06BEy1vobVFC8T+FvsrWkRE3ch2kxMA6KzDQmA14EmGZ6XqzfjC
FtsNO1xs4ARF49di+XaXGmPOi6+WeR4GwUvM1CJ7Hd9bzQuOHbyxNlLaq22jnPiH
RT5PetqmxL7IL/4pzZRSuHohxBz3csYYqolla2RybZS4AYo7yfszRNlwWEtsIy6z
wfhluakrxyopPr3rmOtGluubcEXCPFHGJdY3IgF3jz6gaQM8LBcRiYy/kC9itCoS
oVkfhntGm1OG5DDbL79elAFTHHOZv0Q+W7PzeMW5l3Fzpe4Wu4ITzhoE0lQpw2ur
3mbiqgS4f5gxnf9xwnEkE7bE/315pnuNEi3oRSwq/CsiTD/mmLhnD0qJ+9nMW9fu
a2muFLksKcBTOA3UeqhXbkQT8dw0H3gT9OnixABR2y02tOIPfXwlrOZmneHqCgin
FjGAvMsNpWGxS6Z6naPFEBCitH3A88CU7IEwdr+sfuhyK+URbZffoPv2F379Swzx
rCTtllnvG2brLDGsc3YAd4RYmDy1sMGWJDIW8U59tcoYNEJXlk78BuN/D+vKWada
RfKjgiquMEZSo/b5fZ7Q3ukXB4hnt1B4zmfn2/Klss1/I7pnm7i5CkkPpfr6TbCD
8FMNKq4/WHhX4M+L8N/ULch9yGgBrcsBlw14rSyeqMWD77zHbw3ep66+tp4VnUzm
jB/LtZg6U7E1mBjSZTR3LGARSDvjwRX/cByVhS+5K9cw0odH+HtC5AWS0h+i4DM0
kpGp+CDfEOFnfBRBGReQOarQpS6cTqUL2bvRLked7tBDNWxOy8jIpVMz3fIIhSqI
+K+IA9geXBlcUU7hoO2+OTFEEKsM1OsoTV0SKPACDMahMTmYdzW51oEFUwCeETne
JsaEg0GM7AUPuy9o4AfNaUyPJu4+kLXHhG5qQb1hHtqjGC0+SFBeOaLpvK/OpYlf
lJF5OYdXljaPstGiKOrbECOVGXt56izm01okD2PYml6aO9+EJo7boUxD/bh6/6O8
pEGrihE6DSD0u06MzPauIJbQT38NUmMlJruYPz5ZgfuitwOQDTlP44GXiH3Uw1YV
Xmv7PvAUdWXedmTfmULlTR9mXBuhxPJ6IsJpDObQ+kWtf61r1dH7x/13/88ROzGA
DwteEMUkfoznekcbTOSqWds1+RNoBamm0OI6k8DYl6hqsAmAM8dA3k7aWKMG/WsD
2og5Fsob19/bhaE4op3g4Kc5hWOkIj9W4wYB7nxc6US4VkWOphpyn2fizxYYI5uD
PIyyZt+Rw4Wb77eurgLnTdVdZ/Ay049OHvYi+VogY4g0tcrJ4KlLCpmwtLifdEie
V/9eIhusJ24GHi1hv1Hbi3JB61usUrEeaG9+1me+qiaqt5EZm7vAmFdpDou8iY6z
1wufgiyFe3YPBeisdCpAJtFhwkYYFd7QEWyuG+OiA6SFqzqq2u7jbXa53NLvnuK0
j/ITkyz0v0gtawFeC6qklMXoENY4iR8qu6cHTYSPWi662315R3axU//agLoWXPTT
x1gQojORcwjehVEF9CadcXG1wCJndJFdnNpO4NHtWarbPWCeXvPBikBM9cpS6OdC
YkktS+1L0xky2Z8gnk+smJbFYY9oY7TL0kUrHVk647sPfA+JoQ4q1jK3dSuQ3F94
VfNd9nWoTUUlW4aUH/Oh+0vrUQo+dlLDcrywF0KUQY/O5D28Av0WMAHywYqLs9BB
ipXKBq0lnAUFhiHodQK+j1JlbtvEZ/Cb8Pt8tpujuDkwStoG2SsLnk7/TfgX4XUZ
92XQmltIqHUh+EdhILkiNvcj7o/F9TsziREFCPkQBqVlwNi6KBiO4QMUKcsNdf54
i3hTFq6VN+/DGF9TzW19mHn2wrDxOrCqKm0S5LhIAyu5G5pePaNqC/kUx2jj6iv3
k4TtV5J8U1/xJRvs4hKd8mWalbq3SwuY25MbXIy2razgtOI197D/kmiBJCk6i9qK
yhNVt5bRnPBo2rFmahLRF+fHuGir69EmkRVXmvkjUGfVNm6+Jq/eI2eyUSmrPDjR
oDd/UxTBzG57DYln8Mg+xqVTJlxxXHvZWKAINhMp92Bf0R5hTGDNCOw0BatfUCJa
6TZxcEgINlrTJfCH9mJ23o6KZ2qrCbo3T3E6+HnrmtZl4o+xSKbk6jSrEWi3tC7Y
KlptSG6rPIyIZKKC5SEovmzG3tcWfgTZjPjIf2nwqcKDsBtB83fO3F3iSctyqgs5
+rzmxm4J/de3EyssV1upurv93bitcJTTbKWfEyQLIYSNT/WHW7gGKSdQ9VZkM51Q
Trj7pCXyRJ9DIIHhRSWnf1eDw/U1+pMpRAAWTK4A+BO77SiOWFc6oS4dQPDv9+5B
06sYDxvqDbpAn7gATReO/r+goL1Dz7M5RFwZQhfeT4NVBxiTG8VTXCpFbdmHTKSZ
0qAfGcAjgwXHE56qde2fqMJtrBkb0ZXWtx/P4GaKrHvCG26SypdficqAAXDaElf6
lFQJXqE7ON1Yyww5E+d/p79Lo3f34gFbbITWeXc2aJVZzgTAgKgL201/HbWJEN7R
Je8m92WzdtN1NCiu6nTmfmPlH9IL5U48wj6BURxQNSqiVRYZ1tb64sTvGUwmM6Az
vkKuuryrVuIKr9uBT+hlbYs0GzrgCRDvWzHPc4pn8YpjBff+pNc8mNYMP9LkytmU
BnfqgHY2rSU7Dr2t3Cd8N7fF7d0EEEN3io34SDSUVwhsAu24Nkp3PumWj4cHLfEW
UCIrC8lEVzZ8/bJMjp77uHzAYFbBw1NjQEm8/KO+w355gOVxOR2hFjbDzgeVRKZL
41TQL4fXP/Fm7L+rZJa8bLvkacw2Nh51wCHWuOb+dnVcY1sj96jpxjyba95PHyE5
S0ghKqt7vjF0TiHqAb+6BF0NoB/Ikz73uoyZhmd+DtxgR/S2S+nXv/GyQaF3ERAl
3QwV+RRDt3Oihx1BNkeSGvZvFFngJeRuViM0B2l4QdJCZBmR03zzRtKSdCtzXosY
Qlh6GBrlyZPa8g81sQc+KjiU5h2Gns2AAnVMEq9vY4izCyBy8oYTqB8ahjGfyilf
NbuZ+hup8SiEnN9gSAT10F0utfWdgfqkV0O7m4NIpDFszVSFA/Z5LUUSDrLQYeJT
Yc5Yho6gpTUut9wwdFtKstC38tFZbb+fBaf+lq/gNJgqY7Y7GrOw83oKxlslbgnh
Rl//XYWXzEGcTA7h9K2ZL/vP7yf5cSMxO4ryq+Rqn0OcMNkK+rkaU/W1FN3fopbV
Gib2+4+8gr6dfNKSuBlr7fWiDveqM72/ivQbYIdAE8yhMqJJQ7VhP3WTi74rVgME
Kmzo5HNP7z785Ppg4TiqOa7//YreeK42ZqXHpwr/fzUJ1zRTFTS+eks2jMAm82DA
7W65Vvjn1gXOcIK6Zobp6ai4QQPAqJZFa3eZpKv63ZpI4MyRdDajDPpVvoNiZih9
mOXD3LyKYAa4LliHI0ztrZ8dLYDlguD2BcgiB3Bw+URllVtoS+Q7WeOXWfNPfCf4
Dg4uZ0W2lKrhKpWUh7wVmHJEGMr+rLKDzrJ8stDbajw6Ar7/PujT1AI5GDT3BKu7
wfMlzwp9eqsBtC8nCT8rocCRZiVpABkwwrTZqfzSDYniRxt2s1O8/ifkqb82DLDs
lmKOCPUbrPWiwpxNQHcWloVft4bMXMSHrP3KVzQOpDWS/xSHNZnfNJ2WUu+XqkU4
4ik8R71yT4i3NGiVmF8dyVuR6bZCkjCChlf699NEYkZhmeGTcilqDU/s86VvHyT8
eev6TSZYn7EXybbBHRfUqiuUvXFFryDK6s+0PSJjjo5Por2aedFsEUs4vxobcWS/
1/x3g2JAhaxpkQIAcEjsWW/g5rsN3oOTdjcp+Re7fpwFCD60t3tk7btEMMevUV6o
aD3FsRYA+H3+nFuVZq0eDaWjdHUgBgYSwSbGvpomIFGzwhGiB4Y2H0gcuCKR/fdO
5+DMSfslQJQscJaZFrHnU0+0v1J6bdqC2nAwpionMkLJ7eZhQmOM8ohU20G7q+bo
ePKy5FgEnkOjdQksucuoRYojxVeFvskVuSBJ+dOePui1Pp3hEkS4gFZ3FM45Zy0G
Z58QzEJK9W9/cDJt/T/gRSbvCIjXeqfLYc45JphBd1LW1nnVF55v4AuJ7z0X1Paz
md1+K7dKheb/Ocb7hdg4pj/I0xC7HyqSbTAz7r//2TTb7hZb4IYfeomL920ljboc
Cj60Ry/xltYxsBythTXIEblhmG27/o2YskdDkOKXycgAzlVvzriFmRVsWVvi+VA9
Mi5ZwMGRum2Zny3a6X6aWdbcC4Ip/n/sLy2W3jKBpUMHW71fSMjn39L+qb3YfkLx
E9Dhwq5swyuwxjfRaXmxuggaajc8RFmkcRXYukGVt4fcr2WhMTtjUkT6nbo76ECp
YhDDFwUUkgAGMR6Wd5qkNaKAODpVlLkJQCn7qa25rxCfVg4bKDAKVrBFkXX8zVMJ
wMiOMX7DEY0Gy3IrBe6H1qH81mGgem+SUPGEEisOMzF8bCYl17e1qBmC0B/xphgM
4kEboa/WYa/y6fvDwk3ktYQeloNLpXuH9T4j3VrGKK8qpJYqnVlY19LROW1nB0JQ
TSwqruaW3Atq/awcd5DeAax6m+1FkX3HMTrbqhmltvmNVqc51kp4T7jGWsTGo0lL
StvR1XkcN2OM6ucylvJQdvkvYqhFQJXP7LqvOePbF41wxgZfwHCihDFWADRJpGhn
nCPgDX2SIcfpsVmFtinAMsCGb/Ya1JvFHFdi2gOLAgHmFrjywhVowocndwrr53Ze
yzxqAB36u5S0zOdkzUTy4BMRBHpRsVZQt3EH13SITvc+EUEjRuDwYFGoEswUuOFL
4rmmL5M6PS6VO2x6QB5nj3URbIudQsxduZ3+l/js20+fQQhmAbVnqYgos63mfCaZ
VcfH+19dEWH2noVeDhYFoyYDO9Kgp3Y0WthYVB4oUyNCaSEY4AmYFk2GNVX4x+NM
h3a1D8w22gZeqfgrFe8VIyJ0SnjrtZbgWVRmvfuBNcCSiamRHGhzHN4xAYJ5XeUE
+CDVeuQTIYlpO4znLpJkiDzeg9yPvkKWeGpWc7MY4vQJ8wzCwvc9ZTSS4Bngoqn0
/7feKp1fRG6KLgyUjn8bB1mqJI4hnW0/fel7NJ0709/HFmAO+kWcCAhjaig55Pg7
MCLQMgBLINV3LayGbUeIaXbtLiuaZswn9zEZ/9EQu8mMMFnPxyE1BQ37frbnevv5
rx4PjXVzyCR6n0xlOjgsYhRG8oKwTgr9+V9azMrCsp+qdJgNPl4vmEuqmoD/Mqux
x4aO4q7aHTnBifhEjXg10QHHY9uhr45O8YvzvlKaQgdSrElXCnqWH0Rtx7ZclPxf
rhrbgo+qQDrABlrptAk5dtX3SGxgGJmoHdHs1/Ap29sxHUHxLG9FH3gTuj9gV0x+
q2oI9vnKYa3VQvTHIB6VMogU8PVYHyFJfTQodnz9W5RsMiHLKOsBSPWjAogXVw0X
gUg/sU1Hrk+L3SvOoHT7LWaskUya1Rn7n01WTOC+9pH/fewTgq4I91KHWXonw+GN
gwCx4RYeWjrgWRbnbkAva26ZeWJ8vlGNiqfsHSvtQS5SyjMstd5EbZzrH6U2QiFj
KIlqJYYUpMQN5VM2zCvKRPBlMRfQcUStvbu9TJa64xRG4Ntf20k+gvn2XHtF+pEV
DaECgwVVnDP/QL6IyuJojIYVBdEJWqYKpNhy0FyL2Ke7DeTSIXm19yxNjgICyMc9
nObdATJ3XAF384pXlS7KEhIyimySKgEnHDHAWpXLT6RpdltxTlb0snYItky3/UI/
e4H4O4klht3xhs3L7Ln9/OScqCAWfrvKUH3tsfkqC+wWc9+Mi7xBy1qgGZ5dK2Dz
FaQ63srfTlFAkU6ozi7Tb69rNG2sbf4DlFlkB3awOo+1yCBVth9MxHixowDd2URr
3xR97+VyKu6wrJEQONJ5TT5SjvA/C9ZkrGEgefw8BbpxSXW7+m6mM/MAgAoyVlGd
QrO6+AfDwoXao/8YE3oXI1byRG6itK62kWFDmU+/lISGKZRcLk25nndpAPk1pxXR
sV3y6lbS88M831OVzWKJH24Jn7BVuu+MF2DS6ljhD9DEQ1RmPwFDaFgW/S2NGSMc
We4Ph/q2dlgejrarEMuhzeyIY2f5WCiDQZjnkhdWLRMGtwPJ4V3kdFtRDfKZQhip
np1trgAT3DwVq5ooZm6couylrOabzMuftGn6SMUwanGXtEZUG51cXUANeYzKy69x
a2DtFVEn7/T+QKOpIP+8KYSwFLuaV5PQpB8xxjGYvmbi3NlRLur4a5Ae4FVAZxjI
ZDI/ia+AQKb6o8EiDiOoK82hAAJBMfCjMi+vadP01bx8FLiMigbN34e4TU7m833/
Z15f7KEaDNJkBt60N+dX/h6qQEQoncfGJEf+k4QWnAYLWposLhz+nJ1UsoMMhE1B
/FDKF/AalxpthnNUJ6lH/9T9kaXnY3HPgbRES7hh5/Eicpw8511IeNZTG2PkuBgA
TEEP2K9pz6RE7lheU1bTTgZ/hslrBqNkKjbzdN37nc34BH1Ng/6jKb0H9NT13AQQ
jhHi+1R3UrtLVA6RwQFHBn4wPoL20CQExbumDmtxYyww3EQ30nfCpCX4d7YjpU0r
ja6mSLfAvz4DRLkEa6Ca9EZ7EPvYixRsvQqKJZe84J8ehAUSL+HS0bUEd8C9IxpY
jlJ6FcZ4NemvBE4rvnion7oeARJnLI1AEmMcW5BJwW2VIAxJCOkcH3xnti3ccPHl
6RY+S35uCCyrFUvnaIVBSPfyTe901r1hsjd+iVul829eLYvfoIeorZbnfAYdME0x
hr6rP+ORP0NrrMlJoQ4bAGxQH+h9lCpoLXPNWc69ZFyjeqY4hI4Aqe4BCCml4z7I
rldG4dfCuPVRBnng2A4MYE7X3uaNCvVZQ9w8Abp33q/ljBr0Cl9/D1Mfj0gMltqe
g4TTYkJZGBW6qkzghMOQIHdWzBrcsHxGpadLSyfr6C0FoAGdzH3h/Kleds8kn0JU
34jhcNKb4tNxaKY++/GxtRrBl7YAzRFXXxdHwlKnI5/cpKtB80b8ikrknOGNr9dR
phcsHwDi991vZuPjELulArGJlTkRlY8jpEARmIgp8b2M74Tg+BfVAsaahn92oVQ7
4/hzVI3GUrdTVzO8viP7AAQHPCIP5IOhVeoLwmjtnNmL8K7EvQf+hsOYgTj1FLCZ
b2g+6lLtiaIN+FINKe1bh/GqtQS2vV4/60oSbLhSfsG+O4BrcZUgJWRMcI0icPW6
ku123DrJskYNHqTfk5813l9uDj7MAhM61fOvPbdnJyzIdkSFI27QTat9xPjeTK69
qX1js0DTot2sJoe7iPlDB3LU3WAWJhY4JJSPDPVKAEuy63wz3907ie6eQPkbA6Un
ZS9ZN3OycbhhmPsbHtwZNhUGKwu9ffAseWbmFEh/TS4PQF22XS+4jri4LDpm8Wn1
OCOeRlg+9GQfutmNLJ3BeVwqgSa3j1qGxSnXei8MK7eo4u7VS2Q8oa6n96gYLjZb
KjbUea0xBEFkavdyIHLzzuIEtJmfbYuCEPVSPyU8sU2XQAm0zlEo8X++e7EffX+0
LzsTyLRrr+YknGXJvFGDAfgyDIRKN4kfRU2lCRjfFoYOcJR+CR2jFqbHYIaVGbN1
7EgVjdPK2L/UxtTLycUISNdamo1kgyPPsz4PVLIF5GBnTuWYFFBk5N3cZOEB9z28
imXAmEonWmxVpfp19y8raB4pq5KbVwB4M4SQrhswwPhqMnYqsjjcbtUjDrtwci5W
6C/nHJWy332A9eCUvi6dEsj+/FuS9+HY6aBHYgPczpOKhMC4Ps25fquBxRAlfbbo
RCsszwE8Hbxjbnv1v7XUAtcdU1nYOwTMXwxaRpCUlZ6xksf7eMkWdmNMC34sjh/h
uBPje4rYOcvtSnsv5/UF/B2W1NQ+Wi+dykReGXvbTCfuya12D8OERa15X+2v3E3L
SSHAyjDGM4HuIZXKstVzH8gCyJ/SLfp7GV6SGwsbXE+G/BywlLMZZm4eLbHzm/0b
p/ZKLIP8WSkn+5cEXMpNPuehStIEsR18ghcBdOBtQg74H2WpXzUPYBYoFBhtcqZZ
6OYmb7D3BDowyxjo8C6rhWTYPYIDoK0FgowejVRSSIB4dQ8//BswrCR7LZwAELGk
2fIfwi9v8ECQJfH32OQM0YyLMsnIIjG1PaomS76p/VJUGsTr/7xG77/XB43D2Tvc
Pn94xWpJKEkRyMbEYNDrr1pK7f+qgpkpUtFax9OA8O/YDIK64XER+M4dv2Ej08Bj
1fzT2SZ42rfeRyFdw0y9u8t6bSyi8hfTqwpv60EuypYYISkd08viLoq/EZksaCw7
gJQAdSOkUgdAPs34sWOIg6Tp1wMVsMJkrrJqS+NObOYKBpo2Lbzh5io1HOf//9T1
NqoC+la9eoa+ckUkKpeMbX0/wWcAAYcDhtaOiANtZCdY+IJOCIsLtbhjnj9Y1yWi
m1inzzKH4PZ0chFnvqDjatK8SDNcEPFYOPiGckcchG7giksHPQAPif/KTVlPiOGn
VsTbB/XFiFTCEIngl1NNEnBbWFAYkt6yH2kg3j5WIVJs5dQtjT8jOyjL7ngA9Qif
1+SEr15MfktA5C5cg4coEpdEKoyDyScf5m76yhnA6Bd4Oi4WzaBMW4H/pamHbaO0
YDgyssaxlMySQzPwRm0RQ7o/ErFSacLkZFA8XrGBtU/nSIJfVnjB41h5QUNdHOSN
YCLQOiWf+O+xI9tUfLdnrdCh5rMmy78dzV9A5RkPXfQQjA7pr++V3ZtPayIB6t0G
8ajiaHtsuyzQtzlCtQjApGRwEot+CitvlduSjRXjJxrRnvFoxptDxDUPCTheiLog
2WywKcNooO8Pq/STDquAcyvC9mrjVezj2ZYPI3X4CRLyeydERnFgnAliuXpuVxSj
NSSLjo3HmVGNEF2u/qYNIv8SH2qJG1qBOCwCi3L9qZGTPaBhDpARtvt9rgxXFHT8
R8qmJhTvbxsxTxNRTPcTmPl0Tj9CbKG3h0Hik9zD0OHN/ltqmD/vR8fYlcBPDixw
OMI3wrkJd5pjAucCqqomqsdg1kGshpmni5WRrBVVPcQRzpgpQ9M6J+9Pne2ifu6u
HlXlzXdBBUt8aoV+HuOrW+HwxKaWc0Lr7GLBkRtrVt/qLdrBkcNlmPwy0x9xQakw
ZGxH93BzYGELOzGOIELGHpmmz4gu8hyJ1wh23t1wQOvxPFLA1IXeLon5gSgOpCbB
KPZHGCEiZpz06mTx6Im9VQeYgokOAGTqL+c+QFRfzyJ1W4jzRazrco0T+qWfHmgg
GnjStLZi00/9utL7bgwa3JTPEAyWbBDh7l0ec373xtsceYw94u/QyKlileeU9do0
0pWPcLusDSgi/auDeLzb6/P9txQ4MjRlBYStVoV+47ApNzp6mbMo5wPI/mNWRO1n
Db3TjDYCcFr97oHByPbuMMrd7rRQEAaQ6PNoz9hU2z2QAJMob/OzIT3oKjlTeeTn
EWlVType9pOA+cOs0WencKXJIrefH+xGrp94/oTPg9KkHuMQ6hRPoZOxWZpuIve2
wY9vzkO3TkqMnIgKIGVH3gY6y7/cm58uBUxXTqh7PoXMPCX2uepFr/Z3wUhxsPS2
Bx9Bed6wJrbW4OtygXVTOd0jSmkRIvDgwbhjdtxciIHzVLJ5NWca1zgLWU4LJe27
zHNr3iU9+UNv4QY3POSTYUd7tfeAxx/SJx0waquJVnCRW+T0GPzYVkIDeokF/5FB
V7unzVimeKv+aliyuqo/TvlzdXt9njr1xMOtJZikbeXZm0VWGSIbCIDb4Sv0mKJo
CygQ9FKX4xZ8Hj7/iXfzwKjti+VsHWFULN35MP0xbxSPwIbrPBwSVmOGbV5iuE5M
xPDft3oH339Jq0muST/YtsiJPaiYSiUaVNhO+pewE5LOyIToT0ijRCbYiGhV3GHm
j0Nvw4Nit+vpwAgeOw35UqFhZV31WKcEWjfrGAqwZEj+IOQBhyqhuiSCFP0M7XJN
ixHP7MUAYXS+hNCFdMA/P8rjJGMoCrTO6l10CX1xEikqjqqNMEKP4WHNWfXUEtDJ
VEsWYK6qAKrEibLxXKifoegSUDUR7zWygM3nwsib8fPnIFbFT/JZVFHGs+UBveEU
xyQOBDKJfokQnfXOeNEtCTpGwKhCe1USPC8c0dPtHBlJuRFr6tTydJZjcpYlXLre
ShJCzb+ivhRNcXKqpKQGKW93OxJagC6qwIKAxs62H+lN79gynDiKRwOBFlL5lHB0
oE9dIf3Pohj2C8M1XaStJICCxkCDI4S+VOkG0a3YYdA+mq5LWGaOgyGENDNXD4Vz
dcgmrJhNy79T5FK9eWgXz1qXvMv3CNeUztTPAEBn9c23+7kx5bZjUpxKp174MtsS
IkB+c/mwAcL26eubu0iFkRqNwZg/KM5cZptgEzOyy7MLAivc5NROfdUhEU6Vc/89
iZTR8E3ma0fKHEOLG0OYlY2fADb6eGk5CdRG3mYrLChoK8IZnf9PvaLB1HUC3XrR
yTcYCN5qZvhnz+6b6OhOt/q2ZhLC+QpJeXvp0YL+aFb0QVPZ51qeKLv85roPljSE
Irevm03s3r0BOTJvLAywy7DwNPb0F/dfOQMBO2ubXtuusGVFbYb2ua0gVjSqqFdR
Nu1I0fD3jHGd+JHzsxzLYFWBaeNKQgeZflAGRX7qZxFu0/DeQQ3nnXoONHncw1Lx
fU4PFLQIb13aNxhwPQH55xu4USCjZcGMy/Wg0/7JCEIHx7PhTwzzXnDAhLKdk/Ro
y61+jD0ACkxbuhEDklyRonhqAd5q5fTD4B65rR+/dx3Gmm8M9Ua3PSvDFQropLag
O40roZkcWz9w4wF8ECA0PVoc8WOWSb9D3z4lMW9N96La6IozdWkw57b9DBSL0IJc
7BlMvK7Q0gry6GOxiG5smKRFfsZJlihM/KBhAjouqsZlw6NABnwadQv2NYJlKT7x
eLzfsqwwqirtC6LnCgSRazEPQMCY3KpbkbFdJ9j/AjfiL0QRac+5q4SJOXrFJip4
faFO+J1jteE2YYwpepVqE2SKMvZknWw7i62lsTcCIJ7HO3ODM4VIfkVneKGTQbaJ
rC7L9P7SlV3gbqE/3UvsMTmlq3YqWwjPvNwYa2VvVjBPaMJyJY1NwXBe6TDG1YBi
Smw4ojGB8RxAIsTHF6yOaEc0XslTqoBjqO8vdFJ4NBVreuDuGaPuROkaL82sb9Kl
eugWrjjU7O4z4ktWaJ+kbiOoXTXK1aPohYgxWqngzfdlD7STq2EeHQeNd7l5QxrG
N/HuX5i6TVoecL/6LQ2TR3OL7sY66LyLUvzIp5yMNoq/jnMSvSySshCiW4W7Uj1G
2ljvrnbsvBTHUVl/oI2/6BzOPOjeBNgeHNo1PDkiZxjvDgOf+8KnhQnSZFYJvUjz
71afQL2t7WrCdPrHwcYHSMqpvGGvL1/Yfcv7WZNrboF1TFxgmhyU6psaQGRxJU43
Fx98ognjLBN0zQ/n0y+YdAZpAaqIvmhvbdyaPD9Ifd/9qFM5o5gq+pr366SxpvYn
XeQjycMthW+GvysvmRdXb5S6tgFdS4oMs4JpntdEWIiE4b/Xh1GqPlgw9mkU28HJ
r3ie0Cw+GSIuIFrZf2oGQJIa0yXZOVM574rJDFNR88Ubfw4GACQSFHOBCTVhuRum
bhZXjvY4y4dknl1UAyrr6oP2hY/z/uNL37C8VMy5bvH4gVFtB9K20/UJP8PqFHwQ
3nxLgDfTjxy9mf6qmvmI4eG30bSSxxTY9G9mAmJgxfwLtZDWfHafheNeeS28fXM0
skyJH4xlPLtbshf7diGA2TyYKmQOy+O1HRBeOKR5z5YgR/tvrMzvUM+B6yGuez9L
DalFEuZdosgMO1/2LdDf+gtIqpoXdwmK7x/Z3QOKbZ++zf48vSVc6BgDEOteWlOL
J2jd0JpWKSSeVkOUy0boofvbVegqaitGGIERClcXOAOgwJ3IgM7Cmk17lKeU+XfF
jAUGG7ElZWEfTsVtdWBveB77mtr1rLw63EaTXiimDISRm4au3rxh0h6PCeSws1sw
dD1yvGKqw8lmhOK3rp3j9BDh5f4ep9KzacHIuFiN2OdZuCzCFLmAk6noZ/tA0Mg+
MKOXZYJSae79lTEU2s/7As1PaQJnXjMuTNy9KqH7Eut906s/I9U7+NcuD7ntrrS0
1GH6sQB2VGikBkPOJZ/56nH4jAsBCi1CI6EOZV+87SfWyOSIvFfNdJPVkdwa2fQ3
/ss3VvNqDP6kGinplNLvZFXhchdQ0ylVy3nWb3YNtLjSK21Z7NoQAIZyqZC3Gumb
q6unI78uORe/NXjYVa8WpDG3wDXTTDQ9ChOEFQJyWiv22CXMWuQPrwoxUkz2m9XA
iYSLN+5LFVhwlk6bZVmU8s5ZG0/6eicYFOrYBySu82/fC8QjJVPUQYIgrdEtYObn
tNBnre7ysg4iqtSZWCk6kEiN4FZZf3LNBj048h5ZhCcaVAH2mSdp1Y/uaAOkBBcr
XQNXd9G86knpElz9+Z5vf/xlhSktPKh/CtLT9PBYq+HJPNwjV88e57aCITMVrBVS
TlOGruqNwjaevrNB/10HybAGE0YH14Oii1qkZ0UbXwNbwj+oyUPHmJA4KuA0EoIK
7FvHYIwOZ7z7OCPUyGPCWO8QPk4xKD+pXT51TzXLejux0FrfAVG/Qnwe02vJsQ8o
8QCicQ+70R9IuBrr3WzPqMNdpbrtjj8Xzdq4qp0WR5tgqJ5InSSfZ2dfzIQv46D7
gc5LqvzCsoPWw5gSsM2CdQExNMQtyZHCuhy7i+zjk2ziHOuf+l2HdUO0MQORSry0
kktWwNzyrAqFyunIuDkbzPurd64ze7ZkAIrTckI7d8Bpx6FnBuoZJdIGG7riXfxY
SjyV4n18Sx6EM8eydoj1a3/FTGxOyN64Lv9o5s7WqtYBmma4WKJuuQoNuk1+c47Q
aD45Db5qoSu3dA3S37vwK3QKosUFFQjQVMVjjd2nvmU9A/J6zQhSygMjwRxU/Lpn
A+Vbzlwk0IGXjL/sPCIGBJeaaq4Bf8eJXEWf0DfvexmcsWaE7jGT3m9WmAGzrUA3
Xy6tgpYGcpJeQ/w1pQfqheui9fFQfW21BT5YrtSDBXn7H8tHFsL21YJVTc+K4CNg
/cy1a7+AsbFqIvcwBohLfAJuPnU6gw8o0XEZBW+CkqbjZcTUlipplZf+hYYGJTdU
YEEN+WQsk1YLsTaiwJmDtbL6iHv++P7B9te2ibJztwjMtsIBxIxGrbCBZUe8DfyI
tEjRIpdJJ81K+2/aXQI15pkaplI0ogQ/V/Vs/0XOhpVY5phxVnnyKUYfRP6QIK+Y
giFffUKcPcFeaRYjI3+FRvU1Im6VXFUXUE0Qda/5kXkKkat1qndJ4X0Es7WgQe/a
YPSDnGyQGtJZhjwl4DkPGVQ/GGU83g+tbwye5GaiJp6IktG7xuCwsmZTQUCGbXUt
61e5IJd/3gXGcBLbaN1UvL5sKE2nqGaZt1573xbphLY0gTGH1VDdZ4dsoKHQpMUn
rs/Zy0eAJPzAspwDjzkVEYfvWgJUu0BO/pb7DNfiZPIUwaMhC8trsRZH46CNLmPT
BmU+mbGGEK0yXAHLMj+flgs6ji5ucqr2W3ai8vprvvweUkRVVly/aUJK4DoSxs8b
Hy6DjIZ4CkE4XD9oOnfNJF+2Vokx7nbl6oryHJG8ClZVM80r1zr2DvUFEX8LlyZd
IqQoiiSneEWE4gsz/TA5c6MnjvU4wvKbEh+zWNHCGi15CFG3+C7JZPLumavceWF8
9024d97FlQcMY/iFr4ceoSDNQ9ktze9gERxXnUxOmyI+JzCQdisdWvd8Tc+HlWdm
MZnr849Bp5+tvvEaGDgupGpHhvfbB6XSqIgxFgcY4m50LNbwFTCcTxCqsaKRCXwT
2D/1Y2GiRqiUsprGw8TBPZcaQ8n063x8OV2YRdInQGfuFxsAAOVEJYxSnDge02Zc
CNgghNr9sYWkC4cH/FH2y1cglx+QwwsVEoPEQQm5SnbeVQLbrTwlLfSK5UC86WVO
yZK6ZmNCrOnRRlwuGhc3skG9uoS7B8/xwkVSbx+GyFL2aqXDl8k9EU0x87ugRbT4
7maQmdhgX4/jeDDg+zNt6370J6PpxoTIGvFY9cTrpis3YFVZmYZsYi3JL3UrNXg9
HdtqVRgNRMvCW0293fvrFCT1+mAWGjSroDURKLosFqTwAFKwFanI6r26d7/ypJag
dMza56u8LJJex9I+IBXBrkl2QjTyRZK8uvRFtJNqFUsMBtyRtnaQY2jMA+Rrs+I5
/qIidWlzGukYE04SEpcipC8I7CNHRb/LF7BJKpK1xkymA5uTGnx5aDOc7v0fCM5K
u6emqWBoxwW1vcvkIYpMrNlKNQGV+fqYfLryabDYGyCgepCaKlYPmNIhO0YHpuZo
DpD/girrq8ndtx4Pw6Fi0TqJeAZRuhGu0G3c2XnDSOQtkSdxWNMLjhfAV/LtKWIF
x++TuaID+eLU6eU47mhXJcp9DBGb519pa90P2RMNASk1LSUzPbYGBFo5+sEOunGH
5taHzc710iG3n8394rO+bpOmSChbTQTgsqTaGvZjDQHxmJdaQc966Sas6qx1Tmo4
3U9WclI+l5qTG4IrUlYSwUPMzvCZWST6CBUMFC291Bi9kjM4hdDfLoinyB+R8KKt
JguDIkv0eq4yH1fmoW62spdwFf2Y9/VNatbQO6JJOznLfLzv73sY7TEYafiXmp23
vd/oGUfsjcPpV8s90Jw23sY0oX7wSYruF1xO1qSjHBMaH9xdVPl4SaNqI7wGLtEf
JbdeUJD1e/FIcjNACezZD9hlWyoKyJ29LJXTQJFHbd86VW0u+BTkgcbfGykwXHDS
wPQpntJntqvzbkBx9xc8knyIMc4GNACJjbl80m734/gsRazSKuZ8s/VsNFrdR3VO
X5NM5TL6YxIwMe5/8hSq+5KS7BchuCBvHb/LA/AHRZKMQnMtb73G5Q17kR8rpJP6
u8lEPqQK/OJ0F90xxbQ1odJKjTkHwihcnyjOgf2QihQu2Hufw2kYHxIc9xWgek/+
BdmwlnFziubdVtOtfTX0v0czca1MyFfIElVeTdIA8eVMsIEQp7mWjtmGGqMu7ZEo
uukb2//76vmBLuF0PM6m8/ZorgWXHKWCkO23qiYDN7QuPTxND770YdlkMyi84U0f
kdKMvEvKQMOTRhaMG3P3a1JI+/ReVodKGYEmhNSLlIo93JEJwjmefaCMAvab9ybl
kZb86VAo4c73UK7l5WpH+wLs6I/UREW7DhcnBxHXh40Yqghy5YpxOSTXyTRkFBdF
mP/OdrtvZyap6128q52Eg+Tjq/wmu4T/xVvWKKvO/eQQcur0Kc7H5z3XQocpBhdt
QM9zd9U6felAXL33HUeyNlrhzR0/TkDo/d9LVHvHa9NS2rpCopf/WU73xE8dezqJ
45w1PrazOb0iMnbq/50hBQqJvRKnHAkfkaWL1m0UMybgTT3VpZliEglUyT5gEc28
wSTUXclWE54opeVrXWvZdJ66sVjF+0RFx236Xz42fLqwoT/RUQc8LN/AxIw50cWf
ThSVJxcxHabgbow5gv0pvawwzUba7h8A4quOllL1KjMpx/Lu1KXT0bdaNLVDaK7y
UEtmEm7BNhXZynC6jIILybbW8TuENvcuzqHM5mgvR+N66JsjrCBEcMQTzRQQVOd0
T3WSMwF/jO63GT4APprBWZdbI18YlBFbqM5kuXfF8ccAijeiSby8+ks43Pc6jEWZ
Zm3qB33Yi55e5aSWf9CSyIxcL7vn67S4m2lcwTq1Rfv/5fEABeIIgU79XzNpGH3a
vHEoFOaLfvhZlBUVNlTZCQamHdFeXkg2X0C0S8d5DqFeARDCJvXThqDGcAiuh84A
NuFQAkE2AMrSxUg4168w7/FL6Nllpt5+MM4wb/YF/AN4KKYd1avt5SSkbDmmU+DU
2veQK51Wl1TwkFMYYuIAw1aRRHzqOERllLe1ZIvcqsoceb9I6g8/vWhpZ3sr6r2K
guDsZo49NHBnwYjLdElkrDJ2Qm6HrESBDnE4Gc6u48MXYoSQnvRhS0n7s7T5YtJh
XFsnaXpLdkcqrDf6UXnS5getCx01/IysNqudMcDKLg9OWmFOvYNRVN7G3T0/MgPS
FHAv0ZeiuS6jPurVjOqIUBDH+yQHiIMTUDhKF7X+auMwSvgPAyE+2HI/sB/zsq0K
Hew197IKxV2ueOQASVjXM2d2uLJ5xXSHamxh7F4Kk+crJBhhQopNdNaJZ9nlE2mF
lncbgcumVj4bIQkLwhLhlfVBWO0WH/j7Ek5BUQXLicztpaFyt/haJVwAvKhBJh/b
4HHi0ID5WCxZHBqVFjBHx5yVDg3VbSYMTQvYAuCYxAiUNPZPOx1YEXTeuEwXL+tW
JrUJJkiKGm6Qw1bXhlMa3dq4TQ4ebgFLOE+rVE9aRVxWlFKt5jvcPKP6ZQv+SThr
ouiY9CSpX9d6LoJSe2YJ65/0tIyALpz77Leq2fIidqbQRBeLCymP9C1cv9pknLs3
tQ4LP3pTwq20rEkNUTzGRUmg2n7s1DO+olssnlAFis6m688EsJ5fUg5AQZl7FoF0
5KvEHMvrH+F2NHgbYswFwBLcD46LgsjYt1Kc5fAUAbLgM/XN3W4M9jOjN80MLd95
w2v0slhfSs7kv15lJP7QYjY58Q0WW54tPsDbqAhE0RVLUs2lSPRiC11OpoXJ/8hN
y4gRkIrLLuRSCNbW76gy2hXBm9wE1z5zAQZJNZnp8jQjSxBFegfAYe85VMY4KTl/
lQtQM19N/ArYsYxrTxzPN+7TYa4QQUHk0YGuSDy4lempxCbHMj9iB/xnKIDl/cqo
H/aAJHpOv4Hh70nQvdueWgy/Z3FTnhrhGies97kVErKIEo9OAIzIDwhRZ67pMyMs
esLBz21SbT7UpenNzRVQLjUVqMIkn0m+WPJq2ITIjq/JCt9V/izmy71yxXI4QoJC
E9hv3Cbr7ahiyJZjsVhKLXpIv/vkv9Byzs0dm2EGvRmUeJul37J1fuwIwCQJSW+Y
bu7A2rwGNGpzWL3ld7NiFrX8YUwLcurf1g/TAqo7VY3V7+oZAx/PuxouzlA4VfOc
ojqvpyBMprM272f5TW5l6CiKkaWXvxVx0HxNmrPN4EOCu463spwwe9ZjQxnzLASE
h7PRVxUjReDNmUYwQgNk6Uf7I7bv7zF0f0f+rzbuZYjEeT4M3O9XaJ02XFOOr/eD
1OZLdDdFqjHfVFv6a/7Zwq2BM9c4ZWqxSX5n2ZOV8kkVcc/sYL7BOkA6WTkeZMbD
OsVGW4CGH9PmGHoQNlkRMKDGSTeYcp2P0VX4f9L6BsnISHtSo0rNZaeFAGxVRpbl
Tt5Xt7szcuebDA/jMbwMv2w4ACc9nz8xZAoHqFKYjQ7WRsYwysHCIv65Wu4Fj5xT
uCPFMLxKUnfraDMAEZfYJSkQBygsSskefg5pPQonwvrsrz51rkDBARQ4QfCdeXBG
BtJUFtBbGQqrkszOCh35fajpJGlLUcELAX/wzOIOnMx2zrgHFJ2kxxCIUK+m/res
7wpLHFBWNfa8TahLR4k5qmOfXI4NJDb1jI9V+40hj38q7G9l4EAe04C9+pshVvQD
4v6pFwC+MSW62a3Ei32EAwes3z34LYG/eN91bnklrwveGwyN69mqrucfzKkBHf6z
UYz9liGhgtdWGFwy+rRGd6vniJ40TNLudCfgAYe1mwes6y67zJGE2TC/9JYbWCwy
cTJqh65Oj0eGCztdXoI1CQWOOnEwcR2XNv7Ohi0RXz+A+7PlHmoYhOiy2FCSFz9F
/olYv8DtcXplQzVbqg7gO2eBa/aj2MGL9xo7sBY1vAQmn4r0BjyiHhwJMw40aZYE
b+TbE/rHHuC+2E8j4bNRdxWz9MZiIH+IR1JvBq8lsX1zgilvIL1qu2Ct4FAedoJv
JnvRInTOUl+Q9z2SGs13o2WKFKrG0FTb+fQIMFbNOpJ9n0rYGuLjfY6voPEoGDfy
XPSPSVWskyYZZlrGpNA9TD9IJio2PntcsePNdYWSMGzUnUmOVPt1mvx5T8VkNM7n
1vBi/rHjgO/C2ZSW+BdkIgQ2j8cdb8mf/p7imixZDR50VOyG8w/qYLOXf6zjsy+h
onegtm2wktKL/Nv+azl9BYvKPNpPtmL+OksusbCe0pFzBZ0/wtWL29HZIFgMVrHD
V/OqJw9aA5KA4DkN7Fwk3SX4/ASOu86SAeVpcbAz8GzD8zIusIBQ+BhL0i+pKu5N
SEGTIxrVsTJc51iET86SEcfMtpsooNU1ieuPmRbgEaNxKaH9CdpS0kbEje5ecmcG
f/8DaPOqoPOHT7L8K54M0gJCvmBpcU3FxptFhXKaCddbFbZvj4Hre+rvvEVtQbXo
6JSfX+aI0m723gjPJJW/xhYu7DGiqD+QFweGXCRUO3c6aXY3YxDJa/bOZFWMT2vd
PtDd7b9v5KnILBewdv26OwPgqIxhgLsla/qNLiVCs/OJPo1cOSWFrn8u+nJUssuv
isI0Da62dioTjT1FLMwUE4FlLAA2CbRoBAPprl4aCdV3MZLqk4YvPgjxIZTjCfRJ
DFkL82nvmDBBDOhw/kMHpB8E6zD6Ba85Ki7Swf5WtxV7xUoxxjMdMry2Nfw2HSGB
hDAQB/5u4LpJOqJ4IOhT5ZxAViawNYZCboxb+n/NzFTNOySl4nyF4dGzlED85biY
3eZsAoapx86qdgl7LUU2fVoiSE/oJqfR3fBIjrfJ/HT4aSFfcvRj9GgK5Y6nmgrW
o/qtFHKIdlTH9UlUAsD2zK2CrLN6Lk9SdfvdSepjumdKM9LZK35/V2UUsPgCtLfj
r6VFqeQ/tfBVh6xJcoNstgmdQDR6vkl/RBiDIknc7ysgFEO8mlBQGMphEq2J3Wws
8mKDTQxakV0rNm6R3ENc0L3J95gWd/UOP6OXXAdF5DJ+HAg0wNU5CCqE8zfYT75s
xh9XormVkl87IpUQ3L5tocHT+EFmT/CryJHyRf+EZ2e3nVM/WJL90AbW8zqMl5Bz
mAY/OzBI+lv29EsSdOmiyCtQgOlaSRMDM4H0ebFYGvf/V+JJBh68p167irOauJPs
FwXzFRzW7is9gMxjuH5E2aXA/l4HeKCbRfU/DElJN1/kGAQAt5D79AozIXKH2Kn8
CE9SyQ5z2A4PkCzdhMCg80uLwSuM2yL5WhFZgqutMAbzkYs6ciSFXe+24aYALan1
3MFUsjRLE2m3l9kEnkaAH8ew7mPY1I+EAC5LNpA6XEVI+FidF2oiUsdbh9pnbI/a
szMFe7GD7AKBvvJbVTa++RguKUfu2cgRd3MfWXlQr1nl6tVRlvi2lImbdgBM3gGq
l3iepot7S5GiAQDjCmLSugbg+66cFNnzOFZJHaYibEg19CrXtqbi3NxplOKF79wf
rtunPkJ3Si8sLiqOerlxZ7Gno5UIALDUrlh0Hs5YG3VQS03seOtPiDZCiyAcF66c
JxeArh8eWis1UWmfAxBgPpAvDrws5tRC9k9k3kXSJzrbiiyB3GqD0cbDLYbyiJG8
0/lmFKhAh47nPhqLhfsL1tU0N+15kzrbu4CImtOV8UzSwhLwgYE9QZFo3zvK3Fxs
VPbwk3irDG+JsF+CBdNRwDpuhe4Y8s0uoa8SjbDLftm2OPGqhrBUg/5N5i8idkT2
Zj64tx3J7LjMsAbm4BCqKGSfeYSN3Fk9dB7DsCPMS6m5eNIvigoGi6Bs3D3VYEX/
BqMH9CdCNeiuUk+5w5QYAWMd99CGt6q9lMf4PF8rM3hmfFgSe0neVxHHccyFF5hL
RJV33QVfWzRoMcwjYM/X6/DphRaQOXNcTQfLpC2EJqPThONdbt8M/fke9czR8yhB
xa4hLXaW9tn6Hj4ZSBOkNsCNIPJVwC67AYgXwrTM0dTcNj28v+PiLVH6IoXFQNUV
03qHoog06Z52wHDAn7YZ5859+pJJ/cFiHdMUlM0VvEwRdkjxu5p5Y5mW49w4i2eL
oVUp6NMT3W8ew8cy8ht+aOGZysVLuauXqS3oMrPTO6Gr0aY6iXBaqb8+wr55g4j/
pOU4+oB4rMYGC84xRAw8LIA3owfidraApby5AqTpw73tq6zN2fBUtf7g9eB4weHJ
8V9kA+Krp4Ugq/w3T6rcFbuNDIjhIwldBVlLjN0KVc6MF0bBvS/zhNeHLFAdhmeO
/NGINJTWuwl0gXLcCS7Y9vEcvODTpfnvZ4qRZ6RbQsu3cWXR96ut3xnA+xc90h/F
0bkge/dFbPl0MAHX01kfxKjy7+wzBGoNopOvnfOVgKnPHrikYkDiX+nvZWKDO2Mb
O887tmdzBOq3CWYfi+1JL7UUC9wVNuHV2PyLtriN+c6IpEuHYpgFfDOB5vE37QHl
5RjdHeIhV9hmovN55JiHAigdJe08OJEt1xrWamEdCXT0UAA1XWuIsWNly27WkhHf
GK7xC8ekXsCPp1TrKZc1qku3FUeL2RYi5Js+gjYifAy3n6vA7fcvH8JNtCJqYI9w
IYuQPHosJT6fObSlqPTfHWfm42EI06KFbmVH2t80z8q0pukuQn4mbfQBHNbLh/Bw
OK13MnSuiPa6bCZKzs8BHtZP+7e7yvz/dJjv3q0uz5iaAlMXsYIDtjOmhHuWdUjD
fecafFMfIJysMw5XGYJtY95RaYxRVB+QhpCWXExYP7Fa3iocmZZza0nC0BCEl9L+
Mf6rczPCgsni/X60keWcu3MMAR5W4G282P/oy7q1bEbDs/MqPYTSFwgZqq0Avwsw
NZQ1rk94J7SfYxkBKW+WGYwwkGX1eljpMxnVKTbX6rTTu4a2sT5OOH1o6oVX9JZ/
kZCAeuCckKf13+33uhGTo1WMgXQEoE1/us13dxWtVcJAyOmg0ya/M8bUod9lxzm2
fFTNbVmVTq3ylLbvK1/jO7/detTOx9xXJFabLFc7A4zPEHAGaZ6ENeJ//GKuQTBw
sfalTcVQcPii+jPCK9LT2Xjq9kXCFe+wWFh6op4Zqa256RhweB/tDQJPCKb/0/zE
cy1I2FNEf9AiqTnz1vKPqeoeFBrr50gxST/BKrb/fbtFyE59atsr8Azl8rNhUmAk
/B8RLJ8TqrB6DJX1fBGrZ7Iunvw2hCb9530CyqzVAeaulitigaa4Cf2cmyt4A4+Z
rLCx0YFU1EHSdwJqh9ahT6h4SZHYJPfU0YOUMNz5v9kulzx4wQgvkVvKNuEBp5+x
esvjS2N8YyPc9AwEIius5mspGkhdbOC8RrxuINZXLsnLsog6YGRTsHRHPPXGrnry
TBBgFSubSQgjh+Wjz8TJgegw0L4QLNHCrUHRp2Buz4pncOTG3rdWr9ODNxRZjAcN
HojAImtLb+43KeszrnHG9szb9E0+F1qKqO8DGOn7gynpgMmFBHqfLhjcqT4RjVPn
vBuO8FaS342w0pq6UcQWBWDwIIhcURmm5u4DU7u6pCNQ0wzzZ+KJEGRSe+5aZShI
U0Zl4RPX7aTGlb+XPpQhtNs3dGBsP3ISODGDfItLipZXknE+oCDBDfb5FMGYxz7D
O7WG/YV2rzlu/5QolSHKY5YIlP/3AjRzcqG/I9bJO6ffaEXueUZCwbozm0MolTgg
gThEh3L9hyEJH+T5nax7nvnNdWLAYx5p6oTH233WzX0q4iQhpNd6mXtHrUwe8No2
jArVEutJhPNSwJe/eCzIOKP97YNgFzOWpU+gYMmoklmZgo2osIZjq88iZisVspGu
hTw7ivF2juHDK9BbLBSwUS5M8nZECX8UwGVIDMP25hpcT3mE0TPu2CstX52waQa6
QNWYLmydY39hVSrg3jbac8W81b7+s8rwsARXCdC0dHxNuf7/3Sw+i5A1Lxmt+1/k
QYqTztG3egvPuaCezsUEo1N+3zjQh3NUPv9f3ZbBrB9O5T0UiG95V6OQI2Fd51Co
VK6ePoSJ8SFTFzPjBcfHA23EMtQ/K15mm2fNgHKGjiWRlhXi6yeJ77xyyUAXjZf1
obTS4mJqWsvDYnZoA6Wa6W4aMHDARU1DPCO1C5Mrm95NAOguXeSCxsN2cerE33lu
ue2Q07osFztgkc41luacKrsnfmRST+CE+P01HJZ0IsSiwu3hJdrwv80IcVwMnpqo
Dj1TUG5QHIp2Xuh5h+lVWfCcGNvBRmNtQ8KOD3cWghwXPWUXhyeNmhEBNQOcs9k4
I2sXbgGpSoa/1h1TeFmIb6p8wGVl0ydxGxPn//OQY9HBeZMQnFZ5+dUzSzvapsh0
Jl3Ovo6r2v8toKlwBvZ1K6wMW2SNg8Q/KaRBIYPrw3Ra24RCuz/PExbyEP2bPPJ7
rCSbtw/3+yR4p8psaXvmmEsf5yOcLMRMIiVx/7R/UDcrGy6Pz0b03+lC9d5zJZcY
ZM9Pr3VrpPKfJfJqscYwtw1M4vdBz0KbVuDXhGNx3fl++2hkD9V10m4LX/0DLFjW
l5fy/yc4rZwyzMwICiC7QlX2L/LnMh8C4xMyH0ol4GrkyUV94S/CAnk+9hQwMk43
o8/P8yKFOkNTC4QHlB5kNoM6YeQrg9F/uUG/JaQTEUqg9P3SkiRl5WKgYMXBLstp
NpKjAF7H54jDIZ9x1gsMuuuQtJl3PU9yaImhupfyifgbWuHuv9qTxBfvHa8WGCBw
2YedhxwETpy6XtvNKUJ0cgpaYMI1tZiCU0DdDH1VahoDGGO7BZyYpJE1ZphpYoZf
A/rb/RV3ISDdpDa7bwA5mmwHrZRnWBJzsWMm7nNiUoJupfCibmpqyQYbaDstOfte
13vMaZAkGYOK0YstBKDE1lpRk04K0w2XALj5SgfH9xX27YpBahlZOxBnYn6iimgH
BWcArgvYQWV3/AGd6UYe/TOcMkyJFn9kSIZy8Gi9FXIXEL08tSywu92XOqUiWEY8
+av293O9xbZxiaT2LqL0dLMbT5Fn4tdVMHW/HaBHRHY/nTmingUsi7/fxWdPa8nA
6F8mNQfbdssMl0whXBSbr6R0rE9pOpACdGMddop66o6zyoXBPMLcIjBprZiSmdXz
OWWt+A7jFpjuJPq0f6cV9A+NNbKMjgS4ZnWfCsL3zuBWJpil/HE14Lfb4WZ4U8dj
S0CsUVLRDvuOi8Q2uiKHcLHrVVhw50aIJ2wTrQn6guM4+9iz9GpZbeGhy3+C5/W6
yqQfLa84iwgeqb5Fhdjtmz1zoaVksEmTNKeIxuKmob22ufkysNgletpJ/FAnGaBE
c8IPOMekvmvPudNZOiblJMBiHBnkkiE6JT5TtIzL8RYIK0wE1Jq5IHrWI9z2UGtR
YqK2ZfRu1nmGWOW72Apxl/QtEaYo4XJ6Vl9h1SVnIHirrdsvIhUqbccjOUHDyzWm
MiEhtzEnjnrzk2oh7a9N0BwBVXn0W7K45voZ2czrT2xGqrkeTbH+TJiUpslqOrdP
hu9Q1/2bi8Q5cPqZ1K01M77a19ouzH6hoKY5QBchujRMIloc96QFGphZpLc6jm79
7wDNwVTMIZ/W0XxUuof0/xCp7oAYVH2O52u0oXYFtPjno6+qmIasif5aiPDURkuo
hVGtS7Gs4KSb6jLhMolI79S+SkqJB8aCtQNJBYY19roCJ1JiRE2SfDy/Xk1lAhPa
FLLxnQ8DrbfTCKYXhgbo1lycNEjJ0Z7oB4tck8Vg3D/y3SHgYfiCIotJRAVKiXqC
tbubIYhng32FSDikS1Tva0d6ExMqOSzJFG2SA5Dd2/AyJRl+zS7/aqBurn5JbUjY
sNtVt9RLABbelEm1M0u7VV6jbwnMni3Ipy5QDVXk8/PER0L9bAw0tNVrzW4DVxYH
gmCGGTEjPm2Y5nYIuEMZrBuQYLgTTwV/cZC0dEHjx9y/0SNz6bUcUEHuVmpO6i93
IecLI3MoKxCGKBy7fk/sDXfbZJM0/AYrCVTm64IdH4SlFaGID0n/9c2AHOWU28xt
mKSIKn0dByd5I1i2U6yl/DF4eTwbyF8xOGbfg0PDLgyipBoO/GeLqvSmQeCgQpiO
B5ZmpzKsFp8f3JXBGh0FuIJgLr3MxNsBEf51lyc0tlttP+pXXHATmLQD93xH1I4h
54MLDe5o4ibtTnEsDkYPEHjoX2ioWSlct+r25dyVFJp8gHated1fJvK70enj0w7d
t9Mk5VL1NyIBIgzdKy20RNkb9pb2YhnXYkLKAEC6c3NSXMCygQcRlRNO1TJAKJNj
BJF09cTUNRbYtOG0U9thFqC9LMctysXRqfpnJtPHvSFXZiQuMgw7eVBX940cLGPU
3zjgYKcSAbLz/bvcfqGTU4JfcPsggxs5iQn2A9uSHrxtRUgL11IHHU7WBpya8qFG
9/wm7WD2z/hckATCJJvcHsVTgKTYpKQt64JWxNGHRnIhanguSg8YwkwCihp4Rj7/
Gn1ADXj9+hGd3NFjSwd8pnPECIkdWCnOFhCVmphM6JIjPb4sozWUq2R/BnSNajFn
kLKMRgWKbagL8DyexCZuycgLGuBtUeOXQwpg921eamlwBnj94wBxMBNfHRNW3Rmz
XCbz4VQ7saCKsQsfwNrewYu49BwRbCxpbwdgjh9Gv5F5WTwqmVmeK5C8/i3qjmSW
mnq0P5TQZQflyv47wt1gA8mIExyErnkJ1QRhXUVnYb/1SqUByOaZHGc2mL2dFupt
eXBZdAH8XLROv4QR4iDHEgFBKnb5ED5XzWoPt4LOHmq2SJ6aF5CJsIWEfgYbNWUt
SufHjGzoDfCaeK+iwaNIGm+avo/nJ+I0EApTOY+gPBsdr4xHCZRVMhcbmgSJq033
jm0hMTNU7ow65lUCrGDxNOmijIpY92vhQlPPVIanhosuDqtw/IDqhYgNj1ldKyQK
yKF9ywOBX40MLp1DbHTQwLGv7cgnYqi0q+RcbAXgp1W7xVv+rBfxqWL/hS/TpmDC
guUeAbjhFsL3aO4q/1eV+0OAWsLjKrPKpKGdKYWd3sH0rLSe4r4Rhep5KxDlGbn3
ltkPBvKUDFIeqygA9y030N0FtvXBRBzYAQ4sHQ2FW3MhW8Gheifhf/n6pk+UoBz+
AO9PFUxJpSSlSuHZ0yoFI0WzNySWMvMWvldxxag5YgM7iqtlSz/6bvhZaucGLiDm
RLrwLZU5xaOQI72PKL/L6NomK/THim8oXaK20+nusY7matJlptYXW15N9nsm3JL8
+HOcXL3GSyqnKLTFkUFuZLYbWERmomdS9knwaXhBRb3gHDmVqXMr+rZiC4SDOARp
I6eZVGiSGl0OZ4YZA0IfMwmxpmxaSkNts+FNtQUyPx5gJ6loqyYMHi1Rnm+mtPYp
evW9hg+T7Q0v1EWSCb4uCqTKoDjNJZL7zbq0mC/LQ6rm7AEKROL02lwtK1Wg7yAO
LSazNV1Oghr4z+xBokJoTv/vvdB7auNsDAbt+pXyw7oTCubZ07akx03clINYB113
nHhp92VwwXmjoOV8VS5DQJQiaKq2xrUvI83Do9PMbN1mkHjFqv9H+nNPozoCLrYv
GppQZlXT3HTULSnWmfMC465iECeDnmbSnMc5zl/jdIYAbJK2x+SaVG55oGKkL15Y
rWfGUChkJD4svQW2Qpzjs0vdwEO9TareEHnN5HgYflDczipXypfFXWfVyWVjkSCT
WEf4tEwc9NLHZGEeaxmj0Ji+lNSZ6F8bu05ezgEAr2uVE9PG90Ftb/7wI/OaQI3p
orkjrKv+Wi4wm5Q58GmKZFw6okl8nQVeYjVygtHdk7ypF4SHUkj5OtEQtA/Jlyll
T4t9zKJ2YAT6HB+2edLYSOAxFSxdCUb+nQynNNb617QjqS0R9Aj52AN7MNhcgfkC
MHGbZ4PP/OdkiC2U9LvIeGek4btZY8O9e/C1o1lQ76w9eFUPKjp5tXqxMjjXA3ye
i+PkplMzCMoS2zfnKbqo9uf5pWHwrVyniGrAr0mT67+wSnF+YzEPCkeLvjynzIMx
f3vil+10xQpXseZvhcidAUMNSYVdvRWlmZwO6CGXMNzRs2g3uJ2wXTrrYqeqA2Dx
fOxxqM78eg67+PwDjRZxmO8Y3PeuUGMS5RRNPj9SQKVYQ5t/ebCCOZXzHG34eW8O
2g0FmeGKIS/FdrWEWzOl3XQKZWaHJSnCal4s5O+17EoHbAwGZ8SB4APx3AgD4Q96
qiWdh7egybL5D+UZ6W20o7EWzu8KRuitIxknlQy0gI3T83lfRkXsgNp8i4YWU5Ss
pVZhNcS6D/FQI4C8PDOPHjU0OXV0DWaT/oOXZg6NhnmwWvRjIS7WTz0LZylhZ8Tm
pjOOSpRvH8/TOlg1Yl7WfH/WWfahe6MYvytE9ITaiAOjDVXGe2H6bc4WWBTcoyWt
dcPMnPvbnPF+fu69ZLtXtYAzaC+HRrw3xCQ74MHeWwnxRY/f2qff8cBlbGL3jAKw
t89DB+FD9VYwBFFuVZ1ag/dFRvbUftceQAF2odwpm5sUH6cKdD05oXODKGHu69P0
hwFF1mn6GSLZO6MHiNKeVhuONtLrxnyry3QJRpwOmaZ9ChQtA3G95cZFBqrPCS1n
4giAFOHDQvyLlRB9cTE/+BpxVmiH58PHfCtJ+TtNDRBoNBa6iE11LT6j3og3Fm7X
UJWsl/NoD62annh+qfja936JJLcfQaBRK8rM7EeJJSiy+xuoKTBtH2ESsT9uGsUK
FGYX/mqeVbx0nzGSIgaRE6xIFgXAhGbuNZqXksc+LyniuPqyieCLksi8NBTENbfW
arhO4pXmWOwviMZlelFhzmhIaqtgDMIfBXYUGWoli1qVwx8QCFJQtf3wLGu9F+kk
6wPvad1SUkDF3q0WqZ0FG1P09h0BDQm2iFgUp25pGl5grjrIeUe+VHq9UHa2cdOp
oQPuY8hcshJ3zqkCIh1dgcfE4PPhe25emQ4mmWUxtdpWE38OAZBCHzURLoS8VAe6
VnsuAaQoC9xTne7Q4LjMW09whF0rMBG+wkOHi/1nS0yhKdQz9xI5Qf9FPWoU7y96
/0WNiXWvbb3mu6nxl2kHb+9FkCSRKAO6lLQWwM+jEH3YP7NsXkQnTXdKtqfhnNEU
h3eUC9oAoIJx/5LegJOzKr6idBvU1w6L7HRsCZjnigCJnH6RZjcYWIAypJOxDVG2
paCZUu6/9KMnDmRpzbTOGK+OVTld0jE3oqYbME9AmPHtuEhXkmCgwrEw50zssUf2
mStkt1dVW4eubWEP08yrM918mE6gzIofvBwr2mcsBLTcFpZrth7OLvY6J3lbgNzS
q/h8tHL57xbEDPpafOSmUHM0iGHvPq/5EUaxl+vaaJxPvx+aKNvcDhUlW0LgIUZQ
SAgVmn8LJ0FSrLyOyi9p5cPiaqdtR/UfFr7OZHBWnIPcFq2zMo6Tp4mXxDZr5WfP
SswhuQ152dIAbnvMUbY9puYjlkSbyeoxOtr9iWRWURvMIXnFD+t1k9FA6OrR3Nrl
LX4+A5G/158WdENQ33Db0OiytDu61feKCEbAwtdHguEuitBKz7swrv7KggDwWocg
qBozY6yOPqfwpgJDFmQWrrpobY748mgqwiZNNg2dihlU1IQqYJSdjHG7RLfpG8jp
548XiakWCYNrTUu1sc0kC+T/hcBCCoSQ48xS0Lv5DDnJTaneQIf2mvTBJH2D0y8F
RKtxFWCIymqJ125geI0qbYvyiPdBEClXFhLmA+I/TmWIVmY6qDZmvW4OvmDaUAtG
EcyFM40hC02tIt1KbF0y9hgnS/0lrcA6cmLRrbu9Q8Fgxwm8gfgCcETvgv0Qa15c
JrGhp8yHIBHZz9e/HEWrctNHM6jTiZsn77RiPtBS19blzfbeRhIzBWUoPm0OBhrL
Lm5/Q9H2lDxRKVkcznNCS+VX9q+IuDdINmX5CRd7g57CbOnaSCBYxljqEyaHh27P
5aMYeGj2EaLiMJg26tygIfcgN4Jv+y3ptZpCQqgvnlS2QKBBg/zE+GhSDZyMlAXF
nX34YugpMznI6qCvfg0zftZGd0+Uq9YkcyMAVA1ZqnHr9i/7o/Mu26KS6PulYizn
iXqaB/K0ocRid9SScx5cXjMeT97BXf1hb34M7C3a1GrnbTTvta7fltoTPzNanQHK
BzbgX77FEBDkQ6mL2mNR7gI8yAtpkorJBu/YKVJ2OOCLgtOZrycIW7ckHAp7FIYP
WnNPzfXUsaDiBcLEtB7sz15GFQxllHbijp3YjspX0zYXHcgoRQlbx5I6EdcL4edP
TWx23U7RqvuZDCFaUo8nTvliFlz5kRD0WOj0HdHGsOezaocTizwfm/Npmq/js5an
E+r9d2Ori3RAX3Y700vlpqCxIRu2YHQswxSHHdz/qfzLLsTqhNzfnAWZemNr16+w
Apy4UBicowellSLKILxPCnqcdoQtWwoUe0nLEjFJ+xbipVjQ0xPtUNnxKIJSczKc
dNA2mUBGR2QCZ3EKAnBdEjAtGBW8ZiXROKIalRXDB0oAAFyO0hVoG1kR3Jmo8C20
+46GWTHjEAwe3NnEvK6cCBN4zULtWko3IaSlTr8P6rhGT5LPkUyqktglprJuLSAt
SgD8qcr29iykHC+lOYo3lkq+KHJaUkLus7Fiaodu87b1CG88cnnULEJaMaecU+7d
TW5MNNQ+Z4ImUtauEI+tsm2/dXARIqvY8QhkF1GEX6PVzY0prfW5ciC654pZ+uuH
1zW/n6N4MvPA7JpUUi4gNvdz+BsvEMUR+ENUQgL+vqIRESRIYPlHRMO29gHBvR6T
BS2e3Fi2LRsS0YtXQMFqroI9s5+ytYRoSoJhCGYP57S4+JAFx5iP+gez/xu0wH1r
ofSHG/oQIBIQ32uQEFwR04gJPwj7ko6VARzt5RlJDxuT1rnGiw2RNlMHMp2ki3wD
L2HcdNnUpsQ1rEaPauUFp9FKP47fWa+lv7DzDBscB+mY//tysvRiyE5YcH14xyGi
yRy/7TGSPzHEqIUiIvWmCjLBAdWiu1G5/4tiLjBehPI4iVageaTq6mqWADZSWbDg
yWtF+m3I0j2kmuEjO/2Vkuk3fxGI9B/n9adypYJRf3ukilj1tA1XpPqQueojUSaI
NfiFtemN7Py1rPTTIjlLltHYCUI57iWtUm7FFOBTphQcD3+rtpTpTFRqBuNslbyt
UJ1BMS1++Fv8B89dAQglZhTvMwo/RWA/lqRfgKCzgq0b7Vh9LmQIApkQNlnmeNcG
X8bqrm9MLRmHLLJIydT9a+haVvDQSUTTZRWM+svWmiWDmKzgYmSEVfNShPEZHRBW
t2SSFXj9KOhwr+5zlkbsz+uHj/PvdvrOEPMtcYCTfNY4szMlraNpne+nwLmgHIbo
7ctZwtnuqPQhyum4p1Km5eiM6wnS6avFdWmfBzlvwJfwUdcv0Yh039Y6yufnapw/
ocILx13/DNkU44j8sVAqZI9X/xfrsWO5hOMCEsu2ftQK3h3vA9H62MLA6Tt7eoV9
k63lzPAha1BU1cGc14AUV3ru2bYPdetT2GyRGYj4iBX/aHXuSHjbC7wo//c8zy9z
leewFoySO5yZISBLgFzjs6RnRstAbNdeGTFkWUCxzOqLe2Ho9vCFlIqrp9cqe6uP
zBIssMAMkzICjGpxA+BAWJoWCCiWXzbDuaL4DG4aUINzusSFwL2D5cpTnXzbCDBH
j4jxGQ660uKUbY0dP/uOrCHGN3aOfMVnTQ5Ky//uXHZuyybp+JfJR116Lz+FfzTI
NZN9k1K/A5WXGhSvAe+Q5Bu8GG+C7KJwnAgky8erCPV+D4xA0Rgjsahgo3H9ioYy
ZrVtoCcJG7dCPLZ7Zm4Ut/xVArR/iuGp7jsd2n7I7TAJ4Yff9Czr+9ES8foSVpVa
79bwhaYYwgdIKmT5YElBOS2NjScbAxeiDxganAVtDoqnxxuZ8JJG7w/JQlcDSocZ
XaFxQpUEZJzTbJfkdsLv0GkOx36hSFo/DKzi98GRhw7QGYG78ASBYvVL0FAp7zgd
pa4lbUx+7444Z9Y8+Du1pmF3C2aCPFAXm4s2UZReorDev4hHv4y27p6HVgOXFCLP
1hnJgkhouz20k8iinlXH4w5TxZznOj38dvfLN0tdD6h1wXjQoL/czzAouA97FrJ8
UaVRiuXYqx9E0P9LVjgblrwFxNTzLoZeoFdMIy058CiehgKOxK34lpXL3+NPTPn+
OMnh/yMjs2yAA+/Tf/o6WIn9gTPkMBYXiAv6b35Md2eU785NaYcDBDtPs670raPB
2Ux9WFyiFxHukFuw4pkOtzJMaUVpNbnc3HLKs2BFMXqYVEzYDjzHu3fMX3wrqbtL
zOIlT8bK1fePGra0/OQt/IyJ8k5KESR0efspOgv2EXYGFtT41mrVcfjK3gSLXSjr
8948Cg0LKUh1iqc5HcD2A2RGIk9nEBsXZNbk4lOLRLqyG4IxU5b9mMiD19V+7wyL
h/XLrrNbdxquFrXw0mgHo/a2mBbdy/RnD+hyjokRlm2H1lOItz760M997TsF19l6
h+gL8rvBoH+QE/UmMGoFj82fkBgD36WGzLpGNjIaKpkfICUK8B2g0Zn4XDsnATzj
4cEPWvDYa+E22kSotx2KZ5SYxL+OhQjySbcHhXD813E5TIIKoyK7ZIUaTK8Rsr9N
fJSosb56fArRtoirDet03pG6CZQ6p+lKp/xDDVrmV8TQCDsIxuvuVq19UztpVl/E
ncZjUNeGERqd6qhoU0MObgm1Uw57b9ZztXu1nMHzkpa2PL5koVl/hnheso+6cEs3
Kt0bAohuBvhwV0sL1uD8stVbWv+NpwA299I36B6QpHMWoOEMJUMgjMg/gufS7jYh
VvdAo9ifS3P65Z3iduYFsgNlw76N7YfxzIHC1Or7TOZcNJjCJrVXswt8k9cAABK3
Lnyd7v2qYhK5LVdfFNYGyRXkHrUnpfQv58ETM07d1JMgQNggwecv1jihlNg643oU
gDNBKLMzg6lp6RxlmEIURPF/VqJ8KVaRLLk5BZ8R2EQ677+RwvJTjtF9EZFpNrCK
ob6naxrIqWuaMoDlxjwadackeNZfKdggu0CHSd0DLVCrAERkPfpCXBmChs8kQUEG
NwOK5ZcVz7V8ufjZvXP6o/J72HvOi2d4wia4S9fVav571J20qAutjPIhunDaUFMd
YoDUrjknkGD7h/JJDpKWUJLvOHNDfa9IxWPAFL3xnJn4773id6dETt47gkKu82Vn
jX3qornKKv8tzLn8A5R/KBNGqLqcdHnHf+XmNulHbhqPXhR+GL2cyn2ykXLODI5y
FG/xt05SWZ249xfzaQ2Cfqqz/ICudRKeDzVJsUYfGFhcnfGT4LZDAUfJELtrSMV7
6dy5mpBuh1osWw+/pYi/uhPSn5upnJc607PVxXy20OKsgnwKoQN3AwUnmNcVfXwq
Pnb2CiaixLe5HghjT8FCOrDxuGEEhXZdpzp6QqMROC05gbkWye+N2VvVgdnmsVgQ
K9pD3Zt7kZVmyGRtDbH2LPnOK9BKMIEODadXAUUGerpIottrbBtcREG1Vz8LlOVI
KN5QhRurpctQoMyaRnM7YCwtDy7xrg0Z5s7JGG0t1RMBWSmHVef7D6X+2Lk6zpch
3LwTXkE0R7QDsgDro5dfWwegcQPeTGDgwsl2jjvjCBd4lbXlqDFpFVsUzfK9P2eg
K6yuYjLSG1tr80xLlZ3hIwB55dj9aCXCRT5zHxVL6IoV0CO1r1vsrmPjrfAPOEod
yiExREsv9Uffs5/DxNz32Oop2/uEoL21J9dyl/9bGv2Fl2Rm6eGyQqT4zk3omsfH
i6O/ut+dHVxOztTMX1jqCdjiUYaQeTkaoMH/FBVw9BOeoNYjAnawWZxguIoy0Elq
SQaUQn546m/lOwII9DwLGqYphPI48dIoZr8TB5jRTWYY0tG3Xa9v8JFTg+ijP+Mz
x13KExCyAJUXLFvGWOhT0ZcfCCZkI16PQFzXwKNyfDQ9jxAENIoxgiab5cxfyXUu
HuQB33sCMreBNx5InYXiEfrf32CBusZf5uvARFrvfMUt/7MR7QY7w5Kkw7ZMc3Bo
2AskW9cCPl1OE9V6S+IIjsUT+MHvolpfkS1UVrpR/8G7yLF26aJe6Voxc/rlxm2e
otjEiAiB86TBbbYIjZiTomHcHuypAhZCBel9+bBKzN5S66b6iYoJff1PxL3+Xe23
Wz+MCrufg6vCMEj7RZFJJeizTEUeVzzteysuRwcOZJCqEeFOcUJ6ou1geHKNibQI
GfbOYidiz+5UvBbkThaUtvo0AO3XrZ5Zmy9BZYiOVLYKVPVJnFePCtP8frSmAB0j
sqwRnoaIyfF7sIKUAzqJopZNdvoxa015htvxiA+CxWRMDYgxarj2DwcLqJ6KCYlx
NcEQ/O2nHwwmji4anaU+i0mnl8XdyjXApqhwQk90CiB0ewVwNPvXn8ZbmLjN554w
FYA9bUiBwBezpEVKhZVz+TEZaOPbW+ZDKfz3X1viYBLTvWKLBSbwOhtve6SqoM0t
unertBOeh9kLcpZ8jBm80EQEkEBK+i0cgfMlu4VWbxfeQyyYSLZNx4r2JbiSQysW
cQIFzjJQ1W0qQeqrNbrH8MYRYAFUBZ93E58LuLCFEls1s1yXPCtFzdyG0krsWcG8
mmyBUObSAoedrybmLVrRh4XWgGFJ2Vo8kQfg0ZRvts3js9ttlH82ETDhhSAOgCJ+
JxEIhJjrLZC/B3ZYrDLrk0Ajk/v4Pwj8teTg0jYFmZRjW+b4Rvpo8EhC0jBnsB5R
zF5VYNeMVcMeWqkns20DXSf8mnTXwErIs+AjUyl5tP6hMizfm4Clj9hVXfknRKz5
I/mwKkJJ+N+ZMj3RtvjYGU0fCRHqv000api3Z7dk3GzPhSRNmpKIOqX3/DWwwSFW
wrnGmNl+1yAn1F1M0axP4cEJWRxs2tKmW/LM7idue/m9mKXB9LX70IYKn5hP/6Bm
AXhaqsKfDZuIusJYA6huTQmIynx8N7f2jAu6e6XkEM3UQCT3PhZeLJcBoQ+BhgS7
qftJHqfNfLAidG6FkIny8by13pzWqNQIJQm/GnjDOR0178BByEhNiU8fBl1KdnAX
6D+TFtfX09QNwIQCIZ3o4N2Q64zpkMqwpqLG+0F8N46JjVPDxCQoVPfxvyRHV8Ha
YfhrgZHENttxLFi1ep9RC0w2/TgW8F/yIS2fgUcvKNoe/y/m+fcbjEJyfNZkW8cE
vf9MYf7sYozzGw1H0Bw8pvr22wNw1u4EYzfud3CMd+ISmPiMe1FBRdigCsOXGlSd
7P5hle9ypG/RgaByK+rfIYt+DM36936hH5FQQIWvJ71PAZXi0xGxgqpcS/3nJ5/h
xpT8fxeg/HWx58CuYHEoTN7DhG3Md0tTjGg4g59pRfOTNNb4dm6Lx8JK4pOjw+ni
WFafP52f70a8T2a0azJ4KwUOm5TaYQwqFOfUTTz/YLLenpGjilumLOziFNWaLtCJ
qqxMl+0D9C1P3Iqw+l/Yc8eJuyr2OeXUsn+nHQoHNi3YQO7gfQv7nKE/sS60GllF
5vU9eOpA9UvW+rcXRlhd/RLjmde8pEbIwwyF2YE16PWQJ+EjtnBbq2UNMS/KvZCf
Ke3q4aSYfkvEJ6C1eKn6YekOPP0WwUmx7sW3qwyV4IiZn37HYZD7m5VqxtIxsdHH
YkRDVhw3mQ+XbV/EUpG23f20EGOxjHNiq6kGhLvLqOevPmQEkqXddcsV3Rwj6LuN
HAeg9WKv74Dm6+fNXxldIEpJFfoSpq2+1N3K4+FIVLp4JZZQH9oPIeDg52jKWi+H
NF7gFK+Py1bKX+DH6oqR6mSUmK0TZkDEBB9C1ddqxO89BUBCwvjRQK63bsu3n1Lf
uSCLdiJQgiV9t24zLFOdH80+vD0U3qzKiMj9hjQdnTTMXhqLiZ2EVd6GndRb/RlV
nZpL6U2/jR85FraHAKhPBUtAZuFaCoJe5pxIrAww3U+LEr8GfLXV8lO2t4KdKyUJ
UnYxlVBWOK6g3SShCmgGSPoAAvtyuOgIofvKPoVbAB2BR9jR4IMh/boQKFfb8PFv
fJIuhXGSdphz169rm6uO7SKVMkChGYrp7B/mbSyQKeCCdwWW8S5q+N2LnlIptBf2
KTV1Ig7//l3F5c2kmMCcgaiLzeoxNO9F1qH/CQGlDsxfNdfHkCFD9o8LjqquQ2uA
jv1f6xxbQhnMSewzjL3mV8lH4xJ9KpRg1ASsQnw9SVqUMrEi1F2r1jzou2FRLldr
+hUzh9twCz0HnNOFk1VcED0m79Yg0ArDttaQ+JmVbelLazNmDcVeTcXZg3afscVz
KhqSybto0exnN015SpB2/gvTq2gm7oTrO+TLU+t0oAMSRceY/Gwcuu6UvEoQoIjK
WfJwQDdRIMRyPxDTVzMFg4GJqucXWEyMOsWR+i2NhLzV5TsE3rhdcLHJoUMuf8yS
qAyZaa2/xa/3iCpATe5f4sPoLzbotB3M+13BSheMZqzg8ZlqLO1695CxlAGn+Uh8
6emGRZHfR1X/jrSP6HvuK87/bfmFFJqQHEAOLbufrUUY5+L8qO62NwLGEBUEaHT0
doFJ1Bik3N+PvMNrS24nLoIy2WwtLQ+AcpCimrIIrcFlrmW32LwjHuyEq7pYIMHL
ZN1n83gAa1J0QQp7g3nyD8J3rvMoAU/ngmikv0iSeJwaNFGC4BgmkSd4bP5W+Sof
6FNXBuly50BJDcEmN/6v0654F1Lyn8r6AmXljjW5Mo4tb95eaJLSAOOyt6aZ3XDe
NmFVXf+qkgalOInrdKRg1QVCvB532NjlukCiqfNiOEvjM7lmwMikT1HURDEMVx3a
FQc3B/m8F2DPFPyP2mje1yWyjLNsk/ysYFQJKygpHqPCpC/TNOtec7nTCxj99MWR
MAndC97AnnHlCve3vscIPp8lTVylO5YP4LCickWhyfhhmhGt9YSkGZxP4ocK/I+y
1DVSpEUiqgrD2+GaXsLq/Dz2NjLY1YiRcCSe3AwdxA/r0K4qJS0nKB/HWNkPJNVb
Aq8bk3k9Dw6Z7ZKwwdog0x98+j7C7Zt/rZpSwMBDNxiDPdrAmd3zIv067p7Tj1H4
emY72RR7HTKnzJMgMY25V16BJB7mxaryVOEk4xcNj6q4RjNbjt2X8jk2scY8fJsN
ijoWGM0Swm43DtT/MgvsVBZkKQyNWtCe7PZSn8vTvBr4w9jJzy9Mh+lQqD3JP6t/
FVaZfa9kFIt0UXznsR7yAqBn9Ofx3S9QY+pqNW76eCRjjMuAGe9IoHhUucRY0acd
LmJiVnhD78rIhIDd0hBujt5DlD3JIduPTxUHuWmCSnwnXzu7Tuvvq399ImgDPItT
1Y7Iu9cfvyobMigAIzQ35REysS53kGTk7WxvutiEp6Cjv5FbLs6+852TSnNIWg5B
c8LorQfofV3dmr2Y2JxwkhCg4u4xKzpwgnzrfMYw2WyLXqWhGtAZWUaVC4/AjFUl
IPuhXQULP9esymhz8taTNWG0z9fIDClClUqysV6rLmDUGJNuoCglP+eSJbji7vwY
rQ/cXlbeThByxnWmFbI5q40DcMWaLdrhkOYqSWOa5gGeY23K+pSKJQuvrdOvb1iA
1WZrbeY6xJTlKDO5kDZlNVZzLaJ6oT219sczhfRnWcz5wzyCn1KL6Wb38OzKynNh
USKyyVbELNGlM0MWKr1xB4ba4v6jrFlOq+REGSpyAU9Ry9tBwUYGtr8k/v5+nF1V
SGoLCWKf90dw9QLkkopEh4/gJKTcsHog4d2MHp1JvCSpEG91RecNklew6e08ZsQS
07fNyW1djZjvCG9PdxZ/24i3+w8cX7SaTyPI1Lp3Jv7HuVtgI0AIjbTB76hHZzh/
v8B7FY0qzH9IK3+cMWLrWzcK7R/gLkrFsHiGtu4CPtYiMiuyAFZKGPN7WhICaLqL
GrlmbALl9naApbu8FEvAbgKi5wNOyr7UYij/rU3llGKegGsWlV9Pww234ICZ8PsP
SQR8/DXDyTTE4HViYaDCtH6LbXvwLa0zQm2sjWIFzgyy47I1/d24TdUJaupFxI7p
bl+VR7JzV4Gw01rKqWtm1Ovgaq2/A+tT+bQMdDZyESUAwsOeJV+jhruQOmKvJX9t
OJBEw6yqE0Jq1cfWxXP3N64iZcPtxBMW3TseltvaOvJ4CwzFWqQOLAlTM/hPydvJ
qUzldTK/Vxmkg2PD7H+MRtiRFpgYRlN0SGreK4tO1WWvnEtAF9WSUFpn8/USyzOt
L7ageGE1eiIB/I/iZS/YiNoRvX5yjIiorob3shTKbuh+Kv/7Qr5hoMu/QXT5FOn6
5h2pdKkDzr4DBU0Qb8Ec2U8k/gfG9X3eYDkEPCevgnJj1+Vy85I0Ag4gZsgG6fPB
zJmXXuNAGu7Ma1mBe8wbW0ZGX2Ff00aZdGhzRviPgCNjvBuZMWEESszxHDPvG2eg
/bgd6vIZKl48VBz+9Pu5XXjt5re2AnYWRRD4zVfIcH1kkwoa01cqVt+Np9oHzyjr
ZB+GHnj7jqiPo0CvHKIOSdrxL/Ymhqa4d8qLIKHvr/wlpLSgfb/SyNWzHxa3GhvD
fcQ5rkGF0ShhaMFbgNU1nwCsY5ng8/KrtINbix0D5nL9yhVU1NesXCs4xD+l/P/y
KHEfYUIbitWi+aXSAhWzpWQy06yyFZP5S4Co592UzDz6jsh8HCiAH4/6hkNrRxfb
Wl5j6zmvCcQBIZA/Y2Kmaekyyqf05SVf24x+/I4WQaqkV+TDiu1sihUczddE62kc
4kyOymm1rgBGhNPRqg9kT9KwBPEV/gZyK1u9V5o/kyZa++FJsWuO1k6xk/GOv3+v
ppJZyPaUNlBJo5CTkgDDg6iazGS4syTcRBbKhI0zwGZ4QecgCiv52B3E2RU5bD2r
Ud4DcKevPJuqNQ+OUUxNuPzzcibk6mDFuVbZALBdYw2ta64pY5ttIGBtZHLHzwsM
hBc3Lvmz0zPBN9gpACumwFIIaajD/YUHZoycXuM9TrDTF9/VO1cDw3F9ewxC3zgW
Y9pCWfoOR+vwS1EUSSEHj8AJEgnYk1jI7Teoc9nfHPEziilmjcEyCjIv5EfLD9Ez
hV7e0mCC24CMauA/Y/AyQz2oHw/YhHEf3GpAUK7nehfnPmHc3ZTzqymvMzqyELUr
B9EVXkdvnugLM6CDA8ko9hJq5oka9rrem6irVpae0upKusy/TckSL2m4y5OhxKoH
1Pzb0r88pSF8jeS/CdMEqN8jPlQZZWZSZmRQqh2dY84lx8xBOtYsFTT7abrQlGX7
0aEP4dnrxthXOpLNSVhmks7LtqtNE8CqEVxlYAXBCrF1ctWfa//ogFz2Rmk1KCGV
jl3SrpjvzUUMjQZEfLmzGzprViV+PE6Rv7jF6P+RO16eOwXjP/B7uRiI0pDTIe9f
emwywinCCzm1X4mQXMHrsp3oNh98XnMDJfWNB1vuGLkND+29tUOt8m8wtiFMnK9k
lcDxPrEzxFZ+hukEySazbJCwPC2Pzcf1dRCxP+JAhPmAhcMsarA1e3+A4ciXA4EC
uB0bXRETWfAtuOXZtilOXWwbcYamuVQIFZT7ajonOgTJvgaSVKvmi3s2E5fXwwQM
Po028z689pD/IDXkWcUR5ID0HF0/bKBwDDsKzyyv4psT5fiioMBLbfD4pVlo6ajl
oxajIJazEf6npIO/OURDbfoutuMSSBUOFzaZcgnrNr8ht+WaxR4UOz03gRAO9B7z
MfCp+vJ9lO1/IjKm9fF2rSmWdHcnyBv65bkw7yF3LrRXFhuV4Hu4v3A5kzEry6gG
gQBDgXseOZ78PbaK/PLIX36F6uS6tgF9DcIHfoe0EfjT9SLqYiD8M6kCKNu5gtpt
LnjUtPVggZ7M/sWHJn3KujQUTCKq5ynZ0qhAgFvJCTvuvln1SqFXPQIaC10HSdZ5
69a2LAxxQpe0bE9hrfMuuVkZPwpfe3VcUvzMi+BXVJIR4y0p+9Mtur8RgND9hyiF
Y5KRRUA84iTQMpPVAQ7YAOCQWMKfA+bZApfQ89r+g5KtK8mMKlHUhBHCvDysbgrW
RnmokTVdKkGXfwD6n7Zos2HSpHnRRsVSEWdOVYh5e2jFhpGjheECH7QJoiuvBq/f
jFvjK1nprOdykha4s9J5+8Xd+Zj183AzejfQ72eGDgstPZewFtnjV7pP+YiJ1knh
cvQWsxCEzAP7Q2+ynk8Oz5N9nIaXWxcW0SH9Mal5QQQnpGmkFnUj4Z3/f9ttgPXh
2uRNkPEQfYb/GEAGgo2RqvyRSgo+1J8IeEWEkDdc5iCmSpfkFzevNOIZDJawg2xc
SNu5q9Kt4r2OIAmb0XgwLjRdBBM5ARHNyRE+Wh/D5QmvFJwwNugH+BO92sz3/bU3
pHXNVB+cKuSfifTvMm9a6bKMG4cGuYZ3cK30zZy5LizfLKqdEViYTpxtyBbvDRf6
X2ZCedF5cVtTm/WhNZGQBEsVjBE76ww4T6pYPsOnNbQIt85nXkROJwpeqx6hRY52
AU1H1bQin0OnkwMkeXnb+eK7/DuAWRlIsN8rQdURnY7xXR9OzIW6sDO/ntCyzySN
IxXlcwmuBDqm6ccFnkAiaHE/B0xdlanXveuw65/AOIDklj666DvNXQFvuXzqteMj
kkrtukEiOar5pCRCooLGNAm8EEjVThwpGzg6ze3iHnTXVOhkUUXVK6Qg9PbGvBsM
pjk/8bmNrlDw3YNK/tVCFAGq7eK9vcT019ywrukzx5L3jyMBKZOvc9txyN6ivj+6
fp+HtbZaMXp2SFimX0n6it52NWe6Gfhc9dHezmLrrJmwZan+tiZSQqmGU0gHQIbF
mcXwoHHFGbw9YDmynVaAwslfpGi3AAlwMxL4xfjq2YK16nNpSz9rscnZxAhIyL/s
jWVxa8Kl+f3ePnwqRiHCxSupei5vWzdysq/MN3wwaiDP23ss6CFqm84n79GQUitb
PGkw7K2kmiEgJfb8ym3Z702LZdVtouA3/iF9/WSREkaO70ixkxqCHDGY2tRbIoPk
dQWhD63WNluRJMuTX+4ujrE/fdh9T6/tiptTx6bJa/EngKIbvqRLXcW5MlXQLCPD
yvlSvim5J12OodIRLnjyYtLXXOzZGHuSO5lE6gTFzr5ujr66Dvv0rWZ4bXRKSRbo
9UrDXx/B+NYBpBnpeJErUmHOjT2pJ8CmkMPXPlYlrTPLCsgpPE+nm4Hs8KtbqI3E
SfswazMUpfr4WCO4y0wt2U7+sSeEbJyOJKtN4MShCp57t7Kb3bhVv/IzxbEoxIDa
E3cmOlo93dbXaMlh27LBrWZ/kso9zywjHJD68JamlHKLlnYUdWzCJ74EIxeHrY2R
+mmb4HCMPBv/kzs4N4Bf82Dmn5+86zYdhpNkq8YUkRsGtEtwvN/FU/NdPhqWIfZ/
JCz9PMQrRTqTg8sKEgQgQOjP659i+wnfo19jZrRavtEbQeFwIKR29DyWeqOioMn3
MTI0Q02vCxPlPdfOeZZ+D2itsre1SX4S9/B08tpI4Lx5QrCBWVE2p0+X5tjoelZw
8LMj8SrKhJlNVRJDhXa0LHFzNtZJukrjwxPw6frwrMkFPS/2tGWhPqMuv452uXAC
WA3Zyx5D1uPUtH5qD1oXGBaCZVqDrWA5xGb681TM1KZyAVbJPyHKl+ZdjvLvdzOh
C+UAuU1WYa5GgYBKKjkkulngBy431xP5lfn3kh+znlGIGQzRau1s/dt2lFPOjDva
86rtNcShlMjcus0k+OhxlE7fvYyexiro8h6n/LkEFqLSm4Z/5Q3Z+fi61wmDZSN6
sI77IbXN0drUrDoE3haxSEbDXNp16rAOUxEbx+s6rqCaMPLi+VuYrcfmPmNEK5N5
sj/ekPXp/EDj2d6LVjyC2hLOJQX8NZ2oTcJjBojm8ovyr0IlOMNn5mPunVLQL6w8
AtwC0WJRE4Nfi8nJYG+NdR/6rDE/QItolYWlZ6ixrv6WyE5Isnr7fMsHH38kEzy/
4BWCgKtr5+KNVmIYY7wsCgALi36TpOXxK49VrzCnD+aar3CutUb3DAMG5OcD4V+a
Exx0BQiDauu2yWs3vTWCCb5ICWHiPdW31QcufUbnDRByBtMQI+YP07BTALXPFgrC
g0gwAjRTI2GxTWheAyD2tBlovvsbyMSCMcQj9ZIuHc5PSB062K89YpTPHA0SFvku
WhK/sPJwXxdBag5xDEj8fp/rgDjn9OG78hAY7aY24ekV5wfi/jL8/qQqb7gDJdOX
aulHkcau+nL8ywgBRAWefQ2kgyH4OFm82sjryP8g7M2B7PeGaNTzaDJPpcOpUM08
WJA0tP8ltjY/26IeEyjfTICNrg7+k+TmlIQuowrovgelrIDHTUcqiCMyMLxzHp4v
RUb4sO+8Cy0xUdqpPNieQitn2el8R9QWyCPpmeBMaVVD266Qqcz/vMKm8jAIfF73
BTbUNj9Ae4gfYL+HgMxI4Z5alXdst7tumnNeiC89p/qhpwdBaDi2x6v0ksev7jIf
XpRj7edRCmLrNCEtKSGUhC98ej92RExKwsHNA9pz+E9t9kGYbP2hiS9GlhjmDgpL
Cbjun7Hq+6v0gHfWSnZxCf0Xh7PNca/lbAE46oYZrN40gLb7dpwWEL3QJFrAyMWd
7FGyAfjLZdtY856HGWtbZVKpmv+L4F9VnTwvJusLpinvNVE3+2MUsPWB7JyUP3og
97yk1wsEMAqjuAkZWMAhkL2wgNFtjq7r88ZWC6jdP7de5pGz/goMRNl7Oo+X629I
jlg+mhhF68fKm52sChZtAJeHwQYrVSCmpcO0bVTz6sTQiQpcL9aTX6QdaukEBZDM
z9gBZZtnZjLKNfQljYeA3bHwXqUuaSu2qe1ewobXtAzIF+bW/2L6rnkG5h/Ur79u
Oo2npDzEpElEStOQpfR1PxHXb3NAPoCX+BvgbNNxtLS7+tijCYBlQuMECII56QIe
hVPFlv5C4AdISPJrq+Wq+qbCF0PyWYOS4px1RORKVVX9+KQ0TdByZQCTOFXiMPfg
YRRC0f6MxTn0KkrxhN4AFPrTnCNAxZkSembJL6UfIvPRWw79KF5kDcKt0sOCx18I
28SD1/NC+M9ILVOuud12ieFWIe7rUe17b18GycHtKSn3hw2cxPq5v389ZlPmWeQb
0vefCbkQJndzfs1keqHPrqdSoNRjjZifMU7kdybeiP42LsuFWYTh1r9/5vFbbNR4
psr+d8zO6MWgzFScM/knW5DY2QbKPRBcFdMbyKgpvUAbj4KaivtKBR5yzBT5SxSQ
bzwrtvj51aZsx5MSclBXIncn3ZXfXpWGXsBEgQFNQiTuS5qzr71AYAAdZOce56Ah
gsk+351IKKOiaFbGwV7uLmS2KiJycZKxtWc3zZ6t03sZhnQ5bauedG2bfCqqCyxb
B6gfFxO0YEifEBlSvmOcIiyaQNj1yoQQ5BBzbfMPWZIAxYmtodT60V9y5bFGn8oH
WVPjE02HKv5mHR7QyHW5IqIBqQxWvFrQlkBMtmjSBTMBSb2m+EM/EYtw+crEoWf0
Bl45HQ8mkkzu8jakzLqHdKXb/bs8fjRfH27LnI8fH2tT5j05Da+FOI0GH9XyJvFG
dTLtQPdXHi6PKf46eq3F41ecXhsOHVRyQyYhk/2kyXqAyA6YEJJc4IzOG9x4A3jT
VxPYqpYJ3dVTEVO71AqP8f6hGsd0BUNo59HkDnb0iEwAYM9qBkdaxAxpuoGfEJnZ
bf9Prb92AfGhyIx7bTwpi1SHjjiZ4XZ+raf5RMMrrMKsbejsSfCbEGygwBKGn2u7
Y5zD3LBgdBYtJ7mlCIEaVsbiRmoPcz4Q3mAVWFr/4gWNtjXMjyYCcyfXMBx9V/Qx
Sn1malWIUedL74gUq0EfDgKa1VbfCwGgMB94eq1Ju9QIg+ufESjOiygN1Hi3yrBu
KlrHnmWv0lFIDMKa3UAApP6eTpoIlFAH14gggs4i6NEfBvDDJe6bbawM1XWfUO2F
J0qPwSwmzspRilIO2ZHPxJDE4vEUA9aTOWqj7qDmaOVLLfo2qSiKJ2bQWqnrNtUB
oG8K/Gw+9d06f7gk2LFnGIISpFHPo4/q16Y5Xd45Dd2eROa7/BLOqm5L4r5V9Q5x
ZT0FAzCKsQ7O4N1lm/SNokW5iyi+ECO9aNUUeKu7CM/TwkqeubMvdUS/HmS39ruX
oJMGrwrzzpqYrxVbYxSCyjYujaai8l6EGONS4YRgNkKW5ctk+GbN2DDnK75WBv+q
zv5i5ok5Sey5E0nOSl80YAgHJYLY4mfNMOTw7mYN2ABR3JiApfmOeH1NJ6OJym+7
HTrhJkaiVraep2HxpzHmD8dn1/cLUb5D2EPyTEQMSbd0T3zvA8g9tdzFnQGB7OAl
a0CzrcyPEipbCouhWaPg3Sjo7cqLJz10H/DHFVoMrUiTFXAkE86Gpaaj9VCg+NTm
iZ3ilEUaVsXNhj5zm3YGBBTu1njHzH5imJdbjlTTtBreGSRl0uDgycuSpY121YKK
vWExeSXZiYaQGL8GdLG+AnPCq+M2NRLf6vqZI7/rdjQKoOaUIZzsU800Blnjhnbi
2rv7Zb/1tbiqjW/FRzMJuL9qPBP7Dewi0r9Q7hvVNidum/0sImtz31j/RuhKUUoe
ELgGTYSuweZswJ71OLLFgG/dV2/GUtVkAggog1xFdBAX7yimnfn8spcn0IaZl5bi
OH19kuuAGvT1qeekNbpMhMgzTe7CNOVBzF8K6cQnfyiMz+f/+/ibf4mLAL6nygqo
+2xxF2h5rP9Ous1pJaaCi0EDY8qqQ8CP1Z8w5lQARQrons2/tLK5SLwuMWArXJue
oq2jy9Z26+Cv1ZWNlYYzF2LkI8C25Qcou4De+PFJ6U0ZG5jnN2ppTG89kdaIbpUu
lc/xJl90iKh+msYdlJLPOmg6zJhiYxKnMzNtO5ifH1mAcOuDC6KP3XwDWWkt9bqx
HlnU6DnPYgiIQ+dJ8RFBVWU/+8g6p6coqDNR9ZGfkn6y1Xy4/KkSqo5a/dzLL1Du
E0LVDgAY/rVq8K4TpPPQmUjTEVO9QLizUiKiGcFqQYLB071cOH66waN3aUzCq9gX
a9fl8RK4Z/0KHGBCz2GQrbBN0wnj4GwuRpuyaL/K/2ehsPaiWqh3Pbz7ZiVyhyYn
jlBal9nfRqAXuGMB+F/8HHxQmtzucc/NmQ7t6nA1gQ4rmLtjrdVaZFp1tNPhI2IL
volR9w3Qcny+6tVFtxO57+cG/UdNrIvGAxRz+ykW3d2i0/pMqVrdhjuYccJpjvBp
QWXiDTbzGFkCu3UFORLM1UilG3vBAaP2IyvUPRa6o4PBTYMtmTH7u3e8XwxLqfiD
2wYoKp8ufbJfpLVCZzQKvdy3tu8DiF5rbGRrdxVx+7radpCSnVdAbB9Okhflb6eR
Qo6wSjqSqmWTa61Q/FFEmLJPMCIpgylS56fBrcnl5KnI0ZOPbrUqzYz9AWH5KEPH
j2IrYgNOZdCrFCWBc2rNItKbESiWGwInYhk5HVUj2TnxZ/9tp4cYVYtsw9hP9sgB
RneivkemSW4JkKlfmN3xvq/o5T6TCzunV3FWwKUWGOYLRLLHFhMUwlzkYLUoTw66
KJO/uPRNmuwnY8Jmjp8SE6cpsR7wUgzjEmEKwrgB9C19sAJa8UYyeLGsAJ14EkvS
XnYDS1sypLB1AexID8q+fVyqkSdOFBKW7KbfyktDmOI8GJiwxXBCgczxvcjYd9ft
LNEz0P2snw9YduqQqVjBjuRZzfqnicypR0AzfcOKPNyeBfR00H5bHVBKlJESMaz/
2pQLnJ3oxWBp+cQDDxA1B1BFAquRWDOXL3SU85j9ETM1A+IuMPTMALt10KZGVKck
kTPQ+qLU4NRnzOrH/iAjsaE2r0S/mZSeQUQ5lFSz77roDYTcSMI+b2LH2bhV+e9v
O6woJvEeMB0wojIJZYOjO/U8nWpVbu8P7CYHqyZYYjwKoMs8ESRAI6+koVFTueTM
DPXez2KNNUOhM1ub3cL0JUThw/an0+atObrYu3wvDtwHkfhQvNdxXUz9u2oJcM4s
/t8TQUQowNl+e2VYU1/WCF31uO8akWXQh5+Z+wtuAhQ2BVoMou1fOTOdPhRei01J
p/6YWtx5/CvkIzy2tlZaevBWV3xR6TxpsaKPeNWV4kEz1xZOYplSVQPrckV+sZPk
fIEVqbG6a0qSasJSRkXu/DR4LSvHg+xBQbt8wQqvhmq7zqf9eq3AzOU2Z0XbE1MX
mB7IoJXCkYr1gckUQiNUXiv2jEiRkbCb/8x6kY0DtGBpGaaUkZ/rwB2Rm4uFs1XT
uGcYq2SGLJebJWhh0mthBI25dQPSYUb+txTiB4CZcfjy5OpTAmGcEIbW5ItYIloH
qecNx5EaDcGPubbHQpLXp5XOZBVQ0nztC/OSr5vNSolhWdoC2tFKLr9//1+jHMe1
bStY5Vb5YqvAPEgBA5Mx5hBvR/CT0cd6mS/ZlG+xh8K9mVtHyUBvrg/8yMkn1DkX
0UVFut4HWYmo8eKkbG/UQKk01l22AzdfHKjJIpTI5TqITXr0kLeKPJlO2bn/XsTB
ztYiFSXNbD0ZdJgbv5ief/Cq8MqmOlq2qBM8GcXjTqwhCsmI53qhu5PGotYfN/wG
Xr1VKKkq07FBtq2yHa7U5hhHbFmzPzF1fVprYaxJsS7oCby5Upo0Vi5/oVAiVQUg
pnF3DSyko5eE92CSXIscVWejvudfrpKMsQM7gwT4t1PKws2VdzgMURxT9PrOvYin
mj+7m6/EF9tE+QFD7um6UBDV4t12YbSuvijVYgxSBXlNTDgOtfpvK7SwfxFLqgTc
XpDUIsLia/QG/lBVJ8N6vMCakUbw/ffKQBU74sX9bz8ocrMAGpJ/Lq5HcT2YVxvc
M12hK1lUOgqeZIlMIxVfh2n/AX3qZNfcYV6cBIU2F01D6tkE5N+Dcb/Jx1LtGbvG
cJNgt3VTG5T7XIyaa8R+4V9+NROmaHr2UgZzN40ZVt9SgxtZ5z6naITFbUUbk0n2
drRmJMN3zc1TeRl3bx93rWJ3OEHp4BDxcaEP+RfGIu87l+QLUAXHhQ7H/wgBr3k/
HT2cKq27hDXcmvPsZk+DY0lLwLmk/YRsn7tZ4QbqyOs7KYg8iMtbFGyi8nB9kl57
6day0E9Br1RdCz5wkNOgQzIqHES30qdNcBVRonOET7NvouFwPklfWpK5kJ+QSa4s
QaHagNMQCY8vbZAJ+N/w6eVk3LJTycLViH2T63pVhj922qPuifgCUYLff9NVClbY
DE7t5ezXi94F3vjDZ7vp6/nX/fXkU18TswfZtqsyU2DA6Bmv/cwAC2q5+Kpqdx9h
Qa3TjAaELOiEMi2N9pkdht70feHmQCypRjU7lMHJt8zvHY/QE2UM+in0jBojV6tg
7WWPHuzMau+7biT1PzcVSeR4+CBHiXtlEtKEkW5J/E8PrUx+7oLnEw4iVezq+AON
x81HMpZytwGwT/mlsvToBLSj2VWb7Omks5a/ky1NnW3zPuRFS1h/XS9PjOBEVQ28
3u8g17I91xR7AN4OXoLmKTLJ9nIhfWFAra4KMaq1Xd0MMuoRUMs/1+BlBAtjBzAG
3igKmwgG7FsVlLzjQKktmohwuTW2yE1JXp12gcRejzG7AH9vnNBFL0az/mE+oYhk
q2hkezo7R5oZOlp4oiH4U1cyMl7VHBVVlYxAMtb1jh7fgZyILgpmzqwlfbKJ7W76
qa8sXF67oRV2diBte++zBwV3UUsnLeNzVOaXVZ1bKz2s89nF0qHmi71Rwa63hkTn
/CuXBVo99UjIuDJtVqy4HlBa3+Ers/PFxs7m0QVmpNly9KOHg4V35a573hVhPgjk
Rb607RyPrIvjD0t/nm4/VzFnFrWvMrXeprzbUaAs6KelOGxzmiaKBg2PAwOtpyOw
4u/o5T2AUAzEvTiEcKGIyB0I9CREmlHfOoG+TLlvPG9t2DDPE3ghtz0jinpeHhoE
q7BieYq7i9T0SNOeaIeMwU9wR9Gl7RvM9wSYj8X+msv1YVypr6Ru5crA/Uf5Ngsb
nRAKrK2TeoxfoZHTG81MciwtrZjsJsJ5wsF6mLt1nAHc+9AYNIcyVO5n9OWfMWbw
zwqujE7KCeKL6yoyofJawV2x5sT/1/Hi60nZVTmmMHMo3OihYnW1g0ccWpGTytPN
+r6aTI8cJKSCEGEwG7qBkjW31P/0ABvGtmQOe532zudLymC+QSSLQnuTKQulhtwc
4OJ0ybOQ3cDdDlIEXRDD+2XHVnDGb7q3UpRkKV0O2sgIKperH4wTz0MIlnPiXwni
Bf40VHIbpCAdsddidhT1rdl0999hl2lSOyYPQfCPPTjaNh/xsDg/MIUCpfT0Kjhz
0lL0S/SpQ9+SCwzRR78PKeo0UCusfuayB0+kaUPAfdBi2oavxtTKDxLqm3r5D5mi
2SXqsYgxf21pHO/hBp5vENYYTIBu1OwyoWr5qiuXgW5//wVkZql2rjloAaQ3YkPf
9NtnLX2nzW1+Arn1c0/TSN4t9AB/zMu7wOmiqE/PO7QMYZdRi9m87Li6o7IovlKg
3W8ywUGz7qYWaj6ZvYD38p4JFLlhgZDyWco0MRZJeb9UuOy+wiDg2/J4ibGU441v
UIA/z2/YnNlJi3UThjqk4riZ4GtXqG6EY2QmFt8J4ghTYzqmfKDEjoCR+DStjZgT
cktV9CyB+wYXbgnCz7LzVM74RRfDVbd7YG8mKGOGic3yUyOSDT5vwHUCX5Wj8soP
yBfu7/yUyIpNwJkt9O1IIE7y7KLuf4y+OirQ2QZ2n49ds/O8q1s5K0n92DOvz4tx
vBd9eU/ZdT6xatj4Kwn+h/PCiRurMg5ydU2HG/Di0xTJkX5o/4+3DjvBgkpK6dla
EQbZm8eBAx1Dz8eY2HWmTstuMM/c7ibZEKJ2dP7tmWDugeDGIegbYIWjC1yoxNeK
BraxpJn/VH3dPTgCoR+o59KvoDKb75DQ1OlenIaNn7r2xa68gUsAiMkNCFF/lRgb
DHzA6AJnlBwebWU/Z7bP0fWQhmougn32SYKtaxM7u1Orq5rkZXjy620f7lYrLPaG
6MEnvzbWphCPH1tiplD19A5S9+tAmUI2rjHXzQv5pYQgys25OPn52TO8933siR6f
S33FBwWMPBNgvcXr1eGM5Q03hYW2YvTW02DGvUfHkxy/EO9TlFbTL6ttPiUTXQ9j
iK26zlhVpp5BVFN2xvx67a+nVYGeAWniEkgEp0+sRbxbpgWpdMhdCjHUmj1aAE9O
e+Do6zJYk/HOZn+MvFGXJJnpYPrUXZsEk9KKHDp45KjNp4iXIz96r6yfpPBTe7PL
S1Jg7hf80OQOdU/6we7IHA3SRfUHY11HXGKhIaN81wy0m4/LXOEIdnQor08iPEhc
J6c9l++1Ulij6Cgl38SYiryQknyM3+YG6h6ztQaucQdPRxIkkB3HVZdk8BaZ5Eis
YtOX+Qd8CViR+giF7zC+shDpOqJokfjPE4Vf9ZoI+okj3kMKbF3+C6+IuN7x55k4
ZwEEtBaB8ByzsYx4Je/0Ki/jcyhHopmUjUHooeSHz8IyJCSyIOMgLwqMtkCIs42x
mf0rVdgQHyEbsLaZ7KQElE5neSc1DpY09bZUUyNoVx+8VZD6oGrI0VWzitJsEeCk
+7EWZGRZZ7wB1zZQMY2PrRASgSFE4Gw0QYkANNAxvBvX+gXjbImkrIGqTHw9fTHW
1L2tXZ93In8kdG1VdsjfxPvEKARcFA+SJBwQ7ASaY20WKyLF8Jz/PhDq4KDYs976
zOVQ/0jDsn8SlPriJ+9ULyZAwLASySZDawGRQr6wOFcR+RLeTe9eyzDqBWwAlcSC
aMROdd4OvXRYwESrZz/EVqaXoESrrMWzSfJECsgRZ0GBqyzB0zEoDI69JL+80mHy
xAE95Uf9RL4/72jaBMbctKcgFIlxByKGoH+qON1C1Uigm9VIXGpuaNkY/0Y9dFuu
PXdAedeSVI7+/qJbdgItKsIUhicDOKIgOjCXJ46vVayUf4qE3zLfuS/dx5+GMleR
lawNxg7Fv2CkCrEoqw6YhAfl+CZSEPcRo08YbLPSOHJhmfP9HlxJ+uK2wB319sxC
kH2Y/sF0NtU4b1Yr3DQMyW6PUykEwoIw+FcNfN0kPOyv/17EY9mGVHS+f/GvvQyv
xLVA12y92Cv6MBGSwWD3IjwAkuxQTKZqwHyP7E/WYaDEksEHyz6xNlRrNUifdAMh
gzzD9mN9iBYJBLNuPMV1+49SqFKPdoXQuhOkkMmg6JoJnULaU7RZHYmZIsLI5lEj
pZXeTUnaVU3MwmSRBGzGfiY0JjAHc5HBtrtR03iuzQ99f6Fx1AhUuIJyTX252qQV
Qs0FP+4m5cBvrOL9YqFnqgLtmlmNliyRTO1LxpxBpJZMEOnHNcfWbUYbNjw81Y8z
6n3AxKYUHR5hkUyMejD39p06aSo2on3mNBvkgc4sUfv793c1dQPQE91UbEH8+h/Q
+qTNuBEbRRyPOv3HTy27fYpyBkvqIs3BJgNn9liuqVEVdOseoCVlfIx7mNAZjBoA
1pviJkpaLnFTkNmPEOXhIz5WuL+HsXDZ3DD6SWzmGRlfmg0Eu1hYarZAO9/oxzt1
cG5rvxIXMAM4eMvSQbZIfG3qX1Npm2d+T/Q2D1EUd2yJRuccmxCyNW+fxK2zyFVU
2rWwxrHyYTM0Jg2vCt/9Z+1HaNVDUhtUKBCWHHNQub4TJz/P8QcMw2ck4VF8qwDo
WtHr3FVEhGpV8X5G55ivE8glxHgClWsy7spbQLeIt0B1170uOoqdion9mpqllzSR
X5aBeV5s8j3KAAmRlsqrqGawkGl8lEMNwNwZL7PnHeiUt+6k5JnW81AReU4PfmPp
SXIZa28lIc4pmeUHOZI4YkU8/RyRFtxRyAiR1RF4Ab0f1VQFRXhzBnI47j0BeLQ0
JfHAO3xTl+/LsllU/tK2cebl0trq3iXuqhv5Dqfu6Wk8wMgWKy2to6gT9M789J46
cmmvIJEnCX8XdQgPL5ajWzas5+CN1GiIkPLFL9vUb3CJxaNLDQQWmsR9iCyBp+Kx
VWVSkVttvHAXnz0Dl5B3jtvPNhfla8ZsIFOMKLYOcERf9UpCENuvdL32e98dgW7J
uM/PiwkDFvsD6Ioa/mQEI7hAHSnbnoTZKnBQaHnU8QS2el2/D2/ZTz/Mp/x7VybX
28pe8M4TJZ5nNUTLX/L+xyc9nXRhepGXRv5R034KzhdP0U3/zY4yF+0ZVAIg3zc4
xah5PjERArS9zor0qP4x89tYQfChtvuaIYqpQNCVwlv96B3CVrcg1AOApKLGVH64
8tZpKkUj7Eke2Dz+zmJTlCfdrx/ZVL0i7OHRtFs92u2aDVJTqwM+6P7vdzxxcHf5
22VxzxpaxKOpIAr/w70OJT45USgDUkN0U7l+GoYoxa8nh4Ww4cVjXXxV4H+4mw2+
wLZbQbjqJepVZTSJwrn4GZCCyDU/K2Gr8jGJgM+lMABwGvGiScme/OrSCTIhZSZv
L3EhCW/JcNH/bLMR5AbynEJAy2LT86rZnG7TPYG2UWPKVCtLJbxHCsiG0flxgs0X
VDuqhtgsDRDnCPljSAGlCJL7SGFeUXXVMOCVmkPunclKf2vOu65d/aU7U3cK7s73
XrP2cu7VipDM2B89q/8abFaP2DYB3d6Os5s9FG6MmP/AHeQPnpYr2mgPp3LZYin9
093AFXJQs7H+V771H3q1MpaK1KxINQ3hBA0qq8iiFTm1+Lq6Xi6RbFHmaz6sbPjz
bDgpATTKdWivBLLGotcss7Ul56Yi1dCsOYdgDfayRrwJPnejgaeEo6ltgVq8mxx7
FKkI56W8EL2L0QuWPH63wfFbC9VpQPThpfErOZRsILCBQvxT0dx5+2DQyw29YODH
u88dotlrfngUd+VbIvdkuY7IUNnf6a2w/RszN9AGeuw+vRefKPuztA/2zBmodhnl
iKf5qfMb2dG9ZYRcT6tDIjuXUaCFFeVKbayzKMrQ0KMnecS+uwsPsY96rf9OXSTN
A2tW54u8KNnExp1Wyzmdcl+6v5edqgMDxF6ttLEw5Fzga9a70lfJ2L7fg66TrVIc
R+QXF/yhOjJ0lyYk2X88YQi+QQhP9/7bT+QjEeJ7ogoKXLxIQCfZY+1x30/bVjjx
HQvfr5i7Xes1eIK2SWfAVs3yMf23hJQyut2HlMZKG8IJlCwsqWs6Ljrcv/aJ7SDh
Kt4JXdxIeRB1KtyEOZ/4ywDkDdu64lpSe4Up29DG2kfwzGg917P1u48RmXP1RNLN
chfgEkZx8m/a1QIsSzyRcjwgtiBn/J5eF5pNcmbW5dPao7XpAGdY4+pnEE05/muP
ZZK+vU7Lq8IXeIq6dWrVH2wHvOdT2cc13H3HdNHrIgHeUhrir0akUplj2iCXAGpr
/8JOwewnKENfrORgSZeRg6qwn85l4GBCZXXnFb7XN0mgf0b0QozNLfqW9MpPwvLh
ALTrZHDRHmJdsigmei0L0R022EMaZopPYm0n5RxIC+0NRKCAnU8viaPCkeR0L4Jg
C/0jrMMJi+1sAAyb8/Joi3gvY0KIYLShocqWe7a4Y+cR0AFhh13XwnKYVY95quVQ
C8hK1xMAgqPvdPrfOA+cfP7g5uPpSjv/CDmErNIGwZZaNOSIeUWX+TXdxGpiIX+L
JxG4Gdw7xwah6OqSp083dGmX/gZWgpTgH4iACVfXmkk4c8kC6sSw9GMc//FiFDbX
lnTVpqX8We0RXHtGtQaZkW+KRsiBpHsGnMVoWFG23EMk6nGXBqieYXY3CUCoBbNx
Khpid1ae6GFvY5L5aBX+E2kCC3182EVuDMwl0DRYLZvpXje1AWOvlbezPrL9vGSx
SUNdXWL6WXi0ohtX9kczg1kAlqpIgTlfD/IA7bJ5CltuoyQExeIsgtC5gIU58aPi
6I5rlqteMtZTNi2xGOXLbpi2KNV3HkUIZJ7Utc+ENMH44t24a+adHpT/cXGOwHi5
8mrafAOpAoFsB2CQ5AXN+Zy75vUeQKhdrlynD8254ThQWCE4yZkZW5LhFxYWvgmy
DQ5j148VLIl6evn9nFRpYCo6zsNAwl5+yBqDkBxvWxMdI/RS0JTxQEW/UC4zdTeO
0LX984IGfs8FbkzajN+A2p6nyKnM+gTkxH50NsDzns0DQCyPOC4ue/t4uK04215V
H5qU0vGvwps8VgLtkDmyf6pStxVbVaCMWVoM/4d+a72FshKGRY+p+li4h0sy0MSk
JVhfltfVvPhorP+QZotG1yxArGZupDKIs6BgS2F1oscpuGlRFul4xHojSV3BwqOB
emI1tJtBkXNEJTXcZNc6afZ9kVrz/7viZElz4DQen9kfV1x06QqdTT9OW3kTmMjh
UDGz9CMXCE6PF6i7iSlot1WtZcPLHnbrStBxnB1mcKfGy0R63BVn+qGMsOSENpFj
N+uwNoEu5uh7GNpokFUWatAtW3ToXI/JoWLo47L0d3xaRsz1KUGrzj+EC1dRg4KC
PDyFhFIkUk4T5tRFMvAjRkocFJdPIKFqoWrWS7kxqiFakOLis2X+Nwm6ybarz8St
AyUr26N21xdD7BlA6nmm4EAL7qiPq+jRC5LSSaWYrjTQUoXgrYbrzYJ976lCETrK
cYjLf8jqi4YLefckbU1UZwvKCfwAkRVioR0YTouM8riyv250oT+vk5OrfEO3swbb
y6E48W9cjf2RV8S4euGGjcuBs7crX4EWcWBm3L+cqxDXcTYcf+JqgmE4U2K2hqlt
P4qadjCoX+ExPgtHdYVUetWiKzq8CZMffR9os9DXPvTSbq+ltxmJ7Nq4AYTVP922
NnDUHDfr4uaKzDLSZ3n4vGIxRfnBhp4VQI7pI30hsC0QX06jR8+2z+fOgY0mWMgd
5nrleqovj/3CXT68TPGD1NVYHie8MGEQPVoBEiYLkS4YIqEUKfW2AYLxCkGbqAmO
9eQh7zSLAiO38djzySA+7rPzNoVFykR3/VOwYr2VN7xKQUp1pxnk4F8zNYQ63v+L
qJf7ImR7OIJPbr/rrLsVhMuP9//bwEy05tfc4Bo7CuohrAJYM3qp3WLh4t2P+rPz
5vMzokku99op+3NcSumhQsrOgg81dV/I6MzenCn1LY3DfwIn0jCHr8k692syjGwT
cq0oBb9OeHwkW+eGhTYq9gz3w4Lr7IIVqBDjm9VZDyS3AiUwhwEk1zsgAXE+Ontx
m0USpV4J1L3xWjU6sWVYoBTzhRbF7vFlfNvGY0LMSUEjBQxrSae6kyfDKJVzklZH
ceoZ+xhmIZBkIY4oHgm1SQE3t4NLP6P0ooRu+IAZA9KHWsWVVZsvBoZSu9eYtMak
/Z1HSdgcxVEkqtd7GvzkOijSY328rJcl2JYHG5LD0V0mhLlReJNYHqCwSevAVu8W
RhDiT+hbw1q9w5+VLqi5eL35Shd8RmxWiSbaZd/7JIt6JE72bdwIe/zaqNnxalKI
XiL+sodYk3iJ1RqgM9gYgXNErsn1BQb3BwlilXCE9HCTMWx5T8Yp4XAJmLkbLN05
qh+bDq+d19I5wkOALTbWSRh71DL1ha67jXU3YbaHBdmGLwmiABGQtzZifsDcpkF6
M1I2Owh2goATEnvZ3u/M0iwg7hauMjTdJdeqdM5rCf1JOWAdv5fAMa2/iqrtDQ6H
SxjG07qQ0apW1RVdFGV2SfU76kAL1UdnXRNCFGTvF3s+D+3rWbv7uyqpwCUv0Qo/
1Lw02ASrPdeH/6cFZoqlefFFZWNS8JA5OLZw6ojcr9uPQkhaKsc8ZIfJOGbWUOsA
0DxN1jz7gm/M73CmjCbKIMdWwI8CM/MImq/+e2zAsNJX1+xolsPjDIvRKn9uLb7S
/ISNrXB7KDuhjCVZH3YBABJ7vp08nD933my8xRoZLqmAar3zCkGLoqhXJnO5cOHK
F5HVdPyLGzbr+i1extoAsuOPGG28UpsNun5CeGwBNr0EBSQv3AQ9ywMgZVmUTdFR
9YoA/gIM9Y28Xwto5BnWP7drvR8cwgUynOc+C6GckssCnIcRUKkzMb15QTVHkmdA
xAbUvw7gZHp6tRPBaHsl1mjOcAS7qXT9VZaffvSWqQITaPST6d7FAjIn3p/kD0Nd
OxNAl+Z9rBbamWhC7huEZFppR/VyXYjb93CSbxi0Nw330+iBp2D295/ahfX+iThG
ee0/G4SSpc/1zooxYttHCfPqZtTzWPhOScMXqboz4d2ui6z5XzlKTdlhDw0W16Wc
X1WnzOwluvGqSTr5mrjfbnxy1YDdwxUMUzPK2CQX5NtLsTPlUDADWN57CWC7qD7r
/jENpKZj+TuPT0HvxMjSr8jBuiBTMyXRtWUudBgfTpLV6U48O9cYumvSNikuNrd+
1Es0mq53xqiBZ9ok8eMfW53whIgFdTP4W6dTAzdu0LxR4przLmgvYWjr15N3ucPV
tcoGV8A9d+yBQQHUWakcwe+ge0cQpah4desHFIT1pxyvkm4dotcTOmBQhl4yshWH
+rG+kcFpaVkg0WP4u6mtpYGaByzpLiZ8NVMvmNVy0utgD5hcgQ1LGOV6Xr2y9KOy
0DauzKV3x/LwJTKhv3hJ4hjEtsleoRIkBr17M5ett828AECjaz2Um2Cx3z+a8ois
aoV1gH40k73pQBE/IK8x+kP8AeC1iCOujP01xV7LqX8KBp9oCUrJvWH380hpMyQO
eWxLD+PsTkrfJ/4TDfn5iltff6x0MfbSea5C3UJhoT7SIpRvt7gB/ES1NsEmwlch
039iOJHbpouiT2BV2RXymCvqXq8Kr9vcYkK1fxVpdsLBB+neZKfao5erl35/3A7p
iMtneIQyhhPEJ9MVejkWKh4HCa9kOrPRXKXAZNCpxbOMUnC818NUaY03EBsFeRK5
2Dh0WLjjheWz3fNXumW0+vv6HLMvwzRB9nOnYrPnkWv5CzArpv+VRREM4juaVsfy
FGeHtgcsfWJbU+ZeDJRtkJeLE/BbsIe0WiJe8wKwznMeuOyHYIGdE05CbdyHKnna
AcA5l8LZ6nIfm0uWtOHpIuSanCP5bmPSmXbGIrhH1zzesZxf/yntlKDjHfUdKWIK
UXNX+AslGnLG3Pps6b9UmBzcqRUkOsCekNjjlQo/LE5WidIrANiHPRT93/MzhKUr
xNv74/DHTIoPhTDHTnp4ri8ivI0FlOzdUE5rKADn/ajAOdYb2PSbrv8CJhAXdF20
qo8ks3AF5itpp8Y3FrcPdI1wVTUpF6mZZmwkfZC4+jzJEcs9kBzGIsNDcG2W8bce
c5/NIqaYOrPjmrSgjxYGYxyGX6Rdj/SiIf7cQWu3WjVqe0yJ289FEZX6raoSHQsi
MWYatMRDZUjY5PjwayK4FEWyLlKrSCfvKD0MVmzIQMYc3AIiEgOOIAYqxlzpOd2O
n4IbaORS6d7q4A3qyU6Zqmc4NS3/Pls3FqqmAyYo+t/BHb+4A7gZhklOEztyMiIF
xJu8JGuJapSfF+Rd5cZnwuUtu/hcrxwEi3neaXvYuSiEqBb1p/TAD8UK/5VHk/6f
an1ReFstrjCoxVuOA51Tmc69ZUE17gpLnwkauBSBakk4r1pDic4TleIDwKVgJNSy
qVtNVMCnKBGMCYb9rMpTmCk8/UV5g0hjkxBYsrsqV7GFAAXEX/cyLxKuWDXRJRWD
i6ZPiseOFZIq1Ru7SHb8/lTOZPqOaBA6zLQssyN8m4Fizm7iMSD0SXR6oukAFMYg
G/c+8PdCgkXpD4iNxuil/dfosxrvdGkk4eUnx8x3xn5dxOwYVFehD64n1SWVHYlD
uMwy1mcz94PvsV11UesH7sNjPzhYdHQ7TbD0ezZdQAj5sYPO1yP0lsjxNyo9FvH1
nbzK0Qq7f5qnRu/5SfUz5Cx8Uy86viRGMNA4lj4o/WYKsfZOIMP/qRmA4dKwswCR
KIjv94WAsonEERR4y9yPo6HbG36Va6+QXE+59Z4ndPnT6f1eGeGsrTfLHYSOLpJ0
KCpM2NFjYoLYQzWDMO0oXN5TocoH+iHdeHdqf6uN2hf9G6q3e2m6HP8rWO4bvr4B
9K61x4g/p1kAzGtip+QjHSgiEXxCwea5bNqmFipC14nFyv2viU+NHf7W4w8AiPk/
QsvA2x8aV+aOt1229chlSITW3Kl6twVGR4DORBiCjgILL9fJQNpZoS7gxPNB56wB
v0pO3dz1E187kKH9r8XWyXmqRPVMgxTHOj451OqEGlZowdw7bPoJTEmKnhGyLDVD
fhY/rnE+9y8tQjXcdQzwi7Yg+BalBsrNKzmJn/Ollu3zYqgLZk4VoaAi0QUCwAgA
34cZAZ9iUL7UcetDtsf6LOfmnBxXQG6/9WaPDwhYEKcwPN2GgB3YpsY26lK8Lxzf
CuXZSpb97JyR4VmFzZc4TErmUsi/BgjSGRSEe22xSAfzl95K6eP39x+gtvc4L15i
CCqJssUKjRfFPXYjFwYWK51I0gFG6ywJTOB6HE//7v+f3PhDP7AVGROuVft9ajZw
f5lXEmEo/67cQH4oliyuT9fiRyepqPlkTW9da+CBIGifjv++JXMyuGUig4+APLjD
Bq4TOhhRzM+ZpQOsGRyOVrK4aRQOM7ET+1deVxMXr3QvxvvMASTwHKiudQqZ5YaB
8HP6R/gJD+6eHWh8IWWTbPkAUFTxdM+tbdi3O+IVxjLuq1y1h7HAlz6qouVu0Lz7
G9YF8zReGjLW83lbik45taQZBrn+XKGuyXagfSTkuULtYuDpjEM3GrzqgSLiTNNC
3dVDqi4jXYT7CZ916o7bD4s1A4UZREK5L1W9WbyJM8pIjV31izGH8M//h612F2z5
UFn7+s2h4qbPhUBKpvQMqA3B2Q353cloE+nm13mZhkc5ZxeaGGeEYdvvRUICkfvs
Mq40C4Hvsc7FmjEgvPuYcf1R90cjwiNTqHgpPcX7ldKifKamLYbVwWotBaWarsYA
L7FOYuwj/geh9JAqawKydtIGr24AoHlB/1haCGE0s1gip2Qjeu7b7I5SAXWlglvk
JPV5+04lg5g4Xv9JKEFLaD5vaf8Urgi/9tRBlBxLVIQUqs7InU9bvaLP7m3VXfus
W/FDbOWsnUtTo70R1bHb93/4yxT/Sag3JbgTYHerTIDw5LSx+aMLETkcr8LoX6g4
TiTtGaLlZt3hLT6rSVh4oLChSV/O+b+1WsMswikIRG8mAQHcdP/EzuDZ7rfHbwhY
5tqJxCDaIel7AIV08/Uu66A81c9uxY8SpuoPqWIQxT0WEy1q3f/v8CYq50tferzd
uzZi5crfse+El9+8qryklSZ0twIMgxcMFfCtC+aq7IASOhmKLrhH8FJ6benhxAJV
49bWFmK084ZoY2Fey8C/bVGUvCG5ZfGodoHcIHJ9GrH9SAQop/BpnIZ3jhij2g30
2i8iryyCBqNTors8sQ0P0Fmtm1q94y8zaUJ6oJrm0QGcqjg3Y9rOEJHGgxshPozW
uROoMvXT+ePZ+IHZu+Sg6+JH5YAfSaXNzz04735Z4dcqaGQGl2B/QH+0Fv0bqfV0
zx+X3Aevsjmi5nlVN0WIzWYmnes6bVRki2k6zV3d5yO2d2azOd470WiO0A4ESvNZ
XDMhZ7A9dZ3aeO3oQo/b2ekOSM6dcDbhzLYji7i+MxIu+84h6SJVEatniWgSGUT/
5zx+tyV3Jcgy67n/6JCnjDKUabcwKpaK2N39pZHMhQbZiW01KruDDMV7chhyPBMQ
PEHhNBeoHjkqS+NleFrSFCLQgE41vDcQFLoP6yTwfuWBL5Mxj5JVEnx2OSFwAkLz
2vAZzBR+FXC/l0pa3u2/XfDODtHbzU7XtEk/tnlPrIXFUx7j4qeKahQH4Rxh+ThZ
wW703jULRk4GD18P55L8yCXx2ef6oma/xh+ZJ7uiXrRvYyofvdI2cCpBYPMw/Lrs
K+QCzY+WTreNCbkGIstaD3p/5095hkA/kpJIDxk2DOXVP96yBKGfmL4LBFArVC/W
UsmtymxF5LDGlm/HpvEKK0V0aVXaV9dfHTYrD4uHuVkbX6FVRYDWOsJkUxdZnhM9
rVsOs8E/eaSZf5szK6iyWPEPnlAtc2OnRnCPrrXfNJritnjF8UtqYsqPuo0E1jcG
n22UWvRbzi8hZ/LnWnq3BcqXc7RBXHGIxPVNXdyJpBdqt9BlRiZ/AXDCz0+gYJwO
I66O6QVQETaAO57HX468k2S+Xuc5KwS8EWufGhCDAS9m+/ZgfLAKyGbxPV7pB74V
G7klhYvwlQH1/E2PUJGQ+5KjQ5g6Zq0Q2HpvYyLCw8PfYyvcsYOO99rg5vQfXe6O
9u5OVxJqZt8txGnq+O0FE50XUbEXzVLCihYrxtxKJJoDuIUxQjc8u4owVTdJ5nNw
pnAAMfRgWiRrippjDDXl+XDf9K4Me4WK28p5BIsIPnWmx4V8969rlDuX9L3uirsY
YDPfOELIeVx5DCDfPC5pxPrxniEID//YwvUZMJHeU3BFrbcXJHaAj4yI26ODffZW
JjtRyFzkogM+lf1c/fIRJPQl8f1NoYp/BrSMvVHQArVZN4GsS9obI1CZSCPWWXd7
B1bvItKnrUB7W/bkC4WUuG+X8Cf5RLY3jxvMIRbrj9X4FjPL/2hw8W0xuUkwJJ2O
d0RBeTy+syxFxMgexJ8C4qhzlRiIiUUn6o4VhIBsqQGrSnun7AOH5ccAgyqPGx0V
GppunbTK/SRuyozlSzE2Olf+o+tOebMLU2vql1QWthLGFrdYJqAJUbsuHz6SqgnL
rTJTeuN4h0ytayEL3Bc4UjEkLgDPC7nBA/2q+sNu/Y/+j8zdSW208RYP1YoLFx8O
sPdRDiRR0IoCr/qo83TyAjUMNFXDeaOBQ2J6Ike1/LUBGujNZjZ9jv59t13dRDtr
7qbFmQZ9JhinMLBa+mroiNl4v7sEWPUlX+OEXq3P2Ia0yM6lkh0eKf8tKzPQeOxO
Ig0VBFJq6kYKauL4YF8ONiXJl3ww9Q3kPvJoQLZfhNtkuXV5khgAF3IEmmt4P20w
iF+GIZM20BlSKqxuJTagle8H/DX0VoTr+M8kU9p8Ym3BgLZZiHr/PPPepl86brGf
c/anB+r9QorPR1sEtgVrqK0xh5KQrsWjtwmz9OZY+7Tq3gRoDEWj3ziGxRYhD2DF
F64UJtYc+4NekcdaDaYGm9GnBgizONb2yv3cybZ+nEXCe9kP+rvNZdWIGaDjoOae
65LQgUqE3ye4zjIGq8cnZMWqxtFhvuk3bY4JeTzM3ensAvDy5N7ojz9fybVdM0D6
UEjqqaM1DM5onx6d1hFivDa8a0jcPhxwsSJb3kFt1NSkHHLqF2SupskuQVTEoUD8
UzLlTRJjq2VSduo/RqLjFOnaaC5/iyUgijnSWaWHiAFp3lGIeYcu3FT5nb9wFn7Y
hNnNa0uv46BA2dYdIrrAgjge9zpCpw+tsroO8UjvWhf8VRbhU5G7vawu5h6IJ76y
C2De+O1cRI5FhEvDPxSfoQ54ndDy7SzZP6+3/2iy80OlyEBa7OJHwLZHPZnkeUvx
mamatD9tbe7cR6XmPdwbGbgevRmqQoljmqQ2ch0RoCcXxrZTjZ+ilbJmbaDYDTXN
dQXnyMs10Z3ivr07oleY7+QIgoKAfub1/atevLlK4kmMTL53TngR4ubhlQPQEN4k
MvIw7dDuTkyQbIYL1VxA+HeZo47jnKHxTexbGC9uyiiac4hAwatbbihuIvjpWu16
S01N/6ZSbHl9Z5YQaclhiGVZZTTOQg+WDnlgskHbvLq039SDga1Os6FTPQ6PRdxg
veVDoqUdrIf532qVXVICX0Uz2kXjQehiXLUKA6QapvIW2Nc2841gV0KfqhO7BimW
YxIxXi7yFxZCYeqTMMpkOUKVRDg6AhYsnPZmTBH6M7OqTs8p6xvmX7fqWDdJHJIh
mV2PXLytUXdlGNVNM5l7LMPUCW7lo7q1+f9XIrM5FAzlsp5dSFFdJEOWMSb+jBLN
fAi/tJx1O98K7KeRIW5nNNIb6YiG0d3RWCOwMy1PraD5vKHzKGlPo2jbFQpq0lz8
MULpH5ZtLuCjty3tnZAIdZRD8bu7WvpUuKazDXV1qpvHZaiEHYatlyl3tJr2kWtB
yzrIoduSb/hP+McjbqGigf0z7h+J2xJo6FPrjS211673RfwIB/6njm7+TZLK8y+5
TWJUyVV/rUynJ5dz70y0zcnmdRhs41xUnRsZy4j6VgQaHlz0t3W31eqeMQ0pEIEu
c6ARNK/wcRRfhFTjzVUitbx0145OWd3sTWmdiWwg4ZNXVkLA/hO5iU/wvvMF1omz
jF3q/B0KHlD6KOr5xZEIKVPRa5efic6QSV8nbDw2l/b0cttavR7cLj2F++U7x93l
mz255Jhac5Nk3gQyRQMUl7T24ANowmx9lV+NTaa5MvV5d81ebhntugcBQjdN6jBW
EueRoQQGvNr5nUBjj68GOZob7hHCtx7+i/cHhn0tgqPCbgYNNEBnI66pP/7Tz9TJ
i0UBqqcb4w/lFUCmrcD2oERQOSgus8vGRQoPnzu4dmrHKpHUMaHthSPpCxTgJxqo
zkTNOVWKYGSQ92ZK171kCjKvFxwJ9kk1UEyvcP7UjoKfGe0tDbcPzJdWgvX8L7S2
ZMTiiRPHTt0i5IhehvyapY2ZlLOaB2BQTA7aXAaGtefwDsEYtKkrn5vbmAmRTzr6
+mrHOvPkGGEScURE4ZYTBBCPKnvCWIEY1dt1FKjO34Q4TPV5dGUbEEpcQ+pf/9Pe
yxiHalzBEyf5zsQaYiGYMMY+Lob59XsVW68YI9GdtgmFuEiRRmd9ai+sGm7uxGSi
EUIbglJdIZXwKn3qD4AN1g0ZDj1uErYyNLdR0cHhWG8GyxsNwXsSDWH2qNxsciPb
qe9KBy4PTK4LOqmZp0OuncyolKuNf+XA2+FPr5OwODIIi0RLhq8NGjzboiFGZTWr
cb1RfZPFBObLF7PY5w8DgmSZDqTg3uSmQLICz1u4yqL3UsXgKweiD3oJQeudND2f
QGm4WA76dA+p4rT9Tmf8W9MthQr5jmVOHBb1R2caYiXleW1R46oLLAzBv1fWHP02
d0qBVWT/rPYKIPfOjLnPAzJ8WsltcbHt2K2Y9aD2A3HrEJTmMi/fLxwLx0hNDwMF
bQLQmIo1YUvbQDGeqGfnGxUksJZZBGy/0+sRRBYafIJ+fBWEVDvd3CrZcp4u/EsT
TTCQ4C/szpaWwAxDHyhhkLzTn6DQ8hjE/8pwb/fgFO0mcGdy57O34xgbdkNA/SNr
mre2U1+VhVOhY0yiAW/vmoOA0wpr4eaq5GVgEeNBYkhLoqhzGpZBBwTiiD9RyxP9
P8kW+LKd222Oj4Q8lFwmJek0CJTnWRHE/ifkCNjOM2/VQgwmUSMoRH1CWguDF/th
EB0UUTLR6XweUpX05jhlHH4QpUiin1lUKNvIzXzy/n3E2VMbEmTIk2shFWl6oBt9
ZwOXCLaUeBapBJqEjvFaR2O9oVihnusLw9uTSwpPwpEpn/0ve5DIWXjBIRshCmyS
m90u0Pwy2PyfCKrd5LfPdUpVztUPwA64xE1FFDxCO/OaDmDJFT4tsA3Epg3jpDM+
1rSOiraSBEFVJKrS6Rdr3X7G/qkhHnR+3Aa9j6LOb7/EfDaBW/5c1U5KEolu2XwF
keTt2DbsSGQ7/2bgQxqubmrf1a6jtn9xyCGbZxHjEKe9lwQhZjGa3DhtlsKkfxr6
ngKQFvVM22v32mqFn7GJG9jEF/xN+Oul4uwffVLu9xosew2CmhZ6IgBTD+zvp1sv
82hUp3iPWZuT8VNA8fCLpJGyEzn1K/KTtouuMN2bB0QhiRCFVeEzt+LFLMbWVGVR
IeSE6lDpNg5YrM6KilFUcA+/lb3AfVy5CDbMYqNbTaj40wzGNY08c/sKdpkTRkZ3
fB722CC0JqcdyoMWj6l8fw81mtwXlhJd/mIhyA2KyZa9CoSa7nLF5VtJkf/dBx89
qo3D8PSvYUwsnlrDZUEe6ST7uso5k3pcE8+5mgz+w0c9aOFo948L2bhrqYc26qEs
kROsPsL43KlTzeB8dKQmbwUdqsGnv8GunNjZbLetYzdjHUtZB6kEr+3QeB1Jix1x
ROeurTi2bqxlDVbgAW3vfYURYZiRtaLnFV0Uwn6iGC+RNDF3M/ZaODGM54Sayg4U
zEyyDvhmy3QWDg0pYr9ZzhREnIDw+XHUeYD9Q+o31+TN8+7W/Idd/Vsnxbfm+7M8
S2/noW9bz9rAYhsk1aPYXMblP2zQaoK0tsw3zeh5zgI747H7zZvl26pk5r0sG5MT
0np8A6BkwCvwBgHpxA2ePYGgJlPaycoV2lRhiPMAziST6Up/7r7jNuysRP0v6Ji5
uMfbBl9GzO0+1Xj7XnxrJzFrr/HPCcsxcwXyWbZKb+2yYID6bdWL4jEyPgBVxpOy
BKf0PEXGZsCCTKlXaZQFly0I9gUqOPP6jdoGOYSbNPfJHM0fixCfcN8ZlDyWw0Ih
5VhcnD9PLnHBL/D6PRpbpXXuZxhDyLB9j8moNhPeySPe5osCF/EYnyNfjwGZcD/A
C2P8AwbcTIV8SCd1nijI9I8EHp2nCxwQwNLh+79rTZt3qo/bxszUjn2BV7Tne0z0
yychsg37ZJrJFMzb72h6N2JGJ408SGhOyx9DFmmEwG0XVjLo1UCUtCTHZWMbgpCI
2H/K3CAV5wuOMZGY927LkZnyNZIEefoFLPHPWCoELxnilUHI+EO0eFIwIgiqyxQD
pbYdJGM8uGQJ+N8TtT7aWUTVsrDJlDeoPZL/CPa1ZjXLT1Okmqsyq9l+lSzB3Vzk
rDI/FFpJuHDPFi9t0AunzMjw+e00p8Nnu1yEOZaBIEW9PLa7wUCTX1s9qKQXfpso
LmHEtVNmIg29v8oGtQE08xYuZA/76n1hTojElMftGDjjxnNmweBjwwz17xUFgKTP
06XCI35hMf/hOXI61WnzJ7GxuPU92tD8ADUUCW/q7sLHHshWTfssSF0Q2TCKEN3m
w5ixJ64BNUyovokrSG8zl7wGtX0ZWjgH5rRZDFCe33z8B3vBTDzZ8MXQJlzv99bj
Mq0kecjRWtCCZBa5BnhlSnR2R2SCf5PcYvcC8NA4WlF1odBFAv+ZTneUvTFeBlgf
4DMJ8xieJhJfrlNNT5Fd8nOmgfOWfOpQZe3kvN4ig+AS+eCWzxtRTf6cu2VXzQvo
L/2V4Z78XkpOmKD4AWnrYNdb8wND77SPH/lbRMVvJynk4kbk/1Pxpzm0bM/oYH9b
+lExr9mXfHENoRqRtBhyJ5++ZVYB9TOfOOA8WMr1+l0Xilsyqb/OgBEJGo1Mj51w
TQfgA92uTRst0NotR5+1EDkP1iHtA6YVP7T1Tg29dfzMMvGikjrQ9Lml3wDX+lCb
wTnZ5RSMJaKkXwpmEr7Mx6M7MEYxqFeDdKXFhtnbLXBq0XAdVuvaMHHbaehSG/OS
LlO+V8rEhY6/RgAPpDwi2FL8Aw1PdBbq0oJ6wNv7DS5Et/XFKt4nhlm73cAes1Ec
pRH81UMHvO75SnnmhjITXiUESd9SO68W+uTqNb3xptpMnvpOPpefvH7g4aRrv+YQ
WyMAPr8HiRqzwrKsfQoILqF0tkZwVOXhdD2I6JRmBOXJ/jI45mp2BhGZpQvaZcXK
PZQjBM0Yr0d0C5EsdzU8NqU6nJCrNoSCmEoBF53KLCDclV8Q/uYerB6XekwHWx0E
GU50ahN5A05v3Th8GA67/z8uzECz2IwdElUGqymu12QmQgor7U8MC9ub9dnLOiKd
CPN83qU3fyQCiy3nx9o9JoeYB1kFV6SykazEZS39DtVwUy2JfZGAWARgp7HaP/o3
2OgdIgT85nxUt+eUMITcNC5Y4KZz3U86YxLkfu4FVIYo5KxFbGLbhMe4VKZ/gB8T
t2ADSuh5hDo4LWZg2IV/pcbHlTx7gwqcXlv9++kxd+iOzCcQdgQpZC7/eq4Yf9C5
PQxmjZZ0b4UgYGksyD0jg3qWgoHJBLRc8VbWKUJUAyTGxhSFUglJ4haYjk2l7A4o
zh68Sv6leafOYIetPD7SiexBCE5BitsGuWLij21vg4AGxW6V6/dD5RHjN8x/yawc
j9UIdIiruuhsumPSwPTGvgHjMuuEJYJ4mOqUQDw+ZhoqeN22US3EReH1FmM/EoI1
1lF9rk557X4OxPFVuTofUrVnsz4aqWTbfB4lA70nNCFdKQ3XWWELkI2UOCbsATE3
R1llsQz05i4xmP5+RDC2AKsijdxC/s+CxrmwdbvqkK3pmLptt8y6MHXuOqBXK7KV
RraiFWoUkI4jqhRDaPjssF1hUSF8z9VzA4VbBG2X98STrgVLaPZLwKnVg60uoGH1
yUaxfGGWNQDp7aTl77dNhsg2vjsYWMC8y+zRmAsVYET1rGFEsWyP2QR+3RfaQdNT
KKkd6rAm+4FaEIWE+qWeXjYfrjiKM0djvpzk+RqzOqTsvCNr3c/WEQskApiWmhiy
LbeE5Jl85TfyYIl1SrBvOJJ+V0MwYQb+qC9FCf6l2HxhOv2Yr2e8vD37lV+BWPVY
FMOc+2sMIWDLkytYEt8enrvAdtncoDZuwFt076A64P76GWuh/nKAGCE3UusUWl9e
5K/jwx6HxPViP1isCU//99e4TAKuOtHQ3Q1gUYrmBS/tZSlP+9JSqOG6ZzwyPgPq
J7Bew8Uy30maL795lUXWLEUUD4O1h19inGZTZnurRS/Jyr3gI4gtUoRKHR/nt2ci
B4DcJW8BcISe4mk9lT68K6ft7z3y2hBNU9Xa+SFvtVYdVvqNFFapVxqOcm2vauhn
404aj6N03QtsMK04sOQeC04R821rBgz4S2RsVVW0FWLDVpmd4TyRpU4A8WTeYY5D
OHfOYee1JwCgUTGqZ8VzcKyIBTpMT1Afz+nwBswcAlm4lR/WHjcjvQgYESTIZFmt
TY/iuXJe3l9F1lMqI1lYNE0XioPD0phyiEgoXTYXQmnCfO7do+BeKNtx4diO0cgP
Uw4MFlvx6bjxM1VdBojheZG+CHfyz2UCjCFvWKT3ijck8in3GVUeb01VhpQj1iZB
eaaZN5nYmg+H5w2XlrOwpywettmQ2SdShNsxvDPpn4jMt16Cz0tQMGDpnH49KiAT
+xjnjyokSa2Ch07IHg59jHl+1JvS1rDp30bJy93BLx6onPaoiPLQYdQ4YH5jC6XV
1QQC+665K+sF/UsbXS8k2BafKmSYZTvpcS1gmdaaEQbQAK5jqrs0HrMtYShmZ9OG
kFIOFd+Dv/qbZfLImXzc4Vpk8qjdCALOamwAEOQdTt4rV78ko0EU9pJ0LXcaS8KA
GmUyLxqKUtEshbNB65KCe4Fjozi2GQ3STgIoDkOREKPNfRZJagFuLw6n96rK+zQ0
YXmEAzO1JdQNCn3NHnEvQrlldFtuz0VBBq8b/tUADssLp8Xabif6aGiPFBtxT+us
9PlCVa3aX5mYGGDq+TNlV2jNtAttegmKdbVCSZa/kWlAtgfoDdAAZwMD6kGswTws
l0eKr+wSM558Nu7G2bLLGNlo+13Sro+iD/eX0FPJvDoZcBJxxT+5iECd0XIa7gx4
hmzqwJovGeb1LnQs2cXEnDKdG7oESwL113Da/Oa2rXSl5ijTD/b/IuGZKmVT10RQ
klaBcxWEPCOCGu1nywTDKXi2dLVujbSrrf7SVXBfiA42jelR7/pC8aj80c9fCOBb
/0b6cEq95OhCdJuiTwYfLcZ69YtSu7f8y/ofcebSnhtORHzz3dMjCZ2pYXNljaTL
lomDL0xsXA7ssOhTXpR1IPaUeeRsBQVIrIpaOYj6WOoQpI7YvT56eI7FWNGI64r/
GMqfpDREG593vaEbTUAL828zX+0t2buDUYv85FE+0vs956VOS0Jfb/0v6E0Hmwy/
jKsSfYeim7//lqCgojMZ4+8FptNqH2MzgTUHXFAJugdtWN970a9gTCp+ItUrxVPR
ei4d6CjkFRqc4KZHWmnoxjtk4tuVhN0WfooZzJYtqJatYkD5CUeceuq4l8698Snq
5zScezxI+3DW2jxN4ElNGklKoneKJ/ZV7T3EnDbkiDIJI7tqILbY5V3xR98iXuJa
aft4kw9biNsEdvQ8MSdtKqStKb2gt2r3yjYFYWmUOfDBQdASgVLHWTcNh92ljSou
xiwb8d5QC8CUXPcR46xPON3scbu59R020SJEvWY/QAvaejIdaSjFYjTNA8aZfK3e
M7bqXxfV4kLzYA+uYzZs7uJPIubWIklrDPhjsCXQg52w7qfaf6jyH+kLw4Ub/gr8
voFD7TQTPr0OXr4WeAAs1pntLbPdDMbn79zaFgDHo0VnaUCdKdHUtbU946OIwBNj
mAURuza826+xqSnSv3J6QhlstA4XZ94UDqeYKtYijhZ6UZsomzUA9ZWuqTrzjMsz
zeKb20UXz7av1UMtH0GELrWFmuFFBFNJ45m/l9vjCbMj4Oy07LQfxK7muq3nvkp5
VjN9SLQdTwfEIFDFHpFYtz35zesJuh5+1TyYW+swjiVVNd3xsD6iWNSLKNeInxZ0
zR5mNpqwCu14hUHH0REqy4j8zupnKqJkxvoTkumDPPLWYvogagdfYlZi98XkzBXa
nl0o6cDO1wkW4/z+PYwi0f6dYUSP0YNfqHuUvTn8kszDOePcswUF2IiRfqMR1A4Z
maS2rAWfjiAb179snQBMK7YTHiOS032GKcCTBAgjUyY/mT1NTlKvqz3HyfjJjdcT
nRyyu2J1xCGIZrCbyft7BDeS8Vezmu5LIbdXTGSdgmiqjMSg4jLYOSTc3V5Q0cnT
5EqOzRwjvK34Afqj7QfN31VsxDw8QIohuG2iNLy6qsXUO1U2cDDnLloHlajYIbvQ
k1ki4gmKrYC9zPqi9HSiz2auwq0OhCOXkJ98gE/7dX/SRVz7O6xVITi7aaUa7Z7H
WiHiIhtaiaOEQWbeq5Zt1P8zIXXX7byAcakH1UzSpj1xD8NXBGw87l1olIkot3vi
F2znvjAcXFSF2i5ESbSF8LoUBBy7mA+PVx5sF4kneTu6j4rkBUeaOvGIt9eq8P2Y
A0si86hrOIAyzCz1jKtf976cQviKY4tmkKv+xlC0mkREBGO6am08P4X1iY4eNt1e
UlojgqSzGNVhp76mkoPEUxMtOmp8ODjXzHWhwiEHk4rrXR6NV6wYZGC21+C6dM8X
EV0HagHkpzKg1b2hxD1aucI23Jnv4eP+iuvZs+d7+QRdjF8Toi43t3YVxZitpZzm
2uEqOQs/IY3XiX4wCJzrhzszMzNHvu1Wlg1g5vI9eUojg1Ll69DrA9V6yzROrLxa
+z1FbHwCiBnYlAQhDFBoiMxAXw+Wik6nb35WwxlsWhvvQKB3pI/j3bOOGGRyo+J1
icnlzjRGPWL/glH6BVWAzQ7G8SK3Mjf9PxYsk1L60nRUrKun6S2Dtj6Aga+/OOWs
jRc+DHpLPYi9zAx9U6vRwOCmU1evrg71OtLniYE4ld+x0UiORNEQjWFnRZ1bNVdK
S41AP/4P5MspiqlSA/Yn60tmjwjHNEzrAozs/P46Dwh+P1t8RQYuqq6dolpSWr5A
iOLo3KzDP1pI1ggwBQD4Mw37cV00/erkOe9DjmPC+FocF+fYBD6d1hiZzcdTyIhZ
ipbbhmzCN/BMb74nipheZbb2u5XKgWwXEQyCzk7iFu1gJy+CcF3Fd38tjR59ZoIm
MsyS9AVGKb4GNJNb3Z22PpYBf0BApk7tj9Skx+ZYP+efkrXtPe6oubUyWjW4mBp1
TsdicO3dKBHXUl/jlD/4uci+Y5Dafl/n+OGY+nb7ApkFpELN6ufjbBp+VFOcFJYq
b9rLEPBngIVe84ftLVyZwEiSPZR2HspbEFJd3F94q7mYlt7jpmFMb3vqAcR5jABD
5m/6i8bZjLx9OTRrB9qP2ij11QJz3OxgGYZwX5pI24saMZE+Ov92bmrfz1RomY87
wAdcNfHkTegRhmsYorObbV+9QHFPouqsmzn2q2mbLNMp3gYkUDxPxQhYd3ioNPcz
jiLUcVFW5isVO5TKw5215+vUCBU6Y4o4s/tZm3sAlQS3iOcqNImUPKtGvgMhhbbl
8C3IgNRqhC2OEPNprS4xUuvZvePxjbBcfpuAlimqj0HuaTae4B68hX7ieqwRQMLT
fcVvht2TqWBpuU0LJQt6jpOx2xQcJqKg27XjjoMIaFGR8y36rP5eNMeZMD3rYo5m
iSc85rlj9+ubPSVLGwFlCp24k+BEPhvS/nD3N/n21FitODuBq3bXtejMRbtQYZvQ
jrrhmrO056Jzl76fuvoNjIEVgwFgyMePzSdYZo52IrzRT/k1NitWNiapgiujmiCe
VVUaFAVzxLxNpkJSoIv04/P1k6cSFCMiAKAzK3mHXD3TRuo06Lm+RTRJT3OBGu7a
wPvAQcpFM0rVRnBzc2sfBVV8e6e/5eXgjSp6vc9ANx0ga7EH/L1f8anVGn55d05Q
XTIqxmsUymPyIFlxre7S6Mma1ONPtGawiaUEqkUfAZfp5vtgwH9JAc0LO+CwdUdr
vRmbeoC2HaDh6ChUxVE5GsgTTNFsZExzQrGZVcQHZQC7x80JmqE5jtF0mXHpykDZ
Dvk/Fq83HXD5k86pZuo5RiFYheWc6mEUxYlahLh7xVaDjnLdsSgMqTNdUYdiCoSU
USeO1VGtJzGs0wQhNknE/nFdvsSflfDQxvBT79JvzLgHjmhnnjEAtI+gd6vo7Ybv
4FQs3cV5D+c4B+4Gk0/EwAt25w/DSTCBdpKEM61zKM9GlJjG7F8HpA1E9pD+onxN
vKY7Zy0tpOeMTm6WkoYgZo5XJYlZCUmJ8GCHm5xAE7H28dITzsB0N2EYumqpeBYx
LjZ3V3aGcrRGkz6zrRCp6hAPL0Z2cnPXu1wsnojekhyYPQbE4T+v3AGaPs5eiCKl
UF4UWbk8n9WpK2tdUvfLRBAZxkyYbtVSYeXzTl44+Mnf6u2Qp3467Icb9KbhpTs7
8y2Edkf2MKsu9tBe/icvcwDRBorkPPVOJ0jdEegSI1KUEVGeeFmFmCxuUmq50Kzu
Gqn1aNrz4wh55VyC+iXkV/kxbf8d8/ONykmXSRhrEbFh1s0GLHrIwCUPdLW6DzcG
IUYBKTwsk9X9uw3d5jC9FtFg1aknlGsYRZuDhytpF6JyoPTxuMW76bSLZkZZeGId
7J4QTCM5XytsAgm0KDYwJdsCXSyJlGxUpxyDbCGHTYVm434NTcdFutoMrgwb4YCX
aTnAzjOM0b3J6Ev+AGFZhi1SOuWdu9n/xuz5mCZYtwjsCjDSmfyBKqwng15Cn1jH
bn9mT9YzR1/E8h1nDpM7hGtfoJdl3DxZGhSFinul2eysuZ8MxxXI2GP8R1sx61Ui
xsrx4rZytL7p6qLl0A2KIVg/SNWibMuoa5nT7vfgzMst268tPpIRiwm73E1rMqBt
fqxfNL+7xCtTOvH52+BOgi5vDGRwiaz2/RIy71jSgKEAFNZnz+SZB4477r974k+2
Ni9BA895KIiXvAllZk3qNXv2ZG9YqgTVzJpxmgCNFH6pwtasBocHAcmGqT4kLAQ7
ZBPC4tjdhbxZ/OmJA97Pr3l3X7aBxVc2PYrSk1cb+561GBnFfuE3kxKcF3NC3NFj
nA08JewoXYaSqs77uEf5Gs8J176fGdJWQvmP+v/q1JblHmcXam7X1Vgqbi4v9vFA
asXYw9NecNtv9M+h80KUI0QqnA3CwIIpjYx2IpgzqE4c2UPuKFfN9rL/kEbD2j/i
hZ5EkQMaB0KndXprRnlF51Ba0TuwKXbicVFfpqKMF//nRsxGMuAt8yjVaftCcnyT
nS0/Xsomp6z78XUY0wcmKUWzlYonyCJYY9yEuPdHPEokKuLWlYnvDxnLCP2DIx4D
sRD6DDG0LLJaB4lsbv60Ji2kniWqbEc6dNnuO882WZcawGeJuhYOVzKuptkxmNUi
le0Oe6C7XR9Lzn1Hb3jjEYIOnFRpJSRr5QivHM3a4wcgKE9Gz/sp/pgCd9b+ASt9
x0GPgVeEOGXjiZxKgt2DSgXgGLMAxSZkWN6foiqCl8wRyyPnkkwmwsu1wwZuXdM5
j6TZm9c2Ff5unt2u9Js5zkV3y4l94rWU7Rxq7r3KMZTYIGkWPMZT90YRK0jnf7I1
Z1WTProM0r1tN5B5yZoOAkIcKTJgCQGnzfbzLJr9Ftr36PF7NgEYNxc4XbOuOPSG
WoD+Hpwp2khB71tiSVPqZd9yOPsZ1fP81vX46jGk7tF7x5Sc9V8xSj3ub9H0H1TO
Vgok/aCoBMv+NPelOwmPimPfCaY59oqOj6NdBO4Wgax6dEWmcyx5+B/bBdFvjB2h
xPtwQROOiqcYMiZj2hj0v+GUJvkjbYvLhOduhatF9BqB/lm/OyzBqP/tLQ9Hqijy
lFplb6qX9vv3ntad+HOjabm2sNTjkiyeQ7RlPPKpEvsKu1KcZX9oUa2tBqhOk3Ao
kiQHELPhqwx0Y55PkwonocsDfZFUdJGczF5SVYN2xYYo6xFr2rm/GxlwiMh4UJy0
ZBHJq2hsRdvG8ddPBhd9cJa5g3FM4UekdEl51U1YepWBoYZ/8PEz//taGt6KE96I
WklQsdiVJ6CRowfWLGJYP7DbWCkMQUdECWzVyHYSc+vnPXizJGCkEHmcXMakkJwv
8vpf7yaBds5gUL/68/pCRM5/+Vy/7/TSIRG+A/d3c8EEmhbBZYsBt9hQ4hEbHXbd
QWa1dUwrOts8r8iNkcwLb5OyGOO9a/zrd6uVURz+GtrwFH2XRDfTRFzNBQzlrwBi
/VkYIHGKKJUqH/3IvPRKxtSg1N4WmmGj8SAlebosurMbzQYRjM+JI44GrDPDr28k
719XgIDtdTThs4lYcc8ZtlHgYxk0mFA/hoz5Jy1DllkbNYB9PeLUrrr3GlgteLdk
vZTo9an+QSdp+GylyUJ3+1uoS7i4hpaz0hbil/mjBUq1i0koZkqCrzl6AnarWyNb
3ET/Pr9JI6u8JYM278PLS7h9cdwsPLbPrrJG5Xh36YJs8fHLixJgigTbo6e3zEhf
FYmc3cuLwx0B9L3iyxD7tplafDYfYnMXh1matdmnemXoGJodPJhGVKCJHdK+66Fa
a4lE4m82APgxuJ/3go0IQxxUevFUHxeE6ag6vjr2h69n5g5A3qmPEUIw4nOzWllU
rSAypHJYeuO5FoSgsRlzTSENZ/4Czo0Jc2wNjH9T/kxb2kI9rme6o4dGMlAle/h9
WIE7IrHby1773HXa67EdhpSD5zXAWObkqc5SYpvl9BosHdwq5dJ5MbK5A95hR49O
mJpZn/jnO5jAHPgi4ELZodA+G46XjsbgokJ5wXfdC/6qVh3WTDqKUvhvTRRk5Y7k
W7eW/Ro5KrvGFTiuVaPkQ+evZ9z3Yrr+krBqCfDNKLPb9Vaiqt/MiVAsxsIq/T/8
+IzbVJVCF1ISXz60whCVlVJ3wxmeGdV9+3Dko9mxZlcl7MHx7ku6idVRJYj5/UCc
Ez5pUhpdhYslKgJ4359R7+U3KnrTaNYQG/1X7J6lgGZcdoLUZnz93j3KfnWlBFji
I6RQ7wXrzG/hHYGNKP9enwZKA32qOjXl5LHI4r7bN32caOCkSdPnex9rjiC7z70I
1YYxgbLBf+K7TbUu12PyoajLz0z03Yk4evHfTZcZs1G2jtTJot2fgOAEDiZQ4e6u
p62MSxWaTrbFVkNNHettf2lvdcPxkeufJR4rgpnS4WUGVN3LEEBhROIECIS7AsHI
2jboh2k87+7HnaFjEZ2uYS6pnjdAMjMUJlpsMD8fM542bzYIMw6sz80gcvgE6HuF
PXOKoRm8qMnZFvhlO17Pp1bdyteoj6cdX3aksXosglKD7uLgvLtvTuwcFoWKFa9s
SGqrh+mxMMAPwI7QKqVJ2vBQtKcivUN5GapeyXzv08VvxVpoH2LvOKZzDYElcWVe
0nyfn6rjwa64ldMPVDBsWGLlxlouzta0VN/mnuwuMgiVYtPh+JCo3URHWiYtDTyW
Xl92MqW9dYXIyKXASjcYQ3FMqpwFjWSJkPwWfRnXKWsT6hqk4LMaKHemUCJjpCbI
adhy5vEtffbvp7HMrwJmPBWGXt8m4K//fG9WG40GyIW0+gZPVw6hb2HVcAtr+3Yu
9PA0tbuzT4/BNdrUxtaeObAgNsk0yJ3Z4Y++CB03mgV2VofS3uPvLTWs6e/fa3EM
nN/mo5b5mh3T+CmcuPn/rJ33lBNqp13HTp4YS7QWXSOfhvr13sqJ08Suo59SJ6v9
j5Yq3zQwhfE7szwVSqGoxFY/B5lTj4+YVIE+XMZBaHSJ49369Sfe8P3PhRB+RAer
MgxZRxSndR2r9YBy7ElR5ejNHloZuO55/uqs53erwt3wAnCUpMGmtG/IcTFJkuCZ
uQnEtvYKHSQC8u97EwYCAQsgYQKHJW6cUkGyQsQULFlwH2Hh1ZeQsqtlYSq3dhb7
3waQg0trS/25yAAOLIDISk1HzpYK3tTApDWqy8PJEzIH7LRwJc/3ixNTIuoNB2QP
0uDNjxS6l16fJlGFq2bE8I9JrYnziPjhGc+Otwg1iKIWhVixdJm5Ve0FgBcBS8yz
j+WOMaIiz8fZh7um92HHV4GL5mippjG22fdknCotbFarS3zR8KtmAXHa0TJk19zY
d+2bRJ8VMN5IJ/lvTg5eYNEDefoap7DIJj6FIuHJ76USVz0QL11zyhttUvkwwSVI
8tq3hFgydp4qr4B/pbf0EwdcKK+yJe5ucYnvGu1hFDP82p99JdHa47wDh8lvvAY+
ADRk6c3cqNmEGal7k3Cuc94yeByaPeWwL+DIvlL+ev8PRpz6C+nfhnr1RGJ4/+uJ
bkEZUd/wQcu1/GOLec7Xss+F34O3qg4Q0kYbTw2JMdD8apAVNVRRJw8QG1eWN9Ry
unnnlZNusziuXifMCXqqJgdVciPknYrAZQxpqkjCn+8125GxSj1q/CqEI8f5tSvL
tYUKzY9kYu3UYnwX54MPCW478YWJe6ZwPuwmcAzb3NNJv2w9Ico3rOAEK2t+uxXT
bwKcXJQ+3ntyX33191U8BXXypnldjTpF+9jh+9l3hrBmalDvXOMt2gYGatsGiX0z
BAp/XQ86P6PhHMUuX1Q9+cOE53J6ZBbwF0PoeAtK8GdkOTU6EzNOQXNxu0Z1BXdj
7JY0R/9OAI/J00SgfWMn/uJW1muU5CgeSfwiVuWcdhofL70tK9zqFYS9eHR0OKiQ
d5iv2WuvuZqxb5kRRJgdWj70n4KJGBkARqUsqdMpuD5J7Wcg7Z9lccP882PsxhdK
VJ1BscbnOUjpCz3ZlOr9zhyIQxs6osb4ErtPZQnWSpm45G181XTbAxdwmscyT40n
moor/mNc4+pHOEnXzGYFl562HqDUG08zMiI/G9Zau6QFrzrlm/KCMYbzIpNG7MBp
1VILsSB0qHn+4hdq/FXv1gfj1VPrRd2KwBVCQqrkPclA+MR7yxaRqUYnfKfQBxNr
KZ4hb9rHpN4FocSnHUeXJraiaW8n+sz7W8yb+w0/g3UvEWf2MBJdAp9hxc9jdm8w
5f0tN56YoNwKVunZH6ywChkCRzmQWJn/WJzS+0Yl6dbTO1FFpiD/BHIL9Y8Xmgvz
Db1LXa08GAANB0egn9W6h4Ii8QtcNR8nzEs5JWDJAVsTIU/P8jCypCwFYcvS1QtM
b4oDnobjFcS/58Ia+Ucc5+BSWKaPvNBFOnkwULCxZPBLX5/dbe3Vf6MJUF50zhLF
XskPuT3XLJUN5HGmYnpDlxQjVGe/PnIVs4h6mn0knWmV9FQqmsoNCoKLdAjCMRem
P2P8ux5idWxJaWGc/HW3On3JBxDVoyBqVL9e+g+gR7rvuPGj1AI+BClHJ0tPee2I
9kZbnEu/TO9iDoconlTAiXB5XxXe7olvyqKITzXoDovD+Yq/o6F3oY9pJpG4q7NZ
XOyUo90gdYXKADdHo2MMRA3ISx2uocj244BWKaR+xFVRzxEY7Rk+39R9G5l/d72H
QSKDTSq7BEy967tPTWtTYbqsn12c/AqL6jE0zeV/PvE03xnLJzqztb+Hrz8wJa3G
djr5vj3AbG0Ua07maXTmqqmjRMEDaO0x78pVruoucb3Z/1P3NUvrYUxYpBTIOct3
wW6EZJ4J7m8epe9d3eoNa7ZPSm0tdg4mRBUrIirvJHsrDJMzujG6NM7/1ipdRoGq
TtgbCYvsnJtHS03BvVtZ4oI9LdJr+vJAefnYWsHdZYHi5r9tL30OAvNOygpseydJ
oE1OWe/Qmcp9odOq1GROmnSDeJjv3zJhCXQHyvNeNo4KAI1xWFhqHRymDQulirXo
NzjhjqzInEDb4V0Ls2O1BC4LBGFwbNfGTHKzfP2FuXxWxei7U87CIyam09zoyP2E
TkDloSOTyUVgEpP7njI92Turg2BNofSXWwzMKMYUD95f43i6Vp2znqFKBHYci007
+rERPGQ3aXs5M38nMwbzPTwdaPnzDC/olDBzF3bq4XHTYxrNx1kagUKInj5IXvaD
3d+ayNFXuAyE38EFOHI2jNn5jNsJBnWBVoC8VdD4mu9ckBs1mXKXEn3CyTdidqK5
h4+yKS/iI62+9M3cNG8SyWdQcYxkNOewMuKrqkCBOTyKvp/WxfUql9boj6ryJQSZ
Qu3axmpXmfODbFboQf3QBVGNrM+iCtRA8TJzZyvOt5yZnLXy7SWkBkejOAl2lnkd
6ax7V/DG6/hicDm+tVlhiZ9DxrVWfR8llRqfapnWPHkez7zEqXcCdckMVz6Oz987
c9vQpLWcadZj99bSKGBCN968EBxu8dHwhpxPUgc/gxMqQDihIwrNEqbbs01lZg3S
J97VL/YJE45Wy+h1RofVN2mCXXgsq8pIaCaMR4FtUg943ahJ9W4FX8yTufTJqnPi
HE7Nxy2P1cJat3LYRXKpcqjbP8CkLAcSOdJMXBrFmRz0jyVnLKPONAwTyNQGfJLV
mlBB9ZUNCfxsMHmVmQKD+B8Xlv0AaVdCwsicu4oueDkvgOCHH5hLRPiZHkeSdgZw
JmSUSDc10oy0MRKCe3Qy4dX/dJEfDJ7GIWNG9Ul8VpmJ8ruTcTat6O7+Lic61J0g
l3gVBtnmRLQzJtDBEkCHX/rsBL89AIaKQwQoQqreqj22tgRGngENhpxk+wiREeMm
F1rpWeszBZ4KXFlf04FjHBFfGMrAnoAZimaCZpZgXVRAU9fGd1MOx2ZZFOuA8yIZ
F69MrpvKdUBwnWVPbYIaEYwhBky3k3Okt4LsH6xKHgkRUqH+igy88aiBwC+L5BIR
+qaoqtqxHAaOhsFN9bFKx8i7wzv+mBpxFeBW4Sh/W/zSKEW7O0XXchgGHVACPvGL
TBKO9FhIBQLAp+4QX8yulUfdYVJjCge98mF+m6R1T6WM1KFwEvdlTOPjk24/rNLc
8/5e5Thdn/CB6Jay+9NwDl1Cl070jFTJ3E2t4VhA89y009WaWhraDczZzZrReeEE
NtUJdEclUzjEg1lCjY5nERthVytCoyJN7iYv9YYL4c04/tBP6N7kK2IcY1NwDVVq
E6FagFCRSsp2T+V53b0hG+dy9rYSyov1SKSWdHPltbVcOGwq6Cy4WviT5q69+IGL
Xjq3PMyfrPTJfK+FXtjcCYuhmBzuWLQeXWr0vMa6UV1pmDpOSl97l65ArU1taork
RXTOITRt2ak+EDRq1xt5DX104LjF5QAjKsMWSR4J1tVyqG5JOLUp6ZpVz8rwhThi
3tBn07WeF3A1keFWwc186kLsorBKeYcXrZ9azWAOIP4yjNJpAM1oc5oLKtJXqfP9
us7QfgUN9/TMs1bodN00Nrlkeu8W3Z/GyL3aHFU9vYXxEhxMNo4VqcYcm/Nr9I3y
xAxcuof1SlKvP8/EVuzy7PIR07rbDMQ3W+9tzlIl7Np6nVtbQNtamfG+ZL0H4AtX
lgndmf9GAou1ddMyQV65mcNvaZaEumrlDWuUH+LmkJbAOxZm/n8g5yvWTbi1wowr
Se+l02dJ1qCctvtZAgHS+H+IpeIDdDdMm1Brt19VRDzBZjt6eqWAouRDyYl0h07q
EbPWz3F6+58W7u2YGtTOHwmHjAirAarlMIu7ICHdlWI8l+eh8P6EXOkUAOZAhDH2
YVjXZ6gdkonX6qlEc8hKG75nz/1uPsPys3zSNwFO9xGu1J7+4nF3Y6IOgMWOAZKc
XMbP5XBJCTZxvWQc47PsJmLJkActGGE7I5d+A4SmVbBfwAIcq5vgvMDpVB6c3K0k
4uTaJ8GkvJwN5qpvk8BAM8UgbnulzBzjWSiXUfaeXTrq1gKSq73x8mLyIuAWyz16
gtsEkiFwjcs2aFP83JULWrKSYAkO0SbUOTSrS68BX2AQIJn2zzojKSaC8kWrNGPS
GulBPZEYeK1D8W+o37w5UDwlGDtf3u9odefto+mr6p2ElYl1jlLmms2OmpBeSSnz
pcsiGsJusKeonb5pbhsmBuO30qjqzmS8xxMWiaDOkItNj/NCqlTddK61DFImN9EY
RFdakQffKeV5PMuKc8UluwadgxM+lwt4R2N9OYhM9Cdn+H8xEleOO3cF2BSmKhpr
5F0yuJ+ABGazZZ9wc94p0bIjqbNLiZH/RVVLOKUr3yq0RTuOHuK749atJZUtifEg
zuzKmkrPXy6PWeIoc678EwGIuBuHaXBvvCpMejvMzxD6n0L9ziUcAoS3+JZm5TP+
KaIH4BN1Vm53xqAPeE3rAao/ac4IQU7kfd9qwoBMRVXPUK+tjCxAeZkpH1lzQ8jH
THqA1Ba2XCEU8nvZzMiGgETqMwY5saKvyCJcd8lgcRpS2tvq4FHhcWKlDo/HPSIP
fg0g20OFWcMtUio7PxndyipwR3lfh46xY9eg9tTvbShT2kh+3PA+ulAgZ0pL1S2V
HCX7+ZSjSVFWovvhu3OIkNk4/caYXsMkosXpa3M0Tf97YhlibflhPJT1YGhwGxUe
Ywnv9+Qjza4QFXJ/Y1lo3zom7tBR+h8H3Qeqbc3o1C6OH6Fp+Z4LM65Wfw/BHZnd
LI0EzVFvLQFg6uLkvyFNdU+g+63TdFfHFqoDZ1STCz53EtZ1DXj2XYzALB1AUwIr
+Fo0Zz/El2AjManssuL3OqC6nOJtN34uJTg/lgjuZu6UpoiucUHOqPKyXqOPzmRe
bywllxKnJjtmsu1LH3Vt4aExNpV/mUgF+BJBzbGlkOAzLjuKXNEfTeVGQkrUh1d3
JeUCivXv/RWnkK6FYiEna7MUF6gmTlmNUiBEAhs2aug0bs4ANaKfXuKWsBjfe85j
aalyVFKEISx67/zhntjAhfML1PgVLp2gZoY1voAc0OQ0ocvF4gH1BfSsJ6ntRLvP
QwALeNPLmfiuXtyFnAoIwZ5xUCaSOQaEaOuIYlUW82NjxDDxPraqrBMkeprtwl/a
hbGtKTCN/pK3WPpNq9GU7joruKRGZQRuNu2LZCMQCwz1cdf3eeSxs+Irr+MmfFRl
M6TdA8SDbjjh+HA3WLCycC/btcctw424f4EsDf3MoT62AN7TJbz7EadlBH5zfl6j
PRngmrypPGrKkKQvDEAxzv2YqpWOu8Q9Klr4wwMnqunjy6vVqpNuHW0h45jJAi+j
9uS/MwRHQ3RkqA59PrD0XXp0xETs3kEPsBRCfJ795i4Kh0Ko06/lZi20LRAW6Rfu
+l8fnnjvbda2pHJBxhrIYdN97t1yY9yM4Ew9z4pNhr4fJVl7ERaNd07WXnLT5/J+
hHylU+GwYaqNVugaQpxIuKm3jQ0XX/ABBiR4pp/DsB/UBrHoTR1MKE7F2W3KtuUV
QJKflrdH/rWp7jwhSM5Pa6yAatz3lI8fQEJGJt0VTpec3cq3Cjp8TUh3i4Ai97S1
JVNEpjAcl+XtPC25s2Xn0vHNV0q48grD9t0pL6mIn+yS5NxJIM99DwratEn9agYH
WMxJwb+6LhQxhVu8MZH35vtsftqksh1r4qJrjBXlxqFVAJsIZZWcn8MyyyWYgI58
++85cdISviq04RcWOpzuH7tgbWV4nmtfx7VvKrd2uPMIJEmNavvlI30mlc61IKF8
mb3TMTTCsJ1TP+ZgCfybWnNrHomFpBxd9Pi7IYYx6Z62+dWdeHJ0NVIrCdcnQv/R
doOCfCw3NsLqNW0ffanc7tkQEMupwIdp9P264/NafCkbvXKBWysVBnGJTc+54ASl
xo8S+80DLRA1j+zm6mGfDi32I7s+QVoIdWE8JBfOe7EqRKRNmiBFZuet3xCGb1YS
VsSZnDLfA/GRd0TxCrsIfGP/hIm2exUK1zUEySRGJlomH5HoyvGPyowRHvQg3m2i
2zxeltHryL9dWTOT4UmGkEgY6BU+KI2FAT8PAwAyim8QVcPUElBrDSHTT92UYZCZ
fgt0CA53LdI2NHf1b2eoRUIDt1KHbGpPvBbHDorMse3f2HMbDnsfflUJbrI2pxL7
hKWPuEl5+zD13OOMbE/Vdn9tK2e6so8dUb1YMdCHZxyt4bYsx9t7RqfI+n6Q6N77
g8pf/9IxxHXR/4Y9Q8g6DR5sKqAOho8eouB8mrbvHHJqckUJaIxT6TNXeTVLbg6+
83o8GZRPEM7C/WqZsPb0II5/Yql/0cruxvU7F0J5UPLfe+rlcn9NgqcKS7DpK/q5
gGy017UpDynU0cv6qPjYgZykpUHJESlpM2c5EiPXEBm0YtN2ZaYWZHKHHXHmM8l9
kCW+jjX2rHEg004KyqUKZpZ9gmXWrshQux+7MG2e8dTNUzy1dOZHwzJ4VegWiaWr
RnxljVtJhAXZiCVrPu8gooyjqE2uGo2Z5B5L5jLd8L5v8bH2USI/hidj6XnkNdLi
NCRQ6HHcQyvb95l2mkXlGeyHKyEeh/AYrmMJe7KpPm7S4+Ec8QbKsoke3Df4BbZY
TKfj0w6cot2Rwn2YfdN/CGSkA2E3P4+UCrAjMIGPtePY6zLGuPktGt5FKqTaHYX3
ACX/ugOJAQUE6DES+Poz82Qm1O4WcmZIxt3zJVMICpDsLYt8jD5RvoChURH4v9Ie
+SVl7RSpcpzAA9AWPcbTBPeZm2ei5le+Dti/wboJ+d6HxSawOW2TMzi4V9esAfZs
mBu48soveJX1dr0oHa8yvNvjZ7OBgtZ2i8kf75+3cuGpcNALU9cK8c0o8CMQU6r6
WI9vc1B6l+JHAFsBeAuVdCxVaDh4960ypk+MLbroeWdKzuqk9puuEa7xC6cHLXUP
l4e5vN1dNModHpM2Cxx2NK8YyWXmvwQGiy3tDKzYtKnHi+lEih+dljMLlbf3hYw9
Y7T+fVXDX74/v19G9HGB4AyiG6Vl2ReQ4QQZWLoLEWejeIgZQ8K2Xzq23nCFr/cj
GqQIJFXuKBzeI0KIu1VODxHWCEJvPNnjCS4QiEHwvkv9AVXUUiXXUb1ZtzKWI0dV
LAMUobSNkHDChyxauSDVdaNiGGjazEYLGaHKUDL6HzlgmVVJYDBLVHK2SajbyBXT
5ewd/ssQgH3ydSuq8tdOjxYSwnZ6uJi39+GlZkzvd6q405XfIWJ07mhSay/yHv4J
haxVjomsYAy3Rv1Nf4dy2pSslJz0xbzHm/CwL3qrblLVsZf5U6EpqaFkSu+vsL93
BRzeApMnyHwTTPwYs+blDqkWVsOCXUbHfi3+8aZlKNoURSsa+eGlXU/rcIOujgcf
w4SI2jwvT6YkvF+VwvoBQ+Y00h2cztxbcwqoxrZSShG3Etb6KrtXjjeCILODFND0
f/5U2iimJsoQ5cdwydZRHTEEjutBqGlLjZJXxSHnXbaKO4miHE9fmkwCIWJoL1jF
ReXjfYW2OfaFgtydp0Aaine2c9oTh92ih/O0+Bro2fVnnvgwln6EWokwiKN2XgTc
igvDI/2p38rbZQoesqH+TrZ9I5ERruft+9dFVA2h/pfd798zfBt1UKdLYupBSXgG
dJ8m4rhyXgy2Zm3KMRl3Iz+FHSSi/LemKeK9UCKXBGnlMqoaYcvSa05ZTFFFjeSp
n+PK1YB4sPfHfEDqkw8S8jCXEnfIR4qZyAfs0ppVQCFiIvNzOmKaXauLaYf8HYd+
Gp6J8Kjs+ym3fmXuvcIKY8OrcVeFKXkHCcbtYP6HXi2H95YtWqqXojEHyFr+OwL9
kDt8CgVDoMJAL03cLWvd4XhQROlIXTimHllYsdp2CLf2Vwx3gDk15aWrM5LQe+7L
RnlOg4t6gKFexRQoQuMmwuXqHiWu3xWmWvQgBYYTQ51Q2uVDLm2Lz3FW9pzvfeFf
K3r8dhsLop00j4w/MfjmTUzI68tF/R09li/4KXz8Cv21ePJXfoYGlbUL4RMg/8vo
+FRe9nSdTzhUVSzJbCYYZN2Qo05QOCyfbEne8rLWoPXj3sRNw+eOQTd5ti/ZOTyh
5kTy2e/elyyudDvdQu8ej/4D3F5vu9rRLDg0Bf6g2lquJm0mED2NuCvXGRfYAll6
uxhqfWypmhQRvIc7QQ3ms60JboRSMaO3tfR1BWGAqN6lgo18r4Vlgoj774AFs8HH
pspukBLCztEkCs1yqNm9EHvG8s0LlEgaiOMHEN1Pw/wfyxcPzzfdmUtx4nZXn3Eg
cH0IomaQEj8JToPT8g1kwg+XGjHWvOlLgHwwobUuJWv4whoEW+/p67RcpraaKE1/
8GR5eJeCvSgqJONbEv2qhP1cXvr68v6vD95+T06judhNz6EEb4WUlXZHFwaBDtqK
RkW1cBe/m8019OJ/RKnrf1FSzAuTBQlL5QNMlWSlcj7vofFJQeoUj3fM9FBFZvdh
WF18smnkAiGbxpa6nXxuO9TmqVpNfnKTnRV+tdU/unYlOeNerrKB/nvSptFTjfUK
igl9MQ4P1CJpP1piXRv+JyD0BjcDYsnGTLmu7zKdDjwEdIDNmvAJeH0u+NTzE+sr
Q5M3geQ47jNF3Yj0Mo5DtmXzC0R4AVftGYokdcykYD/tX5/81cZS44keavFhVdFa
gxvYKAZdDAu6cp67iNqHDTJj7l64Q2EFXmuelFIhz77caWGBsm5sY18hH/H0h7RI
y0L2xw7mm6hyewXmxhZJ+Zcl3jFV9AXgDYYtg71jKiXoAs0IkWCVBAG9fCFNc4cU
yodS+gRFPbphKOn4sooRIsvnBWgP7vx8dL+42i4XmIZpaabsAVsuqGCiLdNEetx4
UrwKXgmSzhF0VODr2MrLHOhdDgBoq5UIe3w/v7wfV93coNZ9xUmkoUJE1DwYNbx7
K51s3vecRrFBnBTo173izao+9Wvsk7M92yKddeQpO+jTYdhT1x8o70cJaXIp2dZE
PpL49vxtI20W4suf+nNnYayooqBj5dAtJNqNjVMdzy1vZv0By45ZvgK+6t0GkHsg
Uc23J9q9fm/tGrZTV4JTGEJALGmtBpg+PqnWZ2psN04JGwY/2NsZasSbxcm9ysZ5
d9Wvi8isdQ2as99TsMZES6IrE7F77dyXP1DVj/YNusBOBkg3JYpAzBXS/0UB+OTz
5JnifHjKKPiLCySf3ISa5Coh0y8FDDTlnZMFGOTXxK9qu15JmEvnMq1wqL5TBhUy
VcPK9hw0Lv1gsV8s0TZAG0HW2eGEk8AOgnqAswzVV8K8GskaPWlIhJwNCcGhzAIy
L3Rz8tbrtjQ+C53NfKXy63WjWlfgu2RjN5we8E/+vmjZIIFnWVSwWlLGnt0E4S26
bpeOnn9iGiYwJCjVlgPSvmI7mBTIjQd+kcOsKmEvs4O53duo/2nsmZOA0YokyBcu
B1E9a5WF+vVyki6QXqP4EDeyHU37wUnziKdPGdXrvtbJlacoazNso1x8ceb78tkX
2qKA3oGvzSu0uy06eco/8t3C2lRJ1UfrqeEX5gxPbLKTf4SNSE+LJPu7LMqOcI1K
k+zBYqnycMNxoi072HDRWa54AU13wbEuiQZ3+vpJiKCZvwpKOHo7mm9eKF3LTA5y
MzLljdVpo8ChEwj77NiuZKjR37PoVfa2+tsOBy3nM8M5rTMIVGmjyFJIEIuhZ7+T
2haq1GOJsyrXZ40DxcYpyt03YoWKiXFXuI8wqA52eousYlUWp9JDxzjxMCFcyVXr
8jzFRyDhyVm5ISrqvx3kx6KELRBV3oLgOT5uEzfp3tvbMvoj7vqkbxSA47XmUqRb
X+Fct1pG7K9TBfop0Jam0j1JnqcA7Of1iF5Abc7qbAStwLkWrWrN/ESSH08HZurU
tinvb7G+OQO1I6fYBz8j2KSz3dN6m2bXqOMEMfsqAD4P+yWKOK6TlyYlw/qFw/+K
XzbHjJWSHlbJrsITzYbgOOxrLZuHaTN6fHB9ec04wz/8AJgrUpPleBqzL+vECIjA
9t4sgL0hbzdMU58vumEKpHWUTBM72eajtzsgvo2gX4qSgtMa9xrvMpa4KbPFkDXm
iedPpUngrtXe3A3RQMjlY5X4IQv6sqsKQajubtY91IovMZ26G3MAE1WXY68Q2TkS
M60gvJ0LikOs+ziyGgsohofYymclYIYKJHo6FBIp+uislcXZYLKrC2EP2HEPEllp
YzxAsh4O0CXJn3IIwxslzabW9epm6NCT8MjS4NXo/Uz6TRUw0CPH4D2tlP8I0zTg
uWbO/AovBkJX8Q0m5kqc3g39okgZW4OG1UE3NyyLn0uWFa0s6Yebx2G74WTeCtXE
gy7G411fbzi9uv26Nm1IVFNZUogUnzeIatdTfsmD367njuPmjYQebQFJ8xN9k2nG
Mhi+lulOCCSQa1wfbls0VnE0aU8QzwjJlb5e8AIgxjTGs6yU3+KyE1Qq+wABFl4b
sqrvoi0Nt+fjEVzRW12RzoMnjVRQW30T/CC0Hk9FL1IupMzVBJdAYG7ekfb7hPq2
iC5unxVtxzSGAr9rRtXyIzUrUM03PnbKCdSWrA4HeFwPOqjlvTC3hdLRth9fuq+h
1E+47zO685hf5TfyR9xzUwW61cdzhLR8VCNrm+8feXjcPKIX/55WXCBRUzIaFYuI
/1K7/jdY+ejNiQtBOyCZm6Cvh2rwJYoSv8mfEp7K9WTQE96QTdqsbxA55wYProGT
6euaPM+7qJm7WZ39k/cv75/5urve105QQEmYveHW3AaQOVjiWgQWtN6jTGUghIDY
faNMtq3hfrZ8sHCuUX/9dDZGHYW2nB4krwfQ2IehmkhbFq2XDBXPMvOVnDLPBX1h
lWh0wSlDKbntzOs0Mgm5gGxvwqbNEkGXxelX1UppgWDWsJ1B4B7igP8WoRSRDZM9
9CkQ/o67a/rK1AgpyDAO427MaA5fjTn6/5zR2M7SUOaUuVIX3m4Poq8kC+I9weko
SB3yIxJWvgrhg9A8k5d7tcY3sGrUtsJevMgbJCwDknQpBuH0lKpaIBepq82CWyu3
NpDJJ4mSM9wppIE4VH8dcRXRIUhRqdpAMwVfdVdClRZ/XJsoAlDvqmSVKb8t0cMu
eucyzLNsowDvjbw0G0o+NRTfZJGUOTWvucNuleMh2bQP3TS42jMvl74UWIHjjCmp
2aUOb7Z6Rcv86T80nBFSIHIIAlGdD1R7jykaK8Dq0geRPt2+ftqNkNPjXGsx22uk
wiOPzBKNqxIM9qHuldY7LMe0+8Z4CL97Qc2U2q3fkZNdR5X/jntzlt9uTYAf9Mil
tu3k8bvpeU1/X2ZPHxLDpw5dR0fqjTpOdJxBLEpuvLkvZzK3cDzn+NtlisAoBm52
QW426RhOJond25AkZOlQgW6o69xCDQ8VcZEKBx4RRDtArbbicODV2yAT39OS2nMe
X7mIkQymK+kKoKD4qsCakFj3pSA3RTSGDaZdWP5p7ojwk9K+X9h39PEpJXFwrV4L
gIa2GKPLRHj1YEz31e+Njt3Q3Egv+pHq6MEcXD4gS0rItPWbFOTuLZitXhcB6s/h
H++n9uLrC/+Y/3m/qWbUZUmh3+DC/sRShRzNFBzo90BvlflSuRkqbyPkohdZ7j7G
KdLTN6uqXcZMXP++77m6m9TWiu83IOgdnYQVX5zRqopAUNIi9wxYz3zWAzbsjLDE
pYLEDl9ZFFUfLkYw5wo2tbSExOfbISFRB31DHma++fgsd5Hahpdq/kQ4Snoq8cPs
nYkCCP0Vy14KNuAlYypDBShhTwx6NDt8vlEtFJQaWORpfb4RI3oa0lWdtEEqQLsP
M1t3lvjbMwk9DCziYbbLHLfAOzhoEpwH9mg/8bVSxi13l653SO+iV1TcCOtBK14n
RQpDgF6AJ/H9nr93M9bgnpVXJMK3LukuM7NpG+4o/L6JWWz0/lLTgFcpy0Bv/2Hg
fMlMvglLL4i2OeptFBKyXlOm4Dr8Ul9Wpmc7hp+qZ0+PgBuvdnFimPiJ62/r0SK2
HljMizAeLRvN/vF2VjQALphljyx4ix1qxS+4Cs0nV6QGMILgdMk1269IruCR+zcZ
aLxzx5o0dJEEklVL6TEsWBIlAunIuMjjhtkzHz2kE9nJuPL6nKPn8vs6FiCav5Ly
oQZjnZWn6iszRMOZ25X/FkJs6xtqG7T5TFTgHqnwJLml6lME+5p/RgQNGA7mj3u4
2tKqWU7zwmE3kv6Iu+xV9Kc8gnHQ0FeaiMwEoytpAScOwo1Pwz7L6ljD5CEYbSXQ
iuEkkfKyr+idsCUNTdHj5gGqwrt9K0J1n19VL5xcEltlj8rP1004hYPt14uqEOvL
dYdEVJkm1pn2gbdnuixYNide4ZjLuu2rruKxmwgBDqOy6GolWBvs8lCca5Uqqeta
gu5yyFgN+vW18uwHb2kgWM8+CwjOcfR0Wh0vIkVGb8zH1Om17OXDl3Z1hFAISaCH
bfbtqmZsK3iObueeF87ysCKrhF6rfXY+Niyu0u04HH+107YBCNaH8OzGyK+JGpuk
5tQsp7KyF4/oVJi9D3KqkTEPioZhv3O/KbHPgewEUeljxREGCHPFSm2Gp0LgX9Az
AmMXnC/ofFEbjAhA7YSf1TJ4aFcnrQNos5v0oyZXoyn6TJkNoQbnvgk2SMpPvNVU
I1mtOe7Cc/dgXDMAHxNoBbKhCl/cT9a/GwizrP1SijdicAQuNSLxOS2R6Y+bt3f3
5lUDrlQs21AZxKxDi76+2ZwRe+jIZOfCSkDd093Fw70fPzBitGBmr5b+9THLM6Js
eCT5Mk1jxS87F1kJ+preSzde9U+jfLamFrI7GUsP7prVxRHfBwAL2tEf16o1z2m0
49zsIdUWQWq2wtZlEpiVVkru3OyJ4yAXN1aQqE2Qq0McOkr1tCS/QK2IdtSzD62m
Qbe/dGZVqufcx6DoAgqbxJyNa1bCRPssRkrnrHoEM6S/jRtj0pTJ8PJYIaJtEHmY
2OekZQVXQbuHo3pNAHkvhi3SxvVDf/H8FQ/mXHLUGOyYkWiarCqwBRTmJX7VcsWb
TDv+wcedN7rnfn6/l89Rww7B87DyvZmgkZ/dAa8xu0UdEHYEcZPbpjcoVp9d+Qbx
/qnMgCCvlfClokLKfMn3rrTYKu4ywTYyyKLYvFB28FzSgKiFyKIZkuzVGI+p4AVs
3XrTOjmbfjbRC6LbloOQJqtdXidRlhsmp+ePAQ1viLtiLW8DYP8Yzzyp50i4iYKa
E7u2ef7hFOYGp2M/ab7+xk6tLfHYB3EDzO17UeWLsDmnzBgE1TQO9ia8R7g321Tv
Vd8i53NCoFGnjc07ChLOZLgrp/j7HLbH7hPXwDYTUrCVBa/xcp/bcHa2T3Tm92AY
LJxYKvKcC0PnR+vGVcPExMvt13lgMCL4NNyJV6TOKxhLH/RlgNriKgCsWxFhmb1I
BTjk9PzhhCFlWHPf8mHheNcqWgdvlHpDaL3c+CV9pMVFOkC9IgAhyfCf90pRdhST
iT22ndBA09LrpmdOjqb9VJ++TU3kmy7aYwRARmPmOTI1NeQuE7im1pe9absbEmCF
b1uzPaolHUzWFGz4rlB/bqwxLrBHQBcabh/w5zJ2/jEwBZ8OsUnA9kD98AMm/tWU
8rt6z3//ALsrX4GSAOX6E0UGsEEyYgz703Kg9E4K99fxHxtJJjl4tJ82sYLJmOUy
BdYo0KUANO04t90qjbHiolyoyocHvkAPfmP4sJFEm60sPhkR+RmaLW9gpg4I3vUv
WGYxPaHom4IL7dQkvL/s2TH3+O2PDJNPHw87N8FU8fUL+Wbrb4e93SY8rjb0AvgI
vl3y3ahZFovqWyOTC3W82M44VIuGUu+nydF6/08+1YytIeZdHVebnjxkmME4vK+y
ot/p88Wsjlf8xVwDB6uCpdECjW2rdWv7qSgp/9oXXgpnIsWXsuD0PqYJ4BgBTdha
pkn0xE3qBtTlnndXTuvlS5UnGA0byt4Gkd1ZjWVMSAHZeKwJowyriq5HKF8YA6dw
u43B2pgIPtPFmen62K6+bwW6fXMiwTCq1FGJBWatfGyrydZZNqxic6ASjhTjYa7b
Z6kwz14/7jJVt9imc9d+VmpJdb1HMlXQ1AVxrxiEcDJQpiIuGNTBqZLNGMJetlCP
jW5QuxcovGKysAf/6PHs6oVxspVb909sncv3tRj2doE//cQ89n53llM8SzTnEWWy
W9P/JJTe5viQMXQf/RrbPx9Y8EEIR1Q9aQIMEiF6fHAnY4c1euvonoAXrgoQ9x5L
Fq2txX81lkEdPlbkeN/D2vefKviNhRrt23FDx3gTo6g4wXvGpS5qx3A7g74MYVKc
WStvOiBoDhQvBhEJuvPO1dWgyiUYIAc7SmVVjINbkZ3Wpj5wVuPRzVv8+Vb8A1Ei
s0sHUx2owZ/xhT+iZT4TR++cJbIl2dp53neqzJAmOXq3U12KTCnZDdbG3xKBUgwa
vlIpJQDEeGlLo7ry5XcQqXeZKMkLYVnbtgvKxqcxNUX6tf3H00IB/mKX8jZckRTj
+ok7ehkTT5TRC+KnQrmgMIyls4pu9oFAUOKRWe+rS931k7oMpJuqGV61X9HbXr7T
SGUAWurHGhTTd7KHjcaulHfh/Pqpk8OI9yIbTA1GMTao2ZpHH1H1TMkpnVz+PWJ/
uAEWRvDiw2v+XQGSRkh7x3B3xXnw2XoRkKROJE9HOe+6xbxLB83vCglUEHT26qu6
OR0jxCcpkqMR8dzvJYomz7sKboumu+pL2b4/rsgZnEzB2b2l8nih+d5K4pgf4e+a
M9kSw0IXPa1AWAhTiPClfic8MaJqySUchpBnIxgUZaaM6JC1fInbdy3wBomfMA2N
InU/C+RUayLXibq5M4ZCDJfPKET8UUs144mLy/ImPUaAJS1dgGfvFSplGxGQVE9E
5cN1SBuaoz2FZPHbNVwUuSRJsHdBOkcmFZ61hxXCXBWvAMgeHrbtwOXXvudO9j0A
vGFvrFK0etzPu1XZejah6ovurSoBqU3+da9etKmDCrS0MzugCsfkbLGtqehtPxtF
hfuQeWsAFN/xvOj+tJbh0L6tlKuYgHEsrGMsooTV3Zi0aJh1jUoNO0UoW1kjmKfa
Wc6ZA5sB9Kc7OIfIOq/xwARcMLmdH4MCTbBiv05yVWr5bFcJ2fU/wwlSS7rAVqWV
jSjXxRCM5Qxxae8NIAyc+OhfSXyHCwR6lySuOtwVw5XweZF0p9g6533w1khQpVkY
I2XCOXpovqj95rp1rFfWojwZByswG1LaewjLPdD98fAdqAX6j8REvFjZNfeAjn2Y
TR+ifhsg0Bpj62hpdwjh8z6zecTr3eOJXyygajX+hicAeo5WmhjHfhnvJvtkKxMS
Ciwl+mr9RAY0dxOIs14zg4k1JZFLTtjInmNTQMXe0ZTngIaR4x4dRahgq7/TC6xc
W47xLiLZjU9E0ZAw9K+52izXyIjVCYlARlaWrjKizS/GGW+XWXRCDTu2xFPH+jHA
vgpRv4x0Wg5YgoXpEPceimozmlpG1bC30E8PDOJL9wX2Hjc08kZQPh8f+npBnSin
Pj8+VNrih3KniLtfkL8wZnWoaQJLymFhGNfDxHl7QmwbnkxwopU/IqyaaOur4g0H
4OEjmxHB7D7e1RrmfbFaLIo8tWITHitEclQP3z5LiBy4OVlbhKtjJ2feQ+hFRYsY
itaS/S7AB1Ey2c6DeQAJujHwqGd6MdFfP4X3gDMfuTqomAqf/NR8thKbFTCt1STt
QrZmk3E6ngfCGyP/U/drzFPE6hl8alcRhU8w74aT3hr+5XUPwYgO35lF2V8HQNum
tecBBkhD8bNUxpSfpiJDiu1O6Vb2I1JdYMWDvwoQ6xOmf3ioY4rzPY7Ljcht2haT
n6fjN9eJ+J8Cb71wz2vPX4ldSnoB+MSCTT2KdxhGXyoqSMQMfTl1xSDY4zlxyZ+8
Rv0mz2nlqTozHOkcERFQuOlShI5qAbH/jwjMoAR0AjG8wk6wMz+zK/k6zceOvwvS
XJsWm3ZYEGoQ1p8+NalPPRgmo6gcvfExib/dXmxLv539eaX4f2FLTY9VR3aX0w4/
NEqciCaJqZUdB4ICUIWmiWf7WOS3JCRemkmGDMToOjnyKHCUS5opAuVoIKv0w7dj
VvSIT5VXfyB9QrnhKOdHoWSxTynE2jagiX9D8i5wL3Gx/JrR6vyt8W4r1lQSUotZ
zDduHSf8KZYrAKpXUXh6mnnQIbiqNUqqtN0gyH0xw7LiCfdDOxnPSzDknc01aZdO
WD6e6EW8b+H781tMED9SJ7npBuY1HQKk+StE/946IOjlDsneSMEsrc7qxPzlPI39
0YIaOxOD9ugkqnFMGx6xt+FBT4xfsxA9x4+OXux7xol89owRw/KZH6itLQ6dDeMo
tcJNB/yldyvQ6Xywe2GN13EQmNjiGZ9DuGr+TW5Nx+cK9ppIaX71XAavSokXVbWL
LkTlNmZeqlVRww+HWLB7sMBywfdELBX5tTocwHjWvCxkpuwUkqYcGrs+vGwCVhza
mGqyyelFiRUiniz6wgDqCtwfGv+9+p6owFX6RfvKWaip7fab7viESBBd6Ty+LOs5
ni/d042lxsST6nE8jKnZ5bsi2Keh871ncIuCno6rR0scgDzLNIGvpJ0jTdXYZ8YM
Bcb2HIMOL5R2v2Uon1l1aHR73T9oALlGDhUe+T1J8JvxV3fBwgCXRiK1wj0xRgql
8hOzUNGgVJyIYGfBwtyN9z5LbRgB2SiEYm0WsVw2sA1qP2BATmcqsRR+H0t/1Twl
OUKRHr624iLQ+xUVloC5JgHauTuvLIqQb4mOOWDDCjUQsVEIt61jFqSughV1LOB+
DQPq1KUNSAeFRYVFpt6m0y7LQKhLqOlxIhtl2QCB4CCZMV3uztuUleV63JBSFP96
ijSPz++PG8XkHfZvwxj/20OEtCk3Db6/3eXREaSJQ9eCKXcw6iW2eOBNN0Er25FQ
Vrv0+bWIeiJG4saZtM9DFvNCIkI9aGvs8yyUf76Hho4iSkov69GZaEccVS6Ia37u
kKoKm8c99a9hf15ejxWuIvE0BXvLzlV8vkqUXQWcXroF9A2KmmKXr4DgqvjcBp4I
RaGj1lFbgqLq/sNfhqhD9pFc40wJ9I+vZktAmC5mj8w/0Zpa8gyew/ggIv+//4tq
XtIE9FWy5Sany2Sa3cS5cwGGaNMxYXRgIXaPJw8OwAKKalPEgK1BMoh+lesF0Ogn
/loVopjr8++vKDEQLgAdFRl0flqZZTKsv6OFTp6PTf7SR9HcMI11GE0Rhp6W4M7O
Pk60bQvo7MiX92vr1kNqWg9zIbwdQkAlUGiRANbmimxJ1cmI6exVmxG8jKGeix2u
HqY7KjTdpPc4O7K5+G98bbDnlALo5jynOeEgBUQQRC4Q9b16VQ5kQlnHnoAc8jVv
wTD+eWwjd10SWZDQUuIDuBZcocGIwfSYs4S5W5/IEp7hfVEYdLyaFl3RhiWENdem
IpkGm8LW7Oo0fG+a6g0aiMvbC6FjFgFJuMcdJcLEuJ8M7iVJ/VgyesDWyBULzcKv
EV0G98I6cmdRe/s7mgeQJu+Aqc4yubennjaOGKQVUvLos/WNxv26oXBoteNGIaok
NZ/0g4CBWWJjWftBTZJYphdsrpKPnZAXg9RWBp8yMpIaK+aMqluqTceFYTDG0Mx5
lH/ecX8mlmdWneTDNvjga+IHB91OL38vKQPPuY3gEmSvXwrrIA/xE+Mt4fmsGReD
bBjRlcbssYQ6RFtk9jqVB34oexk5Mv1wJQGvsx2DlRmFLY38Q3lrfyBwuplt66AE
FLtTAgnpaC0huSiUS+MYBnTrD4bQ0PErv1Ro10jjd9FycZihWgSKyZzPYM6lGEZ5
jVnIyl30oT/xzqp+RkBYiHTGNiOnT2PQDc9KNcEZ/Vz7RoaLwTEXoZo7fTwKjicK
xPMowMLzf23gOxnj4FJK/+2q6ihqesXp/SZA+ZLDY1J/UyQAN8U34AOgLkPuZIZp
nKhkazAX/yqfzTCHamyFjeHa9uJodtk8hVfnC3fdZfabsn8+lIHwMbAS+wpHmwG0
g/GMn9AfiACp/dS6GofhbiUI+beqyPLRLP3CwFKDmdGjiP0FkpcieOMN/DWF4As8
ZPu0bCEH+DIHQJt4812dcpEL3yXtev1/0teCbzk0AwQ2LjVXy4Jn/OWsWuyVEvZ3
1jn4/BPbVVPl5HG4xHQLeIWg/d9bm2qb/V5LZYW3AZw7kqRbqANhlKeT5+TtxUxb
qw7RfFjL6lMplQSDvFzvQn5dNxYN3qwETps3mmq/OQAozzFCpm2aMc+KzNEiHYGl
jf53RzMEzPYDDEvmPRO6cAxKWYdP+4x0S3hn5pU8NkfcxXGlrsmd4kH5htkP7zrY
0txV2RWau9yNvVSeUDktKuBVN3NKfL+SZColAIGlTaRU3w3wRE6gsvnX4N4Rv0YX
qTf68o08QUC7qEALdz9r82Orcn2hpGnr4CnUUsPE15u+FB3rnSz2U/sJ2U3jasAt
pQAvKCDcGbJLvsmevG4lVTtVphWLeD2EySr9ozN7f2PdLUTN7nM1b6AYZwmDjrt7
MBjXgBOowarCjf9CNzhOrZdjj9SRNjYu988ZEhApNYkAZo6I98fm4kCqYYP3IcGN
cFdCYG94PcyKtQY2bG1RvsJQ5BloAqZop0SQe+pm9bIbKjZHdt0sXKb7XiKSKw7D
GIZJKbqlwda1NIA7RgM4OAqHBm61BavpgtCzJjfEOdFDMLyzDzH0F++XHvu8yixl
qOypxTsFmmpppzA2QAT6pevfcncnVF4YGn8jjbZ3f+a6xwP93WuSe4rzrqo5KLyY
D/QZjkH5Jm0FmF+bVtQVBeVwsBWaL+GQlgnBwOh+pNG+NF4m3gfsGYmgWRXGuDF/
B1A8BJw2ASwDGa0SLHuwK4nRwWnZM4acqhv22I+n22h7d/sl7QzIOY4WAc6jVKSq
j3XauNEyerZNqzd2sh45b8zFu9Cha8EfTG7Qd5Pwr/58tIzfQ9k4i55nLf6B/6sb
klTGrvyW9IEf6OCzFbn8fMv56qU8Amin2FgXC9rEmR8/eZNDUtkKmS1uXnZiyB7r
bjL6deN07xlDDFi69tmtV9EIlEAxmXANVsemToq16LF04iU6/hAs6zYozRlk2/oq
8QD+jUD0dSSwQHWNhwKa8XS2GRF7OkJPdVllqdiRoMSRZsO+KzZoGuyK/PdfzyH6
boY27O804zF+DQH7wtchoYMV0Q5FvwS8TeQnuY37/vcRkYu89AuZZy73b+rypJhW
lLa1D1t7dUsCSTohL9pMIh4fwAtRLqzMuwgZAHd1W+WDxYEwgCMP5yksNwXYu4uA
ZNcxPlT4uu+oDZ7sf35mO+Mz+1XheWVb6+X0+kAIMd6CgQSr78jLrO7Bb/JJa+q3
rWiDAlC7Vj4hzgeQLWm+mcw93WuTa1/ucZtGcknEW0HwHlASmVmK199/kBEPtUXP
WDI5f4bTgysPlXEdrSDuft8qhDwbN/Y6TDiIj4O/ezh4kQAQFbBN2acTMbDhBM5a
V7f5dD+mrgfc+67vBS6UccrTiQaflnCJsYpxrt7MnEVvPYyje5lzsBQw8izcOpY6
DgZtCniekC7a07jH88REHDu0XQdPhU4HP6xV25wNc1L+5UjNoUxArslMkd/C1s2h
6lhHZ4Uwm/D0WMoEk1rpJ81kjnJ8vlwdPNpyJicwkg4mNJH3OHfDJyVQt6ApvbKm
YU3D5LQN5a/hRtp7uTRPegwKWtL2KnRaLCC+IHkZG8Oc3SIjNyR090f9HSBG3gAn
kZmY0SdELa20WXVoBXzXRDeR/fenck/LyWLiOZ+Co6t5gaIAg53EUBDeH0fnAkHu
DLcq7ryt0eztF+OfJOKO1au/cJ0FBs+ODiGXhhmadJe0JQrioV8pRVW8Fp+WSSGd
NrAoHmqzBrf6SNPg5PwHcsBpodY6e8Wg5KOODG1e1hqmdwoEgEdLhWMimxDrgX4E
545ivkYkxt+JxaVApd00OzONBBUJzahiSXqHbfwDQhsLihvZjzXJIW8P5Dw7OADH
nKkmF2PvmVQXz6B5X/he3Ik5IX8oPN/3UscZ+dXZQa2UmB6LY6twXFLnnhAGtqBi
jmcDctnRHOkqSf4N4vmk77B9cewgxO0L/oeaS7F+YQ1P3sNOHNfjPnOHsm09U9yj
+MiJCD1rcVJzI5RvP5Xc9sdOwO5sBcHCkFh+RexcxEOsUMNVJ8AD8CPXl5qAnhZV
0zLLyd3u9Lt5Bf9f9H9G1nLc4CPMGE8c4ZExfWumakFFB2ufDk0FcHppZt41vfCT
gFMksPJwPrVBM+ZflHFjgYlRtpR6AD4LmXiOEZYKNb2BCNkS0LXFGNibCK256jig
6SN1fSoIJptOGGeaRZsE2YMbdOBNhEIL2K5tz5oAhwCzzCBUg5cX4K71fQKhTueY
I7RqO1QZ2OAVoxnITtTpXHxRg88VxBFJQ4t+nCxY9ppb1/uf0ub82+ft85V5ewPC
qiUT29nqxlZkjBMxqb8xsveo0mpw7MP6UF5K+jlCtdlTNwTyLrVuHhURz9RImbWF
10UpkPFuueLIGgADSxcrpjRMmHtyKGcbsltZNPQH/JV+V9l5Kmq7loEO6y+etzYC
tVKWAKDrVg+qIOMfnar5KhgdFanmyczq8k6C1aN15yWnzdYYiu5H9vXA1FaB0USH
OPn8O040JuX749Swh5jcpenyJeSTPEIAN9GUi++kUJPqCjU1MJAf+zSgDUVIvAjN
ks1QgpxEiJbHcyQVLATVcGoUvmpKs4wGyFb+UnzQhZ76EOTXqaPJKSoDzrPgl53i
9DYTwcbdWE62GO/GbYWaFSTloQ8y0qbZrieE/EZVSiy/CQWniYjzHFzHzAkzUV84
R3jbzPm5g2je5bF0+WCy8EVk4NVMca8ugCNCh/qyd5PYxng6UNrvnuO1vG4tEikA
a9st3lWlMREoJ1Pk1ruqHpr1XCynQPyx5AyuXfNu1e9AfDDmrmrwDum8erGnZU9v
AOfUPY7jv1Cj2Eyuisk3kViA9siivheAEHjT+km4M4qXYOj4c87AQOgfp0m8xnf9
D57nCeQZRjko6tRp6psFcmh76uqCmq1vH4KecJTHe9mb7TxXGQ5+bF+/v/Oc3dug
TfgOPREXcpHVB4LzoeKmzqyC5AEoihDpBFs4M/EunWxYe8ExjarD485r9pOj0z8B
60F3/LMiKIqGJGSOkQ7G9HIe2noAMNRaq8uTcmc3DyhWphpH2s3vYWsCnbidrseP
w3B3ioz436lpI7FjD7aoudvfbluyIXQ7zfKZhbkMt+dBbDpV/vKixhT5pV8gOqVl
qFVUVxgNgmt0OYCvQRyiMdeuEYFppjDQ7XwYGSYoLDu76UimQuFjTMbWXWxBNTb7
vUHTV9CFNd1TJFxls2qkAqQR/f2FJzfamynvSC8j/NO5XqCKJ48bQ8bya+51mTz7
ODPnLslCVGoEp4L/jzXtnWc0pwNnW/e9NUdAhw/ydVe77NeN1bEKOsFFx/yecSCm
HmjVukV/eDdosObt8i55yJ4sAISuZEqg9+p/JqmoGP4bIxE/ewoSRIARCjokgIHR
BmD9gbXwtLLOHHMfwIZalBXWC8oklxBrffynl0kSSw7Ha+loGq2EUsyEQyuy7X9X
KpFaWaYE6uYgOTJiTPmjG7LGvx1FolJ5jc19dnadc3tWN5uEZxceECd1DKs3wyBT
5VcyJwuoDr/S5pwtmCfxr9+YM6arO2quSuuuEJVGF8R11Du87Ij3CkJrqhPv37I+
Y4Xqni1LYk+R66iiATc60lPG5Tio8YIC+BavlDo8gbVlrlyWa90WsvOskSiLJy7O
UxiKAr7O3NgqMmx2PlA26vWR5eNyzWCOtY4HGOdhBx/O/p2PjZaVwg9GLjJ5Slhm
5XMwt+Pt5xPHHUYmhgKG07QpVQcIyWE5eq/wSqkybaBsKwDPv+FTUX/kGj2ZdFAy
D2RPPzpaOrnpsF3kK5Wsg211FhAhL4qbKpuPrUkld23KUoc0h6ufN19I+385pdyU
4b6KHo0yubl+lF3Ah4Y0lU6z1CTG+zwQ4Y1KMvge34MlZ1v994GruoSzXAJggYkZ
nIP6WcoEe2iNozjnhpn1M+0ogAavnvmQzdfkR3ibIEdu8YlWApStvJF1B+53p4cB
RWj4K9W+UubRj84VlT4miFIdLB3N3UTtlXcZEVSAAGF5YHXDzOEXN/a32go4CQFy
UA0B/m3wVzoztt692isEzV3j9VavSwbnw1+pbhKiJDalUt+gZhrpdAEcoUUEK1QO
23wLtyW14r7GnZKQl7cdG9ATKuJN9JxDKdFHHQ7gT4PyczC19lSzawKBKXLF3f4Q
HxjY75FLGYzJ54EgTB9P6dEYpX4bhOpUWRg6AsPO51EutkE+eSK6pTbVlhwYTftL
BeTb7Y30JgR2DKAkOobjeVe1Q03VTjUbgb0rzVPQcKPrhIqP8cRbGVplbuToPLdz
tyYmgGktQJijROJuw21U6GJwLoR/sxgFQTku5dhjfxW4Tynl3ZLm0KrCukZENMKe
2pcJaHgdOekZW6z9XpCwD72kj0wslFED7lV8wodWa/YDNFduSJkAs+/LG8EATEz6
E6c89mSAmkyK+NN1rqq3PwUtjvQQxbKQffpb5MflT6GqmwEfCdBfESERWtS2ktOW
N1evxlmYC6q30oIKtQ5O7PblenmDHVMcSuKYYo+QcyONElrKvU+HQ1m9vE21h8xs
RQIxwjYOsznrjVj9VlIJC+seRpz2l5X/hsz57nCHah6/OfZdhWGUwWwV4lRNbgND
vvPOzqPZny944v5lf21giz9rutlJ3klMnVDG2kKNikhhLy7wXTj+PKX+ElXzNDGJ
CA3vciLOzV5BYZ58jOzAzAR2MFq/II7PzSoIDxIPXR7A+f0rdj8TOE7rPsz5Hlad
93/InuPLuWRRCBd+RnWq1zanhgi/O8ckbHIVN0UrjAk1VgapCHWs8rPs6KujjfJy
cRq1Cnaxkg9FkNNXcgDtCT4vRSLHj90+tLBUGOh8IkArtW/IiVEhGQ0lg00eCTpS
9JADkBxqO+NYS372xYVwJ9GkvJLF13h8W6sPkf3J6JA5AM2r2OisbnEIzKtsYlL+
rBamOhR2zasmtlKQOxTG1/c0oBdtZe4UjwlPl5VJS/Ym2SQ2sqwqUYr5OYO7fehr
QdYYYuwXQi/N6urewSpgaYd4Av8z0horcY4j9/ZBZWs1UmMV0TRq1KGTIEgiVX+I
H2F8K/4DjW3TIQ8w3so4wmxHatcn14Ecab+4sHk6WiFeJ8r3voxpkgq0F03oeGvz
HgGkw9kJXiSlzpuqYDUCLWSrX1uQk95KJzSd70U9oRtVnW4UCUXhORxzPu9h0IaR
i0jof28yrU/2boP9/gX1d0Lp//stp2ayd26KM8zK8keHUV9MZ34E6RlRamGZalTs
YJniLn1X2KiXs7LyhjPe0fYSOzNqg4MMPkB67X4i0dz+UyNsob96jIimbutGPbmE
uYzznYTNRtwavTtm16AMzdwDXLJbv8mjrYs/dAdgXFRyd803B1LD8uVZiVHCRt1b
vH1HpAiw0F7TqJIb2pUlhXr1qKnfuoYbNCawCTSPwBV0ubJ5g28QZhpFyeKBHyzN
hx9FXRdOrxGeuPx/yDTZBBis2kKfzG+TAjLuJGZJCAnBJ2PYEXXIYAs47aTAyUAo
hlryXfFO0PN3rwvZX4Eo6pt3yYCSS6E1WbWjLAF0OBSm7y5gpK4pQQJqDtbTzJto
QcFDOaEIu/D+P38LqtF7j6IyLNy2r1Dtgif1rZJSYO2Yw6Byn26mGIX93Zdpxoda
RoeZfikSd4JWuBdahly7zCGwbJV8U9MxfgStAdwso29Gb0jgeHtf/gfwqmbhlQBu
8qbkWrxgOGbsHFruCChWrZ5Q9/kTe75xH7dy+x9AiPPwCgGmMnJIU31z6Kx6Bfq4
VdJu/kUA5hwEsU8ac1MNNbREzb2HGfAu+zNE0v+lrCqAf36Fm5HT7Kf2LE/69pC6
LlZCWw1yDvQLSndgDEZRUXZ7PPEn05fMReoCqAwhQK+QgCgzhWt2GNvd40aqhlQb
kmCqnSQA9aSzKawlqDq//7VjZKijHT/+9WixRpIQVLNdTdqRTDdSZFGhqCO49go/
aLTBBuskje2glNdal4017nDhElyxPLxRSXdchCk8/SsO7nmZyA5Sf4iTVhozfFp/
5RMGGRsdMZ/vlea34YF1fbIGeM8nbLha5BgFa7v79DLaFlEgLQoFF9v7HWFGCz/g
HMXCtd5BNGIc01A5LTMiskxxyfoy0Qeik0DoM3lXZnnpZpXKC+O1v3HCtylLcmtA
D08TF91yUFKBFapyrxKB8DBT3u2T2IEuWEpR62S5wvULpPM7WAOGyi4uCMDGIcLW
12mmNlSvqoGqNkNvdCKnE5wGRzZVB/13vcYAvkDsDBsgB/4M3GfdH/TEvYBKlOyd
CzvJi62BdeYEi+r/OJiqNYHUw/nAf5mE0txHUIu9KdhhFBFaYxALeqK/XBRSXp1I
GoXPa6uQxkmBbI6+Up8/kSRkY5t4yUsdtjPhmiXNEUb1y5WB1W1pa2+wTKAd9O3F
GsAJ6mOAikKVt59reA6rc3O4DZ8OBv/gD/DM1AMK4uOEviG/AHWWPd3GH9H6MefN
WBWGDuXPR4XdUwGBbL/elgR9CIQhmJS6U/sT2SQj/5u0fULR/h14bvoqlxq4Q3e7
c7WBAXAwf1jS0QNChtOyuQw2FLxqZ0M7w98yUjUXHWk1y64Au9Zue0KAXm/XF49/
HpXA3S76mhhXLLqsxivX13Ek4l9RyqdgQ0HwchccOy8jn0oEVYkhZmboe1lhsoZf
f7qSaSzzXqceZ5OymhbZ1wBGIteawRs7kgIr2hJ0Qi2A3PAdOCtS+TfhgzNqwglP
0+G5woiOh1pLzL/4LGJR3tcPVylxTchzUJJZfKBbYazcAvL6D4+swYOytq1qprBq
UhzXz9yKOBlzkC1+b3FuWKFpZXeAminJcZW1kwr2cnEo7B7jN4MpsavGH2yu/XCF
XvM6CZfdLALTk91JNQvr7ExCUJDHiNM287jLRuBhXh6hevNTPEHgRSy/9Sm8bwW9
siZoPmLHpjbiMidRa1eSkGb/oDDXzLYmRpP04p5JqVQQ1ZmaaC57R6QqyAqjhh7g
L/NchDuT+yJIKxvl5+yqXe6G5Is+4q4GMPRuut0EiHTTl9eZlz8PqawMwCQEwQvU
lumelN/7moZwhzHJ9iZmbZdhhM+mxrNRm54e6AGqWgt2NMQDhqBj8TkLC2VLWEmf
R5pgn1Xa8cIvmb4v9GMO7DjnHWjAdcNmoUXDixChRn0cAM7E8DHepBA4jqqoxSwr
VS8a+rueQ7gtp3h1aV+dm00t41x5Dp6ISKq3l/ERmOdlQ6Qf8pNy9bPOXeZDZ6Y9
NkyLtgEhRZaOvi2F0+1oTL58DM5Apitu4cZOpcqW5F4BbjUxBn2YN97EjM6Fa0AE
Nr88cHNRFgyr9wAU2i/SnPdRCUFzV7IgJJayHW7TeoNqfHtHrN1Z1+PLOXMGkQnH
FqeU5Va1MjEuJcVZhbtrX7bQHiJXDX50hEEMSnV1vibhFYT/FgAmLWcSgsgZyG3S
SW3wlGhvmSufivoCNOebbkOljvAg262oMfvCrWIGG0z2B4YZB/A4shqBJWvehPWE
0sQyU+HWEsXzcLjbfldW5Qz0ovGqSuAEtVa68j3rBLUDr4huJA9vU1Z6/AqYP/Is
5iM3Lz1n5KTfdtZmG4JEzsAOIsv9rl+UFbLWI7Sm1FMpQks3rBBsD5c/kOkgbQYA
cG351CFbUWZPdshSLEUCX+PKeDe7bXqHIKjL5QDOErOy6hIvHkjR1fbmwL50xLPm
ArIYhRAMIJjYr03li1aG7r7DsXfDSG+Vz59Z51NN7tIdRkja38VlcFRm1/5F1f4y
oc+OTD/2krUoFQ2QcW3oaYr39COT/auD3uRffinS6VTk7ryxQQlWqgCkGDlxKERf
nEH6HRZgfb0YWaLzjuR/aWU+b0Ay9wcwjiwb5P/saJ0eyy2npARFn/IT5P1Dolnw
KjBk8yL47SIfKrI1n0R7Pa0z7OkU3WfrIBWkNti0ZsrahGwRBo67i3Ai7G6jUT5M
JpVHbm8APBDU/0tx4RhnmC5LdNcOVbnvioMGprXRYrPbiZ0b31dQddvDaHLxvsxz
A4LbRq1/fuUxd02BvncBujhYiXTosbkq+lVA7rI14y31GTUdge/cdxj6y78nS5cC
sDqhWfbSw9h4Hc171hKZzqYl4HC7UsexT7muJYJ4I9gWTSxAaT+Z+nsUtWHXEoSg
hxnf0qa9JxsvCTMF71Yu8BEdPm1rAYIo+L4n/54GlNIk22PXrxEYCl7AusHFGG4S
x66v3sUCSze5e7yR6wgU2w+Sbh6OY/H6NUlSlYIEEf4lC6x7f+KF42j/iQ0Ygl4E
99/1a583aD+ZxNsCKQnrnSHJvoMKJKp8nG8rM34GkcJj3alJXUyOWrYyya6A5aix
ihR02QPYNFv0RIO/a5pLRSaFM8hUo6i1nHkBBKL8rP3nIlg1Fp1Pyf36Olqg/a/T
BBRbZHAUfmeyCWTBv63ihSc3qPtwLRRKuiiYMOhhUx+rkSm2Dt3kGfJw1l9zhuMZ
Jab+lhAqx9mTdR/Xrzj2RSMA8TmUyjW+8pW70Tqhu0HaDDOhvNVzvcU/4mP5B3wO
F+i2+BG+Yvupifid3vLHGWV2Lle5qBrVmnFFiMaCGFEk2SiFci5xJW1orZ8sd6nB
GLSEP6J90t5gC4butOMqsfnjU8qQFow5OLqiVLJ4D5jLyqd2Lqitdgxw4a7t3Mth
4TTZdrO9uMTHcxA7mNDOTSIo3TUQR5cXU2XaZXhm8Jy2IE9CyvaeIgkCRN3grU8i
zFW7bdCA5VoUfga1GAu/Wo07/f6Mr8v1LXFJh95QVbYJAZCnmC0Lp+3TxSODshJt
0kPLFancDKeNLruIJ5fSi4znJegk1qpdRydyAknlUTYhxPWbIBVLCdr19NPBCr47
wFbOsR/RqhmJF6mdeOvG+aDp0psQXo1t0jjMAzokeikF4L1iFDur/A+4Fcoq3GvN
KuheTpet9Apr5j+huxb3YTMzcX6nNxSK8ptCx9V/7TBeyii5IiVndzDBYqUZ48+e
Y86kz87SSrFTQuegnVB/asV2zk2g+1l1keEpBS8HLA6am1f5gJd0y+QlkResrwJs
VKq31dqMOlWFeGWVJ8vLgHfrQFNGI4vWo/PTsPJldbiHfhoe201qVdMWTnr9bx5+
BCs0awib+4w0Zmq1BBnooCp7WH4HMJMqxggM7uthNaQab6afS620ax8il44Hjps2
7tId+EyClrxJ3c+dq5mVvPq7IeeaSys/PW94JN6d0l0E5mFehIq5aSzjxb4dEr9o
LtQmsZVJ7QZNDpIL3+FoMzVX9cYpPKnzmq3Im3rUZmU5n9xlub6Yu/WCutQSjl16
mH32EqRAQtW0JQn8ahI3c/GDw9n7wmTN1Kqw1p0B9BoZXQmAmlYVqcprVbINLOPF
V2wYSxut0qqby/huI5DoqS5c/fmwZV9x9pFwrzB97maowu8VqAeXc0m2hGPVBIAC
w8XiY/SD3WP1zsTKSXVVydjG7zXuwasm2qSEt6OvY5WCxJk4ujDntGFQvpjWnPtb
eliZWdTWIynBgoiyciGIIz3LTCDPmGaV4Tgdw+99hx5AZeEp07ZdXM1PzbjFKKyw
KBY2LtnAT0r7UPsIDd8MMMWhGqxOTefbnZP+BnUY78WELey6oYbfRDajZpsQAvLS
iObQRUPtrFtscp/A242eWvRMu233IDjhdn+/zLkxMiCqFGmvLmzbP1zEMeTmLo9P
1L6ksoP/gPwysJrbXBbjzFiFHE9/ONLo5Rilx68zmCV5WhRjoMEK8j3M/b1ohhnr
XPeGaVvFS6Ci5tp3Px0Svu/BqW4psGuVM3pEb8XWL+eh8CvdURT2+UW5YBmlpOpp
8Ijc107KpTm4zcDPvzYLZZC17pV0gLJxuDnfQl5dj04zeG5ADo9ov1lIZLd9RMR5
P0gB7iH/oQbyQ6QT4zVrwpuK8zIozO2cFN+x94yPhkqapfVIdtFK5SJwlTIl5zSz
fojBB9nJKyA3aAJReYOLxpOgYiEgPmMk5RotpkPfKWQiSraDh/1287Ln2QphwhE1
kKoq62fYBIt0nqEsLDd7jOOJ1oU4eFe6aRpU868hCtbpeZxjmfggAEteX/sDJb7h
n/7JAjlL4wBPcAAUExpVN/LXreEsD5oJBzHKzwB2VQVW2bIIOurhWpK/jnmgw2Tm
zEEVjo0g9MN1tdT75mvXCH+ERRoHtYktd31eTF9Q4cErGllXrBK4/1vj+FKOwzOs
TTcJ2xgC1K2fFCTIjFOjCEjrEA84Is3GWUWralUJytPClJ/+S4RAMWXdiuBEkW62
4x7QCPDobz0Mk9HPKyrrRRp8eeIg15iHkZ3n4hur4Cji6ANSvFk/RmB1NtM3BqzF
4LxlfIXm5Nhgq6Lq//lqfqc4gEjY5KkkPW7ePCBI2qYlxinUYS6MECHfsihIe/H/
fl0b4/RW38nHKwzqovLLpV36uF7HbMB3dq2YeLoTDXzNngYzTitFWaRCWubJNbPU
B5qqHt1xyAMQBbCOClMIkG4fsdsR/VZoWVJIWofrp1PrLjGTaRJtLX1Q8vqNY+zj
FOcvv56VuSM4o5GVIc8yNXNf2ELnlN5k5AR+rpwa71aU3+jCp8nGF1M8YcaH7HhA
VonE5+AtKfRK5b0TKPzEuMClhQcc1xjeMAQI/YvjJoOFf5qfZhlNop0Nt4jQKJe4
tibAEr8y6w8IWde3KQtGQcMzHndsr8guRBgsCKZQUF13Yu0xpvhIbtqldE9an6Ma
UbEijcFbVIDzVPC4ckriRhARiwvcQqqddGz4yqT3pkYt/URc2I5ucDU5GEXPG5WS
z6UTt8FG93NimCRJi3qRw/+RwsmaucLvcTiBZB2ZCGExNCz1CXw5iWyN0ResHtRn
MHjrVGFrO7Kl3XBahNZkIrXeQsT2/bdWNQWQfD7JBFoL3dg0I0P2HzwUJMCTR05J
OFBC9WgGWJo8wkmsrhEkW/2F/LI8qz8zBwiMju/tSRVRxVia3fDEFs4/f9vhu2Wo
7JTDAEvdFERMjlyzV3i5KRdIPCAUd80hHHWoSS58nFQYIV8ik52XiSWxMGocmvDd
afSpwSw/Zb4gVUkOmGw2teerjGWYeYvjbh3LSmf2K+QEtYSfFfuMW0OiqkUEQtml
+nis9eRf4VGxX1QuZQkRZ0JoSUMonOUGuwDn5JQGrSGJjCr3nsVF6TdBewZ2cIEr
wIHRJj/rk1O/2Gk1sDoJYN4+n+rqOf2+bTSCOkFVnJsh/SL+o6WpyW2i3POYq1sw
H61wNz1oTAuahDoVN1la5qb0z3aaXFqg0g08m79KrKLKiHOSKbUfh4a6HkKRKBu5
mVmKWhWlymjaGx05QCXPF9Kx+hyLYjqBb4KFPfcLZ3IIpIE7l5h77X3SnA3FQmKT
3HqXp3TYlCyKwp+DGFsJpXplyL2nr/FXLWYp8EHmglYn7udsMDvIOFz7Dj66p4L2
/EUxjSbf8wmjgIb8Jwz7wzfVwSMDWyOhy8Wlb0iprY0yPkH4FWod+K5bkUFTYoQk
D5olTC8HR7WdqvNqXzkm6VhU56LaqIk8PkAr+Mn3Blf5W8/W/K1wYMV3T29mmGXZ
9SGhBQwP4v56Uk7t8gUf8Rl4IVnsRJgXV1XLcg4h9quSUNcKiKwHQJPbmyjJduWX
YOUlM6vs4kVGR1m9DZJjGqY8UjlO+S1iFay8rQGLvCzKNavSsVjMqv5+wrAsVtAf
++h/eFI5iniBjx/0B6UG7mVes/T+Aun6PHwmB5TWO8kqI6uRfydMjQEgviD70Xnf
LWFhk99QRXtlFx2wSl1tz7CpCCmTTXT27U/Rhvbk/muGuyklLsYmZnmJsvT/+CcJ
Z+b0tXLctEyHThbtV+eH0ywYXz7kAF7PlcA9fhMaP9IXqY37nAoAQzXv12VukPot
CGJD2isL5ge1qIL3u2J86F+8BGEucNt8p+lWlsqODR5lT0ESNNu/IjOoRKbviqWR
2L3ohs8I24Zore2uBFqjAvYKvMGtwcYxXrCqKsvCrxyOz0uGhuSexdyxEGN4P15Y
tJbK/1Nfe/k38PfEvt9PVeVlSUTeoMd8FKaNJZeATQBBBtUsaA1lLyWLUojUarDU
VeVUz0yzg/vcyDB6UVhGG8XJMawiPlqUX4Mq+BDVdLtp1ZOebPlNaFlm4aantJ/a
iBgEI9U6lfcukX8f4KITm3lFyjAnftNG5Lq3RBnhAmKpI+w5vbki/npxRqK8g5ya
DyGUV/AM7m4xksk40ykej47bqoJhH1ch4nCnrRBA+H+kiGgVyvCRA1um5CFJeyRr
odkaDfkDQSx2pB+mdUTYUppTFBW/J5AESMLIFYivKQ7Q15P4Uvgxu4BzQJRUvEG1
TuYkPMaaq19LTvVqqL+NueDEmZ0iXLmK1QLqFJGAAAyRMA31sB3V3Butpe8fnWvj
zh6V/4DcQ79bABu0CMgQnCgcSRowTVymhe+IoN7nTUgHj/m8o0x76YnoyfFHX9Qk
VFfGonXU5in3Ez40bP71TnPvz5etpGhEXya/sH/azeqefDbOL+Zh+36v94D96P3E
hbVJ4zGg52aO1iw5sYJ9mVhjw6bXVSTQfGmKwVpNl4GnWS3XnFY1dyq6i2mqeULZ
mlRJ4uA3E48Q74KvbiveGOUFwGtmt53PXAeoqbA46Ht2CmuBKJ8+bXTbCpQlZGRz
qXWyLnLozdJQ+Gc9INvK6pcC53JCjGL08CtKa3S3nFCpUYM22O9e0YB7CxdIDtxj
kalXr64e9tDhsLl5DQVXnCTeyhzxaVHg0wC1a6VMErUiFf+vOArIRG5QbfTnmQfq
PR+vyCNXwpOJeQtKbSLDtNNCAVtlwselDQ9Xdcf3gN/+nHKqk9LMKXhLXqsKG/Vc
KiSNDuumhI12xtBFTg278ly5YBO7Q/gvoyPGgDKk2JpazFM49oXjfYiermETX398
P6s61X8zPNmcyYCUwYdGGl8tC/zGg00PhKD8JWNdGAm4V6S5db7aE4d4JKT25hnA
Z0AjuEdHnq9JDLGNL1H9IK1SoXLSk1yXo0nFfZrBWMTScAdvhe0TJQRlruSmiE9e
OY89KeTfCjHlyUJGjYGhnPKSk5/iiLCVw1KBmTI8orFO0F/aEkiVAD54uA73pSBy
Jq35h5K4Zql9ufvk+KoBoOjtkcZq9P/aKKh0myApsT/rPvEEeVcii88auY0FaaOx
/s2j+S5C4IG/MVNkHu6KDZP6R2ZNAfUb4RQnRDcbQOeMui0pLO9s8JmH/RHbej0Z
BfdD5Ve6Q23J278wD9QU8BRbg835KduXh+0PN8HJNoLNaRqWDD2zRoJiYxIUUEEF
+MViR00l8IbnFqAHLT8isgPT/1vK2DyTqOuKc7ZU/8Vcx0p2i+IqlyR72S18KLWP
FWAf5zgNZ17jWPcigm5GmjyKt6ClHk3i8lhZ3RAgIMrsdYV1Rs7pGRETpS5ys8hn
ByDTr3IiWiLlKe/UB2FcrG64TOBDIrZaxdhRhBauyWn82TJMnFHSkcQfCMBh6ZUP
I+pbTmONm8Yikqc4g3twGSUirbeYR+IjEXU4OK4fNExjAJeSF+uj4GZ4E1k19Cdw
HQGTgfI6fXRnOKS4vWTHAT2mqSjtdRwaya5eXprzEO4F3ctGJyPtCWOYm5lS7iZe
cIcqfYC/8JU5FOStdbvLhuHzkhq6uhkwqG8l2GfAn9caW/p9IA0l2z971TjBMajP
AVPXMdpANg6p1480WXFIWhyqoYvsssMR3EOBCOFk7PVtyUZ9QVtUxq9JUdfmIw5p
QFBcWldYC0XExWhtZiwi+NiVAhXmEwiaB1zlnpi05xNiNwNnkGallMDh6xYqzpV5
FL5XkN9yzR8cx5jx6wVCh4h5I8JCaRmYj8GK/atxGw8rdTjZ3GyDf98JgpGRP4ch
2lBi0qQUtuaQci9PO0QDfTKg+XG9FMuZ1IOIuf8XbRX5bY5q70/9KkpLafwpczvl
TZ8q2EHDJCsoQY1SBwIFxDTxUogyeQOvOiCOGsDLsIcwakamIchGev6erDkGrM7s
ZqFIE4Em7U1phCi+EPY62L/5jz9KTFq6yNVgDQYRez1+dwmYpg6HfrpKDRuvVV5U
55h+YxNTSom7MLd725VWAwK4QVIjw0FUD5BPYvQVluvc9cm4Du9QVlklOZaF73lK
1vH0kHyrbkIjlwyLpjaq2SwF4wcuJzRLOSyAujRYRFM28cTHTW0yqTwN9dkgO9eF
nzDsA+fj3f3YYQb/RaHZ7JyHR6F+Ust/BrK8VhKHAGhWSuUJ970x07Hv+RqO6+hw
16XoYELe2Pbl87RWbKFq6KY1UWsPhNUDDlHQTCARGJR2c1npgraeTB9TUBAf3C4f
Z4q6Dzyh/ioibX4yr1xAfjNJQ8B4nYwi/tcYASqUEgZNZB02gq5VA/zb8GNgNHl0
xsnIn8FTR9fPL/owbWoUqUEdq/kkfdLfxrcDq8xOBVAq8G/+o1Regn2RPa+7oIm2
sDWevN323/COuW6egcjo1IaZsE1UM6R5U0A46PoPUXFdrSFOgBvJzIocxDH7LoyK
nUQcdCGNyeLrp3Svp68iN6QUFJ+AEUSvM++cr+mNWzpvaphivfaLlSjHGidJn6gA
2MIk8bz98d/3M1QM1xStHda34wWtYDnOiA6EtWqc0WS31MTh3j8dsPI950epQ9uY
yVuBTvtWknDLReFuR67jAycJIR5PhSvoTM9M5xG2LKidJCK4nATG/MowB+XwkVE6
vvxgyp/3OGen/3IM7Hr/0AnL21nGG+D0CZKmSEz9deV31CsFUGYSSaC9JnnulHHX
rjZq0x2UgltJ1k04SyvqIO8asuiDnbtEC3EduJaXMkoVnO4AthnFa0KQCNL47L6R
wCqBaEYgUuTzUOfI2HKDSqelzg1VlJALeaHwuIIxLeVvBB0FJtF9Gf3hg9YLxoLJ
zQt7Plx/EVb3u/u1Bz8jPwxaXMQfrclKt6tak9tZaO8xHKFh8fh+CD/Z1hZQLOWC
kTcp75yGXoVk3MgbTgLT055D55uedBu4NRRgVpeYJUywVdSgK4mOH15f3MWmOIeS
D5HfUE6jEgj7NeRA2GvG8lnNLIm+eU85xwf4o9NETFJ/7AzJh8STBDErzQHFuuFF
jowO4rMqU09mw1EhE1LFS8uZmb9nlVYx6YLiNZm8T082MiD1yxTCH1fPy6LX2thL
OGkJ3WDN+iBlem3GBUF0gepxq5pCw28tpC8hsSDuAGrKnj2aSGGiUtjBSuZW7dr/
YiDda6A2WJZ6xMr1nerOouRlScVBlj0+3VffXjTQ0jlWekiI8puy+mcQjKms6YxR
LDUuQa2VVvyjxMslFjnxiDzzqpIbfM44CrTl+JdO3lt8Ncum4P2IfnSpUkvGJpBX
GGip8XmWxjptqGLLnIda6V0Cezkqk51S2La5jwFwjj9ztdqLYrpYG3M80rd7Oa6i
GZJvdJcLLZNs8RUCt8fPLJCiYjQZr/yhMd3XZVEO6CEI34B8s1l6PK6c+0AHn6+C
gVCe37gfXZuo28OR4OJ1NVYXySexX4SBlAsDNGLm6soMV6skypM2Wwpe4YFEy8hl
lGp9beCVVwGMRyY8QTUyT+RSGMPIfiRsKM6ywDrZ3J3aEbn/ha5aNrso9YuUO3F2
Pax1BcvoQjUPMBcGJJ/nNHvwPOOIAftMR16m8HiO705tV2D1snkveIwbHwZc2DMd
hxo0HwqI6JSHkesU38YvrUx9u3S5hmrW3PET8pd+KxYLnLgXTOyjz53cbMnDcwPg
EuXaOmN2WesvpHPa8VBWIs0kQscCQobEHVO2L1UcETqcdVDwPgOqR30a+70XLMfM
4Qh7Bb98mSjmbBNVS/kABzhFUh7R3HFl9uPQiuWApboFWd51eWQyf3hOZz88JQBW
kiEvnCMMmpBpM53PTuEUyfXRJLl/EuwE5lNYp4asSzvWuhFl8pP6kUaEDnKngjdZ
KgO9ACj8YoSoTLX0BUR9KweM69AkgPQ0BAnR8kfKpARvd98bKsObaujFHlGJz8f3
cDaRHAJYYwGKXPy52BH652gOlRxL7+sCtvawe0Plrz1KBFa1tDSPuM44bPke81F8
i1DooM1L+K/kojgRNql34DAG10BR1CZgNJdPOHMulNs1FnF0Z06K53w76QJCvcg7
3syprqWBspsL2Q0QgtFaB4ISRNHwjUrSpIjWPQ5ZPs4zXJHMGUtbdRuzt7DdIcFt
D4bFME03tqsgdhpuTMRDS6kEIG93VRYsfCovYCPnD4/07oncKQTl4Mv6Fd0bUf0t
f1ADMpLd+0tKB3FS7Gi7/YwJPiYDDOfdYVAJyEVUmPDV+tIZisoQTd4e7OsZ9BXX
F8r+IWf6t0Mpb+9EutLY3ZaWdmw8qGKWfkjfwM/8mcooCWUMxf8Ehz+JRd929SZ0
upfdORR4M2Z1gZhrgl1ucLo/VkSpQNW3DFBTpWt+STTIUbaq2DRqfkttZCYTE02W
0N2sxeO5++7G/m65wyUbbRztXYNIHPmTtsrsrNI5fJTJIwdMaCEoHazKJfy0knzW
1kfdFPjjfoX/RyFiNxVipdUzzaIha7mVdpShO5WpjTBHz9QhUdqlsnHgKwxwV2bv
dh/U0egrYSiV2bNXk8mjVxGGuI8/sXLAdLEU1ddluCn6rJvP8zh24Z5t2dg60dhk
suaYJAUVLkyEdpHGnFjGlGl9YpKbTPcJLl+ff2NDqA+ygI+WUlTj1d8EdFOSZHpv
V4zhEPrTV8hc+JfHil4NA8EM1XxijE03OZc8lS4iI0Znu7goGlizRG2fZzHQsAeR
DF1MfdD3CoWCYR6MDEXuCfgn2X0VkYw30UxQnZnBz4SqNugxYIynCpSCQbXGnRfv
AMIZhcrzSovXcDxdj+mFtrGLbbdZXewxV4/LCsVrIcJ+hFhyAp32S+SHbVprrFT4
g8CrRR7qI4I4EE17W4Atqijm7rcdEoZbKL0uMs6cJlu5uRUb1leHa9j7YmN7MMfd
jzYHyxDN+fXnTuhoq4o9IeXpxjXJEOmZ71Thq3MBKik6UEIV2lKsPdqkB5w/cOy+
/kvcKTRKqrgr0K5iSsyWfuMQ1YwjvEc3WU7ApHUQZlde8LJGkwexUlOmw3DBuK1Q
sMkpsHpJusRtTsZrP3eASGWiv8u/dIS9TOKgMKXV4zo4OTpR5qb8cXqPJ46kEiHN
DAUXd/qJEGmE0sIJcFD1unAljYJJj86UvJNLnMMXWNQj+mk3O+UHyndcjUizzKNn
41Kx6nf8hfJ28CggX4Yo+dljyqHGlyjgqyZ+D/aurRq02Z7CXfsER3cKUFaVg7uj
09taD94Ufu/KuTIz9/b97hb/Btbb43QLtbN9qvHqsQ9XDKQgcYZFcD/7tTzA6m8R
lZKVmzdG3DzVzkE2nQZ4Smr3L/0tprF+LNqcdiGRUVkgG0pL7OOAMdoeO5bNp0eM
gLmz61LpTLElw51PyAJ35AfbNnPER0PVueH572AKiezerCFZZ4jS4+L5RpXQFlPC
YaHp/z7c9rJsFZIK4ZMbq38X0ESc3C7qioN/2phw2a/lvY/gchQt5lIcLC30tNm2
NkLTYsJyQCQ5CQ1LTA/3f917jbFrB9Tzx//HjZJr9WBnl8OkBisQX6AtekTZbTIq
ahg/n6iiU+vBACLzUMsg/Fj68rN53VkXsU1xW1Pw8Yih5ILLiNwnaiQcMhK/GkB8
xAnxAcZ2twSWdaJdtUwt7lENtPGlhbAGJotzVIxVPUxb0dncOgvRYi7CqxHRGL0C
vU3S3DIQ8OefKom/Eac66gQEU8knGTsu3suxz/PwjWlwHqaU8HVr207oVMrs4KYg
O+2chTo39ru5/0/yOUmC7g8wegxL8oM8c1eWZFb+QE6ElwGdPiqpjGYpO3Pmnw3/
JTKRynr6rLiREqheotaRHXfS2J6K0j6gTrXcZlNLKyJkg1aznH4HGk8gLTLLnhLN
0wAb2zJnqBnDWjIYpXeD/E4gKext6+/iSxoEyDiWGM72/AdB4YVs+BFxUO/f98cW
93fo0gRBoz6WMmBvUiZ1gaJoj1JwWYOknQcXQOK4biuz/xG7tsxK0iNpph3RmJ+D
b3Dv5Uy41Pl70pxaE7A1Y5cQQyodiyVrTMZnhsUzmO+zdS83hNdTWcnE1WE+rLka
LDhY0c3gI61szFVa7kOB5mRUgxRkBGADh9pSKfsK0JVA4l31XJ7idiU+8HbhlgbQ
Z7jxVZcWIF6wzXM8+CMfuV6AUD5wCjLew2wROaPfL+erDXvI3WSXbQEdFD8Ajxvn
MTOdNTWZnwMXng7fqTIX26smaN4C1LH3quI44gHtJqbkVm9zr1iagEOg0RRXTb//
CNMchGBIIPKH+KKh05QpKSydAUBfsanfr6XIXN2mV3mZIyJKYoYrhzrAQqaj32+2
AiWN41AhH/nrXx62w6FciaN3xYA8/sDPXVWWAF+MPhBrb9wG2cAcsK81Fe32lqqV
k+fZK2DzrOBx2tvgXyMmtHWnMvEhIn1H+w+5/M84axanE8FNCvkB8L7kEJ4TvS3P
+IpWF9yynNlbot5Z9GY//XGPk/Uv/YxIHu26R3Ae8VLY3CgF81Unpc6FJyw1yqso
dsamuJqfQMokkw2jfrnQqYYwm+77i2jsUtNf28//m8bvC1aooLZbYrbEj2pov2TI
V/OUTBX0dy9IarDYkWmr8hQpE45SFD/iMKwOrkW6vKUUbEHGrXX8kV9JEyU6MqvC
GS/HgbQ0AgjdQKJLQ0EpzBQOlXJzvRQ/8XOS3iprsyw7D6oEu3Fa/GxE45JZVVo3
2xmM6bUcUwwORLYZCChj/cp/+YmfsoMT4QKt5sk3CAqn1m1QGcHm0aToKY/cNxI3
OMV0u0QLzsTqlnXaz4w7VQ+Ob5KXw6k1yRw2KGjRkYMxm5Os8kLdz5K+FSLjFQSp
ACK/TsWKfLXtPRJEsIYKR9rmVyaGZO/1loJ2EMdNoKTP6uTxCBctaYJCfUubJGnk
AJMlTv1hgu0+H/4CEwLrbfoLiRw+2IvtpVNWAPU1oQIUk5PkB3P1PocSrop0h7Au
Ef8HaIwGCEM6BEKjFFs7Ilm/AqNCzHNOMIHH/nkDoSHOJxa5y8FACRENwMvBvppL
y6IryEVMIsNMfkuRBlMyinJv9QbkkfblUTi4ma/51hSsY24wF6I8aGwH7Hta4vWd
9KNSQMc4kD2n1SnDGMoPLCXckpLn3oQWBCKcXLCRAi1+ejRsPAt+llgOcZh4Hd0N
HIyoUEUfLSBYlQjVBHtpLOnZt//1s3tBd/kpMzq6QgaIpRq9ZS9W+XVbCHrmMGOK
+VEQ4iFjRuEySsP2Q08xuN8clL2EaYGlHD36+SIQZ6g7C16jQeulVxpCm+auUsxa
SbK+2YiOTMwEkiW1eNSjpdJWE4jVIebntNjI22D5ru0XUTYz3E2UupABLVzyqXOy
JQFWxWPIxmxbevYRNl4Cx6DhfMEPr34k9KPxz8UKRrAsLd0rzpeXfEcFcrBWxl57
KOuerJUuAErYsy1aCPK5m7XKHPqSixRNbeg5Oo2PT7b/+UygUzAkb+YArIdsParA
2PjZD5mh63suEA5jdlzv3kMBE3j2+nvTO9/dx9l+ij2ZLsZNgtNEzR1UUm2XZPNP
VYYU6bDRF7ZNLsM3Qfwz8L08aTR2Q3/4S0MHyvA3bqp/WQiDErwDGqDTXoA3Pw6u
/qqxupxiUAsrP+NhFR5/WtERiNvT6ZPpOXpz2k18ldgtRCg2+6Cdkyye9ukLvy/3
BVHCU7hnIaVovQGzVAR+21v/hfQU54QR2PjAATu9jAN0sNrgMi2WHHEwwtbQeftA
wKV8FzMTcbw0cLGahdWs1FRzmdEb26g4ueCh+/lbf9yn5ywz9WYyx6PdKjtGp7cC
sLaORUchPs9IhZ672QEsg1eDHMzW1Sc00MaXH0FTGW4j2AKUNg6PYbTxk7poEwT0
bdKkjedpA5iaQgp8d08NecML7tg7DFEU9+rLod064ez5Hkf7W2JNDiiJtrsAT2dc
Qj6qvfURW6Ddl9n4NYRW7w1mrxxxyBSyv6wiCIxwFUlELgzfUKHqhzUM7NMuf3c6
qlRgrucSStdlU4tt9rBZhbQ2bObRSJN5IskiucXqC/pRKR0uBAez/utoP/yyd3i8
gaeD72bD9fJ4gdL78nBPA8hsrZDd9TgQYrPSC8VyDbIaAcfE2tJ/xYxnx4/BC4hY
gKnUdaNyE0A6GkFRv3TbBGzVgEIsvPRF5fi5UcS8chwtF4rSoF4V7+03pdzK8IpJ
G4vJ5cWORaa0ua2//ba7mgv5/5NTK5CpTZeEk6084S/0Tk0yJrTeH7NPenaRoBiq
YF/72SdvT2ZCr4YD4PTHICiPItXDm7t9H8HvHPOo8tWCsG++vz8LRf5V7Q2ZoMb7
eltxgYjRXOabghJP0Qyp+XMCWL5OPlmLYX0IqmhUJXliz4QRyDOxSola+mUicgXh
HSH5iG/nVMSx8A9GJBuvPvCy6DXyQOJ4aNXPPErZqPalqooBe8nPuyzeZe+L26z7
G2b08gqWf7GM4Mfj69rqTB2Co7Fi5V/GH1qSga8HC/K1aY4GqqCymbb476Xp39af
GT1DcnyKkyYidbP2W/b0VxMhgjdnBE9jh2m4EoBXVN/8M3yxSYFblmCkZJ+3kqIK
sw9eiC29/9OUaulbAa5B37WqDuovjkIgcofTcw2qNrL9VvsEzYvxBFdN6AQhhGca
mQipys/UhoDbAKgz4VKohVu7DJsZfnhBNQYGflLDichM1GHpqL2HwzdBOxjGMW8Q
Kwg8wpT96UQDix3+9vu2GcOQ5/K1LNTmzNqprK8oeHSVuGcGxXsxM7GhrMwyfiem
62XGWLvf67RW+sBmMeIdFUzqRxr4TBwUpOWlz6VOZCN61JqvRyo4HBICyATvAIrH
/C71n9PHJmmXCQjWA0FX9Rxe0zNFk/Xwm5m+dkg84LSciMnzeAyzj1BOyzBaAVj7
NEmRiTIllOsbhxigwO9x/rTlIt3X2XQVFya9kmNGzWcosTXZnW/PUXrlf1M0OEug
TLSE+iVfmXjC+TWNZ/2ZnCj9I3gXaKM4DHZtwvRDn6aw/3kTN7NzQ/iSI4guI4YR
nhG8iytsw1sHMoipW5HkOB2HLOGjYcdxOkUlNo9WxeWiQXy7Kr2O/gMqwaydX+aq
smuPoWhyz7IQ/dR1pg9nkSIN+bf2asN6u1JwvvcZHPBrk3FbHdnPUot1N9NLLiJD
VMXsZXbIuRd2Ao4pZc+sWREgH9S95o3HExCbqisop7R//Emv9stv8sMka56KFqVY
Rr3CZqDf+pEuKEC2riCco3B25fkn7our/xmAQx3NoOtFREjsoB/xiynbQuixgAPh
7U3CmsWml7FksN4WT7vXzAP8/YTphMsrDoj064NuPDgC8ISoNxY70E9WqxoItHHK
7wTkfCa3/W8XMwUIjpzm3X/tE9x0+GO1+TY9V2m8/BHoTJfscyXadlgYnJdL3mjL
6HpcKZ8FwfwxxPyBJx874vawxSSvI4GTb6Hw9lQizb6j/FDh2aPb+7Xnu0fbTWUF
FvDdf3eDeDcY70Q6gRgbZb6ZVw+8sL4HrKWd16JdIN0JDtpzUO5zHXqlP5lL3z8Q
mAdLWD94HekEwC5dBuvNtBAUGaexjBgBqYlujqp26ERQWfmZIdb2tj9WJWQ4/m+b
B0Qk56FIjhaoqg9TSjxlEESCU2xfN8vPeo+TK4mKc5KSYsP+2TKInbqzpAJyX8jh
jjKGfO9PlYCj0gsK01SLBbJp5WBZ5XcodQecfO9zACF9qrCwnz3kd9yo5Gn32kq5
mT/KXWjIbDuPdrfFx6RSYgKhGLKJWIKC7oBKBwZIHXvhy4PbWWK/CaYDOneLHPmf
njRzOkTJ4p0epzi8iY+5V5ReM7CzTAyY8N/Bo/u+QX2KY9Hr8ml8HCo0QHmRUVyu
Q1lMd991LinMyPEx4DrXbD63k/FDl9leeLmRjcRjBO0md41wTcSRgrZ34hDGqS8D
8uETNFx8XwnjB71uJlHqPxI7LvJd3MFXeq3izmqZAgVqt8awyyi3vhBOvfraab8F
4g7HLQSv1Rt2cN10D7FEuP8PYW2weqLsMPgXp2zgw0MAae0SexFxPUUkdRNU7HLh
TZxjCD/0FVDSx3MUc4ypTL+G8MSXEIwxjXrNL9pIPogQLss39oK1ixGJitjGsQ6u
vmfTgOSYw8PWPfm13QNWerzi0T54+V/qtl11/Pr58bmfWRth4ykPUDAjMyWoIxN1
95WFBD+uaMw8UATKLpmarpihPtrJc5PsdJfru5XydxICS7JTZArsDZm7m7so9HRc
mCAVpJMTyk7uzQBdXxgI6iEz+7oFovAJTWhoAVEQ/pAOmWRt3VNfKRRoDQz8kgXG
BDQMUDhrMd6MHksKmfGKDYd6BFWGJ32fvP4hFcPGmeVoaZg7AuLS3BeoKkQBmLdH
IWo8i9gtsXHxnHzxBzj1ppFCC4m7pGZ/TN8gGu2zI5hhSdlsErQuKsJm+NXBF2GK
aecxxCpbOWXtPC9+WaXp/LsUTFwSjH1OmfvWTc8LUGPYwYrPrevGqEbf2cimbah1
eERur7lW+vKgwBlW1r8on0L9A5COs+R+JhfzH3VjFDVsVABelzDD/BZsG1g4f10x
d9MUu3iS231u63nzxeM80GBTht+vsxcvsOKtJThvzRrStjodcUTV68uVvHVwYrr5
498AowPDPJH9Hub1AB6AaVIt7XgQA3pZRrcCOu18RRkvaAE20VcRCQ1AaXboJegi
8xqE53REpDaxI5BIawCPuAGFal5jw+7HzYPBethE2WBTTNO/CqPHSdnUDgBsn1t5
NongPEIH8w45vSoQhVKIp8zHLltdTOMyTJv+yimhH0rSzjB+x2wBjCe+8ycP39ZP
HdjKbThN1uHnoiMTG1DB7WvmkreDrtEonvWFSYFb8mhbPtXIVKCU7r7GYLb3TAfr
RpwyOn1fqD3CNnw6v27NuNjNo7q4H0iTO+Xb117mAQ/tG/LauJ5wZBAxEmB8+MGv
o4rZ/O8aUxndzsZDgwnWs7AwYt5JVzZIe7ocFLcXIhjBzctd5t7YBKAlo00Y4iN8
+VBVjyCM1TKkbauM7ubBPb570hNWeQlh6Mc2LXMsC26AlJJQR5++Ly33srWJDMFa
DC+7l60HC9cI3d5GfdCWWwiAx/RQ8UhVSGBo4hV67P8TczBCLjWhILs1fsk1K7DU
dE/2jdtfHgFCM8mCNbdoZFnWQDzS03WeuHwOu6BSCrXJY/u0m4aEv3iCkY8EWcYH
rMLNoRQXwQL881XlmJPbK26+C0XKz8hPycQBJzQTnorBXgiJtl7y+3oEpB9u97yB
dt6PuWjqSHytvZToKM7Oli6s9CZoGbdU+uGx2C97b0Jhhk/vpIEdlS1e4Qoh0IsT
JGTJA6uatfVCFg6+1PcRP0wFx1PUR6PVokcwjG/tDS0wgcG/q3iNcP16FG6LXEAn
eI+CKvho+1mqwDKJud3RiiL5fX1qU/zZQpv8M8+y7FfZDr9hDn0nd49clcwmxnuU
wsfs35sQQSuBxXINhv5OOOGl/h8D5yhK+kcg0dGVxpQ6gOUyZL3E6pHI78AOFpAu
ZS879ss722bC6/pJBxQpJjxG5iWAKU2b0LkEqtYlAFoJX8A+0Kw+9DEa+6IeJDff
K4hlI3yHcI9vosnOqHChK7EQnPHFixWSquUuvKSkbXErs8jDEv7MDLEtiIkGheOq
CydpX3HltXIhiSQBOOW6l+SzIEWLFykTftGEMThZIPymme1i4DGtOv4h2VLyOx7n
hRAtDHK7A2ydDsKpU4sm+5pMBZEtUAazvCnWpcIXlFadosXvw2n4naxsS+pKlToI
vy3AUlHYY4vtqmwkgnGhz9DyLRTyPS+tN2y3DMlBZ038iJNhL8i/w3QRgGbnE4Gy
oOHdPnMFzK1DJvDnivetDKKoH4ljUVt6AzsVUlXaBeSV2e7m60Nh4we3wWNDhbpg
D3qOqRiZWW8EcMWf5paUHVDj4UNy7i60/JJkF4E1Y0URjYbNABNdHz2G+vrKuark
8nY7wxhcWLb8jgEqpCphCgv6/DjIAFK7Y8xWc/FHEd6Lk3WmVjHvgZbyO0GThQ9n
FkNGz5T+oNt6dN6LNAuO8Z8LaX0PZhVZ+VmPL0OmVuZn9a/s9Usd7VNpIi1xq1jE
ZfQQD8yDeaEZJ15/W/J5BJanA50yapSOGQ82JQ1Rkz9ADiPj4C3s/rBmruIFvosG
LLpK24S93hHUlCJezw3XP6Aw5DtCIB5DDf7txWK0nYvW92+qLvzPH2KWLXKezpdE
hg9/Cw0VQOGzkno1FkNY3CQfIcHtfFh9/N/bfJFuOjNfbWgjkRM2yrdCgcMGSm+S
uXTRwerRmhRArxKY31vp3OuUOXDjB2J9zZcaF1NP1t/PzOFCPPXitTr3tWE/yOjr
GnaSqEdRSMicSXdR8gh66BygV62KvRyYRpHTBRgCzfXKOckmoN5qvhP5qGMCXa0C
TZHnmI7I2qB0zItkDPuWCZWMc3vSZQ3idq2/cRtMo1FMQsPK2akhnAt8+3p81T/F
jZexAtjpoQgtEvGruxffRU9/xafuzVvKnrCHwfghB3R/zGsbRTGSUSMmMwGH/T07
hsfVXN6h0VDLTMFDBFnuWJsNFWL9ahnfyQBduLFxe8cJqUQ8sI2VnwhD8VxzVpgI
IszDXk1MY2ATKd3q0tuNkZubi3QHMfeGYRN90Xtr84wE2Ybw+SDSwa8SwmRv4RUC
rSwStRTyAU6Us431xidXBcbfXgdXLn0IjjqFlnLsNZa3/6gZHMXJ+wgOJLI0rEAY
9Sp07JI8xcSVuriUT+h+PYni9wOVGv9D9CW1QzHNyG49CVsclB/p+58R9QAIKx9G
twdfxgSimJ/C78t5SiBrqLoZEMaZP6NcPaGUDYSAnrg8eItvRACnbwxsttnHoTSE
T8C/a1y1wUDtWrGX4vCNmzjbHjUtVfcaY+9baCdE50PoInZ6DVcWD1U42gV8szse
KDeKGmGOJip4sm+V3cSavUTpm740H5fvXGql6rrOdWX/m4zC8qoQSeVLoLw3Y8mQ
syqgMBJF/yrZd52gpSGLL0xXu3My7rJBfyN7wHBghhwp0oJxln3MoACbe+7zSZSB
3xJ4fuUSuzkgOH1hhArQjWPAS1xHEsTrEwKQYe0XBuKM8dcipi8e6oDCYW99SgNz
BLLp+KL7NfhglE8MgdGVI06IbRDC2J+XyUrS8Mm4gXY5SokQdaN6dJfryZLQeH7R
p5I4imxE+vWgqa2fMAvH8+YS1wz6LpaiE4WZIS88d34gKb4vAyCumL7Vd26Fyuw2
6+pnJBOuJjBCarP9+Z88WGF3oE87jyWiIpeLiNwHT8+U+6r8CfcFT060TzI2lUqA
Bv27zWeDrZBLOD8T+s2MrpzNIPyCaptU+dBr+mxpPCf5BDLOYy+uVqpQdFFGDvIr
wSpYrxsNSxf/lsnDkFxQLQdWST9R8wtPlOQdXjcN9X4q+Ptk+p45ZtSfoQQ8XoGD
dDfHji+SV4WFxHXuui7wwnnVHYPQWbZP5mboFL1kXRgvkdQxwK79CuCGTnrKzCJF
WFgd6gdZL8TVjHZsJdkXLftsRk/HmhjZuOv7DGBLmgRjrfhrPh+bcKiWvjOlJYfR
h2/sZLgIdbynBY2s0/61GdWA7naj8MsOeYx1T6fWxa/OGyJHR0bI8ssFVuqojP3m
sPqt0iaW2WVXWi47O+DlfKeoT1k2o7bCSRJq3unEDjYi8vftWMI8NDX7liXA4GuZ
xZoUyMbMHh6AUlOrFBITBfiOox7rbua1En/QHaS3ZXEqBL5HSMt9UM1BZ37QYfDO
534ed9ex1Jymm2Jl3+v6DkOJp3QyD3Kn795Ib8l/11L6kFLCIUjUAg9TjJnk5Vqq
2iF5Bov5VznLMZzaBXKoTSN2nMjWcx/u5jEgTUys2O4Vi8yJYL+9nDquMnPYUVza
MeEvM35QOYyqT/ghoGvI3/HUpG8KA15wUX25hTJAaJIoURH3x/FTspm9Sjm5kPJu
dcS7w8jHPldBZGwwVoS8L8eeepXIixaM7CCvJoMSv+gpC7dbkqYTIH6TUWM+3A9z
XQz8miFfQuViylNJStGM/ur9Lq1IyMmX9bo5wrBdA7ZlbtCU73Wv5uWfMMQptrFm
3z/qiA/F90iOx+im91SlPkKOu+rsdRewblCX54FfAXIiMYaI9OVGarRaxVmAyJIr
siunRaER8wOyA+cIp6cSoZ+6MKW7uDKnM1/brpWlECD8QTup+F2ei3MwlaJX7jhU
IMrSvVWJk6LUq14838PVoOUMcZQCvuAU5yiZZksO65VGnTH2h4HuhJPnbXG0WSeH
eOeZwzzJj9/r2Kulj/hJVno43OPcFTWzOu2MHGqI9fUAWMmMLUbg6+YLAcLF1Een
iENmMbpbOSHhxhnotZ9ZXWNH1+p+Q0lYunw9RjRb4xJWCTKorwKOyQXPwxrWiysf
Owf62j/d6iYbe2wNNpSB3OKrBH4HzdlWZg7N6HgnkwEXMpYXocih2dvErYYK/E6Z
5IY4lXH9lPRu6dj0DMzVd+XMD+34twrua384bbQ7EGM+AdFUL4xHdOgwTaqcwW16
tiRJAivYsl3C7W3c1rhIsrzlhlpNmXCs9xD7u25VQwS0jmMTdM4usz4TtAQ4zFix
qBCujjLbxZ5n+C/+AxIvDs0nyJY/FPENq9dxzLqAiiJRlSX3xhQPn7rH1EVQPnim
g1YWZ/j5Xg3em8G7D2rdFY9XoM+R5PAVBAXIUN+2sX8aJMEvqhXtNuvLtL/oyoQJ
RlolVL2Cc9Juq0MsBe3DpslVnewwRY+I6bZTnbxPW0QPEwGssiWs/3rRZzY6gqQC
iiwcSqC0teiUeUfIMCPhsR6SxIry4iyUxddQ+G2YO+nXbcWVbFUlUzGOmFCb4g7l
FU2Z1dRHEZbIgqHufWu+jsueLiDAhtd5MR1eQlh0efxcjUo1lhpMA8sYg7iw9e/O
zA/NGWMp3Y9Bl1P+zdkSLKD8Wp+YX17fMrVbfR3WzZU5+LhctpeQ/dE9NPyt4GFU
i7i0XNRZf47kTSlg9r78546mHy9C0RpEDPQfY59ywLAfT1+eLjOTgtwAXr2+O538
lVQAXM5rOWghd9tJa2Hv517V9X3xxVcOMBNdPVGkicS8mTr9xvKyyHUOd7sPWuXo
cIeH1NutZzWTUvx4MqU1VSUSFsCZ9BEa9+tMYcdREYRs0S6zDOsp/F6b38s3Bpp9
f25W93T5R7xffsoS680bL9/Rdw1lcB1PcQwnRCh19nRUqkMc3YjaRmu3TbDQ+Yrg
OidNuVU9Cahcw60TeTYEu+nxRW6vuTEu8HMFuu+DqoIyYPz6LDBnGll2rUIoZzD3
zTMNHObtZ+zg1e2La9vbuhesJQkA/EgK/1gMBQ5pZjK1Udb9CUIaU/XdgEncoU5K
eTr21LGQHRIqwYKClEQ6Pb4qh33w1H8wf6hOMhTQq8JDG62YWR1ITmEfaUh+SHsa
nHasaFwKmlAe1KpM86myZNTPEfnVYVDGb5js2nKR1v2ZeKZoEaBuzsoBZLpwCxVG
4BifHemBy150sOAKFu13o+nIsCtxbjewhTLwByb4ifnaVmBjzD8lT75oqeuVlBav
PpI03wpi3jN8AJnfk2hdgJ4kLYtg7p2hlERO0TJc5dSK6efVOx7EXt4btJpPUApi
x6CMgrldqE5mlggaRc/qzVLQAgSZT7yFYF5g7fTTa92XBmWvUawgq29D7v5WAaHM
LjtKTMdwh1lwUzyHiHazSMAeA+1KEKDIgO5top51I+paKjGf5/vHaVtIpzJWjx0H
0MFtSFohxQjxJJVL6/5z6TDHDdEpm9fA8R3CmzP0GttjoKHhjsoNKyobutGKx0L4
r2C9/Sx7oFAc0Y12mDyF5goJBC1r+5yOT8h9mxU8hFxxeuEvIYvCaThivVcHU3GR
2rRl8HUSocqEbnWVCES4sevYAUJkei/sk/HeFe1y1kW6EFp9qS4m1lVObd/sIT97
LmRDoSGYsvcZJBPG64N7V1iMmh15Yxy+iJU7PGh28UNTuZEtKDz/wgwvLaKVzIIb
mCCrsK2Go/ZeEykfD3VogcU12bm5HFiPL5VHAcoO8+lVloauQ9zHcWVkVEfGF5e9
sds+wBArPjEMQPoXdFPB4sI8XvbYK/nX85rN0IOUF0W+2GVHRL3341XnNlPMgGH/
al6DrNYcsIRk0HBX9FAsRlhkIS4Kms3vd83hQlEvCguEo6zGfw3ITOFovEPRrDHm
+DqtLDjjqkIzXtdBwexS7g2kV8fu0GDVM2JixPdiujJ3lG627JyExwajC++d1QPB
DrFmaQdAQFjsHw2A570JScbbb7ttF1O/1EwAV6YyPAwiUp5+y1XFxGSSx4qZI6RD
mjVE9yFOprSE0BN9oCF4fZ23x3yKnLJpzH+iwmsSrPKZeGRTiFVu4BtMbCREBpJb
LJwXkSiHADJJcIxIxdbSzXwd9hDq5Kon2CyXu3vQ280XuJbFiqb+Jkj1bBY28NSY
xrkGPTEhbaRVViZA4AwwiKn2ZIOfeoUL9vznNa5IEhowPNZjogcqyjiK9WjHOpLr
AvaSynB/nyuCEwHW6YNWy8GUZ6hbrEMqPzgBFDdzFfs8T3ki6ck9W6JFpyovtQ3+
Gn6qwkk2EdpoSj7j8CCWoqUeHayK9KeadPVTyzJGni7bpVGj+CZtc9+PagU8HyIP
FMe1osL6sbQQxUG8wxrUCjQejmuHdVrAwofxfCF52XvoU+GgBRyEK05+XhH2HLkR
Bru16Y53f++FgL2WFGRabKoNooiNx6exseqeYoyQBiEh1tcORMkVF/q+nt4KWMUU
AFubtsWzDxKp11jVRLX/O5gC4szp/v9yV5e1+HBNcO+ZpSbdN0ASNBvKQz8AWgbz
54sTqBdQk9JYdurGZJBHYdN33CN9teiSg8zH5+2pRCOeIxzsfUQW8zj6oWXXso+Y
xQsq89SLNUmyA9VlFRm+7yAuRIXoOjCmyyEgO92pavF78NSmlWpJuUCQgCWZo8W1
mxmy8ib4BEtZs2tlMZ+4WhD9UfNlHfr/Nf+Nz6iFWCogecKYZxDZ7oYStUOrU2QC
v6ZRyLFvCGErTfDsDmc1/8DZB/Bl8vwy8geRllBxCL6bIVWUT3dD3opGuYVAxtpw
u9ff79LV9MNc8DfA+xF5AqS28cvQh3OkDFE+yUxsJKEyCanKKnuL4nO8Vx92UetG
MXkdIgwSy8HaWHH9fmvHVVKE2BqN2g9tFt/UF0oyhfaV3Xx/4OryrAp15dNwFW2n
FAOPRVsROk81OF3LL25fzz9bLpaa9wI76BXDGMgPSRPj0WfDNkVq9VlnYfQguMSC
Z7Xifz/SmTjP9Prm//DzjdE9n4zADe+wJzKUK5JwIs6l7qOSKaXFrJiHgu9TvgOH
Z38PZQpvHOPzV/OuynqlapY8ArykBxoP07H76sUuV2eP4VAIRylWKaSDe2qYLgcf
ZWJJHZFXdZY/Rgb6XrwQonBKSST4wEv/+Vt/4AYlROl0KoQ5MHREtkAOsxkxOHS/
EZB+b6cgEXR0I9UdNz2lmBSjlinLJy0447hNwFhd1bNCxMh8xos+YPhuhxMqNc1L
Cj/NQtJyJBRInjUQa0clgJmhjK6Jy0HApPNMfeQijVcJVUWMkHuB77hZ0ICjqXh+
SWGAG9tWRF0rtN/J18tPD1rmluEVys2lKQrQlHYkg0fc1jrtQrYZcb7JDSyX+1s1
QaNkVz/BSLqV/AAQTAqGjMmhJq1QHrPt670Z1RCziPiLuwzsx0gKLJDsKH2/9hkJ
TcESS97olO0cvOH/bM9MN0ORt93rRaHQw0CblLlIddTBsotd6T0ug3oaR2ru4Smf
1aM+udFOi21MSbnZNfBsaMwBWXO1EYF+aAjwVTEE4LJFQvAtIeeFgYpaXVxlKk/I
XjUfN7KpgZaYlxVLbR8GHQWFwIFZUd4UIO5x0d69FuSmPu+EJuZCryftz77hg+yv
emuP1lsdRCbm7d+AsBagh6NUl0EDgMKukIw+uAWMZW4KdPElWQWcLMBqlfE9V9LH
/cbd5z37X96GnVkAKWrDVCkHvaT6/yKHsPHBwFHtz42PBJLO0MKiupGkmTRrVGQy
hbSegWcm3MbuGXS2UihoWo+If4wQfO/ASOv45I7f8dt1xB0H5xgLoh+gMdrzUD51
43Tdyu8WfmVmx2MQDsR1Iduc3tUSakxpTTUJDcYRiC2OUXhLSEiyUTT4R2csuSVJ
WW0yOsj7e/pZ0Xk+d2lYwXcZYx0SHEa59Ud4OP1G94L8jQ5iDGrz+1TlFQ6dYLV3
6Bczsd63eR040DAQlGLYm07Blxf7Rb99vy+Vd6nppagVXRrJm3EyNFk7G2EBFgDN
mJK6syO70hcxVlxYDwJRo2QrC8zptfMjFyxqLaYeLZl6upARI7fVMzz5yPaxAruz
Js0lnbl5xYbqDcbK8oPNP0cAo7xNERBTMyseqGs4CogXwB2L3IkyMK177t/EMxAy
3dSfv5wQ9gfB/C/hVAWpY9CA72HxwJjnhGNEST0p6GgUdLcqf7uMWzXL5Q1F8TYV
vaSzqeaXnC6/3XacU/Cbd6SAXlaYNSBa64Vi/UewesD0c0Lm+qCyHTvdQ9HBW2zH
eSLce5WS/tzkMZYHskKNJD0I+C0bZ04rliq36K1NcWtS/6ziP8qfwqrYFYiswSoJ
5iJDzUlqRbZ85ZwQ6dw4w2FVDbi+6MRuCH4QjFZ1gR3DR2RJXNtU6hedbry8acKt
NoIM85JWaRfQx+eNCjAQkOUHtrZ6MrZCgNnMRpbOO8z19EwD7CG03pYeKklT7+US
NNsuIKQfvK7Jhx0kCyaarbknmpDrmjGyiMpgG+85YEGa1AgFgeW5OG0RaQsT9fPM
pxXjzynlGtyxch5gNwVzpNFrtY00joOf72TtPOA+qAf/SYLfqPSQUH/jUzCiZuPL
E7HXy3K6rROOySCwc0tk0rz1Ho+/pzSR9RtdI4Xf5q8d/PpqNlskEkZxTLuobgZx
YVLLof0f6KcG+5kzl599dWa6hRmVYqNIxkDfz5ROuxUCELum6xlIYpBE/HII5GJQ
A07A3QyWNpB/Xr0q9sAOfl0pF7Ac5PlUVrPX667AkR5BKc6e1sArdOKR40+r4sor
d/ueAcWMBRSRVU+p1DYY1gW7Uj+OBULyY6RbVRSv2h6cdpTxtPHyapXSYJTGWptv
6kN7tfB9ol/XXbEkrWpV5pwjpPfZxGr+OU4hqRUT1Qt1lpvqM1VPGM7G+irer/4I
P4m/UeVgG0pxqOnxaBASs+MQW6ppmNrbmTYgZqjsYND3TCDG+Cb7TdBmeVbnaqA+
op+bNGfFcfLNE+teuDn+1wFShUTLLpxwzyTVe89UFGh9nNpd1r7cxs5kdl3FV6/3
t1jFnkXZV/zicNTzqBajUE8RyePZaAReh3UUnuPs2jWqt3C9okfRom6ZqDN1zhj2
a+QwjlIgpP8Fnc7f9PxDkiaFlE/4RghguVo9b15jwcaohJCcXxo68dkNkyGVApTQ
G9/37qOPmcucm13CB5sIrxJaApo+iHg+vb1oNbn1Fs8PphqOiib7m5hMy+SGuSIG
LliUO1BmW07dYRDtB6E8NrOkC50BAb/3q35+Ks19U2SCE1sR0zzwri9O6o1Rbjot
qBgodXyYJ4y6WEnMG2nWfPZEMcWIr6nWYgm0ITjlDjN7MEzGr+V9dA/1376X7KE0
XfeWCozf/TmEUAlwHE6IdvyLB8OINkb7w+He+qyHlPqiZ7yRCW1rVqUciEqoWWHR
tK0TqlJfC8uf8IHv/KmV7Q1fXXaLDEIN2/lZXFv+2DLDHPz6TUo6JOxWKAGbV/Kw
wegp53bSpLj0dXUgOTyG0dCTXExp0fwOeZ8QWMq9Gk+VS0OKiiB4xMvmvaFgTwX+
fRPTVMh5nklEeIwomTvG9GJOUl/nHUyO0b4TAEhapRfGl8ikA2C4PBzaE4AWI/y4
72LU2pgEgF3XGuVTdBkEWUMl/TibOe64xoJRfmQyc9yOEbKzV6CrlPmBApv4NwaC
XpyMpve+CWMh5Bs9114/OjQkp/CgidXPYvCd1bYRPDr2zzuB/fafIj7y/LNXb9S1
65MhmWMNyxZwLrJwZC3xzEoG7J5WAOZVLyWwDL2/MIU0JIDZhAvhx1STF8DAGQBH
934bak5Y0SoaVpe7K5ritziVaxSTaCItqQlHzvy3BLR3UUKXR3dpuJY4ZGTfdv+o
VFkHyIg2XWjf4QqXzOiwHq3imdIzgfzU2+P9YqQwN0InIQvCyq7uuV/SyanwbVJX
FaojXfCyVTC5efP5uHyw53Y1aygKWDhfQfoqgU/t+ys/xupY5pBZhY/FTtY5tiY9
wz8WgLoOjSRijCTJo4Pu7i8VKDHFLYl7dLY3BpuYxUhsEnWQZNf+0rUOldope28l
VkBVT+1nB3q2Pcgdm/ptAL2D5Nw2QEpVOaeepGvfs8iPrCntqNHcoxK/fbJhmsqW
DJ2AMg92pyJPWjOh1Hc/YhNfh2CMG70rvLRHj17ultHwgLRo5ciOAqR6ytAhTV7B
L8IvvOfvuvjxXnTxZtJwWUwK9PP1Gd82Z63iOYg38sl9pziR4JLUlyN9J/laT6lp
6GACG9k73EetZgVbH1QW/NZymBuglNfCWUN9qjLKG2OOwTu97GsW/TrwVd8lBEIZ
FZCzr3861p+t88B5LpRV3PZN94aVU6QpvIHNYPPCzbqcyTh7AiFXPdvX2HJDPXRE
zOp7CtYehRQInHmbGbN3WLH6P2Y3dEAqj0sE/LQHHrSPAMiMgkpBtZjAlSec4an/
MGwtfuiymfUf80gmKi8UOdEZX9YnjWEIYlLCyUXMK223rO+giZW9E0sJq7wFnyk5
wfkmGFcDE/4D56WMfCoXAv+jbo8P3ZiQCMhqD+OZ6a8JabooAN7TfUeX2EjhutGc
NNLKPJ1mAgDB7E5jiSI6BNs2XGht+uScQ+ZjwU6O+ziBaVQMsgf+Wk5E6T9pa2Lb
d4CtMWpMon07SBv2TCOenfJc1zPMMi1rMLU/oLubJek3f0SCiKakbO9t808NZ3hD
zscqZ0aTIV82T85PCke2gxy+eL0nvKTMvKrNI8LPu+7gc/p4/1a+GSK0ADn8Zu3h
23Rc9zkwurLMLnhFCYaumCaGMJvJnFzbx4TdUoesbN2mE5JQ3f05j96zAWo6Navd
Ex7UITKzAg8INJvaQCya78r1XjWlWSaq/MeAN7/3sMPGQCklLjzn2qdQVLrz5E8/
ykq5P3qpA4asU5ipPeWgvqkbHvV+3vIONuDtm1G9YBQr8gv7HPP3B4+m0Y2hKWfW
nlxAYXv0R159ZHS3/04YcByMe/TNAxaJRZPPdIaq/uNDQe/NpQnHH3kuOnFxIG4S
7UEQpJkt2bUoqFTxC8Brw8MNvMnliTKRDa/UuGTvUxuanV4/5KG7wFUMygSmbPLM
H0SrtsQr1n10vJGL/ChI9T7/Rk8CthfufV4iJm0ejGHFUXsEFXcdQ9Xuf/0GX51A
HVdPYo28eQqOtUEY8XEf3knC6XSoAhrXQNTi8aJOOJODXQU6QvUJKms3hQ5Otgwx
fAtEHrV/I1H3EBv6TkGPfyJefm/3MuY9jQqU2b2pyylHHwAmo7QbV4OV+mRnyLkQ
O3Q3j1lRNZzpBm2cpligiNBrRFngnkQaxmFCdE7uU2zxUggZuPMRhLmDrpytoqW2
O5wQUcJTq9Urawqo1xtE+O1A8MlsdOo5pCSEYz70W7Kt5G0l8Rj0BpeI+UmXoHbw
W8PPvXZnRRDUftyY0/tGaTb7D5dMu0mC2t+v8QIWDh1LBPPbrpeASPFK4PmQJ1fA
9MqVMt2GR1tmkiQeAL2h7uFmVS8wyyw6DVHVgo3YK4n7eJzMqv5Tz28zOssZTN/+
rD9P3tSY46dgw0k7gnOVhvORDRmOsuGye1x0sXzG3nziAmVMRzptomTjEmrL5Gjw
Tc0ojbXuWlf0DrAKDPPZm/l2s5WUoHLjXXNzkqahWI1nBeTn6VnSTLg2zcG3e68a
kedsEWEvPkNWwhWlO5lLixRC009wRuprjl1BRQdx3iHqagumeJo0Kc4AQZMyOUZw
0g0+9a249iEhcetTWFuyPM5WcpEuW6mcqWc2eymexBwVuBZSeZuk0pAZwc4Aep+V
OvvbdrVvSk7SRdTokQgpG4TH95fEcpTsJERAjho0l5MSkannU3lgyUe+ohqHmrMH
8SGDtDKFxMDJYDaUeiteZO4hKa17Izd/qH5RsbavMYxQ8eCoW4lyOrILbxmfm/LX
K+4zZi1LMQ5Cx58NO5r5GMOOXisv+tYpBeR+5MB5qhGcTSfTcoNgFPiW+Ebv8H0B
o2MR6ckKyOea1lQgO4cP3zMko4mIE4AXICTFBIK3Ns0nml2JKrolQjJ4/z/CKcH1
5lw/XgzVhk07WqsRqhiOxFFVARFa9KruSfRAS75cjri8O/lmkJJYqGh748vNTrIu
if80P3QZ1jU7TKpndCX4YBF7jG6NW/E9UJVV+6F9tD21iVcd9c0xjyZiP1W8AmD1
DKWJbPhQc4DWxXHC+/c1WXdC53x77d7YaYDYMmiT701T5ObqGM8E6MTYpmucgr04
NVrrQYncvugdYcZoFz9a6IFFGAEyHUgT/wlE7/k6//OpIkwIMcsNEyaBX5bAvZZS
cR0F6khFaSW2CKs4KzjEfTNQ/0d4HiGc3nC22tLaiSMgoplAaq5WafmTvCJpj6lp
fXVnxCXFcqeXvxb+KIp34AZ1bKfpwsBZWOr/E3uhoS+WEIxJdlBOHUSlmEYg72WY
vdEVzDSGVDG5pV7hRoiL35O6AP81S+j3j6NM/hYdfznSI057glO3qsRwX2ztGyz4
tmA8E+tikImhQlVEoyt9Sg4arpt2I+oZXwv5nQSCQ+ssNSf5VxtGbRll4OFnlKlX
DDM4XtX5f1lJYaVyOaABUAE9HHTszBP3+d7GoouZkgPfSxFY1zFhOlbyX9+tR5xw
2UNqH55DC7UPJHSaN/ZDTkbe23UpUrjAenEPH4Ua325vVn0z5QmOy69FezKajCMU
PkaYj0usRbcRzh5I0feJviZXI/GkYfvJeU+4A0zldxMESZnydpfxFTeNs6cfM6e9
vIHYly2Qp6XqMrdQUdHLcsg1RGYUh4fi/BqkgTNlpDWk60n7ccWOupbUrFNroygg
2ocJ5WiAfYX/oa5VODiVVylz9dJVkgFxhaNd1Pig/ATNgYlR1ixKyKAKJSdQXOlk
isI4E4s1JgnxWGQIKEyjh8DF/TCIxdjGcsgBkgRwOiL7bwXxt0a1Sh7OpJZ8Epe1
77Ad4MeGk8Lvmpv+uw0WpnLYCrLH4c3Safb4319LMH5ISccC1ykg5GDk44pz122Q
CA73xRxYgLRooCKRSZU9X3ddJKV6TQ0ORwup5eWN2+zwxq+xtv/d5f6e3MuD8lnb
2irEcRMsgnRcYHTHURiaXzffkt3muy3GFeQlB0+fLQ7otQYcChgNxF977aL32/64
xMTKLA0rrFjKng0G1yd06noZR9PzQog4xIHRFXJiYYWNX9OGTHTfHYwAvzg2CAB0
27bRuqPWNCzGUPdVMS8QRiKB6bhkq2MUTi/tbXO51fp22XeKVl3vkAF6Ep4brWfC
e4DN1lVQsTnFydz3PgnojIf/Wpd0suXNjYR0h+f1pQQNaunzZSWCRIbNk2OIHImP
FDsOE4bAhbsqAkrbfrgInMH8aq8l48r5K2VpdhCJVjRERMK61pHi8AfTwM46JTs3
fYW9+OEI/3mrHnNIE2XWWbqo+Skf4IFrgN1jC5skhy1/6I3mjgWkO+/mQ4ZWFom4
PC+2iuRYj6IK/zBSx4jXEcJOqbEpcFS3PFf45IviW6upUDurhUqZhV3SdxsPL0Rf
nidlmHPh+oohIU0OZ5BAdAYUSzFY+vQMqSsTqAP9lbN5LHHyb2RkceULllYxkOCN
ABBJ5aBOCLrFQq8yGfNiOn7wXEKKfDiXPxdzDoZc7Ti7oTFVWkpGLQPkinFusK18
XOkav1lIOTlcStWNZQ9fDPDi5AXn32EurzrMXlLuksqdcgdqQQcewiZu8jOT+CXw
YxVRYPBrkw5Upy1vM/btzNPDaGAsdAgwvO1PuhTsHmyUD6Ain1JvaEucczDXT/q5
r8FUn8b+jKVyzVMxKYkenJN+ujp/AOAeCctSrtKyhHuKS58jt2yKDl6Qx3MTqCgU
vz0iVNsld/BCShTEFzxqXVW0FqghUcRSSpMZG7u+/vMqLwIDucBiJZqQAT6t0XoT
M/GD7He42Ba84ayHpyTynziKmcNexANZ/umr8MKe7FIyIGwRLRQboEQq0Mfw8en6
LwCVVgTGQytHiY9IvsUb2eaZh1yHo4WD5dpN7XKLDb+PPstleNhdXt5CU7czjl3I
/2wM3CmMYlw0+HdIGMLKrxpns9dq4a/K4WByTjjhbJQ7jwlG3SDa9y9lREHLVKal
jrpsSa7YOJm3AonR6NF5ae2PK9RBkF70UhlVp7ng4lwWltqfO2kiI6L2/t5ce0NQ
MtusbGy/QkCoUnHRNM5M9KADvG/Yj6RvzM4QZhUpl4iQb81NG40hoWc043sTndse
+GRVHkzcv9jrbv5twWPwp5/UiZNPjroJ9kpohaLMwCey/8BpHyTiUoyN4vR6kpnI
X/fCRtCu55ri0YZdsl87am2kkEL7GLqJZB/BwBGD4YjDv/uN2ZSygQt9N/tgEqjr
iXLON5KHkKj1DAuwqSEeZ9NPLxPnzaNSYtgKSsqV4qjL8QyjGgR3WgDgXVYN2rZC
Omzc7jCKTC4gCcCTaXQHgg3uypFio7QKysVinyIEN+Y517QXJ6zGN87I18nJcIq8
UGhq6c1sjhgkXgzDLRfDEAuNwFfY9jJIfughiAgujA6UtH7vs6Og9JRTgjD4B+oE
QMDSNph93gSAUGpFE4DpqoG0bmBpoHs+/u6sY8rRzzZTut0q7nd05jJq/iMNbGqm
8rOylC5i3jwZFu+BYaKzgUj+BpLiBPcGOMgb2Zxcms+bUwk/ImWjbhWia0a6ad6J
PtAWME2VdYEQu6PXG8yVlenD0/ZkX7ll5eiC+OtUi3EhGKiCQsNESuwCvm2hSgEL
w+Rjau2tMk+cyqQp7hJ/57iSsKUWvovx+V17NX4sJQZttHiIZun6WIe/kEStOsf6
iL1PPtwpHEC1671dEkgyfCDNxVx5756T5Vvv0/nhwRLnJ9YL5AApSM7oV9dMS935
WulI+3xBt9pNv3PJrYC/hDFrHhXGTCRf1nGnLcQsQEuyFtG30XF0UXJfcOpdkgxH
/3PQYNILdofxOUYoGjqpQoaEb0bU0L2jAqf+KljrpPC2gWTCqVWMTNqJqbYgWvzG
dnHN6Lr7tR1wzBwasqo3tDGg5GCfR8AStzCx12Anvu+Z6YIrsGd2HTssXWJn90u/
dFjEMmACM/TH9NbGCdi+7GufpEW4RUhaLu3qow5kAVz4q40AM7yDHCOvki1xt9fl
0pcZ43gUIFlK6tOMoS1S0puwYa8l6dnp/Wn6x+3g3pYh5Uc4kVra4eooWrKzlS6X
rAqOPJxcwqGLl1xNG7kXNLi2UgbYGo+2bQqkqXKewG5IB7M2FUWHtIORcf8gPevi
OdzQjTvcsT/peeaLdrHFHIrdrS2KmoMcs1cEfV7MHM2f6vmKWb3aef0ip4fKzQYU
7WbmTfFAu2lKJTFvvHlCbOwyTzO1g5DFBxNLgdR/iPOa94v9W7UOR0qkTVvU04Rz
I06ZuKJIytV2ixkR2DNruB6w0rB8HDrj65+0Qi1zfSv98HijgL7mDxklFRF0u0kT
IpJnCKL7pIavzX5uTYzAGuM+LVUatc/Z4wzJMnLKiCqvDlkiKGbrKuHiW8qayiSg
0N1vitPFRpM2GFivEdiBzhCsgFRUIPbrD05gACz3/vfirTLYvHzA8WdRX+257Z80
vjT3Dg/62StCUnaricLrpN7lWLbkOaiHc674p6o7iGM2lMM6BVRrxTA+h/3XP3uh
q9E8LR5c3NFSlqDnnG9mtUc0V7LWRUWu/WjkKX2Vw5pjVs4VufcpNOXvJpUaSIWs
Jx1jl8bQPOCcT4BIO43DQckyVU3VpFWBhAVzF/2WN1EMgvgY0GitVZzqAIlZwNme
jw9EoQ8Ud3ULgcXgQbnCXHgANeG5nh3Y0T/Wx76diZnkDzF7BlNXUsXLcWd+pe5M
VCDuPJY6UjpFhzupGCH+KX0sJ9OwToOQGn77PIU2nr1fDIiQyrmHH7C2KwJ6aX/5
9t42rTDKB2mqfoiJZ8nz9DlnkYYx779xGKRzkosGvuiJiKlTROBo1CPiey0MbSZn
hNez41cpIt+8xd0heV9pOxNaYz1JiI04k/raeIuBKRF/AyhsRKYHU+AMFECKPpS3
bmbKh7HxMP3PkKHdSapHO8LMd3ZeJ/4b8ax4GWbr854X9yx+CcLF3K0mJhY9FQrH
cCPxRkU0NDgFcSAE/lCEOVfMlpVi7qYCuc2jng+u5Hri+B0q4s4N1I6Kwxt6zHw0
D0M9XcEYIVUMiRechkiVZpw7yW0M5xQAf6bs0fgm22OT1KwFhLXmHip9eXrR6rhF
pSagasa+r6BdEjxcX8wltVt0QxzO50Mjf2Ch9VU/M6cGrDe7MH2ybq8iEFoPjB2i
w3yZAo9VUgI6bAfqQYFaXFNZjaay2DRnuJlM69/DFkhHkqmT4d5dlCHMbPRIptVR
bfpt6n8/Zcyc1gm0UM4e/518jVkSRwG4EyB2Bmw9MZDr4JfRwu6jkMUqvwNo1sNE
7y8Ir4x5CIf1QAGg/KiH1dfaXDp+vdKI8tEWrilFniKwYiA60Kf0KW7tgKitg3mP
J5MWIAlKXfHf7xyI2UGza2bpvX1wi5QSAiYws6fqA2gzK9GkXBELxYepSnGZHCz0
4SgwbY3y5dSWMS8LYbFgZpax9m1184EuYuHs5/Wni/3WNZLQTpwSfp21OT81lk86
4FWsUb1QQTJEUvPvCMWCTbajTdu5FwSx1bXptJWSJ/4+jX9v1K09GbBT/hWf6dVH
dXXVnEJMum3k+uMg7PlCyGgvczj9z6ld+4aCJHygvMDNXl7WYS7QVYampUX8PTGo
Sh9au5HXFjvbdXNNuKu3NLSUcP3xIhE2uoTPr5BX5cwJ7bThURUej4CuyE/e4+uA
PFsS06mrBAT4FLsXKhXanlXuzPnuOjS/kltIExJqbLzl3eA1GczZiEjBNFabjPwN
1+9eAMpFnMiNApxaZU/BOFAc06ltqOuk41J8AIUavWfchuyn0QmMuvdICUJVsTsh
B4ykNDCuIfObaVlZxsNlPDgNuwwiMTVqsCe1z3+HnOrTy0WPxgM30O7uI4tADtrX
0kuC/lMwyTB0EqmmXaY7OgGB+Fm1zgMUEIy7AYp96w5v6DzFSWrF6TbV8YhXuWyf
d3QdxGaOZJR/l7VWVa6hD/CwVQs4jTWGq7kp2erveVka/Fvdrew85Kc34UlYsuX0
CrMW04Ut2EBwGKG+v2O94II4bWZEnC9rGIvodAlP8111LyGA/bTHCwWdLwoGlQPK
mhCHnEycz8n2zTMtsvGw+rsthS8XHC9Jg5u27s0SjMAzPmF+W0ixwcJXRgWvDOso
jGayGohZcxuKDGx0h90ywszbI+Bt2X7r/z0WpHZgjsGOt5ApH2qRv6SZniUBg5pK
yKiGV2Hf1WjHGO9kiIyrkN+xHvVHizJ1nDIuZOypuTDyZtGDX/fyrfkRntPOGOiW
eI5xHEZck3a7UsRnMVzfXGOHlDs9m4mxh6RvUfLPakGpUyxosrNf2+GYohx3xBvI
o/CcqCiZ2QoN6kXV6DyYY3WWfHo4rNWfPwrH8r0eBTAg1qMf/Z3fmvp31w7/ujjD
QsYNpjL32mKDMTxSKPLUwM6tIq2k0aTOk7z9uw5s8e2SLmP41Hikw4zUvv0KxA4z
ujUwbOZZ6QcVfZ85Lu/TmD+qonBtBfB87h7U1uW6Do7b77X1FptLlxH29u6gjsSu
oCEgxyAPFkkvI57gO2IqzuRJnYCXuzSLUOUNHRYdqrrR6ILxKoKVCYC5VSDo9h0o
rvj/HVS8GEjse2cDUPiypOHeynV+Tu3AHq65LuM0Sdg840m9shJP2w6gQJSbl9E7
71x5BlvFXdEaV0J4tu+veY9JWEVk9iwTD799nOf4MXGkV76lDGS4PtQ8DS4xALAn
oyDcUHfW3MHyKG7aJ/F8OcZheqzX1Sqd+m3nXPCyiOhFea3XNP48yj21ogtc5/Sr
0O0abFjrAuHeeeOk+NRhtoPSffTAIyjZecC3lInqnYoVBS7pcjpaWgI/8Mg7M6OC
z+FNJ8AtfDWOFAHBw6Epj7yamt528Ay2e+v23KpmMN2X3O13dNQwPdrCjk2AleT2
WR89xxL7N07j1eRlJaavITBdM2AhZ6Djhu5VKrRa/eORxctYfB2TG8wJxMQS13VQ
fn4MVZmrZWpmRlAzEcclcdkPktyL9cafdKWGvQOc7/9/HfOQIQ6L9H5Fd9MGkiug
P9s2CocSSvDbUIN3I8+o8FrW5RGBsGZ9/gMD5YXU7dEcU3BekEwQ3iFQ16pd8QeA
FZPlYdooAdIXLX2xUv2f3nIxQ0AwopkPOn2Nx5pSmz0odKsQCX0hnt+InFOkVLsC
klNlTYus5XyvovWs1YPEtXz+ByGHhZDNjVvNwETmbZgFknWnC3enyhRBD397MzOA
MIIz3fiWOqnfgmuVzUv9n1OI72IchjmW1PEFVNtvqw9vfAHJN8KQDZDHO5ZHTc8l
ChU0gdOtCpFuy9ZeRYMkzoGXUc7TE1Djwh7dHq2OXpBeyCXw/NJnc64TB02x+rIx
Hh+9+ihwOfAJhzllejph+ltPU7ovOb2Osncz3iXlGLrIjkEYm0S5eQHC8Dyzph3X
TbgkK4vcmKSuMqQspLe5p3axYfNUL4q+Dw1odQLBmllXQGiVN01i+Z/rRnRvD8Fc
7digRXARcPfiVwJilPweDuWRP25pzzFzEbsbsSRBQEsqTnFnLvx5p9pXtzCbXSk3
r+PTu0xI5lHiF+tUTsZefHCIbqb+54Kp8cyjf0LucW8zBcL7q2wutN7zVDMcxrUY
2ayclj4fga+UuRVV88gmE6EjXNqrGcA7YbLZ4cmRp8nYXUd0pwF6uL4OZYoAInqu
+ijHemVLwIZ9UWLjNrvTgcTSCzxeX7JTOq9ky3AK6CNIve26iK895o/26zxlicGW
ATSNdTMqXgEbv3KR0lqhP8fAK5Qi1JxdrnBUjub9tLF91Th1DSycAzOz/nnle36W
5tzd89F7cCf0gotcVQIstlVAfHIh49lxBmSTwU+xpISm7kOaDCMo7I2VHsfqzm8x
RC1Wl/+92JYLHpfA0SG3NOwgRV7tGi6YoTkViDcmgFDC80pvI/BiSiKHk9HPzVUI
HSjnhWLAce/pYWYuyNmTPxplLCz5W7RbSaw1Tq+3p6UyEQ5RmLTBaxUOZTQwLeyd
+VKAf8yf/CF1+YywgJ4HnSz1biF9799OMipzZaHWR8Ru+p99H49FBRLN4g86FLYg
SzVStZdEOZok4Rn2l1TAOr1JOsmyka0FNYTP+I3rkzx6SAr4LkbbxPahmzxQmgNM
L82PrgFFGkB2DcAMtymsf5bnWRQ3RNl4MGp3CIhSNtNfVB5qNeItl/s8fwkme7HB
Ndzrh0CduaFfBrgAKw/1Eeo+cgt+c0edxqL3dYW4Djn2Ig7lqsKL09Si7elZtMY8
jnqmiZx8tdFqm8BFc8drsIkgXoQ78mDD0YuUElZeu+mSg0i+8JgeDWo8AJRUgvCk
ILtzkt/W8tdWQVu2ODuv+LJEI/tZzwTKTKYPziXFcNpzmZ3qOXZ8ChbJ1L/jN0O8
JOGe3coHmaxQHJBN8pbFsGw78q87eGDzpMrzf04Ix0gWSEIaOMjckJcJjzqC0BoY
pM8USQaXO3G8Nr5K5PJSHFbBdyojlT9T3Z6MyM5lqUFOHzKRUEbaMY9RQYkR3fUG
uG4SV/F3A7ndHEqNlhSjFbTEtLYrbKKunGRspbS/oylTj2NfWHGo6fmMtuFLxQIp
OtHUwZuhI9rYQ2xji+cr4vnmyn+t3FzKi0a9TiS8we+M5cvhzexRAaaSofrOgk/2
nfxRA/LGqawk0kpdcYqFOWuag8HMy8CGpjbfXoE7UkPDVz/Qmn8yYJCOfA34ur2J
8IK7DvnF0INqq4ED6Cwp6zYmSnv1F8fYgehrMPDQC2rYc3oTy/IIv9Xof5sVoxkM
lkRhJMICvdKjd96xt3HVk24nnEvPgXHDL83KZ3VtstqCzHGXRiym4zzjFvxpfET8
zm4VVBmCR6vMei36/ROn9a5cbwIfcJlkTnG9TD/T5CmzsVoxxFtwLPOlBUJDhgK3
haCXBBJAKostdFRXBdgoHjyI+bI6AxAzg8VySXKBPjeJxcp63d0iufIY68K5Ywtl
mthNDXIivWKCMUBvqFnS4qYLjMKsDYaCmB1hxxVsMfAjfa/KVpxblvYCVykCPNdd
nON8Fobg+W1+7TRj9eg8AQwSFmIx2TRRQ2zE/NrD5ElgOnfPHw1wB1/uaYiRn3Gk
iTrn/sPoV91MmUWPXjWQenZEUy6yHkdLbZ7/+DFZ27NWIPn9ugAPZAzL5miE1bzn
3uEl270etkg2fO0/tJOVCB6m4Wk3Z9aRawurxdvZ03IVIKsHSC5h+Y0OfYtqMtuG
jIPQqUn+5V1K+SrsynCKl4kwFN4m8ZgaXaa5QvTTXh/t/74O32u8ayEmaycb29Ib
bCrJbDWwFbdApqLec+3SGCPQCfxB6mbrJ+f+bZx4CPJw7s9rXkB6qXHQglxmSOis
dTcqZrrna4L4T1o6WDGLWSqlLMBGD0Z+yEyJpO+JbKMUy31Wxl69U0FLqi72v1r8
dmYGmXL5mwcL6BNgTbEl7o+1v4Jokj/hkKgJ431BmpZhx+P4zgJTBzjwqa975RLt
0CsTZ/IqVikuCgA2Y8FOXpRYkmKtuhDxEkllIO8EQk8QdFyePPaUFT+TwoS6mUhh
CbxzHmHu2XEc4SZrIwlQ8rum9KMizjIk/KpsSXeqvW0hDyZriVruv604zcYQDZKA
2gVOE6+roI4/sUWnxt57PSWF6fAoZGBmbwN4hb3PTJ35Gqs/66uSHYC3XtukbhVm
HXGLd3NL3PuiqIDWAXmpzd/lBNMrCD5T1gvm35djgUD+U39yXD1Id4ZgKy7UWNhz
xa8UN1lADSBtbDeObhMmyNQaWaiZozQmQPXsCD7ib6vyptMXDmQKsPyOecHYT6ez
6R4OEHF04PAp9Z0/OlY/W84Ousc7/8rLXWBmWyYJ5Ms4C4upeu8rhaPAuHWmh7rj
bKMWaUpYFcjVwcg8x+P92Z03qGeHBpphceOnB16YX7A0A3wKnOKb8QQfpP0/KINJ
4Z9w2JMm7XR4jetkdwat0Vco2tiofLXgCCqBVkWV6avI+8DHyx2Kz87aGVDEQNPq
QRXpCMjgrTpiomx0GyigE4YO5XrLPj8Cp9EOrLlr/HUVi5FS+/KsTxtO836bSTW2
rzRL7gt7xdOItSqCU2VVmDHpRAVkJKqRFwb0e/guGsqOVX0HHDGcbyUgYo+s7thk
CXEXcRTwNQ4BOQKGR5xAplYmH5SN79P/hJxUZEMjswdXL6XTP6cLjb0hOpVkOvv7
CVKdqGzEU0NSITxOyg4Hw5LMtumoLVEHy2fzQtK045FwgDVH2XS0JqlnHuVGmc6W
BGtDt/v1n2OHqQiNfMKDc/Stc4641OTPKoonHKFtiTjtzHbBTtaFh4ngdt/yDU7x
Lg+CVWJn+Ye64/60+Dn4TBol+wxiXkSOzxWLvqeS2gdWYeSVdEV6Yx3s4mtezwET
5Dgbk7wemxpIR1h77+wgj20UZjEzlC8ZkVY8HNnm29zTAeZ0GUIfceLyNpx3hs+1
GEzZr5PDjGeBRgyKA8naeKoV+1FNBICoOidPFpdgfCdFeDk1KOpp5fXiNY1xB+Lh
aROMTZAi0f9apSzjU9TW+xvxQKyGpFV4RqNSpBFYZedtVaoAmUjy+KzEX7CmJRCD
K4j+HKJrQghnsxIYSV4Xh4mdE2xlzhSJuozW7Gt3G9CRz2E6qaYruBfp0AnDxLkY
Dkmw/YkiVyjuoXO0+n122Dj+Ro28+SodmulcRsRxFIk8MVLFLyyV8tBHLGR8ONNG
UxGaXBN16lTjYNVEgR/qsQzruVufGROVl0Pzk28kuLg0ZP1fCZzKBSBIOP5hRfy8
j/7EzMs8P1FWHKSO4lbjwehVL1EadlnonU2PxzvEas8NDKfoOUf3YQ2RIhPv50E0
8/rbK8v78PGc7C49jkRVVSPo8dPs9EsAPjyWjNoW87MOc71LPFto2DCaBohGjgu4
ysN3KDkwiN0rjj8Lbav0McaMRQcvqKcnkmU0l5HuWNqtNVcMvMSDNUWVDvYN7WJW
yEc4Mg//wyDZ4N+XA5zprqJf6YMurnCdDML3iJlZpVWTTKoAkzTGMx45OhIj2Oy1
LiYYfKc6rLya8mIBakkslPaYyMUnOnPRmWBvNPlDqe4uvfSQv6zxPZBoLcuY+8ig
p7WQ1P1e4K3gpAbFiXPQ58I07Xb0jzaFN4d/xbWjVsJYZh0J7DZmTyxgCkv5PEBF
6YLNQKfaIe5xejA42WONt+FNrneoka/EFkO+Nh1FHnBsjiID6ShfWppUCPLUXgMA
GzogXpp9FodUNok3+JzNAkkxLhG/kd1DCU8BlbM3OpBgAfXFyonvkrLkN8joivUp
XULyFxYvtRImIftR7BOOtNH+1zycDCRt2a6Jp9dIMwYYsHsxOtMqXIwrhtMBOyLi
zknXZu8zg80KAIctRR6qs0iPISVBmFZgjYDYpeovzwjz2QKuyJ3LPgVz+rKYGlwk
pJonWEhbBOTqtlIsaKUWsKyAXFxjfqPp+UltASHeR9G33m2IFJI+6RdWCSneCu5n
8F37uZirCGRTBRj46sBFdnU07uZJdXw4PbqsRexGY3QuMT9ae3X+0uAUst5s2AnG
F0uasqxbmK0UvtsfAqYwdDGN9UhSe65gOGYSNsaoTuadVxjQPBCiWRwe0TfIcBSC
q4XQK81dCJ691Ee/bZT0IlQF37rPsrzyIElEJjzPMiXPoftYXBZi0ktaPjHa7nPU
UFZtz6Y6i7eqiOeqvn3E1PRsF0RYWBJB7p/lr+zn8AIHH5j+rNEFWi1F/ChdRzBu
1inwdnRyEJc6hovd9+C8lhf1a7kSDtRYz1kUlrTlVihefbRnGTUIRmVnfftfygFP
5J0G/vCRZFQnoqtZtNeE3/U620/nKt+lVGBJZj5CLmvvTnF/ehx3OELY6WWHSc/c
VMLJe37VouqqBkitHNB32tkcxQpgT5EoHIvglmydgKd0ogMUsq+lQqgCfg7bmxtn
jlK9tsXHe36vi9icIUfdOGCKGE6M7E7pAN5HAi3mTCppjdOOLbAarxpUlrWeQ3yj
A8h7xvQMS11S5atqp0cpKD7ZGpr7EIvNSTAxa+9Cwly0Hgod91/slBGxJbr/L3Jq
Tfwqg39jzUilHmHcyWiO7aCf257NVJ3ImMffl8GZYQFdsGA1W3Qt2KP3h3VKfw6F
LIIxD/+GYrfytKwPxAlc5o4xbIO4Rcr12rYVxh4FlTLqkjlURCPKXkix+903Fnz3
XvyQfVgKtsLSTfH6gXBQ+1gwarFtyuCX1Fs+wtR9vadAZnbkW2ke45Tamh7EG2B7
zfzeyf6y7CvxLeqzaX+NMwrz36QSw4KHZGkyt+EqzOlllw41B9V4ADhGkgo5s4ek
yjxtob3pzieE16BZr3YOyoFrkpwF17uVeME3tP3q6K1tHXMLv/9IFM+xSk8rP/Va
TnmIMEol4IGfTQlXzljN4okDlWo9yvjtfCBJkS9dwPVEf0MbeWHnn76CK4yo7mgS
HX8BfRCUkJVkmUGoFDV/DsRYs1l+zK4vY6CyGjBR/6nhyjSD8CJyALxF3e44R0Wo
tlRHTmTGpQ+axwA+PCziUqSAA1k/Vxi766K6/RZlaCQKpP0myb71GcTolzjlwRST
AxXgLS/IovTsAeuQzqjlJCAeJR6mKd9iZG3Cv86YYzEJ+qfiQBcKdTqaCOiznjGR
d1CKVj1v8vDPXDM4bpdCVlIDp3iVw1zRA5RtVSicIMpPsA0ZS+qMu6MXZsm21XRL
NQi6cmZghV6wAT3OM2dZ0qzF3WuLHrJO2AvT3AJ4Yw1+mvHfHvJvRuMqf82BpXFu
FOiFhbKym5PHdOf1uJWomNOMPEPEySFXtYzGR1Z3WqAgEzwelXbJ8UzoQBAIIEQb
M4+T7BOlHZkkUpxqlHIOz6+xm85cr3+iVQGkewlGK/rOEhQlj6hhVmlAzOFfo2vL
IFfwuP3O8L7mRzAZ2rbTF9QYPe7LOANva+hueG7wTVTkupsf5ASlHB1u6BMByFlo
xTPNgAEfQTrNXQeMUdvRjgjPRZKLid9p+p0s9QNrwwKsd5sn73+BNvUGpr1JFR6s
UIR7ttMhvPtBBQmF2BR+TXeYhi8NbN6U1mQ80AMSk5IIkLy62VweXagavFHfNLk9
+iT0Vi3Ghtqqd3XdmB/t12Xkr+1blW1cWftZTC1bRB4ThgOSQcQG0TGKtySl6Hlb
aTbiaAeQ6zRounfM5WAE34f6ugBilANCLSEf6FNR5eGfj+XkmZSyqzBzJ/qJOLR/
UNEDuBlSTnw9MdwZlUJW2yYvZDceEIhOl88XdIlY55JXhKUgwTcmrpWXChD4jmW9
qjI9Zk2m2H/mkY8oq/F6dSROJM4OZxisYh+CaAxd+GZ2poqfTKdmGZxUy84Z1Q7i
8YlW0rv7nl7aqJr2gNZPlLqfdirzVXRqMJfePxiqAmDtZATwV6XD/OTnl7nSCsq3
yzY45gdHHPolHA+nwAzP/cNoMUNkLCF3skZZ+WWmVeAQoXyQsTQ88sl9MuzSOUHY
sjMIUob2q2/DZghuXeLWlpyvaS3HYYG/d6Sko+OEA6HOBOSK31UXusv6rczYLWcJ
SBrwhNOIQx8XuAoyDZGEois01Z6qr6dWeJFeDY+XYWw20TZaerUE8c+1eL3cZ2AE
h4l8/MayrNRCeueQcNsuYCs6TwHhLmCApDbUBul6vf3ONlaszhp/4Wbx2JjBrV7+
thG5QRtx5MVAajBj4wwzp/jEBlXx7F08Jidz79nO885PHFfqDWtuo8CLSSSrPcQ7
KW7an+dDgv/BWes3WznjWJvTCK8+JxVsb2Srt0kAQRS8vSo6/Ooi/2tFMUEAD24Y
kV06l9sOgn1NxAB6PQdm3Xb0AWCsO9uq4MgpRugL5Kv7gWy2lBH9xbSzRCesnl3Y
Uym6ouQrCxRBcAiNCfS3scPmUUxdujHtyEezazFDcTbn+ANv9k/iWyiOJpk0DgQf
rLPvDSsvd0udiLMIkWpU+pVD5+dOjDwQ3hmeR2bPKmekVI2YAeThIIt2jgrihrjw
GxZZtKSavVtP0zESg1Gu20GlLr6qcgvuDod6tdbL6AhkRizAxu+vqadgOK+8qFA+
KQUXDaSlWcUu/t55NBfQoqIywv1U5MZDjSikkpZhvceQ1ioIE/8qBTvZ7cIan0FL
CPK8Q1Mfh93I5DO07u36+jln0GXjK/KRoOsM9vySsIgrJ0p9GWcRJXWR2jWjAXHM
N3qMNFL/8lGDMPxS1Q9daJ82rjMedzNV+0wQPJi6yitaP/NgEkEvaFKrTv3VLQPe
8JTG6PQzH21+8v9YgMyX9ih2ntcyI1Stym/VtSPASh/rnPts6qqg1Atwtm0O5sMt
5cqCewZSTqkM9ozhMh4Ksf4LH1KQxrP484w3cl5ggjT78ikQbxiW4TXgEdmBbYmX
lmL7f1xDvZJ6MTa4vrMWev1BOYzLAhoqeEHoWnLVJFy3B17DSfLeFuoby5qBpHhQ
lpCvgp+TML4JLFXorgCPCqivKcaqbpFvBC8iVehlDyGFaOelD5wlpI607Uu5qTkO
oAEOvBBOrMBFd1R8u6k4MYcT7g7j7p1x4+cKxTGDS+gowTjl66eJKlyzBCXNd+W4
5ePlvBq2vzS06ThqKWP1l8dhjTzHvaCWEcr5tFxhCwLWsheO7S1tuOn1cf6i0lQC
MFDgd/hY26KAjRlVmMRwRgjA8kvdFEX7KJrD4aQuzOhWaMZt2gMv/q4Dy2JuFPtC
LEIGTzCZLzoTMUOdub+MFk6GcarhWyvddApC1ljHEmi8EX/Wo9Ilm6BdxGiqRMyl
qgAzQ6vJFB1NmzWN/A0tu6VQq08G+NAG8LRquHgQqPNZvzGX3s1Un9gGPQO8YHVB
QlrcxP3C7qozQ+5JRC55cCa4ya94ztwy0vh+/SDB9b76+FKVyIiI0vBKcFXpSvbd
ZfxoNbw/auKLnY1KZAsm/8PeEv7mK806n49ltKz8+XVppBDuyqpMoCougIdLEKam
/YwQVKYjEQCYTXCqmbafHDSU9wdbjUz3O69tUqcLehqBY5b41J/0hYdbjedBsZ34
ctBl1AT9eu8AnrRMmlcNJsFgUmy+DPEsqFVvmSN4G4QIu4lgUgE+gQWBt/uCQ7a7
z3J7m1FdF75nf0fLiTnSG2YIxzpM04QmnDAQyezDCO6nJbvXey+1NNE6fMSjXzM3
TTdwGfvHYSJ8YB98ql8gEH9Q8Rr560oLHzVv/zGFPuJ6CibaaDhpiZoPVhzc8kDW
vQ5Nv20/Gp+jLJxXYMUKPbNzt2clXVROF+dAeVuSgzFqMxfOtAx15LfYjbDWC7g9
kQ14KQ7Cizj6fNXXEDtVEXp7IuFOok7UjAAo/MNFz3kwYD9sHK8CcUUjSzcRWRmi
9vPVAgqaSevW2lb0hEkFTAdBtPL6XINgXbO/p6PS486H1ESfOyak1b1fLI0Qn+DJ
qEvUsCujUEJaSshem8alqJZ61iwOuT8LxtDMkkHaLuzojN9Ur/MzsMBiejt0LzRT
duCvIbiHZUT7IeeHJHDOSNu+D/r6vNNsI5lWMGsBiSYMG9zzyJNfBxMQWfDMtcXE
sE0QmiclBwHu/1eg3Kx84POg1N4IOosF0M7nXyTzL1UVDy7priRmJjArImOq+GSU
QAeNcknH4JkXhvgec3Wg8JViPGjZjvm530kUfWns6M0DkeCEhTDWggjLrpfgOPup
THy00+ZSZaAqunUdYqFx2zeUhMr5fvfcQBG5YCSx1+aMP7Al3WoVe3s/bzBcNgZ7
Pw6KbxRaDVW/ewUW0ry1xcJB+8KvsUPpQ2BCXL+R6ocutISX2ELURnzWavgDAuGN
6SdRXljfRYCD2/drsrP0dJCwYFjIx/ZPwUvRhKRG0M3iA9Mk/QAF6IEwXuaicoS9
u+jQlIHD0YBz1LhlfskgMqXN/z5cSySP+aMfQ4ztGsLum3rtWjd1iN9Af6ejVjzW
AuzhyHH18uVokuR6iTUd9z2glDXXx5N9vyYf7cglQfu+1wpYBOGjpqq6ZYnO1/NB
EgwkTc82J+ztK8RjdnDOiQU1FrkcI+cv6oT3mDTGp2fSQxqn7GFmWq1IntEqeeiA
8kxc7v02B6ux1ew1bdWDNXjP6ejJNWhMlJaqBT0lC6+JlytlOPhas/XeBkfdOSDu
p9H7xwIsckX1TmWcqtHpZOsQVQ00P3fZHIYlGYO5WxONdrRyOuQx+95pNv7NgNst
Koem97GSTsEgnbnjj2Df6x916Y+cdEFt/n1jPJAQVPsRGwsUu90vYtHjOGm7idZs
4C7Tk4SgeDOBJuBNtSU5vELwq0+6U8+h1s/jy+9SggjsLDdPfZpAniEqJV8tGCGw
NXZYSTwYsIFcjUu+9L/uYWpfgQNY5gx6WWCUOMA0wWFDyXbSqU7R1lwQuVxy7BZM
Em6PV6/Abg8Un8lZnvF3PlUAb4GTCXrfx7IRF65TIPRi5FGYUaabFUzYQuzt3t55
NR89v4f0vsLe8ExX7h/v+U3t+6+LNg1pUjOdByCo2AcqoGPEr18Y12jwNXH7VCeD
WiFbmjWOyGxX5XwgZ7C21n3eFTPKnjL4IZEMZyVJOSrIO4NEgtKls782eHAU2+ZA
qbIN0MRSAVVzGYdEG4efEOyQQ5/7uyhb/fhCptQfSsWWZu+uHjT8x0K4pLiwVGqz
oAyy0sr5CcihbVvnMyKIRByBW8bM+W8Aa1H2KcIAPwjqawsLduCPBdkIGu/niEak
U9XzsA6yUz5SOSOv9KNQkvpWcRj4FHrTVXUuz6wOp4uUxMz7euLoXI32VTMWqnyJ
H5SRs8xWcLKwVFdt/9aXC01KGWsebHgdiXt/tl5LbQfjWuOxm173fO2m6aLstNi2
QpSO0s6vEiwwo+LAScrDbZ50QkuzW64z38afU2pbJSOKLr/hZtIGVHHK6WPhh8Pg
a7e3y1HNWmCJCCkylL1BqWV/R/AcjKEo8aPclY202YFGAqXtFnUVXwCioENLqK2M
o1e43hi259wjRSoqTk2qeywFYoMWInH4B71IRc0iUX/obzd/WeMTvsA7NsS+woXv
0M2AVJ5XOol1oJTyRBn42X3NyMO42vdKBIRHf3DwsBzGLMteMlUNb0EOOT9RK0pM
z3faS9xtWBqWAbakZYLhKDJoYGms4GfhjoWbmN4IWAv8gP5zi0AAElpkyVOYF/Qa
tJQGZ/6ABfiTuY5Brx/joW1zIc0XZn6/XamKjQNeXLYfPE54qM1NaI9BJWDit03X
ga9qeI+jA0vJEJtAJuicLtk3pSg9/oZm2QAv0kXCoFkux3k6byGWdBSzE8wnqpeX
uZSwYK8+gMAYkgGBuvdMGt63W8jNhi/7dHaS7SN3IQEcVR83JU07pBCcWZXmQWT4
31jFkAOJNPsfVXOFxyK31sQNRFsNkpAk9t8vgAvpPhQ3+E/ILIdvOwjuFQwbcrlh
TypTE4KactJw2ntanz5QwqoOO4kqXhgreHORqxQgR8mLyd1sX6HjV1+9zDD8xm82
0wIn0U+6ZjH4t2Z3kIcBS3eK064FywAv7F9qOPk1T53DMQOIVrLz2HdfThlv/pQm
ALckx6j9akfG4ELuuDSxLyFQFCVbT5qw+487pp25Sfda9poSX7AL13c+giq/mBHg
3jbAXwTcRwUmqAnXQTnhtgjQ98xYsOeijD5v3Sf1Z18DbuC5b0cGzISIlqPfdMo3
+ZRlTgnu1RdxoOrNKbt+nJSaLC6N1soGu6JHfbYLSISsoGWCQ27uVPu1hHGJapqr
OR/r2ysQD2BSFuK1cPTLbZT6uY1QT4ay/oIAqZv3ZOFuXFb+o3tquHN0Jk+yAjuR
2ckvyf3pzqsDQDPu4Kb4nBTnFHbYUp7Rav/k9q/xVzUXJ+ncDToQL/huU5U6oI3F
29+gr3N2/y0CarbrWGbaBS44naXUUkAabpeLXC18oDG41ZPSJ3m+dHuSfoEP2E2h
Tf2HaAhL0GXy2fKuWc2NDf87A/dnBjJL8WtYVHLgiCpWcAEX/J2tox6QihmMixSk
HRBUWQmq0j/fatXljtoqBMul192dOwG/azYAFPqU92Ti4kOaAM5qa4mjR1jBNcYg
jtxDjwpkHZdbD8AslhgkCG42I8A990ChkuYEgZNuP2sOUx6xmqDwKypn+GO1ItfN
1U91pMxO/YwZJPtIDCuESuiuTjTrQJlYnnfyei5Kuvu3SXBiMQJNnR8dPZBYW9tt
aF2sHzQNHNjxgD6D0oA1wq7ah9Bkw0SJFuhh2c1p0q2AfnBtOh9yIGvz2ZfJNIrj
eacWJGW/KvbLror6Ck6IcCa7BSPg5IJWbCDX9BhHlchApNI2VXoupwyW4XEAmd9C
JbJpXGRrKB1rEHVzcbd7jOAWLjjjlIBQ9YA9y/8Ek7wmPGb2Ms3nyNcf2080CY1G
bRD8w18oULMcS7JrR0khHQvepea5Coe5tL4imKIX5x+bOI77iTktHkzYrpaqZJ/M
5V1FY2gFcAryLmr9X2tHeqUfT3KpIN09ltMLTwXS3cvyBGtk1qHQT2Hb52sYxIKB
0+xm8tPIvwwq5fh8V1mkkydR1om9cVWXW5kSBop206FIqwUdpcA3My2c80/K+YkG
SMBZQvTu2pSIoKkUfKWYIu0jKnOkS2tC1SvGCwpAB3lD0TdejILWJxkwKeCu3oxl
/qKVYfm8TafUKLQpNkS22i0hJIJ+ag+mXTl9NjZzvQpGzE1hnmC+jpeZ46YNusKo
uj82zUYEp30J+A4olE7UeqWhAO75WZ6XHfs+iKvETAiJ5ufCtrfItHRrmIsJK1gw
TdH00mXUNkJq556sDbPo1GmWrfoDSwZxINGf0/pPrP825Xsqm1qcP/QHNQKEbJWc
V+bocefBAXZRLJSSJtWkolo1Hh8G2MvMCCUkKaiZEbqCWqPzU3FtV93eQ4fp8/en
wzwAaYkTxc/XQl3E3/tkm1AUKpQ6lcWXFyzoDR7hadFjKOgSEvNEBzxDnOEuat+M
BIzm7OE2lGi/wlQzaGlcZS2CfOeJqg6sKy6oaorxrpVHI0DB13vLNafrc6QLWsql
BaDyU6Z5e5BNC7pqIlagtfAP/2eCdzmViCQGP0YqdcQ8xMpWijj/2564eMorXHJ4
CSkc2mlivvFMdI9BvjkXetBkIOiBZGPjsJkEa8vpGasqzIG8doU/wi03m0dd8Yt3
iY6fk9ayZ74raeNTEpV+lvfdERsckB9Ti/lJdMivaelZKJIYtw79OGn8IWLpV/pZ
mSubpVBmoxe7Y4jL6hX4qiJbjqAd4qLXNAxCF33qHPxlaoNbRt7Fy7BKwU5NCHTO
26xceGS+Nim1Pry5WiO3Jdefp1BXSu6abyYtvJhwoqIhyBBxx/NT8rvzyvej2qlM
fN0k0sHA5Ib91Li385t3w9B91Q+Io7W5QLLRjWzmYHRcZ+prJ0sLe6PQX3jSbNNL
jXqzdxMPhDDXUr5X5bOUvSj6c7TdkV+Zj/vNZ4GVvMNy9V2eMAxIpuDJCCp+fvp/
qgFzaTjiCNR1L2tA3SZSKa1qH+9ff6At3RMv4Qw1iuqbZ55ngGL9uL2e1Cg8DNjM
bFfCEfGl5tzpKQFQyeJwhYnCieUh65ytzUmrdVOKix92nv9xyfJU/4LGoPuYQpXX
1WWqFLGQayIqP86JfoVmY11eR0YZSfVbacTQO8w79T7fsBkmUJyoEyFRtAQFlC4w
VWf7Ccsa1ce8NN0dT5pEPM5Pxv9b8YrR31fIpIkVHv77NM1ceW0wyVwbJ5s4dlQN
3V00Bg0YSa2tbCRFMZLNfRjc1wiD9wPKYQwRTb33OXOkukwLpDMxnqPGaEoLekUg
WYN920vgu+FJg1kx3oDgKZ/0FnZ0QXtfylMVflL/RlcGNDBt6+TarEOMlGO6YY80
oAUd3IukkNdA03K1AgCZlDl1mtMCyxqI5pRQ+TzDnasm6SBvUpre1IvI75tCYktd
yA0k+yVLOhPofLE7YbKx0rvkYwxgb/qUTES3inK3ZoFlEYLrOPVvVeU/8W0O2wDL
QGTlvBYHhnEVwFSjSrysJ0HrLDVKtcPmBy2ZDxVzBJD+Ju/oK8nJ3ul6E4Yoj0Co
PU8hxba3G2LC2iULbP0oc4kahXvSGuemDygyTa0Al34LqLv7lTd6CuulXeqte1g0
Z26T2v4OKnH3xEaHSqRpNCSLfGhILw1w4ENqKpmcF1LK9G/1/upsJb9vLOMxd7+O
chi5nMjAQLarwUi+qHr7rQsJvHrfgV0xB/xoSJSXaWTCgtxuJvHsAZ6ENqvCn3Bh
E3K3EpKQDdsml7yvDz9TYHifQnF2e0yMeGYfsYf8w/vmnPL25AnQ4qo14I0cAUR5
NA+ra5ctJQUDosCJ9lXkjZ54BQfxBsodxJvSjOGvQkwFrlUAdhpu1AUaWCp9s+Gv
JL4G4lpCMgdhU4nq/Q8k5dDEjFvnyWwEFmTd70zNZdO1L3tlpzIordDZjhekrYzK
uucRpXniuJWI6rzqWfUc8IZT9ubl+NsKAqGfKM05At5PZHZDWjoxz7J+b2TI6hyR
grFvPdFY+NzXRrzLpnjgX/8dk4nLKfY8S7Ge+eh25cQB6t5D+a4BVaYJHoqj40RG
Dl7ncv8CTQtG9ubpJQGqrhFJzZ0+KHcpNZw3t6+pzpml/tmvVappNSzVZgTUGgze
0DhPsKgcSoGBbmR2MIqb6st9ik+8ZqRsnuBvj5bNwJ5opIKei85AQ58te3uYfYXm
dTBMkrG7dNTwqyf6DhChi29m30wA9pvQ5XAm/ut90Vm9uCO5ZcP9MitR/c/VdoDn
tinUFzv097LLmnKuOl91GIIODHEOzZjZIIRqoxJLIq5ClwT2ATxUFC3s+MEPWmE5
uq/w7aj+t7ldIFkZ9BTWlb3NVorbejLUyhyCPomexnMetHBOSj+XvF6hUsml7imF
deixDrmfihmAWlbse6uPcRi8VD+XYzRpt/gSsNgpJLHatNA+M3nQ+4ZJQvJRMmKz
EO1ThWTMBO0wsVncXDxxz/80crCoavvWN4AH0tvatqt91hkytAZ9je+2oWIwVl71
7q2BFdx5V0ACNTUZlU3HtWXh9uEFUKQ9WeQqDQl8Hc4h07e3veezGPNhGyJEuYH7
zPyiELgrtWSUw11Y3HFYiT5vcRqO/iE/j2OQPYwB4mC2IWmnMS13gvd62/P7m7mC
PNgGCWNUWC/NM+pYOc3z8uLZ0HW3CUB6ij7XId1K4KQrNckKvMWiz7J/G79NGc0I
aKPLz03ceFlPROS/wUo+52ToyIINr8UTcC5kya2J8LzB+bNXJ6SAH2BaXnvaoRdw
YJ7lV3wVH8BE4DlDSxJl2A8dafbM4WVWYMNxd9o8QZxh598zAP+PKfp1f5iFIWNF
YvOiNNPyDPeWB9hf/2MGo32rGIxLAiWJkbawRDHZ4wfUaOZUGOV/lrf5TVkpCn/E
ugudVSayzf41flkRgW3I8n9DF3B4e3NGrUHDHQv9xqbhhd5OX0OrNdVTB79/iiGN
vJ9458w9LnQzBtQlRtFDCs3g/I8BP+QWpg6d0KD/gDC+qDrAND9X7pg+d9/4GwvB
ML1AjWR+PCI2N5mPz3GPH9rC2n5iDPLpBcJ44WuM5QSyBwlk6CQro4iUhOT4mKBT
ZCm+mOxOKV8OSRbt1heTFjllbldwKP3x3VWlYUvvR8WSx9cuFyWWO2ofgB5rSYrC
0hMi0Smr3YPR2tU/zpXiTX0sqp8GR4AA3ZJb7EzEyyzt5lchZbQLjywRoyThb7sD
jU/yokySwqF2lw84vIs432zv9BHQ2XX+WR8dMeRSqAmFQiu0AuS+7bZTfzTSLzDS
HCsJecrn/m/2qWzmB+jjZfq5CuBHxlTul55O3NKW4xkhjf2MEkFkkYiLpc3nuDey
CDLYUuJMvUplH5+n+AMywPioxICM1tmKPFNgevvw3xI+Q+Wggt4VT5D1LAFStmpo
9Z/t6bGW1cLQnCJupw/k7mPRE2FfdxU/4qx5ywyISPz/WWacZvirMB7TGTirsHUs
GBdOI4hYQc4pcoSosDbtQahGcLGnHicg3NASRVdAjISu93rlEONDnXaV1k/si7eH
3o27JW7Kd+8P4WG3kN9G9zQjPzI3UvRkNRfv4gh4MHc0KYnsPMHEJIsfgbt3DR+n
GcmGbb9Xyh4k6f4TYVJIJqd0E3elwvIJYl8W4c7PZxoTZbdCOdbZ4cIY6zHKOU+V
fEjaIowTzO9A5KixG2NZ+zeLKtIjwMif4LzgghUuPDmLkneOin1b4PB4oQZUJ7Wh
dPTfiNfEiFMYShfquCwqkdtKn/Gwgj3IRLjjPKnMFjhFlRzbJFVrljNwPLhqRqCv
rSExJcVs1GJuqpvKer1PK76jRmet2Z3q0Hi4MDGnmSzAMQ2TLWDgyRCCNGCgQi//
wg/GnN578wuggVwTjbZDNJxfPsXpRzqGY4iAQwzAIA/uLMkXnzdseLjAao+VVKkZ
6PlBFHVTyuRv6p/WZMUWyM3nH5pqNgbBdYlhxzWrsZrKjXwQ+1vx0NlFq2e9dCvZ
YQefeynoUuiYL0F0mWcBOWpzxe54FL5Lpr6FZddV1XA9tjc4ieuyF+XFelDV68UV
XRpx2mF4WSP7D0/bsvB0rWe224uw8Fx2Q1dd7rUM9rYuv7kzIlNspJaLjDJonzb6
wmcWLQbWjkc/ELMFaTgv0nn3yicpwsEhNuVrJNySpZesa6z2ILIkAntekUYFCEpg
0q4AbossHsxMOQ6HR3GY6gImTCfKECjx3RMfwkfUYpMX7ETvxg/F6EmnAugVrSJz
vvtgUJRwby5MVibMBFXjYZ6gBNFBtNdT6XYIZiw3DRjInsjAVXMPS3LcUF7QYEL5
ck6WQWMKlzNQs4csN7yrPZizI1c+C/6fFKXwFPYqRGrgTQCKYLzAkLUQoLP6JY5P
Rg8f3j4rBT7Q49ATbOxz9Ubfj8iaBbNkmEM+ZtgPrZ1+LQ38Fk9i3t88KAGp9hEr
hNVrrVsH3HSnSz/nz7RbVLYyHHb6nSOWdkpHDQnmcRD8uSYtJNxMdUnAr1nMyL2p
xZ/d3cf4+MGzf10OPiL0KXxeMIU6EeS9IVu6gFgIN0ofHCJvdrURTuk3Rq32gkVy
A0BHRJJsNclDzdveClnRS+THHV4wzZI/8GzLJsST7puBPNTMGmSGY87I6a7WJ+vR
4J2GR4YO0VKP4XGxWNE9nNgbhqbHWMaPs6Q7ajpD1m4geBUmIWdz+O8So0BBPpLb
cSJq1FrQ17EQZ6NDVoIqBWV/mGPlNjgKDknrNDxEV2WS8X86xOe5/6GDtZGfmpke
zJIsAgKERNlWP40PHcp6F35DoOCDge1Oc8oeCe8DL6366dc2MGCIeVtx5KbX5tvW
vfu9dbNgBU4787Drf/bfPAo3LForQ/+7r6y5LpglAgbgxLqnv/as6INcFiP5Ghys
ywvJGZxAv3jnc3K2chEWOD8+LlLBbPDYURR+yC2h0qq5FBXalCQ9bO4wA/KgtZWz
jMZGemIxajiE8+Hklq+TF1wc6sE2t9XMXwBZBZz2eLn7NMd7XbmVuiI9RLSEiIjP
On76OaMlCkhcBkbI91XXixSYFVbrRa07Kf7A/11Yo17tPfFEiYuubzL0iB9KUl+V
POQqMMrI+VTmVt5acmDAXWQmMQEL0qEu21wqOVaDU3dqq48rSIj0kn27bOH6NYS6
csyGHs5XODfmO0rA7sTODTvBCVybtqU27Bz4jONZV3cDDYHe9YgfNF1STaiOlNsH
+GehxtgV7Wg+zsP+M3xyXh+mu47OQfayZesTLHO4taKhwHdRTSeFBuRN1rCi93Pz
ucwIxKN7YMeTRYp3a3P4qyTV1EfAbYgYaRw0YCc204w1cSjaAFjdxORcnGSzczv4
cqh/+mJwuzA8vEDBNrYn6p2hevkVXyR8Ejh1JDxD+zmDlgFviU2Z+YDYdBWYc5ci
syX8ZTQiys4APDDpEVTzlJQcGtltyqgT8+doexaP+zSamkK9H3TgG7tWmXcnE3cJ
lwRJVlvtoyITamOMSJbXsQNrgDvb1KRq63MSmEHczFsirfx9uUX3glu/iu76GstV
uApYazVSi6U3ll0rm0SdOrxGuTQyYOFFUpEX2b6IMJHWYxr75hiLzO3te6VkParc
5w3PK0lvSjBeYcpcdjFK/YVeTT9Z4mno1o0o2mNFm+niNiSIjTmWacsRa0HCoZ8m
sTqHl0o5VgEPTvnkypoqVbruywlo33za9XUA824R61y9kFxHE1Np3euDjMeQ6UNj
x6Lq23OV5Z0T2faa8v/tf6kT3Il1QCHOzpSvQlRJdUKDaYjSx/+x9N0wEeDHE9CE
9tFhvL75rzQzjLau+1rDUFer1urZGM0hzEn7axaKWEXqj+P8/SELLkkUX0hziVGW
Q67yQMr1TnGbXY0CskcWs/kfKhdK6Qn2Db1pqPfDgZnnxWWIDU5GasNPwgGw93fh
dbIfpfeJ2+n+Xgk72RD3hg3d3p98oagMQ5rISMTAr35IaJmpNOkilhq4hOYWK3wF
xJ85VOgOCDNch+sQ29N9V/78yZW7nW0JB1NTL/SOeOH5hSLpTRKdSdpbf1WcRaSW
igzjEioupRYNZiYeJQgC9TxcO96U0lXr6A8/WK0N96U3WQTiV565pAYj2J879KOL
0LzzfGpXOU5Y9GzkjIv7xJnh4/QpB3+eSG4nq9ZDbxJwEZzRjdqGKNI23quVpfut
bDeMjVpjP5Al7pRaEbHTCa3EPWt1GVS8RYr/KPsU5edQ42dBAeVbEvo2+d/H2sTd
cfb30bGNRylwKPqP1LlGVrD5se6ZnQiBTussQX78i2Wo9mzbgey6RpHzak6UZwS6
oRzrqbQDd0a4gMC45RUVXR3Tg4gw6PfV+0VHLgvrm/LRDynzPkIsqDqa3djeHB5d
iXTxDHJu8QBpzx5Udkq7MqDhFAKtlx+mBO1wxAyZrvpKyiJQlqUOqYN3Gl/cxDej
2bdzV0lANQqIyHiezUHx0MzrSwPPTz2XTMtvuCy//zguRI62kxZAYh8TewdC/sxr
p1H/5fk6dcNdK3GQV+MrtBeNb8vk7IbMykSZQ6AfnmC79mFw87T+FpFbIEnraHCR
GeK93fx+Hel4DgiBfU9wVhESjbKs+xqMvy/h5XnEcnpXc7zEx8DmD+cW4Q+vZR3W
ImzT4r/p4wPPzjrmq7JTyh2xYqn+lhgbQ6jmPFIkz2r8M7snUtPLwe1/32KexIZD
fL173N1PYGXAmPzQma9VmYmPnCGpxmbCKPJ+GoTeyrtzcTYL2uOwRxZnaL1s0xyg
OKn++GQKmmbEALDzjONP/qLC6VdqcRZ1RqsEypxi9+/bmBOSUNrt9EWcu42cszr+
+MvrjZNuiLTnx/M+BXonCFZWShyjuB19hsiADS5HVSY3PJzts0E+y227CKh8N4kx
PG4FRL7uVnwck1o3ZVIUN4RDSPKN3yN6tOsF8x2MQ59Tv8mDzgQ3dyUtv9pcyn3f
k7ytlXuCkL9C0Ij5YxZcVsEG9wlp6FPeG5M0adOPh3p87fTt6lh2l+lTnPQttQme
CBh+otrP0YRTh/PKYqmaNrhPwgDPEE0XsRrFFkMOgAVeQwt1BLIYMSu0318VxiCF
o7NhNvDpDztQcMN7ioYqly/JGkqwDzgilRKcy40Jvu/RM91nNH7JgUcC2jBWRyd/
mdRoFgOjsvcyX3ZTbfO/sAkm3a0JghYzR33qI+QFbT1QgONDVstAGQ12XmHGtr4c
sznDE9Tg1/x7491MxkvCiTu1aNIeNhUPzipm02uIkvqi0smoJgXj2Ve7hxcHPTV7
3NBa3IL8eTrgSYvTlE8wmfiSvUHEd36Tr5xftdj++n/quPY6u/eoPSOeUQ4pxb9W
GSEkqueJ4sQ+bDEzNXoHABXWctn7oiHfY3xc4zLandjo6dxFaIMm0ZkqvTILLw2t
M8OAFf73Dp3oqdNkOnm0jzNYbz9jaYh3/XMZH/ELdKok+Jg8d9W67+phLNUZRoX6
bV0GQ3wEXhcXuZOxxzR6H0aiiA1x6m6dyDbYAWxoDN4zdG0HXJUj9edoqZBn5h29
dWaxLtHmLKQb69Cb+IwfhHCwLXsGqJS5vkb/tCPPkXCVemmV1PSmcPpoZRJei1oB
wG29mVEAjh6kOVBbxl8f3vxXkFwuEEz9dfHG7E+szjC+unlFtFCHdJ8iH7TiHlVA
oSs/NLvEsC/VR3MwSNWXNUD8yczhIYPjFWnPR+GScQahBOUwE5iKaY35/No0BwXP
a7+mKY4eqyiiZQmAFuXbaeVyssTKl1NrT+hVhejaxyTRWRT5qZIisTK9OwCqOCXR
20jcwvgjYKwAHYb3w9uhnJ+wofkzh5YLS2TNOBNnau2K3GWEOEzGHid8Fy5TnnmR
VvknZRVXSHyWw9fVvbZ7fS0OnvbYlOqgRDeu4RjVNCqZ5x83SoUktGkbgKX06Wyv
g7stMhuiK+Rl3uEVH4LQUfg1YrNJUdZjOF0EEOsdb5myfIf8Te4EKVtFvbUYMCX0
OybHbDixciMxxkTzV+IMfD1e2iw5wj2JuJCGqWPYXHfWW59lAbVctW9262Jv9GEm
up5oQQifGCDDboEq+kN2qDog1u8d5ATHkirLgTC3ydbqTcxghVwUO6DQiEGkiwvo
LDfRIkbhrRlGpXOpBsISOt5bAKibgPEkZ7AAWWJ+0KjdXtDKgID5kCf9yMaV0NEx
iCOA7QSgyidhe5AcmL9tGE4PyeABgTPqfYY7M1rjgOoPvai0HvjLjJR+c4CZDv8F
E1NVDPI6ku7UW28WCNRA3YGlddFQm2ZsCmMZ3+OPgWSqOzxA95ru4PN1c8P/XZ2F
Lw5JMM7sKBrygGvQrsEBrLLyBy/QeWmzE4BnKvhJ4gi8SxbMZom5OAid7fZpG8/0
4+opUw2j1STUjmo0SheS0vEV/GhNYt8JaUmLv14Tm9xBeLNQKB9LeUrps/V0S428
QcjV9W2QT+CGihtydTbWrewvPfaI+StI6AbD/AZtAiMJ6zLmh9g6CWeSJaXvH08K
xDji0qXkEvg1U3Pa3rApT517S61uEAwCmbWUJSyD/LuURGRMOoPjJ+vzDVA2CtiC
32Kabq6u4eTmnrvDkn11bz+k8h6c6jkE0wTY30yRcmGYWVlbutuJJWCmHLJKAtfP
/ga1Jrm5O1pcGiTYyBMyLrZZTxCPTVLhdHYwy9IqfLwfpRFSKeKZkMGZrK9KKNU6
pUQfELbJt3F8mHANt9b0/f5Zp0YpdmMYjQVxjrz/HZ3rgBp8692tf4ZVm9KHJ/YZ
beVeqkJ7IN4X2CRCVI2yVtModVBNUWwbQ6FRcSn6njk6p89caQV2Qtr/TnHZVxAx
qgPYR2JFcuycdBXBzcuHaQWYtHu35bzFoR7HhxGsL0mU3ZEFgUC4dglkppYEsj3v
mJqTIUfF4ZebOLaWLDROWaOBaE8ssV/8LOinVqRdfAGcm3GuUIltv7jeGmU+hL0b
QQgKJqCk1IxOsxqH494lYWuaDs9j0e0hp8fxjvIRxjO5s3EnzImj2jH7PwaQp5su
tUw1zkcSZfSQWRQ02FzXw9dCNGcshLRdrH/9w0sCv8m/CDmYZvNDvfLugeA30skV
I+J9YTcvC+cHKK278i8tLmb4tmjIncMome6PFZh6KCoE4okqAJPTXXKWs4Ba3+PM
ORsWij7wTZkIjxuzoAc96V7pE9NHrZdTAB29eeubqV1fCpO2L0zeU7VQgAI0QLCl
7KvzaHkw+GO1oxf36pf5yH1fsCEbmgGRTC6AxfgU+c2COxT9WNGl1f3ErPUHpCph
boa1YN3jNtp9o1g5PNXVLVfZnjE9pChKiOfDU7sa/E+AsqZ4AAL1bzKbWb1psNaw
O9PpKgLyPbYLGwElxrAkR7iRgCX9POSVCJDMi+cTh0c0zoDybiFTSUSmKXocUVxF
dXoXqkauR7nvVXUkK0fqI1LFmcTx6suZf4tRfpmDrzqpObLo2x0zmaOdYgEu30Ar
DVtE6KAcgXmh4FT5xTAAPspXxE7PdVyPZ24DoTdzEKnDQ/U5mg9W5jG+OAa+SamC
bI6yORJ1pRK+P2haoPbO6oOc8aT6cg4TxBVNnq9LweOBtGeQvd1ouODCGXoDu6uI
vltsA+bVxPMYtsmz2WCzRe2VuzA4AGCONiUCIV7lUPQ+wMFCED0iREFnAHsqhfbU
7eGkrpqIxrptOYJh/QesEOC/Pex3hWR2AcQLivWUdGAi9eTXjos027QmqDvAnJ5L
BxLF2HwCb10ysBdjcQZmoNGNrZvMgvfHjvcCj976lsjlTD+lYe0cUifLpSTcoYrX
8UqvlCNfCM6v185T25p4f6lrXd1+fMXK7V42a4QgORKQFAvrAdM6CGdrN5Z+CxfM
tUkFUF2bApTbnBEj7v46dwiQT9is2WjEx2h+d/Rc3sZqbQzXL7axDvFexieU9Lf4
BWIRgDdl4StSSsapVtA9qbVBW4/LGOoNg2Ovbj+IrstDnq7xGUpyNSUlkGv97Y6P
20T6cDJsc9Iprf1nj1tKWNu2ZEKK+5UwbSfkPfsJVRvydB+YdUZ10CP/xe4CRCzA
IEzpgLFyEIrjH1tW4FTwcvoRK9mug3PoGnchUTDjaSoAtgELJ/Qc+wtUFP2+Y8WE
o7l9bEzbE7AxaHgUw0UG+lDdU1shYzTtstHU1EPCdbwqOAykfZg2mocncAIaxOsi
T6KfIeSutFh8z2Smz/ERCmrZrSejogZw+Rcp98GFkWXuOdbusgD8xU5Q3VJwiB4R
+grDy0G1jgMT2AsKrPdqC5ELrqPAUD3yhC6+7f1jnyk9Y7tqYM4OxAE+RZp/5NGy
MsxE+ZBvHp39y8k49KWg/Bd66ZbaYbde9hOzvXDe4pRaVI3yZWTWAeFU5lamKfkw
plLoBaOj5mT/Mu8Lc5eSyOvIMnQNPDi/ocFucy+gW/uSO3iXnkYDPSj1QpFMpWag
YzlFpJnFxsEnEPK9jlopIeErSIB9FZy2R7kuKFHA1Pal8Iw3QpKe2hcpI50aTlTC
Nw7G623nQ+0FV2miCwQywbduZkxTMJbk1XTllDU+WNj/pGG4k4D3FiVmV4igGCVZ
lDgu+V2u1f/PfWLDH6MKPy28E1JSmtY6lqZrxXD+tnnbd2X/aas6vQa/VSFAMo93
ZedlMMlYzrTjfQtlGoPwZTboG3qoWC8YHLKQTuACccOHkzKMX5DyU1DYVM7QAeuK
pRCWpmyEIQ58xP8sIjpGTLlX+qiIFRwCVHWfKdfWqLWvQXrersortKYF/II48uuP
pBEkH4o3Oi2+paANmxcRWn5vaNPpUIDln7/3GCiILDxq9wN3cCP+g7/YjZpRQskB
cnVBiLjKcoNHed/MZga7iqFq3emRYNdjtvTvBRINBN/PNKekkyu1f7teLYgpK7ye
/pMJjRfXMap4mfEBHjF19rpxwz+cGE7aqHgpSlPC7rO/rRcWP1lA/1S+4nzLtGIu
5SvhPs86QTkP/Bx5qnCq4tk8sZ8/qKZJ5uYsoTkUAPDqxQUT2OlSxwrOrmt0lnF3
rB6lV61vzpg/Ttp+I2d5JuoUg3diOOiVO/wQzuzj7xSqWgFat4LiAi1E4pRTdTVQ
d04xkVnDaQj6MkWvPVUlo2yJdAFskZ0K0KsdTx980BNn9QwN/IjWWpKpm2qljcsb
fuUubsYxopaHUYrtzuNpzLxlnz/7RARPS1zqlAlvzggr99lXPLZa5eccthJ+Yh5I
N3yKHZckVTOhWN3QE2SBEd9zhrHdP6yJi98MnIw0G6IH+TNN8hsBt3vvNlvugCkx
WOnPrj8zB5uFGj5/n7xGXN788T7f9jj00N5gupsKFHpeZ/UwhnLvlnyduG+XT6if
pEWwJNqgtiuCtOWuQq3SNU5PH50HYoI5iDir7nogHUIgQkxn0DMTZQog0FpeCnN9
gqQSDoRe9hIzHTPbr+n/gqk3isp0M7E2ul6OHGLOAlInVj5s667wRLhNwREh4e++
Uphrjig72gAPAEzeeJti47/7VCQwLNKYYCn2O/bR4dLHxXhmc+SzBPVE/2dPS4UA
utebCouvpcctZoVUfPBf5DnVjzzjJrBV9zxeqSsjr+NpypFRQ8A7oDTkmPfeh/pZ
c51XnJL2ftsZ0AvRyXrMEC9dA5OWP1wE/Ja14oDvw9S9Uj/o2jdGi/Lb+M74fDtz
4ho/TCuk9CYa0yR6mLLu+/QLNeGkRR3AtDHp1RigBnFFLdrNl5q3zmedV1LoyluM
jAX+Vukwycw3qk7tN5SLb/pfnuMQ8gqMavqKM/hsG99KX8GvQJxa2eiJrNTBdlFt
+k11HNyosfpD4TnwKxkDSC8E1zei/gDg7I0fa7Y1kCIk8qU7/T+J91/Z80hryIL/
xO7TfH6O1O2TdVkzxLdW8FzU5i0Eg5tHkFfDm9jLxdRPzrVAryqktCe354z+toIE
eH5DZZtmkmkSNfvapSftxr9eDCkFf/hWDV1XpkDqOJpITE7/Gkm5Uv79OUqtB3Ri
Sk66Pf7j/QvFncO+H85mK8o10S290We0TqaO+7zAvaAdoWutVbYeT08UXNrfotC/
rntmO6lNmrVJK0ROcD/2wndrEQDgsWndRWgVaXRjaaJZIwrFBLweq+dad6TLCkoG
GTQ15iB090Lzhnp7YczcJ1J0AUQgvlNZ69k8f2Th6Zbq3sGleAm+LFc8T+CG7V6a
Xn3y8mHWR6g6NJ+luocz2glvit7ffsAww2N2gqFAUgp3jkEd8xRmX/sIAn64dDkB
92JStLKC2vLRPkWiVxyfp24BmqqS2NygoyH9UVwHchOHa7nUEei/rFdUfJub20/3
mUwAIGZ+T4Ln4WxcuPn1PfCZYwkok8ECYgPEKw3H3Lw6hAwRmhJPhnK0kZJE7RVW
pWiTr2fyG0aX1YqPNpFdRO6vPvOOeozUjAP98Zgg8T3kcP24/uxGRpBxxVOY9OJh
fBY3CNeDtObdEbxwKl6pn9lrV/F52I3A66rKJ9A/u93crdEl9DRgXhrgRtr1Hvui
LccXEwJcW12EtwDNTbMZFTc2Z+DDuPd3M1SgFsUXq8rytpo8omy+2lyyJEZvCm1E
1VchZwz8zzEBZ6FHmPWaEISg1k16rGibAs/Qkt+jb4nOHA1B10j8kFrXftY0c1qv
Ib/S+4fWfYSQ1E0R0ZQs/TZ4iln8VkappkbTZXfK/bTvl2ed0qi9CdH+JrCvNL/x
LJL0GLkv36PJEjL/xHnfILKCLOeQ4vHsnGA2D59Lamwj7Vr7WLZZeYzGC2EV45FY
Is6r/jEoPk+LqL2TvcAOVEvodfYTNAZ0TXF5y7yvn1DcT3UGh6PN40Y7r72qDHGQ
jJcrPDP60eKFXH2nTK5l21NCchMHxkXxztJ8otmgNzgItQccr2hJqHesQ6QjUi9/
ZR9NcVahLuy3lcUSvi6NWHcXx4Tuk0wvWuzpuuwYt0vExlg2M+Ueg5Md6AHrhnzM
1QTBSrTnFfmgDe4dd6E5sul8aBXgo0vLscLR3cBPjq/3Ttv/tiBsN0yJ+8yLW+bT
QwfcpBYU9Neq8il6JT8ba2Tk6bgFrdnS0bhBX4UDnVaQSaPGRNcYbA68Pt0uanc/
B0lfAZfA/XOnhCF5nnxio3L2RpKAr3OnNvnEX0S1L0QfRAFOULmGXTAkTnjG+G1l
fqv5IRZu03BNMJQK0jPtEwe3iNfg/803qNhMdmKwslbCMGj6y+QxXVXYCNhPyWbE
jLwEwE8T3DCiUlxCfvyUyxmEgxJZsNuTLiLEixSXKLD9aBKFPjaT2Sm/sg1M6uWE
Tz/yfUoR55e4HXV2r/twTzG3jV1ZSGqbKrgG7r03Gck6xPRidMsdSffSt3nlm28g
ndCb4q6/vHBX02yZmZbYHWWEGKnvV79Wk4+dTzRbwFczXabJQMCC3T/rPCQnidbP
1TTmipIR1Y7sybxnSuht9/qNRYOzfTwqceyRhUBlauQyJUt5Y+rCpWeMJk9Y9hW8
4KYQO0JyIgffeNwOjUeXIa3XKz6vwTIKZnDYA7Gzdq8zrIVWjpUZENo61R9vxji7
pqU6cLjCpDeXKItwDalmYCmx9eiboHV6RM4l5ZjmApx++5xm72SBGr+HlGsss4ft
BJl+f5ova8k2nXNiIZUm62YMn7UKNnsxzqQFvA/SScQppUpHJeBMxE0gdDAVOEvu
K3qhO33EukTWuKakB38WZoK7UHbYXj1hfKBeNl6eAyHEtfwpR94qlgD3mcL607K0
1QjBkDQaNzNRDB813gvuJu5v4jgRHbUdxRwx9x+9EaY/tyw2c1oDjO+muKfvJcW3
ZtqTh/47LF47JC+VRlN1l2c01g7DgmtmOrWVRvyzN7h8FV8UgEkcEwUSqgfTH5Dn
1lUaFbq3huOteFviCaJmAdk7pke029+6bL/aTycnROkT4UzxygQUZAVfxx7lv2YE
lfmXxazCx+kwz5ZZrz1C8ZU4Wyte/tadUagsCgh7o4GLAMkQ1jYcmOSphiXUynum
nCTFEkxMlviFQFzAwqXdRtmTrZpOyYGmEYeVdxzQaiOZ1q7by6LTY07O2GrvNV/8
fA137QCvsvhWumaD2HY4B+AenSPCbx1+Qt+jWKpF6hnUuNE7mtNC7pbKj9QwY9On
liuK+mi540FS7DaFQYc1D/oC48Ue4iRbyqXJ2Ggg+sNb9fWpXWau3wfpMojWj+Xo
fGUuHXmfZHGIGQJqB2EFm4R/XFQRZQu6shBbJCeJBxFGphxSz1H83AIKJQSOquIh
rHZ4g8j1xSLVCk95TXLyuU2zNt8kWxQuW5yMDLAT2O9sLEUOrLZfc3n9UqlGiEX6
Nw8ye0/Np31cnXexraAF8L5pSSYHCeGOulHuqaBdRiu6qo7SRM/2wsOfze7NEi+R
QnUghXYZVRXfrIqAFs5/8rr1DWD2BuI5ySJkSfBS0CgmRz3vJt60kUs/bImaFids
r/gkN5yFm5734tUElbHTy9/arf4yinmugRBZX8gZakMrtpvaShjVdXWSRormD4Ca
r1V4DCor2VvUdtO3XGxEoYvod1SvhdYaOZpBb4KW2wiUO0+sHH/f58pLXaUpowRh
9K93JJ9CDIEk8N7/U6Vzzcxvz2lKGOTQVASGD/1CfxZRiEeLlxV1sOGJNb/pTMYV
Sp4U3eQRsfl3sGJcVhGo8+h0s+jxxhpApBPZJghDSJGkL7MmNd8Z4yUAxB4YhHLo
pF4FdLBQaTC9cI1gKCeTkJ3VsDNCQsVmPOR6IT4vHLJ+oGU8TYuLzj5Mxeo7+u3m
htH15FWazvnDYyoSzRHwYJv92JVGix/Rt2rFcwwVCSwqOMPs7kjl5vabiUSlpMaD
TWtyam3ai8fWcktg4OYtp19s4gNPLtIgZft3PFMGJ5cSSrpD4uJFVCnu9XhkPxY0
Mxw918WfaEjqA1F2P/Z7f8qo3XkVWvl+Nj0NHNed2h3kX0Nl0R22K9a7Kp8qKYIa
pyYe+w+EkuMuSKExQIyncJfMhw3gIjTj5aqEbQPXpCD01okLVhnRtSRdEP5rEhP6
4qtJY7ApqpcdybFIeL4X9cX371pbpxRUPCgYxI0qy1YIngoL0mJ4mvvRyPPR5S27
eRmTyAbtlxpxhGi8vZoepzwjKWAQtFGimaHsI9zCq5cuaTYtQlOnLrvJFOn4ujXD
uquQQDZqzBPArALOmC6WJ500Z27APLLGOQWmGy+LfFgpYukCPyNjlI5QRwHplcnq
vN4xYKVzfxjEgE9gk/YGv0jKc1xBYR/rfEMrVGZsJIl52qIb1bhmyU0zGRYpe+zu
5G1f0VxCmXejq3C8vzeh6KDW3X4sFvAmTtK71mcxgAhv4zuctomKuZilXQhRlYVA
FMbS0+5Q/Rrdd2zaeHgRoDpvyAK+Odc3xVRPaoTbvFZTScpWO3H7ppMUaNS0nGXz
v9vWHHcjRocGryo6dZ97KMDcHCyzDlnUM2A3FKrJk/kbKAdba/LUtaJMuuZtxnBq
F0RYyJeNVyAb2sp/+dZoVrW0kFR+cJ6Jn09sZT0+WZMGUkkwtCU7h3MtOwb6Nx33
sj2fvqIkqfp8wK6J9fYLP7c4QDDCEZYhnIRrsqcAxx/8/DmF0KvhxnSOWwaT7SAe
EUpTbvU47pSBLxdDpOCEE6Wa5H3bIwqJFkIJzVaUo/bfqQiKBJV5mSY5vLNTaBnf
BztxVvnAWjsV6T7vyfvxpm8q2Yoq8iyvmdf2feUPispsjk7cb8lWyruUowNO83SQ
0WOT/og/pVTD5t781piLdT9PjGg1ya+0z2EaAyUP6lPy9vh5dRGlPH7f8QQbGBan
bXiVILGLyBNeybdLtlWWCIJ6z7kNl0WQKzdJzsgYkoM06YILeh4CBZUHlb0Q+INF
P/Q/5WDZXjUAfsWVPH6qV78GcuR3uynMQOBUphHntbTIUu1du0zP4rAeGc1tOoiF
VY2YfcsYn7CoYR3WCz5cNuS7DRfba087DnmuxqM2ERTYbdSLmTFa0Zodvyf0Zw/n
yX0xnnzmB1QSgXcO2zAyo9jKbEB1eeZaurlANHLMM6C+FRTDFn2qRp0tYLPfsyYy
unY/+FTmmQscTmPwNWMp001KzlBHVSlyxDRm0qxn8GtXy1RfrdAEUcangUx6fBZ/
Ublr4cmgqxUumDkRS0tUoRrQpgRJfQ2ih6y6xSTLRUAghExNd0BDnCXNcdozl83/
SxpL7O4GbLuFW8rauvxAGmidj60yS8+xpJ/CjCV2BwA+5+Mjv8z6fMGIRXfa5k3F
PhIMJjRUghM4NKHDv7s41DLZ0nPCeCAZp4Kw/KEFK3Qpf6+XCRoCDjCYjnmWJCAU
P0sCDvavH+tl8TPLO+xIh2febYDhatef3ZyDhUN3/M7HgdJbMK4pIYDsOxKjNMLV
f79wVcReNlGoBLUq+rc5WJ4iXHkcu/D4qed+iSmlj6MD9TJtxq+Xa1AI4s+6lwyy
0t1NX4CODe3J1bEb1po/gA6RTA5HifG4MYEZ/DchmHBkciZPW1OfZxhP2aywisxr
Oc/ykER9Y2/rRSUNnFDnKYfdlS9Ti8nccWn/JQ6faFNzna2/yR+So3v+09ckL9aL
U6wYSF8TNXyxllgBfDEgKjWR2Y5BseEOIUE8k8H+m+f408AnFgoAAEUDiQWEURPk
dT4UfSEVgKAbI/ynThbFv1WHO33S8WsuG4FtAdbWsdeC/BjLrR4wCl80ixeHBS0W
OHPYsXm4CzhKdZKjjxwHQBWul110hvuVCQj170ki0nAYLUYCFasVE1Dyg91gh2CZ
ZGTqPfMsBACxVjDsrX790sFaJBZA1pf3WEWWlWdOur7hvY7TLIqYnfiX9rLtFil3
MPjIIyPQGalClwJO/AScues9geJ7ttZKL+g/XgBSFv8XbrxpRB6iIg1Y4KL1KaFK
e91WGW0mnPu2EjgS1OiE6sp0RzDIrmdm0WEelGTpOTuwJjVdrfb37lWjqcbH1LXk
Jn23vA1jkAjY8Q8rWYGuCYy41m+mV6JG7lO2mgCrGELHJg1ovYoT+9ySrA2HzwJY
t7hxJ1xOViFOGm2UF3f4JIYXDzM+O8yMBMVAA9rv7flUKrrPOFA+uOp6hQjs2yw3
2m2CSujWKYatGzBMBf9UhzaSNODb4HRyUKhA9fSnYgvwIgRRo59lMEceSXthAAQc
oSzFiiZyYUA6Ky1S0/OjKLttBb4KC7W2PXQFfoXunzSv8FthGaRjiDEVpqym2/cI
lHoHssXxjoQ1pv2KVuSSMZp0QCie6hotwM2Ne3K+jz8EWwH7YIGAkmN2hLy1qpJ7
pmPK3qrNT7sc3UO4qdK52lH2kUK1phA71F/vAtYRKtxuKYGgYdHDxxAFrq80pdZF
tAOMivQIT/xEoAf3OJ3xl3MOMF5Ln3ezoqjGulUsW2kxZ7T6oqvcjfHoDxHQd7eS
gyFUMUDwVen+9KzRiblHSyGS2yS2bpTZqAC3hWrVhYq0GBYjre4R6F/fFe20mfuU
PMvhYwoffVn+5lIqNdriQDg7iA5QZPIZyxW3M+wGHBHcsTT0RVDmB5K8WzEzzAC6
L1pNbvKe5d+JH2JZUt+rep/nTjznPQHRE//SDzXA4fGfew4ItADFOC/FJPAfegMt
fA26h1QgkocsSVtlCEI0DXMnEQvm2jZOML1muZOi4xaaMZHHafp914KwYf4m0UpF
3386MU50yfas0JIJL3WyzusyY0mw4QEoAQL2pWXrEtBwy8CRLDrIOXKtswSLO9lZ
vjTqBqDN7Valnv0ieDDHR9yWGNNiV2JuSehfrViv2sc8JP2OVM7gA3qBsaH3xbP0
k2BdZqN/iDf/VgI+cMSHVyRR2g+jJpgsLJXtNQReHrSi/oEz289v/uJ8lvsMUrWy
u1jtBD8I/TNRch9ZaFiWEXreQL4NG1zuG42l/poXTGWdBDvkppGlRrFGG3j5CjTy
fK98NuPEJYYcW1lwM0C7o7qFerZ4cfpZ8rHswW++E7lXKnFBxyCeXUqlnanBSV7s
Xin3CgUW9f5IFEJES60NLM6hIzJs0EAO+Ig0oIr2bZXtcTpsSOhWS/qKQcDAetP4
tlFYzjoOdDL3yAtRV5S9Mn2bug9yzFYM0vTrBiZ3J88JaUx/RCJKWYCHPbcJli4/
OjDaNI6AZC2mvHb8ZECZNNydlO1HE+M7fY2D+kgasdiG+fo18bV9EwWwKtD0x+6/
laRKZUT7c1I5F6MsNI299yFQGwWt685QP0KOa+ZP2Adt4Y/ZvkqTavzbOKdgP9FA
YQmxS5we22FP+172aNJ7eFuLCQrhhj0FzRJY4H+XPSwXvLgmrtc5O2ns2JBOZzEx
6JuPBKRCBFUpgz7bxSrouWMtwg8EzlWdGdOFEGpNXI7rZb/utFqqRwi9XhrG0j61
g4rT34NeIvBEkWXrmVZPxP69ixO+FZnCvnS3hxGsfEESZAh3b1POHN8f9X8AhUY2
ycAUC6p588LX1jxHPLZbFjbRptVw6+5deC5tWP8+BvtwAjGc2ikRuGqXqdBdzTKp
LPrKe2P5v/WQ368YUmJ1IfNrAk1XjeRv3NjGXIoqu9fpuEHDEe0CVAJAVGsUpefG
u4v6Ii6dG7Gv7EZ9RPH1aM2+0cjYrPwosrFoeSepbff+SsdOzfaPixQgSK/yA7iN
4hWDieRrAMJLAowqKDj2V0+pmrtFVjljQJYoyzdDAl0WlQJD9h+xTknhc9+GGagt
MBmjKa/1uOrewD7owlouVrsd2oRjPiyEWuKS4frbSNeCH2GJcfNUQZBxJKazFr5t
YYEPyuYbOkBYgFurp4UL961txX8Xz55FEwrLWLMmQRmdUNU0UhB9kqM2ZiJBA3t0
AvLdfEuSkqWgYw+pu0yfGL/fCgnBc0kve0vF5XSPllU9YnDbHulyGWSVwTAkTUyY
khXgTaQVX/OW9fa2a80EODpj7IPyJysY7Qn/wSajX3Gwdcno7tnMMKPTLhgFLREz
fn/F1NswDYsm4HBbh5QRw9boIb4eFsDq4MPRuubwl5WvXkvGfQodGbl0ULiMRTw6
WeE8Tk4CHBnIW7tN2nO61DG7DgsrO5WhDPEeovpt76bY7CyWFUryfR7ir3LH+f1P
XoFajEq8zi7XFqELUtPxUqRVu8piV5LXVI2SdjPR/I9RX9olW3gWfueYK4wtO4cp
eMVaUQaBW17/tyjc4AwZuYjBoYXc29t67PX3MHp8NaMnVkyrzVAnksqa39gAsh5s
oNImCtRXalx+s8Pi7RcdmlDstX5mWffdK+3VcDj7DC6ie+kh7YcyGTFRs/B9O8Wu
b4b9ZPvow4KLoNGosT3iNMAGmWUx6inv725CD9BzDIisQMJxTp24vQ6I1pv3FyAz
RmflJoxCNC0T8Nb8ApaHkJWiGPR84HnUiiLDBKa+clsLJPqdvwVCDynwU5M8+lV5
YkZn+V2d/gLRBgIuW/g2r0DE4CjNkV0Y2NEcAkB/ZBrNqT8QtCjFepju/lF08PRk
9Dd1ES7lwkgJdcdL4A1MdPnqN/lrEOCt4rGq0Y1XfXw7a2leH203mRF3nMjnfH2Q
yALl+7lQxDqZJIGRbm6As+iN8Gs2r7XqYHofv4UJxMYLJmOf/YI8TPdEWG8U+Rje
3BB5Zbe7fT6RfRJyYQd2X3hiaecjDYigqTcNj0PcfJubU/znGDvOTPxzArizC9tT
1fWPlO01xLRppqK8elkz6Uh0vE3YZWcScaKi7pd4hVOcaia+EZ6JoJUG54Lys2V1
MCFVfmrmFsKTF/xg1v0J9apllS8knVuRBRXwtaE4FO0kpUIX85k4v8orzIVYJHAt
q52Rh2WC1CQGjDcdpi1tWgxAJ5lvskPItFLAl6Wm9ppIYEpv71rB74MZ9XzG3HcO
WtkSVTGGccKVdAEy91dRI24O6gEW54mCQkMH1DFQRvVOgX+VrPonHEY4FYU9CNMc
Rrz0hvKblVzrerHMCRSFWs6K37IBgywFDY++baeEverfJBAC3FMdGi7TLQpMhN9B
krpZht/j0P//axONAv9pt0nKSltj6oOXBfOH8t4oVNH4umJInf1LSHrTNWpzExiC
V+wogSBYxlQ7J1tCfFca+dyAmbvlUMVJzbgDbV+dA8aMpuIXsCCYLC8LonARVfnw
dS/DUiKsNA+7vCqDa81z4UIs2dPV72jUwtunvfK8hXM+XaxSUTxCm7f6pJSSboax
gWfGu+XfThMvs3/4xAlucrR0lFjYWI4rksP69S/8/ZwrHhqSHa1ZdFkIZiRvB2la
h0S1Se73Bl2fJroL4h69gdKXB8hec8Ot8DGZ3G57KDZaH7NnQAiXws7wWHGMxE4L
dRVrwFqGksonLNL0WB1DH+yhwpjF5M03s/B6gNgGOGWl8IK5htkCzHhXpfLzqJD4
e4v1JpcvaFlW5ON/cqPS3gQAPJrA5GC0RAvLIRFgWXO4KQjdjxwJDeK7HkD/jXjw
okZAI+u4JrzlSV4FK2ZDMRmDRKETxwtW5eiP4qh/jmvFexuoDNDqIqSdBPnrURuc
XfNF5kR1ho2XmjXzrwTLFgzZL0eZIjeiYW9tCUGqmbS43rlSaR5Ekd5ySnvVT2aM
EMTBQs04/RRwMURvCmaB0c/s/dAeFYmkJZEUG6cIq8xbrv4Slq2S1rKmMUIPJe52
PpQ89lDBEVIjk637+He+xHti6ovEdAYjkSKMcvJq9qLsvSSuZ0FmWM2zeuMJsF1s
H1xFge5wEO+D9HfsaurKwkDrIYhQapQqgCRMrJ7s1VZ2fX3aGO9G3GEYvxKazZ8k
s5kCfHsEXwShbdT8ENbhC9EVNFacOPfBqKnTekhUHW33xZIy8d9Fd7khm45L8KJl
EYvm02PCuQqcDtbkPNaHLVN5r7cm7lipSG5s6FpK1vzHmpVXveGxzrn56bRPiB5d
H7myCiy7V98T/9LB1mN405LoyJ4wsfqfSidW3wuBBk6xBFgyhYf17guppiCM/+QA
SQQ2VvpUNSYoaQ8KB3NEZKv3xJ3Z0wSVZG0a7R0vKR6SiS8B5XhFZUpFS4n3fbEI
fm/T2qe0Bjy3GyWkc1sFsPQoGxjx7Ot0rbqqr90/Gr6YbhASsVYBPor2y48pkPGE
/Qfo0KKTJhr/7dpyDl5z++5HZUGeLxx7sbdWRRvQJik+TglChf3d1/zV229Qf8j6
85cg9Nz+jY97j9Rw/53xfaUxZvPnXcaF/Nz5C/x/tG0PaYmdX1sga3F7O2wKBK3f
J4krqyy5v959G/whBURJrnGtcYFGT4M1/vW1l/4Y5Q39EkFqMnK03PioF1aVKfDy
zIAmOV2ius3oxoiR9fOQ5uzVuWj/mA2jRM3/QZGfSErNhdHe3E8OlkOjoq6fGCXH
/gNrKnTKjctsIMYjwRrhfanJECEuU9oXaUaX/9IZ10V+vjQWwD7fRIvn4TanfT8G
ZT4M5rajaeIzqmWfa+0d6LCBU3dKmxEe9nUw6/SAl+DBMgSy/b9fAhBSQn10x72v
RtvfO4qs9MkkUS29wFN0jKZ+QUgk5HRki704S3RzrS74b4n75Vrfzv8uqEMF1q08
QuD4JOzSDdJc3TFbe4jGDpBHGpKcYvFSE8mLBT8aLivMN/Aoxz4TPsgamjW6vcYI
a2d2X/N4tXjTB4PGv8dWr6m++Q7xKqiJI32a2uLs+rh8uMpKb2uWP7zwGS3EQVJx
7l4iyrhnF6o/tKFeetZLh0M/0BvpmsBf9OnaiaLc30rEj1vs3KfwlK8xVDdZwr7s
pr3dWvqAy/FNfpsyj7VQl/JUDhC8l0czgNTYXbTqm4He5/dsoasZtgjmLcPD4hrZ
RFazOjirlNeOOABWpXyA1adeAUI46vymsPYeZ71v28+X5lW1FqoOI/2PsBU3xhKb
stng7NB4qEY9jiY7e2EjLiqRGjWfjeoLL2FccaKiurI1QKeTk8/n4KKRQGnS4cxD
yq2Of/a8kjoycr/xs020i31yYlDp745+CsbxeeMlzoNpn8V6NuSXFztT05Xe9bY3
I1ictxV5oBTWjtIGJg0uarZpZWH+UoIIAylvmTyCUaSUjCWxMKTdoyQG9sFpI7Pr
ydFfJsKa0OqcxYjUICGxZEgNzJ/KAKtb7xvogiPpWvI0/kS9F0jKq+nEG8vt97TA
e4qewzUkFI34zgNl2FygUX7Iy+fo5FdK3uM7Q+sDxQ5CcHEt6Ezz+E6x/96XJJov
zqcU3On5IbYZc1toqdjC7YGRIPz9Af68sxRhkZ30PQgn0Q41W5i74XITcRo0jaSP
LOR+WFguSx7YZNWZadQ/FNkixyM0DEmmj8PtfcYcgoWPLg0lBhlMzXhp8rknyy4p
JPNW3hjicfHNWzZz7GQcSrfSThL/FyzDDVOgjv/EyPvHNxQdedjWjfgUI0WOMqdI
2Gz6LRa4ZxetnRj0Cm65BhW2ITg2yhVQZ5xagGc8ay3chzqExxUad3hh1B5u/bg9
ongDrSHaqcx3stpxaP43pPyfg7SSWIhKc6kEJzIrngXKIvvhW9Wm7qS+IB05LPuc
NOPJm44YqIxAlLyIYo04p+eEQgPFnqLLEfOy1H0ueUlH3TAeW3JJ+JSKXRUXxgLl
ppa50XCSJThK+QbKxdV9UkVrmFEIaSoQkn35JB5VXGo144qLdDGmCpUITHOgy1KQ
L9mCjfwJwD2dM/ky7OqSJvtjItqZ0XtztAIgjdUsxpiHLQpY99NOu+UhA1RUUuLQ
Uji5YixZ1yS/XA9/7wXL16Kf0kevkL+WtdJngZMaBKQ1vF0v8JHXBFVpiMexzAHn
pWtnpm4+leOklXMOZm3dzyj7q/ySFIfup+Axl5Ja6L6HVyaiqXlykfO6QGlUoO0d
gLB+TR0xHGlhZxv22/MDrnLWQbXaDQRalFbDvqvfBxvuTPb9jCXaC/5SB64ZC61k
XjxmHReHsbT5XD9JgFJQmA3WeWMMs8s3h0s1aeko+5u3EOb+pqAEYBcdUyiCO6Lu
YCif6a5mRokUL7WtZP+lOlODGgYysIWJA1Nedml3aNVp4wREigJb4w49Gts//IRp
TQ3txf+oL6r6c4fbk7HLT7Xt7gPrPEsxvrqrIKMgTNkxiRGk83ecH+0xUIiDZPGP
va9s8BcER6uxEarwmIpCqi4Jgtv1uXpQcOUuVqyXc6Zfm5JQa2bMYXsKiBG8eo2U
41ViwdKpWE+Y0uPr8DCzCeGpnQICjF3TpHHlrI6cgfa4+nvA0M089G2Gh0XaK67e
6pPAMxsZwp7ORgezZOlWMg3nAjhJ9z+mUvQZ0/mblLQgi2vCI3e8ScSWpDKo/NIb
xX7hY5GowvsBw67JEsUgK8iwIurNhlnNFvPDfidy92w3z+EDfPwVx2Vv1iFQCjLP
JVUHy0ocdS3QqaSJuibton148HxOz/pizVPLleo29v+lSukBianM3r6Z51x34G55
NilZVQ+KiAXu7MzkIixWSccbIpevZu4iIC5Tceen0T87HccoYmzQ0H5vE/xHWFyA
xTi+FNRswiJGPAmeFdp2PP7BC3Uuh/E4bnO3O2JuANWIazFnlXTRUl/gEk1GsjMP
BrHT8iSRMEqGQYSTMKXIXpmdn40pLYaWpWjCYkNEl9UJFolH9JPno8uVHACWArxO
v0psJ7UW/c5RHQbcew20yr/TRo6oEEaH7YjHXynD0ymF+7M0zgRxzNjCLJAC4E13
yPH1FHXJjqgWH1cgEv6Nuya0vhh2gEfb8fpNaSoPh56VusmZxfRZ7ttBcw7RBKFN
Y9TS/TUz9jsqfiG/kSt5ym+rgyNLQaH+WrUwbLaN3bLpNFvqaLpMaubU1QkNK1TV
q5UmEYDo4Y6HidsMW3rLr0T+hynXIn6xcthu2rKeTWxlP237vZufx6NGrNGqKXzf
CAWSjDj9HFWTGNCaKbCFtnTBtcbA7SLmUhDaHDrThJu/3TjLnpLuONzpNOFMCMVu
nS2xkB+SItQzGT/0v5726CSy9zDnJtz5qPb+yPtpVIxUqPnn1F7S50hmcKm6x6tj
u7eh1GrpYXDQtPgK1WO79M3B8p0ODkqilPtHCmQCz2Zm3BMNpVJh5xXFTz9gwri4
IJe58thfQ2Y3qnJY36C2W2LPqlvvwpfeJmVQDSWnNgQqobwbfKPfENJyFtwG0G+y
5mJzwhhGpTaKv/d09md6/TcC8fDh63jtT7PWopHLbwGmIArhOyTJ5F1yJf/8mob+
SVIdFOIRvvwQzGvQzTiuJS0tss9eKOoUOGinHKt54+9lKHe1PqHFHw3QT4vJY/sr
TKPR5UXw3gDf3bgui6p5yHLYFPNDtjCym+qj+ErBIRNxzVsbtXpPaei6Ki0wOcqi
dXUNWU0FQvVz/sKVhP2lv4cr1BwHhtbPCo0ZuaYoUfUXZDmH0ymkf/H7jmNzhE7R
/OjC4l7Rz7D/pe91OJqlvznY4RM+7LG1LAyTyxLcrGW0rWOwUQgzzVPIwEQ5VmnT
jQPvrWsqo5qGOjOMUbnh7j3hJBE5TYi3t9gknGZam6Nw93l8HrHqoXj34RoKv+ri
Z3K5Yj+9Ct1VismB17A8ACj2VIR29D23niEiCc0hLxUytFixs7xC5HGY2Lro+yRL
GBn1vDj2n3fq1vgupjVUBflNswPscSrfm6oiwdUWFdjJ2bnTQrTROzMEmp74DYBr
XeHnnHwuRZZM3E21OKq1VI4Lybj1C+InVby+Wd2Mxv4koyCK2zOW4C3LV0lYoc7e
OTGePIDQogiM9E+am3h/PihzZ0B1sxuvKisBTsD0FITEBT8MEbjF05I/DAqIsCYP
MC9Fn0glvXQOhz3V/oXUKVaGLSW1pyBRkSk9N19C3qfbXnKWBo2/rnjw0qjKuvZQ
7rpJ0Se83RFOxVcmXdu/nIT3uyXjZFl+acA0FdVQjSZ2r3kePKExfeg0YEF5nKUk
G6IMBfm333m/Y4OBJXreLT5HG8oCc6vQzNE0/YdhJ/pVkV+UgUkoMy+AfSkEYmTa
jo+jj3QCHYAoTQ4u8suSCJCeaaXW2urlFhO01eqJRB9y7L3OoFJRGrnRQhTqrtlN
ouLg7r3iCppL4g11jvG+8xMjhfJN7GVaulfzOQbhhXZSVCqOpYUpxhFRSMOrA2J2
j8saI5QX4LdKNzZ4mAaiaG0+uo/KTZdUu7832WjjB5LtF9LBZlXvEpH0g2zzQDYx
QUm7Ytim9bzn2pmaeAbq1uGcorphuELcnmSdf0Sdt6jNfo2TdWZpJ+MeEjtKguls
8s7HxgKtUiyZjJhJHyPcqhHeJ6JFVYo1ul09pTv+vHOjkMcfD4F4Xyy6X90BoPh7
A0ImCpIPUppkqaPBJDqcOx97cR9B7Q9CYSWLDDZbHXAXJyRv2gLfEcz5/bq3bbBs
v8i+7OsHES6i4pzhVWAWw46X8WG/nSxDGFpl121eqidZnSvNsQvYqMYAumTYRvIA
8uj8Z7wthaiyDHl2KpGJKmovYmUaXkLQVXtEGHngip5ahCrbZpsCd0RnehlGS5Gu
MQGA3P0M1Dc/mHBN6srYruLwpmKPOWs9r2pdKi9HdHOz/pxFH80MFtKYQstvSa60
Y0t9hlV4vI6NWpeZ+7YgYUf8dBaLUgCi623j8g3+fiS1d9TloUhEXUm7kB0CrUZI
4eKA9sVaELgkRjulOE2u2y3lP01pyZQurmaKrCp8KnP0CseSnGdc3TskDF5y99xY
V6jxGzsBSabZHyD/g3hvMhfgmI4mgux2PLNVmCUhWBqShybch3sRwVD95i3sa0tu
WNTxNvHhlQbvzpwdTFlDSOnts+ffv/uyS1/2Y0NvGAO1+RoXIVZ4zMsw5yV6zr3C
IgrTUmZ3zXNeMmWEVvTNOA5YJdPHLIBRB3353Ws344m5ZUZ/51hXnnz2iGX7qBb7
yeQs8PZp4+ccG/ThaKITFnAoIFYrhVMayAH3unAUCt+RCfL4rdtu9u+VgZq5h8U3
RT2XFMa0c6T5sCx9JfEoX7Yeyc0KvOoV1V2ocZEEc5eOVkM2jf0WF3yUp5rhaN1O
7yjWmCRgTxRxayTXUnvFmnR2hx+UTIZKoiZ2rLy8L5REim9XI66gK4RRMGarOR//
9DeMwWJRhbYPOxuEAGhhvYVvdvo7mhOUzmX9dQaXbhCs6j5qstaep7WKymz9KcuR
RQS2gS5hp3xRIRk9AzJp1sS0sDJdmWlJpcDbw4WE9ka5M8QmF/JeyO5k9co1B5ly
4A3f0pTKtgpGruH1u2n+N0uSR+cNqj/94edTxvat5bz08Xf2Ps4MJW2v+X/ytCyl
LCH+5fx39YTF2an2UYTsAQjvpKsR7UEMxeac2aki2/f5vxZA6KUklqb/rK9LIGVD
aA65ff7e2RxwGXRm4xlnny0mnELpSXm2of5h1G1UBzAucQrTLvhSCxg2bcamCe4l
4gDExf2VjbMv0wKkyPPvuoO7tU0g+AIXn+NdzpioGC5uYAmmpXDqH84WVBhs1Ew4
ZrgpwbMRJHwkOMbWlKiAZuYxWjUneeXeZ+CYIAGgqNZT6XbzJdwTLTpT9HS9lUmz
jhqelbXNjQOWoST/jzbraQpotYbOIwbRlfkR+jUsWGqPDBwejOmi1k9E+WF62f0c
vu9zieQyEirEIJJuVF3sGZ2gs/AtwNEDR0K2EhTqMIU7+9jc/xZnlI9qS4weQVPw
ie0WToa8bXhavuWHWRLDCI+WEyzY8IjvnX5wT7MaKbsqoGJvNJdpOmJn0+5+RQr2
OBNReVieOj6QwpQv4z3aasbje9fR7mWxXG4RGgijK3DJSnhisWgKzMgfHMLn+ez3
jjPaQ0zKFKNBAM/DwyFPpwtlYE+1i8YTrVkByjetesUUYuGTmOd4JeCwVnfuPb9S
NUa7lKx8r1GtR4vyESzNg2RO3jhCy3XAGt7vJKX8iHNUxzsUGG9cvBMcWJ+HqeF9
CIyJ/6da+GS7Z8+RcBzidQ82Yzrh6eofl9ono0z03XCAwjNEcazOIKFhqkzTPq9Q
A7Z8zjgaaaiDCdZybkhrkBs8mcG/k5GyIe7JvemnMcyZQG24L2/H84w4so7aXfoO
8zPHY25eNjU7XEg5wl9NHOYjEvkn1gHR2aC2QaWKgI+yEvx1zWJqBq39isAgQYVi
KoKXKtFrW6bg2p+I68ZrAb81FBgRgovEXSeIcsYxZmfpNVOBRT9pyF13dscdF16C
UzivfbFuf0bYIQCRw06ODybyI8Ywc+Na9rNuBbklFt1BKxjlnHr4r5QgkKSFM0xG
yd/51jV+24Me0v9KvNcT9oBSoaxG/r8L5SUmrQUzj/1aJON8//Ylj0s0gHRvU+Iz
K+lSerBQxj/BpKbXbi3TmlLLPNtMElM9kt8Hg4EXM//FNLYKCHPyv+pP17Vxh0+P
Vk0V2Hm2ZCw5f/jNlNUNOOAe3ifh13X1wkr3i7p6Zm1QiF0fLxxHpRF3cEH5/y61
ypCrWqCv5BagKWsIi7PKy6nUvffQPy6/xjDtV9qhLHxlHjOS2RM74fO+OSfnCJi2
dYN+TvrvJfNtrcGrAs1gMDi5U3KJKbmMJJ1se583+w46BV8lYEKJ67YLk3uEGURt
Dh68r9jwP8qRTGg0c1kQ4j+3ofHlvNBxAJpiNozF3GGQcEdnnzJiaaNiUiYw87vF
DLdVavHE808TMQNHNiT/fhAZykowYvKkuRC1LhP6TTgywoZqqTYb53W6K6E2AhJ0
41673oCe79vUXBdHKqFIky/BH7Dkvhc8TxDjTLxAzZsPJ/TvDAlTvH4qPUuQ+9N3
yEwt7AzHC63Km8Ix/iBe6tezjRA676PI392jZ6YVPWkZbOtUXSuYVkun1sginZW0
aKb9hzWUZhMW6L1leUGrRpOq3NV4mgwH68mnb+Hii7jnBigL6/HW0aoRCgJtMbMy
4PL0/B3jzVdAYnhVj4wwIcpRHDIeUd/ylJGLrlgb4ZOryF+GI3eMrg0GatdZTn0F
+gXj0eXXziX5+/qHVujik9PoWGQziGQry1ZZ0/PdoYZY3XbzkDAgevXKPbwh0Hl3
1+dcUFvI1nxm7qdPIoJR4ZXmly2rIrD/HQyabhkFF5bwtXHryrCi3RNfLYNwHixm
D4pp07H+VZWl7eRz7GyCKX/74WJOnKVoqCjc/ffiKl9vncTcTRnifqME3JnuJ/nx
TiT8M3NxeXJYtERRRkOJgPIv9yTSmCuP4f5vGncFKoowtiWnr7CovzG+HgkzMcWb
zH2dn0avvHN4SXq2N/Wy1XzGp3KJT6U93IqP4BVUq8MDJINPCqAbTv2i+SVKDarS
zcaWYc+k+z/AbU+BUgI881LeLFnw4Li3gYiVBPKFtuqCZOVdyxaQn08RacxnEBFE
aji1ricHqH+ZWbUni+wqultHnONoD3Olf8Xl/ULB+raZOOvhmY8clOc9RhwcFpCj
w30E7m0T96LcLzhc9B+a2RXI5k81xg2d/cvEmVH0JNMJQ8sSlICW47YmkwV3MFpf
+ny6OrEbivgfGo8l1CT7pZ3xEuyJsdSkiqKhKYD1dsldFAFspdYmyxGLRH/vGRuW
0sHiyD1SfVr+6wOXs9CCPoI6pcT+u58DQKajaT1yhvfA4GLHQwpwAAIqgxcjTDoa
YNkd14VjDz6Uv4yDaW3yHBZNB/JX5uQTXb351s/gfq3FYD3nqnSsHcYvWPbXcYH0
N07uzo/jN2gCMrGBvd9vlJoQUEgaoKje1nZG80SNIBU7ax46rG6GLbroo/EKF+6u
QXCspTJ7c/qjgszHYL7XwiVLaYhbhj5uCdTVqZjYDoFxH/2pJmpEej8UBk2i44n/
5jCe7ow7gaMvS89abdztEB8sWJBSIQGpfxGsCLNeTzM4zo8TgPmSdyoH/pWQ+QpJ
drKpuG8Y3/dAVyomVrIWAu6+PhlZfmCnf7LDmhiP4YmcYTNKC1GYoQBQm5wwaDNd
Wsjr86qCw99PYXXUoNSBK37WxsmkdjrppVhT43RHZd9JIPLdLozdAFmii2RJineU
fSnkWMC83gs3I+gwdv+hSZnAww3Roesov4uoMmC3j0wNlDP3JX7CqJmXMlAjfGWY
FVbgvvNkaNrkoWLLdpcf/oO7ydJqjhuYzaZBDqWPvdxm0/udRWBHOs1Z+WpMFHOp
OiCNuybDTC1THqrUv8hr/lLUxOHAMr354E5IciOD14CjZBnXlw6E3+9qsNIHlBaE
dLyZWvCM++FqrP6gfNuuMUtmcvp+q3ISm9SEJ+zdKRD3qtSZCJN2xiGGMjtZltE0
k3sSd3pHyFdVn8zOyAn6jwv4ttu7U2XhVnHw7Rls8yfZk12pWV23rB8gO7FQFBnS
Ed15Dzt3LviN9otS9YftAglit7zz8Y/twAcrxqLkFnWvPUrC6uDsb6Wm81MXshhC
GKB9TRhw+pWS4I7oMYUGmALpclK4dbif/UqmSa8dAaKsIqhznqzujHI907+nr2zr
x7lRpxexWxZDs/yZWxZ3PO27hasC08eBKQssGl3wTy6paInK0WaZ3ozMPCg/7Q1Y
fe1vRqr/b9D74g80KkY+pLNtWKRH/WtXuXAKP8g2pPV2ucAAUJACbRD7z+TmN/XN
b9j9Y0Mh9Rgr8b0O40ijdmzDncU8AQ/SQpgYuODfBDBQ1NHIQH5rsBMIjfrI+2vn
dTfYX6d49tkI0ebkjAVzKKOV16RwS3ShN8MqMaXXdEN9ngZYQUeROfuRVSlpKaOJ
Bz2xQ3DJT6ScA8v+q/OIWAVFgojlth80npz2IynenLxgJP0h5XQ6cPXjKtMuDVg2
8saKnD79soFghvbBY9ddPwYIkNYJY2qCeaQQ9uugOFZBu1ycIEDY0633u6wZsE1n
bAoyLXbatWGwg45q1WXqdCBuw4VSLQrHTobxtvoDno2Fk2REgYFJYc6iXKpvjQuU
39tqd80CQEVbrnYoWsLKpHbtTmAUuDnax1KDQwqj/lLJP9I2j6G/axwipakD6lVC
ETvjQQOSHRBGu7FxD+aiSvxPBAc0k5qb6rwSKjZRQcCljoXdWduANPRvpLJEYVwt
fyR0K0nb7+VGvLOTJ+lnxK/24l38krZ/1VyX9TvXNiB7UyHJTSywCCgdAZg5YCCa
qCFNAof0FAotlpYiBzJUc/TVUMUhyi8CZVcXLknaqccbuj8cgvWxrU6/WvR+C+6C
W0bVNR6SviVhgJkMWKeQv7oqYrHxtBqaKs4h5KlJ2sk6GCGGlyyGcHkkp0F+2dni
/6dkEtAQHzgmUAcBMBh6jpBs8/nqE+4FEey+bu6g7J1NzotgT1IkoVFh8elt8tL/
4lC21NYxoikcdlMaPcPECWdkbX8qxzEM0XLRwq0nioTvO2hVHCDFvSz6o7+1aThg
F5nyvMwYwT+2xfQMGQC4A8vp9soQCPMLbryic4UZT9CA31qpw6BtPqjB5QeWtATF
ddF/cDEnX1XLjW2C2y3ob3hbZdOjyfEnab64ygaqwwtRvwUcDfKIBJhz2SOiDaio
d/J/UCtuZzePPK660Mw1Sq1K9Q4J5t2qpQOlb7ePpNks2n25J3lfbpS25ASDmisf
XOWY0ML/T23IsjwY6UeLmOr56ZwPhyFwXr8LGrr2+Vz7lcbUXgIgKzuKdVBSUZvQ
dlADkefrSCRrxBpF39lSX5u3miaOa2hsBNRHI5miBpyYlbdcyejfpd24/Kufvupf
wxx9LlxsN0GabD3L39Zb6hk4nQOirEYbhRI+TGK4CP5Q75ICsz+dMmoBe3BJN3vF
vznTmyqCtOZu6jsr6i5sLAQMUg/KyjXwvi8Se9wJ+/m1zm0LSlOuVyYBqpJox219
w1bcXWlA4iQWf/UnQUOB6hF2t9iLdFsWfcZ9Q8YI0VErqgF3Yvxy/jcGVko22h/5
FmFkP+jBogd7j5D5X2T5k2Wu8znOQ0+fQLkb3u9XVPunj7BeEdFpG66wDreT4tuM
fEU7g6OumMk4idXGcBfqqgkQC2Qi6hCX9sYeE9+3s/fmFwlw+WDmJExpaoj7Jm+L
++3D9ScnKy2sNN66VtnXcZGAIH5NRVtzEYk87sv8pZTzQAECzi1TZBhoCkyysHWq
JkE3whXvHjDB9huAEVNmQg4u4tD05dK7CFscKC53TBvVBwE15sM8srIZGFJXq9cZ
79FlJc7Z/gTw9HkU9qV7+GnwYPMjSfze93K3uy44fdogYmtMfCgqSzfEAm114TBJ
Z3avCHuvAEyR48O9iaTDZ9cW/2LI75/D2ahmUSd8lhXMRRLX9fcv/F4mPttDQcYq
UkmVQR5aRejAJ8GbM7lxqXRnydkE76sYs5AqVu48VD4KbOiuiYO3bBOsQmm0lRho
Hl3y17c/Nx991OmB18apRFQLlD2in2ArcVoBpAqiAvbjgvSXrE5zSuccBRagSuiG
qfggQYwLFnMDo9Iq9LDNLXxdWgqtKfQoWYnycPwlcIY0ut8PT3tnnvZGjSQcltXu
dKHDKBEoahJvPNEgN7tQOulUxxy9bd4svLFosJU4gtfmy8fdgO8HZC3xeKQ0BERb
ctIZUbZPmKZCO/OvD/CbUkCZGRYDej96SBrHLpaFWsPwTUXmK12S9Eh7d3aQa3UF
ZcFXD08sD8n2z1dlCycL7QLuszhfFReAbuNE2tejYTFOpynDVJrTKYxVn/p4N2c3
oiIm1Fwvey3WsbULsE0uiuHTUqDDrkg4jAPdPHyE9EPpH8uTZyzIP7gdLhDTUUPa
4du462vcYKxi5gwkox0nfvtadM5yM+pdUiCDEICESbvge77ZcbJTJ1B3an7q10UU
fBjmCPawtkZYvVH0B3jrHNnaKQei3Z3qyWM9bQTku3uEAwj8yGAQwzrYBq7NqQOJ
nDc/e6at7hOllfpStWA2i+h1oVjfg6awj0HfzkCKI1GTHiV0HPoqCuTZx/cO4yFD
sO/VtMjMFJzTatzAvVmpznKsOTO+70xWRx2gp0+pvJA5J6WpBJ8hEJRXnaJ7vcuq
eNTXVWcuRzrvspxSnl8tPAHpU3gcWxdOonqpLrF/uZAqgVct5gKEjxeUx6FaK2ds
OVYl87ESuAWvAXyFBMQ2w19+Sy1eGhaL/d2rhmWtUyOyJbWIfVwQuLnHBL6+ONgu
ZsnM2u0rZtCjEHowphYI6UiMdRz3xNG8Qgd1LTKr1grQOHLVtNA7ozj2xeiczrJa
UUtKNiMNOZw9hkmzOkkYg10HNPSHqAtGyZE7kTB4HMO1qyTKYK72v4JAB6wfqrBs
TXNZmjccy92s5yf3g2oXK/OpXwQYA/QGcZ43w31GqHgdvYLD7FmFbvGxGHZd/Zf3
diCGwO/9aRAwwl4PNmCC9+qlwVugSrN0ZAwfUNWxawLsawsykWLVqpjLhli9sHR7
p+3FDzespOVGvR/Neluv39Mb4iKHTAT0c3qtcyHaH3UpXtlc9L/P43vGFa19QCqU
fyDBWK//6F4KxSv3nXi5c+re5/7DeD6sOd0ou0wlxuZVrtt78TQ0IHFnKC630Q0y
yEuip93jNI3YCQGTdbe3w9dJhC5E3GSdhX3fjN8gW3XzZHPw04BEgu3p/uChocCC
bsR44LVTcClhUixtWjtPPG2jj2Cb7YRz4wKswvcOJecTFSL0mdklUB7dHmstZr3l
7/TbiYtBxshEm+OvGflxoiDzn3sY2NNJyO4RzBrL9GrN+SMo/DtNkgoo6odgCxbg
gm9HExHwSj6czfYScEDPjr4IVXcwEg8/Ge3PgNUiByPsqY3tMsBMJqOFo5uYZfoy
pFL9jj7N4xVO9gtn2PuYyWVVega8yWS+0gWLeySgTFQ7f5m5D0oUk0JjbWPkTjrf
5NvOCh8l/ON8l7DBspXl04vz9V5r25lTrLyl7QCvSAGV8AhnSXuSi/ehAfvS2wdt
ahyFQhF3Ioi65pEZC+ljFZwJFDD9AnsSvx9aGVzF70YlV3JQp2VrE0BXv+n3PqLf
WRGTrI8PltRaM60FC+ptaLjXNwLp0hwQxoJqW1jCuNZinmrwGN4vOy23j2foW371
90briYUB2yz+ex0czIgAAytP39v5ZHV/geGaAmiHLUOEpBwQCoDZep6x6SaTv2T0
JdKtqq/sDmONkfHLa0Lx39dqFlSNG7SELJd0PcDT9BREqA97cIL/dXzEqZC91abv
wPqz0pxdvCk74gw/SyNxcUC/OIEG4KO4vnOo61B88XozmdJ07SdfBjiVRhmUOPPl
dvHhrh9Zoqvm5clACJ5Kfyn6vyPzyzeyOkr+mA8WoYFbXzDcDVSyGs1IDhZ5S5bP
gBIMrYjKZyUOyZQlFlU8uXabDkUcFOuiPti6Hu/OW7MElfTJojlzJ7wdtRVq+3Yw
SxZPGgWRM9/pPlBHvywcdz1bJU3sE9f1COXyM02gBcxMcDittLErT5k2kQvzLF8A
dQu8n5KLnoQE0tjOFv6mbFmPMmIa4WQWFoGi8sBkRDfhf1COug9V85rXILcP1GK7
Y5euitSo80blXZEt2WiGYeEyVhtG9hG2hX75SjgDKn4RduFG/ohUTowfvhy/WhTv
F106Dlm69RjjFg50kKWoTTVwnJbWTKaMmk8LzfqI0rSVWWdxOLw4swWGoS97f1PN
iUctQ3eXW50uOFhHFpcLuuZyvgNTcMCRKf4mI0hN6uviY0G40uk9BNPcmzOFCo3r
xF6pWlwPkNKcWFh/ckZqm+cE6FhRAZOAsdxP0sxuya8hISy9IlDFjquFBEYit9a2
Ioor3wyHQV1wSQR4boz0Ux1PbFBAO4ZoTvZ/f1KTs/5W1gXonC14ugGcBpyAWXKg
fgn6Ba3k+LSsuexlEUqF9wZ2XG1alA4PvtAUaPXAllRZKSbYXZcq75ORbUpxZBbh
SkACHXGLzBZ74NMeP5zjHtC794AxSKdVRk4CWtVrOhi+yT2PlXJ4R0/yb6SvgL3S
ticz1mPUOowqTNxztig/4mdn5MuodYV++DfRaN632jtb/YhgOyZTwezxolZHMmfU
7dZHqMFeOkxJ5hvlxzvj+cfG+vufR24QGsNGqfv32cUf8WvL2rybX9UN86X2vhGI
T3qOIouAF6hN3XS1sQckiPw+qaRHM5RsMo8smNgvDkTwZxEWb8EyI9+N1J5df4OM
1zhW+jDTEAvEVDph1dO3nUGBwGu0MDafDTwaTKSGqlYlCou0n42TYO307dlBrmmG
O8GbCa5vDSybghJyO31J5vDJIwNuLN1QTN1zQEhNRchS/LslDfebYx4z6ZSICVOK
rOiQYDmZ3WCpVA7SB+LyM9eU8HiJevdyo7U4wYwss2x0LPoPi2478rawWYoPOWK2
tXANFlloT87jwBUan9OChAJq3BttMT6v6Oj84zIgb2c9XBKqFdKYasCEbOAZp6mF
OzvFXsiNxg8LVCdIkDRJFroFRsdAFftGYq5Abm0QlnNNVu8NHwGPtVeyodBfEx89
W6fEaAh6lISYEchw3xMA0fVR3RU347KMOzG79PRsFJ3DWZDK/Sy7j85eqYhnnwsS
abfZqiEwkrz6D7POmPzMjA6/JA2cx9BpctZHgtuW3PlA5xFX4aCbwTb7UH+zRnJ/
XNUUwKvRjrJWmi6Dm/1rX9ZG+7NrFvunQ7J3uyFGKkTMIsUYfimP08TTTlpYIvr0
JIXKKUSICCV3dI5QGQWVCVE96EHiareVfuO1m+CmlR+Ju0zEDG3dGwH6IO0uJg9g
SkxYBqMFwa4tL+AyGz5Xbce31DN8Rox6B/7HTJbpBSBEbitBpRvEFnIc8Ikmceqn
FG9zOPHtrcZ30b5lFDWmTLxSQAI6sUFi2BtGsL9voBO+aWnC4f3411+p/4JvzeJL
yNHrtXyhvT545H1bMBoK7ziONRrXV5ZolT86/hFL3SzHmDvznnKlQkMdqPfzPRci
rJ7hu2xbmo+AbtfDZ6BFlkUuCbvm7STuRCkA9vJpw7lziXP40fPLdhWHdZNhJPOR
+Yy7AnKZEcBV2AMovVQI5fKhuhxslGNDYyQufVHlgE89w5QcWl7zdgKgoT8wX9te
thV4ZZPaBEI3NG8U4ttn5A3Wd2Bb3ce6YsMs6I/CUDhm9h5/ZUMQLOzqjEvDIi/w
LhHZnY4RIKmUarSuB7sSFFgUxvkDi3NZIjiU2YC3QJmr6lc8fcBFbnse+SKvS+VH
dFJJeqkvfaV0tW2p7jBO6+9wlq2ktg+y2xu0aAWEkeksVocU3MIYnsgJhoT19u8/
NZBRRRhDx7BP/fHFuwLHMEgFYhf///kQKkkI1eLhh1OEUftom+H388vZENd+B+Ed
t/EFklI9kqIS76aT7/275EnGPYm0caPX79KfRHc4vlDj1L3uZvhpSXyNID0dlkmI
oiF5F/sF3AQSDJGVFy+0EpPVXEJHa1/RA5lhmMHfj/WuAdVf93cfBS2FqNvwlMpX
iITe4+JMfA/S8OgnbsTFgcQ8LVD2j2BhDvkLipV+NDynmf3jJ19m/Ug2zb8GwXDC
6oZ3D/8Tg10bhYeGOoCmclrmUTckLRo/ttFF8avv5QA0l22FYF/5CJpZGCOeUuoi
K/dxi9hqBSfcAh4Cv0FanF9LQf6OBLBLiVu/vhmIr/smQa9KL/q1hC1OQJGaWQ3y
K6j4i50RLRMsBFdjdUU6Rz+X/DkFygLuIVWeRLZIBF/zoHXxOzdAw2IrVEoM6ODJ
tVFYlr+2SChNEB1zrqxXPaSbwdMEZ0Z4ShbMrQeISICEMozuKujBOfFMoGuXwiyH
O8vpJGjjkx5xlHMJ/YoO3r2AGF+XTZXFBkemeSiw11MXb/XShTgoAvgqk2JZTl26
N/Zy6kTDC1wQpqVKX+1AJKV8JZFkXPorFDXbtOXka5pruC4HG/E2ymZew/aTZSnB
EAJZyROESX2mmPWWqvwqSCaL7oCMQfGjgo5tJMWxJ9LzBr8BNuqGBAuxImFvtEJn
0uokRkM/bf/O5FO/6AAMcKAYL1CwhkNgV5yvlX7fl6s7BaP4Kt4sR7OI9odAbyAG
bayamBaztcpcgbaBFamfOYXb9TyLmUVFfl+huW4BZAy+OHjr1wE83O8ABgn7xnc4
yBYuy9uTGe/qRrpAFPZv785TEJitpBBOAUcLKXtDn6mEiZARrU11qtSapVwI3emk
GbQOPusq2q1jM315G3jg1y2KtLhoqC7VaVLuscTBOpqbNltVAZTX8mReKrWm+app
Qby/6kWyYRMNlRY1ICoTGqXP1EfoGI1w2TeO2gl+TS46pLcqO+6BnJlqFfoOVXnN
8eQXE5T18/lw5lvM3TQuQqtOimrG268X4q98jFQClOioWoNRkof6PoNZ4ipp6vde
S50c6ViSW1Woih8pnlGlU/OSOFJSn6axodLAzl0pQiYGLTRRlfyY/BWM76YxPRn6
Uyl/a8TFoWqFDdX4lKXlD4h70Zg/gOog0w9Tm4YIAFJKYX1ZcBwNjAUjs7BFtDhE
TZszorfwgOAj/66shSJB0fg8xTj2iZ7P2UNzu7RzMvVomygCCMGr4wjGl3Q/psTO
GvibJXiYd6ANo+qkGmPRdgT92uy3BY/73HKUgnLT8tgeTRZ37Oee/8mg/gJAQYqH
RHq7NBFi/0xPFFKiGLI+b+T2OpcuM900wO5P83JqKq/y/GX81o2sfkY1/OG8slYu
oMja52XzCKFcmVuavCsYn/3n/G+xMKkrihLuMUvZ72qvOncYWa2acKLtde2C8XHC
u6ViAmea02/EWtkD64XYKHsSrIFlRdoOjdWo6UtDMuLzvKN1U/Ai4jiJEgbN4nWv
1JnGDAz6lSz3ADNP+36Z08BrJq3XS2ruOM1FU4l8TVahuvxSpytB2ofXGMh1uGNH
KhZYL+OS4GM6ZIlMmMBD+vSWDmi6UwIk+ZRQoTdjBZB3oCMFtGgIJWY+tHjRkpmK
KElcmluR6yt2kuSsa0IeoLhjr7tQ2kgABRiMCFTJCUnAjjD4aGMzjRtaoptO8BUd
HqVWZep2v2WrBsreLjWcYCETFTE8F+lO92y7RNPybnFarztQMXMnsN573GSWuDQ3
k3dkRtx18GmtHT3ztZueSmo4xwTI+EL5y/3R52iQyPSIlQk1fVsNNopTVTS4o6A+
GUbPknlIv5pAzLzzYMCaPesetJQN2ZPue/wc+n7ab/vLCMxFLYQkOWjGi6l9gTsA
bxJVNqviIEX9laghULDm5+MrHvpLwNOpJsBdfbavMnvJ7NxcBbMgxPWeomQs/BUu
WQ3jqOIuL2pr+2ar00SVZjrrkwGGjd6CSQuRtkT4iMxbzYUh2Zmf7Wx6Ga8HNMqL
otYacKsrQx9VBVWirjfG+fhv2RvO9D8e9I0ckBxhnXHYlFBYCsnrlDSPjBwCx/EA
1+asYtdgbrLtL9wIiraNTfBFosZz8F23l+KjRkEm9b9FJJ2d4UW8+PzJQJI+JJWy
ydk/CN+zmzjf6LTuEGNY9LHsfgraop/hZYtjnJPBe6Y3CfwloBnBG7I8B2WOyiyI
XPBKAECSZsHAWKiaNE9cNUeZXg2sC6VZozjC8+nTbPejnD+V9Ezf3CeWDDM4oB6q
O2HnpwC9SBfa2rb0QWld0dr+8LyF+JIVC3M5D39GDYKhlXBsOjnOH64LS0tzZ6uh
feYMxI7RgxdfSz3l47F1jVh8f0/iwFveP967GU8MfXPxp/rsadhU6ow4IfbWK0Ur
bXvjFf2qpvxsv/+REUHKvAbbUx0UTe0j84H6u7AbwqIV+abLgrGVRGaCIXcEdEPQ
Vi+dSnUkGNC1CciKLTSN3BkzdfgQ41DAMHqHJqgaFJSrZLWtgNaxLHq+1dFF/D76
AeRYOc/HIlcFlPBraTxeHbW0Y9udiREU+Aefzxb1DssoBxK/nHaqzWUdguYGy8uW
fzS6RgQZru34gWege/oBd+oqLVwmImwOaUIGzKv37PJiKwFkwNPNZsKq8/X973S9
5AzS4m6qM3QSlW0M7ERQRFsuwLQcr1Yqby6IxrQTmMxu3ffkOPQbJG9aBm7sDuhk
ZGnCBToTA3hU36xHQpIZzXKB+vEO+FWVlCzatwD6VRfyl68xIh95oNnpzj7rDMMK
uAgGxkge8A3ZDvumP3O/r3FjBE0+mAIdGUmSiuGSWbHDDLg92435e5XnZDDXgkD8
ZLHdGxCSRAYjIDQS5+ImEos62dI+MTM7wWoptM9GCfQErcbCs+gijE2f8A2C3NpA
RDalFdUYDjy1seIrrnax+QPraxt2OuwO28JUPMSdqLSd5t9QkHf/2k9FsSrHjM21
6LKs4SaANKp5T2RXgP3QYczGQDsaj72beI6/R+AvnSpUqIlOzFjtLb0nu7EJfhNY
jbcnSfRoV3c/IA7Sm8oORvPWKzsV9KT2iyMfYeLWPMcvBPyQBh+Q9vSYiFcsVawM
D/1YgZ/1k92c+EJHLAzRkxIC+LfkBI0B4KFHWd7HAtMGouLtSj5NyndZmIRfrGkF
VDYwwomcK6q9BAw/Vf+xo4YTpvbxtwOkSdnmLJn12JQV0RQjrkPk77rWniHki/qf
bX3Abzc5QRL0jY8JVb0cUnA27RoBOFy576h0VUJYD3QO6D5d0PEd6S0j3eGf9851
R5UlKO+FlfvuZDHa/UDqehDvo1FY7uuAwdn132DiBg+2fRHhh7lslIm5nP/661Wd
Od0+pJZNHvWdsy6qYbuASFHdkKbyNJQhm6k7kXmZwFH2OJIEa43sjJWaFoGSJiDP
VaLHdQxnLHUPtl/sOceVFDdIEIcSZFM3GMN74QYpvi6IVYLZbyYcT2c9I3JyMkq8
9l5a7fMgc4aTPb9AWop0b69IpamEWgBZNTgBZC0gr8dzil5u3MPhZLkLQd1B92lR
sLvH7Do95otUIERvUTy6H2W0mIzN2DwB8r7NDl0A3mnnxPviliJ+fM8Ko2tSiQKB
OBh857e3sI0PWX2DloD0WpU2oRTiFosZh7DaNYqoHR5OCNqOQGMGU/D9yU9k7Qrk
UhSFCyFw2+kgSaOopwwJutVWeAn6GRrpc5+ysW8Kvwgt+o+yfPCm3Dh+BmiGa0qT
lp+7JgVA0GmdJPlxtdlOFbj22E+5B29mQzW6+Th9C5lRo8Q098/FfeN+DrTFcMOU
a4LMxfEJmJlJX3cElkAxDXk6Txvr33RumZ9dk9Jilcpn5hBe1Wb9ijx58ff7zt2p
v4saX6RlfPBp+1a08tbVDWgTGU3/eOurdnwaPVLKzEtO4L3AOZhZdyTLk8sOVVsb
h80ga1rrefsYT4jUoCRKKiZPWj2yWTIiV+xDigFvRTV3YNxRksQ5DqiTa4Oo5fRP
FJHQKbzhhPyFK8lWkvrwtYS1QebofRouDrZ/qeh3K87wPeKp2guLxs5TMzYNc69S
8flNfphS0bqkPOIumhF63UEceACtk1Xq4flOpoUla3PQ5LJc1KW+YcolTaYu+CiS
td1VGQsmWeJH+NQY19i/F4b3ZM24RTVVm7n0V4oEEmQ+BtE0mTqx+8Ruz92qx/6E
q4ZppSGMZ8pICHhoZFWyD7urmguCPJnjxaiY5LLeL18lGSRdwgu0rPJ9L9/CvXjO
PSufeTiwgkHs3ojH8+zFRQoKnGSRbmskq0eSKM6poUWqKHOeBNI11ErzvflHeaHj
SwHRXM5J9HrDD+16C2DPwYunfn1sqd7FsLarlPKifKzuK1oNeL823fXXIs73LBdy
xo1Ed/Y/Px096fl7oldhy0HBTmv8kH1IFpXVlkj/pxvPilrIZw33Xoj4Z51/r5do
lg5T7vMhHaTKx4ilR3ThWYUZ5d2zHziFLu8n7OdTx6Nn2VSQ30jv51foWYoujW8N
V1XCdDXp+QpBoRn/wurVYmaSpToN6MW6r5DwYjwltovHZ7HkwttNQywmgb8bceRk
ht6WfyETqBf+wcXCSL89627NzrCyj/UqdrrdX6Tq2w8jrfPKXf1ePVvMC0ydh8Nq
chXHSjRPN60sk8myig2jOSnjKu3mgr4HL3n3ns62PCgLluVebCo6CYDyXct2LSWY
8xfY5rvBhzvtvyEpfJuXgk3wip0wi78W0VpH9egiPTKPLuWxPw6Q1u0ZoqR00Bs+
GErhNc7IreVxfR0ecXiyMdNGQLo3xsqUPQvJnnPa+TpLaQyYjV/Xsc+g02LBYHHE
/OGVL3fMl7cSNOfAMwtp33mgEA0P2a3QDZPFQxZeGtafj+D0z/6JfOisfwafnY4y
tLLn1MEiNBMLoiy/YU7NTmweLI+fqZpd72lct+ifKZjEIXp5u005YcWiXDsEFNFA
WtatqEbehKL6pOCItvYVsPbANhOKCXW6rf07J+L6yQRjFfZjcy0C0pBCTk7h8+aM
opxFG9EKN9aFmcvmkO+pvh9VaTfPTFoIxJds2xt6FYITBV5Y2JVwnByFkY5Bu+Ye
uKJajMNp7vY798AR4XEBbVaIjgu8COYjGgrzePegeb2c4L0pIVzv2jaKPZIevEMl
uajO4/KgXAaEMM3t0YLqb/6AVxsWCSof2WwQu+n9JTB2VGtpuQxnp50KzZQVBhxs
J3HEkIhyUKYYEr5+FKip/WzHQpnDvVTE5x0UT0yH/kUJAscr+BIFRYFbpReMKHQC
KPtjf0ht7BBiybE3V8EO68dMt+6Jgp54nz455OM/lyiXje7jYIF1sYwd3M8inGWd
olijnh9jvzbAvwxx41bgHWoxq88vVphVLbKgJzTJKTJGs1TOfj3k5mIMe+Z36Q7L
jO9pYEjO7CvAqrsdkWPfZV9JxTiBmqNJ/SSjW9fycEcW+XggQ69eq09y+vRWTDAp
z69es6vGuuA3uX4XW+wD9+nL5+4eQCYpZdnslNT/FxNjpVHDpLQc0SBtqlu8SfGa
3pCuWwm8k1mYih4RvSKKURfkAiJwOvgnVTL01KkCHaR20XNDLjQ33t2Z9fMvTUgT
XDca6+OV8p4+9dP3ShOgMvp3073U8atD+aFzWte2qg5tO5uLGyBkcxraInl/pCJo
nOSPj5VSzjPEWTj/Agu6iPTN9yvdEnvkuM16b1jS5iesWsn23HKtmuNN2XcwNtQK
ultt1Sm/aTyjBCWNfDL/BpfuqDoaQj5Ihg6WrO6k09z9ss7d2XnHdNMoWCEPROkZ
bBfhZSnF2L84OktoH0NykrUv1G9paoj7f3fU92zw5ergrRPgisRuRi7ZtV0/5++j
6SutrnYNi73UTi0F9l1cmRG26kJU0sPS27Bq0kJ+wj5V+FxgQwgFOgNFw87uheva
sKDCadfqv5xnyn7O4gc8pMU4OxQfxw+M3s9nQnHj+U/e088IoRO/Ousp1wVKnunp
W86KfL7ytsU8ssHZAW8FfgHbVxaNjMHBHcbeIMtWaAdVX85ylSlKiLc7v3Qp4kVM
smppKVxIfF2Bid3IcOQ68RIpzFvTKVZfE6OczVsV//SJ4aF+zSvStr+fyJePFj6H
BEs6fx6rdRu6VmyFrYZjYNIZ2FI5E7n+/yRm3Pvo+8ENNKa/J84HnKhxi62I5mN7
Mr6IbtRM6REcg+xOUAFAK8jlQUuoP/CsIAYGTGnLqYgUNzzBG6xraObgEDCZmoGt
JZBidoUSCuCPSXKrCjnfuBKOxxkYnRjlaMEOWO3EsrQRMosj2KfTcGrdmg74f6Yl
0VGghQsl3SsioHb1KuousGfU1eE7RVDAhBJr+J3FZbf7wCMTqo5uCdEAgO/xT10j
TyGxVNlTPBJub0LI/t+u4hXUTUH4jX3lisqHaK/y68VEGdaNUkc827x9Ip96qPM9
f9d3UfMg6t+qv9+WkhCTGKAJnkNmHoTVyVaNuADqJ2oHB7jqBski5ZdiewOL2ke+
dNz37pvKlJ6iFXK3SlthB1H1JXqwwL4oaftt2tIJEkAPTJixKUQL9iRmcg6ulS1w
4ByIzhwi/gZ8Tf6L44k0oDiQxagje6bazzkm3796iUBG3wY31ytFt9TkC3smlLto
xz+Lvf8SG7mnOrtBlBEjuD3AUAGDOV5Bfy5mpcPiqXa/eX3brS4EZacqeSwEejAP
bBnm/ASKTxH2grBn8yoYwWditoSU7mC8ATxXoevEptwiS0FtsVbmzt46m1l77LxM
9NESmylfkado9sM3bvHr9OAizVuDHcjLhxXIMBrV79JsGnloOIwvb5hQPjfuZ+xE
Ukvl4lkQSebxazB6W34tZxCMM0pxi1SCk+hLzPC506WiTS4y6Y9ZSiQA1rEt8w/a
7cgbhIXc9Ch2mtXABf6+sPAEC0xCoRRdk8pWChXBfsjONf86PaMVqQ3kHOSm2AY4
Rp/3abtKo1gMbxJqdzCWBujwjbluEcSI7Upp/hRsHnsS76Y3UDokut3eP5L5yi9V
yoDzoJg19w2bJ+fjqS47twJK1QmxBJwqHKUtGRi5Dt1LOYzjHBZOp07J1umf7+2U
7BLNQDhA8j56fYZspMdXY9eRO4y32dhBGS0XVxzbqxJpBPYwYQJ9FS7YgFAe28iD
pDfCyUF7qtnHZxz3bk5iyVLUtwPzNx+uUf1jhNpxTe1IbWFOr3mGK/VlsErtlrXm
BGrEPM2w39D3YQZzuVHm+YwfrTCNqg1uWfm7O7ooIbI5GIIhn7S/1Q8CC19yBDNT
8sIjkd/5qvfvUFHgJT3WsEqelmDCUi7CpR7t1NXW7zCrXT4yGpYrm2coIMlL+97a
UpVA1KxzLB9bSJYOCKV4XAnSNokpLQlaKD+hC5kI+Vm94Qy8YriO28sqBThEPlPl
+djHvLGb4XF1I05F0nc6qaOB9D1Zf2Zbs9IU1Nrg6a/BtlAupZ4+zPhCrFhC8FaO
EJcXL4Y4x/sCUMcf/QYuFAAMNILLzjtu9vPWNPu0R+mJbk0tgDPynmmQdmBGItQ+
aJ+c8k2MMdzcw2BXAWSUyhqg5k1myW5xqjt9aDyaSKQe/FeDEjqKBVb9xr5LdSw+
yi5boYHgB9NjiStY6c/nw79y5qU/gyVaVzVwUnAN7HUkPjfEONyFmQuSxVR9I/Dp
3u7SEJo2Bq/dBGcysQScMBrUZt/A41GcHZTFNwOuktEE1yz+/xKTiM6u2ErH4EHz
1UuGrJgL4Y5/edrwmLS5EDhNsnudNVJKXeTmzdUEhw+uC81nFp4miNiTzTWHo8M/
K5qYOS3Gc4AiMUCc88C4L/vZzhDZf9vjbDvp4j99MXUYesQKQfXOIFfTYUdJy7jA
fOxVqDVOhqN7Te2rU7wi+2utUnmv8O8VVklx7QMVXrjxIAf4jj2UzSx2y4OW4p8B
1aZFWa779aiLyF/mVB15/z5I33xDmH2mT1WXX03ThA1BaadmfnTxLDm8qyyLIqxr
pO+ZI4D3nTJNTl90mfqXP/z98ghhkMmgKO7QWhIjBfzL3HzWU+r6OX/mFvhqShd/
5fsl4TdaY+r0uDtIceyEVrrE4F3Jgb600LuBwmydLsITK1ZztvJ9RGIkLTnseTS5
TVGtUb7dimfUQDMOjFy3A8JGzAAajRhs/uCYS1HYHhUUMzJaiBBVi/AxHMvtQWy/
OnDeR5AFLUK8Zc9E6If0TIqHrofvLfU/HpSpJ/2clCRdcb4Il2mBkI8E4TLSV+SI
vrYAo9gP10Q1M9pZ3+0j1RxVB86yE3RPnuUWYcNPZ7sdpZBNdhqQPV+yiPsmQvKF
DSt3mKRfiJopGjD0Y5E0Uj2x4MpVu8I+fiDmRDU7ws+ZmTfLpiTqUsCf4X7J4eMo
jZyr5jEC5kAkL7vx7mY3dJCZa3RHKD05ijDepE317s5TjZ/xV4sp5n6hSX5m190j
OJSBQL5DrEmu0PGapC+z/lJqa+ZJmBq6vZMV2NEpbCal2qvEyd0KsFHGlSZgRZHz
qhyZiOjet9V4LauvNYQ4zbUEwWVrS+SwSTQ6+694EH6MpShAkBKe1phRh4jPQlqa
T2STWgJvGFbIgWyprFNLdk/gMpylAfniaI4rS5/fRQYfbgTF/G/CeueGrj/SHKRv
R4XOccUlnHqakSThEBxNP8fVJsxwUwxa2iWnoXnHrckUbp5/YH28lA5klvb6S81S
Y7Ce1BC4XukphQaxhAXWzjub3UIXD6KUSilHqfOHXwvp+M5a/fg9TqgEVrMi5uaF
zV4hZ1aABASnS+E//NAvJMJMGbusPrEoFUutzrzTFO/Ga1MRx81biSwCTD+E6YbN
s4dALl10iGt7f/76Rv54GS7cqgMKR5WoUHza7x66YgBqTh+zyS0hbUREa78YOBzL
nmNgf9DbSgCPhdHRaUcI6rYLiZcRwU3wBMQQBt2zdXmsVDpGGe55U24YphXDObYG
45n1CUMKzvh+ZZ4NUW2Qb3gc/1VlvQHPiEE3Oz+RjJsN9VVnrRsg70D5ONERKmlH
lQ/XZ4ly0irAlM9SK9R649SHtNQuy6W9FqH4P2c6+wDLdkQFEbo0It5j0k2IqiI5
UL0Tz8eiSdMGpPCu1xyBS6G1DxqL4QSu9k7S8zJun803XmJAKrKr5gU0B/og4axl
rXSaDkwh7zh9Qvt4seULPz8J3qJ8PksVWXPK6HphQcx0YJ51gUV4B/rTVANqfvER
5SE3OAiXFIL8vLrQl5lYenJcHA9eNHJAc6+zC2mFoVkkr5pGWFp+6qrbfA5vlv+c
l4qEjoeM86+Vu7CiI/3YVQPUqtK4oKUIiNn+kFdjj3cXH7jziWtNhaIUuB8bilPD
rOYISvlwTV461T/rzQ/VC9AExTWmgAFfkiUcmcxAbII3P+wPJpmUEBjZCpQwYgTH
HiAGa3wL2VvArAUSYiJ9L5RPhopYcIsZKvi0REd7TAzB/dnHHW2RP8OcACSWsgYX
A1/2b3bZp36RNNEwy2m6XyPF20dZD1+6Ge0TOzpzET68TJk3OE+1bQ8TNPUQ/Ew6
6OcjT+3KSyhKkg8+1Yt/bXJoN+siTnEiJDAS1l4Ds8rHVho//CEgaZqh+9OiG4q7
0zqvNpB2W19gtFDC/123h3AfhHbfb9//Bcu0EKXtD8G57X4MSoj88PLEXLebMDWV
50vQ4jJbLOKtPjni7+EsdRsULQGxUtPwEeZ4UHZebL4DA+jgl48unoQE+Fm2WzWu
NI4WdU4ihRmmZzugulN50EaRihc8oHJHFQvpe3dt+3mYM4qJ83sQ7Itb3law1iZQ
gpOdgCOf6fe7SVRSM1S2i7NNFTdz1zTre2ekCl+U04K+6edyLJOgs6kVYixfY2Ps
k8zrH8KFGYFxGY5uOsSp/MADkhR8vwqQAZgLoranLnlW63ttPnkKf3bb5QOhnfGJ
N8DPH6nA7S+1ISqcqYxXXUiqQTenVsFB3kgn+trSoaK5lgYHxpRiqfqf0rdAMcDB
z/EX6JT3oGR6VJzHfYxb9VnjrYPWmGMQxyC5Jwx9cYyajj2d+a8Cm6b8+KNuYqK9
iGeZ6YXmXOvsxTTagMxFMqTdPBJE720NY5Q6FcWEqqFcLWvn/dwjwp9GeZzIzp29
fLZts1EkcWbYh097dpRlRxy5FQwZ2ws5sVK/n2bR9+QZpbQGy6xlokYMDO5YF9TO
y3N9qXf0ZtB1bHYXGalR34xPT2mSsq1k41R5pmUhumiFspOUU/0PaB9qt2yo4Z56
YEEyYMVLOAgFrNG+Hxar9a7CAXdVq/dL9nxivDCRDFDLxXBJIdA6N7WM72R7p6z2
5xpkW3+05DK1uElP2NAGmg63AEawUCq+uMEJ5y+Yohxqjy+mLtmGRagkj36+slX+
mLJzGYUER1K62BuKbcP5ifBcmus6bgbLd8LPHu55Q2qULrZv4Mv5YhS3pBSNtkrK
3J6coUNIdJ5yilqIpiGly0VOYVaf4OqOTI2cCVfuYzVLQGbn469aFVyV1QXvP6NP
MwSxP1G+SV/z8Ql0n34DK31GBJiGjA/Bu8tNHAu+PiCEZkMUCk3oWPDSfE/AiWD2
8lxBqTg2JWj240rHr2blAgeO+HQi+5AVytI+i5VPcp+c+/h56d+fS10PPkC7vpBi
6HpyHXuygLZkcHf+XgLXseKmtjsatO4Fi+RWDsL0Adw9mlfvuKlARQp8YbKMdT39
+IyOs+UPAup7CEcFWtoeczGi9P9I1sswxB6IWuXvFuMC0ROFLAoxnIk+BIxxpHn3
pyy9DhFFQ+VZdwsCItHDT/FzpDlwbyShEmiVjqElnuufrthjA2+Qk+Oe+vxqOrRo
vVh/bn6jMTnrp+PfJC36mPN5x4EBuzmEipAVwQIP4p5q68AMdMlmF22v/zA8eLIR
uETdPrkDFd1mfxE2UWkfy6SurYMbO+J0rIbgG1n1Tizi9bNH8KIxdFLq618N3/jE
B5iQgcW13Y648ZlU3r9bFpcwjgNwsolZGrrFHz077a8SVSInMCKy2qMth56Ttmjv
Y+bdM7I0+94AThJTYD+IRjRVfRyxQhRJFNRjQBXqRK1rMxYwE+I8NN5rlvsvmUKY
7Vabhy8Ooo++/wE7PKpC03wGNtBIRH+QoXnf4P62bEXeVt8g4FNkMnrA8WXUQhez
BUpqxbE0oGS8VCoU6rMMAjFrRt+JidXqUkw2JCIG+aFcY5dgYIggH96UZGGOmaJx
Ou92dGB6mySXUvY4F4WpKoi89GHXhztbv7Z33dWap7gK/Bj2hknjOlZkaqul7raJ
FMq+hvO42JTgY9bhuv5pAV/TuRPstGZb8iSuPzwgywJAOCaQqK0guG4JgK8j2LmZ
1fe6WELmVOuSsBBrFmMtSD1dXhMRHDyqqkzuV+pYcfduJFG3+0DAcsP/gEv6UlAV
2BTEb7GnYzgLTTUY9BcbqWTKY3Bg1FvvWPM0+nss6DXpfmhegumK9ESTKErkOW5W
w+th0AZyrmXIxAU+LZN2Ex5S7IVtqU4mFwyz7uBPxgnLPsJ7GrCGUewojCmXqXCt
VNA8GwR1nLdHRlwjItlld1RKHVuPdMHYE1eHS1/CP87mhNuCI54ceFOw9TEDZS+A
37RNS7uaChtlJOZLdQrpLoj6llq7pyakyHZeaWpn7i2OkCB6X7IQ+TVgpTJMczR6
9lUIdRPd8mkPBGqyMP4Syv/l+AnKHvm5mG6+Nu4At92s6bxVBmIk+ouY/8JvE3R8
TItw7oNg5Dwu0zQkajdV5H86q1/gqAYx8JoomF0zoUz6Z1yCLGJh8ih8w72SP5v6
gunsWvX4UiYfC1lIrtauwTMTOmdmH6lqUx5R+3lG6IIxeVdVJcpgGUX3tFCWHdh9
WQO+cojQ44j+lhMmZPEij3aooMo3ZeoJl9FE5WcGWqb6Nzvs7BUAHDVMIJF61XNo
fIcksIefoCMkCySw8evTCmm/Rq2BKLG8i0ovu5K8gwCoj9jhAQChs+BZstx3grk6
Dpwm93BkggJokJnJGuPbQgGtRBxlBO+KRk+dwphaY7oBxu8XuXsSbuPJpy/WKvvi
PvMZSCxRalVf8nG+RM6fWrKpx5FBembdYeJMXFbsfpPFzyrsKjZXEoPVX0KOpU0S
TqZjtf6xqIMV6YQxR2BRpQ5ktso820PuB7JGsp0umqCEXbRWRnVIk719M5ohyuhw
1iK2QCi30zwwy8OGKYyvpm4sdS8fkmiXl/LwuZMpyqahAoGQEFuiel0hBLNtI+no
5nwokN8IEkZdoqPyflcF6GDwjxL17qQFwLoS0OLoKCW9aWc1x99UiPW9dpDhjEdI
ZufRIjyDOpVqnYnlpM+t3SnWvakhOwlZp2F6Qv9okPYAKsGKRw9zOlu3knk/waSw
nDmrTVTsDxuFrWpsPQu90V2qIraoXzcuUn/2zAczaKfKyAmPZ5Pj53MvRJkSFf6i
xFbRwxtONAPzPTZPM00AV/HcXfDxV9A0ub5mu3922bEzkrKbZcWK8D5hlYH4fHRs
KL8ETNpO9nDIJnOLpjZOGsyIdzdLNuJldGSDhmU9FDmHgjBGAp44a1diGyv0wXAW
Grl7n8b/ZN8B5EVyAyiD4YwK6mcsSdvtp4dxjMf4Dk3ddT5w1/IYY7mYRQJ1hIm0
Jvdi4L7yb+0T6xG6Hka09PujdaeWT/hPR9YIfYL/cyJ2uArOU+Bd3MugBjwq4wYi
vxWgOGYBcKNeLBFNWhv3kGZ4GMt8yy8ANOKrCH1QVAf3Zgy07ZRy0e3mD8910Ci0
zGzz9QU3nQ4wL7SP7OfHhkF+1wKgBz9Itr8f6LnioP2TUjwMd//K1ZqwtxxorYe6
on1zjkJma90fRqy8fDX5bQoDWOrcwcOeiB+Z0dhlXaWeeplQ1zpVlzDuR64yUfpk
Tmy51YaptWTWxRpir6VgQuBcnLtoVz0R+GT3UfqNdeub5Ue2k2fHHQ0SfF4t107T
xRfohvb40LzohfqsC0yX8uIoVhEv5AVGORdN5uLDSFSB7LdsC2Ho4kwC8Sjwj/hE
u8nHV7dUZYnTTqMfSbx1/ULr6/SQU1VnIVUD2N9yD7UjV/4iui5LCtk9aprmCP2R
6XkUtsof+FgZvdqvseZXwbjQJMS0AjcfITAohVKLZMgtm6KBJKRexmFgLlFFWprw
wjZ4murFTmdeglATskx33GIBkVcmmN6FqqeW6nGYKl2Q/QOmu+tofYjiC5GQypdr
QHsDsCXURz4Znkx1a99MiNydcqycUIhNlOha83n72XkjQTuG+HPnnFO6Ss5LnqGU
3uFWjsJ6FkaA4eHI4nlk8CMSkJ2MhvAYujTzImXHVMcxCTELoNp2G0+ubzd12RSe
bA7puau4ONlQkWePfV21ylrDatWpH+WeOk0PSYGAKFfXPZuTa9vPld3522LnNcp6
ZN4W9r62+djVL39sEGE5DlA/2VRc4+VwvZt1ZBT0juH4sUkFrSfukUGxyV2CCPY3
KtykPwfVVn+u4j+7ZredudXlpAlCjy5JU158kPMaPCyo+goA1/jC3FRuPkP5xzPE
v2SAXXvmueLB4vZ2qjH/ygx0CWZsKcidablytyxzsWgil/8peuN8JAYKlq19h9rE
7FkWNz8jnqTU7n2tJDknS7JHOOjkbX7QBUUKUm1PwIrl/0NC+/J7KBEmES7orH+7
+9XeQfzp52yYeONARBTPnIaNPSLHxeBR7YtUiBLCJ1pL8kdbCE/L6FjfxvOxS51l
L9J+OUJiEFiV/lTWDb49IrOfT/i3aYp4lT++b4hsRvKj3d4le/Xic4VcfEpsuMXO
66zcvagUB0hP1sVRIc4d1aqXr5LmbJSvDDTMcnXGTkUYzVv1UK9PeyKBiVVsKjnc
DNB7q7vb9B6OUpVU+xapWN+vGo78Oqcfl77wHH/Q3RipNd+caQvfigzdM04FBhf8
mUp2vWRyustC7+LmTw0kFztUhwE2f1nUhI/+Jd+VybYMjDhrrtR76+st640rSVnY
FszFMCY1fRRsv8exQbk+ZRihL2aACEHZzA1Ms0KvlopW/4pUL6TOcZmq+OTM2YeR
oGMHpS7Meh33m2yncczLTj80AFRucB5opXIYPsPpYLvxI7YOn1uDcve9uCZuCr0c
Mx70lK1UBg6jnnaDwA2FFUE+YEIe8tsVWb8RIlCYn6nrFHwHNW2rEKW6QwDdbqtK
BaLnA8Nn5i68GgwGG9LkSwZAlNtUH45DEm/kvxR+pv87kkkYjDW1vJfrHgBSP/45
QUzeUzoxZPgOYiRw65l5VriXzkRp1YZiMMe9jlhCHzM4tLCMJyOMbWc/47WlYBUA
XOmQWA+7EtWlCoPGCijd9lIkXCeze/UyajL+zd5gl0waqbfh4RnWOxnN6voxNU4n
zrT8tB7awZvbWPyebDBSlB/aEwltkIqwERib4q5fMsC8IN1ZumsmCZjlT4qjL96c
9EYybp/hhFXXv6d9irPE9PvOKZXBe1TeEu9fHYg0QrN2FliVV1GaDhfSpGhaBBSE
BVAkj9B0EYA/koxhiDxYuSUg8QfCnCySBWX1y9AHvzp6zqGWDMGy7RtOX5qfDdrw
p5T3mZ4gBQ80vz2oGgxiH87rYDJZQ/7RxEQCMUnTljywX99MhAxmxp7/aA5BxtIn
ZqkoYJ0GALTLXyOW9SbWaWc6mcOkshJl+WlEst0nzxTEjpUmU1c7/H30Rx+VaZHr
OxbU/PQty2m/H+cw86FPEDs/V1kX2uQmxk6nqJt5ibXWzGK2y2Pbrs+DO1uU4gWC
r+h5PILfdNXmwDwhSeiyWL4sgumx+JFJGwuqbaLS91sNSt1dbxls1OIvBxW0fjuB
j40vSG0k3R32oUiLXYegSUpB1jzTejh4+0jgGlKEMxeRHlfXsKgJlvIgxvna6sSi
yVEHRYbXNQymGoKJ807X/cQf+13WVYI6ypdvXffoujhsFTIkl5TrOvQeGwRo69+u
3y8pMA1YLtq8vXfp84OjG8NFjLZOJT35+Px3RTQTlLfZYX0wFMszQsJy79O9G114
NpQnWQ8omPi3/56tQSo1Tr6e0UaMsm0sxSPVVrtbUhI8hH22rWvEvwx9K9jSTyE8
iHKMG9bMGOVZ+2hKSgHBrp1mG3U0BAWXDRTszPB9BElaGwjp8FP1rTF3193R5y4U
Wt+auFCB2WdWuux+6284+FErQihg/0aE0R/AK2gmGezFEMsHWAnnwT8XycaESMCl
xy+bTfOUrbeQnqNO5OjCSokL48N3SnBmHbXjZjfT33wzMB0xK2hvzJslu4lRSCQF
Ns+tAXFxnlU8Jn9JXNqdDMcWEc4fXxszRlAC2J0z95jsA1Ww5FLIcxqC04aJJlPk
lLTTie/PU+mMShibAb4qUbpXSgPJ4UzdzDLx7Yv1OFTMOAae3C6M4bCmOMPD8r3N
Tdz/C6XKb+Ade9KSfgnkFxXMdlQ+4O1/oQKcplbruJwcxwHguyCxsKNQResXiFK0
RdnKTN16aeIBP9GbtgmKjKYvpNIhiG/QKFaIu+jf8XnKpsT3qsSofgDnUfeYMslR
QrkpMySBLnCDrsR0Hsa38gdJoWcs/lntQitW76X+jTZsN2y+48OY7QnWnaB/kIHJ
QKjl26KFOmE8c5zAox8AAHyto4sjpOmkI8A9aL1DLzZUJPBTZj7qKz/0q5SCL1u0
MzvOQgeOduz4/bKDXcT5Nww9Oc3CL46sVIxGzW1TK34Rw7dQ5VCqoo0Z+TfNyTWY
2U/lz+Q+81dcU59vM8Lpsv1gsroRzJ8GTT4E4kkUJRrkGbTMBaEo2gJ4ShFUAEcd
IuLIvS9dhi2U0h/G5dZBnwTxIW1bQzZuk8SE8cu7VrBAvkdVKlhxgJX/3W6s9q9/
/lYmB/KRhrfQFAOUjYrfFX0iv69xnVdjo2F2aJuDE2bdlABwzYDmlQtzwtC8LDc6
gSc9VP0RqzL81HFBXauRQrL3p7kzwA6v4HL1hWg8nslxoDkfn1StxKrzZn4t9LS6
HtUHqNA2ESN8YPkNtXtyDDX2+c6eHTfz6BAHKbRrggyqv2gPRuiROOTBnAyGlt2e
e7lJxmAkbcAfFrovj1xHKqhY30p8Ky9a95VbvLAHxZeB1zf9i9SZ5qhU3D+nTDX2
3ZOJVdYtLYfr4WNr3dYhk0qaUy5660cb4TBH6rYii+fR6hQvuNvZCw9XJ+2PFLZG
vbsOndYhp4PIznBNngAfSgy5WdyCzK/8ThymkB7QyPEBoDEJGagQ5ic+Os/8TD9C
kmyo4tYqnmAaMT8s6QBQhz1FxSs6W/Dv64YBeLOj8OcUJHfVIArEh+FKbhXvBY8t
6Q2uxbl4bggPikrVhoPFlQuLOdI5ukHwh6IUqnYyM3fvw0FqNkehtoOhfXSsSKJD
k0+I8FtYh5htLOQHeFtymDp+1lyDWS+lI6VnJ5otiUbmtvIM/2EG//75WCOs3gkX
vFOGJtSI0K91SVaud4jjzDQ19XaK3Sf7W3+6go0AzwIAY+GUCdS6Ba38F1ZeyNMP
gQakc9HPw6/jdCVcB8rSmk+Zz1Fa+pRvl1x6a/IRuX/Q0TyeAjOREVJaL3INuRaO
7WLRS92vu7xbCTPYR6jw2H1y4+CFHxW62GwZg9PPZgpjzzdTF5WS9VJz+Iiyk/S+
Pk63pjc3V+pyKkpM6nwNYc/QJ9NBrT4KaSx6P9LrFHKeVvTkvTkCcHFS/wVJ/14j
uHblSMVX21eDhxA+n9T1SF5+HXC3gMspM+gaC5uXbjH7Omb+MmwdpmU49wvcBFM6
RLC+laSKDIiI12qkOGN0ySmCKwCvpdzQYqsU2eZF4PNtNav8Ngc00AhxkRooH+a0
HZJ33G/27TL1FapIQe9/K3siDJ2s3dwdWHqrf2q6W5b5KL8Wx/q03u6RaKrQd3vc
A9wkgNJbgN9gqEmtF9gpAj77YSs98Tay6I/Z0Xi9kwN/x+ATlzGGER8oImpB9uk4
l2O0BJav+GOtcbzkM9Yh7E1OnmNfgUmIICnpdigYOHVfQ7EVFS8XD3DiameY8UGP
UNEQ+/BWTqX4ExBdsC1ObTR0LdmO/RVa5KmK6SBR1zFNYMcXQRDSF/Rqfz+clkzV
NsnumNrjE6b8OsjF8a8aAybwQE3MdtyA3xfT+W1VZOvpLB4uDpBHrCSwc+NuSTl3
Fd4feUmyAcq6ZUDyO6smmxU8hjmGp+C/fa0iDEwgbUUwJ6X+7jQG+ExgmavBZVYy
SDLQibCQFGJk7TkjA2A2Yscw7ceDGJgsDwnNdD4DEzYWkPIBoJl9KS/ybSInYnPR
bOXKngarytNVQl+B2pJcS+ozF/HG8j45aq0UIrd3pwp200Ah1gUJsNdb9Xm/PPwv
PRsopSgl1/sYmbJY5R7Gh8lcP42cFv5Pzks+IuxvWxPwaW7ClnzEiU7POoTeuh/M
xRPel/7wKoNYYFNIjgSHC5yy+pgJ8/y2VQ5p0Oj+DkzHrUQuVI6lezht5mlsBufi
8F+WlqUBq9oiGZlSTotQd7S9kff1uyoUoG/zGzc1guQDffuCsolgS4r77OuSX0/s
VgYm2MT0lufelyCSVzw4vw869Jyl4Yund/1XLnrcTjSbbRUe2uxkm0FzgRtdUHXa
I8lLASK+tTQh+Y+jkuk0asNiV/6yDvidEdGRY90toov75vy2Q3MFhxAWen34zUgQ
MFJ5Z30tQ3ZtQvZWAf/7yr1I54RpeKacqQuoGVh5K7dx/2jl+UNMBk62LC5/gsyn
uqMF1Ev2UTlLQUbpGnbxctnqRFdy7bXIJ4uX6Ap70LC08na2nO1iFCfO9LGi9jcU
JCTiFibKl89/aYua11V2LiyY+TzeKbgVyWtkx2EVk2nggFhmVQVKLjQrP0zgqLes
lIqOVyVkXyqrvWgTnCJ3EyfHzaF/UAjI+AUO2MDMxmiLsRlIrZcVNXnxhmq83BSm
Gvxpo0iy7HwTlqR1bYYMg38f/TQUkUYEOu73if2HL0+47ckCBfCqbH41j9MMZ0V9
35GWINoYr8/Mq3HDumo75Osyrh4AvDrKXn76ZJiB9OkZswCqRtoN8UQJ9243PgwZ
MqrSansKDQEY7ChgRxPI3FWL4bOD4GnD0+VIlDYFy5jE4EKzyG9Avxhp2msUsxQa
I213XV6N+IFezlnB6hYhM2C+mrJ4C80wAmOU/0Pq/EBswwUV0X+pOY3HLUKADbSX
XnGcu93E8AytH3uR1WznmPGik7qVolvXUTE0FbUoflwUTcJ7HJ4871tTzHmPbF0b
R1MoMUfFK68C3bGT3olBrBWeYsmv3GheeQFESjjhjD5vxSfToGkZLrQkWgLZuIf5
9XAUcPlyLYNVnmY458sZZFduoySV+2vxoqJjbwXN/5A4frV3vrHxPT1nqpK9q/Ut
hn1TQgld/Gnm/k8BJ6RJVfj3bRuDXsggbZaJ3Ub9RKkCZLEOMUOKlKoCuPskvt+X
0qMbQQECsh/U3oonQ+uQCLuh6e6FwpWZ546An5zkTVCwD/0RCfRhbnS6SuNqP4/S
DqPy1sm9lyPfuN21NOPvarDWNaW4w2n/qcYnJJYfu+Nb2n7ePc/mNbcAjqhKcDp7
/eSqyl+ceH7T+0v6eWRlyBsWPaYbr1yuyW2RKqPZhbGREizejGtwR0B9drs7xopV
e820pxwPuEvz/bT8hODaQgbD4y0U/WR0q5UNMIPwgIK04mIWYhHRFzX92wrM/vKj
VsxJWA1UN9GRgHWuPET07f5Dr99dUc8VL/XHWfDHTDVSZjBtEqRDXf/x2cOlGeuh
O7c1sszCWBX5qkYSGTEDMkYYyNvhdiVg+RWCJE5HgEBRwRT8oQpij5ACeP3qFL3a
FBvMl5rzJseIGuWcifF33XII6eeERMlDVnMpCzvWsGW4+l0krMFxD0WmYygIyzxu
MrpFsBF9iXT/KVWLM/34FFoQDp5LQrQaXCe2jEm9eEjooAL8GqqTkJBaZxUnd212
irwsDQBMOQGIS2GJ6Vl8Bvl5VzZHuHQ1G2afbhqx7oyBRHKjkE56zS6v5ZcO7wXg
Udc6dANBsd34CpRxGxFVTTAP7qlpJyMYd0J/NFHjYNq6x1j0A8taKrP4KvDTYBRq
sg/xMXJ2NqYGt3u+exsUhBM46O89WwX8rU3sHbsKAR/pFKjlX3VRFGS/TRQYV0c8
V6Fw+S5OAKwIks0ztURFoEjXvKo8MBEQ+2M/iLGSkvuiIZxCdp2pk58275xcwovz
EwKYek4n/SF2nJmtfb6Nta153HZds+pueG5O8MIWPISqhQ9vS52QBbTabshUx8wl
M24P0vh8H9JCm2rQ4ljPdkstRZi5t+zTuky7Vs4Jjo1vULLWTCzwaxJcAIh1CEVl
TYKRWWUs18QV8IwOcq8Rp+Yzx+e63Av42mlfWWNke1Akxt2FXvG4yRtLDSelyLkF
+rRlDEZ52bDrLH/1hiQlhc9sUbaQ9JmXRU8+Yd9oY+Bb3aiNb5npJMXYQSSR5hYr
AaBmaVWRZlFDzzZ3ei5fwgNVYzAAfaJicBQQFxfg+HVA38lax2EMBHQiI95YVDxi
zs1IIr8Sx1tBR9SDn3gDO5JrTa59TUfGi4eG7Hwqc7a4WoxBDwjt1zcN7P7wF1Ch
nkzTscgaVyp+xuDIk1GroEvHeksIA7pFRFt+DtvkMjyWsoepS/nyDh7dapZvh/An
5AJFkv9SjUYKYWykNbjLP6nwuLWsKjm1eRR41mHc++DdU3ABsU6G8UQg5Gowrd3A
f0H8j+D/ev9TqZwhl0yupg/Gw2Fg6+FDr0gFwiIRKJ9mCIXEoF8eM3zjsLIjukX0
6n5yWZF49FQZ+9b/af8E/JRK2L9JC8L6qptvb3PrbIZJj/+j54LVVKNpMnK2jaAx
YhtpYfwsKndhJwCMJWfIfj09cZ5lxAiV6GnFUArLXM1I3zybt/5t57pOPSeSx+pD
uZPcG38IcQYAPpvnttzbghDW1ORDUabWNxV962VbKVi7qQc+z+Ao8m6z4yNBoZjH
COu1z8ayB0JMT76HOocJG4b2DpTUbTteI0hrm6UtZwyNF2UiC2soNXRDdoeT5g1Q
rAKDcKh7YDAtrGSazB84vyt3Iw2M+yf44U+Wwg/IfkTdZ7WKaE4MALQtQj07k1UB
Rw9rtmmltXb1njoq8kqCesA/Z1cKb0HJkAZ5Eq/ptnLeUKEE14dJfisvDUuFq7x0
AGd0SThAcAcQdvzJQuKMyKKK3WvAOpSDDnCgxxiXOL0RaWr3xl3puONifaszLh9t
A3Z9/q45bimo4antpZHPr23HAODyMGMdmeP0niEUhl4sp/yYIXkzEmI4WILPEuxh
et4W4CdYEoEQCJWMlVcwqoVNwERUxkTFn1wWb+I+BQdpVKUUgRN89XywKAUvNnad
t9NHmOd0FiDXCJEsvxynXo9CbPSRmqZl63V1ihnou65fX3kwSysVBwoyKpDTPB+v
43DiOLXxW3jnB93DnXXBJKO62BlYPv4U5eRvnl6CGR6csZGjiIB3FELWFWAJ27Xk
Js9914WRwL/WkT3z+NR0XJKPUtj3hL8abX6UMHRuNFMOeQwlZYSrFInpe3AjPJ0A
SVcHoj0LHvuOcGi5TjDDfhvdrJBwy9ehFjo3uW1w7JCiehJsj84zvb7eMPCuwINI
AMIR9rInu0sRMx5aPSAROX3Pi05doSgPsa2+IxTnL8gDjZtKwnikBcWi5YuBeCFD
5sZb0+2G5tbGW8g9VKy132X7k/TDqhva1aHKdaBNCv7ZX2dB0NS/LKubQtu2J3zn
5d27eYOFKi/zLaYS4/BeWZyVQbWP+eifFwMxnb9pHzPGJF8YjD9I9dZT2VumUAiW
xTU4HuLKhSDphkJYNmYO5ZqKaxCWKqAlisEyCluc7gEEMe64wFVXQoP5aSED8ukW
yW2yYsdS0YclNfXRkuMze9KyC0rc0EPBOBTw9bGgROgzbZuDHYlt5gOOrkHfoN6A
S6+cfxnqd06ptMtWI6DkQ69QC8y/If5OqO865m93hnVk5/GkAL6ZJp9A38QobnGt
FT6oUesW/VnsPvK8xuHA7QKxcvkGmgzur1wbxG2ZacP6XjWpjRjb70yYw6WobFDF
WlkhCKdaHawOJcPuVu4ANp1I+tDQMaQ5NYwjPpVMdACasGz4mJmzni9zL5B3O7+G
Z4ycPAeW715/7txoJLCPLvGsMlYv7Ep7QZK7nJewFHAdE4jVmztHyEybPv6kmCX2
gACp2ZvEVJJ+tqc/K8zzbxmrk3ojJkRp4WWwJ8nDnC2PnUFzgGl4X5tFvobJAVAX
G3CUc1KHte1vng1jvGLyNdA0FtQ5CTZAO/FsG2JPqKWaIwxDMH/95VCB/9sGkHHF
TWuf1Z+DZvCxsGBHvNKP1aRVPa4qoi5+cKCyjhfqsskC+f1ejcXiPC+QpQLLRCUc
27sDplQ2dbl8l+5UVgOV3WZhzlmG8FtAqNXF2Y9U8YGvkU9Cq2PQz5mMJtavRzc8
mHaOA5kfVJV8RRYe/9/AX77fmpqZYpakf1iXK4KQ4NZBeExocJ4TIqyv06wyYjgl
Njz+73+efeFtmT78VplW+4JHhl9iOjGRA+fiG5bfJm8JL3lQM7dkCR3zKvWk8y7k
wrUGfTMtCi5cWP3HsxKP2AzYHESI9JU8zOVcdcFOglz021XjmD56A7iTX6hADrFy
YYRhV8BSgLbqdUz0PEUG732Ry0gqAtZTvwUfSvNBDR+S8NcWenFC4K+XUP+1xeQn
ZGQlvcoYtcqL1APAnTNtJ5CqoqkIIef1VQmLP/omYZS1xQTNjgJ9t+rQwDUdUnW9
ow9Z0Vsa0tEM80aHNJqk34ptgq+gwbxhHTU8vatgVcGddLlwsM4fxdy0y6ngnAP9
X43qccITC+izb2F3qztBpRsAlsU/j8EbpnhSUhnvy51sIWVXBggFra0BfvUl1YQl
qTEll+XXcC/yLc5Ib5035mH/WbLByLXnFjO5w4L9oDT7h3KqbZkNJCu2WndInK76
5mf80NvfQTVp/5+rEv7m4q8pDllFn49FuTUbUVoofwJYsTSTiuUyQ64c41qKsTjP
EByfsmgW+DkWLBjZjbj9/pNffVxZtW+21Bq6qg/QcSSeqb+fE5ZTlu0XmEWjeIto
HwkhuWhg/IW5gNy867IJuFeOHx4EvGtgw3+g660gDod4EmK9+/pkNFikxU8yYpzv
T6FWDsG/fBhbEjU5cq9BdaMZrkKAQM9iKgGgreOnTZ6rih6y9nSGAYAT2zk0UAMJ
YeVbqLmgBzSPWa+xKzUvdbKgz9A8PTW/ZHjPCHPNS4zhYMXKdyJsZcCypKUb45GE
umjKK3IKxAIx586Z52x4XgMqygvSmMc+Fyxvd5rLxjoTJMNqCLCIcT/uZh5HYBEU
mskb2rr6AwZu14h2mdtOgcsg7ZtQsnRsDR5t9+5SYrTebfHILkzYec7XaDTpDVny
riL9Ztbwu3Fsl/iz2h7ADtsJl3cQ2knrEdCDEXBQ51QnAFI4l3R9hZe46GbUVpxu
wFcgZfjOOqAOdZ08/KN/Sc9uSssgZJNaf7H13/VJrp0pe7p5bJf3z8RX4sj+sKdv
QUOuKSL8zFVsOdqoVL+OXhh3cQyUlL1wOfWy4xXyCM2CFuVIIA0GB/LQ12NOi6OY
GGszRuSboQfWHq7Zr96AaWY+72+7LjhvXDscNv+fuo2w2Gx+86lhgitvPMNJfI5i
nd9SRJ7hN0+zbMd6ph+32UDlbqW4LRRv6VzF9Lyd3+x8sNjstt5FIM2jiTyU8MSp
Pg6isKx6/DlkWX3sPlr3LS5hF937aIans1s5me5EuERk6B99dQNdXVWCIaHroosA
DxzE6hfxleHnUn/NNGNEEQlxdsb7wlXzbLY91fx98W2FJJUf5WSe5NW38/Do/XIk
/xp5lPXiBJ9BRuAElOsK4BW3ddvdA7IpTJBCj8GX1PEinBNf/tbypZ0xHL6saGCs
A6EZb653yKGcsydIMnnA5fxIgTcrQm3X+gnJ1ZHUySFYK8AG0mr27D8sFwcEpHJn
JMf2vSMzwbhdX9NLKnBdMMuSJIG8W1vSINfTTjE0uLAZXxKn0hoe0T4A46pHprOu
q7hF/WU95UoNSPajP3sHqSZN/8nHr7kaNdqk4uOTv1fnJdrEsKz4quWXZxlJkDKb
8p4TLqcgo2oL1cyE+ENKzKEUy0Z7TJ4Nm7Cl5piYLTVUfJnBmdV8vkqtkf6UM/Rb
lu1npbt+N2obGUISMnORhxXMLxWClVeZLTSMhLD+upjgi/81i2spJlzbn1FBfcvr
k40iglRSTv3YtIHYiGIp2sq01k2n3RmA/GD3Cimu2g178vt4WP9zoHhTUsC+OaGr
933dRYcEnxg1HJk4Bz6vHix6tAQ+05iBCeTxyY5NjrUpIqii2G28hx6WTf7tlUXb
/ktighM9Y2LUTbIEACgkEtItw+6HlO2sRWBZ1vcvBK+YRIrQ28m5QdTRt46U0elS
bf8OcAOqT1WhvivXNWrPkOr6iHl9sWYS1KlqX2jdRnqEEXY5simQv5YAWyy7pBwu
8Wbd1tQ4BAPg4Wk4o0fXYCS/iil9y8kvIxtkIyQrtocbvT2qeWR7oj2VLT3uvC29
OBZXxrDxBytWrV1CjurLLiY+k2ckgCJ3AiIzUgjRKafPbOnBk1ICOmFdRqrxtXc/
40RizzzJ+37QMxV2igLBNEuBaZu2/+vQw4orhzXJyEFk87f9lLZKK8hw5im4TzL/
hpAFRbE6nyvdGc9ZvfuLlafn68A7A7nV/JeUDnoV0rT8tODGITGqj5lykDNbWExy
JCC9k1M4X00sAlF8O/iET3o3ANkbfGyD1nr7p/zrHSEo7s4t+PkhVjp9DYsmXgUu
THlnm220YCx9GVuUu8wMIM+gHjgiAHnM3//xOCgkqsjlGoNtN5S3C6YOfGxpQ0Pe
TgG2TBYBwEs6ZteRmz/E5MkcOWpm27wNQuue2CirfDG+AFlrF33uO7gPbsvYq8gM
Is58mkUe11YHCx1PqldfbLDgvkFOrJHJX1+0ARGHCOpOEM5JPAA0i8E+19rMKo/k
tGQXLetQnt5x/jMwQEIoE9e70xLQfSfcFm16GrdwGqWvurqmxpkM9GSMdqwIvSqQ
tssm5rq8Az4kvE0ldIWBgA/gle+7HUfY2QYHiwPTMok213uXjPGvXz+2sx2VcXqJ
vGV6nn0mBgtG1uEtTgj0TdZj5IhLAcBfGR4cbwQvH96WqkZtJEdiNViMk5pjXLUY
mwBPdTn8z27KqjROBTFKna3nZWiDBZus7v9d1SQwH6N15DHDtmAwkLy0GSJ1Eius
f+etq+CPhN1CWTEFQY3hf6FNSIp1TdEkYV6wiEUAtTnHVyun02N8sCW8KzeHx2P9
EMR83JBTpDHCguXq3jLXejNwmAm52LlM5HQMnsR/nTo8AcXTS9qhIO2lJCE+DdMg
KbgQd5ji+X5EsR6tTyjU3GbDnxpSx57GHIBZIYHeyDjtfxaZYtUDatdpIgd5x7Z8
LT6lu1089P6v5sDKTYiP+2KPZS7vRihYarxFeWT8aNdSFuceljgORXvIm0+LUA77
w7UTvwI8YQLhOsAZU/JcvUF0rQ7oR6iuWnDWlBAqYuSY6QpXOsyeI+swMDt/Lgkl
Mym5yKIOvi8C1kNE/RlPz4LuWQ+nJDt1BK+la3Q+pQt2XSHzxsls+9f9uyYIf2Tq
S4dAr5mfZPljEhBteWhWLorTdVulnwLrKSAd/lTEzIYdUdu3vDadLOIhckXZPRhS
Xl6NQe4I9sciwFRQCRmlhhzU3VGFpNibBGjP3P1ZuvtHUg/QPwlEcMV2e+pLCFPA
10Fwtjj+s/0t09CU//6yl1lzvt+dVsWn4ChR9a5xEUOiWQfIsr9MBIzsh5cYGSBO
0sdEY57pl8YTBokVOvWcKpfcvwfT+IKIAIDCIGJcV2LXWk4cebTGC86lFO/xwye1
/PILlTcy27/O9va3RfQdT2lGhUFeZl4dN6ODQxEnk0kHrMgOlxCN8XQ1N1UxEsZg
50dHxdyT5cs0gZNcAvP9AukUzaRndCAo1lK3NMvKtMVsEQZ/h0fI+yrSVy5KgVM2
cU+k8sk70pFAJkZ0R+8kNVgx+XPbwas6vjO64GLuU54db35KXSodyBwEauupIdCG
k1zG0I+mETb2HBknLriwmI35vk79w+zosGM6TfHxTm/h00dwpS/WUYMYFQtbeous
Njgxk5yLvCTkkshz9+Entlq26FeEn1Vs3L5nhm0u845DVDxPgML2jIhAgSop1G+j
zte7rxuPJ8W9blYBaY0NHRo+vUljWqp+DmcAXnqxSLB2SU0mjBlMpJRgGo94aCHO
C2XqsjcFO7I9keI4YLryms27ntMvZgwo3x7KQ8FGsT+atRfr0EWj9nTp7qLN6nDu
yr6TYH514VIJxcnsuCFQ8o7oqqs1XwCoBMOoYomKJu/BvYeG23NGPYmg6B19SZJ6
6F3e7MWEsiTOtEjVFgVc61TPFfv8Y0eYeGOoMjWJOAQK445w0nIpoyFO2+GDREtP
UNceGzecVmVsRyvds9urHy6ZhrZwwuSjHK3LtEk49+9tgmvXNgAWM7zVRJ2ButdF
MxLF0evryd3xOYtWZPi6MFVASPqWeAhJwcB01MEWp75ICFK5n/2RYLEhB7a+N7UD
t16eYBQaXvOAGxzPSjSl7s9eLd2czeXBokw5fXTYr+xe0XpWquM7B2U9NGdUTSLv
Tk6VOi7p3FL+SJGO6jfAlTxrMhPAaPktUWSUvTSvcxiK6VMMZJvw3OAfzd54B1rj
Ooh/cGxbV4bpEmsqeKWYTdCuoFm7ACaaOGy/3G671/aYjQkOeonzpVOstZgDLROB
TMF1OUnBZk5IyNkOzL+MaAZm0jt3WadHWAcaD/0DInjz7wddwWX+0FfFIR2Eyzp9
s/uiBlB8Z/bIw6JmQNp5xC2T2D4T5zkV+0B9rGJLmOFeCAs3AbAKoVr8pAbW2pGd
I1iyI2OEUlUQkXCJwm1ND63Ab4l40sdoXWgVkoEUaWG9S0Vdd63kTCQ4rEJ+j2n7
+jinw69CxAqzdQxxFxWcEx1++360CrVAeWEWjduPKlr7JjyqLR/fIvFjV7VH8jTp
VhJkEvuu6wwH6njjihr+kyoY3VSA9k+k4zYcx9lUn7faaeuI7K7zcFkQ+rdtzuqA
TkoF9s06At1pjJCAe1rmFzmQn9fndYPIkkQ+mbPnQ31xEuecdSBV2m8R+CfmV3M+
G/rFqspGQO6jGgA4SL0kulKQ6dRqGZLl8qATIKn9YojxUTsVQ/Akz8iHd46MjUcS
NlX2E2omfAeMBhS4o/n+jxBIWTO2yKq9Pk5pn8j+04DbIU+Tp8G9Dkof45CHnI8U
i5rLZ+FDk1gnXOQHZ44vz/MYhwmP86uqo+7vyfFGJPZhbvNKlfNuqSUeEWmiwM9b
u0egMiKpEMt6x5lQHq1fqf3mah9PVMYgUd7ltJ4aawDDeenFLrfv9D0hQ7iPjLpd
A39nkv9uSB2oWkxLy2/dXHwiFrEJmcnxyK9R3464eaoi6XJeeTP437+KmbIm4dow
WBj4QbAWS2ttPKQW9RmNwuLmHkzt5VBddbqH5vcnhHBjz01f37XjCfjAMR3bmNK0
TzNDD5wefM5jofdloah80JBWe3FKymSqWFWsP1n8CrpHrh2OYBY51CBKrQX3lR1Y
crv83dSSBNdK3g/BjEuBrqh7Vg8gaPBu+9grJlEmApnxwwv2pzmxapG/X19t7O5p
huEaSF9aQ49F72UiHGyIUtMSVd/8VD5CeVY4iXNTTWLrpdBi+bIX8dlwP31X9aCg
G7det6AfigtNRA2NFQwTO5fcThxbaHspPyziU+CbQ+luewNrRHmmQZuhgIyAaSjE
YqTix0ugrKhSeiXHemLhhSxMHAapMRelzAaE9oRkpgUuN9/I/WLxIowinIoS9I0G
jhqHwzHIaVZJLmOFEqRF8KKx5nEtFOenNGaEvIZlFjJH1velfMTYdgWwv+E1Dqyr
lZEP3OJdxNLQFBQJtLa30sL6ZBMj090++Q9VUVy7xvIT15/yVFJsTp75Yi+7r2T4
kejeQRbh+kqA0/L+Zep4q1yjh4/GrEEHYusus9fUQPi2kNWYb0i0bsornBiVK6DB
9jsbOeYxQKd6ygGJF5q0tDMwVmJBrt7KIwZLzor1ceiCogNoAk/8plDey/h0m4+e
5O9YHjlYVAc9gZX8mFrbrEngxeaY84pKWItKYwqf6w0Z/Nqfm5kaQXfhhii1A4t0
qXnz/dclHcmtKZwVQu4mweJfrDUA6DdSCGGqM0h9Y8vtU5NjUUgNWaFAUBqVClwt
/vqvz0uFwztudAPytgv496n/y4xDplVdDBNmXjzk8RGpmgw6vuWsn/d+t4Plw+0u
RRj+exg2CmGgVTo8XIOJP5L8DwDNimnYu2dGN6suovJKkOTo6oIEJVSQScKyekZ2
42QVXVvqY2JiWOwhDndtvL0/koF5aVUfZvbUvzH5cuEuzZJivbQjzxFkNTnUxCQK
kkqcPYcec97aE0z/ojhdvQ5Uncw51L5c3lcUwsNN2c/OH1WI28zH4wUTyIKNCZUt
UkM+7lxlbhKH4N2KekWMiEz9z1+PVpMrQIgOEtEBO6irrA/ZH/3KOWYQoSHdGqSj
itYi9tI21yySZy3bkwJzFwaZWmmF/vbjKqnzBP3tb1Q3gxSMvXJn6d8XhFCzOj+G
V6lwJyg6kl78sORZ1WtVsqPI6EDyv+2b1QUON35AtIXKSFbZ2+fXCrOS0pbUNSrk
zCSfFQTnu9961AcDmLveN0kd64BTcP0FWIIJw0iXN7+YHBo4LVX7N0mand3cOFva
8KQJ4zlVoWbsTF9cKft4dZ+TEn5eE35kx5kLv2QW0GtjUCHi/EHOjKYRHc8Ncs4d
f8v2twRtLsdZenxUrVecqhpf2IlUqaCl24tTElPshLYWuHPEG9jr2gmj1fyLz5zU
83vbnotiQ8FF1gTijGPC1TmtY3ZsQnJdYMlMld9J/S5ZMzgLd5Fdu62Vjm4zTckt
fNYb/iHrjDn8wNH3UA50Nj/4A7UDukK60wx/AO5eSELxvkulf+yxt36Apk2FGTWH
t30JIz2IfJzxH9XmzFrtHNyuyzDEqKyM4ga2+Iw4mif9Lyobu08ZuXmAkhlDNw+h
jNzwNR6hVxevTMnMf4s/RvoDPYi061DrfmBCdKD76B7NgU6TpRN75nSfVLyh62Ut
HGScw+GK8+N/cmMvM1zabHC3Dee4FDckHFxdkV3cOZEKbl4dayHHGeK8av0WzeNB
OdZPjbOhonJBYjnc/wfx9My2JPU7bhTTHg9qmUoRWmFWriCChcl2j8VI1b5nJkIP
xASxw0X4uPMFhPWmLGa86dkT3EbkcH553KLVOgrvyyTpfs2hMKUTa2xbX8BBKbvd
n8wcwm4vmgec3GrMUNWtqdlB+pUw8D4dwhHMWorm3808mofhNytf3S5bj/jAN6H4
FMBjOqNzHYcdbsfw7xx4fu/9KInpXQYUDUQK7LdEO0hSM9WIb/l6nyBQ7h99O0zr
x0gLULn2przr6tz3s3wUvAx2p9Zoz76lxpq22az4xkND60Sje8LGf4pK4F1n3VKm
KNu5WsQfTJ7iGUdoTXQ691HuL2k7dxQDpJuScsY7M1WIY3G7aBVwtrcWICe+BNPe
n4wWcLhqOvvph2KXwZ4c28CBTWs/nseu3IdO4XOKz5kROj0HItLn7iuXgzl+JD3K
L9kN8aTDG+24exDSV13chy1770oEzKZ3IJYZjQIY7djex6P+6multe2MBJlkk1+S
0VKeG8ecPsnjSYijRCQffekYdhg4okth5IvMbf34VWs0HnofwVHcf2vroDSnfeff
P6ePY4vGUrvvc8WrsHYriVY0ngun5l+NLb9L8orfsgAg5Ep48f2EHJXx6ePC8J//
wsEUeTxj47Ah/MQsMYdj07eqJzRw5yWE0mDbVSNCmzww8Ibhn7Jh7TXylB724vad
z2aTsph3g8nFXOzAY1SVjjW5VvNLOPIKVneipr5MYvDm+4J7mWWGZEkY6wBjDeHz
0U6PxZg8RDovRnQ4Kt9Jln8Zr2VIp6BW5OiDDzVTP6lJkvUMARJRfdV6kWBqfgys
qPRNoY2Njfd7ehjM8gqlqKXcuWUs+dVkx5G3Rvf/mxCKmfs2WJPiRbxcDjJLv/8X
PtdysM4T7U6RjlWVbVZ7IfjD7YT1qsDhhdMZfRv1tbXVWky1Mw2oeHdJr0pkVnji
pj48NDVGOdXrmuaW7RASCv9K7IGqa2KI99+pvUzWy/2oTGc+DizMBgmMUlQF3bA/
aWSeoXQYRvobPdWdnxkitkbkDiYgw7hu+bEtFopjqf9NbCGtM2EBh/s3NGpHapyN
U+qsEJVT2qZVuC/Bvudo7uhuAhjlwhgLK/uPFzC0w/nd4zmpw+Xgz53yJoxdSAqK
SRhhZysb0T9RdEd+zLfuVzVhmgBc1/TNDdpSNggWHQ2dcNghq6kjfbRVG3LhY6Ey
w+H5woiFk24O5DLOPgWX97BNZeX68NONIrjVPBFsXIsSi/WYxTiy2a/UVkPgq2Ug
Rr8yfVOZroQbZG3XFNMcpx62ZeKVh9xT3yhLF5D4eaIdyPFLiikmDJni4OCFHSod
4PBWyW4/UL1WJlrv8wTHtDd0j38SfGiVqvBxmKE+6CGWZjsxAsIx4IIu7tD94rUj
UGZ2wTdDDmwNGdA64BEgJQXmYJk04/5NT5CIG0IRH2oFFgHajf3Svy1lZMssP506
yFCtf54YZTja290B35Qp3RCbL7C8sMNQr+vUM0uLyXA9OrMrPXsWtDSEMuinx3Xl
pq661bdb6duSbRvXqYaHKQDGDzT0rTY4++X6yYrmohnpvvDVd+DLxyx7jHZUdjHr
+9Yx0lIJ/wiXtLtmC7mHuJ8ooANmpzkO17iJjjC+y9N43nN0CKnULFpOLDPIcTuI
wXw3aNTjuPMUqObLCYxNLd04s23CzguaBUMCFL77EzxsVV1GtI3iEAMqFr3fVTmr
M2p+/8KTxv+ha7GsaWYTkdIYLnPBlUWLncGUreXeoJyofkJGB+tQSMwjKjkGkU/u
xbk4NYTCJwtNQV8jX2ISgPOYw1eDKUfKf0vy6oDZAB3KdOfwRIwhVKCaWdPxZtk+
R89Stdkp1hiY745ZHATSvOwFMcY6fJyGadRU4S18eVEaLbiZ01izJqrYFK4LG8GE
0xJK5uNSs+TyBndBliCMbp0JmPf7gHM2Tv8bgRlINYbJXHrk9WQ81UyblCy2rtHe
Vq0JGzZsiiSESIzrfUE1f8vy7tuq3qTawYX8MTluWNFcOXPQjeWX3KhIcoMn8IZA
0l1LHFsiZG7vnUsfDPftf+rei/TDhnrqJew9lF35k66SaoxocbAyjF/iwrXpuawH
A8tutyOmBXqv+eyadigRAvA2lbgpKlbJ/fF8QBGY4JW42tQYYqfWJtP50EkeLG8S
ZqwHsoxUrStgQ5nLf/Mxzk3EHQ5KJVi/3yycgiLRb7Q8xBEC9Qf25L51Y/E6IpJI
5la5wTNYobd09sOJPy7g8CCqdY0cFixJ8OfwVguJ7No46FoBsOHRt4/5eBFzl58R
kfItICoifSvZepzHgmAuKj0UMQ1doF0ybg66XRqCCwl0hW/l+WDD1hOezl1AOoX3
q+2X4rbn5je0qih17A5uWMv63UGP3VXaQKWpSadH0osd2xjJA8vYJ0zcdMgXcRvl
HhO44UVzoSMvRu5GqXRQvREmgBO7kmgHrX1fu54jQzfR3nSAKX6xXJOJ47uuIfGB
Hsyt6fHuMzHyeYMy78R2zmGp3YW08XgAYAAf95oeo0ZlV06a0kf38/YslXT2yp8w
f0HkjZm+2E/7tBPLf3Lz+cHCS+ZsPWJlS6zJKYbjk2StS9VZIXpXjHV8HSfqAQ7O
zmtz9YyQiRe3BtWQxf6WsSO8mXZTLcNfWk/T/lbmX77+wuiCUh8/Qaydeg3Yk9Fl
BqwacmZi9G0SGdRA4hGrk45aTiZ91t3jH++EvuyIQbwFNgCuWI2KAmyxG0oxg0D9
8Jd5/74qWVGqhUkJV/Z+XgLDI59lNIN4wnC0eE4Y95aomhDjgInyG0OvRnjujCCc
wrsf1fzRdGJCFq7zp36FxYEuGaWbU2O4+cWE7sjrgL7tqnJq6dflAPuXavYrl9gV
9+ViyFvuXLHdrrh2eB35pn4uT0Ds9R2IrzROu5ITHx1VTQcebX+fTNNNiWefEb2v
UsJAcmfA7AwLED6VuaXA8xfHyLkUjZ//7rQrvgmcE+u2xqGj7TsyAkcZFexQYnc7
4xwhetaZksjEP+qFu87P1wZe9ltvU05DGUSVsgBz263FumxZnF1kk0CmfMPIJQg5
yAoiOYkoekNT58ayhvXyoki25v3b4cmnPwfMpMO7TNS/tLZqP6krYSriqEJqhIXB
x2S0NLqZI8682KSM69ADFnoV5GbawUsQBuHqmiVOyzRajKzKagmcWuRMjZdLGxDw
l9WyoSyJy6LeEfHeCNFF3eHMSW4Mxmn/cwanQkSYueKQ7rfLPyM+2htPnGEZEg8O
Tw55JKyidHCF/Pp31bRlIs95jGlfA8bjuVJZQlJTNNnNODSNyfXGyhLURh74HJOZ
2c9JuUc4dMhFwI47qR/gtwQqG4TGT4XpJWrrFlK2ZIQcA/zY/89qb8Uz9EzhcCgf
d6pyxf69lO6PjMJklJGD/4EvXi8zpugpSpbqxtDd+WGQSu90nMYniOQxsO5+WtB9
F5W6A0Oo/h5xuQh5VcsS225k0fkKLfXpM+9fGBmtB0HuoRoAaj1PwC3P+630VG3t
+PZoxVVwQ9U3OSGia9CXggHmKjy5XHJ6JuuvoSW7MloC8JRTjjyAidEJbHZcFbl3
PjoVUTeK/3yOVZkWa5LpC0OlHG8vaIqenHmoqJIXW8CGuIUYrJEZhN675hJWgFf/
7Tw0PwtYu0uF8RsqKli26zov6C9Z62abGReofuaWHYtEh5NBw36FRi9Xzxt8bbjn
BrltrtQZzeW6fKV1+F/y08CvIwCLr3jC3t00Gjh9f2HAZvBsbA1+g8Q785p8aKr3
BydZyoXfn5rnd6sR3wSsdVfuWWTXWx118cg0M4Kex5yRF8on6pdgb1XckI0nNffP
KADC1qqWu26d2UPEUDN9JuTLyurGPBKu4CMSR6y9aC0mpfSh7nyZ/984TOkCNipV
ghHAInUs1ENG5mk81D43glqI5uo9e60/rWu8nwlDyu43r2ne5pX2bZWZdaO+dwow
nOLDjWizDKQMYZgsbWBhWOnPCTt62Tb4EbVI2tFYgW6C/H1qjnztpK1vHzqw38Lp
wU3uf6br8++7vuVfWo6ckXrNTZwhh+Jncs3cNgRV93+IY/7mqv1CoL6uI9zD5CqA
OnwOoaY41Mk6UPNRcp3xhzk5kl6lhTy6WGA1AbsOU80emse8tnFqSCFxYv+AnMqO
HsngbtNtt1jHK5hiEKd8iOFplJv//c+DjAW7jg+5WJsanJP9kRDJssqaQ3aUhRw/
gBlbbrpH+wBxjjcD0bcFBW1AsruqZamI+/reeUqaUhzT1B9SKafOdLFUJBccRaO0
KyZWtYInilZ9+LFWWFvO6mw94TgF4/+XG45OKhy6VqeU2q2o1Px7Cg0DmXxhhcbO
XtoqxnMjRdRYPU8UQ1T37zQ6Ab5sI0pwgS1raPxGJQBYjvSBSe1696N8Ut3WlJw3
wPPGtoHUi9W7sgjFQ3mvnaEJZW6i8+ttIExJLPJipKsSdjXR21CpNonA9HJraJSS
bUEZD9EQoHH4Qy3w8bUuoxOth73NlT1Gr1vUoD1MMNH/M6ZsYta9MavWV1Lt3isu
K5hpfRFbzjB3Xg5syXCia47dVf0duauFZagb7QQc83WpzdYHzv/5qLrSesm7te5e
wKFyP3hpmDVps54bkUtH1R4ajqnUOUhgsuHVPAoRs08Dhnt1d1YF5qXO2lFxM4sV
072vU7uHq2dlilnSC5WzeZHd8h2dysSBzzpIrt0SUoDNe0VKbzjRkW8V2PmCHmaV
3X+Wu2aY61keZsP2oy/9RW5SPp3830nsHJK0naxXSDuCo1dPJOmbs9UOBnyrmiVs
UXzasRkJGx/MXCptxtXRPuYYzb0GWm1kyrysh00w/1Ojr2vlhQtkSym+tnyJLRhc
7TGb+DKYKx1cl8ELJYKphHp/osxaL8cZeIs7Hh7FopMo00h7cI1ITxnBKkGfkGaY
0lIUdCGDCIvhtf+Tvk6QF5LyFz/lpIikpMEYEYxFKxEoBZzXt1TlACikS6ARpJFw
baMfqBeuMR2ADeJy6jc46AI3BUp/8gQG5Hs2XOOxe2AXKzIHgXbrYw0VJEkC0IMn
mC68xXfW2Redsw5O4z48RQ0lqnT4MXAJ5Ek00mH3kIE0TvtF9yCfN+jMDNn74c+o
jvWxxYdB7s6XZlm2pBQ1yfydHhC8qLc0MFAa6QkR08L8pWaeQh4pUoiY2sn8Hfsr
ekKUhfo+p7Xo9/UjEGp9aIysv/2/7GHofLVaVuEgnDLsBzXUzIaSjb+UjTvy/FAo
KA3bpWmk66ocKRci4Nif1JcK6tWEEW+3ENnu3pivOmetzUsf5Ei+i6B0gbqIJ3u+
ZH2TBAReAsqbEYDZxEq13Y2OGUU0YGiySpHbcQNd9Bf7/49ujietBozFa3NDWNcu
IYh21Qb+wiJzL/X6AiqKJSGAfrP8YEiw3aLXSVT8T6UDGLyDlA1sjDMAuvvaIwu4
+5igpbVnMHY16sntMBzncl+YTMGOS6FvBZCAi1Sat1kZYYRbZua7+/zYhNnQVGeJ
Nw5DIsteWLIN14SN11omCHSTlHEuqNaVBY2xE9ncGZ3mU8c+TeGrPfE6V75m4Ram
HAQ93LbAR3ymAv8ePt2D+Se795JC0gGBbDjviQvttjL4aR5qu/ihxIuM5xT34k4F
XUX6OerOXVzPZCQJq7AtSxmIjVO3j7WQkvkYLYo1e/A9ph3Em37NTKzaRaNygY8l
JTYWM+Z0qQTL1/wmlu+7skca/lmjUC0tynolzOTZEfha2IwSE6gxm3NSv73PfDFq
ILfQWNSzvuvmqaJjTKNluc7N1z17DgxIBkTQ8Eq2iPCKjamJXPI5V9RYhw2zNxCq
FDrA02Z+EefPREVRvC6pHgjkcNsZhxkE/5YakkFPFLykzSHByZ/Qq4BV9OvuZZXv
4xYrgeUh46HJPl9qZNZ3l2n6IlqYseGxvwG5if97sOS38J1HHui5OiCuyBa3VFq+
gzwFK5lR+C5TUSNYtyE883Nj0LLoYdx+5PvRV8+WeJqWPoOclPq3XfI4Aw9lR7kv
QWc+gFpnVUiPofP4YZKMUani5usifnFBckwIT4m7gxQayvY8m8TOUPZKUKh1gxkQ
CrJ/xBruEjCV5l9JZWe7LLM0ihQ59cUAkZoSoq8btLqyd4rf41bWQU1tmmKZ8bHc
EkscpIQTJM0LEeqv1077lZkWUpKSkyNlU+H9aPorDw1NITVJbu5B2secyN2qtRU6
GUN+BGBpS0+2leH4DKc9AJymbDDbo/q2t4QDCflO4dqFsWLKDYnLbz06dcYYEGUU
ea+7pGKG6+qa+aF6r45DACDMr0asU8ydQMm0YWFWHb52pTVEmwE5bWSi3Pnca2hr
olJTNPJBGjbmxGXYaAEDacpfUV0p2nb0kYpuZFevYMwdOJ1U0WP9LQ+Y9uTLCE9Z
GqqN0XfZgiP2DNiyquL69a1FRoVzwqdwRwbhfuktIpgn990PGvxfEP/tv1DP/xGE
AHzv2I7TZ1UKsb/6+5OL+s6D/AO2PteyjPQeaZCnxEisP4Or/GZW60f+39Jn40ix
VBekkL/DMRmV7bGvWJI7pL/tfQBKituEjsFlhVUfWMHbN95h6BmLhzLWQEiU1VCj
G5KRP+czzW+2Wyh3MnFDj9+gaE0x2OpETBnxBxT6wvQdueYFz+7ixGcNrHSg0APv
4E0fd4Vzi33cGgsJuiD/5zchnM4OMyhSdZPQsXZJvsbOPSBnezGXDRP3rWfcRCwO
yb8mswoR+pHYJudQ7QqLFTYPO2ahH/IaKzA+lZqt5pJlm0eEFTrSQKeTQdbyco5r
rmYXebBRec+ytsckTMlZZDx/9rGNlL+3r0Ew0jYMRBCFY/IgRbC6xV8EDJFWBEg9
uvsuHGW+ZSrQasH27XjX4hDQS2m12OoiNn98ImUqMBHuOcTdklDWt7jeyz9IcqoY
Nt6FIaZ3gV7EvZF+RfJhwX+exyrZD2a3/oE4IakD6txbi4mov0kNcCOlqthlHv22
z6nn2XUd6GGiYZITJvnlCvPMt23wXDZ7WG8Dg7BWrIPqZ4QYrybWkNXOAzbH6F70
zCwITKMU0Sh5hV4UCm+10ChFDx3hPq3cRgY+Uyz24hHMzzFcxGB6UI8+Mp9ZjTtf
Xxu2ZFVAoNAJsq0MdABekjn/sjccjCwS2Q8iz2sTZIHMyEeh6a4Yzeg8JmWxsWYu
n1BquTPO3/outHHf7Sa0VeNFeCHOG7qvzmclPeYzKpuaurKGH17+43Or7X0GRg+/
zBnoJFUlvFGmva2AAsPuzFY5sFl/Iais01JW7pxxtfZiC2WcYBfyohV9fAfKRGhE
5RrAJhphf431MUCFAAI0pnVTtKaLs9H67ZG5z8w/+DZ2XeIH3I0+eHtuT0/QtsZE
FU8KB7WTKbMKodSvD46SeRsc8qEbVGIsYVuhQhOqQOxiTS8R/+5upEKsbnDllF3j
YqtfuXZxsrQhEbvucpwLqdR0bxtwhkuAMo5syM0SyZV/T/PMnhnkfIiXasMV9db7
vOJgtQ3K+qv9LywZkTtKrWgnF8JBnNxhxvm5zymw47rsQ3Yii2vwqKwPGuIKqUmx
i4hCBYUScsvnB/Id1nrUH3B6DbVYnUyfnHXfL7sn+oQOXfPLP7ZPHxPdVhnmL693
oUf/8nexWr7q4r5ACrLZ7HsifpLjPflbYavhiD7FUU8tJmLgd64cqA6Erq+LYWtL
jATGeAxS/l+n5SnGEJ9yTUoXUiIsS9i8ldd3wUf5Kp0h0MJu5/hhGofroBiXo4YP
QGlaujPAmTuKjf6Yl888rC+Rs2j1bfsYKHOiG4xwr/IaU+k01FclbxEp6vAILtrP
UF1dd8BAE6IbcBWwFfaAnnkZd+xoM4shdzsdEGJnSAZcBmJ4yFOn7nnXJgRFx+sM
kL2I0ms7J41QKwJdn90fAMFLAZkK4djFq2nGPPiwIou8vpm3yN3L4pfjMnqaJ4Jd
0pBKrFgFrHWA2IpmAdR4PfV+VlJY4kkvoAoojrKAMRY2ZEN7pNnJvOvYW9ne8hMA
cfzZf2IpteaSFvSQlIjaSxN9Xy2OyCJj9kf+m7WSCmwwSC9HeXTYM0XD9jklozT5
qrmm51/8/l/82aZn0J0EhoTDXDVK8QP5UFZsNALAulCS2WdKLoYxKYRWslH4BysW
DMeU5UXPFJ9NKhTD8LEbWhtWaWUJQ+1L3pDiFtR/32FoeLRWR4Q+TDogOiXme7sY
UbNkiB+54+a+BFvrmnCkOkkkPo4okuwSv8rIYnyfeSQZ3OzFic7pMZfBe7PKMZNH
w2twGz0ufw3Ry3Uc3LMGHTnI3rTxfLYorijGY4FjQ0Kpcuzho8ZQ+vDj+MKEIy3Y
K1z/GLBbnxN5JeOjrEnGIt6aUS/XhQz3rjBOQKEmHmlFZXhG2jc1aS//ltvEsOGK
cTMDU+WAq53DOqriuxeMH+EySQV3tfSFkwKQon2aathGXYdhMp55yzDOeC1c9XEE
X4VHtmVkfQ63TdNr3crpA/V8OGaiI/tb3pPDoHhFKX3hUGXqS9ZE403XR3SBfJAY
UXpOA8/UeUCGMGilq9Zcd/MwSM/rmxHNv1coOOzK6YwO74ULY8wgkF0NRNjImn94
vqqx94L/N5dSiVykpq9Icyd9HqRv7HmmnCKN4YKonoAvUHkUB4yCJIYrtzLgkZE9
pTHocAHvB7f3jbXzux5YdvKX0+3fB2DsOjaqcOl8X91Oc6cOT6H6t3/9SSXfIGBX
ZnlHS+H0CjLCfTGV+B/rz/LyxMTkZPYKbAzfzdqkUirIWrkLOxNMUO0HwLv+GTQb
I5GRWmZpIfCXwTGgh8yFy/MHzU2E6UmK+j/Jw0Bt1YO+f26OZV//3F703dDEZ9nu
1bx6OHxWjGyYmsx5Sm5PwxzoJzY5DCOyU73hqbsT5LdhgP+YoO9+ktV5xaeWq5T/
cGBEfrQdBYc+GkiLEOP6IgRRL5ab2e/YUK82nhP7bFq9swCSOPeBz7HKoma0s8Zw
QW/2BjabvqVZ5boMfdj/RCTgcOdoO2clKU5Z32bz3+BOwbVVP1k8qaQq2yLQ/G0U
62Hn2WDiLg41pcrLvVyoGhHtLJux8dLw/ED1tAJi6lfmbm5JCIes9h8uIhYQzyp6
meTkccE/Ej9sONfNetM9oYVRCbBX3oc1hSNvpDg6mafuCtQoIfAaIvbvXe1TRRpa
tH3xqFMRzEN6ExOx5wYb7WpUXUpyGnqCqR7Qsugol+Z7qgnm9HaT1u6GrH78GUO1
oWJfxpYx4AyRSuPNVA8+DB7kikY1wbPwr8BOoaT1wbDnKp0bP4c8AbUlgrgUI8Gk
JW5eMU8l8wnKiolUXjfOhUUoUliCm+sYZ1VgyRgtjxFn5T+MxHAC9Mfc9xAv8fOD
aq355iT8pCUYUz/NJ3Rprnp3OvlcQS260xkLSl6d3UOGsLXCnYeHhEYGJfoMjf+e
2YfLWSuLc4igMJiKEY4MtZbUSURq+jI1v017ln7JqVl5tENnz82Tug5a4B4ntW9Q
PNzFdycR8qM2noFuZXKoD51Q0N6GDp67XgdpF15Zj9xpb+GkGNhGgJYHevbJy5Y3
xREIRkyFzxIY4faYbUieptXaf+9xjEZ5fT11YfPYttXQvvmhjhSEUFkakikAlKRh
aTumeKB1kda+KJ1sGtieCN/Djfeq2gDO3IeFVFuwqdB+1V5F28zoRAZ80yLQPcfK
tfOlqPaLngRQLNZMuZeGgiuX06Pj9wf7GG6/3tiAAFVT0PYLMQiLmqTdv7GAJuGj
ehF5GXjNzDMeY8jwjgfHRDGsxOIqzjSz1pDp/xe3RtskoNv3guUQoNcQzovNL14f
3/YkOA0fGHM7bVuiZ33qw/APRkOtndn0PooAUp/cWOUsKHUWDMa2xjEbeBaTRWJf
OyNVZ7yBACCtM81QnzFA3oNhj3BhncuVa9ExgQxL8yU7HhVlmkoFqCB8jH/X0Mvx
dBrY5SDXUBvWG1dv2VkYBEXk0hrXwAsrbRQpzfHQCOJMmqW/3AUMnavbHz670yEA
nyurIN1j0vNvbi+q9isIHf2ZMe2x1lGVrk4uW0TXPuLjpCp43iGEN3TWz4p4tvvV
cBbwZozgdbF2t5jbY7YTAuqRFnJppOTLhLRh8tI27e2DiaBo2BM8mPmlPJMI5iTp
iz6drzesmARZL0YXdb1V9z30fpVDWmiVj3mWBODmFdVeOs4MU8AtqB1Rers8lIZM
pBxcCExAdWUH8CaxElCm7XXz/2XwP90FTyhS4u/f+99XEhuMckRRqM6OC2nG66VP
dsEPs6bivUA3XmN3KiLNplM5xaqDAbXtsZ71Kreu/4ZDmKJwIAHgOstgTNUQNGY9
0WiJoZD6/6ZcS5+og0RpR3qof4zyT0oSNGvunxBtr0Uz1+k0jVjoY0n4uSEA1rKj
IMG9WKt4bK1l5UkVkqeahkjp8Ey9tMBI2Ou4B+eVPQ0nuh9yxCDOxAjohz8a9Ei+
/z8ffpk69bb9xSR1qgkBIeonDIIePzM4re6UwmAMLwmLk8vaCeh+XzQY+PO3wTiE
rCiCzZXQc5C9RlJk/I+38WOqgNULBjbccoc8Hcr8SswawjksFeXDV4YZxGg8ZCGm
Oo+4H2oA8NoCeFzUHwUhmPrBuB895QzP+7O81uzUO1K4CSNz7kICwQ4oP6fKTC+o
AWqB8U30Zw+P6Tp0dghC05D4exzS6h17y27EjO+GpuvdRqlh4O/5Q95CiGh9DwjX
8sVXUBMGiXqw3xdhd/Jn2wyuOOlS12I9ZmVAv4kgA5fCbwM9VfLWHq5LlUEoRTlp
KmJrPeqeiEF1URWbNWmkKjZ61EM5J20jyFMNLiGTqCSKAV6QrGbNWRVwOb6P+pH4
xR/wgqx50iAetkvA3H7YrD/iri6EjxfqST7x0MTH1+1YA0BKrrYwI8aZMIeI/omq
1xRpdVJwsXjK9n2RmdtzGGD6Spmy1wtjZVi00I+W1aCHsUFbyZg3jL4KKoi3JOOc
ItDosT/bcStFeDJtN6WHufc1Mie7cEkJPCi2Nm0SbBBkKjJdrfRMFGDy212aLxBz
gMkJPoMlD/VWJLs3hicWYt8MspNK3W13cvyGnYGVQpBl3J0Tauk+8l8jFRWnjJrf
cNpXL62qx6vMETsNAeAljCdTcKCj30MwSTEe4AUuomw7OPcIfZI9NYuFGNbRENPn
pX2KiSCeuE5YnuZoWz2EoZZh5OvEDKjOFOZROt1oEiJFMAv1jDQQQ1SV8/UOynJx
M0vY34CWFHCbpU6OQIP/B8lXuGKov20klBYxatcQohIagpmyZk3djdfNQPXJAtqN
uAdoefzNcUDxCpwiKt/+WVwavEupurEkA4nBIFAoQMfN73tKBqf7+N6uBLusZHjn
abZbzM3jecV57OsqVGaS2TL+MRLFo0638PceYjW2fd3+0T6YMzSWD/++jAELna2u
TVSfJ6V1VxJufsSXHHaL8j49tAe8tX5yABmbYsPyYOrtlIKhBVrmffMQiPR+qccr
r3coXLFUS/iDqWKhw9FymO5U7VddFXB5zDqkDCK5xP8o48m75abe8U5+Q71Mdp95
aMQ2Q7xKk6Aeleqbc1y0TiFBoXkQrn+tlm1p+V6CKTD4/IodRGtCYOM4e1DE6CzX
VBjuHmpyOkkVQwfSPo6el693J8KcyKmSoYkYZEHwp1ihuOt5JMSWCbJDCMYcUVf2
gR7IXcEVynZMhQRdmqIwHTaV7kaGNOBDSUn7pi8S/kp/iUT1N5klPhCb5Wq35X4w
4706yJgoAjk1KDqiNImAra/n7s6So5d/wPVKSP/K0qF49/09P0zmWCckZwTNIGsR
rK7LHUY/Xi4IWXSG+54utSzMPC0UJ31g0FSi88tRpMipWpHTcKvqoUPic3vZ55UJ
0IUoIUv+sv52oyn95n6eViKC7j6dTs2rpvqP7N3eTHgFH+zk5FWHLUY9ARHGCz7T
aKnyslUQj6ZMjLY8jv5GWHV+bY/lhIVevOyaf1uFX6+8Jsdh6T9h1IdAE4w4L6DP
ej42eVxeGiywwj1ReV3Gtzv1Qz+MdxPZuEzGmhJ5aXSkRI4Miuc7oU0F46Lj+TZ/
TWlBK5b3xf3S7OZZIkX89LlUBTUyXm/iDn4o3tQL+rNLpgplHBrqFmRr0he8P35B
AGTqiWM/CRplQHQKsM7r86KyjK8QOe85AnL50JYxUuCE79gDNkCOfaxShDc/EcHv
Qdyzi15FfGD9m5ahaboZQAmS/DHf1rXzdVwvT59Ux4eb2U9eW5qCgEQIZQFIHtzv
dVl92KwcrBGWCZXTVZj4r6YqmI7h0LVbZGifyyWaXV4qh4CS4XFvgQtwCe3zlT8l
U4UmS7OwOnTpVh9MTFEn1itADQ1sNpQYHa8jjZBe71oIiqEVxgpTbWzuNjB/7Srb
JvKVaj20VNr5lnbdVcODth5FLiGotCzEefPFa26bLHsVGAVEg1p6CcjON56YUs5f
ZpV8NCPrq+kNRPdwwgcnwQWoKMoTWdnjHXZL5qpnQ6UMcygoA8q3RbF0F7+CPc7O
R19MzURl4Ce+eDPDsfBe9XowS7pv/UCTKFb0WHe/zbhc7qUNXnh0vOpd/A6tD4pN
SyFpVMZJd2UsiZB47HjRTE/bz7ionJnLEGXoTw8qldDE/9+Hb/wn0v3fo0SsZvNy
YreKw+sN0Pl0o1HNAdiWpTHClXETpwkphVHftJ6UoUGu1/DsUjKOy6ydnOXbtSi8
XhFkrqWUlWJ2Rhk2DGIr/TRZ18ey7ffrlqHtVGpGo8q2jxFk+plFVu/mdWjuAP6T
fAiH/m68+SiTfBta3VOUxGI7iIF06KG5yesCz/xRpmctueWvyfHaf5Yw8SAHjEtQ
j6eyc6VHR4uM1v4VtyMfoydpbg/r7ObkZwNpm6dA4J4CXRXV/GPCLLAUhe2n6Z+q
7ICbH1W5dvH7vW6Cz/uzjwde1HOD0MKCKL6J7s4S9WFxZ67vAp/0jR6bKNoW9UsW
o4YwHs+Sv+7/UL6/Mz9qSr5VwIGMqJReLpZRknaG8nFJIyJDMhZ5F5SuOwOH52v5
HdybFv7zPHITb52gdgH/6AZ9kwKhnSsMlU2KoRES6M/G+eIJ1r8Gmxr4Hfioke2A
Sav7v8OvQI0xHiqUi4X/j/nhBG4oZVdfGby7/1epXz23MNTc+hDijT2ZzS4xCAIt
NNRlZtn4J6jH7g0rluzSvhuTFv5d2Cgd7Es1C5qUkwRk8MWZy+NJ+++RwzVBBBq2
npf1/VAOpNhZiybmMnEvwXO2Uh4ReaRoHf6Mct9I2xjF+k6r5ulXRRUD1enzwZJi
9GgggiXgA7V3eCQhY2s9BtepzRQH6feq+SnWbr3a0Wd3pLfwy3zF9llQjVo2TvKk
oVbKYRSTlFs+ZcQljKa7Hy4/SmoldHfW7mPuyluchMI9a+eb2FQMtIIGods3UXc7
ab/uksdhI5IVEfgi1CCudVVWV9blHnO+r3QaDa28M08MahO+H1Am0oaMmHkkEYeu
7Swun77J2G7uxl/OIkPQ3nhvekdYmKZmsT+723sBtFfuRvYVnn6jReVE0iFV5nqE
2UsLzaANc6oMEVx1jyH9XVLPzfmBcAVoAO8DOcsK3PEIU21vcGEXJPA4mH/SmX48
/ZalUTch0PI5tgO1iUmTlYrg/SCQim2JcoIpEmPATwAWlyCrmhR9hD2TZ605fjah
xNV7G0LYf43lD52PfQWMBOJgZlyk4LF3dr20Ptq1AP/mh6AAqcvPG1V1hb0MSI3Z
A58hFS8wCI/tGT36fnRlqNQw6hNpO5LLCEzsvdbwYjxsJ2La72QKlItWW8KMhNE+
l9kmV3yTF4C9oF06qngGIe5oxs85siMw9m9vmT7BeEy7FCgcVySrQFmvOeHO9rYN
pBAdtfolFvBX8qUuW1rSHVoiGERR3w8VusZ4UJvq5Q3So9TItPVHNCSFD6PGOIaE
XhYpKAJqxm+MyMJz8oZUNtH3DgyqAPwpf5lUP53OYtqV+Iivjg16dFAYrPdyJCTu
NGf7QsoE7KC2QcxNwPPRnE8eO0dh9oX5nlm5EaR8vD+TdiaIcTYDz43YGsB1h6nL
4AG0uaqqvg1wylSFmY96c269vTeC76/oqcfjp1tIeL8GEpDGCInzj+72XQt8JvdK
E6HY+DHy9ecnKBDBzoKCIypg4kPKzbexxyEbbk7TlCayXHqHsMlEt3mBjSqQrwsm
r9REYCTCvm1+HdB4x3NmQpQgS/ne3S7z1oId6Mwxj5vDpWAetHH/nTW4dJmRCe+D
A2YLNPKhUf0DzqftDoizZnV1Fg0HWrkI/L2aM5JUxtbYZkaZQO5ItZojVFNQ36kb
KR6AZu713htDmF9lHkHUyQNAAtgTE/vvqa/PT8fQBcIjUVM/ye4Jcfx0trAYN3An
j80bsXKxJwKz0/DVARvqdskg8U02QXDvgwnIiwKtMHtHGqczaAm7Fm5Mn2V2mqwn
smd6acIkAC+FOaDaubfXPXg9jNS+ANJyH2AMV5UdY1ufv9eXjBwX35q/agy6COL5
a0YjbbPA7Hq49Epj6k9bj40iU2X/reEca4/o1eyhDhijqtulhouYLfxPDCgUi1/F
YHZZL0B2NgzQwzhlX2qJ1rcUYaZTVzlMsuNJ5bzwcGk1BmMpadQ4uhSXHNqfC5jV
VlDSM+VpRu47fkHlvMMNBm0GaP7Qoist9e7xlqpMP929BuHYaUf1tZ79vxLlrFQI
KNj4LT/PylWWzVzl4LY+bd/CW81qbEKkHUmJr/PRt3/+Mm3145LiQg1k6AW63BPF
GVizOuarRiHdP/7lNcQfBdLjnW54nDpXwKw34RHKAWCRqZMRZZn3hi4lYgxg7ero
28iX36bOs/TGdYkT1krnQZVkbKF3ggG83tt+IrYH6IG3Q4s1EExn7nUggyt6qWDb
5+o2gEOescD9iIPzltIkd4/wPMDD8TjW5v8YNGnTTBUDTpKMO//wgOt+YYEVwI13
ayNdvPr98pfv/E2Mn3pDVekKQWsXgWj+xBkXHKspVTh84xud443NN/9wPLjM6lQA
041tcd60kwFqJL8kpMcf2bVC3kqU5vqcuJLCvpLYtd/z+XasIK3XOJ8EZgAuvi8B
6+kFzuhdR1YjnWCrJYV/qnQU+CT/qCzPyW+tbpgoUDGGdmLeP6n12hmxdNtRrZpe
Ayzay44wwAiHUu2xBzKrsUrEwiXhCJLwOD+C68AxP05jg/vVTBleumWq/siUEvU7
15I3FbwEwh61mxqwaNbeCijYxZwv/b2SobTx92ihFn5sRiIEGsUoVxWsFhUWcp0U
WlXwrfXziT5abrmtRYVx8kWh3kUK6E4bJCMTH55LTlTEK75OmfkwkKWjBeaeRaRP
3AvIzAiBI6ZIV38IdENDQ1mof20wPX/pFVs/rC/n9Ukitj08zLwM64h7xxA5Ale4
84GONSA+dOdRgbzEub20g+fN6DBmiC9+IiVVCZgVZRnTEmrvsYi8AE4YcWCCJMwI
d9vnycaP0B/6lbLT3Atx8aKK0c0JM/hHmPptNojdgXUttpgxi1cDYBvWvRTVyLps
xWGJzicvjx0lQoOKtTwMTHT3eL9QwrG7F0xgmBlcbFpw9OdNCA+eAg4U6wFSJL51
lFBVsWHs2XxNZ6ODeBfzRqVaDPC3u1ot9uyrcJwCDaWWN+vjn7xM7d5CEAMJg0VX
3qTE8x914bJ9ERXHlWXdJBMKenWufQzd254LviTNlECwOeNuiQ/NaIOaFAxX72Rj
Efx6hs7rZzfrzXoEZcaARajrfS0FcRGPjzKl3O/jYj5Z7ewzCDep2HCAZdoJEhPP
+XcnW9u9z3WB63AWvl1XfZkx4veU4wSsbZSZ7dwheqA5jasN5eEK7KSr7hGRu3Bv
Bejk+Wpi9i6yfdSElb2c0JdZNOJ8nFCZfbtHd4wogwh9ib6LCAi5wcb23OOYXulb
n2Mcd0UpsmM0s0c3j5OHPGj1voLusxpbC7vQPfFJOI/8vlwamgpvDoiraZkSNvBL
uGaPUX8Ccnj/WDyktd2Qygx3L7pp8BFQix0B/iBda3aghQNOQAgx/Pnk10h2AG+U
FinjDwlEw4cTrujDuD3dZbfxv6x6f20kjtW/q9VXRdqgmUnubueLC7gce68Exu26
usxPJ1HGY+sGxCkTdFcmU4q2IfRI4bQCgEUcf4w8NcbRw6i9YLS+piNsQiVvrRUJ
Xg5daemubaifa6NOYEdNfdTSQUVUABi7svokaAyqcHlnFivu3cAwaim6nxvSjln+
B6QSr7pRmtEgh5F1M/bOtEGMqxQkV/VITQ8NLyIJsoNIOMsm+Wmf6R7liP8JbkN5
ZORkspJ6RSeCqRuV8pEYDc6XeY6xlOnTa31uTIQp/DpUYAWDKXF4Dz8W/Kn25A+c
YpR6K5858XhofP1FKjN+uP/92SSjfGnl2PM2qSBGcnGggsQtDSkzS3XdLR595qyi
IkxQKPSOjYwV66IQMugmYM39aJcWIeZ78FMHvwkC88+biXm5SMk+nfA9JH8okKiS
qOYUM6VNqxN+2dIdanMeOe9O3yAQKD8Yvy8OPHBl9eRACdPGUb5Z7A4zlu+zr+nB
zOHZIEQOB+p06V/wRXitKJzLQhY6NDDuS6HCGrAkLSBklSXWq3BP8l/2e3gaSXeG
e4SK3e/ZRDD9goECmDu/XP/5RQte10j8Tt9d+O2VfAN5U1tahcJHP+24pWES24Wt
gGqhdQSUYWdZ/Jj3ZJDRAvu9GAo5fTbF/R9My4W+VWFf06YqISwvD8xNy8vgTVdE
irK2k2AbuNrxJDw8r6jsxkDHK0yN0tDrrZ0B09H96HM0rBR7ateSqFceA0tZ5EOg
EdJjgddSoJDDQll1E2ynQBH6ImsvqFnquCr3Ia/fyoS+Xmzz8sfrXbSa6iI6ckMj
rrfAM/wrN6w/KImLM4Hj3b5G7jPKlbZWdTtyOjc7S2VnoEnhjN0i4dd2yING0EB9
g4pbijZGOsSnGuuWoelC5ebokV3IlcFvxnJ3u9uF/CU3ojR1r2a1ndH9wKej25ML
qYu4AHkqpN1DQ13y26L4ESKDM9adhD3XcTe766Xp3SC4HfvQv5h8GNpklW6yyfGK
X//eupRzs0BEYYlQWeVW7JesAvMyhP6COS+IetMTkyFwMXDp6H/j1Y1opH5+ohlg
Z/rB//0P5f4f3rSd432kIgEOGuFVuf4WTP1U0KMaWGynvyWU1Lck3QHalKfS1OGG
ddghshSLUkvBk8AB+QT7TUhsFXy0HX4lyk3K1HK+yLe5K2/amnrEiMP0h78ulFyW
+T82sA/XuhWP64vqtfQ50HfRgSKsWq1bcaqm6RaX9Q6chBsnPfuTYBwE9x02dwjT
cf6pzf6AwYZQotbSE5qWsW5K2nzCQhDY7nU2tQFcBjIdZDMY/8YDCPh7lGMVlIB4
FvoePCY3WgJUnXzfkK1K6VUHLVWQ/SDYapeb8O4ZffGB9a0YW2ykoFV2FYtKkiCs
NxNMxgT1bc/WYMwCkjK8RKqoNjL9haVzDs5YbID7Sb4xTrFYRbjrTxXhYv0mmuPq
OVrRhPmiSbufBYEJcVqNGgcpORKoHoKACr/jikhqmLLKZgVJmVSHXN+2hR7ljFyT
SqET7Mno8k/SPFGnh4CkyAT5MzkDWtKjsdjbPU5cwKufL+vB+GbNufh5wA1O5H7B
C+6ACv+c2XxIO572XI2Zd+ViorRTZZcvEFHAF8esWSSj7S58+VA9x276I1eqyygy
F2dgKJAaEa7+iyJT8nz+R23+pUMp+aSLO1m7TjZ7+/KvUtjRTTk7MDFahvoBZtnE
vGJUfSS/sfAYrq3UGfKePBXoLa/39FBWimk+mziQlJ/IZJI9UkoqdEZH3AjasdZh
ADnKdgFNEJJhtW9AkglbG4NzQXHCQtAODCHn1RDahe8xA/YrsEUoRs4RMG9XiVFq
ZFYJI9cldLvX/Vu9iZHr1IGy8FQsw4CbCH2P3KJH+ZGYnGQ4+t1oUQj9L5LNrejK
ueSlJ2XtRRMaY6V/6wfrnbOeyV0axufCD3URWAHhpTY2VUANkJnwYfw5x/GgM9NU
C/YjYlPVeMHbl+bfBsw7nDSa6AAXTpE+/1cKwSGF7ngcGnOVcD91CQZhJ2YJjRZz
QG2W/mOUsWPKEcI4sJyMSfIFi1Q60tS4xHeogJ4/OXBqOYtXWFILF0wVX9MGMDRi
HTavBBMHEy5+sj2STA8xZNuQhenlOBqL3ESGPydbg/c/XLSlhsVxLOTWILi0vXih
pOoHM70NP3mbf3HJitV7LFv2bw/m1HLJLi/3JMz4+q6ajqmE/rVZdAlilG0GJWFm
pFsWNKN5Zu3jjPrqQdKbFJ96qRFnH1oOONEkN+0ABRrnWEqKTgb+QmpQsMRIu7A2
ImC3F/2EJS1bh9sJ+9J9yvFqnuZC++ZwJqYhBcOucmVf5b/MkE6b/gPHkHp8aCW+
/iwSeuqZkcCE/7ibWKue7K3pdOa/kXb/u3r6mTHlOSeV9l9phoAxyXBuoK111r+Y
/Q6i+oSFHy1SLAzPiwL4knaQP041FVPcovv2AhDcHFH49DNP/MzI5EJrB6mp142z
YNPE2KzezBqvbtazuUb3hwI+XkJA/Q+kbLjzjbM+nfeDCGTyYRP058ongfhDYHGY
MwWlFIvq5uk2/3srC6SJ44UDiXUSgIfSN878ejpKTNJMdbUubaYcrTpVP5mrr6x4
q+zImHt85VifrUkVEfq/Ewgwokd6dQtVagoNN1v//L0+yoK3SLMI2iq8JKfNCHOf
lXGlulUy4/hqiw6mMvPJ3P5KuvARaHWdx01bZQy7Gb5z2CG+21bTTsGeIWqxQxJs
tzB+D7OYGcX2cHzYbkTm5eMdjd4WXLKQU54HMCKOUq2lAibo7vT9Ocln+ppDqGCA
S3wtJcYtWW3bst+fM+9LmJcZCAHI04mLADRr3vwu8PKFd297CsP1bl3L+G0XhBSQ
uIgH0E/DXA4/EVqvZYtff/kugjTvXgtoNLmlJswgP5ujhyF+C25XvC69uG+hxaWB
yZwNquGlRc+TK0ypU3LVc3zKKBN+36kqKeaFM/C0Urn1MPBfYC6ftiky/lPaTujN
ZRRw2IuGX2V48Eayo51NF7WJ+9UgYbT0zCAIFCPJZ6QOZCNWs/dvGxZkFSgbRauJ
0xf1bbLU0WGrr2GZRANFy+Hy3AsycKX5sCcsGFIIj9SRMdC8pgXvfZaVkExC4JYQ
8HLPo07s7MGd2mT+As+P5nWl4PMupWo46bmGBuPZ1Jzy5TkWDMmtI4PzG0gR5A0a
aMldEG0AQJoWn1xo8bBQnktioAcdHTP6rzAOr56Al+/R7QSgov5xkWMMIjZ47txv
TVnpBWkDAYfAJA3pJNEVTO5gIcjSIoNFoEFekVBXm5ARcK2fj8yFiQB/34xmjpAa
jmM4MS8c0CpL4gdAILkB1O/r8oXglbBOTWSxqS5vEoVupeCkm+FNUnRpWk3gJ4Fh
1q+0DhbVvYjlyCe7By+V1gFYMv663Ndu7wXwMaQ6KjvaOkBnUZt9pcO8W6dJkIlh
fr95TdqnxJYFb1k5SLwHf9xNRWn3p0g1pTQ7q3wfCGqlEzYxuf9cxpcywTXj89hy
ScdoWQIdTdz/05UhVDbWf6aBLoTeD4J5K/XgkWV9N1LXSy4KEsmGNerZHkrgo+GS
wXCpQN8CvKgaCB8Dzg7XKTcGu/AHLWrAmWTRTEX2RY1Hizaz05vRabsTYOzAsv1r
dVDmiIVNVv6eREwT0GKau+IXlcvWegqfdIwk3o3mWzpjPEBDUyagtscdajKhSI/r
bmPspK7iIrgPTlT7yacmH9sXwkHw6MDPgULLFOUCeAjNLOMlmJWv31H+Ozu99UgU
8W2b3Mdu0DgZFwFqK4jDbiFeJOAPFDOCjv7RveOlAXPr/yEX5twW3SR/+wqSCSqs
dnMA9068P/EgtrzzhtqEbeQSUvnrbCi/jQxEkRPhiuIKfGQM9nJa/oXSa1Y7iyCB
ddBnYA0WPV1CvLbdl6vVwhJWodWKgav8GXKFJx22BpM8iRp5IhDz7gxzXN2RpnZz
/qVdrAE5TE3uj3cBzCOIcChKqfmZF4LJkZmX3dYyVKE1aH3BSNz/ihPAAVRJbCAc
856VXILrZOFwvLxFKLIDcjYwhaO//sMNuUYBF+yHkOLTc8pFUxsMK8c0f8HS+mCK
bFw6vI6wdjWTSo5PHJHqNQo0Q2a4OD7U/lJRAbSew9s8x/dRcK64E8HafSG3vMy9
0gqHVV4OQLK9fvEPf4h54PtNyJTl55MmLk+hAhMLvmPy0Clepiz8eRKkXOP5Fxmk
i+b7J5Xvev9kYEEWvYS9I+/fnnPBa2E7SG2osr8aNFGnL0t7YQLDCFi7RUWq+I7o
2EcbVj3R+/0+XFrrn0cW8M5it4kX14MD6rhnR22tM37NV45N/I3ywGZxdFYNux72
93GAZ42iv0fCZhJMfwUHlH+lPaEMoohRy4RHHEXTv8+SXs6dPgUA6Cvojsvr7sey
Q/dfAlJXimsJhF6JKjet25WvNWL8rCL/R9CWsqGIdtSd4cHIL3aiSQ5HgRNK7iX2
ba2QY34Yg695zv5mvY9YnuA629L7iOvidgblofUw5y/ICO+s8GLf7KpEHAsil45z
rjoPXF6JeW/WFsIQexiXacZEn3PBoeAeJIPx9e2BLmyrkIAQvlgCGps9G4BZzq62
VoY81Dk7vtyKRqyGrYk9R3Z05GNJ4fUUg59aZX9HLhnNSzk8M91ktIgDsj4Bt3Z6
gRHHLaJ2Nhhp8+5KbBCvImUU7d6ANzjkljzv/kaQ5ETTHgyHiEf6fvQV4e/F3FKt
m41RF8BZFWb4sskYorgQYFUfw8hL+RkaLJmEIarTWi7vlNoz7UWPrOPXXkYiSayW
HGHDQYaFG/PvppucJGI65XJA1fZ+dkYEcw1ZU1br16l/FlCplstNQQlhadUqf5Bh
5eA7So+kb2N6QHlrSnVaKMTQkrhtneenNj7CruVaVQNONwco5ebGT5DsN38WJ03E
PJT+/8ums1ujHHHtWStyQrYuBBMH+3Rxjcq8Yecx0coH0i9QY65Pq73gCOc4HTKu
lkhLCDS1/onNh/30BZBM+vqpxMYE9u9n9jBEHltFaOPeun+ZnnAWpTkUz8Ocjxzh
a+lifYdEe/NItMK5S9Yhmfil61kH0yJ4QNK9gnoNhOs2xifQeqR+QHlkDr7wFzZE
5URmMoslouxVvDykxqWGEPWbFxhCoZ6J1QBPcSXDsb1+13j6zA7eFY/jpONpuCHY
hWzqwZhMQnWA25yu48bODl5jmsDH01UybGtD9yar+y6OUEzmVPbGM9n1D+l2FlQl
a3B+x4zHZA63HWeDUiHZND3c0broD8iQ1miFwX1pW/DeiqXK6npvRuonwj/LmIta
NllfAoxonLiJNCigJlLbh2mxwVHmCu/tIGZJ2pU+BY4XX517oSPNHwvetK9RLO/M
3tjXPJeWKhbdISMny0YQ0u2ZGC6q0kDdxZu5RfOS3Dg5PcZN0IUN2RLxYJOcp/VA
taNyVGecPE7uYep3p6m0mHd4S1shNE2sgxhwmYVSQumMuxa6fXaxrCr/XBMhqwYi
PS15mtWy0nq0INlIglNHgJOsoGVE/8yjCjhSzPW98H1nvu7at++eJmFo7AapXffI
gTxOSmxIJTFOKCY8+wlaD0WiYQ/UAE/z7rQYXyfxfAa2Ohi9BaXG8O+cnmbELgA0
k8IqUFnVWQFlXLzlV5seEN1gZcdiKSx9teajQsEksJNeNgqAdIY3YpYoajkKxC2Y
NNOQ+CwqGUgtzNV26mKL4z/YzNZTq+V0XtYzHUYQ5+edFqnOgOAO9RwkSd0Kpjxu
o1YJhW/78M+dIvhYiM3LKmGJr9lR43Z8p/uKdJ4jqKiMoF/Auw5coc1Q7XoR6cuc
oKq5dY+Jo+LXRxVQ3hjh/fPBBVbL/GyIQKx5d15ktjerUIzfJI7q2U+i58E2A/sC
kWOcfipCiWlndAih7hQAQGeVIcbF3nmTxVhXl3a3XBcUHmZVjTYAEo9YAjt7fQvM
gP3M0eA0pYbqj2TXULv9mP2L9m6X3KmtBBrdNygA9gOMynIJGIKWy/qAOPWbGrGv
i54kOnrMe3PNZGSW8nx0cK8T3pgjHzdhV2/6bxr2w4q7fNnFrejkTLRCjIKVhO4r
BZwrU8kMpNiEQxez3zcaUIUu0sGJda7fFfZPmlu72Ux1WsWjkXHQ2dOYHqKj5fYb
apjHHJ1VDZ3Q99OPeidkp5XSk7AtUFCVhzNYJcJmX0exceJYowVjcICXYjhNWDmF
46X4IZAE8vUNCuh644Mz02Kv5kYwsbdhjI5Ri2oGPdqdUHxJzV6xNbf7LZlLzh3C
SQArNBpYotUMkR5G13Uznwt5gOaTz9Fb+PnqtRZ5qsfJkcYRcVydrktDKLGxRJQT
6Nrl/S8tZ91YywlOvtoesHoGqOuPPt9HtHqEbLe/DQCuspqBrd69E09kmzvCT2v0
X7tWNeE4bgp4vSbQnpdkBVKdRWicmAGGTihF+r7OjFky7rQ6sAPfM4ylyUH1acG9
lGf5Sjwl5IpUsaWA+frFMl9M05J0Y3hoWBvlHjSnVGGO+mE3NNO7FUvBNzmy5rKp
85sYVLyxaf/bsLYqAdbhk2flN3UDovR+2ez7ec1VdoP0rLQAcN0ZetjY6bWJnw/4
MFk2X5Wkemns4JIcOKYYqxhckNvLAHD6CzgmKGTGmtdN8hZqXdGqnRmXNplIJGi9
qNDvGNw6136ZluRxe9HlRx/vaVQxFbQ91t9GLFEDSEtOmN+JChn06Z4TOMlgsmGz
3vgemdhIsLtFshARi6g936ERUbLG0J52oWEDuxwsV/XKm8UmMJ0K0qbebC60PD7v
8xdtjUZwYB3ZOgE9MpZbRp6B6tmy0JKo5vEc4BWMJhd2Be5l88RptxnfEsk/O8GP
ceOQn3wSMlCwD3gfBqDGW7xtZe8gsr1yrO7aIQtdtjWOlneXCXA2KQyNAXA4yzbl
38gSOCE9HoOs+Kw48mmA9TybhZpQ4dIuEyR231epyXY2vAXufsR6S/TqS03YrNh/
HPcfVwkuMmijfUOvbzmeJn6MR1v3AmeNgJZGkP6AyWsnr5iCkB0YXpgZYet1FZpZ
x01QYuAeL+KTOKRVsMdDio1iEouMb1oOUIn2+IpYKzlf+jaJrHHbY8p24owAgZIs
b/7Wn1pYSjHO07pva+cIeqgzIrl9oWnoVsVqhBDAWeWuZSLAa9WV5Sv1kGQAAeCC
AsIPJFwPhhSPBjKSAyIRhR1XT9g8AaBlv4NaXoCMWJFjK/A8u0+H/yehdgdAh7ug
aUbeNdJiEQbalP/dpGcAaHTDfQwM2aQSYWeTDaAqHLMIpXsnAL6NwZhH3vgXCAjv
fVnYuSpzbQEDKfUD4gw3VpVNp1dYzYCFd3bO1U5ZRlKiDO7LfAN58c/+W6CkrRZ1
meSO4ERuktYSXnnEYl+Mjg2lAsBJqsJAl3LZc7pfvsAld//2hCAhINFVyktXm7VN
Z/qQ50xxpWQB8Bk8fhQrCdtoPCusN/VdaSsC7TjE4Rh3KRltyCOkRQJr3r/bjOsm
13m7TqX8MpJZC+UGatJxXRZIO9HD2weUIemVXjwm7j+nG+eO0y2LesHg1HldyS7/
Y//oRy/j3d+XbhGS/ysQ9rh2YCOEZNgOgQw0XFWBu2VdY2hPey7TcTDO+g6WRZr1
OutEt9MrYiTHKIILJ5YkYPmy4Ai+dAI3i4MPDUjByZIyR43D+4PFMNEfmAdcnX5R
NzbNKu9Kq1EKiQ23XC7mLrp4On42VzxOy0hZqhXuPZWYXTn7k2uMa1go8MHUGwWO
ei8TRUZeH6LhVdB/+Fvu3pSZdX27GwgbTNlVRYg1E91M7FSwJiCsOb697NdhWJxy
QPKTLUeyTs8uu5AA8zHetQVR5qQg4q3RnUdGKweLu08U2odmOFZfqQ0CHoL659jb
fA6yJZZHFB2Zy3sXfV0st1JmcJj7FgwGsapkc5Ni/KrmLz55cZwBcymXftsikZ4Q
BnXj5S/cGAJrsOqeykTqljGPLis2fADyp+KLge+JqHqQME35IfHFZCKJ+l5yucoO
h+FMJ2czIK31mqxdXcPTUvaHzqrYHkd4cdSeHLkBHjDXdb4gc1isVqx9Ew8JVcCw
I1NYJmx+99qbsjU2l8hW3CxixEiPm/biCSQ0RTtz0Xv4QM9Jk7qt7YlJX7Ku4wUR
ig3TH0mQ2VEB82UvMSFbvzRsTmq6x1VLwsyTYqjnrF1gEa/G6JUHJrPghzMy9dQy
llJN1sgdG9CUh7u/I9DHJ/P/h+J1co/JR1Q+uJlV/yxnLLbzbUgKvaVBtNmQ+HhX
HcKQHtDEzcDHYZkR8IPf91eLAubuKOCyoYnuTP4PoeS7NRmwja7o4/ewBnENLtcB
OxC4LKmvF1uQUwd1UvZXmG5gaTaIdU4+NBtstaRGUJI2NT8q0pt7Kwuv4KHDwRXc
rbvgxbLstxnZX05IZLklyuYPb09Tgz0zE0fcE7OG4sudPVEFiKKZs9rMdMdgFk/N
xDrTLedet+KpSQrtPLdz9B7EKgGjrh62oIQugi1KHRNERyNhwXKQPcifSOf59cm+
kRbEifvJatax0vy2Q2mAtLzxLk/HM+J7I5GEzMIynwXgJZ0Ey3yLiqKRdmbTuNlN
l/9bkvtTjrNPAKOeN1ebbGGNj1Y3DnzC5oGwfidxtkZtREKFNvEy19judHvhgVuY
UpBQszkgiRoFsiYGueTs+Zr6TuuGma1+pqsbqRZLxsP2Od6TVafDyfe/G3pM4o2O
UH1ypH7R13dDFtaRlMClwIIrRBNpv7tx9P8sQ2QHW/1yDWd0E2SGFyRfYRKp1V7r
Qo70ndmkebCtMgiQXV2WWduuwk9DKEN1p4SmE3tiKI9DfSODuI8idCHt1uLNiXTx
RZKK8w1lKHdW6xh+zqNrbJWX40q9dytMNBdRzK40DDIoshr+/w1wjGWIVQE7E+PO
w6SyZ/LxiwhwtHtDCLp6ojk3gNwFHn81GFwvGH7fKGWyeduu7oXjcverAgUpWfXV
Bzjd6mfh45t/6A4nDODiyn1WpUNxzcEd6MEZr0jLOMMEj3hSiOl6Nqgr/zKFlBIX
Sbxt4esMS3g+wiLcRAns/JY1LISO9vXJKLiiDM1Wmz2PDKO0sZcmWQNgxE/hG19Y
XX39P0n7hXI1PFQRmZaZmdznP/yEDch7PR82/sgyZrxmsfKBMciJbqNS7OwD/u/T
k1ZlSpm1I+H3PQ1N0d4mmvcZwBq6pL28i4vPOOGIAz1v10yoRmevuAb+vkkaYcST
KYivzy3r8RO/6MdMxI2der0DQIVYesBkBCoC5EyBao3/s0Oa6VUuBukfg7NlxcFf
sNdK73NQnfFBPHRyqfer6izc/IlDvoLGfBkZt31Es1gu4E+uPUPtWHGzvg3tyd3K
0rIIAUqyiMBoUzNExncRJeKaor1SBny6DaPtSm2JdpiP9u7r0ajtasYXDur/sDOV
vgD4hLmBuSGZGaJXq3T8g98zTMeBWuhYbfznN8h4+kCk7ZxwbSu7xHcM5yQqAW4p
+2z9DkToHMFshCRYz+zrfle45S643rsCbyb4YThFVOVkItK0a42f8GZf4E64CWcW
+8OMSolsCMJoO9KOgs4ofvzGcpHn0ESUPcZdzX2cN1ubnLP3nwzLViXFYhlhwQJR
Ffd21+xRIqGh+MKYSB0BpXwzwxIq7Zx4LaLAsXrFomRpasiwNIAAhGdnuWKv9KPa
X8HZ6rhIwsMQlfh9b5irE+TkXGQmOPmB3ls68vje4TTl+N1QdOQrO6pQ4HF6x2he
LnC49bJceTMIngUPeclRgcCCBHb+LWfGgTTQGwui1iaHQysLtxns46xOMT+Qx8t+
76J4dzKIdV30pZwjCZ6mwkWM7NlduZn5QI3OEHQGVP1CAnL0rlIAxg60aktDKz+r
cb3Qjb9kzH9KkQElgTg1HR13b20OHxKm/+4nFUK0RuRWrMI5aJUNxjT0hNa0SuQA
eN8m1eQLyawGpzuvXAo5AMEs1DpnWrWfDzAvBsQ77g4HKgFNxg5zOai6npzKep1T
xY+6B5XbUJPYxKZSpusHYZ1kNr45PCMsl4N+dBhxwUk0PdzViLkbFKrntmhUzGU4
XwldKi7xYrUvVBqWjo1V7d06fJd8T5zXj1YifIJXRSx4FXRabDSn4Z69YAOX5Jq/
QppSp8kxGVcJAEzfj9aiXSWBwimE0Vte+TIuJyRP7+juluktZO5GZ+ZFn6nqEzh1
JabNLgoGYUKnBugKv/4JRkDg18H7xq4VL1eRuexvo9f1qfNSVLzWi/LpytOWUJB6
E73t9IJWRieeWlwc4shqOT6Q9SzedYmJXY3SczTizc7dd62uQGODRe26ZE3t5O+B
hEka35+O3NRA6fRNoZbGbgFV+2/bP06Xub9sOq2ARuaUVhpXZfD54jFQd0WrM/2m
2uogUOA+VOpiE35W4klBlVoCb/eXWoQyT9wQqg38T1wckpVhJ6rwUleMfHdgih8l
LUEPdVk43wYFR44hRwavrGX/4sSrekpijCtb+vilFgcizGAsfder9DujUQOz9ml+
3Jj2yVG/g/qMqd65F3wcDgh4lDixdkKvNijMTtRUYi7kmEISYt3SQWJX4luMOsdN
V4ZFiVgruwlaVnNFCKn798L5SkN6ZI5zod9WSz0YS5wWw1vvNbPTfDmBp/RO2cyn
OfmQ3+LfUdJeYFA79EQUcpa84jNGHf4UC2OsoZ1F1AXqOAHE4QWS/ZRrE76Fdr77
UFfPzNA02M+0TwmX1LmPXoD2HYBkGQM7vdYOr7Su61Pm42zPEneEO6Eu7zMoXuiA
PJxWeaVXcpBMJjMMdsAW9/vybBrAPVyWMjjlytRFX36wmM5Khc/sxLjAiv6i2LCF
dE1U8GsY814bgNQk6QYLwGsDD7wVxtwDceukbradtcICWl/7xSzESQwNJe39+MTh
C2cC5Aio+kuWlumCvwKM4Xo+XUhmZg8+MwPgO7IlD4PgxExAiTYzMYlZGxSqCWO7
jGobDz/xEob7Zig69YutahBlcfhKAVEaE+w3Hgnl1G0ChgxBM/DVufG8eUvOb1nb
kRRt7jS9Dsx4NHAk1sWOvHaGGqihvcL57yRAGAu20rle6g8gqM0D29JPzJp3qvJV
VcIjiIYzsHVfXH5VIWu70sYkzEMvZRGjQdweXQzpih5twVXwKIm93KTSQtCEg/f8
B0T8qOG97gaObIImdLDV5DoJMG2Jq6Extm9HCAekLL9UV8SxggvQ7uJXDVTKhZg1
UHTGisOv/dQ5uQinebb6xxUP9TkO7bNOqouyqy+Qq9aLE6eNT9pvK4FnzByKKl8B
JZd8zg7Lum8in6+Z6J/AANoFQYHZcQO+LxcByh0A6YEhm+Eq7pTnz8Q/DUIOX0sQ
xP/I2D06tdu/92ZVjDywOtZ5LGYO2nPn9ydbSPh/FBCzr2dcy1WCSBKTljL9blHp
AEWWyg8Iouv1S3f7+rRaURc/1u6VgSxUZQh1vf9j+GFJGRovPLPOcKrbmCeYgPZx
5tVFHnRcKWNXbEayfa0uuwPmVoXf8yGTg8Q7AD+XX+AoLwtwjehEQ2t2FIUC/AUg
L5aanKsyAZe41TLKglp+K7rkgOFxtB8dSqxaJwb1jOyz4OMzkzaDKkZEdhSIEu5E
mjwPk/i1DbOw1vtZ1lYRw/HGu25dcyLuSZqGSPYyYYj7ABYZmw5IbTexvRAstfWb
hl62iXR2h+7kzUv7LQGGjofR1ma1yqH/5fj5as/99PqjcFO+jHdUNw2OsGsA67MO
66WPII5R87J9t8NCmwCFMuEG7s/ifs2QEQBQbP+VHX9VLIsh4oyo3nhmFnaTokhY
NLHYabnmtd6FvSayFE0BkBp1t6u2yLGrUXGKvsvzj06KVG+V01+TlVYDMqsn83FM
W4RDjfhVPdulfLkGEfmsiGgmvncdMad/AZhZkh/u3r9PN6qgMqR27kCxIRLb+3ae
qcQKhyI/EaFjkeDiep68TNRY6NAkD9gv/UlEC8x0pKO01pL8gGODTRQ/8yxm8z3s
fdbn8is7KxpXzn4StGpJAgPJoJ+KnmdZ0FYdH9gSrQbavnkcQYbugexSP7kpsBrc
gsSoT2NIYi8WoJfeDpOPzmvPobBVN3YujG2zALYN8vVlXrWRbmDXAMdq5HoqIfpm
UMklZ9WeSXDfPMVXgoidR3t7HG2B/Y+zKgOqTSUYZDKTBLIyR3HKDdrC2jUyDI1X
67bPNeMF38nn1+odS4admb7U1bhclbYnnpm3Urfj/jHpPEgA2xD7m7w9MXl32Z/x
7q2+j54NsuyImZyqcyP3ZCjvOOBfLnpxa4uxzye5UjbTAD0SJYEwQS4bsmkCsiTG
+HkDaH2i79IEXkau/STyQnjZE2gcuWpydcjUVE7plhxejmrMvtJDhkCU6avhhp5U
mUo/Fo8Ei7CNmhQ/zuDCLCwmhphsfpgzzgq+BGLIerv1gJMnAGvf0h41Mj0ogTC9
3x2rHxJb2HoUenP11/tDNGN8FoYMAPmwH1Uhuhn1dLAK3SzrVjiCpj4WUaHYPry6
qEq8rlPPiJailxu97CpODn9DDlQBhLvU54zlNlt+t2OXcdHdcxcRRiUxCZTsDpFg
RjrqKl6s6SxdvyS5LVI6I08GUA4hY9/S2jKQetFqPv2VDAWOyMo8LwOVulB09Men
Jo3//n2sjaPll7IOpW1UVYEis7UfnZpgXhAwrXDTqDA34Ox3zPhJXgbnXCPS2yfg
YpX3Wo+ha7WPkSlaIbwiPg8+puUeKjS2xwzCDWZV6ki6eKbFEnr4zsBjK6RUefMU
LEA9tDcOmWEErM4RIaUQxKS8s7yb7Q7UKQAfPbtYiqXY+sHiFA1KL8U1SWy0CbOc
/gj2G8lf5RLzubzc7ZdMieh+c6sIAuE1IlXbIyqoWCGGQaQM7Zouf0GWBojVqDsJ
Dk3ZZ+z2Drj+laHMEtvvuOfdBD0l//F9g7Luu0KQ8U6XdqIaTuqZiR28PdPyiQuK
cUiNGSiF0ksqhZMIltS4cwmKkH+GjgxwvyoD7rtIVgXfImNpqX5BDJtITdf9w0yh
GHlcDApraadNnVBsKK9gBofprmhVd6875LY0CgRYoXaaoaElBjEego9226nUsrwe
v+nopavS6Rra7cE1+94GSp5+90bmcG9yH3bKvB9xoHev/+CZFGlUngYBJJIr4reA
yPYPOtdwczGjts/v1NDX+ZrvS1oyIBJTjxXm1d/NPTN2nGWt5bj2blGrKSTgpg8L
4FYKyXSDxPWDB5iSH/4fKJA6j6lzzFNbXrwRBGane0b4Wu+39rfdZsJ13z3XWhfl
pCxmMSQ2zXk8bBTIn/0+hAHWSNBk20x7UYtbcDINt8+Bg+RX84jvMbQFx5eIG/C+
oQAZkL8ugXVXouxaQJuHvm55MMgxgdP3ZReaUf/ecYSpnve/rNXD8+2hLEWKEHok
UM0g5llziSSRudbWc5jJbx2wxHy1QkaRNNi+6g6YIRPy0njeFn1i/vYndGSJexR4
Bmi9WCcF6C9et+oQzBF8aNoIFyw0TIBsVhldW22A8LyekTLjwu+/3lJQcJrC/mp4
+oFPbrU9rYsMO1E0mI10QzVUimF32HK8Dc6ALzODvME+x3JEe9y8V4LD49oKBspp
nAgVs8tAkN5sODM/fj1f0lWQnYIB4u5XEbp6uzP7wrQ19CRbGqzUqDb7s0lGhJZQ
kZlFbicFf0vnbu0M2aKMn9n0RA9G2X8BLiKG+OWUexBL9wx3m80gFvcwZyJoLTsg
gTFkAlgJPYHDRlexqN8t6wv+P7EqVXYvLhuDoxpVHO53fhrOu54TrPyc2WclnlAb
2AKsEFEn72EgAEkGiPw2uahfZe/UkN4EKJnoh3znAeqhHoIjEsLtNHXr53vUBZWg
g29VpZEfHZ85g7Ct9KuMC4z1bLEN7iYDPG/b8csX4RkPomr01bmZy/rvZMW5DXIN
AQ+29xylDw4a1hGDTeha2zSfiILDG8Dxeu/abr27SLjMQcKo4CJ7GAKiJnkwMvre
MwdngAbt73NTlEZfZYIeyyqCHnsB5edLdmJvOQQwLCR8X4Lc6x2gNRrZ+2siIL4z
mhNJwR83iXvOapxCbgvF41t9ouy+ty0UJ0eBCpXGJS4pAxH8R+12kw1pecE8c3H3
VBEBbnoDCj26dvwVKlPqzjReLX1pqUt4/SUcFRxjP1r2j0rnRuZXcJ4qWeg5zHOb
DW41wjf9SrBxkcZo2UxhWwDW6e2nfD2/W7ONlsvdl4FTcOR1OekOiyd217b939rl
fMz+gORlAVL1u1BG7q0YBpQaJ6EWABogIu6UvbMit7TKDkmnz9FURq8MuRnX3y4Z
SfxK8RQezHi6gpyUscba4kXvr38bZpnBI0Di42bB92uEzMFVNElCIdGkCjw+dVZ9
kNot5lbLeXAEv68DJ5+5Ag2sLu7Ks7DpWH7g6SulHTzlPekjoHQG4pwdBKeyvODz
/SQNWklQGDLAljOW9bMQvbsMnpE1msthCtCmVwLimVCjjz0c1RrPZN2URuaxEfiZ
pHreIg0yzguKoMmy8JfvfF7PQQDp2p2jMDQAh3CofgjI6O3lAWmUu06PQz6hLRns
u0vjV/dE/DXUXxKPmX5pthNn5B+sQ6t9kD/3moG1p88W7EOxhKmpqGgbSZIqFP06
rtxhdMobv2oxQ3hQubLlNkwm9uaCyWEqn+pqn7QNES5kbDzhsxPdiDFChHCHSgp8
2wam2DeBq0PX+MJeCOIfAKd8ES98LDM2ku0lofQxjPWh2K0V5UcM/vB6qNDnfQF9
D19XQ5mTp1et1v4vcDvKbzUbGDxx4dnk/dbOEmfJrtZUm6rnfdEPLmXwJHKRZ39M
vYdXyGTsPJo7842ygagdBz6AQ3OXWc+bU+sdSqULUNklNtI4OVWH02HIuuTeY+rA
8fY7A9OAJN+KluJBYcyLB6KnCc/XPd5kiDliP1BYTUiUvgKa86ijNfvWJTD0JjtK
JwRSynqxSc623Y0NP3U+n0rbFBVaZNRP8zl6TT5/WRgOT2IBviSotzL/S8Stwt9d
JChLaJ4RQeIpKbSLlbKdhJqqKpWepzL61K4H5Cce15Spk1o3tumFyDGLah5XWb56
RqOKp3ojP6B1y5Dd6m39+IQT/GMCzX9ynNdCYGvd2+hLQ1z0XE9q/jYZ3D0UCV0C
nsTcgwjjesISIA2zLR7OCyBMPBrf3IuvpH8sAinz3tlOU9Ib6OCvk3zq+tFM17Ph
SJxGnbmz6YfT7y08Qraj7DrljufqRgKlgZ4V4jUpU5vNAAhZzS1bJTO765EBH9yD
HO6LYlt/Fo8EOD71cpCazSpI9bLgbx6oBWBIGgone8Q0A+LkfKPqJpPdr2xt3eTA
HVD+guGVtj2dpDADbK64QoOdC8zt2WeLFwEUOnpwG1nxAOu4stlAcrZUNdNQsJ2P
7TcCJ4sNOTGAMNo7xoMwUBSBle4H/mdu3ihPSrhDsaQ0G3N7JN0tsZy9h06hmpy4
7V54lLVCPdh5/VSzzfE1TFH8m5lsy5Pj95t4Za7d+HyES+cMTQ2X1knebzXOTJ+V
BKFtXUuPuYGzwj87g9NAmu0zwQPRyNS372onz9O+fUhSaqr1QzAV2Kjg6g1IirHc
0UMYP02F48G1k1KVO2zYdHZJAj1SZQ7+fYLjJfhUvuwC+b6FHmhFRmJKAGXxuCPz
RC5Z83NBiZQFvbDTS0zuCikWeKxtb/A7Ox+KYaOLsuucO1OT1+AgzG3C6OQZ11lr
YPce4mAfioDwHIASfC1DItCDf9o2bKkQG8D2M6KF1qRuJrGKw1ffN+TA0c6ln2Ec
YYX+8gwEvp+QTXrdq+YKpaWXoKRmq01IBlZOdPmc6Q1VZjXoOqRob8g+/HRz6Jh/
a0C7jO31CBaixm/AsLnN7VZosOZJnRn1oALc9DPaZZOp/7t/EpeeufYiProHLChc
4P8JMyK9oFNDhBxKhpXYQXEwR1TjcsiICc4fkEHuYc++HuGDPZ4KvceYFX6Cz6Ab
RpC1b/GjiP3rzCg2UOthyAIS/PoNuYr18u0rivIFxm61bMNON71Es+upRKbMHVMO
Y8vI12qSAefMKOwAo2UI4dgdgA/CLirHJoN2Sb1c7ywhICQuIPrvAPRqp5o+S3qC
hznxLs6lyXBRJwD7VkVGs1ulGNtbIlZ5vmEBfzc6xscy0y289llo63936U0b1Lqd
05oqNmNcEUf4fueVQ3vujjeolIiUbCUB+flQYg2Qsa8+oQSYXTv7BEiM4NN2hxmU
xuU4A6oxdpjR4BI+nv8Na4oZ79gwnXmEkQKm25ITv3DpvEy1OfYnbr6CZBDIkElH
0hS+z9DZC4Wup3qeRGxrxfb/fy310p2wnQHQCmD9pXTFQC/WUYjAtEB2EULoME3c
za7KmegsioG4CWaPadej+XJ/NEhSySdkUEL0q6Mq2fOVq4m0LU+Y/kqfpALdmSoI
8Oo8GzKROd3wsZHP9mUfc+7Pp3G5PJnP5Wq06kJJE0awuI+RQwh5N2Wr+9Mf79Hv
7CKGzOt/wAjIqw0oppumI6COlKiG+t3LiP1Z4xO0Pu8EeQVw5rw8MG90dYO6zH/V
meqyO3tPsirwfKtbhXqyr1aiwbZrUweDJa5ZyF6w4So+4ljstLZLNg3CZsalHeMp
49MG2p9WH1P3jMZTviij6QYbMM+Hsfs3064+jCkIxJP/w6NkYmirwNFMLBbaN+sC
lQQ78SUj2Ya0UnMOBNEmpq1SB3LSmHpB3fAKV0ado81gDaQzf5qBQlk9Q/s2z3rr
GRoAO2lx+Xss+aA/4Et3SLl2gTnMovFzOB3gFgAiG/1mAO4OvivKEEyFodIsIhZe
+YFcP4eomKUES0xJPPshhP+1a6i2uA+Tq/LM/+0vG5tWoG/+KxIwB/iQagIfzFQV
68H5XECOlxZFDGiqYKRCkouSjgpZmCMRSs/jZCe2Yii1roqRn1sm/2a2PbqOcReN
1WHdKBhtzSk8iNYsKxU0ndLZ4cI6xPdi9BcZfY/NqfaS+idisWaw6Ge6SWhXtlsz
aXMrRfyObjeNg0IUEQ1YBT4hNiUlafebbELXUyI7XJ2yljzTBMxQEmiOhmrPRnvX
t8gMA1B58EPqJ58ee0keyORjxfa83MQWj0I/KBjI4PzwrObig3ejucJ+JRG5o3cA
YQzLBem33HymknGueNwDmev2ICI08tMX+Ufje229ngvNaIBDVipflpuTUV2C5kV5
UFhmJBEvXH7JfqTfZIrhDH1tEnTWy9yEMvtbfIj3MxX4JjFTMxiBWlO4MhKgb1ya
bfyU0IUAhGUhsvjUD8s6zZKi4G7tYcwhs9bTmi5kAcpEB+Q8D8PGxWG60gN/aHi3
kGeh6ysJiXSjUeFWnEMDBvLROHoU+Xz6Zze6heql3+/UggFPG6noRnXblqe4dmCr
cgucLEW+GTlWeioFfWV967lX818Ar96kVwa+QqlLQL7wffmLWuD73TcoXINPiDL5
JQ8uyzLcGkFS8+CrBmxhAqe61R7QjqskLpMePuPXE+wU8I60EidhKPGdsUY7siEL
fqBsP0571pKRxtxv6o2GdqHSVmfViXYQ0Ipq2h4SC+hoK0sisnJUZvfqSDQPmySW
hdobJqPM69AhL3QT65LDhl9rz+iiWHAq9TqOg5aszatlO4uvkyyQvonYhh0IVsJA
qh+Qj6CJqKMQwzEQxuidKT3jM8iYl2uIp5F0S8B+X+kiiRt4TB5u80mg2EwCbpTm
hILIhRxoYohy3a1TrD6siciZ67067NMTCsvKehCaXDdrq2YMpjVb/8bGYpvASkhN
F8AUfDDEkdLviQh6oz2fSJdzCOZD+4qUEqDtNT2bZQMJJc3UNkCYVrltD5g0xtoW
T7h3DUE4Um+BhM24ylsNdN/QB705Xbvujhhao0rHKDmNvqufyN/H93T15MP95uNH
HvXdEXRpiSnEFiXTaSS1ueZghPNSj6vcompApkj/Ktz08FM8DJmk50LJfWuO2OuM
GdwhRk8d7j3VJtb5cW2vPFfoVSNr0jWQCtRcNhFVaNj3gclpVVWJpkp4ASnHXF7M
MAOHuSHYlNC9Q/jZyjpGV1AzVL7mZb3WnqQ1QV4GH8b7Wxw9N8+2vcc5e11c/a4s
4Ig3n4Cz0wzkkQzReG7UT/OePCB7xHthZ3gLbS3uvYagB3QnbpFaDBnpv0eVmGT6
xbVUAN6jJpOQ+L72Im9EfMbKEthTboKBLg8FASqoeWgsBOCr9sMhUXC5gKv2RlpQ
KXa2oxAxeLehkg4Jlgc3Q3aQ7v0JjYpqRhERHT2GRIs+gd7m48A+0qrwdLqPXal/
LtXWgvtZSo+nmfEco6ZtuLUDdfX5S7PeQ/pXkMsr4m1t8/vPe2XrA7m3W44NihN+
/HMstbY9fLR+LrB5g/K71mIiX1ua2EPHS8mv41avJuVRfTdzSHreKmjj+NAwoBAu
4eueC7aW/DRehaL97F8RBUGh19p+j1GoivLSF0rWfG3K+br47kBy9Ww2BccvW0SR
bZCLxKEPjjXpH5rYDawyd9GOzoXtJqNvVsIFBMy9cSgrF3U2Q47H6khicn7SenW5
gYd0E2QkvdkdJ+0btBlnzrPt4/COSJpgZKG10vuiiAFC4jWbrHhjCHRlbWZd+ObY
ijlcqLaHCLQ1Iey0BdwycBfR/geGVfs953DRYUcoRMeykpimQvSbfKkufVbLUI4k
7xlcdgHguSjMfqLlD8UkvuOtfyd6BOqgKNs2TiB6+D4cire3ctsjga8nlpUdT3jF
h3lAs8m85pPj+5og5BXbXoL5N9TxWbULwwN7PlLdyw7iDLVyw62Z6KeKhkyKBGcG
2JWMNdeu0GKrM0Nw6QUZmzrsMEwXmqn7pi+tvVGI1ZgHirVoi2vhFBY2lj8T//mh
cC32A2SbUlxk3VuB75VJXuUySfapZ2mxl7T/nEmOw30cXAobsPKrJJCblY+UcTwa
Ed2rqZZnYVx2zyE6Be4IJsO8T8WYiaQAZ7OT5VCgNfQRTsrffbZ8Cz7/MAMGtCid
+Xp6vN7PvUojk8GOPPhuW49Eoxs/lvRTdu1W54BI9cINs93a9gZt4eeMOjv6uA47
HiZL0cIp95+K0Rl7Zoadg3cRSjdGlQpk5vOOQIG2kkt6obQn3Y3sHr0yFVZmpCMM
gFaB4JQ4nUzC3/nkumM1yyCmLlBEbKxB/1vg7IMx+itBeB+JJLz8dYVHqBdtmYWj
mBM3ijiiqcEdwlX5s/ubvsF5XrCDMee0+yTS+rSHkGLckVOMh0NYFt15PVTokH6U
CT4y+xkKBHJPsEmZhhmSVYZQJKZCmUYwj2RVkzmlwgeIZhutWU1xJkmuTfqr1j+i
OQJMHbBQXnzhLKLOit2/SZHgMP4qUcEv6MoRZ99sj8K96yt4eW03gD/jCWsU4VCH
LpsnV6UBF3dELNJx3zY2t0nAbRcMyDHHMHvovsd3vq+vNQPkYNe1jEibDgAVwaNq
uGMsKCHm4TSRkUFbqxUpMwcU943UybdBMknmpbleasfUFiUkb6B2hR+ASRoUjy9m
M11mJlATvHfdiuzKGPC/EqYEl8/aDbqUGYgK3I8yUlmT+/uE8bWTa7IAU8s/Jyu9
qY+1eYZAa3XH2gyOyJs5f7r5+vFsUB+Oi+6F7xA/dW5kqSWdwJqyuLlx9rCb5nmA
o2deeJEblZnb+NnygsZh6OiaUzzq9XQqXeBJgMgYydoXxqGvijIfNB0/x1uOdo64
b/LnrELLjF8RHHdr0SSbhXCA1k2RvNmWRdN/AyN5oSapEvzGbg36VfOkmmO7xvGT
5MKMUg1mSqMRnzlUUzl2P5lfL604XeClK/BrLJq9S7WL/PaB4wnq/z9dnhZULk1d
jgzGfS+kXXLZQoB0hFIuhEq8f6+U3zph1A9x4eqGJ0g+ajTp9bGh503eMKgzRRih
6qLQHWqpxT64Axok+wFhExrm++jYc01oMuDIyGOjo9+exW7kqzA2matSEfkdmDYX
Mt6F0LxCQqDNWBPdnKZuc2/I3CLBOeylED6x7z3pNxxTH0vjKElk0sW53wy+aEYK
ioXtCM7D/h4+vhcuTL6Xx9ubVh6SECnXTNGM4no6A4aVpQ38R+mrERxIoL+Rtj4H
H2e8GVufjnJcY+49p/CoVuN51rL0MOU0IlDgGfw2u0AgB6eYDtn80+7hoYBV29HV
JCalrmkr3hLbarsKlwQGAxAc04TX+JW0E3m8ZHX0T6tNZHM6NvPbJ+30qp5tGXso
dzG+uY32+BY/Hi19gZF318ucCDFzDFdDXGM2239/cYAxTBSQgoIznay+dK5TezBD
HqGqwZVwCmilNag5cePH+wK3HQXT9oWpBJtnKv8gKNG1P1+ztpgLPtvjxeOknDLy
/u1UVKfWsV0JtiKEw1lQgT22ayjEW8K856VCS/kBOW9mtIvX4nHD6ifhdTjYo+Y0
n0pwc3iQuBjbVw9ihhYcJgLUmuzivBSv9MNVUIhBygbRl2eNKLxFtPeREeHbz4ZJ
KeXsVjCFnq6wcd9lptmNfZ0lhO5jcbUSqSB9JuzKucP5m9ciE3gSgldyYar8vAOI
CYYxSO316Y3Yvdw9q9v0Ybc0b1bDeITHGSSEpnzKvfCncwHQeByH2b3SfvsZlY/q
ppEiYZ2BP3a5R/3/fDB81HxIepy0GzqFSAiR9xfd5It+6crrKHcpAFHRyebXxnYz
SQ/9j36GnKd7fbHgvyz+unT5qWY1fMv1CpV8rLnhZ40489PADeLxy5pf2tds3V5M
7eai08+yDdGG18Tf+ZJH3/ehBfiU6THfGRIVs1gCgDuZb9wBa8qFABseZ8g+EzSm
Yml4rPb0wJ7Vp8c+LUdDjVNO5lrJi1iVSe/RBBhSuYG/JF7bTsyDtzmuOej2f4rR
vxqQfxlohcckzZrxot7KtggyZy27pdE4D8fVFPjaj7JjF9xJYOXm0W8WW2X9WuvP
YEPTfHAlIl89NSoT2kVh8TAsNUqHx6opnKC4cA2Jwcu9JddfWHjuoFk+w124ZmeR
cBBk3PtI5F4SlYo1L7cCRg2PRr5CEKq9VuXJTTsUEQ9pD8HFz7asuZleYR1bxppm
vZVG0cUo+fxMUicpub27e0aM2LDq/GAtRXhSXSwKKnFi72wuRfgTWhVMZok1tCfc
25XkJtWe4GTMDH/hE02iETy/4iZD07R/SdsQ74Cne98FMfqVOTqc1g8aXKzZwv08
RG1qaID9UxJ4XABnCcG0tl8PNPC9o7v3jSB2rz0IK6jXr/CwxKufpcLIgNjaw8tK
Y+gj2mAomcOhdg5Bdb/QudcRw1S0icXd7Hf5ndyCK5FjgzkLU3wfBEiFu/qsH4Bi
ZYgw0r1NJ/GLlSTIsHzp+cWXoNZvm9YwZLHnnI7C2aKU21e4SEMQ+9jgZnveib7c
QXjM/nHboAk6ouMa2RnLfwsJ8m0NomJVMVYQM0FNYZk+t/wFyOMgf9zXebTgm25X
DYISfvcTpn+vDvlHVtleWYboIAJQ1zNrz4oMAhCCCvierxfChcTiA+fsp6jT3G0t
l4u9BlmWim5BmajrPfhuHLK/LEFtDlVSiUVfp7V6zjItG9WqEQ5ipvn0x2+3Gnnb
nNffiMW/DrRbEFxl2X1CosyYXtu6yDI4L4w7P30NG7BLIeuYTB2GCnMd1PPDJxdm
bVa9vaaijznmylE/hlyVW70SeLHcy0KV27g3rHstrhAhj2HuWc7dyi58Jajv9LwO
4DMYU/l1ksJbFKU19Azn68PHK9Roe5Qjur1xl/9BRGwicskSa642nEqpCsiMgySE
0JvmALEyRWreiIHvJx3hCfXhipWwlEYNSfJ0kYyxRST2JmA2o/dh28dDHl9djwug
PRyr0UZJOpIvUQTLregOz4ipvrgNZVQuOZmPoUqRPcvq+GVbrciC2tLo6FtVWON3
xSxCpMFBrPAsJso0lXtfU4XzuBKINsve4nElX6HUS4TA0/JGP5fyOICpiM4K1Yj5
wqYzIITe2rcHUwxmu6sxuYQhx9/IVXRgyiWbcfHEc8r3eLZPt7I1IsjjHBy8obAX
TyXBTenm2D23KVtivuwco0JkzfrfQW1geWnZBmTaZnljnqyss9ivQ6CCJQgkbByN
+Te3Eb31QlvmxHv1FPFdLMF3WlRQYg83nsQt1RK2BEITq/egFPhC1kGmWtFDDr+G
f8EqEbIeGPHxiehagT2036NUj611scxVApEIHWrjbeqOAXzntGLnCVNq0cG736Rg
d3uPHQqH3HOiyPHvKY412kYG7CHFhmuOLE6hPFyZ/N6I/dHHTzMtQEaZSFbnp9ME
uQ2+5Tb2CJIgIeD0pwAUYd8Nzn3FvzeEJ8Nbpscm9CFUzgsgLPhkJYoBhA1YLe/W
oXQGo5b2BgN8DYwyxef14Qljy5I7shRskgwNww3+jY9GLEdNcql146FTDS8YCJzu
r4QZI8oI13fBwLMzY9W+vlLMusk9UOVEmC+dYw6wmkiIyn4ajn0gz6awhR3NELkN
zK4FIAOx2Ezzu2IvYVtaal6VADM+hauK7x0cYLZFwllH94bZN3IbC7Qh2K2Fsd6v
xaFdoN7ISiT7GLZcR4O6DcUH195NUzhyChh22vWV+uY1ueBXcUDK34LZXRm4OSa4
FvhtvczLnkmaZkmeEV9U6HKI7B5NOV2X2YN3IdFBPoUIiwwmeir/R4QO2nGM7ALO
BMNNArJ+OaaVb3qTBSYrJ9ycOMoh1HgftejapjUo3r50/iAGYnU4cL2rlpNufMN/
Ajwj386nkSkDzlNqpqn1MO1zyiZEcXs3GBcLa3RqY4VK+wbV4fIuGMxRQJStjfn1
ct76rpi0lS6zc5nzcjSeGOGKY0TFGkGKtBvfz3vuKB6gxQ0T5+F05cxUtW4m2G/Q
wbSpi3FWLS2CTRDyrDbK51U+px+hf23y/xDPl4EY8g2/yTt6whOyX0djN4s7lbGQ
qsmJf9Y7oqZYPV8+4yMglzkfu5yklCHWHK6pYCtD1BcIa2ZP9ki5hSibKVdCoyK/
p1alRErHO1f/glXyUNFqLGRhphnAaJ2j5gwtXXh5Bev7ZLhYSbk3IhQS0d7bBUsL
yGEKXUeKH/9PATJ7D7Eh8U4u6EklfVXlHTys7B4o7zp7KezyksRrYN63tNJbyaQj
L9N2KZBWks2n+UOWmkuD+ymskksInLOMADumeJ3A1YRuYQgdSN5ShDyiGv1oBguM
BajnjEQAFyaEH+DxnyLDghwUs9vtgp83wiFZEjQWLW9A7gjjDTm8MA19XCSeHU+p
tBApH4wjEeM+VEH0G/07FtQ7ec3PfbHGEEhj2w5EtP4kC7KvIE+zZ5OCOH2vPjN8
GidLy3wipOONiSi2EHShPqCEMiLhd2abaV6Q69Z3nhn5UfdpF/esZ/DbnMguDtN0
7vTA/1/9wOKXaUOj/G/0oW8GRovUmMQNYXgbb3r49kHLsWd36cmOshYmKn1Z43tK
MYYBG4MaMn43dlXWOxS6sxZQMZrFfHize3h7bboHAKdqBIwhDlUHuE+w9dx1Q6Kw
Ljx2osAG43NDNw5JMP5gRPfzZ2xddIYGNsL8pgVJojs2j3V/Q7UovKXW9DdwRTMp
H94jEGlzwa9GgHUQ758XQdeWcvy36TkGZAYlZEJbt8b3HS5YT0FqDZ6gKwXIyfPZ
4GC2HOdiHgkwyIFmyWtKQ6JGBW7otZVlU79SIf3z5KaxLdsfmb2PqIVby312aZRb
X/hJEksZcfxkUQladl7iSWiiTv95uN7h+60RXbeKAqHM5q93R6OSwQ+nijZm1HQb
BKpjiE2sVKCRC5twzD41Zob69GYJCcr178RmZIWJasRDh/lHsSOYUHlBDKFJHmWv
TXyxBj7kOvbpQrjr35BEj1js8GJICxlJ2rskT/+HKV54lmqF6Tw53g1TwGKUEUfX
MI4ofpTdADzDsmiEM+RJF3+EjL5hmLTXMuJ2O12RnVU0ntccSFuxi5Fa8o3Zxs05
dDHuHBS7PPsTDxnf8zVmpEJFhA1/7vVbdGKHUpBYZeejRGWx3P5KO67ibSgaBrQK
3TTpZzkG3QDpgi++ed/bF9Gbod02zT40z4/AiK22+DogLtNmyhIz+UGphsmh+p3W
t1iXOsEk8FIAB4osA4NtGQ4cVDa33p0yypZQPO4qrjKojeqVmrnAs0WWGUsPSsYT
9QuEwgFP/tNYx5EKXnzl97CNRraNmBmaYOh+CtfaxBBmuh44MH2bYjEy8UfFZn2c
RohwOpdHvebkcbuWFdW8mOBRWmt+50HeuHhgTyBwst6hcH1wjFSTh4x8g5j17jrW
2icVtquiWyBf/Bx2OThW72RNi3CYq6+MtNMMZw0UiVzst+8y3bFvze5GXPE3M03M
fMoNQHsM11LaNWQDdldNNLtgN5UY4ieDuKb/UK2LmAqJ/DkvcUwzykInL+06az4U
T6lZzwQ5ywRIOfBAedzfSiXG/XVjLmo8Ik0in65nvzK94WEsKAyIOl9oZLUoMxQn
6WXwswJxeYP3h1NHXQdw5mpR4DIVJ8SoJi8pmq1VJ8J9SIFL+6MiBqFuSm+WtriN
B5kSOInHi4dzxbLIq41UF1RUf4awlaZtDdaiCotJrS7nijBIxch8QC3QZQzt/KLH
BP0W5eREsvnX+by7BrKMl0S3bUQn6rqr3WENeGxiYeNQtzfRL4FcIaOxWTA+7apW
Pp8icXSUOkEfH5B5lWM9AJkqsxNRWIeSaVfRYC8rgiZ17l/Q2QBeFz7zvATDazHa
Qk+JwTMf4UtLemgBSG3ebt8pGK0Tuoo/MsvknNGshJgaMBy9PfqGwiP2Ll6DbQWD
GkThajES+QAv2Atn9wkvWnRaIjs7kI9cgTzihkfWcIWEt63dL25W5crQ4nbOqKhm
4pxRclj4i2ajUVsrj3FOhtB9pdFHLMNHkFcQuESGDG+pfNMQHx4Z1EB3EjPVlowq
F+s9Cah/KWUXtXNNzyxtkn0H2du7Xk/DbXSJeJROLrAjcPSQ7yh4ob1jGiWSoFcL
KXxF9nccw6OUx3vqWJmQ9IzFpBWkuhROGxT4mCTGA9klvb/3k7o9/ExhJzUfch0f
6GEnnmvvYQC691/hPErWNGg9kUj7dCp9gmcConCrYwShOrmijYHcX9SswR9R4iv3
9IaCsD6fLOHRMsUELphfCxZpfE0MtHr6roSCXJxxGgRbkU74LuaqWJCbIbdQPX51
JrcKBREvRpvo0u7q0JfyRH9nsrSjfrKLK3whhBj60rnZTgS0dKyzgtQyWYvyJQFN
cAf+rqpiNyNnXMZ68CJJIb5lrH/Ys/Ke3jgychv4uFCEATaozIAxuexJmcaxs9NK
or601FwnrxxxuhAi8GyUd2C1zuLqSwyc6CkDdjcO+vpfUKeSBU2SSnurW44N9za7
mFVb/Qo9XgMKIksR4GknhZMBFPp6Y6l7W5/gbF2Q3RP47zhH2lXJ1fw/n2S7RxmI
KNF9p4JPx7mJr1icxdfNMBOx9WGERAg1E+3tUsUP0C1+SA7/YJH1PGQE/muzHNyM
ytwaJ1Hopi2G1i0Ho8JxLSOZg5liJvmjadwJZIIKOK3iS3cki0zhX4bh3Pld23WM
brxWRvBWbmqbFAlPQ1DrFJp4gaj/3EJhaR4y75Zer9MxEJQC2SJnGX/TjyxV5YlI
vDNXS5L1TEJsSQSpKTDDgNOiTQzMhCQPqnH6HnnlVfzdBNgfeBEsak6sZHlyUdb0
VaU6qhdGwU2fYdW8957QURE7XShsyOo6DXVBDjem6rU+jZEKleAOqnrt3fks9CQt
OJKqrgL50P9RacOOaZqJIbsKtwL0OoPG3MgEcO/apZJThcrIF06sdAH7nf7f5xS3
hfq5nVS5vDEZZtsoGgP+bDNud+2wwx0cMLRpiE0C/1tGLwpUGn4LWyz2BGpCMpHA
T+zLaH33JEcEvTFnGiG7RnMPAPKqTAdYbogX7Mw5Z8BB8z26sJ0X16ZkcHut/EXk
945qqrC0O5cOsRAt8VLQKxI8p8XtgiPjelwsMdcpJQhSq8p5LRE/ZPrP88FEWy+r
WSklNfl5y7VTbb10/oscD/hpMMRSq9tM843DNQTBfKvIec6FK+9m2VOGEVw+JaPz
pTWhBnzO3tQGya0I2y74lHM+UCnWdYBJWkdOh0gErRXwl1eho289vTsAt4MDosMl
dK/fd06EQoWO34sZ67MiD17fquwFQ3eRrgVoeXvJX9O6965WYD5t0G19qPcGw6CG
fHrWRHBcHt8HX6YGlcrM+d0PdePj/1ZyUZO4rK8NiN7Rstj4Y2NANgdcnP6+vUyg
8KAf40A1NAl5RqiKQzG9GGMmXw9ZpPYjYCzV8RJjZr4wRM3cEuHD/gbX4Jg9WxYh
uoskSuVXVcM3eF4I9sPVWhOJYp44HRkkiFvzkooi8TFBDeP4FD715rhloj58i8uc
aBMInKHkunmEyhaf5/24/8GL03A80hqns4EBgHc/mqGejXlJaw7ArY/X/Steyv7S
hgqAuGXxvDnZmsmRc3oT1YbdimTDCLesxO+GNUfPLPVExaZtPTvH9kZ2AMK9mVNv
7aNcIKJkPtd5XvpwjfzQoCQ/hGsZWcrFM2LXByHcRgccVDJmcAHDhvimfz5PGvYT
Be8UcPNxv2ooQLPRp3p+Vmefy4/NfJ15OGcaEkFzK+UzBxcrsbKyD2qzjQCAub7Q
UDYHPHmoLpj2ii2gPaWpMwqhSxsEi8YoGzkAF6jnUG2K5T+kh17czhSHuGdSZhN9
w0eBZYcWEQDxXrdFlok6Y2W3r6EAXd6Xp1tCntdlD3dSk9scy91aU3IxDcKPkSzb
DlNeEtv8FJXfyWd0TW9BCqMgqlZBIUilMTOChoFsyhRkp6gM54z962C4WRSRkwvP
A8ZfhQJegVC5Er+8Yz76ajTPbTIRMQEB0ywSbP2uspWNAR1XkVQMz2omhkYzISGS
fmVddGQIlYiPjweo8Y+2sXqmagj/rnF9XzyCYim0clSDL/WJkFEyGCtJHpSgO1DC
JlFJUxbrD8U0Gmclr/D8L/f0d1AOhzRt7g1YKj57UVny5x7RQNnVG1opditVhewO
70CBcf+2D01C5nxOoVsxu8Q6SVG9E7zy723+pHdPMkXHUoLoHldHX0ab5cTbjEQ6
5Dco6kl15BA7dt5xPmHAtxO4Fus6ZzJnTQBo71jydZIvMhXOhVZJjyytDmv3mpaU
eJAfIQCuDDacs2kJEQvnEM/Zk89OcQ4eKBZbosJ9MrD7SbIlBS7630GxeRe3l5Ck
SK3SkRNhdu84a7BRLQsrZhqIZGHcA6yco/w4S8aFgNfay5eyBzkML0YAa8R3tChL
g0WTisLHRQRkqMWH5CNp/Ukabbx5OV++TqEbpzEDuSu5BeufUT33ajF3UAg8/89k
qokL99fWm6tYyaxQ8gmu6q8+wDEzYIOlG5iD4mXjVxAMOt3WHId0GEGlMs9ILLqu
VL71JJpeZdIeLEVlqHrNal0ZiEaJHm928LDqQO85Puup0XiLYIkIlPM/Ar/xAYuq
Nxk7sdFNz1tEA0G729hSSw+mozbhiBpA7XdU+9qtrdOgq9TD2/9zdattbMvwp31a
1twB+kigghha8mgI3HujHgIH6fQF4Iz+QqxOfrqW+ALiemWuiUAqDEQwzxBzsQDy
Ka+y6RnCu1f8FAqE0G6jaSIx7cBKrdtmB9wWvbDAsDiefsdJlPdBi03pdAmPAW3Y
4LdeQpIWvBEunDfTB/RwVFkVWS5/7XNjtrcUNIizFgExHefSx3711g3ItSjJpNm0
onUadKlbR1XDlcqkuGH+WXH6UdvpLCijXUit6zOWZoJPvQUF+6GQR4D1X25hE5iM
QsSSN79ai8b1/9aqUv2k2j4ffJEnZkoL6+vYWQ8UuOKCu3+lyFge6FDmza5nLuX1
3uk5u3WXnXlSk4+YVFQQhJugbCDDgKmWGidRnZNQ0IVwduOaLv+nLpyjfBolNYsG
FnM62iE6JeFQ4uEi4NAH8Kb6yzdnE9tw0lcf1TE+BVoQp9ty5RIKoTt9hy1mVgzV
DgXrK7Qi5tcsGBENCM2POzeyoCS2c9xEfYyxPKEycXfnfIOcaEjhnX55aTJOyX8l
LDdHLvZzjHVJh8FazjY0z9DK0k6kjVYXvtM3/buceiP9OZ6O+VayktJOuC8eEbVm
2Gs5faR/ZgfJ3Sk3T80IlAqc1SHDY+KJ69S+Qq4qGUC3m17kXM3q3mYzghvo2O4b
dfTf/td5SRxGr4/JYIujcBXTVIUaOjDHB/4YE3gLKcBOkKb2ZQWDmb7CMH0lPH82
e92c5Jehp7uUuvLCtpT/uFebbU9gZKZbjJ1aUUNZisZfJPXW///Q5QyfIkN2TIma
T4lIr0KAswbteAr6rVq1/TnvmHU3XC22wJmF9zxp9giI+6KF/ERHT7bNNllK+n+Q
2yLyK5Bclqes8oGuKUq5Ts3ydIOfLI7qEAqcq9/AJhHy5VNWdCLprKDVF9+oFhfT
PKRrkTwuV17IMUalWZXqC9ZPk9daI60Pt1YcwfpcROnWwG7NcwNzwShhTrYyVydP
2loxmxR/kDb4k+82KRHvxlfbBhVEw8ZDFRTQzpAATZDjyj1wIg6ZAXrcNjBpQwAX
aBS5hxs0rLLOGRJcV8yZJXgnqYDCIxqar+lR38FC0/Mn+Ojii0DMALDB5sQeh5uU
jIbkQ+LXS8zbqwfUwU8OZVH6jHLgcBEVsbHsKhuZ/SZVbk4OemS23OR0JiwB1HgH
oJiluiqAJO2HwZ16vamnAzblAj3LGfhdXoRN7ouAko/yXe/BmE//5ubkrU2BTyyn
gHS7Gt+9XLASxcZffI0sqZ9vBU4W36WyKEQ5+MeHkG+VPw0SUiDU1iFjHMpTXjW5
uR7HgQbNUvH+5W8DYFalfUIU2HYSZIbhULgEoECXPdVebpO9U9H8rtiNeBXmni7T
Iv+vzKNJYTZXB2oVxcokPj4k21s3h4Mq2ctj0GjHuR1DjtaQx34FnS6n9dzuRYMw
i3SqQFUe5dl2k+bs2xFUFXx74twvdB5Ez3PTOKlggTNtuUDmNe5JATeRkou/Vrw0
8h1EeIEN2bHMunkvb2V1Lj6YmGJUWd1gg+bulW1U5pNfh2kBmXxyzABauChNQGFv
dfgb5XkyObsdRwPNeAtC0+PnKn5OpeqJRisVWopgnnb7hfy/NDhvtQFnKvvtdcjV
BgU87aEKjD7aa/uLdkk/ibShJN1Lvh03ldXU2rRpq91wm+HnxLWscy2Lk+9OsZrq
hKTuoTRpXZ3/rRuFPMFqm0fxJ5O7h1wOADDfHbV8bTzSGmavMjNbpvWxnBV7oiuE
KLZ0iOUwcSQPItBPAUnJsjfGB5SnoBD6o17ZRnChKvV4knNfvlrMoJCwJsjARzWp
6YzSEY3k3BGn0TfQOri19Sfd83ay81ro8l55FusKaZQRk/waTORTpBS/we36SLOW
2ZD1rIaETMuTlHsOvyHW3I6Y83QQzqynSbTFabZd9FAs/0nIyYXg055xdZgMABXj
uWAI0GvkQJ+/x6e0mrs3R85GfcwLbZLXr/r3vMMZvCZG2XErD2ZmYh6SiCXaCvnQ
wgoT89DSt2SRr8/wxiT+WJHsacvM/YsiiErRU2UzIhFgxFmuDlhWgraB7TS8JaNQ
fJJhHpU5yukj983+evSmB/ja+pP39rDnlL1uLPqP3huTm76F+pid0b355n3e5KJn
SdpJlQ3z51Y0C3NJL9MbGUf+w2T6AyjtusEWU9VwLCX0ICyb90mUFNoZgSjH3Cli
NoHskKbQy1aOpr/2vAalIOUGYbmIgvh2EHoXTumznqtg8zU4++qXCLoq5Rge28s9
kg12rqZP2JVBhsxBcbh8y+cl9TR6UawYDBmPQHziOEybyradI/RJT4qaqEH+3BFY
McBty9dqay5ezwfdiz0/xyNBph1BoZYwKL9rqskHjrT/woJfVCvjMrx95gie/pD/
vO9s6Der9xZcNE8fQtWn2RSIonvSNNFuJpeh3xPoUtxpp8S6xlgm4G1VoR9WLFRV
2x19JTTHzCTlu92REzGO6waobnkiOFH9Q04tXcFwTSYSOG1hzLBTE/UNVWSiN090
UlwWAJV4/n2DXRadFu6PnDQLJvUQ6mCvFrCtbX8QJQ6R4EBQfyuBwchpIyBCip+z
WNn2FuqnjwvPwREnbqsoyfdWWr3V+xZ8Gwiz7gfe+m3Jij1iE18j0jtVD73ma6nR
Ls4TlBkwBf4W4ByBQ7oq4+maqZ9HeLPgeqaOuFvmsM7mhf1aik8GMt+6E4+UmYPa
TXZuEqvJKwjneE4iOD7t7cjJVsLsh8iGC2k65igD9wlo0PofPUUH+de6HpkkB8BE
F9szLI9tIXATSt1D8gZuycqEiz2b8YeYqmNFvCtrzvQK7GTNUndTeEx41/phw42E
/B4X+oZo1olyT2ud3mR5AhyzLSDL5sRrFiLY9cdwQAqU9lWLa7KMtRWhJdTo0ka3
DkElhkyMaVZU8xzm07GJAekIQBm9EEq5mTdWSUpkFH2NYjaPjvlbfmibNk0xA0Eu
F1FJt85sCinVGUfSzPrdDqqt4gGZ6WgmaxnPnO/8yJNhycfOGZzQfoYR/PO+9ifs
NuvIYmcFbv311Swm/lcCHQsNMGUqBbOYNZkRkd79EPxpn5ahXzAHVF8I/h8MxK/A
R2xNBZKyWFfNhQsH7sTdK9smgRa7Fwy4RR1W9UYMNdoSnm6DIEshePPWkLlCRHNc
tNSZkEn0TDgy+gDTTlZuqxyjp2eESFIh0O/SKnBQmJEW/ZDU/mhLHBm267pyCRIn
I7IDBvrxtehg7O9CeUOklxFXMNjqLbhuUPW4DM19w98KdGe4k4aTWnnZKw80yMh6
O8Pm4z17NGW8uUjnsLgCbWHrbReLQ6PgcyrUdoxnoeihplpkq4cl5KALjmwC8PNc
Wd6zutuWwvcE/HlAXPfDMjiVhBGBQCFhrayVDL/FOB4HQ9HVkXsFEl9a3qMkZZJt
n6ew21aSAE38BxA9jFWzudWfWKw8uXFl11OIsJl71pWEzd0ATa9laCXLejojk1nJ
RQnhGoUEbxxL7PE7JaXBLgfX0S5OXUdVV+d9Y/ITWX+GRHHs0cjlvBcGizaAgITg
BgqTw6HvR51f5getH0GEUVmU/ZTlGmq0rguLL7kDbzb2DiTURBEMCC4bx8jeE4AX
PmBcJXEeZXGFzdfkdPGnluwDZi6r1lxMWE2DkqStYp8uOteMvOvAujLbgvwiV41b
dcWbJGI+kVpGRQI/4ydxG1+zRu2nlVpJuFrbF50qGhEXGb2R1xNS3JG0Q4Gwbixv
Qcead/tg7M4iBX3o64Mw3DaPNJKpdW7foGtOBk2THq88oXw1EmffaiQ6BH8H1hUD
93Oh9+yFpEFOovZFUWrDbQ1J+fhTXb3AvA/6gGc7q4qRxag2h3c3bSVxhsMZzKgD
+NSa1xguyxNTtcGVRL1BngpYbYjCAWIP6W1ywYe0F6p8+EUFr70G8JP6SyayHM9l
uom0LLK5RLWO/ZWxb2TrOTVdXU3q+sGKf4ahdl+/efTEebfo1eAjqhIRw05zfKF5
XWM5dA05kZukh/hy7FupH0vt0A3RubVzDCqovlqKMTaI9/uq92q4qZcEglEduWrV
2tYxyURnZ6f5QJ1CFuclfJGcoDRZUCDi/oSMoQJMtJpp7WD+xYKuFnIWF9LVOJFM
69NxtVAUUaDFd9RseJq/GTKBi6HmtnzLMo9lEDUwIBkPJg9gtqgSyOVfu0aLEIo8
F+qQ081dpaeNOL9YObDsKtXpjXV/XLbKi11v+jRjB59BqbN7GXp+WbWoMUlFnWaA
dhk6Ou45sZ36awnpXbq7WX+4MsTDkYttSZD4S6ELukR8YnLT7f7ptrZQZxxGnQD/
69BEI3qFxf351PjX7GQsQWTncXm+OzZiwM6UBxNR2J40dsW90UHXOe0GTAPMwe/u
gDb6Et/Pgkpj3Zrrgqmcio4AkKmdpeX9cgaQ1K7hi68Kd1GjG+P1YhIIKNJEwmeE
OEktqE45QcfDc8+RW43cLJ/z6Q7msgjAYrzeCt88hUcJdZ78892FG5tELScVgxA9
ER7jsIoiBP+8a6OwFyJmAC9diDFwDh3O4ZQjEcpiij3LlLMjNYBZy0TdjU4CFsOI
YB+G6LoUFlUDneOgegI2giVEmwrrp4/V1bOQFIF1pvKEk4lDeZkyiovrJOLwDBZD
l9ChL0wIx6Zju9HserVMa1/N+RB15E8+K3GuHOju95IqJYffoUu/e9sUblrWSEd3
jU0LwZSAYI5mGw3qnAUVk8+eM+t8vOGPJttwbHByJbwsVza6YlsRR63IpOpQd59d
6JdGkr1X2Poyr1xsIYwdf7/kVP1SyYNv0Pqt/282MZakZzwHbzFynIM2hefdv5Ob
1lPdaqVO5FBGwzOb/k+w8Sn8aWLlW4gntFZ9RBV7z+j5zKSMQvPG9W5o5/clfJp3
A9oPKwk4V7/6qUos+n1wKW2jovunYQtWyLa1tzi8KgmfpNj86CtS/Ud/Pt9ylSSX
T1dVS38MoCTjpv/TQfcpozSzObWnscv5uEzxc/fOwHnqdTqtxIZqVFzHv9qPTknU
7KfivYLzr8IEBCWWFBlzPLb0Z3PWV2bXiksrr65lV2ewit9dBlf7BnVTM9FDk7zR
E2jp0IFsPNziUBYmvuP5HEPcguYh1qQWLm8E7IGa+c0FLVVgBstL2EyOuGIrwIWY
eALOTfGXU52QIH3a2OCPY4SPnC8WEgQCNOKNPn7EFE98pxQQv+Nirw2+mmYoBQ/1
TR0pF6lZHupEBB2kqinxmFsN0/rt4Cp6Hx1x/H1sNiItyyaNviq0MhojvwdKGzos
uSHby1trwO6hC7ehf01ZKEP4yKbtJ3NmX5cYDsjNvTKwJzBXyxu8Qo2YbgYSEu/I
+UT4r3qX0UlvqV9ithRKxEjNmyiF1AN8TXi3uh1KxADQIXxHEN3/KOrMzblAFhVL
wcAKr6K+QF3YjT7EEPsYS/AC19HgHu08+ZMW1pnHweWIpy9aHO8Dohzya/pIU1H1
GjJDDC6LflbXj+in/AcyDScsiPfUK2aKHT17OIFzxcg7FA4dVeLVhHfUc/czuBVf
zXD+yWchfgENHUxO3WLUl6HliwnaClt4tIHJl7/QcduD38HBb9BJZYU8bgtTKryY
OqvVWPxtkpL7lIaj+Wjo76nxJj8nXqKgJvkoorb2Ej52pz0YF0xx4LoJYjm5R7F1
cnkTf5nki6bFbUQ0m1rtCj6+C2r9a/x6pkJm70Igfi0TSB5dQ4fvlGJmeCKaLQ4q
msDjyJ2CZTtbYSJJDPgkeyFD5Ml3sIU/+1GEViioGOGSE94GUCPjPe/hN7mpD8uj
WAt865FRtUIeAsWkQmspJXt92a9AIb6gey/vWOBJPP2+nNiogruX+FpBrq4EAt2O
7dm8nqlJjeV41OYEMclOQyrHKVg0sYiCA9lQmogexxXSt8heOa/1pCCDVdbH8ug1
00i7BDAEbIFoorDjeDQCr9qDBdTjtdU+7kMJjZsE8FZNsT2VL5eJ1VGmJ5k9SEB6
jRGiMyuWE9YtUCFFfKvIbkVL6KtDFRpFiGZfLX/xuc80qqdEKDdjlab5HvDGDNLl
4Er8mu+4n2+jSBBs6ob1XHkMmtXyQiEnpjcoNQenp29AMqpkChmPrIl6tJ2Csje9
GblgfKhXAJnTKJwFQXQIUqw333COSzFit1fkgA9ct37oyVQ/vtstyoaa8CL5lLF6
fXs1iNyE0YB8LyrR6nAqsJFBRoKastNCs2UFeB/Sa33uqPEVb12eOp3U8ZYliewS
4zB5AdbRMPXaA5JXweth3o0g09WVoIQgY8iYn7IZcIKTMGMzFKvu9o5C3uNYuog5
CL3HWUn0YDFhOXyDGAuGAKz84+Eq7gF3/J+5+R3lo4eqRjXsNkeG/iOrmkEgR0WA
MYtMcbYws49jrjA8I2m/tj2t2eGo9bhBaylLuCbSo2e19OdDwqVK2HuULhNjp/TA
cahB9kYT1bGyHJvsg/BWSC7EMmBhtNdOi+B6plV0/k2MCKNbHtCN9VW1fHnN3dqW
U2h8vsucVrlDlKBpLL585gugEhjBKE0zos440DnMRtZQpp/a+Ow5lq79Qch+AanK
Xj9aN6oP9xSth/iaP7WhPahnzvqYAj5Y6wmei/XPPuhnbD97/qgRewK1kBlCw2lU
54QDCYCJ6lEgVRlN+lT26q7mtpxSEWvgyCwUN2G9LRlpvRyuHQizL+6m9tRu97HH
nbjM3Qp1ZBrU6tvaVt1uwc/Fb97PzLQj1W9LRmu3J8drAAfoEE2sdM+PYEMPBXwn
Gabfj/NceTIC4zTeQGWeIFRozNTvReRNJKoAJG9cv9nbIExhzaoNlX+LAI9ptF1p
oRY4S3EmUOnLRqXsSSobz6HEraTrZ4WRNoMTZaWVdZNw3mq65IiB/qowV1zqRUU0
sL8q0iMYeAMrPLa3WnquMHrg96pLdOegbBh56vnvSQdQJHLQaJbHAFxEC4+ctZYa
2TAufmo4ffKcbYPplIZGc5bjMnHtGKy5UYx+sec/83BbXPk2pkHXCDs23K/46VDK
LjyffKariGKrUREUBPqZcj+GgaXvv/sbobW3/HsT0DlqxraTsQwnEQ178FyYrGys
2HKb2LtXxfzrYxzIxhCNvn2atpBifRVWvU+FBZibnNqHlKfrwlaPyor1V3Qg5PXo
txzJwUz3yxazl50iiLkCiEDYF1NnBDwnsjfN6HVk9IGCLnnHMb7f8p36B4Jlr26x
ZHZHOI2axEUkx1+kljQK2rRmUnEd5tV+QnSY4yO5C8fn6I1ljgR3th5z/voJQ+FL
ro7pNfJs+w3KNG8qHtAWVS2P+cKJ9NMNYLmbXgmbJebVDnKLX7xrcW3Wrm5nEq/A
efKOaFN0dXlEQ5WZmj0f7E/583VGhy+XwAYXRq/AQspHJI083+uzkKQiFhRGbvFM
0nZUA2AeQlUz9NQ+ct23Ctz5tja68jNuRUlIY8u3knXOKmGR3srIgIcEYb8oYxYT
u4VrShiHWfgFNDvU5m0C480+EY47ClTFhbRteR2aqjrtHK2kqAUP7O0JPoMf2Mok
O+CVsto2Met+Kun5yyzWKCWw/JyeeiFGZQUIckzf2+/oD7qAvxamT9ncTLXp3rkZ
tl+RJrxRaDaSmC7qh1U6pL4DRF5Qy/idQPOcWg7zmm1u338SnIqJFyGeNzIEIGac
l+og0pU9wKeust/dHF9CYUu21NQvyn1OL3gKFbuWOWyoKPWLeNN609gvKhWewLEw
5VNTMKeM74wWjyPLFWnjiYaaXcRZbrpZsV0U7Jzx+Fx0Pyx4lzCAxfr7GAwWPETd
KB4lyX22FjiqoJ2yq1OnwERSkHX0ipIZC2ScJB1p6V/ln3CPzhHCXELTwRX76e7G
c6SVkYJkURS05y//dZ72SVTcJ7ZLv7oxSfoB+lguP/11vsORhmNpORZhVRcNmbJz
2BgdHexjD58uGIImJUej8k0vq6Q/0nYSZZHCyLR9goJHoWfBDJp+sXjAEljuyUle
JOylOJ/4Xf1ggKvVq7G3n82ffydTWnMZgYw8Mw5Awywf5Niz+wGM63rIyW7xwBvM
wKtyBCtsrEpBLYRuD+XHte91JIFwRA6Iy1/x8HNjpTODGESs3DuU74QJ/gqI2FOT
ExMBsijAD4LUDXBm3xSwx+uCUB0ZBEhm25TGMoLrjvnLDe17d3idJyHomsr/g2Y/
eOjx0AN6CayWfbGcqkRg7e5So9urI/+TNimgklYc0em+c8Hp/txC6RhAX/LUX3CY
FccNLVNj/AT7kP89g5yTOsOlOMQyWvpwB06/dIP08NVJ92Bn2T7erOUXrWQwQwsz
ei7CZ9IoxY3rygU+Qw/YIb6vmbhaTgHxfO3zy5APUw0+V9XMflAjZTb+t21COc4Q
xk9fvRtvkeJrYIEX4qnXBwWnU4/N7ykPiMzrj1pjiI5GdSFGRxpRP7jsntQGc2zt
RSF7Il00hpoBtplJfvAw4+fOHDxcnqwptxG1U0JPDRqkH0Bvuf1kUDORNj/bf0Vg
OqV8s8ZUtxs4FK4JvN8PuN2lI+O7N35YbzLpqQ6wXJV5iVz7K+Uubqo3NiR9lf3J
rXNz1FLYoJtCgyK2KoUToAekfi+mBLn6wvOPDkkSMmUSVPt2hoSW1lK6bwCDP0dw
f4JFLvHemqNtqt/mPsb8Wnf2kbUiLZcNjEylEvSvcno4i5mwpj/6odDGYegONg+n
0qRMvL6bSnFsOsFGrV9pZzjTP3O1twtwFT2UEe+S95wamyCKKqXX1THsxChE52lt
BgZjlnSfDwzOZ0jiW56rS18w4fpW6sa9D3gpley9y7bMnRxhKCeTgfvcaNxNxrVG
WkbEnenfqwoCoeXPGUPc1OC0QmIVEhULmTOJ43ruECQTbKg/VwBfkV0a5Nchg1cu
e9D6oioBs+8+hI9uM86Geseow0sYebeajGtpV0zcQKUkOtFnHG22ahfu6tzFXljU
Ivnb9W3lMGYZ4EkfJnmYnfp42WuQ9xwIrvGrMS1EGK3rEqzwbyXS7L5YttKXMJSw
6OzS1HkRYg4gNn51iPKTRVZQBwX4kyzGA3PgftcMqcLluy87lIIdVqEzEp/yLVSV
pP9QxW+z7HiZGb9wuj1MGk51f8TB5+WpTAh2v7aHWl+J7WDLvLtqfU/7VXq4lXc1
MPCqJTmPPRxPV/T1q36jag0K1nuAFH0FJjvq4hEp632KYHqdopp8hTKshxjr2quY
2ug3z8RAEPULf7MrqoYXZ4udiX2qsp0U0uYWh1lWos+7m4fXF9CdI1fuh/T3SDJH
/m6DR9d78+XpiLS757djZTzpqdZoN15j6m4DNlGx7qE0clpC5kDhgqFB8ewTFayL
GS5ieIWte46QQZ7ScdJ/RwxzFjyQluJZoxbZGj+2joPe7PYCu3I6iJhZHdlkSvF8
8i9fpd+a9SC8VVvtZ73mjeb+CbYoPnhz4Ib7GiwTzHWI128a0NYD4cu9sKdIrU2Q
USgZRDAVovBEATiT9lmRiTJcX6t/e8EN7vVAVJcfDYa/ms+Vmf4/esSBrQX62AVn
Q8WWrPgt4BN2iWFdvQp4GGuQTX5hHjPEU+YufhbabvTIqNZcVd4sS+xXKMXkAmvK
wy/p5C64sMvcBG9B2ugQUew4PI2P0yyqWRG/y8n6Hav0IpQHzwrrch5MGWfjXZRe
l0p7ZesZJ7zV74NqmJXE5MVUs8V6ZmSZatJuT14FeaCt9H42TXTyiEBH5NrnJbbR
2KM8vlhvnJ/nSsy/+6RgrDfJgIWFEoMyFc2Q0kwlCCN4mAkvEfpaXmOXIfGxmQni
w8dPB1brGiwYOXCIpqb5syt6gk6xpv0FIqWWq1H4CIamcyKZv+PH15Esg+vPfO1y
laH2Ws6R2Pceq+rJYSQbK6uOT3e/KkamL+jeMO5a6LrMpHchXEqQz5FRueDfG88S
eg7cpigaauaG29ncwZ9vrFpyfwpdIOxz61+0u7GwWG/K2mVlUY6B8ZrKgWpy/s/P
3eT+CWE6pGY+pluKFLXoCeWbr58Cqz/BX9y0bacTrD8U9gcTMGzCjsezEqChOyWY
ELSGNfnneh2LPlP1+rHTPJDysZhTrOCWNEhFbYTRHqsa2Q9fKB8hBzwgLO08ZbF1
9FR7LX3gfvzutQKSbVDTuL49Z/ORcrA9DIb28+DnOMvGOaUOQSNGhFGuDvhiHPf9
SaFHFh7V2XMlSJGij7nipSvAYXvnfesUjdys4GWQHEsaO3Xw6AbuhB9ErfrTjSyD
uuOeEDEaEyhojfmfvNDRfrH/9fGyOFeeN6P+XS9hQVr/DN8n0CBOUaOGrVoO8Bkz
t8GxBD6UXbfilUyWmrZV+JT2xstFizcLQNIeicPwBdhgvmtHifwVJtkLi3haiBVf
hWlS4fmpnOsO6UeeCWyRsyykrO4QH4t0qkATZCBU0n8YIjVn1+jLlohaEe0IyRSs
mELteT9HJfuLkpD0rkUIr1G5pXj63lT9/hsmIK6tgDz41fFcCZDAA4HM7nMrLUic
dAIwIQFbBtpvm9mYwhCpt/JF8I79DT6ezRfa9dmyPfo3s9WOGi1M8mVFuUzp1z3z
IMgDPpUueRrwztkjUQ4Eoqy2PvyaZWJYK5qVA22tih6dwjonTvRyo9TuseNJEDdL
wBbUP3urVJJ1dOxZ7Yttwd8iHkKuh59lAAHkiRwlSti/IEE3p9sgWEUW5x/Q4J94
8dRO02a3FSvZB2XLivvQ+S2vIIkeEndtXaqodYeyWmXlyGlcinj3wQPbHF5Wn1/V
Zxavw0RIIv4xgABihzCKpask2ecQT6gVU8uM7dovtPvfxz+Gzq1p3pT7+hUIYV+k
7jFGCthrgkc4lVWkQxqPQAaBejipnix+K8GB7dBwT6huHD472nmlbOHwCcor2a8H
RexLxzh4eXuA0iHJ/5QZG+CQZh21h1W1wa0t8LrkQhlDVvJTgFOBnyJOZ6yiL8fe
tol0aX3DLUbTzOgOrmZzDIn0MlamiJFO0OX7H7jjvDqjlZhaY9m2rw3jI74gJE1I
SunQkyvNQAneHNbPdHeTy3JBanUTv+iYSyKdkIqOsIc5l9FoZhhCawek7tsobBsC
lMcxqdkCTewIVyPPCaPbkxF3Vd9nvScfg046iUY25dG3yH0TsWqA2mdvWmlX93pQ
F2pkTA1zLM8IdX+DKjPp9tcAbl4kUfGVqy9YpI5tXpHFEOSOdYv7wVWrCKF+OPFA
4Gp4lqnoSgWLbDGzw+AZQuq3fQO9oyPjp7zX0hMGjKIl+JTP8ncHzcNaZAsJ/XT8
RMo+hkrt7LBSlxHCbojxP9pFUty2X/5NRhHGHNSvWan78LRJd/OsQdIiEOiQBSvj
qzIoPwLvjxDG1WApKl8AFWyrtlKK3rtqp9YVsceOqVzwxw1dCot7qs9tDmxUNStB
D9MM+JsDzJjxG6t02OTxRNwVBG+xi4/chAw55mQithHsrLgfyK89Fudjm2dpuMcZ
7hyw4FdXLf+7DpgJgRR2IHFie+Ehl86qwX88nETzZJxgISfOE30YRHj5IW96LSns
yjLbKwSBDnWapI/d8ZIYJHRaCPePsqXOdIUyImSfKf/eQYeFxS2qkmt/EXY0SJrR
YEBC69sRHt6P2TiSLL8OfFZfwmXbfgIo2F4XlnFzUd7cld7WlBgyacR7K8MxOCqQ
u6Vcq11EzDfz2BCT0kvykBZ8hyMpzYNq+isSIs2ADnHKUPXc7A5sQPMcw/BgexGr
ym+vE+urlYdHu2zxToJcd47apIBt55nqakxB6IO8CguUciYhhdqnrF42OCfVy2Ml
eHlrKpjNYXkqSeYTwuF8LcPfW1J7juYd9SJnT4qI1aXD+n0NJuBjMvEUo0++l+rr
rOqK/6hvonZORRzWpIKfrR/bp1zVCepIo8Ks5U6YlXJgtow9z5xcKXm1/s4fMmuD
BuigRy1jMogwt6emDt5Ryim+hMH45Z4rcEV0uYICraV+EvekNJppSUcorHsYhTjN
6FLYpiAzdQecHsXIIlMAEmsVeiPLZ14iazqJSDaVAxhc0xQ9YLTrlSBBC5KKY2Rz
GF+o9my8TraG0dchj304Ag2p9g90PnhyvNYi1WTHVNvqGjtkVTUE2wAAuoHTZ/Rq
xkgE8UyVqNknOrYnXxzR1Ub1riLWMbLu+0535a6y4ZlT6ij0ac9HlumgxCrjOdgO
58k7g9DB6jkC0deJ02A1PS/2sabKEib6qpWcOs4hdA/bXCWD0bR+/JH2WnzmNd+M
w6kr+XntCwpYi3rknA0NbsYM8RHefxJVLrZ6c29kve0aWBf4fYvGWLcvMJH8BWm4
2xyxlAKvginDNv76Sxi1Fy+/dzzaf7d9S2/Nit5CxU7AMqFRTEjPO8CoaXntm1hn
bRc5kbRgqQczMhiS4Db2x/5jw9hQo/73o0gffRyRaJBFAM/+9Qutkg4GSR8oYq1n
88XkZl7PgB1CaKijN/yah9YCPfkN/FFIWSy8d+hK+hqsqzVw3ERkm7owx6GdsgSv
RL/dNoOJAckMjtSvFtArQn/77ihvZIWE1cUIYm2dBfXVkBzQ8eS91QJNV3F0/S7N
eD3A0BhASf2/Wt7x8ZZjupjX+OSnObZi0KXeCdGvV3GeUy1fvffYU6ruQNb9UobU
SqqzV23Yu8MduKYV6nFuzv4+JxUCCa8iKT8emL6+3dKVH8yyLZiNZM2iGY5g6NFa
/XFdJoBLioOlH2S9NC1Cy326flgezl4Pg8/0sLBQHN/3iJuMivHZlI2MM3I2xyL6
1/exeHBuSWskgQd+TxDvuZu2MuG865LfDwZxTbSVC5kLlK6/j2mt1NWnXp2QZd4j
/k8lUTfudijIrfnfv9rNuks2xp+7YW6QR80ZtkBuPASYJwWq6IdkwMGkgrZqwSVN
1g10hoo+tO2j1h//jviGfOGpggHXdIi2yFT1B2VwDA1rzOj3+iwy4GzrQlsyVVFf
Kao5+FNFDdtYYxPcxL2hgcOmHV/scnQUni8mUczEC+DSeGH6Y4esupfoO8TXJ3k+
2RObPpKDVx0TuAxPfqWmNoA/6s//C68v4yjlAqavEf/ZkYmAHX0Kt5anhSaZzONP
Efkoy4gksxgrqt8ugSf7S3szgMXjOeDnAmyCawEyC40IbaqCoYst1kEyxwdgD8Xz
9dJQmtW3NvSkLhY3HNpwn1sMvI/b0FWxjNTpXLlwN6kTf+ETqTNodVx2HzidnFOc
47B5kue564Fuawh6I62cTLSpz8WuEWcdl24T2prqlbA8jmfP+EKfDi6z1kqWY5wP
s3nu73sPjf4Ej0moKqOcBOjBuFWVsWsBlmQ7oCBpSlFv2z7awoyLVFI003BLlP4V
J+YOCh6c0SBrgi/l+vy8sOuk4JawFCTL/1RAZtK3zxfpyPbyaltdi99gtkERqoNQ
l/ATjGh13CpbdqLNzMQa5CzwU1YgZeJoTt5qJ4b2wl3DcbVts3n2fU8ewKum6Dej
ecVRJvNuooZz42FyVzK9iJI27FP5j16BcuO/lBbeG8jGl8Y61sPk3yn3SDmBC5tG
wbDLS4b33Eq2i/3DLInP/3cpy7zDLBAtnVoHgdVLU+4jKJ0Lh2Rpv3YUiHQlIkpI
KuDE5tMQ44bZnorY40TdHv+fJkRMy8hMSZLIEHMhb4y7qrG6h42AMFewGPY96ZMi
TqfMDPcztLnk5jdaiyD/xMtHu6uR7plxPAsNGvK7I0wh+Pg8PHco9W2a7do9LNU9
QjkLIuwuoUtGmb+rhV0ps4Yrz7OK2KN9qj0tvCNCBsoWyeQ6825LhFj3ZjJSi+CD
pixv02TuIDH31zIYyyk5IKOPS8tLWfZDgaZvZ7XuVCaU6uCLGZ4snBhIpPu+nSt3
Z8s/6MvEv5/mI9Vlnt/oBZMfe6wOnOIX8qMTIS70yPjQBcGp5QBE/cDiUJAYfKwr
gRSRPA3SO5bMmen2/9Ia3gtZRRiUcRigEWuy4jrFFeRXydW3BIhORVJ87c/VA8pm
gr7XVf4jqcZoRJa5C95xHDVzI6Mu7NSwAa8xPz/ESw5RikMT9ivecawUDJppRw19
QXRaCqVJcWSNEm+OkCifxWVN8pPbfB0UPdTligDX2h08HTkaKE01C2AF+6QYRKo1
21dtpZz+JhUQxlG90Eym/R/5Q1vTDLv+DRSPYsPIZYemQtFBc5aDaiqGV1ctRom8
coI7c4zqjQyzyAwuUF7dHPmDKeYLL2nIdw0qMK2KKVkVvSIv6oJk7CUENU80rL0p
eUTurf+CFF+kIgyrtgG3x4dm42OD8fZzn8s4aP2uM5aCKmunW8HD+8fKcfuKva6u
CrF2nzvMv0aMffJfJjEzZGg5qQBJsn/s7WbjIqHUhGW6L+Cgco7Xr5RMQiJz9I44
7ToGYYxQO/YsLpUJkjk3S9UWleaTjGVmV6bl5rrgmFsrz5RVPlXN57KRiR4VUiZo
xMvySBaD2OE5E5QEkKs3UbJsbxioT2xI2lRQAzo9O3z9Skyg/COmX+b5I8qyrQuu
6kU4Kp5W6QeqV0fAXo9FNpNiPPbG6jt3zhvgDlp6K0BtMi6El2ZAGqiG0ZzfUdT3
x+KOyZQJ8WVUQfl+EaPzmuleNTmJ+m1TvxrubHVVeqrUpj+TIXFqg+copfiWG6Z7
/IVA+v4ulLyE0tcPfJhariFQltZul1E1+MIWm05EKZ1K8XzzWYDmpfDIi87uDX6A
uzfggjZU9mYoLFPpYpf7u6kv1H7EpjItw4oPRJUnM1zLcyVL7c/4J6Bal/HXd2R6
3+KSf99zRd5nUzk++9wBIYqyyAgrCx9yLCFelCXNy4/cBD6fgOOblkH/qf1Efakz
FTZ4SQ99KQohuYMTxIcpjpY0rI8uGnwppk1TgnfPFEke3AFSKxHFoqnfHYOdRzA7
XpvIwmV++d3qGS4wHtC4EhCSqrjtuKzq1ukjVAqAAXGqrnaIgl8Q9llkkmPVPL94
ZcMJK0mPIKdC9bWnSKaDTZy6q4FYdQPgLPcZHC8/SZTnIqsvDq0ahZy4WH0zyMGR
DbiEpITeraF85/qyq4oolXAyeEjiozLN2GaQJcOI7Tz/nwHbkCWI8Lt/t2S2fiYL
uvIWES8yPqYSw8+Nq4AKk7ETvLIfwmg6PwCrjcnLRz8PeqRbz/juQyZWleM1G/7H
Y7lrzKjIRLWEwMFvaeyJUXW8+ltJePIMPdeyghoOZVbLovIZTez+VM2WQBcBSlsc
3iMTmoHNvMvhe8qjUTXhDq8YFpU1WPVVW1DwYX1fjRRrDrvSSUYow9jF0cSBs2Rr
7hybykVsIFPCVMdujjhdBfbBwdj7khQ4NHvPYM9EXwiYTjMAHeDv3ShkANehkMns
lMU4pCHeyXV3SIH02DXHYJ+QvTWuVSyjboyEwYxdn/UOkX7SVqAwVpvCfC/kNh5T
uA7Edn2haAoN5ABMSSWwk/5MuJF/jF82A0N0WMPMsZpw3qn9mVu6u0o8YHbvEAUw
QRAyb+2XMBWBJnfaANZj1Ol2eegPMd6OgIHXWkby9qsTbPNPraneyc3UEVu6bHIp
4wG+u8wLS3pY5SzleZaWrAu2vDGsjfd4izzhhXRpLMDpCW3Im1DplVgpq4FuMtMk
Yz3IFL75YygLkt1i5ol4jWLWHVynODtawcPcIkJwL1TnkaZhUlt2f5vKT/wycCHo
02uWHPGt3siDVSsB2r0hs7mt+3gjPGd8s2+kRT9H8kqgEQ4XkHOXhW104JLKTrGZ
POTorYAwVraZ5WfEz2BfYdEmIz5x9D5pUXwMc1OLWiOcc8va4iR09ffZ4qkuUw0Q
YJYqGBm2FoYxTV1etuHOaRGg+IJqYTX3GjnRRAIaoL4KZ7V+oNcBHDyFYRt575B5
+4jKYLQaTc23jyQrRbrveBm+cyR2hFqHX6ilYVfzSgxIoo8l5w1/WF8cPdnqpVQm
htYUJXRhImdM0bEMobn6Gy25b9vwuJwYVtFZauCLjibNCF2ut+fKITCJuDgM9cVs
Y++9Vnk6WqSxkBstr1pSIi6DwAiuTl2/fYfzXtOnjBN9ukYr1035ic9RQ2l67OMq
6sDzDW4dCWiDYy+W4rGleFugd9/Kzcx67SAM3vR2gWpKMSxBQgWxipMpZhPceKw9
usZSM75aX9qnjfDS3G96x/iTl1lRIFRaxhXqF8lisGQaX74JGkDhO0czO8pgKiD+
lA7BfxxTPIi+XYgzhyo5yHXyheofrN2AuBzFo6XBQqyUh/bC8xSSDFTow6TsXY4b
tQnjvIA3bRYc5rjlNHb+KySGM3wSgKyzswRs0OpyQcbauXFHVWMwCeDYcku/83nz
CCD6SlFNduoE7KEQSX9Xjc9xqXKHMOVoUig7ok0tPqDbUaag0lB/6ufgqx0Cy55O
0TxpKbwAZEfjkDwKFe/LnLVz0FfSEIqq/mXmfyqW0pMSHxbfF9qkpoCixzx3uI8R
QR9FdszVREMQPhakCTuEsGzh8h0oZeYXo9EvGXWQrSlycjMcbVNkw9xFeJ2jz89/
QwZL4o7iLlBh4rYEW5ego+lKKMMpAt94J3dL1Ln4eIk8htaBeh+ObEqXMcQC2PIy
Y3bOWTZdy+nfn6UyUENPEMXSVixr19J5knCzLg5hqw6YWMjWeJ/WFmMLGr1gOEax
uVlCMH9B0jyJRz67NYET2vuytzbpn3VRX48/4SP8SwAfHp3auGCT8NmBuSXgVhP0
7GjA1hNi2BHAQo08/VMMUq0tA5Hgmd54kbuL21vIl+Bdw/qSWb4j2mLNTmyyAg4u
fmAfDvVkxibJESZavX/4PYHRVX5XfCFGFNCKnaV60TizZbq6/EiRh2eIXFO72OQ+
tTHex7ObvJuHXmV/mGxJ92hHZWIKgQ41MkQkaBy+54QhQCVlPzEpM7nRtIgBYFUW
kgoP8CgkGxjFvZx4F4rGxLnZr8XV43ITJPUIXxGV5itSwSNKexT85ngyvyaIotKo
7BQXC5mM/2mxLJjsM8NRk1nWv+OiOrK2LvaOJTcXQ1gc3SU5cFSbhVXkvhwR8SqX
NgfjqsVWoWrK9kdZREtVops4y3CpCF6+qTXnr0i9WO1JQMf+mTUgxTh2ojwkMQaI
9wPdFSVTURmk20tFEncc0o03lgHavAF6NhKgG/omdPwMlfl78pQkVIPIFFBXh/Mx
mfKx8WKE1B1dOtqvkfIcphJKRycGQ9SHSd/T0iL1D93LAOtNIhtzQQVdQO1RUFiq
+1Qc5z1uPJb37EZrk8dpXhacqqrR7ONRjSmz/1cUG17kO1uAnQOvSUEVgtINMhxi
H1+QgvZSz4+WITmZzJgGkvZByL8fQx6QYElrRoJNLAlZw9sDOfIbr7+MUH/uO2gT
TX/zroTabjJ28BhUNc+mTQB2T8bAPwNn9YoyQSA6tXPZO0vUbLGe8yEBqI4qK5VL
k824R9Jt6cRuGaihnOZi+22Sr3T7mIGVnXTzjntvPa1pRezGDdiEoULUwBJFb5qN
XS/nzHdkgzceXGMEfrPjlBI77/WV7bOqM32shPZ8UkQKmuyvsJq+vbWqZFKXUHxc
vs4ofv6Q/Tr5H4cOMWjwCXtgq5olPuJdzgWfAfGpvPQQ/NqKr/f/oT/WujbZv1+p
Ofwv3xSpwyroi73VVSU5oegGtmuOVklQ9DfpEbPf1lCU1Tv7k9azzv9PbeKPsv79
UkGyqzjpRXX1m1+g3QUB2TrgIkw2N1VyGnzDJfpLtvFqBWo+PDACnsviPOIrZt/U
G5RU9a1b1nfg2HiNRNTj55QsKwjulU331OaTuYWQXMDJzkBlL5iDfOYm+VdHyZl/
yS1XfEQeeVDKcjFl+kQ5BnU7hx8egDuwVbhWwNX7WlkXI4zyAT8Cl0IL3O3vZsQn
VuckUVBWq8zkUnzXBnYP8m8XaD/ixZmlTLhU3qJ/xRHttZpaMtdzJQ6Sl5xeUTEG
su2PlC78cO0CsXbRAbq+Ca+OVAhc2kzvGsVWpPX5kedy2GgKKcOlEnoCHOX4DwrH
qi2NfCzJb6AMPK1wOi6Xdx/dwJHszqlNUiDJPNaOyBkbjSbi1P8H2GFm7eQutGTi
6dHGcqNVBwsPxIiOHoW6sDiojkcIlhN8rAwEVamIydUAtusBtORJj4aHYw0k8hhr
//z6vg/Zn5304t7LZ9AabeIiiUxDEeDJrNUOOpQRgbvWTBg8//ffdR/hCfdRb44b
pl+9lsDWZBjraWa3T5Z5Dd3PdwqimHEA1jUQbk9JIhbXiPz3AkwqePjjBbd8lrXh
YWHBZTLowi1UYlv4hbjZXQR3nl+PkgsubTFqWSG08CPTHfdLBFD8YkW3ZwOw8YO9
N7tICnl/ajR3Sf1aOx9r9mKv9NFrD9B9oLDp27w2UKycjGW/zYkR6MnorFfioMei
tTbX2f6mxvxxaF9V/8sXL+iyZqWXHUVz5L0t1Erf6R8t9le6PT6u3/fmCpE1+Vm9
XfiqyUATp6t3DzrPX3C9ixgJAlZck5/ejCpFXYbwXs9yFjLOhenHcW9Be1fDTTlV
W88qP4MpHcIA3Or20rQothV+U4eFS3ZHxJahxBa2Nc1R3YaQjy43ODWuPTGycR07
UGrtivwvzgiJtMgGRE7BlBtX98hZZHKwihr4P3Zo6i1Z87b+POI06NfT5c0DQVUG
tBlZkUIsBVDRJHpA2th/6EbpKZjDjslUKlkEQS/sPBF5WJIC2L8aPxfJeGxapoEq
5hzNB4eHAFIQyvggUUC8SPZqp5PUJZOi4d74y0htWyCpMvg8s1Pt386YZ2cv38d2
INygK2aeX3aHvau4Xep2ho3xZPKlA84uycI9zGxHt83r7gOcrgomA9uncM47yjA2
lw7dBJuVSv/0eX80D/SFPyJrq4WFmYqaL5mYA4G9duw2JYZJ+lcpNU0VQQMipkyX
TXUBX8VpwClSz3mKFnDhr4k1KFwZ9bx4sd9APg7ft4DqLRprsAgNyLokoFfIOHlO
/lkV80YoT+Aw5tZuerrnYNouVRT1gzXCta7/XvtWYxmjpsnQGZpt747mBJENRYi+
k6SCScjT8k3p0VcOUQHiK+ZZaRz8DIbrZ0tenOnUnWgHiYCXSNtvK/mwJxWsofbv
bgGWPK9EtAn2Nhuq6JXQa8Sp++1HGeVZtn3R9Zb+wS7/66MFYdfvOZKqZikoYjXG
1U6GMKQBmm3t82t1G7SDFYGZe2NkqFI3SmJm/S7vdZZUB/O3/h2pJDiLmbeivtEE
4f4y7i8SrA7pFdhCSPKmnU0VQz9knoj5jDDvn/XDrvzP0ETqpeX/SyLQfSqoZ6Sc
B+f8vwbOItCTxpfIfpOYVxWzZjTappS7Ula+fVlHcD2v1moJF3WVHmfZakgHBKBi
N/vWYQOmk/TTt5+WI8uBD6XPt2E9pJ4EipuGTf1QCad8vjv4loXwZ7GE+I4jfQlQ
V6Lze1Y4/Z+RtEqKfB5F1tcRM9hd6IcxvQIR2z0nk9cTd44fM8kZaNX3AnDFbZlN
7eiwHpK9IC6sgi7VugJcTkZqihEY0oAuudSdFOnvy+/xzW3jXYXMkM5uGWqUgdWm
2cwq6IOSFyc6rsPS3mLwgdf+hAYK2t3CfTzaXZrb2MIi3RlWr8Uw80NwIUV7UN0O
dnYxJF0kvNMNziiOZ/3Gn+rur8SdcHBg6L9gQL/7nWM2tisuEs36TR4T1Z3Axzrt
Vm2fxNOb+ROTJs9J4Q84jmp3He4PoSykmRvGTpgIhOKJIesFA1xgVuGeCPUImZQy
UCOlmOk8z4fXoUmJyeEyqrBApnpeds6QkdYbFG8URgiFDwGCgQqkc8M+2XPPsmQJ
5QD2d4sOA7b06Xe/iKx42TY9/nMWF6AveBW2piTRw8se6tBgtKhHTCbfDRWZjaBW
bGUM36vC2+LqgeaE7+ZIBQdlcDkLz4g72PpOSYBuFfVlq9aS+4iW6uQnd0f1OjFz
CFUmExpMjp/hbwxqQF6aQSmc6wvkQC2zxNDGZ1MX1EvtWDS1Di8vcBNIztfFEBWW
7OLnmarBlQQcvij7OjXJTGtl4SV+rrh09/wimw5m6utwAXVhMaPWdIsGX4At2MOx
bOVUUDxvmhRFuMeAdk1Njk11R86QMpBGjvxiRxiALDSEYKiFki95BdfAobWprM5V
Obtz7g+1gvxb+x7rNEz1CVHM/YVkjRig6UcWesvCEUDsgyRdyzxreiZLA+XO4MlZ
LlPYnFQsz5ri5S1kKHtaOoiCAwqFfIzD4LUlYOTvr07CQl26cz/L8/ouXD2sbPjU
44SXdhSl2UM+5w7KKAidqh1W0PPI5kRkuVGcrGmw56eZIxKYXcIrUYYiuOSNOdje
GxKNTASQAyzEAjCwdPXWiFxpYjhYwZjAcZKixdXQu63p87kc6nVZy2uHjadmbXXG
pFvjmkIiXXhb+wbzIO59AJ58NEFLv80Bwi8XUchZ2gifsrPpJ8gw8YyF7l94U7KE
ZhniFnouBcozz+08BdlAofMASPz8jZ2POJbnLgsNthKTSfT8YTW/U1khY9bmc1C3
12YALMJNLQ2cO+HPhqRsuiK8xacLtobo8qwL034CJAjLGwy73xBNsE316ZOUKrrH
3nXk9JfwbiJGyxTzLW2fHX23iDr8EuhYAunpnj9O3uYH5jLupmxqRmbFm3oX75Co
h2K1dMxeoaTMrIrwAs7Gq3YCMsg+tKXzMA3BOldDwVb/yd8JKHfuY+FOGeZfB5VJ
ucYkOmtYYy+rjqeiY2m0VlxXezIqDXiY/LQkxsLBXEDSp+77gq4KQKIdpqqXZrhu
UYi22V+KjbAtAR3FlIgFxSqONkElRFRoAuQcZerc/FJ3jf/SPL69Xo4zLNPuWwVT
JF52LqShTZuVIiHTKXgtxkQLN1y7BgUfZjOphkTOCSDqWuyeTbVvYXp2vmv7YDeM
iaOqtISkUqbIeM9kWlXhU6LEeRAybq0LCnmHnonmb3aZAP2nintSzKjP87dvjeaq
1TjwaQL2arbcJs/0rJeb1z/rKDZfHTsbDjG7brp84kO3382P+WnH5o0MrKxnjt/D
Tsts1Vm5cPshcaWnO9zCeBwBby2MvLQCJoK5mM+HCrJfnEmpxXKKOhr7+v/1cuqT
+LxJy4EuI0aFy6Z21C3qX44l3ij9sWCjUzss5AeM10TP+tJguSS+GFuETAhAtBrq
5Yx/zb0p2lE37no8ZBbOZSlYFV7VsilesN555ObCltdnb8FUD5w08TvUkRpUUt9d
2z3L51l+r2+SPDu/X9Co0p6D468072pDmmzLoozqzIGEFxK8AxP5pkXcIac4WNWD
khr4xbkXh8/M3NUPoEtRYOL/KamvWJ9soItH/2/ih+SlFotONr8w2OoKCg6IoclB
BKxbxl0Q4AyU6rhsG6VZK8khERKcaXwvXIqAIuzbGUiZqQ4DDqxdWNvL7HWHFOnT
1MfEEXz3sD7kyA5RI+2nL/hIBc50t9s2augSEebefZvu2VoCqq3tz+ZlTFdSdxRH
+Vup/S6W/qB2p9QGbqCcx2nYfewmY0Zlg2trudHP9NFk7oLomdXdu48Js2eD0i9E
rdhO7+u7iWv5jCiQQH+UHRDsINLT7Vl/tPnYtBecErmZgdXL7lYPbEINswKObbtz
PUmjb1UH2PRXMK6f0jSFgxfC+mm1iTg63hcvk++rXMIpWpPHaTs++KbfiUWI7Wdi
JMlyG+OI/GlERTr6QT85SalLEmBSGqxdnHL3/Arv9wz7rIUIPNM0LPngV1NwE0p6
+WdSPe4ZaXewWOFXjdiDBFuEnOrbx1q+Vo2af1wjRBNUDs3BKVJjZ3AtPMqsmaCL
FksbOml6g3ijN9vmd+oLyqm8j8byKneOejVY99YN/hoANjmN9Uaz4sjswPzMTFa6
S3lSuLrzAZVeuhCnnxbBOVtFkRbS8go5Cgr4FiNxhZFa7gkBec+Z9Ci9K6Wp0FgK
1TAfA+wfX+Qmg296jeK/rFAumQKqUkWyIXOu/ufnADCP+XWXAZKeDw7RAUC8Sq58
uX18uxFZayeg+7RS3Nh9Ci0TKsk/JHEf0JbvNctAZZ2wQ6UMQOP0PCiqkcfHBd/0
gaU6+HZBiVtG82JS7yIVW04lMaaG++qxzW3lb3RnKLRNSQG/tnizwyMOdPm2gmmJ
QODVUpamnI3O8RMuIbiswEbutO95l3cxN2y085Wc2BNBhZ/JCsz/qLaVfLBCApTK
CD/mISwQ8C0mkbgB8GncqUHdM88qJqKi4+9CxPypDkPE1LL12zKKja1bIUzmOwm6
M2DkkQ9HCj/TlCGiFkuwkUmalLkKQnjpUwIX7qn4xqKfCZcPiAyxgIs6DW/pzspW
1M0KeoLmkvVxkX/gljBlcs8CIErPyT4OIdaFuQskgk0lDjfGU0PZMhgtRBN98jMP
YWJQH8HZe+yao96kt4FPEguWhzxBTXZPpBG2LWgu/ZpeP2likH5NOm28slDcDp0y
Tp1lNEl5mday+vVZvK4HjXd2QS6xSYDPJ870BuWo7Lm4I7GDo7yol2FnbooPrcp5
sTudg6nhFCTSBUDZccvX8k61R/bbPWn9aV2k4r9GIiLb7CmyMiNlD0/WRa2PLLXx
olUv34BIP1NOT1P12LOadCBH6M7WsMtzRCzVXksASH2OBduVoVkzo3syYPKNcSEC
JKgSy7Cikt//sAfE7QkycgXYYiFpnOMgTTNZo6z9aFM9Os/2isZyn0pFwPyv4Jjl
p4nGfUbw85F45CIpKIZ7fHP/2E/mJw44SYjUVugPjepRsQ0+6C4VFU3tSxxr/dMc
+pNXq2C2K3hbnG4PBZklIj7BaDmq4XPGgP50N6BlS/UXUaGA5OvCx1rPjQcSU26v
VOto9jK99SFBWMCICkDhUPoat1wwNmbxpEuKhALYiIdGkLWta44c+m9v+jrnMtqS
0pI1aiGZKmRBBqZbFltuCyTdm3ukCEKTctSGoaBhJgnnw2CjHyk7/2y08GJfH8cI
qynLphrWzeOHXWG6hKCr6GraaLCQZnMBlA5SykZ01LZiyIZGbG/y3oe4bS7uciT2
0Ax9N0PmdfT8jgMCMansH658w9s3zjb9GvCMXI1MPXkSEQLMng95YptuGV3T3m+1
7cn2SwYl9I0o9aBteZiyzztgbcIfacQOaVMvjPw7eiMV0/Z3TXZffeVnuWwV3X2o
EhVwwSg+0Xnx5Sz5wmthxRjMGq0NvGxTTYYYtXToTA9U6sMfcCVjc3ZugBWtjGfd
itYEB2IhlehEK43Iy18sjB7/cVsTBLqrjuiSvLjXJVpL55T1xYNrRfwMaSA3Vz77
CTj4S6R2YRVWooQ57RPUMjPDJ0CHE9uJPJZtJyABSwH5ppeZosEdF4HmCeOV47gc
lQ/8e6PwJUfIs5WPG1uK956LCSL5XkiOlQ5D0D04wXhDx2mdXOYhFLUua3NkQcsA
f2XQqpbdiKVIWDvF9x5JOGKoKO8tm61jJpg378iUKmjMom/kWtlH5BPCb+w01VCg
eq5N6duLc+qDGDQCCdYxS2imLlHrfk4iQxqloYjtSqqmCv2elIkubPpNtyGH9Z9r
mk64sWnLhY3VqBnEVI+xLPfxGiahnOlOjA5It8Y1w0c614LbvrfnWaNbEAOXGC3i
Dv32JN0X3oPWY6l6A4TmF0Ce3ni7z/EmRzOkkG9xl5DPSLQFCR9CXtHHOaiYRWOT
d1ohwIpk1UKlU/aBt7fUQO5y+onQyr/bLmK8DyI6Cw6vM+C6Hvul/gm1Lr+umeXl
7+wvv+FEF2ZjGQpSbqdti0mRbJMVsgwRFJSMj3b9l53PtO4Oe0ZrfJL5J8XP1emg
iZxEaURfCC2yg96Kc+GYvBmZRAF6JRDC65UcaF3+KzZ0xhyI+VTMmGv/ae1pWMFL
isgC446GmrLLmYqDQvhbs2h+fYSpKP8DkNDO4CTYyafEODkQDLny0rk5DPbxmw9+
ggvE5EXnNnNG6jF30zXqq0rjh+ASPWNX7wnDL3+dMsZRiFxeso5UNiolCiuS0ngE
35ClKffeljrqxf2Rilomn2+NC/nvxURu5NiWACRj4zrvBVdUIByYUJpVlyovWsZm
0qotzppTuhHxL1WbcTaxTTpuUVQJIxKx/2QyuWzOzhbsH6og5RgzSIj3NSQy24MY
W/I8geOAdXvdu0zWIsAS+B9a7Gde87HkBefhLM9wlyEZBoAb1XRZY5RcagieH/CI
tpCa4MyniQ0Jhgbd/zYOAWCLESV5czYIUv4oUa8tMMAnR0Me/F91jzaP4Yc1VsW+
9amqHLs27uw/2CEQz0JfjeLV+Mq5OEImbc6e/s24D3oIIR47o2WtqEMh2Y2sDqGp
x1FmEkJg17SfqhdRuZLZEgbdx7Pi7FnyfVlWM6VXiFsTj/DzqYkGSyirMRyRuR3j
cxJUZZIaeVqXRishOaFY2fZUv2Igt05jp9CKumkcGqrUpuAepgLXZwZO1ZwG1bxJ
kelSHnbfkzPed6SRQvxaHO4/Ix3xxh3mtV3N6JbrU6sC+k2c05l2fnZPdhKA0Wy7
7T8PwPQ2Spkwu5fiBeeFgb8hA7e4MjhAZqIqBeY/j3KgV4aN33dsQ03n9/Gl2wb5
ywvvnuu7/wgJmA9GmXvhbKU4NOvQbc+1DL6UG3XRqqmhjoYOAS8q/UE02rz6+3AP
Q9Blyntdshowd1Pr9OThUCC9cPNgdfxqbZTX9fB/5IzxtV7ryIJNhqODOOtY4FMK
20/vRAY4ujOww9VCs3UeABZkULVtBo7wOI2TUJn1hEOD8iMxeMgixr903QbHS1pp
zzoGEvTqj492Ahj/taSrJqDRzDDfBL1h4+kIrCireapbH7xPYIP2PXPjnRlk1KGk
HO7I2cBivuGk564vFUdW+YRdWb8wtIVxl6Z+UeaS/wRf2xlVfGeO2Nd61h1lrVTp
bYKgKvDI2UtMtV4pfIjWAJ5+RkBWOSB7GQ0Vgi5lTZIdPNULr1RzI49rVT+8mi6w
qg2qQ9VaWv7X/X9IxwAXIk/oFKpHt+ma+kUB5uePL9ADjPmKmOdotFlA5iHebGT6
MmIcJOsoZgwrH/0FCpsLmpV3GMJSSaJK0ydMtnyg5RCneJAXg+vP+G9rA/jIj+b9
P/A/AfxG0X80Gwp8/TAKEKdtcd7uyaquIbgJYkebxMDPz1va/HdKOnM6I3Iik9DO
KZFtIxxAlCUx1ejLvI6gHKqchbpsDgA1K124CjzdO8lxnekbIYg0WloJcWB2ZlTa
UJxnA1xtuxDgfJI1QRG/PPG5zGaovybIlonShUbPDe0scpyVYw340J5CYX9NEki1
uH63mVDyACAI7Tv/jtytusuXbhpmiIAJq9Shrp7BY1iqNNg1MXRYAMpGbHYJBvxb
hiCXy7qQDQV+anztqYhcvOqEOO7fsthx+n7/WFAJRiq4gZDrOO0WhcphpwHm8uwh
lq+SRegyXpw+bT/p+R3SbqqegsMgCcXxkjDttDUrUOBVwTSzZVXnkoSBIC8oii76
aY3xj9LmQnc5YGcaYGJjgQu4YacpKgG7hZ/drghiy7XVCxCzguLeXJ+i8a+wdlMz
rncLih/BnKHwDXvXLYt6Mv48k/Zl2eGRNaoLDoCo+DJRGK2QUJpGMvMGvvVTsM97
Y2w8uBOvleZXkCCqVJzOI5xLrsT1U9JTjDh3MlX8v593ulAFi9wAWOMpP86os3Y9
zNdBdAxIS1UNJ3xq2eAp5TuAlD+mTzO8++g6x9bTcoAEnC88Sbzj36czKTAuONqA
IHJHXFiNs21DfdjysHd+gC00zfCAvf9Z1MX+XnAjkPyVRFy+fFPBRESPWDKR6Old
m7KFE0MmgqPU4HyEoisJ114gqdh2G4DhRaZZ3GVyRHsg8LYZK7nlDKfygtP2Ozsk
hsOWnG53m2ZTvNyLtqysab3UUMAc9ZEY+LMl0ew4h5cuJmIorQC78yGsdiTWJN3A
qXyCNIq+nXCpitWRkOggGAoVgq6rqmcu7TdgiLWlfx7VUgpTWxomq99RkHJXfEBi
UQPd0zPxPQeKUMktm8/hEaUIcztabQFuN20YwNQF2UjtamedLih8dd2hb5tS6Szl
pI32sbmCN7TXCtCGOd9uhSX8sq5vAoiWOQ0dlC+A+8t7zMkakKSb4OdVje0cO6AX
a4/DW6FBtP7oe72IufgYZatPUkfJAP0QDvKUtWEG6zij4XiLfPFwQSJB9ozSzBOr
D8FDxjS/TG/SeJYtvxyasIiKGcwxOTxeb8I2KQIMQjwhvKE2Gkj+VlEOnUxLddOe
W2a+wOa1zTozHj/dWJLVMODgQswH3glQX+1YECLWPjvAGxZkLHlC2RfQUs9XyGMU
Am9CoUmkJeSAFmuNgYyVTXPy2RKrwCXjJqCl0CmNLS2FR3IMVQ1K2j1N+Jv3GuzI
6WM4hfp/oCbLv2HY9MVCoC6C5Kp8uUNwbc4RWud2CT61+BAZ6VhZRFgLhN8jzSlr
y/fePm5fWEavqxbCOeRppynQ7MQtoUwkQMXbMJft43nquLlf4lSj3zn2Kh0LqhNT
OOBwjl7rl2v9gcvIAhkZNyO7GQTzH6Zo5nZPrCV3rJXKQK11fbdtUlI4eDF6qcVA
KuKNg41jmB+tq54ryi5bcmT195EU5BhVftz5i9BhTleCMC+9AXPbtUNZ1jid5PRK
MvBvKQlRpKGFnkXaVHFKJS1eoY79O/mGcirqzz24kFE3CaD/5VFUBqO1VrVbVCs4
ZOLLpaVUGow7tL6Bb1pxqKcZu9St4e56RXjj5DYghW5JE0lrJhgHT93FT/cjUjuO
hekBARSphCxQmUDJH/BMU6Lb8SGnQvvNCD23HxS/jWMHODnh3lkfKp2EaeJYSGl2
zhR1/ZiJwXdHGdg3FwwKOzPVQE+CK3RXsDoZ5ax+/rjH+/iGIm6eJcxXroMCwUu3
fFyZ3Si6nNiasxdOzpAi3ZNiaEq5oBSx2Tm4CQEjddc+3TG+RAFba/kmj5m9YGZm
RlOlAIdo0FowOAL4pcwd3w1s1XHljHiRxtgpEZtdphuwGWUfuJVBQx9jEXVx2bKO
n1YJAwbhiYm+ZC01p7MRf5KZsJn0k8J1hrOx+VtWCvWNbbRJVpsr8eyCoERTYHyZ
sCmeACw8FFRwp8Lez7cWRolphTStabV8tfDNrRQXSeKsOUmJw/3ALKRPliBgxmti
r6dZRz0x7dw/8H2lkT099PC8t8mORk+Y66qDtbzfKfbf1zgcHeAVAnmsib8EQ7v3
wKUi6xZ4RmhN7jhRg9PTQ0tElHH0BL4JzXGMlXUgE63B/X60KGXYEl7YIBfkp8SJ
/eD71/c4ZksOijMrM/gSgDkeT4V14X68WnnZUnz/MAABRSqSjvD6J9QUXriPTaYm
q1ZbVVik2cTUv/4dSk6Lpzqn1A3SMAwFtDDnB11KLHRQk+bKSaxP0SyYJYtaCxir
9S7hHxpza+NORfusrLuOeGXyi8QYj0F0r+WxBM4+K+ddYP93McUP4kSEr3x9/tnE
RRPAhgzrna/FjGgsHUhJqr/xOpgRtVeTknkUZ2HZIIcj+2IthqTxmnkuL7N99U7o
O8I5ABOVN/TPuTHcxYKDKmVn5vcLJIezHG0FdI+0RnlM85lHzGdEX/BoN3sSzYAN
Smtd1CrVhkbmRJWJG7vnIUIQH+Xw+6XN8CFdwgF9eP8uKZBaFOrDUbNIatAGooMC
0See/aj+VKgD5juV15UrroA4G/bn2Wqh30+efe5lUHNubfonNXPgcKaILmTkO0bJ
0K8/ll0eEQV4DnW8FkBedjlu6UFaVc2BLf9oi5mDTPHVC1XT0PbYhj4j4YSiqg1v
4bhe0ig2QriBGTLf9Pi3IonSaKx7pIGZKTdCxzIM3XLklXUTS635yzwoDOLVeA5x
zkL5F1q+AnnbhdYTwzj3T6mumOPhvIfGD+P7SYAox8RRZOWyiC9D3DdHSgbOvorR
9O3JXiY+RloV5imzlpkWBNhkcs5McJALWJmNcj/C/COwtyZiJFZTAOZi5T/s4wd3
oiqcdEQFGOOyOoqvq7fNtBwQKD3/Th1y4PGKUCXSQvGQSsjEZPS6tLImRUvtwoUY
mPGgeDKuklAxB330RP0SgFLqvXEU2mZJOvDCOf5s7i+EohalayXyMNlsM+qhOOMT
VZ/Om9+9nmhqlu+3XeO0lHB7Vgxsm0amQsC3SGJpQcpnev3pqRs0dc3YoHF2awtb
5ebHXZWyoZZh5aCrU4wRHppXp28we8OB3SmMPrq93pPIbP29h1iV97Oo5q4WYqO0
xKqfNFtdP1NPbZ4RycWCETCM/YpbzN+GXkV9YIPFG0XHXr2lJuqk3eDfHKXLEiVo
mWs2BkabbN6W78E4I+i/IHMl+fWcgmHwQUeft0awkNqucxqZvSgB0ds/IQWoMxEI
bX5jiNohkIW/tuesFBvYawON4OCDGkZLG4lDm8cfW5uL3x8cOwY8+r0T5GqPKMfZ
vdEerFKpQn/WW4+c9WgXjsdpeflYeoFnrLMreNVb/6NkasbJ0V//CYg1gVBaYaDJ
Zv6eBbldAwBAzaS7sFggyM8lPkt4QJUTQIoyrJ9uIaNQA1r16elPMT8DsMaXaZP7
O1G49RgmfZYb/wghD3ZOFOZwY8NPN6z88pcPJQLaJOqd4AQstV38k0+/hqt/5taW
/CqQEWfYPfmMF+MS+POiDHfYrUAo/TY0GQ3UjFRZCFXRpzJOg7/Ris+UZrpiOXaW
jVqH9BT/W5GQ3y6Chyva7P4d7ZA8OtwLI4LrZnIL43Kr+FyjYUzWD+jbc0BxSWxI
9uJhFOSJN0v6Y5Mr6NehOwzkyWS/xLAoVR19rjEKPqq6T1a5kLvrIPkCV50XJyle
7aC7UDamKRp9hRPmjwmUyNb4nZI0uOOIRA8rX/vZLRJngeDwAiYFBGp2x1KcfV3u
fDOvhBD5THfd+dfVymzZ3F6u1/03FxngzwccR0VxHuFFdr7HV5RVb0KFlL40nFEV
Y7It87Mh9w9ndtg+e7JzrDStSSjtlcOxhxFx5kKSRCP77sI54sFA2OhJWzoYUMdU
sZNGHweo9TQAuRUYRFhwdzS7Jjm1khorP91PgCCYVoPYLSQww4tpZg35B3zCwl/Q
XcGqkTEbSCc1CAoAICNK01fuVzRf5tOQYs7mcwq9c8a2Z0pRPKbrypzasmg0Xpt4
0EY19vU9A/P6kAsKhTGjextoZWOaMMqZFUe5/cM1vntknuBwBPS2KYPtJLCZtv4T
7QD8IFPSn2N63mEYb8p18o2h4Y+V4ugqGcjhWzAUnwH5Pp/VrE4cLmPVtQdlTDQP
9CEW34HusVYhlviYtHm6bslO8u+zpP0JuScUcIifZ+jIgdNToCkS9ERQkMazDfZc
GFyPc+6cmfotur9SdSbgPzE1jJ5/JjnHRbv2/zzvs5x549jJkhJxKaL08KbilwlK
lh/Djqu3bc9sS6KT+IdOwydOoeJn0NAQ+5OrKd0Z99FfzBKxYhQ20xQc3+yud1nC
0NkNxBfNKjIxHnG5rf1qj0pFa6Xs0gDOOZkGKrlIr6RXqNFmdj5KacdVyyF4dLTw
NOclAj5jA4n/Ue1mqjkp9wousjUizu29ZVi/Nm6kYR1Ig2UXDJ0Le14D2xMqMRIR
hAJdMcOYK9Glv56ggHpoEiAAkMG3f2ASeGLwJtM2BrgfA40W2EjxQvO0aBAN8KV6
n61DwUyfYg87JkWQlm75Kc74gUMjtOSwzjQ/4RDeieLbP3gPdJeAzbZuXfpK01bM
maOEK9R2J3cpAGD9V/EPoyoz38JVSt4M7qgFTQXzSKvNn6kpLhF+zyA2jUcROExh
L1o/Cv+FAoWc25z5TQVB71L79uYFjGAYsJseiU9hwIiNDWgfRHUiUu2HgGnrseTU
LeJ5Hx8wEETR8svh+Sg6PifOSqWFG8zv8rAn7wF0vJWNHo7yzeSg5ItVuAoa0kch
pNrM1Ga2OFlg+8xO7Wjx5IGBftUMO0+50YMcN69+W7NLpOEwjSIgMAZzpZvJedGS
EAuXcMTSvVhwWj8vCenXY4lmQDiTsaF2hEw7M9zMqXXGkhz+xqAg00bFTeaz5Y1s
SJcV+1ou6DHEoRRLMEIqGizv3/7rxgfTg7wZacmhQ0WqeHMjvZcZhHLv0ckpKA+8
liQ4xj5XXsP+nca4tTQw9KhiLvW+es0vAUGE4YCKHEcykGWDBfw1PODUXp5XZxgi
iNaZtHGYsRQ0nLEVpTIpDr1MQO8WbhPMn8Ty4n95F7C1/o3MNiANbrqX1AIfD//w
ewGMEnCuQPOs/qrlpsLjpHZGADbo6KP3dmpseLgFHPRMywlnqwtycBIf4dQvc2ol
Xs4caQotFaRge872a6XtYkjYgOZErlb/wy1HaAm9fowXS554TJBAOSpjfQqA5c+u
BdidOSjGD/413Ky1QgjNsKqNE9XGAM3p+aQLCE6fOVf82M5ncxxJELUncZV69SvH
vRKAZJj7jzkhBeXNR48Lz68S58zsj1arufZDq9tuIabifV8AWZ5oYDuLw5NblBgU
kCePl1mKk1NvKuIWAIjAGrbQnOyQGLZXqn0s4jYFudq29Sy+5p/lnRYzmziUw7E2
AnTfPWFTAzumG4kRNEfI0d9b6SM+i5/kw6C2qRg3frLhSJOdMd4e9WH2Hq3aiv1L
pLl+/YpRzOuACkEBGOSlAMO+kukAa0HBnv+bC0iFb0VrzI1y2gRq21j/XzKk4KEM
p8lCt91BqWQst+zTXZSskBgmKkwVT7GpEAeHtPuv0h897jsGR1q0mxU91S30emjp
vpK94wCtsdtKe8jVEFH3LhgMcwrt+xirpRNiAbD7IVDHHgQAmRv8rUbDr18Us9Oh
svz4f3n9d0vGiQ5LN+jr3cYjFAiQaB+6S7YEr2vf7Zsw7zX+x5rXv4yT2Jj/wCg2
GbMjxoHZXx5aijCTvEz4PJ5k06gsENW+0bIvFIu4u39jE5VmELJX1dZSWSDfgUut
Qr7pq1eN0yQ91acEQo0G4Emu9aRZRevDh0jaNJcWII7BAm/E699FeW28qQUTmdzt
up6f2gON5kf7DT+MY2ox5AQpwhZ6jfwjD4iGLX2IAEHaYQTYSP2bcEPjniE6xUs+
Ka9CuS5g9b+Z1GOrvnYfcZWC+xio5K82/nriaPIfFoZFVycKNCv5Cv7PqGPt5zib
/XJTsoxN9o5MgynPA3hbvL6GOJQM97sMTGEeNkzihqK2o0CVBRYH/Pr+BsIsN84B
YNIfJjof6768BJsETxfUXUETkXMYcwd2aNTlGE/y+LKD2LFE1eJOXuOCOC0PLY0i
5LLVH54fZXEd2xvXyiEwy8DRVACDKYctRzMfnu2KLls5CPktCCD2sWZToG7fS8uf
0QVl6zkGiH539gjYUzqc4JsN9p20+s1PX9Pgn3YBcAlS4Vlw2LLj2BDjuu/2Yucs
9D0el+JhKBVNH7DOeQmBOnoIAUyCmpL1/bUnN8Jm+wmzJLL4600Tojxg6C9830C8
SOJqRvM3r929f31S+C/ovT8WXz5jacTBk1E+TCiLHQcCvuhjZwzts2vpecZOjAqz
c3UovIZ3aGL6Lbgw6PmGkRABXLkG3gAGI8486fZHESbfePnz1fEv56wUKl5Y5cmu
JqiqlD866kz949WWmeBSIJEZqWO9Dzl7m+LBgGTa3hV75gcgpVfeikBkRZvX+Mdm
iCZOUcTSFjrPiREgfcRvmqTuexu0ZajFK4rWj6E/V2aMsALxe2kKPUbB3nbqnUIk
X/e7biw/B1NNKp/ETuWJPwRZUcg1LdFk1DEc9/IDR0CqM69MygUUODjKkoWvchDJ
jAkHEjfBaK6M6YfrxlexQof10UoKetP8bOfJuZg4Y/to4U2S9TyvN8dp6rvWb6Ye
wxbTxxa+c3mvIlWp/PCsuuHW8cP58BZevOmKCGTyqk9ml+ymR6mWwcYDVbalV1Ed
b9ih4JXJUUid5iokR4kOhQh5o0SbbPTHlsbp+dvC12+KwGal+ocqCPBjrmOIqoP5
/yztfWbudociFpl8trOgkDpwr1Xa9v9+/1HjXvGThkFoURmevvSySe1zpx9iUmvX
6UIU2kaQqs96v3ZsIUMgTxad6s+VdCMSVkFeGHKpWb4e+HSe4BJHHVUuIH7bE+Yp
alQUoPUGRYRfy6iK8UWX/5B0qzHi6xoyaZ64i0IVPNKDLVGt5NcEvbDL0/UDIGb2
vOb2lKItW5GYFZM4O8XCdkjMmqP6+liTRJj5Xtf+q0pTE6p0NoAcyzBJBkuVi0y5
bR4GbpNWsWin3o0EKVwa8wcIdexiSoy5v955DCRTFhLPHYIkQA9QoGzX7tAENoxH
ykjimF6T7W0jGnjuww05elzWs21psh3xcs/BfsLngw3zcUDTXStcim5A3Ayy64lI
nrEVQ0OiyydUEON4JldT2fsmcjWT96AuK8R71qP388CCD0OcqgKAUysG5sqP/PD9
b1dWzbV8GjeXmpZhLm8SHdFSYlQELemFKSe/1IdDQt6gjuCHzt7LwL5BAOisfs/U
nMRXKOpm6jKNYcP/dKFQaQ//ZYl3cCI8bzh5aHTuCnbMM8//PH3wvNtUx9aedJpL
X4XodOw0AMYBXlsfyjeDjJ3qIRwObaXv77Z2vgLebKWZYxJa5u15XpCvuvAfi3w6
Ab0d3Ty/EK+hY2GPt9GQIZOatuOaIeaTmSuTm7tNzrUWrP+9t3kzGaKpe0gXuVEQ
Ai/iIIAnZCe6m+J+XGKonk33IhD+uX3KmywYtl//Af0g61++s7uV+O7IJ8GWR6HS
ZKE99k9E7K1v51E9t4M2GrCzTufUuWR5ao3sZ6cQ1iVqSJOxL/j2frAiPOFs3esG
iVWxfan34k2GY5KxRQaA1OVstbIxqU4Q/vVocY/6oD4+rvsszH4hE0EF4Bwxa7m2
Ymups8XWoQqz8+lY/XN7hjg0CEDsHKWkzimDgYmpWFc8AKX/9hM7ZqSNXHJ9dhw0
LuBPGEoecLSi0xYrqyq97imRJ+wJk/ZooapwHq+hWZuEk32o7ZKILiOzIx4J6gS9
RaNPlh5Ow1Gaihpf1kW+im9bjAt8jFUAydENMnHnfpnmoCiykaBZp4KzHiwzHoE6
3CRCf+NkcqjRqNBoziOXvFg+kVfEN/Q5CM0KvjEmA3P0H5+GVXt4Y2ICIgeepdBq
7d22SFKB9eMgqZMnBYoknKqxt7uetKAUx/kfUBNYLvZyaGspfDUwapWRjzH6ZMT6
zKRZNP/cbQAZgTvLQZ/W8if1cn9OYJta4LzBJcvOQhpLu2mDZM3uApzrV6g98X+7
4hJ6iSq4tLjWZAeX1NIpa0zVM+zmfPHXdNhypxmUM73PH3jdBi3XCbofv8AnuFBy
6kBBgTdODgSCG17MAQoKyG1djf4SmVCuea2grOah2RcAOHzNlcLjdITVeXDaC6d9
6pxmFhVYsWCVPoJ/DvOLLQ7aTI8D4gIJP6dB+wKsnYrbG/qf962eJjzCHnVR4dFX
/qz0ycnOZQsPXPnHXFElMiuXpVUIm/ahKmgz4XqntJM7F38Fp3yLGo9Ddl8QG/pJ
Y9usQV+Dv92k74rY6gox02objrKCRZIYuWnE9fi1CcmWtMo0qBZ39pmiEnkuRQ8w
44WFB1zYHOA6smz6Ni7PIodG8QxZRqdBsraa8gz0dnptb1SZdgv93v4bPkkR70C2
C5CEt8oidLt9b/qpqZ6UdGhnK0DjcMJh6Y8jW25kdNGc8hWtLl/362iQIKfh6g0x
hvJjl38QMn4ivhzmLS79KLlon3v08W59tqcpcKqVrJwWo9/8Evh7G6IRcwKM8fnH
F2VjKOl9t4rusNs33be6Joc8CzhG5xs3FMTewDlwCGL1Ew6swoUQVirDRH9LkKGu
r+sDgdI94aconAAebDY80QrGNb2Tym6V2RRrSfVKayegs4m0NzvCjLD9kHnLWag3
ZRmMPo7FwCXrFd/7zKKe2LkOt4mU1dWlKa2R9wokNvs4PuR4QEdXTUx3bt9PAIOt
2uPXf0wtgQX66UMpf5Th1yDH07LeMR28ELtZ6+mFDN2knPfOQhDeOZUGylgSSjrs
mUEf4yYzDqU2nP1BCS2Ggh5P53EivWlFjUL1aaGaJ9Xox0XdFfjzcUoiG1v2qLrp
/W8LRKn0oUNOHeS8ZhmDBNjryXZwnBOM7XwwnyxEoACHPgid8OvAA9G0f0pV7gQA
MsIZiIagN+4LoZIYG3LtFCScUkiOihcSjiqkqC3H1Gp46n0pT7C7WeOQGvF0CUVv
T2zEj0wTXY0F5g+nFxKcmEqMU2SXNjeX51oXuA53ZwpwFgEvkMGNWYW5YzzsgZan
GlrDSohnlMgfftw/bvHOLvJtmRSXYOFr7aeTYM1BO4ILOAe5Jp/MYoEXSPAGoein
io0j2V1Y5Lu+4NqiOeaJFV0Q+Kv49D1nmIHCTt3njOs972hUOo1GSOL/HpsxLuPW
jGqbuXMJP9YkaP5TPBzgzarMD3nVDCnG2mX9F7nT98fk/qRLa/dxYk4AVLHzj+Ab
JLjK9eHYYl9ewgtN7Mxtxh3pAQ0tFt/JBLYPB/R6lH/x5KqbPEDRJolsHIuaYE21
oAi2E/2Zko6gBVl7dqIw1qMk6ZOZMsCjWsOfvlFiN9eoHf6ruSkG1kctJUZ3kpwW
aj3DBUH+23gi1MMupKNXy3rNG4ZyFxkTgT0M5Xqans29EoTlF3s1UIWp7u56cu92
eWCGn5044AEWXjHEp6qQ2k5XAtmIIopN/6OInnD9dJsh6MHFFkODGEGz7niBBHIW
JXD6q6NMkQgKi2S72BTqFy5fO0nEH6J/95jRxivBt5ZQO5OX2Wviaj1DqKGkCIsn
/RllJC5N/aeRmo338EikE83tcqAX5uuJkZVR+VgBg/IWJe7pvilI12TTe6r1wkoj
nxDjVdrMjS1NQ+OchzsbYXoNwG9wHp9GTgyq83BycwlSqEN/6id44/KjGmVgYGUN
i2rh2s+GJSqM8ikObDHVeuGUMLp44sQBdikM6pGHeSYJKSobPum9xSgJpJ/K5zQr
Pwu1XsBdirrbOydyPFpE4GtedTftQoqC5kvQqolu5m1xMKi3gUKfbrIAMc6HkGY+
/ceiECV0OaX320tGxiECsm2Q94hbdBHc1ja71G98ITaA5LnfDXUcyGAyxSZ9f0w9
AS0rvWl49ykxYTICtRbUt75kkmynxw+k4WrFtAhktR4wUWfH473JxeQcXNx1uEzK
rdbs0QxS1efk+kSxY7ROdFj8SudBoV8Xc3NSmKIuLRW80Xtk1imy0RJYHKXKn3lC
g0wOw32O2PVYyMcBLqXBxd1rogLZkSHdW+Qyfc9wscAPYH/lXgHIKiwEJ5humJPl
/JTd0zxClFS0alO1v2zUo2T8cnN2QpTraSQvjcR7pEZwaKHZ0vVxuUY+vYiE/mb6
WA5n6B2Yw4mHBrRLV6pFfYBvNqm4MKkcSuiX7CiIiUpci+IY93MX8pdmt5owYY1I
y0O2OjT56UjVxHcWqg7iTtZ93QjWjt7k6NY9xnjcfm7wOPpSwJvYkGcGgqCm9TGe
TUYTVCv9VDLxYjAz2g+72ZFg4yQgMxjpTtObrC5Tdh8hg3U061CMGEBRXmgEPe3i
VEQTsntSFqpQWXOrCrKeCb0tpgqQpv1kXvvX4i7SAUtywszOJSJr03tBP/GvFnPV
3D4dj+4+0C0FekWjYyxq+G9iVqTUvJMtCYklNKhJIgOdTum+6XcELzsGrJ6zbIyn
heij+P/OCecYJUlBRmj4WkPCPmX9VTJTNaxNOvUeuDAW5KQyQtpu6sCoW2bELRoj
drfUd3YqB/QloadhUNFmTy7tBHXp1UTax6SLa0DCR8rqzdKvAlvtXgpG9u4ii5UZ
sx3ZjUtyKo8TBgtX5qIF4Zdek9alvT8FW2hFEHONBNbfv5HfIYe4jxGO3oohN4Wz
a6n7DtQL9DmR084g7jMmH1OXp6lJmk37E/PFlL1H3onsm15rg4quSoZ6Zv4mLhZG
wUPY9pLsi9b2pMluUk3hZldZPHUeikhsfhl4fO4D7l+ym4PIPl2wPetGmZZJul0P
cNK/Z9WTMVdfJfFueblXuw0bQptGSyImDaVq5XQr52bFKHNXjemnxBevyQt/XiBP
rojUoVv+vbgtymCQ/zA2wPgap7bvoAQf90vJfXRhPNV/5TORP1NP9Z/R+t5u1mmV
/weMcgy7ct8GfkHLC2Zl2rU4fDr+8eWZ9PC8RrzcFnJQwhw9eytnA1WHscgaw11F
8N2En4kZKRXocpt7GVsiiHpqhrWcC+X2OrZYRtSDrEUNzAJ98DaBhRXySSpAtWna
KkhfN0GseAnNuuQk2o7c7xoeWSq4dG186V8gcv0Far7kL+M2eOAYJ2C/hOTOyYGu
kUudDRC+CRS0Omuo/ZOH7GFOg/UYbjTs0nDLo8GdCQ8YyXjexjYopGvW3TgCuBvn
aqHvy6sIyIKhYhw+nNyUdvAj5ZEXNkRAq9Tu0V1FxUOCDye3tyOjLartvsxVurLb
ENj/0RP6rQWWYqOtjfEsw2SGQQsZJng+GhDNIPvFMhxKxCwe0A8PiOA0ShtCuFhO
JzIU/QTscLL55yCGHwNOtIMDbL6Ad2PvaurEqHVssTaD2X7ziRGATfgL0CoNbcUc
gUKuoXz76V6qcUC5tEzWqTmkR0QHdekgjf5TWL8w5zk4Koyzt+vXY+s9c6/cFpLL
NiuCJK6IwxQiz+YK1gl+K5ey0set520HyZCcS6Ls/u47zsEkr8O0/p7N74cqPeIt
zILMgH9mLGz1XtnB+15NrNtvPc41XkMYGbbnguL8T5h3WEpCTKrwft3Q/HrqL/Rh
LKfWWUpfQFU9g29tcvHhxfLH76qdn/TbXygjR5CG7Bpb0whNLroiLzxvqoRbBRYN
tJxQ+N3C8IipAc0xqyHCZgz4BSES9i2WOsvubRVMPSdxKmefrwJpxm4kNvBNCTBt
6oMjnZbIyDk+ylp8oaQA966S2uWrYRAF7/G1MpfjCPOd6uXmRXu5w/Crhj4AxQLW
n22jgLIzyvinObTXC9wpQH+0ADn+ZZEmV+W257rVlS/dhNzFA8kUaOWprLbpewp7
ft3k6xn0BVFfNBdfNrTwPCgk6FlVKZYqF5ffGIimjTswWRKMfLIGnp1ebmAc0dVu
tchEJKpBLdc2FkcO6sMbQm7Kdm5nr46x9ln3uE/ayuEFoFd9ahvlGGJXbiCygA7R
yLuijVrcAtxmbUd9fPOw4pOeAGyU0O/ja4mcK4SY185j2iNKPB+uR4ArwWOzWw3A
L6rgfZM9Q+1Qc3vQXKFrCYbSDvcyqSfEnt+cZ2evisPL4ZawDs+yefxLT9fxyEmK
tdtNVi+Vjg1ylxD6trQf87oY8l2SwGk7/fnxnfsyVBjpDbMTQhbaGwM65ZPXH9UF
eNIuEr3fhP51PIfG6ddRMOJV5/o+u8hdxra7roPcrLQ/Lnidfd1QBaCYO5UD776C
wBOvlEPDQblLHm+sAuYOIUuEZ3LrgTgwLMOl4ZX+/o4E+VqWWoj1tOwA0Kg/9FBd
CMvjf+ImsnS8+y7e2+iVXMAQ4JdEBzUXv/unFIM4wy6mVHa34GmJliN900O2bFy0
XM03TYW/hOZQAHsY34BZrsREqGVKViEc4kPS6vHqFCPHT9tZ207BYTd83q4+Z/cf
K3aDBB5DrBkOqZRAlhL8/81KOfW50gw+kfSMxJMWPUZRPPGEJQ55tjuT+Ztwp0bO
FXCeYBNM7ZibA3DD0SVBtkMYUUS1JbyeLv1yi2yLHLcAP2fK/3+ZIcbLmtY3YAGS
5iNE2PsqvCkj6Qh9BzdGUyR/zcW1w3MglNRNwPv289Xoixl8uIHkGQceMpMO7C2C
Loxin5Y5Dj46CB8E2+GNFxbF+A3H4rpo/6HeZ4JAyqVxr8y/77yWrivO8mvGvo/C
XH0niUoyBfQ5Cn38ONDQZB4gJt/Ryf/e7Cgb02E8lTrP1VKQDiywSs7ONnvLv0Jn
34JwlyJS7va8rZPzU18ewRrwMDTj6dxaEc7S4lP65lYw1+S7lnTL/J187CJDwMja
4rCHN40VB5OwpJ05r+4PXP8oh+oca5P6aSonAzqJE0W1O/GBg3eak5Vg0gmjdn3K
FBRxrqWZl242OL/Co45vu2H7Em3U+vCG7vmjGYoaEAPKHowtTbfcxV4L0WwaviWz
0YIu9p4O+UfufQ5mtjvy88uhyjcFWnpx637vHLd8NdkdYYltGqw+LjhmibC3Z2Tz
szcgn3Cuje5npvFSJsVEgEXrU9PtaotbnOV4VCOSzHM8zsuBQ2dw5pyUgQx520Hc
pvq32UfC9WpKXpL9t+PV2EZDaKYwFkZjjpCd1bHp2m2JD8fN0//XOIJ++WaqHdEQ
illxBiJBarjyWZEu5tRvxZ6MiODzFo09NwLtft/12zKHDYqYKlL3yjfkEm2gxvwT
3/wCa7ZuGX+JIYNAFLRy2zY5hUxqwO/hI95qr3ocoZz1cqCZPWyDwNjTCiYAYrbY
cSd8s8wOnDdHoGEgrWkftkT/e1pmbwUgf25yn9Z1vLlHbf9lrn0CNAq2QBI8JUh4
5zE5zcredkk4pLVM/hiFSeASsS1bUW+/xwPF4YId13i3hD0y7OeI/kbPQyxceuwX
SEHHiqpI2iOqIj8G6vrJGxucxv1jA2G91VMxxEaM0BQcXAva0ItOJdbAadpBnER/
uvqr+mNi2UbIce6u0JVHxlYEtredtNSLc/LpFWD8DRqfaJ7nt18uqMSpi2JS/ASS
3zp9lNAlMvwkETPwdTnPIG6S68QJ9LkSyKqY/er1U6Y2YSnFdq5bspKcOD7AYbcV
iBmKcjcn9sybaQeCbuqaG0CG85/7jcL6Wb/TysliJDGB+sby0fHXlAt8L611Tpqo
a48GLTxZilnSDya5OEO9I1wEUK3Ns17CVBbpLVuY/BTrTx6fmyWNrZhZpSjK9Zqs
tz17b0AVPprdyj0RinTvcyPLlzQsKHzo5qnCGYDsZGxSTzW8TWyVUnPzPGdjLx+F
h2o0aIztcZGfXj7svccfhK1q9BLQkfZNDMzi6e0CKUEqBMdNtx8+rGKdllOQBRhf
pItv4Ur8l2UFSVdf8Ewmnu5ARGh5phNzDljUMeDqjgUEjcm28TJwn/eBmovsQQlB
9fcmBkTadcO0pqYPhjpGHku7tgifjyTaCLDG5ALhPHnihHd30aPfDGRC49pbhJEP
EiUdzWB9qMQKjx7WTx3/dhmL+uyJcxSUbIl5G21DAOQLT2fVLMx4CWuYY85h7t03
p9abAKjp5C44T8LJqo0gWZ+WTXDvtpvkpgCsghYghDpIP3XQblr/bPAEnsYKJSVa
hBQHp7X3L4cmPuMLwyBcdgTT8DOPKhl/TetRTwFuwyiRFPMJfBrSTISg15aekurt
O6xOB57XNAUJTWSmA+f5sanmGpqZScfnYE5o7XUZco38D2qZypEAAijodftYbyel
8mCDJKQOO2q5pyfSnFepeRMl8w2JbMCvr2J4n5Si1LwJQk6z7CtP8LcaXnC+qsP2
yScfmfr0Wk5oGT/vBDbyinKXeaO3ba/G+ubRX8yQmxdyMYRUhEVHl5+s1lHGgV8l
6sHNDGuOHYVFLMgJJxfwt27zH72PXITgo/zo4C3IOAkk1NRzSOmviZ7ib7AbaOw5
KRhXkPgyFwgRF+4LFYJdoMmr9rV5hWpt9HmuXNBuv86f6Y+rC69RDYsAGv7k7lTX
spLF6Ci7uj9rJEk+nfB+mM6NmkEw9XK2pdSqsMgh8YFuosWDllD1ov/o1PMa8CPS
gtZ8wQ6j7kcp/0N9ZRRBYJohMpZfsBksmwbgDBF/ssgzuhprRbHizOvK5kH2yfcg
OeRZ/H3IKYxAuLWOe12LWgQl4Cfp7+FDbWvtX1GhG+Fwh8K5U80IKSCiKxrNpDh9
AhXxIVMYuvHjP+HmFH9syX7maOPTi7Zi4nO+Jl4gMBDrdMQsyW7aEVp+F9cETLsZ
CMcU9XUyQqmapSMSGOkGdMH5XmjKFhzIxoMKEjARibCShokW41fSPUBHCSVX2HWU
fYbVt4dYHLmKQWwJ9xp+qJlO3ZHG1OSzdq6TTIvdIV1JS4fXKNJWgLBrXM+exbuU
2i4EONk/Ca6sUDIj29tK3lQ5VoKER/7VjzN3GC2fUwCAeH+b7GfMYsniABsoqc8o
1C3TqoLps1cf8OP1Xm8lSxt+vRIzea7GLBISWTn7S6EH79SPGWJHjnc2KsS1nqpS
zLyWSIOD9UuQFb3JgOooPNogMfvk+IIwYHmCk01ALpXhV+d2BD0whUphqdpxPBMQ
6kGyV5XQvTDxLa9kEttW3AnntLC5PI95qgK6tD+PaSLPb2XPtVVPK/dgGamlqptN
kvIiwD4fVPq7kv1FUzdfccAF6ttV+lUSx1ABv7aFn2p6CEg7CE1jbPBTl7ki7sPO
4Crp1JNFcjFyRWoon1HrBNeFz4gJemp5S3fUxaa8ADOEo+JrEA54ako5lsEVcY9g
ygAjVEdpe3vLYxlLtx8BjRflVRnFX3AMFW1ibUCs5OKEfklFjw0o2vIMndjTxXFd
LNavVX5m5pY3VZXB3lg3uCbyb8XbJQ1VBJWCZbdtYqCiftY4RuQt1BXm4Z+Hqcb+
/qKlMTsLLmaW7Y8kt/CMHKrdtH40/87kQ+/+CqONkQ3oharhxodhvqWA3szJ5XTm
JCxUf6RmFMzoEmmxG2ULoX/jnFieMF2Eh6pY0M9lhasBvQFPpmzr9Mep4lKmAv5x
cJzC7zHrrcJVc34GnQGkRTrR80Ia7NLcl2OvbuXRUTY9PQgu1q2kMbt4EyxALIrN
GUPf2fP52E88nT1V/JW5jMWQZicOLEEnXVwZ2+o8ZuoCEXo95l7ZigGKnaLfZYlc
v9UwhSnCWyuy/rUNmXI5ag3/WlO03ZvqHSGR0x7CFlduKWfHH4mUrVugsqbSA6UB
QRj6VWjBXj9NUXeCxSW62cGJroySrWAPj4eCBEILZ4EGqFKP400jL+blqCPMzdkW
MtVbeCKXstT7bLepcglJX+jJ3RZ6vIimES3eVTQYHf6rAbTCiD8ztIrdAMhaT7HP
41bd+QHrRTxxn8BfbZ2oqaql9Jn1XiOpVwZzWTY5B9g+3klFmSKBUFlMbhy8KI6J
V4Ks6NBTlLZC74ueO2yRXqciev/Gqe1E5mZ4WhaYN0eebG36KkRAO8TjdGAr5bpW
+UhA5+3St+qQw3FXM5zYXnV+a6HPc/MF1TM8iho+vfDIAhcMbiCFHpZnCN/y1wlP
7s8vl4dp4QPu+GUsyrhWYy7mBrgkFqTQgjWGLdvIpXtddKu3PpcmjC/0SmpBmA4U
HdoBfkOKCJieVfbjObzKg50Bp7UYU4YhaBlnb0OjwPvooXrZ1GPbbnpH3ixt3aA8
IMt2boEeQ9egWPBubmG1tpejG/u6yCf67EmpiG9BSo7XlVpoznDIPqb6m3NNEBKH
QGRI0SCzLvBlNPjqmj0vWh2G1rZaP20ujwiYdYanNsuX4J3qSc22C1aiebyOzASQ
O7a1MSoSXcDkYY1DdiR2OCsiCi4naPKV931hJdn7v8xr6sbJ/tD0FZTCZNf69j9b
9DwkldPce7kUTbi4myFMVCUmi6mMV4OU12Pxl3JzjpISvPiwqWreI32bnvrbp6bS
v2Uy63/QHqzssXdaTdyMCBJR89LyvX2wohJvfis+x2oNHhyV9RjBvmgkej/ZY/oo
74A08aAWJ7xjQ/lMpK9znfg7dNrdDinUu5EdiW7/tiLyKOFCH8MmNZyCRKMkMKJ1
qQsiy2bUXjJK01W/Dll5JIe6N8Of1daodOzONTnc58dAATcHR128gYUC3pfhFoez
F+/Ns8OuY2t2IGHJLcsPwVNRu/aa/7OdZeZPtaOvgKX1+WMN9r6usMeX400VZ5Nf
PoCKD8f+mXKF/T857hdpP7wK3gqBY0z0+z4ISq613T8Z6iYoZ5MsBTAtgL4Ath96
OElipe+tJ3F429yn2o+w1xBeWf5UXZM8i0gsC6Z27dUmBxq7u1PyDMo9QrdagACy
XUx40R5gnrFp54frQQcoW1JhsayFXahiiRtsUKV52rbQVVSLy29aG3c786W4bb4w
yEtZZTWjTuY7o8dSHJSrH3gipgLjwJBo+/xSYXLsFI5CiBUTryCNhQF3T61wxbOi
iCcdP6P0sII0nYqT7IxqiG8mtvN66Y5f07OrPALfTSC9BezyK6L3V5F520T54p3d
aC/goHFX/mcmx4dnwQsBDLsvHVynQ/ZCap20C28u34zL0/3eFCyQCxH9CqAvd7kJ
z5X2k2D4nIDv6sOiJ/dbA/m+Wrp1QLHL5QPk3vc205VsQFzahc59KzmAE4Ga8KY9
w+CX61XIm78HudAeTyGtX0aeL71/ZX7om/sF0/fGROMYT5F7BysiszlntHXe5LB6
EUy9fncwHDu2afeaGC52f5vwSQzgaGl6iycbH8rQZc/jFVCtGrIGMw38mf1v7Chf
FHD2m5HyNcBUw3YUsSo+L/+b3OxGmfgL4cHsFPGyvbxdZJbqLRhTZRY+kmAiyD62
Y/Cw7lwFQeygr8E0Mq+Nc/n0lGC4qaUErMqDslODWVbcM869rYauAivuYbyqCAbr
Imdk/FxSKzPZV48xp35vjLYUnGj7khlh/WhdzTUHNb6aBf5WJ7+Re5k76jrubeaF
l4ltmXPC8fbjHFCviEMpsk9TZ/5ivpGNTz7aQ9x2/wbfO/xcEfP5eiaYwuLz38y+
bff/kWCmAKDB4Pew9yvU7h21a2vuG+0xIADPhEh30v9tEB/xi/HDW9SfOD+OHqHl
U02fZaivizfsc88SOUKuST/wpw3TqYiG7kh/0/9nd5BfN82yzPKylogmmDyLMKUu
22vo622uJtw+n0eQ1wLtGyO3KJOxomGMn3zxCQ3noNz9uUUcxnRwpoqe7rhOOaze
gageHfs0dSAxh1UlhUVnd8EPeRaiSsD2RjKPW7PUBIVoyRtCb0K7q+G0pa+LwEVb
x2+mEo2IldfF+CEmbPaF8EaM3pvtvlTDkXzgGCiPFeeft3lfJl00bmnPzIDWAJns
VHlnqQ5bUG9jfNwMSrVIIIAxLETOpQWzZra/TzEmVo++ocrq3gydgEStfY2SIle9
9MpVEVW1j7JPGnA6UrQuwgRyeYSl/S8OvqXK57QpgAwp8q8lHIshslUKksBEFHk2
iJQ+QYE52qKq7RFqlqN9Z4GHje/CRfw2NXF/Q6iYvDpbJPsH7JSEy7U/Fj4e0AZV
OLWMSMyhfyAZuLFLMqHxBPn4dXrexp2xF4FekK7ShCUq++kmDxpje691VsPeJu0F
tkXbXOrqhSFuNmdmJ5Ewzg3GFm4esYfsnEwgrWw2WGnk5GmmIobz6B63RnE/xx44
WAFbwwpGH4d7cMTMtfvSQVBunCLG2jbfNzciUN9Kbac+AjdKvdnRPDyqB6dlCXA8
twBALuUeIALw0cESCnO/2YGqB9mzenN4Ys4Q2oLbaBZoQH05+s/SSLMIeMQeWRI8
uC6UWYo8I8JQIyXQEF71IlSshIEU1yyr2rUxdOj/u+vtK3x1MwdSFwp6eJxrYS9X
oWJRcC/ONiR8kq6QXOr+WPtSOofA1XDp43+v9rt5Ghrzqf4BJd/YleLPxmcMOkdS
M5jk6LW44AVKSsgwGBsNc37C4MVbMDDazQr20P0PNhojnrx8dFRccNY1hZhdz4b+
dx42vhwWWwZh855cYjqR7DoGMQ3znVH7TciFVPVlgQJ92KPc4sfts3iDRy2cy6vr
6eXoCx5CgjFOa/9D4kALpNsdshro9MM2x91PSvKlh294PbGexIg9DZBrei2lneYu
Z56zYmmuUULgt+f2Vw/IojQQIihdb+yI7HWED7Qcuy6ZQmJE82UeGHEzybtXNuNG
sfIIGeJ13rqXzTjLFovtHD+zGvM40M5zJnhLE9zQiazz2W88efdGLmtJXQ3AXG37
LvQkcwRfvjZppu+9DGIrIB9A+rI2PbturByfETn27Wdkgw+GoL0R9cPs3h5IQQj3
DtvFKWmNXzuK2Q1VxCeYKFXSYqIZwrBIXZO6S1/XAkCU2Wm2EIZ68s1Yj1FNPGBV
Nwl/+26C61GBXDUkEqIw4A09+81j2Y7U0PIT16XDSePuzs2vswxxOnEz16tgDGRs
gseyL2ao/868+i7OGm/Lb3NBLTu2J6R8M6rlBNOGCE9GPUan8u5WnUI+BZRod5PQ
BUxlX0nkPFiZuhb2LTL9JkyL5uxevAes7GogPoYBl1CC/grKh0z6nCN/dquC6e13
487y5wzz1KDCw+/mdntT3VEUgDFLjj2dfv6MTEL1LZkx5saFnywCvQYU7kDnmtOQ
Eu8ogQoBvUL0mUxwC5u/hkzOZKvN2oBXE1qMBwhopVqJsYrSUbM8D0RxptupEPul
WxPgMJEl+8v7Dwy+BzSO2yOmriVIpRv5EhpPB+v4dRnxgYXsZg/wZauMI4N9z64w
BkgG+hBhDruaZu8gPvYTL7uxBN0J6RLP0u7YNVsypScOkJ8euc5uZ7X/SPgNAU47
IzH1jZmeyHHc0x+6S2xkHFRPTu00rkkXRxLFgzJkd7H28KGMmxu0gdgH6frHmk4r
XXT2s775qGPAbPYP6v6fC2pRJYlhpTHdPrnc41SKbbN9vVHdbCu1T5iWjeLFwTY/
eQozyKq/2OQXsxYA3R0tdG72Lc6MUBJdRH17TqqJVywjtrdMMK8Z6XIdn+YPc0OY
WHZqvnBIV6+g/x44aGH3Qmu06cbMKyA6mD5roqoyzPXVVY72KUATt7IXOfiVoZbC
uHSAfEW4Pblhqtg03CDRjLkt6ZGHsvXJLXGt8X9OK7bbTE1TG2BuGdQcCynE0yQY
IsFYsWgY5ly2ZjmALY1v5991HNHx/SbL6NAWX1xUFFr/jYHsk7bnIcAxDesMzpTT
I20X6PtufxNc055GuwMayvICon3WDHwT65upfzdJlJGN82FkhvYffJiP74orYZ88
/b0OLkiIkRp0TjtFuX9kMRT842i3hOkgjrPYCVbG63TgXuqKMa6WYkqMbvl62+ij
AiWArRUg8M4JJXrbMDsJYpYr3vxYmiELP1y7J8RQK/4Y489+IdQjHNhumrIc7gA5
BOJnCEX5H3pHeyBqqwhcrveCLci1ZqN15u0S5aK3kpi1WX4rxoL9EnUvfb6Dj32T
Tbso/Vg1u7ICCfam78zzfiSvt7HgRH2KeGoBLVRO346x7ya6BHkHzZQ5hL/mLHoT
bTcvrF5huxk0VGBKWV5ZCBCF3Wg1zSfNQiH3mnjjv6BsnDh3UWqgSFORRTmzdGWO
xBriQxo4qXz9lFef+lPTfVhoDcNkNvI9aQUG65Vn33+lz/oUDHzZ3l8OjgiQMFci
X0LCZwOjbgfaA1FW6QXirAzzd7YLeTYy+lZIRs2EYJxIvFk8lLUlxBvPdtnrkMlo
XDJ181nhwUYbVu3cLumijH98jxRS4tCWaHrlItLRO5oczc/Dtqf45uPlMZ41jmdQ
iwijKbF5h+jNAuGbR6HGCjHkB3pwkCHdKQNE0MiVqINdwY1Pg2af+5MNmWjUyUpY
oQ6d9oEPqI4iGqZruonoFdggdiYlkVYi5o2uFgG0JqSS3qbZ+Z3KhXX9IBDTJ7bM
hPX3kqSAO5XbMKjJOtMtCiq6U3TlqruwHb/1UPenWNh56+qN+YDCR63NPQwFZyjv
0etQzHubp4zEync5sJCzG8PIldu4UJK2J2y/RJ6xDYcb7O6oKpnx3ZIxvl/acbkM
eM6HTMnzuQvHnwlAyQyHJnDx4OXYQYMJaZY6tj+gpTMLkZMwTZXsv73y3GUlHjlZ
skbQoAX0fDLaH7GPlKxD9YPUqDObnfSPSo1UqpNcEXDBrcPVK9T9Vf/bmFTAMqBS
2br1vmfHZ5exoaJJgMHolldRK0+QNN+8+Ixp5ypZMxyHSUxTU/cvp+inJvXcEOu2
Yxmw7KsiB4FZRiB5BwwFtzeucGdHVM0EF/kyPkbvbyiM+T8OoOS0oDK3n6uSvEMB
Nho3zDp4JPaVuJhZht3YSBsKncPNVyie0IQ79hvr3wSbvllLfEFw+KCrVfE9+Qih
AyrvMnJIDqGOBn01CFkKSejGmSG94menEVZ6G+RHGEikCfMU0kUsdi4k60IysbbF
Beh4rNLAugbqAGRvQ/cL+qv8kgWfeheTeyrFVI1Sz2EaohuhkO2R0a5hCcOfUZZk
C4Lrwvo4yTyZd0zklAg1f+Y9617n0RgDkFtsGbK/4zbfoXjgGLIh8mawyMMtHBdN
rHZwdYILzoMF49Zj/X45ZXVvRZm87zvTVtIFQ2R8m1rNSz6c/qLbrnW1qZH2axYu
6YMX8W5U8iDmTOZaO33wgYBPuyCgonW3v/5dMxe/+4Fthw9h/CX95hHprHoACPfI
dYjEJuAICyzql7bSMNbZCXWJICRKIC61lMp0BDSu3TN5bV+6hcqGV6p7upxWOQHQ
Nm3uj8r/O7L2YZnGG6Z+mBPZ+TiFp/CiMVnp2awR2Xkn1jiqNiAvXcDtu7wDoSB+
OmRONoQIlCvkrFbRX0rBbHOqXhXkTehgG2xw7UpZEyXvUY7jsZhL1LM2m64zAJoh
zm1tAAMpWoKChDXC5O5gNxgbEcgVJfodYFuvnccLdawqzEHlzety+Rw2IL6MN/gW
XwkTpWHGdtVKWtxyk+q6OilhKFaqgWwB97DIv7YSVW7udFhv/XWXnC3Z4poKIqmh
cmSgklAfMGyVZHVMMK2xjHh62v0g/rkTGbHj0fzGyXO0Yfkn/wDn79EVLlh/IySJ
xCHCtLQ3lPxjyidqxovRNlWz/WyBHWhQb+GkS2NzGdr5j+G/gy89Ve3RI8ORgnrW
FvyE4VsQfhoA7X3nFEOVtHQ2eksofYySqC78sB/9bh6shJ1zjsgdizf6pwr2FnuF
uPpk37X83vGMd7azyGobyLLmDnR9iLMxAorHfv1188wgWS2R5tKz/comHObQaru4
iN4TcKc2ZgY9Ir+t+bbA0uiANBLy6murkiFQHqip0L2jA2hAzVrD1Vgd824ohitn
cLTQlONHVofyDx/qABX3x5kr1p6R0vR0x1lQq7DBx6qPZQtDU1/05+zsqrQmhddn
EhlSiGJ3qKep9YIQcEWYzLq1iajCNHoOtgKQ2CGZEAnMW4N/rwZ9msx/8Sw7RUbn
ySAk6s8Fpx0pevt3178p08Hx28jWx7GC2uoOTS7f/R8kdkbzeziAt20mm4g7dNnW
qm/+5hEhe7BtU5queJki/hL8ISpb2MnJkcWV4r5J/aV+2z7MprmsgOxLFfz+N4mU
6W6oqO7aUYWF2NCgdHe0Pwsga8LVEADbCHTVXBu7jMrSnu86sPUM+LXuvHOY+jgi
OlY7bSg2N/lqgT0wVT8jmX1Se65PlRP0DKgemrk7F1FzhzSXzitx6xuscE1ub8aX
tFusL36F8OBrezIGixAr/PiZZPGgGAec2JXIrX1Cm6d1MvCZZ1wfvTZh6nX1qHOr
S4027DCNlhJtJU5YNo9dEJdbaBw+ScUM0ugwKSCGnKRBh2gAm6mf3OkClh1Vqllw
27cdoMbOIFnfJ1fyuqFXyLp+exDodOi7jMXTGLlJ3LhKXxVkIBigAHUzHXrVFxPi
Uwu1XdtpVb2rMUUpcsAXhPK80j//GOLlzB32UcCgqYWnumjYnRbX4s6nyoYl1+F3
+5wvhD1Zfl+C4P70SASEciin+ihUbHE9u2GekNqxAG6lKKbgP5mOGmXcf5HKO1Sf
VDsSPqKFBpEx9GRIG0W3wmI7AJL8W+UQ7R5eV3uskfyB5fQPDAL2QAWtw19Grc9B
mVVyuK2535gQursPk7e1D+BHXPQ4sAXX1q82ew7aRwKUBtvCpPVjMxx5DQJD81dw
Dhvrw6fTxlaWBxspJzIPoRmcivtdKdT7alYhAUgih7QA7LLfHJ+tcgO/hu5yh8H9
tE8Yrp9ugiJVj4sPe3jEB06DrT3RgGDBL8cS7FJImqOkOEIQ46hz34k/1XEHlC4K
viHrANt3TMs+JUOLalprhsPmCdVPpLZfW7Hmwm+NFVdpbZXhBZa8/nHFtAE7BD7G
UNjFz3UdRX1uugZhQtryICvxZZK7IeBKKEWFMC0wqJi/dZlUZLXf8sIDUiGNnTlo
u7OfRKz3nlTkVM120gNVkInwrDx83U6VjEyN0Cj15kOWkIe0wv7nruyz5Z7E4vag
90wimxe5V/9RJ0uR19lkvEKwDHASp+XHVWZF93N0X2SMSpg3hwVihVeqO/AKGn+4
PZd2FXfIO0/ALHrxVX1lETkkBpQK/ilfT88iZzgMf4q5g2riYoAZDGUf/BNSCKHl
EM/lZKPlkQjEqBI9z0ShK1IRPV/9bKKTcMfblTfbfPIg/ZVdND9cuNCkIYOuJaef
WGBU/SUAhuRnOa8V1QlcF9IFdNQbovoUiFa8TRgVLF3BU/fowLxB8uauQ/uZsaMc
6VM4D7oWUoV4VHMSzi+4YcJzwUSRMgcMj50QxYJdy6BtB5uERN1XuYyKwydqbF7T
6qMdO2YW1dYCnR8Hl0LhB/Lye+UcFWmZBWOrLLOB1CWhEQjgQo+9/5jdAhT0mPaJ
ckM3RGIrI+5f/SqLxO45KXhAtW540f/mtj2IhplyzUciwntEO4RvsJvIUyslJGU9
pIyfQSHHlisB1vDkHCzB4AvLRV/tm0Rzmpzkx8byiZWJU41rGvY2jnT4TSwvUqVp
8bGWvcGXl5KUQKoQZVvuPsKN8j1hTAvAe97MoTEY5mFOmKiZ75eGtw0YoAMabopS
WJPqrjrtTSz/8S6yfbliJTK2NyvZu1UOAvKrnY3A7rZPiwoGQwy/BssC7Im9w//E
8cXvND/H1HK5V+cSP0jgl7PJ8Rgo/lG/sln4TFM5FEhcShmGAgixE5mbAL/2+kcv
f8caQnGJm+y0C0VNtA1L8hKaNdFhUW/1hJ+qBpZoTxFpBcBWE8YHewdEKu71WLuy
4UNyPhucerSlDAVMO7pVWb4t2NQg4QolTtj7sHETlW3iSstg48bxuiEI+nK69L/3
KeJ7zDmmaUIczxVTR7094AURRyMp54APa+HYV5K0XJ35MYYfrXPfFNH9LYjmaMpL
kHe1QuvZmy0a7RGFSho+Gv71z9A6ML808IRX7NXFqPuTEmdNVmHpp0JKvBGSbXvt
RGGOnAWrpusX20wsyqJO+lnyvyiUiBu023EZ2NRrXU6WN2gtWWXYpJklIEXFtfDF
RfpMKGedgjuqyiftPnOPUZYPR7PIKQ/QxAIxdua1FiWYKQlKeGaSw4iq9Wd/zHnJ
JMZGMFHSxI/EBsJqoxn5gMlt71d6Y8yJq4LVtJntVPoTSrjdlpXCwGwNwZZ6ZzAd
UJNYyFJOMZP52ecfCTCXoWSZwkPB+gUJqlDN4n1+ovGbPd256DT5nHxLKvX9BuIT
S8Bh29dnYn4C4kGauS34pzjWIqF+jT7PdNhWCtOTsWn2uvXQ3/dMgX0JZPUiyzF1
e1voC8slKaOs4R+HZeN9FwSGqIxy18cftjT0kYK2p0LwUAlTEpuA6G25Yq1JMXFy
DxtaaqlQ46+o0z8JeURU7bp1NHFoKsnUX1f6QZlbMsQABjmrf7wkH+d2AMbVgJc9
m7/oyM17MqQg4F6jmYg7cZ4dw09/d0Jqgumty0FM1/lSAKtPD0/g41T3tLCkQ7No
zUqMwd29tJNTUkj2h1QbDHcQfZgAZZOzSfBsEB5+uVkduNea/2gApmSkwtdQFRXU
8xzID4Sm0t5jMbVxY8tebRmCjI/9PwxIgLpinr8nYic5h5jLLycqLf0SVEadafZl
LdrqpQjRzifYaY1P83uu3bf+i+QTRXCo/TAOveKbGPnY6yaAB2Gchy/ouVFOUq0C
akwr4UQvyqqrnJ3ZphTFYzf5rr+dyiF6WH58Sz3is6AZeSQea+r/WWtmwHS3bb50
ED4X9UG3lG+3DqqVvh+qGtqyH223LLgibXZ7V+EPbGsW39Ham2FKFjl1EKEKkyJE
PuhwOpB4lVguNH9AqjQ3xuCxaV/VUmFi/SY/RDyN+CWPllNI4vlFTwbXdJ/+3au+
iA0vZP/RqI0JcUgnSaEnjykuPM5vpgzV6bZ3+xm6t4lxgJGPd4+lNaSkpWqXu8op
C8i/rnd++eVTPpz8DgCxcttsH6RvR43wIF7EYBq+DfD+gPArk4EZegODVI4xUksB
LBDeeOYtGyUZSXosHeL5L/gQ4TCBjN1eF1Oz2b0AGdD6GwatJVljJt8/6I6txEtw
OkfXZNTsvhR52vOawSKeFImscA/02fpyz7i7p0k4W/82HzSvTvPxKzBu8urnXJ0L
WLM1vmGiiG0+1AC+e7UvucB1XMknvvUrrqAm+uMTizFn4Le/1IbKwolHgI7+NHV3
g0MRLWgUziJVJA6KI4wmvTJaMScsz1B0U9mlyzp/kAmr9vzau5rP5aooxJZvXS6E
QijOqGY5O8NH2fs2d7TIHLB8vI4ItQo3pDEPNkUGMULJAACE10pJYmicHKcqsw+z
XOis6kZq+CfJdBF58huI4Fc5cjxbDX45eTPYvp+SHPX8VMDlHxEegYibTzyaI8ve
mBWp5xbb6mvjvmKDwGyFrbEjs/o20t3sy6Ii57tHyxo5FqmrxF1OhT4nraQX9P7/
QngyGtUjxnQC6xzN3nSaw7MDq8XUqexoyEGLQwdClK3EZEkJqZ68oLij5gN/JJbm
YaNTfvbBwe7HQLEuQV+jjarLM8UCMNULeocFtsHIncNNgvSyBvSkr5LNrQP737PF
GexZMHn2QKKM0Rx2oM3SuzcejUfYglTNrYZ8mDI8HV2bdoE2pSvcum5lGPw50y+2
0LHvDjsLOLDpuib9wx69sN14sz5leB9ZWOvOcvVsIgaupw5aEYtM4vxb2M6Kr71H
MagMka3yGCzosTwL0dykO5gN8RdkLOZ8HQ0PxIt8imzaUAHQ4milV88WRMkg2Igq
nc7vKmaxPQcZ8aOJ/jzYhByK98y0X7I8ridTC8eeTg0YtSBxw0qQ1uGrzPg4+7G4
ZS2LG/EqK81/a0d/wVTVF9vPz1UBYMSX/NOQILZ/nkU/otsL1xGg02wBOVr0U7z0
pxHp7D0g5eCTgrXLnCDFHjgAcqngTfqYgBOySDioOh6vLctmgWEZ5zs2oMqzAvmH
xXIlN8r52xtODHWPKf/sPXJuuJyjYEX1GjlDdeU1d/Z1xpZmEk9IGl3UORD5ia48
yI7sSuh6bk9/QqBAwTUZK/pFVeuCDj++91HfxBtQlyvReWZtWacUeyhp4xKzCpv0
TBGdRHvO8RbXRFrCeAYTsDeG7Aed+sJ9FKO686QAcFN2p6toHnbmlZWATo9FiJOh
U9FuLEz+psQ4JLKXrt4/78qFr7drRuQYVAexAPaQ1f3c+y0CGzsxe8jMjV2Z4QIm
YMRokvAeeaIxKkpdqDNHjSouem5zfs9dijwMxq1/P99BKAvmhBaFXwc4PRzMe61l
rukhK11HK6ekySsJEcPsDBBrSZ6101dTYXm3wiThpY4jbq58bdbaJH/5Yq7K5gku
PtqzPlPk2mXvpL6Ojeuhu/ZV1On3cGtp51WnZO5vk8ea5nUbhLfuVlW5AcGkXupS
0TTBtY7XipSQ3ReaKM2B+Tsm4df7Q3bsa8qsd/CcPp6zD+I8g4AZ2lU3PNqU6omO
CQlgaKGDcNDGHA1fEAFsZuiJdLn7DSArir8aBJV7LmuXLngQvLR/VrgY7fJLXts9
jFnsHPwawYr47qoP/n8ks24Ap4rldVZNl2KB8xt/i8IL6wW8vRCl3cRFdKQ8BAIp
AQ9jOw73jDxqT/KqoirzpO+1uUKCC05iADeZVmM8zF48/cD66fFMXu2r7iQiBDPm
x3dQp5bekjgzqxsH/BMYmRiUMSA2q4vaSQWFwOs5zz/A9HQcpnijRSSj+CC2yyc/
JMH1d5spguSHUGNwCKQsY68amx9k4paUq3S3BZhRsj0a8lWuFv7697jFHSlodDfc
ftJEZ1kabHAqZchKrfE+OIb+pThosrksboxORbT6vDLkQu+tfvLx0Xufm7c/MPW1
ffr3cXtcG7Xmi1knasPrXUdKheWCyMf8RA9BRC8a5PWky9Lc/14TgVOxV6NmEtN4
cKN0y+Gdll0Fh4VZ1CifneCR+NM5kZ2qEPPy6kVME+yrXuRCyXDPqhbFev9NEKVD
9h/uBA+Y4JacLsLG4IyO6AJI8GVynJtMiFLQs9GjnGiRS1Uj0shoDQawkVkIgLDm
qQXTBQbx7UqLd3+bKjyqfdajTy3cQHwmh1gzZkQgqR9sKuCvbPtBQrTSf2AtWFvj
J83CEDJzBd4HiEJc3URR9xwkE4MFd6ZlaCGnp73LKFfYUz0RpzOOIC7ggiDKxAb7
r91ykih4a9cHXV0AcRuq60x6OAfqaiQMDNK81z5XxxSUUog4Mlix1CbnxEkB9ug6
SZMpPzxvHhKl7odYbI8dDw/B/Rg4lnry83ezGQeEAmytffSXqw/YKqYoZC6fBRs7
0sW7Q3maf0tEMfAdKPCN94ikOXAWqB1JidqQLtNgIr+6n8h7fhlsw1mJ2Aty6TVF
MMRilPWOE8Y36cUCR2UEBLwlOO95f+lLXKHrloxfI46C7b3++qan7CSmhXIMWGok
UlRzO/ZuPFIWV4FpANQxIOPgAXqVvqT2bLQKN9cBo418mHnoblOehzSCvOlJZAEo
As/ojGCYONw/zFTp41dR8ia6o1pSwSCIar/cbTZAJ/iy2NVAlPUBqKa1sl7T9FAP
2Ak5cjyVuu0LBY75uhvt+Fdbf80wRUCSpJ6LOQkUoah5wY/1aik1im0eMBsbmqqn
XBjBpB1fJSi7rOiSf8O7ZJNAOUx+xJ3c+XDfd2XECKXBVDtVFIzvxHVguBcFhbeQ
djuX6XbqztZLjFuDIKLDZkTntj8atxhglZsUVwdbhNI2qhvSwUjy3ZWA22nGk9o1
n9/0+UJIF7Tur5I3LDMPTv4OZ848Q9aNI7u++P0G9FN5F7p0UN6SHlWyt4dA+yF4
2SGM4A2b349koEsEkHqGrfjUm/woISxVrEGoRCDizWplwd9y43JsnWCblosGESct
o/m0HFUalVNU1FpMV1XIapqz+8LRNxTiHkeOr45fj+PFNbtDv5bw3SU+rVXwdFk+
qJa2ykhoBFPGWcGiQ0nt4ilohBidlyrndU+ILGi6VmFzxcGx5TL2wWhhn2oN2Ktd
yh9rIE6hY5kHRndIZvi73zwNimnJOfmsujJvHX5a7ofjq4AYLx5jv22vEKrwUhqu
gJEQ84+U2THugS3Q6dtbfds2R+1ZG22I10mXXkhaltIUz7rvn4xrytRfOfnEErSE
xPA8zN6H7owyqkEuAmtND+ksUiTR5DDrRDNldBjNtDnVZ4JshGzCRkLW8rE8fVRt
YhptT0JfCLDo81Eqh3D0CGWbWc/G+bjYiLX5/EDA7UTXlxBvn5+dPpoydPMCVkWs
1nXQKERT/R2mVyv9swRZkoPLPD6Jr8Zh0BKvLrolYt0gdRWvy5VmArAd9ktL9plK
BYmSpi+8d/BlqhaWd1lkdHROKRRamWhw1VyNand8pTsoihjeuT6vMuEEhOCKfkEO
WH5+uVgi5EDqHpzwOhjV6x4y/G5sG0RWNuSzj28tqqGY0TGX+djx0LJchb8u4LjT
LycwViZKo6OtMcttdhhd836bt4YSOA6RRrx9U54z8Xzz7HW5VY0CwP+ygCWvHcNn
4oEMvWN0qn2UfRlT14O0mkr1sOgUpLhx8YQvpgtj2vKE/gVIxS+DEcXcxLS1NDNH
q0I1HEcccUfP0rhsptMNQX4De6dBgOrCtAS/BIsvbrsPbptKInc0n9RBx6Cz0ay9
4S5nCPwdrbVvEMd1xDBcaC74Br/eUgVFQ7ADqezGbeB4Jo4XMwDVhmQ5pUolNdeo
LreXkwfDJn9YkPtyrNHV4/B46cp1ybjD9SXS7JCOTKzkbysGMPjisr3EmTARHmtq
geA6oNykoQUJcwhk+Y5X8ARB1H2QF0HrYHM96a6CfBafvta7VkdRIBhOfTAhuHWV
mm9VJ+/PWX524SrxRV05aPRBzvQReyboNHRjsJ9tNUcWfT7pHNaG/P2cMLooBkaD
YvRjdIEc0B+/WFr4WgfIh48c2PiNB1L42O3RbIq1YrzAIQBuCFoa3QP8c2HDQRbo
4PqS+nBr5BM0DSTeJfFidRy7TeLFSAF9dIq+LYoIbLV6LTiqPq2iwcxgVVGKqEnP
0pPe8GpIVSHkuqAlv+ZvdRmSWrXOvhlodxq4grx7Ur392TX/TDvW6ZavrtWTFpSO
DFw9CpXFkpS0A0lziDKafyY/cRVHQB/ykX/qjjDADvTxZfR03QETXMu9KJiPWk5B
Nb2vkylUsn1STSPHjrhEpbHeRDsq4RpsBYTT9p7Wy3cLtd5v7YXafBynyn+Tso2J
v7iQZbT/1QfbKZUdjuyNekUzRiqyNxccc3KBDOczqEPZmRWWIZETqYF77ENcoHjb
T2SAqTsiRf5Y4e8jg+GmeancDN773hPSVvQnZlF2j03PR+vImKVqyLTaMkGFUQiW
GVE7OCszc7m0PlxLjP0bQM76y2EVHoJenbgsDlvs7I816GDIdwA/tZRkJylVXxUT
tLbkrlzQBeVGXgm8olzkiz1ZSERFnG4bcAwndkLLJ9SBbcNBT2Tum6TLNppYWuDF
q2lav/Wpr9OcGnmb3a7EdOEXRC8utflDHTzE6Ic/QV2h+QVoDcOOs81RqK+KEHy5
BW3qlmpztk+M7XUoBBH3ewcwqOPPL710kvgZw97snYsROt9bgFmrgAwmuiS1HbVv
CQ7LvZF/6U3cwTn/P5ydsAyTKB8jJtEkB1E+6zt7dfAK/2Umj83mVNTQ56rTOi5j
TutLoemJvpL3G51/BHNMkt0l7ZiVQzyoRYiW01rRWegL1Excn5oqL5w5z72+UxRa
yWm5x2lSAWqWh5rRX/j7GTU7UhWzVbksiDw4IKFwHmpUcYp53wCdg0nTFcszeKD/
KPQT7hxN/D36KDaUnhVn+vzyT8BlfaHE0ttCdmveBx2dD4Bp1satE2YC1U81MfHn
TE+kMK48X9RFM7UG9cPfqXGdhwD+rPHkaLbIsdU9f0T1jZiOswTWYJ2YevuMRy6G
7qy/Jge3ufPGoQ8nNeYbap3FYSRnGxvKROvWt9oirq21ZvBCb2plNwAixMEXgjex
+KzOpS84MrnoYYlYL+C/0l/26chSBpBMdTSfrr02CK1GzKWpKQMNXALOdo8BXTRq
BlXwkDvKCafxBaPzBest2KXXDkLWNnFSLvqpgCb7N/SGUGV+NrOLvxKFrW1nutab
n8LcETByWynF77M+6CBs6rTT1hWIv4bxJoR0ZVkTx6CVoDz+3Nwjz7sXypb18fAf
19XDjwTykdgPGuUxH5jrVmyH2pBmO5kOyZnWvYNulCCImmdzNjWgT25q6fy8iTxv
TtadG9AmlRJUBKlhYTRwO28QIz/6mrpUUSSMK1aD4RqzT6m1It4X4mcrKhvfX6wr
WA2YFiNmcvZApDDDsFpgwGAUcY27DCKYZO7XfNr+8eRbLVBCEVfZM3XRyE6a5xE4
EeGZ7x2T+1kYjQ5boejXG/OoM/M43LklvMJ9ZDn7yqfXqFItCJd0GBVyl+DqA5Fu
tRXWTs6frh0go2dGHUEEIpS9cJL+d9ThdhYjKE+YNMjsOoIdPH2tl3ZL1wCCP+AU
AcXNu0E6M3RdlgUdOhN1l0XA9hKxYIfgxWfnz4i3XZI0XMc8airiLbV6zMnHAltM
QLexwWly712Pf8JUG//GkD0wvU0VkzPkbmy/rxsXvCPTSU0OEyDhUEG/OnBo7QM8
DZ1R1b8M6cjc0IAbdUGSZuZTm33gvPNnbAGhULiGMgl+jjAe+3xe7gL0m0mGVlr6
NhRemmZwt+Qab2Z5C0qPPDKPCkYfU0tIpnuTRHTuYe5OipnqW/ukZsg0KhjARKox
E18qDmC1I5e34sEK6GeCEqi81xnS26sVJ/NZ+BoK60BAm5xsnaYKz0z6EQfOcfab
aTED3g3RItJ/KaLGYaX+FKdafWldsxsLUKdpL+/Dt8xDiKw1pGS+mYO9fWPXpbmC
8GQwjp/fd+5fEiwtos7I3AXDLOWRLYBxagY8xVLxyv3MX0E/Yr8t+pUeV7mPNH6Y
hfQwjFwwnLNoOtRsxfgdDEcVJfiy646CwqqTSG5bivyspcw/YGa2txUgpNt1AKqG
nM9mWvgooG/RkxxtJ9ZbqnKw/t+IOoctlRsSFtscu2vbHr0rUaVkaDRk4pso7v4V
WxGWyK4a1yclpS7yyl7HZpEC0tDHYOOVvTBWENILs4jYNwy+GjBkcblAeRw4C26x
J23aPj3ErNqlh5dmq1uAe8w4wl3OYlAZrEbN2yr0VVy2SwWo20PcytyLuMwWiuRZ
+C3BKG2rqwnc2Qdzkbejyr/w+jHoTEYf9RXVXYBq9bTy0FQN7eHyE8KJ6zeDhIKz
3nkTaBZo4YU53R8YDNtKE15AOWrxQv4BvWiBvrD3c9DVoiwOLOsDCeUXD4PMtDoe
Fz7NVwtRLProcPJMC+gevCM3IBNtolhEG4SyrgH/5yox2ULe9Q0v+FnX/msud7xi
XX0OUoap2Qyix7GBDyX9dcpUmmEk4qBVk6Nw0TAaCPYYjz7WHD0UIUucs0n0mxiC
rep/owsNE96Mp+VVEfBQPI5AdVn9QGiH9pDg+yqry8WyUuYwvTI6pwTKhoN388qc
IJbplisJULIG8iR7sZayXHLdkckPzmGYKdUfTCOLhHDmUX8IOyUnsxpSUkV+9pOA
nwIuiT4PRYQqFIxhadx3W1R+TlttkEY59VLhguAoMTfc7kD1PkNWGDGabo2zhMIA
MJC4XJh/6YiwEh6yVKuDsOcP2n1bU0SPrWPku8gCF3pmDz8xZjZSu2zwewjs2/xV
ehDfvN/1pkL13mCIkC8FljyTMQg6UXd7vAFpEoidfVy3Wheobs9XW3zP7omT7l9s
Vqi/KXDCQ3W/Jonvd4krTcor9xUI+LAo7G6L5Q25aA21cUeWZsKaIMijiFRolmap
Yw0AaMQrZYJSkk04XDEUJ7UPzOpfaLRPUfWo2MlkZY3cLZo55fRbg+MACuKEZxm1
wLXPMhFO6Z6gZJ3xt+lOxVWsFIGuq4t7THTY+jeSoSwxetPQGHLdtnPKSjzlT/Yw
GsyTV6c8BGumXT8HjVnZUSdUuSxzBqUclPSHavRgAJ9NllSXyT8u47CJm/pSQa2J
eaF0G1rQ5uEqisjj44X5Gv0U72eUhN3Lajsd2AKJB8F4k3KKzH8fMg+c5kF/VPwc
VC7yjrMshR48B37pxTn9xUmWiz8V61dlsmj7w9yAyddwwko6bCxQyjvFhlPIoJOp
LSD2OJ9riOhtJt8NmUQYe6WtU4RetZtLdP2q9hEvdCqpNMcwCfXM+bWX/nbHReYg
TFS0NG5dmDIm+8W2g1rruBHz9lLlkb3R3amqWgnzPJfrbbqyqRzgN18+70lGCxZw
IA6YKwraYWihR4vpUiasNqX9L3tHw9BC6S0TIq5AGQr6WPlcQUbeEkVhOhDmAM5N
rVJ++B1mswRBQMu//dfFOSaUnj9IRviJ7RmYc5C98PRScpk9Jor4NljE09KqBHD1
qoyT+tHxCtoDhmlrOxig213Sq9hqHyXGQqdICH5duTMzf7XUr0BtuWl94aYo+xtH
Gd1aMvfyadmJHXJFfFEzB5EVX8Hwb9uNFotuenZ3ptRiILvFGSNf3mg1nitWqpDj
gGAFIBL5zy2yOMBdljspMza+8YXeOweRonhBYmLOCZzWZaihSP7Zg9Jq50V6Znbs
mv7/+x0qILlYsK/PJWaj+QpZYe5g2iFpCxeJf58Fv0HqqKesmR69URaDx8uCEBiO
cAA1ma0FVmFI9o7STDMiXtSwUPJurgDunS9mRco5bw5ALXGVp7AtfucSn58/9BhF
nG1AfXyVE7P2nKA0c74OQ2cmI7cX1IekRjOV2tyoFLViIKmmHiBU/5+YBeeq4X7w
1iwmAs382bi2yfyWw9udb4sDl7J107RmYb57XDI2NhxWgBtHPuP11wckLTQLNue8
RwoOZ9eCx/MU4ylF5gUw1x1xFIQzWxw3/f9fwaIc93nCeXYn4Mzc/e2d75VXrFgs
z1Sc1vNIMjw2LKSZJUbnw5A7QgU28m0NgPBp0Kq9nlo5u7RLiZOMiLfkUCL9/fEP
cGpiT85aBkqujz/K1WigVPcCwa0IjfmBl2H+tvdKuHhTqA50yFXNi++ApUEbuGwJ
/zIc9u0jNyBAMtr1nFF3Qn/LTSjumii9TFowsGegT4EgetLvcpzyd15gwWVbM9Wl
Hcg5DaRBIs2sD87MkU4+hxsathOy/QdHk2dDWWNE209JIxrG294cOIgM483n+qXu
J2jNrpK+SR1cEz9NuU6tEFvkm3JvjvIW3uzuCAHdiNZHy17/za5/OI7oIQptf0Xt
1U3ranUEKBNLtwhkoCsVmTh7IVB1mntsVS1bd4kk1ONeDGEAjDWkUbzlz30NOIk7
Hp8KiBerpTmwTNDkS7CUuzuHNcEctDi9RBtrYObwNMpm6bnVacxmvhOYmC1ewia2
1+IlatKiYiSR+3SqpVJEZy2IrmhCwyzyHy6LoPEeYLK5nvB9UFKZ8qJQKFCp7Skf
6gEo+LTm42BX+I2KRZ8qPI8U9hdPg3HcCpRovagaTorYcoxNKB5jhsR5/F/Q2K7P
pOlKrZM+SihlAR0iWeSXM5+s9nIRSyuezH92U5LbnwaOqgjN3JMiBWBGNt529i5h
W0CKkbc4RPfBowiq7vYozx36LFzVhoaezKca2j2BnMoV7az1ErLMT8ixjEAM3vHS
N3qCGUPXlVCillSBia9O5tOPaI8PJou4FoLZXO/YZ+zJ7BdIL3gnq0lx5Z/E40p+
AqMdq3GmQPBYBMk2XodPj8M9qaZFcGwf+5XRbGXNy7bWzEuaS3CQEDsSJ3MhRV/d
j0Yza0E+vSgzUXftOSOOrJEHeRp1jkEMIDSB9ecljc3nlSSAGwWKFgLOP5rC7atC
qH9WCluda124Da9TDn0aYRguduME8KDV0G+BDiGNUJSAYewU/Hc3mpNjm9rjANlf
EMFckZtuPQ2D6JF9oPtOVd8rRilf7BAlb4fsj+ilLpR+dIGfb36/24H3jHsiemWa
zSDhzDMM9rHC/NqS8B1AXC4urUjucC6+8uKM/eSq3t/UwB6fcbcXg59RmXnJGXW6
qpt12B23BlgG09DIPhxHCcKyQXnAARZe0rRqE/qqTdjedb7WWqqwPQ7ASwtxIa/b
RcWlxCQSfbHNzvgomfh7N+YG3GqEc9Oz65+1d+ZshNUXXT4rHzn/ZJ6Z+WlVzIgQ
+h1YjG8zLVxbAM3Tg9Osb2dDuHXDKZLG7A85rmC5rNyN+22RppNC6zsHHzk+7iMt
Womfq27gK5DWO3RZCN00PBJ7XjcpeUBUKi6pxZjiNe5ml1Yt3uvqC7EwwK2reueX
bVrUVQdndET4IDVX/IrLhCiPHEcxZvhoyyWbsKnjGkmcsV20Odpud+1y7IFjh0XC
t5NxXNN7uTOE3CFe92g1PJSK/w+MRBU8BiwePSRLB7OfYTZz4RJicm/iQHOSsO/L
krMRkPXqjnoOOwdVa6FzT2uluR1rZJqWDL0+ELlRCjWaXHaOg0784HOhHtn6Naye
GjAKIzuBjMOxIsEQyuD5ikmSpelidEFm1tEHesKVzLPa2X1JpPuLVzHAM3gt4WHU
7iOJuULmItADKM3qowIsnq5jV02iLA6d/PDbhrbXgK4GlBDyhKVDHcrkCt7L/wtS
JmLr/ZQNA70DPTlIepwmbvcb7rB4x/GVIEJaG0Hco5GKcDMaFpZrR0IBWNBdlB/o
YQAF69YqPxIbAOI2BGu44W0JI/uviQKU8KBQ69tpLaS44WwSHsoNmVNfyEoDv9M9
Dby6kf3jxleakD0KB4oA/jETWys3j6aWnHvPWnGIOnK1YnJC8kwAoYIYjcoj6nRy
j1USBtplQjrtSZrAlv+NWSPJYmhl9ZZsrzyuSwR0EcmkLKdClFrJnInj+GV3hs8E
ar5POJjBdDAAa0M3tL3VqgAkvUCoJIDn/MNieAlMfciY/rMz5vieSSFbhui9pCmd
6qIe4qFxNLH36WvGRdpKalTkJjHLxx0U/k3gv91TZPXbhSx+vrYlRo1HUsoaIqgo
Wj4bzdHFk1esOw2U06bebw0aPEUpRj4KM+nkHlBsJPRX4JYFbtVPSS6BXd5WciVI
4OL/Jg9AFHSJtgFbsw+X4EH+WcHQ9wyzQZuiGqx9ZTiaYDqMaIFHoZ4fgvXj5Tgd
TDRKcjWl/xlEBL+yp2b4tn+Xwc0fc+ClGhzUfEtjR7LgrfcOm/0WF4Ow497DJk+I
exeWgGZALi2f5d6u0SI5CrRt2M6Y+lEQnG1CgxcWDH6bbwtJRvgb90ZtOlm/9s+z
ovmJ5+TI7pR3sf6CQdwaD/sPiGt4RYTF/bIvvhbsOFM3jLSWdWpAWz4eChXVCzto
U7WyxF/L8Vm8b2HPY+PLxwaRWr6TslfYY9DVcR3VuqtSTUdysITt37FB4uJYE1Jy
V4cXqWuQhyIChXOijPa7Ij3n3DO8snAG/gTnlA2odBJMJNtAshdJI8cI6kcZtBiq
GyxnWIfMTFECJtT+zcM9+pRyFaoRBPJzOcal115u61OOzBktIpNA8DvSrcLuhj+w
IGEgKZXgtJwnHqM8VrKxrn8wMeCTq7pYVWnmixtJae4rfh+WLTUM0OmNzu0O3E4c
rbupa0IeTe9WBEfCb96da319nP/cme6XXf+Lu7lnmkoUrQYNU3rFCnnta56QyBfb
TqEGm/hnpgYJMDl/9Io/GNpA7hwJvV/moejW6lJ35IJ9UJL7cuX04mG4ePgNtiI0
5F9ajRJn+P+Y/065kq5I6iHBP3eUhSkT0AcFNcYMANaV7yB7YbZcyYdMaiOx6jsO
UYSeTR1zY5DSB/5QGk2FDMhvY3mkf27taSgsu27O4qQ8OL6T/FxnFyZnfQaQc+Qn
IVGiZsrw5LJ1kXF/DhTeLuYvV0LOTvyj3DtYwx2aeXH1dr/E72TcYf7jLug0bED8
lhwsgXqoh3s5nC1//PjdMQN8APXvaU2g1Xir0vvREDKc+bmwNXjTPDIwEvWy6QkJ
w9Ooiyvq0UEB4y10a8sB5JKczoUiO8liDyVI43aFmZeTZAyJKCPzQO9VJTpn9YXt
guEe6X6WNd2JZXPCF6r6wV/My7+qqGBYjesfYQ2m3cYADaYrmQbsB6V0cajRYc1U
xTriVdNUJxBDZGSjK/UUY3YqWMpUlpSevIM5xJf0nMItqoNngY0i5MDO2OXvOidl
VAMeW6WvuZE41XiXuZMVy1K3E/mZ3Kd9ovlEDQvf1oZS2PMGxUSu9Y9bClMfeqwW
Evvty/2H4jqe0rYLyzKJCKuFPhHR8fVgSzeBkeWItyV1zppHr5dMkd/K8BCI45cP
L0fh7BmH9vKOTXC3b9o+XduRJIiBKb6yQ0wbo0K4g5DEb4DF0LeDOF6D2Uft4XlZ
yzjuHuZaNNqP53lMZgt2A8nOT0ImZ/amYhuWX6do4CJiEbwhJQoLsaK7NBAy+n5X
J4bRgPqNgMNqo23vrYyjpJ63pqDjw7qiqLhMKGZHDHSImbMFS1VzCBcOJHc8qJy4
umZFidf1NdB/B/h7W/0Y35+2EUMoG6mqnrwjxF9HHvOCD53wpDfqOVBPTicPp8TX
OfEIFQirF7BUWvsiP0GBdrCKd9beer2sgFG0TpaZenJNmJKbVaJcvpYRagiHmHoC
ZtKp7+MGGQlRKQiZN9TuftS9w2w1NQwwan3wXxcsRdW4G7zvD0c2caARpcZ+L5gk
q/X6nB6mYAExuv/AeTk1/1CMOtir5KrXk3ZbfousPcZxjqPTTIfObynK4CMYJpfP
Wuf+dYt6nEWUYTbQkG/aeCI/3GJI138O+vanEO0ePZlCM1NymbUC9VvmVcZ0utUs
hITHmZ7qrkSDOjAKotJnPNIUAlBE9tYX1mVdNbdXwetAJsa/EzkZfjWNG1ShKSVZ
9jieSAOSgzfEL+s80xWtSEmQdnVtn1csSm8ZF2ZetxNtaTUSNwAmF2tQSXTX8agl
gGCr1qH+02wYl95zA6Lct+d4YOuwBHjm57MBKfeBKmeUP7BQFdyq3/FipUM5Yq/U
5b5iWgls/XHdoh3+wobReEZRBd++harhir6WOdp6g9qpJ4IPu6fdkDHEawA5C6fd
KzZNuyxAk0ZwyshSX8qVxdaiTyzRtkoS6xX8sEJYqtRIohqR7W+CL9phjPiXPmbW
hfEQi6IqqgT/693ywwIm4wk0y5DCH0ZKKVUu2u/zH/MAdPb64eBTS58qtLdkh+b2
psmtKCDWlomPSs61zEIHep4v26YJ6FmfQXItwBtgzTrpyYBmy71sy6L5c5GMQpoi
Zun1BGkzahUN3XNSUFTeorgefFos9ErvmV5m3X6MJYRp11wgmKwkIKBSIhap7XQc
SixmOdrBVSHBeHOn5KvTuoZU9aco03Zw8taAIQGs/HgFUe2uYrJRAlkmyyhXTCpQ
sJ1HWV6lrtXtgE6ywLBX9Tz4LlECL1tDboT259/pvrN6wy6x+xy0D7s4kVvl15+a
PpRfvLr/a/YgVxX75sa8D77wixgrGiiK8s62PUa9L16/vQ5T9fAm+LeY60umKGNz
Y/wThrKtJJ7ZB1fF8PQtVWSajsnDZnS+SSxlgkd2/2ZmHg9+VitL47C/ijJBhq4J
7gkPogXIOJbr4xw7qK8Av8FNH/XspHOPyKF9HSuyHt/SUbc87n7vqILQ7Tfe1BnI
GEWYI4VvV6C05aiNGKu9/XFQsPjV9XtFIxWFwS2iSP1Zwil40VDZb5WdDtQA+FzD
tka+YCgWZ5J5WUh8LwSdD25QFQ9d5cIglYbHskbTzmmCDNElVRUoqPLtwgGq2puP
eC/PQcVZd6AZ+wAcrfSXcb0zI0kwe/oKI5WuRCbUzo8BarnRt2P3j4v5TVlZ9gtQ
+m8rPQTCdmTWRvbMIyHj1aeEUSk2LMUV5i4ngLtqxmkOAnxjNC/opZ+3wMjrkFby
HSw0psKDrmney/+PTkWP2rvPkqj9ku2F3oB8brMva9hVYM3EJlukwMU21g/jlRVI
jdNY500Wcux/8lvMq/b6DJ4mmQjZikDf49TlRzFGlbCJnlSllBCURoFhc7yQQbqP
0iF4Z5ZEM2Kace18QiL6liWo1ZSH4N/Pc2nUq4AipFId51fsymc/XEhhJTa8qXaZ
kihd502GmwuiXBKvKEleuifjY9wGB/zYkggLNP0TtEbbAXDLWK/c4jOY+UDaVtWr
g9DjSFYvPJsSBcJmDEv9zLdf13lU6xOLSGnTJvtdwn0OyYXUNfNnYBmB4gYSJ7te
16C7miZ0Hx88lA3wxK0Oa7DZwN891Wx9HJ8VX65J0rIX5nmClnP35OXmU4Sq9sHB
NWlGdtLvYXPsswF2yMvTVfI9MGWpQ8XyeLhZXoVOr/L3N3EI/mHwbbsvSXTUwXk1
yJsC2kmO0w0GFifBv9nACiirMg6BJ/KjTjb7aABgt+dVm9usGGGVS7TRXUtoV4c8
ImQK/48t0UidaKysQPuqbj/Z88LstzgAfwpUHoUGS1487LT1zNTo10ep6ljZUiM2
PsdHTMjj4EIqh9DfeCJ4CebSv2BnkBtldeRY/E9QGNg59Bt47K/2mcdmPyLMStfN
cdctlp9lkRnju+eu/LJv8RAmDw+ixZgFYDJhHmI5uqrNvWJic+411GxtIk0xI87F
oPKXbsb9YdInmGHxmfT4vo0fsQ3knpGCL8r06e41kqHl9j5IK7NGJ38TUgkw9vXG
JNntc0h65ECWR1wuAASL5+uk8YswadbHq0D9fbFsL6frrXPR16n73Y4cjLLwIrdP
hZEpK+SMiUgRYcaeI5Yd/v/6kx4Mc4AA8rbiCblLMSXi9KNa1OWGahhMfITmtx5d
C4M7cXOeBAyUI/767SwvDQH2j7LMMQGVPchRQsyP1ZFRWwiBOTRo9AswBGfpUD8H
ZoCBD7lB480bGKZ7kBur6OBPzUzWqkD8wsDodM8QIUGc2WrT/Scpkpf27b3+3+Tr
dYgARwe/d2cb5iIK33cLbD1vtl/O9xeFzkvXKnzVtKtLmRCyJwx99ndCWUa91l0K
+jIO7NY0cS6O5c4/XTa05h3jA5y9/hSVSV41sZrWjsfrhqNMKFHbkBuhpUYGPew/
FW3weKIX5M2Egn5RQMq9sCKrdoXIweQUOCQQP+kmAjpz4aiJWCUxNNghGbHTCc4B
wA+I1ShQ/xSNp30PMaOD4tJcM1H0p2DWVCp6wNYLhHYsavSEU74t9Y3GhSV6ifLY
ESe2iqgwSp5SeHiraDWifmwxXmzgcj7CWH+wiwNFCgF2s+b966RVAJ2Nm8gC2HvR
33/VQXTGJY47P8F4pIf14pMJKUEM5fBwOGyayVt7OEFcoCYa9FpaFuZhSdjtSTZt
N8V0oq+tpJHkFfNwjk6/Zj/vKZ3Oypq3Pc74TIRDzhA7nhmR9BQmtYlTTL74+3WU
/vuVg6fsVUu1jksMeIeYqepIhHlF4lEd4AzCgzKa1IIF/cXHYolgo44hFk2dBfTA
mqDYPDsG+0viFfCdxA/ZpZ/CoOQ56jTNajQraiMCG6dXnbNhidXjkd5wNn5pToKb
xhi76zcqjw4AuHTTvDyG94zXxZrtTQwYAmKoHie6sXLHJ8VN2FaTOLChaxBewBdt
yLOyZf+hIo0vvNU5WEaA/b9z0oIr7D08lrozZrMwVf5ZGukjpCnWW9NXgGy49tZM
iGGRwEqL2pYZliMWB/76eAMQTagqJWQ6CkWPiCe/lgTkd2gFtO2CWRHOm26DXdqJ
88KS4DHbwvGTH0E3maSMQFTv5yJGWNBti+vFGx50uX3sc0qqoar6bH7rNuwjTEYk
fG7GteP2WA/Jb0JmolFEc60TbgqVeUlT4xVKqFVkXLkKjtdVWZ+FuiAtF66QiC7t
SPtwmX2x9cIn/BNfMaFxyOFrkk5X+wZZdNcHGpZ7e2W2swNaqnhCWCWhpFz+RiHQ
Xs/n7uh8uHXVwIiF8dpAaVV8h4aY4kHR14H/YXRe7ucVGisgrJDqMl9ecMM3Znoh
l9bR9/LEirUIkCoH4/7UVJ0iqgevVcv6IkL3LS/N7GXEfvIsPdqV4JgU5L0ELs8/
QHCQLAzXXqWBUi40ljcKS1DAm3eZKUQwUmm+mp5JWZ81UGL9FunqJ9rYfHXMufuj
gTVpkoH4hmLR8HH3TgMZiiNUqYkcuLTIDII6htR/ju625+dY8mz7X7zGRdxGOb0l
WkFo9JpsGhm/0qWCyYAm7EYf+mExo3eTDesOOeRQ6roFKhNdjq1NVh876Grb3i6V
ZsVo8ao4maxcqj32FhTAksCdSrO2On7thO1DTvReN7PyhReLZskqcBfT19v7vtA9
QhlGTrvW7suX180vD2Xze/uAwpPcHMy2UX2iKZcD2pMCpUkJgMyc9xrE5y9oSE4m
FGdaaA85VHM8c4DvgCU3uSELrJw02iW9+AIzPG5MVBhmM34a7mwmmNmpc5+DRyr8
iitXZEz/WLLkvuwP8WamGLqahkXJTgACtU0ROnwAJpk1PQWcb+R+3rlpkCP7asVU
pIQLlcWcuG6oFoKHM/uiK2W3ZcUrdbfs/6WmamA5eW/C7cQf7DefrWyHC64tf/oP
fo+YUaBM47UeBked8ICmuTBVsC7uFHfU18YIgcRcHoYeBQA0/fIMqCsukK2LTa8h
nIaw5cDtaBEcMw1vXz8MPK9ew1ielGXT53+YeRQOwwwD/9a+BIvOaxDjA/A2tFTj
fjcy3zAy4mlV3qRpNgf3oKheZDdi2Gs+exbRO388o3birFytO+kEJgxbmGL2lqmV
cKpgMDMzsudUNSmXgYWPmKTTFhjxc/CEVBSpxmh7GiC1/UstzY+x6y7fmlXdxbMj
FRGMljSXc1/VcUFuwpSFAT1txG9uQ8XRUUBvuhQ7/wTPS5yjCB2NM5Uf/wX3N/dN
ddVInaUvbzxI8Nk3X9DydH2namTlTBQedL2/7aQ6lb3bKPq4SeGaPfU/q9nl85r0
vKGl2hUT0BViZW8ePck/v34HYEerifmFoT0xKuxopq8cZ7rLAT3mMlCvypMCb5Kb
7ebXnOOWdIUVVbJWMEgMJdvYt33pg8NV6g1p5BnEJ6AFIbWXrfT34UGTO5kdKqYm
TfeDcLUfXsqdKOkfSyIo2XD704c/euKHC8UzYzFBFodqj6gN4sh2yLWkg8rCBwoF
GkwdGSXYv+OL47v8sB5N22kKHruiYrAvJ0N6a/8jj2UL6FRiopuBJkqk5SEyORT4
pJEElSQ7hXSxvw6zI9lr3FKxxW+rSXVdquBdPhJJ7NNtFiFUS10EtPJokWGj1rmA
j9CRMid/Zdea4oX/0ZzJVBFnc9j+vBV0hwwaoJ77jQ1MnqCVgsR+YszyKzueRWDp
TfLu3k7/33bbOWKH7VxGq0AdDR47OdakvJTjQOO5HsOLzCNZwa7OrVFHwxHU7wP+
mwpRwyCaygkYKospDVOzzqHKj1Ye/Op7oU3r7y9vbfTESMRMlYDCMOdNJULGD7U4
Eu94ou9atN1goXLY23WvrDlNRYFkuM6x+/UlDpBVb/ZShOcK4gQKWNKAkxWCoCtr
U6c6wc0Wgv5iSoTQs70WW5tpGMam86yTA7WW1lnEbSgCAYctS60z3xcb9sDK1SKj
f7ubIXl57eaUOImubo+Ew+kxi91fpz/qOXGETClzIQsSqhUkoU9Z5IDpAo5pTSTX
0Vb61GlGNx+1NL05QVD010MEJalgNK9/MPKhD9wc7arml2iG5Om6f5IKczthClRq
0T1oU0wHcHv0qyBtcwwiv1aC4xYscr59Ghpi+G5QCvp/0n5avKvq4ibNTLCSQcp4
Lx6rqGKwI3DAxyzhO197qpRJCZ1Ic/zbiI3DZ9PDxvUIsaJP4kGTgVXNXCaPFEGc
R+yPLAp/Y/EouUNW94e8VYh+jp+yVJ5mEGXLraaIUT49u4DA9Vvlme4k7p72KG7V
lmeMYA6qEQUaOv4zokP1pyEqWn0ETZJE9kKfG4XGYtl4P0HxrDVLzyOB97G0j+ec
5vxsr2kNvFfN6f0dn8q5D/QgmtyQNkMPA2mA/0x0NFtU71denkUO44FawyDXXaWP
AehyulbbYR+sFoGg9O3Yv+8Dq5KXi0XoyulyBgRp/HKKTDCFQte0DiWPZkIpPFST
EfRMPta7Vl4UMPQO9xWmoAyKpduniEZyMncn30li6sMTo39dG1c8u87rDuNAaZmn
QUWdEjuWE1J91tRY6DOnOI9BQcgLBUdxFIymVF2cwfid4UxqYgmk6V2C9/EAB2gf
VApQ6ohwRYdHVTBdk3XCwsLb5zTk7pclTe5pHP6eTgH6C1iktagBTy+Kt67Zkq7I
tLg/X8ozIVM0FZQjavfiip04raxsQ+Y7VyPOJKEfugXafqZDiBTbJbweovs1PxE5
ke3saPkSxQeF+w8eI7/KOmdGLe2nN1kGQbiYeIAxFWljiEQL2qHUw9VZfNbeaf/G
ReCvK+BZ0rNtSKeE1ZHUgjVWGd02ICwRoazuMdtg30vCBxtYZml7vmDjc9e4MIn5
JTqJQ8+j8Z07bqRxw9KeJqc9snigNoFT6IYZ4xB/8P27eWczZqaL62xTbo14tXnX
zlQ/dKIROlo9004Iu2QtsTRehCsZnXl4S/mZr7X7189/mxkqgbvskTfHtuMb9nCv
oZvpgrtYh0Cz7d6YFUNR31khEn2o/xbj0kX9mKiYQ7s00WsER4Om3EsZ3hGR8a1K
k3u5kDC8alHArMqEEb0+6qZ4SSqVX4JsGHdAhcWg5D2dIctbZh55Hn9U9j6Fu+JH
YmJsb6aNeTKATAKlrbJ8osuA4ug/eLEV1M88tlKPthSwQ7hsN0VEJUzk1oIXmeJm
hMsv34+2MgURVkXc57CTydXatr5zoBsuRhtj1NxNWGRUoo9s+YaNZtczc2QzIXDI
ZtRMXPX4CiDw3A5mshGeZXb7VdRfXcu4SLwnMsLK81k93aTjbmzTCnvfTdZedEwk
cIPRBJPJPocFS3EyJNXVljUQ1CNdIqj0FWqEIu6BVzMpQgjdludqUD7FUR6awyWK
tCnS/IHJ4iMCDg9th7DIuRx7ELI0kmRyb1lX2Lwv+AqnMoATOSUhQEKYblOu1CyM
tHkHu0zreU+6c1+Ui+knDVtdZ6ZUyUy0Wt6feiU46onnhbByDihhHWsq9VVkDPOL
AIoUB0HcetlH3IADCmRi43ZMvchlhMntWoBsepPicdwZi/0X+uzbXiw5Ph4BLUer
SPZfg4IcvKBXv09IJjaOGP9VKsfVeE4fIEMS+JqeBs3zyAJFDN3V++6CL/BvrzuQ
LLL5+F8FlrS4U/ueIBS519pmIiaZEmYh5TiEsUQSCR+crEFAshMdEv7EUfzlTe8B
5i8KGUMNmhjBiY1EwqjUruEggEOVdO8ij26w6AYbXFNvAhvpiTHtXAuVxsebYfCx
QQGo+cCWY5GQ8W/8O1v/zGgwkVu6d04qQRqtktvY9ftrfX0zfzcUrNpWfi2ayMq1
Yfr0B376ELUmU7uis4sHn1UZDuxXtkzf74ykwIrlU4AL9GF0lofuM6rR+zVXdueF
yfyfmKSvueQnFfQWsctQ5LX5eEBD/IPBkWNhuAfPKmZz/AhWQ0syFwuwRY4zJi91
HAbMW+Z37cWQ9Nj6xFJ6Hn13TtUyWB9tQ5xMpR11RHpr7tOaqu0cuPzYkA4lgvJ9
3B/Lsn1Nu8hVpZO2ItFw1yD80JJX2qze8VgAx8uPN1YzDy4EGdo/QvZjX8LgQvf4
1Yu8MgM//WjizPVg4ZKvXVWOl3pGU2MPYVdFphx6Kl0Fi4r7Wj5QEZwvMWoirKvb
g51aDjvv3DU7ZpFf7/FE+iOWtXrfjyfB5REgmUyjL1TqT+nxVQQrqYjuFvSBmO6P
ZqhuRIHbQtqliH+AThe69c+FOJnOYgO1J0j0ppLHM/GMuOWXi6gqfyijrgWzN+eU
znWUTNwyfiFreADSUSKP8D8+pv01V/2gin/mPD+82sA1w81NV/PZNx2RAOrlPpfx
H373ZnJA1rXOVjd/E/2kVBJBhdn6TfMLOWXSSlaBvHWVPD8ZbK95vsvKTtqCKuCq
36GvR4W7T3JqBVp73sH1ZG1CSckX+WDag1RKbmT3lmap8wgP0xaTZyFWMktdvned
q/2hX/ogzrLttuvmLwIh2oR+qHvnuzmKC7zQY/lSm0aVfHtlg6Hitz5yxjk6BdCp
1XC4FxyeR/wvrOJ8BmcWjMXzIU/CGWB57ZFrTL0nFB46aeR9L6h9L8vIPt6F8I4j
c47sTuJoMV5mrwfYMZ4voUc28APyQ8Utr+Vx6cU6LHYN7FNdS+DcV3stLB+5jpI2
3LAaA8zREg96zTaX99X6+cFHJnCPc0wvxg/vIdiGtAVj8XuMKzhUXttTT+NbOQU4
4IPGwIplf2KOWsOpkh6k4fj9UX1A3tNfSTO8N/igjh+0K8LuJV0tRQkyOfHlGxTl
tSuevapVQKbjx4ilvjb8a9arfcesoIYUVkvPKtjWe+WhYrMM5hxU8gMfrdk2vm/P
CTEemjSD7oPEJRMPFmmFUvSfj8XgGPAx1/dUVhXK1GJZTGKCk2LNS/Ovj8hgZltE
pg/FLL60HFhNENiXa5OQz3FK2LZ9DnbBgEw0OpoMnu/gj1og7qdwKc/xEjwaq08E
hqyF5QTYZpHsv257Cka8Q7AYuhIkMkBFKRhIJK6qV7CE9VV/MJ2of87hGJqEV+4n
PYrKJ6PCT9B0cSCVgc+D080VmsTZiZJyjOP5JZLREuKY8yU3g0s79xn0DWS6t8YM
Umtfl24bEymjB+CGSsvoFxF4WPhr7ht3c8WIPnkfeeOkdCDr1BctVygHy+aukf2j
KsxEnC48bZvNqQI4OZAY1EBLtDIGeIxhzESGMeAJu3E0Aw7m57bqQw9y+mSa+Zfh
PDEI7hoQn++wWegfHK9OEDToI5AfZtOydeAUdqV9GKQefUC8fBHi0P8O3jL/P47Z
45ywgq2qa9eNAgkOXEZZl+eTlJFy36UsvedYRkaITJssOU/jlXP6PGifyfV+IGr1
K7YL9nBwAOfe+tgoGDlLTw/En9mDYQLbekzMAjXRaZoShitxb0YoADhSl3VZwlT9
VuUvz9IwSQKK1yM4eF0L2CiM7xZ9vJxF2sJewqUHS3gJGXXsw3w6o+ESct9IVW2+
9duPIow7Ho4D++SfpeLTtvEfnMWLlsLrxfE3VIZ6hFYvhJClldYSNXUdwhPm/pjQ
E9hFZPl69WABTvCX1vOGMwZTeCZA1ApbPj2o394qSPCuhPncehWLnTZUSfwUfAmn
wG97kGDR7qCbibHVlCT+Db3WSbDwJOGDEv0M91akcmgOVTPl4GKbloQ1GBZ3cRMy
MGOUyFN7a5LknvmjXl+57D0W+7QAfqqRJjWLd27rrn1NYzytfRcMWvafMwvXenSI
fo5fs37tk690HvRR3UiVobFKMudv1ue+imYecdg1xVUESQumi4jYtUFgU+F0o6vI
6L/GjpMti54Zq2pMjsoyhWebyqvrr/PCxBWXHxbydDfERHuBbTEOG0+jPnv8g0LK
721Frlv0WjeBEkdn3kM8vklkdZ/Yyb6L5JPHhJ6cDI1SowBSYcQ2LNQ0oXmfSMOQ
IugeG2s+QXGG9NdHWybwvYl7z7l9aB3CFee96TtfD3u88xUuHsMD2D0iCrsIOFUA
Ix1kZRDEMbKfdSf3/yBCfVz4lAaMbtdVqZQ7nlWKFtA4POkxzP8vM4rO9c3IoL6Q
CQnwNYKnbVVRIooohYK7Lf0eUitGYBMvH2u5ELX0OQXKy3uhGRepCS9GKmYCsw9z
BTlMwX+RWJGQqCIRfW3GyF47QtF9s9UotZIYvJQ6kuj8Lq/KXDhdAFHsqhLXiSDK
I0psMuTE3I7R+1KMu3RRNbIdpZTmB4BONXtIjB5q7jdxiDC86HQ13eUr6sWcYvRW
pZdKJ3glEGAfLUrypd9O493ufEN8D+rNG6z81DgsZ/z6AWXT1PSxjidUd/29wV2o
9zQv/hGWz/4xD0oiTrqjtVEq1m6EySsRF/CnHvCdkSTSbOvgZIoFe70l5NyJVH68
Be/ruFq51ehvnC4TPoBtdEImVNzsTxvWRFzl603m23v8LE29Jy7aPTV4+My9hDIU
ztmfFYM7y32sDUi6wtJzGddGfRqbB9njFKxoYQBN30ms5Yez5u84t+PGPaMDmdX/
duzpQd7CJgZVKEwuaEYlEwToYT/UwrZPt5b0mzuIjJHML+d1QaDUQFefKT/06ulp
FEnHzIv5XbV4l6eL+JNZQHyhDjQxBvrEppr85f6s+0oFmH9mpaWfDSVSZmqt42bq
U8IVZwugmn/VX+PvnKbt1zOtWjNPH7GvX8EYwlWkPheZE+OcuhhjP4jUT1+vmnZq
llviWLDfovPxNttOKPNyE24MrYXWHwnzjpOB8NCfOhlPRuNgJiBaaRu5085e97d6
jAlIN8a8cLPHpk+xxFbRQdtVXR20HppV2tSaxEkADU24LKfxwPzCAu2R40RtM8CZ
IYb5Cly08alToroajG85r7o1hDGmn52OaXHUVa3pm6hwYRFwIPfOnveh/b6WPpyQ
yKieMNPO/qwDP0klEI5o3Otkmd0ftsvG7lMdK68EF4RwSo8WA61T0/nbDYqXneMm
opgiHVru7sFyKqqYDFTA/TY7/xQwOVjQ5n+J6yTrWdTi70AzW4fm8tySuf+5O+k4
uhTda9roX17HnbmDQ4wYjJ75VCNps3GThlukvyB5g8XtYocSnVk/SgfWaSxJzAO6
E+M3+WhW1fzkxdSpbzufzBMnF7tCezKXjz5YemJdUbD0cjgvbcgkygybCHtOJWgJ
j/4Jn/u8JWkIDF5f5fejon12uuk2CXTTEkK9cMQbCxrDodz9tPPlr0u4r37BgK0Z
NudxVKKpE7Jh83rqkm3p/D4tLlFaI/lgK5airRbD712hKCfstaN73PkFPUhUwiq5
fPVmF1i57kUiAV3KA/rMWhsYFMf+nMgOOou0kDhK3EhFyxim/9D6XXpHVRzST/Fm
RjI/c4GHnMcstUMUqmyMgqQ6GksMAiJGXttqkO5722T1/UTtRN9h1pVNnbTu3lcf
5T5RmcJSP/Rahbi2hGHVmr/0kXbtC5U+zPhL0J/cVEsv3y6DDrBGTrGSFu3081Xg
L3gVGQw87BGuy/bJ3c1PlKgJsAz18H+U06v/qXW99yP2dwbU7o9qGjG/qqe3cbxX
W5kUOKxPM70mxmJvSmGNwcT+jpJw6vHW5VTcu7gAHzxk4c4XNHN8Tk6wriK9/bip
BoLA0syS+8VL6GLzO3Ka0RmxNDIhKQoSr+nOaXMYUC4/v2jPFPUpzdRiqNN4RdGH
dtdjfBwKC0euQ7exmSP6ABIjd0zS6OdDb0ogslKP3iaO9BMVfEwsu8Ai58CjqWZ9
EZUMCS5ltJUE3k07sLy+VrXIxVfAss6HT936/DkPNcgA5DJZzCLeOJENR02dVru6
0n6+/JHQKBYMn/YFxahLgoRsu3r4ICKPAsrfJYpw69uniqTpvvgcp1bd6HpVAdkP
wl6eyrsFwyZA/eqqywsUuwI2LjuV0+8jm63LC42BXRR4kUEE4E7cXLJLNHItKo7R
0Gokt+JlMR+pZ5qlFAbkS34JrOC9IuXwWiUmizm1sw0npbDoNOlYszydXz7hQd9S
YXJdLHvlH5KBQqWObDUH6zGME2sd+m/iY3on2DUVK5HjwdslAJKt+/8UjRwBg1lc
kKMPDSM96HSZjHTXw7o1xeNU4jm7hnAY8r4iYnsrRdCqAwfg7A4/lRALocBmuChT
Y/fJdb5JMCw3OfK7HgIyzMoHBB7MTQeCYg+vgmM8OKZ8dVqr94FW27BTKNp8JxtY
qsXWdf4KQ6wf8Pj9mPfn1DG3tDuiXaRhXDG/cuDDOJ4NPIkFrTG6PSz3NcqqQOK7
J7l5RuQQh9UqdTCd0j7RbWK3/PkM6dxrnnO/fNiRzJas3ywkVA0s+3z9fYsag8WD
9vEb0LnE6cyTQ/pzSARcHR9wytDPwFasqFy15uYDqdg/J3XTgdGGv+9k45TxP9Qu
/+ONhry96lRhf3FUlpGQ5XL1+uZXz+osJHT5W1zyVb0kxV6jduSZYMsLMFVyorPV
bJ2cmZq+T8Nzqtb1jwoKBPq29HY+dmWUPGVfVUELKePSjfVkuxM2zMzWchdLj3Bd
VIlnaZEn7g8h31g4TenyHBCjxfYFyaG1VcgnVX/3SR3vSoagKeCtpe2tKMZZWerf
SBCZH5PCjSehvLX2wYAVXUKTGQ/Nh/3rMN4fMAFhaNl+Sk1t+aeWxh0/aYsd5NcV
E0b5TFCRXwEYt/d7wlOzo6zXlz/tpt3kjBuxn7lhLuU9KHY7xdN1Fo9rZKv6JC02
fXdQarOHlCEC8OPmnqs7pV8KI3xg7LX1dVpMy15JYymLpYhO/ZWzyaInGA2wMCIi
u5wD/EXxLi+Ait5M2dYDS6PudU3caNpZBOAju1QL85EwWE0n2WtenHHL0+C7fKof
gTGmMSryYLBBeBelf/csvQ0XsQ1c3jah9tLvLSlznd/K2SBu+dZoE2PP9n39b7BY
MipjYUdW8eESadaHeudEI27HcIUdflOginjJ8WCa9DNNhRv0MBqlTEgMxi+n2MHn
3dOOuVJBnJjTZPWrhp5tzIdy671eebpYylZtCRSchcUO7BvCkSVOF9SWevlxeEhX
S1sty8MEDVNSb8zVjEgEXnhoVhKGUAIxfRLgvIQ6AMrOlQczdglpsJGCcSiSrVUJ
dUjRmXqCCF8ysTihuNtVs/AgB5b5yeBvwSnQg/YPdaqWPRPeDvecEIh91u0nhmPK
4rkGgKjnlA0PDKwRHQnFs0DgYgjE2wHz6T16zsb0ZjwtXB7UuwbQl9Flx+adA+w3
Q5RYvnlxoJ4jPyxeb9at1Vx6xKEBvSZBJ6QjsYwF7tjuubxfWTmcWc8U8GO1+5dV
m5WTJ3elVoJ+m7BBK/Ez8ck67/TLyfVmVuzbKbsccOHRXX7V/KNHV+DjH2YfThSl
uGED0d9LNujlEUSSJHhEmvWew+Xv+02e8OLIXnI2rnatAEffUkIQJzc+6WeVL75t
JicEvyrwYD86Vf/vMuYzbpkLhG7qS2oMaefacT/UHB2UH8ZabuSPOus40/h5UgBg
C41uxl95PpS3suEseynHt1GH5PdVVQIB6Y/FxhyWrpPOVQt9jWuQ2LDNOGac7udr
3vXacF7KvztWs49fX7ebPZrJ441XpA2c6h4LfPDMzY2WXjCSyL++F68AucXitKOg
I4BoBgmA2YLgJM5Kh/m8IgidHVHezN8PW4SedX5XL+Vns1aDWeH1dtAwzpwtB5bB
F0afiFCMXXrxKMs3wVfm0FIRRmKvR7BAY+Bwr9jlCo0Zcl1J4SzsG9wtYPauM9/z
TlVBGRhZtvL4AtXMtrXarxYyGqudgn4jqFZfqnqPcUW37UNlZGgXLKhKresLCitT
rk0PcHW1SzWiyWHUQdHGGHfcXDxleADDdIrj6wJD/utS7OiJSJJl7dDlFUyIbKv7
xsknvQKeLv9FvJS7rYjmPwJoV7nmxWUGdsZndfyGwGKFDcqkpHosPys/qMUWj19m
1DQ2f7FdpdACov8GiktnJueygYBibazq3jv8WDnKHyuQaq5NaVe77vQRAqlpLtpG
5lOGlYbVORkchMITJtLNalevsOjTi493IorU5h1p9w+9aPtLTunJhN/FDuEp+Ai9
NAL1GS60Z1AOd/wa34PH22y142dH5Hc9zjYbJUI+UEy/s99Z6j4jEnzFzc/FZj0/
vVD7sfUw8sWyXzPGaoscgCoiyDgwAq2RMAcUPLl5TnntPyZPt7koeXPy4nnQ5YrR
iouVYz/d3VauVYcNuwIZ3OmzCST5s3y25VBHN1NhxLKnA0gvdilGjvNDWEH/Q0ff
r2TW0urjTa9DH2uL7gW9blVxW4KV0oj+kpNMD1U8Z1x1eEcDfdcyHxJjphY9ZR0A
1E/qtCpHPGwIYb71ay8dwZsx/m1rXkdwxB8hW9AlWdOIl0/9sCMoKPjbS+NQK62C
Wxbs//ZbMOcFiaQ+dX+V/9DsFvx/4fdADh/L44EGyzF/3MbFSe1ef9t0ose5xL2L
Nll1gxWn496z3sXDrNj6Dax+tDlE5gTtfhDk2K8KNcfmoNpgPamfpO6onSwZnfWe
auLBNd9MXsjR7tP0CkVMgtLKkmrPJ3Iny+rstzQ+tGi7hyQMe56RjElhe/O5XF5W
vywCzPAIc716V7hixYog7V6GfKIVSwIVCHT4JrSXsJGDTHFdpTMVG7Osc7FcO1sG
suPeADKrOJifWYXjH6yOhYLU+2TzSimXy3RrFV+uT2sMwRnihnJUDeq4wyLexmdf
QoSC34RVK89a7/LqoQtmyafvBGCSTIlDlZDg081lzZnMad4kvkffn5mAdgwWWo30
71NmBBY5pILyq36Ku85i3tffiIZZdVdkgXSzmSrokinq9k0J1hcqmm0a3ezo7H7+
OE4PF8e5nX0iO6dqgH3LdspI0l7cZ7X0/NusmsWa8MQ/0oZntRupBqHJermY1nRn
BPLTM5+h1dwwZYDyiPdMq99bOHbWGFRDhVF5GcGVkiw9aRfwEGMfyxUTLymZFzyf
IZjpspO2tkQS7KFwdVEd5Cj6qb3I+greYouQeU5eoPg49kgCZbbJ9lUVRMKo6+PK
ttV2h//UzIm9zK8/r9YaKPJSgZYkxdE97CcV8JT+V/+RbarFFWI7SMCvvk6MuUBe
hYz7ItZJl6yTwHM9gNS7LDjZXRmjKmiq7h0R4MHZeNMYhGke2+t9VP14mqA+a75+
OTzbvL+DdA05eYq7laxtO0Zg7+eO2jSrwv8D9C5f3Q9NweFN2ze5DTveHH2P/ZmC
9TRajz20E5Kh+Am1E/1CZmsB7BWOAWvlQZkvLWr3QbBhUO7L2mE9k2Y/x8G2+2Ny
WmPaKktVFetph7gno/3UEB36NsVzI1u8Uus+KD3UNgM7Xg+3DnCh/c3uMAcawrRL
UCmCq5C6K+1eJJl68MXB5H7TheYYVCXkAeDmP9fASpYHAxHvaxifMiHeJxjzbDdb
u+pH3yrGgSsEYvrsBHe62U6G5B7VgsV4o4Mq/HwkTWw8IX7IqybeZnmmPEtFQ7RY
ZVovFWnZzbbZWWxM3pjDLxlX+7DtbpCpyNYIIyAv0kyGlwIi90R/olKPkHp4HYhH
N0EWKM4hK6A7F2hqm+QBUKHFfeLkdgR51EPrbdjiUsCWGkfCH+RaZ6Ntc+yYAi92
X0l42wY4IZfXUgG9n4bi+m3Q5OV83UPHbh/m1SnXet1Ub9/nAgwz2n625fOtvKyn
1fN2VhE0meWTXfmYCJDwYIo0DCncL+ofSWUrEnRpL2trsSIDt7UGCW35V79E+Dyo
sjCzOgd9L0r8G0Q1STGZovkFBauE9MVrG5kKM3+kc2wM1iXw6CzeayP4iahFrb33
aNRVmsMe/8bjM+pub+kJG6gEPbHrdQXS+T4W0SO8THhDsSP5fMDSuwXmR6k2ZXvK
FX7DCF/aDkJOnKuL1JEZBvZrN1OHjRmZMQcJB6KmXrmp5WnCu2sevrgaowl45kkM
7pW+gXasDaS/m3wquxyU/aBfmXgT0mE7DnrJNhqbDh1ZmyO1cZjz8DZLNIbVbIXr
c6EwsNn/aMxN/q0cPohVmfUQioFi6IZxyLNhAhHz9hGedMEUWQ82u5sTLV/jx3am
VoOKQiXEM8Ovli8fgIk3F3YKdiurUaNbc6RRlK6dx2cCFn3W6JP8A7TVH2Bk1S29
NBkzpyQc83D53fWp3kDOupfyfm+lE6nUoiQkhxHLeDFe1hDa2mtR0c09ZMOcN3G4
IYkI3fdJiXeDkOW5UYq8IOeEc5DkDAki278ldM+qJd3b6dyidq/LzOI5NnPAFAHs
Wm23rS2oby4Sm2yNqJDyXpwceoDtITU3Gh77/5eDcqeSYt7sHQ5jarLGPmT8wN8O
nDYWsD0PwOXqHte+q6HXUCYtD/qe8g04UStuyEtcP5AygqL0hlHKKnYFrdGeDl7P
jOFDKeo4He0TKRJV6Tzc5W6TmqFzgaaUqimRvJCDmF9Crd1D/jMMOiCa9k9eYJO9
hY3de8g7K5vhYdsUnVPAzrdBgYLqqrPnbvsHEXuHCOCaXJSBS2Qhr+mfEmO6XwMN
J7ux6wLPrXTOiPy12j5mZwxZej8ALXC1cKJFdVOyC6HG3O8xUvU7yeVnAyJCvRKH
+z0L5HKFbWYln6uuF3Y9UoJsDfaKxXZU85jGjdtITzW5qvR2j4zuySBLxjDEZgtJ
4q/tzBXFkqmYD34RKyQ/T6/J4PInzXZoWgP+iTA6g1acFWwVjG++MB0qSzv5QCz9
tl3SwRh4dGhvpU9pJlNEbVFyAXExc6jBAB3f0Ysztugt5xjhsRwkxG+cS+1AA1iW
5r0rXtIJC1TCY0wnucI7bjnMPXMOVsCmMlWMcN7XmanugWA3PHdiqv9GGtt1c0JJ
MRNr3fAqwi7YoaEwVdOTsQmuFWh18oaoq59dgjHcrBivocfk6+z5w56HuH1SYWaR
9RR+afSb5Vo303BPyUZ4uCoShSoiJg6Cb5OPbbN6YmQd+G3xrk96NZcFC8jJY66x
7yU4HZfg+nHQcde6rgb22KPpEokULsw0ldej9ueGJvJsCx6nGvF+R3OsfA+kcD6m
Imwb/iy1r/FENvJdAHCZl6hcrpb8nC32sNqdKSMMgffq8ygHY30SaMHBGLvC6rdD
a/ArCUW5rvz4EDgHpF0UCTXJAVdX1sfplXHSbmJlNYRxM5UzsSJkHVILsopYHD9y
vJHNb1n1F9EDjHN986MMzTy5m+phKdzDrjPhlHToQ0YTor2BGLn2uDqcKlkavPpM
bZ5LD5eXG4UGH/2CMDY9/cMbyPrrdDef9vhKwyeAnJFZh14g+b5t/NnzAuOqVO2R
S3Y4m7uLf94GWYio1IpsmaAahdaw2Eo1G0cGyzq9Zn/U4shHLHPbDKGLuodddJ4q
kgU/FyCjAvrtiigSy2mzq4QEwwX1bZtpKd0G7arcN5qitpj43B3XbSzBCJTqtfZ1
R/54WnnL9y2FwgvBwQuh38FkZy/ZGmdkjv0lOZQKYiuaD3IXGpHuLMgi1RqZa3S/
0BatdUsh0wNDdlPwhRb8JRFPBRmYr5rLSdhrWrjgri2UHv5R5tTZx90fY0KMh3iJ
KXqMnaG1R9ofwNoXKzUhBOj9ML5ZkncStXFapBhxyH3g3QDSgAUoa/YWaI7doB5F
ZaoQNiZVtHaWxFmscTcFMzy/HOdPNRwnGJZoC/cFCzX9EiOVpEHC+XWY0dMvYZCT
jyVJvpmmg/d6bERF5GNey6I6q3chz6c1T3orfNIPyk1gOBhAarT4/qq+J9qSXBYF
Nntl9Z9jST3qH1B8SaIE+3U2fkR7fiE5iiTS2P1NHVBoUyBF7bSBDiB/l81m9rTH
gNJJixT1no+tDB0zLooQbo4nfJCMxREInhaM1jUzBpRXHQG1rgBed/ovVggu3Dw6
F1LgKwF0du6auZQmNWrxgREd4ZKu2ch0XxD1U3EeAhIyUmvZJLN1f2ZG6QBy/Tp6
pNjBnXdxY+BJvlqf1JkHAdd0EuO1u7Fuk+Kud5YjkNFGXGf0MXN3QtYuTUqyrIcm
wLxzYoczQ1acTLnc9M/2D7sASL6VK75hxyA/HiJS5kvN/65WEa0l4/GpbtXXwhvq
FV/6X1tG/WUZZ4KSopIyKwixKiQ7zAyeBSbbAjDEPxShUPU1XMs6ztys1dBMd/J7
PcVVbc19qyj/KllBpH684AVMaCiWYl7N16kFrNc73O0rT+mpEUyHG3vtKEIjEpej
BfdVTURxcMfB5PcK2aZdc48w6c8zvvwosmnkMVqtze6/wWR38Do3bZ44AdKLt4+Q
1tyjWbvFwXQQTm1e0SVfVSl7xghjU5Vlaqi0URSrDzP8HRWh3QT2MTh2UMIWOqY7
pVXVPFAnN7FPZYftA2aNMqvHM0FFzC1POVOv0sUbKJ57Df8dWAJMwEcZaipb5Eyj
ZOPfixio3ZyULU/NO7qSerD7wQj1Kor8ZAogzvk9nUIi05p9pp4SycML8jzCEifI
t+S9PuB0EA6IeJXs/akhKBQK3DXHJsTcMacIP7E+lK1p702kq9Enhos7Qo39QNs0
6uPcSJPfIlA8U5x4WXky+p2t23YHs2pQNCWGcBS3I3iyOmZvAz1edEFD0a6oL8nd
hVeEAdo9DJ1eSeNku7Om0Dk9AHXepDZofugX2mx5Qi8K1/ocenKEXut1NKaKoTCk
oSXv+hPBPHdLuvjtkXt3iS6cb3rT7sHk6Mbuk4zcZT0GqABvxBXH6dLBopN/OKAG
vFcMXnh78s9mdEfaRmgLFzvA2VnRVz8zFzSrmnElU+ER0JYufTbeEaZla7TpADDS
diAl5mtgE+PWi23qUC+2QjjHkyHF2Qi0j0R2gDvvEJ9Wp9OMbZ/+Z4qF/ULAbjcI
sSIDJbgUdk9pZdrfeYlY/rcqdncRXPfbqIZZ4myfZcPBZgY0aUX6TGWUvLgr3H/v
BermNv9zGooYUmYqutgIhEajvUKp8AhAY/JFDuUWDbLDn5d3h971Sf9m8Fk21E0r
QZITlU8FONLLzvwGpC0FjxNXJ6dmpUL3nIWGKGUIEkiCU8/aPgaa7HKL8U8jE24m
z4NcHecI03sCi6/haRQr58l+M0o/pdS+Zdd9Axh+8V7x+WQsv2bRHjHShQ4js8x0
MXpDMtUcRe+2Y/rfbThI9TKcacTecyOq8D6lVJF+8zDwx4tAnHAAZ6Ah00o/+fhQ
MT0MW7FeqyGOSfYeib8QPk6ualzjWmX+rIz3zIxGyFdav8F31MXPbsvaeiRksa8h
bSC90lCAb9pU++3yR3RshBPP0Ya45qXmCDekaZDCLlcCQxHdiIbiak37EN5UvUlk
2CqUOm7/RxgreEf6kOOOKmsxtLK2XrAYucZuQm0hsrw/pxNMa4sD8hDCwiJ0l7N3
AYlFFDfGSqm3FjdRxm0OCMvgO17CfTU+kCwCe7BMs9Oa29DDNo4g9LkZ9y3s/gyk
G58PnSCQG/g17pdU0VGzyC7ZQ7NKewFQhqNxjT61DQKmUwYbmz9ZqeQLi7imT2He
x5zDGsTqhsKp4DDcOoOUZ+kv3XDJ/WDBEEVPxCMErsdP33w9FBrScZIBUQcqHgnQ
nssbRklbxBlwWMrzzDjyUQ3c3Ep107IUt75AipLhGt0W855Ab4fBXRnDhdwnjY7y
J9XIS4H7j2eOwDeyqHsbp66E/Be4ys0hPsYDr7qBOV1ykyaQyv81izX4EnBaM2Ao
ZTz949UcyFjlydUQvFhcZ7NLjKEDqUhvS52/qKwzyWdo/cxvax2Ldm0CQkB4AbH+
UzhqDBYE8TJjxryCKn+pNyqbmFLy8QIJswPHsFw7yr/hvTk6+vcFA73PyeWdbmHM
vOl0HY3OniG5KrGTyZTO3oxHPm4GA77LT4wcDo3MqmOIQI1vRWgr2YgLgbxDhIpx
FWFluNIjeNSA/bbDx6tXCmMa5k26ivKthEmUIUM0JNYxIDa5eX5f6TV0tt6u2Qnt
xAk74i5Vg9gIng+/6CLZ0/t+s7D0Zsku9fnRMBgLmO5/iVw3ySd4x6aXv2aD4aQV
Id574hHLmc0Cv7AsmcKyY72mM4GZTqR+KE+lZUYA0es0NteiPU2MtzcfEPUm0Lrs
wjAJLy7agTM0b7KXh5t3zAL+zm9DuZk5LaR4j/lU3S2nsi9QuZyjTRHqnikk470O
zpQfTyyPlq/7IIVjbI5JpzX05n62bGC0GQcq1TyZj+wv6clcvTSapSxa1jVS/fVn
3EhcM7y8ucPUabobTn6I/IVBof3Fab1DkLdYlTfK++2bFtuTNVL9panjHu0OrVjI
RWIkPGMmA3YnX2TvkUsFr2dRCEhkB6+cMcYBDajJhZ31Mz/nJF7ohGPjFrOJsVd8
S0oUKqq9S2yDvCMcwr8zN8dqZkP1yl5dQgbRAzodM/rnT+1H7b2i1hffMGDVka98
SAms7u/Bydqh2o/SoaAmfTPx2Ceaeukk/PjgMBEO+UrVPLs3QRDxtN+ueUbmq5Mc
wSNIcVfKVKNuyidEqN7cUvEtdQKKlAINxbhaf8276uic1y/i7ePBSC/bY+9cXTUZ
RU+PUNS3Phk5my2vo7Z3XjoldanA51AgUl687q2RKFCLDrcpeu6XhsG9mTaxWLG0
I+VmGOSQk3BMeJOnTLzoCYuJDBzTo+WeDxWSAuHzKowPEhB5KQD8PSH1BrzXnawj
jervf0iVGHuqmoLNyjAGvhO4FQoD7dJ5cyygS1so54CrgamLixUQAtnAhkJmb+dO
fqscrVzbOk5ijzYwL5SlC7c2Ea4Q1z4Vte6SHgd5QVk5taJITXsbF6DzCc0KRySb
GrViWxVtrRJ/mGaKqWMDGgZT2+bHci0Cxv/oYDjBcO0jXdm2wWPhdPBGTGip5oaY
bVZBxSCg0sfZK0ewmBSD/DO03Abcc3vCEVIuyhY0a6IIKhe80qp00rkKYqT62v+L
pTZ+HhXNIkmf0bnGlIbpypfi8sltD7mG3FR/sOuU3o4GCxpnm8+JTk/LpSMbTdfC
NbMWLZXpmG3kK+IhwOYPuc5ITNpkKrLQA0iA5EtZ/4WaN6VVHReHdVrXJIiEoQtV
eLC82FDi8wO+llnynnRBKLZWBE2B3F5hhDQ+IwHuCiLD0xXMF5dAcqnbab41Rv5/
06D8O0FK2j2gUy5GBEXWqp9pCJ1QYK+pefQLkQa7ZIPsWLYFonCtLkVTlVxgpnQm
w69sFV5UZ7YgpuppCin2mos+dZWZ/uT1RCR7V8gOqBpoSGnDeoFwAuBlQQgkmzgH
AQaova/bCdjK4szA5q61if/lvneVGcsY6vAHO4MWZNkFyBtXkxiUMJelx6QeAC1f
gMaPTSKVuoVmn9zsEOoWu2tciHrVPF820cZVnYjZ5NCBu0NoC5csiuxJgo4cB38d
7108rSMlMMUgCVarm0SujjQauEss6D3RPEMD6p6wgGkGTLTje/5kPr0dN8hrLZ/b
ivF43jy3npeCRhvGzZcpJvHnzdTshxiLmayKEZ1VoaRBvPb2Tl/DORYj8heEGbZU
gUrpuYKDSfeh3AElnAC6g82NnFxF+L1jQQC770eQqJ3Z6R1ku3IKbaNsknQx3B/1
LcL4NxVdk1KTYbYZ082y1KBAFcse1aimN6dLF9HXLZV/VBWZEKE3ai0y7z7A86wS
WgyZEWzOsCzX/1h0zgI23TR+SV7QByEORHxHv4wz/hS5eF1M9ha/FOV3wncYrCVe
cnEYsedyKQ8QvM3/fGF4HVuvTu/5pcQBUsyAEOzi08JpQ9BbV+Wd5QnJvzDbXWub
bvEeRhS+UDWTaTf1uuU+fbme7eeckLSotOKUb0k8+Agg73ZhE/g3A13AoZmh3Cwu
TPip1E3x3RR1hvScpIuOqJNileoAyxlJ85RqveX2006d4lWXHbciVYR3Klj6mCDH
FeRddcITzEOdEpz46Ib0U+Zcxagmi+YYYp5VB1A2BtAo9vhaH24EwuhyJwUpYg9Z
9W3DBCFa5dIPP/PllVD+aQ3a+J/WvKbT9xGwnFMZ7GmWpfl2xhU7xl5V1pOawPeZ
+64PIDKdvbiaZPQ5k/1nNel+HP5ASYZGAa3AavK0YioJHeRjfi2k0SsV6T3TBGLd
4Wj82qJgp9y67jZsb6bLXS0+gW2abC1c2GSmbNN10YjDCJvrxtJA/lZO/4MSfmHI
OJASrFJPeVbVhOXxc7Ttxr1V8w8ZDo5waemHQx1FX66hTQNBnP2aVJGSSdGHhd/m
qRdoGOUgzAi9g4L8TFmb0si5wcqJBaQAlMs6izKKoMQAHRftki3w11Xi9Z1HjwkD
Iy7oou76NxAAtU9V2R5zX73pqlR2/ssWE04Z0pnvhNqVon1Zpy4/qMK5e+YLSZ+P
K4mQsfKMNQ9C74lPDF8f0XxkjTXw/H+TRYeOQsmjet2+ZWRxihf6+KM+2tXf+d0Y
cUF281TMVudlTXx3pnVkhXlyS+J+gH4ewE12jAFPEsQT4yZMCVeVJfD0WC/+KiRH
wkpR/obxaoR6UGQZ0Gfaj68hA9iokQ16CCaD0uNXXaDJQwyMG5XHfXm10oTE/KJq
BvRv6GFby4l2KZhVV5/ice+MDu00peojCwvnCe1FsNTf15oQJSexVawv/VYYLAjI
ZK8PlYr9OK2GFVfnH0CyjeYXKb9DD6UGrOsuHlK8baBI0aQnT6a37KtPwuGdiDdZ
E6QRq9z1EAie6KQdTAjLNNfilO1sYnVMdMoVEW/rW7zbapg+fppoxwJ+Xto+geNi
Ba1aLtK2NzwnVp+IiDNcX8XjHIwNdcDGIndlggMy4eD0mRPzVw7lADqrTOB9X6TG
LKxnwNvOmgwrO0eN9k5j8qwnnrKO+kaU1GBn3hjgHEean+qeqM5MY6JmP6NAMR6s
RzUs2q+ZOUS6YCot2nMYgPOQ2mw7ozl+qHgeuX2cp+npPuhO5HE1LT8LVIL8EjFT
drpJDwdFTN+Sy4y9ut1MoMTg2HLHim2ZBT1FSn2m/6muPQfMd9Pm8Rx2+FVwBUfg
mKTgh02zwbYdsNJZV1O15Cp4GWiWHHAE3wKEdPiZri6tM/N8nU4nQN+nyX56e4Uk
UbiFndJt9cBjEyU0vvhGgwajUDBuTcF6C2ppEONiix3CwLIuP+JKpPuKATlm7jKn
l/RcFOGGZkj5nHttQKLg5Ujf2hshdScRIvTQQDr6FvenBJtR7bp8z81Nj1kHWe5K
mZo3i/Mi1eJ7j/C4kNY95KpbWSdz//dj0E+SDmE93Ar9FGS4riMcETAO+vFBW1m9
UTN9PPM1iTx4sFstvnrvh61bAfoDnck+EMuSgy6jt7lpQSSodEEhCSb8+GyuUMz+
aFxgidzVVj1hxdW/uHjdYs4xuhvs3/zF6TBOtmb2K/4ijiUxzrR+kUpDvR+vtpyu
GNB0pak7HNvbKMjFiT6upKf1YKaHq5KFRfIYbiVsAPER7dd02Wennbggc4SJvIxI
85zNF9FSO4Ur7lKHfydnkZhudMTdPzxi+BQm+XvxSNCdjfJ8O/8b1G7AGcozAYzN
wU5XbRLDwWAyZbc+lU0o4O1WPQzxwKr5uqO5HX3+d4wzsIFl2Mf8zUJiw6ve5snD
Wg/9y0EH2R5iWuF7QAwLZOwxj+j1vajTR4tqOpVFe8BxBqCdm48BlVz9Xw2cpzKf
CesO0ZgvJ7RLvcnQJJxwxq1vqeEv07t8suqAX5lpTVWmP13/lybVra0FD9tYd6t4
F2p+Ke/Go0uNcPUyyS2AKG3SIq/PPlIWCLH17+PtDSeDYnHrNayysIZqiYwJM2Fd
/zeOYs6F5ZmM8/xAwQJGId4NU+fOHzoaMwhtxOxImnxeZBGqiLcyBLTioHpNWxRd
BPqk+T3owMV9ZrZyYmGoMM6f3Vnfh92fkKmngwJ71QxB6qVJNtSzv8WRQq2Y212L
apl4h10THuTOFbglL6bpF2asaT6z+aec3ZU1/TFmCH8pfw6O4LhnOjj86WYE9dTr
K+ano9npr/OBG21JNWEeFT/FgvBzfShDg0i8z7vc7YJJw0szjLXlzv5TAVUyZd8r
cGZUrJyHU83vieVWC6ZkfrFtwpIUEIcGASA+PznUlLa3h+ucFPNWsBV4N45RUZOP
XMDallm5UshFq7BKbrE5mjgjFY75FOcd8vyQehFHTfC+qOD9uHT2DDH+rwF7FA3X
RbSRdyMx6TyWYgZOLNcsjIv8PeX8x9jubKmsyCHgZhfeUjNryuEQyr2P2+e+NSH4
kawsatp+8WrMzS/z/mumw5PA6dUjcuYZgRXs81/WUwdVm2Q6qp4k+6mLtriL4rXZ
67a+8zZhz0iz5uwt1WTtk5q2HcwM8YmMikcOJmbN6jjAaIxeLdcinxqY61DW6ccf
Z8HgGjBZyTcg9c2WOWuK5eVTt6iIj4hZY1NYvqffHyLHOV3v38E6pIg/47ZV/low
SXCQZZ2EjWBQoT0XPhvBfTHgpfBs6d5lDIwhyjR/zNkgdnkKv9rDKDsUcJ/F74Wr
pdjRtgqXv+dRIPePpefeBIYCtRytJLC4irM9UDKmsisi8rg29kOmr+mev5cISrQQ
v07zEcRUOQ5ofiezBnLfM6eHSa6JjYvFWlEpnaVQS7+N+CSyVVLZOsFJnAln2VZU
ilfLFJjiOvCbj1I6G0LLKTyxQz/WnkwQ7iA/wqKxYb76cltSF1MObT3AmKtCVPZq
DcgpfCs0DNQcL2CwtmjHVAFl59K3fWHEOYKyXYnLWLLZvKwl8eIiMnmL0gyydc8v
34cNwlBo7v+P587zCMcrhC1oh7WCYyCyj2CtbFb3ig9wxYJWiBMZ3+PLqwHpe7iu
drwN9URVYEbWVtGIh6+aDRU7Qt3+o+kA3ko5fVIhRNxqyYAgixZBl3AwP/7Suf6m
QNwkpsn+Agr1NVZM7lVelOoJSU4sLZAoqgTuvqqpQ0x1K1vAnhlBS2at4onNF+dj
19WyjaHQAxS4UomoJ2nqjKjeKsRCMb4CiAhc+1hK3Q/xGWBfKZbxpsgplf3l2u1B
nRJGI9eFH7VguOcnMmL0t9GV5yaeNThf0e35m6uQbgNTN8xXFxWbQtd7XxmMb6Fu
MWDEMcmhX4WmxV7BMkcEhjczAzOHa/FE4MWlNzkQsXb4hFSCaXEfFPp+8qC9LO78
P91dwbQ2b/nX0iTnzin7iRkavLTAtkWg5T4MXyJS8gfRxvVs0vAFFrZtAw9gE5zy
3WcKUS+ZA12B0m7DJzcQeLE7ghgbrp/jqb6zfXnfH5X3tUV7/t6GI6vCgMxVm3Ut
NuuA5Y39cGoZlwrpSSjrCwZ6JXt6jTMlI5AqHafTxZzAUwDEKX4ATVKAgsk1h2oz
68xGaLnbOe4115gXxj6Mp5LRsqmv38yX641YN+EEq2Ulfi/374/q1jlhZnwlbqZK
p0mUIhuUE1uK0IUdHv4onL7hNQ9pXPQT/PuxE4cROF/nK2IK4SGEz29N765/LPkh
MyIGm43GAlpCDw5hbpJL/SDivRumixseUQqeNkbnBn6TD1m1NqRonOy77S854cDL
KzAtmqslxd+5YBjfsEIJFpNZEXATaWQoC5HLRxVz2RRPJL189k9JsVke0GrVO5hR
8NhBWt/mypgUgsjojAEge4ztOs8X5DNJFgr4fDsasQkmtq55R42pRbctex6NKPJq
9c1ehVvWNIentoKmjlAly9VGhTEUdJJ+v3WN46Cs24UHzECZTAge+isx0YVHupa6
8FtRraWt1gPufjKOOds0GLuXzwnn1x15DW3tNQNpXq/jLIYKBlP5hpVbnQomiGI8
ZTDCMOOeIfhqCDyTXS1pIatKbUJx2NU+BI4nFniBfp7+orxnu6xCKxg8C8wwji93
XJ7IfeGu0rMNByHgvdJnvRX8F0eQp4aZ1Q3Zpc74DMxTL6fs1g8rUG5+UiCJJh6i
gnFZeilZ9jnqzX+uk6EVhtgTzGJs6qb4lIQjncInYgWMrHf0gsWBAqakD2AkyvWS
LS/othJqKxB6EB1Sq9jEOfkyk5o1/xvEL0+TNobi9cvCDnQSJB9mdYLjV/jqCyDK
11JMnusBk06+j0GF8eC1q+VSEeRJayePWIJbsUj8iVcPjs+md/E0TN9L95F2JCOW
XoGH0syMYpyRql8gBpHnC8CePfMFJHs1aK9fCOKxtWlyZgBV6qqGRt8xk0vKINms
hRO4ss+EYkSGE3i3ornWWz3EpWsSb36iAVghgE+ZVY5O/v9ysrThW77dB++zdyKT
ovf5AgqLSY3fZ92OyP4W+YVRcbeRaa+Em9qra1uql4a5YsHJKb7If6kmMb7VFQkY
vRLGz/kc7f13mIYg6V2ZiTnRI16co2+IxakDxsJqeugNywbiCzJ4wkhlcVltRHSN
YxGGXe7QVStOgNwTKgKwZ7sS0abnrCFw7OK95AHnaQEcxlhIL6pcgEPGlaD41qXI
azF1Ie1gcKkgA32fiq42c9UX9tImzHqKOEErjRSDnqDFbfDoc6G0l0CnBO5tyhoN
XdN9Wo7R3skrXyJudJDI+RqsyIOEtQbGJqP1US0M8pC7zNLa6VAP+bna8hNGXg3v
fRiUbFEhOrWTJnPaNIqase8Ue52lA+3Se7/rRIelsNZm4wxFv70u0Z4uQeiX1eU0
PRXStRPK5ZoV2a1h559xFc4YBwNHO5ndg8orS2gh5IQhE5/h8CTuqYzWnXFLLK8J
y7zKDWLzch5xrnq3zKL6O6UyoeQ8HyWXrL7lCgYcKLUihLqglD00G5UDqWIdYYe/
69E/cYT3fXM0tE/aVg7aC/c14Dbu6Fe7nz9B5BosKufKz4EMhElJILKjsoID4Ff4
7O97CMIX+Qsyf307fCnoEubjfnEZtFlXupFGMdWAv56bqsXZI13aZD0zulUe64pP
VN8PpVDk7CCa4dOrUxqFlq2P6y4VxkjvJfPyuOWSfBR0rhRIiu2P0IYUt7zBJeFZ
J5h7Tig72V4rDMC5goms3de68utpKMsCZLbsEuLCP6qb3FKAq5O09GDHSpLYONtt
gp30RC5/GfiElKJOKOlVqmpzQbFpAj3V5/KHYpR3HFwq0SyZVDcgpKpnKIwggBVc
L9lGtZgAl2HlXPnMGbjiA7QuLTSk/B4TK5XdCZGLPm8Z534dSpDzgKPvspQ92T/B
Kw+AMisnJ8na4RMlF2nU7VwQEsJ3BDawhzfAruyfw2CJZdE4iYu4TOV3ZozfKTzC
tQ69jTNzsHJk2FbhZdntvF6ASASbw62rne9bKdjUvYnrXgjOrvguLWGaLFr/mjQd
g7J1UhWQRuACsweD6Z8WtLkzxy9D8JfgIYzYiTTa4jjieyHYBr1o+ei66+NZaB8p
xRnBv2fLLlWt06HTUg/SSwvLb9OZBsQeOiGnqhbEo3gfrpdeX2O0yT2p3N2a1S8T
qcI97NXyntjARRpi7VFh1tI6iijZMF0ikqHCKKe+y9jQomqk0EaFYX5nztyZwMxF
OGBuZd/mF0MxXwHpvjm25AeN+zp5nhUcjW3fHWyAEiz9BH4N2AJItdzzbQ8nseXd
gS4heK3Hw2w7/xeabesLZhZysZIxk+PHnjH/MZpKGaPgmuriKCxfbLSo+sf/jiob
qKTtzdXpGvEbbq33zgIAl79li0tceT0DjDTc8XiQD1Cyb+UEf+sket1ClA8Qd5wP
VeR3hTNLsm2gqhlVr+wITQ7tN7DVX7LPjWI+u6K2HVbu0QRjBxKH3Y31boSQ/rjk
CUfnd4oROThW8+XdzlUWrjl5a8dLWsDIB0HoNAoMpqRKbLbpuXNmkWf4/YNWO98K
iPsNQPJ8454cCfhPO0nXfwFgVFy3vptXFCEERegaBkG+GdJBdycBQJWQiqv1bg99
uc2ALEVhJKpqBvdwxAh2mt1op0I1FqNDZ9uXN8A3KoCKmumFrsK6AuZmpKgvuksf
jvUuMSMHprFHF77VWzMQRtTTSaabLdF2SWfl8uLkhEa7pNDV94o3DCI5QG86fMeP
98O8/MQSRhxEU2Iz4XdYQxxzgd7UomAGvva+8rZ1a6875Oj08aayK4HE2ZlmJEbd
xP7sCKPva0H2O9lFfKuOnl/HiZCPRjXYbz8fels4f6jsl87sploN8T9oKNSX9m9Q
0aC+m7y2fsENanfrf9Bi9k3o1PF6aOvuN8sxc8wEFuc0SqDh/rNZ8bmmx/aAt5gI
5T0Yw0dq3DzXRlkS8WpRotb2o/Ea5vLLqVmtytFQDAE21SxnKT7Ew5RTfgr+StnJ
uYNkBasJ3Lq9s965IW0nJYvN8vVFZrxEV+tWd0Hup1Krt6p7f9qGClNW+jL17zZA
3PmHmX8IYlyYCpQn719PHFiyBy/L0MXQiaSE35oTvA2sdmZPdGv9F1T90jeWVBjV
5CJ8W6OkZ5ZHKsrY0lap48kKK2SFSzhIyC+iuFnofLPrLuQP1MOMfzYX3WKR61Td
jL8mnbSZ5XQXexZ0necjndxOgpe56kX2jkmjhLpTY4iB+wxqZS58GhG7WyHuwFR/
nV8VhjaPwltBCObah4B+s1Hz+Magnx2IEdZQwAjc/K8MY412HpO6sXwihPQkWOhD
sF2RADCtG7j6Ux2FOaO3EJVNkrnu92+IDBzrokBL4wvvTfSlsFfLd/SzGJic35KD
Wo86AfTuurRXfYzXezMOWA+ZpKYkFKYmoMCInZgTt6B4w96+VQxkSHEQ0swQ7o3x
yQCv/zQFYsjkbxRkoahFwEfZVxiu2dRWy1HsM307pDO31WKnR2oifMhr99SXS7wM
1l2GtpOg1UEYFX89lGnvNaWkPFDfo+HFZyBoUd/d/u7oVEWSaXZ/jZ6CQk0MJ6vq
bT/bWIoi10LSwOGIvfYz+3k4AJVTad5UKtQwOay+AZB2vl9b313Yjk9SahGw4C5G
JEW2aRSqVhsNQID6ZOtIIDHHlj5VZHKN/C43U6GOnDY+O8WJmaHZHfEAIUWjtP2q
sbQIuQXEYjqQVfUqZOChmWnsKxn0KbbWneMFRgIJs9gjECJwXbor+rsPhRZS3KhJ
va4pMjZmSxTedMDsgqw1xNhGQ3sc88qrQ0Ggtts1O0oK29BO0fhWLTr0outsx2q4
Q3ryMlPvUc3Oc7eYaijaxqbGEQRskea8ICeBDWRkm1WJiRt4TRCqkLv7iRWMWyVY
BmEGFLxQVASXFf4sC2sw+KmJ4b6wdILZgyzNuFO/uf/FkUn/dOrpy+0oVDnAPur8
cyanP/0caY8LIsu+/8S3oUTawcGCdBlU950HjUAbTWlkrOn9fEVF0X5dNRx1Qh12
Y6CfpqklXeCyemtXSP71Z/RMuFatWs0BbTngD3mcuL1yMAOI08s2f0/Wc//UduyT
q1+FO7i0WsV4mciXsElW0pwm/dnftdpMUpbGBmP88/BT1+pymMBpeG8WDmjZCvUw
V/As62zr2creWrsH4RGvJmR0D8J+Quuji1cjSDr8LRHkyNayboh9tA8emf2EKr1Q
plRqRpObGhmhg698Q76k0/JGMQgelMFbdY+EljyPnJSB3pQ1nph/7yyYRdnRFQNm
qtPYYV07ieH8OUymWgsbJzkRkKCRsD6sxFHfpckta4ngWiFOka4JNluE4K/w+VH1
SIQNM74ucYGbQFR23pDovoujSbj97qRfrDDjeG1GLqVRM/QsJ4aAImVKJHddJ8xT
Zj+oJERWA8TAD7+0KlgfSfb8Ve0fR+g+lx0liJqotAoUd3y5hbdKp6cmBkITLvNN
Cb0ClBlNXARwGLwi9eTVGddnM5iNBvSJH6QwFJLZngdleBYnNp3lAP9Np/MupZ0n
TXLlBw5je6Gm5rd0gT5zn9vJeY+UQmhB/2anSjM4WsIYuMU+KhJ3TjzAYdCS5BQu
EbXWafK4grXQXl1xXD1LDTYHULL+WWS0Vak+5et4XlEUdDiLyEOAL+FHQoxBQmh0
My7+ulN3psv2iQSUUqgaRsuJFtA4iXQSBcZ2g3Czx2yIgcskUaA6zJtIJeOS0oY+
QEO5gIjM+QQvmCwJgh+xWZb1o4OGKu+Ec/uhpjRXr5sWFDYTi2N3UqfzaYM0GvHn
CjuvMJcaMQqOS03TO+hecsYJnZHRzBWcPWvuBmRMUigIGPLPg3g5GVywza+TpBNi
F9JdE1DYQ92t2YHMGEIzrCug6cJZN8CwLIFq7COVvqA49f5t2E044enJ8FpWF2Xp
RITQsuzTOPjcNLt++RZI0i8dM/WcSSYEwI3rMddC6OynBwMLSLrAGhXBSOUgF46K
12hJD3ksBiJmIofTXoEBQyXkfK9AsdebVkHojbhNmc6Lz7WEm2BXD5qdveocujgp
uzYAogYynV4VGAOEJpPouZ1/LsGAS4SE5NwkTyeWGwmzZKU/Sf79F4blEZR4fyeG
46s6FuYpYyXNJL/+gis0v9hOrAuUwiJCF40jSry8p8ssVBNtDO9ajyUziQEhhK4K
QlPHxP3ILtRdVHgp4tQYeVncLwJW9i2wJF2xgA5iZTDzdeCe3Y/9qo6jTE12bgfX
mXAHSbhvvn3RvOJ5UA2Kdo8cDdTxw7PnPj5xbDvPqb7SW9OFIHXYve9gMdQI7Qgg
KGotQaPLxA90JuaB9N9Ub37P+B9WXdEzQoK8P8gvs7vmtS5RDtWG2iaPDAESpNmH
Js/7IHlticxPoh87l0WZIrD500PikCiMKNMb0RZIywyIHqPGAEE22T2e6GeBkz2W
ts5yTgCChaRCQ7lw5KorEUVhqyeJs7E8PmJxgBYBEITKixAfFinczYuoNmTaw8XJ
cM321wuteqbQb9tuZpZwSh0yyOTHpjg6iPIP489cCcP1/9FjqI1jzbyKHLurA0pM
ZmkmB305AtOmI82HRCOMFAq23ODUZIZVnOUJ6EP2akQVJCjSBwvfJ5wCEpZfa76p
88Hzo28pUy3D7PHYPan3YQAlSqLLHaT4yTcg49gv/WCf27OroxDeWa/4UQjXXX+K
ZJVlDiNuYcEbXzLe1dWmQvd6GT4JXzWOLfESFIUiX4szmIYQyHccK8gwBsWWqFJ4
3JDW+pORzyK9T8o6mPCtcamibRrMTTGud2M2w6aOtSnJiRlpfztf5tmdeEGVTxJO
9PBzS9BTU48vKAh1VtaqRhM51EKsyoC8RPetSMfc4FV2JvuaeMBHIiXwvicPe2cf
jH/kQMyFs/aUX7roTLLPttNGcqymJDfwM/ssr0FLj1To48+IPSFU1muyLXVEXCNZ
lGSfRVHTlVh1UWZ/V74F587H9RqcZT3UI9iaYUWxzpmDM+7l2heD39OWDD5ojq8i
D6jcxpiUK2P5upE8v6o6Yyq6cK+m+rSj1G5282PWeP8ektvZ1wColsDgsIpc1W3a
IajAH97iI/hAqdPcDfO6/hdtib5d8JvpHXaz53E7K19kxgqrawbOCzhsEFmOZPr4
j9Ka2qPa1vBlpjdqfaOyrjjD/CC08qDYDEiyO4X2xSJJtxs+lgfD3orgBc8j/Pa1
6WCyNm2KHC3BoSbpVcvtiOh6NYNELENUkb1/7za/t+0Ho3LYocc8zRNoYrrHHS7z
YyIIC13W2RJUaKrPmsGxeBYNBEzCkQp59seVdAzFK5uNoxK9Zs1Mhjyqbadj4Wna
wCRqIXkNNpqV4XShMY5xSFHy00khW6pd92MGFxr65yvRVeILrJTQQnM7v+nThlhO
ILLvijOAFv+udSnwuxCUmT1yNTt5ixjSSlXvHWlZMNW7Cy9uIEDOjwd0gyUarVBc
Ld8E6dFTs6aSqCWXNzXvnUOlyWrBSHisuzSHwI8hf+GfGuJBQQ65zC5l5g7ETAsJ
CGqi1dnZaecevZKWf2bxnH6hCMernKqpPhtunh68NwT0/nD6eZHtBAPUBtWvo1Wh
DydRy48g+UUdyQ9jAtXgSkof5xmIjvx2dIQG9+E9/NoZtGiz/8jzkRN8pHPzm9nt
U8aNtq0ANioFWuKdUM2cIyWf3cn/8kFN1YEkv5qJaMwQ0n0zhCFtpA13I9qjouKS
U3d9UT5mg1QK79f0tIdmgO3XaJI2eovT41qxQ/xu9AglDxzLl3jZmkwDrALUlFYT
93yIkF8G3FlemmK5/pypAVLtEhUSMOnENfHiVF4bU+M3ELwQKK4/x8Xz4F7hKcxw
mU8HDKdiIOfvLjMTZt7Yhkg6xSzakEy5OSNpHV06mMhf4Dlo76WtoA4r3av1ii7+
7zeGnD2cBA10xDEnU25hN+bHxm8WK6649dTQpc5R9p+d2I/kv/p7f89XXxLmefkD
mpKa4qIIyXHYvi0wFvUGAkGkweYiwLqE/AjRB4gBt9XhsOPHJScRBrwlxg5Kc8Ne
ijkIX7/8rpooRDFB1wiYeopAQ9oFNGeazYE3BfAo/q0ZkW5+VdBU5AnLOFbEg1Ch
7wiq9N1sh7hWMCsgZsmbgj5GHE+k7eTShewUfNAB/uEoV9fYO+beibj3aCL2kcAF
jTxdAPFr/nD3O/8vgUqZ9QBu+TAz83zx8oSVI4WJELSH9l+WppxOFkZmo/Y3oXvg
oQyaLHi/DhF7pnbNHQRMHDENpmZxKN0ylebGelfMy9k8R21IJgf3/hxFNro0cDrY
lYeFlNDtXWOrfUpnhycA0zrhyCb5t3pS05I7RwJ/W5pqh+3wjFf+rwDy7wo7nxQn
VjORPouNaKme7n6OI0xWDitAEax2aAI4vDkLE3yit3J6jmdHgJVlTZgVKh5JUa4P
izZM0eqLIsLaWdfeh6quZ0Ww2sX3LL+qVND8puiRpc7lqqkRqJ4ey7ozgul5nOIl
lLTuDMcZu3KKNGPt++z1JMhN8VS4ZMdB0Yss5owptDeFwiQV5dWYCIu9nl3IXCeu
HQtTxCAE4Z3+8gFIGDWLzXpZIo5w/CE5ve2O4nmYeYvo/vF6PYOahYrLMbnk501v
dZy0VqYHneYiPr43jvxwjwa63s2THvrbODr/4Mo0T5cZpNcnnT10oqFBDYD1Rbkr
VLSxxAOdvQ6kieom3i5sf7gIQQA+Y8jnqUn25Gq/y34zwVGOg6c8nqddo2cpRBP5
wyNgSYo+4waIiDTblFq/bvmq54pu2OZB0wmpiBWDZjwzcv6vFyVs3RPxig9h4uOO
nDtZTskcZFsAuPNAkb+31SSsoj15G7s23Skh2UnqMRQsNnO29M+zmlYgoteANFu9
R4p81cJMYhNOdKyVmF40kLSag977kbRu069GtC0aLqdNTQU/kwrOWND+Qf/4dxjq
IeStZppSDSIYbIlhAiHTv6ArNfA35cWW1sJBd+YTeaJtFv/23GK0qEDXr4TqmQvG
MeslOGzUCPqavF5ugri7wMSlESlF68Y/HTm3V32e4/BptfBC90tBOTHadMwu23VI
xRyiPNLnmlBc4HLhMPDl9QgsIhmUI/r0KvxTFibYPXxtwujkYZ/Tg6wcJKuN7yQ2
gNWlr7XIsocOWTjZrFysJB1PsbnTrcH0WEh3Py/xDz57akKQqky3wZg5I+d36t6c
6a8yaUd8dEMkw5gdNgTyjGmrKK10zxZRzSDh8qlGf7IEleZTZY+Ox576atvfC+cw
rMh/2xBosf9rZR+HQ58cnmqlJ4MihEpim3qUCzS4u8MLfVQVHXlIwKUg310Op334
yazS+H+VRe5rzBrXYDGap8gpVzT5WPXPSAZyUxVJlblKZ2D0BEcdigLS/bkfgX1P
6uJSswRZl9SKlpvTgBmXWVRu5EeumSD72Gr0KbGAX7IQtm2SQXuarPZ8QVEsVOKh
x7E5y0Hotsm0JBXYlktEh7YVolGENyYgK+BS/Rs+EQlWA2CTGp2fcERAoJ8pDYNm
Xbm1mX8k6eM2Fn0M/h5JZ57avr7pWdxjbOEMDPU1343QjDA4FnQEMvInEXh8bDki
Iwgv1U9ntELrsB+4/KlYqjoTdU2hTv9hDPuv/Hf6TuTgfR4sdbtQ74uwvr4c7/RG
xlU27/JtTzIZ5q2gjwJSSTiP1HBvpkAfXGenQ03odq3pcg0RufX0x/fGxbbXAsbb
35HA42YrA1AGrkoNQW4jHA+NQrIO3sNGY64u5QMPJ9OJa0W2yf0i+zP19A5Ugkaq
3D1leU/CD+MDZuVLtO8R55TwhA5MI+feB//eRdm8bEpXRtXquMtDmAkc/Qh1zPvD
dgGiUrT3kPiqXIwhPcrQR9JFuZtfcrCK93dKSlvoaDJesfLz2Rt8+MLGWdje1KX4
EscfbjTEiGQyrezNBWp5kDux9che3Q4NS61OBlvVi8uLiliccpnZF42Px0qIKe8F
99Dc4RTzL+tJM8+06BvPabS1x2sQeC1zGGrj4fxnGouzL5ckEsnqvXD4LV1Ocy2D
7H0jw56xV6jEHiJRnfmDaRrz6Y/xOo0bNmj4ITar0fKD4zg3aj8y6ypaby3KUaNY
gHux8TNQ444kGYm6vCmMcaNGO+WQYmMczmSvSsJMCdCJ1F3R1t9LAM4/l0ItTd3J
LgVDtVXPBLq0dZbkBjLGD2aCjsYfQS4MSPUhkQms4RArlOBsFiUkkrNPd6tE03Jx
jM2amBlFLQsCbT0jxudvF4e2cDbSOziUY70Qw5ajgBw2W+STwh2z0n/WgFXlLiCN
Il65Z/blkhlA13uCc4fruliO/dAnfGSxNwFnhNWejt42UzI0HHGBt09l/U/RWxHa
EWcm6b9jHrSWkNmjntb3L11TBwQiwzZFapT29FkPLJX8IS2ca+h52c41FthedKKS
syZE2GzVKq8sPGucjbXlb8gA5rastLaEu7UaUnjNHkH1pMaALKe939ynxJkdrAat
pf1xIu2b9F1td4LL2+8e/W/GOHC/QnqE/oYORofqpPLMRpn0pm2UEaytsp5jSLAU
56nshB4JTpTk1FhGTpRPiEJvA480pcHhkGf6mimaD0LlsvsNkvXJ1SdaCDsqkj1k
e1AShwgFEsu5HXumxSWh5T3m9ZfL0DBG4WOfyhSnIKo+YxxfahO8dmfwPdl5PhHE
FP7ghFgQGgtg0auU3qH5JDQ4H3oNcx+EJqQjFtql/WyJJXU3hLwfHmHjpkB45lgU
FdqCvyB3Q8fc9NL1Tb0TCMbVtVnbOquJ+W6M+X/u6roFeA7IoOqZyWgX8i+MC7lG
ugyhl4+T2tFuxQ5+IAbVbscdABFFPziHXRjaq/cjQdaYBCgteI4GGgr3L8FOAqTE
4uaEvnZJqEkuzrYncI/vm3N1fF1/RGEm4t8ppqNldjVsKizSyHVRIUFPkaaZJelG
k5J3dfTraA+K5P0YFwm6UoqUSEwLj0xTMW4CUOR8iSQTbq7CIi9zBeGNU2hrwgnU
X2fXj5pSP1qtYmascVuzvZd7hO45wN7tuD449ykvFcmX+9zSc2R9yf81X9e/Pzfd
Ek7btH8Ce+qRdFM3NPQaH7YAcw/MYidGqjVmH+UrBKrcGyafm1w463lo7hYCKEN+
iaUn+6dMakVoKXipSd40zyzCAjJLlMnIWqwujKu+zeEtMN/kiD9jrZbbr1+yJhMb
QrOQ2+QIPcP63y+72o9U9U9gckYk0oYUJCMebkQ5sP3PHATuZHkPPXuXV523H+FL
1GUWhdXsGwFgDe2D0W80IxYNVDNmK2sCClpMO6C8kyK3y7Sz4mNZKADunldQFv/C
ENaaZW6Fmvj8vDhDv6jIWKEL0IYEAON7r+7INp1gUxCztKLjlNNz2Av0fDVciPO0
TWCYK1WugtKP5IyNFLeKKkmMV/KqBEQ+Leq/6qi+wDUB2myfQhjvTUoLkuYkRSfG
ruDJh1IN69I9QpE+IL94uoC5L4QkixdY/g7VTwcEsITeY3trHkZQeA3oRqCWum9r
wswzZYrsnPZRpojsbYi+Llg5fhdGJRmST+e6dzrMLrKKKRjrtawlUTXDBCwtRNWn
pBo+1rT2wHjkTvWR/4CMcVHbP/IWwhfcaBe7KdV2BhSeEkqNOi0fF0I+Bkk0LbRC
eIipHU9CtZw9VZHio3cTfv+5qVRWEioRgMwpPV2xtXNTxWS7RT8jgsmzV0TKIDnQ
/z7vKJCtXr7zN0GnUnIe56OV9G29x054qoYxooG16l9RGE95DghMtskwpJzu9oXD
HM9TByJynMYug06koQNUmkBL0xdi3tKvLpAWac8fxwqdLbFiGljziiuvOQMfTuNA
lKwrZQj90DnWnxDngEUB0/tTAOXA3lSPVmWsz1exSE6YxLy2r9iY47cHd57sE6Oq
3db+A76jV/sYKP7boGZI8okZnR3ABVsKu5sw9nGQfCZddWhdpf4MYfAXoRphdr3g
mS7x2yNUsL0z3PZm6IGZIXvXSIgIkHQU1EIqBcnvavFY5XmGF5hvTtMtY+q2OW0Z
GLtE9160nq3wchCA6GknnYRyg6lhyXXsS36yrI/pTkN7tonMEZatyXBZY1A0Zwiz
8px8bbPWV0hzrGT0j04C+D6pcLmIWDHCOxPCBsOi9d6PK7afEpu+/Uy2cILkRIwu
Dc3DCxtZVUsMgFWbkNLpCmtDcFilG7CBBUMQnLAL9JhwT7TuZehFpd8X9OsjXf4r
Gej9GUXTfBpv6lg9Gce2UTPg/5oBEuqf7+fnKLGCw7sE9BgT7NKK1wFbQg3fDWdp
7uhUSCd63I1ws4Qy/37lZbeodFmWotMBr8kAarqHvO5FJQr/Lv1yrCevKkx7p55m
a1x7YzenLxP6WQqYG/U/gc1oTtjvI568NHGcI3j1JqZ+Qh34/N8HdnHACeHbMHl7
okYp0XJSJE3Ni+OuE9BIw7v0BufMl13xqtsiR9+sTY5eq6uAULCgZxik4P6GjWwJ
bX5cwTsv68wp2qJN2xRQztta/PPfdGcLap0pls/3WCIxfpypbk3sfCylrJedP9LZ
kzMGU5XtbqmdegZYwSC5dASVptT/FdaaOFSfviclYYl8rIV0N7mf6ZLjbpJxy6/b
3P+6zL/NEmxrJX3a4YaKwOzxLC3hFJ/jW9i3Q3QUbMI1YNDsp8hr+yL82uQi9UVn
pQpsryifM5BcSrDimkBfUUEPjRHTJzTRmdboBnx3DZncWnGGhHg5GBA/3Z/XbXNb
opJDwUr12he1Vn0B9WydGLESWk/MxMrH+JCk9DxKrgZBjUE1eujSCHxHDMg6yRN6
Unv9Um/+sbEgGozTDHSukBp50BWN2kXpL2Gwc/iHog4XAssJwTiz9nAd1zTqluz8
NmGjkxQHLwObiU6OYa2Eg5AjMnWj1ZjyVgTrRmVwrNYywzpb+UFk3RZAU/c3OaTJ
Q92oe0XJZVYFLubbCd9ZWMD26LkUueP/gO/B+FJYdYcL25kYx5Z+31PpPT5FZJKb
5a2WwLj6ynhcAeQ8i2ra5eAIbFZeiaSZI2f13nBtuY6ctMH+JxeouLHtL82V3Pa4
iczsM8y6KPIMeN1UHYZbFloYYJqSMIp2LcPELCbtNpTe2mnPnys/LY0I0Iw/+wvb
KqzninjhVYFLsFWlJDArAZmEeH3qGSZkTsvXi0oS3CHmtk8etd+lXUEX0+3iVRs7
I7BLPbfONUFIQ0JssaH7R2VUJ81K+pgv0QZHwMOaT590Z/PtGmw27q7kcAybwr7O
OrX1tPM1diOzyWdZOKoR9c31oMCafgZdP4pBYZ4YOLbFwRmuh9XSYnMtg8oTNFFu
lyChCHCa62itV22U5ooXbO5bfHhRdh3J45ckxJlcXm8EEMPDpRe8+uEvQf91pj7X
RXwkO8MpOerTRO0u0RSXjtRjx10BHiDk07HEyJvyO76jDWJ4Iwn+F2k5S706Q+cG
3KhjJ57LeVJyWbqtCUVttCD4T/uCKUEP6EMiYQG6PIv9LPZgosuhqPXIJBEC0rz/
uKrn0t3UUWQVheOsyqhSPiuAVEHlLlSmV29JncMz464skF5HOS66BCmkBngXceZW
aDxeE0DJwz5eR9nBolVN7SYDPEH6fywkHuDPEaDSobE2Y0dbY+dMAyd0RZol69cj
/30Yl/m5Sbaikpt9uinP52bQl0FBq/0sc1tLLo9wZ55IfKtNssWHg3VZxktHiulU
nogFm5/vT7n8P55vTmlkRlNwd55H1Z+thf3+p5NNBvhy5EHoAUnGDw91HmZgI/64
yE+dox/lBD4SptUcHmgoMbnnMQnxviW3EBPMqvCUONL9EfMU2PqCm1Nrtz6jwSSL
wZzFOBLioicdLWPS+c3+KnGXJ53MI0VB17/aUXrxn8Xi1nDOtrRUWxqMfx9sC98u
FmcNjZhFQGRWekzrnulwv5koQKGgbuXhvQlMUg4Ry2QL1N+hZ/rZ4B1e19oUhWgB
vrUOT5PIZZjfvhQUZ+zcNSobyMcjXqxW4nOsqnK2wX7/WiAHXcazJzFejSyx0iNY
/oBJhbpdKEQFmqdXkF7nhsP/2w1uJD9liEAx/j2dHTVWiUEEB9HYfohtnvYQfjFN
pwZ/v17dc1Iv6tcWW/2cL9EpKPmjAS3Dp9H6xazdxZkerUEL2akMrXtWReTMkHdd
7ljIXhYkJRkuJRabLoau8Y12YxpxhIzEW9r0fJMhVpfiqeDkKzP6Z+y4hIZIBeYr
1zbsfLspVctj4eeyZ3z6BpF/uR76G/ysnbnNGf1IQ6ZHNFyLwgfsNo4IHUjzNmn2
Tl+MNNHQy5mWlQLkbp+87k2IzzfvhXYxj31xw6LKBa2MBq3xSyvZB1LrHT7UgUg4
Dx9r34q/xGDHVCYZEhnaI8BshdR2Q9D9qGqChMSdz+Zk7PijsowZE7dSsyZQ3sl0
oDosdH9jMhlTdwpwzYV5vIg4CKL6GN/tJHpeH+6j4jFagdVTs71L2XdlsFWwEmwi
0dc1RzBt/0YvCW2Oka/6Cvqu87kTxTY7k1EMHoM22PTluec1iA4X7rLAbs//sj0K
+KS/q3fBm8kbFJx8CCza+iecifXDh8w/uNpnUYOX5UmlIqbmWFfPo+qO02KWW9ve
DwU1xVRlPMmKsjgHsP0JrETKesESKq5VCRYZxk849zDVjHv1lIkPP4ZO7PVNd769
hyIQz66q7TeFREDb0ol0hK6hZtyOJBRtJvN1IoKBaz4sy1/Neb3JZahc5b9uXElE
6+97SET6SK/e3MbQyqXigcLXvM+6pLU2qOfvvwb5TSHv7g0q1kxff3KGo8xJ9g5B
laHKYBEHXi8VRjpRFZ/SV8LxUADQfVBwDWGsmc0ABxaIP1jXIfiDwr3hipEb/Tj7
wKT2NZWkITAyadIm/LIu2yzWei/NGgi4QEDUlcpMuvPq2z4SCM5AvhLE/Ku7SCqM
PXhBd8C+BS9KuSbSL4TRHX9CZ0OoXqeD8iIMSE2vQ8ZZ9r5FU+oVvQEIEioZWAwH
5ZkdRBjPg6w73dQtJYiBVk8o4m9Ne6VwzThmnfXPXn7OxITK0QtTPWLCMtT+Maxb
MPIRPP6qNlm0GYXzuVeewn/4WR4KfoDWOozdV+YDwjnK2LqLMVsCemDYaNkSE8Kv
I66AlNpuXLg/4nQUzWeTVFSrrubwkwe0L/yLXvo4U1Da9H7X/mPCp7I5xFawNGZY
07GxCEXRGM1A3eIJIjDfD62emvli6Xhbtxy1mO+j92C5NU0hScCak5Y5lrCi+3Bf
s0PPtUfeocoF7dM06Gg2Uk0bzScbf8HVuUAjMlxWEwOymFo1Ne7ib1Zg8l+BKtyS
LH3fAUMqbfXuxac0H59HT5eJMOXmc7K8lRUuBIhD4QxmRNhPqYkC3m2MTrppFs7h
4R3/Iq2My7yRGFeRGJH7Dwd3Nmq8iGJJ5W22En80lqQbrqfDw9HYtE7m5oYXXo3k
H0te7FmiBdeJFnUJvOmVPKGAWk14dXjUk35x2RvID7NqTbgq6mJKP7YJL6x4AxoO
x4vQLoe1mlXZKCNXwDPC93SfKu86VBRgnfW3R7EOxTi1/YVhh89x4mPRdnRkqQEn
d3PvPMezXDzpl/0jROpOmD4kPuK0KqM56iJ5gTJy+A1j1gt9fOUpTsz0jmIJM/YO
IeH0N2FrE2oQ21bfeyC8m9TQ+lRAQUyCw02QqqU4WPP53aFl+gnarJpJuoGYlyU0
ZI+MamJUa1dkBWujxYbtLhBajh4SZwIHTu9skeQsGut8IMIN4FnI3PsROJ+FVT71
1Vca/2FcK/QEvwMJzru+RMSH6oOh8NM47p6LAUQGgsZygVMQTB4bH7Rq7HSoBeX0
bkjauWI3qc7Z1X7pLgpOXdLwuBLSdNwpDm120FmafeDiCOJE4abZvh5xYh1G/lVL
TSoIAp9te9PP9fk5oCJu+yltDeJvzFn/iX4NMXzVOT+9YT0py64ZQanBW/ywni6L
oqAUCCMp8Am0g4YLt0TJnn4jQGQ4VUzWqX97ngIt8E4MWaXVvCKJ2WKmn2Pr2maV
hIEpfttab5L2iQErRq35u8tOeGfnQpmm45VLTMTnxj7q7DaatxZ+3elzb/t9XaSn
leli47RrK9z1ZgCabLngy2gv6POVA4dd3u0WjlVoeOIgjalNQf0jE9ibOeTWk58U
3N3dqdukVkXQwc3S9jZwdBaUSoOlBGBejGN6TMkrSgOtBvjqaSiocj+nN4p9+im/
XAxHhHiCHc+9f6ZYXJNSVbHhmFBYWsFm3+nT+PLjpayqc5o00nizHqvWyoy7uT43
mFeoGZWQARu8KtT7ZqCXJ3NXik/qia3oIFs1ebPVMCNTojVzfAtj3fDwCpJD8CWy
QcSmOorVbNR9SC8wiOFzduoKndj4+hWQpBwRHh+k1eYX/hdauNG3Q/uMiY1TTXdA
FvTD7CKRgCn0GibtZ2jaOEC0KRQV/Ty4AYrUliCiT4OXRcwDo7uxYWmTUTFBarHP
wHHDXNYDprXa5JYDzcdMNFqEWc5GIuCielZVaXRo84BFWNPbyut98G8zWRcmnVzQ
vMNFcA0YdNncqYevP5ctb0/0M6ebV/JkqnxYPgALEZFEIczZjFKqdbHyehaFJLyr
RQ6sUaVhCVsWxeXAQe6bngwqoCFYWtUbeArFNt3qIhRB8cFjABUa5Vv0yj/Qo6UD
IgWLD3w5DwzcGqgXJKDmWAYnH+SOj1+9trMNFX8UnxO29S9N/xMreDzvYtrIVECv
Kh0NgW23BGjJhCrp3hzcjpd10HNGnI2kvWKyvRmYZazVzlLuD3pCbGMuonsF4Uj4
yZSdI0rbde385C0D4JKzAPKPE4zEs+Qk/CJIGePr2/2Ige/qrl9mn29UrzY2Cc0U
izafn+qmraOWz3cqdiHLRjYdA9iIhBbXSkBGe6MtVacLBgpqYd6fJN/WAlze0eta
xRkwbWI6zu2udZQLhaIIkHFcX7IRjwImnGnefbwrd3Vo8R0yu5Ot/f/o3m9bdOec
e1S/1tRaqyq8GgTcnoa/9bcsHds39J/UeYiV+of2EwW4hwGpP6EQQ4lfTlNBpsj/
YfGWhEODhk0Z9OmL5YAOKAobIBuj6oiO0RURbDYc7N9wNM7bBpnIbGcl4KpkOH6j
pX6+swmfAwSckskbmdWVaLQr+9IHNwGmcKjLl4Np0cmOVviwpS7Mq4bkMzI8XZV7
CsjuGg270wZdHD4TyZnKsgK3ITJpR9c2ICBHHbTWtWAut4NYAO/WDLm+zVMSk722
sDwknCek3TwqQInxJ903l0Hl45LuyIAel/cMmRreawHwaw8FmzUlOoeH0zCnqo/u
daVRZwXtukWtY+mLHSXqQ3kIIJZmnKyCXj7dymaAz+qHoJpj61oPsDwhJe2kLz9y
bn2u50JMX2gi/wTfF+7LjAeSjddiBDVP7YafOQOSBeR4YSHmtcIKq62IKSL7DA5c
JRbWoJs/P8BLFzQNQ2lMqLrO2T20egryQZVbFRbqMndsxDHzm9mblE5aVRCD7T/4
PAhV2k33iA/JNcEGmECVNniAE44yxIZu8S1oQhhaPyjIwKeyNeS9saUxHm2AhR1N
vUzQkHRqsF+jeO4/H4PU5Ged4jwW63PRY9ARLho1rMZ/uyWvbu8c9zDw3tbIvllx
mrwBKnASDgii8yN4/T7XayaL3uVewMFOTmMgM54zMK3zgob8/LZsL7Pdr2QZ9lZJ
bJhGiN26Ch751Rs5OeF+kTHyfYnV+VUfRN98dD0AURJj+zEdBiu+xuFij1RugyBK
6ocDEWbhV4I84ujgsDUPaGs4NjyIO+WPF1gKuPAW9Jeo/xiMc/gaBzz75SzsiM9A
Qvkqv8Cowhj6M0nEUIalGMgysx/0DV22U1rgC2MQYibzwSw2IWJ1JKUzkwS8num6
aKhLEhr7rvEvl1iUPtsKrWTKDXA8/RKMV6IF3yAgg7D7B6C5rlEsUta+qAPtBgLm
2wuJXbd4UfunsluKIn5qCxC3HVA6GuwHx/P4PPmMjWzJ8YlXUyzvhh8AaaXmRpIr
ktDy+0p/UMj/XqYiIIyrf3qsPDwrs8i44Z0cTLnmCWmUQBMoBFyI4saec6vo1gHp
x+5Q88LavYUopJaQWmDxLIbIaeItUrIHrM1CHX/jKNBblLJ74ojv1yND7IvHjb+q
mGKe2ITlyBp7dSem22zmQ/0At/eEDTDxEU8rcJhDcYC/w3qQobD6CKgA+wXl69Ra
zutTShBbiAjxooYlwcTm2RTcEOpXYeZxTeQzWFPZog52BzArF3e/ef0TrQXeXPwc
0H6JRnpAyCeUPWdBWnM4suIVYadx1C/H3GE5YFIFnxCKi7CyGqP6twoDkp2zExXf
RBLPUVOk3k4HXxWjkQ6TRjHUwD1gVw0goQhMNPn/822+He/4X7JTO56v1If34VVw
76jqPKIFvLMzka7fTuCIegzn61Cw4sEjrdQFgzEMNxV6Ykwdo3l/WV4eKeByrpgG
qg9N/Yt/5dc6EZDN3VG8DFqo59RlFg3S5+mE8KYx+L8NeCnd6zzIyOGDnSk2S2EV
NSRbezb9rOCQxHy7Zgom4/fDPBJ7WT+g9WvpJCA50Od3e+xEPPzaHJDfEJcHT9AX
XFJJElUscgqBZAQlzbcE8CLi7LFT9TC9LPa89DdoQ6HFGRSuqwUDVW1sKIdAEPAw
qv/L6dq7xKq0ZrGrrRVo/RjfjsW1D0pG8hkfrM91aubrwgn9vvKhFZpfgfoSrusJ
1azoxNjQGFX6fZ9pLH/Md4tdQkeuSlqM0xLAtrLlEtsYc0xXE+eDyEgLDahxKhSb
0xBCQldFstn38MMo5cS6nY0vx4sZIaUkl0XRtFAb2sCyTF3DEYtUmeEttVyRbbYl
VOOTQD/gJjqKlHmTBmPM6dOadw6HT3HvUHNB42H1Vv6C7Qlnod8n68EZLcnNalof
mzmbDvFHn1yMuGJofGkQS66E4aqddmxeakyLL0/pJnj4wMi5NsMDpnX6P9wgwbHF
3MXd7fuz9bYKOKPxw6ZQxaY7HoNUP3YZeion6TN3xtf0ktKtcMbqHlk4+5kYrEww
0HUdl9JFG9xeowpYDPd4lDsbo+O03jc+U1zcnbP9iDG4hLtjGWX8rSSS56c4RDw9
b5UJpPXilmmWY/i1c5aYKFKrAbiQHPRkVS0n0dOx2fGo+UDbEFJ+8IQWzg9rLbGU
5aYYBca/lLlafPq/7YHUn0oZtCiJs0sGMsAkgvgUxoDeUyCGMKqYdyyFKYBE3woX
0xfRGYEzYWolZFbcYWnwjyVsG9rgkvv90sE6s1ak0NdPt7l8Pt6rK2Wk9Fs/w+eN
wuVGJQgXD6lPDndq7REaSyRLgmK7zzWhCk2xj/NpZ8Q9adrtW4z4owigv07cW/y4
HLdY8WMjKDO+tUSW04BszOUe630NJot/1S2o0HNruslAx17ZV3zemNnGeImePGi5
uewDnvULNFhovvfdv1GgvhI2XDXW7wRDfDtaNGicP8JsFfM4gFMvkRAexA22qvS3
AoV0WN9UiMRU3vLI1OoZ0TnN0SvgTlKW32qvz3hXY/QHWJZj1uTpJtkKkGk/VKpM
K7DJlnSfR5X6bzTwxP3ZN2EpPvHjTp29yESVFpe9HYal95C+HsGGWiiNZOzR/TwZ
yYPqF2tU0W+1h2mQwBmeHCW5p8hL18IPt9LDpdxVLYaK2N4OmHwcHg0BenHVAT6T
NFMWqtX9nwSmLSPwgbBLvkj/XV90GrJGidoUGeDNgiAdG+1ldvKivGGH4sroGiZD
/6PB1ll4W+vn+mL6pvYRojZKNMQ64IOEeh2gkYgdDQMX17kwlpKS/J8gLeST2qiz
PowN2HiUZ2YKdGMRZwREUM6aIaUg7ha0V4lXO98cPTxiNFiUAs3o626I/sNRG4Vs
P3UGxLKu3449D+7SHiFsav/zauIDED3SmqgPwVAz2zyPq9s9S9RvduxGh49HhPON
ziMreHOhxZ5MuFpG8oAg6MCBWPRS1ayoQGojSgBu81Bc0zjV8NvRcDVMqhqBi3FD
gM726HgLSDiq2A6zJUD5kRMRK5Ls/OS0CrRDjvJ14wTE21NQVFQk+LusdKcXagsg
RdrYhr7L0jdhWPFdJ95/Fv4SNe4cY2e86RPTwX1Sy2MuKkinv0Lw9afEz/oGTb0x
97P/h6h+ue0V26rBTgiPzaKwONiL6wR1QDgGIAE0C/bsULdQfilJgJdtCNaFIPs7
S9YK4zvzv/27/snr/YiNopl2YUMvs0eSOBOpz/kXMQd48i1q9qFNvmNoc8BXHgTo
N9G/ywZR+WGKuS/CCJeeUKThkXDdIkYBSALhaOOVtRDSKifswIM7PsrLbAG7kbCE
UPCqjsfHclFB5dM/tedU7OyBz7w8YjVYG1pH05qDDoQiiDAHVr8Zu5FKkktfQfGd
bvIb/1IAaM1jsU0+6s2VKMIikxSEjcL9cZBXzoe0CLACG1l0P8h7LXRyjOXRuo6J
Oem/EWJIOHkx6Pnnt3e5LpUwnNmId+d7uRC34Bp5yuhQEm90LQECKD48Sae1iFrb
W6t4VMC03H4LdSXZCNCCjnmJSBeBp5xiopSGWK5ctesEwaL/bnTwkzbwi/xOWhRY
xNYY8C+ok2WiOJTRg9a9t4pv73Nv3KekAOJaLvMUhvJfM3kH3zg0FjP5e/WjFS0e
XNf8ijaeuFh1q+3m8FMMZXyNAki1GgDCSbyoA49PPnJtsNbWSYhr8O/3Tv+vUC8p
HP4oApSKqMa+oDUe96dRF6J1hDWLRcONpFve9+kRh/1v4RyrvNpcUnMHK5yl01Q4
ncmQ3WxenDMYvb5Ix7luwJhNLLFsYK+KyebQirPlBrkV4xCLJhVj16mAlW49aRj4
dhCD2TGRiLKQcLx2XFNEKduL1jgNH4bCBUhQvvbiDRCyxv8rq0bXG2u8qgrUtTeQ
YqQBGKiUnEeZVnnsHoz2leUImWLCx7LqvweGRnuYDp6ZFZZMZfcFG2c2h7yy+ejD
+b+dxnVVyZioRwu1uezhP57W1nHvbyUZUZopLbhZ4tRFxdXqTQR1s+l2aBvS1yOO
v294tCQ48kRo7Sxk39yh1W+8IpZ8OcjK0da6xiaAxMFccYw/acnKRmKCkmGcAgLp
nxtc0EQNstV0VcWW4VHEUvlsDiJrbT2so9k0vkVpRbWAWXR0RbzFDTUpSBejV6mp
NWffSMHDMqF85zph1rR/NyvvL4qGDvBn4UYV2kk87dgZRzK5JSS0ebaN0GS9LMkW
p3TUY7VxFExgcy0EEvz6gT/hoHVproSWlkBtWwkoV8YNBXntA7bEKb75Ik02k09Y
tQLvbbCzu6LPkKegdQ+1oE2YqvhFv918/sJ9JBeUyw1lYrNZjevI4ypyXOwZDN4D
3If2Ia8R7QMR5VzotJkkQHP7XdKXrGqCY8nWg7XxBdKxLYVLcCx7pAG1MGFcoReN
GNyegxaA4NuKWW8mO7tf0iY/JkHLoud6h9tcOemwOn6Z9tLx90FFzmKHZpHgHX/N
8tYiFLyrQhNULz3QX+MteL5fkrQ/HE8FegqU7hZpb10S4kU+QAl+9hZS7HJO9upu
OMnnx4bdWcQc3GBxYgwnDhiX1vlMoxXduswpwRgO6X0tzx2jQqrIcXgesrMMpAU0
zDPVHTk1Mu83OxVVQWIuhzdckj5yuzC3KLVHxA5Ndyrp0ulqURotbpWwLZcfCf3i
0AhtmHo1iesCj3YaeRoz9G7In5v4qPVJkWKGHjvvMvaaTWYxTIoY0/ILMNLgLhAK
PBj9SGbCboJs8hDdUSFHp1P5adtp01xGpvMYjN9Py17wbNP8QxZmZOFaflafMwSc
wiNFK+nG0oB/gV6MTXH3bU/XODwFthFlHqf4Q6Wa3i6L2tkkabvs2rmammbC1Z9o
USI/0g6hZyRKpSUbmXQ1y8Mg3qQIUeniO2pzNn9+Ykc59D/SZDL8T1szIzZZj1Le
1PiZlpnvFKtgQ+1L+bUnL8LTzxqLYHHk+jKFL2HzdKp8jFRsQEsK+1sjz5APtp0g
c3Brx2baZG5zWfSIVrFKi461K7u5VXIrcNDQUgtMTnRX7lZgzr8BnCOo05UagTX2
6Nb69AGzBSHPNh0sgb5/ZWVOx9moCfSZ+UQl2K/TUyk9jvg1uhV0hacC+fO5OkHr
2cL09fckA7PfjW5zIDN3U+Fw2hmqMP5Ws1o+9U6OSnlvkUV9HwdgwWJ7psw/u46J
1gM5F4eP/V8eHSp0DFdhod/i1mf2WAgcKDBylawxwkFLce+0eDBwJSSU9w7K8PMi
ncTyaZtolrcGNmXjXfk242x3PO0lujb70EpGCNVS5C0KRIoqSd4peZveF2A1+vr2
u9GT7ZOvnVpmES3g/pZ0YNmgzC9/wQyCDVoA8ow9tuIhGWS47ZGcecoFMl65ctIt
NRY7OwRqV/gxk4wwXh0faFxbM+ujvz8A3aRBuX5NZMbUa4o0F+NLMjUWS1NS3Fxr
FWhFJgXOp6fN/Hkb7EutugSz+Ojxjw1BDKzhHb/MnJiD3m3mt/FPvc0Q8LbVZuBj
TAcUq66BKwCnL/gHHqUaKvWKI4FTzm96qQdWM4wl4+8mG+aFdw+tZwX+7xArDGEv
5wbUE2EcJaRrMW3/TBgGmi5ZAHhE04hc4xDYNGN9un8effIsohZVsN4XAhsAaTim
s4d2xLMBVGYBYeaghPLp1R5FDzQ52LBNmiQ2bEFhVtwPW0lKc+ds+uyk4Q014rPF
RRdfTN0bs04Xd1Pp2thGWV26d/NXqBCY4RvOWh44B/jXB4PnwB/o8x9pm+sXGBPu
REbHbpB98bO0sgCIRJ9nh7j3N08J2Lsy44SRwyO18sWpZGFmto3kd8/dR4Cividm
fX6CwkftUMvTxyTduH91WUborPlVs861S/mOUIWMt5d39mdrG2/zsjaEpJmNtAVb
5XqdF3yHW2WQAopboTybn8CYBnozKXcCbXuSEMLLbcquLJmF9SdDguOM42BQdl9f
cvtKys94cNPSe+uqx33pwb/LGJ9vp79WDhE3nGuXspEeDt9hTph1iwosTG3C4DsO
KxRVyWv4YP3R19qnjKLMxscSq/pHAhcVQrBb6IHdzDqm4xFUEjG6D6/+e7LXYWmF
ijv4HxRxVQsypIANwkqU+HEhFkfwV/HocPQpCt0swUoNpPJ6piymtWFVjE1WFORC
zDVAMUD/XTrS2XAnNLkHRoF+hZ+S4fkkzgJgiX3dHj4I3vdIRuljWtodP0LR6QQe
keScMMkzf5pHiB5IaZSEgZIzusCAbTDRz9EBT5eOpylJ7rA6M5wvlmQhvuDn6sVb
1+zxetoknBosXWBZkPGzVy4EgJEBOpShTAqPuxcx21Wjxngp7pXXpYyHexHEcfg0
k9dsQXyHmIzaCoWw3dSUGnnHvjaD1NapzQSgw52VACotQUK/P/LDQjB42KGr1WcI
8g85XvkU5SfEorXUNprwupjBw5HsHpEwuq/VTxYsEzSIRmSzbbQ7Bs2jVHBOmZns
juF2DumeaU7inugB6D/TYbDdfa9H5lupORGd8pbnHTFMGakovegHY+hilUGTRpzf
fgDZHQYdgfb4BypxYTk01aXBYR+8wPLSQiz/ILzH2CAoBT4igJkCzgQxnrGpfG8h
jB61+vReTUbPV8mth3O99jUlQZw6+qtVN07Cvb7lktd/NizNWV7WCFrU6e/zr+Jk
4KhtOeshiJ3+PQlYyX0ewxwuh/A1CeR6xbzFfzr92P1LtvVffLYnCUt9CVizNTi0
WEO68uburtTQBxd8vboi/aVXLvDgJkGxa/mw2Gmqxn5aZLWd3TL2t9shfBcZyBNf
oEPTyh/6idsxgMQmRXEUJ9DF7hip++XFez2uSWDMPJ31dFuzlRimYoxFR+wHtwb6
ReNYZKRAaTm+YOZOvwa1Td0stfxR5+069GmV8vy0ww8B8n0KHCKR7Hg4D5VcsHne
lrDx9FbPhAAt+wcsmx7+BdCvlRabY2Hqa6pAjeM45DpkCko160rvDNvUnNklRJW+
lzM5KKDK5BF6kBmW3oYVqY+UzhjZFQLcpgb9s7kV8BaVswIsTE7yzGkuxVUTAawJ
I6UauBQd5CaSxnWeJZRkxxQO7rhNQrNTVuOsPE1ONqpeIeU8xr8U2DpBABSR0SA/
R7oi/NDX/aiipGhPEC4l7oclzZ/mAaAAK41awOx3MVE7VTeci1m5cAK4MWCt4YQy
e0T6qV6EpDYmifcUeYbcpW6dbd+QQftqkY2luDAGyJP498/USMu9Pfddq1eRRTkN
FYNO6JrQOZOCRU6jjJs7iA7gyjNSVEEbrKQicJ2NQKCdMcikaMxU76SuKJ3QZuwO
YQzsoHhGeJbaQpb6FqWzhtp2vSpl9LHUr5ME3UrX/skZ4gQ4f8aviR7WsKGou20N
vuuCjJWQ1cV/FameAgivUuJzpCL0Rahz5zqnAQhu4C+35p3Kh4/q/DXc5i+1zSOD
Ih17/rXLkSPZaPtjCxMs1YZZRwPdfsUksBXdeOX6m+ToNqX09WfyZDcLO6xogO+d
UbrDmz326rwCdA5MyL+dcu5db57sD+RG0vArz2euivgyrSnsHTJvqZUXvI0ddxCu
hKR/GBzpvfmdV5FPVy9LrBJpggmZFq/TBnJ445yp3pwS0QGR2n0nryfDCkfN5nkP
LuBRB2Jb+DWTGGR/VfZYZTZyxdrROE92ySw6qYQnuL7sVnGzA3C3pPDQ411PyzxX
GLBK79cQYgykzHrUEZCHWunUhUdtEFwxR1U9k9xZIbHQOZsRo+j/uvMsuq5qm3wk
pRD/8IJPOHB/YhSf21KZW763bmNLfKGIJKvpRrSIzm0LewHYAcuTOcY0YxeAot46
F7x5Gr1ePRTebznTn8f1OqDGQm9c/iO1gORbE02E+SQwoYlNUjt7R3o9liouZAuR
1oxLt3RrIbqDVXCmkXoQ7FmMncs+c5GFCiu2SiyYBpGmhWQN67cV3ZX9O8xYwhJL
BQ9qNJWOTEAS2qaCLBOTmQSnuygWqEHDfWVONruth8iwx9/nZbrqPOEuy8Q/+cOD
BbVDxPipPNwBV1kxESpX2NPo4gCkb+sNdSNgP2Xb/q8TJdgXXE+yNmTawIEHIHih
IkHxZALemlkusrvKayYqPTp6C+BZ2vHMfDmLwDUwyDB4EFzQoIyo3CeYpnWzGO7H
CmbiKvxtl6G/1awxrPuWu1IFW5kwtbO5UTX0SEcnmncharqNw4URpAiFAnOSUJpS
9kabtpLT/3JjAYWxwbuIAqUXRG0kjEeAWGE0TKQbwo+znW1hsES7+TGdEZEE4nVe
iqo7iIZSbpBypXDn49NLHEbn/Q9Q/LzT1k/Qpd1rflEqpytWykVscZM4qMtfDi/X
cUo6BzLoTMURJjcp60JAatgxAcEK19JAQEjQppyUCUe9xkoEz5sn2629Us+snvT2
uRzLSVnGaURmiIX7ytklvp144y+D8B/i9jk7IgCV7xh80/rfO74Dqb/lw45K1GPx
ixD16+U+kS606qvJfvAvdOtJxKvXIpNa0KbjWE3s8ZGirph7dxG/xtIkqWjyV7wq
28CHwf/wO+/vLlG8Hqpd2Xb2TseX6qjfjsO/7izYkWOQmUo1iHWrkosl6SCyp7xK
N7Jxks7SXBsjGYsRWX3Gra9HhgNYeFL3yOV+zSRt1c/Owszg51ekuZARAn0otc4e
ipqDLSIXLo8FkmiwtpaM+qwXyMACI4dMN4A+9hoEuLCoeaTfBUEbarFqc6tXOcyG
VQxqpimmD3aoj5nxtQ6HK2l8CInz785cbo6mki+EnMYViNOHRKwLAfywMgTCW8UX
tb4cfk0OnD1a4g9auflQGNJE+ej0AHNwVYiOmzxBzOx06nEDh7y47lGDv5SfCQSS
8dil99cUBr76ZxVPNpMnBJF9qgeF6eBF2u/E0xpkDkIKgnLTGRaIzvgAytcLUSY3
SDYHVqn/zrc0erT2ZICLakd+K/o9wKm8n/x4muuIAooCJQxcOFDQ12d4znMdTaHZ
8KpO/BMuCCpqHPwiTsLKNPLd7Ww2gWuY5gQS59jrwv8Ki8DQWc91/d48VV88YlPo
/K4Ro//8sTQ9khC8zTEZTvAkOfjnhhkgwCuq+R89B1wELoO8VMzD2/lowzxmYORZ
aojEZO0HWXy5VDX5i9Qj4RiavF/SO35+aMAZnGRO79HXiyuCPdb1yqC2yCHqwGPX
3mdV+EUMxGOwOvT/T1FW4HmdlBdX68JRJeKuFiu6HZB4mJE8KAg9YA9El7fLnPT3
dYFZpzPj0YB8g2NPVZaQ5loxIz82R1bz2AUPLg2mIqNWV/N7hYaM2/97wh5zherW
s0DfIViz4VnvfLwQs4GoLDRhTM2rL4UQLQG5axZNTLevKTUwVvERXE1SU28NOHM3
lSTiM8IlCnkG2W9o9qbpXjqXG8eVTxYcC9ismDQlFdEOZ8xuuw8qaXqXUJq/rwWi
APSoU1xuphHxGooRZtNOzYnr+k42UwGtHroW/yC2NS7xuPNvQZYCOsyAmoOFJjkU
E/k9KfJHTwe9164PxgWCfXCBjLj4StThqW9D4WWaZe6V5J/6PF+ZgO6jqM/c4/Rv
6CREkq2A75g4MQ47p9cOJO6KOkh5ztr9/rClu4QOn0OD8SABNYHYVuH6JAbkqgRZ
jBhYu1v72TNPy6Of5jMTrne3Mr4ktPvMmMS29O0V1kysnJfWzgAeOXQpGGu4Oo6B
Eh2D5fTOUqSRQTMBcq01QsgDgQDy1RbdlRLgIwUNfb3Psknt1tgtsQbDOAsu1hK1
Lq7eVKFeCyovzTnf8ZgLusQ9P9lngOKgpAm/p5F1uEvFVK9TZYsjAraBOShDT3fn
R9GS+/0OIjywjgAVvP5d9OLXWos8HTN6pbPxcNY69Dcsd+I79VjOLj+l9D+HPNsM
f8fdre4EnnpVisMJp7PhmU7j8ob+YGM808s3a0mmJeJZmNTeX76gW/fQVGRIBrf5
RT8JZqjrc8y7tcoSfGMs5hsHPKzZqVYIzfr4RWgSz0cM4bxYYZwHcY9mBxdvFuCx
WF8mSs5gYVu9aasn61nMBNfvSGSTdQGEl1JN3vdQa4g+gsrvrf/5J27/e/Tn+IsF
hr4tSj2bV05UaMjyBxFCDda6dOeeKDIkMCH4VH9NbJUJ8jUe0rolwtbbjZpGpADL
xfcjEDAGvjdEHyxEMVrrD1o3JlDirnaWKhIpHPWnAQ/Dwm8uLGvFTbi25oveSgmh
8aHMwaahC4sLwsrLGHBKZ2H4BY096joOQmBVQsmtkcrbbxn2bhCSXdUNzwNG7BZp
Mvh70jILve1mO7MugfKyIPWdVe7DAQ8rpOSGQWGHG8z8SjfwshEIs4Ob6F2HWqoQ
72bvo3nuUVPQunHMcQ6oemOROYQld+0uDFxHyDlnQ/dZzOgJuGl1V+Kzo7cBQMT8
JU7onQRvCD8W3jvzMqxzfa+0yOX77ZYh12LNknWJmJt9VOSeK3QTRoDShYxibS8m
lK2JlL4Kj9uB0uduc57G2d+DCkKSwCZXgCnDWHzNhbH4kuuAhQ3OD16zn4n3lWZm
yUzdTM96+hx02gGCExqAbsJb98kW+xG36vKgTPU3r2iCTCeLA7dalE6m4+pAMpFS
Bx1uBmrd/AbrKUsRc2GXDZ3ecmiT70g+2t5w80MiVquWETvrVigIpXA8VzSXm2+k
8izoGhQtXE40FIICM2BFlRrRo5U49RyZrnxMS4hFtXbdNbszzAsFhTdTY0Gk0CNo
Pq3bRHKBctT3prtqfd+CFzmbtNwETJN0KzVwu/GNz+jw3caoBduTjzKAWPLDpd2E
tNY96p1NwlpOqMipIoZbOHchTx/RegH/PJMBZ+zVoA81/T2KZk/tgGxfF7n5Kapp
xxpQemsixS1BYlS31jxCzo/XOE6GOAnULF2UnLM9vQDx8lcOQDJULEgcIUAvuR5c
GFEK2e+fBV3LffQcHCt1q3U3dgAZhDOey2TJoOVd+uGfXcjTVwPsyZLJsaSKltEv
WeUcSDDZfnwbrRVfCLLPZtrcJh2c4AOxEFpXI7iXQsJQEGsM24ls8lp1MuYf4JrT
DQm0u+cQ0pz7TUBCzdPeo5cS8LltYPPSWoSQzryZmr0iWJTyV3HTWSANRz5jLF9i
Nqntynrp4VB2JxyTb0pz2rnD95RihMyKTYps7lB3NeW2iciV2Tu7DGAsG/bvFzHZ
4Yj7tcdCpRcOv7zOBeQRhimlNM9DoXZhIZyE1h0qaDQzfVzZ5duE5yPkiLHGOzwG
BMxA1Ea1AbQlRGf5q/V5zYLRG9cT0LASp5kqmAnCCBtdMruSTpBxVR9/mNB8cFBG
rQJCdgcom2hOx7v9qsEowqHIkpA0rjmczMMjEiqaKmz4aoqnMx+kLKB6A0ccst+d
2AzesOySIMd3DZd7XjemUKWqBSWCROk8D1ddP6zt7qf3qk/LKdIo303o6mfwvL05
jL1LY+fq3ZSC8u3AGB+1ipbcivDQsy0JyRUGfCWsumhoEvJz4TGZJ0STI9xAfLBq
8DCm3VcK7L5TsE7IbisaR130VjfS7BnP3i7rzkCPIKMUkAgv4w25eW+QpW43E/9w
PmwjBqRO3KCvvLKtPKe5YzZXZjb7d8wXF9flBVSJzlMcj6jGtFOpy7J5NqVhDLdI
ORFXsQ30u0QRkZx0cwkDFNcGniYGWmZX9ppk+nrTIujpNPAQhy0PmoVBtbmyuy+y
icjGVpxqHCq2BcFkEBYrws7ODzK70uXkDE7A0YWyCH2HYGtfd35gKZ2BU6gwK4jN
/VMHJ7oj+3NoR4oCsSeS9SElYwSqnd6wYaaz/FulS4B0Q11F0rCBiX14kmJG95DP
7M1nTmCnU2k+hw6GtABdBzXlV/XA1JqRDhhvcA/DyKkQxA/itAV6DnciyqYO7akx
WxQq1Yz4O1EfZsSbLyNKc68kE1RqzKddnAf82DKMjVp+Gp+mTHZyTvHgesGJUd0U
4KGDzHLZm37NKnaJd31pWEIfuLxNVEpgdYpjp3xVrPPTekqhuntwQJOdGogOydqK
bFNrvWtC/q7IbDeJk+BEVDLIuJ40tAJTJ6C+9fgEyCckZ65c48k8HbJdAcg4l65u
WUPtEw0nVGsNoJSajdJcTjKGpkCima4TqtX6pCiEnaoN8yU+EnNUvEVk9bsOxXxC
IRBwyRnCHtUiLG2HRxFS7vhQr3DUotsVE5w5YBPcH45rZM6TU+bZKes1kePwowvT
QvA0sADK/PF/V1KO1DRd9VwR4FlxM/BykSLhedcwpnmSP64lPIb85LVLvCIqQ5sp
vBah+vjVbnBdDBucE+4JU8JlVhtVFmzNhgVWWcszivd/3w5lbASq+sIamSFpEpPb
CfKXkE6S9CNDkti/rcTjIOQPDXwvr1fU9feS6pvHdv5acWt8nIv5P7mUWE1qdBY5
NOjesc9sjFJnfGm+sfA/zoXwuQqm3dPU1oTckMdmf5OqZDavq31Ff5W1Lxkv4N0n
0Txj0nLdi2njjH4NlTnjA2BHSXoSQwKjcIjgVgPgsGRxC0GKngSsjLDMiGojweYd
RfR/tan73kWLHP0vNmEI01onkoNr92wcNT+HCDv3vCW+T4yp4HBo/kOd2Xo0wxyK
nxQu7XERfk/VsAL00GWKoqxzHSaoQOTI9Coq7K+60JKbC3B+02UIP74e/pawjdGP
ruEtAgWLRpFsigXxEvTt/BJvyeEm3SUgRO633uF/jrXcEUqznLw6I2JqXdMKtVtt
K7F/CqRw04gBAApOZfifwjzQmOuSXpCfz2aGkWHDLNmfNi6W/Saj5llWncfQJEXc
Diq3CN2Ccy9duPJNSjWUxExLeAhUYqvrklbAOJeofy6X1u4kAxe7l0vRadZyZvJr
AwZdT6iKQit8Y4msTCzp12G/GAb8W9iLEdbSRjP1HNmkvcazAzPzJDdDD5i46uaR
/QTXe1DXhscjhwRuEdejd0ble0sWJFKB8QovPWS7YyRLf+XlhGIJ8Mn8BEXn7Aph
3IxN6LT/nrIp0kW2dhSsTE8BuLL9HS1Qk96KaQLmWvgTPTzZNZdBWFlRfoENRKOB
lynZgvz1fPflb3cY4jvLRZE+F2VivjCzMNcb9Y46c+kCqFvq/rhItKNlNyZJD9FS
KSoUoXoW1te/VjNWuDGn/8EANgLfEInStXxs5elZL/fo5Pkp5KK++1lS/o6G6bnI
QQli9TGKvUdoYE4ICrS4Ao5094BmFaEzQXPDdV5dcSdWCSzWBb20X8Gebqm442H2
k6qsfFkFG4NyzD+2KdhqrWbPyRoFwDbOpie/KOmoM503KLWAPPIa7IjY4qyIGk3e
gLWVVmudhkpvik6/tOaGyNxVt6aNJ17DAUoUh7q3qFL/9MoMQtDBH1iIKbKciNil
dEGK4z5COh5AJugBP38kg7djodQt1HupELJXEb3uOeiAdB2ltOXjUJsXz4DfATGr
lzp1H3TDSMOX6EJm77wqxgsLHiSEa5z5srBR374oS3H9gLyGzuiEoGN+AkBH5JCf
FM9on1KuYYvt/gbEGV8LzBzw23LFkW2UoAtM4QFyimBAa0x/0AOeF6a3izBOyen1
Mpz/HZZ8atZeDdvMPV6jA6rj9FV85OgqLwCKqNTsVm0FeXJEDn331muR4zDuu6EH
h7W/ePni7EyzDY2Bx/txrvSk2l6MGdvQBOXKb4cGqi4Ifh0fql5latW+XQftu/IO
b222TuUoV1XkwhNfk02RrpZ1hVY3kavRkrpsoEIGfM8fiBGJv0LYxotV2yyUrZr2
NZidShMnwo+2qyS8Ep7YkcFQ7DEon65rO73aA89vtSY30snED9Yf5CHZlSf2ff+I
tEKOxJ60crJvDwcbgbRMMkEyi4bGSBKVgQGRt1/eCQLuDHytdMsUlN66OZh/DHMV
DApjbm26XcM5/fc5e9t710CSh521J9G/5BXVmc5NlE7/xSHyr9VNmW/wc2C48lz/
VrI3HjQx8rauey1habCZr2Zjj4ziDFU2vKsJX50krYs4T5LTVP4BIO34wRU2bvgl
LqWSBunaC0BdCtu8XlnmNvSmFNxMIWpiG1M+BmVziHzC6ohJVXJn+1hPEwfHUxkp
I2Apka7HmYNg42eeVMUcmgxJdr5wadU77CjDXCV36PPkPRLgoktvN06NBzFFxtRG
lYOudFcnshnfiLBP30SJn1hfrGNCRlGytOv/h9Svdb8p6uLDJ+70Pn2KCNh02LFV
wXb716IcfV7daH98SDFQNjMptJtRbkgMjZ5vDQWNxDtEB6xeTHVmsNIF7KAWRSn1
GIgBHonk78ELnDp9QVUBIQykF1qcrCV0nNZmKzDHGMh0bviInd2x0qHpth3hI1nA
gsxc3enrD4VBD0eUNNkDvqWNpf0aBHdZoo+eng3Q8zYOCG7AUz7ARJD7qEZ4cuDO
Rv4LLoa1oSAX0daifBInS9O5BRgFMMqCGPH4Lp8S05nBxgxYoE3ukbquSeqmsEcy
/UGZbcoAmBLYPHZpspZkpYizZyBe2HBeOtVBI62jnp826RVcFf5dPfGu2xYZdoEh
rr9vXyPb6Wrre+pBipZHjMQsiVNq9TvM64Ldy3yiBt4zq9RTKmYsPqXQKnnteuoy
CJewlKa306pW+N62xncqssKHYl5Y3iKiyahNq3Szg1/cvJB2jon+VI/1OtPtTBVP
gapcvBdm1NRvnTCYlc0KXnU17Wm3qAJafhAzwj54tjiMEL+oTCEx25st9Bm55iRG
RRFvG1xrLFmBhTZLU+nc6CUxh+KpDy1LIHVxRJn6gBS5Eci6LxW9YXxiH+foaUlU
hc0eR2qfN8OE/qixr8NYScogPuwf+f3jkkZTPc/i0GD+l9pn703GbMe0FyWsMYDQ
/PnmQqFgdzi4QaxdMhm+q1p1o1JJlbW/2sTsa4edo/c2Yo9itWcw00411AdbCu2l
CgqlYBDw+m3Y6tY9OR/BbNEvIXOX0WbH+27NBAr03b+S5LAFGsMJml+m8ERKFs92
Az/DnnuuADJbqKiVm/vwLqCkBAJFrkEV8IVp4k2TyLLjWh0YrwZYcie2iHdLkqM7
ODWkbtTGPw3UEgaxiprw//sH2VjU8PsI9vRcy2FtvVDs3wURzy8D9HPCUumGf2kE
wcYLH5mWIqP/4KiQhFjF3ygf4adwaorD6TOOB+4xzQWznsA9oiUJ7EiIY2qx89ud
Scy6zeLEU36DBbY4QwmmATOGvbnTiApyGwv2jWd8dXKA/OicsawwlaBXsG5zLpoQ
asdzK09T1SmwyG62YQ1cwxX+DZ12BBoTMRK+e/NNSg/l9wEM3mnfhD0SVHu5oicJ
IwU3fWlT8J6GPYUSvHVybhSzvnaA/QYWSzxEk7yNcCSCshD9vG2bwAIP8l9YCR/l
QeCC2jSGhVTvrVazvykd4N0SwnBKACd1dnvnUE545K4T/nZJYIbvXZ0k+tVelsg0
DjOG5qilG/B/Q42ONjfow+kV+wO2QXQFc/ErDmDmyd0fLVGVOIe4Jv4JFXJdSBAW
xjyHexYt5fJhwtqMGK7hO6FNJW65i6RFe7btPmv/8HEnqXvOU/wN7aJYQqAKORTk
w0b3/GAq6aYPv/wNeaYWyNK3FCaC/Hmt2NGEiQdmIDZlD7XnMZmsBwJGwLwBjzoU
PTXBRmOumSbYlWqCXdJ2HCP7e42TVyma01rnlJ6U8lH6tINLH28RJ5vl88td9Yn1
V/hgsNBD/7wkN1rFYuApXawlnSp9sQppCtS3XTVU2zyaUV6j32GOYuNIqrdPX05S
0nGKb89sGYJHgUbz/zA5QtrYsbT3lw00otF012/nbu19yO8R4ZniEnE4WP/51nHQ
le2/dv3W37Q3ivxPE/1TO0ObGGN9AxkiAmzumHSB3qxu04EhVqDaVfr2B437m99K
pRsviwqMCiVwB68ZqDnyAwcKSSxQp2hQ+oY5DDxuvcx77rdW95J5ZNMh/U6Hnt5p
Sgx6QUmwQTuUp/hOdofshT18dMHW58wkqWjI5trdPTQZzS4eztD3qULuqJ8wMt8o
SWwC9MKCMvU/iWDQ50ln9wVId7JevIW6Hmw5dNsqZ3vzY5FltZsN3js8VPTs7AEr
n9vZlYnTd4VwfaZDSuBd/wjWC8at6DBftgSEyLk1iZFYHcE5lvGrEqEuu2OqKR4C
4TGlgq+N5j49Xy+Vh2sDIfri2QwCt+W+MVKBoPxILC5sHDHWsVnu/nJQRRdRYinq
bpYj5gTjO9nkP0ljKfolp2j2kEmBsWRxlGFPEJY/njjX6pJuZrvrQPnQT/yXGSj5
7qsfrat63LCRxinRbYCZdBsojY+lOsYNM9M1iYzGdl0hcQIecBvngw8ES4nK0zqL
YrbX8ryCWD9IddwZjn1dScfXnLsRsI7y5V3JRKY4Sp135jyplketCvDnPVa+cWFa
AGE1nxoeGgRIrLOJpMqR18Z1qHNDHh3ZqPy28E0rRtwECTHNMItL6NB6i4bJ6L0F
JqCJ00KArpSeDrA2viEy5gjFAF05Y3Bmnqsc9vYV+SrYbVn9A53TBdoibxVFDX8i
Zkn1MzhsJ70q5hEyCbE4UAHnicahlKgwEPFRYtV94GB+TTxUL5/sXcRvpCZIrjol
EgERhJT5GX8SxmQ3bRVewFXqu9Ec3QUrPYjWClPi0OwhhU95/G6qOdqPwkxth+Ir
NiV46K5BeDhNaTjXc1AXPYSHDKqx4TIGKjpvtWZyuKJLIy7Twwo1eNk/ZBfZ+/E0
u1sMtPJ4Ifqg8iLDSuqBDdOl26/kmo0qHxtTYRnft67EeduZGJAKmE0/tYyYD1g+
9wM9lwELprM13QL/VTiGaAbTgzN2tFHii6FPM9TFPH83r7vQf1HFsOG67w9Wgzef
wtQtF5NK6GJ5pxAwOK89V6eJ9P7f6UowDlOh4XgTqvguJc3uaCbP0KEjWOu09Brd
3j0e8YLtJSjEcf4imP1lMKSME7hN2ibScVVnxvm3gEtD82RQT5l8YoVRNjXer/SE
yi2PgFnbBlcxUv3AA73bfCxnl16cXXwsCP7+BUppsQXIPDcqpqhPs2rozqzhjfRl
n/rF7gpYluZpnpIMNDzoosEZsy3gAIWJ1mfkr7w4bweqlLmM2XWhV4iaTpd6S1hf
UOG2+Uk8lnhy6lFj5jhzJNRuvo0HIsimr5CqWLGg+0MkE78cF6CVP4TA4DddfBTD
0dNcxvHwzJa6Xv1qaYsPm5TnS0FVi+K1ku9lC9HNMmslU6q0ZJDDbyCb1Ujx0igl
UKLt7YrVxP8pJrlc+mg27WTTVtnis4FXVHrx65pQYUA+WSQIbCmrgj2gxaKjYjaR
7/iNeX3BoaUr0g/sUVDjQyW/Z1zSqDRVTGJsNDCv1IlO5GDqH3se018SENFg3Wai
o97PSSxJZq6/rAdoQxk/YRbhKTj06J0zlhKcN5KPcn0CrNF19NrbEmg/0FB3Z74p
QLL589idA8TwQ8jzKoBliJp1cNC7y6r9Z82PcEtCOBokgjK3k9PcwTCK6sbo+tpZ
EYZdBU47FVR2CPJna9ii+1DfrLvsAqWnnD9tKLNKPNp0wEaQ6FCzEhfUJw4l19Ng
Lt1jAcIx90/K6RyK9UBnYh/BJQo7SM4GE2rMm4V4ixDv/+7cJlOxW0Sijbt1acbV
xFM2arXUtVuD8Uq8C7+nUFGxeYQNvrTfZEWsnuTqdOdBrfNBWa6V7O0zpe0v+nsT
WZ6ameIFPHMKaMcNGnxrjYYGnfmhvDT0ixPDl5535/8CURUrceiPY4R5zKHEvE2E
QMKzsy133z/Odx+vIPhaRxpv/jLHwUqloUUwTUGlKpYyOPLOSl/44a+kC2vSxiz0
4xyVifkZfU7EgbX1SBoT276sG/QRY96/wALWuRM1p60W/2TjZVam5B+KxxyEsvF1
EUqbVx3BrtgApu/LcLDXrS8Re00oBAv7/KNAU0zwSTwcLxX2JG3WEuDGndygLYZP
9KaipwX5iAb0vZEFqUOxduXfvyF3N0rQZakMaP3kaTD1tGDavNF9A6w1TS4VB/7X
nAiBGr9HcDOt+HZJ0jut1f7+7AlRbjTdJ+28YTKuqWR9VE8U8AUpIvg5iEZGVJob
IeZydV/M29SDr48d/upkcW0X4tBPp8/+O67/56iaC/rARkn1mAHVE2AZMiQ0/YNz
lLuy2CZqtHG1b4ZgAq6JKtnbScCyiJ0EUgXTY/uDOt0uTfDFvLqLKQZwYGxZbWWA
OCS3zHjdtWLUFTH/M5U0AQ1xHGKqcVWhaULe8UJ+qjNXnftixwr9XclQIId9qcK0
tgC9qTmpGWEHKgMVhtVk4K+kpoKsMWnOXxJZciubP3hAzVGVdyTgRGtzI9WuDVJR
BsLsz/Lbc4Cp5Xwp+8b5jItTpyUmP0UXbFeiJ99jPhkJaWhFhIeDpWPHijxAvxYq
wi1VTKBRZbzrHZS9cercZaMSDPWAOsVDsR4mxXxnjEXS1kH8mDLpRb14IUaYEgVO
soVAH3G4shNah30r4VDfr8H2cNHpBbrTddlZcwEuwaPHNxwW22GNZuFYXcXZGmNs
vF3O7dylgszB3l1jqH66C6mNsvMqrwYRF08OXfTe81AstW2gg4GKQcHPgzNBBs//
av34bnbGGS3jpgrLMivE8xuztGcKgqvJixNao2tNAmqYoej1rEGQaw0qvSRjQYlh
nLLl4xmjxsWaaa5Sl6oGh84ESNwDfPSdLVu45pfO3VqgmBAZSF46XftNaI4HdVzW
rYMguJ0GoEGIE9pBGNpMCy9y585TIWgZpheTMx7+QtITLNgHFyh20jWNkt45SDis
TzEc3LUmmfNdsIXfNwwWIWzgZiJm6/qvZlG4o/MQ33IOh4bK0HPIHaYOIP95laws
Tm0JGMHEKQlE3N/MN4vTXJBhkzCzqFBmoUvICKiin/6s4LbSgmhVPnLixdOhDFQJ
vVsBH+Tri/EbagcG/S+p7VupPAoLBoILyaA6+GjLxXBPgjSJnUtJbCHkkdoIwl9C
Z/uLu3MSFSlIHWzNJwmanQ+sCR8Hwkbi+W6QjSuUDdj9CYck5KmeAd/yYSOq+vLv
JiVm/tVTzGDRzPXl841w0FF+eG8aa7UK5uOt8WH3m/9v1f3+b1tpmsxxgt41D6sH
IqBj/4B02hk/kT7BsKWSXkrUN8VskaE/oy3QvU4ExcOKVkWr8HgHNBrRuspb7vV2
wh5GOuVmSTx3Bh8nFbag/Ndvy0C0SwJ1ieAbH3W+iuEQTQl1pvqviouYBPjGcHPK
E2nAa+HlF0snsV0A08nXTtrHRGuxpf9z0IVLYXcTcROftMd/Xgf8gl03C2Ek/Q83
dR8oWULx6qutYi0KxY3r7pp4rc2VwSDx+yI29cSZcxTmn12wL6T3an6+Qmz0kTkN
7MiJjBAU/xXDs0QpekGNNAdzy3/eJtiFX9SZYp3rSQbZR8GZytnfQSoK0B4AhjDw
CUr8/yLrKpbwXqTh6GYHHtjRQUsRSihG/wN/l+p1Af6GX5FNGNduupsd3xAkLyAj
N5Ink4qWQVlxMSOn5V/AwrGIJxUlNV+aMFte46yJsxMSDQssPdmLMplFhHXA8JZT
CMGi4IKnL+uDZjJkETt7IYzE27a5dHzCBXaHU2ythJbX31HP3TGscVy929bf2iyt
ylF0/V/cOnZ2WNorupXIwIEx0QrorqVpPJW75hFHkh7/JKJF1+JI85FJFaNOwDbz
4TfhS0ww7mpFF4EllpkNqCMTNIV1Lq6ca7kDXMkGgHmVeDAUYblV9OpGTtr1vj6n
Ayiay9LOlA61ZEzCyM5PpMwI7314zpDGv1tKlrwDDjJexJ7t+mhYf+kfUbWXCoDp
ZSkytF38bShDS0FeVNmIv4XgX8V2qA3z1alZRQQtMvJER15QABwJ7e32pnBuGHrK
VGb8VfTAJrKVb/9n+8ns2zumO1m1tNYEpXQsFr/OzNoegTMxQFQd0nGR9t0+mGiu
LgdKElV7YfDYwip5pVZIue/8teHJIDbnz4y/DSrBYETFm7ySriu7y9DZX7TuEIeP
W5XcG0GDgmBtHOuLIQipYh/IHy4daZJTgczAZ2+aD5H9W38beok4eOSCIrumUZOm
46MMDtPwYMvsO6nTiKzwd1wqS2Syi/bvw3n34bGlcSTwDO6jD7+I3BoW3zifRnJ2
qypynwdt6j5eaatEI5HzygvpBTcW7/IenPJ7/GRyTmUUKniLw6JUwO0h6iGV5Y1v
ABmqzFV5guk5xN9UjPmdfEcFQFQYb95g0uS/DQujx4CY0usH9ru1vsjGOhmBZN+m
l1ncowLmk7J5w5TfQW5jfgmJB+wDy4rXk3Ow2GSdpfH36HonQTVrGyghYC2sbgAh
jnKqP6STLkgLu5WsEWMFx1UXX/DgummMn1pRd5HYzJAXlYXmuASLtJsu/yOfge5i
MNNxP+78a2OcP8EEt4s2W4wOnPt6zWFo01aqWYAoxy/8TAMG/WsaWG7YBnhGEM2u
mFGqa/KIemjYgon/QhGZnZUoIKXduix9ST/kpUruzPO7fcVHaCAV+GpwYu12Etm6
Ihh3sG+4reNncQgNn48+8XcqiVYGb/UPtQA0vh8Iwe8i/Tdyj90cyAfsrkt6qEgy
rsdRHWo16tlnlG/UoMvH2LkqPPjbnazFv6VZhKWxqaOkox/yNOUbO2+RBWfqSCaq
NJKLOpk/wjypGYtG/sQFnSTEPR+y7G1748mTewaTLSQS2ANSDvGXWNDBBC6WSmhG
bo2x9Z7jr5Md8G+0VU88K7Q1Cu3GgKhDGL7EgMJpIbqW1pcqwXb1SHMPIWidOVBv
CqVXos+oaytwwJssUqo8bX4I5X0fE1rDzfXKjqcR4c+VSGClmjuv6n80nF+o5lDP
4W43fowTYPpFhYnrJNs9GQ+V7B6YlSHixcjN4CmUiuZmHQ71H5/WCCRMwdOj6s7u
s4lZjvbiKLCL6faJ7Ztc7qku5jlfIF4cxdyz2kvFtsPOW+x2SiRBr/DPCb8LjeJ8
ibCGCSsVEYyWFYwUvLu1JbwVoftS3y8LaQsq6PyOgoGzVFhsWqG3QMQMqiw+dhBO
0WewRxb6o394OxqilGYdHAJB/00QWuMi/mBoglpbPaaMuLntGvzTz8xX/jE1zBHd
z2a/qjicTy8PTfdsMOFCNB21bCUYc0EzkKQHfpAV0TPd+qMsXxwpOXuztMFQTp3l
hog1mThVtQV9vY50H1XNSg2xC5RCjyAmKykYySTkqd4w35H6fp/aZ/fV5v//Sp1r
GFCbfjKpnNTTLF6EvDHoG2EyV7AS3KA/TI33FlE21R4HExjdMqgTz9alkOwssa9J
N16MmemBZ2HZbTNVIDgvnAe6WRFtGpGhodT3zdxxWA9/c5oAcexKEV+E5Oe+xAQE
JcgFpFxrsZR5vT1VcQvuZuwNiFWIefOs5OcoTh8Uk+BZMAy4vzKpXm7VDEAnBmY/
AWwy9GFKM4zkR0lSJS4ARu0rAVDMktbewcm9S7sechudt7C0v0eYFsj8wpTA1VS2
M755A4id4T9snSbxG6RdmhALi5SU7msWqoTfPnUNAe/4AI87GmAN9mt4x0922JLy
bqOXx9ELTV83zlDgy4qvTx+uf24WxHIkSP4PFW0+3ZVP3ziCK5xyG8lNMcwr3auR
Eb9obVi97pzIHy7Phh2uJY0Aev4nGFKu4cZVKvar991H9CwhxseA2i9IAcOZzhwE
nBtNyaXSaYrahQhDrFGewP/XEiA7QC9ScmMm7s3sr/ckbhym2WMXNXdK+4ojjQZn
brMYOWqX8DN6ZW7Z2sBlT+bWYk0MJDluKzSUUX5z44g5L+kJXWr67NA9daVBsZJ/
rBSGK+L05BUJPDpn5Jxx6SHgNkiRdmc6I9NJ2G8wTbepXuwqj94gegBrYzZOZODC
Jn8ae/JacvC9zNqRTaPzhmN2lA1F+XR4cKgg5iYYPJ9lpI9169N06NrRji4C2MS5
JWFPJp9oXzzyzWBW7WrJOuy4/2i/NMH0f8GtxYnevdVsyeJs+YPdEGSV/TdVoO6h
JQIRDjrPqMBdnxzZhvGi7PoFO9cEdS0OJVnOBiay18hMtxYaU1J+GsIVpM6D+QvH
3u1ULsFfLKny3+fsfVWXGZ6P8bmQfFFJJQ7YDK9BTK+msCx/72uCiqR9dfzaYreS
RONufvaT/iZX7XlQuNusZXBnKO1CxK+hUKjreZNbdNuzx0siaRJPAsH/Hb4Cdl/3
ZTSodymyzGTM5t7MvkYS/FAIHnGBS9nFRT8BJi3AWC4/yZPTInuWRDpi6G27WhF/
7+onKIq4abk45DFCoGDU5MgSMlKOjQi8ZneX596EoUpM7/xc+GcxyQkiUmWw4D7B
34Ce5+K1auUKHFONZw3K3V7K7BTONbbl/chD3VUugFAV1+cwS/WET19e5qlqNKPN
3WhQvL5hpMjO5m2QUc4ETILZGZvwH1w64vgEmRivPNuftJ3xblDh7xovTcoMOO40
kva1Y889ELmK+FiCPUwYG5DX7gYg8bGx2cVWuAthZsKh0atMWaERL2liIsEB5pbh
kLDbNBzxi4mmrMouqbq9Ts5AgHZk+1cv4yBmAPsxzPEs19gnwAtasshJ7Ao7W8/S
lz9h4d34uGpWKCu9+tgh7OSnB9Hh1+tXLtm4hQSQdnhuDN89/0ZC0l1RWy5+kbIb
Y32Bb4kE7RUWWIqnszXRr74iiSuo+sdA7F5r0E9USHXEFtY/GRetBubKuNu88MXw
7W85SKcWPZPzSubaQoO5phRxiCBbx4QjPlKRq8qoFYuewml7vuevC7BgZlX08MRs
Csg/STj6jbefFHGHOVqXZQpXF75+UO2ZDmDlxrDJHns0nDnK2WqKSRg8pfh+zPtW
+t9KDbjSFrHySOdNkRuWz3sFtTJLJZGK8wiOdsWxy2z+nDpohGzDxj4gLITWWHMu
74VeNkfn0xUHE1gGn2f9zoaDKp/Ef5jwwXBb/jcj7T9mqrrRnBMT3zcGt7Xal0RZ
NwEmWnQZoymNGv/c1X/w7ot1SR4gdi162OiWlLoQr5ALjDkTxhRaG0yOFsx1u8kM
CxerxTq14ddkVknsxeh6e+L1BCU8p6sRrAGUhcpMzB96Hb5UOkzND/wIb1z2zxOU
skL9qmwRkZGeo3doeiFu/pG7eT8dmxVip+s5se3GTBe9Y+DUhqlsq+VONi4isbJX
Eh11m5LISeViX2C4LZmdSP9l6otAKOH6X8reF27UD3eLCCsN1pn0EU2gckhzzTuL
ryRotxaSLsPnDRaTiPywLyZ5Z88NZvwy6ZNLdLjjLFCi5z8gKnwK7pGBYeS6ON4/
uyuztu3rmd2FmCZULIcXExbs+lD8hsREHEkZTMCk9vTEKBwTLEG8JDlPk96rRVjq
8s8XRhcOokf/LpNAQpcZdeFZAXS1owhtrvR9qhndNWd2jMqlwSWt9j/50+BdfjIl
jbYF/4OcHRUGGqY9c+kJDmAEroprddPBZcJpgVwNAuKBY27z60KpxsrNOX8j4cAK
ZCwrluGRrDQVKxEKXmPqBxFcx5hclEMjY5+bUHgA8Z8Oq54p7vJC1p2Hhc/EwB/Q
+bZmCOiwoR45lDEQzBvvk6fxpZ4Nb3TxovWp18fB22xI3sIZBofwi+WsaxwLPTgO
bQitet6NPR2HVrA2tGZF/IkV5sGuwWVN59UXJpHqjRR+MpYu6ZYUQNeVeIZiNAm3
7EfvK/5UNy66D6hP0pw5yQsFtTObGihcL+T5/MymYTfzKArDgkBTqBcpozBLzbpq
k5jhsUYsQNlurCSj11Mod7fmX+4lJJO0DtCWpvO5XowzpocTlWDqFUOTJrGe0O/e
Fic0DT39Czb16JcJDwXVy0Qew/jdtq9R65UOno66mK7i/5M+GJcGXzB+3WTs/+XO
Jupv1jXuyoujI3Vn/lwV82Q7LkJQ4DzSDIzFHuVyQ+4MMYZOlleVjLVtLkU8BKuI
RIU69x23PaBfihLrS/EBcT7dRbctv2AO/aOGab9y4d1jmhZqc4Uu3/G0XXY6vQ1k
r/NRGAa2EpH/sfgpIbFYjoIhB9sinFDYRHD0GIW4d956K46d+S/QwxALDV6cKtvK
2SIWWSvsNOnx6YmN96JPcM8o73MpTk7nWE6OZzPLdyegryOLMsxlmn6MQv/wT3ad
ppoprtpf/YsSjwLWZRy/TOOp/qdjxgD1eCXwZWUjKrPvewopsqi45v6hnZmvZnwO
DZ8poyulaW/xVrF7SXenb5xnNjzh9tRmL1tp+JSKEGlPOvs3ebH00+RlDxb8mlPj
JU830L22yw5l4z7fDnQpzLPPBDgANuL35Xfkox54O810ccbalzA6w32U0bzkywpW
lcqq7aisLYcHVdjXPrYDbYRbmIN4ka9lPUoWDOGjitENBt7ssmRTT5CF6zQJoiAQ
EhadnZALZmhYwAoktd1flaNXOj6dXKGQeDCL11DFkiOhKLdxXnUSwWl3NZXUjvp8
+IMl+r9jKT/MMfDcaLzxjyFftGMlwo/iQjVyYCwqzNLUJH9qcB4TRbxto0wA4Q6s
bHqnNrPJALwoYBPdE78CZHdgIkjb8gwwNQPb8DE8pv1FWkFxIw+vfeL0QLf/7aY+
LBm/l0gMTPuasY2MagPpqxIP0Zg018gihEEQE9TPqvBZqO2nE67sTOt738ZxHBwh
5d3+yP7u9Xw2qGA2m49pTYP8PDq/lPtST+tpkFhv/g+zHjsYIr0nK+uqbBVT7vtd
5smVk3Hjgk17hUDOWELy5j18U4fuEeDYBdqgdtwTTKH7L8hso09Y2J++ruGyahfD
zE4i8Ek30SnsiPs9M5Gid2z9AULvD/hl/fAHE7EzlAicjhdJncq2dB1LxkpbamsT
rWHwFKnaoCw9A7zZsiHnvhUq9CpX993bXss5MIxzdQd5IvzTQbvUUPxMIMO4B6xE
/IUy/aJDbr5S+VwvqZH9BKv2kRmmHMioAiipPu4k1T29u7Hm1bZ/pyg5/sXnTQBd
LZYcqXqtyN6sfkYDIHNpi2DCPs0OUynWdhoe9CbaG1Svd64tlyEGi6ve1D/BitQn
UBQAS/Xg7IpJERsH1ty3jx+0BsMbPKZGiCDKQVAHpEOyZ3BBT4wMosbe2zzAoTuC
mBWHq86bruL1OfcQKoS8oH5RdxuJ7GCDxYUfsAS+SujAXqNIlzHW/oxdauhXR0kh
JxQp7UMUSnqVMeXybkt8Sgbj74jrcmyzvCzlxUhqwO6rMWJ8sgkbJ+D8OA+klBfA
+fCM+VZFUkEt1uoJ2Sm7HM8OOhl3GpX+5ptTkllBJ7N2DDMfKjwjlH8ZPPgF9q37
sPwr9IQ4C2wDKtYiPp5IW3kKghp6WlqknPvASjFkL44QuCOamRQHzlArfDK/vooM
uR6AHukk8/iFNAvsKJXyE1LPXwoqB/nM38ATD6lUE/mj7ajeMxS/kxkOAgA/5OQj
S+kJ9B1FYQPomNNWL3vCZdeuz9RPyRlObaiJeEXin29s3h0oTKM0ImvB2gLDPhVZ
IbOXSQUqCDUTthV6vqYsskI/IVlTjy1tAA1dL4q5sCCcBNVer6crmFDusPkt4GFv
0oQb20uAGgLUJUbeTtCw5jw88CUFow2lyqKnPtgK1WxUOcEqD1A9imDz0hLRE1KZ
k+CFKR6sj3/z0vY4uv2K+uznDawS7/WSgc/AgiQkzM7qr2sj95s8/xAta8nny8VB
yQjtv7K1ZRPfTZL1fzOb6XVAniM4d4YdyDSVotoBSdy135AoZA4gEtaHGSz710Wd
hz485edyjBtez9MlnqP+SaCJ9nTS5tq96lACrHAWapNdVw26Se7R/x7eRNi5w6cF
YvO4TtCglSEPq1ZTXww0qZOZQHO9v6ic3uRQKKO1PLjYSDYY7TSM88tz7SBE7ZJr
Mq6PtkhFjw55/fp+NrNYCNrpfe8f9uq5zoZFWQqMROmROHzjZHOtBg2MVdg4v3/s
PPmBJfAcByR7qJxWGg7XN1Nsze7z63cZoQFsKfriPLYDuLlK10KlFyjqbXhAO8GF
0UGa+kywVRIyDrpDNn6pQVj4xQhZijefjVKWR2kmhbC/mhviHL0ZPrMOoZMmXVwG
pny0qdaYHKKrvdrrMGBT2l3+DSjVKjXut5g6oz92giPfkm1+su2BUs7x8cy9VoRv
28eY+ueUi+KXH4EH980FKN4hAQWzcAVlddVW1EnaxVZ3tqahFkKdXjJFcFoeY5xx
l9zHi4w5KYkH6bhObMAB3uFAq7G6jh6qYEYnkGki8Ga624W+TYT3k7rbRuBW/4sR
YsF5jcfnZ9p8Gi0MS0B7c9EkFD2sd9rti+ar2OQ/sWguhrbEMVpUOc9iTCmOxl4L
7diCovzcXaupLJ5nMRLKinBCCbE3wSsbCEa3IlXT23n5ezy1Wv4UBp4XCrGZl9Qn
cUz35ydtDxuTv6Q81obnEB8ZbM+rt84gY6YrnTGyk+ZCWnNy1ODrTeNaNO2Dtq4v
E4INNwjG0Sl9567Ewp8c9tyw46cdFN46sRCKTcB7sPe9b+XvYvI5+GDS0aVXuqis
3ldRcbDflq9gCsNUIDi/CBB3SbJOBwMEfMjlmAyxasF4BZz5K7AtqfDQZr/BAeTn
10w4eUid2OW9WU3bAwE+lx8Zc6OljMeKabo2qh046G92O6O1r4Q9fltDCULlIhTp
9UQ+m5DiosOSD42+USdxor3chtSu7UMxC5/MBsZReOvWeswhzkzSnT+VUJ9NbBIP
O5y6U1gr+v7k5ALTo+Ocy6Te+KRIWshucBE+8P8lrDTWg3MT9S+IskZzfuFtUxZb
ylNBwCkfkLE0NChq22ccPFkNDNrDcVEiCtBvuyLdgfZ7411RPEYC1i3QNc5JTbEs
6at6lZ8jfenyfQMUdEdL5LJXVmJcjRtxK06dcOpga1YE853ADXG3HFgLajykOuJ3
KSUyFHq7a2hzMqjVjfML/ZBnio3b2Fb8W9Yev8b3jDp3JMj2unhapD16uMyTKBGk
9atSuaDsyvlef5gAzQ/es8pIFbJ2G+BLYlfcg/ea1+KmA6nUbWuBj1E/oRMJQMfs
P8zcPKUgli4XeHb89Imd3Hv7I/N+13fmaGlGbcnEHVL37/eHnQ/FE473pP2zpsea
fdZImAMGuE56KbQPaYYRAq/3wS6u1/LNMj1B4SFmZqpIZQM9fKi1KB3a2sDUGcaY
3vi8ObqKhYt0Ksn6/xJN/mIcPtoCOlXIHgkwUWLOy1DIBinZf+tJJMWbeI1WMpxR
f1XJ8lzruEPQavcx1Id+CNmh/Lre3ooWZr8S4qJbRUYeRWEWzA1Iw5b8Q9xUy0AJ
Pn7EW7ybGFKJ3mniWbAU66ql9nC2nKghC+VUuLBiQSQWqYYX8pmmErhvENeIJt1H
oAe8DOyhigFljt7fiEaaNwWKt7X7SkKgNXszyURp+ETKAs+JCxWu/og8Ra2sWXVX
pV7TDh2IeQjtpmVmql/LIOFXvWWdgI4OSU+M77OZhPFoGNCVFA/vdDnAer8Fx34f
Kp4qqHQ15l+JYtEwJzMScS1HkWkFcy7jAgJLGxegLFuioiTvhwBtMXnxVDoMhy+e
CmO7vnkQlobHY5NwhBHJF9fxsaJtv1tjsfgk/Ujp+foa+PW0ThoyIyw1VkOi2ou4
1vhDHl1xotpKmjRapglN2VY2JibkaONEmhwddnRkW50ker0QNQEaSbcQbNMpujny
7G9FLcBFI4Rscy4FiRao4VPtXoQBbFVQvqz3t4xsUHCGWie+O2o4lV8K82kPu0zy
5aVCZvCE4sF4xGcRkztjWKvkIcK0uGD0WS6xR7G9Frc98lDDLGLLS4eIk4TXT73b
tnE5u0liM0rF/v4alIEHP59mj7dHyEYfsZYp8ZYdPZm6MayG8oyMm1tr7IU8UASW
ZNzcvCXXfwZrkbfg5Wy9klNqaj79bBXTg5g1E0Jd6TFX6TR6exhL2yQ4l5BFuy3L
tuhf7Q9LKQhSd7d2PWT60/vgZnh1ta9DpUz5esbo50y7j4Qqr04UspZabTHbzDqz
hHSBZxliwjOfbCQZXPPS2AMn0QSS1pAYhBLT273JoMKaiDohxyklEV2dscIwP/Qz
09m9jIVX/D6XNk7L/jfCoWkqvxF6k0LyF0zKbomdEL1dcjK8lEH28nsLzpqDO9vj
MxOQafpkrowp0pF65Dqbdl/Jw8Kus+jsfQA9YIaC27Z5c3AUIunh1d+0vgA+rVY8
VAhVQQyQgrl6Hfm1ochofv1dXiDiH43/GMBbnomvl5aOOLh27DzJ7CNs82gaxCta
QUF3Ju2O3YAfi7O7oPxUtV7aLBE//GxG3j5Yaf16UbewkS6suCixilMjqa73oqe9
ePiqPbaJ+jL/jWtKpPMHdz78meeaR/f+B3JmmjYny6nreyFyVmDcko0YGHl3QzpQ
blUAP5FsFfuJMKx6AyRTMZqcz4bXqrr7+EgJcPWmZZK7mnuSwTZl6Q/EFqgwuhct
rWg/FFbMKTKrKKimptSZ3zB8ywJnkQUfJSsUsW3+fcvBDgVoTGNrVzwV+i3NvMs2
F7bVtJraNNsK8oGLfsgFjm2HE5Fj9CQHrvgGWOeCPfZCaKOTMMM9SY78t2BkRhV2
SeoF7Z3Q96kG9tfvMVsRYW1zDbxnCIIau/VoYq4kxqjylu7pzKWbDu34uLgHtint
1NceuOvslY50NmWp4yXd/PdpIxSs1TcOyX+xSM8qhQ1uum9+zgePNHq88xPUKW15
4M0fTar/ArOkHPfqLKcHjYj0x/za75DBsavOTgfbEKYCWFu+09VLvvzZi0tLcvB7
zH1s2zSJBBk/NcX2L07ahAPpQX2Xpng3GWVMVyR4YNJsM3td+Z1OM4sSnlmJRw0y
TpMe6IemcQtBXt93g6u0BdnPj3uNL8nSjHC8wWbX7+I9hMUwNC3oZvxV09G3DhSx
Kh4Al9rPcwOJ4kgmdZziQYGKxd6kcq0OdDHKv7ndhos3/TkGwesHv+VTchewvTwZ
0Fws3aACt9Q2rP0YDjM58T0mnqXf4K8w3IIR3yMi9yOw1sqo150kOCDSh6UJouPy
YR1bOfWZhVhCEOj5fvjEJC70lw34GqCC/tAsTUrfanEcIYEGAyg/rVR/g/WPA8DK
IuuVLuLNPtMxxYXMucyKXTFYtb3rvZRNNe7Y69pTyWfb4W4eyUNbBL0UAbc5Vc66
nx4AinfN3nJa9E9WMFh+AsYTW+uFJ7Zmiv3GN76xZ+MB8kjruABeBWtGkvvCS9AY
RJsNCw3AUu6U10SkZM5yUECvTOLH0+K+W1TowYvQi6617rubA7X5IC9GcfrAgrWo
FDJL/XbKpwWgoDJhnzdljHJ+U5Zt0PlC91T59KM8nPCWZXOUd0mVBx0cs8qTgQXI
wkErCRTDivbGJAUZ6tYNWoZTNpQVun52hO0zrRCk4TB2H2t9p0kQOUdsSfNiqsKh
oa87Cp0bQHeUDj8bsFhYSfhjsTBWoqgU9gr2t8ZH2c8nXlJqIRRmgCyNfa4gEg2n
bYl4ms5+LbPf0XDCf8LFcHSd/aPSZzaz8+g/extbROcmIJ7DrngX6+fRmKaL6BzH
5bkToxQ6VokBYLgK/IglccMEwEpezPyDkdopm6uHEcNuybELe+sLZzYFN8GVUAKx
rDu2hgdZdB6HZZS+G2NSQE/KXGH3szPgFd0OBbt/+1nWKuB1hoPBv2xeJSCk70w+
ZJPstOTj7EES1apjiqNnBuji/UsrnytgUCzvl7f2UOtSh4yo5npc3vaib4NTlB12
VNxWfjG1d61snYSFtDb1t0Di161Z9qMD2KdPlq5jeNCpMzfgM+Br4AGxRm1VkDVr
/aauZ63pa9DQSH4FsSzEgQiUOEBqoqYp2K7hIifUmvPx4LMfXyajmfaWRXEXfrn1
hC+NFpz8m91tyza3UWcnylYwH2LS/cObsWXkCDxg4vuPe6OTyrtWk4Ted+Sx72o3
PpjWvdFpjiIE2Zol54AGLLolKneco/NEBivb29n7cEJU2Iq3/f7zEx8ZvJz5brPz
x/D8jkqC4rlMSSWOpFJj8bEx4MeT0Uxsxg/Nf53gbbcLR+XMVDjsqGIhS6yq89me
a/AqCKd2lsQhtijyxdmu3TYZNNzA/sVapaI4U1YbP1I8QBQv5G0/J5KSeGl1vN+K
TLrYbogI1/EXN7H2twJZ3Anu65eCxsH7tRtqZFTiU9fUn+ED6WHEn63X6xZUaQ11
Sp35Dc6gQuMrHYelvk6QnprPgHaTMUjCtDeGNTFi3bedA58GMA24qLAd4lU2culi
1K4/yAIZLBt7sDRq6RxAt1U5HM12E7N58B0R55wi87b7nXOqHqNfoLd8W/U4HbS0
Wvb8osuVo58yw3ujpWWCPsW5ttlJuZE9l3t3kRhC4kQ8DV63VqVIQIPbXB//X+su
Htz72HpgQEV3k1Ir5ygEv6kT2KkCALgUQl+jS2HqpwhkcYN7Q+mFJloGUgYIAyM6
ZsDgtKfr8bSw+eZ09jf2qFmiwBHVIYfFr+hpkKlDw2y0Hg6+SZCBvWNuf37L5ztP
UmtMJT7uy5Ju/r9vqIVN4AyD+iGcPSeIynU749HewBL0frIKklNM7nd27TuVb4So
WltGMMFNWcGGjMz/YBYxTwWLRFGKTiwxAKGXmFD2543MbIzLjG9PsTObMF/um3c9
tH6F+6JtuNf99SjwzJNYkn9TtxQfrWzO5oajUP8AigCRNLBU4wrw1gyKQw7fnEuO
QmmXO1B5piHVEl1lIyqN4GfaZynUOSdiZ072KKk4EMVUwqR+l7uxRLNe9QUvVJtP
EucuVfVDVIuwjRmUY48s7CCjKguLi/uewnnK1uvHxr2S5bz6JjbATyMqKKcZi3lt
6UiDOLw1wTB1wst7NICzgC9vT0nNnUAm0e7JnwANEgVBqzkKb8txqduPFCVWyg03
hz+Qk9Ww9eiQAMX+MOSrdAbi5DZxYZgk109yFA+2Ut/0e5Q2tv75s6Rs3fTfZp0F
32kzY5gTyYpAiv28/WS2LIn6xu7JW1pfeMYandl8cxdYoqSy7uNWrtSUkjJRSnTn
BRT+irSP+pXQHhQeW4ELKoTjvy5RKPLV8Frw+ww87R+lN5ZMeHItOZ7Se5pyeTGp
fFvgMwFl9gktpQ8zhuphBG90vDqzr18oQPN3sFWlIHbGeHRBefuDW7ZeNsRtBJvc
NZnjI7tuiSR389qeI00rfnmWYefzUnlTI7lkjoJnCh1y8ciGXPEm+BQpIFJivlIP
j64eKRzcoxgMHIqAXVIH0lchKfdQUwT7bajQXOTCx0fodpafFOFiNLERDqFPLA8O
gfn7HxS8DAmGRH1WRx0SBWsDRonjgosIgnbV5NsJXAIG+dayVj1C0jVdCAspUBlK
/1TsGJwEOulskIpybBvtxs10kkW7RmtFVA5WlLoCgkdfFoE8aducFrGKFcvGIbM7
2Gmw/CTjF/uA2Hw2hcDlXZ2sTwReB/DMvzBSQ4QxzEGItPrujhwLLlgBEN7HKycj
0THTq7cvymkrnMvHgyOIay0XQ16RSKx0rdi/y74CWdaBaDFRI2IbgcDqKM+vis0j
cQrZypso5C1UiF6FnPtxRd32aL85tcI1wxwX4lDQqFLIl+i/E0FQGpnjZEHE+9kM
B+rBln1MS6y/eXK6ECE9H1zQxxFvMPIzdmXgBCoq6N3Y/GgNvFAeoUXSFV9GBQHz
qMe7wyDO16oB4rEA8ySY6lD8WuhgRE8nwd7Htpg+6fueQccsTTJCZbf2BTCiDajW
AzUOX19wbqgezAQi6HmtqxKYs/ArkZ+/EB5qCuFii8h2cL1F+nae27+c1he8jnfZ
5qEOnNZBVHa8iDVdKmg5mpfIlczjU3E2Io/NgqVQbAzJuwveWxZYbS4LeNs8jL+g
anJLQZUiSv07RKbt3T4xSBSjVyUV2FhwO244/m1niPXGn6kn8MBaTNpB8D7irQlp
m+o7otqtoIIdETKxhPO5FW96PwoliNXiZ8dxBtEqEfSQnE6+BePASYsuDI7FmmEO
FvPl94dW7lznTwUoRUZGnr6FJqTci8Da5nO/uE0UlzwVpiN8RHdkGdHoX/lCdb1Q
Ud7a91vpgPgh74jKnH35oCUixliuKEBdbcITR2k6PvsC2nqJWg7b/hIR/t2CBzeK
Tgl4915WhTltm/QjKM0CbvUQW318MOooOknestzel9xvCdYfw06jb19JKyfyoiY9
fQiuNCZ4ymqOFBErXdOd6Zyikq/OwzaoA4/Bk9ir9MCUY0lJq2j7gZV0ZwdgI3Nf
PvkNRNxKOz3rRGzwm5CerQ27Qr/u7bHB5X1pM0O6HX7yZRF0qEC0Y1gaPf6ZuuPR
MoP1j7+PXdXQjRyt5qiGOxoCPnQFr85vabRtTb5WrMvXoXRIfv53U0AgjixQ8h1a
CSLPrvhszc/Xwv4NkU0bAzxz5EXNeDt29ASK1mbn5WVJPsYztwMGsG0cNv4NcIuE
byLFsD8Gs57lNnafQvEMMoQCLdyhqb8JwxaxBwn1QHgNNYIpelBV3AZzY73mcd6M
IYqLeygYMiWZTXAFhAIdWjCJn9NWQD1TQvNHWWfDeJD9zfm+t/z9f0bX2jE1BM+m
57LDHxu5NHzyruxiYtOd+gqeM/Zy5nyKhvq8IhLYM5LE7TDH7rC18PAwJ71AYNjp
gDkVwBcBuh6R/3wEgch3oL0f6A3BuQh1WEKq28YZiFyqkDj8xOiZZ7nz/5z31Jxb
1o7mZmY9aOpACV2cWZZ9OF2LmnEJjnNtVCvI9Fzqpz8x3rml9V6CafFy4Lcp3TD8
Sklrbn/iq/2tyQ4BukmDMC6VQTyYEmNv2UvVpQT/0LL0zKINyu7PDi0m2pP+uVDz
Od9AfSsNyfj6xaM4aoH1J16XFM94GW0TZep6jgACyuaYymrs79xMj9Zz7u7TrHgr
wrHp1RI6tw7NUyLFwkxi4WDCR8az0v6pR5ePXijvlrmDub7WipcPZaeRa2m52XrQ
ocllsx26akTrNEA1ilUs1/iZmT444vxJKJSxXtdM/M1+13C2+n2QSbvcS7xrfKSe
CxPYFrGB1vGyUOw7XsNEeuwhpJs4Mofc0YPQHtpAzNmrwjWus0sGViZbiyY2arT2
Xa/cxUSjnRtbJht4fJbR5GpWW7zzWKVRwqF4MVZ0BXqRRTFc5m3dyr5s2n8m8WuM
85GpHMdD8mWZdePA69cHsPm88R4OflFrkFNP2m2RptcZQiI9mJCI2RsIbXcy38I1
+A0HJpmWcAM2OuzlArYt13BCobuonwTiUPS0nI5r7ktMGdYuXlgPJyJ4wuylVWbB
/aRPFMDj5OvOXvj4/NIzc+S6LU0HibdMGz0z4F0FuYQ0MqufXWUrjX6C+VMb7pp8
o3or5ZFm+yXOAhlZlBekTNVyjOIZA2selzpuwMZKejrMDkkXzzstNwYQi8Wh9xLd
3SdIHZ9Oli0Q3dDNktoZ7F0ifrTU2+RC0C63QaEgUnvBOIOijuJmEsyL5uzLeo0O
H9O4xUKHDur7bedqrzZMNt875YXzffC93scugfunBCBNSKCjp2FE0JAookn3Uvyj
pEbmd/ghnu++Q8CW2gYJU0+OMjo5Vat7M6yP+gkRsxALBGktjmE73KAzyQs6qY0d
jMAlUKk8wjy8zCPs5kzZlBu02nJ7fmlvkLAiwX3g3O4nRnftyXdxvS5Os7PVcCOJ
VFCDI8+11QRbgsr/1ex6YvFhwqNUIIvV3veDjoGZM04Bgbb7hutAo9TNavL5U6zH
ioYTienpe8lZ6z8ErsZclwDdtczzlK+OzkhJktM4iYaIaiWoZ3UsJg7DPswAhB2v
n2UMFn67gIyYJyiyZ5MKmi++mQuvEsL1nIAm2ai1AXlByEuxbYL/b6BUa7nhkU/E
QZQA1DbYje4oDn6o3ZRy0BocjXk1XJuzx2S6HL5lkDJXnqbnL+KUXMzcPAslPkY/
7APIqJZ8vzrF9kATBcu0Jv8+TLRM8k3rxvp14NyspggRins2j/VaNt0R6sALu8IF
y4uYjRWTyzVQi4qMgg+MFmOHP1vAhshG87kxN1UMXXVzE3sQHe8/ZkMcCrKqODed
duhAAOsxB+18qomECFxD0ynxG9WSf65uBiD9nxjGEfS70ZpsvG1pOrD+F+NDk5R1
R4/3XMhPVB8X3q08kqQi7Gp1qQy158a5SOCutW79keDHpxXGHZnbM6g7EbI0AK0f
EvoGzHgkkxxlQ5Rh4FZvvtzJzFWGZzLDwFUOjxPV3Ei/V7mAtBkyhpZ9b6kRUBrI
2nOHxpddwbpj9DirsgLX3RO+c6lfwFv9NB5t0qWPNkIdIOLfQ3ZY3eDz9urwXcs9
PdmZq3oAnoZwE0IVK3sZovb2Fl5i8g3T0Y1HAaP9HtTLBRZao37nhJrdzs+6qJhg
30IeiLAe1eKV1pe5Jaajsy3NcQVm0cRzwalzbQhVzoPxnMjK+GShi4rkI0CBwFoT
TOuKnIO7YlDFlLwe1yMGNlhE9Vl2dcowTIm000nU0iYPpYRVSaxN/5Ho8/RE2uTX
dto/dar89o13IKGNxN06cRgQ8txi+RsQ2va5L3Rbthifb1JL8Wb2Kwklx4Jr63G1
roUiWSiol+rbXxyBANmDTbhsGPodrm9R15CtxarEyP7vbvZp9lkn9fqCTHW0uNJB
LHCpTqzjNmfct0OGQ3u5fe03GQha9geka7f2gvSxsoRx/1X5mVqiTQT/BGTkUrZU
T7GNqANay5ZcnorJ3XtbQScrjEBgAWcp4ey8Xm8qDqkqiY80eXmGKw4NRZESZLgf
MAiFARHzqCNy4L4MEpi0Wp2hVz8hmWeCAXGlbqobER/zOPmD7RV6zcvjqKUIP3FL
Id37XgmXlp8KN+qG0XD4b5W5b4SxJl1FtIL4oRzgAbrCzwCxiznIijSE5cNjRZAm
gilqwWnEI+ItvCQmFkhf/YgBBLk3ZzpJn3bplqzW153fzybtTaobyp5urX5z1CJQ
9DHcPJpwbHu/vuVFRJWHzDh/Ll0qB8dN2hHkxNZsW/sy0VBZAbWILA6c5yJdyeDS
zSULiJk1V05O2bl2jBuk2OMQ1uKOo74GHicc5zU7x+qaeyrjL8/ZpVCgMvCbRMFg
MG9d4RXxmXBgw/Y2itX/i6G1RdfxU4Y48TwqZcL665X71tBD9EV1IljcjvOZMz1f
D7ABeQfWun0xSZanCxwjUB0gjlTMacDp2XJsHzIfPp2GXelurv0b3IujdxAjfYKt
ml9SlgPfKQN+mbde28Pucr0bON4gXHZ8ZslmHF1jJbd/vUqLIDKNhMpLxuktTqsU
kCaVV/2lQ3hMAAQu2VfUpTRzlZ8UVRJtdd8dGqNeEVj7my/0237IXpQZbLs16t4t
RzA73MggtLbMmsqzbz7cPhBgZMzPz7P5+5ROWrVwANEgPFf10coqWNrtGQneFIuC
x7bqjcuwffABDOR6MShW/cFt6iaT/IGs6ulq/LJvPt3srMmwC9H82HbGMWoHPVFW
bD1GkKWvaIjdCTnKF0QHvdGPeU3pJ+lfoev8K9qUGIjImIp4CUSqeAVidVc0PcZN
zTz/UbvfpRt6V77kO0t5fzqozFJMPlGZS6Lmsrni797vKQDd2AHTxnC95bmUFG2T
7N0Iq4CzlqCnASBQuK8zu6/6gtz6BRTcs1av+xqCQQziWqTlMPcjN9w1qb4IK9aB
tLbpRRJiW7FaHddVARGdAXe8URVhbQpXp4J4XnfGhCis+8Be9C+VSklprUN5Iqt0
e1ThNdpDMkQQHP7y/hT7K7N/cBc3OlFmCr/f9J9YChKbI886dKuE50d5RzzlE83n
SVHyhin2uFMswBqwv+Zsc1w8z/kUWSGe3NsPhHOnfnYLXkE+kac2oXg9tpByq9Hy
iYzgLnQNTgSag6v0hq2C14WjEwAfye24mBKErA4zSOOKtsRctogvpr+If+cMZkGU
uP+yv74H9G/EwUxbK5x0I1eXKWsngoUD8XlVHUX0ALl2GLlAj8EfPkKNW/UAbPNZ
Cjnziik0adAbL9S3Zs0HSMhg9a2xovRb+cM0kwbVbqpQhcpW5p6TeYGPxZU7QcZr
uzrvQi5wOty45rHjb8u4nZ4X8z5zikqX5PhiXKinevQhpiyRZmg7AGXqbGiR9j4y
5dW4tZp+7vFt3vTZX7hg55DDTEfjL2IKlmBLfzJ++lNxPD/B364zlIo6YMAExlZw
H1T6UU8mjQgAvNkxeSB81+MZ2boCvPHC5tQGXKMKKUHndPwOwBCbKHB7TSq93lpt
HUaNaTDBhIGohD1HS9D1+70mkK4ZXwNwmOOXAkHOPICvcDPOPUkNKz+yCTapO1xE
NK0VzTcBA7sbTA3M/SeGEfqABJfQLHnRj3u6M47EFIByuZfQEYIq3H1a0+J3C+zU
1ViXemdULYAvtlzk5XbfOkCw6wG6oDwKPVbijvDe2YvsvydLd0fX1oG8eUdfrnU5
sUxFWOBG0J9mEC3d6xeVX1Jd+OobxDtn+hi2H0MYqAK2oELo/JIna/LnCIoY4cXk
nm/M1DLtXnoEKQgkIecGBfDxeDLXL++vDOZyxRWnCp6+n0EKp6BVVJkc1DXkOiIa
v5mIas8azgHVaIyQcL9yhgaAcUO6Qq9+X/TVZHpzR5FGFV6Ip/HJjxopETMpy+Ol
vT+ocPFYYPRnjO5c/zCVHTBrGXyuvrip/ZwSJUpCJUzySdDpQjv1rjzF4sFa9KKT
D2K1/ehpwBdkMyArZvOKJz43OPKuzjXva+a3HTeyGtaW0BwaRoQKH2bgoP5Qwq5Z
5aOmQO/aiSxxA4J5zpK0t7RNiNKrBK04XEqqrzWsregb2uEe3/HrQYZOv8Gkg+cC
PQx6behcsUoZORfVi9ox/e1pRqcvmAoswqQ7Lenl2Z6JRHpoqQgXLtY6BTtpAEj8
VtTZiWsjk3lz/3tZ6knqD0bioYH6ytFVbKws1LNBsZAsKDLUetAF7/84sg984HR9
JlSt8+OSOtzwVujMCI0SxA6HNg1akhxMtx2FvECPlu56EtijhQLQig7du9wD3VEO
G1SSwcZVSgj5rdVt6NkpJAaUMM7fIcc7kwRhR/Tu2u6QVijSPNBfSeGGarWroSGD
Kv86oocUNVWpJLtyOWus3MKU841prLjMviY0hEtQN1aNvjyn4W/1u98MEXMUkPdX
uYgPEnNZVDlYascgYa5l9v97P7tY0WPrp7nqmT0FL8AiF5Q0533n+MWQvrePbnKY
r2ScEAqMAjuRif3WHnpZrt+Cg2LE42AU6a0kU7xOIngTf/cKxdJL74mQdWtbScJQ
TrMZBqeaBCRjezs5LwQamQks3+PbTaoOwBA4d+DsS5/8yzPLQhjWUSsUD3GJZdFa
+2yLqWY/8hB9dMnIUQZdvO+Vwgn5CVzS8aueBhsboOvBIFeojFE2bnG05qv1r8pY
oofizaa1Edyn0YdRiJ03FLjL+Hq+ilZ00YzyG0MUFMH3fLW+E2yuqfE29U+j+3cF
9k5y2K4t9cCm53SEdQWJKhZ+/pc8TanIKW2DwzQdDywp5MLOD90MyQwJvIYY74i1
HmtS9MwtdCTcQZLWoMQdsVcAaGW3RfJlw/ogKBXkBCO7Tirw3AuFtrRjKDchV8Vs
WtyjNEgBV0u9kRTTgx7rflIdIjM/dxCGqFPQP/IK2VP5pyMNG/61ioavpV1NdLon
I4HW2CLjTGpSbxC+svrUpKu7cm9zyvAfYEvwCYimWE4/y1DV/A/720zOinc7KT/M
j//urd1Qo74yNxSUjs2XqE3dAGPCNp6VcY3YORo6wyBdwGRFlEnXd1M7AK5GGyhP
gN5FU9nREOSsA2D/h3ycOP6n2RxNM96MDINYfms5JlOrnb5WYvNXWQCFANVNqBjp
+lmPglz4JzMx2+lOqp3Q0WcWAC5Jz3GI/VUj2XsLa9f1S2XtvIy788yoGU4Ps2nC
B0eMBHyx7eakCgIKG8ibeKUHyrGIPC7DzckJOLPIEJKytSuNc7urCrtw2wbBUBEq
zop6nPRsdxhXHhJzj70DY0awtkGm+jb5Sn970j/EL+ovSx9fPwK+olcW/2fsWaY1
LEPRu1S+R1VZc8jPf2NrAiuOCIGrPAIJTDbbvbLRWNGwxcZQXVPifOb3D07YjLHL
8ozcVnhcx8x3BL9JTvPA+wax98GjCVbuykBaKdM4Jp9dRAq8C8LUUFKP94nlhBD2
QelIy6W8X5HnCZHCHK65tAtCpshMHUQKHqBU1EdfrkHWSgEeR3RIQiMrr4H0ctPW
0vScZ47mgATFsp9hd6pI4WXRBkYrnzYiYfTdAL8KEEtpVRwm+vEPCrwsLkvKwYYY
nZ7jxxGNkhxTbRjzLuWFOjbBJHhTMV1jzjKIsrnzq/GTnciYeFp9zWi3i7NiS+P1
npBOEu7h7fKt5QmcaTIeZIHP4Ss6p/Iq5F7i2BBwR7/w9BKuqFiKvCgxoR9uYFEO
AT8mlvOOGrbJUdWT/zcLUQAOxYPuiSNW/bIUlt4gm0yEDxnkyMnZMxl2c8Z12DOG
tsE0YQrzvavb8UdgFnxpRSyzvsnBbMm3kkLK7KWPpSLhNNM7Lpw3Gu+0UKAp8OJ4
82jlVJJVuQ70V5nbltKIaq9+dataDD0zLmHJ/aBtNRidl8Dkk9xisDM7K1SnrDWC
A2BDcGOeqgvdETVChoawvqvS1fLTnCMpaIgKI/GiLlUNWAaisiFwZUIjbdiIRN99
EaMSl4zsg/DoKudgphhp9uRPEcjIWwt+V0q7/b9WV4jJrAjCs4RbPRr6kbq2tQBw
m3pjrtMMr4KM0mIFhlDPBboItX2JyUGV+EqIPUTUIuWfEuBNd5h8yPc7hFrH3c2E
nRONSkq4uuvVAZpspIY1CX5SWt3BL8FcQ9F2ERQs3KReCClris4qrdvQGvhWO+ab
o/mX8l1u4g2O+HTIeAVeRcSQAHftPaANunVrrh98F3nB28s+jQXwUzDRYsSdGlki
JkaH59x/ZCQkrxZ1/2npgDuNh1PWlAHsJfn4qzIN4HKdKUBiPYVsKv7d7MT1L/z/
BGPPRpTZPwgZPIHMep/rD0SDuJiTVW3Q3glU1s99cuGwFyPGBbH5BT+RH10zq94g
iDWKbz2pRUvf/k6apBhDGDMqzlxgwcJ0X6zo2+Bvvfp3I/v1ZEYz5Tcm5V1G2Bsd
tE7ioEeADupUaqQLZMfaXJxBQ4JNfNUrXPbaDMVONP3yVRMdDIcos0hLZhz7hBTl
jGZNbVI5VB+Y+MTJ36DfJynN9RI2XxInIz6R5er+KfGh04QZ19J0hnvom2O7aDj+
nYITq+9k8M3QiJs6PvDSRP8j3IrDshZ14nvPJi/t2V3w58XARJqjhj9T1xUk76zv
lxusbnimqFsrO2r4Cvn6ryn+0lwYFneV5V0e+5xMU3kskDL5tHs/LU/Z8i14zhzW
1h8wCq3z9VtAy1yDdFzDfPNSHDUYa8WzmzWjnQDIcAZFeuIEO99ZS1yeLPY7hyuH
TIIagftuUTQ351fcc0QukSzJJH1A7nw/ilB4EHtCdLw3hRhXAET10UZ3YfunN5z0
0eiPtRjBqNP6FQRGi5+HTGNI4i/Z5GAJIPstoDVdVkCc6GkeSf1WmQqVZ6Vg2Ung
h8bo0P8vfSwLlKRNJpCkw9G1sDw9sGaPqQjS1fzjSGTRa2aVQ+4K09Gr/R0/KU7V
IPb5NerX6UpbWvzVINUpPnwwnVmikFHnpj940kiTa9PEFVaATxprpNARw9imiz59
Tp8+gmi53q/3J72ge3s2heDFsmF9CrzS9QzpU+8Cr6itMjOaeBbWQcXAOYoi0qD3
kV6ZtKsAccK0mQwl84o0WxO/2zZLgcv/GNDYuFOw9IMZR+Bies8WIqP+04L0GaZA
5msIWi3DmbRCncFQQSRvXtF4+WY6x8hZSk7qcpqvBqg6jCOggMHmFAzgrfClfCLi
8IXA4Jw/+PAGJKQEJ7qH/05aBwW1NBocryjBU+6CJKARsqwzsgYZ92upF/ZKu5C4
Jbl8ILpCSZoi6+T0rhs76/MqyknsreF89RcYgaeztKYvd9jAMuoiunjkiQ8smk7y
uSDFF378EFc6mSOrOQ7QweNDkMsPixB0eJH5XihRKiFrKVfK/RRwTvbVyRjJCx25
9rdnTx/PjDit6mNWgv0g3fG+rBOjJpJ6V8s/kNLqtUAS3ywri4xUQSXDxRtCCLBz
qeGSN5d6rlZrKqOAUcz51HWfhsmoAcErXSLymvRVeNgTHrVzM2DQXKwLy271bObr
ks4rEfds/qKWjlDI+daoz0J+ht9BI2X60nu2e0So23MC8ccurcgzKZIVeB93lCdL
FP6N/l3SCjjbceTPG4+qufdCZhCZF7pQM7medOYeNG+mdFMqe4fBIcV56Sg5ztFc
PNajhLx00m7CnfkaLZa5cqFScfO7RI6F6ruBHD+Kqs0zE4doujc4sqh9cPFWQDK+
eMWcoZ4ESXgRjeBnJHrrA+sn8+wVKQ8bq+STu1twqfn4Rk3VqsS08Uu+ZxzykOBv
sOHoBcIqhEiZKI452tY6xdQ90AAJhrt/nLXEkbV07I88SjpcBhI4oRMdCqwVQWiH
K6L3mHj9rue+I7fNZimKwpy61J+Y2OM6CzKMJCsQMqon8cDb1PbBfxjDIJGhZcem
hFdsRbYR4efpO6bSAKaW5PyhN0yOHmLnpaGSmiIsIRbqfkdAFTFunMOV24eWUZ/7
dpBOLxyvCD5+4cD9L2o4DOTe3rRFRBN+kJahpcOS8glMu9ignp2yXguv53HzpoF5
gLqoOAnSjBqV5kCMZM2qV75WBb8IGiTvDLMp8zoKmKHNMTiQWxByOUSzsSBopwoM
OFSStvwSANrg/dbP/0NAYgeAbPZw6KWaJm0cnTenu9oNg0fI/G1ZD+HAw6DRiFzo
rjVd8IWUR0T7RyiHqT718uwkoy9F7bixQpLrad3SHyE9Y+QHqmsDlOzJJm3XLtFf
LJ7wEtUmEU4X6Z+cZE8TQX2io0X/D585gZQFAxR3vk1Ce90oZyNqdm9NY9pxYQCP
YDolPpgZbc0RXwPKZy9PYySdiSraJJRALclgxUFcpuGoq7V0YDb1krsg96VVOq67
bgEGdW08pr/KvEct4fqgOLgnNWC574U6Jj3BFDSZdurScNpHQZoyngKfFoE49B+X
fVlZDwvuvKkePVWtNvk/7zfrYGaiVSQzjzF776FJRgfFeqVzdXmW/2slRw3f4GPW
zq1xQwqAWUhgqj1VzX18FOYvNtKZ9kOhx59ljzUKVrFeUeN7Mz446dSr46jH0ozR
ut2cqMaVNfkcLsc0B7CH+uNBQSiUl6BupCTBP6cVq0+mMnbClMpHeLkdZiLTWetS
IHBWW20OV/pZf5DUAp2RJz6UE+l33dbnSUGWHFUqqO520n3ANnv8PdDdJFCwJzrX
nV4q3UFeI3z8/oP1KMEfl9BnFHOi0xLir4TRWxOZnvxmJIutBcu6v7gNbjLcs8vM
xIE1HpgPminnPk8z0Gq8UCfSMkYpOObDlfbtl7ydmAWxDM0YwTJ+fk7mI/DKuNMo
sPmzEQWZL2oI7pdzBL2hiIwPSPeB6gTduJe/Wb+EZw3tUXmg2AlqBtpy1Q12efcF
J1AjevdzTYzhrpXBI/zRjaIu0d2HGyTcd3fTJ0B1u9Z47NY7njEf1t9nRR1PFE7+
9nFp6Rhk8yF1XcNosVzZhTY387zWRbkk7LoCuoBt6lalSa3W/hiOmzuI2nf7P0Qk
cbT2uKJr0Qe32zVZIu5pa+se2HXSX4/mPjEgpIJRSm82R+Wf6icWbH1T/NUJIMvd
TkxSp+a4F52GNzCChS1OkcecP1pXvFTUZH0i9nYUDhnhY2HhRw8mS7mp8MHjze2d
YjAiNLLKfGuhy4GTd6DTHHHF9BhZA7YWwlKl3xnY/I6h8YuP9uhyKnTISKUjdYzz
l4j+IYUI9B1E7AJ5/9ozghVmrpij1XthiqvGzXhJcSOXgepGiRh4w02rvoPELhDg
+hDu608rAhwbMdISclU1g8ccWiGQ6NFsRH5oBWN2XxbA7GZ/xYTUhJ0Yz3nYkzUU
DTc3lKO6itk1AP7IsHgdFy0+HYdvLKGdnIXAx2ltCgUh3J7k39y5eTzLQ7eBewWp
qsmzdR0bCVmDINho1nHhsU1bhL8bNfVEFVpuIs00CGO7eoFysFsHBawuHVxplJdj
aUa0K1OPawFC38PAG+mLwFVbwbf5eMr81U4KNAWSOvRrt1bRkuMqMvoFTaRcKCCo
F++QpUTfrirYczRmO1UGrmGPwUBNcHwhMiUTaBrDD1XdXY7DMcA9uKwQp535A4V3
tQ7eOIYyN4qBgyPFMOutVLyLtRcoTxZF5g6wcxjw3ZTFd2gFnP9AgWFI92YBUVPT
xzA+o6+D5752bqc+FohCtKpiNgdxkkIMhLYikd/IjymbNjBFDMBz+WV3tMaXV/3x
E4/FH8qoscNPTpYzcXsY8Q3fi5BRCe2HldCEAkCYVg5AuCM5sS/y48ldsVfIpxCz
ec6uhztZPM07h+jcrIFuFFYLaSEZQAuguAcvg2Cfi/fJTbF245izIahjpW312jgm
iPnFxIFI07lQ4Npn7okr7D7Qlpf8o8u6P0oG1tc2KKBMzI+A1zpwRSKQ2Kt8jtNm
OuIq3aKBf/glwUbFuLtlNfgQWt3JisMvvNLBZaeIqqWlidKhYzN1swr3/UwVeDxS
KG1VSYE//24N0TiyzaZINM9Sc+uwjgRi+GLMwaG3iqj9VLpCjKivZOdJBkGIVjAW
Auw2kTSbfCcpnqmKI8Un/FXpK8LHQMMDbCKuEhSyWEc7/kpUzfEdj8iPK3xRMLYA
lzFjcwbGbfRFrqMRv6h7mB1WjSHz81W/GuXp3OqjHrjfeR3P3AMXXBwzONnvPnus
wEDZayHzROh38eAJdBL9D6tE4xFvUCUTALjyEqXa/CK2aGXfx+5cJenP3efJWicY
Loqawrdr7UWSxEac2w2Z3n6FmtHvb4eGUWlx2dmu/c+DZ28ePOrXAqpN145DdiN8
V1DebUDhruReDjUjiZQHp7FHgTwiIDJRZWHO7l5UdFtX7Utmz9NHCsBsJlvFVZ2C
d07hJ8w8/nK0FPjogvqaOymSjjLPImg/Rv5LbhNOridv0O79hzGtiWj6etK6Du5y
CvpESa6HoiPQc8VufvF2MPSzgQ9oHUS3LPnV9p6zJiswLGOnRit+bIahQsngCm1E
5D7dkZMv8NP6d26dap00ldzL6eMne9Hwc1kIaVMr1Jai+amuEhwvGI2WxNLTVPfk
5zPDpBkhDrs+hD5V9sndZ7+iV/hAYO39m/+5ABUzuD4KgcthmTuVca76vGUXv5tW
P+l+VD2dwWwYN/Tf86opY5mMt2E5tjkcQpjejqH82odQAt5jgb7G0X3dWK7IdHmX
+9gRtBZ6j6onA4p/8v6efFO32hZtdi6ts8rSl+BzR+rBAH4Pb4dtFCyiGxBW37Sq
prNJ1eAuS+O64pe3WXyCnlHtBHfhZN64Pte0zUfpWgraURuM3VCIqS5wI63ezf+e
JZJDbNk8LkdZcNvuYaQTR+PUNagdrMkBPDLDLEMFisf4O8NQpQlQKaQLBE31PrFy
DjniYd7zCHqmLOviMbKlZ8aMgSSZGlLmTtZk+GZE1d6ycDJQC9AhvITBJ+Qulmr5
43tPP2bB+PtHzqFpmiMBZysdlOcs+rgJzTZpdd7ruuYh4uI2MnxVwzEnrvSE+Dac
DS8CMWofcGkvfcTJ7EL7l02XccGi5rQUwx/+lPaILciyR5YgWPx32wNLKr3KeXSM
pXoOuV9jN5ADhNVYNtWdNky/xOA1v2kxwbn5QVZ4bt9esbvc3BnU62gcEb872kxO
svVdp7XkPoI7Apfu1LNopeZCoNkxIf3I0EyQiScEXGOxCESeVX2kWYhSGo/nWnxl
WZHjP7cj6eCi2s1Y6lgwhzXcs+BYqnlX6SwksFGjMU0kxhS//ts4FmPlWS5JR86u
ptzRTh2ih04tfLTz8x9/ANzMTKxr3ixdy8DT7ab4nFU5jFjsh+475Ee6JSyj8/X/
z3tM0S3Nqimnp5EFSg8bJcThS0TVpU0kQ0A0wvBN8qPybWHy92xO4ZNfchjmHKLH
2F5uLhkZCYPQcfCh0On76iMc8bHFsyVs94RpWJyUoyXkmfhMs/XPnFyC+X7KepuJ
aqLSwfbhFFbuMEVKfdfOdcBkCKCX3Qu9kp5UbklAW2PZTgInyk0+aYq4nlESzQM7
sE1rwxIQKz+3k/mS7+TzkipyXd1iTU4+d+lmIgF9+z61oUIOqB5OCYLjbcBpgseF
tRm1frPsR7UjxOZZY9aEfXYzMRmaW1q8+Bc2rN13OmNc/Mom4D2UYidT47NuxcEO
KujLkHLSqpYlVwYxOCB1s/faHhEMt80kzeET8hGyNhqmlv2uTIpCdYERIV7ovAVb
uYe36ysMWbKVBaXJueBf2Byo06G73qm13ckBhvx42tsvAuDa1+VivwMpLO8X8N8D
LeGgC8n9YwMeuNSX7iwDkIV67WBV7YX6ldJxDd/yg5jpiVYNMn1rqhH9InPbuJfW
9bWEV1owJNentckbKQsq7UNMI5QXg+CldFfQbf1Y5uV5hHy9V0HZf86gv7FE10I9
z/Bb+qlKhQyE6Ges8Aoedj7larlNXhqNsTJqg1p288Or0AdcnEujqTMRZggR/rF4
caxBUy0d5MQ+aY16YugG6QQf7TpJGdS12xNCotRtG58ObrXcN1RPY8/1p1eKMqUm
hWjldwKUBJoge0XisPvoxM4we/0bGAd9LJzFXEZqPlDlefoYXIsrQWtG5DqtTQOL
qx8qn4DHwoE2PBJ8Y6OSSuwkVSGhG51FACN+tGsFvTp+UeK5cp3NbuchvkjVfYTt
7+YrV1BfBAi1mvaR6gifNEr4QswY2K/XZ3VwDo6xyHoRNvrxcwPY3Cz/V1ELmPB+
g/P82G6mIWw75UJsd4TYYZNjlWXzlWYwaZTrHMamxjfHLd1RfsFiLLiIjC9lAdMX
7M7f1bVhW9dnW42iJ+yIvPAyZ4dn4O64TzckFMmwArD53mCQUM8beXahO5fQRyA6
l30bQjbefZomJZbz/PZrsRdu0hBeqEaLgDkym57/D+MmXJK3BjbtSbgxIVhJaCeO
DaaOWJOdACIpGG/LQLqmZjM/oIQsLh3WvAI9sZIFnoOOICRgzysk7o2IA1VzP7qt
abG2FbnW15cugYhjfRGO9tT4NfIMKSw/XVnmiQPrP8QDLoLa1n6tiT2X3U8ykuqx
am7sQzyea+1RfW9hiwe/Jb6RhM370jPDYnyBkphYXh/RkO9O95qXf/IKZNLID4eA
mRjeVq1tR9oWIrc4dlVB+C3W+HWwOIbXThiMqbMUY5fr+MFxCoAVf/aaiN69mJkk
1CwO1nT3YKk7p4LWY6jJLC5q+3v2Nmh6ZAPWvsyATCdjKeUlkzP5QOEOhk8l51+F
8vnFF3DA5NDlOko7S4X+s8qd/dmtu8JZ4teNjY9eOAgc4T895Xz2U1z6Bd27SHJF
PAo7J1Y9dstdu8+q4EEWK/tNJBJQbGgVwaJrkuqHzyd+ex81IDShur7AjqMTitna
5yyPVfG/gT6e1tOGQxEJPGrJotIC3vgVS0xLIOEu520/15hxRa4EM11fIjgQHPic
sSguNIHifULaELuJ62j5uOFynYTt+gH1qpBM4a1ahWy+UngOU1GYPZL/kgOXb0K5
v1asYZjoL0u/zI2UAkworcZKtU0rhhiItTyWeFo8+ofVnLZyORTcIDVxC+xq9ty9
d0MFl/ap7Y8S0BoIufA7Gq6yOetsxKo67LPZ32/Jn/pxK7A4iwMfhXKSpDsYXE3h
cBacLTD27oVPPFJW7XnylECxUHFsc9ziOpFVjF73KlrUMI/pMYMU6pFS1zqSowVZ
h4MFmlMjtlGvIcC8Ia0jAm1urAuyYoq5MdHb67xP1iKcl6nJaHUznTVjWfVyvNnJ
TB0HU50XAHjUbEG90DJtWwhSpXRBRbEP0WeKJjpffQtrKFZXF/uiG6Hm2Db0nHsj
BnvOPKOFOd/XhlLQn36nBCE4dSup05nJ6pe6X4LU6lPeXDh83j58GyZ/oFOjJC+k
cWpQ9TyJ9IoRWqeibNKw4DONhscN/P93R5g6wKn9QXnQGIRAkvsrZ9VXcjk4RRYe
PTgTtpx7KPhYQoDk3vVl+f326QnZmOyjAVhzwGyn69l6kCh4Xyo900SARqPupfM0
nwcRx03mWtalfsE//9uJ6ueXg79sg+68U+cF8AbrPV5XIH7hghdsrFjILF0J3vN4
UPKaxR/jIJwm5nb33eTZ7ejlrdt8WrCxM2NcywhNif7VZbP3lt225n6UDcw8B/ji
03GNz8MxiSu/7yLzXpDkIOzk7hB9/dAxA5+KJbBTHNxamDSvNReLX4xMjzmDUnOm
5XAKyU7DCg/IzXLm/z72qEi8CRMIawetXz8EX4mM0pTMha7uwe0AcWxnWm18uCc/
0WnycNbNFgI3qDxuWKlDoOV0RyMT4ws2x1YuSM3GQ71HDGOvTel5vrkW3Hflk6WU
zshJsQPdQ+I7sTcN95J8ESABmYW3jPhh2SiSnkGvPDBOj/5U6PmsbBh/tNr7+eMo
SjkOb8gcXx2Qfzm0GtGxY1h5s5AJE6txze4JUaIF7+l1XjbPaLtYc24akKokSADq
7eBiMZVETHQebh96h0AlO82+wLlWL+lWfHhDP9/aEzcx7qkqAL6FZCiYN4A2fAcg
+4wNAYVbrhiLk5ArrogW+0+wZqeXvYHcjh923eii5q5iF4Z1rjS7dt72jgiXaAxV
yiGK7hnOHed4dqLE3B9aoXkArZ7MYEGI3MWxSG7DSVxuIwKqE+48Ko3l+qsuNLKG
mIzi417fjKR4HKBoV4fe0avumzZnskTnngLv6cuREXkE0I6nZr/q3voR9hemLJek
csMaA9KTiRQu8DFBOgQo9xQSXIP5c57GX9gNe5HSJ9JfM1uzBhxrA5QYBbIW6dPs
oCk7/XcJvoqtIfLD4A4Qf1nfuUKEsI7rlix2e0ZCS0UxfqV6QUWE0QMw33FM36LN
T4nsjDNwkq1tHjF/44f3HsrkKnPzcR2cfNuAtbCF4yXkRFBEa+1vYwipIu21UqpQ
HgG7WpJWj/M7jyqEKfbmh+JY8FCQRO9m+B7Kd62CntbJnB1tGMINMmkcktmI7Ow3
rCIxnhSDzHNUUMDYWLL9hjJBde6gRquI6fGc2PAHS5Z9sjheypJJYF/IbmUMs83X
aHGjdeWDSFVf47EdHWW9NMfK3cPgX41/PCdKwVH8nC6EMuxBxw36gjKhZNFrmBtQ
Wp7Th2hsEujZQ7WNtpvnblDtw8bSIbIosmmpG7e5j3agOrNDsd77cg5HvNbg4ouN
pYREOuYKa4PMXqDeoueJj1/42XFNffMKX4MarVavQBb6r1JdiIbtOPv4FKMdyuoC
nCgnC+aFInCreM3Ndz0bsue4G+0KYLtSGpK6c2816IEDIN5sGx2BwEjUOUTT616/
GezrQpMHuNpSt9lpxG95a1Jw1c1KLb7uGUqU/dvms8W/goIA5L8gYhmlHRBt/d8q
dqtkka1Zg1kD76J0tmt5fa3qptnsK80kKRV67s6617f3QOSLtbzS3+rpLtABg+4U
Kc3svRTxA5G1WnXJ02lwVf4nb0ErDOb6dRmYyqCuXTxCo4P10EFbM/BDMiSmUT3F
txlpq8o3+mhBK5fngRf9wAjkrScW6w5Tnvj1howkKC698iIfbkj0jc+fnFiRNSSY
N5hmuHBX+Rw65s+Cg/p1vOuItookgK6+bw/meyOkDP0Rs7ZOfV4ZjN81jpV2iR+0
HtnLDUN3Efu57SEf+Bk2svMFUTExtL+joH/603hZ/KYm4VDvj69Lk5ffwENMcTxu
c0OUSBcMVWyq4MxzQ5M1W65JrD39QjhIfPPv8s8Dxz7hURwbML/sXLiBjvauS60H
IQeWw9N4EGsU/TxWP9TbWXF3e/+qShSPTBW4wSMTffTSDLLLgBlRuLBUba4QOxn9
yabhb7b9OO1SkR3IQWSgvP/vIWTmx42tSpdLOdHjv65LqmxNNJAGEcELZU1WDdtu
h2h4O5BbJVnaKnr1SudI0548yTIFkeoDMEOHNQkcUyHd/0RGwxr7Pxp3XmGt6Hpp
6Tdd6JUN7JwzsNlc++n5iixjZEB6iLUwau8thIqjGKsuzz9Kcsr9HVG4InoyqscO
iHKCtIEvD+f8uVBPUWaqakP6xzBdyBbrZL22iVdt67QZ83xotOzufdphRgyOBcPa
pjCkcbQVwZGEymXma//HLZYfWGldMJSYkJ1SgJF0iKrgMssnN8Sxl45N4CbYeYS6
vN4TTM2sAEY+bKxQRvE3PWdpFTcjmM3ppbJuVzJ7V5J0+ynG4Q1r6ga7fK/RdbeQ
2/ZNHH1qkN3q7kwMZNYgkgYuuY86GeS2ecBd65sDxMNA/c6sSlABV1N3MUIh7jsY
i+q3u7U1mXWDi2LxwdDq2HB6ymvN/qjNqWknnAxkgZDxPMQHOV/Ri6EovWHhRIMV
T13rhFg6C+P7gRzi+5b4tLHvj5fPvGPkf+coz/DX3OvEKedd24EiRjN48ioagFem
J8K/A7fVXx+4ctojEWS5OmmxfClEgu3+rsrH1be0lJU75lU6hII9qmREdmMNcCDi
xCjlFDO2v8q6nGob5ErXU4Zl2ne62La3lQP7WdV1l4l1g+lLuFtDJfgrnop1m9h6
7LVEzCLksSE8b5jwqmO4iHircr+JOa8ua8PH7E55oszXt3STHZJV2ufTTxudcdyC
GgVZty4R+Wy6VoCUESxU7Tg/Xyntg26/xQWbHz225sjbNaCxV1n7BwP+ANNqFZJy
xn49UmNbMLNKoDTvA3hGtFOHc29McexYaGrhyTBzi8ZTFWRyvfmDA4WTmeiDccoF
AI49XpbknWihRih/LUn5uI0TAZoPK41qSS4QHu8eE0FKQdh7XAwGMxQJruPmTkOp
p9+wHRfI9mw8cmlUZ23tQuD+BHDuOvCR81k4KJv+0qSmY2/0H5PqroSgpcW681Oo
hSPh256GWK63YiKuAsITcQUextxyfLz27Lc++t+wPEdyoXukoFi1QvBnlV0fyNah
PRDmyzsb8bgtQ7kNaNFBuOAAn517jWDeo3TLBY/vWeWu+GL5AxhSZIrTx/JfOtEY
v4awclMhYxMnI2E+8J2jGe7KoBcKDtvD4kPF2YcQYImvLLyrqdkk3COVDES9wZv4
G7OEnCgD4ehVNmUtA/5VzmtQkCaEgxHO/y8nG2rRTB1SzxqnoTG+AXJuWazLmvD6
7RH77pcuPgEfW7Cl0aHTYbywvTkIJPQpsKbB9QfrMo7iISqjmWLq6jxVKgfbqoDj
Rp2lSFZNqBIdoWPfPhmADhVKRLwyQ6M4dJlCEqiMVE6/kxxCclqhvf6scV+/FYuP
+E8/3xN4BJnwe0WZfyF/sfcHIDFs5cNU9CatQwpHigcuKdpdQsHgWKLVJqoJDf/5
B7Jz3OR/o3RPwBqrIT+9kZyfW4wCNy2mDKjpMky1CR22w/WTM6ohQKiuXWvYJ213
x+Pv9odTKYXgh6LtlOXai7sy2txJq2lDRF+d+6CIZMZw7mMEG1Wu6BHUKwHypZGV
hYVvMW71vP0YHMxMYl+nP6ta2gQ7pkKlrP4JT4w8UihDzw6dd/JZkjZ9fBmMoCcu
Aj/isSMbfrWalmm/oRVejQnFoEEzBOSuKVlNQxBoZddPTS6+ecUGm7QxaynpUqdF
/4+iLK54f0ExSbL14CLPlAfiYIxJuj5meBSxM08rQPyBWkF0OY+gp/87o8q84GQt
RlfZX/YdlHdZcv5ZSoVwJEy0gFQmTr14akGwV1+5kpGaSTljPNOJY7kDVF42xhKQ
HHBderPNhINzLp6Q6n/+lyg0sElN2F93aXFxxqRzueTFYy7JspboHuzPykRc1rkc
VKoRDpAmfVS/W9ZiqFFaF4mcgeH0tYyN97e8Uc0jImn6uftxZ3LLrUBMVWmNiZ5W
HFTJ5Rl9gixuDzIX5vfh3qGedGflZTYBPjpEfxFLshYyXiqPTFqoXdeSSxJ1zu6U
bgPalfvBC+hMeqGX+2Jb9wKJ+wtXR0HDl9cyv3Lwec4+w7eiY5o1dTj/9oxXIybT
AHCslq/xzXkAHRLkqtPAHFUDfTloq0WjUvfqr58+cdhZVNpYiSfyhSXS0keODoZH
rbLNA16WQgqkAE3IuvGh0JJk1Yp/1Me000cGkEvFwgredF8CMmi25ExzsS5OKCaj
k2rPla7A6TG71JvHl6gvwfAbCu8EUYDliHR+j+Jx0S0rr4osCwx/MqpXBE20b0os
J+KxwWCCS9j6tDAgKLUuM2j/paxGZxiQmbgzZ0zWeXpuJ4qm5mUs+L41Nm9mMkrK
iBjfq8M+iZGfkXKDdWNYrt8aCp3z0UwqObMufx6yduI33IyGsx+m6vdII55XhDPq
xAY6XC4QTSDLF3PIJsQrgp5pVFyox8gQsUXsIpHT+asAady0NOLxU/1tj+MteT5f
b+z1LPCXV14iyDk0UUM5FpGnAj/go0KPkcb70vA45pUCmcYhvyAUDxUT+VB0eIPL
2+CuNCBBMNtmIG30T7B3faQxrmfT0vZXs+29jj8mQNiumGzA9rdiqycIzqdOYH8S
aqfm+/oQvITJ/Q8inaxquKSIMnxbXVRRaf3qIiK2qegePHm5ePcmbWxsbnQQ5kBY
POZdiO/5Mpfmvi/gTOaxyR9BAuFP/mP1YBPCc30U1DS1BaWd5IfeAx0dEua8OOVn
aUDWTHiZZIRTYHEcDK0fHxyzFYyVCx+j/EofE7uIgQQPuXsxLUMqOoOuxezwOYA6
Y7CXOmxQW2GWradZb1QWVZIw7TfR1Is7rxwZKG84CAevTrHsnhfEDE1cmujW38fm
mZ89SnrsrN4ehYgFiD1RnV50Qpxb4Co6Sau8PTlA4AvmKwYjQ80uQzw1gLLtpLIn
C5ijgYJkgs+dB6VfgFjAilxTpfDTC+4kQu9RZGflJYFkI8HFHYAi7susy5Mk/dL+
n/GlafNX9MfIVQLwhSLd/8FTISR1zGCuzxpJqvy380aY6CnqPLsg+A11KRocoxUu
FEzOF5DB8EwEmmN3/JyQUo0Q0LIhVXyLw4NL0SCCYruCVq5s2AJzw+iwBYMeq7bc
b8xpfSH4ble/kDx+ukWg1tZMBfkDufOnxq15rkOIWXHEXT7OSdaSBQSV46gAbCSK
1qxJY9n5tCYd6hDqy28UGeYU6ZNd3EWWXvT3DdJ+GNGfsCxtk1CRxou8rKEzl2RL
KaY3EX34qUSiqnuNl9cZi9UaQLUsq9/KoPCoCRhu9O/xZZTZPaHD/k5aryVGCmXe
P8woTTP7CPHe/dLssuOf7xJul1V3Tog7DVYDx3pOpTDPF2OtLxOb/wiWJRFxAB+y
JZGbpk7F1Z+vS0WXK+RRs7PZC75e2jDD1qdxhNmKIKc8orkYaG1wGOSr/K5Uh/+d
F9BFlUd9x7VloIbgrE4JjkIJQ9kTMfIbcfloO5L64psGyL+6bPD2dNgqSID9sgaw
GI2+f/KDgAUOUcJNwzaNFtf+8qPYCDnouRZLoGiLCUfbRmmZfHSRpdSY3TePtdI8
vlqm47u8zHLQoHLHzw8WjSUyA3jdGCUL1UnY+MoteQlNGZsp5caoBDmnPsnkuaq+
K/6iz06Ol/Fo1awPHmOyb8hz29t9g242RwzWSOm6/+UjMCQoPpWnd3HwrMoKUOID
QNQPor93B7pasJkYgVSZWRhh7IJTwCSNJm8Ec+nAuAwqtFGvoeueouvDosNPIdWA
gNX6rs4NoqBaNvS3XuyjN/v2w0ChmO3GPQv9f+OptSYaCkCL4pyiHPogj+IFzr1y
bKPZAF3sneeH7o5rDQgumKQKm1OgwLWLEP8iFKA5h+FHgGsDp0myR1wRwI9k+aXa
/4WibxNcaOijgGQ/NhZqCT0cXZC5ko8uJV5xiUvcS88nxNBhvuGjoz0po1f0gij5
jac0G1IitsSeyLqeXgs1Tz7GEmNg+CYjMHu+NIroe+ITtsX7ebbWtwEv6iRHKIIm
eSqTK13YMWobesuG4WspSt9tK8mZuToF/xT+r1XTTJERpXzpIAytYqsfnqDxHAOs
vkqlLMpfNSsO3pBwQaOmbOT2A1zvkPBEXNYK/iBEN+m8eKpTQNvwaK7WIv+FGM8V
gRK1hNmfBEaMw0WmIQnwSyb7Bukk5paSFeRh8pk/4iqL6ipPQvUBS+vtxnPzmw08
QLxoRVQ75Y/2wlhhWH3+dViSSQ/e5TBuWjieXZgsFcdeJtAXqaEu7uPcXAImjNMB
n0RpI9l+6q/QLGE++yJknWe6Tp84/204GmhUuQtTPQlHQYdglDo93S9kYhvf344e
lN7P5OrtPoyTBnb9q5y8fl52CpxYcU3cesFh5O5E1iFVQHRkL2/r1cyCnQGLzkhs
jeloXpSePC7Hpl+ueQE8UyeQJlJAjFtZPBRx5o/MqUJp40/vKKo8DNTCA3S6IT8E
Sle5amHqKMy0NiqqvAwQrLzQP7z9GRc6KB9V0evXr3JMonMa41DTJBU5XqMKRiZ5
dlJGv2S+MdNDxUzH79XTPsca86mTpokWkZDV3UvN8f8KUlVlEUhQg/7pp2SEZtg5
rUOgUpcoY1rnxohbxD3x6qmeHviVdS7oOZW13hmuEl0jyXPLPJ0xYzE9CFmU9/Mr
K+qvGhFDDLSEOExaVjV6PIjoI0mFOe6LyjuxCA3V84MdG7iQ8OmKUeQQ8OAXLeRQ
OlNcWlVrafv9JpROLwrNBxqtc48zHh2vIs2icT+iG/HFt9JgS35s+2RGMVwNoMN1
M7rctvgSVzomPXvIEYaUGyHv9K6Ty6H4szVbrmGu8pAcGQNJfqOcCMebH5Yfn2EA
LtnAaOQNRG+q5x71KIQ3knhKo4CnHxP+7yVE6gf3STgoTWSP5Aud/ToAtyVplu02
R/o2cAfU/dbi30guMjek7oivBd4GKKnoRGsRZp0IYf89aQWlgY0oZgqioxRoqOOq
AK9KEZ3cPtje+7D7I6Mn9eTmOsNKILFC+Vet/sSLCf2ew0TlLMYzKckUz4/QcTht
OHCj21zoHqGcYpBfD/i43OU+/DOJlLHTFVkp2ard0edFxrRB78x8fhknLfR6ZcZB
aE/YWUbgvIw3JkR2mvCI4lidm/K3znmXi+CeqMOWhmf3ighYNHi9QhC61WR6OQJf
wx4IOVN70EqrFbIU5FJsvPYHzbKar7b8GpeWDkvfjx+7KFTFq70EfO8HdXxFyaUc
CwBWPbruEr72gLZJzNQDcP+d6mKeBclZhfTAz+0uQRSZeh2LT0XoSdlOl8+avYKF
5IRZ5A7xMZ1GWBls7q0cPXBVzsmRsLoE6xkGmBj3JTEtYar7aTZw4I7G/dyJ1hD8
2YupspHRu2NW9iW3+rlu/B0c7ZTW/+aUmOHFz2n1PqWSuL74jDfbBbkZQhpQJ778
H4dyH1jOPTScGOToWxPu9MnBW2GaLnBrl4LDd2Z8rnNiY+gRJ6RItUJbQkAEwKdP
6Fq7nKXHBoRpURfSPXOVL1p1diWH7F2DbmLWdZ+wg5e++qS0zF2TCEiflBzpEG0t
BMMloMR5YEhovbRiEI9PCraVa/12rj/lwDlX05SF0L8BUPfiztaFb1VbYQdW/7Q+
0UJyb+U5aESQEJOgWi8Na9ShbxDowuThNthTM8jtgaqSOfU9tvMMAFTFNASFMUPb
iNFO8YfR5YZOiKvVIOc1A3lyBhZJ4aBItN/4hm1SjwEyIVKuiuqKUSWpeioYgVxM
6x66wvBafj21q87JBhdBDM0SjCwQ7mNiYqKQt+83QdFpyss75BQ7m6HrFJMwluTw
uCu2eDjZHbd35ZMSzYfLiAegf4/gFzIfXYO2aeHuHZsCf9pj0rrJwnvHufqAx1sk
FMbM+QtxF6gwIBvPKIQrMCL+3yKWY46LbN3HYThPt1pdz5uVqSFX7M1tgeGO/4jX
wwDv7Jiqn0v4rVcN1NDVN53fwZT2U2rAV8WeAnDME0XHr1gfHBCiSsgxiLlOxcd1
Hus/DVSP+SXxkkXctsh0KkZ9C2YFMTYoRs6za70wWhMcn62nrS990d392hohIvbK
D9ydqGcxEWXkWwiuxWn4UIrf23ve5+lKAFrz/rJiRrRWI1Th3uedDJ2aMdBSF9fH
3rCJrEnmzVSM7NE/IOaiztdquKncKGYhgHu4WYzxSHKO+PCmGwItmtdQylDSmM12
h37uSPAsmIpqY8hTMqPStbHfJ1SFlC98oDsmaA9//fO44o40JxPveoKFQRtSE5vS
N8iNqe30zg+8T/6Kf3KlfjsJZaXQkh/9GPZpymnJcy9iVIfncg7MPDEQXvezQ4ct
ZPvEbVO5QuRqq3F3LAAENMOn4Z3nrdwrKw5sCT7bhfMwJSxyUuFhsmteTkMBqJQf
PJGTBjOZgu7Pw7+KkCEVldeJnipZbcKKFtagaDIADJZqHNG6qvZ9bD7jg3rvFDi9
dditdPBDeq82uVjDWFPOypxKwkDMVDHO8hOSRI71r/1PIcBYOFMF0O6nQ7kJfp4Z
4pnziTOmLzfeLee5MfdAJxZuZogeEhspxAUW/PhE4xoF5MIFlwlT9I1FDsiQWgnz
q/YOGmWkO8XFxO/f5TEvxBReZBdLlrRqEu8b9yw55t1VdIdwxQ/3qmUc51dwIYqw
5KeYtezKOdPMyh8pDD0hMoUMc2PaLMvMDuwpg5EArdAZfGaAOYpBAJ3Qiov9hDkQ
5/hBXhGoRvLy8t2Gyt+GDefm/qVanxucwtyrRF/L4JG5Hi+1fqT9zgtJppc3g++f
HVZP4xt6nd3L97sR25XI3+WzHwaKNUiEv+3a2bcqKmXrK5yf5WfLInICvf8kJG1J
tT1s0BTujEMWUuVJdsPH1XYfZgO8FkLSRSWUOJOzkxRO5XewSwF5IxiKEe1QvFuE
H8jcdqJ/pAgMTqNbY3Aj069xm2OobibDqsLbc4NxL3dSzxocaDHx9k3qWh18pJAo
t/w2CB0Izfzgy62ChFvI7kGglxm9Y7VRcoxShsF6bJ4lgCKRsORipK767fNVbnK0
sH6Gr2HVtoUlwuPwJwpFFSPOXY3y8oKIkBNaq+0Tl03LmAxIJLqpbTetmWW37l1q
CPqaTi9mDfzY/pL9qhXWNV+tC1R6eInRRKKH0GgTDknqCesFJJFgxbBBv2OYygdh
0Ay9OzB+OUo653WoB/jxxsLGQlluSfgDJj2gxN8RuUpqMm3HvwRXRllAsb6s4pYr
8lzEe/yd1yI/sLn9e6zo9G+Er+2l9LkVbkTbIa+klG2HrKHyh22CiIE4jo3nLd69
fmFI03qrpTg+c9ZKnZirDJne3iLACXnuRw5UEUNSmNCFLqwjLw8kAQUpS7W7/S73
UnUd4TCkHp4s6UJk7PqclM8INOMDp+UL8fb0VIfZj20vL/gq9feTvWmoiT6+kb+Y
YxHAlV6NFno8Qq9RAqCkkbHmofWUGJ1QNORG7Zz+QcvT6LEv80mSx1nwVksagZG/
17FWoxU7GmRf2AgWpbNFMMmInw8EREINcuXW/qcJMxLIXfxQxYh4YBxPHLNCfBaX
CM5XQHi57BE2jYq9OeU3naO8AqW+o8Ug3S6VF5zFZ6zBP15VpcniD6W2pOHkBqkm
nfNzw5rEoe/fkPPe1OTrRwd8KmlrHnFrD2vRNZ17n/yefw7bWRQM+Tr0q+V7LPck
MZjawm/W1qYwe2SJr98nddvIhKpBk6jDofUjrMSEq4dxGdap7cXX0HEN/ObLzRYe
OuOVxfkCtWuX87FIrqyYNjBo0a63ktzAMbu7LX2q1QSbtRzLaDKhdOviUHm0fbF1
Ki7x+dEOIaRetZiuUXjUNrqDSxWlYGVZsLYkawJFp/pHHOMUJen1VtUH9uw2ijoY
hIdnpeOhEhJ1men27GMqqedLhiCGllvjOODzUfUZv1ia1WJ7k/M74Ie2rzsPNcPW
IZbfG+991KzC9wRysCP0pSueioUbjVaZIh6Wiiuy1AbOP4CmcxRuk6ThzmtpKbl5
GYGQSCCjXZZLnC6liVjMTeKi3hntJiTmuN3w+HgXv3W5I72s+0IB5MSKgB16c0Rb
VaDiiTiG7dnqL5BI/2lu0t9auGOyZxQ5yIxjkO/R/QNGcaeoNxKPSGBVAjpLLnlN
QErNieVs/d4Mz3WN0ksAzZEwMMkMUq2EIWL1nD9XEzhHbV/tw/5lNr/Rtg2zy7J/
Su3Bl7bGRbAANMc5epHNF3/GLyjaKW8pm6mDCuP2SBcpk4/3GNFlfWNWNMUQuSiT
Q7Pwh3+kStMd+tR5iMcfOqf5Dyl51m6MT63FPXEiRaIH7oB3JR4YXO2dHAfHBrYF
mZLlrkpFHxLjIxQ5zQs6VA2SHs9l/+U786JhcEAU3xUzP1qvxaM2OjjnOMmTV4Fm
og2rDHndv7/Bs+9LkV7lPA38KCGXNrqP1nlv5aGh3IMJryObfwoGzBlNy7IjjW6a
EmPT41FyFtFJMXGOVvfjHVGznEIGuA3iGww5eqwpEqh5Uvt1X5Dmx0mLfDJKaOKL
sSf5WxBN5ISnXe3rw3hGoqjbcLlrDZ7wVFToXF6OtKllmMy4P3xMy7zS3u1gbqkB
BKlO6d4PWiWyQoZqIuGIRj3khoNp3liJmXaBQ+SPRCq65oPDEv7SVGbLQb9xVAZD
yYDkh8T/rGLDhINSoe3M12C+j6nHDZVRQdGDwwDLZidcYLeF+m1CzyPQS3F86CuW
unbezyOKHIHLiJlPUWCghhSwZcms54U7R4XhynBIoDDTHfABIiuOust+v9K8K0cj
Ye8GHQxKUNBIJIYhl7dfyw8kFKeTXlFu0p9gePvsMaHdkNcY62xDaRzzfPSvg0bU
XkXhz8kH+PwrohKsqC3RWLUMUeqLbaBvjoiWcmOEXbbgr3l43iNsDbuekh1dzRu8
l+QHm5h+hHu4bUAwyx5eOrunmAeeG4q5yrGeEi/VFFr+a0AApzojeTIycerjb+bn
BrrVfx189cH3s34gzhkrXYTcaDBaJf42u3/bVd/OlRYaoC0wWozFfcbfwaOqA2wW
5URZk61zwWsGwCMjegzJHdaSjxknMwxnnebwoHmpyLxV1t0YZXw66o1/olvFAmcv
B0+bTF0TjMl75z+UzJBwXawZ+dkwNDkakYi0gXPyAALNwAL/dqLjgEo4OYM9ceJO
pyLdgjItELpvKB16kZ9sIBNXBlCfWmjE1rDVGhlYzmyOns3jPlwqpa5jP/fOm/nI
ctQKUu9cASeOXwRiR2waH3L7I+c5BWqlilHiqHV/u2lcS/ClSQfIStGh4iBP6BTs
pYUZTPOpnT5vNifio+9B4QADI9aKsRsgBTBQ3GzMShl/RvFzDGLFS8NGd6ekS2cE
eba6/Hb6NVZww4Fv/OC/6yCDED/YWp70+u+jGHvQksJktW5LBIbervJv8U3ryMkO
aw+NnDKhLYftBM0GKMueQKbasubJOcN8iEIiOT4c3/DoQAwP7A2hv9MliOD287AH
iiD3i/IXpj8yRFaZrygMP98ka7SrpbsWh0WB8xs4b2W9Hu8Tkc2RGnQCKxLMEII2
utpxWKLHh2fT/ZSrVhjCXjcU2+HJkZ9Buqfp6sq7746bAc/iwFmhZcdA3IrFGcY4
BlCnfSCGwG9F/IUSce/h4+teDxCV+g62jQYKhj8P0LytwMESNhJCEoHCM63TD5Lw
0i0TZWh3ueN2PiDAHkpyC6f8Y4qTtk5Q7iplh2iVIImd9Zi+yvl8IZo1ABBPW4J1
anuG7yVoJdOS+dpooGXKAqbSc1m4IDLWHqCS6YPq6goazFYhRjZGPhJfDykFiAVn
OlLx4d1gbaNfTQTeqjhy73CFt7GjSLIUizBjXYkfb/fABqNotWHcGa+oHf8VsHpw
edwHHttBk8668M3IzWITmiPjHMqYz/WxGHeb7Rvtq3JBvyTvbxmxZojlUbfcLHDb
BQ+PLWBogxAPpt/VwhyvvD8vAoCvziVX3DErGY/kOTl3RdzElHSBTDP/Z7Ibbn//
TyRS735F4vUaEKkHxR2PZ4bSnkkjdghlrjd/YZfGvXGhHdNCVkQD66Y4tEtWSHzm
1Ehmf2OuEAFlZW2xS1sUcZGlYZi+L11Z05fzEQU1/ttVsKyLWu7I4vu6JmjImQC6
H0Do9z4keerG+IsCKVbDAsE76YVlpQgb2VdEu3tohFiQuhW4X96n2GNRhhGCrIqn
4qF2M7QIetlGvAAET5gGBjutEYILAXP1naGHQ2dE32zi+CtV28sGcddUh7krv3Gn
SKmNyPRPJBINrjpOCwQ4JSjUiIbAIGwTNUeQ3hcARFJTpPgCIO4HdMJLNllM9tbF
UO/qP7RzHls7SC1mjJw+Q+xoakwBla5xDgZ7pulLL/YEqNs/w1lCd15XJaL/X8fv
1b1+CdSfj6GnXpl4YbI32Q6y8BGs818pVYheVOdM/DZGhWmg1OkndP/g/OVBFAZO
6L98SU6+cZzqLNukC7t1t6UZEzKsau1rT7S6I9VjHYKvcN4nw4YGLUEraUHyrnI4
8Cx5tWoRBdqx+vULOCS51xA3id4TvVxeu2sIGe0jeISBe6tMQXCeb/95iUNm8Z85
viAy3bdNm1JwPGemTIihQzU/3z0XXchlxjR7xng43ztAsEpiJ9IYimLDmgshdSnd
wDrKH2lTz+mTLX5fqRtEOQvuxvipqNIjxaOpbSIdry7L7jxE6e6dlp4s7D7A51R1
fBxMKMyb85inHdVBPAkBdT5TNwXcIorrtAiREY2xp4AG4Hv/07gVcHEZqF7XK9LR
tp3hfW23+iq60KXpVznNI5+eycr4zek9prgb3DveEgbKkcl6C9UNg1ACa1LKsSbo
Zg0yXa70j+YsA2vByqYwNceHyXi9DSJAtQK+FGRT9EEzjFkuVCilIWlPBLit2Qw4
1L0oEp0Ysn9iKfXinoccG3qVJnW96IxN6O+B0FKYxpTLdcqVI/s8eD6LDhklQ58M
PsAkBKsbG20xt9VAHuw33jYB+MF6e/PZJ9P9ROI4t5QSA3e8KrC2u7/qP93InmBC
51dmg8mWceTV2b9pNiTPeaTInUJ4C2wHRpynDPL0VvMnoYfIP60GKq/JFDO5Jnyu
tAL1dn2Dz+TKmzmMsgEdoRqKhbysJflpJ7KQnrHbo8QAl38iKRjQMtwAzr2aSe28
gBNROpWaoCj491S6/shpd7Et6EDZdL96uxPB1/FDqF9xqQa1N/9bPaWBBUqZihtv
xrmjKSG/5iOERoYgXE5yn263vmvzQICUXmW5/S/xui81AkG7vv54TePAPRrSnyA5
GmBUEI2lPCEfT+2uR2EShepjtAzxjc8GwSFHllWnPBknnLffK8bj53W92vzCekG3
a0Rt2aIxS6dQLi6Umx6VcghaGprYerJJGbxJrXF8LoGu+o5jgoo85tPjVk0LVHqQ
kwztIg/cMvKWDfndAulVkCkIdY/7oG79f4ZEJTjHQcq9wEYPm0fXWg5sq4xoOB4O
O3v32BjsRWXoCNITAIl7OEIiTfmpB0tid1HpAkkIg96RHuNXZxChxL/x0CIwLW3K
eFrXENdUOzD3ibDYCZ3Foljdj99C55mvsspjhW2t93+VFw/+jVsOX0EjARZfznG2
tFwM2DgliVHijye8rX67bIege9QLwK0GkqPdAzWnt/6WdKsMd+xwi4POQcLs+TgY
AGlXxYB1QDzItUQWFidi8gEhmjktQDc7J7YKn7FB6rDMhGL977gjcC0u8D4BEjKL
h/hGdJ659Y+lgWXHaEPR0WSwgP3ldXr4n82lvqgAOI3y9DnaRXdetXG2Dh9jef6N
y5QRbaaTrhhvk49+Q/kLkZ7BUlHeG0GFffGypd66J8MGFiw3LqwJDPCnMzmzuv5V
Tf8r1HRmQtJIWR3xkWG46jKGRjxy40LqXlrCJwUj0BcRKUYzCg/qENXq9Ii6Xpvn
5Tl6dm4AMuheYFqHWSEzrruAfLxLrHeQ/vBqEYQt/+C6M3HlgUP/TAeRadhU0WiO
tkpmfqQY83661H5AT5RfWZde1JeIUmhe8XHafPavI02DlzU+tSyX3gHjTM8l/uPo
WgVO9Pv3ZMoAUzbLMrLCY/5Zbqrzy7wAtMq+/H6zG4n8aZk+quUMA7z88mhX53Fz
96dd4r+kJh1QSYXEhxVx2v5XSHITt7Y+sDMpXu0NCPacMAueJYc/UX15ewO78FiC
tTUTjnd6KBF4rypMSKGyaO9i8cqwOnoc5svEQhj1Fd7CasEj7ouEtwpnqyD8E4lc
5RtHFuixi2Pau9n7tc95F2bDE9zbJQD0vpM8JLrtdL1/960UVqm4Ulq/l5cIJTGx
rITJYozCDcgbXKYWVPNHtAnJZ7mdi0XjsHXwY6pSLiDhZ7dmptDm2FscilFZIyyJ
3Z2j6fU45AizE4WhJXRVQMqMzX7/wUPO2ST2xrqdXSqJIXj6wNxGH6plpcrWUyAe
NwGh9LiXo1P7SAc4cSph7YVAErhFPYKHhKkez5iGPJHe59bbu+KPmrwrFEztKDRk
2xiUi9Vx9JBDc0i325KUHFcCCAyzi8siVtQ53IhU6n+r+zi/8pvu4AtQwMO54AGX
kptokPipEFBosx9hO+hIp1RxkJvWBl54DjJYAyeB3Hu6hRec2BXKmHrpdXD+Hkcd
8pNgaKMwqnaoiIVyQLBJW8vkRdpoNaPx7EEGpCsWqq+IhevkEWd5rvxi1ixdNivl
xtlHyHmTF4u2dpj7VDFBTb/rp+d0l7mcZb1gtVQobmin+u+Kfglxhb74anSlErxK
MRnIOBPmtyzx+lwOoxFFsDe8vcNEW3UdTVnQJtMNR/dvN9EA4mEzcpZFYTJhsgig
VjROatgLgGBNHK8ZQ7WyH/F1W9FaYVqkqh/FHxfSJFi4pmxxpZKTNfRfqHBHyU4F
Z3qwpZCD1LcVnjX9cZ6MzkKG4p+kYgdQffoza9yNjYr+8reUvwYJwtmxUJYF6DfL
IkZQFpBZjpS2ZKRCjyXiW4VsYHrdFgzYpoOHMqjKRKB69VRY33G+5e2TvNJMLOz6
bNQ1LoPIBX3+9Sl80C4Y3yknAUP7MfbdHXL023YV/NUh+tqcBGSHjMvp0dVBGrj5
DrPigBRXTPZa7S+AdvdtKkmGBd4XYE/Bfc4S2qKHU24as6SEoZ76wUs0v/uOBWWA
o8+zixyJmS/jccv//EQH8ixBJWJOiaBzXmQ5RRMqxX2MgQPmmnnLlAOqJ3rdlpgx
vJIuN310crLlAYxkzztl5ISWfTYvIvjyO8CKLr+qGsg56Q0BYtGuesX1eMDK9hG+
c1gPFaXP56bAt6Qm4UCPjU0PgFAn60gxzAJMIfdOrRlVDHk0UskGG/ZiZodH9A4t
fYp26GB0UbLTwdFBR3zcgNbD0oX4FVZKtMVCWMvOSKjUPOZ+ddSNugHYzZPy+hh/
R2bMD4E5WPlQ1XnyQ7P/FWsnUXUtfV7/875WnVoR1vEy/N5A2XKi4WKShqFu6O0f
PSzXspzgdcBF5mQsWi97XtkcHfz75+fOQSk/9IrtKAJsFHIKOqYOawaKbplPTqBE
KqBSB2I/p/GrJdqGqSFaaXTSOMoNNCNMSXctgsireuAGTr+0G9Iasmjaxl7/CqV2
TDQ/xaNtxT940qzIHGLsx2vprBsLn35Re55IEjQCMjYW2FiZIsbkkyYduVeybrbr
Fzvn0Ndn3ihbRQfacMrJBc/QD0g545gxiF4hj4zWG/WtYjSrE8YgGB7p0dWvZvK/
d+PVHQ/gXBV2b/HVwFgokQfsizdsUr/MyKaLqC3dqYzb+bvLtBwAx/bjew5s82C5
o+4yqIYY10gyldpDqKJelY99QwgD8QIfoyGOZuvNN/g4H+sVEy9GqvERw/CfAWsJ
5DWRtwSwpIC7jwL7jDldM0naGB7wN+PCddAweYErRx64s/36dwoHBXjztSN2or9f
NvjPr7pCQ4b4EvTYTBwBgUPxzM5DKp3kDsM5aIaEO921rH0kFT84AvVt85NSymfY
PjIzr72bgfokaZinEpXwDFvs0+Gs70wV6qOBfCu4ViFFz+3/0PRWsieSroVgQ3Q7
WOmFqdYDPzaKMhJQnGb31o0+9F076jfkUyn0p3zchEHxsLD1yc7DoURmMaMbG0W+
kt43VVUL4RuWqWYaHQ/6ey3SROSONvIJJ/WSGdPd8Oj26Hp8PrrdaWMGB6ZEHODY
4Ws3BHeizPcEnfDKCGBchWjovJiWfBLZvh9b6aEYxjKUQwcJIvsld9Uh+I3JecwT
tPcXVx6ABSJMt4eHVlVwhRISf8MSqgQi4QPzyFvvxxeGDWOC1K2tAp80zLLzoW9h
wQTKGZ0j2wDs6ilw7ggydp6qhmktxyeu3U1wJl+HkgdpGqOe6fBOfSbmc2Eo1005
2zUT/nbthvOeB67W6QYKDA/KjllZIqvsmtFM9xpANIjxzNC5YWzg8jECr88Ic4yR
ByAaapVgwazpyHJ/TXAqF9khE4f8XsUMeQ2pfH/QOwXuMVsqrufKABaBp25ZyPm5
DJidIgN0EB4uoaQ9HwteyroDAJ1OBobbWau1LCqyd1cEcqsGzpa88CYiVXvHXxs5
Fpr6YTPadNBfLRCZggveqiv05WsbpHRDnVkgvnp+f76VK61CgGFUwpvkMHpPwutj
BfjmeX8r4ae3JSbANwyipEpobCxFCnUhfxsU80yO7Me/2DObEX4u7JZ55kFDtBW/
T5NGQJx1OYRA8tvcYytnSLC/YsqVyCVFIyabhvNlQhu+iJ73yzoW3zyT34/H1X2j
I4OhI/nhL0SWMR6pb3XetSW5+HVkWyYjTvcZLTXw1BT2hn6quWyvnF/nq1Rzq+6Y
EynEiU3dOqiKfTDUXYu5niBztKXFTbfIMTYXBM5vmiHjF+u3ofFP1S8RRhPu4amx
3qg2ZLFdK4E/SXj/PmLL1BsW6iZxtgW7I9ujPIM6mdwAPhH2L1frESj3bsoM+YYb
4X6M6+tvD8uZjrlwPgGJ7icCgalN7fHZoJQJBvtTykCwmKtpHAaIAXfVlB7t4Vxp
RqSG+PluZMYkbbVIuPYSfdIFT/oQsmrQ+ojllMsQw47yoJ/sHSKlkt7a+4NUxd4h
watDUMXJZVgdbZu0rhgns3oRFef/lj8h2FK+JHuJ5yNvpCyEVDUp8f4GaisSKvJD
2ggJRDUKLFxskgjchcBxqXI2rySSM59VohjhUJeIY68PmOyK1MZCJG94wzYThmli
mr2p/RdGRURhYb084eYXvFwwkg+DD159FxNK2ln/0dRZVZ9CIHRhhs0sTabaN15i
d668Yl6KbIIQ5eTv/6dj0/E0T9jxEkkoBW6kVCW3/fq2SK3k4IhlQ70E7VXGlgv1
OEnQLqutlDww7BTM1mmzWN0ZrcGRiHK7bQHxX1fcE0RdhEZsbNZENdKhoHpM2gRQ
a+zcUvK0MBAuKEejUsFP2UMRjkc8LhOyh7UieGfKKUE1fXU4FwopO03APGBtN9wm
c18EnvVkReZ7PaYSST7u1c8tL9EFvMVpeuUyGJWQpdM8u2eXACGm673rQo/AXPys
zPLDD2jOi7SaIumFPbFSBa1gh7y+O1XqB/X75ZVxA4dzMfdT7uIKWzJh9qdqI84f
vqWz6oo2FMwON7rImeuY5WsMeq5/6Kkb9s7f0MxV/639DXdK7MigmTFPLHqaGOKV
/GAaaWC+1zFZUQc7v4PECneoVskhE2uE5liF+ehISzpageAPhmEmmU+VrgOvY+iK
9GEPmI4fNd5cyLip+uopZ1gvWVzX6kitQq3iwwbEcZyE6NQ5lfZpBbZfHfgLoY6q
X8E4RLYEnl5rZ/TtVR8k2IwwbB/LMI4rJIoZE37Whpw7qAB8zwfs/4wJux+ptrd3
gEDNpAYT6k3BwDQejTLtD5zaIRpHkFYM3J+lcZ0JNiPbEJ3qkOKDfHWcZSCkXQC8
/EQ0hmA+v1EzitsrX1IwM/lzRhkmmifhpW+wGVnkbiFrAfdxiQpezP7pRuY9KcFk
8I2ofTC1ua7p6kpAIt65IxOyDdTbHdjLxxcTLOZJ4q0aJm7+hzWsfFQQcFSkkTo/
FoTXJTkLcFkJTXhT6QgLoq1rk5Yq5oos6ehyQ9XlMRjrAT4s40hdIMivpN/aZfNL
T/pDmKVuvyZikt0qcd1ejFPSJ8m4xowTwDg8p+no9JhycDrQ86kC2hsmaUVwtVtU
Q9iqB6eAlv8r5LmwYP/k8Km9n78FNj5iBjuJr0Q4QKNQUCay15CijWYa1TGeLkOW
4V0XSCwGmSAp0RlR1Z29KjGhadpZVq0WcEu3l30qPGIIQXbNhr4waXyMLgOsHRiE
7CbQ0zA26mJHHzka0b7QttO78xq0NDia6kQw1Zet7MWHeEgYCwfiJ94rBWenQ9fD
V7vh8GsyglRfgio8C2ByZW9LGJjWk468UqZrl5Mu6y3iiFxral1w9SI5GNwSqeyQ
b3vgWPKRoBpeRsamGTc198Ff5CWKZsLFL/f47imUsrLfsiBXUjpELc6BsUHH97WK
IsLFrBoAMSP++zWc2mDNCb0OMxO6XW2Hig/klzTzGfr9Bg4XupUWeSIVlURAUMCT
pZajRhwoOMFPjsz7ZWx1lbske5JSUEatu/KV4R76MARmcC+51j7pba3AuKx4iImQ
Va/QSrfWt/OC64JPHHN9h3u9w79o2RVdX4A7BOmJNPpslKTw4xbfmSTHn4xxT4SQ
Y5HwKaKuItfDuToqwbOSoA3GNEPDbdQ79KhHG+a/+epo7Jse15rN3Xm8USUzTJak
KVbKgGmD5PN6ycPYH9ysfo8vjNnxFuW/8dEhqe6YEbqQL1CnNhljfF3ztDTdzNhE
/Pn9MTi7nIodn0O6mz1qe8JIWLWfZ9hHv+bP/rPO4dHbad79TzjGUSqKcfPwQkuB
RR3d1n69sj+3bm2eKQhgszY7Jc2QZGrL6q1wD6MKHvhYoAo6vADwDl1glFrwSs9L
ZiaMYqBZ0h5Qi89HJ5+Pz3zWfFDGmrL9E3aLfG+FBLsRE8NQ354MyyAi5AW/ZZ9z
Wcx6jB1GEGagydNIvAZSbMNMVfrkE5HOt2wE5RX5gKuQ6Euc6F3WDG1i9ztTgK+z
fk+rfEf4IyhL/EbUPddf8/y3GUJw6gwVF+eY33+1+Zxia+mJMnLyRtsfCw8QSeJL
Pq/4Yt+/yV/g5Y7vFFrOhR5v+D4PhWBOar/StDZimasLXlJeuKZSDm7jYa0laRjj
zkePoVBZm095xEdQ8n6sEdAIXtxDNWQQ3a+VhN3Hyb3kJRHyYhGhEpnPSM4PUgr8
B5PUumsdcdvptvIdEqRLvhoQdBWfn652wuj4OdGRq6lPKWDUgYWvzYMbkUJdnVGX
14SfNm1/AW4hID1RrgKvH7oF+L2jkOcxJnG6YYmHbNrDKLQ7up158p4ZvyFwRFGG
ynOlqM/qRpqrzzzk3XNEG7TO1sG0rSb9YrjfxWpsRi/JiWfmbWMqrK1Ye1pgFC5I
/wZDiKGFvsscWuE8WC0MQgSyHDfwKf/wBG/Wn/sqI+CF2Ehbv03sXci6/IzwXOFt
CRO+P5nYIngMSI9OTd16vDsXl7/CDbCFTFKuXtQCDpqX/d8TzSFBsvvvU9hQB9Nl
ZlbKGYxz/DuTwUpdkwhuYLca0yABpyBwiJCzlwIjR3qWSYnQcv0eF47nFpt7+FT7
nt4ZlOGrNSCr3mtLPG7vHBWGgo4kKgZNw+CKOuC2sSdFVDRQsijwRvzhr9OXOfAY
niZJhknrpGw4QT9vNCGfDS+gIaSRBud7GH0Ckjj4D0mOvWHnptgPW9rUq5yQ0A2v
ueZHUMAbMtNmpgJADx3Ou9yJZVXFy7IZQLtFfQLVrtnaUGhbmFmYXIlbJOBGbx0q
2UQ53m0I4hnMcYO6BivEB6gBkx6pIskfNsj6OPgzqh5DnVDG/5L3PJe+U2LVtBRN
KhI5zEc582GYna2TeJ3JMchS869IPw0xfa/+PO4a4ejnMaD9+ZNMlZfVyouWigHX
2QxcOb0ijADLcUUah11Sno45a70gKAKEi8YUzStwbQ0DlTJNwKzWYNbZQvdq69Hj
GusL9z7+OPmajWHxKfDq/75Fj4yptVdoZMijXQrNTsY9ilgM5oWxnypcBjPNqFcS
FLWyySupMU1S6kNQgjKRby+5ibCR1LX2xdojuT9kNqZqXIPso57Kf5P3dbSHLJxg
wQeUzGnfxF8eMgUuD6nT2qN8ahLIf1pA8hzOKxyTE0CS5LcsR5x3pRs3nLLB10+W
ZMZRYSEAPVdfUwhcx+xghFTrmU485ygCFGzbMpww6LipGbMKOO31sYwAh0cX0fy4
CVY5Eo86X7x1GOqj3RDETHmpHxPSwm1JFVfPP4rtwNRsb06N4eJRmmOGKnlP/Fj3
i+VH/5d6bDw7/h9FpGMtXWFNHV6rXclMecienNoGloFBs6Qmf79hLLJCpYxMzlYK
wjBzdXzNBa3O7rTMkoofmU7zrF+0wJV5+ALEm9XLFQpgcMGdUfFskpG9hWU2NelT
UN7tb9bV2BU/5Ot+RF4yNHZfZaLjfvAsv6SeBaKAMIjmZHkFC4TOjHNQXIXltsuU
hL+hEroWb9lPEIg7uOgIBJPlpo8X5hbnSuIOwWUQzbk31oMsg4HguERiq215rIDz
yHY3ylNquvCetVYYipu1kRY4lOhtWetk8LtFeYrsBA1lLYUIXuXVoexge5WjlKMN
cVsmPA8o/QvmU91CsZCU/NQ+GAY+SEX7QWVBcByZCHG7o0BoWL0evIab1g9xIG58
WrD3ql2yJiHmb715JcHFG5OsLCzhsX56xUppefkIjZvA7hqgWr9Ftj+Xrp7jeKtc
d34YsFvRjbveuKGzyg3FDt0nCRSsLGnxMOryEVfEnl4nh6VgWBvTX2H7txcI30Lm
bZZsg4GAkSbM3md0rOBmGKOL4bMLvIdKCuiwTH6ZQ1+xMmbhfx0t4k8WqxijjVnk
nW7LobnicfQ0YT1jjPbeXAjFQUdnwAEtcGlpwZZF0594qG78PY2rS2kS3eVbFrFC
JIvsdHdWr06UscHGQ0Q6pzwNKG1bM6ujzjkOsZP67SFk/Sm7gEWs6GpLpywnYHSq
jLidSwrCS/n9kPo7Qpimgj/c80wGqZTM2WpTmHv+NqzOptx/ve8b/v/sYdmI/QWw
wgrNqJ+P9uwbjL5uvSXBjwuTDN1tvjk+AOULj+0Uo1yvDmYRHnLx6ZcKmsbUCkug
lk30s97zLasKwj7gKfS3whTi5pG+JfTE0DwW9La6xGe/kSIDDi5eunHnUyYIz2vF
FpjovEe4MH41B5KEKM1pD3PupIIrKnr6TY/nOHZOwZWGgPwHD/Zp7KNfWvNGX0Dm
l9buJY15p6zpNqatrNOoxvGZJ+ovgcd0pClB2sox1xfRBZ3pPSM+fTv3PEXO3zyb
vZhaGkIGg/L2r2L/s6PtDPbbCfURWIoeQAzAKqsOyLXLXn4IRDdcMIl6aTJNDJDk
cmQQU4IH4e8cc+Bo0aaLn5exteUil6mFWhodByjffz0ERwGnjYxUhBXj05LZe1Oi
0r0YooON5AFpa7LbVHaFol6mI3O/K25Fh3YMTy3kWKmtNnJrqY0xTdwtdzJDzZ8J
ZJT5BjUJuYQJJxB80K8yRfVcJ5yOdfsApEVBkal4tESF7Vac7xi4KNVHNjLNk5IO
PTQByi4SQp48FWz9udNtXACwMCjvSkl3Zius3nNupvOETmyjyDYNq7xsw/+pQW8V
ble3NRiMvwyj9ctXa8xYCQc94CA0ooWq/6fOBrCZOSsK2ICNvscsviOyEho0eV4u
i97Mi832eFFs67F1pM36kGrmGb4K/fB88SVtZg2FHaNlqxU6hYNJLt1p3vYfaasF
fVrcVPChr1eHZDWSrHKEGap/281P669otPM9bYyLRqFe+gWeP99EWGuGR3WfH8zv
fZ+/2HSrrErsQL6a9+2WOwesPvJpd6tzSumN17SEQoVtfXbk7h8RjmvApdASVA8w
zfKV58l8kG7uEinknnqskZYmv4cXShKvCkJyU5YNSOdozSi1bLXKtLfnLKmMOh8B
EHehNEXRRsgdrSqd5FdsKIgoruPh3MaZtUiBm/Igy7JpD8LSbYeXFWzLje/sZU9b
NM+ZTjMHRsfvAZQY1bVxd25TvixiRSJzomFGzaOSZXfaonw/Lr3sSGWHp5fI79US
hhlw2uDh+DQLTU4ouJ7sV4IsqVi71bMp7M3saHDGGnfw3sTjSUTAOZ+9nIT5lNlR
8cgq5FSQTDKBA027ZhfxNURQ8o/BliHXiaya/PAhoSa0nwwv7x9Lro9owU90FtR+
ZUgSGxnN7iBXSQ8vpMEa9edkOTXZmHB8eEZJGB5IEz2uU3xCFr3yusyhkxj6zl2r
0Gt48Qfq5r2JHCLP+TBdXMZe1S3AT3u8HVr4A0fiUDZwhsO453vE+GJjE5lgsL3u
Roe6P9Woyoc/S8psGzH7i+sxfqVJNSsK04aMgvj/8DdC6lMgiYEvT7IQTiB+TRWL
zziUXDpAXOfmEG6WhJN5VnFlGo9VIT5rCFqRM0sQp8279HVCFlzC74VJ+mKQjWML
Nj0cQx8us11gh5HR9bK55wtTkC3h5Y+6BrKVC3rvu1FVH296FKqzOKduIRKLoqfD
MocGkGOhgqSDyW7e0UoTX4N3ocOQ1bq/haePtJ6pJ5Hp58N0J4JT1A1Bv1gMMVam
Fl1Tdc6wCR8Hwj3kgt/du4rEGIicPFgcs2KTFy1pe2MkdaRzMZMsj1uECMXs1SvB
5tqwQ1hZbOSLCwlEZmeCDMwnNHfhG+6QmcqW05tAlwV9pbSxQcd7k5YuSM4vVMu6
hPiq3pFCKrKcvdzXOJq4JdirgyfQvgMJPsbbrcbw4CPM/xHN61c6H+CGuW4dba3P
LWI87PmgG3KuRaMjczMxRiRiXGAD0lwqGKbzfcEeDanY8HUhc/QsM7rp3Xo4z6tN
R45rDp2j/LDuH/lpnYNoi3dKJZC2SSl/hkDYvZTPqVNpw8ALOOoj1e8D9Zao+kg9
niKo7fv67JuIU+Lib8txhavpYivKBS2iTTO72j1FnulKim8F2gEsE5hKWMXsvzsw
bKVPRZhNQOZEXdvF8FZHwT9hlyH0VMDqzJvS+4tRLStvkNW9yXNfpa6moKq05ElR
FZQ1mRRSf9ij5YRrVy3BU6g5kuEZCVDBI5LLvowIr0dAJrtlihBRynoHbIoh+1U7
mBr3OHzAt46qaBJ5LgVwOGpEZAqoQtaeEX7pncQv5FbsQWdZ1DRKbOnoK/JdTKMi
9nFqsh3648dc1j7B9IfV4MRxlu4nhNsWz3xllis0JNSKp9meuMLAlhA4IO7tKLNo
5UH/cWOoRP0zq9hJwJ02PmIye7Oq8RBq1xuHjFwuX4Og1LV905B/Yb7k9XSIUpOt
zG2I5UU9pTEgbLZfmCc2LTr4xd+sF7YQ/hVU4PO3rWJTm7zbRJ4/+Orr/+gAW5FA
9m+Ie0KodXHpDOd4j1rlqu7/mdzeJg6brGHD228IiWFYISiFdZSGzGk0Sl7R6SJC
upcgqlX367dY4HML3sZVJ/MftW3/x6gOWkc5MSze0uTb8K8bER0pIqoBJ2To+M+J
CawNel9lR7+YGx5ZMMMv/lvdsGGYFzCDDGvg0lp61pj2TAhA7DwXVc45hx1caRmt
vcMt5blDZiKvGBd8oOgfvAAcp/8RVV8/dJDiEKDBV3EE90fN4jnrspt2h1f0svZ+
zUqO8ppiI54uNiDlFSnJI77Siaq/3myTLJRvW3GEY6uDfL3pkPUQsGrLmgL2GMmo
z3yBewtV1KTSF1SL7Bblj1Vq5qS28lKsrLFDJ8ZQhcw0VUdN1hefql2D44Qa00TN
985nqgr3PVNTOdc4utwzZzbfmeBH3+jD2gH1Dg72BrRNJHiSJQaSsTR8D0HBR2wE
GmMBe6xT6XRds3pOuvWVc6S+hnCPxyKcjBNoIFBdSKIr05ddoFMYYtWTf+J0NHFl
ucbLxgvhc2/brdzD5XKfDf/x3jQOXrfXQDXKwf6tgPMKWyeV9MDWyVjukWpEDkjQ
1xZJSef1oC9R3J/Vgf7lnnZ253E01H+H5IlxNxYt2crD3G7wciYJsYHNPKjdH2Om
rUP1kuWOwKBBqXEOcIDy1RQuK/QB9wnu5nVSfgqO40dUDljXW1k8ODsUF3v+BliS
13f8CaZdBTai2Bt9hyNNhW0lZgsZpW3k5KzpgwlmU5yjNkbedgTqkALXyhlKxFfw
55zVhBvJeET1yrOJL3AOvqu4ss6SxmRy7nD2G2OtPoQZv1TvyOTqpmw4ejRPwUDI
raNH2q7dCIQ8oVlZOw24NDHFYKSxvRb4DSfkApDee5/5XfymIblnBdk1I/5CopNy
E4JKSZUIoHt2geo/JtlP7z9ig/VDW9TIlFpQnoJa1W4aIqkH3D/pfAekgVDzqb5C
iyhAuYBkrkvDf0zVrq4ggChUFVUnUuRhcyu8S6VW0hMYGXQcppu3wurYFjMtBFAR
HVmMkdCG5kWVzk7FWSyjQwqSduBJfig9ba61KoiZOSVWV9zwMPwv+9hhyr9vWSry
AUtmEUiwENmb6pNZH7zu6cZouZB1t2U8D2MvDhGR8jA+WN0Vi4umBO3UG2HhzleC
bM2nm7vCqQ/la96VxhnS7SfVRefuFOv/BrFBArNEzAA0vEwjqQm83XlaMKd+eGNO
r4Dd5fcKxnNqkp9PNwPMFnxiqcRj7ZfYnW5f+lrnwt5vQRN03wjeTQQAQqinCVuE
n19DrbrD2BSZF6h9DyDulTVEE4GBBq6s2kuyT0/nhCcjpB1zt2VeMqFAnObqnKlK
3vKXTgDlbFVhHwFr+48kWV6E0JMIObf18zaYuSNhSGbPpwSPHx9eBELab9583AX9
4/wtg0/mob2YsCD2mr/thU0PyFF0YhIB6BpYpWWMJzn7pJB+mY15C3Wf20hhpwhA
paY38UjjBmBVIFQXgsmpCpodIoCV5sY8tqXBcumPRNuTHDMjvJBEqu8PzqFDSfng
WELIjzGmYOP2AmOsFZZwBK9qKXNWn7kEXMkHvV7zuLBc8KA185yM2u7lE0ga2KOB
05a8IofnsB2wyBwosDf2sVVEq3MKRimiVLTjlQzAG23eRu4qiavo7H3iqtlJDkaG
vPqXls0uZO9/WgNH7AyoBetxS0/42KryOW/Ag1xxl+OIY744IBi8wUT+OnP6I28G
+JyGGU9h4BF2N3uA0CGaCsH+NhTAKvkWsG/1SNqyAwIScRyQBeLFOx3hzDMRoqL9
PDY/TMqM1NZBu7ms8dHf032ydjqkEHQcSizZZt7H7J7evAD9vdV1VIBG1LBRkVS+
5fyurkhZewdp/AJUMUv1LXtYKkwOjO4m9wLoko7gKLLZ1N2TOnfhMXKY1x6/ZZwk
rTlNjbDqTGwNs0bXpA3RGOmuKBc1cogEUB3hb8or21qnES7HOh9DyIomBKagStDl
d6FxBIaE3PyGWIU/EDZ4zrY7j5doGAAaxs4s5JEcxZbNXnSyYEEM6UeJpOanj/+H
y0gVy4nhThSY7pq/5k15KYSIupMHbZYaVS+HJFBA3KB0bb0wdkvysAGGEo7H2N//
1MGfoj4DI6zMwHSMsD6HQLeFac3Gvv/Wk1vV1iWMwVZhnRqqLveDug8xrynKwdN9
gufdU8wTJTyvI7gaKi2F9NZIDVOURFAUwLexa1kZ2PjxQsZn15YEwwxQNZZLoIVE
qMHviwAJ4fbkpDQwK3Qngdc65WR9FnG3/KnGYgLG82TfsjNOisx1HgqWNiM/izla
n+BZh+rEnFlKa6bT+bJOEXhF9gZwKfj7gWVw71qlIiMa5XltJiEXbL1Fv05n17NB
vsVVdu82vTOoea5hSXjB/nIQ/cEqd/xGXEhmGud+NRBP64ZSBS2BVE0iloGkif4i
5NWVq3KNlcB2xYpBwf5vq9CnebTe2DVoUUImYaTvArCGFFivQOaNLbT0n8pa/0Fq
mjxKRXINrjeGxN9s5uUsyzizrQd5BtJgHZSLCQ2k1aJrzcqRLhmUCXzWP1+7DIAH
TDaPRlrv4U5oazhqqldqgtwsqouOKFMEkxWtWYBq1ugPea3C2ZqOCwUJfYjbxP/i
/6pqKC0Y6wdOiu4G3DPdx8ZAct8pEisNwyOz0vKP9HbwSIGpvW+EIgCwLdkHke4X
DVcL2l5UHfG/W7PqXevh524VhXHACYCJYLmMhXHNC/saiFkX62FFb9GE+BOvnlFY
m13tWeGk9UU5ogcroVWY31saFZ0peDs3E3mzeubZmd5qwxz+nsn6RZ2Xf9D8sGDt
h2fzUAkHUNZ/xHItIAkaWiPdBsHuoN1JhEZcSPRVSD3H040dWBmmTnPkpPA8BJYx
ycHccLgWMuu474Z9EAFJ0RziTwNKBnp/7RW30tFUdjsxxUD0f9/oZjZb0EUGl03r
IyHExtuU/J2flKpHWIVDqN2Bp0Ml5cWeF2unHu1/eHefPtXDRlAKnyOp2jQ03crf
g8NyrMrn2BhufjpXqn/h65BJeSvK/wsFJI5gahOU8C3daTHIZrCTtXMiW55xFXHK
q3gQKOmq7W+yWg8LE49Rq+nPXmDm3XkULPKs36AK9UyL0BLVRj/wtgWVZ6Z/gbPi
CF4RYk8pADSMtMjioaOh2OemE7C4yVPUaRte0C7tTCek8X7NbGrUoJkL9N/9Y9qE
dL7Slf6p+Q/pRuJPGh9OjNUXhQkwhJJRyh3Ruvv0uO0ba8/SQ3rJ67L5t7TX0qZw
ZXFWwrxWNNBjrdCe7165eG94lNjjv9Ec8Qr2SMFojiUm13hqJQgijRUul/8QiElb
BPsoqZPLcRiEdVIRnECnohdk7dAbm9dg2LWdIhCwXjHqEqzbJ14/7dr/EPELkkAh
wDn70DFgTNT2RbmlWgYesmgQ5KfK4URuNyw7oJ2bxR6Sajh1UsaRwnjsgGJdOyc1
iFPQmheLXQ64WZmFSt6txqZ7q7UKbRxntOpD2pjjDETTvexsLlH4PnBMmu2rSFeS
vPV7YFggCaGRwIPn4fqjYYFVit/t7iMkSo0K32TEX16N0xhu5HYpNB9g5NUZxwvO
Z2m1Kpd5g3/P8lZ7rsTS9ys2ePZuDwQhvpUEZdGe/5R2asEARNkNqB6Eov189gDH
Xw/TMHsDIODWJU0ZMME5lqkUcM9eeQKV5MLckrpWYpTJGtF3WDRZZRz2pNhFY2o1
CmCOOpKRvdqTHA9JPLDQdL/zBei4WeCS8xWQSxR2LdTZ5PBqD2yeAVkxidRmUIpV
+jFKRg0+F7MnQJj+G8xjsFHZ2WU9hYip+M0YWh78JF6d/dllwXF4eRQ7yHGj8Ob0
WLKPArAiallus7QkBtL75prUMqkbJ/qxMpzlNtPLcKNjepfBOm//IoG6r4uuDfsK
ymuvcNpu15wQYGVIdcdOHOqtwDvH0/Le90ZHWx68Mook36n0+WKS2VBFexDBfDeJ
ftib9b2ccdzbl9LdtOiTktiYrzAtc0kwD+UXi4D+Sab3WMFaqEjfgkHM6UQ8tJS6
4MlQYZeYGNbVga74Q9bj0R86iZLNtj2EXqW8fnU0vThRouf+hlsGLLxBS6RhIo4P
Cxx8xF0P+kMIosECno97GL74nJCAFCQSEFbV3AdJ6E8WiOB5B4a6d/+YHmUMeovP
677q7TuqYZisj3Hhg4ev9Pz3McsPnGfj0iVCv5+b5OC0SkaVFedVlF0Ijfz/ISHt
smouVlSahFxp36NHunJNi+CmfpiJ5DTQ3xut9Gj49toqWgIira7VDo8iDDSkJVae
HbEhdTldGSAluQYB+OAeNkr738DLrNHnHq0YHK7/9/dZyP050G1qGqGnqxkTcGBu
5ESK8WrVWUAxhMrKqDc6BwOvzDLKfszeo7YgOLmMTR18+5pP35EwdCvG+wa6Ic60
37VUsc9pAP2L4TKrWKffKBOHPQwcXxYgivDzJC095o8YhdJh2Tly6vSgKSItlJM0
ljP43piyDJCKuec3RehpiwgUNncSDHRLoyyn0VN9LYzw8fIoJBuKC/MU4SoSrd1t
SRX1iBJoqE/3f8RON2gSYGm0XdP4Oz4rgl4tHYzT3Z0ckJDApD3/6j86VbOUrQdn
cZtqMRlUtdgdwye1Oq6xWluyMhsGIw4/2XNJRaNtpG80+ySP1brh4IVQW705YqjS
WMuzXZYh0tD11Dw470Hbac+cUI7dohbMIdq6lC1dSQEA9W4IJgSft49L2G3bXJkf
0W+DOwgTZI3AlMZvZESynh5W9Enw+TsXVQLSwsxYxqVnth00LSs4k69i2YOwTyof
FF69REOmDSkIPPjtEIptNy3WB0T+oUmczlEFxH1YIZUrdut1+ALSKpWzpyE8QF40
2wW568XufSkWCW1y679IG+lgVhrKtEH6+O9thAK67oBRQxr8hCk6anrEfCPff8Sm
6sTjJjqBMme9zajiXRTmo3iXWebf21nVJKPS3pmn27YvntW7n8nqL56o0VY3Yhyp
sYiLr0lW3G/feJwzIebrkS6AjS1nUgPy6gK1OACPDbCibDozBOw0KilOy/dqTji1
7895d038lRzTTSNo5Wt3V66ONA/HGBI9kI+AANV7dXKMstcsXBeFKUYUiEDIb31X
KVzVcVrr58Sa7lDX1ACu+4o2nJ/KU3AYT/8HJxteXUvo9sNDupD+7Kvtg/zkyNmu
mK1NgEZ/AKV+df1MHUEbReKIccxOzEmC9Th8oY8IwWMyqTXB3binhJD8C0HhnhXY
r6zc9j1zad6Mll6HI6x/dLXXnD1nlWKe4QuxBnBtJn51SeGimhhUSO72+9vSb0ZC
uj73lW/LjoSbeWpLnXRL48NkgcvOrH5ksJRavOP6nLbuOlqlkeQj666s3nCWyH47
hGssAQNIoGWthtm0uN1orM8SQo4G8sFd2t8VLmctL+oym0JwU4TkfAS1bX9gWmmZ
TqFSlY1mkfSbPwLLv75wDEoXi5Ch4nMb81CmLZFdyPxvsE1pXZiu/cgPRj4UenHt
5iBJ0vQN0DMAjOSs5ejoN73UZfokxvqw5M9fS7sEaDnv34CwPaZlF2dmJp2xmG81
jwHOaF+2W4zAsr1plFMsqLL080soYimVowKbSzHtSzY68clKcsSot7uGJRHxUCF9
Rarb++iAJBg7X207Fzr0zp75v+Xxb03EnXOybH1N+sdfhHNgaN5aWuWTlJJ9E4Iu
fgpSOwNEFQeNeG4JLQbI3qt+0y61K5tNr3UEcwbAeV6FTbW6c1zk0EVV3ud/zfBZ
gjAVdIsynusVDA7hfmazstry5eNpEKFYMkknsfCX0asB8FjWNRlELstlaMKwo4Qr
ZoIgY4ypL+bqLjaPgFl5MGzkQNDF6zPXdH1Y5+Nf4gaEoBRIJTENOgMQsVdrK6n2
pSvpJD6Jcms2OIPIR04kWSvD3i+S6QckxhuCxrctn9bO0kN0pq4CY2s8VAysinFj
0AmGbc/D/3i+IoQDQgwc5sim10vnB03G8HaJLDFlM6e4bhRrc72xjYaUMey1S3w0
LBS8Ck3dKrnRtkN23svyHb8MwmBM1KrGlJPrnFXgqVZX2hC1fi7lc1OnZCH+9LMt
K3fnMxdXC6ssnd8KvR5q8VI4JFmDSURp0g13vy8+LbeDZrZu7DvuR+8WL2UsAkKL
87HX+JSFfu5Tix5qKWa7PfCHb+mSO9lnIYzuDIEHM5EFJhEImMQIWv8rFirGQTEC
5BzVpL+YlkbCUUOrsjdjVl3D2bdubEN0N7qjpWAbDYF1DTh0j5EqEwsm6n0LA/p+
ZuvHhrd0znOt9XQxBBhDfbX0c7irTFE4JBZEyYtyKHt9+dUIawYURrW9NRQjFNVO
umP/sKvKTZ2s5XV0BWfY+Bl7pFuJ4B4ngJxHN00rtF++wEw1UPzHUjAVynsOHHGd
664pg/TLKpTBE4Q95iid5oKeR+Nr8to4VW2i+7DP1XWU17lrcp8WMLHms9JuG04U
NxIP6AjbIoW0aa5jU9Ed0NKqheKwMg8utsIj+NKTg5+WQHcbCMD/sOsCqNpDv025
9mtlJWTouHBe2Le54EWpNqWQ7OCtpj6zPua5a+KGgB1N48zN3h+Pe6GnqtJYZmpk
FJT1Z0WHmqc/zvpB/EJOKOf4kXhr15QECdITnHdxj24kUH/Ba+PafUdKdNX4hGw6
8zpsdC3O+gDh5fYjs5pFz44C/MlDKKbtVKmb7VT04u0fXCd99bzBihhue9P13R9h
bgNrVypv1uNLPbe5sfRT/7RwcF6YBH/9tL63MG9/MLFXk2/my94+MRuvk1VgZ7vN
5NIQg/GoshFcwo7PyGOYTpmLj2DcOSu5smf7R74f47W1ekMrYLwdhd3Sv4d6ftce
YcGqRh6QuhIIvAM9jOy48FQR1pKr9/sqS2Cw1Mt3W4RD+lqLqFCUi8e6ZnxLSUKS
PNvODoeW3iHVik9xJcm/hGO/83v/wqqUahaqaCZh98OSApMeHvLH5euh4wq3uy40
UX8CtoBedNH8SuK1i8xoezxAuL+uXDG3zzaHhvI5Vj70G3MSS8wwwE8xQ4Wp6iMY
jaSkC5Lh+5yUP3Sr3VXe6RQQPRgAK2P1eeHRO+lV1miu55u0u5Vlt3ioUQyU3WNE
iUuPPZ6lmk1QTpamjmUL1tqJ61JtTgxCRzNd/lHHi1sRveyoC21VonvS6+m+XU5R
y8q31JQqQYtidqPw4qbZs0OqkJmp/241A3wHnC/WuluxZwD0CUX9AJODa6TVdHaR
uugxiNLbHneqjf0TykN8qLc5fGDFvCYRPkpbuOFXllNgGwmbgWEVFwdEvnMBLq7m
y1pU2YDvSyBCz5Fg7u66+Roe5p8IRgEVQFjjIWNfsCqgesi1rSOgV4f+OBuJaLs7
WROb2C6Sc6itSm1LYzZerC7LoE9llWZZEO30IQyA/Hr+Xx4As0V2EDFAFgdN0nif
ell9j62m9eX83fkLHd1UTzd+xFMJCrY2ouNkAxjUG9rGMxYmpedTJOggOxDjYgyj
sCOrASx90h5MOI3Sm5S550qdarJZMlvDZOmGSJdHldWYh6/DyP5eQXxMTkuqY/9y
H4xw+e5hnudfZqWxC7uD+AlaYB3P+eAt4OcYG+mPNNwqecvG8/8I+tvTFxAf2gTE
zz3EdfWohYQSl6ub5OKr3+SFjnUffJLa0lqFmmAgQNnO+04pkSyYakJWVE3uBT0M
G9J3xilqUKDmyh6J4JFGnIGmUzGBGwXoU90KMvooHK0AcL2V0YGJC/Gje8vtkeNf
bitU4JazFIwgSDd+It3o09o4v61GiFdd0Lv4Zf6xPkeURmAP7yiobZLyrEA4l22Z
f7DkqLTQoItQCruSyp0Bwt/2JAgwI53o7ts+4rLS3g577+SwQn6IDEEcLV69sG9f
lwYt1VfAzybUJ78EjrnomDHOwrvKiDG/dcWpesQVI765qiySBhemCUAorEcascjs
M8jFAdPILImQeMULBgNCgXmpai+V4aOQI4HEuyCdzwpjYt8XJpGe7Pl9Ytaj0R40
cE4Wz5F+41WlKsIGCC8l+PpOScWRu67F2TMj54IUd7KUf9DQWTYiGZkpyOCO4ZF/
On4clLBZOeGHatraH7MN0qTNiaRRCQN4rTJt/Ec1nEQ45kdY1NgyKpjuIi72+LeE
PyL2OyQCkhr9+/UBDNRqiic8j8c+wmbUIU3QX5Tn1IauxQGgYR8FW1eDF/bbKGdL
JrO7XjDq+nkhCuPvK+hKv9+Cb+A/u2wJTiA5AnXNXes3p13hJFrOVk/Ut102vBva
o+WHmm6N6GG3DbHjL5kmLJrlfmHGVe4h6sX2e3jyFd7ibUZVwp/sU1MJVuCVDj/8
pUihZ87mh7qrl1XnLDsGeW+dJv2/tyMdR4peyT4POwg0BInzJ+bJEd1YWGvrEA2j
xUs7W91B8+AyFAT7rVbDkY145rNIbFcJ1ZgPA+Y5XyjpZv0j8voZMRIvSrtVPXWH
00xVKEwCEGWotIraAiJMgfGAqZkbRZtHcAebpOwtBlTqpjJELkpPgtBHyo4QL3Fe
/wx0oFGag8e83N2V1+ZprJb+x57eMk6cb8vyOT/3IjKN4N1Z3dclzwMw3+nzMOdN
+Tk8qtnrLPh90XzwCABhlENYi3XjA2zRC8tmA+BhB2kdcHLsr+gJXRSrNnpP0116
HYXALgoKDWqhkvEkwx0T2oj73ETUN/dlfe4PL/ErTB7X+SIGNYapuy/jZItvx7Q3
oXMPc/830zdcqYxXkBKCq2Gkn6VFa+q46azNtEKyO6dp12hR1zwsujud6YSotl8x
qt3loa112X0jkSR0SMHO35Aj14y+DPP0ymUiOkCb48ln+Am0Sa7KunOy13s6r6UV
op/ItBKKa2R6XnuH2VjU7At6Zu2qjuRNxcgJbA5ZArVbcKyUCSyBR2G+HIE5HTSj
ip2N/XKy32NBCPQT9Ol2EakoGfcAO+EGY/a5hPWp4Muhm10pG9ezkPRk2FwBe0Fm
kRZfVdWjDro34CcxtmchJVRkassjwRdXZ6mDvkPY/9dyxBOA87ij2rFZKVix44dw
AM8GE6UtMNW1ln7dapj+xrKSQzsd+u8m8IBa08zc2YhfTjrRP1Ui19VKbHL7U5Vh
ZRnl2KroROl/8zIVH63sEfU0ia3b/JADilyd8zNScuGi7Jw0TVKVEk6x6QdpI7Y5
yHUqVKeTyUUGsGk+9HYA147E6pPtNGO6aca1p7J4BlTGZKvWpaFKxeCqBUiJjQAL
2ti45q08Aog9qRpaVAeeuEmhCDlZrqABSUeZ6d37FKxsPp2fK+davq81t9qSmvs4
FLQFUzqVvjIyAD3G3TEKjw2YNTmSSU9yXBQkvcLDhznFwcLpmUe4mfLIiww432Ja
ya1ty+yD77H1KuQogPprnwZnVZRH9OHBdPwHNn9RME9WiJj/NQndfy+kGAo7nZ7C
W4Ru5FMlbK6tQS5mdmYXAHC9TdCdkZgacnEXUdtjaG0SVv14RDHumJE8v6VNUuwM
3WNtSsWJ8PSh3DV0zRuMkq79V+lchGKIo2RfpEcFuRmgPjrc79UoCPXNrLn9ou5M
WLtC4FWnZc0rj6hlHbngeRPdxUgS2SGfU5Rx8sW7kDHDFyvQ2S02deCZc5YeytyP
M54Lq9MrYoibvU6G2qzc+oUA5P5Oy2reT36gGeFpLm8nE6GxqNtMTTeCty/CiU+l
A8BgQR1s4WFR4huWPBQFRdgsycbstGpYDeQ/cbyjuEyjk7d5V7sG5yErIJaI8BJq
3odIfQIBikhisjE+OKo1/DQhGskSDHAUI+C46zhxRoCSX2lqlq+nGLWmCJQeHRG4
Ic7Uh2J4jhqUzEP8VL4LpBWh82kcopBpE1OsxRdiejys/HfVWI263jnvvpnR8WVr
AGjLCZwNuT/YCy03eHkXra5TyQAzD9kijni5d5Igu2BiNwCgP+Wbsw/XAYY/2hVB
2UJrn8YAuErDnQKcQJ+3HXsRI2na9+GDL9tcwXQzRdypdMoURNBPBXoMGcEw40nl
Zcp+Toy4XXjJuQSrCBD6yZS+YscEvZjCOEFH4Cl4uCTf9E6TMlcgSzQIRmfSUATS
SKt5fox08dcHyF1dNRvzYgxzwbBLXAMCjmW2Bgrh8pFv7WFQ/6x3/XbnoYfaZ5gu
nRX5oP/h2m65gN11Di5aJW7A7giRrl/x3lmClmccV5vL6EwDvl/vZXZtakakfw1H
mVxJ0fNrw44iQBSQr/LTvQUJFQr3JlLLeF3O+s24L3+O5BsQNv7Q/jd6chFbumMC
pr5DMEGcyOY3DsITCMJEJq1WkRKa2a2uSCxD9ZP5YXnwEAJFeRSJgv72DdYpHPrt
0qFd8+aP7Gwvx59V3QD6k6UT81JDfEAzxrY5adu3jqSNUtwTsL25mzRIVhWMxSuW
NxLXxtoJWIU16am54xPizIgzYlP2EePqNR9nMnNfLGVmJGorLWhYl63Plj4NGBxK
lya+JLG663acN+EFbUru5q1f+/8yHt2cdIdhvYLlMPT7e/iMMVtqumefmZHAnC2g
1PdBgdtz3CnNcL53WPYPPIsbUeh3795hZRbOym3RiNxm5vwVCOxsD8lpkKg3ApfW
1fMMuK5azxEjruM2Q0uNd+Ub3IF9m7KHbzzpENVi6tq4W8qRZwXZSyinQGxkVWSZ
M7+M8tmz91JvpDo6VuNDydgPAkwN/z2AZEw3le7eWzhiw+tCny29zSDC8w0LJwEZ
brSjfJcuM8Dpkl2CjNEAevswA87/nJIDW61CcYJ/Hue8rY1dKAWDg2/imfFmCXSc
7zu0HNpXzBRoAWWy4nCQqoG/j0GPVp8LeGXjbMzAb8NpwN0lNaJQyquV15Uv7MOk
uYttI8OGhvp5A4IrIU8/0E3Rj3af7b4/MVFUM22D5Nz0E4f6X4ZMV9mVubExKCz7
0CBwnJRszpgHSfu9QRYMQk8w1/bi5fctiL6qpsmJuGZKUtFNpVJ5hnb8w4hmajsC
WmP8ZOf8FZeESXWp5MPe9nQjuq+mI0YWl7a+xZq8BqzbYw5U1Ir5NVrpoTz+UEar
FdU44bq9sd8mA0u89XFT8pJwemmiv0AgTLDQ946HZoR4zVIJE1P5R81ixkhsyTRJ
MNXNMU3vX2uNnuQexGSIWEh8SMTQqYm0uUdWY/pr/tSltCH9FgatDKmEF9pIGEOE
xsm7L+YcsRMNl+wCCvV9vWTetV/uVFYxQcA+YoXFKW8F0GDhbNHQC4NKG14k/tLX
Vic9GTZ2bGzqbfXZX/XPmOd8unK5YyBvxx7Aha47Hng4ksOEZeulUcGl90H1kksr
N3RkheyFEDrZ2s1H2GQV6fR7jCaUr8iyxfPfT47cCM+JN/Q2aUSEELAWGcckpct2
2PQG3i8OpN8GaJTuUUFbq3J3u2LsFuM6onh7YkIHXCj/T9PrDp6tUPCvE4S9biSz
xs3qbgUVp41YxlSAMhBHx7sFp2fcok3fqYz69W+RYouGq6tcD7rPW4NDcyJFPcpJ
bT7RFuENR2nWxcibBjbeEdhzZzD6eiLoHm5XGCRyk2WTwEa6p8z7GU9EZjafXHdk
sVGp3dlPscKlrmi9s78CzvZH76p2KWEPFlkRitd6S/TS8aY+T/qAeCc8hZXs502W
Hem/GHU7FZRtOlAJdjGCAEcuxuI4dLinLPzq6uk68jNWVvxpUFdhfCfVwkttjXCt
BjYbMEwsGvfTVrTyGwH7sGdONZW+79OAT3VBnCzuXJjquRZRL+/zw4+jeyYKecaX
Z58anr96t+lz0pCva45jVV3bIImQW59jqhooFblrFlEsjxPYbMgOesL7WSzVetat
Y3EXPvLgy4fooU2L3C29APQrv9y892CTISnVPM8UdBNcvnxZiQRnm1K1tvDCoxbR
07dXRqNGUESPi+20D4HfRkhB74IUpQ9yRrJe5Kak6jUEF3Ic6LFS6AeE7r/qso1V
dL15u1k0N7V6CpYj+tuvuXJFyYB3aEUHgBxC6Xdyc8gubbQVzQMx1EjeaKQMAuAP
RyoCvDujAx1GpP5xj3CwO4qtOIj1lvDXD39JGXxZGURFMTbgtRyjbCipJevu55B4
jl2BWVdLZLTyxObr2XFMdpdpF+uOgg85xM24w13yUF/9n64MReg8rtXdtEsav1/F
ToTYt4weX+jl4R318qeQiXhFOFlRaXGiDuW3GhoXi57yu/A7Z/6utbA7ztx3n15R
M9KQIYmigT4/tsoKUHezD5QKUhKEeKO4l1r+Z6kXWf3ltAhh+BVd0HLVfPmdRAS7
yiZ18Yl6i2kg0CoXqJJiEy3dh2sFEku3IPH9eS6KvKRp7dUg4aVp+sEaKAZeesGU
FWOn0hHIAFx5+LkhPBjyLUGO7xBSm2B/Gs6/LdQJpriXsw+bOx9xjbQv7kHp2fr6
XV6ocBLIisI5XlrXKNr2F/+7n3PaHYM2zYlPxIMIDjfsj/S4Y9KrC+vMRNwuKdTF
vdIoGOmNOW8IZGVXHHR0JOkZUGPXfY5sTiDj0MEanwQPsJ5i1/yXtevQQAOttS9B
W1LcR4A6CszSveskALIgOraCYkmzQ926PmRnvt20WH6SzAW4tOCkM9UgsoWDcK+2
HcUB23b4d5pyE3o4v0jg7+k4NJGtmVbUN5Hkm7DqJM5QHBzkhUyWIycdw7jmxfV/
ZdsRRfjeiMXc7cHCU2HGzDChY7yzYx4BQaO86Q0ALcjMJJSNFaO2AMb0BpJD0bTX
1hifucm6lxBSEQfhLvwoS3wbWoMgoC+meKAdURhXUwTaThxIaGxe9Ee58T5TOb2g
L49AzRhTk8JCorKIuz0Xpg5G/iNDeprVl8UM8Z4WTvj/ZCSbEJawfVTgBIl+lih+
99EVe2hHFIP8SirITMFGDwrzdLiG3BGaBMxZOWk2BbCSuFZt1DoHz0zJqUqYaYod
1THOHdaxqpaig0JTLN9pjGzNA5tMdz9mev3FX/rSyRRgS351T9LrMm/P115Lpw2F
/VEE747CSv/YD+E22dA4oOjqkoT3s9Rn3RLuxjMOedbiVE08ajbtKVkiLJlMe/UF
DrSkkk/pZDWVkwGC5Xi9g+VGUrXVCeekvDSiaQHQ8mjSaNAxCHhQM4FelDb9aFnx
OILyTy+HO0V0txlpF09+Db3v2RNLger891m5GNd63Ai4T/QzRprcvtczW/YzyI/B
66wkrOIDDEEOq860EHIXC/6Kn2DyvPCIagHTfCctAUTPNZog8X3mj17fmqeaoY5c
kfAUCSo8MNc7npPak6n02t/Ak0GSqbq0bFVBekFFiCIvfVZqqXIav56qaUQDq9n7
GVCGNP9B+d0nay9dkUCE6zz5wuwfpqiUwxOvE5AwwHhiaKKk4svEQzXFa2UFTe8c
JrSiVInaLiZhhdRc2pE3WpiaNqaVEOEYwublA5Q06A3T9J/bpWQHRdFi3+bc20BO
LBiprdVQ0B7St9MuisZm9M6EmcdQRst/dDT2fGybCEtHJsZ9Qip4nDZh0RbK8ftf
LkhwLf9Eac2Dfva37Qh7RC8f5lcIFa2nvvq+kp4dH7gtcL93ZRZZWUG6e4ePFvkN
R9OY5ozCxfsz9D5ugkXufwkq3vEoDbD0g9eoCZ576BRN4X4x4bwyFsAxgu1QSPgr
/9vOR/o3a1E0jkUjZc4c03SrrLIJzy9wR5RIoFmRjN8yOc8BXrW896s7TF1eTiln
wu4V20dnnhiyWYVXmfFy45WPAc9r4KcX3MlYyZKlifPTSUMbnAs4SA4VsGCfGggz
I3JBcqZPATQt3zwg9V5+ahdCm+0+w/JsHIiH/mNcO+Jbn8VnbjsQwhIoCqnp+Etp
ZLjxmGQSV5LTZdp3j9Hix8BfTNF1/q55i5EGx6LgI3yJs3fhuvvAmQRlRrWGVxZG
vFIrxPV9brnSYHaGQ8Qddu3F+yf0S05Elj9Z8oCNP/3L5AYE2PNcsHxr37JggjZg
iCGfaCrjUyuGiazYOV6BE8QUq9GUSqGm8g8ESFIreW2Hij4FrusrXWnw304s8Quz
shMVr+bik2z0aFH7VCqBt0+rGcizFiKFn2hqCEdtcWcRhNP89ILAQdJY6Tk0hIyb
jprEFVMgyhhBxgFX7+DTTt7CeUTJC+7ZYB945Zpcp5VJmhKC1xlljBb3WCObpNBx
xdv2G3swum9oHC8xh2RVpkdUhDkfHrqPYIUI66o+hfi9bwghfERaS0VMYJAns6KF
1kPMWTUvvmrlSK8B9uE9URpBbGJkeLwgC/iRoQlJYzTDb772NB/DlO+Fad8x2waY
tAKkc4x9rURhlGIG4g/k0RfFuuuiI2S8wg5PUjbLbaqs5wBGLvmkf87qLUhZ+Uj3
wKDYEqulE9xLKVIa29scNcNNhdiNsijiT5fqdVQ9aVTfvM8ApX+jx8FA/q3NEYpb
+sPjpGpxR2+CqybZU3jcb4RHMRUrYl5LUWdwtHh4tUI7QFdwUwLN1MzRgrRS1tj5
0U+1S0cXqfMIBg3VoDJP3obl/BJI7ceZBHtwoL2XahUrWgHsm/iO9DHBbub3UCoX
PUH5IDu1qYcDM8nkMxzqbh9fZ+PrhscDeNV+nLCloTGJBNB3w0lVaJy9qer8C2K3
6VjqvR9t7yh8CTqF4S/C8w90/1sTT1afbyZkBXUEsEnOixbTUqbZEaFw9cdEbbC4
/btbFoPHLuKDSFEJCocmXYneCyEt9p5llylKzRBz5xhrAot7vGX1mcJ7dXNrjRaA
BcbjSoNu/DZ1WoTU7Mt9iScIX7VpteVrJLomNoDMBM4YxnjSNFumCpHQsxveKzdr
yNV3ieSs3GtBdXtZ9w8TfMoVtdsf6xxN4Lx5DmFPA2wNN9OmrS6EaWoZ/Nw5nh4b
JCS0LZSMgdFDHe7rbC4BvGu6kQfo5APxU9TjTDdHBpWEXCzdYnK6SPLBR9eLxiXa
TkUyIidNobARYosCdNzPP+iLITL2gCX5KRazlkG1xfNgJ/vgzC5Xk6AqyUtETcK3
lTUwH72ArP4yOou31hx9P5fgZ/xETEU3fRRdiQrYLUvwkhPxjakwsDhTIg9Gim25
4GTp7KTxnMhpg5BtrEyF4VjiCEi/czMI12WwJyX7sKLybOhbftaqu3vlQEnvMHR+
KE4Bkm7QcWAk08JMfEtEnsDybc6OChXq4syP1mBD8C2yOVOZp/ENLbNhAlCIz/hB
++wmQlonSfAgvwcy3XMj6xKBQOa6g3Fb9Lw4Y5W0CPvRntD98Ja5xnfDto1QjRST
TY1RuShz/yKN/OSGdjb723NLoXWCt93iqib1alF6HeIJXYAI/1FGplghsw+8/Erv
lwzSu7nyxiy0/+RGeUxZ9+RaGI0iSI6DBMIc5ytNBIxYwayjngzUOk2a74A6J0cl
QG830C5D32aRlJNONjKwTaaMuFpYwGx692tXZCjIQsVhapnkJF14eoBFb+SNezac
tKOqJ+RBaz2ZnvfrwlDz/J2h1vNIDj/qX5nDoN6IXe8ixiGnrBvtUToSST1FrofL
cpTORCnSuDfKw7ir6I9VZON09BTyHOMW9hB8VsasBRcINTL0mOjIMeSj50T76ZA6
DLStS1VJWDlLuk5wK/xNfHjw74Ec/CpXwdrUtEJ7mlJNBM0wmqskuuxd0OasVxnI
odQqJNEFN8we++I6+X9TTX683fWNwn8X67r9dVCvJzkOAg+NG8XXUtAXPighmWTK
nKe6mNIl/Y0HZKe0U7q3X7GJ0CDpTY+isDlbeDVxG3t/w8uf5fjLbXvVmhJ3M6Vk
CvF97iwkZ5RryfTwI4Fheql/W72Ml9TlxybiLbIKQkZ2vp2kh6owzSzjo0hliiQJ
fAGzsaDJeUdvzJDqHNiizMo9qCas6XLGcoC32BW+wioXxn+csq/V7XlPCq5Ia/b3
7rN76mtNNrLAEENFIWnF1S92vMPzk4kiPjQcFVn6x/WjS49ZmxaApTtD0rXNd0y4
LciXvKl3Ge82rmq/rT3VlXzP9R9xWII39XN36amaNfWS2bLM4j2FATjygUaZ6ogV
VDpihqKkc76cxDbEulJ+F9BdUOUoXYIsJZpgUcprowH3A0W0V01khNDHMp42ja/M
oSWH4+fVkmlxL4gup3s5IshFFmKRv96nxHM0KT89ryGo6Dd07ur37wNtUMQLCM3K
NsdHD27omgfll4F/FSgzsH+8N2JfzHNt33IxLt0FqPFf259nP9MFBguMMiaCKKJk
am3dX7c81BQfj0Q5iqfJXs5kOHwsdIry7dBWJSCHdrO+MeLKE755SeGYLiuqtzu3
yH8MqtvpzTxBlWWWFemB9Icxcj028mc576jtilX0CaKuXrxIQ9zl/0vNXYm59FtW
wyvLh/XqrvoOSxmIicDlwpksagxqxlikc+2kLsn6vjkvnKWQkEs7CU11/ON+fvyQ
sqz9acfkou1Rjbuy62g/UGBtmdW8aXOJaaBqg4ovgM4fbtsycViIPFgsKUoLkyhD
0Y+SeM3t0bvmOu10aVxqr0WJfPyH5qz7fwD2EIcFtw2ROBmRUhgTzbgY+IUOWVbN
SYFmnuTGorDmSxA5ohQYZFaNDvDbAnwiGG0uzE1saoV7y61Y3O5ZEqFqRwrR0DAs
Cj6H7Pb7G+gZzktYoRviFycu9K+gaHnVBJGw39c7gXpuBWwBAUqqHykZHXOjT6Xp
sTOuw8U5paN2NXV8L/r6wKczsxrPmKI9DGst1vfMsAUyc/V923nWZuL5W35BQp1z
f6YSgN3kieIACfOMvryZL7NguhQ+HJU8NLNUsV5Si/tINRCiDRsiyYor53AP9IDJ
78Usy6BTMb91U/S/nBbyLaEKmmg52lnEbT8Fuvh15+k4+Pq1yizWi3dQNEP0GmpR
iODY2mdEQ/ZTX+5vuO83UrmT5xsQOuoNjsq9Zn2qZTf27v027vHIvHkV6gDQCsMc
iA6Mjf5SIZGlRIH2sLx4onfMsgoZ5rbaunYlr9ddgbJI9/Lj0jLsKs3mtsAG083Y
O9+cWPM+Qh1xbqC1WRCpqECzD0+oRQ3RRArlVCBEwJ/wNyUsJOgJjB0VzwLkmgPE
4KvP68Ga1daj6+hHPczBnDOq1URcqz31NygZMoYe39ua5g3hVbzgqWPlfkprg+I2
LQfmgrHPZZgDbTfx+ZMLPCFnpYOFTFgPJH/5PjcRR1GQQU+Qpka4LxWu/EYYTZga
YVlLQn2v8I9Z7UGd0EKUouDmLoEuC9CMxY7dFokYvSpHzReRMYnv0iMI9xnOoUrn
IYJUoqbNje579iYPYHRtpdZJds35GAolUpaOSiYNYvYGINfs7RK6J+ayxQWAvK4K
5F6SaUNdaMV1Lt44ikTsek+z8dP/Npy4XZ/0RcUOYriVe0Taejegxbc5IE5gGy0p
jEwclkThqrqQLCjVpsDZrNw6vZmL47SMwaJmAPvlhRdCkNplkZ1j1m9IPanW4BwG
w2zG6qvQFY4fbmTdx7JgBs/tQXPKAVt9aLVFGOQsW+v6jtrhMVy7rNZskIglbZqp
cArxhvpoBhBUpK31G9t9aJSOog/b4Eo4c6D+Bri3QhtVrfC89Gsovmzgq6yNAMAg
gS19um2gXw08oXu22nT5HWISpf/ibEbBrc0hmxpB1CW+G5UW4UDZWm8puYFof8Tg
onXyS3/aC0Zjnb8mF3qvxVXF/BPbnvnI7sIdporV+A9q7Cc5mwyA+NoYOki1J+Dv
EQ/YWK1syd5JktGF+CKEz5erohKTGzBkeG9k+EJ25a/xko9hKtFFpC6Q5KkDpgIU
uJcwYKi6x41xuCKQhRK//Rai+GHCM8BbFByw4t/+uCDT361AXTFZSjNugIZ4oBVD
I3xNREfcjxENay/kJxngoYJoaqpMZhN0xUovP4eZmHHTSWIAGCZZwxQuRnxBDvnW
ZbbcrodynecnQRDMLUD7SBDqPMc9X2NbHQSc8Fo+Co3UVav1KcsoZxvYlMWKYNxW
ObSiapHwB5ABSj4dwtgjhlKtiHefn/JhWABIpFSRjeeK4pKC9xV7oqG24lXt+ffJ
DShLdDD9iw92QayQ5u9TgELJrbYk69RJvTLw+M4/NNv0PmZExam3oG/03zyQKfC/
V2HRRE+lDdtjKl8e/R2v/FiP65fZoiiu2PEO9cuKXuuUuelIV0rJ0kJlK78ALUJ5
9vtmM4vLAt1l/iM7/qCxYkYfOkxmcMy6ALseUOm0xx/97+i76zl/Zwt54R2CJiip
XjFaLDy++OxNpGaACxhZwqGyRQ0BE6VeOlVpGlzFUIv5rRVw7TmreEhr2/moKIXb
WRNDktaBhz2AfWS8rT47sDrLN2vb7gZYJw7OElSTQMHNFRLXS4AVCkaliM+oEDN3
SbFvcDxFWnY5ur7n4sn1c+DMxhUJC9y6IGjbmwP3eAPBIEfyQK0sbytQq9lVd3GG
PUedOUTOlL6yoEtvJtsDu4i3VFq8c4PjpHkWLMN2DFjRnIKpbku108faJioMQfKl
QyiJ6aWn0Pao/7mvEvBkM3OnGc9QEthgNClBnfpDVrbrohUjR0uVfmPHiPM1L/cT
bu7ApgyAeXGTdXXLyQclVC7UWkLPzTjAj+QS9uA3jM45HtTDXcpRTYxHz5sXbnix
UgFdV6OE6hlIieMAkSpiBJ6aaVxIkxms+hfm2P8ioyq1PDVGJLDanrPhrQ46ew3d
PNkjaeW+g+scu17xS0ZyoI+FeoaIwa5iMIHNCpirXtRgx6epjIKPFMDXOWt/OqT9
2menQpw1JgI3xEHcslW+vAlXOP2yWOylmduO7mIu1qS9cy32gkqpxFfCNd96sWEL
mNL9yLNsApGTqTdvfi3M4TA1z8Bn+Q4JSJiKXpWiWYrfIsT92yjfqWIl8Sx5iB0X
9Hm/ekZJauX2Y1B06/XLXyTEv3DPTEArCJrp6jp3o9Bkf1wj+nF6ELhaHu7ACk31
0MaoP/QbujL5BzzuO2VUjGUFK+EyD9vCzTWpdUJAiZHLCvCGCtlOPcRZBUQZ23Ny
5BoTTKKBlEdwpgdvu+Q7E8QmnO4kyT8Esai4A3mm9K0lyfAvlwg91UTnDhhvjR3j
42nTwRDceqLKgiw5S7hogpYkNjQRdx9goSoKTEQPAOE6bOoPngIImeGbLlM9GW9o
T8Ce3L7lKm90E+5SB2sGXsySG4ypUFd3KTtv8bVFK9QepwmgVA6upzqVKTI0U+zo
fVNAL9sG/FVr5RxRuTaE5TMtFyNaNSY9JOPel21/sdK0xOvwQb5sU3O48Tn7/oy7
uova2aOxbNbNcjAGuyTSTCbQjRSLHqxgYQQ6EwX6CTp8ISxGa1qd1LIgNpNzPQry
5rxHAXFwyITvt1sSOR62yir9q6hKFrinvvcZ0ml69k9Af0s0p50ejAzJD1+bAasU
YSGdHnCtbqCn7N1LjCuwrFlJPpfez/jvUBkLKtBwZjVcWec5pjqk5NDEQAN9uw4F
dEQHLr8rViGYrjSLXixNBGMTyRgXMZ3yNH0ISZrfOhfg/akiE4IvDw+8o56JIQHw
AylCrEmtmzPs9987jnPAF//M1WxhPHtMn87/MR6ibIf6hdLbIGtj+/fJn+3NZTJ3
T6QIyJgx+8FEEsLD33s13ZpIaiNGm55gp2zUgey3TK7yB4B8BXLfEOEPdmvCImnh
L6Nbwyeg2uwWZLXTJo+bkXtVY08q9gb8KSE6fQpMtMjp7O1DSOk6p+YXImehMeuL
sIRRMCJi4IvvULwQ3TzuFU5+LK3SO26AfVO5NPNc99BkvPnYjCSRbtgkYG7SfMFI
WZH2MiB3bCVtQnsoO8CaKfLypIcvlXPNKGSBwKP6Ys4pit9WIJusZsUVJQCnAJwI
C42/BViuI/lCQwbwMdukR1nnsL6HyAvGbm8B3kYTeIprzVsy8Fij/DtRpxL1jpCZ
hiPutHgGscmN7ZNabABL7P5WpQ3/UR18G2CUAUBmUsaSu1jGmHu8dYZSeRqhibcb
16Vu8oWEEVNh4UknX7A/pydTpDNFK+94RymKprEdj0IbgeYYiBIM8mQbyOjUCfHz
QtuhLBY3kwWoH9pGN8oBarI2m+8zlSqhl84io1RtG/KJAmhrVfc3RS6HAT1jPTyy
H26pFQBh3DEZcNNGMIGPA8O9VK4yyJnKRDSK9eC+IkXhCB7sRgosKr192jfg5gG1
L9V/EP2e7TTAlCfTUzFcMfEAcu49Gc/29lq5tFs2lNp9XxOPzWZP6r9Cwmk5Rftl
0L4NO6gRot8st0ikOTFDpb7fCU12tS+CiRnPlIXqs2IDM9tWT2BwrAvDK0MFzddv
T1clI7YZWzb75hP4dP608uWR0TIwl81ygYvxAEysoK38M1/74n4NPbuLpMXj6Z3M
7AjlMOJKL1YcpNkgMhnWjM/kJeDarbQNRcSFvDCrRwfCtSYFGxiJ9BNtJlZqgVL+
dMX/UBrZZK2EB14YFxFOauzqwqYwrBGJrcn6DvMnF1n+SxjGPS6zNRs2Ti9YwOlJ
RWR5hGjmYLxsbrJzWOmaDVhkcPXthWEckMcmhj3Ck0sylpKgk+yOfcEFpqh9NC3F
sI9plaFn300iyjpmoNf87qidTqijEnn0Z+1XjCEcmO1JiBiyxncuITvqZ/fOXm2u
hx4NXLJ+gKTlN+nR4YFeGxUMa/nKpXPVfwMUorG7fovlnCm+SX2JDQq610Nvwoy7
+adYvFIxeWfNlPJOE2cfl6ODyKP2KKhNCwZzC9N6FiRHYd6OMmSWxmT2Nq2Il1jN
EVBH3WQWOIM74mrghkL9B5suWCCCxH8kDUDZ6yk+9Gdbyb5wTUnHrDN5JwgGuFL+
/A4jaqffzv2zV86nNw9Dnk39ax5YeDJaqBtzo7ti60eU0AtWXYe2aIye3FlIcrjZ
JAQSbQnbm9MzuT01Ew5NRqgVlye0M1iAksriWaKQTSF834PIc8Z3DwJTfWHOfSLB
PKl/Js99A5wkJ2dSDPkGKo4EIZ2kRhCcG6HsrT3j0ocW2fnRsiVscq/g7gizwlwY
eUVrx1PZw7t/WvKPqg0f8AtaCGoe0U22FbRtl7Tzz56q13BgR+foj7WWG+eJGIRN
mLGZ9e6zVxqPi3S7JQmZ4SYxYwCpAvImJyEE5r66CaGVLheAaiTvBl7FicMNBlhr
Rg2D3F0vL40gyl2FBQaf5IaG0ag6W5jJ74daMuQyRlJbndQrPyC4sianm10ya/G0
13JZwLtZoaSn6BL12tHCc5U/lottnMuO8kdmn9K0blEbB+yYGT9g3cBYJ5LKrsfE
kmKN+Y1GwYU+JY1ULkL4POdXMn/CRdVvxmKxW+ybfB7C0Z55nByOQdBc6DJJoLA0
StPVWjKC/bRp8NkW0IQLZJokE0kcMuljG9a/Ut2dF6rg1Ej9M0M8IeOsLM3khXk7
nAMKeeuLpldaRDT2pI9MhsC7JWjXV+veJTQF2+hqsrkZwQfbrWJC7cZqtRSmXXBJ
9j5oiah3dYuFqFGeib9FKAJr0ajW1iwsXa5Djty3OqBgxfnsGb0WXciyHZ73bGJe
dlNmW1vuBSWogafrlv4113c1iq6FBxVd8JDHUWGvqhmr1BmIxgDS1lhrapBjcPDJ
r1bEJPGbrmVUgMDjBq7hsM6oo8fWhvoqZau9xAFFTH7X3Vtb0dK+IOKK5JYOxGba
RGwfQwk9smZ1sCXKo+LaSJNfhQMtBT9uCASua6+dnc/dl8PSyLzml8yGeKTqNQaH
646syJTQ+YK0kgMIKRXZoXzAjyPHUbcJiJQe8a2f7zAjpZD/TvGPJJ1jaf0OpObi
zXkeRQgw00+r2N6mvVvejuheT+b6JHmtzD1HDK1dmyQABGNdZeyQURuTAnR9CNTR
h24wI/+mMzOyYce+xFwKbq9FYu7QCC7xwftDXv87xMZLoJ9wpQiwgZdgWTOy1Ekl
w/L/R9Y2+zBM44mAAz/7eIr6Mrs1wX2MAjzrM8QUQn3Fkzgsy44NdfjDx78mEYRF
qNwHsbi7tIxxdu7Q8xtYi0aLQcfw12PVdp7fWOAIkNXdcieIN7oNCjMCNL8ozkGG
z7nu+cPOZ4mfq55/N4mkISlhJN9pNBr5MouLkU59KTF/woeRpPct3akl4y8Ejjke
raLcIzvYeTbjmSjJ61A42NHzrf67MOD2JG34TQyTtnKuiIvSZ0OiSRk0q5fyF3vP
qUVBeBIKoIhzgWirOfzVyqWBViekDuuBPG+9ZP+5pOxFwiD8GPZIosSJD2Td1g7r
Dmwm6bXk7RzZz5sWiUIJudArnkLDhglp7HpBhbCoiZbDGqX30RC/iW2mfI3CkBYw
Q/91skBacz3ptNdotepZlRlGbpp87SOHg3Y32R1bDPXlt1CgaiPk6pKEEWN7WdzD
jCvaEV659LXY/wW1AgpZ+k0aTLQo9epMFmtd1AIeBJc4VRDn7hn8xeuEnjNvkh4o
ly4CbTGIHJ4IBmXhOmOy5cDmar53O+sC2pUeDCfzJMmaejNGEYc33Iu+43y83iLC
fGJ44vNkdDxnEv/2Psy0b7v1YlmiN6A6mSQqr002kYAHlRbPonq37VPBAdTTaj1H
ShJ5vKOgwvxGmLAjzQLGZumLzI8SpmoHg9L6jKgpWIyX9evTngsobHQiT6GQie4H
ZRJJ2pGXYDvBdT508QRkFxdg5hJGgU3IUqzV86ijo3+1VQL2BW3h4tJHGOq/5gwt
YLx5IIYIPAYRUt5s6yKXtw4nNovY/5e/a/y1AN6hKScuLaq4GU2O2QTjr5i7Dlhp
vTU6/xTfAqKmJROCYJso5JYoC+Ohu3fSXDYO9ybFCPUglU4oXwcBxPz9rf2IXyrC
XsJDVZOWlhPYu6hBTcuBwUqKBoIOKuAYnpqokMGJiQRe3i1BswkTLMCVf0eepz7f
GjjDh7A3KSaiKe6tVI3lAFrgTEo518WbgHRjNaX3T4Y/hIsRXkLWsOVwqCS8yQQQ
JPf954TDWWwT9qwwlhh54GcBdhxY/5OaycCHf762cBiBCusnlO7BG4VR0iFWFusn
pyD8vJ305upWAR8ILGoFboNRksFv5d8gpNtpvCGN0RmWdAeVDzL0rbtyVIuW1lBc
xZkvZx2RtCMDssNNKMzm13ypxSltWxUj5tz4SfJdVk7TPn3JEV/9zakL1nyGM0Re
4Y6Rnc5lQXdFG/zyqLstQRkAd7bmBoHi5ORQTagoc7GzD1C5l2wLzhzQLok4WIQs
HtYzvT+E3LYn5+LPPZc2/i0N7kcTfBNEal2qOX6DP254PoSDppzZtKcXp5uXIoRJ
rsvMvt1OUuLZbaM1I/v1fChmjwGD7yZ4moWhzRDR7RUbKHC1J1Ws6UmYw0dPcEMR
bLLgAHCtPTfVKYe8lEQ9nKUDEw3u8Z9hNgqO7lfaKun8yxxa908jk0Qw63uVIVo6
tyczpHKMmxl4vY81eIFx7hKvFzEzarRzkkxbxsbIvIAeVkrEOFKeca50zwlUIwQN
ClpPwJxg8AO8244otax2chvb6lcvsIBt/7Ooq9ewce6ptasc0/MWwhhsafY4QPFB
Os0x1HwIluRpEzww9JE96Hue0/fv0H6GmxW91eC/akR9oc4PtP5TblrtN0E0CfHx
DskAw1OYcuTTsMp/Yoq8kQ6J/eNmCbcuohSYs3mq5UKOhxxfkV6f14sav5JUyMOF
BYmatTn2AiBhVFGl7jmr01z3oa6YpNnk5IZWS8UkOVhEq2cdJeTCH7OspHHarcXC
W4j7haiwx2xIJiG7aHMf/gvN0I1iLGquUo736b144uHzfvGPc5GTNcJjZhEsthFH
Wn/D431nPsCh4F19uI4NWdE8rkZXeHjSt80t4n0kJ1CysmZ2vEddWhceCKlry7Rq
5ZMZfrzKTZs4tgPhLALwptkKLCAegFPzI4KXUaK5JuSX1kAGD+uEBL55aGjGOTFa
m3hHbzIGqEefdRnH1tlrjTDwn68Jv44z98h/6bfsnnZujMRM1TcvRv/YJFhU2cv9
V3djpp4P/7op0wEXuMIJAQgSmNPPjnksJcigWRi4QvNk6ZlQEC70BrDVSo3NPeT0
sQNvHhL3CYofwS/Ojn3T5TDgJiZHOpMHTi0FtUKKk9ViSSNU7Pc6/ZEIoSb749YM
Un3Q9qNUvpInAYcrtg6/Nor4ZzaoysTfRWDyXLZhOdfMAVbyFLbidbGl2YAW/W4f
fKYm/K5BiZ+YIKG8dH7ITo/9JPEjbuc8SBXCmbDLZ1iZaCOo8EKHT3dN2L8M/iap
Q6eBSIsoJPKZ9vRs/zbR4uwbIfy528GdPRnVBkHOi3PG52sn1jswWi93nBeQJKz1
GJjZsd4RXs7NQQvlQ0Yu2ylhJxZSwn2NTSMoP7kV/CPF0+fBBAvB5p6tADQdewXR
h6wCBte4BS/xW6SjkY2Am9/Z/RxtLZTdbfARw3RgZrOD/WDhOTZfxDefl5MkW4YI
0WM7/E5D9r0lv6DA/G6f3fk47yzS4/8Js0fZY00GisvjUMt/aUDi84jI2CTl+sfa
IqO8+pP/zW68gBGt2+uEybW+QsIzdT+OdPvpdIZ+ZJsU3c+Ci0Krb8umgNXOxezz
Z8fzj8SNzlW653KjT0NrgWpiylAhvxGCjkBEoA61HrZlpbh6i4rsCNdJxRVJteu8
N1UhEmXfbo1GRFxz1x60Irlum6o9F9DDfuWdGoJT0Ii4sBiszwPBD6tCbqKFBfps
OxkV+rN0VHws6Ty0y8PrLvnsiwDL9XKEW0gdw3eMVdRscrUM0q+GeJoDPRgnH4mO
quLW84QrCjKRh8m6bVEWrQFcywrgh3vEt/e1DT7oR7Vde81ca4vVzu5+y9s43Yo3
7p7ibhXW8F0YSSwr0ijszbEEEDFKWf6ekbrC+EQCLihn9+YKFE9vqJXgzUrxvpIV
QXUesc31nMs7s8fU7tiVcN3Zbd78i6EDsxPMCYdGFKusN+g81FXf+pIhBpQOmsaX
4oapzCOcGIsKLEt0SLx/TUzyARXdArFCKPZ9osmWucPHDgLvaYfHJ0XRccE5ExKA
NEZ/WXeSEX/cqwQW9ch+QqQMbb3PRHGbgth6ti0n0ZIxwxdHIinzPY8d5priqZnh
y2Tr9u1dFfJ/9w9EIs11lyUgCI/98bOEVhdH2DmsiSP+LO3fhU0S1BY4j75UZTJY
Ecfu2MoTOa2rUL/EuDOY+2DfXOtUfVCJBCQsU5KWNoVCFR53GdS73Etu2rCP3MSa
N/ZFukffmg6sohaW3uHhgOoF0HwKe6f0tQV6gaES1hwb/DfXNdFGfNPkM9bjA5Xx
HSn0oVNsy0zgT8hLVEu0I/lNwNNmJJTZ6tnpF/Bvr+I4jzgNN0Bb81wLXeU4odhh
M0rI9U52q44ARkcGu4tj6dbQM/omXewZubHFLKA6hoGRMty0SvKjxPB0wMLKfFzX
1fNM6GFVzmmOPbzYpnjNXBr6JD7cQExmPOixY9yNCoFoxhgTxkjJX4V0ECWqqCwl
TfzaXbNXZqcJGF0edURjnp5qc8dmKSQMsmKnYq3PKjTNdwV17t+DrbrLOAWE+R6l
yXVN4x8xD0D4Mnio5W7aOkdCoW8fSEj5+I7ful0AzUZDUjVM+B2PuSvDJJpWEXD9
7TpH0sn9qqQ/fsXMdw07Zc64qXEUz6q53cNFBWanblX5aaSr5HudaMxUezxK8ONo
SOJtSnNLGvigefDhNlGLXbxXQHYnN20daISxUeZ2ov2U4JB0TJ24Ga3nenmvuvGz
VgHyXQmTwYc258NPk3YSpWUZ5IQEvgTrpYyflgn7TthpCDSArwVIqrGGAV2Os4MI
fb4nVdo7+J/0zJS+2hn/ZmuWz2CWZiYV86sK59C860J7Kryk3UWYAeDpshRR9G9o
BQkWTgxWF+MouQAT+8yOKjHxv7SIb+vtuDFfQYJ2MqWzUU4fAHsfdAR+EeqiIMj2
JM79AGA4bQLVx6wxKDWy3UAokewRnk5RIkhd1NdOz5Xfox0ziD6hV1Cxl9sa2feN
YovcrroL+ghPetQTud/FM3IrenL4yMioAQ7sGNORtbeV16SeEuKeWvpz9ummDVPT
3rPgbZbPVEwtFTENiA1iWKMJjrsGtfUZEiW2KgrBmVl+Sh2D0uklvvGK4uOKX3cz
VDOi4lEoubdMcnaggut1ekatA8AS2ynZilNxdHForUTM8518nqE3Tj1zOjamdrSm
mzbqYc31F1w2OnR7kMeuOIaczgN0dVm4D3ShGNTY47IHp3RQuDeSyH08LqKEL8BA
bn4i0u7MdTmVA6LQMiuLBeeDEgCfAw0vIDLCmgQuC14sLbHoMF1laNco1EMd5ukn
21uUNr3NeEHrlB08d8T1RokvjKQWa+h7IamBPJkj0wtv1xxPDwuIS7nr7XWSvYgv
yVs5UFppJXbVN3XOThshYwZ0657sjfaBIWOT2Mbs66oXLEPdRz+L6Ypl/X3RfSI4
cQCC8h7CrxcXkletSVq3cPxeXj1Uhyl6PmSBUW0iC1Qf9kUYuTkxpdeGsbsT0IPv
ypGKrrBSr2iMi7ymRP99EyVLC5hZI7H7tqqJPkcKnzlp/GgZyj7S5dO38xcK1NTB
C0wn4o/ieGqES/Xhw7iBkHJG8YFI0UH+TilmKwGwvNKyGJiIPqDE3YS4zYDB7Spv
OSg9rW6AHGV4IX0sftJU0EKcDTnIMBVxgtXuojeWNjDvdDDshbpODS3WrOrMURDz
G+G+1PCoE07mvd5yPfQMUpoL0kwyhZS6K6bmffO1IgY6gR0+/u4wAlPFjFUqqHkm
3l3c6avfMZ2vnOAD/+FY8UzGi1RDKr33hAS5YG4qB5z7QlXZDMmMouzdHa7qHe9/
Oiy8AV5Nv+Ow58nalcoYNuCbzVCy6/puVVo+He7LbdwVLdyDYR0X5dwCoIRAWLT4
3pefbwYstG4tQlz9pVAD6Tsx0egml50QD5EI3QGhEj4O394Aaeh1tsf3BxkDKYiI
tDhADTMC+4oCJkFNfm79lDULIACfTljoW8TZHXFFRtS1PxXmcBgWzsUnaH1BfSfe
wgn4kkMuz4qu34zkcCglhBdvc3Q3Bkrd5Lua1DzVM1zsp4rIdDeW4p5YCC4wwGVO
CfKfAbU2y55Oyuz0lZuq1pXK0egdxImmkOGxORubKz/VsrQqVPN5nqf7f9HqArfK
30TiNgjnmoExpgPwrIyG5uDEUbeSVaJ2RxdHHimxHYRv3d2ZgIs6yE9zYHjMhaot
qC1Tc3BLQ/S1Zzl4v8d4r0btH3xaNCab4M01i4ivYPK/mf4YAVyW4A70o2h7DDtT
LZNXtvVnIHPwvlsui/xUuSGCVoerf+jZ+Io1EosnlwX5WGQvZqxla3Zrpzf5WjNu
01UdUKzV46coRP6O3YPkbt6x2Z40q2OGvMosSCNA688ss4SoygqV9TsPU5xuLm/Q
9PM3ddZJ+iBHrZIXdo3gxs0sARgb4tsY5J9x1Di4owkxPeOo6/o93P4Hm4rITdDP
siLqfxKElKY9Ijpj2+MtjVZBGDe0I5mDi/xuZPfOQxgaBX262uDr0a2R0rfkn6Aw
InaRerUGYcL7bnKyY82cHHb6c+Ih+45w0kpnY1QI8sso/Qbk1IpollKEe3Sj0Bw0
OMKG+f2928hgHnvwNqJUYGW+dPfxp5KJ8x4NYU9RJ6hH9lKFVqdi6/S5PPbehAUs
UHyB2c7ub3BPito01UK31RqnBvdjgz5WkrJNV1brXVEof4QjLYahMZnlUgPshCcA
LWMwcXdmoxw+Eh8lBzy6BohjezQIzMI3wGoRp7LVTUP9pYwec9jolrfeuJwC7mvz
PI7pGZ+qatVkFy5BOIhHfzBbJJjqXuS+Q86QdPmwy6bFuAEQh/Awmh6hVNtKJgXG
xadLXmVdvFgX/TWSUkZmr3xMfHM6U5PF8Kj9zwZjFgag4ILRYRtRb6DdIhXfG3o6
BYmLN9H6b8WH7y/ulONcQZ66LNEfdi7RhFGwhzvNcwuhISkJzz2+BriDNBq1qXjS
YWCqCLY/hOWzAvNL/6FKdwZUETRSNtOvMk10OM3XmShzsWkoOIc6dJOguQjbVu2L
g8kQIPGHRb8tlW7jNe8JPLfzBV6LMFejLtbIbdHcQVpkw8+S4V74436wKUPk6jXZ
UFcV4h3cy499hVI5Mo2t9Yzok8Ef/sBx5NM4GOFDMmthbTJtXaegCo7isFsb23ij
CacgST0h1KiGlKrzJLNnl9uxuXPFYTWNeCQA4DYryt3UErcvHqbJG+xHnop9Exk9
GEtQN1Ugh52O6QTbDYm80k326ytN29WTl+tFBgmgc96sotaB8gnwYGN+GQ5h9Yju
if4RzEqsEIgKaG2WUfN1+uf8js6oWPvKoEtwbT0lSWHUJzErE62aFAA+Jc9v4qOW
MXSyRBBa8P67K2ffXFD97mS9orc0qMSrwXAP23ET4lt2y2yl8ITmGKVzHhWl6vg1
0fWF4KdQo8T889mVbsrsWd3Noa0wuYrL603dMSnXe3zV9idkM7mVZGJa9W06CVW/
nVldXVw78+YzLLl49jbua0vjh3NjFAVXQPOGc1oD3K32ikBAM/SVibyqtUqkbu6w
3JPY0pc9eSmzriO4z6yOESGPmyCbwcqwbUUtZlZDXcfP7bbsP9ww9T1y48SXgPQW
GMqoCHbth3d3XWNxBbdcsbawWzsEMG+S5tE3VwyZfmdu1m3h5t0gsNOr2W/eZ0ZP
4isVm7FgUTZrYsRO9ea6U4W0Gf66j8ry28LbTfD5Der1w2MGVFIrWDnJMW29kd2o
ZBLJZVPyvU0Z2S4AWiXaHTYlX+HJp1YOnPhYVsI5AD50AHfAPO+s+mLhdVL3dMpp
Y4Ojd8JIzvTlDvfqxeUuAqqDKibVEligYV7iZakTPZv0g4vVGgD4cbX4sZ/wL+23
d3bP7vFDlVVqbyLmVM/WUBP/hj81w7CPlrWhjGebiv/Sw2Lfu994jg2ng5vKMw3Q
yfVxHHzzRNt+wTGLmDGRpmZVoJyIK/41k0jQe/M9XaGPuynYS9/xljZLWKmMXYV0
pPCwEh6R5IilIjFDGCPbMpRt2OkhBWdrD2v2QhfUKlDsqDt5jNGaUBOFOcUJpu+a
cXQWgMDJO1BWLNCOfIQmZoa6xGcp43dgxxiwdqTRd7EPYB+KUWqe96x+aybKanOr
4Tm6RHvxA64DV6VwUb2QZrr5+wWnYFWZXlJUMtHNOvFRV7gNzgYDDu4DIGglnwue
zvBo5pt6ohdLOpcb9y11r7Por3/6EXInZ7xDepqUPNXq6V5+J7PZl4vZDlzOYGYu
v7wD2VKgb7ZHbZmmwvu96X3jX976tNKwIcUVloq0WRCNSvkWMwybziHPQErtiAm8
EaqekDC57wyezL7NMrwtaEnagVoEzncFojFMBwT5JI2ZLJVB8Iz5cYY384dvpbjd
4fPJ+ut5o3TLGKuq+ovW1ct1yY78kiA6Ti7k3wUGoxaocjDsQCM42K5dlyDiy2wY
befaAz+16uE+joUvbSrTBvyVZ/xtQo6MjwPpOlQpW0bd92rPtcgS9y0rtgWRPU4O
+nicPhw40/xRFtivcyDC+ageGLfQbmz+VOAK+m2p9Bmeh562bM56LFEIHduJF/bb
54is/YG/Zt5LnHifx+TIRCx+KDvsp7uwI481jQflPLk98QhNggQcp5YxooPmvORN
zgqlaeHa/e1gO0Ti5cquAanlrfI8R1y3BSM60MLnHh9BErSORX5TqCVf7jJOIsBm
7yda9Mm2+fcGh9wXO402prQmMFleb6v8pfm72BxNzReWPgkMihRBcfDREH6bAFZE
PslVftHHCLAXhpyGyx9GpyJxITQrRhbtAbLurixorxEb+wgVYsWt3bLusj8SAjbF
q7NguAzNmbn7h/KWI9ZZClfd/WVwl3U3kTJ4HXzYT3vwERCsD38JXaaVHM1jwZ/k
AManotBbF5Ku2gB8TlUMniK55rxkGZLxki0qcyaCChsWOek9HHAgDcE0VW7lVR3k
+SdayEgVP2iR8IlW86SVVT6yHOjbWwnazoxztnPx4cYVImtM3sPrGNh/W9nmO8Hi
bEMTVO0tlDn/yYcqL1ACC0294MRRa4uUImsV9C76Rja1k438L95nuhe0bLW4uqyv
7ornAJR9J9XZ/8B1P/x0NNHwWWPSbtv0Oe9hIDK48XniWR41sRux6LTbD2VI5LnS
7SjqYLLOuvBDDbzI2UzeL9ArE33VuqDWwF1JUpOUX4QDc4sFoYkBuDiL/NvxAeNO
NwnjLypsGJa54fp5iXnHoIQTNQUyoDi4ahTxn/GAIrAGrf0ZVjBvZLa4mt8o4a5m
qZAuz96PrZQ1SwulE2FZH28uH3i0KrwLf0Dce5QwgN7vOhMDXJw7CjjgrO4wVOwU
1J4hbTOILn8oOOfRi+so8VjKD1WDArRYxow62PEqCYP9uZ6IFkUBlTkWzSAsg3xU
yo+tUKE9tlXeL9ztsXKabF6MwiHk9tTMszQUi8iNt1vyV3v6FQ7EB8UA91+FupKa
pZmdoQGJmdT4r7OiTqdUJTzTb06B+DomAY96ZX7rkpW8oS+6dkx9ko/xhxfCITue
Jybeo9XXRmTg8R6iOUp/3wjGSmz6shgp8hVbyQAAr3tO33pSxRdZJG2Seo10ENgS
OAAW4FC0X63L29ki+rD8GdddbMCbJ+aFIim0HoFM03gW6JVCeR001cLd7ZkOuwz6
bSJ68Yi2XwpJ2KtSns5etvZCpFhQ9ytoCEO+F0lERN6bvihykLNSDP73+t5br+rt
4CtPDkOvjur3Htv0mxL2yb/Fg0vAYcZsj/C5pUa4aX3SoMgqtq/FkV9BCz2fVeZp
cLl/CAi7GjrQ6u8QqGMGPTDcC29pW9pk15qs43Ud9BpnEXFiKUcNYVDKhPv5dfGp
XbKdscArvaTM0JcBIKF5EOcR6Z18oAwjhzM1nybeHtQrOXTPXEq6zTgHyDZIHEI1
lQUaOQ+E2qvcdHX7JvKgnGMh/blBxvOyxEmEAz4hTlX7Lndhbp8comYGLsWtrC+s
JjCjhUbAluWTEJ5Q5RfqNRQAWSQUMxqeSJ5qZisvWuvquYSnQrjLYFgGRiVL0RHA
s4f5kyKgvWhAYJAySjXcLNqx+MmqnGsRdywdY2FBgOhR0yIqP42eO15nz6OLpmB0
qIf7MHGPOWl2+vAF9IvR4uq5+F+bL0BBcrfcutayFQ7ZlBpS2hr5lTDm+CpLh8R3
82yS1zz8+wzcEuyoDexoJpg6u4BQTidYS3+jOTbvulNptE+ehRUPesRgN2qclEpH
Y/fwna8af60wEo1GEkqgyOROU2ruuqVRlYCfdS84spvA2PSJAAiYfXUySRbwNExT
LQg63Kp31x8b+6tYqa5UksJ7Diuw3yUpPnoWsmgtDmGb7MgfnELtTcA/kivHGCnr
dWb6mw5ALa8a0FzyJdYA9b8/Z7Z1t4H2GB233Hhkhgs5RPzpQLZ3Kw7Ydnx01iv0
zYkkaJSUN7s4ncjq215Cy3d12ml8HkLI98DluT1url+SbOLmmOh5BLvbx6JdGNpc
bWfxLJ2HFGag/tefySDJ45q692N7MOtEfkhGcbDTFmVnaPUkEy9Fdw5egxqpaUyX
mJRqk7ZsCmuDZ60uPFsQ8x6Pl+QyyZbCeEh86kPhT5eVCYl0P9csdUnzSZ9Ou8gQ
GHk4WKu5ud0kz42Ptta9Gz917N20l6stY1Jg9hg7wOWhuzRkJSnYUdvVhyUcUJ0v
5GNL8BEajD1//oYmB/sgC8NW9BTA4pUf7H/Xs4oF4KOiww6WqXwE2hT+wCPf00CC
+AGIlPPm2CDit2G8TW/Cqvb0ha4TO4xolqttBl9cRF7wi3oE5BRKq1wiWw2dforD
I3VE79II8X+m+olhxwZCFNWuCuMacnAoL2PDoD4KSf54JGZpmzSI176nKL3mKpSa
55hGgxwSetx6dgnUeE7XGnmOSSPu2j69igox49oceG1k8qJ7xXjC0lNfHoDlp/ka
QR3jmhoIgV9OmxqNiZDcQOfkt68XApfnPeluZHaSnl90fb/GlCUIa1uwDq0z/eYk
fu+pVC1UIuOFIdXG1fnnLf3gT7XIg3x/s6Hu7/I30wcN3V90b9GonAzY5g0TxvCR
uVYyXitR5jP7XYRIJQpsXUYJTtbHOD3jkIaWheeLk9oPEylgk80Ny5d23siNicVd
uErm+NJj0KF5pZ+RANc5daA3iPO6aQ8rtVe6AwgE4EoLRolv8uo0SXVuUwAoz0sN
gh/sVSqJlJ5F9YsQYpeZn1fhqBnYVo/BAT0/xm1xU1CVOHR3qw+Uq4wLGoXUNVVj
+YwVSeh0NBiX0wozAXJk2yCtug+DUi3cFqHa1VqwceWWrVKUoC8+h48AXcBZ89EC
V0AaFHDTcviCPL52Hcd+ZzlaI8Hf/kcmiqO31miwPqeMVrs+QdnilZPCkZh4O9oh
luowtM1Es+YQJ4ZhYxlEw0pvgIKOOM7u6YaLPbIJerYkXg3gV6SOn2lOAUjTSdid
zgxGBz+6Vn2ScgeLqUtTVU8awC2WUNfVUXIYp9FtWHUBvSq3j64NJdEiIKKwx2FY
ODSst1kheQMvTw5Eq4vk/DtHVa4DVwcyBey9oZUVAK7ajtIUVQ5VdLaCsoIGpoux
QGJcU1/WKPv8tvRoSDd+ycS/Lx0LfX3wBcC4RANOovpD6e3oDCPhWMph0Myt/oCz
zmTO8LPLzldZD7eyfsPytCKt0Kn2A6dyQkyNEJAKJYdapjN0WdXC2C/3MnSsgiHU
varQ+fKSisHRFSuLoJletfqJh6J33uRw0I4BEqiauOBlVa8p/KIYfAs4ndC0vHMm
YjBd5F6UtsOc6K0PqFgz4mfIT8k66UDsUxgjTpN7E5K0Wgrrv0gVP81xPNec0RLh
V+PAY1ZWejnLwPTzwS0ChnOcRig+FvIXoUW/hUw80dgcmNnOHigFxFHoXGy+SH8/
exymG8QvMs0v9mCG1TLRJsR3u5WrH939Q9FtFsulnCLsXpHcZiMrA+2T3VtS4cyi
9qCNHHLf2exyNSJnbUIQaFV/KrOSupxgJPrA5yXB9P5kANeQZ/+cyGZgz9MUbD6A
tHZ2v5ryYO7k0QZYvynhiXH8TZVvdMLg17VMCnUlHMZOnC8+RwnmcjT6j0lcbwqk
2ghzxuJUFgR8UqI76EbeZG1nIwfVDn3C/tnkKaZmkJeBONc9DSQCtzeGdP8Ivkuw
iDA4lM12+XxJPfOJeU/BKSGOLjET3XiGBV+nP0CEAppHBr0cCHwiWmY8jKT4hpjR
H8NLMBdAwUgzDh0T5lOGr94ZZai3y5I6MqzkFaqJx0w6qGQEA2fiXjpaVylZcPAv
rL3h9JjHchiSNwqeWndN6YoeYxn5QajQvPdyE+5pfFdjQ3BkhUemtAVfLcYhNsMs
oeqr74JzuCZP7/zWvWFxIPrrhUgiRnvHCe2XSKDQ+SbIEown5oPyr4AAEmQ/F976
+tmcgL5r+trVXB+JKyZkSGQKa2rAWhHMKWTkCRRKWUJ0yhi8aY3Znh2XTPggMQjN
9i38x5np1b8IyHiidlHTCCpd9sM0qz9I9vhtpHtbR50lMB687EPo0+luuM48lr8Z
xRYXpnw5bYfkGGG7xDeyD48n3/UQ+AF9py4LGK2w/Zwon/OztwJ02k+Ww72B4BHr
LFaJ9LHrp/AZ3f2uExSlOAWIU4/Qvw3aIwvQf66aRY3qARiUESJR18PUhBr7reRx
0EpmNZjoeLpqGyr8FLm1KjQaZnywBU01wrBoIxdEgo9K2JsdVM2TAEoCH3n9bCxH
l+Cs2zziwPUF8+T+KJzzTgxY+lr8kAISs+x3EKpFR8TXFpbsKZ9QXTV6EOSrNnNP
g6tuFplSxMqut2UV1/rUAg/Tj6M3RH4upRxPoRse6IIa08sp/r6iJwNJVs0QOtBT
Wn+IgNOpOYhidOdjSx1bK1ZE3JNcyqzw4Dvc/4qEAaGzstbH9E/TN8Mntsxh13RI
IC2CwuPeT0m83OGJfzjFvYWuSDZ3IXCSfaZB23LqyrL6PaR4G2Ke5enKP7flBvK7
xdIx0JhDmN6p5QbhaoLHIoYFDIKF41W4si+2/3Gm0S8yn72NTS4nqUHXEWBPc8Bk
dpUsNATv9RnKFFCyJYAJYGmCc3eibo4/h48JDnMnuXUAVOsymj5W8zdXrM/4+n3F
3yY6qcl2JNGv/S5Du/2tItUmP1t7eRspcE2+4Nm1uFLZ4Yp15MSFm9jo29inZF0s
6+u9Iv1t1zwj8vdKwd+FpZv6v/l7LMZFoueJ14aVRzlidiVjn5z7KoGBu6KQdQmB
hsBydKioy3h2EsDKYqghlZu2TPlGUM9qx7OdLxt/HoAf4QL9J/fTAX0PL/DEUNEn
ze4Hpv+u6IpSfbDqCZ/cdETsYgNzcc3sbNjPuXR/IXCTNDHlOLLNMcR5xW+XdYwO
umkAGdyIToTKCi/fXm5UVGbHePFOiCvwm20Wl7RDCv8gujgFL5gfboPSiIZ9p884
UcHz3A1Aj+aB5Fzs8lO7j93i+arn4nUnFQeIouTiFXs5Zv2cdZ0xWt/pKOrEA1O8
7D3MWJphsNN30uLk3d0p4jebfFSK9q8ajacYzGWqRRY6hkIXmbcmYrR93Me/7+cG
5WIhKzfcWciDEL0GuOiQw/PFGRIA2EkgZK0v56NVo1k+81DVEgACysDpqUdk1DJ5
BbkHCJMx2Zfd/yXwmL+FWCVtJRyTZVnBa9p6i60+jHdL365ow7zXJrwOFD8SRGry
2XxuKIsGb0fZFoirNjRlL4acV9T9+aEEnz9ZVqaadzftxEgS8IZ66EegO/X7K4C+
KSUnkb8Qu/rLVy0Izk6vN3BRink880IJZHxAtFvG4C2sNrpA6WjBRp8cFv4oPXIj
0AD2RPOx2rAdJeOvk4TYnFCV5Usj0wUcT43z9Iiu2N/VkY4aN8on4jkOlO4zkfiz
l3oxSj/DAQuHkI6zgM6594/s/pCkjQ5qwmAAwyJ8//1D9OhoCzMFdub1jCb6zNAw
nkEJgKVKyCi1kbVKlytN3wen6+v6dUhD0b3E5MvMIcuUzuPr48jDgy7Z43Dgypro
f1BEunQghTApKOSROnGYnI7yB9eY6fR09Aiy/kqmwI0UJbN89Y4uRojoxS710GkY
rKsCw2CvlDEIZJoBiB6rd996bN0/oivA7mQLALACRJw/36PJtICkycIoUtjiBul9
DSHWNMjoL1Z+8DchLTtaU1x8shY1n3+YxPLxSBJMW19k76/EvZ90k7PmFxxn1RdP
d5prRdFw4NlZfUsvA0sJhxwin2qovjvSRSwm8Gc0y8/jqhBWH/8dEha6LQ4rT6MQ
IpTtiF4KJY0l7Ly831kGh9z5yEIF0H2SS3Cn7Pqte0ajk/1oDdmJQRbS7Lk6/HiV
nEcM8E7fciLaH48D9i0BsETD2Vbg5z1k2ewI1dcL0urOhJt7r/eLchAOcaZ6nKhf
RQWaKfEBuxAyNBe/rdz6E3w+/tdMhqjfQLRVRwPrM3FqQmSf6kEE3NgsZN1y8Lh9
VmJOBHLyh7SNXFmM+XbT+jJkiNuyQ9t/qVhnSskO13l0uBHiVxR/wzRn2aVThXYT
kNpO+9otKK0qlaLzIWEm6z1/w90oITpaJqf9EpiRaH8v5eBavpxrHK67aOkvKNiQ
tmi3s4+few7MlASM5ukms8uCUPfxE/TE6KZfvKryNcpBaUEUFakEBJhGiZDrlnOs
oyI2WWOtFn2bg/KKbMq/ndMB1W9DYnWjyIFEtQgEr781XQzy5j/MSADQKv3uKYiO
NCOnEvf2ctRFH2w7n4wwFdXHRgMsisC7r6nHRZ8Jp+j9Iv3Rjhx5G0iU68i++lm1
Z1kAER1AlfKxm3xNbBWPjVbrrZGXHwtsPrcklKXQDuLY1l4SEhp4ytnPI6thUIeo
2kTiTF92byLxB4yUh5tOxr6wvDyI5++xSEDTLNGOAVSMJgwTX+Imybq4yrA5b0B3
l5La3VdHhSk6qHf28W0hlCIZl+n3hGi2rq70uMzU3D2zvOdMfTgDMufxRjKffZdL
bLwfgs0pr2H7BtkykgDIPs87ccpdqhGD2mrDrYvjXzF4iCsXMjaUP5NSQ7LRpniQ
5Lgu7dmwSF/0V7AQ6pdb7aF79hZRBwtKfWwya3vK1duy/rfGgrblHoK8fwLD5H/Y
3eTgE3lzE/BZRTG7JQjrlsg2ayQfaVC9XD3vlh6qZeAjVouq2OmbTPu5p0EKCTeD
u6QcQWx+NkDtT/1QcO/dnPc8oDWz2w8wm0JxWh4JhR8Oyo2AmHM3nd0pSvfKbZxj
TSN2NAWwHSYa2pt/KISjNPd8S4yg2LiiwhTSC+5usrs2g+IU9upazbYPEKnrokkm
QpBQYjMK4phNWrGAWH+8JzdqrKePtVH9nLgAIYJ9eq2/qDYd8kGQmoLKieH/Naw6
rno0249lXP9k+xO7+wTnnB6gK8wFok6qpcISD/JHzvkpeA47TQN2g7mHn5cdRcIX
pMfh+t00PsIXGoZRB833AmTee8uJbILlt5EV4QbA0XALmi06oBj+i1qbt2YHwPyH
lcltAqyxGGWwcVC1O71rBfoCMmzlynMmCoRBuLvN4W2bMBl04RBEimNoAclj96TN
1Q71XPdC9DMRay1rQUzDSt2Pm/wuumQ7HE4RMOanolVMyrx/zuch8AmojLsJ4Edb
lCjKI0rQ2ESPzuaYD+7r+3PnrZygT1myvHhDinXy1B1przLjlIrcmq5A9CW2SMFH
RVqlXomqo4UqyyeEHwWfLXtbiZoTOOFTHZYBjRffh4eH2kCtKuZenz7ltC1ZwNmW
3OL8WPmO1dkxEFetZUSjUwFOmXtE6hMO165QJYHMhgPWSWybaa19DduEM5pflI2A
bEkuN2uuVCnUVZ/js63Fzc7sUUVGPFurBuFSdTHeD2wlbAOBkWhEuSc4sj7XijrA
Bi8aN2Zq4Ma19s1eCVcma8hxbrjzeXqwcIYK4iRdCmBaIri0luQzBaymwVar+gG9
n47gH4MzXlfk8JuTaDoG5E0+NYYKnaDGaB07p2o/Dg7Bw/Bu910C6mDy4zIKlXGp
IjSTPZYfD4K17gv5np5Vswk/x13y0IU9Qw7/E5saJFdQ9pngc4HQMUwXSe+B67fb
A6rWstmoOWU4h09DKpo98fGthaDF/GDC47etcCtvHwjTN7Ns2C1MjIq8XGzWllC8
d6RTk4E87h8WUAqYX8sTa7gFk6qzpubv1BoJdS3SNb1zujqBEFeJDA9BV0D0M+79
GYK26qqE9YutglVd3njW5T12Qv2m7y4RXobC4jpdeGIkt248U81uXrW65FjFrlsK
tBt5W8t4mSzORISlNqOLTeG0RPdw8Y2JxTHEZz2/69j3SsYHJiEy3CwkLDP0nVRv
wKyoRjABY9povMpSqdcPa+OSW9OD354Nw2u+koV8nH8ZqAwNN7xh2WYk1y3bdtOp
bUtE/JlX/14sgXHYEpUbk4FzNoD/0NTbFYMuS13nw7uf0eCro8GYfedTygrl5kfl
P3ieUumrbR/UHwk+GqhAkGRzlkXlfSSCaiU4bd/sM4sdb//CtBhspTD6NQ+gnYU+
m95UOjEGmcaIJUaf4024e9cNE0v8jkCelxPxC4JFs4M3QBN7xG0zyEAtIljL49xf
8Ke0ogUiwDll353QYkY7iYHYFbhjhrA7V8S6NMlQtcRNK8NRtrYDLibVFYtIDiVW
di/3j9whjy7ZQeSem5+0uHFohBS/UkTCPNlYqap6+4P1+IdouPOBtUGHbNw1JwpV
V4t9evGk6ulryZ5mG7vek1Lf3rePvy3WMf1tLxhzxl0bgkls8iiTz+3SEcLoOfeX
irwT7pPfHxXfR2jTpQf/zWkuXjvnJVmMIWutgXQD1eRT5jkf6PoNkW5N9c5PO31G
Pk5UaQR+LIJ4kWX06GCjx2+sASOPPPJODChrCp2MfVux4TBTweDyal1c0vb2CzpQ
3m4yqfXNuDc2y3+IK+nu6PUGQOgqNARx1lvryPUI0jwbIgN7xAKFu/bHR+AYr3Zq
4uBxh2QoRBhZd9oHPHPPLmY0iqQeNJ3nV+WZ23SkeIDUvYJwL6Y00OpFM87943U2
6iCBSpGtqUpxrHBK2/n1B57xLdWxHnXZ1G7Sv8efP8vLHB6zKqAHdX/9qJduKsCv
6+ViTaV4nx6fr9uK+HN0mKe4O6DDcPBUBMG2v/8QKn48Fo1lu8YhZrEky14LPUiD
YovB80A7Cnk2XMX8Gj/HgBVI+ZKZ7MrvBV4H7HKa0DIz7V0eAWjtM1VDAXSDtJ4Z
GqAIQcU5Ogp5m2MNfGyGiNuwBIk+VfuWFXkOENLGeQATkgtl2BDPVG+8ZAxK37Dg
4XuMJUQCZCMFjf92mC155bOtfelhBp6wdeB9mU8V3bpmP5ir8A0eRpImqzlzGLIN
smY16j2eHUZpf2qRWbFgpt9vPUMmfLYkH8aLve1jzIcsdKQk2LlAMWTYAvzPJnk+
1zIFJZZeISH1nLzb/1z8sF6f5zJljCFd060mrr01P6uMgxHQ1X0kj0fz3bEtG1HX
5A2jZ87tAxOQg9PhcwY+470yph5Af6l6m067V6qwNo5cuipLCdhs81y6D8hTJauU
P7iXVOh0LRlbheSgXyUXeuR/DKNAQ5LnVKzhgRh1pyTAo5Lr5P/6a81xKYidvxTU
uRIfHMmIo1aDuSacR39pbEnvrpTPWx3GmvATAlQAiNw8aCqecrWoZ3VL78Q+OSP+
VWy5yWAC0Umnsv+i7Mqx842/e1mz+ALkBl5hyQxHzjfyfUBh7vEYfCLJoL3l7hb1
viLoLSrwzW4E9eowmCE1PZFvEL9ThTbpJXQUUiHi70J8tQd1gjg1Gs4LZn5B2YWW
AjKAxeiafP+rglLRxlhb9mIcYaGOtCFSnzyrJYP9NmKnN49lQrEKYXLydW5Ix65r
3rww35IRzVUVCqmfEr1881yPtP9dK4nhUnnTyZCK+GXxn+NtT5Ajw0TNma1ZETWh
tg5+y7ch0JXFjdcl9lBtFA5gGbsrLfAaWe1oUdO5yVYTUxCyJ9nAW6S4KbOHkEdM
eBDdLcMmp3hv7IKjV152YqXwWavP/BYeRdUapAPVwrtcqEdYYm6J4Uk5xhVjYebV
mFfiP4D9nwsOxww8Eppk0toXZkiBhZ2WY84n0psgPNmAXPiFBdX8UDeEGnV6U6Yh
g5E0blfYoizCr5omJ6OYQAxzU6UeUkAHovKmOyWnuL/m3o6ofOb4+3V6zMr4XO8a
PvFgMorGifUDcId0jhJQ+5XS2klz5adkDiArx6ZoTDoPU0raouaIQMPLGcHIiIP9
sAYE3mbjFwEjs/pF8iinaKBD+jdWTdrZWNj96DSR/kEqphI8ipSXQEY70pEwnQ0Y
FB+d1DkB4RzOU3nh4PdejnFyExaKqIWwpRE07W4ZHXf7Xnz4vdF+yROi89qJRd2Q
uxmTZKKhcXk89wWA4+TlVM1k5Lw8hNJWCf33lourm1nztyCqgf5OpLKeuGWCykCF
IINGEWYlBNJQ1s8bMq5J5h40jNGjyF5qInOTmxbaL0fV2ohJ6fFbjdh6WtF5InoB
yQMH1sc3JzOTyHPtl+62wEphWBlFlSPNJu4ADvTAyjiCWUYAoDBaoUqLA/b7yHi+
36Ceh+3yTocwTAK9VIKU0AC1XPoekIRymcbiR2gdKGAxgF8i1Fu6cqC1UXL/+L4Z
+w5bdComPS4ge7YylStUZdoOCgDuC19iQtKMre9LmF4v8x6G3/M52NG3k0ZEZGE6
r0ETdolZSYF+QPRqe+6aocdRjXodxZlNNG+x8oOJSWbFtYqlGKI3Kr9/wgXOhg+U
dYQkHb8i8KQFLYAVvg5gA/EuW510RlOQdkOpjizGDsjz15JFyayZkbAVF7cBS2/c
ol/UNVhzoGpVVRh238Sswe3CIpvBUwzxQMDeiJAiSPUuFc3LEnVgdCqbyIzXXmxI
yS2ps81GzCxaSAHfIXBVdOqeK7DcSeKY+4hcMhT/IRIQRbI9AAz3SeMNwLjnV2I3
USvvQ6UEZcnl7f9b3V+nZTGWMK/SAFe478OQnuYdP7EEPaMHS3eATsofYNkJHVR/
7LzxDfxZ48CcT7YeklSxJ3vL4uhGIIBffkIFbnyLCvo30C4YfDdwAaD0txIkHh7w
ddbvfGumLDnzNXiWYfGBLyYsyVr/2zAC8PKSGjNBJQ92ugTVl3Q26zDZI8r7XOLx
PaQZSJdbxnjzEya9hm5EdHV37Af4UggasVw1JTpDA0385I5EmhHsSv8Pn2W7nOC0
nMwkFwasbnl14ZUjP/XgHRDhc9dCTiWi8+n1J7Xt45DzagSD0jw15xfd2U1Qj5mh
So116MKo23w4b6tEeITrft4w4rfcKmehpruKdSRJaz9CR8vl/I5GSMpI+n+MFUsg
zwWQicSFVsYymyxX4W+YDz2ax6ivpvjFQUyiPZ7AXcNlqxkx12onOXhx+MzEa/NG
dyO5x2tMH855JueHA9PTef01zx4H88K2jLQXjTuTFW5oL/ZVZBG8CK8e1X3ceu4a
jtvNS8+ximOS2f6IWzctUyFg/aggSs0GexL7K6KFeFtPo+GPT+DywbcWwjYIs10Z
+FqYxzAohx9ezJoqMR6l7HVg7Z9COgF5gCFg91cg0citgqil32/VMXVHQM6xu9XZ
0sJ7u303/lrZe2SWPjQqSMtCJvjlVPj684kgC+6mjgFCIoR7PR88AHEokUtNuNZH
5UgpmRJPn9GnlusEeNbXrKN9HDK+zVTnaMWkcUcKlsWyUMzj+q3Av6tZOmwz/Pyo
kr5IhIAxMUKsZX2pujF+GTGfYbATv+Gaaa+WklQKInoGtagKNU2X7wNqs1NqYxNI
Ht94JX7oXcbc3sAyz2cRLNgV+7XqSYKgGp9kvJHBa/8t4FIW54zYeIe2egADG1RP
c4pc6FYe4EAcf3aLrsr6fUFwpqZ82tItWp8epYEsmPed1Jme9CxRNE9zky3ZjrM+
2KQv+jCLaNrHoYPE6X8uw1Hlw/cd252inVAfgOj+ZywEUqozW2WWhJNXwAJXOV9S
1bI36YYRfiudrmXmt6k/8sFlCDNtH4VVwX+2kn2I2nj6yt9Omk1oD5JKIPZeKcPC
RiaeeBNHcmgfZ4BhVyPeiHsqAVHGJfrRqTM+2bUEBhiClsF40BLGbsSlwpqRtLeo
YICEBJ0g8hp2wkevJpXPmoEw6CPvQouTCTFPPjfsJhD0fuUnI1Nz4Ns+zVh4TpPo
sZAq4/5HDE/gZT9YpS6yN44zIgd3mxeEr3sRJ4FeaW4cYYs5JC8wY8WkTlM5Bo06
d4DlI2orrXwfTdv4uE4XeHfx/EcZAtdf9/fkLAQjme4VEmMXe/rPwoDwGVniYz5l
pcOdsBXvHuSHpNehpOGSTB1N57aFbiEZ1q41qV7tG7KBMRB8RVIlWv2Pox3ypaTa
nFaXG5NoGf2O2jtNdCzzw0j6T5wzeG2t1+Qz2AEjHlgqygBah8hokCxd2gA05pmD
oK+974xGG/mnAOCKGBMl3Wvsi417CxyN5Y7uxi6MBT7khMeSB8wR3RwXuU64NFK0
q0XOz8PdnLiZKWP+Z64uNCGWKKrgLLIV3UICQkeZ3znm/6dH8FVumo766pNOPcqe
AdYk94/JDJa4rBJT/K1XO4ZMp35Rv2Sk2gG8zZipNeSJz/8PTszRU9RGY/T4qRJZ
DGRtQ6BK18SMEDNgA3DzA9qyhCZIMGcFQZmzSvgFd2DRoZXjbTwd90MgG3H7Cbj8
HwWYe+5cr4m0ROvRv1OHfIrwyLE/i3gUU8gU+DrU/xRWro5MO0gvnxlm0+0hcdct
BCgqb4C2lkytCFI0ET3fwkAHMBQh4H12DYT6pw5IJ3PIPzGMmY+arYR7PKrHR2OC
nnLDbpcgXC2a7ssaBX2pgzYuZD1wsoCCj/tbxyRHh/Pj0uq9lIUe6232my0xepGp
QR75JQswTQfzvO6PdKboLC1CV39ZaXkvVS7CBtnNkXbwWqjDlAP9CzPkfl4tu3vi
Hgt8QJbJHwfr5dRDOyfT5QL15LtuBQRo34AKzhDTUgJ+H4WtE//NZhUqpJzYPXBA
+ZvcNNDPbLYuN8+PAVm9rSUdWz6M9Wfk9h3IwBCiMhLvS7q0vwSjPYevCTU/BuL0
l2c6jLVBdZShmmR1WaqPrX5Pvg5eP8eX45k/J2LGMtuZekYqMqLNdyFmhHnTPZKj
19tBf1IXVhDdI6LkAWELs2d17tA2mev0aOtcwaWHv4I73uuSpeU52X8dgSkHiTq9
QxqB2nQ0rAFHG8qlfoQpH/ReHEhBq9fPKNydUbzLSp1PrUmx2nMu1x8jOz3phSbD
Bj5qS7hACpeXtsOTBUmIRIVAzM+sPporjkYVsRnHMyRmKnfXC1Cb2k2udpIbsC6n
wYdlH8pQybVzRvF8L+diVD7u+PVR6sP7NmZlKLfjiittd390LplGKf+2ydwz9Jmt
jhifbOKDmeTyVL11AupQusjNuxAVh6x/I/luoaebRRUkdFtlC9pW5H/0mtRYX7CR
bcf4D9OUsJYdlDha60cSjplW+AeVjiGNwWjfPZUFqhzHgxMRgOSa9+wI4G4for2+
HQns1AGhAnTgmZavCD+VjYlX0HobZCTFoy91PExgLK/ZRbnPIurYjaryuW/+u4GQ
yrRKwBdCd7wHp0L7yzTYBc1tQM8Sz9EvTXAJ/Rztn/s+dFWwHJLiuL7PWprDD52v
k6X4IL8s3atClXd7AOtFq54ofcLzXIIQG/kdBsnI6CPRRWad9ul7tOSQErONQDS0
Et4SCJL1RidfJZg51ezBVEedWuScMmKEM1NmlPYhsE7ubq0HW5Cg1q4HwyxMGFDr
IDjcGRt9EdCSkFJ/nKs1jwF2e9+JNM7svaG9SrsO/GlhWut8Y4FdiZ8stSBtm217
2bwGd7jJxyJtKCTHtyqZpAvD6SK8zIj5JkScttUlpR3uIQfKOJ0kUH0whF0ITUqG
7wIT4nYKtkZwozASqfl3Cz8xAONX1H/dUQu8wxvDrhjufZjJFm/HTc1QvtUO1Kk7
yaenylmours+arbYW71cvFmEeJyc9nsaCTmmtS1ORiOtk/zqezUeq3apnJ6uHY0D
xBR/iuv+vWCfulG09a2rjW/UsMAehHLNVzDdre1yQh+pA4w6109j9fytigpOlMCm
XuAzC00pIeeXUFFvvkvR9l9a+dkQZeW88o2EFVQKVDiAE0KmXf9AAszaov83fWEL
Fz3kx1OXLzWy3F/1oE2yr4GfGlMMZAUHj9K6WBtxPrGk2/cEX60pejV5rq4pC9rl
8HB7/H9Er97z4B7SQy3lufoKU/KRbHLUDUnt289bkbvdTkNVbr2ca64c/jL207D/
akqGzxBRNTSbfbNSTdSZ2rEZWGLGIsYk0k8d/dBXlKAtjVSB8IbwMB+qMl3K9LBi
n5nSEljSA+nm49jFPCB1YWvyOSYggtuO836gadW6zfKMuwqphPH3aOLmSffs+Wm8
8wEazJIMSxa4LR41VUUIQxS0fZY8rAkS0eUrFr7d66EAfgmEGyoBpuileMOIsPnp
8tVj08/3KF5BREPLAMVV8ILeAFXGkjW/wElyNTJL1xuaNBZD1IC5JLUNV3msGn8u
zg7mDguDCQptv/ssKP2YVP6T9ob0Ozb8+UnUhwXZeogAZj4Jfeg6uwPrnIm+HEDB
Bwnmrtanv84zAgQHlGJZYazhshKEaoqJfA9NHfAVxaPTWf1tRxQ6+4CxOuVxyQwJ
CBWAzt3sC/33uqlyZUu5M3/yCePpxifoOkz9tiojhwsRm1Wr8G1SkwyV4EZAlbn8
+cmqOzIm4nWiZlkOMePWEnhU2c6bEIqz8Uz4QH0f7ZrlglqNg5/EB3JqrbvgSb+B
tl0NnU96c4T713nfF0CB+457D1r/nbLCsFd69YiynEz9ExEF5VDpPiuJttD3IqVJ
VCvz+5bPpN7sD4MvE/CTZVOmMAswTo8iTVylRWx90eFbscc99UXmwBwIv3f5UHX5
7ot87kT3BAzK7ZBkXjEB2XyVJClN0ZGwx+XaRk9Es5cU/8Ht3qlVclbleq99K5WL
SNXPoHElxEB6Fxxo6j/kPvFEC61/kZ/VF65ZhJAgSZ/F3a61SpwM7QmlQyEsfe6J
Db2gQ9OPv6EJmA7BGO+3kopbXUEY2p7Z96lx9HD338FAb2Ot+pZeWg15t5BARVkG
zfg9CFRbtOolh9rpLQeIzkC/NM6FdQ++B0GG9Rw59D5XonFeaMQKv1wMfpagQZNh
lDo9+doS27WqjIcBBP4zj6R3KLIRj2afChhLcjN4cdyBppyaIjj7hoQNpPJj3AwY
EeJMBbVdgK74Rnt9o6lSYgzuhV1o2u1X1FgpAWqgXXICwpdBns76NWIDmOcjziA4
nJ6a606QdJzqf8ADxlYVb5e97YIgAiN2X+8rIisqjm98RZP1DTcLP69FEsVLBGDW
MJKWnrnS0blumCISfu61nflGIaUSwwyCy6ugBVyPZszpR7p/acpZ3k1Y9IkePMHD
JIocUwv5hluCt74u9gM9ztpzKLO0SkctaCN+lJTNclk2IHP5T/P0lcUd5FBH0w4S
kd7D0fES+7XVOfJOWECD1ZPBHaJhiTZSfeN3Yfsy1e6lKE61Lfj8RW2p6MYv0Vm4
KXEdJ9DERseIr6JpGoJYv1WgVGnElLCeP5t8PzhWyqJwfpMnTPmj2Ooo6mXCf4IS
qdBlJ7aBzUl/Ei3vNrDB/g0rHnkpmwnrBp9ax6ZKPGabgjX8o+a0TltcqQjuMnoI
2cRpAGUiKuPoPKCl+MTEtyv+fpXh5XeweZCrehMne+JdV77m/t5QlZoioOhzfL8q
15m3HD2ArI7SDwAnWOxeyMszEaYvhIh0DfdxpJfEKUgra2J2frudNW+NNUlv13wi
brzf4yPn+iCoGX3q9oElS1q7LlIAEYUy7Dux93h4sywTHOYw4jrq6FzHi+ZPtoab
e+GD/KGhOYipei89OESCntJzDyHs6rPz+uajL54gV19K4SiaihX4I+6DsntFit0b
4/fyr7+hbye2yi+YZCbXNwtizfXsXPWF7we18F4x/sw+dq76K9PcNlHacn794z1j
XJeIRaAv/e37xL9CFoS9enLIEAjoPugn7XAGXikrZHkFTnwyIxP41lFicVXOpvCj
iLbKqcR5MUszvTwSlkvnOmx6FPgjTijK2aW9HPSsSgsXxiMXzHZmlDIGKmYqiZ/A
6D+SBI+8P1V8IHB2OwAPqxUdrTJCFaM8zxgr/MDXlC90yVQ53vUXfsYMQffDBFki
1LxAz+3hyuF4mIDbpy0SckXiaplhkcBDPWD2g5cjnE/LeYr/wg6mh/nsBwIxM1U8
zFm/S+WGR2h5BkrUli2fiN3XgXiDuofkd69+OAj4roZCfD/lMkPKB7GMmSPH9VGk
03A7smBUWaRwPvr4pht93fr7d3/+RZXUroQvjFLe4JuiLhGh+rM1GcbuItz3FU7y
ORYrYKFSgmKm4hMLs+U9+mGL5dT97k9wXJ0BOrBmo9bCWBqL1BrJ/mzgwJNZNuLd
WNymM0/5j2MM/qwGIGbOp25V0auTDJqhR6SRsDcBC54e/CqCPw0lbjCiKOhiiV02
0wl5T7tMb4eXXKlsjy902KJ7SiWY9FadNDE2CA2cQr472HcuduK0z0v38E1cyW93
NTOVx/vyr1IlUxLKVrMQlIlRlMoD0UClCddHNwZNAueL9BhXt6mQug+9XitaP0G5
um7f16JBAzZ+03CUa32o2wBjO+/D5m5S0zbWp9+zx8RVhHEm7OU+LVg2ir6PLVDx
mErCIx6ix+MHK9yGUlUYbKMREInEgZKs3UYYbqcuMB66UcFsszckBH0xkO8A9CK0
thh32a2/c7XMIt2SznXh10FtyZ6AuE8Fh7tLNBtjm3s98SMLlBLeLQ+1R7uMjjfB
9oYyeVe/GeMkWkat79C62wOJHX61F7WqB7IHbFm89lAcmiuIJ9pJcNg+MZODYOgL
pHhbOW0N8dGz5nEWvWKg33ZEgQslk77a6ZYlsVzgQ0ma0dWWFAANmb/8d3X/dzGy
pf5iyIRqQ9jKT5lRGj08davpVPnwKAv/ZKD95b8efgHl/bknR7ASD5gp1RpkxRW6
0lGNYZiB8QxyhHrfyxS0SO/ECBdjPMh/wdxXX2/47qFOc8Z0jIH5VqOiSbs2TFWd
cUp5Kl3rovcckslYoN2C7mvCjqEDMHdOSAIh4kObX7vLvZXi7K7xjuE9bu0QVHCb
wDPpzbfYdwAIiw9QD2Pda3KSThPBLBfB/ai8nBEa0cvKGzkFw5dRaQquwQOKRIyX
iN/lo/wTh8GsNPgMHm3T4uKf+cbC9gmot1Hk+yqvNd+Acy8EhJOTtV+c3ApBzbG7
ANDm3HidI5WVWpGNr7KIcgU+oVOu43HZY1LzaPIVmrM7+IfTy3GHFf7jIvuveDvb
9HltxghyhTzDuSx1RMdZo7GoEvC5CMFm8+LHVUqW/qJigwRw5kE0WLVA5C0IwG2F
b1Ga0q/7FESq8tv/3YmLWahu3WPyOW38pwHQVbIysyEdBnaioIiUgFrgdxMa5NOE
tzju1fT4U1DoPEm8v6YmOysn+lvJwSrhyypGz6QHz7Gc17Q+vWCe8rsHhDc3yMUW
B2v09zoHeitae1sThKPsOLDEhVNd8eTLgJIndI+Xq7NLxxGzkzVuUseYVgJRPqf+
TtNHrTx3AV7JKij937N0VFmQrlesPkJVhkbe8yLXAU2Rjmk3jklEKaz9xSZueXE4
jsjTAh0zJvA1DPT/7P5Lo+miEscABlVwRFcC95HCGvRJfNVQbu/dCnGNsjDeoPRL
7fK9opfijWkr/UjfsBPdxPLd7FSSIrnOG2k6JwJriIGX2GxN6483tLlpWP+w0Cij
KIoW//ZJzts8dK1cXCGe+2viPDW560twbbLSznREImpmxXURkeSRCNnDtN5qNHoo
SeKCU/RxebybrC5dLOUuqEQK8WNHY5jtIpw4yKuzCyzA9EwqF4mqq8GNgeXC7h50
uXJ2u2bAaPlBm0nRdUms8ann04q+Vq9BWvm8AiY2LVPPxc4oheHRM8EE59CVTM69
igTVrVyDN89PaD2uGovDpL/rsb3QL9FOh0r9TFeD2SkQVr9zrV81EA7jXeTLgAtH
xmkJvgFW7yfpAgRP3TDMd0jAp5dikBCpwTe2IA+ZzW8PT5fFUA6AO+Uvz2flT8Zb
jAJemE5jHud5ZCEvq8sk64B/In3UBWNoxMuKIRoidEmaiTOYgGVSTEdrty7EAUrb
bHX38tlxQCMs5Uu14xsuHPYBRFNbFtS4mNMKpdtX4K8/LapKtbXdUSTrMLtVsi+T
KrlyiJuk+pkLGydXJ2DR6reaeqSFJWOMvtgle3PH1RX7EXEwtpEwAS+hcBLKlGIy
VESq8twbam5geEcYmm9GwNsyRF2zV2jM/E2wLPBms/h597QrK8IwihGKF5cPqL2u
JeE0esi8r2mhDivRqiKVUe0Gocw4hH2+ly2afnfxDYtbs3CZnn9Y4VXXubbpUSzj
gHWL2ytV/Qxb35VwTYQsSb6/emLzJXWDX3WYMtEJ2+lemWyx8RnC7zIluMIw9T9K
DdKg/V2I6dHZ5nnILY4r8hHN5ydVK+2Z7voq25Vk0y7ZqfXunbXdj/2zdUFquphk
R6gISekPW6Zc8YBi4JOkBXXAcxJfKvZSG8VLwvhjRHb40yYUIDe6+p4woTRxAxRJ
fN6COMfQGPzNwZNIl028OljokD+hGyB3H2+5j9eMahvU9GSMXBfCDwvNQxu97Iol
nmeV25OzjmnowiM8/XGJOCoStJSSnYzwRas7eF4RoKCDv7qT22UV91s894YmbZXr
8OCyLSSZWpXkQjBEOV7JgGn0K2HwO+Wui6nLlqlDbbZyDck28VjujoseEdK+Qrrp
7Qy7Fjg3avPMS4Xm5DIG+i5o3mih6EixDw5Ly9x1N9dj1OHhcU2nw7MYMrNqGJ9L
w5KDxv1mK7ndXBSlIXfwBDZw+PDyYRnh4eCQ9y2dQoL1QCyr4LG+2BwVO8iJfmKS
ea5hDzRgeCeVPX4JonooPCTXmSZHjglQgDaQhnflUgK/GqiGMB1WGg0rPdiV+VY7
2LBcDo5rByvJ36Ga/HlZgOhc4XF4K/8ieMHb7mKbjv9GVt6nNyMnVYQTkNhew5sO
f+RzYYR7jItBfPuwiVLFLZyXzL6sSwN6O9vt/ZDScU1iK/JleuXoXQStZ2PagvUB
nwgPH/e08KUoJYAOF7PNlIxljJB2EowvfCPg1lsRqmu7EGha7jCFlcXXcyhCgEp+
2rB31LaPr89FZH7ojqufld6Dt7Ty59hc2N19aTFfo0x2MtDyg+yWiNPrrGRdo8jg
cGbHxp2iSVg3Z+1+gvQ2Eq6mGXwMcDGTLqh3INJ7KHMGF2JgCmI0XRw6BVEJCZiS
6UpwfDANihATqRbhxtD8MuBwYtUBeyH3X0haQe48ZfUH4wCtn+3vr1vgl+ZqdOy8
JaxPZFvmJT4Oz8izhcutMM0artmn802JgyVmqvond4fC4Ek0Dw6ZEvsrrRBb+oRg
sbigC7RYg4SRwJViF5WwEgAJLpm/uqvaeDGS+vMAXvgD3Y+gYuZ0Z5sKrxxpVxje
BQMhH1kjo3EOHrmLMC+61X/UzaJ8JEPZyu6cjTaX4fUIraq7xeZBjh4GeFzcPqYI
UChxz4ZBSvMTIH4uHxNw2HLGxgcBq8d/kq33bUCdEDpyg2Pu+WbRY6jBqroKLUNj
SY/nS1Q3nhYnCqScwCJX2Iuvrz1yBE/VTie609vQXw9w0nVDvAbFRdHGnJwuWEHT
7PsW5DDfyageAhX+JxHuUkLRBTdH6x8B7DNa2Wb03BMrGkIeUZR+ASxQ3YXdsdGx
l3R+0/SK4zpg0b5I11haTyL5HHwOir/BhO1Pz6geGNZKi/6mDkuBBLdX8PCf4UuD
TXw9xoNGB+JMABDUO5pKvPreYtih7Zgyvm867Kb+anLnjmsZwEeM3o1QqihTRvx8
oSzJaia7IUNfO399Pc7hQn1sV3zkXifX5lN0dNVQxOGa7uwasYesTTZla4P3ixly
bl+Pp87NnIo2BiGMh9shWwY3TtHwgHn3nYN8bGAU/gtElvhH1DOO5VIrzDA5sa9t
fPK086UR6cilpavFZFuMaxHkXrY7xQpywuMul15KmfJRU2gNw6+vRXt70avkLWX8
wexOcMCUXT1WoPs6q/zkwWw6tH2AyDceSaOm85XqwGtHTMssUCasBtdAeN6fbZNJ
5lymIgKdI71wDOZ2v7AC0O/2vZTb7MREitbnIkcHy1i0ctzwkzP3bMDo8k0j5U2T
Fgg9a3NRtsKEP/MrD3Nj3eE+Ir6AqCcz0Ovj5rV3SEghAtQAkypTo1ww6/vU3clN
43Z1ucyYmKtO+XG8hNgo6E1L6WfRy2llgGaFiZPVbnGHfBPTaGYcj/XI35ZOP4bf
Z4AhZtqR4GTDO4wWQ9FsjIV6xJ7gzt3vhWXn61O7TxNWL1Hwaqq6LCYoKK2Dnez0
+ZKgvEWV/Y211pzXXvqAW6Ysr9N2mUN/u/G8yvTRHT5or14v2y+xE1zvsE7wMzwg
RKTeDCJqhrxzj75pEijH5aA6k3y943wjVduw+6V/ms4fJ8ImRkxuTzynCUsZDg1h
ga6UQSSkucJLgEYEf1ezErMNO3f4/KyAWlpFQ2q5HDJQPWmqfiWjvou3if/GFtxC
jK56k/qUkC1xY3qgr4eK1GeweXAy0mFbS38E8m3V8e8D5YyRLi/WGzMsF2Z37NMz
qdfN5foZKyCh56ro+VRIcKV1N9VJpNehHb0S7ZIKseDTNxjHtSxHp7wcdku6Hgjn
ydJBS+2MTSIcNcn2LMiL9dYlntVIIavmNXyEOYOKAHGs4W4McWIwnkpiaCdlsl8D
b90p0Nms/vY7GUKSsRHR5SUY7NlrcP1OuEqOK9688uKhxEXKw8O+xByqsuibWVSS
8+guUDpHYCLeV4pI0n/VsOAdjLYgX4f3xmKU+ZsZ3oi9Auy4Yyys+sHEGCgi+A3N
cvRb04f/LhnmcE2bThuWJC2pAqzaUL+WbRc9+if4HcfMAUp1a4x4kIOiazEJC8tX
G8WQ3ipu5Oodgj9rtGJvmZg3oXryU9K3ykUch7+ZraenVGumMzj5YoeQnHgtDvha
RcSMk9Pfq/pmAm6Fz5A5o31U/4qcVn3cdCa9gLrlerW4eV2IxTAXPVBmQT0GZMLO
Ca7XHKRCGBTdOFm8XOdN1eua5tOyHebwxwvYbnN1I7A/YC1IL+dn2xmB4qAtDa3b
HW9AIULVx62+dyF0ifNsmdh2St3qdL1eaP17+scXrNXlVsqajoYCUwwEBpg7JNAk
9F/DODUZTtvHlOeVqt4p2uY1iYJo1zT4ONd0L3wUMfELoGki1Ix7Z0RLdziCwJTx
LHTBZWncVfguLcjo3g0ph1I4ffC2DaRy1Ua0ZVsBHp4m79z6O2VCAkiKsMpdWZYW
ZEy6X03K/CWNUJ6ffCzOYldSFkSb8/R9QDM/wgE11Gt0sxu9BWUUHOhpcu5p4nmY
RqKQA6nbItDiSe1Jf4YX+4MaJrrTe1/XV0QCKff/IypxMUao49aEQaczO6jNAv1T
jV9isYqKsUIwfWuZzPl2/bhtlsh1orG0B7Cv0JXZTpG9fCzXRglzFUTYpD2eKPt5
aPSlgYghL4yrW35ZzCYJlQM78NGXh+5+HBW/ShawJFs8BfXeek5vutF0NolSbGDG
qJDx1FYG2wRR6u+pyFX71jfqVCNZz8BEN+v1ck00K5vTosLavvxM0gBv1de/h7jr
N91SYu8gzz3u/qEpdsnwPWqzPygGF482NpY+2yWI7HVZNZGiqeQIhPJ46UiHAI1w
QMYO3xejc2gMArrzF3Ou813H3fnYZZ6TFZa1avyU4H8NBzifH6jdRjzAOIW2vHxF
sJHkSsf4UqJs3oEH8I2psNOhjJrJLqVOOFQuubDaw3gAyzQDqkNCmQ0W0Vemnpdy
GOY02Vu8RAHa8FVu2dBSJjYw8a1ahvDKpVDc/uLcOp7pMB8hD1a5FfnfImj6pCPz
xEge3ldGO7CtYEqBcPrHvI5mp90KS4oKtctfve041kXs1qn5nngzSuEi8JcrcFB7
qfFujs8LIQG2131r72AFqMc8cLCMbsJKT1RHPx0hv5O6f8qBXQ0YpMNwbi23rpkx
oaTovrE/a02kX/GOcPaK/UYrPJ4pYEPwCXDWXtB4MDWrEPjfh0La/QsjJyWEsVZw
ThecRhD+16HFXuUnphRMl/3Q7sZx43uemslLdbiqxZlDEYg5I+IQnsDd/gzTtFJY
7IbvQ6kSOfLNoTUmE9ignj73y4paYxyceh4yw5LSGIjVrHyy+J2XR36+nSKWnOcV
DEP/C96Yh0melv9GGQGxASS1F8l/7iSIewuNz+drTSTqzM7MUv6QcA92Nw3TNUhr
nkznn8KYvdMd5PG6PCe8CZg6MFeDmqXaqplmLr7Y/sDdFeW3PtuNaYvjdih/r/Cs
AzGTZOig8NLKX3Aao1rUmKTBEuB3pDUDpJpmdOpoHH6KXoYdJFc+NGjKUGstXAuI
ERBMgWj59Myxd8dRiwnA8oN0Pm++DEbHiy0N55W7GhM3sxNS8n18CbSYxXnd66J3
Io+VWRULVL7uDMjKDfj2CtyQRwoRVSZpjgjDoJ8D5yeGqMbGEi2nRLolvWi5P/Yj
jeVqO5c6TH3+xYI3D57mJCHUoziwYRHnjd5FhrWODdEaAouODewGqcCxgTH+UlC1
Dxdb6JwIwp6TtjbRQW4rhcW6Yi10K1Y4f6TYLQrGop8xVfw4Qn7q1NFKmX+G1Lv6
T2Xbj9G4BAwf201sR4LcIPxf39JViaCeoCu1nngL6i7FYSsAbGMSGSKEuTSoDGc1
KAts0OIaeM1vp5aanoQsFP0hs6tc9GAX8cGMcgANWTB6jFGN98JYGbpLMS/dwPMg
UgPgS9iZTeoLCbMIyxRTpXVpBhgX5+/NOW5Pipu2YgBZi80FMyOgs4Y0n6cEe1pE
x0xdx6+TZZufJmhzW6GI0vNbCk6ppRDHsGQuPzXEQ85D8CAqE+4OMncSPFsv0mAi
iTtzk7rVOAokTw29nWnpMqkIOr6kKwYAWQmbi7quexCJH2ns+9e0CC+EIoya0DQ0
gQBjpwvCmffF1zzJcVqHofNeSbo0cyB5V8vy+HrM/oPM0Aj+rsogSggzyDnqdQLw
RgXW9iCI/PQ7e/kcKNOktCWONObeU7mCGCwEOyT/k4tOO3dFpVG7trfJBNjw9p/J
6OHP4D9wRhNKtNfAZRUXigzPkmb0CApMxYE691nb2yrCwP67ML8JDDntAkkj18wM
1qlYPN3hhl0pIkvTBUKRYnOFJrt5htN8diCHZYf7dmzx8Mw1+jcO7pz2IvbnqQXI
M7iffwSleJWOX17ARIADvXbeoSyAjWwI3CTQwVzOhipasNEPJgLj48zcQ62znS1T
1H5nyt8hg6ojRCM12P0TVu/KMQ+RhL6pIg4/A/D66YLywEQ3wpZ7XYw129Y91YIi
1d3t4VR5mN87+CLRXDnfcwYdiJG96OJn88xPzEld56LafK53Ayo3nnSmz6tHjaOB
EcGxs2VEA1L+JBospCi6IeE6WEOgA2OkE3/xDas/khGecRo+h8XvyH4/NEfzOGEc
YRbeivQiH/gSSLMux2u4BF5FcDbkWivQJUbuOWUDVoCQWpLpjXGFMfZnMllWIt8B
xCh+YxuD1/3ECRVswCgfflHky5SukFXZedmODEP9+mNlT4spLQLYNzGJ5bKS6NOz
q9oxWXfxXzwOV1Isu41iU4+76tHzcPr4rmezMXYiJjtQCGFGYnee4Aa5yawSt0Js
IjUL/5hejTT8n0idlQji7VMca1CzIntMgN0T2p+V3XDZESr80TfVajyqssrTZqV8
rvpbtK86CRJOAQVfj+aH1D/03rCl2J6LaEn8wfJmmtvF95U0AaAAc0VeAqZRyhLX
9dn7FJZnhDzTkw1KOc8Z31dTZtD4ieLh1bF2L6xGB3V67RN6zz8gTYO1P2VDbDtL
17/uWhyF7eo0DoUD5rOLa5RE/RF0iMANIDlcCW8a1PfkVYtOa4e2+bYR4OuIzXSC
GFOMwvtoh4mnTdol2C23x7+yjBTKd7w3UvVVZVvGPhFhZyN8wbjFkIhTg3beXuj9
0KwgjOzfDlmG4qIs34XddPHTrlafjtCYF7XsNO8ojjqmf6lIjK6MNbx9V9Tud97O
pdDUmfLv5d/l18Ca52/V1KJP53hlERUxLG33ehFmpjIcgisIaABFYQ7sgQYlneNw
vfxyAk/CQrUjeoOKbmPTkHckicSJ1JJtkXPxZgWZ7z23njox8LUwbFfdNhVUXgGQ
57vPleokgoiwhnACXzAclTp13WTJHrC/YNh1fT2wnxzKDhUQz+NrFGygWSBHZYHc
gw24ySNrfTTB4HFp8OHpqg4IiKAnW1BF21hdO8reBdsvlZtuvz8rIADazVOYNixY
W6e9JbCl7FERZHFuk7f8hUaMCXuYbQqThlF81jRpXuwSJHEkZRXg1THfP8OC8FLD
n1fnRuGk8qG49sKNJq8WHM0N1eBy6wEYuUY/WuK5xtPshGQkdOYJ5+0mlPMNoWvC
xs1OWtdTNWE0/O4bOD6aukCj+kBfo6AZnRZKPWF4frSKT8YPsFbODnBW0e4EE4dk
gDgrekQCMpj7GIa/UpDbQBZxQZZ1wCmYTNiNrFWkG8/fieH1sDfNTsfSt2jZeX6A
oLNLtOWtc6s2kSHlwf8LznCwup4sks/+34gmvuWJ2SjB+2d4cVNCPlwHmXKzDl8R
3Wsa06vUTAcwhamNwdMJY2StNnAk0kMAzoXTR8ALMc+SJyxdBmhqByk6gweoZq0r
G/eH20DakJYM4Xn7zi4Z4UZx5GeqsDncfMketFmZAKc2VWxGQkMbH9Ty8qS2eOEu
eWn1058RUncNovJpnA0lBEXIwPoBxSWHmQkzeQM95eaqQWw23k3Eo+VC2HDdACmh
l3uFap+9HAJsBzSLGZCDRYCH4gd+mP8TKaFdW78mVGqhy6Te06GBxSHQWLJUTJPt
4yKyvaigJK2nXuW/KHYMFn7ookFJQa8hCPYASQirwiOIGQhdYrKHSd0HzqF0E0aw
zErcd5P1m7yGyLFGvdAkKYpfa8tO2hZY5K8hV3XzF4HSC6eIKthYOK1xYb+bHjTS
hLQJoKct1dryL9j1a0ibQlO4xI57pbG0pBnkcgdTbTpqyRCZqPM9a4ivjD8KA1g8
dtAtrvrON2eL5GSfl/J4CDhEDF8lLCcecY8Ozv569cqCQ6krIvR0jRv7CPJfdqmr
sUIj6X3952GEn6ElJW2vV02MC8htLKgCHbLKckx4FPPMLT649Kl0ErAYu+I6au+b
7D4bydqvbUOMMj5FuiXdBbYF6SmWVWzq1fiOk6vtA78hLI5fZOoxfB/u1mDwVeI9
MLKNyldDBLH4KBXXPCpYeTeVxvM69QGTXlfe6oQuvJeyA/PXzxmXjnu8onwUkAWr
JmjI2fPxcIL1fM00hhXU4At//DSk7h8Rp0ypf6FzrXEZOv5S0aH/QSbPhuWMVQSp
6+r52n3KD4PmefAw/9rIfLPTlEibLW4JyhJdcNFyPS5794VOPAz6513sKbx6xumF
4EL0pfBYEuzbYytdm85S4sW+BHQF9gZf0msp6s2e1HPvFGQVh20rF/o7DwT3qdiB
TxNtN+bDpDNashcr0n4hNl4ITxWlyzOX3Vth471xSDydy2pvsd/epM1/L40gCfNp
gRNhw+QCm9zUkHykxmdVIrmKABJIq9MHUkvbNLocppnMsHvEI7rRtdUXeKB2om1H
6ZsUTQJ9s/0rc64iOfBC+mncOISBInhKBHZ5Tbqez+lbCSGJGBPTUDJAH43zxR3Y
AOwvWbyKWjo+0boovnUivRE5F8DDQ27V74K1A9Lt1PPCFqIYq7BkXohypoiPqX1+
I99WoKpvS8RxR+07sJ2dQvqRbglagjPUmf/xxfJIm56P8WajoUZn2IUD12Iypeli
ZhUOHsmixmPSyKwXzs6hKIzlzMY7XfxccM9+qULRw85u1ZF1TM8t2d2zGmB0YsiQ
jDHdtpYbdp0brcPKhmOXFuCSVZ+VkgxBdlSqP962DKY28PlARkBVMiV2bdOT7yGP
356dVjFV6X4DwKmQnuMRiLDInIowivC8oLDk9F/ogTCphZyJ+h2TFKRsNLPJC8RG
U2AUpJIqfHn+i83rjlLAefFKIv2VtC0NPpnn4osZZ0BTmLX0vx97eHhtHDGY1OoF
ZZMB28y6jZK+BmONetW6K0DAXWChQ+i2JSAbgPnmUIwdq4xpU8IC7+FIz2/6jRcj
0jIF5uTUHSVMqXF3SFqxdxD61+Y4Nho3D1yXjXT176JzjwAu/Fk6y4n82f5q4M41
3/Afr9gJGthZsW10I2auBmXYbOz7eF5AgqEcVp7+93qHWQCYY+TF6BNQQAMHDWbp
Nh499jkaLnslbA6qc20DXgEMDNyiIAADqE3h1YvW636Rvq1u4iWXJUXI3tMz8JSR
+tI7J6eVzNt3Wrnm/KGk1IGHsBo/PdV6zCeBvsyQ1Sr2Mq18UN0kIVEPJ2nh5KIk
s9nNCTKzwTx8kz/MOwOvMlD73RntWPmWA6pCkAnHkRiGM8u+/xtf9auyg/q1rCMd
I2Ag6B/UIBMzZfbSBtLdkJU21Vk8dcxDVq/IwGrEAjuBjEYsUcx89mgq86qewz9E
56uFq8poeBBahlsu/IRnyL9pO3mzCyMv+bowPSRIYn1S6Z8pfUCpoP4MHwup8PXq
Ki4O0qSYlK9g4Nnp27EhvEGGKq7BN1Qa4403yG8dO2irQB9Drb5P7gyQU4H0ndke
PeuHEzTLqeMY9BKzQoC8uhpnCfrLj2aAvmo6TP2r1k/oQSnndxpBDaP9FPG8NDY2
nfeUvx4+gFBvok7C/iIXmlUUPiQPgxnKx+6rLbKnEjP1Slv/9iJu3wpelI9reDRN
vMHU1R1evdcEDAYnRQv+d3YhDZLlB2OjiqzCkJCuEgRPNtiWBHImMjr+HJPyXLmk
pIKOvufFPkK/Tc1bGbldLolNBX95W5vIfVxkBS2VYrJqc/lDwcmaCiGviz4Dl53w
x/qWHjHCQA8yMSI1DgeOxRIBNHnhmshO/MTSyMxxz9f2C9au4tGcz4M735Ty1W2v
kY4iD5DLNgoD9nC4r1+etSq8s8vPfzYfU4UO/YJmc0c7eYnhMZONBl/nuAoQ7wo1
wsbBeDMF5MdE6w7T0mSUZ31BU1orF4nEW6vNkbZsLs4TXVMDOSLnQrNEggFpwKUG
WbNcvm1hyc/xuZqzYy9Efj/IY6u+7EKIAN/Hjf33RTJ5OK+YDgNF4CY+0em2tAFX
oeoAx6GclGbJWRVbFBsmzXIBncYG1f9wR9+7DB6NrQww3jGhbcr7XjtSn0Hy2kUd
kxij9TwQUEmoK49bOzW8XTTUm9NusdNNAYsG8fuUOEKsTxgW5Aq1hj5BGHWZrqqu
CG3jGfVd7h1tA7KMpq0kwrC5sXHkOF+bUa/ER8TEzv6QJhc1+MhqoUoENSrMfpql
+nJHzMXvgeKms19ROUfY0xYWTiA82TdJbm5mIRXuAGPLKe2AUmq5XdSrC+fgAGTm
XtGL2cjUk9YwrwJc6ELDU+g96KsIdwhGEcadxuP+SS8fuqNFa1BAjjsTHdwQq41t
pI4FKL900W3F02HuqxskAtLVZAioDl09qHwjxGRayJasJfIrNEyvzqJDat7xEHJj
4hTwalChK226OT9la7HCssXXVv/YNM4FLSUkipYVBghtgKJWumAlzaZmGtaKvZ1d
Qg5hwba/1MSPsoKYpNIcrtuyCI0GQ6u4rkVGFig2Rjaa3ylVNuI1Mn28Gh4aiaLv
iHQ4wdQn9bWljvh4AlxU/Mzol9YFD1nkQ7KMJwwP1hxdZYJpZR3f6g9wCyV6VcWu
ajigf0YVbADHxvzp0MG6NfnSe0s0KIlkqkjsZuCQKquA5nIuVviBMPwydj4GPwGn
ytavjlCfv81CtIhgGMiXriFaWC3aVqzKKHpRGN368GdFaiopiWzPXS1+8yHeaxXW
G+1wDA5cX73XR8ldD32h23+iz4B1Zp+YQWSkVJ9WVfASZ/Wn6Sk+rfvcp9pCWH3r
qo0C2BqRu1cdkLEisijITUxHOwZm68qgwZ/hhce2poVcYp9103bKoDpUEHFjM4dq
+m2R3TjhBf6oLyOCFqSfJAXWAslFYobMMZ2pyLyVSK2noz68A1EF/yd5bQ8xVMHq
+rXfykSApwE7VSrcdK7ExdpEDiOW6vEyYsCrACtepRm4g4LpFOP/Pgx4J8fgPoWu
aeTPRbTJ1UQ3wRTB31C/KTVLP7sDI6YeK3BZGGoF8PLYenkiyazPuj+DdDR65o8H
3gxtvB9ynoqo2EXZMK3Er6T1+GC/21n7VMxlngrPUpi1Yci2Yzs+FsxkAJSic2CB
sua25aZueUg8fBkJhHrcHlTIL/3/Re1JlpRwPK8oEX7IfPO3pdYothoQI2wsmLbu
d4lpqJg0Cdti2BmkDut9L7MfN0MnsQUDQrwwrtnyUStCbQxScXAbjfc4H5oqcOZj
kEjG1++yaivjbijzAOB1k6cfQuQHgOj4L6mcOmMMc40gDLW8mMkzwSqX0d2onWhO
xGCMKEQHxCUD2C9w3l7IJEjHFEBGw8E7JGMBeCtFn0rdfcuA2ENQ8TAlcFYzORJW
ALyT2ZVx9Ih5LbswfdljLENxb8j0r5oQs6cwGFmqJB0kXcLv/FY2ABkhoiN92pqW
wGmr/scc15kdrFeUxNhs8HDelCSv91+0J+vwjUhT5Be+tIP16gxhqUcblBJSAPW+
9n6Ka48yjy4dNI0Df16EbmCNWeQgl6XSa/1Z+GmkGkFMSQgxEuiPNwRoS8/asB1N
gVNCGiNMRqCkM+hoSHgrqla7rQHH+93mJmeh4Av5aLVEzmD/zT04m+T0eF3RQxji
Q8S8Er1lNthvAE686HTr7c0f/KBYXEN5UMxED7vqQZD7iaiD2tr440I4Pdn+TDvn
h23hvZy99Ha+PgzTTmu/ZiKlJY+aYUXnBeTA7Ufm7aIgTf6CFTDkZg/5cFhqV7mM
g6z9XGowMYnNUwEQmJh6PRevLVmpHeNtmcHY+HaFaWAyHFdlrCtLd5+ktDrREg+J
cGEzN3LzNUHs/4tSorcrubinc4D504uRFo2wRLjg1pTXHhczrjcW0iOWYJaKq6se
uA3MpDx5gYZqk/+CZ8t7e4OL+dvMn0N7CRoNcPzQM/IUn/a55KYKp2ZC//sJLVJj
3Ql0Bn1DoIoIwWYYJ2Z0TAuJ1w8URGGlp6FDYjuMgd+p+bJvtdXy7fwAFK74sU6O
pus5Kt+yS0PE59/bBnWZd8pzWWq+zWWOysI1SCqyAKwRipcIOIOrSkY2um+tTx6O
CszHLPZJ64uAIMzKIp5nigeN6/EL3VOLxF9ttW5rQKIcTqughm1ZLf/3g6vOQSEt
28PEPxisc7Tlr3zsFKTRDN0HGeWQe1qAr1U87maBWvfFRjcX2BV0gQHMtWTV4snT
+4KXzLi25YPfzW7Z2ymditfi5enZ5pGzbpNZSyNtjUlxFLUTpFvQl3mZe9b4qEUO
iMbJAwChxcmu+nYKkzYWuMgtwHkhVZOmEbw/9pFN+OO7LnsD+YFDGQMN6pOvVv5l
T1oW1txseWLh1cuGT7DIoxZG/vRKyECjMgUHwXRnybqe9OzDGLhlpz2DT+0YBgqv
aplxqhMSczvwhin4XAz6rNRp5sBtxJjmA9Tqlu/U6rjX6NoK5plQEnCI/graXVdm
ZAJxAioifU+iaD2pEaHNvprztblETSFanazt5ky0a5xennS7ZVv/1+ocBuiFddtD
xRSq0LgjuPgmkNQywk7dn5rEZ4CAPUc9BhQK+Hp5kDiRgAgO4CStQ5oQ8ooiJXVk
N+Gg4uiT8ClThmQRx4fqlXtfBJ+FqWliAEOORV4eyG7t2VYWH2Pnbh2Wv3/jPAu3
yxCFYevJPSA2fr3tQvGRfuee6LDmpm2qT9axwM1ALWHEAPLcgcvvuXvVtWgJ1y9o
KbyC3+HNWnF3rOmMZNkhCuuSKs70f/NFQ1dKg9Id+gVmnsxszHo3ha6uZSwAtJdk
Dbv/VeFDhYlTVO4MS7GJgZ+yE5F/hmJWTPzb3zhMvoOOLn3GAEAYMXC91vUXf8YD
g+32sJ4NpRpDZHtIdLvEGO3fuADaUhVPvAk/DXrA8eDOwW53GL2l1nh0dmwoLkNs
D9vMSGYh4AnJ1ampPVrntd+lAB0211CHacPdobeS6i7/+3pbRjtbSC5SbY0V1NMJ
qUNBVO1vigM5cyuChaGaSwiTc9ZRf80H+gKUSkW4Y1H1t+oVgwLOuEhVxSURAMEM
6DfvfsoKs/Ebnp8iWkRE+x23LWY/U1ejCYuofN+XfOlwV2hz8CiO91tFh9nKZhrC
jmXZbG7iqV4NKFjIr6/bOtgc5POkXeSkX+s7nzrI8E/+3OiWv0ktZ3b2Oc/BWjLQ
J6i+2kOMDC9PHDTTgsZMXaIo85OGvk92aKdgTO3xPjVYUVDSczkagm/BNBnk/qzg
mYyOS1EpJBZdQPF67iaQCYwgDv7iDqn66eAZs5YQ0VoX8uXUJH3TldbHGimKA5Ca
kLDNblTUS6ShzLuJdCgaojCF60Rkd329m0Y9u4nZw2MxxtnYTC2KcyRrKhPy6X6O
WHEpmFtEeojQVkXQbCyUg72gIZcJDMiVszXLlpG45YU0EtvkeIujM+ZisO/tpsJA
/xF6jvgTHsb/tRZiU82YcOgrgcfrJDPHas7BSSRgwNhY3OAxRtX8WZwVhV8a3hxv
vxf16bILMiJD/buFhbUhhzxI93aI771w6G1SZRITCOgP+LiZVkQd55VP603oB/nR
9X7VB8KfCOtBHp27eiiLesqn2LUQPhcDz+nvbh0GXVuQFZgqukNARGVx2KoPAWeh
ViG4UIOuZHmOrOA3D+TYGSpIauC7TR3L2W8aWwfdmPicDYjf8eOA2Lj+Xo9Q21bu
2F23BAcguOyFOv1ACUR90FfqPUU3AL6d1/EO0sAoDiPgYCnoTP7R1U+2e8T5tTsX
oyV+WOYwCFPjO+vwkLiteTatmI74mTcWjpeWCTI4cJILTpcLJ5Yky0h4FXJ8TH+o
0QUeFKzZ+jRzi1bbMFe7laWJaP18kWXJvWcgtCUfYqUSD0GqGaroz07ssF4B3F9e
naIDqv2+mi5RpLgQt68IbqGjg8lHtv1z502+E0vrvKAF8UCRzN+/q3rc9ksowajU
DvL6j1d4h3qVcPDWdZxiiSephKAW+yJ+3zKTuD41E15FHrqMAJqSfFTMNDMsqdB9
6em/gQrxh+1oYdxIBwdPEvuGfhnb10VeW/d41TUIniJi4Ij9qeh+SPg3fXAQwJ7/
M75d1SpcQVdiOeZLOfscYmuC77jkGiPF1fS+hdYfuM5pLeHIKSIoBXVS3YdiLcMA
7LDs3/Jl8jpyoUVKZGKg6m1kXkd1qQBH+v9+MbQfjy8vc8lvp+fUVkQKSLy+ZpnX
5Tin0456lanAudhiAgLvQYqIlpkwXLL3IbEqikBVeNclfVCORzFkZS0dsxMS3NPw
pVsK5yWUMfd8UCXKKqX3LpyJxaWDnJH1cz1/fPfzFLCvWn5F1kALYeWrikuRGxjt
Bln5jtyzLejM+xPx95qxhMJ4PPv9QQTDyFZfyT4Ggn/sdadGhZWokW+wpUXBF+yo
F0tQU0HXhtlY+K4E0NA5QLVZIf5hIAu5tMtzlLEpuGGApvB+gNYRxgKSCECXXDZN
lZnEo7nX8PWejknx8LPN4S6PEsgwcmpGt4kAipr88+mF5/J15lhD2Wj9Dq6YO9J2
oNpei2fm33w6UV3FDIaZPsN0RSCtJR1FURlZKy+JcaRTCOZS/AYySrjXG7TxtrbG
eTf4TQj+c629hnqfD0ICZlFIsvflmo1BOyP3C/7IbGzGPljmwkTTSVofkacwwGtv
jbXP9OYsVBfTKJ8FGRUA04s3rbU9CTvh0OSVczDh/YR6Iwk62me5tbEldpMRIX2l
D4y/yOGxdf8sC4WaiUiQqNyU1IosE6moE3fgUW7oOX+wESnQjlrmz/MErfuk+6yK
+Cwo7juT4W8ap0Ghk54gwFqYLpZpdth5Yk846fPsESw1RNUUFu0Zl7j/7xtEHPJi
2TLjHuIxsUTZz9WW5eVitDnRBxmAy3kWo+NyfkiaI6aOOH/5hrf/89f/DkpGncVO
+dV5z5h+BYT9I/3iQHUmqoF6K1ffhWoOmpbXUW+gGCIwLFh+Q6/DMBP8IeINqEKh
5oRNIKgU9sTalnSsJxdECxWPotxkpFX/DKJ+7J5qcJfGiJFtlp8QiNmqxslo/BRI
u+mC1YeWMDpzusdfbLMSsG+lE/yYM7rtc1wPj8cPgXbu3Y6eCbi3oFWa6cmlJQMT
bSmLffK7ObPDDQa39dDE+oq2Lt0wNEtAdlNN7ysNf8ZkwzEiuVdoHa41ivVMO8EQ
LkabVPsp5nF51vLGLiupXlh3xnlCwhn1BPaFVfSlflYgO8Zn8nnuIbryq4HCuSvJ
NKO9VG6j83VnJXPPZy/7qcL8vPgJRNH55i9nwfD2cAuFoSrR37u4YNw57gj/gikx
vvRBTUXZbBLqliq3yLKfPqzUAj/ab6SfPOH0tFh3RuWR65C5T5IuItWXNEDiroab
fYXOA9jV6C1GOhP8eOBqpq522GOGrWRuR0pLruBJd3sHPx1ajth8XRazkPe9jzzK
oF++e15GuK13GZYH185NwJ+xNfpfatXAdBAauJlJLnPl7Q3mLtYw6gGpY9zaXKZ5
TMuJtht8Whqu+s1BUJvd7lZM1ns7dn5axB73x12fcERPuUj4D8Gzwecg/i/HcLfq
6De00bFM5/2EFVP9Em2yr9Sbh0VUssdP9ytI9jm/3xHvPgovXbxqg3yvE4KH6+uO
AvSpMBtLSlgIRNRuOans/oNk3kTkHLBZuNNZ6mzmhpgPbI4VjBfN3AOk3RzMUZur
rUkGhznlEX3jPo2hnLifxXOtfefEpSKuiX+MMKymkTvBPrCB992Jqu/94rletqa7
Ko5iCay00ToBh9Kv363Pll1qEUFR0OZ9ti8CPCZGK41XXIepm2S32XET2zS2nL5G
r9rrb9LBFAisUlnMpHlKGJqSeIBAH4xjZy9lh5K3zibEQ03PUhJBcdVVfe3pUE13
8raWtz7k+Gb4A1ZMCp+Q8wNBI3JZxoU8cFaU9qL/O4Jv/mH8Yx2QMO7Qn1HiDDdd
3cW6rTT9OwTnwP+pLKgYWQ2cztrQOtr9MdymRJizXgGjn74L6tWuoHzUiGmK2V0k
S9HNZdmWdAxmzd1M2r3C8lroYzPgvAqiFeH2OmY4iwh2IjgaPFwaVr4zhIeaRGcv
zROOe6rCgrzQnrs/NzFN1ixBTQDaU4/jwZmjvPkJr4Sii6ncuybtKxu/0CkmJRFT
J+2StH/VcrM6VCAGZDrdwDO4MJXoXgFCzDhk19Gay1enghUPT4cE/5YQ7R+MN2hG
Z9GmHq8uOa85mrBAM7LkAoBAQDuBspXNDzTqoL4sbJqxwvyfsKVvrvTuBI913kzL
hY0Kf34FEpCNkCAn3vxPDmKhEXFYFYrD1O/QftaPQf7N8VK2FwZO6AULBROm3oLB
rlDxas+ENmPWkw+Ll5sHmkKTSjgp/7n0A896BqdSiKXmYCWQ9vVCETvr1RSfPvtf
OCF2Oflx1Fs+gMN3BJ9TwuTb+vBDQewsAo3TXapUybcV4OzHMkrg6ogejdoZBNRA
x5A2rM5lUfBMqZ6vEBnwBDgqHNwb68SWjGl6DNaiqhpUm6Ea2NcEswqBjz3WqUWA
mABaQw214FyTf9wvlvOlYWXEhHjGewC9lp3myIdLfppDVEN5IRxb7hIvfhriMvGg
vJajfCDJRUeqvwi5brdnLIqSvBAm2t+nUYbHGMLLGrOPbyEUSK7fcx1m/x3D9/qQ
vE51JzHEAfYSFEco8FpTZtFiOo8RWWJcaZ2E1qYQ3mRF/3BZMgQVvJrqKWWgf9SE
X1ICUWQtPGPoY8uBdyEN8AMVAIKr7gFIMg0Ys7YVgKbK2AiTdYkoTYhEXLmYLxpU
djOWDFxOiUBdypEqQTimcBqP1oPzTGPzK+NrXGGi4Jj5F90szClosNDfzer9JVzw
KwvXS5swn7ktzMD6SBC+9MEfxcMCpm4nrbC54gdWX7YTSPoMsc+4vcxXGYOUNCS9
d2psCBSuV+e4PymXRbBvQ6M3q/KBAPFyV4B8P0YubXtzpEoLlWKqsa2fYiNyQ8Gr
lzh6bKOZyzmzlZPdWsI2F7EtlfThOLXUSg1AOq/V1qvLbCY+9JzhxayNw06mBK/z
vUZZYVz/in8b6QP2RKU4XcT9xAqsZBpk3xVdvTYXLjGs3W2XmHbzumYFS5LOSpYu
7wN7WLWSsiWLYaTfue96Rx3E+aSf6VfLZgQTjVW2xJsTqO8wPscm6ItRB5hPgzl/
RKtc/1XFaET8KUJPJxjcfZv+UKQY57OjYfvpmgzWwe0vqM6M4EyK0ekmwzR75p3M
D/UIcTTwuQdjD+Lo+uM9AFBSrsRPPMTFeoqu1h116BQmb39IgrA1HjTtVJyf8fd3
fAl9u+HCcmVU/1JdkSQp7hhKue8iY3LoA0zjGckNaiDadZ2jIaaG5mewsWQD0mgU
WWmbLbcSKnq6rVBElFUK9+ju+8rbd8XZXu4JpMoqhw3Nys0pkcZIYaVTffk0t2Cb
t4OOU9TfyJElv9PVHeSYhO8naGPUB7SbOT+D322Qfffu6cmM56rfXlCnuKAnJydw
GwQNFTYtFMo8DqPB7nac1mgy58RYyJlzqmOgp5Bn/a3FIpva5L9wOwYO/uVMEaQZ
PVazeJRN08Dgq8YEehTnzrlNODIOSfUI6oLuspbzNxUCrcQs/lqd3wlZKGNcczeq
f2HI0Twj9s7DhnxjKTK9ULulDvApZwl9eHmqjPhUVB37usfqwoPAu4IL7v0B7eZu
BF6u3qKSet7w9c0pp8U5KMLd6mLn9WBFxgWxdoi91vnEkSdRGUqle+Teo1RTbqr4
sVixhAa5Mm+3fHt6ugufhcUhbPuHJlDnKTEMBTaih990X/WlDe4MHc7oXJonMuGe
QcQH3bT8GYGAMjl7PhIUk+hoLJ/NNBhnOAIOteF9sJnMBxD3Qqom4Umf1wIYqMoS
jEzGXZLg6CFry25YVBJE83Wi2ti3dqlKQGZubsDcrk8zEi2vc5kgSKqzuuA/Hma4
NmFxNVi43ZwuX9Qxknz9IoQ2kPmiMh2iXdmSmwhpYEiQEAbEJh+X2GLgdzWwQwmk
fXGpAI6kkRxcvEMv4+Vx2L8Dt6gJFhKA+tLv6Rts+puF/dOD/wOr9lmoYjc5g+2Z
26f70Z7VsXXBQJ5TxfeBJLEsxIJkcN8GZmG6HE88wfAEtj+M3qHHEyA0VMB8EmlG
W3Dy4nc5zd1ZpgcCti8hEQutTy+/SZdU39dYdmLrePkdqdy/G5OIkpdE2fzLDVTc
xicJCasQ/D7qLvHip2+pUb5cIBrJLy0a6U2Ccf6UkMKHPOmNDXCp1ZqaocqCh1Lc
GcYcwJOA8IjwWka5zXAflG3Py8i1hJejrwSNuKbfCahcfvCO2SU5gHvgHxBhXbVO
trX0EpQE2vK9UJephpln4vr8ei8BmRx410lY8ocVHV9FJbdSw1aGq1WhdT2mdHSy
Z0vWBMdBjUrVjicZwt2FlesGVvnn2ExQnNkllOeaFukJsz5CPDw3flufHq2em8eD
bEQbIkHbN0q2etILObUB3JR/e0e6bYwF7aLxQy7rSiFn4pKG1q0lzVAbSbzLuCn+
UtI59Ypz8Fc5G1rUenABbv04PFuk9QBz4P51Op40pG4J1uRw+AMgq3ql+2nrcUco
PQF7hu+8PLc0tpEfA9hASgB1dGHtwEakv51Hid+Bj/WMSOES6aNmWjCLhdu/8ZT7
JUsUItu/QgLfsfJSgQ4mdIyJagN0LO04iIURiPn/SzEk30/GRNTYLaKWf7ItuhJi
lMlFruIzjNneGlWjk95ECLwuDjqFJ5d3/vCDakmQUZuHCA+pmlMv2oCEDp6e1MFC
F55ubWGCmKLOb53juHCAUed87ATU9zHoc27OiGGUxZQM70T7LK3GbZQBmwRhgWgk
WNUCRHzbxY1MAQ1z1uW9gJJFtAYgqimEQPVlwS8DP8xzvRdGjJYv4qxFcOd13l52
vxijBwezHS+RMZsVLU175XqRXd5Tu8t9wOKmYZYM63UYTi0NGrnkYdncpLBbBJs3
5KNOt/9yPcQPrL7BNBANS7g9JQxbkNX8msZtnSq4II+aZZY8hLyJDJb0MJ81usrE
b8T67hFfiBaoTX9mDdIrgRCduRtBfecP05+jedH610Gt/quGe/Gz5OvR06sYZ2I8
9zMsGHAuZ9axPsLgRBNQ32veZHSngWY6qFe0lTOyZY+n4cTa9FtLdr/ojJ8q+DAk
05KO9yuNmeXSEIA+B7rpYYqKNDh0jn5tl2p8gP6jFhCesA1soVZ9rdbYqe6adIHS
UlPcGoxFnrerVgrMyJ+OjhbY37Pk95jBRFNLYZvoIalqD9c1HO6WlIJuGldi8SRI
A+c5sKn4v8S6tdFcwf3Cdme5T4Urapz1e9V4QOeBNxkQO5V+rYlQDhFTgafbUFsC
JgnkShFH8PqOas1J8Qdd3cM0aDtClWPEgid7dVH1ratimeIrka40UIfJucSvwBI1
a5t1zgn9zg4LSfOWz2aXiRBLF7e6ZUK8Qvha5vCQ3a6OBLX2V9EFmPpELgyci0YN
+4ajYNA+x/c73Wxjypz97z4rDbx5E75EIoorFttzVVKxowwLcAYtA8sKXMPDPTxI
iDOf77WyVMBfRqXlVUAhNNUAH1GRNGC8UTb999ry/sSaQ66PD5/7MPTPoVWCn3k7
klAnK245s6xP3Bz8N5dLlfYXXetMRvvwcg5V/Oc9Eh6jBdEfWIu/5MsPgM7+oxY2
DqkfCbPiHG3AscDFlNwiuLGsmWDnFVOLtw36zjWzKb+xFO0jIndM3vC8sx4YCOuE
c0QNEFeK/5ubs1k5V8vtOEn4cgDGiuf6XE0VcdR0MB+faEkW5m0HxS8parZQ5cd8
msF8MtFNEDaZf2SUMW6Fal0A0lk9WxB8Q2ux+WWHg1Bfg1sHEXbU3MXgoaAOnJCY
kdUjIF4aVcCs88veVybtOp4lt+2oIsw6CgdtXZzZJhfDIFuNAy33pgBmzrP+WeaG
oWBcIM/d3sw1261CGNh9dvsP2uqi/6piwVp4buF5PyiF2iCcFGdGOWeMI446l/Pp
WysUEKpaE+MYsH3EhYGqNUYLR1Oj12zR27fJAftDPW+yPRm35TJo9zR1uTVzAKnO
eN3w0g2NU1kPplHcScnzvJIHa+sdjBaeQuPT4gxGyQ9Ajkwnq0w8l3E4I6O/v8xt
JK9fRlXGrc02a/owZTcvrjDNnbcsKsGt6pogL2q+9vDCzVzBgiIqpiF1cKpKzU8K
JjEr6qo8x2vCT3i410sQlMhBzIoo/I6c/e5ZIuMWfEM/CJOcm50NpSpQrMO9IM05
vIg01EMhev1d/Z0GMwXFFD9MD5OmLKJkTL87dDuuaY1Ic8XWJYbLwQFxL0ETGWc6
ThwSDOyHOLYkOIK6JBpcvnFoIUq3p8TfP+fi7AUhUe+a/ugp3s41O9d8nrNqhr0M
Kp1gXxk1dmsyyUwCbVqLkRv8eQBauNoZ+qF+itesZzB0C4vZ6pjXmVSgkL/HmDwD
y4LaLwrC/lduDPVu+a+XLn0ALpb+EMpagysKJbLdalFVh1bXkTLR8+PPRXLUVibA
22KymizsmOBysrBMd/MS21aUGXKblCr8iEeH3kyXwyedV08yORI8BN23VeqymKx7
AfSOaaH2v8b9Rlz5tG4wY/yUNMlmP+J6oFyh4q+ChX8qBolngg+1FFlcIUztKJfF
OL/yW8IsyrBd1/4l4NtraRYO9bpg0C9usHcUtV6kymegLDzYfYnxjoiGP8M7hF6K
JjbMbQT+o2M+R2JMdIv9bhb1haQv0qAC8YUlQeypMskln2kq7/8tcbBxjYkvxyKn
Yax31qqXuUi5Q/Nk2Pg3J1fl8X5IlqpHUaYU5rS4Qve6Yp/UZkViYZMU+y/3LBR6
aDUX9J1mhsf+mMi1i9xRRTSxd99x+Lwnaf0cpbZGIlEBeU1go4Beah9gqV1AXtl0
Y1lcCx0PEJfmIe6UmOTGHg7HRSgstflFJ9tivoPQaBwsfG4dgBWQAvb91Y/iEtDn
k9pXIG3ngC/3UcD+GYT0CIc075/L5jMwbtBFRTJxNKg3VD5AX9hIe/S0iq7nV+vl
UnSTvjKkB2c8MgUlMsKyVXaWes8bR5luu7huKulbJhktuDlV9zxwvG8mrBiecKzt
ZbKPXLnv/vDnT2pYqGsN7xAdK5AyYWKXiRJx4J3aJWmGj0VzpMDB4m5qDK7QFDOx
t0mAA8oNy5w9NCBcQpTjtmXLOan71AOWwkx0VcVSbABfLPgXE9Y40sSIpgGs3DL6
IcNAC+LI2yG0RkkKkCkkLkk5fjRzmmHDhQykqOyPAsqvQAfesqYFTrNx/TQFJqjW
yePmzGruDzpa0Lcs/b0tCY43AqmOfXg78TDR8VkP4rUn7uzzg5CTHdKbXzCRlyuK
RiaFEnMjQq35DC6eSa8bqk0tkBM3Xw1QHwv2azC1cmAA1TOoHlIACdYUAvnHUQNY
lufQZxiFPQy7/rrLfQGdmR4uPWFg6QXp8atMA1WJID5hoCmL+kTmsYzOUaDFn6bM
PsEQ0pJvrI+bcrx2ij/VLLAotEfkhGiHaZLSzSmupKq6anQpGLvZYc8ryW3DcwhA
ZaE8nGiDJAcQhRkIIioaJVRR/URakgGJ1Ieselu+UWzPqYud3s/79WLSyBn8nygx
U7xyGZDjn7eHph47ViPleDh6VFdiUwSZGBf1ZxVqTf+o2bZuR+4gFPeMHm5FSH3j
9xl/wsLydiRQN7YJDHjm0CoB5ZX3Wicn67L0leX9crEnDDQLZjTh4DH+cOaTZ/nD
q3nBqRvlwrZwzfsNaFruteKsx/IsBcA6YWa/z/A1GZOzZJKySEVddckG2gWtQtlj
xGzwKF7lu9L3zMWygCQhdne+E56FKIYzEIlOJ4PZxo1xx0p3gjgMJPSnyM4VyHHG
od5AlJ17RavGJaU6imFFQ3MSZVLb42A/UFIrt5cncCuEHU9Hf08GIDhb89PcNv8G
3e6les4J0Hy8s7GYTaY/bK+LcjgnsCNXv1RofRP0Uxpseizu6iD34Pdn7quKKMPb
YF4OqRKNb4xeh5aY9gqBwK2ltG5K4SqAFbw9LB6+XUFNdqxbTFKg4SrKYhDlFmH2
oaOuUhFNWMYea5j2cFWUey/wTNejFRBGe1QU/XbjcuLhklrU3l7tX8GMHo0rrcr6
SIAUwUaKkUPg80aPhNwysAiJWdsAdRvd8uKqxwf/aNTLk2v0+OKpWdDYKykkJ49Y
Fz9WuxFMHjhZaL6LxwN3HwYfzfAC4NooB6GcyhSCtU7oPwZ0ej3h4MSQQdR6ZDpY
+mYaFLib3y63EAaJP4hK8Syxwkc+InC5R8epgeHZSLZcS8zrz3ocv1Fg3VGRUsbt
iwtodDEL5YJounrI+f2BjGJxRKn5okQsTzuTIvREUfumH+dRSIZTJPKyASYX2wIs
onVU8beE+V5IVLdPLF70ZdJdxQuruSZoOvN6GzeIHGeDENGrwwwML/yToSjE8QEQ
4x16JYbYQBnPryQSqSqOtv3tYAsb8xtKMvan5x0jNwfkJdz62HyLICRaw/SjsAvd
VOx+iAzeeLQXLzsRlFujkxQZP4xaW7IOirCr0gaEEOr/Qw31S03zqd9+CTTqC2xI
O5uIn7AKBJAYM4DV3ycSIPzuSWVMyXRbT6eqr5lLtvUJUPTYr9qJ5T8FODjLfPFF
MGwHGfJ9+YUJOr5sN8bZO0X4Yo1gBfFqOiDwN9OcCtBpzw1ZzMeA6zN1DKZLIGUa
5CjK2B1HSg2U0BhKHpGc1ptnYhZRkYVyDjH1OMOdvC41+nksMLWfqLC0ABguR9pf
OqvDAo/1EVHgvF8vLpfs2ph7zqtR8uWDSi4/EYkpoFD2tnNkQxfnfOVln062ij7W
djsmgGt8d6fliM7vu93txy7Qa3Yzs69VieyJyJEadwc4XtoGuImo4esPoXgERlpZ
aK/r8ipUuDdwsf9FrjfbOviAL7K/77sFpqim0CKaiwT4udZOHnadcvFxFZ+bmN7U
fN0BUgKQHHgpspRdOPDPIVse0S4ERz8ps4rjRVtuIWJafGSDQJXZfPvPmh8xXNCu
1yalRj7AukS8my/0Ez1PczxV4aQaFBGfovthZRSvY6f5HTN+fik8BQJxQ3hMAhPh
zKJ1miwO2Zj0OVEZoJa87Io1StnGCTybiQNO2QbxpIyxuqRvQp5zEOW2+0Tq4a0t
5zaluGvWrGKSCjMZxptE669WFSGEf1dMJnh/sB66kxbP+33Off1aj+5UbLPdtjXh
jmDo6Atz3GZzaXGo7VGJAQhLBLBTOls0/zyYKp6t+rWoGO5SCR6XMb8wTbm2dVHz
Y1m6b/DQVMka2NTL6VQAXjV8tPCyKaL9BBACsADvQ8IQ5y/oJv/cR1FrF3cXvQ+A
HINgrJVb7kNrsGgKiIOkng6XySM7hGS+F6J0kS2XEXEtQas0p8/76YmRMhS+gtMs
mKSI4hnfuqnRcseS+JfXjOztQoEtngKPEp1EMp3a740oqIGbu9J7WUEHua3x39fE
4OeVXe8SFOTB79QpW/bYb2jTFqNZKfTBP4MqDYt9UMkMqopHFCJ4/iP8PAlKq4fV
S8y1wUvFVIApmMfHZ+/aI/eCV+NPtmwrK959GKtrvFnM5PTSxAfp9SOy28D9OxSo
ubreziq1t9K2WZeKRPldv1pvkKgA9mwypwiS96fIKyKc0ASTtjwhVLLPsvStNZ8O
xRzAte8QyhFEhqX9XInP3dUi9PYV1f1naYNgoOGOTsgTsxITHOwm77o4Xw/uLu0V
9mvxrLpyFFC6nTA0psc7GWUK93a16ef7+s0SpW2v6DHXUt+I6I0sMOc5y/GjNVqY
Qc6TrHHt2cWizaCrrS9EbVYDFR0tPVKj9TGXHUTzVabpoYjhMVJ7/AgQtMneF/LF
1xUwZgMmPUZ2DitaNIXYQsnxIhLWGZ2PE0OJwv1He4n3h2rwhM5Qt2ok0oyY/BDO
dCGgfoJOzLtDGrSWvOQ/E8+7f/iYQvQvSvjWB99wzB+NNfVDydql592tdyXZgQeh
ZZJlmreMa4fVS2Pamy08Tne9kQplqs4WomB+qMWfNzyO0YikDtXRf5v2uvLuT+CK
CKR2hoIv5mM5sDWopba3N4ouDx/ZVQ9L6/+UMf84rNRg53joQrlbwIvP1FLUWrgK
Rpx4Lc+0NtMcif7IkuU9DjMkMrEYYuXLTBGDA7KE4tWnP7+UCO1/ULZM/+t2js6d
3++Gfmzw42cS79O/EM16VXZEqfq/E6yog6KiGH8/iRem+axPbF/aE7sly22xfXc9
/qeLRfpDRujXdxQWqSA/Q+SW1ffq+rnlC4y3fWnP9rTqGIWaFlARZxADDWG2ZCfr
aOsKlWp2ggjqlFn8XCctCX8MI2mRs5XN/JiISz/ZhbJGslp5r8mX0UWa1caE0JTL
o+5SsD5BUQkvT46MNibAIXMmDTibWZbGmW7GwI/2asFNpJtGmIQ+dF4t4BrPUzaN
uV/lcOrNAy2kzpiVfz0t2mMJb6gRVqjjU5hiFDE4b/YpnXTS/pdngcQcTktnDHoD
oh48uNG/tm1rFbagwIfJ5jg9VYk+dELcizCP29W2393dwG9YAUEC+VNQs0vmIy+F
xZPPuJroMPbm9dqSZvYweG113ydmk61KFwSuVvADlycIoB4B8iFmWFAjA7IU9q9Q
PlaPykS4MjubLC2PVuXUv6KA/8M7qGV/nDGWUZpzswUYc72KBeAaS+zqvg3V3hcb
Djf62JeeprcEEl7G4u6JqZnE9SvJsYYtRYRXPeVAeNT6tyqyOLUAkpWEGPP0kKHw
SUJwgNfNjQzKy6wkxLdlh3FhE7yiPME+0CVHPIl2Nc1wADBlxUQSVU2zflBSwsCR
SuM5l10+pDrCWIbkJmD32EsztldH4M1cTwluPal8iJMKOXBnbQcx2LDLlVLFRchR
yeaXNP1FfkNPs4c5FI77MZ9BMu7nM8Pb4VyYoxI5rHJxcYHrnjGJY9EWzQROg/hY
tRxmhH0p/dY7fnGOxjrrQG8yQwZI2jwCcR6XgXxhbID0QIxyub8DtcLUlpNvogv1
VLtQiAotHHUL2B3SIMH2BOUcTsu/PTi6OA91mcswesJdC8pBAbA2FiHRTu/HC3M0
I3utW13wx3TMCjF4132mu2FeFASGTuQcnCzaIwitdb7qesRhFxIjRIA1YtNgQfbK
vGKdVwEu33Sy/rCNLghvUT7+KvXsL9aEGBf5mKVMywG5pMU08nmqVQr8nJmX192K
JPLyeaq2Im/TZ6ianbMuIqj8r9zHNCp7y2cU048l/f7vmhA12IL0MMQ3cwk9avpV
3x78xGFcnxlncEnGZPjEFKQBXG3TDnu84rLkhLWXTHuLIyyWOEhRqTpbc4UlSiLE
6jp1glRsgTB/k3QuzUXsJnjvNqdTPpKUZltpXJ6wL1f8qYQtb8P50cnHBvKULfnE
ZM/Z/wBMBwJA4WpR4VhIIobMs2vZanOumSB2crhYX/N1WhUJDnrDU8H+sGC64vFq
Dx+DlchDSEfmqeTO7t/s+rSQ9i1GmfILbCh/pb3YnR5dgGQaWQhmVgWQVL//y4Ww
D2Z0W4Kw1YozVSZ27KLj9Uu62oFF9KhXCyxI6SOZ/9cNtfGIDcwedPD9XAfaAgEu
HWjF+xyfSmpVNpDLMcDphnUn5LdxULP9vGxMkYJYJE00T8TQBNLAbl98iI+vrVL9
4k1LqTz/0XCS8HarsjqH23cn6uts8np1JTZ8dP/RMu5gKSP1LYnNeL3gH4nKkx8J
uQzNdLvlB3paM3DSy+H4KvvOCuXnBfrx8ZDa3hmPxU1syBGrKJgvZb1jlSRnV4Dd
QeYWkdmb8qmMdgfseFyNmtpE5MgkXURwO/Ecbxc3Mnx6C5SsFd4ca91wmQOFUn8D
bf99pT2px7uxPaaWdrPqu8oJbHiTEfdO1i6MON+MBEN/UerKNrBBIPKlaTG6mjxe
LWcP61/I3reCIdZeiMji04v4Z7Va1FJFYClnSJIPwDhDhdyxPmSp7BXVym85ra0x
KSHCawjbBhSIY55WV4wC3RHo5oTNd6vg0eggnPcWBSC9rYRMXd0GscyO/+4hC8In
IYEBAD+GewAnV1wTKIMPdW2Vw3BNN8FTKLrEiCuYt1MI/UI6YzlBZsk7y3ydo/nx
xoEkCuv4siHIf37y+Tb2xLsfsptHYlm+tIPfxVC5BKno5CvIVgicmbjv7riDjqZr
5ZE8hwoWXCklR24i3q1Bhbts/IZz2GN3alssHWZEU7SX7h0GAABnRhTQ4KBrIKvw
/O5ZRyi7dhxYsMIPLg92MBJf8i7HVDiiFlcKYNoZkqne8GA+7PRlNcvnfAZB2VKa
QccAHnng/OiJY2RxyKcIzZP/cI+7f0U9VW66jA85VE98paQKJrq9GXycKUJ9ogVI
hoaQ9DVgHomxQ3v+rle3aVmeUcNw2mC2GBP6Eo75mUJ8O+W/AvlN1KeVrq8+dHwW
nmgcB72vHhjI36oGXVYJpUDLon4NQEdJor983Qh++wSSKpyGpl5R/MSN9P/YboOL
nlOZolqOfOmAPSSdLtEiUSu5vau/8RSlGkuEVxbM1QzDOSD0CdPEcj34Xwd4SDrk
iz9w+nr8uqKCSIG5y4/AMPdIk8mT+qpeHknnfOh6Vdd4nqYsqYhwt7+GQ0qu89RF
E7i2GCYA0NdYUqd7J5RmlIp7M6lNi0Ha5FpSWaOOEgfly9FwKCQmTf73v8S3pwfj
qBCn1+DoOcuDFltJZ+j592iQ0yFEKQ9uXgIbCp1V+pwbFgWpZ6uYzDy5lNtKA5pD
Htb2Fz7wkHxIn4VGR4DSkzr5IweJlteZBGH5ta8V7flpLd/aOeE7u1zkVhI6o6Sh
MA63cN/pcKfLCYyl7gr07CYG+TWL2pXXz2nStLjAiDcBShqm7z0CNTRUg+4rYQWm
O0zMe8O1GoMhpYU6+2g9sSWDj+Yx1IsaSugIo/ok8FPmlvh9xfa5cK+Ujj/MdZZm
8kfF1PNrYvtx0dRJPuEMQq7fwjOprPvhQpUzkkwl057oUqQTmunl7vwip82cVX5o
4Kf5K5fMI1L28tdz61FECX1Bo2brUjhcD3/X4eEjk3Sw9HAJGCh3Bp1VCZbPuBa8
GPwSuHwZ0CdGF3G1L+i+31ASYAwYpYYFApzHGPKXMjSkYkDWiErYuQEWyt6XBkwG
IXEGHkuOLk1ZC6+VEOlMbJsB0xQ7QvBX6vBWB7l6ei/pvLK+W8powD2SZFNGZ6u4
isq4frbcKYFdJzmyguxUisohCX38/FMpWLwNtTI4HGqdajDV0kUjkTGLVumavGvm
I0tVzZ2blJ7aW47IviPFLlx3xnitzElGtgV1VG8ttBtpUbr1GD6cN/B/lJu2fznN
nNHzIPPfKhnKCFAF+9rEQpSBwA8u1cUmf5Ixo6Uk0mD9P4USwhcC8iy08LVZ6fGi
ChaKbZuxwGmrQyGwp78bQHakl7DAe1xphGdraBkF4tcpbgCNtCfkmrR6cqHBL0GU
CdCZMD2IpKtFOg8vMRnb/vZ+mIx4xAEyPGFodWBQNmQv3veSVAX7Qkr5PSTQQBjK
mOJ/aIqqk1r8Zuzek+i/TPojwvh/ZuMnj4ypf0PmRVAskSLSZJPrj+H/WUeKgVOg
7qc/DfDImIhcG/394k1K0L1q6wZlJuNFHbmOVJ2zq+a2WqsEweW/sra91B8tW1jc
lZBh6uKfbyjUIBJW1UtgKXvk8chqAvR4J9f8A603/2QUqLbk5dyXhiYnTQ6itAmr
su7egBfiAtlbEXUgF030NsQo6eQ1RuvLesFD3n2Dr1slg6U/e50r4vE5wKV4nWOP
1Hf4oYV2W2pb9vLf64bDtFpJbVmJkBecwfaKVzJaJOOF/ScDeze4JxpVdIbm8148
QZhrNuLFTiNRRIBafq1m8EKdgF56hiru50tc8uX+abNafgzGhknAfb8siwg+QnEg
EMX1clojYmie3czRCYzP2uhtHpNc9GjP/TuMoODtX/aKdWuKgQ0wptAme7c49vvN
EtHStzmBMDlaViu88OGPoqvVxCBb3coQLG8i/SPyIWmHF20MBYFS3s487eDpTtwC
IkOOr2Lv4qv0dwOuS+mWyVXNybm0SQa7YOP1hvbhGvUTwUMWVk4Ki+kDolrH66gI
GTpW0kU7V7erTezcKx10kDRQQ3Tq5MXuaY2cO6o8UguB5ckIzV85anQSApBxQZAn
BDfKR9KdWwY+HFBZEhzr45F3ta7594yDekOInpSDWC2e3R6pCs/lEDd+kvXamhwv
oqRR0pSLPvRRF92n8BifKBPwK/CLw5xe1BvGrEtYpv+ZuiCrwUvJc2GBzSoDfvor
9IudAb6yqeiPZPctoVkGquvBrU2n4X3OY9B6FE8oI+W9Vz9NGqlI1+xhTjDrqXTw
RqbxcdGn0/ER977wYGFej+00e9QgTPZkMWwG05PJol40E8Q/olLmbXZf6VeP/oGz
BsvEmspbJItsvdIVVD2ZFndR6FKszqrrkdHNtkx8eWWmxP8LrtlgLK7BUUtW/GIz
YSUNUQ3wPje4XhdIB6461zpVUdr3cjMedkfay32evZ23mmLnmVXlLVuhePwkcJw5
Fk/zERDkl/DpftjJOzg8+r+v+M6DdScktckjUhkILPqD7cUGskc+KTq3MLfgUBbE
7PWfeZ2IIerAUV18HQ0SJpZZVRqUq4jk0/zdPTMYGgBlDnZ1g0se0mdiMQe79ebb
J1qWkxTv3zGfrPddKbsL+VIbMk3V3D37Iq9+1uKfaDZLq4p9/Sk2Zht6DhxaAOkh
CuY5qF2SsOYQM3Z35XUoBSHwSnDa+YrMVGkQAmKODH3BCcoK74AHvifLFO+nCGtn
KWus8yY7taBQazD3i/t2OwdIInMbHKxMSfZsF4IFWS3yym+HQBuNtAtqgkSWp4Zf
AM1hMknmbPObqoULchCBER1BPaiGE4cYzZbijBVyhr3D8ZMj6D8vqUa1fj0neKqZ
pAcHuJs9Ut7z2A/zL2nNtMlsqKX1+qKzfnzoyaOHXTDAK0FnJzOgDg5WUsyimJpY
jLAVJeTUBaPnX/48RpgNglpm4NpfpYFxI4cD7sEmnvs0YODiVaf0s5JTYXf768OW
n0aoSgHxOjuPnu3/R2px0jTTUkjjGOKzYRoQiwyTYHg7VgWc7NVGzG21l2dq/AcW
9AR0AkeIK9VHPhec/BHLsY4Rwsjd4ry+RENzrSosVw1vkn4O2WCRIEp33YhuRdAK
mxhi9LU6oQ3Yk5gtM9gYkcw+OY0ubnbhR9/kvYsGDNjeqcGkhJZNk4USDchfowMm
sdVB2onSoQyWXR1aoRQA+WHf4drHjG91KieaUAgW/PiaUU3N2MEIT2a1Z1Vumuh3
GtGganzTdnqSb7KAi0cue4uLxLWSX1B3eYGBsIO/rQ1c2otsbgyXVObqMp25jt/9
m1TYCb9QRKK1JEE4CzNsH1bS6Qm+S3RIobs4Sgr1oPXP33l6D9nn2I/3snQpoRVM
6ONUby3t28c6/3WeR0Krj6ZiqohpZ2thQbsVeogXZAGm7mnrEw/tzajsCks2OsQt
FOsh5eNLYtTtdsO9EZbYGK8/imnl6ABsK+bxCRgGc3zm+iO6+lF89ZgtF05efxQ/
HmHIULR/stNpYNRsGB0W3ONxxLQoH8eX885Max9HC2+aBQv+prayyXL94EOVHdrC
TLPvh5AjPLNYXTkq6Gv/gJZcXrGatDdVgOifHomhbWcGjMG7FTaaXYTx7GSX2h2d
Bz3HXxYhZWxML0wy66E2vKWosTAlL8tgs0w1jeUSBpxVKqg1H8mO1/d1z2WkJ1MQ
LNo2mGybQkDGte2WebgAhuFxXuqs2B2fbbtSnExiEJgxTkL7VT5Cw1F2U/UiFz4E
1FGTIhqC5YJ6Bv+2s+K52a31aRTFGIh4A3TPLiViZoC1v1PGb+MaYDzYCXEFoREE
ndgMf4laaG+61ce4eEUhioVjaVo7nbk1NekgTxEznenkC/eNYRcJ9lrrIaqZJSSP
qU7WMhtA8zTd0z7dml4OQcEqd3LSlhrsQKJKs3tQWe9vx74T2UTcGvOuSv/KmGo9
c6FbEekVSH9SZRWvIK1Ugyo8E4Pf73++Aj/TuSYC0urpahfYy50ppuyL8U2GUaXT
E0mHoMcspaF7MvpMsRXBwaWOX68mQhaZbLi2ouqvajJxOBxAvj0PM4dPotsF/pOO
TzxkSGFkR6t0MRUJBH5vFEYo+q6h44OpNJTTu7e103h3LDYcdVDFr/1nXb8Vv3oD
aE6M8WYwkO2i76VBvO9BGVqmyYmmhSoSwEnSyg8zeSqTIf9SW5RMoBlsK/hAPGzr
izC/ci4Y8IUtcbW2F6gG33w0PuMn8HH+SbzugSwrobrIoWm3KNbxXytfg+SqpKR4
gHuxMxHQy1sdAHMcHKa/IbDKy9BwDuyf89+XEhkm91rC3gSfpe5n4SpBQhrnZUUh
JZ3Ckp8ThDJnwvnFNy7XRgyu1RRpdvjkx7txBWwzuOknvQ5dphw9FBSY0be0m5Er
0JMVaBTztmbAkAsUC4NpsOb2loZl2yCachaTRFIMSAbGEWIzuvUJ37sp+mt5JR6U
TTj/LAHfW/WVQTamJhYE/ccT6MtvSYIDbHKCmAWyiwBuAeZhRWSGxhAU0q0TADR9
SjE8InaxXJY42UiewpUzUgHNi1MO8EwVjWjdafr/7IYvQ4AkeNpdbnBC+9GybOxX
9NYu5lfXKY+G6QzsQ5Prd2s2ie1ckaLSyH9hyavaoYYydPWgeNXLHOBnzOJwtZJ+
ZCJ1zAqUKb6jD/hZqjzRBK3pqB2A37fdS2C1WC52X8pw/xOZRw9LEM1AEthPC/0y
AbCx84vbOgJbfWPpj/8thU/UAdR+Z8Iu1ex1X8erhEkCtBoCdLj+zD63pEjNgMjc
CKJv/jNnhcVP/xSIBmZutJm9Auc6XAhXeEdvMQRKdl70Ix/pV3zBr6/NVYikqKd2
1Y5NKHbVWRvtB/lMCePLfQlTUaN/Ra1UGWspHG19GUnEw+3RaCXvvzHp1+QBb/0g
58M/gPzpCh3uBObShk7Sr12FPqMvcGftA5j/gHqTlkQWLnT+ruq7jan7iZJll3NW
Z8xMjuyv5KF04nQz/FuLabLffxU0thGAKN6jXNSTElbQOuOM8Sk46rKF+BIihoNf
9336WNa5elWPgUnNkwEpFF8fWKmRepa4h7vqrVFPv7PRQv1qVR+dHd1itw2/olVB
payesvdycTKIv6Kc03rCksoTJWgrjzD3+31JICRZooNM5GdEjuo+/sdj24SYxRqu
2Sl8VkHbrKKmszy2Bjw9SXzVF/eRtKXw/KoodSXQWVXb91kix2qzqAhCVYP1ufsC
OZYEXxacar6dogeDYaGDgCInMrE9UvPpk2EpvFIKlMfrn5q+xamj0SvCCcC1j4jS
BKPvRs3PQT2N4B5Oki3uCBRSvkdDWfgzGfTJrT7CHjTiLhQbj1goELcG6pDFAbi+
Ua3YeHuxJGHVq2x4mdMeTtddlWwO4pRs/aJ2dPWTEKsMpNLSFErVa9fgEF/nsmos
Y/Obgn9YDQ7yD0Xi+Pvcp09Au2G8ExOiUk1aatE4j9r23a6hIyJgb1sQ3QspTKO3
Jvuvhbql32eX+wazcYbtcPuA9VGQTL4yb81vya6iuJj2SUgETE51d81B8It97cI3
IJlkC1goYjtnM5L722InXyJqLyIdS+G1falDky6mMnYH0IfXWnq3ZMlCFyinjN2/
YkU3iAW4Jdsm/A6UIt65GDcxN2gs+Ah1kV4ythgcUKDofwNyIfZzJC1fAZCGPq7c
lbTvBbmYamAzvYvmKSrhRYwgfoF9HnkUOUXGjIcaKEVcZJuV5T3RkKq6TCKxuSxD
KiJXKpV8NYCGEBrV8EtijDLnKKDDbRevShcwRYWdBK6ZVuoOx5a95TqAZuzDmy8W
dXKcNfz06oDqyFNZnE44LQQUdCkhIT7XnBg/iqVKesNxaT5Jq8xBg/7t0VABBVJR
EehXZHbLdE3OSREopHkt8ZJDKZdBMDcnx15TN7j1fKvjnZ7P9q0L6ozCoQ1MdXwV
qovsVnQkZe1G5OdPP4l5IiyFg78zki1bKXCX0mBevAQRgcBhiTHz8opM3lDqGUiR
PkDvuomcFToW6iGB9aICDPQuluBVNDbykA3Q2Dd4CcmvsjWs0+ByYy9gnV4plKI7
SfC5H4b7qzrjiW45dZsb7IxGIqs0htxjSSHJJ012+WZAsqYhFEoaGw0HInbfMKHc
q9L2NkCKIKOUx1LJT2sO7ZOlRgII6h5kNOsd9u5cqixIRWq7cF+Z4HOSInul2Da0
yeADfZnHzupP9wdtD/8V47F3Sw7KrdD9LMXD9b3KMNRFO+ENm02rlWp/r49rhpDm
dCkV8OzA81BhLCZQFc7PnO0xnUeeJ7ptrqtp0Irew5Fz8n/nFtTmatpQw01AVMtt
x6ILbkjliZdhP3W8oHBTrESfSp4nJpgNgK0Q/FxD95g4VgnJqV8vQ4FsGOf2z6yg
WuAORsSqWnl7bQ+OrhiR/8X+Mmqzdc3GCHpTcjttnsxmZMxi4Uwyk2HcF+5NKKo3
1hJPz3dusoCT+UU4H1PABBai9SRZhQ84jntUfH0TIfmHjpum/mUxGvQ3grt7gWKd
ty70zyuzi2FPzauaWRtmibOe+d81eN8GqKfWPoQwE347jtPP5plc2FTG5GXcIxmi
84l8pfamxQCO+GmIBL12mu6Skc68qb4vlWCO8mZbs6r5PBltneVnSIXRqCxQ/3Ay
tpfs0GlFqhNzSbQrtUXrbXzP01XMH2lBPqVwXEz9HEI7ZD9LoF3T/Mwols8KRNl+
o6eVQ1uwQLN6grSHndzKglH1l5KK4U38k5qvg4t3fZTjIuGXwhX4xIPUNvNf7nCm
Z3TnmYwufCRc8WHZJ7otsDCWoW+fhxZbTeBlw9JO1PYyXlXwwMgQtkeHgVtbc9Ri
2O3w+xShVvqvpyXGBrVpxKp/cdrTQfiDyv7FGbgNryGsKOWmZc1D6BH8p3VTk7y0
cr31XajxOw/CWL9P1EjkZPTNp2odOambuJxH9zIF7buIaW/gqiDbkEyeDcoex6TJ
04tC8HTyYP1JLBXQBQvL+JJs63l/5NisHG/GxVWECo+7LmNZIPT43RGAtwafR1Eb
b0awIb1gvX6v5nI6tFG+rGVIi3P88DryMd06SW7aw4Q0p/nlv3SyXGEtmNXGDWHr
BHc0BHgpvDb7upoYZ9PDSsmRpk2sFzwJwwsDEzMbzOT8Kur1H99vDdfPGCqf7hVS
q0x9/+cM+ngsZeHaXfqUbznSe3EZT2FSU5JnmMTrr0yXGEuG5fWRye/mT1ITzM9u
mFmfHVz3psvRyGQEtGHbdBmn2PlW7bueSfF70hQHTGB23HmaaQWhUDvojosi8QbU
dFlt9kTENMCfOF+esZ5F2BiDX3gDlPYQsUol6ZbRRJ8wLbXJIi18C+Vt/BJEXZW/
+WlN3lCxupnYKUe/nPh2pSaOvCyvKLRZCAJbMFczqKHct5cBqHEpuSXLyZ9c+mKf
AshDOg7kMZIWzSuxjk66sZ8GAtIIOoR4+BWbWm8+fohaVMuqYgBW9kW/iM2T6Kp2
pEbXTELfDwUiC4ZBSQfP7/YCv9sR8bUf6wAcPkKCi7TQXou41neF5IWwF7wWGWAj
ET5ILXgwtmHWkHhWK3vyfNDugYRTJFmpq26/BLztqI5/0MxoPUdsRqRQ0X1JQEuU
SogYzPGBtT4UhhEQ3TfmABxmsFaoweecn+ErbAfrxhnNsXWPdb3ICmSHsDkiMHHx
A9nnXqUdMztiHT3BlieQL7tvJr3+R7ltC0zxpchLjqYXA1vsAjBSXDkuMHOFD492
KFtYm4hj4irI3l9b2zvMI566DXYuK+M9ALtEahnQqXSHkP+qTE4z/ONVCtej/eSY
vyTE9kdnVXYB/f2JpecoyQ08ybwErYAkbY80d9VrDWVUk6jpcnYsr5jc1qsIolsT
x0hSJpin006uNMp8vditIIWimTqh+nqERc2zAw2WA3BcFolQf8kiskq4rzhgmMJT
47JE2ewU4CmedW+N4Xx/VNX/DOO/cSUQRtejVPwHew8zVAI/CevayNWYy2Wx0Edv
vkpbx+QCo7KjgXQEGsKvFuhnW8pQjoIKaOppI9fC7ydlV90cpm3Mtf7D/vz8sM8L
+0bajI/I3V4XUq8Vc+1kMRA2T71e5MIVunxAOBF0BVNrcivCYyDXq6JYL88FEvkg
wDD1P4uVBqo4de5YE1nFShQ+dml6w+ZKwa+XbxfpstIqHmsyJ2PFVdkfFJKMeJ3E
xgNL4d8PLbVgTzGsZQXB2vMPlCSShUNZBgUzAkjKryGdd8dyvHw7mcPgbaw3mQO+
KIv21CwciPDcZNQW8YgVbW3nseQ1i3UbxnfVspzvg5UGvMi0CSEflCYgQs93+7gy
esAKrP/tLBAZEXJ6jF2lLzbt2ZtWYrnFTYzzhNC99slrwF9scPB66oPYonL+G52l
y18kAkHG1YZdCLgB0lRaBQXMxbGAdv6i//wiDlahOoPdBG8GdO2OXnhx0OOwH6b+
hHjUr6eLVJmIAfyF6W+2mEQi/7TCgtmyVeZCWMs2T4NgoAQflLiJ+myzc//sKqrV
1ilFB8vNOHw306vPM98ijRsb56c0JfqMzg9QhkBPk000FE4S9c83fckELT7JKB+O
3kXeuOKKqfJVOKZFc+yqrJsZAAgAXHw4ntIIOBuZWs/AGIxVeB1tOh3XJFUh8XYe
JXtP/a5y+dNSeddFuXsOAsyU2EMwenEhMsKEVv0+3HJakrIIg7NK/tpRF74vIESc
Cj73T+XQFcFtEonyOcZvXbyEUGrTU1EvmQ4c8uDQAihDuGRANQhe72/N+mQbuynO
s8IQuFbvhlusC5QiJF5dHatvaUPZDgHqwHZNq6qrO1iqVgTVVRSytX04gvwJPvoa
DmBicQLJ4QmgJSO6Ygc5r5tV7QqxkJmXDw9+LVzfUku2R5hhLt1iGOR7yQQo3n4o
1VaMJZN4QoSHABL5dQ8L57+tXtX8cqNagmfkougpv/ufGrgASgnJRhOjWc4xHBMq
QqAcabfv254SSuEJQLk2GAbVqj/guO+aW2aCGLVEsu1jPRIFEQgkw5jHyrbIAaeW
YIt4FncWWWSesS/peH7gc9sOV+4XGFDWc0oF0vbM1RfleoHiwUsmOWgsp/+s3cIk
xJYA2h9v7RsTnP/Ipec7AuMX1MbRRDu3aJ9hsjA/ZdvV9u/hmkLh6JcW1u23Akes
6jf8nMPjf3X4K5QNOwe8NmHZWFhB+Eir6NwmffqTWa5H960VLQPRtARIHISB0seT
N9ynXYNpnBqRbGgQy2z6H9HCGRWYiV/bQEAbTWBxFcaUNFKna2ZgdkUdH12Us+jR
xtEAC7DuCCJYrtAW/B1eOJRhnNyifR5irHyVNTTr6adHcXlgGF+WXKl2xXl3TmxR
c7sYyCuV680l3b8KylGYsMUqoux51+CrJUduyXIUHughbGfjfyj8FtLcNV1p/l7W
+CAkCD/Jab51aHCLymKgAucPY8AkR4cCiTmkNZ83RWfLwpLOzbEXDHWC5wUlS4WO
jQz7kHGitxVVJ672nstp04uAC2FiGR79Lsq83EJRpmEw0nLbUfaIBlUCkFKGxR8L
G/vBf08T57JAWEohWbYMUnQZyq5CUAsMfpOoDFG+S6JP9q1rAQA5zG6LnExHBTht
lnr6e0DEBrAiQvbwjaCyZwtOi0V+2Xxi3ITMyZIVeF6zHtXwRoigZrsqkEZO9PuU
fXq6dJ3PP+a2PexxPXtw2Yed/EC8rCGgsNZyS2vrqsDzytB68q1bC47/LXMTeVE9
jamjo4M1ydpQ8s23raK3Dfvuor7f9ZV0NCR6df/g0cBClTfbtJyScQIObl3ulihN
Bke6Gy3fDvg18o8CQbHrHVp2o1Hbxx0FfExWMCskqzOFR+w/d+So9/sRsba/guwA
CKpo5YtKDvRdGppz7GmegTGZS708yZqgVw/zqxNeYnHCgudnRm9UQwV11ujiU4Kj
bi9c7XjqpiMCSuW0JFiC05F/vDyxfB55+ySz8bL1//5wj/Wx1mMm6vD/GKTTFS3n
Ywg8XREgQiC2m2u96noyy2kiukKfveuBKA/+wA8hRTyV3zAeyZwXI9tvh80OC+2Q
oFW+dJIhsoi6wRfh6R/A/GFTiXFBwc4tzZEBdvQBxR9CZVlUGjYGgODuUrfL/fMD
QLZ12/CojOgD7DdKKF0HTLrvFf7VcXfP6eO1n5gd8q84K3EvfYGXcIuPS0p1s3Fw
oNgMawBrcdm4/+eP+5tL18OCNQ4e01dkYwuNz2oWAqpAjWfy4Jq5T1BoV+Qim3eT
5ZNIDfS61bBx1COJ+yH84Nb3/D9ODbOdiaNQJcfh4IAknp4DuiyfWEmXtTmeJBaU
0VuqrJ+3zYdQqKxPzdsZbJpuW3qMHFnBoS3ubrF4giJWbwSTTcN63ofMjUPjP3iS
gs6v3owvg/3OuUejNQHwX4EkEjYUtEF5jTvJ9inwcaWPVy4CHcbk3Ptz+M77GvjI
EoH/wSWvJqJZLXDmJhdfw4FUHebEvHj87aw2/aiOYi3KE73XEG6wyiryxvJkXqgV
HcxYkQbyCZez2ig4655tX2AZfwqldaKWAuKzv5GxPY85jWbCclkaIYSqi0+BIn7c
VIVz2Io8COYrYyHRcBEAQ4aX/VnNVtqwgQj+/snBPFhrlMn28kQqarmM4v/HMXNN
KLoZWQ6dPwnLVuRyqLi+dxx8Fu4jIU6aVRMo95IG3jgDTJPD5W64DlOa9cp/AF/+
Ls4oPWd5FlMnn1gnycyjNMhmcixN8TlLERcuAYsqAEO38SjT8U0Nq4GwfX90BsK5
/VjQ3atA/m3hK7swaZdezBstsMp4YN4VWD7+HwCzWhC5bw1fvmn6B1ymBNLhkWl4
2FCatMCYqpynSoA5N4WQ9jA+qT+RiGGaq6YKCVLifTEb6EHO7nYxHdTnsZ1tgtbx
HvMaR3GqNJZmDALTqobOYpV2ywLKiaosxw6zWHTxqggY8p7JUzMh+O32BNljrdrC
rGm1hXzB3utOggIsQZQPZSIjW+UtOyON8oCx3RfXxOC0q3IGkv4dUvFec+K+7LiT
R8ZIpzWwEPHeFBaHxDu7//NdTWhfOJIxJhCfSsoRTZn3LbfWgLkbh9v8z4In/Qpb
Wi5HloPpT6xWHV7icfuaw135zqTzAXshlC7A03kMqslbU7IaRLYoScEQ27PYKR+C
tOEvcJTKd48noXMr5skonih5iwozhGOxv9zNVosii1HRbMafV56aVWPSZXrz3XEd
faXDdbDYBXEQ7tSHOr51u/9SeTkWKwuMGpxv7ni7vytA/o0q5CEw6qXSwDxdB0kH
Css2UAAulDXonCrzm5kL1KoKLMyaJvbqLHgVgivkF4S1UYn0iUlls3+UmAd/hniZ
74w27+Qb2ppBOGrqikJ9PRAfgHcaXA30feWubA0bd+293pPlzJJ57TAuYo2Mujap
8rCfJqzZfAGZ+goWFcaDM4mjK5uAMiQFhdFgGq29ji9Kh2IC6UPpfBkZVA2xkAja
WgXrolfQg9KYKJSLqSDEDdCIdarxgIEyqDsdQHBRssgzKFEwJwkIzK+gB906pdFN
1MBmrB3EzmzmT49gAWlUJoADJswtgPWFs4IcD15FtkGh1yaCfDerZsiCuvaPxWY+
IICbqQEwoAMTzKcjk4yziyklq8+q+pQLNtoB+TqyuCk/d/BT0fYMUEOE4supCkfm
xWJayMwnA5IUefp1RO/1Dqy31BnDHykkoXfKYeuoHuM/ID/Y3ZyRGoKs8aim0w3P
3iyRIOmZ13VDIeDAHTX4BsfMNm0QW424GfVYKUnmfyd8UFbTYkKG6iP3E8Ew9KbZ
HwFIt1buBWajNbCXojhKQrU2eau8qx9xEGk9dBd7cjldF9V5ot6XFWwUmeMk5RRA
ETHpSqlFZfKMHviAqZzKRKRbYa6c6Jr3LqdnXq4AQ2W1cru85bMsjjPWIa81MIL3
pMO7YdyTPFcCZZLRoJqvKt7XZTCZq47jrNibWqwWOuC9kkvw15OCROzS+Xd2HE4a
gXby6JJEvW5evfKCroTjRovPG7X6oeE7O8rZud4MqtQPba7DbFuhrzSKwzdDe11D
oOSU1YB4TITWS1MRWd+m3YfPy9PeY5GgmHy1qsN+Sgk1Cf0ShMZNpaLoVs0wrgE0
5eoUcKtIKTa6/d9qXB/cZW1b8pLlAR/ZYuNfFidkpurXAfLgqZSFHieWmRq7kwEI
bvP8LlesgR6DzmTh/6yvEwv141Cmnzr8OljUIOImvBZL3dDEPHXGN8s/pl+fTkTv
p/mKjIylMdWk8J7qyvJ+2h0dYnn008mRJnstjKI/dNZ9spPxA81ksa98pHb282HE
0MLA7MZnNB3Ob73/HbiZpfEgHIxpB7B4qit9orpxqfZ6FcBZ9EhSS96MO0mgp3zT
uXLmW3vuPyMYyjSVvorIjsqBEwuYKc/Cx7vXJbpwOJRAg+DLiDFTIOXSoegKqVga
qzm1F9VENW/88tb0ucQzjRO0AVatHKv6W68xp1B84utKft/9f2HEaJLdYYYTCnq+
MQQ+KsGw+Q+FGZRqAJuvsn0lpzTK8DKSucCJVC+acXtg5/vMR3ZBpYLSxdbgP3Y/
dRqoREcq0cBs7Xh5VhHjDtUn+uOp8vq1uNKjwwDG8DH6QXP6Ge0DSbBQy+OxeI/K
qY4rq4BrMlj8IIcCwcc2eF5UpRr8TKmr2L3R6KTpXgW/aMYumyMbJMBsubSrOTF7
8ZvkPZIRmN2k0HEuyKHBoNorCzSDZe4MkqUx0R0FzmXiSl0lWjvJMzxijCVtfV84
BUnMl7ojCLIicbIB8qDBElzCU5ujD45ADdjua1yUtTtt1AvXQ63FjG0EZ6uGW+gf
5CXyOedxI+4kSkJaJkygDRdnjhk8MgREL88NJxMehy4PTxDywx0jhvYAENZyqUUO
vtMlaYF0h1TNEFqLup6yYYrqLqv1y+sQ19jmBHf6gYi3/0qkejsBl3VSgk7oNvvY
e54kaO8ioHIeA9GqWGgxMB9VQB4nXVS/LjPkPAn3E42yi7MTAHCz/OHr8/hX7S8/
19NC0tumtWps4dLbfG9RtzMCcIFDaDzguwTW1N6u97fmIEx3zkKJrjvQ72IukE7o
YMUOvJyAiOga6FLmckOLQhKd9yQD8u4Xrmgk7vbypdE8+SWy62g+37lOKhR/faa0
xTU9+brKTrQRhJuvWgIYnKngw+6fgcbQ4w+BEvo+bdzSC2DgDPmDCifc6GmeqxBg
4Z8amqjaAnstHczrkkL8yksQqedhxTMCFQPhk0TI7xadI3/f5Uxy6acppdMJqRkI
G/j/xQWi/IJXprZ6aDFX6rP0erS3C9f4O1WRBUXjekIP0jmT2Nsq4MuSk4Ug2eCw
4uHaePMvZF7Tiq70skj2tiowOqLTznk7fk2keICYReD64CfnrlXd8JwPE2slr4pt
HOdsSzINL629REGdbbcD3XI0DgLQD+kuGkK5zW294UyzhUijquZLVwC6QtSar6NB
hPpjKMf1ei7OY7YLJY8IgkitaN3KY2iSjF4lAZosYRyrChpCbh4e0NK9wDTt4NPM
CVEAzt4bTlSQXAcnhqqOZXrS9esFpJmpmz/uvbwepCtRYRLFhITOPaKN1SHZM+0u
GEMa7VQ4B7/HbRwmdcXRTPdrhI/NtmA2v0j5tmbsI9/JrLGe+067xA4cU3pe5I0N
PbeGToG2GDN9c7EolW9AO/po7RK8QWsn8R0Tk8jTXbdna0pFAqBTNFClbDs0H9p7
lgVOU7JjdVOY++D1NbO3T9loQvm60HPD5BJLHtUbwUYGAS+TnUsC7oPDG2h36VVe
N5GsWVDjBsSl+W5/YG+Y0V1k1csc3p1CU2yTNftXV4edqMpMz4YJ5+i+PMr+ilhR
E75l51wtbEwdlyijarHG4cJDvYAvSxSKkouM93ybTvzVf3neLlOExhoelbco8dUD
SiEGYuBjVdfW/PMTu0LF+u79t1yZkV5twtR3idShiE0k7Locq882h2Ea9OTla4W5
TPfbmc8vD13ZCBdjQsrxnfHlQXzaQ+8pLiFjBErJst6G10cFxYnMb1LzrRq9LW0/
QQhE+Z6jSgoRuJ2QTQkl9O2VWP14+sur3tCPSSylPSykGJC+9yafdyYRxG/mfTpS
e0VdbI/OjDFr+yh2mxFl7zXjaZBk7FcACkfelluWL43CMdtt04pcX9sMZiFclrk7
ogEe4SvaW74VK3NEMa8WGMjn1pY9skpsH/6v5o191ER/5qC+zdN7Ma5SWqUjF84A
/4EPQM7CqoH1uRlHGvCNwl83SKMXynAE+5QcZD2OREPTYsZYwEzYHWZSCnJxVLi/
aGtwt0KnzBxaVmxXi48L16p+Y6MnBozLvCVy5ZHTCYxCKzMcc/cmuA27cmwobXa7
yPUoHeDthhKzl1oj8B9vOGzJSgg8EwPK0NhmX5HaXAeOwAC66QZlg7h3t4/b9c2J
VjN6FAg/AxFNxnUhrm86nTKF3CWd5QiIqRKHEJNbT2X9Cd0xYYOqZ2ZhCZ5GrHWa
sH8UvJX+Eb0HJ8COGXcmNscveg5Zl8I+rqz8AhBFWDnFPOqqKL8BdyQrO06E4dZe
YHF8kLyvxaFuhFepYkZpX3G2QbV5nLFqAr4uCeawV28q2997NFCNsfl0V37kCu+X
9hT5QfaK+Pk2J22OcZUpFkertXi1Js9PcGxiO/tgXqMoxivHCBNk3etX66zBtGkS
4C1mRK19vhPNM3v2RvfmUJDW0ZOXN2NyPtkPGkN6SKPFEs/Nm8eUTuPOpu5ugUhi
DM0TLkDNuLXZS1t/tc8cOhRABQDg8I/EV9WoJry8LDIp4rqPb+Nl9i8+1MOE/ixE
BEeEqsjA3pJ9gORtHkpMS4OyneVyaWzBMOlqQOb/E+B45+ZNlO+C7eFm7RLakTKm
AGHKhpCKvtcGKbTmvF+dfIxLnyCRk+eB6/8+7no8soH1ObdOl1ZtlefANYcVl8bY
NEJflzDhk9nyn6PjyRZrTek0GfkwTWwKt2k0Mv7z3ApR1vYehHVpWNo50ZfFW3DX
rdls0AuoCd6eN5R6JPP9LqckPgnrt5E1mx94kDsn830bo7vVl2gz1y22jBHHEhxK
8hm+B+ZTfnpbCIeycmG9rMQ6D5GguamixAKjcbdwdG2ZLwBCkO44wVfZMQReCuIQ
mmgHSionncOyUegrDNwTpAurXDHWaIGZsT1WaZhIg8vnKdDm+1dMIsQnu95XL3m8
fX+OVAmTlA46wjHjFypIdlMe2viXbbwIU/vVz3I15HHoJb03RUoPgaEsQXoJu859
d5YUiSVFFIbjI6UxHsbh2TtuHxDI7ewj5KeeD7Q/BYhGdloYul3Mm0zcchM4OPz1
6xVTKPQvM3/HVfTFTcB5+EhOulkTYQwMmph7aueOyEnNadfKtX57ndCfbwGKELQH
r71iVmvpVNXYnLkIJNSzivyeGVZJh/7IFOkK5Ffoorx+YoKSAaDHejRIrH2ILpl0
XU4WMsCMhhZQDihRePVzjFWxO/pzNl1qP202EJg/Tw+P2AM91wXtigCTpZ2e0id4
PUWLHT3bUX5qf0DfmFKqyZcJVElIGDCkwOuxx9099ssMjm+AuoZPqOe/pcRR6op4
tk2kU/DKFO1LERIT/FoCID4gwaGo/dv2XLyMLSNplihXRq+k+Mez6Jaebgr5ND2e
WnLbYHDla88TnHa+LJ+oNNC2Rjs3dFukoiKP2gPKbng+wkA3FGHK/8vbKESGuypz
MLd9S0AIEyzIUDnE3zjFG2h8Q9pGuSs/DWkbNJRJDD+KgTrD8vLolbbj4LRO+4JK
+rgE7Uj/RkExuCez/AjMuoKkaewIsj0oWrOpLbxsUiEEmN03+qwl1TrUkFDx0XFP
Jdwl+3YdbidOUoFbzeRN6gkd0ud3HAaokLBHwObm0dH6rk3AaZHpNYf0jHX46gqy
9dqHJm5+pD4zV1BO1MUmTA+KlbX78WVyn6i+1xl6lEYLVPRoJxOD6MZTtcDbNq/C
DgjhevtrN6dkL0bQKsEUMDhQu2Ov5P/fFrvfFUVOvi4QNerRIa6pLqqREPfA6JUo
A347p+0nMdr1oTCL96g4NEh0lhWbi261U3ov6PpScfjNqd1l/VtFqUb/pO5Hex4M
dnZArm6tkEF8jPY1txnv69nDsGKhLRsnZiujIdKMHeaCrmMotoeSfa/KY1oSWTvZ
8VwZyjRgC3tO6qPWDyqtXfwD3teNxKPVQkCDlk5C5hExzBo49cLuxpXWms2Pc1Mk
NaitPROcwtmTtxhFXMhWj3FOFvFZdXLU44gy2DOs2eg40j9QeXvLy3e1apz4e3kE
563H6fOVDFV8lZRhaq/oPP3XboLwXkiWHecSDjVaa4CloPin+0Wk82jhv1/6WTmC
S12WTumAqWBRrkLFVk/zTgINbjjBaH7o6JQybUDZFWFH3/LFQWpvsl2dzaDeiWuu
RF/LM34OlERGed+pa7tIDFZGJE6HgRueaVPoqsAQVJUe3TsSFwSzBwQvddF4AgPs
xI1aOQmxTYfcbGOX8TbYlAa5Vec+kKQjBNNpvbqpdgq/b1bjsODY4hpNNrQZthFk
1HhRHAfcvdvJYLd3ftiwKiDpx4oCR40NhzmW7k7KdBGXxRQ25W+BIW9zgc66M0EN
kLbav+50qoa9iMEO/gqKpOv1EeJs1kaygOnQN3MzPV8gvYe7RyXyJdvWtw67Ihzo
BDmhuaBnhaogPbRe9qK3eSC7FLlC1HLhQ8m9JwpUVEyy5hv+VY6Uc+Sx3ZDR/0dD
RYNwgOW1AmLivrSxRvBC646DRxc3ZjyKKSZOgUwQL238l8zur+qiak8nJr91OCwq
z87ajBhK2acB8R7m1DdOxCPl1+uNBAGPO8SX9V+briMT34+N90Bla7KDz2lxuLII
CN5picPqOUC4rwDD4s3w3nIouIhhaZ6dT5r/xUg0C2VYJJZYTLKrV++Op/jD6AVB
dG9mMkePqOtd9nW7P/veyoe6fIZLdxGUx7U7DtbLPLOPA9UDsLUEfk9AKekxiJ0y
LJQwYihjfFRotPzHeZVquPErEsMHs0Awu9BA0XIyFUQ5Uf7b9iyxn0tLby+WAU3B
HOyuYXkm8DWQ8x0mP3bNJYX87DUEqReTZt1n9DmCeDwak3Ga+q+PfyF2rMKs9DXq
8GUXa2+hFWYqf/qWg2BummUhVtBlsO53rDfF3IA2wdf7VxktnRMGl3zliKWJZZPR
M/X1rRDsmUEy8K2F7HQce/EXnD+itMfw3/EftDXmYLwbJj2UbwGev+62JKhLWEOb
0HPN43oIcu1xoXoxjr3KYbaaVI02VZhfm4MgmDg+v8u4R+C86srJU9SvtM4ypQ+L
75qNxObgcIMzcz4SHZJpsUL0LMo/za67j/l0xpqh1rF05PyBRtmuHvVRPcFIXn7Z
rHqEH2TyWgIAgZykCm8M1T4ymWf0M5P4cx4xypN/OS0wrQVzvEqYmvw6m8zFOpEr
gFk4dQYCthx8FMptMrpjmD//LwmuFsiFndJYE6MkJOUeTflb5YpHDhjdl0CpXzvv
T21OaXkLJfbY13/Q+/Uz88fYxqaC6fdzNsdDKN3nZEwDhIYK8eRk77Yd1weLCUYX
D0p3kaGqyqLyRJuZHH5WitbeemSKzwcv9g5f4i4Frl+lOqrVflWlqfmDeAkdPwpz
IhQx82pT10qmY5IUW89drhuTOxr+E/HHvNxuWkfuvG3+Dg+V4XvupnqP2g1ZVhhH
Vxd08bXG32OVUgy8U4ustB9Fpc1EGiIaM3RxZEEOH0vpjgBPFgJUH4nY0BVQ77CD
KILvKC46ukvSA/kNHba9u8ha5TfQeq4vgQH0a5VGresOXwd+0uxSb9EDEpu4AuZB
cxU7zoWqSM5mmDkYi2qnmpDPJS3vSyZYmPyEa6U1L0z67nf20vzcIclXcB4KZ1+Z
+17OnU9wQXvzJpPGKWQfxtDglDAEn6kdinMMPa0SA4lELFa57k7y091Skbe7SYkT
NjP1M9k+/YqoIhCjher2h+SwvwpYedYp5dFEgKWSDogVuRbMTKfoYUvqN69xh5qW
rwW75zW/V1apoKIuv0EZvq0QKI10jQaIh+rU5MOTdfv5yyXJwR0b56BMgDc++L7A
C9j+WR2i2P6oMiahbkOjLUayMbSDyPsMl/16BTIfTNsl19Ek5U7mge1NZ3O5aUU7
2vfio6acNk+EgbKU9OI4zGLTeJp5N5itsKJsex48U7zDiwOk3F5c8Ds9WJDi7lt3
HXw33dHfvxTMhxfG18TP9xeE1aUN2AEkCYJFv8M8s1e4tFo82l6qVZhOdcizUszM
idOeIBNQZblsIJl757cten4rGWMc4iumWyWltXafcrqS3cHoH2ZUbAqKAYrKkxzB
2cr9Js0GHSDrNoUJx1ncbu7TLZbjD7ll+3U3zGSx5PXI/h1b6eaGyVFsJy5/r+rQ
JODgSp5n9Z50MZm07I8yoz3exu8IsyfNDBRLL7/kfGBN8IcKz6kRqOHExvcHYSVU
44XXK0WIIi6QtlRafyxD+/7At5WpGFdM7WmIz40WV5BCF0mzc+1mlwTt7Ugpjx0N
8qGrgtmQ1YG41iVEpzmV9auJj6JEwzcOCE31fIdezliaB4UKw+8Ou2lvgcPxi9iu
BYFzsi1KY2vHtEGMkGjC8GX8ERFskSi2KuN9ArNEUOxWSD0tMvxuriSBXQvyxuKL
Ya2vD8aIGOTng0gZDrTmzO4VV4jWHVFv+8lNheRxCMKUDEeEBcr7VDGX0bO9Vpny
5x4lmACHcURK7JHBHq5C8MF2yqGTlOEx7Vuqesi+JEpEPZMcr2AsXgrjtTjPUgcC
9F7M9mLTfN1LvvXbppUI/eG3srQouotaRxLLuDexLhkmHvZRD+l7CPkb5ax9M7c+
92gorvYmOJsTNyREcP/dOWBx67KC97O3TeLyz/IADcIOyFMip2ApbVYSkxzC7bzt
3QIycJpjDpBscTiYiwt/2nABEMSs2tIA31gE6F2GG4ZN7+VOQTrVjNANM3kIHqKz
E6NIXxJ/tWVOAQZMZUOny7Uk06UaHDF7fWizxROkhawUuJj5DMhy/mDg2WATUsD8
gCjL8TBDEYdWjt3Bcfyme6IzUtQFQBZi6zJBsCNm0uhi8yrloThM9SwwMlZDvhff
aU9O97x3kRdq4nYB6fvRQpp4y67m3chaVzN7+KV3hhdb8hROgRSyLzhQS2XChvFS
HcUXSiBEWOEki38lNUZz0n14hKI032yKPNslkZVXVH6u667NExuL9owHuHkMqNZD
9S+6H4xniY2pCbq803kv8nm9rD+0QnpHeekZPuDZymS+pH09Q1Py3V4YY95W2nIZ
7itVUHqNHda8UPrMhwu11fTy4yL/VLHY3RhcuDFEU7UcPED5dZuhtywCHtvr0MPv
TAAmmgv+QWM2LtV+8z661Npmy5iF+qdEMtpDRzMLoe+LSDJpy/njA1Y2D38PRMnC
M0n/cQbHaPT75nTp97liZQ1RSL/K39A0ot8OGPFr7P5Vf3uIGSZj/L4zQRa7YSSP
6J31vucURkZKmD2t52g4WZ2VLS3NQODvpwKx8C4hvp4rhEGHmIaxxkUFIjCS/6CQ
xbjZfcIfqHm+CAy5gN0XbYkZfcDdvbXwpXXRQPN1CPDPC8DVVaU9NXsD8T1HoYhs
T/UWC+a0bFfVklZtIVaSiZY66ZFYF9sKH60BO2Is9woZpZjemUZA3MD3EoZEDr46
Ey3h/6whyXmEckaQ029IpaqodfU5ieCrQadHQxBT87PFD6vTp+/1jv28obLEJGhh
yMoVQ0g0WWQ+VHIPC0gxrTSL1YKfchy3i0p2J5mx7qRTrBlk3LyLHE1He5b//5cP
HCnYWtnQAguXsI5eSa+av2XdrHnaFX7WWgBZFjGaU+0AWbse0bdw4QIuySrmqzrX
QQ4jmJP45Wkf6Wf/q+wlYantRtjdsfdRIit2f05+YI5MktqSEuGtpVeXa33VY798
SrSb9GMiXSuW7ZF7S0fge+vZ/pxDtC4BAZnxq3Hmd8RWl/dybZ7NyrWhuKTXhwd9
n+fq8nYEn7llaSZhy1G5XBmf7b1B8olskPR0wLMs5HxlzLsoBY3MqXUdsgwVXXul
VO7rfhq2R0wqgcY3qbXBsenrIlGdQ19PY/ZW0E2yNT37v8pLQ8ey/ntB21g6iuSm
ptIiElgnoidv9KkmkwXjvlFZJQHAM7oFf735gFeClxzld0z2HGYwH5xQ0VYY3yVm
lzBUG3JhEyH2fvB9+wfz1yeifup3Kw5xrE5y1RSfw+JgZApxC4NKR21LJteOHtQs
BGATjIu+tVHQw7b2r8Mf6YU6zxt5DqAP2Tea3dMiLlC04DmexEJdu+BJhZWYcEJE
YO5hvCVUNfYdMud6VRIiUmlqvcPJzbXL4DIhgtFGZNUC2rDU89HSAzG9W+gOKguk
50S9sq40SfIpwUeW/KE8Ybvz7DyA50QbGWIuJghER5JiY1rlF4oYwKAUryO91YNM
709mC65GIbjINwCuIxW/8xzW4NdPirU2X0PPhw2CkQgY8zof37kVR4owZyvSSxMH
NamdLgjJ/rysxF3m24d1ZjmZmU3nVMSrvaT9WA0WybpPaiKOSX/3d5lXT8aCCI5b
9oI76RA3FBqyH2I2Gc0BEIpAbCxotaiJK94Ah9X9CPaO/cEM8UmTiAhYN+HSbF7j
vjOZbdCSQ++fT4AY4Dwo/BAeo4S8lZj5ABS/gp+iFzqGPqX+sQ29fIelRfC2fx15
Vqv/8mLvAQBbi1PzLukb8qhU+n9TLDsCvvIBTPwO75JIKiMIDjdOy8hglsSOsSmX
kmoLR1VjtBjzdKRTC9x19uOy7RoKRWJn3wkYKCQt5LJwpZ7mF6sgmZukRKkr8DJi
n7ShTVcSL38CJ5/6uRk7XVf9xQKMuUvMfLSpNSaGcOmkQ0rTkrqgirVNY1pgdcKo
VWw5VrAz4PztYL0m13g8Uf2s3UEVvhU0HZZZd912lT/dKMFkBzQr8lwEVWTMh5JY
kXAXOc6l546EV2KglMSc+ALN7ykhWidUnF54ByoxrmrAfRxM3sJhsG1medLZoD0y
cdPzlJdwse70Aj9Z803Tz+3H+CO+tpXsLPKu+iMWRglcxWOgMTp2D+PQ6thknsGj
J7TV4kO+lKw688XNV+ybbN6t9ctoJ+b0wjfFa7bDE8Tn/PkxzQHoXSEhSB2BaRzZ
eX2rADtnJB4byy/sD9RYfMeNAtSn1gVGmyZ4sRA3yCr7DoyF+GDXR22sgt8cXGgl
Ea/69O+1GM4WE2vTZA1HvHxgZH8ntnsiNss8ibY9vWdb1asY6C/5RkD0l5DxWZdu
MVOZW/wWqsKlS2Ik+ZhgmzSWHQevFJSlmEFumQJS2Bd66hsOlaFi787fJC8h/sXC
tUXBfHNXZm2gn2Z0D5nWnAGjJWL++lyu6l3D78zUqVRbPlpcuwMdp9q5veOGSRmz
Cy49PAQ2ntV5AB4oAGmRhjy/iAomsmpNX6EVC02MAHMqrb6p/c3HPVO3UbxJaTr6
uDMjwHAMAVlilGzqcg50gjDhwlEIgvaeOx9BecsCQ+wKbrEkDzkeoIkam7+aEqCA
vbh2Rz+6uExBsu3XGk7XmWHLv1ruTG8wmSICK1zSuN4Fc2k8dXqksafePfjmFmlc
sqkROKLeGU4lBl7O2WtThQYycu2DeQR4hRljnCL3YhyojXTc51oWRwDmV+NjG6a0
jNRI22B/IsKi3CwbJ1j0+ciaO//Jtf47NA1R/apcck+/cS228XKbZuofPdP9AJSi
jS9YcX7uO8qYoeUXhVwahHeINh95JUsg9nXoQdmAOnJvQeG1dzzwkliy3brhIE2N
yBkI6m7jsfWXbSH61nkfSF6+i2T8gonubMRrULD0mHHj+yrU9XHtAZ/LzHKQ0+Oq
K2k41gq3d/jWkfM7E1TJkAUlN1FM14yFQ+dwJACVew+vGsiAbw55+LLlzfZyMiDb
YmP4A05E4rNFu3E3WWxXuXgkor1JIwDCrnz6fVNBA3NDzmcsyXKthACfmdtxOENg
eXH06fsC0OHBxZKaDoO6ywIUlJYQhw0PDHOh3+zf5DyRkYQVucuLHzNfmU1ngnPU
EEzeXqBptrGHm9cx7KLwRsaZFtak7el9tcUgpUe4yVNNrA//h08qGbAkPXeKkbIv
YHEmz+UFosTFsaqm10c3BOzzru/0sHooONSJ/ZF5S3SYkkV9J1o7Xj2Q9Alg4F5E
mmng1UeSCwXsL79wkpP8oxKl/DWThYSydFZK3OehHuI53ISOlpzb84BA/gJfdl2c
N/MJbbSf9ihTtV3wvV3qf6WtNFbS1ztOJr4cuJdEY3rlzLP7M1mpq4nufLk/TalJ
0nuxwC4s6wNRIk0oansvXEWBmd4VI3yN7GT6FtsN/SjGdJ7I8U36i0k10dQftvR/
MVmjt+7NNjHoOpns7mpAGFxLLyZX9KCeKfG3EtQWYXzhVMRTuZg/YNA8DxgyruWv
TE53yefXl83R8CpZ7BRoJMRCvkcG/j3axUVKBJniq7p+S6OwK/DcSIvFY6weHRH0
vpaavjlrQvg4HYlPwxU760dd+F+Hkhs/TxaKNpV4gGakBDCWavPzSiziVOOPuduO
p0zX8pTSnG9TNJFp48bfSG3piDfwTR8REDKsMq95+Qzz0BKPHdfzIXFTf7HI7u7q
AhKINfiIU3Fp3WW1BUeQxhfS0TF821YVgqkLZFvNghNipGsfTDnXcZ0QYw5PXntN
b+NbnuREzFpb4mqIfEHL2DT9k2GPHRhDrI9DKnVPHgPcJ6y3T42aZ9EJq7Bva3Ii
e4mLvhXtBto/MJr6oaoZv/ajwSg0XJZY4xBhmhy65H3ZXHA5Usx9tdzXxp3y0/I0
/Sul8qsM9y1HplmG2bTmSj2n343Rg4lZWi2qBlibmW74GAG3cL1VzXK+L7z1K33d
3KtBMwYuUpDx1uYniI1KkYjM5ObMVMVY/K99MktZ40UIwkTVjvifpZ7qiy1MHLo/
eSwK8hGSFNK+hai4moQgFIdxBSKxjAF/+R0TkQGkY6uOtBY/Z/WNg/TSb84tWmwS
E8WUYaGD15I57AD4az0qeaCqwTF77hiCepmIO+g91t6ehVXTwAGqkzjT3ME0Nwtb
Xtnx6okWkM9u9pr2pXsGuh8Vv07ch94TKlLsu8am4ob3l5/0RucPOfobHQ8ZHLWj
CnkPeHR0be9GYd2Kh+RSBvW/2KCF35nITdJHVac/hitlhFDTJVejwEbmXiwQ/oPx
tIT9L33leP2+Sx+oEj4TF0unK8ZIWTWEViP9bhIrM/2Ev57d7RVxhd0d3kzsjUot
WYX8413o+1sdPM5Mp2XM4X9tSze6fw7jDvIIiZEXxj5k6P97m1zEJQMVO43KBT1W
anz3u2l0+YN1iuVJz/ErxmFEnBlyHfaQ+ceWe9mL7/0vnpBHsk11Y2RAOs7WEmNQ
9roMgxSzZoHeIrwOMH+CflJ0M/oiknhDgQx2cpNYgSNk0BKhiGfDUy9Xy3o+Ygx+
aFg7vV8JdGq/ey/e19bNxbWo3+8NC3xnJXOJXGNyCNfQ7gWWGDEQ8ZvI/CLeI1kZ
B6BqvliIK8ePRHIPZwhO1XITILPBXWO9KqKt96FzlySIL0gxlQ6XgP8RrARnzGCM
Sj3uU4NnnRA/UJPlPVoZRe5hrEzFo2e3o+VeVxfy+laObEOfiCKb2k8imskJ9wow
WM/TLLA0mCzH1WcpM2vfhd97Qw0Z0mYLUE2giXy/AgMFx1FdcVFYcEFNiul6/6Pn
6RsMLh8Jw3UsEbnZsi41+YrdK+0f4wyrWrRbRX+KF2qVh9Q2U5PKwA7C25QtvHX4
jhmC/jP9eNm8qrpvX+UZXo55/pHz3pdKnS/YqWQUPjH5pVMwHL/TtqSOMsER2J8W
YG8WiR5yretM7gFVqEUKaRdwjXbpXGnSxqjRViivnOWS/TKQTYJrGErad0kiaXjv
JnNcwgrZK6CUFYPwCd0OsKpmS+lphVFncI2WpElGsZoiDNzH9FekgmXYLFZ1zLl6
pV/0xLRsc4fwtXuRiiuRvSCz6HrFz0f4XNgZrUWU+FLXcfK9F+//lEi9H/eRqIWN
+s4tbdix+S3whvY0JymnL9vjw+oEyez+69sbtrqvGFJXY5tpFPhTDajJaCsIEB4H
Ol9xaMyTL8lIkOjFhImLQ2LrcPhICXEhBgYBRue8D4zpAKp8gGBOzvaaviVNyzM4
gPULk2QzITr8DdjTGTMuX3dD5hAl7D19QePAN7KEJlrxLc3mN5CThNF++cQX+fVh
FfHZa/w9QkZRIaB90fkoFMZpJUqwQZVy3IHRJ8OBx3ohDfMsqJ5UC8C5iXnW3sf7
vfn9ppxK9Q60WrI3mfSjMOeXLSDYcuIalxPLeybU9VEYlM98B+txhXJ/Uj/rZPuG
ZqdLCryCpZzAxeTdfHbW/KitrNReTW3kEV9MC+2nlQcR9phxaMIaHg8aii/sfu7u
eGWElnr5Tr0kuYioITHhxnQntm04MuVJ7mHKSGIrtIwrOsvWGIjpzY74jRnKNC9D
govvga4TA7vbCQ3A+l4u+6E16Q/xSnnhRcunwRu9MQimIrVqusnE3uZfhDTpAQdU
At6sXPJtIFtW3s5AA9oY2gUpsUu1dEpmztZAUt7cXBWfbHbCmYYqZx9VHtWfLo3L
0FiOsP8/Wpmg2ULr45ySU91fTHUk4caslTdznKGeMu8TmXQm7K7R9arlY8GFyvh2
qTQHbQtqDBhjzFVDWF+x4OS8cggSIX2UDJeoLB9DNTPOCWWWcB+FA4Sk+oaRgYJd
5P9il/sq4QAj90tesFLbrdJA59z95ZWAsafg3ERAFMh+OofcIx26hrOWipgRGTin
PchQw+BGgChCMSh1XcTL9AHb7ehuck0OcY0c8YKxawuK+GRpufZlj1cCb5XYr0Sc
tNXEouMBilxs+4pr6hFnYiY3Z/qnkAZSAXYEI4GEWShjpPbqVU/a393J15pogBOC
/ZkDPxbsgGu1Ok43RYRZkSPNaM+8rXbNKapOck9CD9c4v46t6Jrn5VBjLWDM3k+4
tbQeAske0u3yi/qqIsnyn31AFcq2js8+ZbhQLbMBQcMe1XrobF4RqeNhKf7PLrJc
UJJsOE4j0snsIEman1lB8HMEH4iHqLPHas43zS/h0T4V9EwlA3D8AyK86O32w9Hi
3ef41XWk9nrRFo0EZfqqdZCxPyr3MLSNY6Zg2Nj6umy35RMIdtdvXsGbMQEORQR6
J+ZEYbf967qDhHvlvCBt4L3stlWgkSj84GUi3TgJ3guR9PSydm6jSKhbQhwTLsEL
Hvc8g/8C+wW1EZZwK5VYnv4KX6GgPrgSUxGJ7bC07qMSjUf6RMe/BrCrvsmahw6o
oHtHyn8Zbls35y2MG1s9aXutzZv3eKTZIDlgOog5KCODYWMc8/Zqtzl2HPWBeQel
WX+YuFOnROtM7rmFErg4RI9OLNgGLz6AYeRq/sI3OJh1miKTuWuYcYExeqdZaNc4
Ggywgasau7mYCCh54UMmiGmkMrfWM1mGXs1hES994VFFyTCTb+1HAnrwg/PeUGvQ
NciR86Hnt/iI8uxSdexOI9xby+cFrrwNV4BDhg9YQgty9iV4PzWm6+/T9tbSLzYS
NEzY/aUBgWh0gkJ3/HTBhy/2bEg6H2gvRzxFs00jREdTmo4TA8IhRwUN9Y0e+pst
KNk/RTpgMDTJ7P1mAClzqzFKYN8ogmUjKea4MGe3bct5eDoo/fGthliyhmzJIllG
WXLnViAUC2wMt8d5mgl5gMkGP4ExCZWdfUT7h3nQivITxsP8jD23V7FnBwQHRWFJ
wHcEDuvYjg1C7sRgnCSumXuDeoHxYUJ+ckL5O2Nk84K/HcFJALUt7ycY2uVl4gve
S+uAiygU0fPmv+hkbKiyKtrQOYvI2UUds48MzAfCJknSBOua4RqsaGuCHGFdQm7S
Cch9E3RB6p9HGRkwEPTQOt4k/8hRTg+ceHGfcFRmZtKw+WoDxJEgHFENFfPQtZ1V
zi40eMfzdwO/GdwjdIyCN2JToSPJXM2bINEgx4ZGfZgbmEYyNEiNFua0xeo7IzWq
foycvjsZvC7GUJn48dV2pO91AtHvph45fmdzuyjfWIhB2zgneGhAiBPF3+afWVyV
fbtpnJ4NRUPUODiTrgzjknUj/cR402ZahGn2/oZzTkMcHWdjtFXP9ka5rnRF0wlz
wC0Nv5skx9Lw8sICS0rdmJIbic5fxiWjmD8e2afTmZsWxl4qNQw6fit2zroBH+6s
KQP6TuhCPGPlbutP45VTaiOCsH00AbYekphf9ltMPv5X9JAXGQDYFe9VX48ha9gK
FYMRvzf4YGwEDRDRc6qWi1JPQmuYWRCS9XY8oqROnyQhCbExE0mxZYe+Ia77YKuM
ghBvd7z+0Aj0lAsea/Sp+i06tr/QNrrcDnUuH3RIm4TM0euaW3q+aOUdPsGwqu80
jsHOmARICL0+jL3bw1O2UUmZHxWoKKnWsGwcPIJaCRlD/eUPX/eLiNX5QNTSqZcz
71Ahxwxr95/AaXVQ1GoQBR907Z068PabVvfKSk1z9pbzajUziazpxcUYUMy8Unza
Q4T717L0lpSYCSp4KqY+vPMlbaznu0DlGmkQlEbgPFyyg9a1hH/Ja0a2NJ7/BIDl
7kw4f3mU/BB9SW4v/DyIyubuj1b94ZG5ogdj82f3k6lKkZn5KJRnJ1D4XFUOSrZG
Ag8+LPI+twTelhWsidCGF7Lbd9mLMTrNf88lZkp0+k1iswI3d6sNE74C5LFYpqWq
LPc9t270+bXuAuvrkb8YYZ+iAZJjRxMTeULK0MhFSsTUWafjDgeWZeDJnqgbp7pb
T1s89xu5ciq2egLHyyy/NdhtZlAvSumukhV0ciLADq33qth0eEdXUe3wHE8sNw3J
+IdL0QuvSemcvlezi6X91HifWOoQWyJLLNoFDaSNeDdewNWC+NHp7zwrfaFZ+Cey
67NjGbM/bzWg8/cjikXBUpnyscDT7gvDHbQBEm0u2p702pnhvBAZRCIuNG8/vTO4
LYhGyGE93kW5A+bGHIC2PUifjdpBFA9N6mdnoFnFnpcqFOuSnsseURQiTUMDdzAy
5dH4grJRqbDSjIMXyygq8lrBGs3bUoM9fH6bXkIipCL66ZbtbEPE32G/oe640inF
NVqn8e4j1cuSg1Un53PNu729KgsnezUdtDxi8IQEG46wbnSiRWo6/fw7HGrf3apu
vnRN0A7nBGiuct8xB4lV4uWfUb+wa3FUvdG+3V7+Vr/ZCw3Cx6u0XNsj6uWU9b4U
vX0jm8HmcERX7sBPhpU7Fj2iPeVvRKiFujvmGYnwYZJxEEDtOMQAkN/qP7devdTK
aNTGFJch6DwkUf37cchf6yTRzQxpTbwWlafmfiQENQ+/M0Ri4eZXBICrrRmy5JYb
JlltZBL/Si5DQ9k807jSlSVYewnTI7gCJMzDlXfO7E+1FEOaQDefl8Q+XxWUM0Cm
xMqw+55tgq44u42r7duGxR9CaMTd45A5na4UAbrnZklcsLGujvIoFhxvhAkNc3H2
gvyz7KQkNMBdaQFQyBf2TiA/npK9A8wQjaMEsQuZYQb46E825LiewaUMzKpQWcyo
2XavaUSVIQCgU6BST7ZQZAV7WEbx5TYcGpdBVPBRpa8I1uCpGp2uuPkdgDUJmTs0
b/GlP7c9cdxXnFiUcwWf3ArPMDQ9lVJvowIz/FVip9ZDNm+5ym18wv2PIMOmhioo
FUvdPFf8uo2TrTB8fYyNdxKYxbvJgeY9PUYkAYLrAcQdE1cFJhmDa9hSQxg0312h
NJMFtVnKIZXpduo1wzurS8YFuY8D3EUyotN+rQjfiy587/PnEc0dezbgCwJ0tvHp
mfisSBmJ6hFplVv8WpqcpyJOZJRZWm/liwr/Jjcc6eADkvxRBAtiuNyHS/Da1zWR
PsYqEYiNLaVXUVNyGexedp/4k8kUC5tT194DfFCboS/k4c+SjN3Mkmk/tWE4iBmE
8/wFzRPc1a7Z28yxqOWzu09CufF6lfoZqU1DNARiWygSXneffHVBa7qdTJDQ33wa
z45wukRIyxGr8sUdwV2LE5lpmHcE8Png6DG84l4+iUKSgAGxUnp0acz7S0E2eS0w
VuNIQO2rpOrlVafhprMeLYs3eXS+zYN458EuQ08DZd9xTkhbdvf6up+qT5W16EAK
sdpQay04UrzzmfCkdq0fwziUpJFSKR1A4s9BTZeY3QxQ8xr0AbMt26nrQU/DlUlF
a3qp5A/JYXAe3i95VvEmd/cFCIpaqtEZVJ6o1RFlNBpXJfB4HZSsirNpF9/k4qXn
RihyDoExJ+uNm7Q4kDmNvlmu7SzSWNskut69uPT7cx877t7okMqDTR+usMpzfQ8e
yZfjsRvxi173uHJsgnEvCeW/oIKA8UF9Tg/aB0jl5gefq1zbid3x+ti4ym5XTHFa
kEEO2fXozNafFaY3Wm698RZoHyhPKgqpLjs8cxxUFBUhIpGlwR87Onqj/FpJxMqg
nBfXOePotv2BjOpGI8tCUIG42ICWddv4W7n+hkbnGGPR/HJl5Q3Uleu3ssuPxJ11
pMdu8EtCCXRDKNh+OIcMrBHa8/gXuoECh0/LWTnKLVwIvXkmgGB0sbtrNoFslYX+
xabDVRQclm2B+jWdkIBwZrwWVjFqQawD6RdaWWXZWkrxLeVPwYf+19s4hwQh6IyF
m9HOhUdjMpJhyOynwMru20LeAmDaadfwDyqmAMCtv57pafuPc7ieJGB6lWl/6Qql
UFx7kztQXqE+C7mlXkE89nsZi6Dz+SvnDMhdU4KAsa1+Mt/3E0PLlgzgF0HPA1WU
SSd1b37MhOe+ueC7nQKVKHr88XbRbihbeXcRXcX7PYrJpUSC0XSApslXOyHcC4xb
6oyKj11jFqA0ydncNJylInf4LG7w/7MZZhgJ6BhxB3BlFZ9onBlObtLh6uFX0nDM
GgurWMuPFrW6Wy0bJn2n3g/j/efdGfspTEUbKznm+5eUUeQdHPZTIzqkjdHsDrgW
JVJ/ouMQnnqQmwLzUTaf6NoWh4LneBLghp5q5MIgRnbfk+mo8gMIhK10hK815KQw
vVJInuVs+xqeOgPtGKtIlA2FSkqtIHBGdvcbyFWLBUbNGEt8UgNTGeSHjBG/98Qw
oY+QTlbBRrOMZ5eQ+m3Atxrl9DQTu1vuYh0xnvwhhtftVsel2Q4p3Mf3BT6BQ+jR
JsDVmVKm4QXiIpE5u/JpkKRwXQxZ5Bv9tPOtb0eFFfj/VC0ZSrkYX20ABFqYFsqo
JxbKHihEJO4CyPlSOZzCqskxlFzmS+irWUKaX0i11y/IofsiMfWVXQT9gzd5J5UD
QQY3lgtXH6ITj5M3p1XHb5LiE682Z4y7M3meCt5Q0I4Hg8WeImFIWDhVGPcubvE8
sKODUxJsig5YQEbeQZk9NLrayZUZJFS0HEb5TkMn876tOT+/sfKtdrKntzMOdMpY
K6d4C9ldh8HuInvht1aAhK2JQovzbOKOnW/CDfnBzV5Vyog68JpnymDHzGMMAvmt
Y9hHv0WmJJa5tqhobfQ5JGG5dvEHhkXPIb6I7RnMpSeuZHDbPoJ80rnAQHmrKonq
S3yl+6fS1HQS80CE7VKTVHKeB7aaHDG8NXolUdm+SbjA2oQC0QrcCXX2gl0AE4aa
flxNwTrepJZGELjlHTq79CVOl/KQ8DL9F0j11LF8zv1myUexOA2QtnPYCVn3ooZh
Lk5vgWYHLgPEMIUkSYTZ0UpPTbhcwzZ7uN96xNHMp6QLV1o/Ex+6odx0ZF6q9oNV
eKjgfBJoNBze4xHn7twBj4/Htb+h+0Ol3tFT93kprCFwyHu84c1Nh7xUcNcKZ1pE
tZFISm0GVgBeodb1iPQjVHsH4HN51Y9GjbSPqx0WF9y9r5q5ef8EyKm4uFzqQM3C
zK0C2/Hx7GCqFqJ5UyVq/OGq4dXXN8VHBR0H/73/4wcB7X9iFDKDuY1336i6J4e5
lTW3wMFlcLzeZ8xTJifYok1d5wU1lgyKd8Plsjuz8LWy00lCqOJjJc7dQwqAXR1I
8bZgQ47av8TDNwtwIvtG2k5D9VaGKMzw9PFx+65bBTDYfi83qPGMOSLCg93BZBcC
ZvtvUBkI5K7Q6H/Y/iuu/mX5UshMU6+sgKXaQEHom/Vg1zPLzY0f5nQTfv9dVStm
nAmJ2heoDp2aKzcNm0ZhS0U0iPmOVumyAapE4yIqTPHeE/itcjEX6hC9zWIdKhU3
mEvg5lGfIUojXcxLqfRzLV4qSKFlnOrsIZ6f7N+cy/ZS3v/JoJ7N5jTLZQwEXyAh
90gkcncmU4R0YFeWD53wIqzTyvg47451pVPBnPwDZ3kfS5vhg7yVnwncSwQGfbNV
yzmfDGs/UKrQwVu5bmflWl26fLPiG+HbGDo+G+VgOaxfGsf9H1J1O3MZ25ch0qXZ
dXV3tk2EvviWmiN3cGrqtCGQREmUxIHjVrRxtB3JzK2UKLKNYaERgAl/ZWwBfypD
oY3eR2I/Ha9KrAnEmi3zQGgZlLirVWA3NJf3/LXcyNu9mqbdCu8Kt8Rt5zmZdxOw
NLIWCUopiD7u9Wbnqv+lFfmcOl3EmFY0EWXOObcTUy6O0rkz1BIhd9mG2RC63j6x
8yJbmVigoxcMRs06mnPzaoSbZd+n6K5ohZx6ni6Ub1pSC+RIL9rty8REvSaJ4lTq
3U0HGlYDlHRyFtrfyGSZ2fEUOjAUqqUO67+4Eziu+91ue+3g4AJQvLQ1/xXOtkGJ
k910Q9b3SKUG7GDVZHtdRLBh3D4LTQxv39MvOWKVpZvGxqwTZAA5IjiiBDsQIwbZ
jekXmkUarruJgOlu0UVjl1b29lc2PjUpha2AOu2sS8Z4md07BuZy40OhyKoIV2Gk
wndFqLX7nrdnI9m2YwuP98wAzvDb30v+AXdelJY8E7o5vtAeYy/ua3iKKnmTof85
pFyDKhBs7aGTlEFPYdnq7TjcJ8CRxnrbcD6dR4YXTkDLGLHh6FEA6QdsU+uQIVKf
RvZ3SUWEvTp3jL1t5VQQW5NvlcX28veCORpgAHcRbqgW6rBFDXztxucdWp9x/5Lm
IFOxttnv8Bbxm7+xoK77zyggGAjSK6cnT1SbnUOdgIVPbos/zLhUiY2lACqUMmvg
eFKXgwOdw7FCrVgqYMXOqN8JIi/vsjPeViraS89SqsBt8XwaxJQ60Lz484BKGqhe
eayuc+cZvIRIh+dd2vEaJZg7WSBDfMg9UKQIEvq0CgCRZh22QclFv4GTg10AXiwB
bbg7Yhgic5LC8YAZHhsg5f3hKf4ESjsym4F+/3Z/gBsKIjIe6ghKD0LBqZztfsNK
3JQgUORVqro5zH8hJbjmsEtXEfROYcty/FUi35AsZUHeKvhRK1/2F6BvRw0iXSoD
p+V43V5Cqyn9BxSYP18VuhxXmnIRFYwy1ejgPnsnq62GPaHEz5JFCcIyeTPk3Wm5
FbG4ePhsvg9Fl+zSUqIhwfQFXJzV4Ma/S6+jetm2uFiAyDthl49HrNKAM508C5Jt
7V7ZYJS9fjnmIx1+LTY4Cw7U7ycFeSrvdg80rQDQwil3G22npzbE9hwC8oi3Qxob
SgHTToj22ZkvNkcg93VxNZjEsInsRrCIsfMgXqapZYRmF943ljOJ5613w4b4BMPq
7LXv01h3D6kcw+iDT7T3Sf8qZmphuz/5DVb/R1qulZv6qThyF87lWDzRrjvHib0W
ABlFwKVjgdKf7m89+tA0xugkImfCyztvUXHlAk+Xneta6VDINmIV4IrBAHQM5CJz
MILugdU8dhoSUQcljuKhWT4f099QXFI21HxfuTiva7KQI63ZDZYM2zWM1rZf1Dys
L1meXCobyFVGYrc0jaTTvZNKZMGHVbppag2msNsJOTCalhGzJIFwIh0xi+swTMEY
BAa06kcv0W1P5a3Vg4kM0Z3IEPuFBrZbJAhC0gIAUFwzpJZLxfg5ND1mm2Wex6Eq
6BHBHaWK6gHmmHlO/jMU3cYWx+hi0ikWHU8LQJl289QOrRxRj4w7B7WPc8taK+bf
AQHBd4MYYG+ypqhAIkmyeAw1FAjOTcJbIPAv87OA8FQeanVLhzqoZ0dCu0USvdfM
G5q+by18twGytl9RxvjNvZv1bP5Hokd/lB8JSdAVDBVNyMzTzEvLJg2iIw9M98Kw
ohX+S25YIFeJDIVisGeSHr7qHahxIF3qU8rzsy0v+l517v1YjyVWd2n4B/sO6F3X
5Dmb+ejFsDYlYff/yNTaXVz3mAfodOj2nT57Os//82uTJ63SJEmLL5t6AnkXwNom
pAtl+3VEl0oms0YAqn+SN/WZvBkXrV1zrJNsu+wXAiQSRR4oUkC9zSika6yb8z3X
afd8P6JMce3Rl0ZN0LPrqAqvfZeHiEqKJWWAhqdg8fsPnCwmh7Y8HLu31QVJYiRZ
QS6QrkpjTNSNbEPwbMsatoUNxoVAnkXRxERYUH/g1HYh8JWRwSaosJJ5fzQIDqfv
V3oo0u7f8ho4pTeemXcR9Lal2e61o7uDck5RbPHHe/l+qTL/Iuz7xxTFSQ71A3M0
xqRQrk3/qswaycK8bDf9ySyUORIyOgSac5TqDGnAV8D3ZNfEb9A+l8xC38nbLGhW
j2zwHED/uA39r/ar+05o0qYK8adx/1xgwbVUYJG1JFUTx/46xFHdlGljJ7+3MP4M
M9L2LmtNYKGmzHzH1Bhh4rir7EdUfaXRjSn9H9ajumd1LMxgWW25YwIenlTSiNle
Jg4mXPO7psZt5o1A0tB8zJkXPNpWryREaqon3Qb96UvwRgrKQmUGoRHzbZUeFaz/
sshNiLeVK1E6jg7EjxW4ahtFlpnRoSgGbNcvanDsEbjw8KhT46WszvUuSmNt9qV5
YqELHa5ZLbK4hZeGYv9zo80/qAOPdNzc/qnTU9RXrWePF3tOOxsAzPnBwZlsMoIY
oSmP93xtHH0COsd3nxRWX+6dYyTYKtMfwDDu7qWro2LBA2819Ke6zEojvZGb5EqU
U4U0diLaaVWFZcU5/JYPC7oBKHVAipLKOFTzuBn1oIgcgShaa5qUge91NNhiA7Qt
Uf2TOcx4bBUTbduBoM4ytHLLCbcnRsV+d34i7mTpNoFMRUwF8CqBhPu88JNxIU2x
MNQ8q3qRfUXeBjGGYNpCjOaLQpzS4LKMNebJdwlCUkSHccY9A04DnSMmeJtcQrIu
M5UHmzgLtQnswKNf1FecvsPoZWbSGU1QjeAW8ysG0BMxnJqZnLzWm5bUoFlbKRIy
z10qa7aDFBw9vXtoHN42Mxso1f2lngtvrIdP+dhSUWA+2uUrS8a3LrW7st25/cel
05R561MI6sa57ygyIwrMo6mxP/EKdFoJaSdTBeGNuTvGBS8x98/5odSeQemlwtkj
GLjya39dpfhtoVe9jBX7s7U6Ne6/C3FlJLxujsHd/iudSoUdSSyvAB3qAlS7Q4hN
/MRsCqGyMyfrqFNxahxz8ZnRKUJNKXQDHzoRMnLiuV/UQ67o5wAlTtN12FKJUFfK
cRumFz7UAvRppGepyxc7T8Gd4EKTzTqGctNBm+/hWpPBPiBauUwjH5juomO45M9B
kWH3dezonc8KK2CO6eua6a3KLe/UKF3M10AR56aXSFVmnzLG8aUM1tiLSdPWdVTg
kfvYI+Eq5AacWaOaRj31cHkE8xy5V3YGqVmPoFpUoclNJIaAzrkld1hK39hIyvCS
0jRa+kN24CSOVTpkY+iHoOM+CnsD//YZeFpFfmKWHdRraVKR2XnsfNrRzK4KSdmJ
5J7qd793DfHmXP5VL1Siy9DP/V4X7atRCHflDAU+hJQkKTB/pNHTRm0bjF4akAf6
2zBs77GMSulZnbCDUWOsfLnNLw7bNHx9+6zraJ9A4eZn1gGHk6fFxLZBVk8JaFeB
e79+tzxTAJT183Ix2AYFdBs6+PBJnaCLWFBByXwcjSO1+araUtcbHlx/bfC330OA
Tj9KTS59zsg1Fqf9stSs+G6l5fU48eFJs7NzUTu4wZPDog5EwemFHtE3B7i1+bJ2
CpAPd0uO5IEpyD4zro86sIjgLDgpr4zPR6Bll+1c/7zlWaW0jYgrtHO3DydCqGYc
SIn5NA31y7bVOD+9//LLLF8qk7lb0Yn9SQJ6k9NEUlesIVdbAYDvUK37qrfKLHrg
rwxK/zIQtQmbBHlE/xWUbkeIFtFJmXoK/jEsmfNaZ1uxiag3mQIR001uGJQi9n9V
IR1sTF38xrAaQLM2jUWX+rvLrBOP+jq/6M8LHi3+xQRRKp7Rcw+sbLrc/ZfVW7mP
ews9RA93EzGghjZMo2tY1Il9e115IcvizXt3QNwG61TddJH0U+/b44zK7fZ9Uuxc
CEXqAZblofdn7FJOYM7imV5mAWoweem9PWo88dOINGSBbaoKllkdFobMEeJyXpkg
pUDVyKDLuIvW0kdU4eMdoxYarfsVVujXWvjR88zi3ggxPcefSculK1GuiUgAd2Tk
G1xK4iiDmQe6Ot4LbhSM0A7p8miHIQDuejfGZy2tqw1cHP2hdkJZvH93Ijx+N6Td
LYkXLdhl7qZKWHIPExzV+r6wxHqo5Wz9Ci7/IIz2SF4PP3D+q5Cuzr/49nrGlOlb
D5xz7WbhW4jm9P5oV3pKHtCFkSzQUJP2pZUPnnZ0o1Uq94mf6NCsZ5zYE343XG+S
mLFqSidBdCeHJ7AUeMSnFeVpCcn8sf+WqQGdxe+494qWSVEI+nOYUj29T3CTraME
c8zh3Ux6+GWVAl9K3nn1Q5kQbfwo1OWUGcDHMrGfq0WTfNX+9zPUKFDmD1okKiP0
syad15iXkE4Azsp0aO/CVfIALvYIFKuawyEJ0V340bGFH9JrSoATQWzKSW5N2NQ+
qjIk1w9D5cy1S4Woy+x6Ib7ffxBfZxGAWnCSI+S4hBT0uQu9k5OgQMr2IgdS7mfi
wVhhRce3ZUXgWOs9Zi4uyiVmPqOg3pSTHrIn6I86PSN2SrZdcQIj7RDg26n602bH
biwcqrjRqUXKSo2cAQoPPxs/KgFodltABKEvyDTXzSUjTHg/PARUlXNrP7ZrG95Q
e14sECDH0GzaGA1CXRuvULRAMIcsh7gIazL6Swvd2IZRTbqxC4IdxKi5RrOnK8Od
EekoS7W0b6fQ3G0LVF+XM+IMO538l4Wbr3WSF2PIWZNIYLwfSswtg3WMYSpwc0EF
TjsR0vzdjIOh9Hr9W7I0oGwnSzwbvCE8oVMJP5xLGLsh+/V0xGYnd2Tr1llbov7R
uE3xCvIu+YvU7tp2J2ShAOLZWjwg4mRnhIICETgJUxFBT3QPV+24ERRjm0Bfa3iY
NijXthn/yG3HB7hEn4bgd+URJOoRpW1wrYxmE4yZP1uzjSkycGC3JE0RpAn5d+B5
WMnALj83XWa0dtkPEDG/Suxe7gw8bPt5x/ocvjCJGGOceq3dnVD1UKBZeQggThI/
UwDPG0TuPupxuWM+t8nHLGuXjlMLPHb/agdPtm7jURmF36tKbrNpwRLWEO81+RSC
+JbWjw0QftuBUF09qfOmEcrxAMlnQLpxEzW4mmxeuDCBqeRvliVKd0GsaCNI7/WV
aRkYafM7WNu0L4BY41zGNWg1SQuG+pt79UjNNN9YfbP4OQV3cX31S+IXMmNYNGjy
jZOB+c6JMn6ZdcDGtyAOst8F83suUGqTR4uBfM8w46q4Lt5CZwT3TT7iRV3NsdI+
CsYoyJrDzXD9pW2dqXwcxadC8/rsPSB01FAwbC268/LtO16IaIw1pE0SGewz9l8N
MOgcnETdK6JtLAQqQ4e0D8IuX8p85BlGokyCVaOJQ62/5xFP70gpBGP7UNljN7zS
oyuhjuq2FgxgeO8JHxJZsLaegWl5Kkeu9t+vkA0aFH+b8HD0nlo8Tym5W27x/C9M
M0pNPx66AKce4OmZgwlqRsiHNiLw/O146M0DTjrSPYVb571h0rP1Daz7iFy6WnWg
bi1laORCJCdvUdOkAREq7Z/vpL63481Jm2eOfR0CpiXVJUK5IzBf5IuKU/1C/+A5
vCcLIiYcVuhWACaYrtgPEwf0XIEVHtQvmPx9T+OxE5U2IqvWto7xNukhA7syiMlr
7XRjWpLk2c16ddui8k8TGQ/ish0GPBAKRknasSEwqBdk/OVD2WbfoBcn1cf0aESL
MbvBTqx2UpvdNSHHwrxBHqLlUW/zBVgpWFjd42CY3xt3V2ojvu5VYDzfmDJY8o98
XL3LR7tl7amq0goUnPS7u0HedXmTENw03KWXCbG6CGj54pit6pzust7oYZCLFexr
+2BkkIQ1GqyoonUycK6chYPEh+jghGgmrlbneGfJa5SWmYeKt1FnirwYnZS6Zxvv
qjHaFCXPmASDoN/0xkuaKk0Q57QfoZqqmdHPyRoWEJxHzGjG0j1SiPpuB7VB/zIy
S6SREWSxnstNN5j6+dccX/49j1c5BYE5jI+y45Db13bMzizX6IoPuDDEARSe/rIc
onKvOjnVsrQcOP5Kx4WwdTzQr/EDz/IQh31ry9SurXsAuttYXxgpzYT7ub6JO0wa
1Kyapyn2PKSOFtIR75UXYB6XTN/FWywNBgN/SffASynY7wG/cQ6kA+pWNgKJfuMc
5UyfUeuE/b+MF+ZiX2qTvd1PjkpH0d9XErxJMyrmhqDEJv9R0tVS3B2xINuS7Jlc
WysifvctfWAQhH6Nc6giFol6yxoPydFqdzInkKQrks5t6ZmirhEDT/nZ/qjdjaNr
ptIrQOtwlD/2njUUoP2nw+nCeseklMwaEZX39M7a20eg5lKn2HXfx0ZyEuVyyxUX
9DJbpskrvQD4pHPwc0JQDVxx9FjkTFB+KnbBKAa+SfIiLxyA8Bvk6n2+f2iQHgiy
3u2sEW3J68xj4EeQq4oUkNu0iso7Hy6n2vdtYso6T4944BQdPDW9aAKrraXIciwA
2GRSpAhVnlBH2b+yFzXTM6m/m1yLGBL3IXzEJ0oxlD5lJs9ZnUyT8TkbHJU0AWoX
g4oI/79gAtZTO64hHppJBuFf31Iubumdybc/aD3nMQMZ4T0rxA2JsVxpYOjRf002
vMF3VeSDLbjUFzmJtlzJS6njws7idOWTug2U1mWFsQSFwHQqnlpLyr4sHD2GmR8j
jC6e0VZwUndSPKexYuM3/FKbdknNaT6WPKZMaW4QVPYrYZHkZ2QRPk1kDZYecVcY
r98iIlAiBOJX6YjXZ8eAJQKWZqsVbdissgdXttb6x32iPrp0XSLl1xHXcg6VA4EU
EGBXmMwX5iKPNewtV0FzMaaCUjF+Oli1LufrtQ/SEOX5pk7JKUUlD6KwHrdydWfi
hRi0K8up0eS+dqlGEQrrFm+cREXwgYEQy1w6ACU2mU3aMFuL2x8dzxiJkAj4DCjM
n5LwEyQxRKcAk497EzIXvF12l0xVRVmFcbqaIzxXPH/Hxupc95CGuK+gQ2XNZR7y
9wko4jIReUD749dGlfEb7iylgVRw54v5DgOhFX3KjZyoqEJ7m50T/c1MSH5koSV+
2cQCwop1Nomj/HxQR1tPjVx/M+uPrBbdJIGH/3KjC6Zmla1dGKB+dtLPl7bM6fVv
52MEMPWOzVRnnXqEBQWPDDstHxnHjm0f2QepvBHyaa+pDmd1AbwwJId4SVsXNALs
F8IANXr9MBL0tnm965oqJ3rRaUV3b05zoRu19s1cK1wyv7Lv4Q2Yc4rEFJTExgDW
468cBIO0uBAYll7WuKMB6uzJvTARMwHRifFXvOMexjSDmAuhu+cQdonFmQNjA2W2
foGQQZ2Ew2jD8phztf/EeE5O/WfMeIZECWELimW0N6UrpLnWgHBtVaxwRtSrcBMG
MC3LCBIaK+GWbDow0y/C+foRz6ESuyNIJ18An0KdQxbvwTQUNpMt4PXdl1EsjHeA
IrISE8uJDufOR1JQ71v5huSh6KTgp0hgfFjJ86+PWucwXSYx/YAqaeNupVwe458m
ugwpPkp5ohIKnj2MICpWL2JXpIy+3Dym7ntaiaLkEUVNGmnxm5gCFE1Ij/U6UN4C
ZkxpbbIvXg6Xdsnu1Svdc86cokGS7oBd7QAzNeleF/yq+mCq8NHvXQUa20d08gB2
XVMZmbTN16HI5q6BGFm5s2oOMpN6fze+fLyqyGuaa4ZSblnuA/vFxHHQg66JkNb0
f0+P9l9wICTSDw/Oh8U/xX0t/oLrOwAxdWxjVbfo+byJryqAONDWjyYuI0s9VV/v
DQuI7+M0IPO91jrqVKYCDlmTjLS/VvAFQ5Xy2jcEYiBMwP8BGKd54ExHwxxdKpDr
D9Eg/iFkkLLcqfnqg3dlwrGCgQG/KB481H0Hqn5uoXZk+NnRp4yLFirLU3weYfBk
QfhudmU8gGDkeKi6OUmmzOnFRAo5DtmVHrbDo4WHKPFIYja/GRSJwmYRCZuZmxUL
Gu95AhQCoMmmxNtuyzahLaNItE5qIID3maft/g6HfZXMTo6ohpK0d2kTBRzSsKmD
kKKG2OO0ayc/qMH1mPnubBmZrX62IHE2SwVfYhR5yfEoFLPttCCN1BLxt5xwNX71
UrlsnlBL355q5Ti8fhRklwye9ibsPUaZygw2FHPE/h4WmYzYWw+vKj9mDY9MIyeK
XXmHyX/R1z6Q/WFEV2AvlY0Lf8QqKTsvv68ZONRBagXCsGJJnxnizv7E68NUK73T
/gHqq8ORL/Jx02z5ckGoYKkDRaK43l/49tXcVfzTKI1yM/WjTnZsmnQe44eXZxmR
Flk+4/ZO0ITGuGwUH+G+1xyRuJONfnwV9wf0TuiUHlkr7LMRrVIlJFhw2MrCCVc+
Q0hwAhSBYGfllMulwNzeR+XGKWqy21DDc9PtoSXQuTmJ5a0hUIIcz1LuUMbdFVCo
ybsyqqJLFIB7UAAJ80uDFgmTG6GswpNIfmxgyCnoxMHiNLfP+bKKeXW9/En/bXAM
mrrY7UdAk44VVxxtk8lNdiCCDxW33wUPuB2cigCUBUfL1MY45gcb676GmxW26+h9
0tB30SI0wGXzwsLahlW0tE9uh5uhaBS54yN/yO29raPTrL1lkcjH0W2/kkoEnD4Y
XyEW9AkPy7fFI1zLuUH6CG1hewy7kJJ+T6Ezrjy1EuHw9jB5w5wMRPOUMEzoKRJJ
ArZAFx0jMCaJfewAskNS0x8DkIcwsPTjmlxFpqDVkt/QqUaAGINodR0I6m5jwKZu
UYLpdhBqk+VLhr8i3Muc+xDDKG7FzTFmP/+WaoXhqs3gjtvBZWNB7uKNUpHJNzWF
DL+M5VZuBfHJCiyWBR7J609QpyzpwcQglzc9L96M/IiGK97qtk+IVx0aJ/rOwkuN
8rnB7b8w32LvBOeaGFoLr2H2trAXszyosYJrJKdKdwC2xkzPBFaz0bVQddtzolYd
sm59UcI8pItTzuwbDnlLm1TwKdc+1SFDDdF7+M331O2HbX6xez55O1qLTJ4XZ70J
Z20WhvZw7neH+Y8UtH7JcIiWHWUkqYIfIchdZDepVp/YBcXqsAX0H0f+e5pA4pm3
tZZ4Z/DC1QThkIwqVqhkQbVWNJSFcSYTYYwvH7syFQDi9EAEx8AZPpIhK5SSM6rH
/LchUzUeAMGDTHv6R/zKQAeQncV10RlKojeYizYJgqd71fuFLpiam+1xl5gILQi6
OPKWydt+pF9sW1v+/vORjrVmRUcO3AUnDl2pNbwOTqLzmcxFkXO2L32FqMAwPL6n
TJIBlVQT3yN9a6NyzzQb35SEk8hTqdEY2ZR3zNDDtxSDOt579G6nizFeUDmaC7rs
i1rbKKN8A5sip/beLtqYPvA37Frt2iXZn7w1pz9cjFGk9cAnCcOtcJet73SqV8wf
TVVx9LgD5IptP8bqDLK3RlmwSsFyUcyJ+3RPOxe5Od0fAagaXKR+nsxFSOksqDVx
C+aKNpLIdh1QTve812fmOloUiJCGpBoBlZHlpuxUE0+2IwUN/sI3TXLkW6wXuZEJ
mePtlt08U84B2DWSga1kaRatKWSFpe21lXZHUFTZCQ88DyrFdumkp2Vl/606JeaM
K5gSXV+oI0XmdkUfBVRvYDoD4wshYkWfKto5SEIWjS4ePjVnmWNuZx6zSSY4n46I
jiUVNqturOLzAuCZq094Am7sacrX8QeXGuTODGR1yxMnsBxPTW+jKGALly2Q2tKc
vdViQ4sfV5LGPtvuLQP5/IFfjECvxIfXskq1MZSF0BuwFZxiXWsI9I5Qw4n/oaa3
uyonq02D7f7Y40/3Y/s4sLqjeraxJ+wdygg4PhRBYPWTAe4tSE7cXeB6ZbzN6SIg
Y6N84IpRr8+2ytbrTc6SRisjnrLBno0rySeh4baqyoUXCIJHR+BZ8bTPnQ9/Vnyk
qXTpMiKxK5xXHLbGturYM5mdjVXxYDP24+k0jsuT8nmQc57kMZZDhu4YPc2jL5ro
At0G6SdZuOGfhiWFu5TJ1p+wkVa5xrs8d+I+95ds/QRGGdhZ7GSwO9RgBYWAZLgv
DVL7xivQOn3MuULI9BCi9anjBFtHErv270kDdkJu4oXKl2/mbBVf6McAXpuX1R/2
zIgJUttN2Uz3P/yUqcpX2byrcPsm7p9mG+/l2v17l9tHmwktuvnquI5efdkem45p
blVbF/Gnfo/4fvJ4tUlRH2fQbkVAZ8t6wZwdemo2O94cTmvu2ugvUlw/rdODObWL
w6c9WwEA9UPhetkPAtaG23o6ZVZXrcEVyAWxiOw6+6H8vqRuBNkmxxh0MJvr6+Kt
4bQKk/j+Dvs6uqpekfri7sx2TvlKbEWFFzBI3buuxzewPUUFUlDJl4P5R2rswOQV
wGupX2NqqQ/N6tq72weoAqC0EyvVgUwVCO4cIPJ8xFhSqhLNpblSe4hc8V8BgZVS
y0gCDTkQuRD2vCySSaVQA9DiAFm1f67EpO6mOgflYVBn/8d0+Pe0Oc1dsSORqi+V
pNN80j2vAqqt+zYNaRuEVvR1CYcqq3WZ9+Q5bpGWwwL9clhXwkt3lj8bpN06KhXs
ejnaMb3LueEmX9/lp5leyMXsgolnwZ7kBSokXI4DS60QwZ+U+p9O2eKFiZEbsmZj
hOuy3HaQWOWNbSYVH2+FOknZFpv0DDjqil/hlUaZopUmkrda8ZCmoIb9CyLX0TTx
mkTKjl3gqaE0Hx38an+O3ZkbUtdEsFaSBKz8ScouRyw1UTDFHMIJJvcFpBOOfPlg
p0H1IEiwfNzqbhIT82EcRtHi02c4JykRAEFEYXig/aORHHUoXFRMJsr40/1ZvT3o
s583d/uNovEthSLvFE0a06o6uU5xOUA+46xurtuqbr7+jcJhWsacSZvDs7ONUgIF
WyZPbDtwgVHdFxuUW2LtDlvZcX9BOruM63S+2zEU9GTfBwBm0JL5xF89FE5GAI2U
aMkDanRHup00N8Fcu1s8HAwwnbLNPTU7o7+4236mHjCpWl5kiejoS2N407e10oCi
925oXRBxNlASU37JawXyAXDEkg2G+ii/NyP/Ej90BEAkraltYboTUHq+U+lDMlgV
k0t7l2hwBVlA/wW2x3tSQ02HybFR+mXXLmXFXyVBemccV07npdYunclQq3Iz7uk+
fJb+kazQJj+4UU0JNnbY2rHEIaPMJ8svg1DR4R1y0ty6zA5dPmzVxrc9+b6kCuOJ
qHKPEC+sJkKjElRT77+pCCr+88y5Nstiy7mqtuB/fT1YjgJYQ5rq21zYfS1yPgQQ
KiXxMRPp0wbV0nc/MissC+3Ghc5U5NbEXiekRZ1KJMoQt9UhCYxJ+cn/M3pAZtxJ
CvPa8/4yaNyHO6b/nuVV5fqW4zA5pVKGp2M4M6lXeVTYJVFGZzbAeMaeyF1MZXUO
rhQ8SOyMEjWx5ByhYH16CKBixURG0ZlOlo/0shVrXWwIBePiwGjGNqPVaMeM5/cM
FIbbEpug6842+WvbQ9PIn9y8M5Opg2EMf7rH/jow3UdxE++yFbWfuwKsoWKaRPWq
ZwQbkmCaX/Lx71O/UpR3l1cGRviHxLwq7h0ejdbCkAiLngQE+Z9kXrcV+NvPBOg8
TsEGQB09VyQgMbWV7ujfx5z7AePLzkkfqKVFMrP5Y4s0kafct/1YmYKIv4WjM//S
1VgAHwX+UWEc4+rr+ZBbp8ajrbgdTSKVGm3KOvRBlhzjrW4CxH4S0cZVTVZpV+fw
76E7ONRFlrYP8lFssTCGyu2jDmNAVqIKjwRfHfGwO8JJC1SCXY755myBawKKI6IU
f51m0vUdYd9yeBJI/pDgK+Ux4gcnYwelaBayjlnYxGuKGmEgJmdKjeLLtkAqBrPC
gfjpI14iA03MOAcAbImPrBMW2eTtDI9SnH6UFUo1IaSFm7ba1szJB7M+ghiocndI
Jwdqkz37LhjDpDscIuAlGGfCHjbU3IIdcTegPI1ifTBDBJ9dBPa53cd90+wqNbc5
Qp+Lu5GTF7PEM5TALG3A7/G9nQxJD7VN4/276a+epXesKp7e6M0ZENXQefnrs1Mi
i7P0Auu4E8B+6SI09rxzyiW+DjMlblH6sLiM1Tz0XlGTYsj51hgZkIXrGkjLr7eB
NRirO5xSjOvWZ/94oApu/zqoxwRU1N/Q9gHAoJKvV2ZXyZ8Ujnod+MPBI+pDX0dZ
CsvPj4NBv2MQTYLMGYUtkIO2qCSVmhVfM25XE6zpduMaUJZxLbaxhnRd2VJ9KC/R
zR9YQ+U+qopXSei8y/kD4VA6ZPRhYgd34auSXxb3nrDDzP/8jczoCKAPxq4ujQiU
1lrvFrB3Tj8BgjW2V9yAkpBMf2Z151/uY4uJNVgJsoIAJIC8ueFarpt0ByMGrLHX
JovyUxZzWuzdAtzlCzCq/88w+x8hbAqFVYsxT4aSR+nhNpVeFPdW8RRD2X8yBuYz
o0g7VNjxYcIBVwe9I6+BSLlw/Z3OLFutNvzeWw7Teeg6XIZoWZEoHbs78CDLwPTY
3nPDtyICJkhN6aEbwqCRlJCyXEb/p1t5njsCuny69QkeP12ePlnhVty+EAUud4pY
5pMTq7zp7+Obj0Fr2Y4ALAciSJoT3FPq49tx9b8QiZLr1BWa3f0D4bdB8kBMz1+m
1ph6C6PeT0Z7a5gFeRe67xZ4Rfgz7MtqdvDtPPo6w4mgaYFvr78aGmi5R7uvUMa+
BWWyrzb0h3fw3cuVPs3RSNe4xxu8QFzaBH5iuAjhpRHlIniX/4tfswkgnQ9ySLOp
NEvviDRMAgWA14J4+9qSqf5H89+e9PTqSov7iowLf1oXtUqRei4e5OerNJCheMU1
VHZwbNvE2lAenlYe/+X/VqUySMGFyb9xafUthIUjdTPHkWicDX8quOfpennMX64U
+YPsg8Z6P/+ij/bLJJqII6MpnBmDV1ALMP0N/UdBF7ffDrCu6ievajvEHwKBEiKQ
ok38l0Ka187P2+Up/p/voaiVzFril0Y5b81OF+qSe5HEmifd6FUNwvO8L5K6R2BF
PoDqd2WnfBq79EqzlD1mz9jI3GDT1UE1MJkJT2MtQl0iFAQel0CeHJMG+KFZBsl1
gLXHXU+WU6AHpcbU8GABOHtLubivn8Hw/bk1WE8EN+cvQDd3dAe8iYefKCYd47Js
zUBJ3T6Ho51EImyCnAvokScYY3RORjUPVcCxueNL7iVX8fPWAlqdpCkTU9Fq7FA5
QpLQju9T/QjaAUHZaL4GhgImSLC3wR/lvyBRJpYGHMAN+zspqaLSrvXT8sWlm9K0
pdKzf6a+mYP5efoRWPXd7Q3TiN/kmbIoZ/TGNtHlunQ2Mvk2PA+nF6nWOIwl9sp+
wSBdmzgRwLaUOrmc0NkmlL2eHQrBrYBZ9hzFD6h/V9IpUcdObgdABIkczM6CPdEo
nblPKKw/O35fJfsQPRIkwOntrT5KvRzuKecInE7XwRaOtw19htjp00jFcTBaB98o
dhJQ3B+t4oGq36qsPlz5w981fREzsUU2u7CB7gOxvbSIttkMGIvmgzscfETWph+S
qVGMDfgK+Rr+mT7n86foGfccLp//8IHRFU2lmoY41qbJXxoL03RLhoV9HbqlC/bJ
8nHrj+DN9TnnzlPDDVSXgKvSugbphM6AyZjGY+o/1KSx8ZRs2jd96XCI6UBoqCuy
5sJ//suMOBYcNRa26ZYQV+iXc26E7kbLpYA3XDwYaQLhyKsLMG2Da7HP2obHi/qb
kdPprJauxgEkgotJSqBlkdODzuCd6uccasggv2V16Ne8v/NVmrseTWSnVqViPKuI
nrR0qifIrSFo9he0hlbJCxfPNn6ASFVhToyaKSrBZdvYmC7tA0UIJ8e0x6SiyQTf
vF14w3En9xfkSDPe9LXbMw/mspF8E6uyal2xFAug6cGvm1ewWM6eHAgeaCfxVgYV
9cBXHCsz+gbt4UrfgcgxoMkNjEdI9TtjDwVh9zaSKq0vAXtPPNFehDxG2bKBOXZM
UNBAHX2KvyhZe7f0goz7KL6W44Z8UcJBk/DvsoNymcjFQrwjqKH6J/PDWpZh2eDn
XfUPPkZJDDUl52tpDcFnaKwxiQ80mI7oS3Sc+TgrbQq1BfVSv6MsjRX0JRoe7mwi
TKQJruFdvl92wbzh+2whdVq3WYsbqlvosh8LEFaB3m2M+Tw1hZf/j2fYyPcgeWjM
AHixTrFrOjbaCCiZFRgvJpAIxzsAGMVYbcEZ6fwEWi5bGPKeLPXt3g2q3Meu7ZdO
XKe7Khri2n9tbIpdaFjVGNLBD340PL3TxNWQPPupTJIEKPDLOxPMa2x9KI6BsMH2
GrCyVVnSCIu4TZ1fILxXUv5oKPenpf43CAGRNyKMZbK4q1M9Ma3v/fqrYyD2ja8k
a2XyxjPv+4buLcqwm9mOJD4OqTmiuK6hUOcWz1wPrZSM31ODr263xKiDT+tUkATt
3BDwEQNMgmrm+fmXHzJ44w3A22QgJlC2pnGK3N735uwEk25vH1+7xPUT7wM1Bbru
EM/kehMaVZ/LCWpnf/KE0iN2rlouXABxwfVYyixw+dCQ76aktyc5rOnP/OqS7ky/
GNe3puQKkShBKT6twyMjU1cMLPFjpPYs3LZyGvCd+kF3nGABjRSYBzmIhOCB8X+z
/GeHCdqJNgH0ZsW5STLbDucwpEhYzW9T32QHEkvtAlJBBCc60WDpIjLQTen8UCKw
SmG4UMXXNMO0W3VuAezjSYU5ydGEImu07KBuyQ96FjaGGS4u1iBabQVTMVhiBTAh
iDB75CTZZmP9HDnQ03VxErQ8Dfw0qjbUkDcLM+cbT0C7nWoCLlPuxhJgxBjRr276
ADnIEWFMHrsHPqKOfvBOB3A+v/V2M6F/Mi79L9KTbq/XTz3LdaUV+tKltjOnCS/+
zUvXIKGTE1jOMnVkUur5yhwdu8AioHZ3CfpUCmWCYYJyffOndHSXQxjnsonXtAy2
f5MydXeAuioUZ6XolQxcqQzkhXL1MtfqNi5flSXG5G2nerc1DaJ2EZTRuNDG5XJ/
/s4whygO662XD3/x9eum3li+wBGEoIerWwAxJG1roqSwreGVDE4dlXAkJczEFQS0
/CyjitcB1sOHvHam16CMFp/p4n/vKcWICpTucVkKourzAZIEMhcBYmXvcTrO6C8b
MmIw1IueLm2lPzwTOaJkj48XxS4SF5bwBIo20svr5jzmkKnIlatnZYOomPg7mJaA
4x7lecj/IzjHtQEI+vfeFjJryXcCFGb2SOCUAjzNbbMY/ZWYbjzbBLyucHi2gOfc
hk4lC54DLrfVG2v8vjMp5Vb8LwtIkoS9uEDw3WONp/zkGuaSjMVfGzwRZzNYTs0r
/uYPs8ARAnLgATXwqy0Yoxw68/i0LDqKfn8xxj+IsfEsPHa1O7WlaSUC4/2l3kF0
vlDz2wm6FJzJo0bK43C8Yz/6SZZsVfW/KE6mdBO7PF8GQlWroP6DinO88LpXyhk6
quNmttE/s8xCwu6wqlp1wr7koIYHJXw2td2yqV783VqnN70dyodnTwX4OiSEFup5
9hbw31LfXYof7PxuTZSwYWLHyWm5Lh3g9GzWUFAXToJ3jJW9zVb6omKGd/zoAaS2
d++u2/IbkX085i4n7rzL035Pzz4Iga7QoF8hXgHTSr4bBH8r892wVA5a23bHBFM9
8XxquxtaKqDQ7Kz3rMUkgMk+v012e/egnxVP1gRFKcdQEQ6wAHE1p1y6Ny3Jj2dH
Zi8NnWEXOG9V9jsRo05vBDqRBru69UjKzLxeaefgjs80xpWPLZWCn+lgE7ClcmkY
hAHK7D25ABxMf81qLf60s+UNsL0xlJdfSxRMemV6uVrS+htsdBEt8WExkvyIqwuB
T4ZyMkpEdmKkGzzfkJlM4oDfaOEYzUGpJekJdMaQwl1wGnbg/HdIrvdTB/DilUPZ
zyd3YsQs8g7TayhRoTPDgxF/D8Ks1deFOh5rDUS53dnCOMejbYOoXB2s0VDc/ZMN
77OCefdWIdcQp1a5bgbudZmYDAnHmhs8sx+ynH3R+n34+YQXg5Kuhw837v+cLt/J
2fKCGulIVOmWWr/2h1CASzHSbRBmcBnlHDpPbe5V0ZfGFvePe/PA2X8XOwlyWZlQ
xRysDu7CDa0oZkG1vpZYqP+aSd8bIqedEBa7LzbjpKd3TjTuXEelq//BpzCZcGay
L8AMGgDFbKBWSnreqIZd8FPVcC9bOAlVAK4AWAkyS4KWpsNuMYurVkQDpJ9lixRq
+L9v9OTMi5Nq7CF7yCs5+bEj0MLO9Q7ZGL133FXNsAL7PcA0A/t12is4bTh3yDpw
LHZ7FMmjB6dvK6LXeqUWGJI6hGkhunbXgHYR96DlaGUhsrmG4CXXmghqJxObtElf
1IIjhjsY+/esO7KcD6e/TvOb5JdKqPjVTi62nfEc0ePEJCPH1hB7PCDVzXnD6o/Q
V9scwS6TS4LzCO1He7c1TOu+DlU7o+y5I+LG8AwSqNNHF6DNSOQYxkzp4KxQRZY6
0yn7quqGyF9wyZ32tmOPhMeaddLrJMAJ3gzYG0I0RfJQua47GlxcaYy8k8V8jiIH
ED0vEwM4Yy+6Ih39suLCVmVhiWoBP/RI+rghHlK36xxTYRMLGQVS6eByBTeuZ+H7
hEJY+j317ras09b+lBFD5kaNy0jzNZ2uKjm6RI7AqRK4qiAk3vvJj+VOL/20XRW6
DsIyKGjqUp/wfQd2xNzWWD3zI4sRdSzrLj7ZdZU8LDAKNClwJPhG8U0Pf+WNHUP/
LrSQt5GlT6ncVNKR9zNsZZItKZrg1vvfIaJ0FpnUgJYSbCi/OB8c5+AbJMJv6fIo
6DORP8BJHg1IKxHnowr6Xe9OFSDy0nSqemvj6J5qQbRrWhCv3/ZPeX5GT7J34HQ1
7SFwS3uEtucpYoV5xO31VWiDx1L6Gey4EmaT02akNSGHVgX4JyVA6Ig5qMtn4hpi
ilr+4gHaqICtadXejXcGUGazYvzLFcCrd2CbQ6lc3GI86KCWD5bunY/7sCaJz+R+
PSGlYYY3wiH4gpJ+Dotq5tIFLTiincyMC2kxjqPEgcPU4sbcMcKMbYXxyS+YzyZB
ZFBH9rE/ht2J2ZFwBHglQ+Vrea38BeN9/TF0CHuRUaQW2YbIWKbWcfD3zHgAksgM
D0Dk5A57ZZAdq8WbqBVTF6aJ5R+YVwPFzCix1Q5ocWmg+2s9lXLoeXheaYFXzGyf
1DLDeZKCgIAZGNykGg5RBrLWce8/N9yV73UGd2I4ZpL7kRxvpnsyuTeVK2iW5iH6
JrhvXEAG3c9b0RspalHhNG3iYUK91u6RZVe1HJqmCmrMZWOebnOmtIvJ7bmvDUEC
aqM3k3avRH+J7FTw+sHN/KCH4HC+qWmaJOvPzL7NiVX1giCesJnHepeOsnsf0WKA
RgrYL0ejZtwyzJENMspAmuz2+/PTEmhn7AvAYux13f8Oan3KfqPh25Pr/KZgdY07
7qdBPHfPwAZ25xyWjJRHPNT9F5UP1aG+ZutiCjGIiD2XVmubdblGsNc/Nw5q9hBl
XUgioLHFjtsCtXLPF7YiAZ8Grp2ntlbRaME+SXc7d0OHZP8cBV6NiQnX+mstWzrw
a+/OK+SXcoWhtMQU83oGoMx85rZW8fcLsDoZuNG9ng3ty5OhEQIvZ5KZVgTv99Ba
bivK2qlygFtsMuwCh9Ylzt3YaCAou/PHDRZnOMrx9XFK/oCZL7H0fLaMd6WcmMkV
JEjO3nkmcoQNTcYILIcSbecVgLh5PwOJb0v2LWpQG6hd1i89uXVunAp8WinJRZng
PSCjiT3F5KRjcfZA+NLiw9FoPmtk8IVVw1KcymCI2QvM4B6ZA+BFMFcRr8OozqjY
BHMLwJovz7QKBUVp4MmVh+a9h6DILCKC05+HldaZQfjCfunGXhveahE5p5ijbaLD
JkpG5zokQ9uJqSfH+6QoapXJtxvCvghvFiwUNkqzZawBXrwRUI6ttZ/MLWKz1BW3
tjmedD1iaC6gbVNsu4OWULJTzy0F8408VtyL9RtdsaIsSkcidCXcPwhZjgrPNgSU
yQ7G3xZ/iBfJsAkdtjP37m8UgJLElVo2xZGySE9ag61uW+5dtv6S/CQR+LMDJjSW
Z3Kdy7BOcqdBLLYdH/T9scGYmhaHRNvTlL5VJyIIhqAFby3lv37cJEbz05VxWyD3
siiOKJ6PeP7a810zp2P/mqUWM2RDQbyhnWsAlqa1kMv2cXXTb8QtmWlGg7m0pP2I
OGJVd+wXSJDYkxQ61eFgRiyz+BSdwlLsIh8jeBcW2ZDcrb4ph/4ivb/xRDP1bvDC
73N1cCYxmx+bcTVe/Xnu/AzqS6zpXtJf43XiV/7FRoChs6CuUI8eAu6v+Zl7Aq+L
vH5oFidJIWBeycI8liXqbghOv6XdDUEtmyO5NBMHmrrtriLbww4OeF2FWk5tEVc1
LG++99Lb82sh5Qd3J/ZExWiWiO44Ohp9PMdaR8KeyeHqEeuMVQ4SF1wFsq3d1WZn
l/Vu4hOUClxOZMhl+mlsbuNo12nXUYzITITUUxeW94MJKtDRjC2U1YwGGlFBjqiJ
RXqXv7oce9YFW7+Ld5J6ec+t4Pz6yAURtycO2/rhQrdgFN0Uo13aXICdMcnhYN6z
HaxpCfGU/MrEJ2plApTBDeb4QhKsQ+xr6bjgaICT+oQsLQs16mksWfvMV6Sg12b+
bh7j4JcdxZ8Jz2B/n2qdNBSSDf9W0TjzYGbfECH2S+/yrgteACB/KwY5mRdVMgi+
CIRO81nWRlweXhLu9nCjmKblxaiJU1PACG1lkpcjtiYFM2wF0hT211GZtF65J4pI
C6MAwV9aB4ZZZmFHKJ9/fqMB5C33HKb4OwIbBNxLVgUhUtBRXyhi/n1vF695nfcH
Oi5SCK5O0mejIMtOy0RExtGOUSjK4wgDo30etolw9rXIxWQslEqe7AOqZx0IKHzq
EZCauy39g+d0FKqqdRGSSdqNEVKSmvImjTYZUuDP0JZGXL8O0tiuAA0BALHnGSjc
eM+/orcyCWQIz9zXwKPJukRxwqHsBvL569TMK4CXAaouC5s9C7r0K8xsv1BqQLig
GAr438Ibyr0M5+wHU+VHLFh1RvUGwaaQbZhMBqQadXLIBlX5BUJbNul5oAqAhCWr
POjeKtLC1kVVIBkgo+nVF4R08PtnLT+JStRVj3IgL0F1LQA7Demtwp4R92ZWNouX
/MWxYRFTze3j9+bA+NyVwlkAlu/OcO1egpjgQ++nbWifawDZg0ld+CtlUSdIDwkH
TAvUILz0UAOU5dXZxb/JKUHf32X92orp9QMyy92gp6QV6OgBaGSqX4NCM/4VQsla
bQVzmvM3bFwUYco8d9szK8awPhxABx/1Dl/2ex6LynZ21AOo7bAwJp0vYwUL7BKd
K/6pl5qo16O5PpZhMf7/BqvLrj4tSosOcQ0UMwYDwP6dx/Bbg9z6gElTErV//OaL
6hzHvG0rBQGCSQDZQ8XZAmGx83g8FsUx9rBZSrsJDgvlE5OuIjKT6EGYJ70ZxUjH
T3XEoyiMzeJuPDngTRVOQhAsyf6yu2YvXI9UJiCikYSk//ezsHK79azYmvNsdqHq
HcAOp/d9YFNbRBJ22dw+6dyehTlwKU768h8nj4DnzOWOMzxkwuwkXhjnbUHKBQye
SAY7zXN/NJQ/63pAPQ9lAROSDfs94grtO4JN0QS7OhpuuEd3n01PZTiU3yWQbvRE
C2C7O8T+GBYBAFl6/cTB6x29dF9YDFTR+TFH3fOv4w7CyS3sF4c44zFj2Eg3ZKK8
ul7MxEGEhgqfMdCfKYb4pSF9rw2hWC+HSMESihVYMOGJMpIuCHphQllye7tGzyp3
AuNLWbqKqVRnCP6JSBESeyyniFWIf+llJaJWKY7MzN/7EmU458il/JnkSfa2mLte
tUIIpiKddCjrGHmm9cozvWKw+VcbVv4btoYifTvh1ADAgYaigy3zQ4C640wiLGNc
FCMgf9WjtijGJ7fEAKDLjDT04z0arSCLviRY/8oBATmZSKXJ9miLcmIJfi/g8Wbf
PeX16yMiXf/7+sLrI0pQOKZn817CboPVAs3BXKZYskjBbdbYrPCJEwfgrQneAKvX
pFmz5ffQYt6AXzLvxzEum65oazm6S2PU/b5exj6N/4i20b6yOcBiORfOS4zzjvD9
8c0ix41pyt5OzorEFWtd74OPKDf9MyAXa/IBygnoRok24oQDWJdS4C7XTJuXIWFu
Xpp6OxXoplA1FJItzgv5oWLssj9I8ggRwJ0d744Wu5M2X/2NUEPerCbQS1OJfO3m
w8oyp3zZYorsYAMm4s8KYjjJNuYVSo+ZtnS7kzh6xwRmhu04ti/tTrRmJigKlV8L
WLLzD6WuUnOeQbVbfXXaa9a/QW1ctFw5ySV6cJY/YVs6XOcJAOPIvpGVQj0je46r
DixGHMQ+DwlIbRhlL4ObwNWXvEZIA0pvA2abYhoVVLDX1vtR2HaXXTMb1ipIrilE
oraMoL2rKv+FhKaulhY1UAZ51JLmijNUtTqZsfcl/cqOypiuVtXTL2CUyO8luZPt
ITBRhQhc9scCUd9x2kITHIuuL9E5WLtuVC8vl1B9QS12oGs2lnDawuO2/6uCbCL/
zx81GHVzgf9pLAABCtMkJhgT3BDpT/Kjs1rpsqasaswsV8JtFnMiVDf3ksoZRLCr
kGoSbD7LRlhm9RawXsnF858HdUV11ndcOn7Xaq5sDOlsN+jHdD39uH2ee3rPjU0K
cPsHCjr6R9UAukBP0Ml7/quIca8iYn1CMvLpDO3RLS1YRO870asYtSwXTftZykwH
WoRxrJ2PyTlIF7NlRKjs5msSjLATIjsmdb0D74XAwjpyKXdBtJXg/LUq+uXbD+ZC
qGo5oi8xO0lQegcoIYROYAXZwsyNTGupWLukYQGLe1gufL13YmWjUfK0HjvU+uE6
W/CDUmnkJT3ne+SRqIpqW8mdYurcEYuXZg+rJQY4x93oZPskZ6QwaX5gJLgWOrmF
FdKgIGw3iqJ9ZRch39pvuzaI1Ghc4PkC+HvFTh6gIGv5+lf7oy/Y23C/uTJP2+Vh
wcp3YYOesjTnScl1K7mKxiKIUxRszRQC8n0C9J9NsKkp73730P6B5LUJePxREGIg
+muZWt0EX3PXzEavlznHd+aDZbFCLhhIFDZ/Hba4SNnA7OPS2WH5hgBwPJNU5vvX
SmrHc2L+UUw9XtvwMgGtgEOZZG4z5QR/tssybe+Yi/+PgTfgiupCNwHU09qDY1wS
srCjh0dEeUUwUMPOLRs0BAr1IkzJOQxSgX27donWwvHUc3/FkI5r8y6UVphKKiO/
T5zf7GpUSmBNTTCIyZ8jqalAyERMPwNj36XXCcFBDDO1JhWnMMrLjvdYrKLTCCx2
9sEDPQL9hUGFBJjIPkn6iP6noWqyUEhAbQSOFOJFpIkaA5ffh3D9JcT01pUsRfb+
b41UsQ9Y6zXlpIUL1ypUHbLj0neNB64mjjZkPKIs2KTMWvKdXNpwdGcsTjKLbKav
qLxm+/dbU0NiunKrdr+afkLNN3/7AYROimANLeRbjLochvMq5xOQcvySTAvi7GfG
UsnmBEuy7VEnaxBclLB/gfslFtiwR2hhhLLJmNtB6/9E+Oc71RGBxi2VFN9xF6UZ
jOqsiAefo/YPG+Xl/9iOhOKOhaUBdvKnLGYbTEI/xgmAKUcAwPQ2lB9KcUHHjhnz
AEyjtevDw4QdJje+tfWEip4iRQiKm2aV8ahJ1Y3sun09bvl7eZXsinVuDbZEEVXK
LiWV95I0HHPPmlhlQZKUYGaAjXxYaQw7a/5bXivS6ErXsFkrHmvI67/VdB+Z5a54
8TnYzLrn8Mbm/84mRMtd7FlTkCyH2PfrZPVEKyqaWFV4UNnEUpycmJvN9kYBxwva
Ou1ZIeryzgISIkrOTOqjBdtIM/cJe8+Zsa0eWRjQg0K2q5Bfd3uOoEZd7yuDSRGL
xnqYc7cP0VOT5Ab8tFhhl9VIMMNNylAzDALPT19lMSXPGEV9Kw+oaR2LFjGFrAuE
jKZiZs8smunnpMGt6uBTpXPDk6K3v+vhl1dWZ05R2pytM0rRphKkncpKtYDHpfFm
XalsGYia2PDtRJO9bAkFKZ/RwhDsl8IEwYgKLReonmuXbzS46Z2qCb3XwVaO7RNY
FM1xiCebQugH6Kl3yk41MhHEpUVA3ITeZjbrE1mDyJtUr32Cxg6RFeOlHYQtRwTk
34pIpOWBYzlnwW4A8/+2gNSC6tjTT6c8igG41pUHK+EJEmCyLZwBvGo0bAe72vGn
ZE/Yib+MXBA5H+wYfz6f7P5kPREjnFx5PaHXmSG6vjT5uYPBEIBn0KDBK+E8clf3
9WAdMlOvzkOScs3/3A9aX6QDVaBIaKIBPKH8h4vkmjonDN7x4mmKceWdn1HVvE11
iZn3f4nwclxw9hgxQLUDz2QsT9pavqA5jNxlZXXeCMCLv9VDpJ4vJgY8IsP5fAIA
T2T3IfOoBY1dxoKnb8MNJOr65ALUOlKsIw48KTIVoLNjOjbIfgVDPKo418JDHpYH
SClyPMX5nhlmJBWjc73FQSDcSkuTWNwhwyzu0HC6SMKngPrnmxcL9ESTvBPkTwgy
3dRxZEJxyyCTH7DO36IOmGeFcAobu6d09ruM3rN3A9XEBzUEHXGElsggZdiV+kud
8wpaQee4JETIMFEWKhesRpQW9C8D13nRIHo/qEkILefq1KKzasm7fgvACd4ukkTR
g7nBpDfJagbOuD9+CDRei1kSyf3gJCJjA5HXlm62nuN2e+N8xizXJppzfRQI3r3B
10K1ubXvQ9D4MPlLBjz5tAHo8DFhZWkRjVpD+/NcAb2Ul/Jh5Yxh3wS3YRk9UGKl
E7hTOugrs4rTBwwXm1WgzRj7D+icJZNULnlpFxCxqOZSn72HAgPPEPVTXml4islg
CxZ1RdjMFTkNlLX3KPxOYrYkOQnswFpoK/8ADTgOC6lgxI7L03zAcVMgr6Z7rKYK
x7AvHEX0cP5h6MDBvactU5fhWXlaSxpcY+ZpMH7HCO0JKrSbE3P9OEC7A7FCoykp
iVSjLGy8LFmi8k5ENtAE6XEQZdQiEXkx0Nn8hU7zqQgeJsQDaJpFgI14Em47qENW
OdBWfpUMemT48tfbQu269XoiSg5oSemIZhuu1oLm3wRsqIZQXMA4WkUYMeo5XNha
GudfgU0dwvfaQfdE81WUe+oqoEZcDmGIJDm2zohNGs6MhMROYByCe6JUDiDEE3UV
Dwj9dsFEcfl3HJDyayP2hY0D3uki6QLhaXV3S7mCs9ekpoyhEyHRQoAiHfo99UYM
sNQ3HGdy0bIlXPj1WiySTiCy2su/Ntl6LofUQwE4AuUY5p4/a5OFYw3bBrfb8PXW
iL2rlNusi0foDf43nTyfwvs3AhcatiUBabQ+Irj8lf3r8QZtkU68LIAFgRO9b9U2
MmHTO1kpDIC1mqwDcDKQ3yWa4J7r30uJEZGTU/jtKemzVeubnzqG2gALxZzPtvUU
u8dBAhUUipnS0eYXU8tzEfoIREn6Zj67QKxgxJe6FHtTCMA/MbGU5cIkVdrIyJFJ
AdMq00LiijLcmdOHgijswWsDIJor6FRN8aLb3wT6czyzU6+F/EbmcmalW96VO7Hu
5sESP4iM0vUiVrhXQJ2fnmj9N9qILTQY7PJo0SxRhEOzR9qsbneCKUjTJt8SbHkE
aND+Vt26A9msJ/THoed+D7kgPrHusIEegmnNCUzoVmCbSZn35a0P22BaL4+AmxSm
9usnmvz+R60pbbWE6K4i1hMndXc9BRbK3/yqRxxjir7c581TciojgK8xrUkO5TPQ
VAXvpS95UsuelhhZ3KAU7/9+fdxa4F92A0eY1h6xRdIpAR68ss+OGwtSx6y+OHSe
fnbDvNYDXRlNH6dVvePbFnhl5uTHjsH3xaQB6Z58Nl/9qiQHX9FNJe8ZtCP/atmU
kTO7V+UthIKBOddY3TppBqs0L5yvxGuWxuvqdaL42Z0HFui7Y/Nwncu9FPW2rPCI
wGugiUTUfQwD1AyBAsy4uIBd69abpJ/z6sfyYliSqOQXx4cpGkpGuaKN/FL3nmmo
tIrid5lBVprDLwgUULI2xo/jWgBSOSnIXBMkCauYVbsQxFpGTHEcx6Dn3m3nVG7L
S2tEtCGFIlcZ/VzhG3NcgJrIqv1OhrNibateiDc0nqFp1GHbWhE4wIrAWbWIV+UH
PXERiZT2dvztueJTCEdKwMYFlot80nhC7k+l6th2sPTVx/2dbdfxJ7DXSFyxTngo
rZ7kaJcG0skHcCa1vU/6sMrtzOm2TH9c9xz+2mYU2gqoLr3njQLW4So8HHvRvjA6
fdIMyRcJXWZNzQSmf8I1gzMR7X9AsTfiVmw+RxY3jlW5PM02KKkSoLyM4aj+N/d2
NiwVRe6WIpo8oIcAYRt0ZcNEzwg6D/F/DiaBpS2m1HhfKkvb/k4fTJfACyhaOv7y
AdNLRf7D2N7BB9OY+yWD59DjrKzH37soT2AdTlcFRCp6p88ghacwTYSCR70t7nGh
MBUY9fp2RMCj/18TTbY6jVbF9Qcky6qdGSc6SW4UyQRIad4BUDhsPTdLWn0Wqclj
uG0K4YG0LDPrbN/CzZ0/FHLO2JkcZMlmm0codwEmeGESiQWKCogWtpC7zikxb1Cv
jRTUD81UnRO3snoz6KHPHCuI8WE7Igmq3kKf3oJE0pnCEjYjkr75Eoi3mdTSJhVG
aQtCVJizsuaQ2UKLeUxncWU/gr2hsLUTAPH1tRCc6+GKi3OjdHZ/pwjalXiG4D13
68+BlpwIutJHJp7kVteNVWmdcbW25OXBvUpEt8JmU3Ynag3TOEKljemhV4y2zBw4
csQge1Vn8w1YIGLt4sU+/j9RzlOOMIp29UDJ7xwxzviFVZucpk0qu1MnHcyU9yRU
yO1CMLinOSI0zliGvAHaGmvjXsexbYTBFXe5ZEwNSELFV94HbGWAKs9iXRHJhyp4
QvX+D5/X2jj5Al1tEOKUU+37uCCk50TmdaxRprV1DlcMruwy8ono8RtQAav+q94q
ojjQsWxORdbrzaNsnB9TSXkDA/r/u3ztzEmBUGqpqSCQjsQVQ1eiqToxLTscgXHQ
VWTjlPA+fsHUT34ZG4s2nUh64ZobDAqc/+Jpg6/QoFm07vyiJ2ppYUgME1j4eufR
HQsR9fIkcMu04PLymQQCGIxm6fUYAaBBq2DOSkIUd/BscKF0Yn8RZdAc015xiMoT
bZS/WiY4Ui/gA41QWsTaiIdwKpPe5HbQO2agSjd8dFOY3wfQjvoqpCu0yoo9mCIG
dhNfNkv+4VCVrFiat7HcSdGA6dfKzMt3IFvkqSBXvwmy+q1sYBlOjB5r8BPWGJMy
aZahzQo6FfMrV+1oAy6fY5HFiz6SIfPXkCLNgQWja3W0MCeb8dekWkORnEa5oK05
0vPAwA3cr0YgiT4W8DaQ+ntHpkGQ4rBBUMMKlSyocBkj8Or9aDp4UhDS2fuV89ax
37/WnAi2TbRfKa22CrBBiqBD0EZfcdXNZiSwmS+KOOqbWS3Zba1SFzumggEwC2Ef
G0CIfGoDFXsW2XtkOTNVIvjiP/X83OoXy9kyZkQ4N6fijJZbgQUZ3vI23eYLiuQe
dc2MxN7yOQFZOPujorkuYYplLvbjHgtaWArm+O9w54yHYqN6VDv1VPbvcPrle9Q3
YAYicNxDdbj7x4PLUIRW4Cf5V4CQh0BO/IhALKcK09x3h1zrA6rM03rQtwpwaLkL
uvFp0fC88sVEA6XrOT+LQzL+FbqR8909xxKwASy6zbLEs8Rx65QJ03l0JRbfN4Tu
KYwyyx+ApSieVvlgsv+BJVT+RW6cFjNVkLvBwnTOdsf/1B1pft+qsSfFloq2+1fL
WMk7qCWMVdrjEhE7fnQuIDeUy1FE8EaQMDO164yZRtE8oHt8+/GzzE6+Ch4EvZS8
I96ln278gkpYEeO8rDZYKWCvo8OGhHvPrdQN23L9uRYb9OtKd6y/0/AXsHOUWkm/
b7s7/iQcE//L4Z8r0YBF2axm2FSHJ3rydC8WhMGIDgANOxO2Hp2XxQ5doG2BFJC7
VjK82pQ/kYNGuQF+Y5y+5ALBqrulMEeHBJPnLTj0kTnk+rZgz8wxlRUZbq6sZLsh
ynCHoivcP0DNaFuJCVqFj+jE6xVK4cqy27a1jijsrhZgv+nFK1IMC+BLWQAXPLpW
cy8gjd19Wr1PMNqIueXYvqkaC0djE5PXO93ReXrRf0/F5z3UAe7eWUxgGor4QaUe
C/FG3OLhb/xD2DThMYzMFW5BaXbAK86EHlQzbkNHoJriPiK3TtefyQ4yc9UB/Qp8
LH9t0MSbeLm2o8vBe4tGgdiEBB7UNvI93HJ4Z2xCziRQ5KZ8eEN/UyWuWjLsO1fy
xjrwf26slnSl5yP2jgxFnYsfonIzu0NXhQQ4KsByUz/2NskBPTA92k6Ob3q4QEac
NBnG5FpR/TtNJV1+POrdWCG+UNnI8DiVzCN/CEB+6oBZ+EuwkAayhdao2q0njFFO
pZmsjPOKP7L8C2X26fuOXBqKvEce4BrC1wze/U7iakq2ijOGFrETTB49GQcVZqUl
JIyNVtorZzpf2GWo56pgfpNwvQNkcbaYwiXCUNkQqweeCtmF15b/YxF5fHcrRD7C
AnnxvZznSo0HMu/QjCJmasLLyrKjuyU02XyKp4jV6ZZIl7arpYiMAb5bh/w1USTK
pX0xTSlgERYgf6lGztl6jwdEPq/75lswmQV1W/eL5q6KhG8NwEeT0bxKMrytGGo/
5/I57wbACEPDQS0/MEjemY88XgD4X7E0DFTnyb6pquYYndHRMqiDFQxVaPEeXnZR
fI4E/vRGox6KPjhG1WI/HO3dvCasjnsMQ8tDVur8RqPLvoYa+EJSfHVZqcayAf17
IOfZk0HMuGatBJqe51KNoN+lsVEVtYDz3D4Uly3DTd4/vG8on0F4Enh9QTFhh7SQ
sr3d9JNWbYmvLMgANlrbwz3dVFiZK2CegGxUg6uh6lKtC5vRIDB8XniGa6KFGu4+
wugbXVyAfiaa+rrnJxZ9p8AF3+eLiI1wHUoieEEJC4OSk6WiLgsYF+rfM541UIv3
vh/+4FmANgdeBINa9AxEsqJoxILsSfxJWvDQvEj9eynBZoCMxM2GTzPYRUBJmlPB
AsP2k5xVwhR37KsPT/sGtsE172YTnVXFPVg9Jsm5+K6NI3EYvQZoqdvjNwL1nZjB
gWNJglGC8iS0xtq1TeoCAIDMtIclgDnEJmxEnPOYLhR0gq1HJphh06vw36Nq618M
teXWQtgeL24fGH+73hVB+PLrweHcxNDHVrNIMNNBojCEFLjb2MGeTJ6OVy3IXfNi
Le+sbsZG2r2/gwWeJyxLECNfewMMevYCqcjjg7B62PtYh/GuWkX+PU6Cedw1m/lG
b23zzLlEyEbDoR7dzA55UeRuHephKyLztqWiRaOTTx7SYYMgss5FCveMFmdNJ+sx
pu5fMYEmhj60q9jZh+o9I9v4CkUkEFU2gOJhpfG4RRyN3tZIYN3SHy1oo1tZKZC4
7ZzQz3onpxSIicXfNyXzws6Q075weXM1iOjWAQ8CHrUE0eXoexnPJlJKn3P5guco
5zI/qJy2njOzBYtXEP4bdJmpXkAzj3p6s6UW3e2zAi053ufHuVg1zkOmVwpJk46/
Q3aZ3DgnFQXNrI4ggVDOzt7zuoRDA8tn3M+xMB7YhhgbEv1rOeEpacx46dCE09qZ
g3aemZgezgtv0UtZDGaScPj1k/wGIGoXAA2/Kp+b8XyhIfdHddhQccypvej1g6Gw
0Jm81CVnNtJ9vNI3UCv74zlEaW5kjU9fGB/A/5umtC1yLyzvcVVLZA6KMbJkNQl3
JFO1KiCUCYVyracKBATh6o11FiHCWIEQBedsafMATltdhhVlQ+n97JqsIC+87m5e
HFGrxJY5Jb/PdIheVfzvLML3QVUZsxW1M8cZ2V0+VD81NMSzX1/qHhmc1XJZx2/f
7GA8A8kfblENxvb13paOOWGwOmNXRxkWCPYtd2b2TVR1SXKJzuT4TIp14c/Yv+QI
qtTTGogT1c5epgmYW1wBboPeRITyQ6zvAtrrrqtrBwkznu/1U/KWDQvUUDFh739a
EUS8tU3oykjy13lK0ZlxohfV/51znfIYf8BVDio0HqM68Tw6774D75VAUvUdC+2X
NAzyGMkJfxUg4q28lprLrOHaLfGn2kaiaG0adO4n7TdZQUZhp7T9duot4ZdvkW3s
cgrWa6mbk4YKAv9fGnxQEKPsR4pr3II7XWyLYISi1qTU63VdoA77QSbeqcb/S2Ye
qaCjr5VQQ4h+ztpYpZyZ303d3DRQ7vUCrPyPoni2y0WUIW5+Eq+bwLfiBGbjJJoD
cuDVo1F36naBBDQZmBts+eYZO0irGok4DXz8i4C0aJhNFC7NbuQOQa98QYAFQj+2
QgR6t3ZrXVVc6GuLDZTouor8d4EATvZXXPWLRmz5AelboB5wgWtUo9dTBiu9bPBr
FphbT88g6ZnRPbDR0uBQAOL5UPEOYy5PtoyHr1Sx5lfnRX+9+9jYeXicnM5fOTSH
/YDIzzm7d+Rzgp9tExvgaPxLE7HBSoUG9WzE0xsmA+n74GQsLpFU+Ip77DSmz/Ek
MEAdSWJQ+i4ybroIxLWEqoYW2oTe7axoNXl2QCqcMjYrYSUu8VnT9/HJduRadtwW
ErTHUFkRlW/L/pxumbPZsD/QCbraHLqg9TxGk2yE1mKlyz+qCq5IyvoFQ/+/PAvT
uh74pF4kL45VqQfCbum8p7vfv6fOm1ICp3wqB4fAdDb5d3Ikmr6a1/7XxPKWo27K
J7BZmHKXbazNL+x7jQ6KO3DE1yokh6D5MUwP1mMnUFZwpRciUgXcl+KPjaOd8TPq
wK8HF5xb0oXPA+rJmxIVbLTQw5JnEgn7MXVuUg9hTa2/aZjC1yyuuBk8GVa+YeQf
sx6POmQKwrQUJZ0l9AY8eh6pBMgYXOb0TwHwjTG+AAngOZX5R5iHn/ZOVgfdMQSK
jFY4jYdZdXkKIAfT6aDRFHjnqHcj8PUGMh954w3pExl9UDTu9BtR9jzsL61JKjsM
YSno/7ploZDd/ui3cHMeLCbwmr2XaVRnLJZEX6v6gKXH5cwm9KM4Wu8htxJU+/Yr
svNhdz9qjjPcLH2WGAtl24qjESEdRCt5z3icGvEmA9OX31Ikep9nlWtPTjXTIzhF
yWMODQ119an+sheiyUuVTfT3732h3R4vKPM8B9Jh3SeJSPDruj30lLNtJcoTKyVA
yZZYGT2Qw/3Yqz7XAMP81qrNaWCLQdni3y+kO5nqs5IJ4HAumLVd2nSoaU1R10Mc
vPNrIdZXpYSMZCea4ycMvwdujkHv7lJMP8f7kx3BRljKIuZQ1Q4caVRnDx4gl8rA
Bg8QczKEQDrzwcLNxZFUPvOLn9wmscFSkKo/P7ThssGJRoiIhaqMc9kUKvlXNtLE
sWIotU++USjafNsF6paWw0y3KkuDHxsoZycy1xUq9WcmfzIyVb95ozDToy2eeqOu
QUNBzFYt4ThAKAPIZSJNpD4Tl2UjdFxoZlSMc/5UETKCLuxWFLLX7nukpQPL8/I2
qPZaGRwNFoqDVqTeJzWZfagd0q9Amnn6mQplgEnuRvRKRZCL07q93zQ9nTfiKJMp
W+KJdGrOhAuo6ZWu8x35wdQnMUlcmVX9gKe0spmn8WRl5UvnjKAniig7is26ojXB
NEVu4DkRfZTyu6dAimglI2T+Nen/tlkiwUN0IF+00a13i17vRoorNdq5xe2U9SIK
NMW7tXTPbvlCBq4acopZVJyAcbxsNXwedBVxMsaZW9bkXoNtZIUePVO/1lYWuwr2
vJVOtUzspIkw5lT37tKpDWfBtiyPOY7b+2zHTKuKz6ODbAUZbGyyGLxbJ0xHGNbE
/e5VC2rRQhBLV/Y0BQQwTO2GLwImxq59eD3GtBlqcmBKOOhhfJxa2vmwUnUYOrx4
p7GEWp0waZKTNw8qRlh3zdT1dOk6sprfRiblWiaDgvAf7ptA2w29YN8OllzqQFCt
Arm8F8ErYRO3HFF3jtAcmf/27JyGLL3YPJOi3ITNA+m3R1Va9GJMxV0+PykeWBnp
D8gOfhsH7BpE6+klPms+oiSj1zn9viImHYDlJKAJG7+kpfZmI3lsofbx5Dx4gtZT
1PbZivZSNAmUsNALBbOSQB/vg2a4L2aVBuFH2/QmJwwyzwuN9A95hhToAjKx/Mbl
Q4iHLMT1cdwmCnUWEkqVpJfR/q3DZWyCi6WI+05Kc8c2ek5zbfOUR57BOffiK6Et
p4ZmjU1vxvtfUyvxw6v3kc/tHFJGG3o0V1VNdiiB+oywAVOnqJM2UiBymArn3aqp
EoOa78AV4t/5KuHzBbwBfK0txpDVgYu7Hn1GLNt/Y8dGvyy4HaJ0w1rF4Wi1Q35H
hwzH0dcf5oXNkU4PWVzs1TD3uuyozdjs7Rm53pPr+kuQ6aFsslo+KL7ZMvd4nYAZ
+0VfS3lfxnjvQXApUMV3zw1yi3UGNKTmvDLZIDSA7y/nGzX6NwCZk/d7dn+OYA4M
3djFQrksf1VWVH75SaTKqMq8twUVxDoKklZk3a2nNEx8KemsZHQagFO7V3fqHAP2
6Zjk/JsbCZf3C52n3LDCb9yK3Uoj2aBQhVwTdp1CczuwDNx52wTsDNtdmRVi0dpL
fOk8fFNEBTvLCf7Dzh9UzXu9aYFTZcA8LlwGuPbciCF9DjU3nOvlKzqrbya3bhkP
UBkJbgFDy474+QMHRPO16ixWb+1fr0xySxonEKRQkuiKTVVm5mg5sIfhtYD5PJcm
Cam2nvDrbyIpzk46/ilI+0TBHRjYwJ1QklII8Xg2zoa45h1+RcKaVE3eSKXuwFBK
H9PvLLlNSFCx4ywYTwwb01RrCV5zq5cRBuaj3X3Y1ieJKoLWRWhWHmCooNXG6o88
NEiu5JzbZ2bsit03s7lNlxow9E9anV+YuTHOBjW/m1/wg+FkBe3Y5ZkUOFFp6lgD
ed/VXf2XxNwQCeo7Ejk85SD1ddTwdXrUqZQNap6KUv12bbZx740A4E7s+Km4TJq2
Ax5/VZNGq9/mr0LNSHEIBzehUf2ZMu2RWczK5PcWtDkZEakzUl+GBhLz2ubKZ0NA
TExdGBOP6ME1HoQ2JBqB6Y0hkKyWwEwv1hOrx4zAqitjuKkGJ7i4bV2YyetLjsNY
CFB4dFDpiLKsEy1rWeDzGi0dZSZKlNcwP5/sg9xzhFmSVQHEMActLNRAk9De7LAF
XXYghfsHqMSPNW86u29xSbS/y8StjuUSRGkCcIq7iYV0u6CdaZWsYFxB0O8RHkyu
eS5cUET+zYAJmKa8kfrmkGcBuZACd3YQljmeTchefGYoCmohmvb99EZSw461j6Hs
4yL0lYAk9FazA9l1aumzjNpWK6mq/mQ/n0VTfm/6w49S/A5bLsCrXbt36/RZmYBn
TLw5ZH4eu01xyauSmktwLcUsiAVvHSJvwwqd+iB/a+F/O4AsMsxS74dpzPbv5RfT
d09hvYKXDJAzCuyhTPv4ZyLbuR7BnGkqRL8Vt3cSwaMi/Ef7gMCMdw2vyNW/8T9p
1qB5aZ8qFdnX12jG74eUiq47BblqqHtuyBKmNb08H5PIovmQhzSrdJgTiIj2TSJZ
J14zfIg4hHqkuDBHRHab4e7cCVaISFy6J/mb51j4oq3W/HUMqCbz+UxNMIy4FdTg
ZhoNq5n+ovvDBhlw9MBo1jMpED/5yEFBE2VVgRPHDh9nRRQuQaNkcg2xnA16oMou
zB/DdvlFrweHZLx4f0fA9RuxsHuWDoiP+kwhoVW+puY3lIsEnwdYKhLh37ZqqCCW
4Y89ZJMzSIX5d/A4VX9n1iLj2f8WUOZ/wNKvYWt/0/bTCsLyJaakxksHAMF/E7Ni
SF4HcrqHppINqPN3GEN49vwSjoU0Dqn8VOfMFp2zuydaavHkKTZbRi0aa+AYJf5q
ChFV+/eri7tMY/php01Dd3fpA+MaOIqbHwoet3VfAxub0VEkPaDZ/Qxk0wkjeml7
r9pvSDh64LIoWYOAyknFV3y5zOQUBzFpKJ6HOfCwn/2CalAOyrO3/cmIxv4kjduo
sCKATD+cqErmdj5gHEvRmtpAcK/bxsXro0OaYnOMHPuwVwSc6usiFWNkdlDg/gHF
kbA7T4q7jr5s+ikC/EeTvOnS4sX2gnJLz/wevJ80Y6QTlzahKhj7WwOYC1UBevKC
8cVUDZRgB+NON9Dgcj0JPTbwWWlGIK3IQEpqgQZ1muKCrWp/y4VNfjxo+pxkqZ/h
yNs6VGk/MIG+v8NTpSTwsTHMvcy0TE4QABvo3GqqCb9dJQ+3w6zppr+3UeWH/D9h
0aJbDqnxWwkn0bi+jyi8ZXCnQq4utPI6pBYFMN5aA2WwPIug5PdSf82bWBnxt2ef
Nizj2wOsO3by58N6a9SKNd5ZfLh343WJtzoQJVjn+UuJZRw+gVij/1kjyxiAQQC/
L905mKg7//XBfLNQUlVRXatSmwwtUa/4lyC/bVYOPDa4z4aiBan6xFlGvnp07sAl
RzUzdt6car5zblF//8N0xuKRL/XMaoK0Dpp2s0DG58UiUj8Lx20EmGTzmyrkwb57
Vkvj/eBA/O2+PnrpVM712TgJ8RH8VA4pJzaERCFX/7WYm2w6+YHw7DJc3/zKgBJI
sswUD4tmYuOL5PJgJzrvbOK/Ak0QN7eEDWbP+8jKwBUt4NDux9G3bwZdfVLphxb5
L1SIWEvISgeEuI9ONwfnUb/rFWgGG+rY4Q11aF20f9ijXTfq2Qbwnm2NxZALVQRF
1tHZr8jC1tG0+6QhcxHnx1J3Xtm18MI73jYgv/Ifjjt3x8nNvA3EjTKXUrXxdjO1
aHgVNUOQpqJOBLChaFFGd9SiflPnCPy6YZu7V4HoeoZyqT77h0GezErQyS1k7sVI
Yh7PA4pwXlcGCcnLzS+7uAcqMjdyTm3Chh1lGikFS2DO1NVUQq++au/KJoVbJAGh
Fm9CeVCA8LETSzcTHIYlZTjTzyVA71a7/uLMxZcEacbdibjJrk78TEUdwV+ZpIjG
y11SSTPHUjNqyAG3mTRCYNjt5RM1LA2JID6aPRY6pSqOcqx5ydNBHO8kZgRtW9xB
jEoowfMMqhR+n3PqgeWvREqIBrLo6fE7Uf84h+DQpur6k95bgd59ENyMuHOdl5vZ
eHr51NVE9ss+1yJtDnK68TLIY9ciWjfCDaY8dXkeFxpAvyBnVilRWbjphvLYq01a
K1MzVep0SAeD6slGLCTyRXZeRarBCfsWnSdlwhSOweYJfHha54aDRDCM0hPM8qEY
rn0Q4UI3HHzOZc4lY3JT57lfi/pXeEqhQTXz5jfIEKyH3VQ3/UjAddrjOq8Hg9L/
yei+ct2mciFrXvsrFPFEGhbr+cMDuZkrmdY34ZrW2QcrjMcA5BHt1QXj/ZUXZZwW
Bwb8u9HMNUitbHViUY0YC0AO5DC99lZY/BzlBamm/bgpbqx4nUOJ2hC0HwT15vYE
m26G0TICKd3C2gtbCcBFRfKjXTk/UqXWRPE9+jt7uaAG1mE24A2uq9QDfixKbNe9
8wxM0TnoCKF1vh4rJ7nznwnVCdzDc7WBv6HjDc6BOUdch9el/gX6KwdW5UcMJ6/9
1pyY0sn/oDDmNj8fRYJDVUbGl4rM3Yj3nDtZRH9FY3oPdYXsyx8NcvDNS/jUp0tu
kJBx/XCC0Fx0qARopBhaa3ldR35GouYl7MjcCHDm1BskouFQeJpLSAExggI5njLh
80NH3jechx7G0UhuPWYWtpgaioeBwYoN2W0X5mX2OhcZD5bZhzbPMwOE9OcykvkE
KApLDAmnmtPCkCt5Ak8lNjlmPGD8Sr7I/IXo1jQluT3e6IkeL6ZWdl7oqg7plOi4
/sZp1R075uhupJXHy5jv8a3XBkuu2kzoIABj6vVtnbH5vxdIRy5RyoJ+2yqh+zw2
J089rDqyLZ3iotNZmXZ8XbdMQJ4zJ8SAUhcbq+37SPCTUKGNcAQK5UARotWN9QUp
qBbckZfCBSm6UPSXz3sBBQnqIY3OZUiV9whXSbLyasP5U20AGd6FFxC7mcKCY+cy
kP1boZL5uas/asvMRuB5RGOLMMezngMhV8AXz286hETggzKaEoWXR8XuY8Fs6JqB
F6td6bCRC9PiQ6HQ8fs5AjedUb4iSopVfdjXk2OW3hKIjwqphymT+SURAIzQMsdM
m1Cd0+gZlGnFAfeCPA7jhFudSnqum2T2eZFTBemcEpDjGg6lboc+cJEyqxIlJdui
1YfVIipOj/R4eZPg/Xy0VHV0upPsT0/pX8nl9l0lF/+dU4dnuvq0gmrbJkQGjji8
zQoeEjjmK6yl7NnI/9FOiaDaLwePVbamkAXTgb3dhAmP2lnYvRsn5a2nS6c9DVcc
NjEv7Lk+6zhUp0kk63qe1wEX+Ye19GVtQAROunlW71Dic0F3m5tP+sUL4+F8utN7
lDsN5vUWkuyGZqC5BWNrADT2K7RzNjW8ugKISi6hZ1qCLawZst3flFMaPcXxuL2S
EIeQajMJEMZpG307OirstIt70SUT7ht54jjt9nP2t/Bxyp9xBU7Bf3OYIl3D8xXk
c2QSTtdj516kVAbjcqVXlGwXUJKMl5nkPd4L8AHjuim1BEdQDMZFzoe+LYZvqSPe
AkUuwNy7R+KZeZD2V/pCLd8Pk1O2b6tt1wVuOK8a4JJzCERmNMpypRsUR1VmwYvu
lz1vjkqkXQpcZke9xuhLw6yTMR2liCa4C29NSdw04VyNiDNeQFN8b69ckTJ5Tfoq
QzdlT58neIN80nwiDEMLEIgVqAmjLnyGhgDagATqbzf2QIvKCW8Oa5nWnQ0fHGue
uLCWerOvu4xnx7L4fR1afGqwd2OKUX8Gx8jn/91CnCfRMSUKLvcVD0sTXI0ONWFd
fJiTmmSOa976Q5wieCltpXqzRGvXOnYUXq1Ejb/RkXr5B7FQQRkq5itqVW4qK3N5
/0Xs2rJdLfIBFDtO8h9hs6cwZnU7YJNe3on9VrRWAIBapM1HBzwI/GaZv9fSmBPC
/nR776//w+UV3H8xMWtFsgQGH0jhC6kfZC8eUKtf/ebHAHdDqlUnC2jIt9LtqK+W
/jhIcgU6nMBjUTEC2uKVv3ZAMu9rk29krzcJwwM/yBD3nqEIE9vp+RiB5dh+0frf
5g5vcX01f5Pp73xTFcNPEyuxvlesWUANnsiOGhdEo8hgFIyJ2uzU9Wxh7yMQJ5xX
j12a+Bc/HhMsDkJFyUbFpvHbCle61oc+wfFfp4/4t8xnOrTJw7RYMbfUGwzy8zqp
R8RoHwLFE8ZL9lG9XajGJIcJluV+HGUTjKZ/JfdIpIWzuAwKr25GKNgmg23hX1GW
IRPLiGlDAIApXV9IjYr+b1ZGOofGlykzU8ow3Jtzgd2neBEByTZ1LOHH/IzcwyQs
whi+c+20v70zq10W7vhnjnmQi/CkVYyso/OCjdCxJC1Fzags05YAf1zAZ2UXZoS1
VwH61eQ/kIQO7GZG4vmxJvSempGxp6uZrBRxW0lIrtFvagF0IL/IWUcaSWf1vdtb
mrbBDlL+F+dE002J9YVL09Pj99hiqkfYTOnyBob8B57uz+vYwUKdx9OzUGexJ/eG
B6LOooIbKPmUmcrPC4TjNa0Di1FEMRgcaoJ/eFRCGr06F5YvPyS64cbMFwLxlUzi
u+uQLKrqIKHtiWggfx30J1Dl8KZyc0R2VmK3hiZpWTtU7Wyl9fdSJ+uOe/We8EjS
9btBxdYKxXRzwqA9F0esWJlVrysF0NARutMLfs2/OjDyIq7294BqUy3Gjj/cl9eT
YCv+TlHp7zefwqHe7qkXRdr0mvoq6KuXdKRRl5OTxB5FkpzexqFSTDB3S5xPPNxG
t+M2gAj1XvGIZBoay1t5e89W/eGrg5O1n1YJtF2GsZnUe38o5V9aw4xAAGI3Q14n
AT29akvItWSh3aHfy1Ich+CPJNsnYUpuNQa+aGaOUugvwSaQ/9cInXVc+sxOGdIk
OL87WalBpd93QuVB0NhDFlnDDcH+NbjuuhiRL//getll+x2sU5OSHpSxS6aaVCOJ
TFqi0osfG3HgBFTh0psUuy8djLUqJXEB+E30LMadVjjGrnSuWXEQXqY3G3Cxj6Jr
jqs72iNczXSDGJbv5lFI25AvS6h9C3e+c3hpFEiXEzlTdg3kKpA7omq0mhAPZGF2
lbeBZ3hm7XGr8HWDtAf/yOzGnhVxqLfqyKSbBZSdgokK7GWBSIw4bQm0h5MzwpzA
dUnwLQrQEnh91V37k8UTBqlaA+aj7X1qTSvUQfW7F/ZrY65Z9OI/qiLwBlrdwBFU
D1YjhqFl8oWdz7yIMhOye2/jBwf2HAhmVbKtQ40Gg5HJf1VseQkdtGlZzFwh7JN0
55/EkMCkixya5HezqzadVtI1vqEYrZnljowNRlSUFdq0/XQqHH+Cs7VCddZjFcgV
NtLOXj9BE0NQe5K6imBudW92XQcBfcWwYa6gnhM/1PkkxQVpoLRS/5RCbrqsyF/9
S1Qd+wFJYUNFc1Fn8pQ7MypW6HqaAkvfp0Yjmz3Azd77nAJxFrH9X2NUFGOoSIZ7
I9fFBL8/H9ytu3rBq5ERdHOYIZLZvNRtvS3SCAMO1NdIXJxdP2e92wmPXUNoWr53
uMGwiY7ctPfO+W2UDfzYYHXPB84tvMTXFrzgQibh4RC9tdUvtEGVaoLu81VNsuD1
8tmu03VSCY5fwLTeccQ02YqqE0FWb6E/V2cJ2y5ouNfSo5f/4BB3DVZ1LzfODiZd
PhfSqqfP6jPcNdiBqx1OTsGd2V6Mm0N40BoBpiaxIMgCTZNEarRvGloafGiFiJdr
aXUi6qCThvAbsNu02BlqC3Pmhm8zQHm9Vzebrr4+9UDEgzTXtrfXOT7YQTqLs5wT
H5NmwvAsQHjeqnznxaJo6+zsaXgtgYOi6rTdaUim3NoC2oAKMurhIhFdwW0wpF5h
Ym4yFyFOnJAu1eGPqS4n8cBxXMg6H8xhVi2apsuS7DedtnocUOlMrlPPfbjB+y1z
befXsjLgqKFQ9KX0mRWnsSUXZfmxDtHfTzNrBHXS3FlsMzVRGaLPxudOo9WB4L1v
tQ9mAbDPjiXTsT9I3mcDACjgKjAKvA6E5Fk4J7jkLlu5ie7RxYmmdBWAUqbJlDT/
MM4xsCeLMCAqDAgTGevF/FqPoKmGpwdK3HzhKf6Rhoe290pSlQm37GlpOq7z1YCL
y8yeFBXFGz++T1yJ0jNPU6wsqH+ShPK9n01Lmi7WKtoBSuazteBcx0Nd/2ZOsp5D
dU4dZOiqRdcAnMQzV5zXaJ/4XmwmKkt5kz+kis+eA8jKQ3h4gd10VsLMpmSHGZXQ
wqtIKlmuxUWz6MBCF8Awq4pgJUlWHaMoof9dOj5KtZi3P0PdlwISglPNqTTAd9ez
dMIY9F+iqIG7qQtKe4h6oic31F+PosqWNzL0qPiV/0j7ZWn514guG4rkR1RKaGLP
iFctag+3/seukJrc/rZtDWuQS8Ql1s5B05x6HrJ+4b2Lv9n1fRi7iJ8Ritfjn1Lp
vghge5AQR6csXTks2J3S1jZRUKH/iy1UgqHhB3yVSzmOT4tcx/4zQu0H3CklooAV
dNd53TUyJOrDkxdB4jBAICjr7YcggZFS7vvc3kOOy1eMZIHiIh2Bd6aQ/dy9Nzsq
4xCeOh/QtBeLcssQMIm3P6hWm+5iRTe3m8/BH1iyGRpvBmUc5slPKiJw6X64rw/a
ZUpr6AcC0Vp7ZSsAFAFP1damgJNvMVN1wNy9rHHcU7Q6ubooLnpXfmJys24uP8aC
mujZkQu3ams+d0oz4DbWl89aMXMepMr6DjybKNxcdEujoQIPqp2DdAiEpw+kPJNV
mVW3OTxiGL6Q13oCJ32Mk7G6F/r2PM5eRVQ29wzU7p8ijNrp8iv7ZO4m6WM5Iwfa
0H4IE8ArTbvKcOqgKvhV4Jk3Ze2yySAZrDIEvvXeNHvq9RQl+HmmjsjBzUZgavC6
w9DohOfs/AzUji5P1gHR+yyN9nmlFwP8Owfbkts6QwRNrYQ5JdZI9gvNlKAXgQF4
VxRtFPCNrltU+YNuIHevSfC4vNGSmeZaynGnBsU9kqZi+Adm8GZaHlUJE0h+PKrV
K0mDFzE9EDPtr4zigEpQJdU6lXwNrNafESNmWWbkSJSWWjsrbVCbkXvjc3UAzuut
+pOlfeW98vLGRfTp7o5AcYlDm9+cHmwYaYRNN6Kj+wvMTFgU/5SRxBXCbwGdBVlf
JCT+5Dfw9BTPy8n9vLQLkjqZOh30HW2U7G2APkkTmOvNnDgurdBFPkOABxkyuIB/
EsLgAR8pQ3yM4tQMcCA/E2W2jz0ZS4qiGwgd0f8p8PAoikfMcZxCxz7qrSYyqGza
0fjTQ5VbVDoxvpFCq2WJnQbu6/2kw+UI6ujIUgwLy1GDK5y+1ub7j3l4rKQqFHy0
IjZ73uJ9TPKd4vu6567uINT5EH1xBb4so0LoC4Q573l3DnpfI0jmxQobz/9yYEod
vtST3w/VOYuXkRgn7uO7HuRTXp7a1oSfjpyPutjq99+qLx1NorY/hTcwKvRe0+SP
ZOCGIuGaOWnyHphxcrZZjbDzGyS3IMarAcA9QXs2JGZT6s0B4iODVibtgeWcRsDe
SZjwcOGpSOe2vyW9kzPtbPgsfFr4koyAaqt20VnTTYUCdqr7tsFJ0Mba+dlV+W2O
yg6Zk4xfvEWTqfwqmEq5FDgJIvFf5Sq8Y4By5wEEWD396+HpQJCV4MLCxjMPTsC+
pMnMJfPi40zdaGq0t9IY7CApkz41BvgcF/g3tqOeLcY6u7IlkQgA+m5ex2GYl1gK
h2n63rsgGikvdp3ou/4TwOYGG8G1Kn5AbjJ2WnRjiomI+hb4sHqndb4oE0KQSj4J
hluTGaZsqo89MqHENf9U6T13M1kvxZLE/WBWTRG/z0Z+os1USATG1PuCQARzJUSE
n4sy5OybdqKPXBq0hSwW2gHRUTvW0uDFM/z9vm0FCufpxbjtAyoPMo1EQd+OsqxH
hDOalVnzMLOjR2beeQlmw/CIGOl9FN+FhdIxcoWg5ghPqbUbIoFt8asBB22/tQfD
Qs9SBOHMQ7N9XKhQLmPWA44fUfCwVm8ISO2jMNiZa3UE0yuZE4lj/h2v1v01wSZR
F38Pt2lWjMTCuge+lAROngdwghq2G4a4CDxbEWBVAUoGJ+mPIcj5EpS321j4fse4
4sxOTlGDqed6BY7RY8mkFZlv2k1SjE7F4sHFdfTWndoE0eTi7TNe+9NhlH8PXG+6
cmwW9rDBiqIiFCtwsTXkgnxvazQz9QS0jIiDJBuGdQR6d6ZHqPhoRAN09dLCHAaz
4O50xvn9ZbJ/GclnnO+SoMWL5Wjpq+4N0Ezqw0xovs6qyvve9JD3fgL9bMMapxyf
wSskHPizyqhYQr8d4e+8xAoDGZTdoFyl1IDprmICZGkQB51B4z1Pk+thCooaiNlx
+9HAbtskH2yVFIUfM2+ZY13Tl4y0xSPKL03oqpBPUImTOs+VCObiGoYLbBbIKhM4
GkqS9KlLSDMIphx+iefEkwr31JevUSCSlh0TCzELiHjFRsPVpDIowbIE0ZbpwNQ0
Hsb6KYOnnyceQoCp6M310PkKZBnjQjAxYqHCRAYzk03eyCEXLuBxo+buP4KTtYun
PsZqhYBYmZ2sZ3I7yd6IGjym/N5+LkfoFG5QeGz55yd6bVxhX3gQdg+7nIvT8vwt
QAC+/hlNrzj1qBpxF0uWu+89E9SyHJ6+HVm5AsH6uRltgxWQeoPFkRRmNZeJ7CZX
MeqX4hcPdm6HAgdwwJcxFcVAAF+8y1SCd2xdIFkjSsGiFkQlsCIW5fqIbL0JTTLV
lhGbwDyfcG8g+LfvYkpQy2Wi+HiWr54TCq033vvfNUQo4XNASiCDvrK5UmOGDyFO
MJMrqzAllzJhjyl0h4LmH2u/rT4bjCfW59hgICRYLzgIk4YRpT4h1+VVV+cjOcf9
TU4+1NL6qqlLSYZMGTFpoOIClqxv4vj1BG/zdG3MBortEmRKWBaaeQwbSSALDf6P
7oV/RGWI8R2tZSp3e91o6jVrtxSCEXQ7YQUtsMpOAvgNoLOFGd2VC8QPpAKW0Mep
L1guzonIbNu0JyNmOXf6stHNFfCCgeUa+vAaZ9SgonLjMhTqGQGaMc2LgP/kQGmI
WfjkJ0LNKICoRIJkc7z6BNOpee7dLJj3hh6fQdewGTcNiKsYdxOcHFi48a+rySMF
0HVoGed9yM7zEWW2BpKCCNuFpA7W3piLKsiLEhn9P+5PhhgsVHRN1LMAGFZLjhc/
4n/y6DVFpP1juAA0icoz7E1QnBjTsv17Y41/KFCzM8WbkkIKo1xfXQzJyghTdSpH
G/ZGS3SorWF74gIJcRnBRJlAn98PJhkJ2KqoKt5Muwk49EN5NA0Gwm/85JYxaYaK
n8NPHmO4tti/2RFEtqcVcs9addcqBM68YWZQz8ns//X9nYmEzeDM7s5uguwp55Qr
ELIC94L5H0gOg8Zf3KyXpOW+lM3JmGa2GpMBKFtddFYMY19/etC2ILhnABVNN4za
f6Msb+BUTBhI6i1mlLwMc0bwfylS+mt7HH3XKRTLZ4sVgIup+YXnbRLYcCXofEfo
wswKOqNiVJ5c1PGBNkv6I2u01qGRWBv8kv6kztJ9KxzzE3tK6LtDqv+deGdA+q85
LV44FPcn+F4gfsMFbxmrmOnKIiX+DkYXZJiDnKCPWYxBS8P1aosNem8I3Hwvt5H7
ugwict6VSHbg5Jarr7pUKDDiXdBhrF4vz+97aZ1DKm+p+SFxL3Nge3d+apMhovib
Tq2FT3H23PI46OD7j0eO1xWz/hDv+u9sSbRQ6SckGCsxFpQJYoG9VFAQe2lKSkqg
Oeg1u93mbN9hhRTrIJ2xwcAU9DNEE6eTv0+88BR0th9ZB7fppz4PXmS2MM5eWTIS
d60X4FzT060IPlsgBYZzLD02I5AyrAgDDDtg/Yh2QG5Vp56iRaG19veF1897dqkG
j+B1AWsS9lOfuoGvKtHFG3VCWzbARmscM3xzceAocCUxj+9dW8cU2sjbZjxTgQpk
EhIfw/7D0quUUemJ3F3KVFccZFNbBN4s9oL1D324PBKOYLE7TZbTBMmB2OhjpgWe
ahxz+HGcc+mt8JpMcklVHrEklQwHYevAa0a16bueLMwdBkDcxNFte3CZZc3xOayb
SlGR6kHT/Q5Gp9vFYMfIXJpa0xeBiWriRV6zVyj7cLurislnEOXkW0lUQWOlKRbF
NyaS9CSYMu67lrDlku9k+JgcSAloNkxtM+qUB7mIb7bSpVU5VN7DHmtm6CFVtoKW
OSt3uPpTiPoKazVjc1Ff581PHFk4OoIgKdqvRBiyepa0DJqY8TH3DGI+YodXMnW6
jv96Bt6ghvqbyP9+NXfez9oPNzGsWQ5tj9y5ePskgICsu3DHF69U7AiziUPCaGHw
Z5Wf7QgHnv1tKIR5WPBdvbkvo/tfV1LHpP/4yCHU+uUzq0+ISFJfFDeVb2AhPMd6
+69I9keX6FQYOvPk6j/ahsMyHe4+uPXpN6hvj5vEO2CzJyBQkjB61uPDJ/wwPRa2
lzdW8TU88jkTHs31iRwN4QtSEg9Dn8PbOh00fEFEOLGZDds8fXip8V4qhDHxju9X
Yt1RfT/Fcn3JZcWgLyteB7dwVaD24mcWQQZXV7tUmGftsmMO/uiXLVfCPIN5RrmQ
LewsdBxOFj18d4lmbc28U5CZ2ZFLiy+CKNAroLr4wrYxC625XfajTrQofcF3KVyz
u3bGEOevdavCEvDSo4bFlYgHBgXwbH/6d1X61+oAba0UOst561b+TlmrFodSXmUg
+GlgtFW8Elb3x4YAOoBDlTPhgsh8mBXPf/Swlc20pq7Y/aGGXlNNTbYSWhR5Q47W
ZtE4/l00fR3NqJvpsnHsznoqNAK17qVl+msLP/+NRUOJ9pVffYIQKJZ5qXmh30vR
WeezLo/TMkZDTR05bhZ7lQV3Co21eWGUN2n9jSqNOGdTaKNXN9wJ9ndJYXdciY/F
nv+X5Kv+eRoGVJeJpoyVX9YNTcN2fs895caTE0PHhIhGyxyIJZZn7rcCil7Wh/K5
UsSykjkPmqyGIb6jJWDtvJRBCLxLstLJq2U8CaPLSPfFrxFoTttKSN0CKdhFV2ud
J2P5jlXgLHIalKGhEi4xfGReztnWVCOdOBYuH2kbdg6QTc/mPvEGLCw/LxZQiAcK
f2HJqyxLgy19423PNvrWvwJ/zyJQDShKFqdkaYvW8+sXKk8dUifTzGQlmHwCuX2Q
16nTSHjuFdFdiYWlZq5m27Upp6yJYLknD3eNqa8+giUdK87BYsWKOizZTkyp1MEF
QhyaulQVA/bzpHdSUA0Fm/RMQSrNE90hZHAO0pH0F3eE4GM3TQ2oqYTJpokb7U18
mC+GWolN03lgEz7lWQ3mhb9zvYB1yJNeqxKB7xnnbR4bZZYcDUumC9x4GGErH+QI
jiZlytywDy8c5f2Ra/FGBIx9QBlaJFQAywJUNRSegSnCO5E67o816jFTalI3Maui
3Xb3Rsh6wIy9s9JIi7jSkQsiPiW0yK8NyrXFJ+gsVKSzmunVoUPXsaYKOJIz9HY7
AH7jh00FAEGVnu/MB83CkY7PN0Z/pLu3l7yVhRiMufWejDYJf5Qkvww8+502763s
w7EF3O7WpJIvBuH9xB4Bm/0NTVkycp9CPYRflGBeOQOe4ICvQGUDm9/WlyFSB6Cd
67D1pNUg4uXdxZITllV/ZaWz48UcI1rE/a+bHARz3hk2HwJLjQgPUHosR7OWbdc0
G4kr9RACJ7wDkzhYLtuWJl3aVhgYmtQc54nUasJQ0cIYsvVoL2zHxbIDt1dc2xRM
R4r8kcs2T8YfV0sc0beV7m8VOfCWnT4I8gzj2Dq98sxxp9Imq8bubOArC8q3k/Sy
p3Bbf67zCUNp/DWTNfU1vslPtXTatcWd74RRLnO5AGsWu0p7tSUv4/iTxB19pgy2
bt4gYysJBW13jc7BLbhlbW2v7tSParBeoqRFkWktsG2Awy88NIDP7zRvpnE32xS+
l735fkUdlPvwN0y+bvyEa/WEYvzX0HLwVVEqnaf7/oqfHHvU1go4MwwFnCHU2oJi
SBZt5p6KDQBEA/Tne9kOAleHz2apU5nZqy9oUg2dn+j6Yxn3aDQyCo6qHwYKuLQ5
zc7UyZkrMwygqiBOEOOJRvc0D64t2naAMKiChf7ALaDe2YSOAqh1zlcKzHgNofeL
k1rDbErj17rl0CuQ2Ct1VqYCCzkg9giKPWLPca4RJSxYBC7vyCKhohGvunhrKmLy
StzXIp6eY/jdtrUJ7Qzcm/4obx8ZNcUjGeqFxNxMsPdx+hn6EH2j0TvGKBjPTpNd
IpfLvazlQkDrkU4tjK/4hrRpRR23fD7VirjTlbAdHmLcpzIsxWkZso/0pkxscbJM
sIGZLYgsQgHOKfkHC00IINGSIVw01D58Fd7v7thNkABQikaD195jmqz0Te4FgXPz
jIXHbguYqJ5ouDEhaHF5oudG9dl4dIOlslLTVFu8BSqBmr1XGuKiDPhPL4A/Bb8Y
y3Nh81T/ePO6bOU20nsbqq0WaMWDctCjPX0gTfm/ecydY0hmI6pTM6V7PS60umKl
8gM69vtX9qdKC243wL6hmWYNG1mGtVAyYZefvss1DsJtwoWxaVUtHg/gVneQY8eZ
llc9pRGhk+3gsRlqZlptGkcWMYN0YZMTDc0ME/M19t+Nv+pMSzvQAvB4SOxDQuRx
ONhYeiKNL21KjlTwROTHeVuADB/t1ODmM3Nx6wccT3+Ms2YuFzWcsT4tPFNo2OM/
uO5VLrXz5HyST6BT+OunOXsa4ppUcAcZ3fRyX7CFX7JDAMqud3kWuKBOKFFxwCw6
vU6hElyXom9tjYBDwND5h5m3PsHcaDhzlmF9njSywWx4C/7nLZj4UPrxyaFqqJYi
iTp3XJWC5UbWQ5TAgKt5+q4LILBWcra6EZwYKU37wTO8sHDkZmisbn4f8Ud4e1IM
u52cowto5THsKLYosnZjnj72wP8D/j1HR5afedMajYQSeKmfDnBoR7mp4x79aT0u
po0LYXXVNET8EwrNcqsvn4M68zZQjMfgTjdC+xgGGgVV3DjFYvdZ4TjcdsqJU03K
scZVTuvNBI+PuKl59h1hXvLzuhjMEooeO/7iWxAhOs5UGcWHhbOtHL0Tcp19rjTv
OO4SyhHoXqlPHKyEhJS6rCKs6aDV3xsP6MbEuYmneTcTmIo9mq2CVWzka8u9AODx
NZIvyV7gLg9bVuWG4QZoVShCmCsC1Rx+e9II53/cclO40kDnXJLODFB2AbbILB86
K1TZrrf31xCfqoh/6PG0Psr/nyH/WJ/HT9vIz5WZJM+0O0OziXGhdmlcYI/MqBgo
brarvjJK8b4jfQ7VCTb3UUZ9YGgaKic/eGYxN6sD1hYNBi2EicI3BbuPnXuMafj+
aOqfl2Xx09v7t7ta5qDWxeoHoJ/1f/PT3Z8S50JDPlgyYfipR8EupbJro2GRJSUK
bRYmvsgDPMwdK0v4obL97cDK73erRoLScXxUSn4TT3ZOyKcxmG15d0wrBuJwks5H
JErj74Y0Bs/PweNOrHAmJATOxe6yn4fZhZiB8g/yAU4/x1kV8h5bKevvbKpJyDhs
mL2M2R1DIi4OYgjZmlpgzOniiG3lF6ftiPwmaOG1MWdRQTIUjuU4HxvEgsiK68Ci
oKC605O87lCqsthDmQHGXM8s01zmoDXCU8BPtc/XGy/20C/h4728d4ngqN/+4+UY
OJ8y0u2KJyrimbu12AsMQ08oTOZQ+jbq/8+RcMoVmRPJSbnnxdSizilIaH0MPuTV
aT8st7Lv0vpIA3QHNC35m/1scJd0r8vV8C3VxJ+3ZrgdiZAqMzixqtkCWUsAXqWc
Mq8lqvVOrfuMuCw1DN45u4p5ShLXsIMqD29N55mwp39tTpvaSQUQSkSrQbn2OhaM
WDb6fTimGwn036bLVJvgty7AvX3ntuJQswCJMnxM+P6f57lUQtTOXP7EdE6XufKl
OTVYjx98gf0FjL39h8mPHpL9mJL+qCc//s0Q7mHiACzhMcLKYRm4ZuDuDYcClITR
ojGYzkbi/olFOvLPITHfc0ycWmn8E9ynzzwhUnt9KEA/aHuiFSizFnu3c+5bv5YQ
XNg/TSaVqwL8NKnGWHoph0vIkMzqT1947mHYaDhIq2TjnMHdOM7iDeT06iaNbAbm
g+eCInJvE40IB7+K9aHkk1kaziA8EtmCtjvvqJyrCG1KZxz4YYjOiUl3VW0QYL/C
YebrkmUn3Y4gPmeSZq8cQU1x8Vt58/cMwkYFlUXuvTnbrpCyNW6+1k1wOg2V7Hpx
5BCKVZrNnh8I9TQuTl6UeTdy1q0cD6PsxyUXjFvpoixhTz8lg7HF7My6pZ81TTBE
UtuTA2yyzhn1i1ceTkIKsICmrg9Ic+8pPBs0JpIOsVGmTglSFlCO2eLs4z79uI5h
XVWGMfxnPDHqaRsqCotGg0w4a2Ujqwns1gaY9YIaRugW8fsFpfbcB2bqqkbpJ/1p
yD7X5Yy1y6HlXpwzqWmZEyj6V19SKpYqt7uWVqAaKxgxUXOheVSLQWSU9OzhiUbV
1YsXjZ7yjaKkJHUajdsMbM3oCM8JiFBlH9jXOZ7vHwtbjfreJmSEIoGmSxPAQByw
ySPdParSX1TbtXHuEa/lpe9VuplsJy8UU36x22DCcIZOSHBDg/WU9YFyg+Qmh9cb
Bnqvzem+q3hP1aR8CrZbS2uFWDIwuyR+WwKIAy6dN/t824Rj5mk9XXTO+e1BVrfJ
UBGO1fCQuiBdxbijHPdnB3fBdgVdCiEfV7OsMJUVDr+0uh2foNiHbB96PxiRVinR
JEQXpmkdqFgN0kHBN9sUqcGmMy2kVBtnxlQZhhqOUPp69okl/+PWauBA0kEZ/MP0
C2oauwELCbpHle0kUrjAqD819vlzQIJ1Ru5jJ3KEXta7N+neimr5osKD/f38XR6I
4N6AF09ciFSUO3JQ1lUkBtT815fKuC94jSyYANygwzSHq29uWgIIjR6JLFhvP1Nm
gPEZhMeuv6yQ1lURO/VHp+WPUM8eVnORIdD7JsNbKQJuPdMEbYOD14jls9/vt7EY
k+NY2VYq127MuyLYF4G51oqeBpmthZIMe17I+7DQx8j5MnQ9Ji+hr8fuDNPznzmt
DHU6KlSamf9iStensJbg7w/BYZIP/iy2GXZ94aYBn7JX8FsKfMk/XSFho1dupPS0
WbPjRn6iTJnm+mWsmr1kYSUpBK7P/QsKbMEBqSkYxN8zlZhsauL2HPMlwftQ91Or
1SXutEmLv2WGrBxY7lhOH/RPNNApmwHjS17lAG+nCRc5OeuGn1sDr2CZZrNELRxD
4TKiCqclj3ZAI5qG9MJrm24TO1z4hT1jXvAWLtz+xfLBK2Nz4s0HuWsaiwQssWE2
0s5y+C7sqKtlOEWcEL5XWrfRFaJ9bRan1wNEZvKOGBcv+n3k5mgI1h8nJtN+E876
YtknHeq17t7NULf/aCUrZFUlxeugb2Mq3b9fsJiM9dbKgMGX0ydY9/+oR3+tiPEF
xOyuyZkudpKSO+EBmCfBS2BBlRjJn1j/nm/jxhCiz/PBuIuYzbZb7+cV1UD2todh
Wp/Vsbn+hP/6wMWr7MCqRwsoaO/zIiDsHl6AF7mSwe87eSHMtKUL7tkn5tPN+K8k
d/el6my480xg/xSYbs/ydLYmxlbiDiV9vQSXI+vCGUsvtULYR2cev21U/cOkTqIP
5kLYyFRcV7LWQlaLaLSelV/3cWbi84MBPnLJ6OqHCc/gCLMRWp4NLygbCGj8Mp2a
lEHezFYCkWh65925+g4d89stWfkDTx13ltYYnxbu7rDbLdJSI6whmwgQIA8bBof6
4fI7Nx+6ZJKADALMXzVU778wHjN6g9ijPJ+so7X3jYXui4HeB7z7mgfsx9A22XZU
mm0B2DUdfrlGBjH/h/8CtsqyxEpimEp//BMyeMzbcwcdrkvsV3iKcGYr1RIDf5iC
xEqLqc1rJe2Lqs7PxxSPRJHI8t2hcz8DBu9BGSZvCWQ5MMYpMu7+ls3P2b4iPirq
b9orup1yQHzZ6oOVyMsdy2rATQfctYHW+jaLSa641Jt8HzU7eWJgd6lPe9Q6d250
cHO6I+wdHXghFSWKsDWgeNnWa9xqFfENeXFr0RRowICh5VYqPljBauPPXnwpOfEY
MvW4wepx4QSW2TWrhRHCj57nyoPpFIEHiXRfAWHtBAw6KMZnutvtnvAq1z4TWhFA
qTfzJS957pr4JhFY+CflOaah+u3eg6GrP50e7qW6CEHZUUIyJ3tV19ooEjD+gAA6
63Fe3atZe3P/GNJdq0HKoFVADjxCnY++yFcDLp7QnDjK2B1uGj3WBAmVzliJoK6R
5CdYaqVIW2DzYvDaFdKGbhZgl1JNccn2VfHqRlScZqE8eTLBj9IJJRP0bEzQuO6h
p6XAzj7sb883kl04JMQlYoM4Pf1s6daHHQmo0llBpgba/fbZGZ8OVW8nysstjfT6
uK+z+Gp/ZeGADCSo9wZutDyih78e4chMXlV0ZwyIW6Ko3VDxbV7Vle8Jq72VJ6Pt
hRkSRUygj/+RlZVzOBIl9UPNuqSoWLL3viMcGik7xG0YG7M7FtCH3BEx5v3Q7g3P
FusYjJyDo6KSe2T5OeL2SSe0+dHjePMx1nmCVZ9RGBHHSEbTlPlNiIzTEMwhNU81
OPBgva/PEj9hFjBTEJVk6/K7X6kFMX4p8K+vakhO1xkaAtl22arob1upuqOLylzd
LB5Xef2nvgnk1jKpywz9t0c2LWf3R8xU/n4vTq6dS2w/UHB36Qu10GKoIQ4oWwNd
P5V7eYwG7lAfDQZCJD3MYDWAgre44o2jTNnvuUZXWCa2NTMkFY+L5TuNrAGgZELZ
MS8OIR4/0suRow4yE0832YHeu/WirC2hw9C8BWTZDYqcUN1mhXj5cu1NJ0UFR4Sp
jFbITZgS10XW0BsSlZC4MvOBZSFLai6o36UcHCwPOe3QiOui03rNF358Vp5VMOib
/IejRJhCmDWt4v5Mpc5XtlNdjYDLA4NB5LDN6Fz9wCUNsYUmduseWy1H1QzdMKep
Mdbi7wacXNnf5CmFXi3cTtAHvL7R7LScq+2DzUt7Djk5vM0PV+84Dt2j4V8N1D1M
v+PqKPLCj32QtNlUMaPYgw6R0dnn2Jp6dm76VtX6QDyZQax/ZAgKqVNhtWfZGE/W
HECgguyD1YN485GzkMtr3DHbjYeNvY5e1N8yY3tejZ3l0C4oBsM61WCe3Kh6y64k
Jr5FJFBNCyTYfl/GHJlvow8FLObE2MFo732V4ullHTqMfU3HE++wS6C2o74+KC+8
rXRsSqmL17gjYkn4X86iY+vO09OecSI5UJLrfhhxxkTZWIddURp4OyAdQC3y75er
c8R8oOj8ObIWTklifavzBO8t3uMjMhORHYOsl7JT7vCnFYcxHOVyqUKWcgQjvMz3
q0vC4NslQJtusohFbMlp2FcNy1RR5ICWNFgKrf9lxXklCWNdszuZQIJMc5R5Z+SM
mzjrB9rs2mFq0/QtXO4TSs8pg+dVx6P54DDd+NfMOT/4ARAO7iPlLdVuoZDL6+Iz
IDdEkF2WDM+WIazE5F/L+r6JizvFq+CMAWJ/hKH/FlJoWLonYfNbytU8l0DQTPvY
Ia6m1icaeU+EdZ6j9EGLoCGg70QDQ3vuezWUtKLcrXXeTx04eqpdbxxAnVupM5le
IoswEepzVk2OI8Sl2JGWFCJ7opROg9nTkEk4hx2HDxCUzmBm5JCh/u7gpBuLv3TT
RKsTQPmcZw74f7xQGoh0LWNw+sWpw70gIS+Wjr3D0peZSH2+L8hD1XNf5Rft+950
+tMVQxkqBAMcX81T0x1A3gGyIupXoCAqccWwCYPCAnmK/NCyC6lizzIK1lqGgL0P
JXd4OxYJVIX9TKuwIk2fN3R+j1g+kLcvlOFjX/arbI5qm9wdWXw9pWxMyuFPv9kK
IC51wOGq7aDwrUGp5wgSJ6zX2aUV2T/eqa1mDRavADiej732i7C1OaWOPPCIENcA
XvNXhsmdO8XUC3GgNqbRYWjdOZEW4+QT5ZWbTiAxbGpxcsebJNAIyW150oX9J6qf
2csjMIQ9xKjiXX7f0sZnxh/UZDKunxCtVMqEW7IFzAEeI6tt4P/3OECuSdPZYlPB
cR++58em0R1Vvkm8HoyN09fNN9KJX8AwZb9jL5TSz5BwqmGHKGonhM3ENPQsLx2m
ZOYBA0qgDMupuszg3DeqDVKBfVWpJGE5qEuvGAHU9YBR8gng8J/pbjl/5KZrbwKa
jTaO2eNxlpZWrj66fTMMHTnLDExWzIxgmKFbYqSdvR0vE3Kh8fQPGxhiIDnCbQqa
QwIuNGGcAJakiLpcJJ6bZuSFJG9N/krMFkj6Ga4K7z/iOfS78V+xLV7yciiTaqNo
m80+NJ9l7iPZa7iVTeBag6Vu4HnWS2yQrSzapoVTU2ZVwSXtR13HEh9yBCCWijJU
q8RaGK1+TPnkZDhbjRCfP++uEiYBFeOrBFTJd9g7Sz17UlSRp0xNV7FD0+haWRsv
xOttqlyqKkNL/goHdBBdg3MNY8sAJfJ0t6tik0aQYR/MsDyMkO93Jm0NUJItSTCa
tyGzeo8Jq79x9gqkGy5ebb+VLhzJKVMpldfvf0cUx4teU0qpBaQYLgQ0OpDcjiJH
HAqma09aHSFgrmLtwVEr2Kdh17Ag5GPZYdfXDSWKWZadxSHmWqx+qj7g5PQq288k
kdq7A8wo4fszIGRuDHXzyf5+FF7od1fLvy6prRAP6n4/SNe7yEtOsMEvIycuvERH
A9p/AXmTgnQM1EOt7V33tOHagF44SQ0Flv/mv3EpfCoeb8eZj038aqQZ5yEw5geQ
vqaLb16+SutVe3mnZ8x6rDBrCXiz0brwUoVMsWYC8LQ2d3gF+UwpeX+DMSLw7BCX
q3uTVL2oRWlkuNk6r2LwNBMxn/ADPkAhr7X7V9kXRXDBL8n7YD+c6Eg6Oq/Y3vfs
C2D/DeTJqbQeude4sm5V/T1nwCY2knD8jxRYR//Ix29d8Lkw/NAfPi8pikiPbxkD
mlazMdEoZKWNWF6oUGaeN5QMOKDm65fpfPL4RzFqIhcCODtaWxaPeXto3WtopD7P
4WvKZ/43a74rZBPsR4wsdcpToiYXN2exIMefWwOtQZBTqnATicXFYxlG95IYXMYb
UgNiG77QfvcBUbbCai4ro7zUaczbQCzmRW+P32CBTIO8VyaCB5P8zNk3/4++LyYw
zDmp3DNoZan5rF8G+Fwbr0rblHRJKQDEW+FqVef3Amxbi0cTHWRwo4MZFaDJiIFt
pCEz/GEH2ID3AE1Lh6siHULc09GHdJJhr4FeT7Ns+PBxcpPFzyOkgG2LV04GD6OR
ZtBbWLxnQ1lNUd+35GTc8KL0Ne42IkTK9o36hyyq9Cuw71457GJ7rgKnk3C57nTf
V/oKLY1TGspWDXcgH2DkFgh12VC9J/9DIFNB65mtPlZ9zx94RRkNHnwvgbraHygl
Ef09YrQFK4LK+3Sw81PWSU30P3lezcDpIbbpBkfZeghXmJoUh50tmg6ezk1ImCQz
1LHMBGNhH8hdN72kzS2crWzYnkogxnZ89x8vsXfn6NkZI3+PNRe+Z2oPl9Nhgywj
/+qRTi1tOGjuO5rZ6WKurwrbqqoms7nTazEfkqRSPMiT86qFtS5DsN0mE7JhIrNV
1OKLuq5/ZYk41GDsFnc0X3n2JvPqqW7NsIfi2x2XmwkghEH9wXR80j9B0gdGq9tk
Vsc8NPMTGnwDUkpzpvgB06j4UYf7/EQ9k805e6rg1VGOmiB6KCaCuun1bn0Hpv81
QtY9oTSe037QWOLuPJ5OROIWJWR+tpSToRGkXJnxd7x4BqjFxm/oDZn5ciGJfxii
MMPFF0Ri9DlNbn6Jk5M8+kU3bhL9V/JWsEGdRBZMYsjzcfDZoaGdo1xJvdw2iJ+f
dUBYpzPoUAeblkwaQ2vGxuRixbqSay4BdFykfvMDGnuKUfwe2DtGjYJ4651xVSiJ
2rU8MNpPhB9yna8sHCRdHjXGfgAKtEKmxsh+uhPnkQn9zvT/aedeHc3ZF7XdYDbV
Pdh2IGMIIIK5UCYnZpSPjdaokcBxaPUhWaf2q+o7lg6aJzMmKW/kWIZOFsQPD0c7
hmJZ8cAnt0lkYd/BS7+EPczv3SUKOSWflVSpmu/1cBuQ3a8Xhi5wmKXJwE/gcHVZ
/9w2i8pYvEkIBuM2PknmXQtZKdEMcksfzK9wFEg5aR82UOrFHN25YqWnyA3y9wOy
e5NHNN69Fc53o7Ll3VQvl0ULjuQWvJBZCjzvs7AQUq512VS5o+/WfZRikSkekqeB
z5xqiIFUiRLuQ1Yti0eV/PVyZq7Ax48p0X8ZFkJOOEQwoiDTVzU3Fqkcua0RDcVF
lfyO0xfRBUigjXcCFDs70lsY9NAYzSV9sRLpOBZJxP2KzCp8J1C01IGJIlDSr7pp
AkIwHxzbtYPE4jPqni5dPbAkJcOmD1MtjIQjC0Mlxhf8IdN3e1gpnZ5P+uIRlYEr
nUxAEh/wd5lgl+8KKltu8sOL/b+H7ty1G3ILf63LlJnWvbls920XlGbMbnH+r50d
ttt/RABLGLSjBiaskSocOsaFbyln4hZdsYBWZxNJvTyNbTAGq3XQ3D6NMiGSRGii
xUSACkg7IJTeItRbnbo4oFYoHUBxJfPAzPf7YOWkwlCI3/QvQvfCbDqMDBknY1cc
sWLrWJuUfEaCzJMczoMtRBpsJZiLvZDl50o4PT1/Wp+rgLsMQwlsN6/MRqGVyPBX
Rh622NjvlzRm+RvgawzrHUV/3TRTUhYF7FuQGP/brRmKsBKkJPpWulHqluiIMHUa
eRwJlwASEoradcoFCo1HoGh6RedITW04rB7PxKQXY3hWw8dGNt1RixK8Y3SgMQC3
gdYC6+L4MGzn4K40SZLDiIUqWyrZ1LiH4NBBBK/A30Gyxz4sndkwuhhIxnjQ5Wy9
1WCAXz+nKcy4B66c9b22lPMgJYfTFzn1tk1lr9lk9Gg4Rn5jU4mq8UpJcsyp/TrE
DhCyVyFq8NBNpsKzFbA/yfddBykvwGCfvPy13y9rkSyaCqOk05F27IGjBzjVPOfD
H5S+oh6e7LhglGJyr0ScJ1AJksM7VOuBLGwoR0CDj2EjibdnYwxktkgbU3nVnD4t
f0wVWcmP4//gv3WsiZw4mEdvR0TJ87cB2a78vdizUOg/RfRWWu3t1fxsZb/IBCwM
/TM37bi/hnoK/g7qDSF+J9gpJn3L3JCN4AYqxRyguatW/I3t0lLAeeYKNgiAWNlW
Llc2g6cFnY+z9mOMMNRqG0tqnJjtOB/XVfKSJeYnKGuzK3OMgENTztXE1opkD26o
AffwpA+RvEeY7YufokYlmAnru1h0aadso3S9H5ZrOSw0TMMUa+hTSAVpUzFInytf
m/I0lJzTCv7nLMMWwnRPPZ5o39ITSWRop5s80fQ4WnOa4n7323WrPVh8Y8OKZpjZ
HTXBtM4/Ni0TF3h/SWb0y1sfb2l9TfFHM7nklIdD+VMIjzU3iXuuYkeW2I744b4o
t1AbY6P8jm63OCTJTXZ6+ITaFFU2iuoqGCphGT2XcdOIzleZz0SHJUsqaE3vdXQp
N6qNDI2LF+E8cLlkWCIWD5PBwtuy1cKcaqP9vChpOLoYhY4JyPyxFFNwnCcpGg7V
5JZHyWf/yQBuZtAj57QGp1pD3bcU1St2HmlOSExu/SDkQHLeGP3NPDU5bjVI1I4B
MQInETrqj242CzIPeG8JU9XKeydIV8HTTS3HTCJt6tnqATnTZsUYcTLPAlu09KHP
0wVe8hBQggtUfMf9MCUrMql5Whn0lVt7eA1NJ0mj95XwLRafpaYrY869HURUvDMx
2zKzGhZmlbyiFI3Gp0y0T7fQmkLphEeuZU2uhf1FVdHUqshsP225Io1XFbOyCshb
JtReCzqrq0WaXIj87dhp6w+xkm1PqLSwiCnzdqF9RRAUN3HXOmV4ZmkuNjn0bA00
7+4v9b1eXhAo1XICva1R6OfPJ2X6KXRqDW/obs2hQ9Ef8+bJf7KOODelCTq8S5EA
f1hJESgcL28uELfIh2sQBppqJbI9OviJGYdwVIP2GCmlbzdvbNuXH0+w+qZS9LKN
QT3UFTBOmt+AkxgoUZu7W2GM0frbPnf/E4xOU2gejfN7ObScfu+ZY4zOwXbzWhBR
T9qqo3RIExHxbpmDaJfTbw9Wx7XEd9HDrJ0gnkx6Vdi6DYNEYszBfcNxPlI4NScs
AjVGtWlyQTS0PB+C9UP4y2uOAK7bbNRD6LVoysx79QgLGXABVQRnf+ZbZh9rQmlf
23i7wlT4qeNhyNkXxniUDTFemJH1OU27sMvIzaaLb0eUvCGZCQZq/NGRgagFyKh/
FbytQy+kotdFvtmbncaPa5Kv7bxuiDYU3+Lv3n9ijeS6L3o215R0UKZVPKnh+haL
MB3fkZkdIUtTnkDQOziqmOTaS7dsFPR7wZsmTewy5gq+KU0MtW+OHhnv9ndO7bOl
FKQm559ndwD6TxztHankLM5481Td/JlD+WRwDIEiKyYc4jADUKGvhWxn/lNbVhOD
2tuExmhKFBSuhW9pkaYzXtnnKdwFAOHQ/k9J/GngW1+bRak+YWK42T/WVPcOlWMe
B36rElmJ+RLx9SsOMRXcdb0/MWDM/1YMcze99L0j6BYx5iIUB6YX8qf+qqBy3jbM
93gJq21AUq0pjzdf9ZuKXpReSNw50MgB439NmgdfQdqAAlgPS7MghVEKmfxKXuvc
c5nDIMNJEozWobObcjoqSI3uKKrOlcRquGuhthQa8RnPc+dS9R78QETSeqasbopz
v6oQ08sHJwzXK5wDSfqXeXjX2GXlc+ltCo7Hz6EOAXH/IH/3lC4YilBACdIM/Hhc
U33LDI8j17qxdHFaU59JTqf09oMxbPrl2+XG67RtSiHP5v6cxbBMQWP0NyYdDZUm
DmtN5UNXHHCa35/OnxY2iVlNl2dyUdNXUwPfEAqmQYsNyWR/nIuq2PsqDmlhaZwC
fUVKceHStJd4fxNGsH6McYO7untDvAUAOf7PVytFMQuvXdwXQa+iDTrhtx+oAPyf
6j9t5ZQsJkranuBrblDwAzLJU2pjnhf9F+OWYACG35ZlJS1fFE6xxiWEypUnAkez
wVjx98LJJghaqrVK8DuXmiNGyJp9scLj7fkZAYPBDst04mxhyMDLooQsBC5X07R5
itMmgVw0kmlP1HVFP2GCK8uRPPofW12w+inowc6xultpkiOyBYNGBtdrE834T9tY
vOuyeIxkff2ta2BBqFCrcRgyg81YUq1et2cSkiuukcnoVStGdxMnAs/Lbt1pwrBL
PuLYMYwPdBoDp4cg+XuB9OcyuY+HoJsLHZzHgB1x7ZDeNZb22SZ/TDMhP9Qs6ARH
+zjfxU16EYnZvX2XV2zcPh2BoQg83HWkgwFJdpyz0n06qtc84CuT9XmhMydnSEU1
W6mM551n2GH/SVngVuOKCDmR7NomLjdwZs6+Km/rX1EMYWkcSDBgTcHlqyQcFchH
GeIXDetjTs1INrX/hL9eaVGiZgWZEjVCGv28EybnTpCAbOkDUMkkejbU4DlHT9T1
xj8HdTttE8RPSSoc2BKl+9M58NslXtU93xl8ux7xdmOhsFdTVUEUHmdEI/9vVMyF
kxaVhw2chE8/6UVamwKlkcR5366BYznm5lT5sjKB1W7uWlX7zeQG2FK19dbqP2s9
58Jc04i7VFXvthoJPZYqwEfSqttvKyABggCTbW8qrNqvjcpNnbHrMzRXF40BI3Un
U5VreEbWgR9lBPnpMnAVn14tkPzVrDvCGRiKqW4g0ZROED2BWtfg/fIhAA2y8VrM
qaL4tjXBMIqDDyYFwJMRzVvaH6INuhOrVVgnKgv/hDDylO8Xn9ayQIsCmaHFfRVN
I9xol1lRaI2c3W0fyyOi+++4QpXbonJzSXQpC2nMHa63Y7bg7WzmiCJWfBfJS+rM
HTwD78spRpQUzE8w6Bk1YRMdShSOn76/7v6eA6Cb6QsrRWx6LJiRAqz16m+D8EEd
l6icPr4Uv1ZKixw//8EuvzaH43vPcj+WrY2rkXawdswJ0FNF84Qgaop2QtqGkiH+
CTHkHRxIOviWkhZIsbwcIGQ6TXQN6avTwEXb3f38NuXG5qV6/s9pxyFTe8S3R42e
ooNdDqCVLSQ05GfbydCMgECx9v3czW40hiQJjyJllx+Gg2AGsQs1FExcd8w4cGMj
Kh4ZxGSppq/JYQUhHW0ztGwRgem0mAnZY1d92Irv9dEvbREp4ig/X8KWyVM4RXZO
mOrEVdKO6Rm4d4RDHhVcQipOiDKPkysfTRHUjCArEpaYSo0wl3iZEX8CZL2LzMts
k/b3PTL22BsYXR8x2WkMamTUvO5p3rHoz2hvuSbzpWYVNB+zp4v/Q4hKEIQXakPx
gEf1X8hJT31rYRztUBknzGV8gAaZBoVWpX2p/irWLf862iQ/1uf9gOgQHCqlY2QC
leP1HmJLyEbI2RYg3Znna5ONGdB11TQ76NenxZ+9v3OXYe2SixiZgDbqv46hrpm/
GfsDiDD/D9Yj4+l+21xtn9MGMyZeO16iNRIUtLL/hCxCPTExkITZc36hf/pwZd0P
W1epGsLMcYfNEtorZSxFxxjZHZJ2bsB0dmXe3RsqB2Fnx+gbpTjD1WiH615aYqh8
0AlcujQXUglculoKHW8cuxdnyJA0a4nqxVZrdbPQCHkQoihWy//g4ol3KhmP3gJt
MM3UYIi6uJaf6OYT7nPUsfn97m8K3tSWKBWJva6ZgW/kGhtBAQbfnL4O7oeKR9na
S6vaDSLkM23qlt5vEZKAcHM9e0DYhIJEeMahu9L8r6WXFCpfduwzqVlkHEWvaTu0
FzQfySg9kRXUxnj/fsSJfu3hrgcQOBXHsawBmL7FAPxCMSbgdw6wL1iAMm92bhWF
0I8MBjhn+FNQgvPbH4DEquHYSN8ba60M0cKb4NuBs6XySjd/qJaiKnmD880tIld5
l6+Aq3nY3xLdGRF6jy/6lpkHmaDUS+WqiTRd8vPqw0+7KWsv3SjS+bXEe/haWCeb
u1uPaAaHfgXuDDQZiO9xtyJYgWoLIW5J/uZNgK87K1l2wKoQxBk2obWHXmwIBlzv
uqi5dbqrcaMqZdeHBaguXYC3X79QpmL91iZiF4OghAGWMxzd0OiS5sCVmLgNAElb
wY3OTe+MSZsQvEbHFOiGT+XElHcnV7SoJrnGvLfAgnmx2Kjs9yMfD9ltYnqli0A+
k80sYfBievzUxRxO4+sm6jJu9xAsvD3rt/iPhEZ1Ed1lPbucykN+q+LrvyT4h+Zn
kc1YdxZSP6KS37n6AWZwze1PWz5ccbX8jzVXHtB1IwotRbuGKfhRyhxr+RO7jb94
u9OB0G4cHkz20jyfnErf3zNTMpdKkJ/N3J4IQpj+at3k0BfugBBJs5dADW5eP1/2
OpGgcb2OFQT74hVz4qDkB2sGaxNKzunDsJClPyC7JU4A/nELpbxz+3vNF3DwPjni
k6R3wrcWT+kfRPcXschUtZOICwSQty1hdfWyDKtCD3c/uiHN0dURokMfRPZ1pvh7
CKNk5l2EUmy7Yjaz933VO7fnGcbQRyaDXRJnmxeu/+c7jQDq/d2yGY5FMAMIgJbu
Tu7atVbHLG+8hN5w32pD6NWOJ86FfUaepVcVQzrCdE9Irr45qnuSXCcCG2K/4wmK
9Oi9zhwZhnBLbO3J7WDgev1H6SFfXrEdVZ/XiOUQzyiCbBOpJcqki6VF0d7847vH
M0XC5kwCtsN0NMtfogBkXWWq81V/TH0FF/S0RfKDbttWNmxurLEoMGKC19MdmQMe
nrgiihPVT9txROXGcqtVqiWS4OprAv2HSPdN6IwKYGv10/eFZWhyXvJaLcPrl/wH
LCSZVeNJ6CBMxDl1dVdph4vXqCpIn+lP9AiA0QapaysucKihj/NNH+LoZEvX9hoi
2xd8hSCQqZvdvHIN8yp8n/x9kQ1UiYew9Po2rjuQABvMLmfi1n4UN87jUGMHhcFW
wbAFx/eJN/3R/WColyGnjSB8pcZBv5zVKrXSVTB9M94UdiQw/1VhaPxWmNiuNThp
6riE7hiQjIKYmxPLIbW0tLbqRfrorOFTCNU33zlnkWHqPHjULPerdW97G3n0pyhL
6XpiCkD6qFQA2rWmwHtwq7dlQm2MEHFEemllfzBimAY0+U0Uhw1YJbqFbM/8dApu
PXXdGLIVpwVxPpZ4M3O0i0R+ZEEJLNGJdQgkeMaKECbWLG4PsDilybwMPjce4Stn
S67gsaz6LebP82R8HmrCsdAY+Crhx/d7zAUq1mXXuyWba3sNiic51o8B2bLgNX/V
+bQ4/hkJxdqqY7/Vqac7SBCRcCaOZnO8gscDZ8hKdg6D6gAASc3t61d9u/yx9O2o
xLnSqM5N/jQ3NpAW4SQ4JCvOHi4gvcG/s/K6Lrd843UV9VYq6hiSdK1uwupQw5Gu
7VA7G40bDSC0ZtPpez8+FLGgn4UPnFdQs0SfFdqpmsr5vj4/3qS5BxezHH0ccuBz
aqmm3IUvBfvenYaG2x9PWfsGIjcQ6bXm76c6K4a+7xTZXDEu2otwXtbYo5wqd0CS
Mn9SxaIySovB9W3vJnHaXrxWYyTmZHOHO3u+cOnmyYjndToTJLN7RTwJGtsmiB4G
g6W1Y77RtrzhYglHnlKUH2q5P7kQxLzyGM9TmQpusYiyo2CelpKVEHm467DE47R8
aifzMHN08e9u/wxS/0B/FG1+EBdtmz7JgYFW8HcwHXpOYic6WthkVURrvS2S/qH2
EGW+77TKUL4Aqhl3f8Nm9ywsgCcSZSQGv2EsBoW3mLfk9aUfEo6z/1mpG/L2j/TP
2NXKlt7SxW5qUq+rhrqYz/9InLt/xq2nZudV4dqEacDPgrR8l4DsO0C7xrYGDJ3W
r87/39OCWpBbp+ErMaW4FIxPoGzQhGhivoTknAR7vncBQpoGcQQPsk5+BXgUHjQO
fjwK2c2118d2VPbPJGDajCP7+6FqiV5JWaCX1UBeSrD8sTT7BEiqMBZX2SdkF519
ydeH6hzqMlyhROy6tgCvj0eI0fG/qlVxqXo78dVMZP0d/15TBmYuYAaKMGkCnNmi
fZOn3b00ODHhQmgU9YZDCEvAFtffn565BIxowsAfZAnps55JT6th5NypHmKL+7xf
rN0pp6H8wUHXXgN20x16SS3d4W4Arg4/rcpN2G4hb9wBTf+5g0dlSSh9knMf6P/t
3nPgjrTrbzM0fZRAh6dz5cIIWq13j+1oUNv9fOae+Koilhn4akz74C9vEfkARn3E
NnOdEDGNJobmDqNy7eUe7HohwNVcRtKgmjlxm/Xd5PAt9uh+NxD5JtB++YhRjEKv
CS4+7qyVb0eaH1ptQChqNho7pbbn1E7Ikkz/OqkjoTXn338Z/8iHJbvLXEVXPwql
sP5lH+f+4ST4SPl+9o9f9aAUvq702zqpKK2x4YvCbzv9A0gtsmtFOHOkQZDguF14
x78D1mn0p1KgrZlK1xoB8F0RTXPCi4lcIa9LAmyiiCbZCVumUgN/qyVyLnpe8bzk
03SYiw8zKj8y/m1TFvPTxuMeZaVDniabPrEofihjxD26RLAs1jYWJ+3aIOjeaDKl
inyWNN4CNUjh7YOp3T21aIOXGPh1i7I9vqgY2nY8FaYRXT+oO9N3LQS/a7ZqZ7pS
gm/wcR50zUp/nw0opHlhS83acfXQVyJwlZZqln7I72Duq4rOnfk7nEWkg+w52iPT
ro5KSA1Y+usjQYilnS0w8uZhiVW2sUNYnbDQ7XPfKM1HfnAggUYVVvrSPmtXqzz6
CXvm8ZOElek5PA0c4OcMjjznniHrEt7pGg71bhOXpS2SOBKVLnFgr3SqmmycHIF8
KpA9FfwA8ZkB4bQCEbc/8lpwtxJIJSGXb+0Ennxqf+nrcdv9OXgToCyT1w9aO6fE
TmnQ6/XI+l1l1ighb3HZIAtmadAmtGfYgOtUA+qDQktGDxKBWZlKFOr3YnpORe9X
57wndVVHXkXL+XEDo8E3giq9JfzH/bueuSS6C8akY5zzMeF21C8+hYAWfQIf9LNq
bf87whUNaMkjG3cc13/1rykz+qmgqduX4Tqziax4MVkx8KVBCzpAppLp92hA3b++
nZPKNdR52QN7nZrT/JRfrt9ypGWTxW1Dohk5ED854146wUP+tKr1eEUoxGc8Z4ef
TglqpatdFHFF/WBp/VaxtllnfjIBGn3ik4DApvJw1m9KoNaRzl0XUy531lEPh51T
9ovvMg3fBDimRgeU3Qi1kjUmYHwvreYzr+mueMDHvRWvrTyOt3w90ibGDUeFq8md
KGWJemFPu8VkSWNbnv1zMDBQH9CLZRm0hrHoZBBoxbnubSdF3rIELkNSU9+eZ+jh
megmlCOsZ73nc61rBv0tw68lT003S28kj8JZL5CzvLH3qEmValo9uuPSYzXlKfw7
qPgdbmE1gjgR9YRD1IDqLqSdJ1Lk8ldqni9yAHu9QHlL0BhR1ja+26qqOh0Jz6En
Rhtajaxnax71Agsibm24l1PJHuKaQA0QxmdPbhL5jfuw32t6WL5/xfnjuNrYgLDz
7JQcvVKMTR/LTd/Sbu5yxtCRtrYE1lE0sbcN+CnCOJx+IIMJrK08qP3cD4iJNAO4
FuWAfkDneRt5j3zJFSKDygf/YtL5Fa82XpAyW+emlMupy1P+RDDOn2+KLwjjV9G4
Dm+My9vJkikDYrcek8AdnZvhIo4meCcnjvILbqftbulhk74pOZYVIbRFbHvM0EIS
z8FOfvvuYWTwW5sLBu4j5pSuTynkiF1tVjLvYI70VP0WpujZlpFtnlza0Jy7imtq
5X1X7af2f2di6G8YP2LujYOecnf0vytTXEpLBjy5l5LI/LkDS2S/+UEFV5Ydz9cI
4wqcx9F96Z6y2jy49l8+zSVjiXQnkdRKUGUwCmi8FXuWbkWOBJuZqUnIEIzITs0z
sHZ/b7uLY3kkHE6KI0yQGxFdbiTZvmrf1KHkfaochwbxMmHiR8k0s0MQ7jGOq7VL
USEhq+ACZLeD4EPqeKgPMfT4uJGUnWauyKDLDXVyP+Az+slTE/JJJPS4jrNEbh4Z
vl+LHbadxr/FeijmC3UU/OqO1FqSEFn/c48JPbGRkSuetrPXfYCb85LZjqtVSUH1
6Fj0hi1gH4ZP2uDIdvhtVo39//23S6f6gC91Us4n13cP59gkRJzIufgCGXTjn1zA
VbOWDOAH1PA7GW7eeGi2SA0GFMgByAAM/x9hUnWaeybnbCwyZOmQZqUBv8UwiuGw
WdWg1sgKZEkDaXt8bpYZQLGF9296LX7ELPgeDLIKhs8G/6/bA8pltKBlGc/RU2Zo
M5H4/UE/tQSpaysDJL4vbwgDwTqwmkBEiFa1Luc08SKBJ43NAKY0sy/Wfd42FKpl
+ZsZTIwnLS+qzq5NrxcIq41wPX/40o88sEIBI61Xt5NJiLCRaK5zqlIB4cZ4IUAB
qq0rAFkRJU+CUbi9dsI0GYcjZUF9rrAA4ayJr9/Cg9eGPsfPH5A4STXq4EJICMUX
5k+G7lLJki7ECyWlDQWHCpWndnq07BZq1TicXnVv8yZVqXSDOkDUUvdD4PMlCE/K
IYkjH1BLadR4RDbxvPkyA+AtazDoPhu0c6kyItFVWiMxjlVGaHKV8aiFRGoEiZ+f
9A/w311ioArmzmH849XwYEs0IfD9yZuiqwYhmwEpI4oZ/QuYkht6QcAAKQhFTdqr
I64zeJRQRRvpnUin6XqOvO629FszKpbsJJgG1N4Xwr5MrnyaHgta5sTzPIBhd9RH
Y7C8cqBh2zLCrj++ksnb6D1dAT+0aq693PpsBJP0BEZbcs2ybsqRWSjReRlIftq1
VKfDywlphNovTZwb1pBW+G2n1rV0pqSV0TZY34wDpDR1f2XYVQaXMqfgV5Ifc2FO
20MRjDN0h7qpTNTd/XUPX3Wc/vjaAA4qbXbkp0tquNFIo4EhjXs4iic2RjRT7U+s
Tu5zCKN9ZTxQ4ry5yav/OA/mBj86mekExE/wCMYNCdTSf2REXne29AqgPlyIXTkB
YTHzUdT0VOv1fKnIr8PuYJm3f5JVW10/uVr0/U/wDfgSC0lsrfeU9pKOpSHROQW9
Kj/VIeVg2PoKRSqiph9sfHTsoCetF7wm9yDo7OlTerEcoXpQPGKLR7IE56pX1O/G
0uDJI5v48lcb4QUuVExcJsqTgdoycLk5XjPbY9KfDtOlfj2F4PrSLCKAtVTJ3Ech
2jYBfHSmApOzUtKQQU++t8o4tNIB3BCsgGXmjWmIhJEERkN+N1s3xqaLCZbVAfeG
kZU1o2NJa+1U7bx/gqwyqUoiuHV9HY/Avf9tqOmtuHOLNr/H7NAPHSpPBba4myJn
i/XVpJLYoMx7rlkOKs6UTuMEd9D71AzJR+olNKs+iMeA5rHmfc6rcr7rGi3rtO90
g5MznxrEjgsni25xfCOF4OvYKp/jgOOUiDTFNDkM3erzqQd7LEWcBlkYAq1X7YtE
8hGNRN0sH19GDVAyp8F5Qn6CLhkX18uEP5Z6ddeM7vJItp99GxJNc3MpZR3xXfZI
b89INbkFt1B9rJB/Jns3vNn5J3BPGd6bPVb6JyNDBe67M059jdmD/Kout4nQQnVj
iKXoVElRNxpkThUL/ctPygjk8ZSkNlKmrx6vhSH9sqeOhqqFs6kQw1v/T0m9Dj+f
4UOKLtvM/HSs+XbtSLZ7aYNI4JhN8TRjAfR5K0CGBxmXFqywHA9d+CD+AMitGMZ0
SmfjwkaXtlWoAiqv66MIcLklsWBdUAtE/nIHMaucwbxyQbCaSQHPcRW4lb0bGBFg
xZJKe8rdLcF4oSmRC8SKcIPsVm338safditSvQVDm+/xonhT0L5nvtBuynDin2oX
vf1iXxaadRp08NXjP1Hie69aoHvsqS34og3n3R+PUX5mh4KuYAPzhs7no5wzPOUp
ZAXGwVnp7ew/xOB+Xf2iZtSZ6CEfiOefEmYwtnE3FK1AK91ip5s8Ak2eD7dVJcUU
gktscwIvEfY55YUjPFsvgx6q45UtYnwsqri9O1PtLfG1XARP6BRYT+53SRWDZSU9
b0FbGpWEf/A7h4ZZSJqP29hlyiBxZ3J6q7gCE5vBxnE6UVy13iye+ULDm1fT+UTS
O3z3fyEOfBiGhuxP+wMwuqxbQODOXpLBnkwKRSx5AeJzCvfnKzAfU5K4JNnZG36Y
xX9W0LSSKpJJQ2DWCo9LYlZc3sg/84UWWH4gL4F3qocNNTFdxHNdVZVXSULdqzrO
XilQrCBy37rlijrWEJM/Ui6dnwaJHBzUpSnTRF3nQUJ2/G5AcbQUCneFvit0te9S
VXAPvnguMPJ3XNwSaQZ3izdWS77kddPkaztRhSPJ4m96fVjweSxgveEAl+IhwWNr
dPzqr7oIM887TD7755YYQvWZjMcQPfMcJB4wJv8/IFsiB/VhTAHuNa+7PspRYGdP
VK+Oa78LLXbowoo5SMmL3apEdjoz8OHi/0Ay9qtUiM3nPQiFBVFlAGR6jE3Gr5E0
j0XurTPMWQWVmaDWon5rxQRPDFKcSOHOzfNnJrCnDI4WakyLyN1ISmjaQxNSNtBj
N1RP/tInei789f2QUFTWM5cbxftPtxuKegfupkqPqW41VqjzNVh/gesOJv3zmWRf
iMsIToYRaZixepULOjPiVHiTEt3JVgYWxfIW50fg3gr27wB1h+z3yQD+Ffq8jxic
iawjn6i/No31RGsnC4xuxxTz/7GL1hGAjxXwZ/Cui65MGfj94UweBdd6K+D6QaJ5
rpSjogOeoH6vImtBjyo/hLCcKiZl3a7xPbEjr/Usoip0YUmrz2UYVeEpmw133XjU
VQzarl49jfFhI8H4K/2YfzGj38YD9ZiJ5wuRcM/ky0hhHevjvAjIbxgXGmvRluKI
sLFc2b9pWph6Qq7JjlFzBqBY41P4GZxkxAp4gkC392eXtLmDMwK5mknMfnFiwNMv
lUh1Fhn9ZY2jIlB5LiJGak/TsX7fz54TgkWaJKmp/Tf7QpLV5dlCAEvwY2iwooza
AYe+kZ/DdQyConIJLrSL8AJBECdPP+Pn4H0QmgLrW8zz74d5XlyXAoM0TIIs5Xr1
QlanS2zTbUsBtVvKb1b+63eMQkOJVxYMtjcBbfd9/CSG+0Rvz0x4kjM+CJMeYnJM
lWJGvjT21lEiD/dzDyLZ9M3Z5lm7+ecZCoMp1hVVlundTny2vvJSTdPcvN3EjBbk
ySTGXZQHIRKrkXpeRk0zwRJ9z1X2rQCW4LCXJg+ClfqMFSojpXL/1pDZGRra4S+0
0c/BIQ8f39KLZR5R0JW8f/vutdtW06uq7EQ8Z5aHs4Na/3pgF20VKcuDzzdZE5yQ
Pq1uS2ScoyojjFgd3KPWEpEb+L5iNtJNNdSW3de9mOL7TUAIFWI5TKuKIj2zO6jo
unUJJMHZYaiSj39Rtv50UXCtZdEnbzXoDL9ze1RhuOxwIyJNRNhhvpNMKBxNmt0W
bTMZsCUS5EIspp3VA65IkAqECg9LQnrZ5LkRdOx54ihITam6Arse5hdyT05fD5Gc
HB0aQZiL6paoZ4e7594ZMlZKPDpSVYxTru9a28mrGvVTg+ozyaSYYxzhvoIcHKIq
+i424X+QI9/Ip0Vn/vtrRFjSsg1Z/w/rt0nfAtZaJ+8kAbpePwTMEHUsaFqFJxBl
a2U6xYB222khR717nWHma84Mdacu/XdENjsllbqaRzHKUL/O/cBhffXSVCExCKLM
bpMyTtdPOSMpoy2v9dlhA6k6zj0rleqluvtAPmupfq2Wa7o6TD3YjlA2euzl9NKW
bVWfME+AScnW/lteTDO6PGAOYbelihjnyqjhGT8HZnwDC+vCtgNMvtXEfDAzhmZS
BTvd/BPVl42j9PkFsm2HhtWdqOvIeRxYdDU5/JlCFmTWPTWLBwKBYiq8vKdMwUKH
D/I83fPuCdC3dPjQfJ8G+c6RGbfGRZJPBz1ol+NHjPnFVau0uTwXQl0m85vH9yBK
rQ8vt5NCZOYNLm51bF0M42a2N6+daGD3s9p/qc30168+wevvtbdZPqrUOEix6kBJ
G7j42QGBPK4mJsPOGOjGYREjt/LZJIkazjbNbtxxFugYhXo+DemdWDfZZN/YbFWl
Nrb/74frzRnojyd4Zp0jtd136m8496ZxSu0rtNaSl0FukqlwkmwQTJPDEq0vfeqK
lUt2w0FdHFY9GCIu0qaFFqjLmaHRMe5mGIbgywpTmbSqFph6NaWJV7JZzqVoGUs6
LIWRvysvGgS6J/BTprPBAO69oyJGHhyyUgBRkR5yyZ5VSOtXbS0QfpCdH+ICoxaX
vEnIdLF3pOq3Y3/fFhsFIO21gSQLnr1m8xzvLfOWRusRkbxgsvcAlqf9wLLGXlEl
Y/ryS+n3saEGSHMEJFSBKT4zXK7uqAlSkzipybzTKZ8fp2jJoN8SRVwFymd3zy+o
6xOX5NE+8mShP//2LhakLwNrRei4SVlIVb4mVxnz46W6KvoMHdMxf4Wj0huZHC+6
h/ygnQowP9C6qE3GjYD0tct79Xc+hZkZqhZXixNKLq99JB3S+WDKN/HrujpPggtE
Y8MMu+Hypj0e2CK55svUQ7I1WB/2FqEe6yFZLX4IgSVpoFuCSaSGMQeEKu4S0uvy
2SelXVxvU6VCJNO9vfzyst5MfHG2Zb4A6kxEevUm656K0mloHckCRhYo/cqMTpm3
ImLwVHTP3Fn/jAbPVTIZQTSqZDLOdnLEdzqQ4C+Kt1KrCcFEqwDxToVTSLMjPmWw
QR1gVmmIwqQf2iHSclvtP8ge+Eta91zSIuUdRFCvi7KcIBzFljX9FWur6/Q/wLLy
+tE6vXrz5T+ag4FTX3rslzLgFJJLWcYSaOvPbMQkfc7hoqkeAVHFf7jFUVfYqzJ8
8VYgz9pNYoFCprSNOaqGWk0j2+aG775bDveQVQZIn0+fCf8JIjCZ2ahmCiVdmFKc
38Yau2hPNAQ+DckiKbFy2IjYAUTPyDMb6E1/IW+Jwqdg/kmAxSEtla3y1iSMeACx
pFZnZsboqX7o7IjMCPLkZrbMSFmC96T5DLIBlXuW5pn8OpsK78Wb1arQFtLLG8Yy
3D1ctS1D0v762uh3TsKV3FkXGjIMZzyUIH9ny3oTq3KLdP7hf4OReVuHS4PViHKa
7zklKVFpdXmpAdErLMh0JA2Daisur0YRJOZf1LSlwCsAhORwW0mWvanKk4Nl+b1u
BdbPKhsylfjAjvop7JiTgh/+6aGauQa2rppgW2wri9eKvPgM53tbriN7LRBi90wC
K3Q8lyHnIII3EKOsajJVm5hflLXzC12HSyI8A4NwqGf0isVNxOyyIpzp3ieIvsJq
hzfbkJlKzl8sWBU3ZliV6XRNIGHtoyt2JHqJ4I1zYAKXf8xsHHw9z8zZWCpx57pa
9anpA1qeMOXQ0ktsj4Pa2Mqa5qUVuUbPmMHIsqtyLZPdghhTFrW5XJtD8uhxpk3K
glhGDOML2jsO8QBy1M5wXo1uB3/Tabolf8E4DFZJRapNYEzLbtghtslOfgrtuxPh
QlJzkX3Q2CKs9MMgzBseqTFQGN90lyqQtWxjwRirTMXUtLx8b2TlG3fMJ9tE96zc
+ReS/ZXsLuuXIxlw++UYyTuH5B3sDlPZl+KnGpWA5rzsAp20nQiMVqdmj1Py+byF
klY1LdRLKRfazYM3IE0Q7DpZWpf6C4v3T+1/VYLvHsJzI2r7g9XEokzcywOZVZKq
Nut2EHph+GblkCnBgiY8aPyFx/fdQBW521yc6f2kXawk6a0XOB8vZz85nIAMe+Zg
7SEj5C/slKkOfl2JTZsw7BWpuD4dkbKajV3r2ugH3KNeC5NoNrnyCCYq3j2oXY+7
aqYhPjszuzBAldtVkp2xDRtWmKKMwxNd3hNg5YbkGENDJ6C8oUAp3R5oxBdcytfI
06SAEAXKAq3qU8IHDw4tfj8oxzAyyS18b/DhT8OqAlEo66na2rUNBd8Mqy6WX/QP
xBF1g1knO7QhXjRuSXF2u7ex42xIjyucETnv+riPS15RwRg22s6YJPtIGarkPlp5
dHse32uwVCBUUkBwk7ilX68tYQ2NaXbZNCIOhpiUQx9j8zvX0A/i5xAIi+HSnlxr
c05qluBTIQXT9C9/6sp6Vm2YY5MGV6SChnfNTUTg08+xs34R58j+XhF1zPvmCQCP
Ny/4R46Lvx4gKym3elbF6m01rCyUEwXFjK7Wmy+KupWr989y4gX0a3nKA1BALPwC
FnXZCtIcBI9nuwjQE03gMzvMHUtpjZorQ4tShcCuUabmv68fHo2A8MCWxi+pPvG+
pZje9d/IoTGiLwB3s0RoeZEMoK9uX229rYnwr2X3Sf1RhXNLGygKZ2iR5sTj7b5f
s+u5GoDDiXNCvkKOrDWHgqCgRhMBb7ePSMvSOhJiWKniMxNw+y5HrQl+8kVm2udD
rvRsCTA/y3BcllqTaG1CT/nhlHqTjp3YNvFah6nG3JfshxDha2vdIlS7dAkAe1hc
SYUW6Y0mUuoS8zZuyM6ZUc/k8X+YW1JsdTrt+/WcftfQNDe2QIizUnyIlXY+8qf7
LwVYB9wzSpM3S/v495eRNWChsSFfIbEw7lRxl+hmjC/kWCsQFdns/eNNY3uX/kaO
SUOM+6AJ54b8bUG3wV4Y1idxTL2PQQyvdC8X8chqIklzDaRWnXmVGV9VV9ZAVPs5
IxPrwy9Vn5FiKX/208OeKmlusCWq1GnzzbYyy3Wgznr0BK+PVElbzVTOcZcZRBa7
bBxyUpt0OO480krFn1kVW7bAXCDhwhf8A9qRKE5Ug8lQcx2B98rdcpcOvOs4Gr2b
SBYro5fsJg81SeRX8xB4Xc6KZ9CcKMOuubmvWdn2Pz4cbMPXGkRkvKFQxvJQFVK8
hpcXJiAx0PlyH7zkR290tQyWUYtYuaFF7CpCpKFExtCUnDrEowoJIVvr2bNC7lEl
mFXUevBiZJVsmxGO0xV7BWIdkGrnXBhIxHjbdKIMaawJAKPxVxvNHT7NVdHv7QMT
ju0OxS+5K+Exgajt+1URoCa+Lfoqvp6I7vXM1NhEaXJa6wpCYY0FAQitEWx1ls86
WSu5QLStlquXbUpC+srA3ypgoY3UNM9LGO7fBrI1MLQ0ZOz0zSuHaqwkgmGpWPMz
OCXdWzv+0DD8V727X07Tjw57XQBOBtnVnsBvDOPBlXu7BhcE/XAKeUihvQXm79oA
sVrlOWE1AZ1BQN7FaNSMXzVezRry+2Gu/ettikIhdAi7oSFrXHsL8lNcOpyC4PYl
5WXKkWy+VxHABkzCq1tl9DrlXxuavsDCAwcKmuyCBybrirTUHkN/2pNyqwB1XJM2
LQO79aKdvGtl11gBL3ZUoUCqB1vEtirkxClvbj/IbCb8jSGrLgSlljU3ZdylBRw4
/BsdOr28h6bTc7+TTKIor3Y97LnOWuEOoEiaKTPeLW/HPqAeA8rNgnhRjPrwhA5G
5O9IX+kbSgHSy3aCAsEQvVxyIe+ndtYjOen+i2Y8f8WuDMJ8aq0WFL8mNvACD2fJ
lIp5d+ijE6Uz7iUsDNSKooZzcvF4OxrlPBC2SJEPSa20YJXkLzCUwwi2F2jvJLbt
aMSLVNw8pvUJWhBr81kBR+pWg0b8qCJtY/zeoSYDOmJz+h1Y1HL+HwH3hhOMnU07
ALHESqNGyKgpI2aZf1aJ/Qzl+ma7Ko8hzk8Av5dTDQ7i2nZOQMhYE+zieTkgH6Mr
6C4Fg49QK3zMA49J3rSTLCSjsAUqdqmOki5eMkXOPwjohpt8hX9dPO3knTabwDMB
uG/nWZ72+dOrWhep8nDlN0YUkBFFTfrpS0ny3GH5z9dPmkgv5ZfUPCLT/+zXBogf
OAe8R+k4LU2j1/guOxoKcI8nWxmYyA7qO/C7gXRTH3y1MvMqHJUpjXtRgdfpuaiO
FAu2MgmseDaPpbBtw4aLZMEmHK6vcphgnwylQGXEXl7HGkX3fN8OfSRRM4AeMolS
4sBVjZTx5Ih6deTxZPfGd2dbtB7WPusNZNiO1VN9FuDIW7GqfFmDjvynOhEirOcv
0hXTNUGAGWaTgeWr0SCnvQtBVZR1a4i0/cTX/dxXWg56LUuDaJavNrj56cvKQeUn
M8AQeye614+5InJfcZZ/Qv4MMZLICRk0Wbt1GIOvRjWDPFpNE7JdIFITKkoMKimQ
T6DxnHNyCzAcxgfFwwqmcHvuGFDuid3gXcN3wERYaI9zMMQfOQOSxLxE6fkkaywS
6VLh6yoZZGx5x2mFEdGfbAiCh1t0nTxUNq1joPegBVZgkMbdZr6h7wP7e4anp/fh
Ho/5LfM4+7mEMlZr1GnptPLAWo2a7tFsGM95biuTPAEtf3A/Gc9feAL7MU+mpO0d
k7rFSTi8UiM1I536TCMEiso0L2jTD+r8+e/uUKhdxNkW3dWGeloU6ySgYd/aTDMY
AxYe7jw41m9JbEIwk3cEs7FkbyPZk+1Lb4TRXgCuk/u+mh7ZAT4pFQVkXWGQmArm
PJFX4qEZ71Oaz6wjOKqKmWMkQKEF1JR1toClfVucivzgI4SV8UctCFrBgsXRvJjC
7wtkeeVB2ISWmflJjT8q9ELX31Q2eh/Ajlwg1SOKfpi+B56CFZR3UBm2q7BEPLcZ
mfN6HtUmt1NOsdiAnYwXpOMpDSopUWeyEy6dGbixLwvSDUG0WghlnOWSe+mybyfP
2XQzpEylfSAhlXdggf96yFsCmn6P2eE0PFOqqBC25OUwzVC2b9JuRuttBY7V06Hr
K2HV4Zxx36nfUBqcf3tLam2DSEgNfyppGa+yMSZaBEXdkakC3Gt+K1wxfplcu2GA
XlR5OWYrq00ThTDIDGpUqfBZwBsvC+ldXWQvN8SSOoOJEYK2gnf6QcdqDdPNgPaG
W9Xm8qYs0SQjwzaZBd8WCYybQrhjPykxd47dbxefVuwNrlSQpJhNUNg2XoHLZe/3
enTuNNiQaGkO6NUc6e425EE7qJUnwC4IfyVqY7ZF4gZilz1Zj0djK/4DDDrswbPX
eTvdLOFKCSmAfOTit+L6i/IzkwTuigEeUzBK7R/65wpeD7OM5mEL95O53E1oETYe
laBYN4C0GOaa5YEGBagneKncBi4Rrmb+wENg2/GWiyrLuUDBpBd+GzdnHsjtOIER
yen8Y6lUVIDQhvFyMeeDjp5ANIRohxkfvDqdfoC8ccbNy3ab+EzYsLxkM30TjokR
WSBLftFXderr40au7wQBnPfaq0snOIY+hv/QGNRbZofLNOYyvWLoJ+GnHjbcwHnV
HpfcRNx048L/d2xXCbX7Cwn9Ru9lp0QL5kyeWmoaKqis23AbEemUb2ys2Vfq70dt
GASEhegWRbacr+W1DYRWkZmRzGUhVz+skRJH6ykScT63dTqeEYPfsW+P2n7Xi81o
srOt7qLDdknQ4//4VTTg3DzSTKZo5tv/so/jI2f7wsXkBDX5p+61c/AlbWx8vscb
LzbfmLXmP3doNYzUFRH0wY4SKA4CFMYcJINU0GFU2i/uDhMsLYTa9YJJkkAMcTmP
Innr+DGrARV+bhk8hTJQl6D6jD+AdKLXxFUQv7rSpssUTU2fZu1MjqH03f0L5S4W
Zt+9nZlLIcgYK3T5f8dSmiRBJHSQjed5pLWxkOA8CIxQwNUQocKcN8J2PQFSY7aP
hIxZACkKwz6AA3DvmzO0frXCCLVvHel8j0qOvIVjO55N/8kqIJlGIA2wZ+H/vy/T
xLsOezzM+KNEBW4PQf5xgq7iDCv6HD7pYsPxPlT8FhZ19tDd6beo7zqOsY9mhrl3
D1FCKL0/sAEW0cE29MoEcrqxNxR3IbJmLv39pawKD+g7i+EwIXuiXclj7ItnbNxd
7/8vHNnVL03ac/5o7D1trViauB7LZFPIajJLt8RXc6wdg+XKmjQDwsbNsE1AxtRb
EoMzdlM+dUQrRtqlwTyS/gySlDCfT4ODkQD4wkfOEdihxRBGk0erNPqxzJ2CO+Gx
YrmABb6o+UYisDUz2x7fvTk/SP9C+8kkQCWh7lrexBG+yS8nG8jbPtVaiz6xipAs
NTnpM5jSwDsPqep+14YGMGLHwHk1RTn5w1BLavECUdI87mBtMTgX8pCKXS/qJAiI
9xYDYsgcIfXgqDJ9ebFD30uzEqiaSYkbakgDjIx9Ed/1iQcIbPt19zyx5uJNvkUp
/+Ky7hlh6C9tosXQw7irmXb4hUxqnnJn0ED6bM9fRrAgYG+PNwPj0C0dkdEIJzik
Du0xG7+oziwNDe3gpvXUTQDurG49R2Drc5e8wq3iDr6gxOfdzbBPUtQzL6Mksf2E
O0GMSv9DtbKKsOORg3CzRlM3iZPDXHuNe9E+8w97VImsqz25vIEN/DN/wRKXzNgC
nUKRUrpLlkkV84xeT8nIRb2O4PmzEAlONCKpIJPX3IeD4Z8WvYzZMYnd9wNSd68Y
L2HNcIxZDl15g5b/lM45KWI4cGAyMDVkKUkhFJejypAW2eL979lLaCJ1EKb2dNns
IvZyi0YGp9404cJuiG5EKsp0vJCYI55XFx+YhwkPq+8xQasDQLEq0YGQGvzJZM5s
wzBMd3J4GSfIa95Tcjmsb3yepdT+KaH7B7GPaj0J1NOPgw/rszkN7ngQs/qbHs5F
+07VmOsC8LNd1bO+xxfVLWznD3y5ix9LjRoiZgaigjqJqTV/PbdLbw8JErQFwR8/
puNDguFEk3nXoFaAEs9592qK8PyXaWng3OKJgGwL31IC80QsLb/0PajVBGt4LvvV
VuOGwmuz9ifaW0KsBZSZrnPlk7K0fBnaQqK+4VSBUmwJq3yl2QVJLAmSvttRLMFd
B9K8RKfOpKERQFvpuWfHe0/BnMEQAPD5/Xw/PvaugZVBwlxMJRZxg4XdP/LGW2lG
8fwYojVIGpjnupnu4pMmaaHvOAnkCJxDDJv/KdXfkp2kfIzPVwpJY0Ognlq50zO3
gOUJsc14nvJGO7NZkYdfJvIWI5oInDCr4mj7CiF3dHHoptdfKLB2fimWMSk91EA9
UWh5mQFTmsODgJCbM0Tj7LORyNHW86cAL4w7RDnunoD3q06uEyHwSpN3T7nRmK24
2HyfNv9Jlc/VHI6p8CsUjbH884zv3qRH0IdNXT/Q8XFvT+P1J81SqKGCtvPrez4M
e2nmGLi5d5FGkwMnbo4EUCS17O7YSbVkE8frCUwDqaP8GAajddVIk2gir4Z7g07b
UAFUECyYKpOMe82rz1GS5UzKwRTBL+G5R6dLIGElGM7Cn9dbpm171tBfxZpKaC6w
krP7U8K9OXTpAec8ZwWi6aqTsTkjcrNa9fOtag8qItbZlzYF2K4Lh3GA0vAZ3xxY
F+jt2uQF+p/HVR7pimIeToU+fokuTKKlQJrCHf69kNDF4tS8WjLOJg9whYfaEfB+
cwoEnT2FSpL+udo6GySHku3YAG9pw+5h+6e0oY3uHtlLay6dhzI06riJiR8V7EH0
BYuZsl90ptq3lq0dK/NK0qEAOTpq7UwptvOf0cjWDEfbIjsYeuFNvIwag63Lrmqt
DXcPL8YMcmB16+zmpIrIBGpADeA/tkM6XUzGiOrA1Mk3nS7lxFY+D4t7sRhI0crS
Djdww2Lj+Icnl9Zi4qR3RptuplvTkNB4kkJ64LQYz5P8+KxdubJ1YWUZ7NA5685s
gol/Htatl6wtyx+99YQVNZnwGHpONQJ+SiAZHN+/yc826HBJzXjz0hvqoGQlrDAP
OEVSNHQYHViG5ocVKhV/TQNO1mQ7OF63a/y6vLIkOPpJZzxDwYImjrT0XZOAAIIy
qrgjD8wF9MtecMruf5ZjTrGJzTJSHGE/B4rSu9CKfJNhkP0skAV+JdspgZ43HL3O
n0GZWoCljlcpcX2gy+0oZfO7+JxUkAMjzgXLlhwkmcFDF394OMp/WpKJUP85Ur/l
rflQ2f79nbRHC4yHGH6ooD7zDYRoT0jmnsMa7BufWIOVgW4KtEGq4BsqNFH7UWeR
WkDsLi8VCCpLfYwPc2nRmCQkd0LwKWawkCiYYPUKpc7jrB4oyb8KaKxy2h9pRHnn
x5WjX96rMG8cAOkSzHXctM7UTlmbkIz02x2J/Bh/X4Wn0o4VdJvGP8GPpq/GPm0f
c3b0Ata2lAxTaOiRz85IKKb/DwAiSMnrnpr0u0PnVKcesoWcmZOlinTmR6mKqKMN
mLmHtp/a1zAJygAyLrxYEQBSzQqF9rx8g0LOL72L/JL8VAh29EsyWSahQW01XOlD
hHB3a6xQ+Pgn/CqmHXxUDTGKMVbKRY1R10SzeazD08yWHuYxz402u4pIXFyb3Jiq
1tgybJzedZUhooLcOWYRK4peeJf6JW8SoZSKrMMYofF3h/2FhEfP62JKM7eCmcbz
Lx/EQMz6SmRE33igOdPTYaLXhH/1ONJy2cj0mmQe2EgOikE5W2BWO50Fiyb1BmVg
L1XpWPqCVNpJYMR8cHtg7lNYCX+bcigDI+MdA9P/bbHMykKrKMXKX18H0IPVK2Ws
/BiKofe1tSn8GrN9o/qlHoYHqcAIqJnmxRlsDsr+0aPIlrVXWsck6pQGU/g9FVnd
mSwfbmGJSmuXFILI269ugF3ewmZdtZmzrTb511Wj/Yr6NWLUln5jO+aPeBMCeqIO
HXtZnwTunysKtqmilgbPs47dpseUZuRGHcc26rm839nyssioz69D4S8DgKyfrY5H
xcPJ0SUtn27aO0PhD5mtp7o5vrX0rSd1ItFq/RPxDiUqSGnW0kQmwYVWvtb4++KK
aq1MoQ5a2nyOZBwYIDnIikgL2mqrFMa8Bwa79eiPaT4RhWQGq4lPPKtXr8GSCITu
tKGQ81EDf85vZrV/kSPsdwIauD+M7/ojK8pwpLsd9FHh1JJCTjRDEmmDLdzKS30L
03zgk0OiYYgcqN9JJ4KFlwrjkkc/JjE1Ztym6SJ0ZRZoDrBAJQyHBOCFfjaCZZ6v
6GG4e6BGJjUC00TgWS+6ZxnOUA/TcBQsHSi9nceWkZCopTnNqxqZxa4BBv92qa1X
qw3ie4jO92YUNH2ogh8sSYwOoFW+vT/Ff9Z8Q+5nSN0l6pK8U5gbU8SR+P9f/fHu
8XJDL2h3obf28zKymtqdd7WFxt1lhEH7vQ13W7RwAonfJsBAfDm+cutC6cEmZUuE
WHZ+NaUpXfiQH4GSM3GBv8i6FkM8s4/ewmqszhEbSPrRFjdgKmkNPiRUi1UasBEu
TIxnoAIwmwPN2Hf6hyMb6uvZKzVTOmgm23+A4FWuFsRjiL7sePQ/cNmPTDOw3uRP
0HOszkViXXArvfogu1bGJ6xMxFOXOv3z4gB9GWvWvlWjqp4ET2GWsxaFctdJUi3T
8z/O079y6YkLS+jfJvpyqiGnqmHJaF1G++JnKUx3S/WHmuSHM1aSKBOrOgwBa897
rn6XmrtrtULKue9vbDA/lWkBAhNWbmSzq4vr3SXQm0JFhdXClVxbVVdZe0szez+9
9CyPuFuUzm2g9qyMECnWmXlNrkhoukx6NFzBcwhsLfk4BD594aWI7P8TxLXr+WCx
AynGZXEiSZ+FP+Pj135Op+6cZ4kA/T6QXG8qwIeH42n4V2wjoBoYsuoUd47PnsJU
vAMcojYSE69PWLjrlIN39VC5Q0wI+ybcypk8fV9jWibVQXpTKhlrSeBHpL5NKNfo
PXOYtxe/o+snwVA0/GYFGWNhWXiYb3bVJ0kl9KmiPOpvChjEZTcZCRqDEGuVqqNX
A6FAfHmOfXspgWnJzVkN0D5BNpIeqUxWUT2wRqabCfTt1XxySMTwTLG5qWYheeo+
m/k+naBGOxIT1q97qWUj3bowUsaNekTu0ZCgs8/5zLFevFgSyCFtsIKpoPSDsmGI
0ndt4aKb4FoPA+wo1neoBs54yagZIyX/JElChVuQIJsIitwjYl0xHoS7soL4PkM5
ul81lfpzWdJkvPOcBEPHvFcUXbw3C0IbqC/J4A0n6BGvjXSo+Zr5dXexRaq1wTsU
96E7QW3Hl2XxTulznM52xvnq5KXYPT3Fj6qTSgXq4lQC+52Uta+5WVNbhJPgmqeO
rbNyoHaQxqmlSgFkprB2yvS2TSScpk5+gCBh8NxNg4fwxyzLPUq1ogzNp9Rngumn
3lSaTIrNMWuGvw2eKJFpeqsOl7685tY8yxks0s2RbBwwUU8NnKEufVYARHX+Sp4C
pSsj77DcoUju8QeXJqCelbgMRqXbGBeuUa4yCpQ0fAdBxVJH0VL/GrQiOGNtyWoA
tPYWo1I7QxpRs09JLJnrfyKQtBmVEtk9GzLliMS9357k4cy0yRXFN3n8F0XrTgfM
rfRbGqkWtWFpg2Lpktv32S20XuMBYIB6sOXnP5s0+6RHINtr0Je6sxzQoKFaZIUh
XI4WTQ8lcjlJRwIc6Qex3WWLIXccv6UwFnR6UtX/yqTimmOFTAqKBv8L8PajlWpq
tLCtpBanmQhgUZJCA34aqraNF/iEKOzt76HImpkuq4BV1S4qxJuJxchYH3+6JwpD
ngRWWKtFXC1faIzP6q91vwXmK9HaMP0PE4hfU495g8YnDh3ysLaV2549iOESv54v
EXJtmA8CmhMAhrDehtQkZz2mMB72PguTEiWHTZo5eSJKS5eVcYMFs7/yFe6vpFA/
zcLx6B/tfBZ+wW08+kM5ANps8qpeDLM+36bB7EsLMlNdn6FzJ8ZkmV3vWLnilS8F
fQUI8T0GuPCsCQRl1JWNDe+LL3JfTqgDuN2HGdkey0SFPVuQyKattANA7l3YDYDf
cGlTjuueGx8yyDglV3bcGbGVq5VqO0sNfnPXgXGP4f+juXcUP1BNFrALb1KDH4yP
Jd+Qqal80ayAmYnrBuIvS8WJ9FqTjbi7MHpreWdgtbMky0QtdXKMIdYdMO6pLSAL
hPP4SR4xpEAuCL3sxsOWkkJos8E28mkehGIrQjzrKWu4g+P7Je9MHRXouVbd/pAR
nE75HFKPRSCEduz3C8rr19G7Db26MPkVIcW1f8NeeclpkH1BpJQfMV2L23pyIeJG
VrXZO7vmjGn+p0yfxZ+RVb8dgAbFqG3JgtsUStdaj4ZyLWpKvgHZjRqDEldKHpbp
/j9fAcZeFIZ6615BQ5J1gutatJ9EfKZrqcpB3aMDpa0qOBY177hwEhxQOAABZ/xf
3o4l5J+AiN4H09LbM5UCAKWPqfsCiX5VshvllEFYoN0DS3aa5of8JwIHBbKeXOPH
jwgbN0OuYwdWfdEV7MsbVq5UlhE+oh+YUnMgfwfKvkg8S3P5F1j2AQ9sm02fwHeF
AMCIdLlKOUqn2GKJSrgQ+5C1dsJ7vDksbnY69gqGeOtCNvgzn5yxVHH0LXUiCyhu
feHVRAMtF8pMcppzTY7gvz5Xe/XJStMSPNaCznja7hIM4oKT3Jj5RFjwz1vi21Ch
fbw0xP0t40ZIP1YcIDVO2hyREwZiJL5O1/ASNrRQ2ku1RaolWJF3vwLcjS3op1nE
9cMC+orGpBudkYOk1Qv4wlFJ63MZEEBBiAIefKJwQJl99KcggdHjkwGrNToQA8n2
xhqUPMP2Wk2XkvAdVNoOcRM7LBDNquVy+8Fj+c+MFdYqN/NZn7jLezE7t3FTKGtl
Kzygc1mdXK+Op4fBeC8vJCoIi4iQdIRKH5+WtMeo8N4N1Q7QDt5DR6P2V1MF+i4n
xkFe7Hmo0/io91ofVp9YrNhBSqlV2PTYy8yVXrV3IfTBCr3e9DiZ36pxexJ4m6yR
ZTiV5HYlfWeHhSpEM5Kyk11+5jeH0j495Up8+rLWfQvu03WBeOV3srDxpPR+06Za
KRfGLhW6geGZQJeOBWNWlHiDsf+U83U5YDPYynW2nx5qcTyXP2f7uEYmigVnKjv5
cL2spdDT03dQ/bqUrXEaWXPWYXRgq7Ls7E5w8aVm1hGCaUQ2JiOf7fRizGEDh9w2
CcPIiJOzvk4FghegJicfEBsAqMPDKudHCylBvA6PEe9y42hz3tZZWpo1/cxFEfg+
WrQlgL4Y1wmAsu//jftuT59o1Mmwru/BXHXypIS2oJ/fIqCq00wspatWL2Zt3INF
LSRdugK5d5XXOJCYNDMAivqDg8fiYufkbmjV9mJK9DJdhx3oOV+a8SvV9L0yhG4D
ABIyXYA/629rUxCJ5mWD8IaoTt8GkIhx9XQ1/k9hTqevAMonDsBnSTsGaM15qSkx
zuy5ysdp/xv3BOOLJQ/2s262OiD9amgczYgZd1k6i9pkkW9rZ9/94VENYleGxZka
IIcZ2YOtOnVHzkLl5Uo1cu9mlUpePGjcv51FoT2m6e1du4rkJVz7Mlj2SjhHzp3t
VDWz0jPWB9JJw4XCBvRew0Lhy1OtKwYiGKnvrLffnhieg4y1i2EouDJ3s7XHbjgT
QFpsh7fUF0VD1Sw2iygHbLbuv6SkxbAKzFKtHlf3IwAXZLM5bw/s5TEsV/wHZmsO
vtkslyZDQoH+dew9aasYd696LHUh4Ko6WZe6t8IyVNe9fizc8VMWi+jPXluGjj0h
u0IDBQt9Fzsoh+PDo5yce6NHFfdck2zbmIVciG0Ym5HNxd2xmifG6l0Z+bAv/Rkz
Ju6jPe4GoqC8V2bdoMrngiIgG4+Zdwfcv4dV3pq0WDczoMgXdClitGFvEHWRjR/Y
zp+3tcb9csgUuH0TAMTuKEOSTH45fb3d3vwGj2Mz3SEUneq/fcuKO3iEW9+VSUyK
kA+CEHxiH1kLJiul829JMLDGo+uSnAYAprxJk8CwL/7yqpC2nK6ArWDzZSZuk0ip
/EXZWs/denWkVKXbt43Y1zYrhqIR37Rf2IKlDniKwP7W+izpDkK1Zd/7DmnHMytC
x3HtEIUsWPgvg4G6ZmAH6xXWaoiA897Gy8rF/XecBBWArqgw9iEqDgkYftJUvDyl
NXbii9J9TS+LFJ1/qlkBk36EqtD7yMTcBx+WmA3bwdbFfHvAF+5pISnGyUP2cnR4
zFmIxDyhd+4xzVPH60T6MDC05dd5ho/gNLPNSc4z/JNvWQY26BErDzKAfsvlzrNc
qa1ialSvSKW3NHPjKbwgL1TIeiZfBfEaDOjt676CbeuJJyWUfT7MHmK0kL13v06o
nOLF3JLr2mYiNkIzMachG+9G0qZ/EFZXn4vQDtZXxeffmy6BlykXY5P5S1fI50WB
FT3CpxQ6Yj94Hy55lxnLk+nnKiQb0jlTeJjaWux33f5XIEZZUYGPeHW4pxJAXpeZ
2Gw5ukGegUqlSzUMkj8Hje9Kl7xzPlO4YOT7o9/MS+4j2fv90UV6fx5Rb+ad4I9E
HGI0w2CO6xT7higfjJA0ZGpx4sGiIK9kcIoHZ6MKZhfAwEmslgPMCGSPNtDcanEm
ckGrTLzU2uCDM80aZ4oJHJDc83bA9L0XUA/kk/NxhWGesJKF0yJukilpvRjl7rDl
ea0XcJL/fhS/ppNqLN9h/AKPkjcCz3fX2jK7brvShUcB/Fz8/DTkWOhabqcsmfxF
UORFgyc2/XXk+hpOat7F0iawf0C5hJD4p1rYlNXYFB6N6Oz0PK1MkspgrpiXAb3G
cFUHGE2AWMkKQP32uE62KsyIu/ph+lqQ6sIPjirxBTgBufGrlA1eqNz0yoZqq/w7
kufOY+crc26fNmo3ukBCplPyKLyJKtEWIvu+pc3KvYfN5A8+/Kwa0XzXSWCfnoAb
JPXdwwwnREnrKfCMzDACLB8MU+Wko9Qjr1BJMxKxSZ9e8uwyrD4U1jhJ96v8vmSN
t51tYK8vNChYPJxOUVW1pQHzxf6CAmzaEIgzURhEbdrAN/dyfDX357DuGW/zG6E+
xz6P/vHaQZUdK8N3idxvEpn9eHVz9sLSEwDiKB4e3ti+OvK7jRrvygoLNzjJ14w+
GlTZcq3nvIJ/0LZAeB+cm3GGrcFJT2nEipiU+mCxljcoJI8qh2E0MnxxCe6flR7j
WEu++AN1XSsKSDCoRTXTQi4ASOQCLeaFNNkx1lvDl7XAWQWlFquq6pCpmi05JDlk
nVw6uqK1H0oGWWKWrmMoYA72rQhbW1YRjRYnreRLQxsuBYIiqAKDqXq0nhDotPjk
E9VuO+Z1zW5Ao1hmBO3kCIi044SOObVlz4z2EwM3yvV75aZLvdVUq4+OkgAPslkz
kQ6l4qQotnXKrwAIaXANbBwPZSjm0epJSVlqKwN6nvDwAfMIZssDEtoU3mLvSmYR
kPzmQTyxC+QeA44JunhgnO7/BihU6ToljHEu1Q96nNE9NChmUd8BfOycKrVpWd1e
MgeDJwOvVMtoPp4V2+wVsZ7Bbbw2vNYKYGdCdB1hVwhuoA8DbHoRFQVb+PmfFgxZ
BKTSI4qaKdXX8N4g7nPIVXX8/65XnzR3B/w28oyQ6GGLdF0gcgQebW4LA7Jtxu8l
0RmXoD9p2/7ATky57NX+hHvjaWYteBAYy4We+F/q1t0I7OGXSmKEM2W38FKQ4mzC
Ut5RBSBC9MHkdvlHLVy345lSInBVXgoiDvf09o9NcWtVJ4YVgiEw/l9YIhZgjuuw
W2FrR96lYch913UbPAVX2kPbhbQjoRfxWlOg/grrLyD+itjken8380AQ41n8LAW3
tTs+2uhvI1Ad1sSc/Q+OM0ngpDKl8iVuGppdR2oKTdk/mxEF7CnNvy+RS8GX/IIX
qdnAbiZ5FzqNpY+zvNXum0TJAJAEVzIW2zrPuSAbZKwGy9jt+UoFbF8tdAfs7X0Q
U71wDogqGcXSKoDshpdX8iLjIKpiBDZG7pVy61kC1rCcIJ1aFxzsdl1rOpK8oTnK
Ikeozj/YX4F+zLZ2O45IL08eoH68ext2GYlJ0nBwYkOMmUl7tgXdAikP3Z1KWg2P
Be0guMJs3ADQ7lQrrTyxHMwDPsLPiDjvDDU+jddh6Grh7z8EosBO+U91lutAovdh
vH9uqLpv5BaCUSadA03roMCPZ/9Kl/s5SIa5xguMsx8UZqvytnNMeX6JkqkRRkeA
gkpWdrhNPYS7fwA1gOBkiNVXBZe0bpMBfTSOVnV7wMnlZp+3G/PId6ruoJ7CxBrx
egGVhXvRJRkLV3/m6s7LaCG4Ftvchd42NhcWdwPQNqiBBobE9CK6MAVhuZ/+7ARC
6Njwcx9oJgvjkA66bAKS91bhEqJ9OsF/o0kAzUYjLyXe1UB/1mKADRAWp7dhJHhd
O0FEwszW4aW6EZwCMhYfO+nAlc/VC4IIFZLn6q8/tfs/CZmjiOdDJjMRt27xfnO8
oMzf5MDuOdUEHOyiEkiGkumfHJQd7RVCMeHHqJWO3CAAOlSt8YjpYpl7SnmOtXn5
SD2hsVnt8cJSon+WppF7mja4OwvFfq1ftKty1cDsGJeTxVedjnkVdSmstfK/6VN2
p2pSQukkBugkbJCePHDNeNXEgP2yc5b5DCaDkYNWen082P8Lf5n6frYHBz0j7L49
Rg2057Eo1uZhmIWgaNItTDKzEO2Y2jieebNGdBliN3jy9HhWMqB0pdWNJnm4Ip33
0s6Jt4cOK0SkpGVTT4qIbmF9uAIsWBzlIIqp0EP40oiVDkZganuSustSYL79R8hP
4vvpFO9ArwQvuGC9m0w6jy1UKpLjmOcCbfveP0OjRe9bz6tHJ/+eIBQjocui1S+g
LOuGtDLIQGq1xtXfuwsD/cSao07cVDS/cxATbZpTRY2q/QyTZ5VfnLfUm9yhPh6V
49qaP3t2UZ8vwiMewFRR/lwSw6IIt+6Tj6pSaYJpQuAmluyslD4yUIhNXVMEyrvR
ZU730OYQndmZjJqNIn+3Ju9bGhHW+F82ZSWBoaFpKA05JiUmaIITjs6+Mo8ZDpdv
EKsM0ioytfKEZCSQ3t+tM3XncsdPt6OaTvxa2R1VJDmA3OKEdVu5WmlTzvjNhgIG
6VkkWddaW/0AtIY5+MceIImN4Q2yAl1p7YifSZ45uLg1U/XhI5EmTC2F3pmROfFo
uS5aPjBQyqQWzNIC2FiYKDz7muSrG1QqUlsaW1KsfHpaR3VRUG4UV4755L2UgFtt
2pR+VAe14Jf6z2G7VoRThUSuawP4soqBLPfcCeiiQdUR3lgwwjnzhcVJgZ0iljni
DwJ98Rdn1LIA2o47OCVB2BFzh2fO8ctRXLUrez5c1MfrCjErKYra7UA7Eliof0WW
f7nX67XSardAaMR0Cf00cn0O6HEoWVvGu6iefKItzaBskRqqHj2xrq7eQ0zBwlyT
y7WwzV+CsCtRbCow+QRaW/mhbTt75554JoeCysT9CxnK0vzPT2Ovcp7010q4gc24
YRN/pIxNMPecW/ze8c+iy0NRY4XSDXLNT6Zyf7M4AAVsxl8zViocRKr77Eqjzghw
e4uIyKt7B4VPXH8M66ZWIxW+H9yjnJirsl0Zz8XWY3klgbuvNfNuzsSCPUCE+Eic
URgoHkRO7VLy0mbW6LcIAF9R2JS0kwWQU1QhyHm0uQXSVLsPPSDCVQM9UUZVZ9Bb
kDphOJ+ojp8RtLqqJ656tukMXez2GODTh22ImneQrlDAmJkXDEhIk4Wz+2bue1N0
hLmEMpAWXTRbc0XeaRQfE5mw87aIlsIAtjKTg6K8TRq8ckKXRcMVOQZqw5dq7fsc
50ThYdxkPKWJusQ4OnlHICKJ9Ou2eu0OLrkhvwmY0jc4rl79l7ttk7w2/IVseuO6
ca9iaTckkxT57V8tBqjp56KoytyJ50//EVa1Ia/+BGFcISmiPyw3qB2/LltfBmCz
IsQNCPSJkfh7tmZcbnDa3cL/5hO6SRFy0jzwGxFQngVN4qwLNsCbJuIe2QL+M5OG
uh4rQGXBjME5O5g82mDsQSDJwnA6jDJvdQlQ2vcn+zuvlTsz5PxXXqxn9qOCdjse
tsIlB+qV9PeigJFhVGrmDU3cT22QW/lzYPWGWuJI3hpkkPbNCNHDOk4b/S8cO1ha
/gB0M78ro6Jtb97zDLDbessHU30p4rnDTd/CksCODZYlq611iyfwCBte15ns7zoT
iaK5s83bmfw5Kr9RBMNOPhluHS+v+jCG1iUqKeZNM0soicj04ONifbZfQh3vkqkT
LxhW76deo7YttNcjICjUuXwJ/aynTnpFMCNwC6bKReDR1b1YvyY98XIrzEqc7df5
+g5WK+DuP3scx0mNbBpeih922d6gEDT2ZKk+tKKnAW7NsbfTzYioCMi8/lwoXoWk
HQpIOtJ00PjmDM/aPnwLlF44zI3+9ro/ZjSQ+eKMOSiqjva0XvrfrCixvxekSCrS
iuq7zQTBMwrAMZqy1F8Ld4fwjAWpPvpjef5F/pQqwauLTPHGhvsZOIzV0yAKvNgy
pgdtUAy9nGtNJ9Kar/3xNTEYGZ7i9+3mSgfjYRMOAVl4JYAsTN0ETJF+F1Ms+jgd
iPNP9HwHxR6e1f3pl5lQoZnboM5Gd3ofZ/83j3ung+qGx29zmFHxRRbjjlG/Q7RY
YhsYln+481FHlW4ovphc3kpTwhan9B2h9suz0liTw/3AnXOBFCVq4VNYeQTqz68n
GFY7RhB1sgYW7i+DR1jAtPkmsWgOzurch5KwUciEPc97OnBBpQl/o5w1UgsX6lJY
qqhRJ9fTVt2eMKlPNbmaBarTyCWk4kLj6DwqDW55ZiNbdlzskUjxFrATxGLaiHWT
QKLvJbDgDyUJwwuQLn9NhswFFaVeOt9pO6cYDhx4+cNJnAm4Rm7DyXmxGNpi40Bi
/3vBu1R7FAOsh3ReB0pZkTPcj7rRUnlMkaATsIlxyVwysVy0tJFPB5VRFyQ4r6zI
fjAaNkqa6ZgBpaje7obaA0jTcz9cGnwYcC2vS6dB9hWXCn+fMU2BddrstbtgXJig
nFESqGteD4Yswx/Bqm1nIRzeO89cAjQr5ahkuDpyFto4tzh3a/BiR0IMnQDm8wCZ
M1D/BBFgKfzuYP9ydT5s84ybr9oCTAtlpnCJsyzk30Z4+RRShZcUSPp+1Ri6T5J3
CWHD0tzZaIKEBpuBBODCM1mIHnDwnKVIJWRtlPnBx5tc21FSlac6IG7ne9nOPIl/
a353qu8vT/oPdGEmddURvGsnKkHG5/ZYJqq13GUWNad9FxuRlN7U4E8lLvl+VFim
N2fkQeRIyLJ/pEYBVJEVc+h78gXKvxwip2ucukZ602zXztoDE3jbpcB8zuKbSOsn
wQEZrbWB7XdzpjjRXuGtSYHPv3nSNDq2sk0T/fV7ft1sKYnuYn17fo5zBtJsxW6l
dhoacmaE9UkfkWgQpGCnN7u4avHos9HF5pAOYuXRpy319I83y/8qb4rnyFoHFu3T
DXkey44bj4/i5L/2wQiUDr11sS0hbOJp51x1epaXcPD9A82H1qxXFtFLRdN+kLAl
yAeaoRIZUeh7A1azW+C/HuWveOWpK8gm828mZrnArUu0hzOV9Q31CiJaKxZLFA9w
6lCpguywDb1DpHI+oAEk7kVDuXjeT0qVtUk1OGrqCKCGo6Y1jnUbRrxHNDJVqtg8
iWZInFSu5UhfPRk4ONW/6VoCCMiwdg9K8Eg+b/79DxhvEPhtWfp0cJDaLtbaMHr6
4Oj69b7xYGGSkGp2uSYO6w1pp49eNHQ87fMffmc2PPtRTzkLwTCLmWnP3YvXge/w
nbOltqgYxb+7K9ABMWbP2/vMJJDQOGTpqt6U9N5QuO1HH5wghtXKtQHENUIsu6w3
L/ro2/x21a6AcRMt/p69zIff0CfkvQHWcTBWTu5GRelFBj1l4FEInPvQY/U2du7W
y0H6Kp10l/6sPZpHMt7WFbD/fxALhOVFKquQ77DUZgiosFY7+pzSwYsuYOrFY6Ly
m655DQfe0IFXeoEnBxnrR++FyMv//4LnpSxOE1hjqFqHMGLVhef05qoD5ekfdyb8
gECNGcJ8mGPZxZeuY6tLt9vuDTbqEYbZrYiqZWlohy4YKLLWOMMhmdYEi128xZgM
KU04PSPWss1Xa6K7xlQg3vsbB0R/dQKUetL4fUKvnr7XResRw3DRu67ZlkZbByml
c9BQYBsSXFataYGVPS3vSePyJ0Mo84vFyN8/fZyRrLkVw/Bmjwmy961l+k/RETVi
iAs6or++f392YYJ3fW8p9sy2X6QAQsd/uW/oWxqE2J17cUaUpeVGDWb8V0TrlOmo
Eo8zWnHuO/y1pZf0PnXMmuBsvnCsOqHU1uFCw//xjvNGw30VDElsAh+JHVq9wIt4
0cXs/sTKIssys6spC2U3DmOPu6/U/h0JqEMChaxv8H5nscGzEYSNuKisQIN+jGt/
gE16G1c8ziQXBta7tVxzM6DQKYq6QOSkrixQmHZ2F2H6nlbQDJk8S8nKqDGPsWtR
Je+WCG66PhyhDF+3o6pXphKuKo1aGdt+Ez3KoFUGTonu//RT7lwet3QHDy88w0WS
5kskpq6e+oT+gOUBuegh3+Api4988yLytVZ5H2UFhidY0GoL5b1etW+aZxQn7ZgM
R5jcoefJAJXAFQRzunAuoIWN27ucQrqlkI72G6q+YEPgiAm1EjroUeKZBYbdJUgb
tMz/y1sd3nRn5VuiNJ6mPqGuz9wcPs94ALPV/WR346tpWcx8LIJlNOZdUK747rqT
jK8HBBuJq7BlYnoyVsKsavKG8N4ZmBfN3fuwgNKEc0UbQf4lrPZDRVEuWdhHPBPY
YIjAqmfFi+nWVxzlqCwGqMhsQx9S/WbKZzWx4a9hUBmWgCF7o1cGsSUw6MbMu628
iPq0zCjXY0X+EgaN2CyCTbGUhEUYzimzxFxHmJQS2wR+5VUrVx8Aoz1AAW2K1TMI
cwuRyLoPukmA3Exkau4AZ4H8zW1vayhingTuzhbbCMfCVuvaJMUqlFQkYY+l18px
AiW0xUw80IbR6EegKfImVE6H/7oe/TLFDeq4TdgRXaiUmyVycvoDSPeEJ/+dOxLQ
RuwOmWM+IoF1dz/mN4TbY6JgQZ7t1eT2SaR6oei8gW0NrixjhHOMKBVfsMlCRqXp
e+V8jR5Q6E6SqjyeksuHmMWnKSgSDjJCO9XR3QMKRcZn92EEc6FCCOZwIStQy69j
FyHr8LsZbo0+Sbo1+sDvyeVOtRWlPVEm5XnDa6T0kartthtk7ZFQaUhdw0okco7V
NrJVe4/cRAplwstE1cge1tLQyODCBVTAEqP9KSyEmXAsteKy+qfjftW0xfCeJjxG
vN3qr+sJkYsahopyWS2qDKr+eQI+FTnb9fYCbFPIotQGFCYPSzMdS5C6Ng3ixgrd
31uGjtB5L4u+Cq9kqCihmlgnvRwLVT3wxfur+axiKr4AxY+gv++jR+uwD/amg9pD
K5xmredhRKPJpBgPDpDST1LRTFbeg/ZmAkiDd+bRqGbM/sIVplzBDGUVl+3+pZK7
t7A9Xl8FHXdMMX12G+vkld3wWMkRAmzfzmsGTcU9e3vnQzHISY+sKXPCWMZw3Lm1
B/7/aEJ71uVSPxNueXUNBEBHxd6m07SchkyPTfyRkfh8NstiQB3U6OoiFRoTWu7I
DR6QO/mnfNhQCPjTvOots15FIW/HQAwDBPOL/dgKZ2VOLfjgZ5YvCzkFzak5nZqO
+LDaRzOfjf3d/pnob+Lq0Zd+05akqKBUQhuw+ZpEy+a7uecl78onJN672cejkvzE
mK6lZ8g3ONC0utr7sLXhEqeu1F+c4/fJHjUbT4RQiJzABE1Tk4oeH2z8VnnswDOX
zZJ6pXzWnj3aEY8C1IEDH8FB+VCVuE8bO4HCFo7xU3KKaj0LBPQ3T9pFqKSBQny6
dIhzmCPgNhVKR1EkrwO2kNHpGAfBEbMZ+hwqsMXAT9tDC44M/O2lNz1tXmmKh3cH
tk/nEZle3mVXoj8J9qFeYvk+ul5c3+Hjp2M9SoFTO1kNruICh0Zlv338xBfC2Rf2
KPrKjB0U+8uoIPk9eY5JRflfX1vI+0W44TtOv2jhgRy4Y7PZduBK5mReM5k6Kdz0
J1Wnfschz8VHuntBMXXlxTDwZC0YL1snLG+XHmc7c9MNI47CqF+FvvVz1TyG5TFf
XwNLpzXkYaI2vt/WA6N6E3q5bLinYdbSaNt4t/D1eOHUV72auuNK53KYynPgDwTj
7e2Mtly+QHOloSqlqwvAzm1i0xvc7Xg7GOg9/8b7BjxYifogbvqsJl1SkCJukwF+
DykIph5wwDEg3lU5eJz/Rq97MdIWZQnttomdjub10i1JF8rIVXWVeW5DG/ek1SDQ
BVCRS40CscoVVMkZzZTGIBZS9QbI4lYkjmnG2lxx7k+pH+jX/7wjyE+icEkEYCC9
4/dJ0fKWl1I0XKxS/aybRO10hO2b9Lzzq4Rztgy3eOnCaYpj+4G4+3By2NJa0VUP
qvv0fj+GFOXlkC27kBFeklk2fg/yEfkO5ZRv6Y1gU2BKj7lzaO9B3qkPQEvw/QI2
/WlL+QMhV8X7Qj5gRqMJnrfwEgirFQ8tgyoUZLNSPXSFdLS9ZQWtn/ayKP2obc1Q
4wSEvL1OWFvec0q3BM0FBKx6TbAr71+2bEtOFVjbJZZWDEq2kLAEW5QxHb+vewfM
+xm8KpKq72G728qsutte8XqCQStzr9Rl9AABwOTEWER90eACF/PkSgwiDboD6TGC
ewAY/xKHcKxZpO3b57UsWj3EMtlZkd+dPspwkSJBxabCm2rHHuSq6L6AuIY0gegZ
KN1qKiCHo+C5t9eAKQvt0t5lZyGkiBmF1iCexLlBmd/CcvWcN/h28+wNkj8ewU9i
5r8Xs4vaFUiGjvtMUNm3Delp+Y3CeLSZh+vqef4JXAxvuiS+21In5xMKCSUprKbp
DHBbJ3T/ptmdGHm5QM7vWJLQp8pGK8gnJsnRY1RIv8NDc3OF8R+uouBAj6XzK3dp
3zMSMjNsRtIMXuz0TL8q2TaNE9Yx5KjOwydLLNeqpI9IUOiz22FKq7LJWo7sjJsB
2xA1hXjINMa10FOvkojV5qB7B+xshlrz5/slrI91SOq2/DtfMG9OhKUQAloKZPqM
aElVtz/elzN3h5JW2T9NqZel2V+knK2iQj2GX7Mtc1e5zdHd5nNz1bpoVg5BV36F
khPYcAMhiiPefuV8QyyEelbgSafQK5YmTgOiIOzgYKfSE8WLblh8UK1bt0kxNqz1
WTSRyjnhEQJVRRe4m/pnNfbNO3q6uQEfXIIHu9WU/GtztxLObvEKkcm4pXfa7hxP
UaLSN+7v/faUwNF7C0j0AMpYt5vE23b057X+duLO3si4nFqtGxqrGI9n0EZSJ+4K
bJVRUxvOdN6QK7nnFNR0Bv4AD1cZU6msTrvkAqHAIZ7W57pa2wDL0NfCm7uzQF0R
fBIwvySqiYce1Jjalu1Vyy5BvUW3Dumnfe3BOvuc2TQ8mu63wHz5iskoHV15q68v
T3Efw0tj02yaVYVq8vP8qz+i/nsKkrlOwrq91CoJgdDRyH9OHY0IPtuTMF1MRRL9
GkTbWVO29lptoQsAzHk62uZ1vbxO4S6X+4l5mFd4YqXMcnMpsMeKm8sTv+TngZib
nldWazIBpAz7vShslrGiWbE4M+vAs89vPXLWRuIAFF6UCaIWKfrzhcLgsQ6tPJPa
cjoQYEnXdvFrS8Ze6KThcot6OhhSvKc4ViaJHJ8aCEVSog95mlbGYUDXchUIjPil
T9epCVx2ql5rpkgUrLcMBrRwyzG/16juFnpQOh4mSG2RA/nFjxA5scz3HfclygXi
7CEnYuG8MTxnzeaVUU7NB5FFFU9Zbr3jtPSgafrIkwYTS/wy/qUIVTlJJbYQSNjC
6JtB0k7rYFnBqcF88DuaBmJEy6w0D8y1dHBq0aSWhO6PymNri/yX5WwrqtjuxsGp
rqszJAKL2mJMWHf2ZHexw6hsBWqZQa+ABxZg8jWh8bluvsDJP2SxaKtpnG4hfzmy
WAVR5Gotu0MzBV2P/Cz/cA/V5jk/cU3w92Jy3sH3GPpHBIN+P1TuNWMtaqPJlTBh
7qlu333f8ulHn49AhVYWxHQ6zZPTingbHK1UWXZOkPpqfa0QScipUnKAlkP0NiZA
KrJJHXvEMg7E/JSKK9HqI94KbVBLjvVfJYIKJau9WJHpY3xjhIbHTtvHSduJiV6b
pCgB4RyYUxwkdTko+KvQNo6IhCGZJqRFz3pv62k4zJIIlZ9QddZGUPAmPVQAHE68
7/pfUGG10Li9yhYieKnqww8TKPSxa6Q2C1EHLNBJA9dP65mAqBqWpmCo3NtVxM95
8ZAKhbsqi5rrkIu2D+7kSJhk/6LJqyXHVOFu5MDKQaukVBfIJ68/m1w1faEhB+CK
chiiwc1j9lYfI48wqtg67DWEGIIQ4hrR6wBluK59t6DEx7HPCODna1l9NF3Cr0S/
fS5NJjzIeTNRWdqHUx+xptP/1vmlg9jXp6O8Ai3oNKk90f5LfC3IVW6ewREyoy27
Vns2yqOjGq5E1C11EXbY5orOigjBZEPQ8HDl1xng1RJvImoOCAVoCVjGXlhziGkw
yNyF8sSjtJRhOuplTWlep131gZQI4imrss1vhZ5Fc0T/7deiIgQxB6RUXSWN8cuu
TH2FSxEjU0aGU+cbRSnBz3VSPbJMy2i/k6jMHqSyWeicawBuGXZfjvfAOqjPfOJA
wGKYC3cxvAWDKwA3h8hQ+eW7w2KBL3UTZOcukSOkSEICPcN6SMgXaf/KjSJWRbSJ
AP5722IftUEfn2ws2DBNIAcr+hskYR1JW0GNXgJw+hR4eqa8Af1irqaAQHErH24z
D3V3Vz/j57WCa7YzFr74HWYrB+0xfqJD+dFqK/0El1lcmq/sw1V7CwXu678OgW/2
cBq6v+Jtwx4t8A+n110Kez+utyUqWLt0trVqORlTC972Ob/Xhf8V4PZNpfAoVLpm
ah1ftWzNS59cNSXgQKh4PDFrzauhpiNRg0aaEu0KaFdzlmwJTsOn6Ti/pHih2wUO
0/H+1s/l7hrjRLAV17l6pfXq4ZNGzQ/v334RqcYBq2hCCMavqa0VQIIm8HlbR1NC
QdXW2SSyCrq4Qulqmu5F8LCPLzaUK5OnmRKKqIDL4vt0JNHRZFRWHKbk7Z90ZeAP
lmKcCEYSNCW+bSzRN6myoKaN43nfzjLhfHPJmBcSrY2KPg2KzuDl+g0LlMvb5ZWD
w455ZRMe+kEdIC8ffe6Yzsd8be2otLlnMKMXNkIUYDQ8DIkpulw+zXUGeuViCrh4
a/bGs8aedqlym8pyEd1dQtHh6GkPQb1iG9q8tMjModUTcYT02UOSa0Mzg9Yv6d2Z
vCLQZXr4PrLFhE1AQYTOYeFWH2QYlKjWXHoI+FGPlY9Uyyzv/RhcYkpcat1Ez4RI
w/ZM3/O7eyo7zlDVcI7chFp4HVC42wboSUOK7DPHMAMRNetM11zaVDhBnO9L3iqT
PWC3TsHbnJNZmJYPxSvEL4+9qotfqoy2yEHC0OMZ/VtVE2zLM/p5+h0rDyunLC0h
jn8KJE4rYS+V2UsIPT5phXXr7viGTQCcpp1sO+FssEZkC+dQeUDNPT/CMr84y7xd
W2OxKaj+bndK+ZKhk4VTuq/MiocYFueiouXtprjbkjLWQgsfdp8e5LgyKWyLUszl
Q2keihkQWCWGUa5N2I+pqzA2vT8QKdfJ9qWYVrFr4nBn+IvPKy2ZTs8bgrpwP0Qj
zI6qHp8wGMGL36XDZ6NoNgUSKa86CSZxR+pCCfeJs+WAeo+tiiXFQzrbbJZhfj9Z
yWT5m6LfpwKbLRJccAGe5X/Wpt9haOIBBhDHBOXH/bxcyYa/t1lohfX/GL5yv23m
jyFEunyLaDSBzcVOkyvoegQxNkeDuIRvqvfLjpneoCvtnjcjWforrR6TBc4F1BiF
VsrOdhevnQMiYsiWkcU5K4FtcEkqdoVyVzsWpC6hcBUPH6uOj/gYttVfdK3qXPxd
4qVuxqLV4TtdJD4avNhu40/OKCYWifS9Gjcg6caguspsXrbMk+lSIRnTsywpEs5b
0hi7pSz92iK7CtW5ivZexQd1ZS4QTWwf0HrKioIb6kFv40eZnjHiHJpHGaH/dsf5
yPNVWeSj2KJUe7WGSxscIcAuhANyFRlidt24PdzBx/WBF9joux/dyk8VXZXbXLu4
2pBXEjHYYXpzoy/b0dBtdRmd45UoZwIriDCisZxDkSqjns3A6iiW4JXvxpx/W5ym
KIoAjYkUJNncPpv0wHrS3LhfPUXxdkY7McyskW6sHIlZfdo6vY0lGHyFvVpC0yCA
PzN2qFKLByupKTnQfNR1qvAqbwQQTkD7BtyyrlUP1RVtUnxcqM/dWhCKxGfLYUtx
ekhyLMGQYH3EqOFfQUkKKDiJvql6d2FZ/lPnacVCB0q+LnjESQl6pC+veSTreVhI
0mNNGlWIHt6wWLjVrn4lGjOgP7/fEolV+Upnn0rmbvd0INYQT8ESCULHnlrYoBWh
GwlEbnwfIOfVeBchDsFSy7MJcUsjZu+UCvAYYIqOqEPrkAR2mZDfDXH9L6Lv2qut
u/ORE/sOgc9V0VL/UysVJPvSo/UfVgDF/jGy1de7HLe090kcdSR0f3jEWB2JED/Y
7NHtTr4dCMSwciGEbYMFuX64P+b5Gjd1ZSzJ5fCl1AJOfcWX53Wi1Ilt6HOhxAwL
WfuhGn0MhbtMLv88oOTdcZcsOcijpWqUSC2ISX+5R3jwDjDeep4wn1gn4j3dUs6b
xvC0Io1QVhMYOTFmaucxviDbKF8eHlrp+q53RYQ8MneisMEsyzHf7/W7AXLFAI2b
8ApkDpEgJWEvurLUQhZSNkcWZRH0WU3ekq5Q07e54PIR6nDbuBhwNwXj7r/G8it/
rGDf7OAZzUoyXpQ0FvblOBxRwoN4F7gzfWhqoR7i6/poY4bpMrsoykpjhXVUvvHL
RGa7wJ1T/otJhYXO7jfNbbU1VuwFworYoYM7VxPX+fKhbAUNBdTkl6XWn7QrSXW9
cOcb8qKndb88EI3kx/yMM6e2koV+J0/ptrMMv3UDbm7Q53d/FkQQJUB6KCc0T/lE
fkWeyKVOrW0iTa9aiF4g+wGLqx3/H+SQas7hQobNEZJhHAAaXqrUqFtOE8fsUKLR
gJH9b6sytRv2hY7mRkecwz+oLmF/YTZuCQW+6GE7C/J5XD38Ks4/sirVR1Nq8/td
YxDpEI4igSLYrKUZJJYPTQQGbEHy0EjXUATZmTNfqeuUZOvxPBtu/ovfdKryjVvm
wZVO9IAvKMkfN5h+clt0xKHSB5Jxib8Xeh1jVMXlwB4Rt9Zu1cvgqgAT3pg1yqCO
YQ6rrFGyix/3CM9Uy1jBBAFhoR1fye1a2iH7yKa8kuE1h2Wu+gXeoaiqTI+P4v0g
NZGIdmJ9vS5fOaTvu0ifgrioPpCUcKxCnrrdf6NIogcfYNCLHAHkw66i3S4waY7k
psaf9FBtLFVQdetAB7m1k6r4DfJmT02cKF/sAXjLDnvzWbzNDu3Ec77NK4JbGNLw
ogGg2QbuJtGGiAv/mGJHuKjayVuU4zglLaP/wVKUHXaBilJRmHXIyWoiawo+GuDa
EfqvGmEqdXh1AgMbDjenG13yu5IyALvl3/nnHbU2o93QnQtexHaC1Ol4aY7Kzlhb
h4xdp+IV5kticN67kxrCeNibIUO6tc/YvSZaz4vMFgvowDWW85SfqT7hBKHasdQF
C9eeS5vx2JZ4xCGO1tzFOWkHyJEg/M6JKYjFLWJbYmnHb5sIm9doWYlBdJc5rf4Y
slpJsz2IAsO5QxNmHM0gDHRPyWB7pBvphgRWlv8e/L94YLAvnfTmWzZYtRB58jyS
TcXNAMmjy2IP52n0XZfYElTS3r5yneeN7Tq56Hrqmt64kcGVUuNBgF0aDTnQnlsJ
eSJD0/ydECgxaDPuGZoReP9RhGPC9JcjNIJxE5B6hZ9oLFGzPfzxI6zMt4wW1vNj
nbFPuPme/C9b1mOdPD+kcYcfrBOlO6e9l/tmhfeuNZ+mT0yndBlGOMkxstb2rQLt
beV+u1yg+3KuIqsQM2gz10v4/aZBA56vK7+Bm+HrgcDjuze65/1JGIy+tioz6Crv
/nE7cINeBrbox8JVsC7JAME7/bpYffmeZNhaw1X6+nRHNYEKnckyuCufR4qsddc1
+b/cyNHW3BiPANEbfcdVe5fl60UZIBBS40yVzpAubPtJWXlOdBpFk9AllW+TiOU9
P8MY9OJMoOFaNZOnf0Al+4jvLS/ASN2B2W8IzWJ785rrvzhDV7dp9Kjll4hy4A9+
K13VwYWUgkJMDU+T9MLo9gx2e7OIuPRXyaMNfLpx9vmz/0zafpRSFw9+id1oWm+K
r56t/eBdEWwbTvA9MEglSs8N1lh2eDVQFl64YFOAfD4WHRnbI4BjM3paIzjyu6Xu
jWzwtYbBlv+gJJ99Bcfu27z2ZSWzY3ffTgHhSwqLIB2LmNT6maBXgCw9VwBUkKe1
SE3a+xHRstnqJCj/cEY/61f2LwLtxf2SVl6Zpb9sKP1F1w1n5ihSGckWMq6O9B5C
7WrICMfLJEOMBe0UHOA4Mj5pRz7iqcJpAy+hcKTAzuJ8XXKgPv+Zrh2e/eFubzLa
LjyajF3m2XCKVOaU8k1VOXj4OzOKP9rf5mfpnPqRzYLmJddvLVxyVVPVB93kDK+p
a1R7BSaxQKw3PslNlefi3t2obww8CDHV/kkZrpMxgVBWy7FTFT4cajZWhaSVvKNV
M7SsBnTjMg3e8nMY/S5V+gFp7YgAbLnMbWhIPQlBcPP9E3qZCmy66ZeHSa9Ty6lS
5y1dPeNy5Qr7jr70w7+BHTriouIYP8wiChgVoTgsZ1aRzRljEyslgOwToNDJgeiz
3NOYg5Di627+MCwKzQpj3IOpGgmno6x1Wbl5z72CHf4q/Zb1dpqQ+FYL6Yu5Ygmt
kF/yt9xzAKMw/vn2fMQS5XntlLS2ibtVEY+UdePUwFsaNG6CL9hLj9Xe6IVHfB2J
+5g2yMZIDvGrxMa85cMmctQLP5/qchZdxdK7cQtnA3J4XR52yXJZvx5bY0sfmdEI
S3Oc5friIk9vFa08fURp2OK0EvE9sIvM88q+nsUNcgVPExPm/v7HzuerGrSHg1aN
JJms/+sp0JOUQ5N8d0TZPMGITKwYNUEzH8mxTGlIq2BycSraJP4QFhryO+vENX9p
bNBjdi3O6jZqb43zD85FRtfheMfBv1yW3+wg8G5cFz2YhMn0eNGWOokG1IzDl7CY
tjLq5P5/finIPCWxp5U8hZuvh0Mg8ayAxdlifjLYdiCgz4r5VaL4YMjXPv+SDBrW
Yz1hPC7FYLMM0dRFnkWLokOzvVUjHmRl7xTM749GmaLq/QlRMIXhOlaTB6fo9IPw
qAHmsciLVOEDFBb59SXYOzAS0dd/PqWVnAYYWCBlum7jCLpKqqxM3p9VtF0GA03S
fqPe2qjnAhGdjllHSrF54V+qVEWBe/B8LOoauGEN6zQLg/kHWPt/NErlWJAGAMtc
mu5q+e+i5PHbyxcW8z4Foxw6ioIWpUdVGbMUv3BLQ8Rrs93vKcRyOiRYew21IMWv
4nUAXa/4jLfRSqM8jEtQwNLwwIgx6hMwXYfLetopN62Wj1YXdF7nvevrIeSxgmmP
g0USz3woX2rupeM1hUHRddFa6ElRCrYfTUJsZFXmYIvIujb4wNXaB0ZQofz1lvzt
P4lM8Stu0McM417IOeQCzQBmaIyBDoGzXWxli2DH4R0gGsFd4UBk1L+M/wJpGXG2
VE7Nz2amb0aFtJw+u+rNqGozE10LE97JI8fMnS4lWuYGy29tdAVnMgdD3R0v39sU
IEMvfa3HPsztbgisu9zLBcEv4VkE+mkeBIYm68QyvQTt9FmCRxW/clOBMQzLpnWj
ijMbvTao0U3gI3kLIbjRMm7uY0ptnwpQZHiMQS1lKU7A2PlCHgTiCU8/hAsHF2jV
Dmj1/WiiLp/Sb3uSDNEt5l15bCOs2IfjisPlTUabBNhCcX5ZhiO8dZUih0Ae8TmM
xNCVB3lAlmWhQk2SC41egxT0TQ/NuSxqGX7MuaFpJkaDywPOWnsqY4Nlv7uMyykb
P6O97VCUqhSwzROY60Xhd3OM8IRBiOBmZoBOcYt6yE27ikW0bqNE6WRLiDbWJURy
vv148QmKLWTNgBUxXzP/RuYe+G2kLChGxhe0JmDs8A0k4V2gFGx4fesMSIYjOiH+
4V4r4r2F84YofSOdGiuh1al5qzuykex/Xe6OQm6zBcaaUXJPsLQJFD6RVjShjYGJ
VKBVUxPw+6rw/iAMM7MHJWTU4+dinQOvUSM/RGQ2edxV3Dvd1jXGPChcsY622XiU
g8As6zPgSMpz9apyOaBXOrkKBUQ2hCp8CLGpkLWBMmLxvaFBhKFTxuYGkAJziJTm
92Nrnb4qwGckZlVmbSU6+4glTDPuqHCM/MS+u43yWOk6+ORc0FSKIcEkFt2Jt4H0
g/GI+yGTTkow/HZhlfHbVkV1Bpytmkua1jWVkrf4wMxK6grANMm4ntNhti8pX3VX
jb/6GdbNboFx4gf06v3Yg4nS7rVI1RoCpzvJ3YLT1ULY9L6vF27Me7LyZvv6P5+X
4WDBJYNv5imegMx251wn68aPeDL5ZB3kQM0KlvEu/bPpjas/mxFnC9o3lnovobkG
Mw+PiYxh+Vpsa0VEzl7kgN9WZXKLoM2t4mJTNmHBcuRWFZiwX5EUMqry7nB7OVsY
S6P/FbvR4xphAJRe5RuGANFkWxDyTDtAeNCEVVuaiTkjgV8GBbkx6Ihj2dsu6H9o
vQjrSZpt5/DoichCOvxtjXBEruJAOVSAca0gh/HmSZo3GMOIEvRx0kGb1jLYWNGP
kH+12sP18Cg7PfGHbHQYx6XJxax4TGgONAcUM5z8fUWWur2hbRs5uVLLj1wOPvoD
0fgDm1BQN0gxjIvraFDg1rCL5qKvlVCCwCFeDeuHzq5MnyaihBeKJqxYwHPziUa6
YlDOP2bI20FX98ZIe7kGDTwFb03/kRQ9EQ0XjrYdRWD+OAB5rNTdmShlP/FBNScn
oInaw6jkGqPQzurtrQah73xzhHXpB60nCWGvmTI72pg1AV4//QPvIZgYNBnW9ELT
sd9HDsweu5Y7gProRBVzLuRxJvK5H/qiHOPJ7hSLsRvv5FJV4MnJyOeaOnq9f8G7
R0B7XozoD7ntfbsBh2hXLHdFCSW3FTDl4SD60pTexoOtso3H+jLYaoqaYITdXs7/
XkICB37DdRg1IlCPb0VEvSc5syJQVw1ZIX00P0a9WVLNy623kXfe2oHI6BUGuMum
df6hXuEXdwu1AbjKOI3yLmHf72fscouClOLCbizMx9Nn4lMZ6Ge77x9MahWnC20K
GE5ENWqEIwiPj+W4Uk2ZNNN36DBhTh+y1M2vfCbsNhGzaa1a96qDhW5RDgsyAPrS
HzNMpIVm1Uk2+w5nmEzsW/o7hf5fn5LZz3++3Zfq9CTg4Eo0yRWgRK/8pCegx1Wj
NQFUPmNtcguY9KLxoYzAX6DOvfag98guI1TpbZI7iImHh51HsUFS2QW+Ei2MS2gP
s7riV5ULlP+ay5Nyyu3EL/yatQi/QkXWJyE5QHXqq8bAAGtCVfAEdolnXOAEVcsV
SubIobYXlJ0Mte2rh+UasNVaKqkEojXlzT1ne/jFxG76ntblH09q+YJqqUK9yFbz
pPUv1NUlbiDQrUkTI/BYnlVcDQrV7RlF8zIeqiAkCzMdPxvK9yKrt8r3SPChzR4s
LcOT4zIVYAJvo7vjJqcbVPcVR23VPjAQ+HAg+rpwW9nGBETvKFW1ZVjNTnfsKqkF
HiKxUQ+palo/ejfLLB8EyH/CDx1Zn4QB420PlaRcaXkohzNnkXePUaFreTO4BqKK
+b88YCfJGo94eb/jUt71mJnHHHTXPEdgDm3EmFJBca2DZzNAYIP85B/11UrLG+k+
kIz8sr/GrH9xKerAbbOix9CgNHkGKZChKRcaHps5rucXRLZbDvI3yLh1v/rDjIXY
UZ+MIJD19TVXQupyFSzTToIiQmrri8sjCBB8cOzB0BtnPdCohHkhabJ4RUxXfsE0
HCCN8KGY+H25cNZp9VG/u53smT7CRRNiewMQfPQSgtit75Bvv2NLIf4R4cG6c500
AmmGzif3hTVpRf0z9ngYfHAlECX9R1FaTB2I+aN49ecqFvX1V0O9aQwdXX98iJcp
fexaTL3XU5ca46W0usJU/iwgx2FwTsFELvEe0vgT78FME8zTH7YxnCATt+idifgo
KWMtbH5z6eVG9F8aV23rPrTOq268Gxw2HZUIBLWap4TukpkBGemnkr6D47NrAAoU
AlvkY7FOyIKhwfY+nNvwzbu314/tmb9QdyKh9Z/YO84B/AQ65J1T4XzCh7O2S6ms
JByVFId9WktORJzl0d4LYwgVc6Oq9U+4WMb+N2esMV7tLe+iNV4AxtAOjT6FOWi7
WIOmhJXgzFJVPNXQx1YNf5wgvgx1n/8mNOcAVtjvmmF3S21blBzF7sfFqNA01uy3
170253Y+7Zqj4EUD2rmOcHTm5gsHAS8efOQJKaUie574HzigXSZuHMvzzlMVZLl+
4X75WvWOOaI0Cl7UCQrVd6wul87P/3LWHbkfJIdtSpNzk4E/XKUcBK1WGFp5cL6x
0m4Ih5L6ZSeJiWlYdwraFEc+Ds9w8cHkVk5CtorAkJvqhGQNZOKz8qR33oPpOfOL
fp/p5dTDKE3LzzHLSnxPbGilGzi6lw5Eoym6F/2cJHOReVXiQ6uKDaXZjaErxQnW
d0CESrvExz4TdPW6sCKSDNUNkxbD+pG88pbnzSeRa5tUAnrvNtQEJaGrqQiJxkyV
VvtQBbcFkpfizFdS394IsuB7hD5opZm6KDiZXG7lJREruiq0HGFCgouJuhMpHB9O
okuwonNV2X7sSuT+khaRDceOjFWNX/AtPrBErgFG+RuGC3w4KhVXVcOd0DIGPk9t
pbNfmsZ0PlZyXlxlWHkZ/E0UuYj7Mj4uQjf20ry8PsJmwKDhbEtrWaThjIH1S9gm
qUQPnXBskxHMsckqe4t9dD/oYH2Ww+SnwWfR4UAHQPvNh4y2TeFwpBpeSA6izk02
4PxXvIdvqcgs3Br6cxgP0ylnjnEEOGIgOeL1gMxScQAUC5sadDuqBZLpJXeje21D
MXDNz/Y1hPe6dflmtRXQAsAA9O0Hdpni+fwRDG6y0RQ+sQJgCuEpdNniHOrPJUfs
fnQ7D0MXO3JXmgGw7J2XXtwDPqIIG+0QB0HuSyut6Py8lTOam4b82H113y7VRJ8S
SC8zssHKaP+Nr6Nz8K648pku200YHOWKEnIC6zqDRliOruA5Tf52q8/qWBtm7yVg
XqEWp/I6jPoy5Z9/TDXyG8N1FrsUSywLWU4i/CydPlASrFLGY3xJQLKfHNClAXn6
M40FhWKM1+nuGRNNAalyTN3ejaAuK/Hn7FrEiaWS5zTqI2cM068H5UofXkWPb8fi
BQqETBWIuzNkfd17AFX8g2natofdtsY8eDScwMzJBqRq9SBvY0MtM3KgAwhoJzhd
WpEEjEyw8jIeX/1Kyde6MufE+kJEkGGsmuMqKf/7k118BU5EVo2MoJbta6i7lH11
KJm/udIG1weM1cu62qYC/MlZvfGE7KRPH/OItbf2VW/fEjMKPPglKr3ZguMeuCoB
gNhnGHVBTQfYOL+mpzymef/txZfDFMxeOne0t1y0/T5xWsiGOs8GVVSsPlUgfyrg
UM5HAFcxHhKTRFqId+iwb12ic92HAE5UJWBXdKK70wNDx2FJmpA3kyinKCbQ9ceO
mK/+uSXGmQI0yOQNfd6vhGxeeK3v5tBIy8rQl3/guSiWMSxZLGB1kZ0rbTjOInhB
FU3ff6VcP7cXW+38AliHMscmkJwMEtH6RHDEuN8HshW+f9r/vFxc4AnZd4RB5FuD
EokqxR8s8IpBjM4UrV1Xu6sAIT4ZPjO+azLrq8wtkDTLuE3zj5lWqLtpYPMFPZR1
OOoESJZUuRxk4AjF86qdNUJ2hTfa+xZkZQVuCRtdoETplLbDzfp6MUML6jUMFDbX
LoZosKPtvQSseR/rW6OjRJ2q3vyexC01CBizvdmoESNN9NjNmpCguGQLZ05wTLdO
P6Qo322lt2trQLHj2umKaWKqXDW32kHxDlPTlPkuh/OGqAdkenmTdYWIE9c3mKdR
fYw+RUKWrf/VqYa1EgTm3oTZvLqzskeq1debNNBkdOUDjUZi35vONIPzgRG2Dqud
qgJ0rDeCDDof/29BKUyDcZwaqVeasV6ZzvugQNwKM76aCs5vVMwqtO2cW0M/3rXw
BfpMdjl227AFUNlDK4fx4pcZfQc7UzYyOzPy+nEYjC7BuwyT9kuXw6RSiEV/UEtj
11B8Kq2/lOe4IHUZ8GmeLUeySsLt+B/MN3pvLlQ+xrvWyuWBg6/b+OB7t80+SdVC
vb164UtdZyVLpnzbSR44QZxsvD9COpJKgaKtx/UybOC0yHm6imNy+x1vErmFN4A8
Wsfq7Wn3l/FoxPqEY/x3x1ou/eFcZ6YW3epS+j08h0NWZiOpcjd6RZ49AO57dKRe
BqF+Rn1sP5SkJgsMYINF/FGyvuIu76VuuVoUhFRGywlAarvjO91rLzcF3P7Bx92/
//Lu1S50uQXdmelhaSgOA9WcI2RbTG90V5rulHjupmePqTgTnjZma8xKTTv+zh/D
CqCkfJNvu8Gzf44ut3LKTEF1KKoyWpjJGLrS1FYRy1ac8fX3m6udt4kdNxyxKI8F
+d72gOr9Bw5zCEHPsMHYqvD/M+M/VRlggYGDgn01oaF4XSF/Iq23epsPvAnwXZpo
1x9bJMavCalWWOpwodFsECom2rUFuWMqCmMSQ1AzbRmCSDYw+4HSkF4CSMUevlsi
X9jCgztJmKoLpIkUNewzHfwmxBpmMP5+yxa65jDSMyUQLdPwauPkJtyQAw3pG+Bb
hd5+1vNXMqL8M96NHkr0MeTGHwFSpqWyrxD4HkRIn718cec1SqhTYwJ5YnjExDCt
LDOHOYlK8kB0GxB46V+ZXpWITaAgFJGmGFDqfjq4aeTuaWGLEVhs4czVhw7bKQ3Z
hFWT/XnRvZ1Kk+spHufYnm9TehDwH42Q7YoeMPxexstg73BNin7DNjjRhPkDxgF4
mVtNVgjSKzjD59B7O9kFkMnN5IfprpOYPqOIIiGK8fpOyKDdZH/1+KFo3YOWl9cW
InAkLke0kQXIE/FKw0IWDXhmwwcEAJbt8yM2NMMQCCYfU6/MMt+unMPznPJbO2Mn
N3rygotNx98DD5T8yIvBrzK6vwdJkDBN2bryFJVVWotWvNsyC90tNsTFzz90/WZY
m88T0S/nNOTs+wxuyyKwu57irabSYJzouEEPPDk4mMRQ/Nzct8KUr1gaOW3NNges
ews8Sm6uuZF8ZpMlqMJ2C7l8KL5qRGtKyavDt4Ck71xzFIboDiS1FCFg6VEQzJPn
2J3hrx+AjsOMT3tnifIwkAljTSKd0LykSh21oboa4k8ZBqGNM43OiJvORrsc+/kI
ODi8ZCybP7mbzguYraiYR2hO/eK4HWrCsc7HLgwm06S/roODMjANafBxiGn9WyEk
R8dDTUnxZw1XFwZfrULtC/yWQrBxBKLgfA0tnZfnD26A/yXqTNrvDYFGpUW180M6
cjHS11I0ZG0Ms2yLQTKeLRfOhePMgU3bjxeSfUXk4rpk9HRnCevVKAmHsHasha7I
iQ95j8m/yDNh6DUYBI6Fs+ZAUul30zDzu1EmvuNiALdG6uCF/UuaCWPwEepdEDHI
aqPkTgvsiwjpECmBTpwZ0ex598kQOpSev240X2CT+LCJDUF/G/RLCuWkZDPbq0+s
LsgETnsm28f56usHmjjYnavpVRfhxBhav1p+HNTB6P3ion23OgiWkgr7tqVhCei3
Wl4rNkcxeyFIzaXFXUXfCd6+B8zpxk7824Lmh/pWh1i1RwdHbHtrWL4zOZcvt9kx
gWfeOoA8XovwPz1EWFGGJRgxwrepQDh7oQ+UEp8E9in7AL5D4B/QaPOW1qsyN55G
UPONVHVaSfzJ9atduWz7cxsX6JOmH8Idh1xK82/GVJ5BC5sCyIpDzWQlny7EJRqF
tWWG459Qi/AYIDbQ+04DXiuyiORwSELoztZb3IFY6vwFF33fYZOETcylLbTq6bwV
k7Q2ZG/vSPRR3/m7RTUmODCl79YLrd85gQE09FR+8ovkfv3n1YxTB34M9n9l+8IL
yVKCYXqtTBpZd11nZVOEKSQfN2X1dsatGRG0WHfcTFfYUaY9xjyfQNVpjkpErCBf
FSSf9vdKYXNtv9avuFzW/ZOSihxAmkzUMiiQmzOz/ZANH3h9/rd0wj4VDIxqXim3
vK46PctsUtI3XcHKBeb4GGrH1XlYJF3D6P75HEGpD+H/txo4X4CVnX7AwG/fys/S
r2U2OT1OXjIuj58eqRigsapOsn7s0X4tSx66Cf5N4YTWJxlCVOkjkypJBWcQcuBS
mZqw0lfIl3YPbvVkowyEbHrkvODx82TPLYyG5h3m9B+3wi1ZJlQEoTl5oi5VmwXU
9fzU0ZCZWhTJZ+4FIxBYt57vFXKa8bHuLn/VhZiJ1dQANQJxtigtE/WzbZN0SfCv
aDjRAtxDaslH/UaSwOxvPipqdHDTHJREJJbqezHd9yuwAP7Q2hacOVeD0QL7O/wm
SHMFCzGue1reI8Y8hgaojqWubC0RwEk2mZZsCd+S/Uomim8qwz+4edy9SYJjPyPo
9UwtKvdmNmt7OT+29vKpIlmqSVpqnM2ajSD5wiOXwYQIAVgK3VQivvaleky8VvW3
m4OELzhwisKoLKpsqp9Iji9CPJwFSIYptPk0JH8NrGOaUmncmNUtpP8QVlJHp5Xb
b0ekYIRxzHHuNCmMcQBX7cN5bFGxgdPSxRastAXurQQSlyg2PAuoUhpL/Gx9v57Q
0xhS8WcDpvxan6U9fKx2bvVcnd2+PFSSVHnefCSlm4I7taOAvlYAF2EN4gNpd6ZO
fdaccAObMnAF/o+ifVrUkjDzao6ZIuvctVBEABD0HbkjdKVSNnLW37CXQjkKYZr8
jZTMNNz5D3AxyhAClB2+lPmIQlO9aq27zxOGV3WT0pe9Q50PF2GlXe9kZwN8r9K4
qcDpSAbHVtNq6/Uh4M1INKIu/UNKT7aOIRpMgGrcbhDjsaoILlJfRY11QFo9PFcC
p/crB9Gau3JI3t4Dh2vARWwrvd9q+hdtbIpVcLmZmaY4Hf2/zGUy/gKhco2t+QI8
c2FNbk/ET4fOXFq3oEL4xlwcyxFyte095BcogyNBTIHA6VhJiazq6Nzu47n2GwpB
4+vM2bUhBTj9UMinK5yf0golYtdz0wak+aF2Yc/SqlPWP1ZAkBJwiaVAiICzDsxU
rAXkMdZv9DrjrTeQ/kYSulynwR2Iep2u21PrXA7/F3YEH8/cKiHWYY5tcLtrQ2yy
2qvs/G2FbfMbzM9nQy4ayaGffatRvujgDAwAiD9EX2kUN7SZ4iqZM4Sent9/r5kN
t5CwhN/cGV3cwo0mPMBLL2Vxx3JnTJiOaSs5qKIEmv0QInFjHAtPirdfMFd+2fz+
ZzxC3WmEY2xSwwXJIk08wnG0pGS6jj9r05Vam9H7xvXYIOMVHE6p/h+rhZl3EVD6
T8vchECT+wVDC1lKwFa072zRNd39Q8umlv458hb1sw4wJe0/MsLLh64ZL6IWqkHZ
zW/rNmNCPZ9c3yxWsgRVikz8hCwQfFW3A3BTavS3jvo0w+ug0UmsT/KEehQSKk/5
35fEQn+lsex9AXC3bfjxPPc4Qt9BafTUGA+H5G6DfqlFM92wZ92P07cQXxpwuNdg
67Ge8M6bhTu+N5eDQ3L21p90EQtT3AkZV+E25eYY21oQrQfa2PwelFjpLjxFSmJy
o4OiNtEiecmXrGap+AI2Sm4Pcrt7tDR5j81WYwCarosEMLikRPr74vhmTZu8edYA
uOfeRV+McZrArKDClZ+mmCvQI4YBb9ZjL9MUp6FK3EOINGpH1bYHiHXfbLnRHGwh
OQn1369DKJw0KUPoL1OibJHNwrVWygvOlkP8h87Za0yySHc4MMz+lUlUZSVOm2Gn
cHhiyGOW0aJHAW/CxzpavUT0FbwmW5FlCU19SiDrb5CTBZ39dNJqafpo2wO79JUS
RY6h40/SRhakl4TFoGomjs3ahcaLhJMdvFD5mXPMk08RJJe0rSg8caV1kjX4HCyW
aYC0YnwFihmDKhJgTJXzvOuQST2NZmOOMdyPVo5ih5PnP9GqLM8yNFnjbSxOmr4A
CMd0kZGhgz82zsoT4MoCC2Jx8aHeiRnzqhjzvqNBYVp8RiuP7g7sEFIr7LNr99Ry
m5VJP7TYaAoCnPeeuKwvlsaH8CPGa9WrFflOT8yuPQkUiXf7cgQ+hR6RCmyNgyvl
M6sVjNzWEnbQ/Jdv45RUqEBhPQhMFyjV05taeDD9maMGfVSZeh463qgF1+pAd3Nj
0U2uY1qUPmTMGDNb+1Ca9XK3Xi13W0Zv4NYvyPOE22zSXEWngAi7cmA1Alti86N7
8VhOLXEs5+CsjbIuejLWMa8GlDkuhHwBUlRavwnn343C5x+8kPI0017dBFSXYv3j
V4v5aY+GJ+Qv/7KqK9Pf/Z9G7mo336GBmTCxGAvG3jprP0ML1x+X1CegPRcu/6B9
YCujIN1plv2ARzO6q+D85DbWBDyjzLJFT4so47ALeo/hOMpdxrflsQYmK6Rf57HC
nsMNyNyxuz+WRFmNFMwZQtLMOVk0DccA5il+6zver814OicgfpqJsVQXt3ObUOyW
Yq+1ltnqlzXmpdllhdEs++PRSnmrP15aWfCCMtsb0wEBhMtGSOMczp6L9be4aEGc
NMxvQX1Oa2RWCLC2PtcpEngaDdom72dhvODdSLXNHDYhS3btV1T3ZHEEryMebNbu
afkvD0hnGuzOWcm0tzGlwgqj+bRr2X4SXB1jrY/DYF2G08KsFIUIWUkAJiNkIbeT
3W0tY+2498MOX6RCD3frkaF7amS/NSy7SkvseieqGx3uKBi844qwAQYBfZKeVCdh
HNxWF5AKfP6jJ3Ze8dNAuWOZLp7u6elgDrwYrcUXdJ+ga0OAii/vYa/YzrUZiUk6
sn+y8hF/Ibq2ErRaQ91mesd+2EwdDmEquIvgSHSZVF34wS5u5unBcoYCbZn9GSsM
N6jCArPEmkqwTFMrIliRejsjWqq7GeVZDjQTNOoUh3ugHA0ArYg2MG/1SQ336/i3
TQcWdCcHqnrDR61pKrqaUhD2WeHAw2MkxH0fvglC+X1hyYRgNZ9ewDKZ6F4FmRy8
ZWPU+CVoXOfvUXORbIi6Qgg0fW/jNlygF3uOupz0iCpHadiQWNi3qXcWp8CUNBlf
vXFSpnAqQO3qbgpbL8p7MffxrSFRGHChhnniecFpxuq5ui9i+GTuCPnhRZ5afl9k
NXzGIdVamZoAYVrGArgCldHJdwZTi3heNbmR64P7xtJkdRoRoyeH1QvVWYemfjAl
eWyYlmO7ZSRtrAGAnSKJ8rHoS/AlMIZBKeI0LG6AtGewmAXtQ+ub5eO3EH/0f6+I
QOToVXqXEzyrD/6wWLUAPy2AM4fgnbNLL2SWeMJ2fIhrCprB8PYDQ4GjVoS5oWfK
1TsHWf8yOQYn92YN6zswoHaq8WQydY/UHwoWlcqpmgKnk7d4UIlghT3hXJdi/D+s
N6GWlDmuFwdCp0ew4DWXcarBGk6iFosnh5ufw5RX8/bP5RzXE8FWomb188LLwRqC
Euz6/IEKR2Jo79gzLgwhfXGlN4vIcG/9pj3mI2s5upAPu1IxPHcVPA7ALPkzdyc/
tzzvcVKbp2ScIq3ffRqhuia5FaBwrbzUhju/1tWug62XUYlvq+0f7kR+mNQHsO0j
3qyF5VyKqOXeUZtcdHWKXPKsoeyjsFCX5kNZlaLwJX/ivtxljW43+MQpT1lPGUCK
gab0vVuF+XsSymCAsTzZXownDNAlQFDvyjs9WDC3uLlBdYf72+2WCpySE7lhNRkp
2N/A1j+uavVfxYoo1vUAmhuvmJxnsi62tv13gk0aO05PrAlE/f3sy1GYa72tDB+9
npZQTZ+pzBMZzsbPfIJR/8HGXwxyeckWKT+uJj7iMwZB0MvW0pi16tmamGJhzu2K
8MLq9XIaN3R87d02XMLEN4ptyrxuM6iK/fb8xE5UFLc5kWIV1nlb9ZPUGP4XCQ2J
P7IIyeafV5vOobb9+yYpiIMzmr5L7GsPwr+cqLuIA/T9vdb6pXmNZvzUEG9w36aG
M76IPUXBo610ql3IVRZ1gjrfoz5RkY8bVPOVZiciB5/AWgkAhQ7aurIX0nI7fu5m
cFhk4XcFFgt6TBSh63X6OnsSWS3kwxDfw0PwsA4m1RiPRtwojxNWepNJaXMcW+9U
alkuZ6FVIdv7wakMdW+UNuQ4+KdxPTB+bKpqlMY4mLjX97y9h3NbVUl6so0iiOO0
WWK4XQCS1+Bwb764h/ghO0CWWkC467Z47WanpPhuMUrJrjQQg5RDHOzKpEu+7PrU
EClam4FdTmKfg954I0EPVzw8Qm26em7uW3UGr1KWalvVCb+rmktbinQMoH9tTUEd
Wnkp/3t74KUYg+aGBVlMu1loovPdDz/IKSFmGzhTcqDEMEZIPy5Ec5Aq0qwzenbM
Sf2E9v2ZXN+0e//27Ie2qdHeynv29k8zfTk7ZQAqNWuBupInmVQC/4l5JMaM+OcS
coqy7+qiA9Tr8u88+ShOtm3MmVSEOgk7Re6XwzG7+Hd2tsk8PQm3uH9fm9wMd1uU
3bauPN9HL3XUXT/FaEMOhOaTVihGu+rR5pb0uGjq60o4I1DAv68s32uUqC8+bGOD
K+K/pYDjBWdyl26x93MR1P1rvhV18M/b5WQ9d2LGf487957L30HRa1fo3t8lqznN
IXVTC5Nt3iJ7wUAMdgbiKpcLCJ/YfhvlCS/vCeqR/sfGg34SENOIUNwG8ZLz1roy
6+DkRWlnd6cxSUPXv6sOTcZc4guT+OBCklINGCSWA8QA9959774/PV/OvxJg3AhN
VSNCdMqOK3O1Np4gUygfwyev6pzDb07rkKxmmhWwMHBcg0+9XGyi+L6/kFDfH8GU
oSAAXfA3Ei2mzIJcKwuIaIGM96w3Dys29lWcq90iyL0Zeyo5oEzrnncxZZEgci1R
ZUUccsVr6Z6zivPaHEg7jC74UYmJSKTkpQHgnc3Aqk+aUCNdyZ98GXu2nnRvtVOE
DOhhQlIIPB6WNhvKCwsCXUlCkKpSRn1LClA0XSZOtymcV31feAoLKDQRGdEAlatl
3hDiXNXS6fZWQ5kRJ6w9BE5fTjV5drTnC1yir4jPhftsvLzqTu5hjHdkXqkCUKjJ
S1D5+MqD+1c93SIvzZUujcCBCz3trjFEinLVW6q9OrRwJbfAYQfm2cOcxUKZTmLN
bf+gVooVPwCH91lb/lJQmZxhjm/opys4Me7oGXl42LLRHjaAACdeRiNRPwUGoMDK
uVjs49cGdzDfYaKNfDLwA2Q3Xfp/iNHwlnRNXBFcYd/ZBlSoGdpVfHgHh4XiWICg
woLzCR7MHokVaPkiTfi64kHO9Z5jV/3pm6BUTMwmXbiPzwZv79IFnYgA6YgmDulX
Hsi0M5+nyVv8D1oVGLHe3MIHwaKXY4np/NlWg5LW5bk8EZKXhG2GfZrk8SC3BG/6
Ky2cr6CuAo8K2vo6FS7ejl0s+6MK6/Eo+hlV92eiEzun3O/Io5PUq0fr4FGIAReu
7RkzGRSh7MXHLjaqMa3BEwoA+E8LvuZ0bzo2VwkX0ylIrSGSGGCczOS8rpxeb1N9
930LDpGQNNPTAiaYAs9VzaNqbNLRvPKZaBKUbCX7SX7KZH53If+38he+FR1UeL8F
8xAVAf/JaQx6i+r1Lcu+E4rhe2V07j0cBV3fzXy9IXwM19AAFdZaiAN2Fdczjk86
B3hKqZZG5tjNiAAaTc41zjz72Ip10XKw32JFLoxwbqshZV7nZsxhNLgEpodT7+z1
dAnunLOq/mtbRQWSRBc9MG9EQVae90Sg49dySgG6ZF5er/KgBeigYncmSxNo7GYp
tGNJRfqHScxx+cUoV17x4wQ5BwUuYN9dFyFuJ7E+o78iGQsu8SCt7cxZxUXFFCbQ
Coeb8Wodtti6ND3t/zZIO5YE5DBiKgXb7svnUkLkO4hpFWBL3Ld9u4hat93X9BO9
W3JrQTUvhFzo+CouN9vlovY6PTqMfkJorQNT2GSSThAxvBXkpXLlpLehsmThfJQz
AWXOzwwvzDowgrh3O8ZuIMJwGOl9k26dwInUKOXKjtYDsm+UEFW8yJsIr1eQlzhf
rW82VWod4kPBvls7GSpKXpZtcgW4dhM/W4c4YhHKGn9Q70yn7z44ofo3E0o1o2GJ
zHM7xiUkzW/nmS6Yy68BR/N8XzCn0fhOsqZ/G91igmdjA7SFlc7eTWg2MwJm96ZF
mpTXJ++cfB/CFcHbIWzotpfHISka5SPoj+mEIHy/zwNPbOlXqBhuf6MqV+dLlz5O
MXK54Mkd/ugjYdmBGqA5hob/CmmMuGo3aKzzgx1HkIJwoVEy0yV/pfy5gT0790w9
ON/M7rRiQ0nlDc1A2OW/op9Gm7AkaNpWsn/j51laxfDJ8x7H5OAg2GxOhJymabQL
pfMYdL0KxAMNHQSpA+7ZNVPP3bhDEIvaXkfHYR1RAyI6i3f+5bF9AeMukyE40jKM
U3DDj1lpomvFRXWadYNQCz5m3AbOIcdYtCaoMlsdj8pMrbRE9ka95wlLlLWBhKFl
NbPqc37hzxTgT7+nnoFecyQuT6mglW5umCj5opm3WJnor9KejFipYPv497aRugZz
ryJb2AdaYs6AixIO18RpDxjsu6c7rZ6jwtKjstbA3mabUaY9bvWGtO5hbRHM8nSz
HVO3FbEWeeAK3Vumud4FRUOHhHScQy4SBmJDZ0bCClPYyE6s84FFlPB76d7jeBjj
bukEkEkoJpTXhCylBhheQL0y3DPYj6RGi8ZWifR9iWVAA4WLosdU6ISbn9qvXW6Y
FXEckzfmezv1ZSvYPiigQhhmav15AM5gfomMlmxsONmHmKj6m0+SZJlX9QeKfe0p
rjoc6AWdcBYEEHBCwJiEyX8qJ2gaP8sepQBfB0LSeh7vcJJkaM2OqsAKjRcZGiSL
l6t0DbOJrhdnes0mXQiyOIsWsZKvXHMVPAjvyZherFrDRBQh81bUthe67gSFZyOP
8Fx/sg1ko1DSc1CIq7VFQ2TFc4xYqKIZrsnHvTDACiNdrIMRbzUL6oHijol8Gad4
fSP+5Qo5M03CqXWtYPcIr0w9kvCweWfffpZqkN1acrZtPh7n2A1Tpj1FiIbLLNxy
c+SHgfWfDYtpAUwTWicmLpHup/R26KvBlCsyV44LipXGv54OHwmIwPg8M8K/EprL
KYdVuf8fyw+98dIjXi8wx3IOTZkoNw4T/auIO2Wp6RD56wD/kurp6s9XTecFCnb8
dSp3wwKuGeYKhQ+sB4/OFWTA7LFD4AIe7eantUAhXX7PwPV186wOf8/usWCdSxTE
r5QEpqTPniaS/eHB58tjhqghSGF/rxnrITB+basoX45TArf3ZFzm+ey1yGGYEnHU
eHfii2zgEJaYQ0X1t2nYG8KsvrqGWNNr2eofo1nNwL0DxzZ4ON3atJ9ctRHiA6Bv
5HeD5HE9zpAha/qrUx0nRKh4zUlCpIo0yfjdzhXKzZTnb0kwahfQeCE2McO+QCrm
uuwLModklLTzlBnr2y0j/M0fyttZp6BKP8ii5ej8vFMckCt7vRE8ytxTlrXDOjh/
3lujgEwWk3qC0Iydkv3UT2suMTdBfnni0x/yWzFJoG3XFkygjLE16OG8eHYtQzav
GxPyGEKiPPT1WuTA+j0YFCoED8KmrwDBoAhE+33fwe1J43c0BBKuthpO1wwgHSNZ
OKDkHZKMSyUy5ArniE1vcAEkeUd29dxbYiYSFU9aFjlrV33kwHBUvH8YU2yKGHxs
5mfUGENN6yLSqPEBMZ2Nj75YDONv+VzIgSM10qgS38L76xhpmt5/pfhYStzby4Xb
LKcuzMeuPKVEpROsrNimjQm1MSJUBW35Ar84q7+8AyXEeP/fjh4TUfD14Z2lebGl
6mJ+Q9MOjiRQPf2kDCy5xiypqohOPHXXgMGIJnM1fiI/lNaUmGFJSINmwRxE7VjZ
EyTEnnHC9HDZRCJqHyqb416kqoON2bRK6J+gaIaRlZ5pDGikykmqx2xSbZPAUEei
DTCi9yr/yc+EztcuAH0TqpsKvHi1h2Jy5qmhjAOhH+DkpIFEjIe7PtlpLnsMCEFE
+LFFU5RAzZ5GAmaKP+lDXdywkpRMMypUOlDi7AUv7Oza2ER/y8hGi1kWaMaVs7ss
nMWb6t3VdeaJfkJiQe9sVdUQgg4sFpUe1EZMrJCQH4fxFZlEi29e8Pm1ZQjCxlRv
ToHFiDQ04jWZoNJbDEfoprCtvgkM5amY5FmimmD9nvX+Zico3kWf3o+hlJdTSjPI
cZB8oF5G4b5yfIj1RbnRvSuYl0iPeEllkz9GoxvVcaXvVKs9Ww1ATkzQDyQXhb4E
7Jf98UK4jmzdBuPXjqDTBLVjQ15zpinZVA7WlCtatW2auMxhj6zeG6Snw3k1tK3F
8y+oRx/Ido0c0JBU3d08w7Z1uAoD45a0AVL+ZF2PhB+nvdgRuT5WpEOkCm2e6WYP
bL5+ZRc29BlFccZNPKSxtPwtJFeKXq+S5xsTLARyvN7HSj5rN6EXFjbf3BchBOpc
8qMFLPvJJI0TvoVGYXbILUdaxWxZzUSl69KkZrK1zJu53S+HOcRHXDXSl+duh0Yx
Nh6jM88k5hBs+WGq+f7BEv/pFei5WqTjGqCrHWSGAyAr0jtok/VWEtCbrVV5+FhH
elstoK/a/kUIZIEiA5lHmPDzwcoTWkM47e+iSz4uCinfbts958nmbPrQevfvWs9y
usCeRcdqJ0JFB40gMPdKhnCjvtdRo07r512Bheh4Hvw6CFRr1Wt6yErv/d8gV5U4
uJNQSlXetnTMLlOeeamTbgaISuPLp4QhfOQC6pWnsA3p5IDYH7sR2TeSTGFcWzx0
Lki7hm9kf/jZgjkwSiudJHWP0tt/g5QjFtmOpOi/bZXl3w5wBJk5jEaA8lFnaf6k
ewr6UNqPpxA8Kt+AskA/VE+Cjp2LmBA13q4CNZNnxHP14VQ+gmv1Be2Ve8fIepud
B+vQn2+veCsXrQ9v0smNm/4ySySjz90xQgFVHYSGj4ydnBBxMQ5F3P4YswXr2y1x
lo+EJoxMlFXi4MOpbru4d0kjDYSuq0xl6Yi7XTRcyBaMo7nlIzM0nG7aepeJ3Z4o
RlTs8Qq65it6MrvvC6HKLEyQBo6sYuRzcV+YZP/+apgqgEKDCW4cz1XDnwJas7xX
Uso4ZiP2RYXSgDVCqUaoBtHz4QihmXTGHj3y3AHCz6e2TSOYDIFxbUifldRHLVBG
qZpKM5DDAwI9TF0C5lr2XLzNssBi19otQ7DgFbgss898guPYC4M6e9WfQZ1MA22S
D8akrhhdesWJJfapq6mbJCO7Py1iU8frwsC4g72Im1LwzbOVv3ofnGEEPomsTM+T
oGXHjgOgl4OaE2zKkQD9FRj5T7B87GNhmPv7vXQ24RJ2Cx3LrU6m8wNPeN9N1fqD
kOzf/hGIyto0eEGmFRkMY+ykPy8E4AseJmHiYklEZGoL9oc+X0hiOhn6BKiwhszs
iKM+h+FDpVcd6ZQXHhyr8qZ4FTdgvzT7G4Zqx2lbb+reK/jBkRdfCIR71PUchaDz
LDwVIa2JS3uOx4TIqtYIP/OeZF97ij84t2Rt80KDJFLLos2B7XBikhuWBa7jEn/B
oq2oZD8V7QPn4eQqKRCxGrrvI4YHxro9lCm9Pq0HCewaT0voGepBLUNH9sW/mXLN
KrCGCuiDB6AXPCnEiDwpS4oziZW+E6adavJQx+dvzDQbl3AL3oGiXB5CLYGLc90K
6Uy1O/81iBo3TBnLSN5MUEMy36VcwMsaLNzSihD2DdT1kqrxNIHg4ElujC/igNmU
fss3SfMTp3vH6l79ITSQNwl9B1EygDQu+cSi+pOxwe0LRJaVsMMwxIC59lRubfJu
c4VZXx4AiFK1vLxyouptPq7WjQhqiNRAo78BlGisa0cPcuJ1QG0oHUZU+lqy4J3V
IFOdCV8xRl9XRGmlQYYcLyT3kKBjPLSIOtzB6xWaHjydvvZnwiD+upe+iyML1t+f
5UWjAwhVFRcZU0AOc/1S4nBtMwuN7kkCBnfrQuwPJQb4o2K5RfXMevRqrSp4Duiz
IEqvzc4InFa7mSfH8tBqapeEOY4KqEo/LxS8gEq2XnXoV17IzDFJtkfw0D5gAyJ8
5Zu5WbDDycaUysFJ/UhDCgjyveK/J9FroR8BRxZQRehGqcQJTXM9O6gc7zi54aTN
jEkeyNXOCforKvSD+k3re/8tmE59VNW1lBGNk/YEsXIQbobe5J9JvvQ3FjQ9qn3p
C8JFMGV3JeA7sKtTBKo1RBb7EznulWqLZHmTO5PtrnFxeimK0XZ3XRXvc3eojzBF
ALG/SdVcKeXKNBR45qNP8S/n637X6xXADKUhS3OKktxq3EMlZzJ30KBNRkrOPNAD
PTmh9RSD1dqBhOyELFSHat7euie24SGu10byOmBXabicmhSL7bM7LasFUVyFFMke
8joKvTOC/+Pk7YqH4f+uZDnxIEFqMOl2e7P9RzAcq7EmJNxnbQJHbKwPmrhrDULq
prnwAJLuf4wyEd3ELUImACkHgRpueSb1Gf1r8c5OqiRPxCV9EPnZPCBfVsOlyMvY
YtOqL0NKhqxBPfxSkfol6X/Uc7ZUyTi+86lCZrNFQGy+kC0S71xCyGTL+aMHJhnA
gvLtamhy1iiOBQycX6cg9zKDXPDtY2k4DCuuWpiUEnq7VmPBN4azCMbVsYmYU/rj
oLAPNQGGpaYbK+hVR238RxB/QPRQ6pSlbrIvIzCDJWyzIZYgbJFjNcq4ZEYtkp6Y
6Qb3DJusx6atgffyf8IpPvXW8tuV9C7mcBsEdVJxq+xJkJY+/CnQbk6duRKuDDly
tm9SOGBYxY9Ief6sWr+op/YcUWJng10m+QIB62l0N+Yet92F812mPdKkSAL4dOyF
aeW9EcN1XmPchz032YyKnn4lZYq19UTkyMoVZuWj+0hqtsDbXmka4/FZ3SdqkGT5
0huRzSk47zoLmRFarYMK3UCCGQ6p59wAV/9lDNpx4PdE920EFtbzGFLFqE05qHm8
2bftfhsTEVqBniSE0QsTi8c4Ug543kiwBfiCYRpV7saBGS9m98vrs/WYqyj3Tngn
0i4q/fzekOTdLbF4qQDsDJGoM63BHznMZAcMMXC7fGRwJ+ApjPUhz1hFbRD9bKUq
vHUa6NSWua2ER25jPBIIcO/E10nMQNmq7j+c75JJuWoTZQe8X5IGODdA/bq5FHkN
cKEYA4JmJsubd7r7TpAVeAyGN6NLNqePxlBuBmjjfetOnh3gLJa6Q+qUJCdbLIXd
rmvJxS48wsGG1HroD/HF6mfgA/G1GGcBS+nLQHSdetfzUZAwHFcEltxYYnnMD6Dq
cLk3yJoSb4YXHgL+9V9bZDmLZhm347TVMBx0fLVLuA4HgamhSqSUY59t3HNXQ3mZ
3DRSqnFQ+khijqDrn39YHhdMSCaZACZDGbX1apA6p6IBTS0Aqhey5YA+kaH94dY2
hxcRj6rYsazNIhJ90FFSbYF5xsNV0A+BpewZFjUtL9PC0PmU8wlamGhTR97R+ic0
oak7qgfKCTzDX8hoQNUeRSl1LRHR952IOSGKPjDPowzp8IfO4JPPjZimQonTHZ2J
mEteozHSmxoBWySMyhbJT78FNkml0hCbAcw9qxY4VsaLUja7ip7GsS7MxzUfQ2u6
KLxGUmAl0hkM95B6f6EQ0FVq8uzkoxti0heWQPgulVbOHo9+EBSkgCKL3nvek0Yb
g8YWqezAUfa2Sb73MWo38q7etvMiA6ujagbxhkJM4/ehE4aN6IHT4Ky4lNE+1zHE
rlo21KWBpEHH8Yrt7fyASrPpEBTVLrztb4nXHlEq7CDLrhIqZ0BH5cyc0dtQSqFs
B7JBhQT+HEhjvgLBw6s/X923vpWKrDGU97ytXd0G4bSwS+dJCb4rR116i0Zm4grm
vf0Ca8GMXegdNo3UXd0AqQDPUzE9mdHWY+iz06M8KgB9cBmVrL3gH/VOvHS75or5
SEQ3KhreyfWwd8g6ajD9k5YEBCPMklyh3k/1y2QnpBDtC2LWPiAPJngL2uJJJPou
FTLbrkFkII6+yY70yWLaVGBXEofNuz7r5kTG4q4GfFwDZb0syLd0Rrh15WDJ4O+E
XIWVEdVPSvou29xNtk/Vyb9WQGc4lQwrrbnRZyuJEMC/Y4W+WSbE2EELpNHTB5nX
c68az+rWB1PlZ82k+kED6CiGNvgjELAySwZrC2IlVJ0/wHtPqIQVs+Vjk/2u8ko9
nf3djO3pbEEcYjMegh1ZDWshSp+y7/wjCkqmv5zdNPwgFo5cwGFaI4+tadve+Uj9
Op2O/Y4Nh2Lg3sxK0nZF1uaAGMPUzIcGWgTqxEukVBj9QGuboJYBR+/ABjwilNNS
smdU+bfnNMXt23sRkjJeSVNMWhoRABCx+jRUnoVjpWRR2aNPIjx1BFLFoR6ZcP0k
WEgt6I4W0J0xRYTuCkMkXTBYGQWC4A9ClNqAS5aK4edd72qR8kSvWjeG17/dJe8O
r363suV4BG5c8ahaVoXcVBJOqoGvBnsLXplXVSbFAbtB3Tz5tUyFsJPP/kVcOJX0
RzPuN4OZ2ZcL6Tk2YIiUzhbtNeXXeVjwWotYJTqPMzObY3c2uZNojklg2LqGT4bB
KKAYjKJUf4phEg6xAo+jnB8FHhHpaPAYUJnHbQ0CfiE4E+9HhoTGRvdWUW4z5uRc
7/Vmj5bkZqVjGuEa8ORQnNUsGt40QH1IzilzNhsYYwhwCSStvI6aRCqZg1hlMvc7
BhkpdURSRPa9nJKSOtt3O2cjflW6IC3a8roycbUafXxbBsQLcY6MqnhiltxVdbgH
Caoe/b087O6jzPsO9UKluRfZGykRZT/YacwATdbMaeBWGwlPMnng5oSs7Dz3JGWR
1FE2SuZ8k3NBH8tsn0erHVKIMUHPzB2JGpr0JaZmS6GgMhOw7el20zUDDDLT5GOK
HXR0W0kJag6lfdL1LIaA0VYk6oLpuUjSZ9bJvKVtdwpEi+HW8Qm2zKtE5e0etqqw
nCbudCLwmi5zphK0UUlAbQJkl5O36kgTNRHohP1BgbHHyiX0sfyUMWRq+VWjCzc1
HJ1dL/Dj7P31E3OzDTGZnIDpT9B7iOYx0P40NOF5iZKIygodS3vY8UlPJnI3n8H6
fpNpj4lTUbqe63g3ofcdBNHuE2h+IQ0cAVFZevsI778gv5fDqnGgSqOm9Rrwczf+
lJYCUkQxFWCzNCZxnGfn/iBQ2FYgcwKyysa52ZRTKqSb33m2jGCPH26JzfMQDgSG
eA/OjP2cTgs3mLRaBDjTbptZaZSYjIDroE+zlO3kbJyuFdWDA61IlFH+bYgnNNGx
Oz4I0zpe0HrCTp96cyLOkfuV/GFikH/YqUw7co/Vz/qFL0RVZRlfeNuSjf6g/cpC
Z2RLC7yLVqH/oMG+pbiHaBfm68HZ9DUaPcjVj3Pf3UeGOGxpu6L71pVAVsMEpPr0
4AuXHFzUfNcKexdRkry7Dzb8eNyjBZE5WhB2lYbH5d84MxYytHQATac3ADSkGiHz
I7lrPtzPlqDxn9xP6ByCDNnoI69JhnDGz0GMbHyTfDJaGDP+WTd4YkqQJBI7ZNq4
NqwF1zOFUQ0Cfnl6REgL/em8ZBrXDwM9blKq79d+WigRKZmnjPsmAGaYQeiKG2f3
SA4v/73kI0omC5A6auyQ9JRsCAP3sSTA/wf+tIOM3zu+0TTRq6Tb4yQFmwnN3rg9
R2h6ogIIkXlWKya9jtOnV5eJXQ6Ar+OdVEHMgeSXf1yQ9WVRwDWK9wbS0g3lgRLx
raotoIT67FC33QGyR7/SWQXFXn7RwhRS1jctYrodibMeyosFsisyOsxw7qyd/Apz
WBSLVDpCPfQRzJf8EIL3ekWLxD1HhV6WJePoyropQ1O+fHKaXcLAFEcYn5I75659
SnvE8T4QSa+u7Jite3YVcO8P90ASvH187C+plhUqmXxQNspFFD/lU3adZLUPo2Sq
6p8mPtX7rPqLbXIV5rnu4Woseb74nTeHA4Pj+6/W9qKsrQymQDdtDYGliEYkjBzA
PXqSS5jD3LAZ3EQP7N9ifc9Hw+/Ik4BshWEPZzdApllc8XzXh7MPBZCJvuwakuRW
KF1m+E1R2rPfc3qoPO5JgJYNaoCGUlaZoY3t7JjWhjfep10m5TshTQKHjkgVhXDo
VnybiH5lGVz/DRNJNKEGPnYZYUY1ouCPe29NZCKnnhm+ZdiMf8v2pUH3RWOmkmFS
xyvcLy3tMPpsPwl/5xj8QrM9QANJkv6FOXMOqNOs9HioRE2ZrMJt6c1ufHDl5QE5
QZ4RDKZIoVaQWOCqtbRQ2t9+SLSiPx2GuRa7ZbIvaU3IP1k9Z9HFAK3+ouH2jcoR
To8t88vWdGQ1i19ZEPtw36s+hIIk4HbBgEw/D8B4eawe3Bkwr+NcK7+39rLTki9A
Cf8hbWEF6VPUbF75rNorVg6QTYkhOxk57LWkIhYCPbjwfldxa+zbi6pebEG5vpOZ
yG7i9+yGOUY/0rpxmLeg9OqYhCECsS4IrNdo9cezb1Dpn0U/WNrv6NJdmIlq//AT
EMsdcZ10kQjYs97gR+oSPcU6vkTxXXFiXuZTtdhE+e5sUI0e2xSEK9ycUw+FJkKE
I/qGwhAsVS/FdXDXYJ4c2zaz5cADXsN6ncf7xkFKWEh5998XuVH1e/BprEhYQljS
gVv++hWy3QcV3eZ3GSxUvZOMKIRNnrlq/cV2lT3/iou1gROpPA+NmpeJ3Lfd96GY
FvML6HSIXaf8ezmH7rZT0fQHJi6Vw7ILy8L3Y1h4wZz/06UcqrqOGhsX0Ay0tN5r
cXUwu5eCRRsw2Ah2zCqUhI8ex+x/la1ZaJacAN9Gr4NR15AvhAlOyCUml3V7L7zV
5793FhMdnOpTa4HyYr4YOIUtyTT+Y2P5YtroopbdyDsATHawdSuakakLXFcwQLlW
eIoCXrfyv6/+5Bbb8wgqIesJ93702dt0nntkunVeG63awVuuNM3GoUFArq9EGRbD
S9ezFF8Jp9q5c1MPNehkXuUvLnxHVTNJ55NxwnoIaz2ZkpKtJrNE2Uhxao/wYsXw
bezDNCjhcOFT/P1duwcnDKzURBrr6aAZM0G3dUF6XWrQZBYZOXOkVBPIbzAwt28J
z9cbRpZScMFvhkW5I6eGl1pjTj+xTSmxOcvbKxUj36KwPoMiQbsqT7fClESOaoJ4
heomwWdkeFZOD9vAXJFPoR4hXXYTTzWNN6WAeDSD63TUJHLllkVRsELl20Dl/Oih
w/ezkZcZuSzXoLCGk8jvW+NxaV6THkoqS7fHiCZUEvwDWAaIfhe4s4HUR+ohfz1m
MM7xUPk5yRcZqdyE7FgxlEh9uMugnVAi/QdgrS/3mgGDqXIprAbgD1BUmJfeCZ/X
NJ1OJZ1ENnTmU7saKoBN4zAjjQXZneTP4vxqJiFrjGxyRGmq8lQELuo+C8lHObM/
OrhoP12DSlPIrucR5muPRXqM3joQaUfi4P1jb1VPsKtAm9erSB5vx9sAD25dN1I7
AikTKU7d5scZYAPfcBkO9doanUpmq54DHZk8x4NtpDa5vAAbcWKrp+qQdHNmkHi+
X9U5NXOhqc+5t9BYmiYX1LhC6AIB0E9QbT1+c6ee9yeghWY6zLAvsY9wmNKSh41C
5QNiqBUvaEEF0iNMQHdXCsoPQtSMxos2iV6rNphrggvQONuQctDI2SyB4ZfPnwkw
U8dyyoEwanFph5PeAhzNeugxcj9/nr7VVzdabdmFsy8fY1f9igPwwow4dU/CUtCI
TpkMjYbEemAcRbtibc1vrOvUQAVapdNOW7aS/rFElWCWNcYN9yjqhCOmpJyb5Svw
4nTI9UDUTm1qmyO6HGw9+5mdSFD05TA1Bml3JtIE/wHFUONP6ecj3omFCgtj+RBH
0Zusb451iz53L3N7UQ/XEVIxjVHqCVnqmjiKFGnyE8A+wpBhHY/Y3LvNKkLBkjBj
aQ/UwXWb+D3A/bLWGFeMnD+UiaPz7M4CPN6N0nOX3yFq7BQ+7z+twdfR09NdRdJB
Hxdyq2CC/9ITxMy+2Qbi6gK60fZWAuBUQ887UbScQ+lCeISYx4hhCjtkGtKr0YTR
+CuQ2jB4iBQFdBYYcb+7P9sXVTLQlZ5CQJqdaqCwHIy7+0WTT2pK/G22rdavrxFb
nknGUsVFy3crNOZ8CiKDBLnWcTPNgpDSz7nh0aQlY/M3rJ1OlHjXMt3myGagPuCU
PR4ezBg84dsLCvlCOkPiExMlfiIIXxwyXO52d2BZOO612LwDRLGIGBxic2gcum8u
6/EVWT0sLS4CKDqa5gpuMViaaawDQd0VFnqbLdT6KoW1vxXiR7mdUUUuNUB/CSTW
e4bROUEoPXzsVk9Z1RLzbsyZlO0uyUtmepOalg02sZeJb7sI9meKqQ6o5v0eERkL
vB8TyivolxXZ/HgFUsfJsBtOeLjnwI3B66ZSulisIehXvDIqmbFWYJg7737+JgrX
eEcFFcsC3MyThcNiaIc/h8HDkbj8L2HfCbStTVZc6K65vSYZ7Hjz7YcVCUiSx5p8
beZeglqUCJ8K9l7xFZ6mZRyekd658dBqEo/Yf7HJ3XmW+RN5AdbtQzkPTHNfNJTd
9wg9XjIc8iOpvFcIMSYQGy5m0QUL8Oiz+K7qaccEFgCtlj6Njfk/Uswz8UMLWwDC
URskdHc5RW+cB8YMYCVxOXqR61HcksWO4EteuLRiLdExwRp0qwLxcJtoI6TYKsiA
Hbvzb3oAdIxp2eSl/IxHMryLHMuUIvNd+Mb9mmTqsxi61HPyMZi/COmvBbTEybCL
A3DlGgT/+NHR3EnVkBsVAcBz0AnoSxePHoB3go6lBtj3fe3Z+sp+GM3L5PSdKCsg
3lBpwhSPIAvKhNUrIxJTYyFtIV+vLIQ9K3s3eTj5+RNWKERL9IpUncRe3026M+Gl
iW5B8nEjbs35ZR7d4iFh362rjt5I84L17KS+QtJttdx/U5rCxUp4j6bsUFXnIfsE
lpGJn1+yZ4YsEyTeg5zwJxPc/7ITWeL9PEvHGjYc0+QgWCm3QkNyjJg97uTUJP7S
Mn7csyONugdz/E6q1nyNU83IZ21ECdi22rWpxOMeAhc9ufzkcOCehhh3JQMK7x9F
GkAdLbGJy/Bfv3RZMkYc7KAAwrqlbkZR2cId7s2rM6B5Hx+mL1n7vHEOIJiNd8sm
zDT6jDm1uZznWMCJLCVz5nSTTVmTpk6Vhlqi8xqOS0GgTpk1gp3ledo7y7Gul0me
Xl2UDdIRlc2XYqLcTjpTmf76indPxOjOI5vYdkMSaQK2D8m0/IcJy6kkQOKeZqvV
K+fFgKj4mLglgbURW/xgwyrgWAGcGAI9PGXwEEN+behK2LEh4kYl6cK7Qt1t0fLy
Ajv/EPiTg/Qrvw7Fs7MbPDJ+zIMQJlKCLT5nwuHIUej+6+bRtMRhu0YwA5X44sJ7
bnEhXYmBv7ChdfSUQa/vmQSNSweO7s5bpKN9AbP/Z7BENGxYFKlpvBI1rITQnlnm
Vn1EaZOlzd/gjeL9QInwpPsijbSjKqIKB4aZh0IjDW0ytspbakCriR7LLsAb6E6z
eQuC+hMqDKo0vkZxKkQECsvHRO2ITYF3bcgbvjFR3YjN6yMvp5hy/oA5emFK2ucn
59iH18zHE5TtF2P/5MBIAJHzYGp9MoUMMQYH0LhJ51nWe/EeptUHHONLMtkso87s
Gt5g/F1WOF6v6fcrBAX4ZmRCU5Ks5te5KR5jstz4EPufT7aR0SzDKBhK2GDcjOE6
xnJaE+LbqpQRRtxUtwpeWrMYw5Ywp9x1PVmfBsk6DevgtMz6dO1gUdmkDaabC6tU
PTfmqzSKZ3NSdsWg/qP+DEpsZP6gtbviYH4b3pysvUNA4ZgHm6PBFEPLiDeJvzn8
7rixTkmOeb5bvyL5+/gJNLDePtbmeHyvVQgcHCljiVRiewFZACsxi2EwRUbTIFrS
1Qa0YbjTbjo0Pp9LMxpU/vt9XcrOAKRwvwnGzbHXXH5Thn4ZjlWvZvqCUHZstqdo
nMieDnm9hrMdfOgCIEgpuHA/MVRXonXlZ8wG7Q7GI3eZI4dVFsOuOTC054a+bAo2
84imkxKKcUwkwSfLCmqGElxViXiuBz4SbfY6M30Ajp9/CqMQla7K6S9RvkkVj7za
7FLiTMqwNrPWJhPdN/n7pRGyvoMJvh6Yy3mafae0sm924wt42ZiozNH25VVHcKpe
QpJA04bLux/44tFLn4PQPQzhJW6iqpwHqPns12JRi6AVu0pKIL11zOruS+SIVRNR
j7bLbD95hX8/eC83cSpkKMlTjRCNMzsGRuj5X96k8tig9bHEeBhOgukr4WA3zr2p
/NP4ypvRe8mt70+kPHIWvvFspzgCxbINGVlwqgxx7p1wLJcEkbQx8CmAx0QYrqRS
BJ/DWSPzpbR9IkMsaiqi5lAZ/Qm7kSQZr2arq9WX9GmFwgARxTtT0zp5e6HkeGu6
1vTmUKg6PO/cWmN3Q4MRZrJMQyu1AdlMSCKvh6eitdQe6u7yAwSc3v3CfqFpPci0
ewkkTHDg0Ex0wwMvxU/qgxPrYmp3hktbs1oyF6agjlKroTKmMSwNOUpMOwij3t2E
ApWpv3QWlyfxsJr8Lv6h3DV+PxbQQYm3DeVtkEQtAp+kzm6Prx1LSrIi+5QRrCGi
LiN5ul8qs2V6lPBTOJazIrT4zW7aPPN6Y4UYRZX3KoBUqImCWCYaPgTT1ww7LhjY
sa0WpA+FiS1LCH6AiKuRDxEGBP03rWA+3o+59oDtj477nro0iAxU6ceaXF1MRoQC
z6gm5St0CYiLQUz1tfCbMD1XgIkuNhj4gDLJbCJQmfBn/+jaY8rJ7f9WbMzdtxRV
/z3+ayKmDF/UtjlyEPgoWneyDHqcHiwXeDAorQX7uC21QnwRvnJQ5knUpPg+83iM
QX4Kychn2/xuMppkJ8TN0SRmkLXJRNjh30XmSvXTl4TZR+8Z/QyORiWe9IEpfSnv
/PzM1ftTH0lBl6cDpVwnP8ZWkKgenB7GEwjN8SMRSKoIvP6NPMz1+z0m3oZV6oxu
KvcWIl5QugS4eLDgatgdBJhuQoWgGT8HHemMG92vTFGbmzIbf/e6Y8VKZwOp3sLq
HNz8LMAomFQQGx09G5lf+/TWJ7CBnKA/URlWFo40yNi0TxolSktLT5jIrQzJmLfC
J8PN23/yfl35KBCUsEPyO4wvlynNCwjl24RX6fLmXnmru6DitsThaAyR3MIY08to
G1iCAi4mt5bNunQ0FPiJPn/QC5JKrZslkO+IajXtrH9eiyjhDZlfQZqWJZQaYpgI
RwxIW7lqjXGsRBBfoJznc6HiNp7D1DFpI6U8GkkFuo8GB9bBItIKjxojTfDas/Gv
RWOOlZ0dPuGA77UAo13ylJb40wUYBjt5cP42yLWfpNH/cnjxNLfZr9CdR4/uRMzP
Xiwc6iyt9YWDBEFTzTA94bc30o4ClPzsNkICoIpD8UM2zeN09fvzLZMVie9tR6I+
HcdziiNI18JdoG8HAG3kUW61j9XZUYqad5F0djTs/0n5UbC/p9dptbWoZYH658+s
GzZV7d7FmMQhGSmWDzpov7OI1j7OXSCAebSq88D93FIGmd9k3jqyghqKhp8U0ueE
rbCagvRIQn43ojQDJJjrkyDYTZf9sPTufVn9oc5HM/04NSF68Omb5a0D8M4OnWVB
oLnq3L9Dm8HI+j2IqCq3GOWd/5tK+CuybZmI2T5lCbzal5a09/fvq4oTjHIRpcMY
XcUWlrk7sE52SlKiXZkJIEAfyB+SQAKqh7x/IXwBcudq3XM31C+c8HOq3FpOrmxL
4R2+Ors+oKBtrddQiPvfuI2VRb4GuJrDQy5FWrJEAz0TCPoAQYugD6HGlH6ACHeG
vYeEodbazS9sUKx1Ih9YiZUxnKVgFMd+JfcMw520q1wgXgWcUCV4FlNZkhREy55i
PIY0IU4N685L6CiCv1POt30Kte8gmwkea4PB8OskSQMZ0dRBNuSC+YIf+aBJrndd
TwWIgJHxe/fs/BColzOaiDhU2C0No5DlWW5pdBIvygp8Rg0rqHNuyukdyQ9Awcvt
N25MlzYDZVzZsYPz0jhltuBWaaW31Zlx54cBCulYrFE2NkILM/e1RpWbcWiZN452
y6ZRuo/TFOhtiP0D7zzla/PEUvwTyI6+z5KiX9CLmCeDO/Zgi21HxTTkBADUo9pb
Czno1+Wa7C+6FyJINpDbuyrz7U/Ey7IsuGI2EefyY8MjH3Q9AIpLsTX3CXd9Rcxp
4zPKOFcK4Op65PPIjEWoAyn9pbCqNUMLYPtqrPnF67O0Pvc+CdpPrHbDUR3yAY6M
LyT4Lum4RulFEEzcAOm2ZyVKTs+s63fZMf2PY2YV2wo+lqevL6lUR2Z3ChQ4s4Nk
v409fM3I7aPNgXVJmiDnLjtmyvHw5s1n1LnCHzzFxW8lfBF52MPWqq+M6qUCxHNZ
HCGrgvtfPb7SLIlcYeyfStktfUso8noF9907EZkF/SUS4o/yUoIglMcRsRtwP+BB
jqWM3x384yiM2edkvfiSpt2WeLcfFrgl1iMBt3ArtagA7YAPvFg6UoHDS4c7GsEc
23nL0UhWEbzxq6Eek8EOkvcPJ8VxNs2JV6v5R7Mosd3dHJpMPsjKgHum8pda5jWk
gWxT4tAMKc7qaKzK/sQWLW8YEcNjDmJnfkfj3tD76o2XDVhAUk8X2IAxhmFHX+Nq
RryCxIH3jRVHCGxI9t93ZO0xplnlRkryOr/4B0UQ1jHfXyIFctra4PnXRhxC3DIs
pdgqMmwtUNAWznEj27qoS06sjoX1kHl8kzi0IZcgIHhK1643qxnE9RLc8dlQ122n
UTMWrEvdhHPKRexJST5H5vcV5pZFUJ8ottdeNqZZOoVdxBkeeOBJm2mOm8FUmvax
IoNWhHTFbsxK4dKEr1eMdW5K8kzORIpzHoKDiqKdKgeMQA8embCpj92PQSKmF1xW
reHNSAQrS+34rO57yIhmyiO2Nn6CUS1VpnA4pH6c4e5l9QyyjYb4MOsLCC9txLt6
nf+xgJjmzswIYNt/Hb5aLPgvtYG/ytvoiZ/XiCv5gideZ+QPFOe0uR+13me10uFy
BmCTjYikbMN7113pBJe1g40jbrrlLnI9a3ny5Q3BIMZMjDWIHuE9eB29r3usO/8U
mFbB7h7Qg20QvlzeCfLjtfEz7r+6AtwhMs7lYSXPsmb5kFNUz56n2V0X9KZ2zLyy
pLZwx/wPFsl0qYDWnizko/Tuz+CWUbdkh8iSHrH8+iLskg8FUNe9X2zkRsXch+xv
r5gxJr0H2g81jHpIQycmr5Sk2szsrPB1l0RkaQ7QJADvRqzpjsX6Fc/RfNAbwNYN
E0LoV5ms21HDYKczPNHCJuPHM8p4GcjorhEFc8jes/gCRpSR3ie5z51QivW7DTLM
KZjJ1JO7GWLQMBkP/VvsdHtuWqcVP57CKcWmUthmyCdb8lcFEtzD1uzNb1KX6j7M
PKQMj6IdL3/sns+stSRWXRhSIZ/NPr8ubMAW5VYP3pVDvqM9uZyNx8CIrjCj5ElN
10avg3LHtuXw2TptgsYekh07Qn2+qlNzobeXkA+xe+jnEI2xDQdMRzTu7Fa6Jsg/
9eSPWJKdHrgpCGOQNWvjelWLFZqpwyDhzZ1Dqv0FM12O3l6m7fcZps7mx0HxETB1
r8Ve/gfXFOAn4o1SsUAQvD0mHxuGp65V2QNoGlpa7RMtOdsRA9kKB2f4Rxcqx6nU
3IC1CxWun7/DTxD6OqMbATcyPiXZFtxfCqTlF+QbbixX/AV+WoyVgadguSU2SdWP
Uq2qb9UBTsA9U3Jwq8k9gUmQBH6g23+KyKJ5UiHzCiIQtgydgNdDkpAnU2lwsKr5
Sg/Qs88Ryoe6p/qdUkQyVNeRQWfPUHUqXCfJNwc8flWzjoRuBnhRxwN5WI+dYV/h
Yr9VNupMg07AVl/AxDxtNdCBL4sNYfM/76T/HoTxr98wEDbm5i2oEI3BWrq0WlbK
Gz7TU1BuQl+lsemlnoCLqaTjDd9aUg7mBsjasYYN/rGxKCa0u+B6WbhM57o3nxeG
NYQD9ldM6Lgkcpq2qWS7Z3YXnozFrY6JPtQc4USMocuKQLI8lwJRK/oaB0rMr8Gi
lbftzqd+NKFjEF2EWqcvhnJT9VBwUhpjUftX3mLc6/mZAs4T4dND40DLMXoI18fk
8Ru4jJ6N+4eh0Qjx8CnyNwscM7faDBjSqaR4dOpMj56EFgj4FX1rzqBTs7tAd3cY
xCW3VyjZSwtSzeRqI6C+7YV8wE8o0XHjGDYzBTw6Touw943T5ImR5ovIle5J4rvb
gO7E0uIJZLzCACMLWK7YD/08u5fQLgDsLquI62GVJb9t6jZG8Ab+3xgdRGK9zsOF
d4STVftuv8NlSwDyzfCG1dU7zaYorUkaC7Is7sCn2Wb06dUvGDITwRaiV4jvVvlr
8Nl2Eezy+YSI12nQ9txdDhukvqKmZOMRbWk26ji+X1tmboX1QNmS849kmGxd2m+8
4c1DRvSZ8Qdc/jiDJpmuHYtk8b3yNmeBTo91Iyh29m0CLDiM7u9yKmzC0y1cmbtf
k0wX+PcT/ifk/yavYEijtGonLcpgx23c10+RcHvFE1dF2bh1U21390f+XHhIEwh/
cJdJwzNlRqLt9E4t68/PgdWreOWGQjGlstzlScT5o9omM8vKhP8c/eQXHNH7pBgP
jstNqZsjtHSGUAknY2uuKTDZYjihA9Z5HUbX99aSFqzAf1GR23KlBSQbAGgjuD7D
jzZEoaAapon06h7Lbab0+DF0eEZ08IY1RTWPbPj5EJko1O7fs3VTvdvIGpGaZxqp
m8DQgv1yXPi8b9PPm3CZcGjqCfF/2/0ivPD2/rCqaJnAKZaapU1ZfTRtafJKaRvZ
h/fsuoHZdzI2roshl3/XDM01Bnjo2dYk/oFaHkKc0HpNDi/PlNnyckLHKaKuRLBZ
jrmotRBU3ZR55Aq8h4OFT0lMwJE/uVXkw6OMenHoU9L0RY7+64Qy6+3K+1LRW5Y5
SmT9fwoqdmX6GUfl6jOPRm/EQngo1Mo2cB9EeZ11OnF9g6xYjXU3GSbRZFdjpGtC
VgWWf71oY1wRzLItM1qPCtRahOiCNuYeboiNUtKpRyy6QU6E9XCleGbuXhPLZvJa
FShcsXT9Zpd3E1iO0KNumQ4KyoRiWFtaaDHqlKAOYamhnX/jER7/PpRsJwQWS7F5
u4+5jMV2TqdXpFBSoarzQz3c60rbQivOhplfC06QV0VodiA64ogLhfWpVFg5pHDk
WD5Q3q5t8Xmc9BZUdBt37P4Yi7omyrX0QXeZpOb8BTfo6v2UHXhnVrtAF52XwW8V
luCurWtLpf47D8V3DWG4ZJFg1AHlf/VTsc1iYUBxTRaRC2q0A8+rO0fTPJa3weQg
dD0MlruSgNfWGn9DzqRHwTFRPhDGFoi9bAmVoMiCTulNlupYvOQxwooUXwJ8G2o4
yxOA7bEosWoCRGBNnsOIzwnyGEx1yRALGMWHj1nMsqQN98NHcveP7btjOkEVBbC1
8HGTT8xgh+VbXtjzpghrF1l0NAO3oHQ5PXECe0wGEs35h2uUo3HnNoRLz9W7Zmw2
Z1yfPF8u5+0Wwg9H3Ac9nQkuQrQ1SGmWu1AzX6IWx5Ro5Dew6RogaFxCW9ChriPM
9EpZTzKPujipEnJ95y7U8yMKvYGGYBsqQxL5gaD/SwKDVyvjFAUo4MV161K+t4eg
QQGLRn9b/tCwp0eS8mZ7UqPNBs05SLET1XzOgiJU/sCI7ckb3/uPY4O9LxmBOQGD
+Ji5HkjhtCv9brh64hMEcXhmqUMrxjPvmAbXOillrksazzpo+1oVTpxSAi0hSbqK
PUsvCXkLTJ7rUAYdwCd3zgaoYWg//Xd1OoT3OjcEI13ivURCBQcPuw5YjxAFdN1d
0j6c+JxgxRPXtuvoJR728It3CIEvzYy5QDSAAOfX7RYdGzqPaNRwNBg5vOvSZw94
Uec3mFcjTH10n1+H9oBtKMoshIbMq/KId8WJyU9Hr/kRdaqvlFv2rbLl67XCQ8bw
ngjnMFOdVZNP39NVneWCta2sNhj6szfj9wz5Sim5ZRr47nYAggqyuX+3Y5bVYbMr
qBiiqyJ0AKv3ZHviWwUutgkB+dduVGc7YaOnpFWqXZAZ5YiqsbeqzLg+OrUMqeW0
CzxzpKJUkkavsvLNJyh5t3SBHCHCf9W6rriREEDokIrrczSa2lFAnAwRwfoUL4P2
n3JfRvvTnFZmAHnwT6Y/98SzQ57rAzfnrFgKGO2gQQrR9wz/2fW0uyr/iISE2wi1
V1qekpqADJVn/FWqQg5wGFvac90sHuHlBGRXs4uLMCVXZxSxWUaPL0Te6j7PUZRl
w1WoB618DY+1ZKd3ftAo7wdtTgSiJdKwhHC4I5kEwoYNOyaqNdxS5HWv2WYjyeGp
98Z6w+QDtYOvSFQFbLXgRQdb5D8fRrMSGG5fSQt9KXuCJ2mwLXjKBpkIxuGA6S34
FIA2qGfU3dRJM9KRnxxC443O5clP/kiRCKLRjUOg8RfSCEfG6Nel8qRcPSoF/GWw
j/cW2lV6MW1+e+RcP/6e6LmzJa1DcKrTluKsJymn0A2suHpdoyXngk4HMnCJsdvS
JVP9dfUAm+1lZQ1BVubdltx8/IcDAAXv56CQTvvpl2BDhq502vt5a3v3H5cDiAtk
k2CivaQoDs416X33IRgcBIusOnGy0WwUpH+IvX3jnieaKnTXrqEqqcmu0V6gyd6/
ODn9gxe35ic/3thmtRh4lWwNY/KN04qPSUMzwfhXm6FAk6uMRQQkqznsYWfl1M0W
6fOtyTnmuYz9bxMibMVgb3kSI55XDcfT1Nq71GK4E0UQmlL3wx0vzeK5RiT1cXsO
FjeZZSWvGf2cdPuQHE74I6cFNw5CVQgYgd7gojPaxxBhZ+XtO9Rk00L9Efm3C7mT
eqhrzZvdeShgF1+kGPuoqt1IN2KKFh2aJPicLwk0+nGh7zYuQHJRxUUfCUSi0N24
anS1Jhm68cg/P/B4HC+wDTMDwKQPjA22lTLbYItlM0C/vq3J43+3qDIuAwbad7fo
RuRLCdKtushf+C0ccmI3wLnsVvath0np+zpCyaRRwYD2YZ2VwrlO4EBsfFEWn0zt
gO+HG1zwlqQP8+fUvpsoO+u4pViJjrZYCpKTZwpmWp5KsWXdGLmdcZnt6aqDohcf
5zfJ2ccX3mA/SSPjejVUTQ1PTfZHZhOhiETvn8+aQNTVLMh2OLkt8GupFminOGAy
PRj4iejZTYb5iu9i0C5VVQnfuF+RbqhE/LM4+1ArBSC/sta5UqamWBTzbWlqbl15
zg1fmanT4cwAFT+V6q/xJtn0HPJMY7LHNRvRxr0vuT5nynfcCp4Ju6+CfdmblEjb
OAs6mr8N79zvPUSKqbmkiAIqTYJL96DgbWVz1G8cVK8vC/wNRj8dybRCR7emAPHk
CUrSZFXa5dupNXOAMF+WyDQ5t00aQ32+lVhR5YsxFoT8lDZZOdr9FRii+1q4N4U8
VY/Ph+R+xrocAKe2yGElIucm/d9usYsUQ/7CT2ha9cz6akyf324hg0HRwjLfIUgq
0edCNC31YcrBn/TLz72Drn+8hQEf9+LWSRYsNp+d1VBisIpxj5IHT4CfokXJulwQ
/+84tllAUOGEqGIVA/i2cbPtGazNEPendAXZqrsXLoJcG8W1nV/HSFFRnzeoTD68
11DFxMxJzf0aqe2hJlg6FPVrjCDIlGH4Xx1lTgbJoEeb1aiDi5iMEo8/DmiJT2uv
UVEMKJNll2IKWxkmTOKZJGY/OApmEPT1rtZeFk8STsn5V4mjpmf61akTIeDGVcYr
QOmcfHdLrTxGoJ+3EMckfueH6jj3XPvABB3QlCgc4KqAeXpk+fRWaj3rt14tEojo
FAsc4uBzqy7e/zSpSOwHVSjNI8CmziqfsMTz20A5kYINGvWryBBKLqm5E5xRmfkc
veznXcTpDJTleZwzmWR2e8lIqsww8oq+NTq2FlXfZ4AW6hh1kbEg2fZmNURszKGL
HK7iCHRA7UjlHQH2r4zg2hYivfduVZ5px5cgCH8BqdKaralws9xbvvyI5BaW0INT
nc8ceiMiE1jElG+SZ6Ry2BoJehUDD+TP+ub0P3ujTK4Dv003L6Ue+ABdBUTXTaek
YFC/d757Tk569N3acBZe4cZifI4pkwK+58CGJuRoDNjilzq96++JEYAcUUZvg0Iy
iueeA04FfFBBuKQ5gJ3KyBgUs/5avlfdQNsX59rkeMkcDGchrh6TbPSCaFFj9kuD
2d9rz1omr6GRAtxVpHugMN919CQNgHkJpXHNhxdkU+C+MNtTtzf5bYmptK4QWW19
l+zoE1e+/SHM/4o16N4xvI3BfnTZ2B3pI+WgBYH8kx1wxfl39yNP7G5O+eSaaCXR
Viyn+/FaY3mNCs9wInuvLfM6S0Vu9yAC204bUdUx0NdXJ/z/zVY2l1T1sJHaCSpM
qLiWPIuJRMOjHRS85emZdEGGqrB++K6BzR6Ez9A4hF+g9GzofqzDrmcS+5xWI108
rqJQlDtY6Pj/osAZGUleGFlfiUXuqqTOa4w8gQdifuYRqMgsdbMlayqgxo5va0XZ
rI9uE0eTc6DnlLESDtbywp/dsqX6ePet95oUzk1PtQyuEz6S/f0T1DKyZr78lPwY
ah4DTmXuDkPl8/gv2tXzzzLSoyffAJl2yJcDOQLO70k1Sns7sOQ5/SNa1h/D/xDh
SUojo0N9nUC39010xsDD2xhIcKeLzz/vhNBBlShURvk60tm7JL8yjPjz6642GCix
uC5Kgd7Cz13k3BoiV4uq/YVYYDuQqmum2Zr+hPwfyYAshVGihw9wfV0MzHgPp8G/
ur6EbrgeUOniCJnkWQqRZr3aNhgqjBoFQ3TR+6jaNyK4dMQY3Fw5az8xBksXlgRe
MXlh7Cbif/R439+LpXUxAuZMWl4rF2JPZTvgGPfD8BkC1ZSX+X2fPNwsblm52wtu
jLN5RfSCCOg0IkopOgVtnHAkr6Hi4yNwZ9FJBR/G7blrQEb+hlONNs2DQVRsFo0O
Frr6qzx6W4GDHAQaymUz+/VMdfNKA4rlE72zJx/2swbulCBfBE3qLdRTVW3Ow897
Aw5pRbmCT1vqz8skycQp7Hv8QaoMQLB3/HF2J46i3Bw+NB5zDcQL0lkwCvDjqSsm
ErKfRP6jeh83W6ds2FdxPIlDcBGKyVUgOZ8ToaBp0VaS93zFHLijvUNKsK5oO+/B
sopy3ZjNMhDo2OeoUfd9yhnKGht/rNXomJ98d9ahmNM7giChjcpW1AFZm7GnEbRw
rOcvgLNJgmVSbkjCEASmsTE1Hhd/MzzRLdKup8nnrUrggAI++IxVfdmlEGBWUd1W
lDDOTaOHqWBSS7XM7mrko6Y1tw9WT5OsR3IICW2kqGrDB7qh5hK33O2p1ee/Qr+T
qsNg86h1ilMGhqyMopQ2nsgiwK2JT/znJH1N3S62nIsjKxyStrTaocLkQvZme2ZF
6/1rrrUanKJQzBS2uvJVX4EeQL+nUJC1ynHFWf1RenNFsj3FoNiMiloFWTkbqHDC
XAvF+vNlBpfmKQAojhaVkNP+0wcS6s/BFN4x0FbxqF3PhBbB8kG66r1Jm7d4kfj0
LuNXQZ/W/JQvBrXcb25H0DpDZNp++tLeUDppmfwnSGQgYtarO0ikUZ++GycnMHqw
s2I7tK+tiiJDJr2QAHk1uMUjsgECdf3SYKQlG/mM9PzH0MY4QcWHQ4i7zO/vV199
bytKmzeCgJBzqOsSerXimAO8hZb2R1oqy4djUTJNZ8S9W3pQup/XFV9DtQfh12HF
ivw0vijzl2k6h7d8+tnbyAZJHNHBfoIHFddyg5PAq8N5AkrHYauz3elOKgtb23cx
2xjYi+hqpNd53Vj/uIjWJSxfIkV/900Vmj+kZBn3w3vQIHFaru+5O98RTjvEY8Da
B1PjbAHKtkzaZsTj82vrxxMVEOGqzcMgwkfH/Z+uUQg1Z1EA+MR/dsy/5iaaClhB
A0fZrw1WENFAiOlkk+kr0V6wx/Mtj5qc8HmNH+dJq9AW31yo+hcNDOon+nk6bO2v
tfIzmu30MUw5wfWgCwPO+6/HGwWJOdXEbQ6FcobZH3/zEkrgsf0vnwKrjCq9bpt9
XmDaXzFVh5EAuxPejd03P5z41z6KuTZg9GCdoyL+KA1BU6jXoF839mr+OQ4nc2cO
mHWTb7AXBZoquWyt9YWmHlTo9AVcPyEPYWrHtiYHoVJbxFYlh7OPmzpc+6AEiVUB
dLBYD3czzuO1jcx2hI1V2CxP7p+73i9Gl1eGk7h4/7svDopa8gZ21SZdFNENAWZs
w9If7Ldyjxu1fhDvngdwxjgP053QYNMWEx2ST/sQojQsgbSPi3b+rmQizaTYXsWG
s5DF4qvCLsShXUJ8ETz8kCpDzd+yQKttwbao3UXZ8DTqImDvENeBPvqJ1aoN9Ehx
XRH2oB5meWXSVd0NXxitgRbYvc0iCIpA/Dq8pCNmrR/1+f3mBPhuonN0+nvlHUqc
yC9yHJuwebaG5LwINmhRoyZKv8Gvy/slj4EBTcxyeeHx56zAXsZqLlwA9II396vT
6Gd4BJKh/FrPgtizr3H1GAwqXwDKcSi6PTViMNiXfYx/bx5sksAY/oc03PUWaBHi
mNWweozFtWTN8O9L1GsbIFvynWHZtRO59YkgSmU7RipfqBqu0IIaq9VLwrtoIIWe
NXF+FtoIErpcnSzTVrJWHjenpOMzeesILqAUohnuBUUhuSFzWK5R3aHtMpAX9ORC
Undwlymx9ZJ/IRUWmwxLXnqD81VLoQakGn35uj8AFSK19EGSfVletQut8OGjWalE
7tEU/P58/EOXrcsNKJQY5u6dPdSjPmfJwC9EfDurzDaJ3a1orwPhCzChG8arYb2w
Rjb2f6sGZSMBfU8DJ4sr3w7NhNjw2uF6JENIpgkBmiOX0Gt0ooGUk+7PRm7C0aH3
S3THVkkf+pwEY9JJHQUqYA0gowoGkysvIYNj5oLJwR0L3iIrZpyVEGn/XNEnMfWq
LzkCgd51z2d1C9O2LlD84mRMwa2Vpy6AVcTNhdMBjmOGIWz+oZyl33jBYuKZmaf2
zD34MwwqnJH8xJDFNf/MhoihoqopGuE9SWkAxW/OSQgw2PweG4CRLYGc1AnXfmOY
db7ZHcunkggafFPu6ViAkixYCfZ+tYSrFcIy5frCZjoSkNxMHbTeF6QezVlWZ7xT
jMAPMZ6HPSTyT/kXF0ABPvO4T+mlqdSfmunIqFYoHu6F+YWfJ7Kdz8YS+T/FyvBP
3b6l2KH8Bmm28BGY8CQkpKAtGBtoOif3r0BJYCPqlRy9YTtrgTHIhXIRJo/WS2D7
0pVVXH7be/wRj9Rg2cV0E6gStDeu3xpg50PLHgbPkhINPo47MrmzrjKmReoJRdqK
w8kdwq4ckMzLgQ+rYy2E9KFcksB8bdrBVFYFgB1+lZK44tsYiLbKSP4GA51v0tiP
HkTK3m7b/Uu2lk7QX9flY7jx0KHjew5bDmt8GDUxZAtyp3RGqxOTGt3hdaP8Waqk
FoqIs2Lzzm4++isp/DL/Smi0e9lsf1MwspKf+NRAjqvS78Or2KhIcUTP1m5DjGkr
O9klfPsHY3dXKklrVgU7Ze8dzLL1cB+kgWZN1ZBRxB84CuIWY4xHsym6SLKmiClS
A7Rt1dUsvNLB102U4NrwMrKhsyNLncYR2UVgPyD5lxCHyomRieL9g+8ZvdfL/Rqt
mdAO52KQpf23mpz/qya6/8kIMUFvmAiek/1YcTGoFP9vrz0IZngRKIrzbKT1+Le7
sxGfhecdssz9c/YNaYU6Sr7iWx5MVC28BC0aFxZ83kaAhdV7GnLBuC+vfibB0105
aDUPQ7TjxrlaoY+NSidiGxQ3BkMEfZVHAlTlT5qvMxD0qOw/mTzl8NgWP/Rz+0++
xPyTWCXrcemoIOENBnP/O1QmLClFzMxmVMIyxwmqq6ATbhApsFDesQtfdSPpdS/U
5ZWeVw/btKmb61dD23G55m4bnOpMHb76Dj7+1ryOxhdTWePauci9UWd9LVMO8ouX
abNH4on2/31PAC2HmEDbJ255dpzW6f/2PIAdDa/5AcE0Zu4NsmmRi47HSbxQBOwp
7gEr11fRE06XY00dD4mpZvsygyU2G2HnkgVSOsw00Evn7aErtxoAOGUoETmQYTNa
fYizVxaflB4VOt4X+NI+UesAsYJKGjTGbMv0aq9tGmliSnByPqnANX9CcsQsP50/
4Yto+3nzlSSzDKe3v5mDeKURkcnN4hzIu+O5U++b+XfhJmERzhT9Qh5qH40pPrrz
5mLFHMKdwu1aGAYHD/0JTEHv6fq5nesJihPS5428xHpWdBuE/mJYrc9IQOH5xFy2
nE4F24WK152SIDF0u7MXCKwJVm0uU8ylOig3V8+Fnf/mwHFdhYHr/hGpQPM6n4s6
DfnzVXlSG9sojgCMvmfLWhnHE247WRWloWRg4cijYD431KUEq+c1OCSTwBsgkBvu
P7+GMql7wrVF1EShntYeu1L+MVqZ0YaewkT/Enhl9t1QEAN2rdOT1aOyNcD4MVe8
dp/tR3Ul5ib+HFsdAtIqy8SzDUX6l/uqrGuXIJhtpxhZ3s9CDXQ2lzBT83qyav6s
0YW48aew0HiuqyT7xPtklQGOfzQx/YTQZlnkfqXo0fgQ4r+hije/jdNblk3doKTw
m4wNde6K8ihDkb4MJtCO34DHzIhKti+xtMhdZ1dABzvJBhEbzKcR6T3e5A7DYgn+
6ze/6+XVWWRVl8Z+0RA2Vzm6ghKdc8xtEhXpEPCu+R7FIPDVIhOSXHeljysnyy90
grkIoUs4+Sr041iFpVya2zAgN3gY/MjI63tZZxep3++tJnzaXCkplc2Ku5vQwQ18
NJMwwZU3GUI0UYbY/giYq3k5p+Jc1e5K2cfKBtoba1CjBNoASV2h5plWAJg+sUF2
a07PuGe5I2VSjxAiSur+yMvIl6LZfvkon01vVcMMHBXgygm3cL1k5lguFtH7rtcy
fxfABGrUc3wIrCJVepYM3LQ5nLa1KhcBoOzRsmv9PrnRHD23aWiY+D4dPasxjc12
bByojlF2TqtH0qYgntI/iduBfShy6EZ02qlBytfoN7W5r5VdsE5qlpK9BpfrUi/F
TAAHn1llAx2mYa68e4HqEOH/aqLVh1udu9JMiPpdhtvSWOoQAgWCP1pcdRXMQJuV
CREY9lfJMCoNDeygA/k3OUiM+WyekCyauXxldVMM5RQCvOf9GmhoxdV6B8bZAT/r
AI1kEGIsNqBuOoYrHp2ByRjvYnWyP9Sw8DvB1Meh3lJuYHGJ39QRSIP8IRGHicqi
v2GF5K/9+Vb0Qp1kRDmwMNxDAADAR+LCDue2UJ4V56P+ExI1F3tQ/YlALldMcRbh
fKMzleqSPBghIlvIj8b1UcWsIqCGpF+H9YuIb5f5rAnJAIuOWURo0qFBdwRg9wjv
qcfaL/whNYaa8tTswcffpnRtuQ+AG8WxZTwXy7pMiuv9lrSHsqrCLE4+QJh585eo
sQm8ssbxdQYDwTW/bm3hdrGnXV+KEUGlTrNHFOx033MUAWgjDCUiRYw0kU80Xzkd
gNnZj23+msELJnbwNzyikbpuFm+/L5/Zo77fNFXIQiUl4Lqg4vJb0z4GGgguQfeI
QHnKNVLJU9ZWYTudEXUaygtBPHpNv+3lEJZ5ga/FCR2sukUsH8eiugM8tAjd1i6q
gLogOhUZdO3Td6sEngmkM9nA3BAedLyIMMtMPDnQAj9kt/PbcD/5SUpSPGi9mje8
LfUM2MqYvPF1qMyBDb5Jfm1E1lY6SY4ZZ/Ml868496756f+n2Cs+6ZrKazLLvyoL
3jSDdY3gwh1zSufEJVznnSxmZ10LTeBJXono2ywAzYA5zBFwlLnBM2mEbjqbdM5o
rD2G7edbVBZROHpuoNs2ZY6dmO47wLS5VIHogr5mkT8P0cz5DV3vg5h0kXXKI3P2
Nd8I68vgZrNbxtwMIpVCO5NjZuC2hOicy3nk8/1txRzlrRwe3lnmPkYdsoQLGFPO
xd+V7h/qmyp1QGnuVgPmWQDHyVS0WlUz13X3ohL7CZMs0Y8hntUJ0eIkokPyw8su
SQd3G8GJhzRPtpkBWsCjfkCSHgiPy9bnRWATcyH3Gh2rvYzmYl1Ir+ACWE/yhB76
/i/izYtBJas63FXRPIXZUgrPD7OME9+fsD7kU6ioMeuvrHbrIPcSJiq3qOMYBCEF
oEkc0iCCnrT6m/zKKP6lPd6CHw+ZjLNdCHoHkogDxmsTFrvdZU7XDR5IVkfg7wks
D7P8sIgJE1JQvYhHNk5uYhmOOCJj22FbyKMXh4GJ/sGb8aEJj+1gzepXfG4+rWZY
zvIOocXSGb1VZoGlDzhbi07QClCDw1C2alakmSlBkZJcTU/MKwkZ5OtczUOAFPyy
wbSzyFKoMvWTUPBB85MD9oDJ0eG9QjkDHU9gtJ0wkBXjDb8D8wr/5Js+ll06/bLZ
xrHqgg3PCY8QYg1NiZxs4zhj3K8XRqAodxqdRfLavczRobE6leUYkPl/cY3TFrz9
psevbjGvyojlFtTBDjtPP+Yn4l04lNJynh+bz5M5GqsIdmYiSbXIBu5/h9wN5Vxq
J0o9PNFmKlUWfDU4eoQc81YjXoneVIoJQ7wMT7iXsrUOX5XutyJ6H6tKkaD/vzvB
8Xxsh3OG9GSGhnYy2k4bPvuE20Ovp02zwwrBwBMQtaT9KefMyi6kmM4p/TAj5P2M
bTwp1CumPxRARw0GyxcgulPB4C3BCFbZL2yjHCYnUUiEwZ1vXbhaoNHNpSl1GZww
oRbke9nwN1f1o3EF24bH2pLCFp1Xeqgl1gXPcRUfoqmbyfpcdVKANHG6Sds9AR78
jiF+UaWOBvSzXsVbY+v6PLi5bMgfb5qSoaqy1SheC8BkpY4eKY/FQtfcbt3B79XM
EXr1J5wvMUUgjdBjUNF60584cWL660WvCvvg44IJkWYvLnPNJpQdZkDfqU/ca3AZ
NMREBfRjhaToLAUihj0+W5RuSIo/Xk7nJ0e+pj65eHCfiWcel4fdj6lZOsHYiaiG
EZ+3PybjWd34AOhPFX/zNd/HSDXDuzgMpq+NMvMY6mBifuiJx61R3IpTWrTeRiVk
WVdaUmD2jXJDRwS03hkDZUbhndMxpQaRWkPf5PpUw7Y4GrPmRxVpQkM0J8qdZE11
2nETj5cmr/U5PI3mIKF02TL7sZel+oiwRgE0g/fdou3Rc8V7cSdNNyZhCkZfDmNV
RxaZ9Y0UMx4GsunPKSQDvtAS1V7BIHF/RTh2glETc7+pEu/bOt6SMweaMCIy4PHE
eEK2gxOdDLA0kYLrg/33sVIEUuEBl4HeWEKHm2whv5M2HwlHs6CFCj+95ObZzrQR
Sl/hZehLbkL6cEJXJWOWel59AGN4wc3EMPtOMr8at8naRFVk+wZR96XHFc6TC6S2
25GKC3yfZ1IPAv3luO8L6vGe+AOjqajOLCA0hp1kc2SmDtpMPEkRBGjtGReDWMca
x9tf4gEYvIZ5ECmqHiPCjIn3BvRtwHLTYjRw/HTtYVkl2ahGcpAKxKzAYBWGUJdL
xwnc37pyr8uEpI+r0NR+iILAhAfThFv22bDU2hzGYfKEEIkKouCuyHo8svB+GFU6
cVNH869TbYjTrsRQuciAIGHV3bcp7gZXOhhX2ndMYHUlkd9NJtlMZ3Zc+ArGOKTw
A1779Bt04biYFdTxuJfgj5vCaOVkH2FxloyBAOShDLMaiu/PQjjkK5UP6LtUlB3j
3/1AUeekLS91G0XY7ZfQMEFBtvDHZa/Vd3alFotfK7/iJ1+Yq0yxC8HFEivJss/k
goHvcNz55H+RoX8m6fVjwVJ39LTJvRE8Yk2cWt9Nz8VMt4kf4Ouk0ELsEGVmDwvP
jNEqKKEbbL2fw1JkhbVGzQ22AxVBA5xPP/BIDxD6jaoRqXIZk5xPW8jLUKwrQfX9
3+Jq9R+INMCkHapGXsGVzamUcK1SV7EJ7Q8wYIt/fbQSLo6tYVPSB5rfRgKYfU9b
q/6HcxS2XtzNqu9Rq6Br/Yjz2I1uFnxbokkdKnyhIvCCp/b9z6NwwPp/5Z7SJGJl
8ISw0z2A1aH8IhpH2kvpHDr33aCqNIxvC/gOJqyj7uoCkS3CR9docJIZrRuISK1O
013kUh5T8S53fws1l44+mliHKrl/fTDW8REYCBEeQ3IdmlFKd2ZOZOcbTLfCiegf
tOPvnp6Kiu0Wj9zIKBbNZD+tYPbUqGyvXs42bqlTxuBZifatR8tGkcwhGbSubbGf
SZ+t3Glq0VZDhZsrV4FOTdHBHiqo0atyreBYrbvVW120JMPaoyF+DRrBi8MkvMkd
oCBFKfE3LPeFP/ARNoIs0z2+LV4uF5MHHAldiDMQDfYQ5BRnpXHkfunu36xvccSS
4hTPIoQpRwKz9iZ3LI6c4E0wqJeRdYc7oV3Uvpo1Q2NfuD5A7TfdQjP62ueriNTc
ci4BxAL84VaQKJONi4tnW/d32JP9AlTucVZjV/TTyCKlb/EGvi5bShZL1lzKVTz4
kf4EpDxbjKwh9Jl4ZAY9A7WMnY9zqr+Z0ITcIdeIIT4U5Y94WlPlvErtjKXj4zGZ
+TF7oeL+2txejDu1MD5GJUnZYW1BDOWj7N+mzurleQ8rRCvzqCAtNrxPcmEa8eOr
GVaZ2sdUyVdarZk2WYBdLnFLUuxRuHTnuEew7s2qmHlcdnitwm7wKYPEHx+rNbBV
2TN4FWZSyQlW2a9jhAqyDKJU3Mlr5Cp4fy9Zxu5w5W0y+ckuifjbKrxiLrEw9zKL
c4wzMgK9CP4JbjY+OmTj6ah3unRFzl1LI5XM9Kp2QBgZbogmQwVe8UHHvZ/r+dUa
QyN0FZRdFdPreyVK0LaMEmAmznep4BqkEEE7Zagv5bEBu4nFJdXri1WEBCB3mgd3
U86lBa3+kn+se5GPpnKYDnvifBUojcYOQ+n/IIHj7H+q9XT814kvZdM+UJiqU5Le
MUR1ltO8g25LsWWt4GctECbOrrAmZku6J8U17vm7b2bRHqi/cKrool0nBOEKJ+Rd
KNgG2F/+k4Z2zL0458GTVPpOHpf8Sc0H9rmcQ2rP8/YEb7Mu4zWMqudBNSwhAC6S
hYwSHMGTFk5YNdQNE5hYAR1fFMFIzTDzjW+V9UmRpYW/+XFQMlQLF0H4NVHC+1q6
EnM+spX1RUUOj8wIlNL5jcVdNLqO3k+YnVdWgjhFXoNno6gpHfDuu0Lhtkzuapgk
w3S64PHlU3fd2Y/aSo90wDkC2UUYDTVv913V4Xl3L0PHUMMxFsb0nl8wtmweA8jq
fisLzC8wuMohQpfyQ9HJLXAuYTBF+vI/mJfxLbt/vcU2IEa72WKF5Ayzzh/LtJQt
FKy1wSyBg08jMgyeVYcVL+lD5WCv/TJLbiJTtM/ieqZ+Jva3FUuMLoLcYD0qBpmB
M3hxEMp/qJco6MBCUl51A8PMysNVw/FKYdXAZxND5ZUVlTWmVSr/0TdOwdmfDVPn
NJEMtA0HmehSWRNDW2gAj+NOGtCwihlWUFZK9V6FQBOZjM2s5v9a10o/cGvvQzQn
dVJu7hV698aO40NqZJ0kxdhyJfjBCTtqnY0izOiZS/ykiXbzVgreqF7nCuOBX1Hw
ioBpLTq6xDjS7k7Dl9bXTvi8pMdXV04i0E1PFABuMrw23gb69PoaekVgID5JZsIm
LeP3ErNZ3WhqfLK4h2XKcghY5Ie33UkKvFFoT38NFLjIG5MRHQGQOj5aOvcjmI8e
EaIIY/xEe+I7Aup4VneZZvIQYcjSaKUYxzehr9EgYh+ZO12BsL96cofpj0t1S8n/
/hAfUMorEeoX7e8FaekNuy/jg0GTpEVlSzft1E5p6rBfjWPG5yym/C2IjI99tSI+
Pr9UQlVdE459co4MCZZXxiP3y2u8/VIgh3zxUQ+opqcoKXUbCMpmKlhPcVlx96zd
9DhY6b+PeQ6ipF7+K7GaJ711sp+29au5CTokeodBZJv847hMm+dnrEH4WTslTXKw
Un/1garKdAmCUHtQrNR2wSrCTSZ7zq9YLAwgoor9woBBsXjXP/a4x6SXTeg0OkCA
n8MgTHbeQTEN3JDpXTATqE02Vou+sjrPkbjtWBhhtLC7VtOy9t+8HNipE5nC1H1k
I556R88ay+0dYa8uUJhez4/rG6B8ufUJXQQquVanRY3nwtGtS52h36JQTaUtEHnB
eXf+CJ0RXLr6uLXnN54JseaT+KwJxbEcvpHsDbdkY87/DKW0LlkhHn2pqdyt8Ocm
hhs6uuoRO18ITtSFxHCJF5B4S712bmU+7qaap3KD9ENGeqJgfBmQ+sRNMOGSJdT9
a+eSGdxVuiLbUUyqJBuIlNQlTyn/+oNnyBdQ82/9qoVv1Y2hKjCxaappxY6naZgL
2cbWsn5IUPmTf6D2L7aBqUtiZ2+uthTqobIUcu31JBeyhhM+2sedovBW0hNUuRLL
FTNMJ+hQn+MmG+uFO89I3dtAZS8VNkTzT1fNKfka4Y/rbzbvdqE5esnsok5e1ZKD
bHMvtrsaZ7FnwKxgo00Fk91z36rFCxJllGnLp8dvDE0XT0KVymDNuKT2UU5Ris9U
JJdTI2ycgNuTv/wUrpvPD+35TnVVJ8edzt7eXjnWBcjAMvpc8lQWrmX8LBZEfo5W
lnofcGG1W/9ax/1EkAPurvijbaKM2Ub64C9tWNT8wnsa/baPQGFXeV+e+nCeyOid
YKeRevV9BOQJNTuP7AHWaGNCjHSvoJhmcw1KNNS7J0ASJU4SKbXAiLBgjwvE6dC0
TGuOEFUha0cAJrjcf5YU9lzHWp72pAD0JEI81d+RzGCuBxeUktIQZG90gNsdKDi5
WkQjRF3MTMHYdBtU4KLWUPTVa3U1cn3Ykh3UATR/+3mKdjNV21PcVHkd5nyEspAM
xGJBP5a78JPUpaeW6qld9GC0E7ddo9ONIgUM3Or4ik9UvAaCNKis/6wFGvEC45fJ
QfbfI21sesimuv92rOpkaKonJIBAhhp21RbKJthSigkf5iWZup6rpYCblTdV8kBH
uy8IMOWYfJvPmEDp48BZNGdnmszH86cx9NcXP/KXcAxnN86ln018GVjgcVEPu+8e
SZNp6YXTAxbjQq+QxWJ3tCBeIPkiRFkFgsI/XfAQbc41ZwJeQajwaWCKXAx6MncJ
q3VF0ElodVpNCeQqAw8md8OtLh0vovGhyAb17Mp9T9v/5ONGB503S0DeyZnoxlb0
fFg/8EX2uilVvRjrXQblgxk5ww0YiVi2svOGhAsG1EH7QnIfaNPY+fXLK0K8bVG3
MjjMtYYkHkuzj3yemmFmiAigHg2UetANgPlokqOsFZLzo17ptJYYkGGwezzmBsth
RpPqU/+vTMn/55cZMGOcRSykGPsFbJtViTJCdjWOL0Xwn5LcuCEOzahsZx1bhOY/
IO7Tmgiq9eGiEeH1qe/97jy8m+0JTTksFoedvKNyM4VTUf1/wJHloUhIX4vUgS5E
y+Gqv43H8om2eXjVZkZ4WzAwCSs6eUj4echpvXrrmRv+snRR4LdTiqa/TRCJm7UV
GFDRF2IS23ZBaGV7lDwqINMAoOSdIb+P3ppDz2hQYQ03Z9pOtKyrnt0olhDSXBVI
7KS0turzp+pDZTduqyECcogV5TxWq2JaXyj20NQngZ4viXFOpLdXSg5lrkODXbU+
ToHXauhqHERtDMW8oi7iVFXncKbPxN50aHvopDi2TIifhpzqWrmdOIGaNNEMM3sH
s9it6SSI72immER+VoXYEyLEFPNUAirXkXydiD+Z9BQXjm6pfXcNT0VKOM+GIqZ4
Kbn1iV88Ez3vK+wwvKx5YbcR6uFkr13RlydVcbT/yUix390tXz9bQFn1PENm4lNH
Zz5RZf95BZRyxUwV9DkrF8jeRywuVUuyX8Z4Fdre6iH/yB34W/qGRScgfry/VCAy
xt3OD4g265EhvgwBHeCw0CUsDZ4uxOTEJxlO979es8WEVhcX3XegUTr4Ed+HkV15
qMQHZn97Iy4nlKo5rE7wZLTBuvqr9pjDO3lPe7nCIqyJVxRNe/JkF7Gwa3UhAgK0
R+b3DwotL+qHs1NQC+1L+/Kli86k+Q0hVDdYiOVy0UtqpG2muZSfhSqaqEzyOUx1
OcmGuJR7F39BFBOymAC17vw/YyqMgWgG1fWCkRKN/NhKptH+B2pM5eXxrC46Y24I
C5zhs6oiQx1ImqJhQrXr5QBZ93phE1JPSB2LKRPRhqi3V6UlRr6C2ZpQ2kNUYyBz
7TF61n5hPUCew5gXIW83y+T7MeJH5BRlpfNc3Bizg23Tui+NNnWrJXMRYQskWUkU
B8Rpi39sFfCXPrRvJU/A/01zhq/sXM5usuu95quhqznzOghCCQ2Kk9WHQrKilHeZ
uvTmqBaCOVdA4l1Xwg/RdE5QYvWpFr6oomtRuruToIxB05iT+rI3DtCXUQvEc6XQ
hpOYN1mCqh/MnmPXNfrwHPo4Rc9QfakxnOCbXl7ueaYsOfv1TgxX8j/BRdeaQVan
7Sbln35+pFB27ZSzxAonCDYWjygxiXF3vxp+TNk4HaIVf0c75PZE7fHSASVJqimt
HkyeO/Yue3WLaUnLLXcO0RcDZMu0e+4hNvHAlpGIh7vLm7gR11IfyzaaY44C+e+D
gTY0nbopUkYlOeqpNWjjoslHy3vqCDUEAEY/5q1GK5J7OnJDJVhWs+JqmWQmullJ
D/0vqI24WtLntPN73hw2VJdSB1JTrq/zdAhKbZw0S5bItDEturFpmkxJoW0jWPG3
OxsV0ViTlRtxVAvGBtJTezcp9XOH/wKEpRg7TJUk6WX97RXaWSdtdBRQtG30in5i
zt7z6lKu9q1wmhyl77KYjsArvdO1mBwadNRUMCVB9io+NG2IfYjGcp8jDOnqBnXl
RJRG/rcNUTB40wmj834lzLS9+rdxEwwQGdEt6DH4uY6KNKJpQifs5Uykq+Wu+tAz
rLBkEsK5VyWPssghHVslTODy6d9QkcYuXzZMO0Dn7d50AAQbBoe4jpdYoFeM1viU
o7dLNhVn6uBjn30UOASrg8s5ilVJIVHe94W+HZ3nj/pJ0fh7WJZ6VDEEtomdLOh2
5+mw32DVJyeFXWiWdotsLNYuy411s5rZ6xSmeTVZXkePnZ9H/CEe7xmweFa1Qm22
kbMHFgUYqW5Y4g9AObSLnB/2rsUAxRhAJBmz2/W4quZ03OAKsCFgboFEv6f2+96N
DyGVJVlSBsZDIFWpC0oNUY2OLsSasrIIkeeMWJPO5UaroilXw8lt3UgwIkgGjxNh
h4B5MezZfrwF1epJHCMDPy5gs/QQtz7lhH5n9jx2VaE86hnHzmKFxTuSnCjGHwOL
7pLkT5S2vdnWq7YDlcLQAuxFHXAe4FGTjCEbUcug2QhRUtFrPNKWpX2YGFtP2nnr
Soh8ksW8mcAvBG6GE3u46ao20n41B1zfu2kcccpU9SPaNMrDOxOK+j+3J5Fu2pvw
6ee4dbX1pqOnDLRRlMS84BA07FaTe3C6SfFO4T0wQTAj3NjJOSmrQ5CF+DPsRPkj
cmOiLlUfpS/A6zFaIbPq593coZV9zbrguErldCA30FeeclmqEgvcNJm8OAqRjToo
6nDFYfQlueiY25+ODkCs5HCCmdYfoAMWm93Rjty+JDafW83ONZtIeW3JQ2aO1M4j
9NO6/7lPxv8mnjKcr3zVlTBjaucljp0jWCy+oCPGR2BYEXmTVEI84QD/e+x7S8Bb
3QbaQGPHnC1SeGm3rUMjvoXWJQDFuBq7HsYYBfAX3wWrdRNsk/9kN5hycLWzF25G
F2oLL8WG2ZzbqM92QW5nxw15uFdVfa/h4yqOMTXu7mr2KJt6cqEl4mEbMMwmSiAZ
1+rebyaIBzo9OG3SanCB0nhWC6mZxVfd1vFZ6BYFxHlZWhiGKO9K4u5l81FirVTh
0TrWUt8tiaUcufq44YQZ2FKXQhuY3l5+WJUJdoANWoxgX4fl30afzRGXJoI783N9
irQCuhwG5uv1Z5Dzln8wBcNdBpoeWx80rstvYNyPmE83jcclXITRIzt4nISqjRDh
0K35dcGFoorwjL6aNZORNeVzQBEf6CSnKRy5Fb8wvdmjAgod+z3gmhueoU5anhcV
0KozSse6SFKweWzn0Uc/FX85OLI+rBAJqUd0AUbkJE0jVsG7J8J/O0ESGuHJCWi9
P/w/G2+YohVMSAUCd9LGMP1nA46XquED9wjiCD3kkQG34LW0xKKN+4QSgGgXmg24
q2pJM9d9hud1CgCFVA7Q0RWhXNDYnEJsvjTfaeIVgB5QM/w9yMdmUYryQfj03RZv
8BCF+GgH/0vMqrK7O4nlaK42pqoJTlSayLZsc4ZfYkoO9Lxmr8wQmXd3eRJg4qAI
P+4RcbQtmSWeWBeU/3wfwehJUHblDgPJkrh1VRaIOaDH0RclV/kKcSCa+jx9W9+x
C/UkE5cSSt4FwoH0jQKoDr2OIcN8GmEqOzlm/ZlPSGpdwBZPG4oDVpfGJsGgz67Q
dnQ9l5UiL/GzXbv3UVRsl73XTALlz/TRtr4QgzyzyYw/301wM0eTwtx2ucr5XZ6j
nHn8+dy2dZ8c2T/4T5qk3zGVunCarIp3TWJlUPdyW6fHTc3Y5ZO1yst30FxS359q
mvrTw0S5bo6qg2SAX+a4L2rjL9fisMU0CaDIBOB2vdtO9BJDoGpiMw0okGY35by2
RKy2fO1JcBlLssrhIuomtEDU7USUJ2C1fXK7u0zKLF1jC2qqX64WNL4klu93JMzY
Lm4HBeFNCLDsKPloAMrvaOPHksKDP3pMq8/LLa0MuT7Kz3FYcmbQA6gSZKIj4ueR
00hZctRNHMNUL8eE7etHuiKQVnSvs+XdU8/1ecqYxSeLe6dbEDaZmlLEZBpWlucT
eBEIcgOz7OPahVTM3vfDwnIf4CNEk7Ua3E+Ocjkz8d6R0MwVgqS06Ynd15Ue3vW/
4hiUNRk2fyCsclhulZehBnebmEoKWotSVHK8rq6ZDshaYnC2hhSvzlPpCbaFiTsE
+Q1xtGSxeg+M3jsaDverHKDLL0BWTznERCjMkIe5hwmeoSRaI9fyrLXEmnfr1rQk
33Vl6AUvFTaXW2K3jO8vq4NiOyrs5RijCCmYer8VkAgdbbOinwK+QrtnMyOWKG0o
CQ/dUbL+J6edXpF+qVmMBwEDHe/9L86AyyXFfgrXYV7YGcZ5UdhjRL0KdccZrHWy
wuoZsmawDsDIHq/OHG2K0N/PUDHgfTNLntAihmC62Cb2nyQ9VTUVrgArRSFuRIFW
8EYCH5spfwED9bdfLBKlzY9dGdA3DBhzDns7Sf2rvvz451QoWw+ZoX5TOIHxwPIi
UWYf2swoJMjQcVeK05Y2q3aHhXXYpWE0Yraat4rmCZEFgHb6ofNeMAY55tKsroc1
AX7FsNs0DB75ILou7vcxwGpufkPwkdBlGQmXMjjZjs0PYKBwdz4A6Z94r6dzxrS6
4k34/ovvowe4Zo5wDWgXmhcCSVQBS0c+qUSGQIwuA6IB//WSYiKBlP02LhU8Rjv4
s3yvs1IfyswJOHnDKjC+lg5HrMP1dYIc2UC0E03pGHvT09WSQi9dIW6SIF2D7uYu
3lZr0KCcvSKMwcHZ5AXtN3EW3wt9T23G6tGSUG4cpY8vYBjpp+Ta6Og+nkcHK5by
jxNLcNlGZPFaTJn7+AILYlnu2ZNMTmzwcW7YGUDYssxEozLwUvKCT12a+O5N5/e8
phjDI8YLZYfpnESmC9WJ3o03jBfrcUJ16fFHXT1uuEjs674yRmmqjlxe94c66KpQ
6pn0tLiDW4LTVH7hKVbbR8LQNwh8n5Lgn0/sK6IvqpvkJy590IWEfXgY2C4v0FzT
HFW46KwBp0EyfRvroEPq7itB5gaqO6bG0/znQ+BV3Btq0frO4OXpq4khKrL/adxW
m/4G4fC7yTs60Ol6mj+xDUaRKmWwFJt7wIh09Fa4lkd2eTKIQk5W9plttFGkSKHU
hcdUbHJKjs0/SITaLj/HYGjfCMVX/WfbzNidXp2Ht7G1pprxxYsLGw5sXd6z+vYq
XpnvtqGNPOS5wkNDfgCIiLlygr6NbcEc+2+JiMeXsEBMaU4Rr5r1zRHQMz9NaII7
REuOsBgiHN1c6THXMruRGTuBwcqRba/wgpL/P7aj/e6a4tTEOelgk7vIVSdUIGHZ
euIi80Finf7/Rx8LkUKl6r/PktrzO+getS/6oN/ptx0p5kgNzuzwEmQGuaFovsI+
fFoUi8tNqUO4PWK2mShmPEabv/XvWLx+VwaWrwYO/sMZ22b7w7NIFpYmszMrWMV+
ne2IPvx53SpDu15qAcUFA+B9gqjSFB7mztpAC9ua52llCGckYplP+hP1fnwRQ7ak
67j6XnNy6HCnzowuPh6X29MBIaqf5Kwpp3p/kmiENkIbQ3rU3liRNJZEWxoEC9UK
P9D9slmQHRScAZ+2ZWjw1Id+NKxaTyEX/DIf8gsLOJRcdjNVvdwAMJYbgjuVNk1R
/ALTF5kWbGd1Zq/8wahRsqi6gHQ+MDlnSx7KtuX+WU7rd/mPe2ZzHQIeMo7MOeS/
+74JBHRQJ+dl0/F4g5Jtgj4UvgZKAWmndO1HekDqGv7wT/keWwQLNPR0TtdMfKYE
dfkbiYhwWjZobS11PBqJcJzdyhqF4aLNY6vPJlH2/E6Yp3AKOoYnntd+Do29FcMS
rbNH0D7VelfcT8bp0sDrLkm+SLwjIx4vospwG40sGJtbX6TUXqOokXmTQJ1ndqHH
tvwdfhAeGCpA4or2l6zGizNMtW9DQi8COVdBOaZFdj+oDGqPzhF0r09wn93vEW9L
FgVnvAI+pDD0TfretVpH/xOMA0TwV+1Q14hmu3rbHgIvPhGFl33i3pG6xa8opVy6
moDRmnYhmFtF1JkzhWFl2kmFUEaDIPeBRjUh1SemDa+wOSZAFbVVN/WqdQgjcADD
AECPxigUYcKIQ3Z5qmGFQa6mABeqHuuec0Sy05uwZfR59yBRHpKivCfdzBexEoJU
3AntA41WeJHED9KshWKhEbWno40LjHJULiKcicGVFyjCqYxZYCI6RPXvdgUPnFDv
VoMBewZkNJU9jo6Hs21Xh3/feQDh8CQRMD7K89Jg+/AYjwMA9hKbBXsTqA3e4DAy
d/ZTlUk2W2h7VU29borSw+GhruAi/D8kxqew8+FacIhamkfpf+ExLumKBg138b/P
k1llwg8/HBfjkLhIE6lGxKr7RwlIp6bEwxoWSCQgT/PHfqnJdkcinaHKuBOy8LEx
TCSuns7Ea3a3dmOsgu9YcB0BsQnYEVuaIU+yV0yEx7mUfDhMBrRmmHy2+FVCCzli
mUrSYfAznuLraBnd3XG7ZVNOnHtgykL0kdtIlQRNyX8KjIltHErXA/hQse10EcEw
vcbDo/BmzW/3Fw47zvc3p+PrdsJtEuldHrUE38yNXKbEl+MxZb3p+sIui9gbRYrT
hWKuCfVA0D1Rfu3R0SVtF7FaqY8zCX4rDu1zFGXxKAkmAmlmXR4nUErKp8QFu/eP
Inpn7y3haqiUssntJfhRPRt7dKk6BGM8zfmVeak24V1WAQGaPnyRRxb6QSmS4C1b
O0Fr4IS/VyKTZPWkRcamJ6QdvVQzKBeF/7jCH/alBqQDERTMJjkerKOBgFJvr6Fn
HQg4X/TVFIT9RCeEfKZSiL5q+UlhDaO8kf+htuexq9Q1yf7P0OATqkBUYCRXiLBE
oGsKTYhc0xoc8BK4ZTwdk1EYKoUbNIvfLqT6vA1Ed17gtXv1vmAak8AbJ3W+N8Ha
nYNAqujRvLruMSeCWJHM7keuBNgFTrBmP32bgUfu7bERrgFKfFLbjfiJZzsZSrfx
1zfhWl8mNIZfF8Bnka9kYorczf8bxPcJNw/1zyFkSoXAgGko1QJeKT0SmpILDYnA
v6NVawpgH0xx1qbUVXfjKOlKOLty2s3c5zsk1VufH2NWZRdQY+boiiKzWVxtWASk
pfgHyziSv6h9c1jqdoh3PduLdnl36bR+2jhTluE9FGM/XALgtswmf+IL3ON/xIil
wnCBfDPfP+vTdW+pv/FTB9nhECVn6c6AVLS0t2d2QUhHrQeoNH0bFLqyicXVO9jb
Hv6xbduavZCUmlqryH4DvTGlnVp6gLkmRdzSDofJGr2/uKDMARDenSISakPFe8VI
ECkxRSgthmVnQy2xf6vL804O4mDx5CjMq0/aq+V8o2zbEtQnaK3ktWcoynvlKZj6
rgan/IlgVYZ+qv1m6+Pc5GmmnHQc9HSVsworAO7fMh6OFJljTK36b3k6eiROM1oU
mVA0HWfnBM88QuhymSm7x3YaK9PsLVOiXGWeTtZX26VfrFqHLA1EgI0fWHog+7rc
42vvxEhsWDPIbq/6PKhshCQdC/VgSlIN/95XOSq9rinInYuv0/fLD7kXx3qbgA3c
ApNqFy6GlwzqXVBlWCmHLQIseAedx9o2nAzU0xhGrUWC7LV/RhbUNebT0cjpiK6i
WAp8ebJGHpTUKJGJxsxiKCWNvFBTrO2iCWBgfRJYsj4RcZkRzoRMmLc1GKbb7O8C
2vn/ompclJ9XDxN6FugYqOED48aKwIa3DMnuq9/tNK1OK9sIoIRNgjXtZqZxttPd
WFljQDQPsu/8VGvqb1L0KEMFN2CfscRtwYzcsK8EU5++Q6i30JdTGo0553qyXMWQ
T2R922BSp8FVa8dL0GkQWmlH1NlXWbYjzUFKNQJOOdN1IaX+By5jVAdWx+/s7ESC
0cYUG4rTiynTxxn1Oc4jlKXE0uV5IncC3chsE1wsM1uDxFJJp3Zl5BjtJIHwP9yB
V/oummsGDuxtqAi9Rybv6ZZi0sOqYjxG/HkmxjODF1GRb9fGGrf5LRiRpxuL7hjo
8z2OI2FswseZOB1Kz8zzZuxT3ad7IoGpj8ODfYiKFJcxPjmM45nk6fi6kickh5hI
TK8QeIvMwcdxuhwBqWqVGSR72wVfJk37C1LAVQXCDh3g7xavo6LvoSi1Yid9AehQ
Vs/4jcHHQteUcRAJvsYZ6dYPFecPF0cmsATnVgNwHw1thgaH0xcZcqwPXvpxWP+4
KrV+3BowcIE7ExkQ9CaVB1TIsJKuykt6I/aU5gEbDzETl8AHiDbYuOdR8hSCIkO3
ULljkc2c2ONSAeo9lfI70jVy1KXT+suRgWSdf9LQcbtTg49y7X4ij8+tTxxSIrtg
FXFLje290Z3P+Ksxg0c2cu3XXVgT8rlev58GOmsYb00uX43+swBXHhJcQcTp+Cae
zvfSXKQ3/C0inLPZ1ua1auDjLHJm87/pBbV/lCX34cou4spclgrDl0ZC9DH113LE
JvSEq6gkrrlnFSdeD/Tr2w16ArN3E6ROQE46UkVrPxhHZA+xPNNFDI7JW7mTHHW9
Q5exUfaQV7j+gEi3qbuUmZYq4xaSkmpZZnyF+tuDGESCQ+joUsj2D+hRz9HKcrZs
PcEQdpNzvvZpYHWhrm9b5M4U4Mxk1E928t3X5f1/ttpFqkBkpoETR5rtsLI+F/9P
E7y6fcRmfMaxKUG7aJbzt5NSaPP1pnB+Xj0dkaBvGRbktDKhP6m4EehjySS7G/1Y
OX1mndasUdc9DYtORXbLh2TNNy9NXrI/9HMTf6NtLn4+zQp4tZgKGhoc1XqmgNJz
JYnmj+x09o+1hZ1V1Qtw3N5p1/XLfJujCua75dI2zOgFtkSyfg8Qx3CpeCtdEkbd
5CaAObBQ52yeCsisLZRrxtH63VxQgXt4tCohl+VR7nyJlrcKSaFfibWdXEyNOEj2
7jyXmUBKS5U5JVaU+KI0nMDqwieBsqzwdCXzb/hvSne4c6wx2KCUGfSZK8CwLCY1
E+FDbY4bjRCxXfLncsZgb0XKDRGQr8FFV8UtdfxhTwrURMHjUOnUnj5H23x/2M/x
euutoYP9QvVOdUZ7DAeLaCGqoOXqLTP+T/tF4k93Jsf1GHtWAThtTIt047+Lijxs
vEL/CNHuYcrHcXxesJgHn2+K9VjrwFm2ZyciT4jEddUtx/qa8VQhJcsgjRF7MYst
ZNaKmpmbkZHjk9ledIjeALvq3bsO48XDIiYDzeKkvxLtoe5C+MT3K0Y337fClu0m
az8u2eJ8XmDhI9J7ashkvdA8Y44L9h6aTO3on97w9PHrP9Md8i0M1mnl5+vHk0Nd
FnAwjTJPYcf2nnUez+kun0vSHxw/VWz1qsZSQHzgm9SWO8jfKk+UjsLXdJ2DsyOF
GtJZOc7/YrCOWQ0tgOsYyuy5mswGwRTT14pobxRzs7/B5ZnMd42MjIjwsob4jZ15
T3bntWNkmxNOlTylm3lt3PE00dbUnpGmZqP/AyBSTwqO3aPbw0UmTT066mtKCX1b
Px3n/WLOpgU+3bZvfmHeOwHwsVa+u8+pTeuGcm57slLWx1b9Yu1zQ8tocGGbu3Fk
Vfj4aPio0nKx+lV1Nf5sBvyd26jv9MTQALbhkfVKd8rArI/2zJTL5f7537KuNgei
sqShmWOQsIN76oTwMQkxPElq2HPTC2ugOnyfQqJSA2ZyVlUt4rzKC+CiS8u7ms9+
5gMCGyWzG0YyCXI1mskb17Vu1uw9V+yW3WAebfuFd0+jH1sxTZx6ytXFlgnq7Ay5
Dj0bEXTF4O4aTNb8VmQguhNMgoDqwQ11880mxUOzXKxDF7S0pyHNJsNWcGdrvcNN
QZKpd4vHYDjOvZ/wOdpMqoc2vVoZgKK0gyNzb+KR44ozkvDOPC3dj4BTM6+HfU0L
WBhLcQXuzwo72lUOqbQAKE9CN+jqJqTSSoIYZWV+t3dL/VvaniPie/I1y45QTdSq
BJPO5RrABvksMXXCnA+O82tdToy8HeJZZmS+07uYtDdml4f4ofw3KAbiKM5g2mgc
xhSGLU20evVnvlcdHyjGsF+Ryr5OKVqMgSi83RqBB1YXvoVzGZZ4XqbLRWkJPU6s
vm6adl0VkGRmfsQwVenPvjnzU0TX2sXnVUjg8C/pTkjRlmAZdHZJxQnOQ1iP++ET
+D7qgAA9rO5Y9qLtMUwAobPJ06q31RZ9UXmNvpCc95oEQajMLXVDvyJmrNWWFy1b
v4fSOYiP3b6GjjA8ufDN4dw7sEebMPKjjs3NtYbEI64ONs/02fR8aGKgmQgSrmI5
Z61bHJlaa/XjKpEv0RgkutWWMR8C5fvdkRfAiQP78OUDx8uyaSJ3IpoH9BoFPO6b
bosGqtDg6Z9DVVYmX0sTiH6vc6xHt9/AqzjOErP6l3vhlnER/VYKdJ59mhNX1OZP
rOO0YidbOHMT7xtb6XRPUjpGaWQCOgxv6xty3XW8VXBCsXxaw5fObU2P2D9brLaj
dDuXrGk7QGPzEVP2Hp4vYFxoJU1FbMQ413nOM+9xwbXuz46RpaQuBssmnXUbCNN1
lsxqrwhUq/fIobLsFxXmU+YFSCypH8sYuhTSDnAL47uKSHisuD/aq1MgjEVvAPqw
yyL8GivNbiBMCv6/Yfx252XrfQtNlCejQqcssZZtfSrRM8QdY28uEY3aRhhT3R5e
DrB8uye2qHsZvZoDNIE7yhOfVuXT8Yzlzs3D9vWTyLEtPdPShMIhHWn45Yr8YajF
sqJxJwE842dVWAIZWqgCh5lO6zHP5RhNHtNuG2T07io+NnuhOA0ONOqpZFXoeOQ6
5nSY3nIJ1oVrf3wqLWMxYRU56+Ss3wwgz2Zg5B6pYdwpjDUcCL4e6RjUIF87wfDJ
8dQ1voxdEnxf9yYezuJQFquVhJwNerWo4kDhSBUygk8dlOYwp5bnjMIt7PcpekSc
6JgxlJkKrvqNXtsbJlNK+0dmt2ObklRrm6w++IOphuQMog7lSLLdTagp1K7QUqFf
HUxPKiJf7sKSM+G1G2BJXpdh+00W1v1xVbmWNjZqaIxzFDorFuvCRXzjaj+VZGX8
J0zkUxC5OrUOm13LBepnRA/4xGW9Jr/BtEw6YXcyg7m5yM7ZOQGoL6hLDNYczqPP
p34AWRImyMOUz5g33+E0CbS/78v4w1+2XtS/HH6YIaRy3NJqH7zCE5+T6L+phRd8
Bg1W7mG67IMhauHABV+LCnyFydn81Q1zdJagY0udjv9au+5iwCm8AIHsDWvhGG0/
xAKv0Zb33DZOOjRJuGK0FYuAheIAZEiYzJ9OEXHwzITmhr+LbCkf02fO4Yj2DZUg
V60mYaIZ7AUJlWySrvtLxtySzn5hU/mMw+b+bMq17kAzEJzg1/G1aT2hXtm+33XY
yrPJWaNOW/dsP9brlgmiIj5LwOj0gGZJU3iOwNGnY6NIzdtC1jqiifZHWitfWYTt
J9hvtJXYF+9VFvxWUWFeFbjDEbUzdGpWm7UGq3TBbrxmxJwhBJLv+N+ZgapXZ0KH
oJx7f8VdT32jJFbpqoeWgFB8Dm5NcZ15e6muptD3dMCt/iAMEMT43nVjj0JI3Bmo
o7+FBhqkbGWwbAMQ7mJFymuTizxBunwiCYwNMZ42Z9oBoQ/jT4Nxig4jM2DAaKnU
sY6AsAM/2+ftnBvOhE+UwAHabThvOAIGPBsAzVurETPChhjnt9Lgk17sdILEUUX4
24U5+0dQQXpLfVPO3WCdHbC3gpN+mHADGeYwJyDWSBUU+De3aT+FZSyXtwi72PBK
rV6rps8TEMw82TRQwICuvx6Y6YT/Y+GYegisHhRTURgjHl7V5U5OqH2l0QMd3i3X
IKGJJRXzeKQLvoFiozuYAyz1DJGvxFdW1d/bGoHqCVBOpsnimzdwcmZBOtAQryMW
pI8S8FRolMigHDkzpBgna5lq/pmo1LrixdrLekZmcLmGKFAqXiuaqnxuU1FjKJnc
Wy5TG18pl9K810o55aOrVuDJZ9HE1fz9YxKmZ6ItUBNNnEcvarZKXakauF339Tyr
F7GpnRs2KlpE9taTT66wxtRSaKWrf1BX/WkmYAg/+PrTqAY6c/CyIbwvjJs7DrRb
lxiCg88harB7UpUncL5toqn8sp4OZejQinWnaeIbppQvpNrfYcUlqSOQgSRxPD+z
DJrQGkKfKAjAGp6R9tsGLXP3wA3V5Cs2ROaladdN9X+tlDoug3VzoPuJoMfz6+Wu
rvK8e15GUk4pafHBqYJZlQb5/CLEqu80Bs8gDUVnT8BehjSlnbG0afR5+wyy1AON
8KFlZMXsNRXZaUJNc/i8iRg9baAgOUBlfhcXakB1WdkvtYOzBUEBKu+0DruCO0vw
K1dPrTqaynikdp0+XgN0Chr5FCoJi+d9L+yjC5kbcwGtjvPCLWDvt3HQL9dLZ7fE
pWwCB7Y+cidCNHQsZDELN88K06Ki4pMsB1JL2w+lbBILOvSJxKMuFpX35vo7bQVQ
TR6Ek63CBHnEp3QHTiB5Vgk5ELMc7uxm4IuhyglBrOvaV7xqIzijmtSllJ5Oi2Qf
vdbKvjKuDmD0EN1HL2A7c0ODNdGWITdjPPBnK1xG3oQYIik4TPPdEedfDMYPIJ9L
I5Mvz2Qp1M6qUt3EFFnSrbPE3tKlkr/9Cgp8eHTTPmP5L0gaNYBJviJXYZKr4bUf
zoR9x2SsfQLrw0B8cbbQ/N1A0+mPoL612Q2BL3TgFUPzn2LVtZH/ml10dNIIFVnq
mY3fmAAvUeadHxej0g2OvoviY+WmxWhWGP4yrL8ns4kBHtEHarOPGvFWbreoqXWs
dJLH5V105kIdg5ppn9WYfymlPThh8ry4K0Ih6u79Kz+Kp3g8V00nWe5goify0u/w
GE5zGGy5dtLDGT60pMc/Uhw6rlRBY2V4oZ8h5FZPsoMVC/HQvJAWSZiPN5KNVuWo
fG3ujYW8FAZLOyIh0gXmQ1imQhF2d6DoOHbELky5Z1qxGy4uyjfry0gVTvra9rOW
3iaVU/Sx4QOb5HJLfkYVpMgt6YnWcyPBWr6++InxVpfCVr3VsM/c9IOUACXmW8xZ
DTuGvtjR7+mlecjBI6uiVMJCHKkf5mDtmrL5Hmxj6bqEmb+PH7bfRYPsAHujunB6
2wuUKCzrqFSDQAhwVPi9nj2CwDTJ/6cuDNO2QsUQ68umHI0JRL2DS6ypUMOIcGqD
8Sm3psj2vw7W2iyiipdzIVN8n/8h0amLoDrksSvUDeoJRnmPiM2DBw/ZoXFUCerF
U1OaaVvg1ooVqvibnPvelbfi1dhJ3p4y4LXB3C7sIKbmz/67N5wKh+SEiCiRO4Tb
LfnyolN6B/sYcPkLqq5tTolJEavhoKoaTMh/cBW4k3bTft9xcTfgAxDRTCmcNEcx
6FL3Fdclcn3cGUyeGob0gVQLN1btqqq07A51Bw21iy4jwyi7AbO4CcGy14dWXYJU
O6Fjj8+EG1QkAp6FvorWLjFafm1ST7amKOaSzgq+O2zgYzfMOO2azKZZk3g+XLQL
2LURlrCWKAlB/C2mg7WI34A2jAzECB/zurOkIfW3cYgKSgog8CnpwGXanq4P/OED
zZfyVEwrsazIoxHdDp5a/pizYy85ZAOtm55wa+rMGvCFeeb/WqsiKD7sQM8/bps3
X/39OdoftjmskeXZ5NF6jW+jI2WpQymA+QaQFCscTZlCtKxAacuz4VYTliVDpA/v
qoxg7VLMP3zzBOAF1Z6QqTdos8jXEj+E5Fq//4ackX/c4/mihST65AjHguiA698G
awTl3ARNAg3cHfb52mrvppLqut/LHAVFtZWYcKxk8TBYu9WVXM+ceoUbbJVzRrtu
7CSisFryvgZhAh8zgnISTuEW1NH09tkIDKGKO3OXh9hoNa3wNJm+2xnPl7wimvUT
fbuhBJiryEhsAMv9cSxaCkvsbsTD6WlVgbKSujlABqVzvb2Rq+Zf2Dp6Nq0YtNSH
h8984dHDQHz98yWVxB4JrcpLJaENJQvwboy+yHZf00lWFYwHok4F2zEeL3fsdeOA
ciBuu5RixQL11QEvOdJS9sf7vwXM3RnFWfMuP9YbMnUMnGjjnOhHGNYRWqm/Yx+/
YyJFFLud6/S6I3KEPFsz3eMfGIGGOT9XK3EIbbZdkm0R/lz6nSPbQVBb9MXGUZde
10wEXuEZCThvogItzCYoGy6iiTJYAe2NbpdWXyuJ1KRzI9RsrSBtK8XxiGiVBlYN
Vso07crg10hUaW3qBuSUSlXZtOHte8QDYqdCWKXj1amABtBS5GdERdjvvIfT/YBY
o+whAFxRkf02MOr2NjkEY3YvwkiOazL8+eM8Up4o0Pzhlhz0Vn6qEGvgZCx4/bJf
dPCWtW4CxaZCwlmk2nQErKceXNH2mq0xz2KhSAod9MY8KOunVUIAWSHwT4ayDu4R
ioV/CM2iFtoDPzEbZeeEzeC4/QaBHFF/c/XjIkcULEYPJHzCVT6CB+/SBsoEEo+T
NlUv3EsUX1nr0E2tbL3eIaJXNOLZQvFlLMUnVAZdZddI4jG8Xq2fWhPBes01aNWX
UaamYQfjdsMKzoqNWD/BkLw9l+0Y18nl51Be1PH+zmD8ZEKBrv3n0BPrMbYtaRRC
bfRx6DkXS7W6mV+WXWS53V2IkbNmNN4Y7dRDU8no+GJaO+N6ZYrpKinML/Ncd9W3
lc2PQadrf680BB1fWJaAbFNDhonZWfNo3cGrXNdE1AOczNE5fvQox7e6C+xpVHJ0
ws4+i8ZrPNlHyZ7XoQVlZv/woGB11Modow4L/szZXV1tGdAfjylOV0gsi4UQNXKl
2iVAqpnwZgDm5jHCpqwgsFSFreGIl2MhWgUnaQ+By7Apq5H6Xi+s70VpWHyD/zZq
tO7HSSIs8jEPntDW51nm9hyJ0nAsRsWKWCUT7Qt6sAKlA6Adttv8hw9GiWfI0JC0
mKa5Kd85/+SUAqHa/2vAvPtzUvR+Ajh/98TR9MZLtPmcUdWpNteu+o++PPq52L22
aM1D93ucgqX75l+ljOPUB+CuVbKTNJLwaTOUmUD9aRrc2juXWNp6oCpGIlVJM7gz
7yMyQwkGqziEyRX4lQ5KZd/BsHZh8uQEQelax+qCxh5N9HXP0qPicduTd2y8jQGr
3omiSn7uQZ2BoDJDqLy11vI4aDwq4Y0Bc8zWj8lT+Sa/CgDCqsOcc/uL5mptNnrD
EJ2lW3zN/zSoisA6ASNaJEKFTmV9L/zs2FE61Q5kGTl1A529meP7Qc7yzPLPplgR
Mq64leIZUHsbMbIPt6tqblVQqg/HRBzY3Eqch/qE0KsKOTCQZ4BraQr9LCP96lSv
9WRkjWaQG/ieVdyijE8OB9pwxmyV/6jE36xLF1LOAkhK4z136Y73b5MGE5JKWrb9
2yOvR8bSWI/+LGVjhFRrQ6ENewwJ9XuYwBsWY6mXRuvSFf9aycDaSIsH320/4P9+
ggkDx58R735qkO0i4JzCd7ryJdBmgqF58ocs94FrYIucO11SvIRuKjpUUnva+dhJ
b3qg5TFJuogQjtuF7AGOH51RRN0N9zwvFR/y51VRTTT3VnWeQCs6FcQllLpNeis9
5p44en/tK1VV9XChtd16w28uswHHI3core3BOgF7Ufsr27N69uSWKb0DgvTUeAcC
YKYvMFupKjxaMVvrvOspoDatAOFWacnUWzneOplrRVvk6w5+6uK6bJU6D/5eGqwi
axWwcyLBJFQAkitqzGMSIQ6kxubRMbDeCH2M8wKGkSuJXs0WLNJPjtiFpiXul1B9
p5cWlNztldv5vl8uDtLphcvXuiSnQg4H/Fkz5ehnqVn9k8fEfLEPv/3J5yXisgK2
NkrhWng9+PkdEKfq/wy8isEaBqNWSWUm92JsS/yV/GPO7wnIhQJEzAtA3fjmpoVq
yMxVMnv42epWNI76hDRtcxtz70t53oUccu6t0dZtdDmxjSVrdTE2a22AoOgfIjqw
TQWzGW4P2tymso58k6ZcDHxF9DYEqZRIKTKpJ/U5wIDW0l4TELvLe1Z4/LvtGDH2
VlFZGpge4eB7CWrlne5fJjQrtprpzqmA0+OxnCPORaOVBME6EXwgeXCFexTgrqAa
uPwQ1cLDJMIugsnTaMJAA0fDf5MMAt9gjSY0jF+7P5CTMv/wBsekq9AMP8f09g3Q
wzn7IRV1MkOoWii/2zE5Pk/I/7rZet2AudnpYFFoEEaxTWxHxzMebXGiaFiY6U7T
VWIRNPASs9JPJIcsvd9teglb7vj/aNfCK7ZMkPW1rfHRH1BsAGyhGtSvRNLOCNgi
4AgnElV93OYn5iddEXnXf5kEjjCDiSJlukUNie4TqxDYrkPVzbmEJOQD4v5f0cCP
Gp28TEeThAEkxVaydOgWCCu/e+ubT5Rl0aPdAwWvcPWRvFJNeprFxNL80mNhc+kb
y1eNb/sw94Xz6jx0yvduGSMsUGfEFYBuRx8WcCHQgjZlC+jHUMNd8Q/gpj+bisdX
ABXZ5CUT8s1onEPUM1oS+fCxfRdSrFSCS4u053OZrpdAgeSpR9c+cEjvGarvEjJx
0H+rq/0QxyZ4DllGADg2Ftx1KO5ywLAxrwrQ2BQeeNODClM5C6ftm0rDIBGFFnHE
6d+HXcZeyDUuK2wyEMimNy9f9YMRHLOPzND1ulJoQaconxRz78GTeWzuEaHNNdUS
qy4Va3ANHBvIjRBBon2CPfvf3ZiS/O/MDg7Oj4seIQ0v166mwYqyAYYI62Y0raOT
2vcja85qhWsEGxXCbpFOdvB2Ojo48531HbBqUrN04RYPetVF8Up9NM3G2pOnJnh2
UFgI33QajA6LFFlaLoFr/TODv5uMl9+vdA/AkFInKlII4HL8o5x29SI9Cn21zKwy
jdNNFqSyb2//27kh7I+b1BBQuUoAGZzBejDrdWeETVDtRdc5scIdlhfJOSLWKmr3
XQ4e5esXJQgDw6/inEMdzVC53ciFUL9ka3oTUdd9t03R351HGRE7zXFbB+3OuNvD
skDPCVNNpRbRJ1YidpPwVcuZiWZGwNuHeXiFn8kqKIOaNmL4shfGHeMLWxcfdlwn
rTDoOVkn0U/fVXpbMV5GcYL6OElCFGDBxQnGhIxJtuL6egZu6FeaxvZ2vlSfyDxr
ToayQTu9V2PW8k+0GASKx/dyFpUp+enV0U2RvnlR0lIMUsyAxBJRTzwJQNeh5fB9
+cTgTUPGMHnr91y7rlT/mlz4ljwXOB3zdvNi8AsdgenRkIBw+M1/ZSLyd+N/MZoc
30WZ2UCS6C7nK/fO9qb4m1wQjeJQKmSxGD1GGFwyayu43tqNP+A1jLRJTaYWsHHJ
reN69AuOmfB3vBJ5LNLL2+Lt+l7ldfolx2xwh/29nTAOG5wNj80os+uTsmwrcW2W
OVQbaUQnkqHVxTatz8urvBMykK4oecmCQKU6er8GtqhzcImbG6IC+K3Du2cczoR/
qmIm6+O9CMzzZ3GhD4ohOAuz4kG+ZS3ZnVsfZ82VFse7KvXbohhhg4W628AP3s0g
f2RSIs8QvozYfwMKsVmxWVpNXRuoxc6GR00kdKAEeanZxLpsg2k9wmnmBsEfZR4L
5+b+ZPOhxuUe4xOatOddunjvRMD0hNkWXX9MnQ4oJoRJoBk2Flblp1jzj1xLA/fz
SwPNvge/LAFluN+Y4NzLYoP497PgfBOC4nT2eK08ctGAYMnrMOfVB/Uyw6bjdNPj
cJkDF+Qr9E8BwV+20XR3IOa01XRrZ5thBdTtB5HGtwsS71+1rX72q4WRmDvlvZcZ
eDtTp/yrwwh7yGLa96LV0lQIYG6PblOUc+6CkuWwUIZjUA5TH4lVNdCZlmNKgAZu
Nr8VQ6eUUwUQ2vLSGTJn0QXJX1Vsxr5AunU/69PcZuH21HLpZHlOTak2rILg/0zb
PIa/oD+O6r615jrKZMdfuZU9YvB4V8JDZiNS4A6/MrV/VygLou4TwRiICL9s1bhS
H7UvfDmxKXCnRGG76/324uOdUPyDKbb4Oflynd9ns6MvF84Rero4RTVOpZAyY3Kd
3ONke5vbQOLXuUifFlWjAjxY0v6L+gB/3Sa/EitTOzgW9GwJcO+ei5kIE3PiThQ7
d/KNdAehe9nyWhqY1dPqvewKr3WgsO6aAOVUHu3qxpQZ+lABq06Q1UVMi578+kwI
zZ3jDwzHomjAvEODwIp9gSITOEq7CfZC9TUGdIb7CuQajZegGeVyQcna2HAeW3iM
KlO532gj5PG1NagDy/pIZzjJ+YQaQY1rmzIUFBfU+5+RbKCNmL9hptzL7irt2mDt
LSpOOe9Amm+5E1n3EIl5yfw563zwueATyjFQMLCC+IY058e8PZWNEOneXfamM+bn
z6yHzMLYx5DHn50KHkcFi4lmzPmuyln6p92h+2cRYNyD+RrnPoiMg4WAxVQ1uhfe
6yp89Eioqe5INiUByvDGWLNTCoC+pOXVNlwYnIfA7ituo1MPaeE8mu4j9q+lJ1gR
Vrftih5i+CZZOpWO0v6irv07mx33nlK1BfGPrkvsDfVR3Rce5TQijKe5lqTZ7V09
CjB0CSxktV6LAFkglNOYVAEOJHfRAaoOxikpZzmv2OPUuTDg4cz5DW+rjaynNBwW
IKd28ZXcIrV4Wg2uXCwmoiZphuSUIq1qMtLEgGFjO8GubyS6j9CI15oCreL+N9uU
8uAIm1bvVMGKGOetjfqDgOQyqhMvHBpFIFNiJ3V4sIicv9JNEubN8qC1B76uWzg1
w0bCBnWRPzPiI6eU/7Hi9vmPvYhOM4wa52pXBpFcNux5o1jep8ro6eIuSnCpOrpX
PMFjJOlEmGoFGwhViLUnq3CwwytvYVD0LFFpnUHxK8OXkdk/qkLY027P4T0ky7J3
ktSJ8I5+mef8ADq9Q8uphQx+c7YadFH/qcwpqLeAvzunO7v6yu7j4vk5KN279qYY
W0fQhda23I7kouIywd5Y2kD8VrdguZZ/lCagHJyWzL7/UNBhfsX1b/DAcJbOI4lk
T5VuyBZYQ1yf7O1YEVAN1JF56hoY57xuay+6vDZLFkVCyt3+1ceOmO4uN+oc5+4f
9NDIx0JKtsdZRD/x1mF8H2tugJorQ3BZTH0KcMoOwkDEtpRAoUDQhVdRegSJlLOv
hWheNqaKTv/dLKcD0mRxF/on9dGOjl9bqjxY9UbLXsCinkA3olEhDOGhpWNRrEdP
0sTCmr/edcJnj5KDZIJQkFcqKSnjmg62TFVyTU+4y10VMTqgJ45KYWuP6JnA1iGz
PpFB7Dy8IIV01fYDNLv/74xisGR9c0C+EloDsNOCKSGpRogN2IirR5wkYHjzkRuX
JVYk7eBCXE1xGUVPjhjdrOzA6BC/3gPzhaYqL9htx04bgYxDIZWspRj0bgLunirk
qT1VU31Qq1ZkvzESJ0zjE0RvnYR6hBk9SHSzMmUJxduO8wUW0m/WE0gwF/e15mFi
gX2F8XPU4qw1WZdYptmwgZ9RzWQ73MQxpRdRx9rpMw7F9b5d+LQDJVfDglqwISf+
qRLsDFLYjxs4smmCbCA3/cgSuCxXju0gh3lwZAFhpZhK4JI+ESWGDXtpQwFKllko
TxAoPLlgAGiXey0bvRVvYZj2PKPxTq+NUOjWq1PNRhv8MmL1JreOnNh1erqqGEky
uZtmWyOaeTU7qrwUT8mCjcspKIQoOyDz60DTtIMY5jmV1SvHxXseOeTuQ6OZDltG
a/OIjojmhSWD2m0PptAwZXK3xNFqQPxOU6B7uIwP3JcVq50Z2naDY3CL2xZBlOOo
0WJUer+/6uk3V4Nqqu9XhedUdDuQM78tNmYJdpyWVqKKdb0tUgV5El6Ty8bDjwVO
oJ8h8goTPFXLhueysccypz5ypUAqvg9N7sc1XQTx+Anry36Ab/EfWbTnMWzJzxsW
Hh/nCaVWr/AxSrGPg5uGNwncWKGCxmYE+LxCOwSmkUDzUqqy2jpq750+/5IMyFH8
laK86dCnCqah329oFFQtmV1duEG953/91S8fc5Te0eN1PUhBsF1PnFVU6c49vKUi
QvNLLD7mOKZvKJdpf6UBGl50hgpLB7XcQH/wi+kkvFI/c5PHR93z37SahsJ9yowc
CvbvxuoiT1qttDGI9mRAjPJsTmF+rpFQ7J/l6/y9cpjit/Oq0sDsas/GJMcVEAx3
h7OGCpYjQIDv2ddElh0SWvccTyk++Gr8NepDOPmmGt08oHLi7mZwAj3sD2GELqBn
EuxLMI+d18Ug+M8sdYL/nX1AMOryGq8tmXG/8E3uu5+xvnuBdzj+qdUCoM+SiD4V
BzXtRTO7tYy/v2AyOIS4rVOPga1LcXopPkgVGqplRGVHY0XU4G+cwcgJlKM1Dpuo
gtGq90Y13Ic45IMgEsVsvwMhNLSY4ma+//EZDbNcvuwjfZfQwMA8wmfVWn/EWxrY
gPc7Yy3K7LI149tokdPCws5nuXksQSqBnfhsqA++IYeqXSrYAuCSulfhZNXsbpQP
g46Q6iwhHoEUUonO74Oge2gfCCnJZsD9EBI2Wy3OeorMC/MUaByRKI3wqxPCpdG6
P4IG9QE5zmLLztEPFm3afXLkJ1UPYvOB0QRqTWkySKgHT94jCoGlamRa87yLQD6d
l7JptNQmB0PxH3GpcsmgNpGlfbCvQdutDRfPq7ZBTPIn4aZb1/+bthwdA356/m8L
Ndd/qPo6eY/r8bejstr5X/sZQ1xGHAyeuRg0cvau3F7+UvkHP91QNs1vMXao5y06
45wS/13/x5UdzRnM5GoRsodQJfWQnkq9ZLba9/Iow2gyXaP12ATdvsSc+HE7pxVo
ZN4nyr1k0HtO9DBdBijH1Ymtv5USp0FrFtZR0rnVvFXka+1OzAEffwCv/Kyzw+II
TrArai3jRAJM5jRjK5TTXm9xL1fOLvMNqRap04XJ8bkQSdM+xeKVZzs+UWQe0bKh
SvCrRmXSx7QJ04hAl9LUagKMSILVTnoomK7iYGxkS95jfcc3K8oThD9bthg04UYT
65c2PjV8g8LnVRfvLKy2MYLJ/89mTDnFu+X09SHkeRRpLf60dCJBQP1Y5In3oXwX
x9flynbXsAe36Vv1B/uJLG8ljMjTUZ0qNJii3PvNPqO/OJXRucwfKcbHFPcdS9lA
ZRAFomU3YBSpAbUQ6b07afTft2ehXE1NNK6api8hcxmxs5qqngx/UL68clFAHGM3
jE/SQpExcJ1kD61cRUA5J6hhBGkit1PohvI00RKZH333XIo5wdTaQGGmEZ+Y+4XQ
Qp7Vz8lAuFr11gl5U/TqwlT9zIwEpwaYoXr9U/DYotrtLomKz6RYaAlYuBbgZWT/
+/UVY/6elbwr8mNZlNqFeWhLLgu8cIaumbVZYgZmf1vyYnhzMoxGzzgg2Yq0lP14
Rn/+039dcb93ntykDzzOq4kK6LK5mK7sTeS/WziwTJP18Qivc3q278UGJ17AtdyW
VeP9piSv9ISBz4gS0xnZxp7tbCGxo0XwO3h6Mp1tWS4RDP9gqUVNCu1hYP16WyqD
PkedVtKuKXbwPBrBeDIqN3j0eFixJo6fBE9eimJMHgz8sWqBimAj6pMEWexoh2cx
54fM2Fm09mfZD8WQSBlQkFoKIVK8lB/Txkt1WIc2F6mPd0r9RHl8H1G9LRKR5VEq
Mw935p8cmJDT/e57lhbWL9TAhKwK+9ekpOQyoXrdoUyz8EXRL2PTo3RNabjOWkgD
kvL0b03gPqesWEcZyPVmSrASbdm6LflhRuMcchlJ+pHT9L3LRs4MS/5ybnymvsCc
bihq/Itiks1ryXM/xBFiNzvQsxAfqQ7HINDfb45XHyXGhYDbdV/JjzCGSb+RNXBg
swKoXcJd/h404eU9XJnRMQQvR1o5htVIkRdxrjpKEp7VhmzABMS/rzi2LfpUxbg+
QYgxzf2Vj2DbKwmyvTvJWm4yzvUzRb8ihq1JZHNEizF6UwO6dRNS+7IYfhVVSVV9
T3E+tp7X7MU25MmELK+eEqUpmdmV+SaQGX87mcl4Ybm4ryVXu277C+jLCll3hwSb
PhTB4tCnytIEu3xlYx5ReC1CE40kaDUsZ4FCrmP5ZPso2c5cu2XK5CBOWz+CGLDk
SOvbUWbxxqnbwu3XivcjvKxROPzZJhNNpDi03VFbnfSsADqdQNtgnIZYd5Stpe9/
ULJIlHhCjsD+kuZJTGpgHvhqZf7dbLBnKoSwfbBcTvV9PwzNjWspJ4TAVEoIsCNb
IIbGMSoemioXL5D1jynaZasGQ6ZZrshpFwSnVyWKmLhYYUQ2MgJJ4n2+NUAWfAmP
Ge/fJ4j6F4s0J+xIGG5EeWdDVjHf7+9ohm2WJi1le1CIgRgUPIDdGYZlIRu1Qcj6
bSgTUUCVuTyinfVUauGK9u8YtKfhss91qU0MXGerkLrz9OQENQ0Aeq+L3whIBXhV
t1yvd+zCnyprmLAxjA8l/mfa1ZofZYEKRLZRfbXEL5SSRXc4aevDIj6ev0GdOeV+
RDGEM472oo/Mtz0Vw8WEKfD8HGeI8ry93UHHetrQg/h39wy9KhWyvWmQtK861UHu
zJ3dNNfep9L7qAl63zHrOswaV+xLMeN15SvwDodSVlPDXohqr0YFlQgRxUgJITTW
4IgS4dIiqGkPE5eDt6FRdj6Xa3rHYU4C9sPHbQyaK2NnC5AzFjNUrbNMnRMm3vTo
cLxOKAuu+8cRXSLRWW5A+nQwJLXNIBbRwrQ6ZhVbrBmJIJtnOhKCcDJ/IGdJ5P4I
MdcvBIyorp4zoml4IeoEv8TGbhrgTJR2tVE4Vgpb2yIUqHGlMT2Hjq0MihrDa9Rk
YzFIa4sLQLg4RgdtikvkgcEHMr5hpSz4vZyLf5fqiTIwXeqVY2Z1318Rsj5FWEhh
TsRioRy2J9xr/pghhTq+YqQ3Ct2B1FZNzIFNwKRMpGVvrEumInhUMcToZuUGgpD8
rDIrMot0GCWVt/ONzLStH1kAAHmO5/nnQTT72uYt1qoCQf/4k2lS9jvkaVLQ08F8
4UU0ePVVrmMGCSNnLdQUzmD1g3vqTMw33PPlzLetGp3bkHPdyNo16IrRF3znegDI
Z2FuJ0lD2zfQETsLoLNQ62UON65Jk6iCc+XXBAMLknmSduPB49OwdOy+Te1KJTOT
4p9RGBuiTe51Dg4NJ5VdAKa24knBrPtxhoHuYQamcS5JlwaWIW4/xEaFZ14lAWQA
/XU6YjEJ4Kr3x2BbgsBPsbr6oL+QSjfjPgisYBq5SM3LkRAS08ORsCL3p/Uq89dE
FsGV9JPrPfKC8iZrxIOAmL5CbCOkYe8EEe2GUOm7ANCH58H8GjWdxjgUUVE4/s5w
gYaYS9wP8i+AaUwmY7jJ5eIIQASyjNkWvNoVOVY+om+OJSouSCIbIl5SzEWLi74o
xWfohKIItb0ZvA6jv1G7spwMfAISrBvNxTpWTZN1sO98YKdMjJwx+KLZJdfMUyD7
GNhASzNDLI3vV4sqnK0+xcKsRXk4ZyLMcRH+PgdoXtakXOuc4jumvN77+nehCVxt
RK4Nsu8/PfHf7tKykUqmC8vNy0QdRJ5sYWold87wOKUQZki1U+mfaLPIydgvBTWl
jtBjHJQPWpe4PLdls7ufmSwsUUSZihj0o8Ij6B7Rej0vsYGBEtynniJlx8KzxASD
sJv2r0v3jjH+VjinIj8kswWVIcMhsAqsU2W64H1Ks3MaaCfiV3ae5n5qKKSjzZ+Q
UvBqeIpQG+LEv51tiZoGLen4CgX1ACYKOrMGW57UVHZC7IBwqEoKRkr9fwCcp+bD
ML7WrUr4J19LYDSiTT8jBv+AbY6zjPHboNMpp+IwzCecnC1D8DY6AlWBfg+98x/Z
lcm1rUQtJ7MbHcthjYfqibsuPnrm0x24e2IfwfrNh8ttDgn3tW+WjhYSa+9QUEJC
u1ea2dJSKBH26mLcqh0zsPIrwXavoqsYeUJLfbNGEh0yODtLVc9/jOYFQ25syFyq
mWTwaeQWieH6BogriUFSqcM/yijNibpn083p/SC6FJvbUG4IRbjTMyyoDelCrzWB
honzdkkdxoHNGztjwfIBy0IaWdTo/zLo9JO0dfUEtp4LPzIQk4+ChcDkeg9Y0dtX
/hcTP6wgG/AKU3BRds/bbvZUPepiNbE3ipoAbZnJiowYSI9a4YNoHyNQYLp4hK2o
eFOg3hy25dNvwei3oa7Jeq8mnDpHTM5fq0jEdl0DD/AJHuLebsyOA06G/N/50LpI
whqAUtJP8fHO/V3coSLjsfBYicoFeYdtKG/JGkiZvVuZRxbSqo9RaTwi/BCgqHve
38YHby/ldGmIh+Vtag/TGYbb+fBxu0JZB84zaafoiUso8+dLdn/ypS3jUN0ZfhQW
ZFNY6Aunx1Wukc3jxFOaUCJorNDoapmn7raX7CuNB/o2hr2xQk5mQrscUbZkhngX
cxWO8vWY2U08yxG8JW/MmPKPt2PLMZNLGiwY10JzgFPTbcbAgKXJmTBqjJt4wZdR
cq1LHpe7w4X7Jnla0N9YWjZsHJHnJ/QovZqFZGZRCHDqXONVTefZ0TodOPAW9O90
eTAihQjlMyiED0T2giuLhYBEwd3acJ9E5xs4KCJ6qmJssqd48omhgykx9qtY6Q/Y
wtdG0XzidTPn4hjEZP4AbngMHE2NDZlxHJxgv8jbgBiVXYH0epPdTbjmQHqVkliI
44mLwNylD+VVIPwa0CUTbLymvMduULzntAWqccpSUrm2Iq5T9gZiBxx4RjoWdPbV
u3yN52H2EzQGe0J7JVeXolETeP/DVw5PUAxOBh566iOErlqQfOVivrGtVNukyV9N
ZrIUAcmN5mQ4ObFXnMjAJ518VbPwklqW3PEU0/JChsHUKvDoU8yHbS3bjmUX4JPf
uexHLVmT4/4vKAlevr3MAkF5VarxVVfBwP/bv2X8FUJdT4jWqHyi3O+WVShtbopX
q4iooIwWMB/0Hz63BowuAw5yR5DE3gkuJ4jr6jYW4uNCLJ+hD8hy+B/9LHt1v9j3
B/9QPShq9r0QlVRefzO5TfQQf1Jv5mB4m5BVuLIuifmOFgF62pav/FJN6l0dgPmf
in1M59RTIRmGI05zAN+ZXeBJTUkAWl6jd8zpImKfQX4fDzZzuJVrx+45WC+wblIy
r54n+OsEhfh2O+zBg1e9vaUy3TFGzc6MsGtWLDVl86MaSExbS8l1Rqj4sutnP0tM
KhFQ/IBL3K3yz1ffZHjgti+1BXGnXnZONGuJlPwclrP84Qh9iSbqQKCFqveegZyY
aEjGSGcjR9mGD7X1C1koRsT8bBqTHUW4emBcYIwdYSG6Up6rB6k24sBCBp0NLCYC
grgd8EHG3ofpmDF3shc/jwWFZBlurE5nMK2zO7Wf+0VloqJqi7EjNHY36nuIAHVS
v8R2oN+kkpSecsSUYNSdyikXMvlZAr8r88Dy6wud/859eCEICR8AgSpQtKWWymQz
qqk48778K4dwwWqDi0937d4HIb8LEydQ+apXSLC1LM5udj/LeNTyx0D0ZVBAUppS
QiReQ4wBR3ee+QWbm7i0eD/HgaYGLAgoO2QHb5/15iGs+VOt73HiaT21vd4tRBFj
0SbGTiEjbOkqzeFY+VvR/kieDdIf8G1uz/QyayW1KfIsYC2eMQgmHIlJgskrATsE
OvT+uQJ4ERV2Bo0c0tvrucyJyCtHLVga9w+32AYXGJ/62OEN9QqCSmfYLy9gWk0s
Hvinru7ZthAkmTttWKV038dosw44TsxudO0GGKTIGQIgRtuUpgvODVFwuvr0s+sk
gx/SPuiegzTb2P9+LfQ4yAk0hnX+yFE1Lllx/98B3H0v2yKhoJaE65wEvi14oYdc
9Ppcxu9XkqJ/8TyLu2p1p0mrmEcXMQPvZ1k1ZS7e6DNvVDcHNMm+qP0qjTId3Wn6
8gMOMEAq8+dXdybkD8KyiLS81r0s4Qe+SvCgxgfl8Aj0Byw/v1Hig8vC0E/u6oHu
Iyi2wLymlqwo5wDqlA2h1B3yadyIrlqKrN7Y+tTTk0+9ytagz6hEynLUdpVMoOoC
AvzIYnY4Qr7d64keQP1UcOfStMuB3EW94y5ynfBIpCH7QGXflFYbF8d7QsEN9Cph
OvGMYM5EIqc1UucccsqTDTOcWbdNoAaKmu4E+eUOcioPDz17WQ+1qI578HmEZTIQ
tg2kyNpKduFKCXHmUgGRfJOgdhHraORbQgj+OO3ZhMcUjSXUItMIZ4MlajN+6TPK
nzFTmPqBG3cp8WwoqCFOhQSm2cE6bGNfdb9uCQLkgU7F50tyMh9Y7E0rX6Nqsw6a
xEcRmTrwqywywULk+jvcG7seZlPthbQDWB1ZZU+g77unsMXXFD5GigWsxgPMUwmw
0tjaqcRGSaLTadfDjj11WOYqY1yAhYDG6vVvMiTKIdBqZtdPf/NjYmueVm7Gqq18
3rEQesSaMWiu+EfhgMgcARa3LfGnD6mUfYUzMBdEek+nH9Jl17bQtUSAVytyZSsq
Wco/BACGFNAfuA06CtYPEJr5JhRmBjvBYWz8OiMTkBjTZmh+hRZQVAuZiFrei83c
Gc70+aYvw0vpXuCcXfi5L5fcl8rpyvWWBB3KE6UoMKoDAqlAg1p2MNJpDmVKTL+z
gbg+3PACVoaPkrTYyVsSf/IHbMYpop4ljUWnYxvV/3K9vpYgnVG9En8qJHGBf3ar
QPtzVgJV4fDwuEszHsRDVezNNAZrbCSDUX0EWl1Py8HHyXjvzI9XVPEgti7OHqyV
TWmIPHraXO7PLrvtW+Q/ajvnfTVO3YtDkHd79k3KMtYQxfemake5llVj/GIhvq+e
j+riujHlESiO5rnVRGEFVFGM8/Cqn9iMau6TNeLZ2N1MPTxSKbRUYJojUoGQ2811
0JZAiaTPpwYgoSp3S5/t2WEPl2+f6DmCfNHA+7NLlMFcHgmSOuqfdGZPq+1tfwTg
Rnneptbaniyfr0vOuoyCRntboFrCipru8tBqVQJxF3Jh2Nu/9yy5PBUbaIVWmjZu
oYObT/bGaSSiy9xTlgsr1Rr2CTAvpxFKTgApskiSYy24oHHo+j7/7pxV5A0HUmRp
t5P8WvaN7vKS/aggxJSj/B6umNrSYmb0seC80IIO+KfnAlm1md24EmaAmCWSiZyE
uKd3BC+n2Rk2SuokQy7gTBZW4iyBqgoJY/a2IVEtaFOw5tSB/xhw37tBQUTWttt4
2DGHwZkdOSy6HIxG+XCK1mXtkZqfdFZKist3xMuOxJqipTI9K3g9+Jht9lqSoIVV
dCezCLPp4I/83f8O6Qu+AyCHmrTqlyx7Xkn7U6egMjnJFO0ozJEmJk9i9Og+AXAT
B+Lzy1hFSTexMFDi9XHsUlo5ekdVVHP3CudMjDIlzfbCGG68ImxYlasvYi7KzVEP
akU8C6OTwm26pfBGOeDrxjTjDQLV/Tw43RnQloDojUzeIttmlENPTlNIz5b5T1NG
6Iq/TNTbywEtxXNwcAMzHr3PAzKNjsCf8wzUa3N4D+yhnLRKgRjSh3GhrPKdg3z6
cS0JAZvtQxn00r8yxyH2PAchDaMIKMes+ZAfbnTYUgihvDGvf0iZLZKAenKQBNnp
wMs8EyAI1J4vfCGc6SHtO56pJgmA+/7U88CdNmpO30ydk76pJGCL21LVj6NvCGRh
LNfFkvkGsIWxO0H/QMU7nelHT/GVw/4fPy4GLs9MipcjYlY5V+xoD1UzI9//pxBw
xILfkboJwmCm2OovFiP38DO29IsSIDz62kM04Ev25303/mKFrdL5N9QhGuAUBUA/
lQIwb6eOYwtSl29RhpMi1slG55q26e7gsKpsrVEicYRjpNeSMmwiwPwrMJthq6B4
LAfCTOd4pKwB+S53eJYemz9uOJLwCFDxXwQFOjw4bDkBGMkcIc3DKoNdoTkn6v2w
UtVAg5LMim6kI5Kf8jxXAy7do5vBDvs0qoSyrPsoY47nZ2euk9K85HCk6ZLlIrda
9tnlqra+JMurBjC4FXN3bGyCgsXvDHiw0/UfK1C8piaFbxPTGOswrLcbvL3fnExY
0ob+qjYL+hYFQi2IAAVbWZI2ZTIO+WA9HS08M69co8yuvOv977lbtfEkzdGhjZPK
b8RfKD/bBZZU2PG64mHFFrlzbs1H6RjaZVNsnE3l74WmTvf0u2DK+7eCZSee7KSQ
vG/cCvI5CYwh8srQ9puhFmNxQ93/oPGgyIJGo+5oxrFKKZW7uhU7SOYPANXqXlDI
H+cBadIF0sg0jgdiUHJnQl/4FyB0qwxqGJf3azQw/ZPQgsNhwSY5ssk3ivwoofq/
qC8UjZKU5Li3R25txaIQ49sbV5Qtt1RDKDz3PY1ZkX+NhtBxH7jIDmSl7BduCYIo
BtPEALRPb8B2QaylRbO6sD9Xi8K428m42p1dBu0wbkDQpszV3iXgk1RAhNoebQEP
hbdXjU9GWQ9TtFH/J3YJ//FsDV8JqCwSecTii3xtdw4kT04LzrYloDXCwFL10T3f
rneNClKtEW0XoMxpfa9DR8X01IGg62O4G+7gxdUZC6Fg5S7dBComYEr/uRyJURE6
boFKD7/szkP5CxUAwtPuIRbRU3c2b490qT4ipg6mcVh53xzIhkAcIcDcP5VsRK5W
MbnfHHKIktysj60VuWfGD6QtElmfmOAZPEjzKNIyrsbnwesjROXixSnFzB3ZW0zX
gVqgAh5f/wpDBI3S2hQV7ZkYzQEJfJrcK5p3OHMrO5EmzgZ3C0k4LmGyS9cED7rx
gGp9m/X4edXhxCGTR3bIpBGlMo/pvWJdtrfTzL64Juiza+7HbpiwcMzy9vu+Mz9v
ouT52pCnjqRcbi17halkVXUGqtdeOeRy4Ya2s4vAVyC9gut98lCM7zI3oFG3ArkJ
6FajdS64zrYMyt4qjX1t9aTXDIDNAs7sci1dbrQoVjGCollenH/ofDJN1syWOFND
GVLL4dG4V75yIV3qQ8vfsisPXABoWt8UA3JHm5IKzZgGsyme4souKDvaQexNadif
sMBhB4SuvDlwuGei+6DTi9zwl4Xaz28toMC19TJMh17uDxifX1c6kgjrdJUreO0O
OMZE150cjbFMM9kXqb0J1YOoBTJqPz51cV8wMfQkjr1U22+NCxxfi0VZ9xfhXtwS
vJiPvjuRcTQ5HJX4otiWo6oluMcVgTZqvl5icpFq+BYoDxc5cFpcrJDCUXW8bvf9
LSeydXyjTkt+lEYnQ7eA1VDu+FPpM2R0mwsrh95ToqjRyrPLfIR5/hmUoMhKHq8h
57QxcFe1tGq/VJ5+d4kHoeE5+5ccZvGLHVSAf9gBSZMTlmcQuixLQGZNl3pg9GBd
OKrz261t42BfRNdpu2/H75yrP9ZleGlZL0DMmwvG0+R1sGWKc6aVGObxSBWLOcym
Mqa30d90vnraqdYenAUCUNs+9r4rt9uTn/HM4vQ5KNg4OIFyoVf5+nxhmuhKBFpG
cECDq2SPKiGvz6BUgtJ9flt5fAfHwknsmLziqT/spck1c345B3wA9bjrLBM0Ca59
SJsQ3thapRFbdyt9tLafdrIkVLYcAODJ508h2iy2ww7vN8qumLC1uTpFTj6jr07t
LJL/4OYCPuIRkQyf0z73wCHjdRu+BOXRQu4Ue9uYbVdZuBQU1M/Tn3o9F7ih1HSf
fM55IdrHYxucvaLbHMEu/yjF/cTSlBqnEPqYBakQVu21aBNCyCNBKvLgIu3uUv8s
gX4H3HEZvHiyRbovJW3vQOtxXWESdGyjDK4zsmIovLDcCp+o3RK3kxQsychEA89Q
YT7giztVZO+1N4l0fuonUL+q4sfpUg73zbAsine1WFJtuJ/QagkzrqN295Mmgq+3
TdIo9efZ5vvYtXljW1VFyM5YsLlplR1Oikc5Dk9TW8xb9v1FMzFGJV6H/joLFCzi
1aT5bic07JMVlqi3NMG3iILY9IoQYyFB/gWxS3Du3nvenW2jqkp35SjRO+lyy8lA
eiu60ZfZI8+sgFC9OshnRXnOD+EyfrKO8Ul67ygVydWtXFUClV5hEYFH2nS2inFI
qCgxAKS4yjPqCywPs9OyWURiV46AxJVMaBLYuyl+1wFCOcjuvex4ImkT6LyhUr6X
x2IZCIkC1reUWCyljbI5jPmHMClM4gCKtVbUVa3CnC7ufeK326DIvejTpm9FnCSS
4S4Dc0CIeiIYuzQIzWpi/AATZZtplAnwuTnwOySob7MQ9cCMk6yRXvQXgtCrdl3a
V8iYJHR1ciAER+7BggIQSShkI8qIlPm3COKAxdS+fP3d5I1Lu3jYWig5Ruq5Xn4D
U5swIcuE0bevxsHg+8uj0rzmt9eCmXB3wAw+0Z+u+9dBUKJIhUVtmT+Pmv7kNp+6
xa/cgnhzdw7awlGZS/+lUAL380JhckE2wksQxvjXYx8gUlf6XAe9f34mvRX8JKKS
fzA8Y2ZPXLkvwWYfgfzXTKXbKNOtbIv0rG5Vhd55U4J6AsEgb6dM0NZei1YDaQdk
6WZakIJua/0x8lQmgZTQHiroYfB+xn4nlBYVPTQTzAZqEO+U8TF1ygF3/gmXCQjW
d+WCR4PFKuyzh9jpGAS+TZQF7CQ3+6tGBxt/2MG5JjuuNg1djBvxoGVmBw/c3/9x
DSi/Lk3T6tAkN7VytwYz4ksO9x6XwZlg9AF8I9jO4SmsvQRIYqLbc+kJJb2mj0Zr
/xJH4uehT3WTsaRX3cUn0DIaDGtI9c4f/Dp3yslUs3Fi+qusb/8UG89CWNIwA1Hg
hfveekCJYAd3YLFhc+H8g5d+EOGcuimrFZmCnJ0Hg+pKy/zCMwxly133ILBqyZqd
nRpYbWw6zUnm714x4p0HA7URyGK0cM9sEP0GDIdx40XZrjcmrU0gnOgeQmBacOFM
hjE9cXr7Hgp/WXruB8EzbcpuICHiEuDGgwUjVcM7C/myTloyVv7ILYlDwbAiN0fz
ypu7AnxLUYYJQt9lmdrtaSJkDOsAHH7CLLlzavyg6hv9aHzwFI120wsXo7iJCIFy
PRKiy1wa7rGvihugVMYY7vrpMkMQ3mBRGGjfgkvLtE+R9MfGJVER6pg5D/7rMtlj
ef+PFCuCnNOkWB7DKksIwXjb1B0CqjbCpRSA52YaUQ3XagjPQPhIIkjvsUoR5XHo
Qycp5qH4AhpgHGhjFLPsn7gv8LUniLQbO6jgXRc9WH/Qg9j2JzKHIwH5KLDj09we
yfTFLomJqRRk0iIu60YXj4D09uNc4MctnXPX5b+vm6BNfnDLIgOi1lzpKb/tTPv8
wxGRHjX+ChQ4bCfvMQM1wCu6tN/xNbxH7Kdsjf7G0x6++q8fnK8rbD829viUJUQ4
X6aNv8EsSfF0Sq4bTR2b5eskv80R6mXxPVoJzLSxRc8jk/rauFlPvd1qhWOTISxP
M5Q67utvFK36J0Nla9WAKQohLgUdEnZUlW2Ji1RtcNku8eBP9md1LVUy97lc5KHq
6Fv1qs2jvbP6ZYUMfjqQKGqjv8ESUVLEkvkCecmk1Dy4kJblosizLGRpqV5z+a5P
eh21HeMbVEdbo+szXi/R9+wq1hrnlA8CCyhpE4c/LxNkHxz+Bga7oTnRzBtxqFC6
O2jk3RgQSDfi0XEwpvX7qipt4zzsou0Qevt2lHc5Atx+/qdV1OHlEYbduZfe78Oh
b7OYBBpi5gG2ilkDGDQH7oiieBjM+7oJzMamzd7DXPv1gwS8/F0NYelBvXt/nnZa
b8JqJ9MXpTbGJUxUfvop29dZ1yaY4WPDuYHjpfkyZsqAPhyv9f96yHbcrnihLD2f
NJLYCXXoyXoHDo1JCuiAq3k6FOTjaLDkSNyWN3JdrPJBWquFy08U30xnF3YEdpol
68XGpaHtGwXCiRpVm4kGWsUMx1JJuVGPiC22OesTf6UNg7V1G31y/SvYn7h2WhcS
Y0lodTCj6Z/DrVL4RqaWgNJOMTAgLUR0tCoRalBy/bgCMeoHEw3BJcHBq3/Z7R27
gI5n8FVQ/jnB/UaWcu5M2xtQXTMvd84bRbb/HF53zwe8TiJFfadxcMRUoEdYq+6d
kbMmhW4zKzcCVcYZHpe2OepY8F94D8fzwdm7/44DH7H9UyItcdWvr33CePvQ20H/
ga55TgW8tlTEdwQnEFd+OVycHcflgllgPclAN02ImsBB533PduQr9e6YR3TZPyWI
JgpotNlSF49j9UwH3WiDxJXWyHQffZXlG3UAovVUVMHEHWwoo2vP+r88k6FtJyUp
ze82cgY423/C0I4oV6JAAf7tQ182mGbzZB5n1xaVZj6ZU2p34yEiyyW8SumrR8v2
AHfPEwRHkvlARiB91ZI8j2F/CVllnPSQ2Dlyy/K3XxQ7Yg6N3ZDwpNDxb9QNQq7j
4Ani5tMN6xobObhhvUhGvvGOClPymLGvBbubKpQTT9nqOnvwWChqKz+5AlDw10qv
0/tyDPXDqyqaOwKTjpGuuZ3b4R7PvfXyqzkLpPEVtv9RnKnLLVwQTZyyEDUg9o6c
1szqhl01Nnss2heMW4hEjm+CNXnUkqKaxAZUv1V2TTjIdmWxG/92TPPPZ9cTExF4
aSf1SGZf2PQo4tirdtJ9UMQgAcUcPpEndjYRs+YO55lV9kLEQfdDik4UtqWxeTFq
VtIUrPZ51Cr/3hNbUPGR/EVwZZUNer5w3/b2e+rYGwoWneKn4KgWonILhOsBhJ6a
yblIRMjzuaFqS79ulsHqHIA4IIuDTax42CE9sVQY1PxUil/t5Q/C7hnQkEKaM+Nm
HJjGsW0+p6W+a6PSoKEj0RZO/O/cYYzyPP4WwYdOXGmp63d41zlNuKeJLtN8fz8N
N/JuNbcnH35u2bzSXNcqMGh879iaKYu4EMX0IDjGyFLcrtgGqWyFIMhqWfBS7IF1
iFYGJym1RLej0mW5ZGN7GYIq8Wpd5mYJ/tvEV0OZxmDdZmRi8VvSFkG2Z8rwSpgf
yx7HmDQ0V1mFK7k/cKcWDuM9pO7wVQylLeyeMn0GbDgDdYA2FyAXl4UQWdCeLuhr
M34y7rSnsaUdXszZLTexMYAkCgBYlewqigpJLzqfIX6uNGNQIi5hfPc3J9QWx/wC
VCM9d0/hbQ5X0mGOBjIHXmfm/e6MgF1pidm/IuEG1Oel6CUjHhIGKHVwTIgumNtE
ORB/yiTgZSDeORmHO65mr32f0d9LX9EdgwpS7x5H6K809Zo/z8VnKXxgcEBiDwKq
nims6lBm3tj613YY1zDPamE55eEEzEIlV3w8Snv2KFezHKavIdKVbbAxFnDlve7D
L0qDPAXKri2Lz2rnPDEuIjxBAsi6Dkm3hSTnRQ6I/m/8RxhYNi19EfiHsgOw7Eyr
LDYwmS+FthpJAQurpWONjuKRe2lV0lVMONyqjqYodNPE6QxKN1F/pP7zxmfdDSKZ
3HknRZlHdLJimOZmhrn7nhggXDRNWzUH3M9sxQTqxojFbh0OV0Vt8IEO6myIVIns
OpTmewCLZsd4Sd0YSDFy+m3wCFY1i8WUUYFVg68slHXkN5YTpNMU8NziU2RbDozW
CTDXGXhceEDMWn/KPnElpGZtcgX1f9ccfCVEcer6G3KysYyKaSkhh6HXRZEZDodA
17vEEPimckofxJyIL+f/D7Sg6ZkLCS3UhGrsdh92Fxi+gJZLtsdJ5VH0eo6Whbuf
H3beVpS4L4pnrTMBGfXlC9jhYFRH/whrlLsR+2zmwYQ20aXuhSSAKplXT7BTuili
m6E/mDb4VgcOGyLt/flXhT+No1AsRWVtNjD+lJUcuN+Xa8K83EHr7gVmLBDrfgbv
q47EoIkRyoBJb4nUh7r5VbnicFqXNjDPEe6YzqeLRUhr3T1agO6wNfEmkH12hlPY
ATkFf+VY5EcbF8tHUgewLEcvq0nlTS0Sh2w3hr0Ib48zd9SZgzd3iaGWwxpg46T+
J+VSI6j0Ch1jy8m7awr2dKOSBAnVImXmocULcGeYUhsRA0IOjFPGLDXgiSv0W9DU
xleGx0L8tM4YOnrRD3/SUVohxPrXjvaIhUqlH7WWeNFFUyl6nxVx22ea1x6sej2o
6vd4o6hsp60nW4saMMK+5BQyg16EluJpd+H6zHLYKOcB47jRXBDjRXPHIuQgzgQY
JP6YEROe9skq227L4A2GTNm8vaW6mD2uedPN3FHLbscRnLyU+G9tHqnv0Y5urWL/
h03nUu1R7ZkZf7JsoofymKvM1VWgoTcUk3uDNGpG5zI1o32D9NY3fgTHl8xyCsUu
FpAozXYisWf7GRL+JGcw0lpGyKIV+z6t7iNlIwaLVQqz2W5OaE5HKnh8WUGUwca1
azlIPkunEhTu/VIzQB6T4Wngva8iTXHB67KqXK7jFGKHp8ElQLBd5Rezln5/Pp+4
72s6GR+B5ZVURWLZk7WaBratL8X+G74Fxker9R12YpJu0LzN5/Ptw6niDegq/59x
kZ3HCrONStT2p3yCA+x/hKii0Jyd+de/gsyAUgvCdZOfb/8FFgpokBXJu/4E93QK
1DGANtLYhDbuIc06v1uiVW3SU59KVJO53vkK7Udb/MP7YLL12T533DfHYkqJQnuz
eC4GYKvn3e2y3OvbW4s6cL0TpFCqlzu/hHb/TKJpu1+TVl4ZQXPt4c1xjYVn9v1s
LskoThmSKaREZyJ5RKFBQsuHZyrF2Hi4ri88ry8ciprvtHXCg+SHq5b7wAZbyWug
/J7qPAL2Vgxm9Pgj3YNJuvGOPdDOfd3ceRqgfIMKHEOHzk3spuOWrE7cAsFlyRjm
+b9YAtGFqbX5sIEcFZaXH0xonKqypx44kF+cGV8k7tnsdLOdPDhJJwicl9q2sldM
utkFTAJdoJ4Po7CyFJcHTtIX4wEZ7CdmTL0I5H+NLODgivRZEptflwrza72ep48h
vbSL3DsJmmEFANODVECO4A+jK0vo8SSF4qkUMOJfsGdFIsyz/GrWoNi+voEY9af0
0FmSdriIkOs/1W/As8IWz5hvzU4/vXfp2M+AmCC3cOs3uufKO2Z7koBLgGUMqTPk
03WDWBy4O3UjdbWNn6/WHNirzr6cjjtlzuChWw4FKSTwuDg8kvv7QIMtGqV9Q4Rl
DKeUvcV8AdaG+D75Fw8DkFxFALMHN7eVUDKrqLPg/uMx2wSm02sm+40ua1hNYTF9
WVr38Y1Bjv2S9jjUBTO4EUKlSYr6ARgoK/ceHLSk2MWA3ZsUQiShmZy8y1qN8Qzy
euHvGTJArkVEj7sxe4Ym2zcc8rfG0VxGw2sri62hKjengxq0S05xkpmu7ykwsXSa
VpaKDu7DHj/5uon4UH7w4AJ/7LZyLMJc3ZjXLp9D1ttO8qGL3rAD7KFdFjIiB65B
7fgTi5CoHay5vnabcYnFUUfxmOg7XViXy/KQZ0M5ZIrOUyWOLjOGYNERYrbTJIn3
VylWuc0TvO8cikUxI1Ssih5i3c8oOX+sekQVqjztJrYHgYDf2X+VHxBFU9rWHbni
1gh1zb0BEicM6AJBClkNcBVrtmZfDrRK7th95lZGN43TVa5WL0bkBLEYUCA94tRt
akGEbbRlL+oTJrJLcrzBo0kwiVYt4qpJiZGHLInv2JEdF19+U9JjFIyB0lgOYZ98
WLp0ymT/s+mCgcBG6Y1x53sRce974WY9KLSClX+V94y7gCkEjFVclSF4AV4iOlaT
D4QvVw2Ge8m1XV9jBQGuFslRkLc/PC4puPMkEi3eXbchYheE0JiFJ9gx8YGh0Qb+
CHKjsd2RPu6RRc4Je158B3E97stKVk2TbewbZR2Z3plpyvuRMiO5QJya1JPntYot
u87QngXkJJXaNHlrk77M2kD1yUUeSXivDsEilyfm41Ijc4krtQdicMY05WjC74Z7
jZ4PPLlyxU2lQff41DVkjxQriAdRc6H8GF0Ubgvtq2FM+Mnj3j9wW/Yg7xsfhFd1
GuMGto/pttNUtrgF3PeE+o6ElRNLBucAYM2+rQ4I5sMItskhz0EWHgeYRsGz0sDH
oVas5SH/tsnry88l2AsVywOifGlKTaf1AdZ6GFPor5B65q1PmT6VMZ+G0WNF4RXd
nAsS0VCE8KrpvPLTT2XEZJhszVsUNo1zmzFe7JNbjB7oEc8OYA8CRojJiVegbLNm
3DuYyjVmMwSnIrIBsvzKeDhZPNzcQgj5wl5DXFki4jqk0nunM868LSMgukXz5Ehu
IyGyUvcaulBDB+t88yRnulITLwLCbkszc+I/z6nfO0ILDzwN8ZBb1oepg2CBdiXB
GWDUAcL4MWyHs3isJ+yZQXSWes7Ub76onc15ecZjyZZtrkZa4R+mUTZRQ3kWdNJj
BoZ6u+zTctl9l+4Yr1tw3oZLAXkJ9brr6BZWhl8TYoupHZ2mRw1iBwz60banl43S
j7tKvfx4muQ3nCtNrmBHAfOsoxZ8HFSkG4aG12MVZ2NwiWCk7TEwvyLg+KKL81h3
bz/Yuve9n/yIg5O4LYVkwR5/yTlZQoPC+jEEobtqI94BoC/QFeSgEtaCTqlUvOLo
Z8CIIr4aUAmklCQ9qJl08wQ+5Ql4w1rCs+kOyIRbkWfcpOwwv9NhCO3xOPdIfN7C
2//mwV4Sk92Y0E63WeYLvIyESOmPw7Lt3kkzQ0zUrriZFTeDJAQuyVObBuGr+UK5
4bCUk681sZopxK1AsOFCGG9Buehw8F0I+Atsd76rPaOWgc8bvq376KXNxkP0NGjA
rcLRQQg1vjcSD321h571MLKcymTCsV1Kb3Q4YsuHDB6Ldz/IUVNZSwZMEFP18d6M
7/RBwPS/gBiYTyLxs8G7jb+oMOzLTDFg+8q3OTE4aHV0SfDr9WBVUOtPElBBjT71
VHDuZFTTps38vS+MBE+ff/FLPrI/7e1zLVK1KC/3iDcKPD7F6UJHHGaRZR9l0Eob
gR8a+z6zGJUqqrYYNf0nnqXxklN6Rw23nwToG+ivIN5jXFAAYQ5a4ZoIwVf5zbpn
AaygQgbNzdVW9y9n51Z4yJx32V6vaq2E57TGQBwzCq+iZ2HvSb4gw4SVhEvnz1GV
c+9yXOTxZkmvGvefRG26UPQOhWGaJmEOMGBAbLSrdJbILpjXOuM1YhWwHpRTbMGy
Zet2rf+h8g53TtsHcRQPUnTDpbsPo4Dmfi2XiZ414UejsatOr/MERQ9gyAt5nt75
76JAiKj8+nCpheg5CRAszrVrW45ueXsdveBebN/3jfOlDWwFV3zo4sX3ynZ+ga5n
Pg9Byj51tN+B2+QMzrhjAQ7Y5JdEiDK6DEM6G/TO9+Ez2ckeOcmeLXe74f/aLoyh
IGyQxwzxe0uLY8+P1AdA1yZwZXyHFOQIdIVUYMkD2Wo4z4xOCk8xx1PcZJp/8F4g
WFlMp6KOCbfb234l/QcArL3m3TyRFCi1OEPOK6vqRA2qnslGE2WNyMpcyogV4if1
sXPDJaqOf2OcAYAULSL3DkCakDVdmKZA8k3E9qfieIq8xyd7KVGLLV7EiS8cOPbM
IjccU03mHkNiYYf+VmvZ5HyYYvgoF9eKiQ5qmyymsUimT40TZGyKh81jLmYs1kPy
BosvWBqNAvxUzB/75ADoZOBF95i0y09W4Yhpjb+AX0WDav0wfuvGhr46YBItUgtH
LHlWWFSpzZcEeqKAyA945QzoxOufvjJgSUOlO4lI9MOMaSuaYGJo73LwAueTxO6l
3TNWupu3u6dR8lUHBdC9NLl5i/miSRX0uH19422Sm0/invW6Y7VbCkaGRr4ppgUp
tbKH1YatYgNMU5SOlwmt9RKcbkBjs+rkTI/3WxqWJMInZEAUCOPTBDukpLacKnCb
No0W563ffOVZE1HKzpgIUZWfdHbhmfU1QUBDXYJ9DByPApjC40yDe3NMW+k2jtvy
k1vmiNHBUnv5F3e/qzciA1jNKMdnIMqE5PqV+PFhBKhn78TmmPjfKErSTomGPEdQ
baU6vqHXbo+La//UNCAz7qPs0JoWO9gal3bD+bDQdFNMQ6adgTd5OhdONmIrRyBt
H7DXhjnjVr6fV04BB5o7JcjSjYN85h6Bj7uF1PptqX4y8hXBWmt+EHpDk0PxT9ic
ONHe3dy2jEXK6Al4g1WdDaUoE+CTkZo30tBcO6NFWfx9QsJWJTK00DE5Pf0xA12l
qhxPyTq6kc7HZY4LIIUuSA1MX7pNvrJWJWxkj1Ej+xpUg+5ElYL2jZg/EgFp/+6K
RNbfCkII3dFppHdWiF5M6qFx+yDOFoFY2O/v+gg+NaGTGFz2asghQuKPKy7M8p/D
u8iNNSoWvoXoPfJug6s8LJZTBzgsfv9Owj+NZo43kKvkL57+C7KG+9XhCF9sGMzw
w6kLcPj4rSB/rHpKXtvB0CV4o2JS+C/6x3bpp/vzskMQw3VapqatEon8c1yYRLyF
GZwbz6VisinIBilA8wA6vW32PPR352Qe5NAP/2tpycq0fdDbz84p10IdBBpbZ36y
D3Chy6Vty60fSdgpFBWp5EY4NWgqpnjNsDHKHs2evGLpyMtkXi+VUtZ9sgFFzIj6
qi1p+E8mNY4yfEBQN01IJI3vz3Fjn8HN7Q3IqGVMxBhDiwJtJWuHxrUFKUHBqJKh
R8InFwCyVan93ShNflYOrqKlF7F8hLdrHWf3DBEHYcqujXPYOpp6htlBMlUzn9Sz
l/jMeV03JS3kYLAqRz+gZqicKk6cQCwkWNhcl1GpacFtLZi6OfJvsC33gWwGa+cC
9oGfIygadt6RQhti2X7erhzEkRW0y4HeUdD8J/lmh4NFGzgwxfQwNqxU13+FoXcJ
gSnoRVLy5mx5VDBpDS/2u6wtfEdX6v20ZvAWeym1TYoDDeztCjQ93iDs3LvuhaLe
w/s92J5attbKCxPCCgYBgcQ3MXSjsebqMb5yJ1meNnH8Ok3XNGkj4eN/s5N4oJy3
Qw2c1AfYOYhz20p2/D/5L97oatQSwSKhaJpgAqq38yipsX4j3E9E+ntMzJefx+b2
kDa6zDvSAUpdsIjAMCRK2RagDUHVcopNP2+z9k2KKVIYe6GYRf/NfByb25JY5Dr4
6K4vjQYrDg2EtkG4dRbNtmkqmXgjPIjqOuN9gHEZaDYqtz7LNP4HEVDoyTTd4JGX
O0/q9RE5lFcRivoi/3xNW8BHPqD+te3Q0M1PWGKVNV7YdwqsrSArRRKhFkWm//2s
dzIerloCeHwEm7lPBu00iUHe0cbCfvkLMKOIIjYXwv4MrkjyCcA/zZoHAWtn1dVK
+tIWVz4xms5hqY6x99lC3BPC3SOO9Z19wNjlfzhGYWjGCYEChpo+jFMnA/niHoVi
AW5+ld/dQVD1dYbswq2BqjRXE+7bxnwsQ01X+k4KBb/2bErI2M9eUVNC64qjthJA
pTjl1/15775vlgD1tc0RL+xtLixaCTxT7VUBwhGaV0SZUxdWsMMeqOIGFMHp1WJY
M6bjAT+iIYb7lrJ++v/dVyPRVnKRilBw5cVRu42IADkHXFRptDG8NfTtVavN9dg4
aFSh4OPWcy8bNgsulLb2tmfaaw5sqzAASZJD5tO+K/A4L6lM15AQuFk0uyTClOqt
glnwvPBQmBG/NkmoPrX9Vt4HlDW8/QWGQk85HESrYvE4bKyQ1CyL54phK2ErxGyw
WIoOzGwamCvVZ57cQgXOpdWt7GNcQSHmuSMJj7IgT+4Ks4rPIZ5lcRwIRcTmmHOb
R8Q6fe668myzFs2sjLuFOlbLj84o/4D+WBnO5G9rlN+Q0ELcJK8Oc/uKeiVxlOwg
xf+MKmr7OHQpQjhBt9KO5M/hc+iKZLq28yvKKsgxvDvHCLPl+XwTG4Hy6Ot31Afx
2FDSItkJEdFX9g2fc3s3yZV71ANw8E5Di5qdmfc5uhotjra0hb/CrqxUwOTmy2wV
RbJB3FkiNdvntq5BnQUAibKf7AxWxAAcjgbZ+p/TWovcixaeej4r/5gC19sZMXbx
RxOdBXpK+/3re0aa+h6WWUHPpMmRcgqOpYz/hKrhnPYGHqLwbxfN5OR9DzD0jEUz
93nA+3H45ziki6gNzOSjEXv7FwiPnbVCQrW+SG66n2V1l73+/jBY1maFclXpU7F8
wA+/8RbELWAFVQdLTHJU0jGNUCMr24CNmFQKXaWZravD97Wio3NB053D2c2J5TDH
1UM1D5xjWWR+973GP6zqdcQpNI5unlQSK68MFntWEEW4Ydm4FjJpeFBccq0L0oMK
IbIxwt3Qmeasjy2yL0gjLqCTaOvpGRl17VP+QGCErgd0lG9wa0kRBhaVTt8JpWoz
U7Ljg7iHXgX4o1Fe8YkFvZskStQy56Bp1/gJqJolLkGXNENwgU+jG+7fIk8rVpPG
nNWV0IEBQvRmPbY3QowR8rjclvI28urOZe9aHcSAT0uJeKPpCNjNtUoWjEPNICua
2q3Vtm4UTS1jL7KgmcPKY3Xb7o9MteDgIY6Uygrxmh5oR9Oe4A3fUTuOomBqj80h
tF6y0Fuul9mOP3MFqkWgQedXhTVJ6Q+NXLJNkcc8wRNwmgZhyUreoFh7rBUtxCJy
XiRxNvov3rk5LQy5Xl0ioVF+A7O1ecM/T2s79G03bsOqNFt1LjRn2Q4GZ7djLJrp
rpWfq+eUbmXJOcRn3QRNnAexP6aBkNb69Bwvek3GrliWGXQHtQbMePPCclZgo1v1
gaxuw14bt5hV20AcP5m3ZnWXf/p+bLrlXUFdAk1z2ENn9dPKh9RiWWCqZHlJ7EOP
yi6sO6B78+kPF/o+jDEs5yxJS29MOlejqlTfi7yuEFlRmEg/dDE+WpQQjpLoCM0n
eCnuGbRPXGWbjKknSzrbP4zWK+5YjDqfwcPapzZm2+D0dlOElPQmbdTURopYZTRq
bbqzZtO6BZ1jhidOU8YDZayZUR02cCvUhFcpCKZDdfM8BBrpAnlVUVY2Apd+B3EI
BhjW8iq1ZfKcR4gHrZo2SNYyKOnFJdcxG1uI6xVamlSF0kpyvL2x/d7IhBdhhuyW
lMTe7HqHWKbVDAMFX9W85YDsfXnysQeFfHXku6OmfTDwMgbbXQH8DJfi9WXRnIDt
JopgmryY/3mhPVuozc3bF471AEET6qOjcXVHPGAEm9ExcFB59Bgf6s0Wu7l9eZhO
gdVkNqxtJSbDFzVGtjDmcmnacIECgnNhgTpoaOAk3K8e96lLm6daf4ewJZzTQujo
u4XCIbpzdW1pMhvgPaU6HF3KAEFFfYFeqMmcBf+J24Uy0AIYLwxHC98eM2ZARzSG
u5oyFG4XDxC0WyHwKi13vJtFE6xuixVsWzsUXDK1yxpcjY7/Feq4dwyJSmjVUYgV
Y8vypcwVqNvUimqXAlN6ltC3CTxtopijYA3l4hrbFNIf8k7hoKaCzGJVKG26bGTc
ThVSlB7wVksJlbeqEQi9DQ2aTYrIoKa6L6H1KeEvUfPrLi9ZgfBiDozHUPw8RbIF
3omiTCNt7K1YycVipYP3Ht/WefLXD0rjYSpj72MbeKhPIyQcxBFYY1jS/udHzRrA
WVqgHUF7th1sz50gqi0v+Hs1a6hXzRrflIcj4D0H3pxpourA1N5OVoVufnJHfj46
P+rdjwbQIhZgPBOsMTuosCgUYyAc9DHWSWrvSNtIwUTEiw8DNiD1eWsPoF+kc1Gj
zTFr3oDEFErWzde3/ku5uYiJUWvQGnyDUMdWYsbSUBSc7oeaZnQrEYfVbekGeCbj
zbRCLSD2ZTbeIQBRw2xMlA85XokmFUC5/uFDuCTVR6yDhgm+96r6YjT7zQzN7+1R
H/I9fdHGWminXerLk3YJxsnKvrUR91Y/hz6aFYk7F9sQIZI3ewC9/iAo3L/40B34
zO0xoabsDxY+/fwBlx3J50pmoACvbAnghIJ5qVguh+oV/2RVCIG39xG7bv0cZXGo
cVMkGWx1MmygSuDPfBQC40CUw5xp4PqCi1lDeXp5ShGFMVcUugjZRb3fi7klWAFC
geN6ZtbudfhM1pe31MqwQqeYzBB0+hz1swu/LQYo+duCP8QdCfGEWQjKqU8oD0xo
iZW1S6t7pYIuzS0c4OLdMSV/RFzKTuOe3KNHf8OkkMBkTj4ZNsEEY804toOBHu4g
6Rk+rdWiLbJUHI5HvE+gMD2BLvePNN2loiBqAOUhrHJymd/D+h1aS8eCfSZNVjix
Cdyfk4H5humTcg0g5lIiZBGGMBrtlmU2wrMpooPZX5Sun2fcZs4KQbMA2G3KENIY
a7lkn231KuAvZTz0VewchNmg9zWwDpkpaXLQ1WI+2CsQZtPgv+CwhyIe7OdHxtNP
AUOpc51/iIfI6zpIGVbUms6ctu17KB5h494B1vLuBifBGZpPjtjsyPIYCC30rk/O
a4o8PktpaaevPGzWIQJbae1mB3S/KQrOZrjFd6lxgwWo7RO6CmdCq2xgXEf8wFA+
F3C+rTkxD8FjQ69+M8y7QMTTXEeM0pz/ybWKWy5vRk7RRySEZzQ0UeO4HaOwWLS0
jd8a8v+Qp0Wg6nl1+EH7g8A5KSCF6C9CBfzrPMOEETWDX4wmOw4wOXYN7buJoEpU
rE+2tPuatVV82rqKxzbH/D/bi3vm4UUEB+xHw7LlzMI4xARCfHCB7DIbbzpAzFjq
FPNUzSJEjh+N3LlqmdTfPb1/7mWxiN77NfiJuPvfmbdILQCFiyP0WBwhuWj7+13n
ThcdmNYItBrSTDehV1xNeZNUKVY1CoT1T7TAL4ahtec3y8+4ZE73v6926lhMrMp/
yZLNQ8KwUXoRFB3aZz2UVmncYEVoEvVg0QQTcdv6/RtBm+b1e0l9ONz+0CMKc9LH
/qQ4WBYtQ5LL1UGSrmy+KXFtnXru1Pk9jCma4O6sz3cqgMShv1FDFv+bB2idNCNA
EWIVeld6pKh39zAKQsCvhKQ8VbFcwWhRpzgW4SgarGJOf/fAXR8PsRkZCbdC6VDQ
UlfRBMBV66b7QN6Y0hAtLaNlQH1ifDPncpnLRajgw371crK8lSdBO0jw4CRSfY2a
vWj3yeHH+NFXthFOc3jvja/DYS9la9cqP7BTbjKNO6q2hRRnei/z5bxqG1h3gKzd
2bom/8jJpXENKXtHRMfc1JI1lEr6vuUbEXzbiWN1Dx+Y7nRCk50QVtxO0oET7yBV
cplOB8eZzMGu+P3BzLBj9ZtpdP84iklt9yOzhQdVJSPunbEkRou+hGcr3z1jmwcl
bgTGC9kO+p4wjwNj4rmqN+HxKDgzH6k2eu26h9litjpNNgRFC+qiSGX7cn1PgAY1
xc1ExQjKlMwLdRXmup1ME5lwniFgjFg7zImQ7fi8Uq6Z7sVhHmq4Tfvbb8GaHIfv
tIR5Ty1pdnZYgAtxb425pWmT9eTd3E3azTLsnh9cKc3oYIhbTPzZzS7FxKxH03vn
I0/T3lR+czwsSDsGv8ezUNH/p/2fHueSQAPT2iuFfF3E+W52fnavmSxjvyD0Xdkm
kMIAugIPWNZST1A6lMFp4PbGbKbNPJViq4SERM4r1tA9L57unnkoftwvstAa6ax/
wFV0BAOokY4BCOfq/RVzWszSmlUvCmMdiv3ScSBx4RRBBZLESch2cpCgkIbP0pbo
ovx9aX/Rjkhmw+cSOwl5NqhuBPe4lffuIbdQ+e9Fi0oJ/o4Q5c9mBwnVAX0SD34u
ya8IkfjwPSZnFdq1ZWsCmVarb93zxY/1LDioedlZOxfrfEklzsjyB6b1f5IoBhTu
AyCCM61U8WZYZiZxFzxA4KBidkiG/+OdYP75s//mzKKHBuZ5YfaTiVjfNbY/IA0+
Bd8qDRfXTyr5Xhlq5WlfvT2Cx/P/q57CWv4foTq4LsnB3Dkb86K0RdjxcYAzH1cZ
6mmv+3IfiO8KGTfr4UdVeXn3o0icO6gOkAf8W2Lk7xG/aJxw92DJhXwlM6jWaLBg
u5Mh6piGKNbLcZQd/FlAxwjV8vo9dNE3PuCR1LKFrBrhrniSKIST8zdMIccJm1Ol
7ozXCk4qCB5LP64s4ahI38qs9KAKNX4JOT0wp+0bPd6d7Q/2Mp+oevyt+wBsjuYR
zK84euIM6JB9XQXMjjLTHU/1wCs9tyUzmq8okzmb/JrqZoKpGJS08MunZrjfb+XR
Do0+1+NK3lPv0c73UIZFz5+wwDzd/Vhyzq1K+UHvigcLBs43r3kSeWf39HCLVLUx
xKfMem1sToplT4pGGIYjjpHi0WGLmIT32xHM3TG3gz3aIjaDvdKSCAGvOiHJP/c0
L+fH7TyJhLMUWEnXuYrRmf8oO0jcxBtK9myeHECjB7MAyJ0aUHOECBwBoZ+m87/5
uDvjfwV4Fs7DMpPsZSLPdc59Sj6/ZQMnigbKp3/ejEhJOTZyo70uXDchDB8kzgJY
p7Ysz38xMHZlCSDuUMPm5YM3kMsyD22HcLM2zn7k+9aLCax9cEBfZZjrZqI11m0I
A2Fmi+Cfz6uSbmlXx82QUZkU6Nk1EfqTwzHUn+Q3lXW6flVtAMt+Iukaic0JaWVb
mM+Z4bduCOjVhuhsxtYJLxmzTCs8VmfaIrq3wTszaJly4xcNB9Q5KbSkAWsuJB79
GsdNlcf47hUiDmUWlV/F3p7xIc6mD62Lq8BFfdjJuyDSAMSOvqDwcRdpw9MlVdEw
Z+L32U7RFfNsg/ApD+jXvD+qNcGs7yar99OGJj+T9EKZUF9ajwbs+PzIYPa3rflv
dYJSwTuwxcEQp8UoMdHopr1LMVGCHL4fehS/VLfR5n9tpFwgJeLddcBNGgCaui92
NvgYiaoImi3HTb/sHgjBL2YaJrSLPYg2Eeo2mFJk9muw99x+eoAFKUM60kUYh/Nd
7s/rUZ26JX8vitI6+SQFaX3QfIZW64TJBtdtHls2Axrgjvl4tOm3PSdIiJqg9N6J
pegLHep5ZQJCu0lVK+9JgvDJbVelHrZ1ZxMQ868EOEBiWrOUrL5CvQEDzMQMy78b
4AOnJ2RS2p+hDY+fkzvr5O4xn6XfXbWtlIlqvHTx1IJiS+OOwa3IGpc6TQwqMUJo
bOaVwD0GUprsNXwHEHZJt4LpHFep/DPLHjurNgtgw4BY0qzxD8RvZoEeSnD/rLCY
snH6haxN4nao0p/8IPoPwCUYj2KMhJFOSbICxZjz5XHNiNI8qMi5hyIwIdTgV+gO
oLObKY8bElTB6DX/9oQiNGwsV1CHrjaAEW+FXE+49/NnU84o2HXuxoPGDaCf4YN5
62vuiTIesIm/OETXnDOZG2cGSK0juU0c5odEgXehvm8IwYp6haIFvUW3HWJV7d0/
ehqnLcgk1zr8lUL6VPWniI+dROBLGHcjUiOV9HZjMU0NdOCwuH9VL/QkKuI4+HGt
pbgFUp1qQnJ1NVzpWlBcmOnP3lNBdPgCAGP9K94YIWOBFnphi5pGryvQi131EMVp
c93CWRN9bVXD2aSNDywXJiHSJqRcKzUMjTVzVp8D9Ac7FvD7xnoblnMptlU9wskE
24rSdzUbwwLKuO59qUjyRL1X4nmvL3PLhOvzV8a/+3z4op/JI6SDs78LI09fkLKK
RgMcKlDUHC1NgC1ilT2cI8GJWfei+vCqHvF3qUZKAB7oDkS4uwbiGXBRk9hNsXON
ZFfK9tBfQkr2BLMhMxyWOUV8uQD0cgS2FqbJsRdkkCMZyfuVmabamLEdsqYnnKgU
z1Y2MvtYD+/6Cnw58SG38kbelxH1JVnSCkUxB2vAn4V1pwuT92zclOZYIYu3YTvL
57w7urhwlaZiz9v9khV7nhRR7iSN4+m2NJ1dHXO4ucUFB4ajqEncJXdm99TZ7bSN
fhVzSbC0OfSe7OISRtMmg3Ldhv0+vXTL463mgw69SHT5JOmXaMKH5mf8t1hilgpi
UcCkDF19UIInkO4yB96VlbI6NKtGqo45OPCUq1/NDP+m0Mc/xTPHcyhelM7MFDFX
xWYmZhsfNc9HYrpATCMLY5l43f0hwy218NJdaEESq9ACiTrGQCxTM+yJhYsRUctM
P+/C4sCgznlMUeOzPMmTh78PL5fa1Sv3i8LFP8XvG9VCkmUgHya501u2gJe4cJz7
OouT0MZ7yYOv/C2TYaUJ64zjwt9RW/DXd7mTYegGB5kFOyxkMzs+bnX+UsMyps/a
qSS5GDcZKBueELlk4I1auVGzT8dG2OWxnWInUHXVyUQAfT4/l8yv8DOadvhWFlod
Wpw0yQKtRQ7bnIUEMpu+pB6VGGkN+uyq7zeyi0nISD9aWeB+aqRB9hg4o6L3/d6c
wvDl6PYJFV3eVVIVS21ymu9yEzLYWlERAB26OASgMSTSDtJLXf1Hbl2KjCeExib/
v8MpT2wUyHc97fMvDtHLe4J9CTHSm7KdNAZA7WatkhRLivOOhr6o0TbusIij/qe+
KaDz7EtATig+AeLTsFiVE5I1IfG6WlR7IluqzBSxmjgeGtDn2eX6cq7EyzXq10rI
8jsU/ey+eo5XEREZGcTi2ujXFcUPA6sVqiPfpMRc7J/gQIKLMXmM+CVRdakq55M/
D5awDsPgW3ZgniQsILI7eD47FhlU6LFQpOCV8XPxauRzMiTQZAZ5mP7chhonyvW4
vwY8oizplyZccIEiBVzryOSu3VidOzcCqxHlamTY2ushOca46cnfyccYXxZTc+8+
H9ntnD+jNhEQrfFgzF0FRRM1c61Pu3LOvmhIxpkYUA898r8cfATvFyXrTAgAPTxp
MHaMaAMjG494YXSAaRQwaacwOjjPawGFceW+lVH7+K2c3VurNYE4vLTZUyn+XKdY
Q10QeV39QrIEfdpYH7WW9eCbsVowCRL/FWQkzMB2ygUiMshKfDX29tq3y1NlLaV5
ApzJ2GTLY8PXplhDM7clV7crpoe2HaUUbVik7XwsolqvfSrH3ygLFGdEwSRQGXiC
3ZvOwGMnVpm9vHRw2nNOrVzh5tcte7zW6Nr1dBOvh9kMiBQ8aOOJxFpQliIt4xvc
6op1GDcTxla2HF+gJo9bccpaq9+dNQC0KkEvPux96Wkf6VzZVTMU2B+jg1a8Jk0n
eCjreR8A9OIKZ+ipVX/SzRvqXZkdsHEvptb5p+qlPTnSZtogLVH8+ZaikhHe60BR
iYcY4Y6wGG+tgafEVBEPl81Or8z62OsgayWX+76QsgoNPfSr1AEtIghuvHD1ZDJ/
yKWxlPBwc+uN4BymsTylogENROJ4GwWaDO3PaqDHnbH83AOgmhjk1FrylmLsWG82
mtMWey4pNJohSjlesLTHVbmW3XU6xiY74WYOuBi5jhIYTtiyBW3xJTBXxaS7lHhH
h2UE0C9e6MU9PCobxNSuDKGpZEh+oyvQQjDF6sZg/S4DO9AYG95wG6Y1T1SMSZF7
BmSCZ1ehCUULaMD/pYIVN2XJs8e/q2660eZMTJfzkKCzI3lq1pn4LWVnvl7VC1T7
ZqHh6Rfrsy9hz/fmrSv1EFL/3+O1yD1mBncEXJ91hOy87VvJEvAdxpnTHySFoPN7
JfoZMK4kwQqiIePNL/DJESC5TNWghWYYuOFbYQja91BwbcwjxusFCDS4TH8b0YZl
HPQjQj3o3Dw23Bk/lnfKwbxBZ6aHtMJnXr1olBZISe+YGADOg6F6Q+hMjE3SmbWO
8qC4b1sWzRxm4Y71iXAdYS+HM0i71qkE6PXhjQrmAY8uXoDhrRWDQVeWLsOVdeXn
zJeqCRIta00ojrendlNXqyLi8Meg0bIlLN9J90uUYFhEgnnF39p0Ne1oDq+vwmur
1fIny1L90ehLrNqQw584AgwsQWhIzsue/IRjTO2oF1kjR/u5pBwuEJWROFWnimE3
g+I69IjXOUsZvP4O7R44ge8gMrS1Qw/X3EWB+jNJMFJe0cFg5pNxTNJxJrcR2EEv
/aPXaH8Epr4KyfkR2KoDq2VgOWGRvVXtTP55kzezQfEc9YqpJOEx2SySIRQ39mXY
TQ88GufXOCBONxTTKcz/JEV/nDSx3iw09SWqBeUo/z+xWMfAO/XSqN37362J4B6d
gwfnSQZY2cS9rOZzNLmI88KTeVlzquRtGniVvnTvZKhPfO2QDb6ITKH3U9siwQh6
ysu4Mzv+yJQ8OK6lESB8P6665H0H4sKKtn+YwpxLNuRloHydgIDv1UZECNzrjWIT
GEgZnjiT3GRkSz2F181oIHYP2ksBAEWayHdWWIgs2dQhzg549EzsU/WmDs3WlV6H
LrRTm2kD5Y/NUw3oSyivyNzojuY3k/3H8Prlo+EpwMVQdx4xAPFF4I1dE7QNdE92
2fHzNc8GpDcOtBzkxjNNkg5Rzu/wvd+tQPXJvzmo5gv4cDp4IzgXJ5FzCY4nYP2x
W1NNJUY2Xkb4y6OG0D7IpmhUhpfP5m6Lj9HCiuaJOUirYbwAT5uq8uqedlrz382N
wtmY9nmBpBqffIKSl31AEHxzpO7xPJbVLsBXBCUUTS3Nck5wyUBO2ewhjQDkR45P
FCQIA3r4j9s3rLf1UOTfggqLqbwA+w9WoIhIY+Khy7VOzBhOyn6ClV93vOgm7qrk
cCfe5Vrt38jmTDeT2v3IOY/mIs5G9UsygQmy6uQcoBmGMf/a0aeNF2aNUd1axxiB
1XFK6b5Sc+W4iggZLbDbvjK4tvTCcKGgYWWdksZJXZd8KUYhxqgD2UxhLjJTnR8N
3mRwWhvceStp6UKlpkVrUBiJmQ+f6/L6rAqHKs6mQLPoUOpf7cktjczqqvwRn2li
y/X2sqjpn1/m+S5K/XhxCO3UTgRWn1hshlDn0RgqEhb8OIhB6Vhfx2qZ0mgbulxH
hUQcGl2gLcv8tBtWtsjK2ssMDQrP43yJvKm+MXJKxQ8hHqycL2yKCGo5jmpD/R5X
ulGa8wPYT462fetiIjEOaIQd760/QRS82mHIFUWDj61A4A5v/NYRWPNOCuAaZZXZ
0Y+gMNLBOcLWLAlrd6vsTYFWedZv5u9VOBeaPJjrdM1O1TSEhUvC8UW/korAEen2
XEv1rymAefKGFmbneY9Zs0QEfsHYcJwYiEoEf3fM6JhzI3KSiMc/Ktv4ZyNBEXf3
k9DHkcRdwGe1XKURrSnCkw+EIfltSOJDJhOYAt98UolCWYe3cOzJqYSsO7H45VXh
bsEsKCoIdW4kG7Q44x37FHhjQtIGwmvl6Wa7dLt2Vp3LIGsPrxfq9bapqh5FP5H+
kp0iQ0sMWLFPAItdix15ESQhe+AQm54j5HZLaRwTKxZ1i24grszulDDjiXALVtWZ
1ZdcZpyiVnMq0RHDmfoIfdWpOUszf5Gb3ZAoTx1kfVmti/esx+Xuu6uW2sM0HeYQ
en5qHhS/9UQKqozNEaDaV3Sif16LlmZLNw7F6YhP85nPINGMOdIY6GvlE0MjUu2U
k9qTMM9B/cFsvWeKt+FZu0bVoXSnjGJ2EWTjhScdAbo7c9swCeljdqUvHi98S3fm
GaUcwp24ky2qXjjZbS87qBF7w5MOevZClFJx0H+akiUaa8cx4HqxBNszMzdVkzKg
J9prMiUs1dUeiR++L5s244dwmQ1Vv2uEc0ZM+s+PVpSs3dKyLjPnrCSpYCsFU5w7
KEAbGZ3WDD4weS37PD0ef3Jvy37VLpKmUW/dhkYq4bD9NaANf4KNj3qi8tokDQvA
H60oGr3IFgRzkSt2qtjSUApq/I+JGP7k4C5M/YUlZGjpuyZW4agkkB8eV5li9HwY
q9gKLQ9geeHnPvltcb76Q9vT9XLlofXAlwlr/nOxep35eeExnRUjqHz/dxW8j2QR
epnGvGndmcrn+8BmWq/1CvMNqGycXfkB80lyAm/8sJJyUUZAUe498/RQpqG4jqYK
x9ZQz1epiYg9NPfr4yhiKBO4MraVMTKghgf3lFKOgMn25rCWiDw4Sq5mOZQmHDdX
bieTVVPLh5gQkJH3DEpu/iYCPXGe5X89SW1MGG3r4fzoZeZm8LAvDqy9shkp1db6
tVLYn/UlozEkNzHfGC7c2hOp5m99Wsdey9Thv2UmY/ndPv6FV0GwTdgixuNCc9tM
Y7VMw5kv4gfZp91ocCewpLngef8BVytOyEhdtS2ZOPcMka17MIPC27RYDKzbfPv4
U22eO1LLilkiKbdxHUEA6Sz8aPVJG8m0SV1OzreTV15WAvD03NYVuQtWU1Hb4RAg
zhSvu8KKIBx2a6Cot3koJwMGCCDPUuJCkLRo/7Tid6UDTK53QY9M/u2J5D/JxDz4
gE20By4Qtte7WwAFghK8X504e3+syak5ZCmvsF5u/ghH2fT/ub71oU9xw7hA6azJ
2+S1n+3KgjmkAxpIcSQi9s34CNVap393WNQ8yKDVRxHnnPcYfeLpTY5TkCJwv3dQ
b1AF8DqtTvBEF2yaNIn0vgYPR6/5Jr7/HDLawCRCvPa3lYBGUXZ8gO+/h6WQucq8
P8PyAVZhIK6RmK2cG4fsht0NL9PxF9EHxqWhG7STwxXuxY6WcSh+9mMB91mDEdHB
YO3DfxpNww5WSboEnywzqAeo6dk57+dQ9vZdNPuY0r21G8sXdgGScLA3dnHpQM4E
5HjLQh9JZy4f4ZyqMLB3K0jAX8cuIqDaxy57oxMKDMLj4K3li+/Uo9PR9xLInj/i
V4q4Ub7sJffwOnJ1eL1wRAh9hbgTUYxVDNeNyHnPNhlOEQkGivQuLuNYe3AUP11+
vWYS+X9rLEXYNt3vQWOYjiCTJm2eGB2BbkqT3UckKmGmWpvt4QI9HMJ4vQYazPfX
003wHkyIssTLwlL/NPuol6FoU3isV4WM1vmUuGT8ImBFH49Qh8sKu9WuSFQH/HzR
oJJzODppIL8o72dxscbUBrh61tlH1CENmtoUzcpXuQKvrFaGEDVD415rDm23IfGr
CU3i/I7VSpHytqUZloWpQ1Zu2fRwwQneDRHubMXBeNIOVLmYYx5cskHu//Z0w5Uu
82viYImV500gjTNlqRIutnajBjuos6hdvKuxuzon1S/DZvpqcmaqsCBz5lnhh5SR
YJ8dX+v6d6zE19vrGdZe3E00Ibn32b92BkW8Lf3p7+I1sir3FV56XUcRIaoesDji
OSVC32Lh7lXqKE9fMl0TTlx/o0CL9bW5bErEnCzkAuMNkcfwyFg35wWWBUexmi0H
stY75zc/DYjIpur0c1X1yl9WFxpir02WHInqaLfSYTrWL8F1VoGkUhELsF9ITpTi
4g4nS7LCqb6OF7MqBwDuKNvDEiIbXVbChKjxOJoGoQbbrmDltKRJ1S4afkczlxBa
qodaR+lPFeszc329fnU9+y1gMDQdEt8WUnGV/JqLUO/Of5I1fkBa/qMxv0CZp1DY
tbg+U05QgDX+v6d1YmDezB83veEI6EfrHRTmLOGufUnr6fHCbzHW4hi6HwIa3lI8
iNhTUgQQN7T+pIbPEY3uVJpfUmgLINMT/XYz83XGApFWhmhOSBaB6ZKGklkNJhj2
uG8C6f1mNdWoye3LvEtsxtwHG9BLd4qXPRvqkQXdSa8Lu5Pw87GIbtZq7CkbQs+d
cHdECvFmXpgEO3ySFu9DIBp7PuKkxiRJUaO+cM+30IDLoo9niVOKZbVzsJ9CJdDp
tvA3cA+bsYE97Rs5zl43lwpb0GmoWUtOmJl3eQtRI/zG/vdT+um2Lz14guX/zWLQ
dJ/zou6VbkZjuZjlskC/cyd8X9tR0r0DY4Ra2y+nl32eljIqtABEg91HVM6C8uBv
dP0rmA6IS1lWjgsbswjZX2nU3OvY5ZJ98tq7RaRcKLhM2uVddjMbCtPgDxvWKZMh
ZPF/nQU0heerQzRkdAQkm32K6+tPn1hdXPdqQ92ejO1DLWlmRB/w1CoiAcaSUxyt
v13UV1Ik5ybgOMXHZ04WDl/ElRZG399T5ajPL+bj+YtPUurhFB979x4mMuDqcdIL
CadIBJ22Mcxk+PE2lP6xau5w4//2uUEXW+pxXTgKJ3pnVULLdYG1SfoGvUJrbcYB
27NuzFIDqJCs9lmvXOEMZecBcG3feN9QJWOqMXx3cRK/y3f7oj59O28KBBRbxpUd
/2UpjPnnOgbTVdJEu5Pi2veTSoOXJnulpQuo2uel8P0TQBBoOhOWF9K0zVjXnih7
p7jbywOWEMjS625N+WnQnaWggKRj3zE9UH6/66UpDjINgsSoL8wbNUUBzGDZI4Qf
o0kEc8tSdrXYwy8dlJ2d1KitG7jpRd2qId6Jxy2Mg2yFJKrbMeNb9Sp0LDAAVTvp
FQzGk8rHo/YLWYFuTWCmwFPui3GA+WPtl7aDM3FGdsynauCWcAXFdMZz9ZahgFY5
BGl94giHasv97TJe6sksXyUQH/3WIOkMm6apQeM8jDznn8TloGeD4dlG69L8uwKI
PSxkN/aEViV2rj7VUdZpY/CTAK+xnyVPKIxhoHWNO8fcEbzV0xHILrjJIAk3ugSx
w7JukrBaawpExgn79LR/CyGYKBdzNez+g7KCO5eRvQ3bbVTTYkPY3OPg5bTCfRFw
QyteYvF4M5lEnCV7L5DYLJ9+EFitDteJHmsR1sbxwS1tlmtRkYW/U1ag+tA+y5lJ
ZgSi8Ed/Cx9BzMo9CZzvXh/GPPaAysdUxCUKW4lKEj3WSFD4pUve+y4bv89xoE4Y
pJAEaiuF1eluVQJePb1XkVVYJ1NEssQdQythHA6Kl2r1rAeN8V53/kiaXuAdEx0T
Yw0XIjPus8FJ79rQ+ayIkfvodxyVfx8AUU6bjRZk/Pd94NwrG2m5nTORqoClqngj
YNH2m3Ss+8dwU/S1CphHjkng18+XS92G/rOx67fTwUr9lIllrJKzWYGC4mgIP519
SfsIj2OLvBo+Pg6yAvqA8v7YWsK/ikdb1Na5QQnOTJanxmBO/O7pVcIjleC2xpkH
7lhvub2eLVj7vPeUDpMLFQgykquSv5J5V5T0+EbiYHRcYfGfHpQiHB+jMAwtPYQZ
c4LygTZGZ1OvLYp6QbyY4dPOIL/9IilHhwsjb9X0BL5vn7Zizr6eBPyd/J6ML/A5
VVnZ5e3BLo0PsGhAeF3b8pWyAeV9bPpzCdbKNiFwvywE1saTpJ2plvAiwBuYdQeV
e015ZswYM2MJYQiPc9u7rdz2Oap+Upw+7nt3a+UMczLopzP1ukZe6J3j4crDxFJK
PVGnu1LPf9PFLh7I4TNvuYgd5SmnLAf6HIaMxPWC2OR/rTK62v8Bh9MO5x2u/UtN
jS8v5Kum+AYsJEAtXVN1kgpU5NJt3au6dA4j3AyZ831OaV6WIlcS9k08C4Z6ueEv
nE76bhoxYShVweuZOGx7bfQD3WEJLCc3hjA8dCoCU9iYuOVLPz3844o3J1+idymK
3qnxdUXz5nyHPZiZ95LQkgo8kjgtgMmuKK+K10t6kMPdnTRKv5F0PeKPLeqB1kUF
hECu/gmAznPNHVa+fOs2VhQvwSDYj13hzsm1qcc6HK2NQPfKASmHMj+F5p04btHh
B+Kv+IlU+CkaWTZ+3inXA/3mJA5YU2HEK1H2FMfpcr/eCw5AZBuGUGmab+6sBsKl
zFeJrIMKOR2HfHVA5+K5pT1OG47bMDRzU0tOL/WMfXLxzB1s2LjBA/xggqPTiyFs
hMtydLlO6WIVo32RZdGQJGxVMqvD8xmeAFBgOB7MeioM/CRhf2eb2AjXvpSVokV/
oCFty6nttTw6vtxoRxKD87hVDNm02+jRw5EcQ+bLkiyVRcZQ0+7RiAYjNyy2spb3
tAfkVYUDfT1fPzH/ddlmosQIuc1Uy8iCSA7W6tWK7/rnybXHhoPVwdIE3jYKYK7l
ez19493y5OOFFuY7f8PoDDaou56ZLwUmFPeOCpO1Eqmmh6HWpshijGW+v+ORAtFg
2y9oLWoc9+6jfDB71qalABjjdwmMW+mTKWvp7xmxCBo9ZCxhGPbVZv0CieftZh76
tUGOiCW2RmaYnQMg56V7gaSjWB5YPoVME0PGx8DQm660jUyAVpr/NKMBTKisSjl9
W+9kMCEmORzQQTxbU8MSHTAxYtB01AH8KIv2tfxdzms77ZwX9syzmh/rWrZqyfA9
zz/eXMrcjwArM1DYPB8lAWOm1lOgv6QjaCBiuvImEwTWE/7xmuRWBASpzlew7bYe
ZM5+eXu1pZ92ZUiFiWrK3ygG79yd4colxkEI7pglFCOVdAzg8MnhAuPQO3f2N43Z
nV2t2L9ySVPr2rE0ob9r7uQEcLJgmFWFX5lzB51Uovlg8nN+puSptX+Al9R3M0EJ
F8+9+B1ltpnzokhmFQphm6HTterKbeQfwFl+8eKkkuSESp9jpAS08dOxJ3ieu4TV
1KmIuk4wMP5O2UP0MbA1THCP70mihIoRkOvDn/UT+EH8w7ztCSATlwzidI9Stt/P
iALprnpJYF9x0zggeFbJxNHfGBwF8M2oIh1htDvMHwkVPfIrpLAUPnLykG2beEIP
A0rhoL0vS7EDBCdA1UJA4BcLZ2ZN0Px2F5ZWKR0FN81nE3N6qbDRtR8VWDEPTdq5
1sm2XszIBRXPyBdNeDrbVjUBcWpqn/BEE/nPGfQsoCC2kdrplSUfr1EEFpbQkJOu
PvpFwsqGnB72+jCV6y/9FirwCb6+KJopaPUwigcfDV/1Jz+WdgFl9t8i/HnsuYAJ
SgXrXixpksSyJKbKk6iZgNlHxxJbabF4Uw4Kiu+ovbMWOqgBHi/+N3I3OdhLZRVo
VGBCqEfoVHc3J//hlmY4jX5MyqKKJOr+BbY+KNsPB195bygKt31063CjK5bGeube
W49nfWp58yKsdiVm3rmfYHCecviYw+ww8Axrq8WS7sWdc7mOlTpx0OL+MbnI+uBO
xU7wiEAqQ04nvZJqGIM5XFJItTKLrlUkf7CHgKwU1460Cm5kfs2yPjd141ss53YX
HeDQUiKjAU/L36aJGoz63F9DiTjt+aQJlXVij/wPAaxah3aECG2OAZyiqm9Ijn9R
2+DldfFNMngF9UnKlSF1RsmC4sOtcifi8CccyB+7RJHBW8Bn2ObbPfFAjWijlyHG
wYYhabafhc7siQP1hDVYmkbcKXGhTOn0ASho0d0oGvxY1oiQEbwnhSHt8BDdHVId
v5P5oRgFBWTVcUnje7rjLyVjGC7W2qFtZkeZLh2jphPYtaipf/bHRNRMBPp0XKLO
d+AX4O5cH+8CaVTaKZETVyFq+zheSKOzpWS/26ewy9Y5rySvt+sUqu83r+t7IDfC
f8+hWVAR9IHhi7SKyzKXiiSlD+CfhyposEHnANRdgmIOpKTPPh1FVtdJUrVtIc1V
cOKJJH/96TRYC6Xf54hWlSzvZe3uuS3gHgvvD9ilRrJl7UJJADOZujRztNroJFYX
QVrQRcQA2e2vndgqSSQWVCBXDQUZMs8PDrZW7QeMeQ9gpnCF3LKqF8kC7Awqymex
f4ZzQRKY13irxfTpuGQbCyPHQ4PbIGr8EA8feGL4E68Bc4kds8dSH+LyCpvmrp0M
1G59nwPOQ+fPhTaxVLMR9A/HRTgKK7FjIzhFCrC6OtecbHTN7kfw+RuvZUZZFptp
hB0bbVLG308AW/Wc2fZmXKAoBed1lTiECobwS+23fpFgVV0tbfDB9EHfqy4v0YYU
qhJLpSGM1XYIN/vuZxVm5mRU9pm5umN6B+SqUL3VkhmuU4ry/j66dph+KzuDxdar
kUGihmOGipnovOZWT3Hqadg2qFno0/urWQW0zJq+e+LVZBTiisabHxqf9S+P4xgT
aG7yDXCDe0T0L/EQ4obAwSS1awypN/P0aynj6esmH0Uqdblol7geoMG/dGv9KQ4A
bq2nhBFci38WhT/CCCc8arsrngqSZ23W+mEaQ9ruGYApjaagkJbCIt+89GsNF6KH
c0k+Azo8i5lQ5JBlVlNDVcZh3ilty0ZV+7343nUVXtA08571CS9MMjUvDNskeCcN
6EFoWeLwFL+fyNGWRUOQsXiMGoRc4DNH5QPVgW6GkXeGa3KZPYPBehHPbHxhRLTY
nFbvvSfcufgfczLnRCcK/7GQj9RZkHJAL9V3tEFRWOMPqJwVmpgs4MK1KoLQdjDp
YpIlZOF6w6RJFQuTVouQiGVxuxyAqgOp856bmrcUWUY29oSFpkuPSWYL7FdC3Edw
4A0TYkUWn7AVbqtw9xRyzAcpLMTHIpbfFneSuCX6YhLRRYSCdWSTR6b/p612YcpQ
f6i1Eq7qvzgYrKgAtLpty/GF8ut+khee0VyvBYJFcpnMh3YhmDw2324veBHlgwIQ
KmkK538rJ1UxPO9aS/tgU2B4rtyBmFAeZBg9Nf3VoEXoAwIt39HtGPYUmZ5PqDAL
nBgShoobz3ADyIf+tHNkBBJFFMLYoom9qkJivPKi73axqRyHczZAB5pRrFohfXmC
KLs14Vrb6XyxGigyZZCP4/1Rl51ejgBbuG6kKcMeakFgk4Rx/kxj8s2v8/itZjiQ
INIgDneT3+181KASb9NKzlfVNnytZDOQjisC6kU5R1pWORIWfNSgbYW+PlmCugs6
UO/qXHWrcMqbyIdWJujnQT70yKthG2PyUN2fnXzuOUHUPRdGkMaycii6LmWUtriH
aRhs+JGV/g4NKT9GfEpKBtcMl0n7Vm9plfcraRyY6bHvwz0CIqoObcM1KDnfD6gZ
6sRwOWYS5H+ZfYJa3ZCaTfi6IMNQAZ1GMzB5JtNCtrnwAX2Sp4oJzadmz3Yn9puo
L2WzARlZb+txcouHigtKwCvbuNAPsLPafIGi/62vscSL39/Zo2PKnr2oc6AnSB+s
cwenf75vjJWYwJqbNrutsXgsqVZLOoqwQ1/DKrJQZmP2gUvPDvTVy1vMp9j0Z4pj
byu6Ia4XMLlOdpZZPPc7+KyhvFkvlcD3nOTDS/76oQNiaLpl7QDKkaM32Mes3r54
Tv1ugpKMDDvEGnQD2ZDIli6MgxxkxczplXwBQ5fhvaJ0kXM2bv0LRRhotYwXhLAj
QQYUzHhrB82NcKdjT2mGLi6kkOiH0ynhL+UW0I4VfhEao2W16oh/t8MMdpmZFhe5
2rsmFjEvM0gC2Jy7EKGlHebpL+T8KnGdnhylQ8jx36zkQdF0eDesKUf9Nl4ZB3uk
d7YCkCTUbI6r9lOqpi8CXt4+aSNqqOW3mcylzNFjF1kqQIWlfkbgDjongdPXeiI+
p/ikt5U5DFL4xCE1FRbrJnU92IvJVZuY4M1ErQJzR8r8q2KCVdKiRUxFpyi3H7Oh
j110JPZgbaJiK7sElmk/baw4Ieoxvzw7+Oc1Ai+CogtGTKDl8GzT5KCb+Nyj7pXO
fIyDgXEJboAijG6blVkRQHTn14MYYjau7AfyGl2eb0/HtkhPQLYziz7PNKsqF0yK
wUnwA9QPOy5HnGgzF3IkEuBgXAd5w/vy5nbnbnZF8CSh3Mj0dfRxzaZBWJ/LPxX/
mQWOw4upllJ/ToLkLyVFiuJGV5KXEp2YY5EOePP6xbdS6sSldxHIxT0YY/CzgPyO
4Ruu5GGf0gZKYSUFZ9fm3W7J371owgluICSu47NXQoxsDVVJ2UBL2x+QWRMASDwa
XZhFrDmjYI+eAO6w7V75uEGjTpl+pCbNp+KGjUxQ7Qp74pHrQukXbkCr8piEQX55
PcjByqzrxqvzxuyepza0HMr6GdaDVdVO0y/e4fpSIeCb8hQQUrcbQGV7OhPL6IEU
8T07J108x4ozgYFS17iIkFCyXIlpflcwRz++oQRBySsoy2xrX0JZIwmtm7klKvRX
ugIDH1wIzVY9VpUrb/EdVncbDLdiLMRyVe+0QoRC2lWzp9InjX6cgiQxJV5roqQR
/6G8fznROTqMshXhF1oy6If7cs58rFoIVAbsGngw7+AThc5dTrRHzqJzSzZ4X8Hy
w2H8pchAkQgKi7oOWlUcH3PNNiHkZ8yAOxrzcGl8mNk6a3RkfXSSNTfAd+KqrvUS
nN6yZfo328K/YVgDWVxX4f858sAA38XHq4vqgDgGlvF3rGs4PnsJ1IgXZ5T/PBMP
0PgUdDXV1qB0MvYNSNyPqNk6bGRweElpyIPCXT2lQvPGprc+K9P715kd+zoRTVOE
U6gN++jycoUo9QMoXOEG+NZj07w6cb3ROeq4GQ/k220BCQM91B8UoCooeMKA3Y2+
feM/hywBD9cFxQuIg3xDrVvitS1yCcnNMg/JFX2e5chwAL/MS3VZmWpFdgBFC9QO
c16JXIrzIwuMILWH36visRINYh6N6YKBjLuWhbOnff7s5IG9nRc/ACanSd2B41ox
nxUK6+grGWk8FiOxMjJyncvkuaFKTohMq/Y4y2LvoIsqDr3x8KTmLMBgBhmxJDbH
qR/WIaKLa4jeT+YFvXdDkYp9PgCUQEt91SgSEWyA9kkMHzJxR/lwdNeTCJT19ii5
oFPzNYGGBb3z4tGCbEYhQPRv3oFST5FXLr3j9rd7YzNeYdWS2yKPeNFbONF0f8zD
WeYX0bO5PN2Pj1GKzGWF1DbKOlgMckb8O4SC4U9antss3/hgQiF5xzgkEvVxBXyd
DOWZhrgBQLmdcIOUWsxPfHGgjh+rWM25UPbgsxciM8umOVKUtmT2T7G7wqyjL3AA
BGjUQRycnwvf1XqtqA8OJ2VikBSLx5iT5MR0jTtP2czd9NFpI0+Qn7wgG51GRsRJ
sdj0A7nD0ijjtUTWHuH9ejAKhp1TkIkic8q/scPVe37ZGzU+Q3Za2TAeECLPS0Uy
IyxEOLhP1EJvZ4qvn2mVJEgNuOzCXNTBKy9vrOZyhyI53PDZEHcKhs3kDD4fnZrp
t2f9TOHjVg1Jm02OSFBuWeBV9s1GTMBMylHSp/HieXFA0WiSiKMHKmhSmPcNswnk
v2RqtY9FQ3p8NyyMKbYIZtjLpVEqCh/sIeHaE5dvd1xAplfT2b2NvhSDjmiEXQST
lliK+ddRzmiGILerJCEafRbzontEUVGxmkjsup4V5c9yRRNhmooAwBkridKqtTeO
p0+kSpyepOPDNKmQq556p4XK00fdTY9Dbs888+x6YtwDCc2n0nDZAu3LOK/4h23b
XLxylyqBHxdub4nX4ZHpoIZ+evWUTkjQ+/E/LKu5tb+lRaK8+ZsLn1ZXVgthRGL/
TG1gTw6J4D6FDHo92/e/DqTFwB+pwZ39VfcGOC430ASJvyqJ4lwtlbJkbN6eWN4S
JQEdYc+EmAT2mRxkUnP6tRrlDo0Jb1l/Tx4NrkDYkvwRgbs4SUijGbTklOlBvNH/
le5eC90qUN1X09UVTp7IhEG1atzHMwLqagexKpygykKpkOA98pCd2unNDHNEeiZU
+R6znqFQfEWTofbAcb3ZHZdaedCs6TH+wKM0//0bVE2sgGh3ITXfubVbDu9nGwV/
/hH4j2ineGcIEok5hifxFAGseXXbWyriKZR5WC+K4iwqYGBc1Gz4hu9gfPoIImUY
rBto6G4bI22I3N5TgaRINDISUwc7YEffSKXz8UP3fz8zwqAmv3dB+dJcAaHa5TUS
ELytj5xHO8do6+TF4euA38FWYhzgH2L2rRrDH3GCeQB7CQlaMNdGxQ04kC4/GBeC
FvFGyNPzcOLqGnskDJHrMtEogzE53Vu7vJvUOVeas7bZGS3spXFcidMm/UCYUkf5
uDl/yENvn2qxwVPV43Lo/plyNUMx1HJUlosvshJR9S5OzrChU7rBcO2++9kwLhZw
mbbLJlxv7wQNDsH6raQ+Lu4syYPI6nqfDtvf2orEUrcFNxRroIEvHMg8KqrP4Usx
RcxFWsPsmtKZSvz1/nYdAh/OprqNzcQSPP43Ccx2Sc7lCk9cHrN6zeuHtw+KjOBM
6WneIUcEYhWwIYwZJSnlwYhdUZ++XhH4t1gx+D4Zec290+Y0ITLaVrJHC2YkVYAR
e5VVkbKXHMFJ5psDm/xmnHtNP0iP3qFrN69wR418I6LTwGnUXZuxT7zqzFuzWUfB
F46BC/wvWoZHaxyxLo6K1CrtlxZdfdy22U3gUqNLCs+0UT5pvYp0e3nBMCrXyHT9
mbaBFHB2hdvi4K5jkqn7Im6Arx10kJE5JlQvE4D6YekgC0s15TgCSOwO43WVGWFd
S2c5z1qAzGtS9IiWI0Ngh3qB5NTRntSRkY7ho0gkgHs00+ZCq4tbr/8N/x3mWl3b
5bkwPPbFnmpsbod5oUJNNZ/yVf3Mmti9CGDqd8DmFrUGwWm9FurYh8ZJffObLOfm
Sd1cLVZGGvDzPSHSc1YnpCtwlb/w582voPRUDnOFBZSbhlYqX6Sc0ugO9TXJzRis
zAymkFHb/iYQqxWSS7X7sV/0gnW93bqKWX2UQ64AEiXpCgpKY6VQNUx2f9PbVLYN
RGwbBsBRO0O743aIxnZC4ocFuzTLrkxAoCDIPRM5xnex73KxZKwXcuaTEJQyoTAk
w/VB+I/t3jQp3NPSXM33GnRD8GuZF4Q7FvhAOj2xUF4OePMGD6XYd4DDTQcMtjkT
VMGq9hravFGK/vpbTt+C92quELApvQfB1X78eXoHUPEjSAJb7CyYOMtaHYB7ABw9
TrSVQtG6eMUHnJdNGEE8+DGbmV+DH7WKvXptkCsyGU1QRnY8FYWQwJ9S8InfVpSs
zZJW04OJbO1zk4qy2tpjj+yE//GhAeX4sLcsBDNkGnlN0yiDMnvg/5YjufVvTbRN
6/fAXw5KbUeRcoUDyIUzV2UcFdf7IxZ6t/3Lyd1aLJg23OUXHd67Chc1Z2ROIQk3
410w1upYVsseWWmKIqm1FczTjYmt8lrolShxGR5uQHzYBgVYfGY4n9nQEOYNd3fi
+tzNZL4e8v36OoGtGGsOFw97MDc+Tm800/OFwP3eZxQDRKTb/ni9AlqXwvpqf2vn
0/P36SEp07B3ER9hLJy5pirVJ/1Zv1m2zdN/6a6KEhqc9RxIzCWMxCZ6764PC48a
Ggo29gZE3EVhYak9D0xkFTuotmJmyggCkZIPj6B4AzVH6S/5zXGKh4HJ/l9/2p6v
vWsFp2FUHdX62EjcmfZpoh6ooWstCkiHeJw6ljDLEyFZ6Dbix8Xt5XtMacnkJ8i/
LQBdTjdhgV0sj3ngFjv0u1LMzsu2NJhkglx7nXYpio8wlX2cb74mo4hKTLd6IxVO
Z5eOS90wR6SeFYWfMiBwi2APcUI/TJsBvLm9NNzEfhzRZn5iXyCxp5ab9H6Fgv+Y
b1wGi1fDWuTTLMfQVKu9COU9m4wjnxOiNTpwl2YW+2g3+uB11mz7OLd18aMaYQzR
WvowTifI2EOtyo9eUzP1ptdfDH+wz8YbdfmAr6iOtpSJw7ncVhL2pJhbRMUGk4cq
/AeG1HiWlTxlESXGzzDRT4pF288s/NlyegjjjqO5oTOEkG/HBvPFk+NXXAYczY7B
fOm0O3eJl54O6Zru2iD1UqO33l1l/JsVJj5RCHLeHznC50CYCFvTpgYmNG0aTuo7
kK1eEFXqdbKuEGceMpKf1cKZF3cqUJ5Z7RkzhVASjF1Ie0IGlix0gV/7Yq72iJt5
XrwiTzLsKdXxGMkQQr67uz78SATEd9DuKgOYAZ9kAC0mNFlHvGguu5deaU1fVaf0
zgAMy4ZPXoTWI/TJYvSfNAgodpHtfvnn2OsQUnPity2aB9Ny8yWBwiN9WgOXOzbI
Ud6MDyPW+ArMHcTREzOOXQM5L0hUaIj2hEOTFW47NBKQlRA6SoJ42xyoTRxghg8R
kpqHx8PADkAAnFRL+eSnTFUvlaDleoM580Eoqt5NEdR2t6XK9VJ3dpXPJNq/NctA
Td/eRUbZCtTdAXarrqCn3rzjlhjdqsZBIM2EF5B7ftrC9wNXedoIf9lczqS+7Ykc
c/Tz3gyPjz+bhL4heSWSl8iw5NUk6sF6sGb8UN+MCyEDFTFz4pOCjQAbH5/FMM6E
j9WP3UPngjwNwIs2mSOmuT+AMr6sV4srBaT9GZ14T8zVSZ7HZZHUK1Ivrkw8EH3c
s1X/u0LMe6l4PVHim9Z14B9sua5cphgZPqzuHYZ4eena+i5eAh92nnmkQvStjtdM
XZUKcISRxgybHO7oocCvMGxWVvihoDnF92SfrOi0ZlT43TRUglQmCYiqO+4/abvh
US8GLOzgk0BJ4HUx3KkmRGpjgGLJwUmYutGJRapGdNZNYS7eq9e1z7IUD933C5SJ
W9UqQw4Hx+1Hll38b6iS4nMd3Evz/DER9bHDmX4/DKJ6I8BKykESfVRoSju3Sgj+
8789oOdltqLOmTyDxWf/Cf8uIlTxM4DQddP3aMmOaTFBN78YHuExCW979pfKd4Nl
0hBQ7zVWQXs8HTu7cBGcpKTJy6jkxGqfBoW37OGxXqwdyhJLy3XnT3xm7bP+heq7
SdTAhwdq3adIrS1EPkuTQKHvtZGx/9PsZUu1+SUxHtSKYtbRh1iqcgWe7RCCibS2
/b71iZSxOFHhWRzRAcccUSjkcUeVzLnR3DWh1ETHAmG3CAiiQdMkSt9wWJJnHEUt
R8zanLFC+t9qu5DLvaUmKBOUSEk3ZWXvVgXdsmM6cyV2hDLM2O0V9eoLiINH6l1I
vnyq++cVLQCrkoWBCrq7BZQq4ztg48fWn8q3WgfnhDeOcibZ788tEgkz9QMupFBu
CYijGQYvvZb3bXjGmae4dR7ayR8tId1B2xYzRUbgIeuVA0dOO5PSBeJAclwT8xor
rprzWjiMteSEcWvmrFyr+5lldVHTO2tDKTtnXvx4PW0ffFXxqxPMVtKQCcakBL7y
K9MnqoCbudSlLqCOQ05AnQ9BNJpz32CbfI/r01uaGVQKzRoBlK50SzoKCn794+9c
rVmq/LwLoPpTUZpf6LbBB92rd26aeHuD5I16Cx6NBEqa7RJyxRqumd/bHinG4Oz2
FJKJOp3LMIfAsu2M8vyBrQtUE+7j7ai3UV/wzoF0kusOzwfXZ/xxJ2+aqQQDxBPV
jVjGCO2WL87b4a0eKid1yqC71qFpcDBhBEFQMUC48/JLpxhCTDwW/R1s1blZ3j/M
JhyF5NMWmtzbiK4C0u3uJC8rh3pn668L9p1AUti524UGP28ZcSy+3nv9QhlWPYhS
DkGdov5QodJ/4XxkkCm58onFE3rNHsWX2pf89gOHhOGVgqWvKEep/NSnkoUq20UI
KEexTcofUanEHkZMoheW9t4gYoU6Y7AS4x+xtYEQ6wUlLaboW4aYqnx7p5U9XwcS
o7x/TPq1E+RrxjCHmsrt/f2QlsdSXwSu0VWDTUCwXMLUtjhm4YdBjnHq6lZWgF7/
xjUSGrDmf/1NZz16DqPjWENPIz6zDPKGjrEDXfC1Plh9A91VpiIRTL4tfOc3ct9r
QXUCVvW1Qq/sieQZZmYLQGzG2LYEvBUzF2pxfN+pJnL93qBDFrRPccN7iTw2JaOw
3s4LEwHWHEBWLa+KQ3SfmTtcJ998fjKlaykhkFQSAPO9MDVsmlfss3X+LnUi8VEq
AyBVU6n4nI10xjJ+ayfOfH0GV80atf1TQRBnQmgQMlVlBcgVn4tEGOriwPwa/Z9q
5sm7VUa8IuHrkojO76qHsTnGVD5nIqJ5UNmGY7IqW/kg2M2sV0MM+Kf/E6BYt6vG
94W28zOAfojfm+o4dj3enHdKLLbQy5kMt0dvezaVGTsuJehpi4pWdrMQqNycSEmR
Rj2W2H15ghysSGvmj8xIEsk4FLXg4tfohxiE2cLrRf2SMf2K4/cc8LuGOqrrPvJQ
DuRbJ/LPI8y5xSVffOY4iQDbBo2WYnTEudlypsfBJXbZaRKp6NQMRbW3cGxo1Ex7
7NYcyXkllZEinlOBE1NWxkwhiW2FK0O0IE3K3xX45cYdVddca0iitFZwy2/L7BIh
6CTUBewbEMyBGVMkPYrU4AtvuH+daO1laKKPOXepck3ALLuRY54CgTcNjjhOdez5
b8x4B7ybtOjCSGh/G/eDrW/ogmoLceocdBXQHdoAOMRIS9OIFk0FFvzuatsoGxE+
FWPo5qM+glthUjJuaXjHtJR+hQu1LBYwqIMXhmEt05JW6Rfp8wkofYKC7Y8/cIpW
P1XU+DxlrC9XFDhy4mOdzxF/09A+VO7tRFl+dfv6g/9nKwiieexiWpXmBQOeon6V
bWFNnCxT6dDRenSRubnuQpuic935w7QRK9dBUeXyYTOUhayF55xa/AEWnJ1BIEGW
+xmfyK7RL7RgrUpb/h9zTWf80zib47YFs9XDDa6M7upGZJCy2Fu7gmla91x0RoEX
9O5CB/HaqOL35dlcNgCJTdO4Q1rSqRLH9tz6gY5H5w64fXY1vptcJ4wx9/BvpW75
2ZJsxAdR5UDldhFQCYGw7Wo+s86h29/iT7Ah9RnHdjIhfTP6DoER4uHwLqWumZSl
1F7wIB6/MGJeHOkfYivEC4X0TcCrUAW2R781yxTCTPCInOkF1gVs6YosJLae6afR
w/pl3gMZcq1eyeXFIrPaS7fAYxoEDPMXpJs9mxj+kaVoCpp8CzG0srBSBqTaHw6u
G7icGu0wSkUKNvUkIkbFKKOw4OCXhW9v6QlHGA+U11p1dGill4ol9zmMgzM+/P5O
idKqXeWy0+EgkOn5z1N0xyUNrG8wVcIJe/lZwbBqam0QOq7Tt4g4oqKeir1FSdGJ
U50AUH0BW7whwDvwJKMWwOFncIwo3XOlHG9zULSki/DhlKWaCj+RnypdZSDAf5/r
LzYknYDjTNknCarRWSsZkaDqSXMr/wcGrB4sneMzHNfpBPaq9B0k2Xw5riPFTHRo
TDiDAjEJmABruRxd+9diinnG1am/DCzSCBGuHTmrngeSfJz4Ph/UJpcme31OCk4E
iw/+Uh/aSVsgd+g47U40AUX2gguzw3UwEU84quJTRlWi0LrX3fn7lcatrTyiqYDB
QLCtLWCTFEL5855SHEVJdt3Xp9bzsA/a1E+A6dDjYE1cGTqOGD5FMeuSrS9u3j8a
3nugJg6Y7LF7ZZe/+S13sS2hR2x+L+1SYlkB0lnDNafl2Acy4LgjRNmHLzFhrv4v
m+Y3nx/hnJIywt1CPCarlIjAec+qQtfCC5PP5L24HdgMFN7+D3E/xBdd4WVsDkqo
S0tCzUoPUfA2l5dNvswcp5gjG9/XcXuoJAE9TC5mOGTJIyoYDsp+IH4GVnfOQyP0
ia3Cyee9SNrT4PU10zqcLLHwWVnKu6hl6UZqE+wZJZpjcnhuX5oHVIJ9fb21VtWt
6pRfKCI01hd4iHxJFULS1sn1O/Z3U3KsuHFubNLBMx+PxQjuchn1YzvhceCH99ka
0Lkoi2am7Br54XiS7mus7RxfXT8O9ZmsactI+90jPClsxa79H7dzUtKoOZKDng69
4B8bu+laFG/sAd3hIzv/QYt4w5uWP/3juGxyG8tmHlULCfyGFWYcEkcv8UKouZS8
hz6mineF0aUF1RZHRxCvLfJv8j6Jm6ag01w8vKXTif9GKNOFDgjMaHTWPSUCD4Bt
IEoMT+BF8S45rNRrQrKgIIn6ja99mf1f/q1py+OUFnDLluffn+q5FNOba+ay7I/c
8qAAWpy1EnNsXSxwPXAd8RZcVGkkGqpdHwRJ9uQEjkb6X9LeYIxXTA1ygqD3jbhY
fqOXqvJ68Fe5Os3spsp51spi8SjOhkwnnYcitMulz8RQm4XOsYQfdopmKvuuBX4r
LK0gihyoEW9GWuLu/v7wAATYyXP3Gz6z6C/mSMtjX5OHDvAydBdZO/CYljjMU3oA
t2tyYOjDjEYI+w0OL2s+rXjvhkaPfN2ZwR2oWelreAbEEYjnMAZhvTYwq++yo2pk
q4lB9Rx2nF2BJymVeiLGmkD3XvajPSc2meMCqbVpWX7KSTYz7DW6nDoGhLuFE3vc
lM+WVLQ1D/py7I/wl0KO0ppyJLBkBj+i1PGxDhf97DTXz8s7n1LbXKogkUmYn6Ho
f0Wg2WfA+T05pA/MMst88BUL4ymQloSMZs4TZumfUgvij2fesI0uhEycjWKZYrj5
xbW3O313ukaHINOlKJGiFXI1xlfeQR6jU5yRsRs6KN2wJn+qE1F7WWE+aoHL6cY4
ck+Dvps+Md0yHDd5fM2aEdByMsVChUSY8a++1lYRpPhFOVJ/Ph24SxnGb10AEkob
fUe8u//GdtDtgHfxyLa905Dqj4aPfd8QuZD/CYO9joA5IVawOAoimcqyQ+KhiyF4
CLqP+8jG4rtX7tyKoIaQiN1bCaxEyL0ybCcrMSj47sT3PhiMgyV21ddPei7RvkHs
xkDIRZ//u9VqFjxRCHrOzEAzRtrF1zCT8Whg/pWXU9zwrXQQ+yViL77hIUW3qq4y
3cVXoyCNl9eXJojb0VACTLcOh5NyHguYnBJk9PvfS5Xh7j7AN9uuAdg3A3DDBBC2
zjE6qXtxWZc7zQe6j/D3g/YCAN9fvcUvyGYwQ4kE16kRqwE28kMRK+PFkxGXjqZG
e5URL3wBuGtBbKxv75p8VpfKAk0x208z/t8IC2bluNhWcY8a39u9qkn6WGkD9Bw+
1tUCHb2eXyM4IpcCAjXXVdV70BRuinVwuboFEGKBvKCfgp1PFJUv1M+FY1v9sFQX
6UVQGhnVLrqX0FJpMFL22CR/mp2ycz39caYXQmF4pSJ3qta+p/cTfKkKLQgBXxzJ
sVw9K6I+Nw3TKrNl8cWUKTwv3cq0QoPlQmRbDzaiUENWGX3FzakIIcScIEDRvFty
7ctLqTBkHeSyEbhsu54crjeRH4xU0fY0LfDKXQP8qA32clqJg3BB3i7yfgoMw+V0
aoIO1MfWVRmKQXAQh113fBzbzqdqn0bzJSzw9xzAi0beNEIuadh8pfcDoco4GMjQ
fVhcclL7gVkX4p/k25dJ9CCBriW5C2GMoi6xlV6pX9kyvHiviGE/ylg+vDZB+ANQ
hZAiJiaPxoX479Y2h127QuqKe7W1U9JlpYnygNjCZU3Si1z+4Z4gJdQR3zlhBEiC
IsszYGSLnsO7xnvQVBSNDk3AahqwfI+ujn78hHdsSWjkCgYITBIuq7Ci1+2AcXEk
qDr4tzf7UAo45d36rkanakP07CK8hUYdcNwhtQ9+4E5/L8uTx94QqZyeEve2c5wX
EyWSCcFU3402C+7q558NNGk99Bue6/bVgVBVAJYTs7UW60j3SGZpevOwy8N4jZRN
notVhat/1keNJT+h1e42NdppOjDmJgCPhILZdSRYhS8BmBbEGgkBuaZYD2FHHs4W
H21s12LFVJryIywsPfOkW0+UPKaSzcCrIPrze+JdRgGPTn0oTxHzd7UoqEc0ySCr
P9tF0BzdwCUIZWLIJwMybNfVP+Fz5uFJo1UI2EdQNShIPtJlA+8VzPn7qWduFVvx
gQom7+z9WjxPnmepIS7lDfb0OcGKaNppgjbcl+7AnaTrhE2eeALGO3apTwtnUxIz
A/9EBuHoZfZNWDjy6y+PBcIUReXRYEbcJXTe/BfNUZ3wRm0ANTAW9Ktxkye03V0Z
RObou6FG9mrGhkdoZCCcf11vBOHsPwmS7PXC8EqB1z3+yuvnZ1NmqgwH+TFKTrjc
WeJ/RSYTw+ygdAnfl3JXMnt+x3LHC1Cfc2WN7R0fpIa3Y4ECsU/TMZKYzjfjgxOl
9KLSfrXEaL368wwFe2eS7ExtdP4Yof9y0PpVMYK3KVHPzx5QRxlZNerHciMZAGsh
28ikrH8zutB+LlOC+arh6TgyB0lzskUJX/Q9qByexOsS9xUA/ZH5qeTkgYn2mZPX
5K43kyOmaRkMjNyaverazicNyDYJw3kXDaO1uMtBOV5nUX8v3YjXfdjBx0jDAPEi
VkeOj9sMgemh+QZcZnb0LR9jJuschCZb/D8R/LhYLXM7TidhI+N+eNTJ+vPydvYs
H7V6OB6cgVoOO/jhD5nc5WxlXzKPl6mONgrmap5Ps12C0Ol6bnc6mQIcH6gFtpXJ
ZYdF3H4ApJiFd4XoyOyaHsux212b3nxnsrc3vdlfr3xQMn9Zdw9XtwgoAAS388Mv
zB2zqcMkdRkKTeSKA5KNHgYp7ls89bjr2H+y4qisaXcbhEe+iWjmbCXrNUUofUBX
gW/zh6j/ddV7bQhuHzx/6PY6HbZgJc8EMam84WcmCpStoqMy94zsk1MtgO4t9kVs
8e/R9xoFXgxUjQnw8sMAjzyCQtPNeeMbiMGt3g70l1DSvzglMnvj+B4iZjLyiNcH
ziXyrfo4nrY8te2Xnj4Ij+g7nIAmjgo1BgmPUi+HArpf3fx7ZtfnU0nvCoqNsPFQ
8fvsNn0VOR7apJz6lOdF40aIXp0K4VqAU6qW6FXCCS1ckVVG6aj9XCCRrCiiZoWn
IhKS2TCKMXwoWBYSpw9eLJM/0wYI93vJC8ZRjKJSkKFGcx8g1++ZwtLM7oNJ2kwM
4lPwM1RNF9Ee9WnFa8dYExz5L2KOzwLdXQoEvv6Kg9m4M9yz//c+KoETy57/9tk7
7KtvAcrnnRPYL8s3Ur8soVWweDWDl4n467v5pxeddz1YMcw7HHkqNJRTJbZ3Zf2k
uRMt1rpZDPyRiD17VL0OnDJ8mkfQ+BOtuVCwXI4O5ePiv+pabL30WhynhCg+LWb3
y6xZu3W13Omt20f7wscf9SaAOTjb5Cpds+K23j0t227BUTDrv8nY7cZ/AUH836+7
fUIey6o4srhUC0fKOpVo1PwVKU8KBsQqjgwZENZTIy7l/zab9tCsS3ZbPvSJRYFK
bnllCSDMtUlxVkneLEcAHIDy0J4SoEaXZndSrhQYxYVwk2jYZqNWfj2MoUC65Z2O
UpVsuF3MRJvgxRw7bRCShRMsidm3+nx7gT790/om6Mo2rjPpzV3jz3K1F6vxTOHG
a+KnZKK/EJS3WOGqPgXQGsKCNe7d6R5tEnIQ+BqzCnOly+div7JsB81ntRcYGF/I
gIFeenHnCP/Qn9CgWIs2UFuQPTjgGuFdp5pRDFYa9ZrSnq4bYTD5tOju5fhqMyp1
jBGmj5FkX7Z58zjcK8jz8QVqCCntZjCl3d525qfEeSUT85M22yc/2N0K/8o/N7zB
CnQs5N8j8Bj5SLkQzz/jmTDVoXJfdRrovVsjt9WxGX4k9u3B9LmGB+Cines7epWQ
7YDj7bjqoYULe799DrC3Lsj67O060QlGnFFVr7ln0dfFXK1jvWUP2FxyC9dtS3xm
ytmXduiuFzFZcVgcBtzv9NyI0iBmWvnLFiMp64UTfg3PAk413DtawdyJa6bpMzxy
CpBPVaNKlE+X6N7Cq4qLi3TIk/vDm0LwDhL3yjQ1+rxfVfQBzOiyrK1ow3u+gpn4
5vPfwSZ9TOr2tjLmcfUvJWhlxvxXx/XYsamae0vk12isqjPDm210sD5KvFUIg/Af
sw1WMtFwUuzBtCFm2qIS3Ac6zktsLpcrsBOW+G7WRIweLHKN9h0BznhdIFLt58Y6
FyEj7EAZBI89uiIr+oYQ8Y8NgQ7/Qh3ixF8+3vlQ5r1Cqm2eCPZ9Mo0TVUeyJkZw
2Lzv6xm/CL2FDUMbfIo32srKDOIqtnHpJf6VAgDAkEGPx3H1PaOJDq7UYLDpr7cw
Z3SRKzgRv9b2T2Xynw0iSaeclgu3hW/nmWXPsUyUxaEV2/b+ZO5AigJBzEl/Cffb
zV+wggRIVzSzKkCx4y7FJxZmLE/ry0AYXlKEXfhi/clVL3ESdhj3MZyxVcU1Yhu2
mmT20kfryZ8L3HlVTUjpaAG9RnAlBJEJFmoXJmURP/mInPn/Yi3X5EyKV3AkKG29
UVP6ROVxfXNLhU1nx0FDUDVdmQcmGeMvPKQ9tBhx5I+McUkmzswYFrRwh52TkBJB
eA7lHE73VOERk1vc8sJlAazjDPRJo1p5jUeZ3RZASQFPsTzTl1OU0+/34B2VGCGJ
MWIUMSFLVEWgcfyaZ5xkvOdBefacSwtHE8hdCVr2iBlDLRBSl5VxvPm2gYOnw2Yb
1JRNPCyZUljI9MHo+qRUcjbbdWNWNPpTUKZxyCdmVj0t6Qy96FgK8IaNu6Q7e1e2
9A9JeiwpP1CFLNvT1aUnTzAlXh5fG5cK8a6KAbJGmamEp0Hueoyk6SH2TDo18e8x
3vLO9gVPd3wDIi5NBKyEv5x6Fh2ZRG2gIQUYbbeXP7zRLAT0f0H6apX73dxtVpfc
i8i7HuB2o6W0UHmSQoVxcDhakThCEqCx9xhikayoPvT8bABuengp+q+uadSjKNL6
saV+pfkdMdjTYS8wLi+2laZv4VXg+f9G98Eu3j0XEvq3dytN94CNYpG83T98ia3v
wbYsgL5sGyaAj/sYduZwYRLCQA3QV91qq0B/oQ5QN0+dtBKVTovj8/L1W0B8iuVA
Qb0gSXqKxbZrVMySfl+qeDUslUm2L6eC180Dm6yOWXPJHbP9hz7t7NX5lgYESwoK
J0huPVvbq6ZuNoVh6BCcNBuGiFxFeyoTZJu4IwjeqrkO3P3S6vhlLkAFX+IyYkqg
JWliTR64B8TvHxcAtbsrHrJTrCAJNQ4LnJFtELvFK1m5C1iIfqlmSVOH/P0zc/6a
ntrLpG6W17EIyEQFf9lsO1spTGDs7+pyTKbbGtipM7NjAgSrIULvOlsAv0XtTk9Z
dP2tPspuuCOQyUHc5gznt8/ULh6J84DI+eUw6UXzXxBNUydl3GFByK3LMNo/K6oW
f5ypwDlldQNJ0KrZjFhdBtOPAWFItRqdrV95KO+DDjs0Q4gJyI8vWkZO4dCli+XP
vaWyT86aGrho5XCFMO5QVEX9+KrF1G7YhFrIhIYLOSL2i8yMSQBdEd9jYBnih2qH
GBL3vF33NAzte+C45kt6lRGSpDHjyGGtGWNzqm6hQ2XxwkHnaiWKpM6VOG3dRJEM
c5cl83N6o26H646Nw8u4SKXep0ImGu+iQHUYMbmhg60lJDxPRCxmlLgP0B1iyuQ1
aMxAK73IsmEL5ydUR9C9/cYpRMep6q1M+2hj31WzF+iMwa7NC9umWtXdw84iO8ak
HoS10m7V6La1PF07/KSA0mcmUpPTV9YH+0oVTHv/d+yeLewujca7V5+QyGUMCebG
DZ4vJ76vqVtbFEaglEz829sUS1oqNeD5GcdLCzdM8gGLMPE+O4Lw6ir04CW8FS+g
mWsdoP4D+w2xoj+rSKBdb2PB1yJ/jSYUF4XdXj5o2XIq45N9+a1yt3yj7s1Y7AgM
kv9snPhyD8TM3cECExGMRHQjya73S5TwXKcashGa7VmVRfRIuATBwRsaR8ljrg+e
1V9w7x5virU8yp2TvK8jXAJq48AY+Xo9HokotWXEKmseoYSVpyYN7/StBvG+Akr+
c+EKSGILpObyM8BvOPDfIvBePuEunRKvv8SR64YL33AtMEZ5kxGOoucOGor7wgW/
GRbF9+/eaUA5H5fjqPoOKGUGv/ApESbXPytU+Ba65qEoLwIHq9U/TSBP9qB58+sD
g6+KFgAlW3bdTz0JJ6sXK3JIKfNfdKX+YLzmLDyYtixxsEKkV432FOKvaFlSRixC
OKzCmkbxxDXelAszJu0C66JwVLIRS6tmzRHNp/kvN+P/Amlk4AN6xjm2jphhHDrd
l5DrhnS5+8cXHACyTnj0bcrp6s4YRA3nVKrtgylufPnRiAmKSO9AXOPfdxxMTnID
1vcXbk80K4UXRcRg4H3q7OMt6D0SNJApO2SJ2znhCSoNh/ymIzTwd6X97TWhuZTj
wbzQLdKeuhHnSHtNDdYlCURGlRKnia6HDYKYRpkYRICBxX9hbnikJZvxV+iyrH9S
NKYtTxKv3qkWdDSZq9o95it+hVW2R3ROXrM70ZuMTVLsCDAQaUo5FNDQX9fJXGLE
iU11s87PONKEjPOSi3rs8MsJhhz5j5VPAwnTGRRYnuQ6VYqYtw0D3+HAn7zPx19H
PhFKlBFDAn49e4XKchq8x9xKowe23B9MfosfBmUzkuF4+qHLbKvIjpyYWecgYgoZ
EYbdjSM6XbaurAaR02NuhEoKdgBbAsOXMz5O/xozqNHCWMVunuvJq0gbz2ULg9Sk
FDn9w4TUwMWc+J8ksTmqIwguSTKsZ+Z2nanqWrDXAKibvlHhCIXSw9EnvRGjj7wK
EaOuvGR8qKyplsvZex8FYy3aOtYUpOTr+zF1qczDKtO30BUpXmIrB7l5g8ZULQYl
/KuKOkicFdgnYa+63yTJpJdqQ60vJ0XpMFI6BV/Wq9gQ48jof0s7isrH6XA46wv7
KCW53oFxLSRZUqLrxnDrzl01Uq+EKuiQjxEkoidhg98VWQ6WvDd1F806MZp0Kc8e
oyzJyGUOYntrWKI6uxMr+mVWIsz2k3tJRSB71HzcsSlWdtx2WHc/En7GcGAnvXhY
Aa0rYNeCnT9IJLb6/lpnfniG55HK4+KBGDHIQKDo/lbxXxZIiPrIENI5g1BMyR+4
WOU/3eU4UnVr6Ku2Apv2ACWLqwdwTxXAFeqXlprcF7BI3M7VW9Te3dOvBjQac1P0
44keT4XHBNztUPPJux1WYI14LNmQKD6mTardmWv3eLMO9KnpG4rgvi4DAA2Y93fL
Jezfa5eAnA9KTwi3y5Tkwcgb8Wo3t0pLegc+TRlmtJZ3F0/OOEjFGZNMsnuPkd7d
r5J5+/UMUpOk6gu60K997cWzIgMWCEi3zSVGKZbCTiHoGS1pGfXO0putWTu4WHst
EIcEi9c5vTY2PSlirzpYwKBYxPv5pjevWtkr7YEHRSFCylst2AjDzb2bKLAbT2t8
uSWdDOh6Mktd86eYoxIk+K0Wq0/1PN3bRbsJMF+mYp83xdvK0SsbEBD840uNHL40
PI7iMTiNMil7uy/J7pNgDiA3r+2qbUjdLi6yI8kydoeG8Qdylq79vWRv5NefjF7Z
JNRA+T1WTXW246GkIrXIZjmG9+JptMvM3nxPhYpDe1ta/SFyPSNF5y+6WK1Ke0UB
7Ig95553J83z16NzBkyqD4R2PaYdLTycY6LpcDKBIb0WrNgYbBdjZkk6p/3HAQky
KFQ8HOSFOMb1qNfuEiJ5cSH/oce/jekA4uUWjyWRduDAZiYH/HRaqff0P+LLS6ZN
b+nF7dq+serqcST3+baSSFzYZalrN830UqkhkNkbQdRXmdoZlSpPjU5PMoD3gYsX
eoxfu41jCEE5dqiXB5Iqxpad3r1woWQwnSgVcb9fEKrQldSJxM7HVKadTkYtLjMm
S6573uSvMui1jmCHfnIX5g46+UGJP4w2wT7+axQYE7/+iouGPfSS0KNUuvoBhEiD
huVUbyY97xIbbB9XR1L1jYMjj+SOZIpNOKCBUUslJSwZEItcD3D716fLQrZHIYuK
f7K0hnR4UU157ZVq9uu5UEMrtUNVI5nfBZe5sKA/qzlKfYW0MKHt//VFqI2ghxmr
1tLtLe8uxpAWCgooHZg9Juy1su7njjFfjk2E71nC0fXuMmcTPOc6IvAKWWlEvpBC
UDNcjmFALpN8qwFshIGvuPUHiIv64suImRwh9bPM8t+PcJsGvMWhLNq1VNc2xpl6
722d/m2GvI5H99IVCGk1u8BWyRORHEWpTtgZXbgXGp2Sk/1X7FdWt5VGZ0tzg20R
FHLpVSMe2dic05xl9r1C5qG/VDQ3ZKNBUtuaTMjKk7HC9w7zJNL3hqs2YyVYFbLi
V3jQ1pc+xKMYSI9TSON7eoFXciT5Sky9y69Za8NKrq1uXs0xGEjgPkxldQYWjwYZ
sTSzYMlf92/Ah47NB6dP2uaZVpb+WeMlHpZ5mnQjvXCP3a/K8MjSoo5fA5Nb24f8
8UBkmoWMVHBG7K9lGtmOiNuAOQsK82mKAHS5fr5xsOuxrjSAJaMFdz7/KfnzPcQY
A7rkeVRQ+RIK2EAdXdTlGeY7JjOg3GB6uf0vdTk3hb1OIlIFqgYDkpZ9FyLNxZXh
IVDuzhyeliAsuwPYX6WWLH9gjQTK59FNi9ef6zLo5C0nOY1X0ekGpuf54Fl1nzn7
uS+UT6ks11Im/ViwXMCiocMDccJs4AU2oUuW+Jcc/egd9esj1nU8kn3xpluEJqiD
ndT5rYUwZZKX1i7C+lYUpaDX2MafneBpn+audnkW5THLqkMlTikrnA8zzOI1eNk+
Zlqa9jG0c7QlOoDZQ3il/6ovUnDK0Bl+CYXbDvGshAzlTzhbKpMqlPe24spiiyxh
A/U5rQ+vWLVUk0MX9XePurgxK9g3SdMtb798ihZwzU21KUaD/qEyQsQsTI0+RZyg
HxSsWkGtAMq6s1ZWbw14q5A2dpjHTA7rgz2UJyE+uf03Ijke+jr4JNgqEoLra3nL
mK5EORxB8IMZs4irpmnyRqo7ZOHh/xdXxQUk/i4rXLa0jutzLt4ETAeWbl58ghNK
9DdZH775p5IKqoS7/m1EVudqSc+I1zYM566H6I3ZtfyajY3rV2u2JIQHipWD+scg
3Tb5oiZmm5xX1Z85aT0DDujfhEwZ4OCoKYB7PlXMbd7DVGhELVqGcQodclJaHCNv
QmOSX5777cIEBaTGGfZyFfmLJo3HZFGMbVrHRHx/YlBMEw/SaUkzP+0uZgvOez0W
ATLfoU6QNet/VoE6q76mOIq7bocGoJo6SlJK0kDZO1kqLONCvEvLAGvOm7j5QTa2
UQ/f+9iikJf7oPwWRsMWHVVODaWhpLDkaPi81WFUTDIXhMWtydcPbz63m+7ktTsz
X+BnRY9voULYEAwdbCbE6IByWwz/CsKemtccdKuARxwi10uNZzWniEe8v+BCQtl5
LBYGtKsCsAL1CBZmIYdA9KxRDPxXGzzhBaAyttoY1yUxq0idpMaCDItrOlMnGjKt
dPpGgMy8Y6ZknRfXH3eCmNTDVr8+ove+V1/jOrQOTyzEwZ74sk/NhlYG4ktVzsPA
iNgTJhj0Sbr+xYtB6H4FfXw5upw6kt2EV9j7K8/BQsrvjiwcvfYaUG63pp5EZc6q
yOBys6xn9J6jbZ8naS7V2Lp48G4wWyYzxqoUnlW7MlhpfNLmFM/TGHqzkxL2AqX5
eV7/bQPVsH5+CW5i7y0HNIYu8jswTg7xLE/86vjTXeLgvzgvOyNwb/VIf+2Df/OZ
qcPhKAq8EObInx+oxuztXuShbvetQ7bt2sra0FeoJ5jZyhb+6SowUFCX8QcRU4TF
OLQfsMiDx+CN6IlNDFHTFyyhh5q0k/SUsMwuZNcNA9H1rz4n7XhNyl0IU6pnjw94
RMLhiUQeZNRiwpCiWlU4r+VJWdvTv1oacDtCMq7ZPhaKyZD4h7YclA5MogdTd01j
xNoSdzXRGU84vqkxJx38Y//7ImbwVeRHegNLJa5AgXUcn5U2aEfCTaPcAeT38VIu
dNTb5Z8pOTXbNc18kILpLVyRJn8vFiAw/YY+fzoN3enGhQhFuhXjZkc2L41OfPWF
RxpRpVfcvpsZbekyLYFKB4I6u6RwHpe3KubciykgXBwIU7vvDNX299sL5nhRVCY3
294Md7lyK5lrk/YT/Ft2jRb0iuYX877fcTGBRMNapxxDh7fzBMRwz2LrZNwJjKHH
z/ygCyHzYTg100YL+hnuvAL5RS2vkLYXeB6ksXIzIgCOOTKkSJ6AokOb4E9IQpbR
EFzoNA6V/8tm75VKIpgP432PKokVZHKYtGQH+i+3ymwuKA7EyqvQEd5xOqKR0b/B
8wb2qDX5PNljmxDEl9lsFHbUVJWrRtzVb5eYVs3BwcqLCVDgRiDf9elKPOenWqcx
n/DS41g79zRIn5xxVUXWQPoIFHK22CBizaIUQHODwd46zZWd7AteiVvsCqKA/LS6
k7QIXvkUpdhVwZHnUPcopoWXitKyoONiyoWel3kTd6cL+TMRienbP+NPJeeHTba3
WLsLbnfnTXQWCnio8I6d7gaDnzTmhIjx2naTRodEHTI0z4oEv6SbxhxVfPdNy6qe
XktbFIgLGIT4ZeB/7l+JBzc+XKLh7ZkayMotyVQs+hEQTjTtB33uXilFOHcZszGk
ML1pOlvDIfH0id1QtNlO8GjIkv9s8+FYC0+ud+lMZJzGQjVWDHOTais/C/oN3ZaI
eT7ORu1TtyeNARNrobY+NbSkn7e0mv4RmBzvSVCwDLrs4rEQJnI/KFkpzmS2W77p
KvnsWXVbsErk6dH0ZTqpnAfufwznLsuutBJrhqSxVOtEPxbo701njlQRkxobYmnD
13afNcHlcPfZO+UJBrYIH6qPKFIo8jzDmHttd1C+Gk+dbEZC39f08Gw+nXlfNCuf
OSAgObSa0pUAC1KZKxLnEJcS5iKwR2/e0wLmAHpiHHA8ruJ6fmvMWLgqIfDO0eWs
VITAVaBm2KixkmW3KM6GL/WHLfjIZ33STveo303io4gYpaq94eHkQAJqipGuZDeQ
22KssajMQc2O3uAiqzgOegDFMH1PWk+1IYflhbxUokipb1fmih5eV6SnJ/huQePz
p7Tdq792VMN+Gyy/t/3peXSSyjwNXBabjaPd+NHRmFjjmhtZGRpNP/LFkOJF7fLp
MbR5yRpfmh6PvXTmAEhC3oQBsxjYk+pRFyygsfKIkozkGGnpUCMdmtndZnKM4+0I
iZ2hO0ShSXgHgnBNFlAttSRmXqN4oG47osfHI/olwmaOqF42m64RmSPzeCH7iodO
941gm5SOeB5d0R7XjCZ0HijpZIGkv0cMSAVuS6NYDxVQJZInoM5KGPdL4dhmuvaq
B66CtGQbRMr9TTcv3fh68ELVIF7mpigbqws2Sn1xS8ERBqIeJr3wB+lKZuHEoUmM
gqTN6R0kfp01ZrE7ZuVj2moJPYwiYOKQ8MjipIpyGA8KK/ARGDaiMHoy5O6QeF0/
a8p0tkdO0tqHW4i826P84ri1OqTTwSaRMUqwMPmD9BKm7se5cCMdtkRRq7cX/OZs
/RncCEirzvXSef7LDVa1vmtZUwfzvNbzehLKVH1wl27brZTr5bry1snvGM/w2r3X
3lzX1CK+1z4iVQ8rvfW69FvCxeHkGi18ODCXgpme5uGeO3GYKb47AsEDkY6qtRTX
bLGeTpALJcwMBbGuh+WI6S4m2qASChMtsbHHCOduCEDu/k7xuHrT/PH4kYmy0E9B
Cb/+hHOBkn3J8msnbDqcvFpkpMrSNbUeOLYEualC1gyfotINomYWhehG9N0CW4Ak
XT9OAngwLfQ7SB9FMP7CCQn9oyEL59d45lcw1tF+caTYbRuBNoBM8XaWVlMfrssH
HcuuegNy6nbT1OTLvu3SaoUG5tVmMEB4tuf4dZNV1afWPr+tbaLv05l5wW8hOkbo
AMOIUJfbIoP2v1umAEnDj4lEzRpEV3eBOMf+6WHUESKMW+PLkONVUrQt6bhVPiel
p4h7h3Cnoyf75TgfDDVCz8g8RUpspFBKv9gTZio9ymm82271VDZ1ENjYfq8E+hjB
t8QOs3oU6QzpYOi3B7pCBAHC7yzAsqOiTJ3XJsDRTbevUxxm3mGtuO5EmOddLmum
8UVb3DF5yRE+KE3WOQWPUPKymfXFtj7ogdijkEBlAs5F04+Dx5YLz5zGnnDQXKHQ
RqmNPzZ7VFf5BH96LXWiZFCNQ9EbHzrRxPQuspyWyT/BF5lgdkd8c9G9tMBh1B9N
PlWmijack4CizoqBo7SUtQ8VKnfX+FPuOWoTfvrYkWcGI4XxJQm7gtnewHGv36iQ
2aMXt70NO+WS0h13aMdXytrD8R962HpFKWm2cEI/gtgC6Xh8Ej/YlEXHMBJKTOyF
2d1yZF8PkLvdkR6lR9GzTbN05R0YfRVm2stl+WHmoZL8GxunwyMPVAvJl6wfoBiV
7SozaezDrlQKru2le05IQSYtN0oa1ZtPYmzLIAMmTRR46tTExn1+mvnyE1IBLjbB
1Si9t2bpZuAJDXeYQMpYKWHaTpAwoprxnZjE62GCBygFGtDMuK8q1gGlHBkCIaJb
UhQJfkEN0TcOJRvYTWrGiIjX0dxoH6KwXcCvR66H3DcoY/oOv4bNnvmm0XIy8mNa
RHapx5AuCoYZKKzAvdHrzrZnp5G66orqSwaOPgD1jeaaNSjCb/8KMRFE4wqCDLmf
90FhEqFQDqIj9tPyf8u7lpmAjjBS6ez1Y3ctzjFevBHlnHjohF1GY41/zXWU5h0m
m9nyDoG7uNAfGObI1D1roJ4hzSyL8Hn2fPwLs7+xwefrpv9DrJfw3CoruaOkF+UW
ynVy5ehPNVaFCj2/yWHrJkR6EjzF/GMZJpRns7DzEVbxCWtYolwV9nzYNC9Z4tBx
D8ssLiOSo0JRgbhvJV3W+K9W6HkS/6FB+mN7Af8oCMvuQSJLxhF/keVaHof5uRm6
Fazfz/1Ig+2mn2Yp3ZYuH8KTTAlvA29uqAIBTxpRA3IhiysnKVrtyJZHPzU97D4u
gJbrAa4UnmWpqDr4BUUYooEQ4p1v4mZG3D01pBRcM0oa25wXiZ0E0BDP0XAXYHyK
fFt1/R92h37UtMfONRElHYw77dTefxJYz+/tROqWShyHZPCDfmJo5aFexWD39e6a
DODIpOcNERm0ftJ13X9sKVokpfHICdOBwbcD+7XVUuK5SK3LxFJKeWu7GWpgHVYR
838FhVoqVdFp3W+jZ43hhzZ6ySB54ZdhFuLgBOHZZMqI2t6hGy6FXmf1FHfpDwGg
NtrXb9xuD9Y6JX4Ay1sT41W4ILZO+DjHhATa6XqJKrzkJ56Za+lO2b9gpkwXu2gT
oXm1vfeKawa2t6xAmaA0c3207KNi1fdtnwyKxqywZqLjUBqdncDjvnidOAFz8+1w
f+l7rzV4PCj1Umnv2GvXC1oNiTR7GI4zppA926/V2coxts0jd1IAUeZVJt5ZGN9z
/eOjApmZ7jTY5+xCZIK9e75LnjsHmH1dSUOJ5rEf0DB5PGskl7ocgvanTSm1uIXi
vEWzEgHwa1GzjuukTfzj03Vnd5xTRzYPfecdUdMFVc9B7WHcpAIbdxQLdIcQQKqc
Do1B2cbHbdTmjhxpr8NYe53QLV8Tg0zXWFaypIsgeqJLV3W8qhrY5PE1ngElxs9t
QjQwIaBDIpxrMgO6z3UiuIzhsbmyzeugWUjm/C74B8pc5IcF/zR34Pw32qBC9/Hy
nYwcDte5XiplKVkfdb1AksEg6NbcYPWT8s/ZU8NZLyDODSNPepVkaq+8+KTmpnzv
mIEiZ/Go1ouj/FO/6K+hfk4/xeOVFHIoN8aLY+hH6dJir2LKikTZzmc6ztRld0+6
zwl5IPVdy0DBRsFdeq0qbGF0zDG1r7ynjJBEiKDYZP5FQyTU0wGs9nc3zDYMz/cu
RCOlAZqNfou20f/7a096UY6wobb8H3caC6SsZIMN7+bVxgNdFZU2lI2wqii6oBx6
4aYv2fqOpnkLmT/IhRQJaTH6eRgV81hcILboFTZfIy32O+WXf7ViOSVrxZ9x1OG2
3ZpqaNVnhP2ktzCT7bZsL593jFJVfiVJ+l6PTBIpTbmG/j6/tO00eKZ7OMHFNRdO
mXQsIwGjnw+h9n2zK6UK/P2dyuaN73XA0bG2sn/7BKWe8Pm/emnhiHl9Sp9iNI25
AkfLHMt6RFjlNMHMUMKILdL/lPLZkkwnncpnzi5ZIBFc7MFARAvbdUJYONRlamZD
VPMAajcjg+7k9gjofvH86WtbXebp5V/fZ+QRCvbPLmOvdKARA9bmXbs7dTB4TrTk
iuwORyMKaPiAPOFXeRLnUaIqnCGZct3u11ETCbwD+VUhTQCjrHGHuhFem9Q1eohl
NoTPGahRUIxAPNkP/cL6n4UZgAGX9QHv2zE9p/UchpgHPGZh3WX3S1GozX+ix4Jz
JMpORshRtFkwsPOv9nljnDV7y0OVjaulzqxTkFusszngZdZEKM6LZ19bqPSDkvkB
UDA/QXc8LFj3D88WweqWpdMJDPkQb7OZ8vHyFDuPoDFytAmuztvZeQU91NAM+jwe
6teMMCL816DnjWs7LUhvp6o5ayfZYH+XH0hg4a3sfRqzkm/Kj/4ELVfHKAFsJSey
gWdfI8ELfUyjbWcNtkXx07OD5jxaN1PAIXPSHonSRbFQo/8KtPQY6LV3lWJqcL7L
0X3MPyrWGZ3eEDErIdp7tPJ1i7PfkkNWQRO3JdclB5pkggxvGFzKozbPd5d7vDT5
Tdk5l55XDNxUgbnw8SZZmKL5eoB72X72RyPB+iVZLDD46be3EoJNvXOw/RoLTBc5
t29BSejWIGHfMKdD526kv3e3vULyRKHZAHFARKqkMBJhuVc3X0Mt8F4mGx0jEbFW
VzoLIZObkSfu/cR+qYGI+ne6Kk4pRKj2ONRTOCvfAhRYu7fIWkaBKb6uQOCn37I3
RNaUmHI5pPc8B62RaNhNML3TeGIeWopZ+ICgy/JsldiozsVPOCL0zNhC3T0Lf4oS
URIPa2gvxlRsuujkLpfMKSkJzAeK9saylmbUzGpzFjXCkaAn79yX6KES0K4zNhXs
5kw5rEyVMC7bckMaJXdXGvoJHHmNFWMJGXssWNTYLHg5v15zbOu59/P0wvOjmQwy
omPopkBAnn+DfHG7zph01QrqWA/unbftgSrkcK6h+adSb+12Hi3dTcy2MvsG0uFf
qK+tJbdfJXaFhjJaRIjIQpuTlxKHvcQHXX4nY+GqFOg+ASufu5LBVlJGgHOGACCQ
5KfyjfNzjWnRJcKJo2dQD6uv86im4FexvwN1oUdUeFCH96GYmLQa4groMbXFIZKe
Vgx96XevmgQZ2VHjIxlBjJyPKw/pQiHyPqp8gGjfr/JF1Pn6FFBl1usKtsTtpNbe
cAd3ywIW/uakIyXdzcKRZBd/IF/mZFHhVQT9bSlT9vlaH3mWwyYBgxGNXjZrusJP
oTpIG0eZgw9Er3lH5l8wVhBhosSlO/liSMcm69R7lrzcLmUp9uRD3FW7quITb7EP
VCyVm3J5d8KcK1bHrXSx8RIbgT9UkAuLm6HbBgceBE+WDHzars5LIMFpavZOJxA4
ltGt2n9FT59iQbpSiLOMF6C4jZR+q36lXpuzjo0nb5zZ4HCUAWklufNkxBd4iblS
0NxhKcR/lq8Z7Wqxdk5w0AgQpNduhZH0vZm+gH6kRERHPgbTo2fay5VqoaUWAGmh
IC6U0iZ+SKw0dJjvSY3nrVBxH5TBa2PzpL8j2aGP6eNKAbbB9eflKmJGmmv1hrzz
pzHEjVfvj0GibDGw1XK18Q5wZrhMKTzs4b811Jvw7usOSJlhp/LMXs/qQUB0ziPQ
HTXCCG36v3Q+9E/1rGFPl4bglpwgc1TUK73/T2g6ancOke3xkerY8GKdO2cyy9JB
myj9yNMz+hwkOqo3MYblDQKse98QPnB1QZR94Wqr5RBrtPDVMM82kqkju4muqBPE
BEZXJzn43vkc6s5aj+VacLc9qGi8XUd8wW8bDSkm1mKo19HvBRjox/jXSpkr1vzl
r19N7TIpwZbMI07UWQDlhdE0nXc7qAKWWDU9a3uZJieKGiIrUjCzMbJV833kJc2b
MFkvyo6Znl5gO/lz3BWjkL9p0U3eqQGVgta1IYkZ9nDs65p0urNXfwW+o555D/h0
Iip72qMyTBRG1+k2OaaYWDPV+1ipuWHeYVJIBuvMAeg+5pyYqvrmxUobQX5DvLYC
huD2PKW51IUEZ0Pultwt8hhR7q7wFUQYFJXWLXqN6GcP23zi22WESFQSh+b+QGiK
CYlKPKzkHj+trcewDUxz7RsDVmCqlApx737VlfQDdJRoJv1Ewnh6mLnwmLNm2u+Y
WeKuimWmBZQTlOgKYIM+5TxzCN7yKvjYwblWUQfGM75adMQ+zWL7lVUI+iLy6mRY
e7R2QTTYnX+loNdAKVXNsR2V/PWHxxA7frgo8UBPXs0VjCc6gxE+MWeWTCl76+PB
3oDYabrBke8EnhVX/2nyuMnsrJ/CY6WWpOs2glDxsEjhNf1m6cVSIQJnYZt6YFnn
pEKmX4z9wIsQffXoHuKh2/87xsCELYc1Ya2O10CauF/5g4J8Vf6bmcSs9f/xU3ZO
pivbp3mL9YP4RCpoLyXUgJ3rao+zE+nOtjZPVuZXCn/OB5pf/Icyyn6flTiyngnF
v+MMn6fcPVQUPyNLRGvhVPkOcweERZKByZWPiSPm2vIPNGfSi3LHR/rkzFf71ocO
7nPFXyyvAJW8dwGOJaMz+29XtBD+jo1fsQDV8qEjilm1sJZLj5iJOFp/G6SMC1//
AhBJ+ZTqOo2XRCe1eBeJw/Fh/6THaHDo5kUEK4fj45BWRv4Vt6+653Nsw4rErY3O
UZCnxEl7+L7rNCE6Lgy8hgz7bZMg+THgD9sqma0QoQxT6ql1zzL6A7QmFSJXMY7G
1BqaA6Usz+QdhV31GMHowNi9JqKXcV7TYUy0gjok+Xbjdb+eCgMJyQp7u+RDuUx1
Sa4sJi96xDel+W8kNMHTTD9PtKY3tDk1/BaxR4wbZdTLr2bdPzm0GFdg/ppWAYff
SJ5S22+B86atuhFtcm3LWukylm1RKLRz+KPax4O9K9y+VqzZy4nk84imnp2hTyFz
aSP7Ki8jFpzE3ADY4TWV/xuiGUZFrzfL5n9RR/qRi31t4ZPJZNfi2FPfMLh9YfGq
q0yqo3xYwQA5cO9c+2YJS10KlwuGt20mmSSH6u1Rb7AKikOg275Z2SWpdMj7qyDn
YH/JKL45HINlzQzxszA6ThtKZSWBdV2BYKkY7vTI9o505ZbTrR5EA3lr+m5VLn0Y
EYlhxvfXxMhxmjzqECQD+h0lHDJjle4Ox9MNw2OZMzH6WDWOii10JwCAzUF0h4NP
mE4A26tnKbJ4f6VU9hzTrKZyhy0EPtnWeJ8zWGfailxF4h+Nns4LDOWhRi0XulzG
TZSEgU8YyEPBch/xSrvbrAd9+6+aB4H/LEr2Ukcm4CgdVn6aoJ91czTnKOkxYL3R
Y5DWzDqIea3uTRXudBRyg953vj4/In5Eo9UtGAuq0Z/a3u2tbH9mgrK4U58/UUWc
I05xgVDWL546xdXvMpdS9FMhby5kOA5zh9kMYhV+OBULtSNyQS2Y4eKcbwl5ukOZ
K09XxerTMuirqGWwFxtFqYzqmRThEntr4tD35inoTQlLoVpfEJOeFtXoK4buyj3l
AeRIr8HEAs1aGvp5oNR9NPoiegP1EXz794E8BpLqiE7sLuCHN7H40FkFMcHVj+o0
dRJbgHqh143t9+Bvtl88MQF3XgNSoThfZZu6IH84/9o0ZTnu8cdq5ou7QirE0+DY
hJUslgWHZ76W5DSMYWRcoR4RUPu0vsTkr4acyfjFOsZgq2BPFnorLsD4MpAc8P9c
AeH/9UWlRi7BuczmM5vBPTOTLyYrBhdyiAe2PwKtbpYY03/ZYj7wBELgo+v9xTvO
CGIVhUZwuhhb8m6ymOtWdecX4MBBrv1LfDZb587RwVEhJfn/aFk7FLbtrpT7V/xk
zpYfZFgjwDZaMNP2HcR0pSi3XXx+0yMQXOm53FQzO0SEkRPaNAGM/UKTLOhc6uBf
bBhRkT0dywb6JG4MfxEQcA59/CP/g5bal/h9VHRU6gniEYtA/9TbBdoE6QYbi3ah
a2t321c98M7Z2Zq3On1gpbBwhKsy0wdzDxY8thB4kx55+hXelnNJiPzVzJMqpmAg
dwav0rqxS86YsYQWk5yAsHjwQYhhSho3RCvv8OXVpIlf/ufyrxgrUIOnDwI8ArjP
ZUhNC82P+nIGEL2kIL12wtx1xMPZ8p4ikHqDVv/9tTK0fkarTO+4CNXrEUlmYGua
WyvwjT/Vhj2thehnHj69W0Ol2hyz2xXUW/XLxEaemOzaqdLgjctDYbcQvnqtfoKK
IyNDLo0UM+VbVOQ0DniijahlDPvI1ogtBC4gozIJH7k/D4PZ+V8DXor4FIIQRb6t
H34cJwsebMLNCdQzADCLPXf6IcIQcN9HS9tFTJhmNVe2gALWXuauRTk4ymIC0Zfu
Z9W/Csc4L6pHHkCDhwDB4WvV8+iua6JwButM3kKbZ7bhlFk1LJtaX+nZ5rBJU4ar
pZ///pC55Jjk+bqsCPRegzfssYlTwFXP8OQi2WsgC3JAg8/am4nrinScgRUZGsCd
Mf0NZSQXgCocYq7ol0FCDle5IVnDEYIMghwPj0r8K696ZXjAjlAIY+xLr6QDE8qc
PauOs/44OLbqYDTwTpHPk1kj1evh9qw21utspk5D2TeWc3vTCVvY2umTB4R+UvKK
adaX2IchY03q4+eHroFmY/P2QESDLdmY6085/FwG4CMKrZwzEucTvhUA2li0a1Wp
yQWFovkgurMZnHX6EZtDqnOerF33QHO77QE1qhXe+LasGbfwVkqTW99j780Lzows
Nd5gdNKwZ8E5md3PvX0l9ynNQpFqu6JxCSYNA2ACn0P+71yfK+hCEU/qd0i2KS/s
vJgOcopZtZ4mowH7WUoBYJH0PU+CzpZV14q77s8Fgwj6wfkAUgjHGcDpxP3z3U7k
obBfl9R7lyygcFbrn+8iPvQZ+0z8lwCNt/rmhRvOQsLkaqlOs378QSyFGPPdQBIQ
zjeT4NyRq214Bb/kYoh7DQaPBH51abMt/qCZTAc8IYMemSeH/CqXnMyY6oMNHDm7
AIg+HbYIteMKWlPefTn5uJwubQawueoSuam4aDUAUZv8lJT12j5ShMVixjeaB+er
ypbHLfYCoxKhiV3xlGftH9nrxTVeC9aluDdj5ga8MoZZL4tQ706Pg/iiBjlk/8/c
RhSA2IBDwOJ7jvyI4c2NTKGNb5uGwwzjjjHdk22BYuDX3/xdYeX19teDNxi6oKLz
n8fRyIEAMbemNuOJoVBbqPJ3tU9TLhi4KFLRjRvL3O8/AcQV/7WvDgceD3gtOpJH
W9kBbmAxjjsfVzQM/vuqt3FqrSvxoNCyXOdoUPKxQM8h3FJi4rq1ZVVwtpV46dXD
Mf8di1hWqjEpQeXFmqyh1aiyFmwjeuSMrRpHj1cI3KxZn8MG3oAI9EHy1l5A86cp
xzjU5jIuXY/asvwk1ZW2YBOTR0W8/DojvEDOXq564l2sLrWqDLnSD5Jo9r+7+r5S
FwGCymivbK7D+0Dp+mQUoWaq8RZ6aZ3h4VcCS4FFmDAI/53zZ5Ulhx30BwATN71V
apMnvDnQqKKHfhvqmMGfQhFHzxkqGX9s4n27+WIPudTB4JCUa5cYJucMQ/RW0fAa
zjX5ED6vb/oLEIdJXlU3Sp7C5m9HL+xBNfRjmqZlta0iKHztfJaH29nvfnZRLkKh
1eISFKNcg/TmWC1olzb9KVD7Et0eLnPQd7WDbTRV2pyiluTLq9da36LaPLcncCp3
HOqceKD9OEdXbRAAF3+FOhsQUTJVKJVl1aTNI/YoDj2G45VdwCOZycZMOeqGAcuD
V1gU6jjVpy48pLX+J55EbD9bTQCwzzLzVe8/GOa7PAeta92gXZFoBE9uQh5Twt5x
xbEI7zbE/1OLLHa7SijagXMDezrondKdQuh0UGqZKnhftzhub5Iegn0uQrvoHCc6
wreaPLmgNocFYUv9V66Fw14DUn5Lp6YsKiRFQryZfISGsmDvijV4IEPOlnwDSbSx
5Gewsz8nIMG6qmc59ViLK9PSXVtQEKbH1S59m36QW4R/LQW1VSM+DQ6+F7ioKPgl
Pn7l8WYEOGYUU7U9GIeoiHfJIuoJjNNNmkCEu3wIr1tHkIn+tD2OOFtHKtGyn8wZ
BtAVrEBavraN0ERkbPBoGBecYTgdumq3ZOS7O1p+LreQ2YtMUln1o3zkJWv32P33
PWYGCZ/+YGZZAwb0dOIsVHdO4dnBvGVs/yA6jJILr12pbCkLNGaUwebJXjwNUXRZ
L9IGUeGJY6Azs75mZtH6QUukDYBrIdPJnO+QPDHNISfqQ52gX4R6gXPVxK8sU8at
YcXSZI+baWCeOdJUFfx6fwsez3A0vorL0wE2q4Xsat3txk5qSJbATCbIe3d2xhgS
mDYcIkQwu0wfFxifL74NW0sP6h0IjOqTz7AJ2iOJZ8AhnWxJwxC71Ayi0DMKBNnp
N+Mj/6nzivsQYon4TAneBKZwnwOpjAaUH1udKAMr6MPokCBcUts8GtddABpj1U+9
iS3RyI2B9LGE62TsMxxm6ReW1NgbXw6wQ4wllUiVOo6iyCP4Ij/T2WcHILE9UR+W
4+UGtW/tjBjNgbHtbS0Qdoj3RB4GqDeVb8ZYD2lIVpUSnWNoBX/qt+UJ1HRBgFda
xC/u5PRdkDjKprRB/C1GaU27iFBatFn6XPLt6eSL815WYuctFfPIJywtJwIfznIe
94HESsPopmVbJ3Mp1rdgXAO6f2lRUnp67MxTR0WuLeM8ukTf+NfLnzmGEkYdIDDb
FQ9FA2c3sH+mhj8wOgGvzOVsUSOI5YGXXTUhGSfTtTPEv6BI9PADaLL48/PZ6k6W
ZT31BZNb2xxaT5WcD4znei62ouXM/qdxeehsoXocKXij0fTFkExdvCSPKGJTDnp8
pvL3+6piW1CJr+DEEah91cCMm0sy6jLuNGRq+G72iepOJxe8z16fWkyG9sEmWkOB
gtTNeS5WAgx317smupoQM6BWHnYuBORtnJiqEj29kSi16NV9ooJl/LFq0zxD1CTo
tUGGe1UTQMKOWdbs8BlI64F0Min7ojh+pKWqA9V/A3eF6igm9bFaGPX5am4uu0fF
4oh+yRhA10A3MzehjrGvsbZrPKACacO9/GctPohqm5AP1/Q7p5Uzje/Hl6i1j6xH
f5kf1GK4DTGquUcKeXv/MmeWK7s1W7Xiyr2pY3V37kpZTLl085XkYYWDZ5q1W4hC
QR8u0a0DFiTEFTdKhqOOP8oD4KQA2bPAEnNWQEUjNVCD1G5k3YKHYsTBfSwm1eKs
XTgII05EpUS1GQF5Hwx9Qdi9BW+aHpKJ3lSFrSCxqTl+3kM1jqSkOwWgahg92jrs
FenZE+dt4bwu0X5m+0sh+JcH29tAR3DfjNfzyaSyDEuQIRY85QMDfcJz9p8Um00I
gg1eC+/2GQWRVRlU5+9FGmAvbXl48LaulVhMN6rZsSroqJjdA14AU7sAZz8Nj34r
Ro916xnvjM86pmcZUCrf68WlCVGLUZRUkp30NlGqBRFBoJ1hx1Bt/fx1Iq3IxOGZ
AoeuybdmpnxC+5AL9qDkn4WZ9JNxSiroKwEyTrisHQD67kHffLAHcVJ2ylvH/Nhs
hK1W0iYV3MH4Ko6lbC87pQ0C7wD+0kPvG3mRx4DrGIIVWa+C0XHwSgZgTqK7LVoR
ywHLJYPgSWnctzyqwHmVO+QFEJ08OJ/z6E8yyINABdITQvT035desw10GXh53kjk
uS0pSpY9H88TBndTjGGY6LSilBpiV57Q5Wnyr3rmrRXVxXuax/7bijZFZegrQ1Aq
W5UtzwFh6K5XES4oF/NQWNRxQEpCmbfnm3kSF70YR5rOo/kP/7W/wDTjpjzDWapT
cXyvFfL+/utqQ49vqPVXRi9sNnRiQEM5Df9tNgW3DYQtfVg11hDDJV0b51AUQ701
NgT4IK1YNP1xj6Z2bpNjm6E7eMghEojvvWaFF/rEMxW7rrP5NsIpoDVX10GJ8iLv
8vzJi2lSFjiSLMpve05balkpB+lrMq2ySNpUmPqvxgZJAmY44MUw7TwlrS7zgOcu
R44Yz+zTN0vjTOPfqF8/5rjOG52oYnitK+QomMjPZIS9DtvUVcMEmblrPmH7BKyD
2rcfsrNXw5bplHY4glhdWjkbddwNHy9XZ1XbPDQI1BejR31C8YGYH67mzV+PMbSr
LNI87/sNlIFTumzWMsC+S46l0fvV2Lo//Qis4cmBE5VKGR1BTcbLSw+sECk03Srn
+TQtuSDc0pTObyMFD0qPhBDnclihfnVZAUm3inu6yuULRwwFhh3c7ns1nnhHDeA+
zRlE/yOW6WA/+39vzGVC1l921YkHp26R7wdzr/l0lw12kjwTpXUes8ZfhQ0U3rg1
8ZaiTxVqdxYOJPqgWJHNP+8PMvaTDRgTvbz94a2Rxy1j4wy4enouvPPKt9AvBpop
lilX+b/ywi7TKumGOVjdQ+HmJRlrs9ILL8Lj8MU2lQdLxiSunACTPr/PXLrAoAIb
mncz+e42BGasSdRhH/sMZRvGhP5Qkq9NaE9TXPvqMPT3xSyQ583HjaPByEZCHL/t
10X3hbqI2mwToekOtYKzcpAJH1YLA4LqI0A5wZsHVcJc9uOvCqO5GRDHv+CEq33X
aWm6sN9iOPp0nm4598ACYYyKExBS7PVBGQE4kEvj1CFpKrGbRe41Vqe5kULQapav
Gh15ei+IEIYGF27Zd4oWLJLGf7y2kVxJgZPabPzkC7WGjFpe8/IskoXL2nvul3zX
jJN06nwmZrNEOMzTIs/HH3vQK1h34T+kv0WYzC35imoRDpIqJVGISK4SicynFC3Z
N1G5IhByRZ3257nW8AYhHmei3JZsGG3FWyqhSISIgpITiIqj6uuwgvpjLpqxwA6h
4vhUC49Ppk9C0ARlbXOug+No26/FkCidQXN1dzh6l4uzx+fWNPsktkbGK/IcrXWc
Ta+u4BQEK3rtTXevvqOW76U/Y5oq5PkvtboegXmyz4310qDVFJopUF/ziGNHQU9k
Zq2M629NLLyjW5wmJKw6gZFlykufqMKYeYePOh5rYL/MGUN8XfCXqWXpNyoqSxoC
3SNnKyEh6VqkoAIAURH6jChA0bPrLYfYPG0/2Aga3nh/Plz1e8w4oak4CKIfPzQ9
t2jszodEJJoIo83qwUYV24Qf0isc672ec9YzP4XfHXz8aKrG2kQKaGxrbsCpBTsn
/bEQ/wue2zIOfee+2+KY0pYN6PRTbturWoj8mbttNFoCeKeLCvIjZsEllt/lHeZ/
vsNrJTYayWJr67r82UOJRfgeQ6judqt0T2rqwOfdNCYXK6pqIL0BwEzWzuBu3dhv
BxYYDrzWIkhrEFiC9l9ldQaL4sBnFGufUjDMO60XxAEAYqJlbzZznV55zzOpNVGC
YQgoCjpbHOxOKgWTDHjhTy1v6qmQpJxa/jJIcJ0jcMjtA7aGfBTP+0I8q7qEvKKF
Q1lxbiIzkRvKvcKSQZ3frK2bZE9P8Sacfx8Qdwjik5xaobdWK5zLYpwx6PxZdizv
kcXdIdw3TssgGUDLBQmWCyDLvxRz40OEyl2El/tOAO/ITfTrT/1pMfNrjA7pg1Zy
krK06q0rF1ZGj80sd5biPfUDCdIWNarbSL2zzkosQlTShRKdzWNEjcjCbLrquYIR
cuicJbXwcso+hoHJAsjggXLGD+X8laxps6U+TdgXRqAJ8icjZeVtYNEhzOL0c29I
Bxk5Hgti4mnd0K1HsNf++dgtLcArUHlcL5UW454n07etSYoZfwm4Jk/EK6Et8N5x
P1z/A2v4YlIfTwd7SxUAiCM+SlXfYF0e/CwSRV3Su8BisJz8tiEEh9QR1GMwZyFO
6rnfENlYeyx04qDhuHhOUI97cdUCe06wfHCVFsLvkI8AOvS2veA3V/CXEv81pgW1
Zg544BNjKqP+DVAiOktyrC3+5etwbDIW0gimJjuujBLryrJ1jSOhHVQoi0dfP528
PQadTCEq+z5S0oDjyYXvLn8SxEbvnqsIqd0xOz9p2FQ9M3Rk3pvAZFs2dZhtU9OV
yTobMOPNPXbURHK2vCdGFSoQ1106dfwjL4AaxoEcM3UxkS9CvJ466uPvKW1xtxXL
4mB9LYSGqrOSryZSTOGE1RENTa8IGFvtsY9qdPMMzhXwnex85XMLgkRnYAnszezX
lykseanmoxX+svEJjXK4be1i5CUS7dMQt1O7/o6v1AkChXdwsTE+V06IfR32H6ZD
HzvZr7IM3igtSgkJCLmBM7c2CRx5Cg5HrAm+iyDf+kumHq/T8qaexTHlrYeNdqAg
WUVJKHkLP6UnKmcC98vcBM8nlvo3H1+MCYc5/BNzy7yFwlGQALI34lTa/D8JgxKD
p9Aj/BVdfQspbDY5G66E7N2m87lOqaotJdOKBeOMtmv5mVTbQc8Fa3odlx2VIPQ9
rGqf0u0Wcx8I9lkk6teqp5zql/Nu66TKNwAVrXx8zAbTLNUymQVVqQqbFxjGMx1F
Ze3mxdSAZ32kUyK8O0zF4ditn52VtW3XJsBncl9KVAjw2iUYyxkCWSVeaSgv61uM
J7qKpHZYhKzwqXzfS3+X2dnLUy/ofOMO1zviebaLJxd69b+HXD6iAkkGF0hKdFn5
+qYr4301BHn6ZNErFjOnfImAqBvCWoUEktxHOFfSmDsM596tvYYeamPjbv/EPQgc
lvoeDX/wO+xkVECNnyqYIkDLsdb1FnX6P/q7bIR+p1Nyg1Hob+m9dUsBAZb1c2PZ
Vai71ywEf9xw71H8auxu0nEuqi3Xvgg2Wg+NrIfEpOz6ImXzcMlk4clHOTI6rmpB
EmNifia9jb8XOvzdzdRmgoqp0kuR5iNXUPaWIICtXULaD5pvcyIkXhlGsjdURsRy
wYuIezCkNNcyIjgqLGCuHpJ834gCXIPDZLiBCIWsBBYOJaXpDIJMA1YkoNHgwfSx
IlingB2HY3elyiWWbCOalQXwDLSDHi/Ci1HoVPzgjk5/l+J0345lB3a8Tx/nVmZX
BdNj0Xqu+0RkAF6lIssN/vrLTsiMhwIy2KANiHxrbo6NzpqzBLyS9fShkMbuhGeJ
kzqiM+VgxHVzy1kn9/Nu2KJUlkqPLw0fvVnvwIe0uLVJwTF8rt/8mHzsea4eLTdl
gihxjBx+PAVL0WPXBQCg2XsxsXTq+Ds5sl6br7caKsHJKeEHzqdZ9b3otBtZtKao
zAumD7xpcA6aDflzLiYEBiv7/xgn7Rp/mrm06yQnsL9QRQFDa/0RO+eVUfX1grjc
ie0N/1y05cuR84uJg5YVyOAk8cFHOp/DZtYNLYCcOiaQ+846jsDcWztYNZ/KHrnZ
8I0pF8i9i25BGpcdTw5CznY8SHhmptxHdi5z0IsGnjIaAVBUvs/YJrrYC17erPRi
QiL8upgrRPpBBRCR9L9Bg2Id7Q4XeLPxuKbkRxIEAaufOtkTqkETole50VjV8HQw
9SOv7bhFMBmj30qNtv1B/92m1JGaUf6ctH8y0Tru6HzBaFGMZePPEh7okwPdRVzH
YA7Gl4QH3HKru7QyD1sR3rsQedxArcaS+csjxgFCPkLpst0rzNJcr3nlXskKI4VR
tfzRbuzmAO84u9hTh5p5F0QIf43CnY7srxfWatbtQ6Gz/yzbUweNR05R7XF9jtHW
WAIal1qQFCa0/JlHO8UeDhD5DbrhCBX2+CWkN1PeobqY9V4AKPnjobuGnazEep7G
JoOdVHvVix6YpzDG3Cr4LC8PODjq+K7RBfdUBwL2aXmxec10vbYnCOsUr7grXkag
gayixUsfeOX89t3SOy7Fko3RA+A3kHJi586bSyKO8mqz2SZguZfPddwhdXQi13p1
PgyjPPmtHgwcdbzoKWhW8Q08sjPiUcP6/Lk67xRl65CaR21qa6gcUNe4AkXvPWcT
sdN66jvuewATREkewlNcAG5MuUiFcnZ9p/SmzE8D0BXkv+qPt7uU/TgnEilPD7S5
+z3MxSyHPC9wM51nU7ng4G/a8H4WeLOQO2OfL4rJjHfcFTX/H3oCKNNUdnCxNZY/
L+EHnfo5pjEGVkik8vJkDYmN0OdK+to8JaIHJUtUhOPWhrxfxJvwW32QKkuBOSMX
qz67TgO1F57eb2OtNSl49BwoQJ+UWDsmM3hjXvFPa1tnComaFO/lT04ABtxCxfCW
zm3tWOcWlT+cAgiLY4k8Q4ozjjDT7B22pvQ7i/9+qBnuY/D6xi13FrPKXDaSlq0f
rUXT1mcCDFQg5z7VPAW44tevM67A4d5s7VKFXp/NRrkxIoIqtUBIdkwsorPVNpGO
CxAxJDupcfU0QR0dmXdYapdCtfG9rVJaLVn+RFtaiAZ21eDfyDUpGHIvh8+AX0LP
XHXLbCc4F8lECDXI9F7Umaj9j5GNn+/evG4vOiWwP1TccNjvJPTMpPn31AeSfrd1
8IBypSzBYT/FUyuak05ORIm4Nviu0sMFlkmc/L8yTktHIOzHRM0uTxvo1v9VuY/V
XvuIW7k5pGXEg+jMN7CquLU1jBVJahnI7wUR4UtPYbt/OdcxSssZ6THW8COeGMdC
y3bbmH8+LUBle3NBWntwR7xsEitiX6skwcr+d/r2I0RWv7XZmaRc1AmhFc6l6KxL
1KtpsosOLqEKl4eJVsD2crBf0uPvxQNGQe4KVo1QGOMQFymiGOK/C30OPzm80YZD
/RnI0Bch50Cmvu8TQXIm79PIhjBIBce1xR0u0FMQxUaMc6TldjOyp53QvqtYWGH0
VrphXylTDBteBVtm/UvBabJ1/lTPw/c10C4PJng3GIoFYtmu9IJfSlcxwCXRjufn
ksgHnIvUlJPZPEXcvjZSA5TFUpp2/Mfbob7NlEsqC2s3+xvA1XN+L8xloVwMSJnN
2ukgkK1qz6VEeNATS65FsGgZueICC5qiYXDzpijGhU1MBC4+P92EAXS8cYxQGlLx
RmMiJJpEC2MYln2gkBV9BPEvPoZz+2bc0jJ9Hlc7PIKK2+IKfCmtP2XyFs8rdyHB
+3gdpcoSU8Wqhf9mOFkD8Dgca07HSyf43aDWCJdeyj46BwkvTU91Vfja+Lq4VGgh
QF5BNNyJ3RxS2EZQ98bzAoZz3lwy1nfihT4ESSOHdRTMwy15nQD0wflSBObXIuFi
V3lteOTKqgTRQMdqDgNVsX3vR7Lc8NQt0FLdVq32qOxVVB5ZwlMcVkJBbSSpY6U8
LKmKuxBkqZBUlKPbzA6nJl0Ihz3S3W0zcqAdhk0GiER/RrqgKex2bh1WFowzIzwg
iWqLq7F5xBMs8HRmXDXK4WTU/RF9no9DBWSY3ua/HLBZLxbrHnRfPN5Syh5jjn5G
S1iNIZeASHZF5eLu6/FWPk71rDQgv8h0BvQ1h2qS+9k0cBhYpeoZVdBKwLW+QUSy
uVcvafaOElDco2FsURfrtZK2X3Tzwf8Qs1eMiDgVHea3Osekdh/U5ugJBkyRTUX9
OGcSfFwLDRQkEEqG10k6bLQNNKCqVERgsHWKhsk1EMKGcz6lGH4YCU2kJeulV0bZ
p7eXoeBkn7izP/jzRIa8q03p13VdQq1jGKM6gE2PXPSnSLy/KAXNtjMFnRQpTfol
AoSBItsKo2BSe/RNHZYlg8Rggm7ObB48j09CZ9OyW8sIHCV9cEswAtYA4A9+jhsx
QqEaX2nwyZ7AlX/mM+7pS5AhQEhMTfOBP45YCC2wWZz/Z2NjGUDramdGAmaDedj7
cLcaAeeipDs40QHcNn4lzS7YUO19UYKxCGl37k3PqFxzcz+rfBGbxfoFJXodIufH
aJv7M+aQKb6VBo/ZMRZX6lvXfd62cX6ntg+gZEWdMOvnSJ55P/YmOcbwV64M5RQE
IN5umW38FMpNrY2Sj4cI9YohbSHzvnAoO/fxn80mmBUsvNfWYkx4PdFUn9Uym/lp
C2qrw1aqU+bJn4Qfq2RnJe+umx/fI4nNHACHoGWOB+R1RKTZ9ZshircD3pRw0UUW
LSbGmUFYRz7TFc7BNeg/lokVe7oAc7zX06d7naQ+8C3zjWzuD0ACUw0nJ29VOT1m
74WzUcalRJxOJ2akx7AZqBpwLMhGfn2AFktID/IBBw4wqfZ5BqC02eyM/DmcnTM4
ZNtVd9GBgWTsAv6jG8YQU7NcLnkAihmwKd715R77FSROFLdoPz+XvD9iOhGgC3a1
y2+T//dM8BrzYyf8wE59u6ewmDjysIDW/h8/ENeK6RBaEtQ5dHEKPmhgU43EGa13
FzDEL/LMjPnDIDrFpUvlN6N+lH4gPFGsL67/bT4SPpWywhP2dLQGUrgo7JysvoHB
nYRanLTo/nF7g8LVOSDTpsPCOgNoNcxPwr4vaAV4DL4saXsoEM4TBf6Y0VbJp9ra
eLTybwnnqOJEaQ+C8CY09qPsOvi6WXfrKqdylOJSNbVGIpvPtyHb4sMvQLEiOXk3
3X5/xotDOdJHL1kvd0fGYrc5qdhYeAcgFrEtG6IRg2+hDjBgc3VRdNshW11TRxQK
aq4jHT38CgestjBg9HKEN6ARR3LJBBL6oq9dl7thnmZPQxPGTg24QP6FiOo7Ebm5
l1cQHkdA0Jey//+ioti851AyB7MMJ5dzpVs3R3jLTSriY1ElEk98YU3RxP62Idqi
shwJRxPmGgnB4LWrLemZqzQOegLdEhyw5t1zNqfYMypK6QZBhGjy8FK1lhfzU1m2
9uN8Lsq2e4APG2yh90uLsLNSzlL1LK9/DeFByMy3+GRYhHGezfvhHr//z4Dnsg4J
P9TXSPX9eHzeFg6u/QvFfRCshYR3VR6MBaJvmHVbwDxDikoK/oy7a7quLRqPdHxO
FaojNHblqRIH6ZaNLZvkY5Lk6zn07WI/ekRL5VQje6TI2j8UK8aJ7k98zmnkoBnS
G/Lv0YiUdmrFcj0zYRZcyoqrC6f41/YcyXzEEMuIUZ8GCESM17tjlaafPy26E1K5
Awp0uQdlyLUjvpeoPdA+36785lXemG/ZGH9E+TWjK8dwjhOpjf7lP4c4Ogy8jGQ1
P9Vr6oJKkDN2NinBvR46HuJIEPW//WLXNmj29LyqeSPS6TbzlOFY8AKVgD21G03v
w/DjEuZ1Gjhz54Nv/xzdsu1hD1e7W0qpx7ONNW1r3JVYv8oBSNq/IvSdGFzFhNcH
Tdv7uaII4Pg18IXMMLX6jRDcinGxUTtW3CaJm7trS6jEXeRKYqk1xY3s4RwseZfo
2ui9oNQWnBPhA9iDRnhwny5gIAiDthunnJ3/tuUa7HrSrz6R1lOeVWPH5CoURysy
YcYgQy3yK4vUpXIMs+ep76jcA8cgnDTUsmw67gA9EW6hLjgwkZTL8MZXu5m46uVk
uOqvlnNAD2+zc23EbnczbkQXLMtAVZnw0kFXgaNYlcIun6Hh8+IaCd6piOH+LA5r
bVzoaP6qPFFVZXKUWMle3HaBqXjNbj27NcDjIhLMQemag3oGTq1FfS0G+FBRE+OE
7aNgQ0qbtd6hrTPiKWoN4lyUrr2RON9ot2OG00TGDLJmdbCcKrAlloSDnnwPJE2V
5m+dsie9K8OKU2y1SAXoWhMuu00lBBCngAnmiFOn/QiFWvTR58O50eik5tv3Xa1J
uWIkJdNfw+JPGhakn7Oxml4lhFPLoTWMfZHzin7AIQWmR0aHni/UiZ00LBducgSL
dKVEo7OuziIe2cAqpI/f1RzXfYaZFIBrX/ouZw5G+V4qIzx+GBYKfmScVDOck0KS
ASwN9cAJJ7BRkuJ4Vpi5lkoUTxPoCTutjSeTIDsAKC1RPk0cuID7JnZGlFLA3gYh
S50tbw5VUHzgCwiSAIkO8FhhYiybSPkLCODnPGNqumGI6Lthuj2YWL1SqFfqFC5K
tfgqAUocGDffwiLI2xyyZiZrGnl+mM4h4JmjWqdY4vbWwgIh+xKU4sYulSgHmPgx
X2yEIVHDSErfO4OHnvTGp3vSah55fnigShp5iG4G5ebmIoUmf5cGBtyKHIBEUzFU
IBNdbFhUQ8jpNg4YGsZ2uOC5ljFM3ee16YxxWsj95mqV+QSK7qj/LlS7kCMWhmjS
8PXwKtU1xJFmk7e6H1W67lWdKaevlIgApZm6YiCnTiB50cMhDQv472k4rq7LwIxP
IUVIcGjqPb1njXlGamz8Oc3fav1WIq6YFLVeJIV9CY0QArnUbpxm0L+BejtmJap4
4furPljb8/SlG6gFj/KqB6YlV0EAWREGQS2fp+vdvE14Mw+oJEHUOI7rQR/x8kt+
F/SLHW1IbWn5S9P612DpFSV3fin1d2ly752zL1hB3/CTaqdUGJCCe0daf5Ln+g3I
PC88xd9nEYO7/VmlAR/SodTmfq+R4f9qfyQRyq4qdNWd1W3cbh9WIXUDEexkSxBl
bw+uMVyJoqlAqpUWW+F0LUJlgfLDFy1Or3YWat8h5ma4x+bn4U8TcHwnXZPCBcEy
b5rcFCp6Bu4lqlo18Mdq1eftnQGGQ45KZyznYYOXdG9MRkwe7CCfYDoosvtVyCeT
2oXwCACPmyfx+SVRI0dpAzypGBUEeHNechGi6JyzhCdMI7Rqlp14pyeGyzI/fZbU
hGbONxufMToDH7PR1ylpqgoLZB955tUJxQ9+T4iWinfUEKH0ydtIBCM27R2wWYa0
KJN6zECaZbsJN9qsfFBylGkOqipMj6B4xp52o4BIaKpKFDm6QdiR1ELmupaeWPtx
LZ0ryD0i9/XyXa8e2XwFXMkTsErn5xicDfZqOjR6a5ulPgDODJMMzzQVNZND4k3l
/IuvjIhjqegPNzM03dboouOBZYZ6RslNCjV3c0O53IDv/eO7Xm4Ta4r76pXo2eB2
jamv/tM7Na/qtxzH6szOQiI5j9+6+RUIKhb5a2M7HzIiDDHghvC5BVXxNiJFaVsL
E0ojco/ZxKUXqVw1Urbz/FprrwRpqcLGL24Iakqp/AWSk+cP1uhnV0UZLoquyb/d
MKfYoSoK8ole9TrIEUIhgHh7iGzwS6nIkyINwCoxeEO1jAsEmZOmIXWJYYvDa4vn
kARP6zYDo/iUGfnC0qL77U31sIN+3OHP8BSBisXBHyYe7OH0/n/ZQZH0z2Fx2mgI
JWqQLN1UXZvHl3ChTW6xPSbxmJa7gUIbWXI/JNpWzdgXDuYym0Y3NYARPl6mC4vW
cf84Od7wGp+4iRUoOGGYt0jN6g2lAnjzDY/wV+ANXuIWuY+ccSpiKeVVv/qo2o98
smz+oTaLm0qVtX23Co8W/OLCac2HpXetnlbolZcDW0FOPK6mKVmUuH0793CehFX+
Tbq9b333ZPfb4CpVeJ4iT+nzIL2LqRd/apkgqFTypoGy/VDPrmsRYX9qpMF5Zm/7
yk5Kfqu0RN10+UWDPw5Dy4a7kL2Ejy7R56n+FSJI5W7nKYfFHc2dguaVGU1iezUm
wilbX5QsE76nIvMCpD7wKbY1Daj43xWiOlqqSQvXfzvkMklEuUVkuTjJdI6D55if
qAN4WgMJzY5JqyxXNolVrp+KwUFFek2ftPRfWgBHdu/vnCNKThCjIh95Z+Gt/a/l
77IzRowWjZKh2zcO3UdXu2Fj7alDOmjCv7ibm8pLdkXeDE+klk6GraV2DnpiMcxY
Tc8b06l5ICw0Sl0EZAuBx/BLSofIG08maqfrN+A7xsts7hSljM/1fFUnDuOO+juc
+aheFchaWo0Z1XHizigD29iA4//wxWt7WlOGUAgr3kqU2RpSABqhpjc2/S1Hfts/
m4yGuymrJB4b0K+RKeXuCn52sVLQc1q1/QYWn3HNohVR13s2CiRJVTOFJgXmwy3k
Iep7ohDJgQc+6aY3eIAXbhvgE8gywVIvNreC41XBSsg2EG9XfdskuHHBP9QySD0V
fuB1wa/JtNDjsWIqY9rs0EP2Bcb8rSrQnKsLvfsIO6W9IjT7CkGSlhtmDLKVJJTX
Lnr4WhN2ODeXdOhqQv+h8c+qNQ83PEVGQgeZOE04TDf2Qz2kmibIXT6RuxZ7B+/W
62o+qPra9zilOZwYDKGeIT40GWHasMLRcVCw5Nx23xvvn617lp1Q/dSBeL3aqLSL
jCEe/JErhrG1UQvKGC4Okkv3llONj9/zi7D7N4iOoNBEMbur9b1C+kpYKlSsfdYN
tuIFyr1lmLlYGug7OGjH6ryDiq1pGl1YMtvz/1Vu34glYxXsTlhp9UkTMc8bjoCi
jvsZcnTJeMq9BXA/bOvrrcrawCqGGtgJeovEU47/inEdtVI1zqE09+NtuzCcbpyN
CDFAtDndWtyJQSLl48X+5Oevo9Gv2RfGLxS7+IyeaF9Pum+GD8e0c7DdCkygChBm
LuVt8Hj2gfrxSXt8wHyT75iWZZhreaqrKgGr5eIsOjn6b2q3zAuMFx//oqfZ+zpz
aHudtOie5StntCcNQXGeY24cRySc5lo8hVRKZbjKUjXFCI+pDqU10QvWh9z8190s
uPdueMYIz4ET/HYPxWg/0eVg+P+YEQj+07vZ84KOMBLb6t6/UEVFIDeJlJaPUVng
r91TcFWNYUiL0TUxBzUgSMmmWh98Vs2sj366zSkBvcf/VczpJRbxHZWjRNyXt0a8
ZuDtAxHL90H8YcvvNwrrAus328SvawGIZ2I+I3q2sGU6TPzq3dVtf0J0Hels+pRr
HtxlMyfRrL4gmte5yEgoHjPIDokSrbjWDetnEcpj1Mza1nBP7njX81Vra/zfxsjR
mGbbxFRZyYWrLzwVKFbtYabbgSBgewYneCefx8WXWaYXx/OthoEm7i5qTYJBcU87
K0TenAgBZ2gCZ5AqdYXcZeI1Mncvz/Gb0HaxDZmA6/iol0rNdjVRj3dDemmPzcHh
gqiijg7yk3f0cRf1fPbmlIL0HdVcdMtQPQgScfE/IPp6XeaB/F47gDp94MgqUMJ+
Gy2zvccDYYn0Hln2huEdOcMOuuq6qVQNTZW1HaDtmR3ZAFcL8+lXuzkLbC8nszuQ
yVaJRUuno0e688rCCepYNqKOpx5HWqaQEgTAPUsjHHAH94RTw/o8m2FrTmu0a4s3
ZSADBuRFckqTdzid0spm8QhHTAFGGAGgMRSYewMmDRvMgjFm1SeO9mFzCqSfeBEF
u8DrFpAnsv5+4TJu1vhBOmkrb1Lx3D1SmIhI5WnBZcs1UgsN5rRM5cIaZlniJQed
lRSyXKWO9h5opPE1Z8bFFV7Mkvjjv3j4jfNqC9+LuMTN+JhZoCfkrUykS/3lR+tw
O+Xo8+5mTCNle4fwqtJfDRIlPAIqFQefyG6mok3YqPakFBQIVKE30CmBu8IEnd08
r5maGozxHQ0nBn8TZ1a6ZnsjKNowuJCZfLr6UaO9rULuF0XQdCWsf5kGR1iVvLIp
tbPm9pSKSDMO1rOaPkLdCpE4RS/mEot2shYTuTAUy6xk84WOAXG6T8K3Tsz92Itr
x4ifMej8J8aelSFY77IMT4UYU8S5AmtmjBmbNg0IICkpypxJJo+naoLoQKEKe14E
K3doIZjC9tt8oB1VV4Y3D2V6+uFJ+Z/OQWgOkHIX2NoTzTcraLoamWejRcuR6zMA
Ypw1PoRXLci/qcW1z9GP84ywu68uim9pRv2YV6zFPzvE/Q8fa6N6IokZnOzK6gGO
xtg4aphIe4nbw5JdD3UqX5+neUNjHjUpUWLhEtexRkeWB2OW0wk/u0ksuuv10Gkm
0jjq7bxV7BEfNpFwTuRMNfg7WzGIsSiNkp7g9wIUN4fD7SEqGD2itqHteaqFhRl9
rShACSvnJbW4G5u6I+TUMe+TQ+o2WiBlXfoGq8qX1k0vduUIGq2Bn1vuGxFhMYCC
DHJtcAP1u/rHGozPg2DeslH00O+S8QVfYqWWuui0TuduueiweiY1Pi33Tey6i5pK
gfpwXWssg+rqqhZVcyPiU1Y+VTuFak6ZwmLwIbyA2PRI7DaPSLON5T6xxE6XX5pX
6pLvaqcwBD6ZWa28523g1nsCaYJEQlLNqj+e0gLtk4bLtQU41daupcre64GuEo7m
3YtrGxE0ZdcFXbKzOkXPus9wKURZqAjiIewoxYTa+xEULBvtWcDSJWXjlFNZCmrV
65DAnsK6ZoraYM1VWLNgANtyu56P165J08ZKF5cjJQIh6SD8Vcu/bvkDhFf4aXiD
iC+7fhV320/cODhZph7XEAximapYpQCuZ+eHp1WumB3g1ysFKRwy6CfKsoDKz1Gv
8y0q2I8JKJAxdKoW+kgQNkwcE5U5O7uLTWsMNhxOCX06iBi7nfj0wI8b4I6G0cV3
q5OMuezyT9eNIjrqpo92dDss1geCj3CC5T71uid+OFLPkbWghXoOb6eV72EZZ82d
edfN97vpASsOWZaVtCHRBBchXqtTNvpH6WOOGQjDfpRStmHfFwWX77gE3q3IfZOY
WfrtMgcnNnCzqPTuTNEJy97kVm5eY1TcAWbETtM3o96Pg18/5RVfISsILk+VyL8m
6+6MaD/81n9k3Jpy9thz7D61E92WFhWnnG7kxhpmKB9G2slgpuzAoZ3EY42tOm5y
NpZ+alkMOFAdy/kF6sYAB1yhgr7fqdnABGDq/gPdOU9EBZkl798Z/raxW/3O1cFI
ECBw7cVF78ACUr+d0BvyasYNS0fsUKDmdN4mOTUCRG3W2g/YsdV5Cha26+5QDhSf
4ztGA/i7qNuu5HjbIPW83/bfEmIYRIq30/yD5sCSDeIORv7gz5OPT8CcPNrZynuJ
VZmy1MfFyxWwK5TAVCJMtT7xevPwoMqRYCwzA5bYPs8tnegrIFy95ttfbRmQPhpE
eGaY+m9diX3uxR8TSxd0Zeb1ZcGWTEMWXWcx4foW/w3mrJ4Ax0VC9vrXHu8N4grz
lxiuoBtvV3H/sgkuM4DcYDFKOY+SIL1Vd/NsbCxlZqVstwPKlkJsk/AKTTjzAXcs
V1GJpaaCzL7/VzsFkPTF6s+1/bqDL+6wtVdJi6poXistfJBGG1vqaoTVxpE169hl
fj1NqDKCqIYtfqQKeORvfihO5Opo1X8NMStP2OkDb6ZcDpjonYNvM3YY7vYkahIw
0n16M5ibhmhaFotab2fvJKOSLddSAo6L9gN7+vxQoRlo2o2qy7aQKqKdQ+P7ZCMk
LoOOERzfX3oh2on2pnQxUdDPeVJlmb2VpO8Il9Zf0PhtLzt3Fm1seXuMQ3ZeSKXy
MfKq7Z4ohfy/2BPkGO+p+HjU/EjNXm3pwz3Y79pI4lK+ixgtCDbXUDhnVgn8hZBM
2oV/2Cn6wYuLIS63fXluGyeD/1r70CoROix8aCde239v6A5rlwaUxB1qCiEl73dG
OmSmPoZOs3tvPthtoZHuAwrlHXTA5aUQmg20HwOurIcgDQ2a2wYyoNkInabDm/l4
sOxoJBdAcmNoDLsrp/hiDwLnhueM0wkvOcncdDlepiHm7tO2VQ0L0aHXbdKC7NBM
IS5K76HBQ2YNgRkrVplaOepJo6UkkCTr5XUUdKHxczZciSGgU4UJ+x3wWy1/Th7R
gzhccEOkdCnk8YEWmeEQNQ62ryd9y7cbUmxdYNsP3Qt22PRdUXHiQPqnGAtH3J6x
1I9Ir94Y7ZwVtvNjRQOnLnJAOEFl9SIGwXv9+nd77Y8eefX9RnobFR8G4CI+Rjfn
aGJph8N3a4AGSi1INiPAkv4R0om5s3YGf+OXsbEavmqluFFevZvsz9ZBVbwTaU9/
WmtA6zZcCGp0XTSSt7mM4srDbSSRTrQoBgHVHTplpsGsXJDF4lqpDZOkl1RKMngs
ZBFF8S+RJc9FqYbS5zfMtvRaH3v0HawanbLxKToYf0lbwmj6FMHCKJ4Wf/pdD43U
3kEX68Q++bszMxLZf1XX09OR8oHSrfQeMAQa+zGF+dUV+kc+BshVqa1oG+7ha8Gi
X2FN3T2OMV5gBTroXMQfFBh6khIhWEoGUcL062/btfcyLxB14abf8UGGF14zV5MZ
8uAvLUGX1Ij/+rJJE2l9D4milCbSXrDhc+nE+/daGZjOvM3c0lbv17G+D4w8VRk4
zoHqZuA+Xa8trEDKSojMOjXffUFVFE/cgbQ9UrXbvWPtld/d18g357WnkkgoYeGU
AJVdUCVL7Ew7NRXiZSjg6cIWpkdwnZJQN1LCt3liCgvvHVFr5wpLlnmTdh52N/W0
M4oEN/0Y6/6AiwqH/CNIWkKUIGodkeDjcyYADCEbPQC7HOx9Wwk9ufEAumqh2uEj
HG+mnwu3qt7Gyv1PEA2l2o1bRJkS8mvsGAk4IyB5XUJvHoGU/xAa2hPA7LqDVai1
23DTqnaC48AgZNCSgrhEdvvlVs06d+PxFla3+eTa8tBY7snF9z7o6Gu84uzO5X0v
XilvauekLWiNA6fDtklMaAOO9OVKQ3YGj08o/vzEzQtoFamreJ2dEi9XPlDIFFox
1JetlqnXxLCT55MkjGuxsPVtoUNz+nSwNfghTFmV2EhzqfjGilT8mY1DQCK4jssk
QarWU80mpYIPBf+8xIcl9Tff+jV4qfFF2+k6ypntBl4bqrNPqupncENE4Md7hENy
cRE80sgF3dvcxuFWQq1q8eX1zrdxqpFWIY/vadhVrXkRvpmpcbvJnEWJUn9rOgza
lWWgiZbi4CPtu/J3Lvz7e7m06puXCab2NIayBw3g0ua6pVW4vDQNKL+H4IqNqMs3
BNX4tiMcrMqjpNun/lEXwGwSjcQ2lPcM5IxxIeMgGQF9hpKt5r9glvONkqAoU/mB
mnL9sb38TBnNHh3lzYqq86VF0ju+i96UmBMrXAiTOI7YLNXSswp0RqJk/tsI5kDD
mQcJF2YeSSL9/gJWzky7P530IP1KLMcpcXfMoy70HNKN1MoCANgJ9f1BTgUOf30e
r5UAEujoiitn5wl2F3b3l6O9cGHckSlOCj1LLKDFM7Pj7ibVPoGr5/Cm7BKcnBEx
eoZoayH04Yu59ko3s7O4Eh0tkgfl37IbskXoZQ10/k2KYxC/lOVDau0cEiM6iamJ
M8i6/ToIxh0UPbctSe6SKYylR81Kbsy34UaBn+C0qu53iDvXfyTvZcUv1uy57qHo
YK7UsFvJDDtkhu5lHze34hgB8/mtxvpgXmOBMzM0Uh8H/jgOuyp0dH5nVj5Nzg+4
zstUpb5cyV28XWMRtgYAY/AX6I94PW4bbsRniCgSKXKWI5MM3AEVcWEL03HP4gsV
HsBtJTqJvu+/6bIeohPNeuxr3l0ubh1az/ozlrkV1AQTEJrY0vG6y58XY/JAmUzy
OYm35HER4lJdXTjnZs41Gs9mqjNl9Co3l3l4HTCcYUfxLLYVHka2hVjgdGEdWylv
0vJExUBBVTLsf1ybp4ZPD1DGtRNuZ98ARJ2uwTjCGuv0/2V3fdue3R0dEjxlutqM
JWyeo/0E5J8cIFc2zDY8dcCAHKn6oo2/bMAfZsKavrTZjCTZ4vOuaJM1ejm9WvXa
A5kHByGZROuK6WuBEzpxivzN01J0jhLp8SAipDFanrKAYBOvC/SJeWs+NsTVg4Lf
cqPNugZgzkLn8iBvoIjYnqWq4b8NxLpLDkTQ3oP8AOYPDluiT0zBanTCpMb6EqL4
G1x+lyQgun850YqT8EKJnK6v7onyvuiiSvx1cHcrrIkb1EyZTVoyHPOMYRtz/Jgj
vWLQ3CLfh1QUecSfrFPEk5UHxbV+Ul2BTQfbW2VSLp/Ci0TWAm+DumJaMdPt6f3i
OnM4vbYhxSw6oJeD9A0PsQRsj4ATfff5v0UEhi4B4hjHcurXvWjxe9S39L0kF+jd
GyA1GIJsmbh9PaPLdZHjW6TyGyNv67vVrO0KlKsBlOuW9ZGO7kNXKNBPKHwCOeAC
NRHI+UjK1JVzZCjYNcOLPgezkoKP+/xqrRnIwSgcQ9zkRlcath2TEO9UPKJorUUk
MxMID0wKEd2F5iPM69Ln8X0tBNxJP/gB+tpfZq0iHLNFow37QA9FbAyKzFgLSKgq
b9+384oHxmETTBigcTMcmlnkGYZC63rco/mxmuk6QpWSN9Tf//BTu40rnF7FpGSs
J8TkO5fOiGDfzXGVgCVj58GPt0JEfo0ukAHdCT2hbHP4+56rOA3ykwf3y6wqZ2xO
k0Uwqus1eJu76nmS87Q/qlC9GmaT+Io2Djko9K3k47URyrk08rpeORyXz9FDKw9k
DTMrQWCgRZb64eN3Mnu8NAJjrAo0WZwZtFmnDVJ9jT8dcC9VaF3CLXvcV4Nrg/5v
upLCAjwQkd3DJWWQy+4Pmqw7NZ+c5YBfAZuwxLcB0dsA9kRL8gy/O/KJZXe7EIgP
XrMr5d7Kt0t/7DwH+LAVZdrISKt4ELPqzHx27qE/DqxFl0qXqI073E222Qd95z7k
l2J6W+fUURG+kx1AFUqdz6Al4DfLBbwKlCOuP7IKhx2WXDsWHLzTlnZz9SWe6BWi
jUzqZevNw/Z31SbKBPx1FGDbOOzWY44OcJva7hxs8ASir+a3w/bM6xWS0ZAQcWG7
YuQakbDYD3TXZaA9HTLFtVkT22QMIFf3YjIpLL/Ff3nq5GlB8Yl5lb6VxYXE8QFM
aiH5WV92A+gy4vZCoVpNzO+t2QlhKOi8kOq6rZyblsjiowujkbBnJXRoVMm5W4PL
nThaiXGg1c5CSivMG/iNJ5TlzuggY3gdkky228aGw1/gRKD/VaV5FLu9Emmc6Pdx
+fupaoi2sNdabeK2r9kszLUXEkGpb7Y3WWvZ/Dd+sn2Fbad2uJqBpGR1O4Ro4wiI
OTPnLNSgV+KmfhRXM6kfMWSqvgTwm32BNGunWSB2ZMGzFfbTZ2tobSnZAHutbK6A
sZjCZkPCz4bhaHk1tfpNvF7R/1j1HYd0UpYPKA7msScwjAClM85VklEPS2PyGONt
jZashXZAtUNWgR96C/+dHCxjyZ8Y1efJZzHsfIIEuTdJn5t7Iz2It9vaVGlKBmRZ
eRdGJPDbU5hc9p9n518sOKXt2cWurSJVuOQuRKM+D7k6NMUbS8iJ7JO56RVhRlU5
GG8m90oDDrW8Mdm7BRPXgFzzRxRuyBp7dqNp8FbMofyMZNds2UCiyP6cG4LzYTy3
t/dv2QJAs0ns60PHeOy/ULxgiTv829jz5Cyka/g1cImGrJRXl9psqbXYD3Sm/t/X
da6W9eRgS1duMexjd58Z9bjb46/HadjNiRdqHie68+V2sFT6qvvaQ9zguFZu3EFi
NMyDuHZiTeAWZ70HCqQtErw5JGWUwX6vGlw+41k4DHL/q4g5e2/uIPf7vkYc0gNg
gF7Ne7HF3WDdEkujAzVaMIgB+onGLFtc+hlHgCLySiO7venP3wqgOJaTtILun0pe
6yDFTJuikW2mnXO/DDc1A5gyBo3jUARbuW80ROvKRBvnEbtCTbq5N9u8SC2vz9/y
DBA6ei7wcBjDb6VZ8fdrslnpvkBxZ2GC//rQ+iuL2uJvkvtJTEOcikyBqbKg+9Gq
wOQOFLwNNsBrKN+TW6LRgUhwz3/pxjkLdoVZ31A3hYj70dCBMBGbu7Tw3SbTYVnP
Js5TjEKPGW7EHjet9s11OnwGsl0ka+syY6PxJHHbrBd7ttua/wuEDhLB/X0aIi9+
DXzoy60BDLauxFi7y77eZRRs6K7coU1dicQh5H5qaCZb+/3F7Mt6GCklWgrwHpw0
XRsN34Q5Xh6rThY0jA/WpQG/4/BTnv0COWnM4ByOWicryY0+MZ0BmBH7TMxmCayZ
6ScR9Gb9LWzHx/+ZfkfchL3Feinxq4usbLRGXuqFE9ygJ+Xjt163aWCkmPqx9sRq
xdu53owENDJlUu9nzLUlCmGV0pDynZlDqkwFSoNlh4wEtSPgIuUrjgHkHmi2DoN6
PH+5tb6bALSiKEhJ6UL6HOmd7+B6tIpCbLtMTFxBxH6Tc1APaZCxHiMIXGX7+0V4
Ym5I8s4Q/a8zRLCy2MeBLirRwGAmJNvLlhSn8tP4YHVfeGWtoFiyO0T+1qRFp1Rl
AVQX/cu/raUGHxRTG35h5joD0trz8JVLkF7jE02sxDyYp2y6/TY6+HjPprl1WR8+
YIEN+Ooq8FhVCp+ZzERYHwVKl1Md5ld8IWsfoKssJpHrUbJUzJGIVXTA2mK9Kcf3
yJGvO9fsj5e7PYs/vPdyUvOMjImO7jbaaoVB+UZ9qz+wtdwHvAY9vUySCQbQ5E3q
D4HBFkJZSdYH97hkoUjKgkRl/7bzbSHoY9qGGWbh8Ytgi4IkSeOBRb2jz1Q4Ca1o
W9sTWJAYnr4zRh1dpxv6HT3v360FKzn+jetCn9dsSORqg74NmgcdBtLykZCIW+5a
wg/OtL/eytNu/n2HRRKxi7qCEqQvhe7JgAm1Czfo+uChATsE1pBxbsQ+8c8RarKa
0HJooegJlvbb8q+b9PzUhCabyMSbTR/7oUNFCAJ88wrp24cUMx8NWFLWWk1EqMKv
cDGdj7+A9tGoonCBDKYYICP/RpsloGkX66k+ltwyMsD+89Nxa6XlICzolrfsKMQH
8fGJZ3rcW2JRt/lHa+USYrMbEa2ZyPSbbxZmNmeGMwLFoUtt6pi5L9p8CWh4D8on
4WnB8IqP+Dl4z07os0768bxAIc6xbfcgCOMBC4pNL9v70AF2fdT+9KAXmea0qPQm
Jqg/A8z9+T4eky9bH4w1jUgZpxu5Q9ZZqT0SQRGuJl2yxy5+U5wN3qRMklCI7BQJ
grbBXoFSllEhgsZ4M2BdGimo+Aknj6+q9Mr3/uWqWu8sd0f/fQAOt3tnpawZ8JGT
QDkpQ1oNBeOLuYwGpqmXGr7ABVNAiWzJg6GHactmanSUVuP23ECZyYZhBu4Rq3RY
DA9cfc+OksSIucHhUmCQSco7dhj2VYtf3FslmeaJj2Qm48LrMSgG2C05n4hqaFtJ
CQRdHKcC3bsttfeOlOujZieGtp5iKThTqo0RSN1rZHyIUCl5FNzyboE7sxXps3sX
3kO4DU5KLL6L2qGsN4gZC0S8PjBKO6PaByDDUsJkKR8sNP3HcFYIem8nxfhzEwWv
E4TmYxWtnCFsspPaRZnwK5s7YOqTfkxxYDZ8f47sMCvmKUc7wTSiTEh3HNYaBQn5
1z1tLIX6zUgZRI7DVGbcaV1dR3pba5WzLmjtcn/6JcxLJj7UYv5KmzBwJogQMo7m
CkkfeCuuQstwg7IcSETwiJNiDz3mSLgKSK3GzjSPWj8Dsu9rMfr5aoT+4fiy2rFT
J10wcGenxJFsIG4Cr55stCQ+wBDs7VGXkg2/0Ky/EsNijLIgGXgb/XfrQNEtiipo
vjlf/votxCZg1snz4dS6rdK2ZBLftXVUZIqHhCxmB/ZCIXVZ35tJgcahIGUnbeud
1Lj6gCVF5hi1LDhnI0cQXngCxco8LNR4LpXHufPeNOkPdJkhCNafKBXff8o9Jy1Z
NB9x/73PxztnDnI1AKnsdmQ0Xx5qXUvHzSgyto191cQi70sLsLDltuooKRsSYLWl
+wYbwRD1wGv5WdKMvKmAg2enimy9u+fjYmncsALFGXeWlEbzNDGrycL+TyrCFWQH
DOlYUHqQ52D4rvu/ZeeGM2AUEzxhuVq0bd8+QewAsjgKpBaHbCmfTKa5aC8T7VMs
FnN3Nx/qow6Gh6cgvbcHGKcggUlZ/cSGGhfXN2eC+5ceC5/QmQVgPk5R66VFix2f
Bw9B5fqeE47Y9NQK+EX03ogU/ovOtRor/WCIEJ+qlO1DWt+Cs0Rd3e6p62QIz5uV
zG2HEo63b+Hbrb3kdtQYiNlmPusKqwheP/7TyNsmP3H9xg9qduiCt/9Kbj5nIetv
d6Loca9QlIuwd0wn5F4PPReuYePnUjF6vh6lOdY0DLfxn7UPJf+Xz3LOZq2j74Sq
fftI6lhxLSc0XAI+z5pwe/4WZz0IjDZmXipXfZcGxq4SbiPJmZTAOk9eYfzS/C/P
KlXvdjXPuSRM8FP0odRb60BIHYc66oy6ccPIaSlWppt0T7WMtp26Mg+oeXpJFweT
lOgIIKOnZxEoDJzpVsNxeuwTUSk4GdMSPdf+vZOrmEy3NFaVP87bti241JcXBU4V
x+5CDupJ+Vucq1OqCuDHVF8LU8NU+Im6wTsa3pa4HkvOprfLrEzvOSGCavHQ0RDk
tLfO5dCJ0ddFfXEoqZO5tcEtCQtUYGDZRkGZg38jKftXOTKpiELOAASCHpTIW4M9
R001UetVgoGYrm56wAMgon5qmJX79gtgWXH9zjZ57V2VrcOLrSBNIhUwctFW7pvr
vSofdwadoqHaevVpEA8ZMbBDThDN4ns8tN45/tH5U2HlhBR+V4A+XJl69jhdofBZ
TWGh7OjU81vABsdqnY3SBWdNkef5mK2ZSRz5DO960d+TjqQ+abHg87yDnbpWAKc2
JCY/NW7BvXgaj6MCHY0gk8huBWg9aBd8C8jJ74aM8eL0wEdISJOEAE/1JG8oTCai
sVe0+aL4AkA+DO/1s+gKsHe7hefG0Q/H59tnP8Q23QhshVu+0/qqXURlG03pr7mz
EQNBm/VUYq0W9cjhqmq9lps19Fy57uVnwOic3plYZwCA+XwApyhgLlQSeliru0WE
YjuGBL27c4932GmXKL5K83UttqdDj8sl2+KM/WrpSvWHdPQYtrCu7emH7St9Nr2C
+UrDebeLGHjIFyrkdkDneHxTYAa0PZLrbTRoiFhAlNwCl/Ubx8edwFUO+8jVoypJ
6JC8sBfX1L0cZZ3Wyw2H51tLuZ0w3wmqI+eHE9DcPQ42D4qL1VeQGDVGxHliSWJA
9PO0uDh7UbR+RH/zrgBqSD8qY+RHjkEvqjky4TeDFuPcacbeNZQkTVSbKItJXs+h
JkUG+F6usx67yMTMN8WnNVh9GFo9yW8qUVlLN03OMrKr3Ozbm6XUtn1XeEbS1Rm4
P03gBtO4uV2CLQEYg4qZTaY/Xdwj/xiW2p0GlOvuO9Ppfe45qwpB+JtmwNRVe84o
b7a1dDb4p9D+PVHsNQFHJ6yiDOSavUu23yZLlYjHF8KgTuJHgHVu8H/QF6gzjaCE
LEzIaSfrSy4TXpF5RhezwD1EkhatUmidoWok7A1cMMe6Fxudu4Ev1efbTdRwUv1o
gEkBmPa8S+SHuoougM5LIpGRNZREcX3iP0S/VyI7DmldUhdRESxS49nzZh93dTIX
UYH63PNSn24yDZt8rg7TLJJmdFOBERw9KeGr/QdUMLqAAZI3bsvnZVLW4UkMqP0Y
PI58Yd8pdx/2IeQXbUxop7h2JD6HLkYaGrUEif8ivRQ7UoNn62c6AZWhW3f0BIxf
NNv1Hco1DuLqeCmBGycOJLG2UIfca74FCBSxw+/DTe+Wo1flnh1+h/hBCSn/EhDl
BNEAOdaQB4Z3NvwfptfLQ9IjybPp7j9n48pwSuh4ZGox/+q+hDliQHnEo4AsaQTc
tNgOHPsIg9lM4cuPruN0zNpB6hEmTpHI5gojAaY6TSC+NR+nTJ3fhhS6WKPwONud
B7EepD88qNriaQv7fnAfqxnZPIrWR8VAcpz1kCCPBuILsKWBmokWdWF8qmHFpjoo
PqEvzme4wUp/iZ/Jv2jtduTinWQZvIC1xi0kNtAKUTTgkpQtqXECw2KWj33bHGB1
Od0rNTi5f2YbjXn4aRGOH0NkFrxyXJNW7D06JBjVqtE6UNuyPm/xz3nwaZ3gLXdk
/VSkHgDC7nuj7YVjgzB8zKN6+IGFTYoBo/z4+mW3eT/zGZ+VFk6d3CEKs3HIDeBx
KLsY0fFbPCr30X1O9o677USYP8kXfr+iEXT6qSyB057HTtBdFKWgMccXmgnMzGR8
9+uSuykfb60fMLYhJvFnHdu6tZ6zpxJnk0QkJ9+IXksCqxakEBUt1NgAB4dmme5F
jcErV9UHTBVoR5GLGmbGd+HAIgdFUHTCG5RyDk4e2gZFUiz7rtrMuePpg/KOZcBE
TpVpYcY4xTQPNDCTj0Isl6K3tZj5s3KCEv+26MmaaX0K7DndbWgbBDK3tcs++MBN
Nw1HVTw5UAsneL1OA2idMF+NpSoUtnfQ7yP0thG9262x6NOboQFCQBS7pXnma+rS
ihnLqPt7KSn9AgRoLIbjEZuOKJZ9CgO3ly2yGtn8dJdBXMTSfnsd0K9C/IdDgwmj
ilJQln+YK14COYyvdZlil4bvHvwCyjfT1I4PvGjjqt4O2ovtmGMnzAPHBwHHrnV2
uR/mfP1t9WINMQ1/QDHMHZOZnIl7RMTaDeKnkmra2TM7tzDm/LdYO7A0E+xk5EPW
oy/tR3zsvchaQzmnuvLpjg0RCfVveq2hpd6G2Xkh3hk7MLWEJ3b+w0NdWvXofiSG
LRAzrvUlRa0gcnmts7wSVKeIjrD4/ygfO50GSwcOUonFWwafeo8lxClow5Ld/AJE
Mm+0eDdMrr1qLWTpiIrkkb9TeiLcii20FGQui207/8x+9A1Avt5nwAJi3QhKa+O/
Im0duj9OQCgFHuiEbCnyHZsRXnsrIxqHjXQgRTrlRBfJ0JCmQq1ZDXVdk6UhgUpN
0mrrm9MOR11CGvBtzcTivt1ynCw6CYMCtRlFWpPmIqy4ifWRJXbinZHrI9FLdkZ3
LIzj4xwMXjN2OZTlxcR6U4Qt+FAJyg5NL4h/p1n1TfuvTUMWNjebM0XhEf9tRLe2
0A9Z1AEH+LDEuVTjGrWuQ4gzOeDGBs6dgFr0/CsB34SFtSuzc3/ow+HqrflK/P4T
GH4IMMwU24XLRqLsKiDJFUXpuD2azKtlEdPSDJOnEthrGAaJpTC8MtiwRmFbQdRW
dpUMxrj2sYcgAQsexEqNxDY2TONELzlbhVN61yLrBKmrz36mgVYYgaxoyim8hKJq
KM6vGx3v0T+ZRHEjhd27wCizO01GQMS4AnCEypAjEwoX5W9IieaqbzQpj2o2N/qD
I16aTc2XawYt/Hbq2JFFYHXANz7k0TPZ/ig37gJOZ880SlNLpudfVRpusozCxBpX
MSTzzdnIqHx8dU0wbrwrnB9wTTCB6km8UN1qWiSkcm13IAiL36TVOsOfiPd47jrC
9x3hk0GrA6f142vNB9WS47BkZ3b88hL3SqjvV8FIQhfGUvlyZFoIFm8wLjhEDp7J
t5u53qDmntDwMquen7+yylXSyAXdek7iQGJCHBnUBhJ1LBO1+D0AwhNooPXGQmpd
y3ce6PBZ9Y4d/aD56io91PYBNepDgqWa8wgUPnAoJJZ8R8hkETAYrNfo8N3l9XDa
THL3rhIprWpn839YCwjZdBK0cPTvZsUWrpz6wjmE1iSyE9DT/Lony8Mg+mshuNFl
BgYHH4/7QkweNhLRErAMhp490v2wgyzbs8PHv+wuDHm4XaRnVhsbQ00Emd7xN9UN
9EYIpVKi1aQwPniCdZHov3tvik8D6KYFrfp/g06HY5shkCxp57oQqh/BEaMRuPvk
7Is9lVwn1LevcbxCLD9bKk5y4P79qgkBAx2CevPVYeDVVeX8VmCgKsBga8ArSFRC
dtvYhGLXBkS8n8lkhchJ/1NbDS+sPYqIfP8LqVlTLQH5NqaK9mRh7rYhIFVdsJFn
6++EsY2WePxAV2lurmeGDvCQVu6f3+TD9LKBrMARsy0whhQGhQ7L6w21oiGtgB4r
YCzFYWaWzzv9/blRWprmIIIspf1vDLe3JxKWEVuejWiyGX4bl4CI6Eabg9aWvZhn
9mos5cN2OaKMkU+lbRDkpbGWMosSfUrPpdyI+eXDaz1yhCQ0LzqgB8bSoA/IJcZI
Qzcd2HGwRyqk4eH656MiFXB7+w6QbqRqTYDWE1nF/srnzTAS+kF24I6eQ7SOArSq
znALybh9kByWZuAgH4bHQEOtliPz3rX9dsfVX+DKV8aYKCw0XzwhHRJQgRRCwU5k
sMGTYImJCqcmmDnOMvusW6CLNAiRrLcNkta9QsXmuZroxtRf/EoFUDD8pW7nIgaL
+HRt+ya9BEQjl/hEhWO0JSc34W0gwYf8v6/ol23biz2YzUrfWLTGgcUafDecgd1U
99g0mQK2WRe65DidN0GT107lJQEXs3FcLowuIJjZji3KeHZNbEn5ALcSa/OOBks5
acH+h+rzKnqdXKkOVxhgnZcfpANzndEOBQb7nE5gP+Ing7f1X8gw5FAcsHmM1ErW
XCers7bd5i/Z3vNZ01+0MTo77x3KX7bZqOA12HFlznw+s9b5NXqRgAKxccy6MIVS
uEb0GXzbeQrUfKNnXksdt8r/mQMnuYVmq5vGn7j8V+twPM4jfYvfcDUpOV0mtGmB
NndqJmRSHjeYWN+lMXyhlcjdXFcINSdPgwmY/ulaE4YnSsbfvbssfAaN0tCqikwb
Kz9WuCDevGsPPv1cwuoXl0WKbNxnYzbqJEeyDY95AYNUt3ncwwOU3CIbtbmUrsJz
jdOpcdgrAsvlIhbtZPEfD25Z4f4U16LYf8M/UVfT5eaIHzjyzRrACUpH43sy7dVi
hFiFgzdx2kcF8NYdQm0lROr+j1vJRYcZhcYZydWy8NK79fiEJhYBSPrPPQf0ObCO
dLAeEUYWhEAirNVB7vc40qXG/7AJ76NhDH1lR/MfCnSG2FvoHcp1SemVj1m1Fm4I
wvQ/+1ts5BNfvjV55ZWpNGTv2zw3URTJg7RBjKqWjlMKq3h/S0YvyiZQbQEAlJX3
K8mytj9NaBJhnDZy5fT//+KxdWxON2XnqHnDyni3j/Nh4CkXAoi3jZmCsrB2bNGZ
hMnW5VoDKma8FNHCwdak/SyJrzE9ui5uC84nyCy4Ahz+WrIiYexL9iajdNC9ebtW
9+OF+Sgs9LvZTjgIs7iRdXWBF1gLAG5XUWiU+tLeRrauAfMBsyER3hY6uw8gi7jP
W/IKh5KRGuJGPkopVmBoOanuN9Agt4nCP77N+qjPMyC36eBdnita1r7oyZuNtztT
7NsvUWQJ3Vtax2ZpW9O6QWVmSZ7IBRZnVG9tfCdycD5yeynTFlcvk8A8Nv5mduKj
7Wm2aKiQ/SJrow/ASdfWhyJ1sA1FviwEg0LegS2N6ejRStEejv+i2NlmEjivv8u1
0pWi/+ExR5cmrngd2iqwrRHneDpsJjKRu3BAzfobDbBmBF615MxH2CHFZcOX/eQV
Le2wguQi9D8KobzkEgGankbFLjIx5Df55Q4rp+I8bUMCp2iycJdX91e11qRrc30l
dqBamp37dF/aAz7Ppf2hX/Ii7OPdbc9anhdgrKlJ7FoCXfRl8EPmr4NEpXujOfGG
MbqYzFeI0il8IjBc2rsj5S7RyA0sDuVG0L+Qk8KYxOMH+XqcGRxjYQuDAlgiRv3p
ATY/Ek2O0+BIj9e4KvRwa4eOEaf1ktiJQkZtq8ZUgPuhZxoOS2cpPziOIsLubyXb
02kaSgpSLsCgwrOfKwdmeCfXk8ttTDOT9LmycSRkRZyxUmmvHHh56gkXWO0XZFcY
90H6zUVhwe96GjIWFwQIifphzX+lFlz6v0g4etikyFDDR5F7eSZLwqsNs0zsu7eh
FJDHTNXwGdHcCroIdVQmw6n2k4oEgew2tDiSC4fc6SzW9nAGv4hTGtqksX7+x6gz
NZKIOfOnu18vJbcFYHxC/xgNbBfdxF8hmDjjlwjVQEuAp6THaVWYh+Oe2qjqkRSx
m+8+9YutTCQUt7VwEz+Ct8UFMMSK0esn12rCqaQFNXWTK+RUD1BLcioEiKMcilnO
DhTSdMRuyzCQrqH1TqHmIh5ptl2zyHrrVJIS4w+1QPnztv7C1mqEWwkef/yfzuf9
A1hU0SXvjfygCnlq7SL9sfQHJRQfjBa4orWqYgn1fIlbi+Jt/fJku8ObK9kmd4wx
JZhfI3JEQKP88wiJK5I13vD+Z+XHMr+R5akgBOuhMJDBXjp2WXPc1fGneB1Rgyzh
fujf6Y2rD61XYjh95Bj5dANC4+p+ZRaDNRsARXPs/WJOsEw2gMu4g24FzApV2wgR
1P87nUPNMn83/03TexDpzvXUvRlzUkNZXloL56GeJz1raXEUDbqAdBV2mbsw5I4a
yDuY2s5BcwS5n5aR1LwOoo2YlHAGwt4KHIH4kUSOE4u5M6vqmkkDMXcHKTLhj/gi
y6cw1dJLn6+eZOjvZmCpCPkpc+4rDjOX/b1NtBEpzsY9n6TWGvtlI5srz1qlY6Ek
wXpL79D9NNAzZ5wVDiN4jSD/EoDh32Mpkzp4bjRjsTA29OcIwMypB+vTtRypnJcd
AauQOFO5gybO3QcUyy8cjzVNGb/hGruFuPQ+GuShegs+clG4mUJfoPZZCJ4eKQYi
3hJ/o6V45LjPdyERvaNc4nNYgGZ+wI3XYGc+QZkpfvHMnB/uufxBe8Efuo0J8MpS
qLuVS2UsiJChsFxcasYUzV6Oy9sManjc/8feIsD2xQP+c0HqWeQRVkKKXwCZwizf
HXgVT80TW0dTEw9OdqBBIojASm31M0H74T7wHrunX/CxIBGc7J7YkXSTO6Cm1i7v
li72vqOYxTriQqm4ipls9FPnhXtAoFBDEspKJUMdKB1/l2JEqDmM1TbBq5VUDhzT
tb5krPUkoRpdfSd2jw5XMJP4WEvHP/K5IhdQdfRmcqc9FHQdiVofbmTabT5JC03R
7Qs2NIbfvoDEblJbPRFBv2bqCPkDhHnv+CK0pRtG6+aeBVh4mFOIH7qviUTOyNPQ
ZdMc8spIhDaA9/iAQYZysDf1WmL9VGfAl+6dA7Zlcdn2hl2AD5MygJ8IczTRoWOk
cjEvDEMIwdpPGnyFXL28dnAGeuzp4coeBlCojJuh2D3ONO03mNlJzCINSPmIMlcM
W0eelghw2wWl1O0EEv8SzMXA+Ca96Jmjy6wLfrLxKadEA9dvK85r5SB0WF0c6vR8
URI/DHy0YF/NqNItJBZPgWhEekD4TMVSqb2qxjjQBfkjPtL+tjOzJD76RV5chyZm
ZL+XhzuIVcvS/MLJP5R7ImAd50Uh8MLkn4soBPgUf96bLq6p2ZVXsM5AcWu2Ss5H
pEjFfh974bka0GqjrOcUnrox+4+UG5MuiC8STeEots7ILemVgVg039Jju5nu5C+z
G22qwUiKS0yprV5Mlwk7+DM7JLkeLDD5dgMs2HE1FHfmGAdIxjkKxg3HEXYpEZhG
Ri7eGhqsWlJQcfkRGdhGdGAtYqfyFnIuQWk28K2smsoeNPxBHPYA8HkAry+275dJ
DQzMtiIICjz4ScOexT1Y5FXmVSiWP6vgGs0D/wun+O90r0WA9GngJGzQfhQoZew4
JwBFqvOkSnSL62zZN+Bi7Z5usfG53AYfGTdsZoRGTvlOPlx9KKgBRFVx73LDGFn5
MDY2mZT/SD+ge7XMKivd6Vn/FnqbXr2WbOBiqWI8JU5e+ijZ42fA/tQ7NLVtf4Ed
4QzWq66ZQ4r1EFF0lMlWk8yjofc6I3Fq91j78m0kG3VtBxihYGViOZIdwkcwlm9e
Bba6SipfgvtdEmyM3Bc1OxgWodvw4Mw6Z6V8Zb+xsrmf0N6q9dA0lrtuFVMQVhXZ
3HhnBUXQPj6W93PdwYIz6/RW3rOTtMiJZNRznCxuPES2p5S6/e/6cofqrFuWGllm
RMMAWvVjUD9T8ZlerSZ8pNb55lH8U8NKWD0PbGXMXR0GOUILVd6dP+hpiBQ19msv
o4h60miMuqc/tieuvYTJkCCh3DF+b3+HU3HXjBNoQk8g13C7GszOQ8uZfzpUc5Ch
oqUvit6qmiPOCqdvn5uiuXtmOout5KYJUQWkB1bivTC6nlSdVdP6sO5v7/AyL8vF
zkHjv+DbW/9JhtNaM2/PtKajvhj9uyVNrO1jOLyBVQZPqiTEVzCznF/328v4PWHB
KId+rAZT55z900O+++FSGFJSL1vSiTWgSi9alp0e0V2aekq8qm93Wl3wO216B9uy
AtmeAQa56HmfLt7CE4sCYOQNjlHLBrz/p12VfRx3eaug8PbhIN827gxBKGlym7jR
ElASg0SebPeun8U5h9IRSSOMdQEEUXbcOxIRsOZS0vBvlCuxKphBwU6hwtNcsL5u
3ZE6qer1GFvIntIjU776HeyaRS1Zz7EolH68eaIsXAfWfj5ZRqRPomMFbiJcrWOu
LCMidHDyQ1QdYbc89UP4qWddr6t3/ZbCyUL3ZWt70/Y7ZhBVStHCo6Zhf4jL7PiG
vfOLfzvHL4ZdsTPuZBzA2DztQCCe7VwBbHrUsdZLpxxYotZ6t4hps0V8bUsZ1lwo
o4kMoTZGBgbMhjLKyiNOTysADFIeF9xNG1P9uqBqX0r7EQtA9lS+i5HTIx/XspI6
lPThFuAzWYKY1PHZ7tWj6vjqA0xR9u1BDv8Q94Zy4J6OL4cC62cvEhE6GXsm2FKs
Mg/z3Sz3MSYhFf4vZwcsrhmh4tAu1EKzjkNNPLymF6CKq8Z2SZqBbPtmyN/U094O
K2U67B72RXwhj1evidiU4dYtOt9U0V/aCDgilJBbWbsVZEGBhJeXqAsBREa/RiYn
akGdD8/UdME3BxA9hsZJIE2JwMav/1/hYjX5A20o0uqynrJWfvTjPm5umCIKLDRg
+qJ2uLWQb2JTajIKavjuZU3J+NuOiU9OmkfqkmbQO0giLKGvxiPG0ERDBVVZAiZy
Nqxpvk1dKEkJzOS6Pz9D3/wimXkHIiqlGHnsO6s238/xBhhWPfWu41rLIYXgmYHM
sHhnQKv6d/CAmkm1+c3PQK6IplrX7296kr2VOMLEZRbaUgqKSjNWdmZH3Sx3UVsU
ZQ6JIXpZtV2N1ab/E0ora+7ATy29F1IwsAU4BooTgWkFvBsUnVgEkAa4Rj4YB4hE
s0QW5/TDGfRHkXYFapvf7MJAyDeh7GyGgmOvwO1ZscYkdcSTTRlcp7BmDtMKzVHL
hzAgAumE0fZp+Oc2yOnxKog8cMhwpfAfWtf4cHiwhhv5qYljjBbeLCAKd8IxdpUH
xgq9GLrpRvVJYk3JQYC1U9iVCBlyqt7gZ8MlSocV7MSwA6RQINDkUZh/h/uCg8QN
VMdqVn097ZqzU71e6crC9YS0iS1Ped8gHXtqCllOH08gVSI9JKKVpl2jsbS6LrP1
/gDqkz/ZZRiwP05NECiL47dVlecbB9ZFEVG5MDnjMrkpt8OcxGz6DiEnb8sqs2iy
G7rs7YDyIguldiYCKML3/t8WFBkt3qCtkO/wltfAgMAfkj6gNJiRxTLWKs1+cL0B
c41aXPme8mNHthhuKK8+FrjPorYvGo+g3XjhHPtGsLTd6Q+a7h/6xkmi3+E1gtNo
GXnhOicqCLo/KfCzG4y/qTqnijmD6RPO+kHqwVA+CUF+l7Q1dgEyngaCuOkPFh+W
uNNPeMDRff/OhdhELuViXp8fwEM7WS/zXbTd8p+S12e1W9orglF7gvUV39WwRohu
Y8aChPbqyZaO6CgdQyi/yms4WfQjQvViK6QOsJaFITr0zCSPIgAlaUU3v877lgpZ
WNsXIsoxh2N/ye1l78Vr/q5gYtEoLwJ82Zv+Or3+DpK6dCsg93WX/dRxyTy3aDGx
EKvtPRQe91OqCO9O5FG2YYfKarpD11muf+aQ+Di8PKN9sOAY7SZmeUIKQPLAAMZH
SSvYHelX/2cB8dh4Nf3lATXeKtrUTyQ3xINSNH7t4sxGcTxJSIbySSp3ycIaMtD5
ObEoarfFEid0YVzOW048Kl63K+iUFgOUhcMdFUqSr5l/xvvNOZNmxCfpX2ZwSYva
Fd/LTA+NZdqXQ96vtFOlQJypUjn5I9dAL0ljlF7wB7ZzOtvgfH8e0TSozHxNrtog
4GpY3un+oXnVlpf+o83gHY4xu7xpI/6K0IVgRioRVp317whS/3BRr3MU90V6FvbG
WSKi7b8PA3tlBsYQ0IbggJGTC2ws4nurIvfffPrraIftyZMa6+SYEtQS1P68+Kjm
ztupM5dwaiT92Kyjlee6TnE8amOCybmMITHOjf7vlU29fVD3CoqAqjrOBBpAjV/p
gJTn+KUGUayZxAxw9Wp55MvaS/IqEYz+5oV96Wj0oWoubncjiQXRuyIIclt4at80
dlLQ4AdoMiYWN2GgMBZe04shRgCN04Mmg7l7qBX13gMA0D9yoaA86X+Y2/CDKajn
JhIWhLAggqX5DfV0q+opTgBEJhjZNAGQpnCoBncxVr0RAkt6d1tPiAXQAOOTQHrG
xqJ/4or4Is4ZXTuAGbVvqCBmbrUy2hsbQa/5p6bqQWUouhqwmwTeiXBGMgaF3iik
DW9bd5ya418gZz3ZoQwvm52dxpLR5NYaI6aXsQx6uBRiDr4mRAYMbq+aGhmpDlWg
0PAdMCWgFPWnxKf7KyDRNuKlG5wQLZrmLfymudDB7PAH79f/6xrA4KjLqy+FJ0PO
/OCmdX7hp4W68Dhtt5lVN5CSUsiG12YRm0vrQOz2OJ1MW2/oxWatOYiJqXJqzM2g
Y0itNgy6v/J+fxd7KtEq4vz4XJy/rlCpbt/wAajHmbLQt37+f16JxTnGIOb1GoFe
a7OYZcMgQjulkyvVixMuYdjEz0HWCEPwTkB3tNPiOMYX/BS0U5jDQTFdxJSvix12
vA/gTjjX7E/C3liMgK63YsGEmNrBMO5tQNQ/F3ZFZyWmI9fMZQrqBFg0qgWFJowl
Q/WW3XXQfu0sosk0NTtlA59BA497ewQ5uChlWfUff3incqNdGN8u0XH6mAcK09Vi
he4Xgs/vUoe60UpcNGfKtNUQWm0Zl5R9J4ld3QKrx7nZJELdY47LXniGPePOX2d3
0gQT+LsKPQZIrYKSAvdD9/aflK31G+WedkYGZhr89S8Wnkew8IH3R9r3nCx5dhzh
TSfpnoV8Y7guCeYRlmLol4PkmwXiLaDWQvcrP4TQz3eIEhZRFa2iA2HagIICX0P9
QafnAutXOitV6kW7+VGOIR5DKU1M8JO5waMKn4cGGe7h2WPQJBbP2wYqpZbbxZTW
9ENY8bDA82aIvwJy0mkyHqETus4haU5X7CEtVpW601tt2P5tRJxFM8Gd3MfvcT1U
y/kGdLxPWDMiSEbs+wpiBwqg54ygSquIM+9W4riaR6EQuAWiWSzVWM/1IrTqRB9P
+VenG4B/8UpGSMuZzI7t7jzM6hvfP5B20Cw8UdszWyeHRGnRgHgkNP8rSfuBI6wg
WUmsCaiDllthtpeein/ay8Z/vOboZXOQ1OQcJzQAQFoQO1fyDtuxb4wrUkrdySr1
P2Ze+sEVoH/qCjdlkq33BIUAqNt4Kqs26FTQDFFju0O5NQAVb9LfumpbacTitrpK
PB6wKoOukqYXUlQyo95K+bnURdtaI+UnL2N3wwzDdmIH4+2TxgwUQzwHQg2A+ifU
GUqQ1ik1Isc7VgmY7gw5tGZQC+LTbfCDnnx2sjCmJXlhlIa/7rwiuywLQQnlvcom
Bz/qq2t25ByCybF9CeLr2Ke8muFC+iFpkAtf1MhiG73SazNxmhs8LTRiQG9zTUPV
bAuWDkJCIk1tAqm/uRCsocmFGb9oUsmURBun4IU6zd0oUg+/vDE3h7jN+mz9DLaU
IDICwHDYxdWOW3WRpJdLa4p5NgIiPwnJY4ATlf+KmI1vVDiBhojKEFbSUa51UmVa
u4yarzhAdJhuEDM+SslQjEks6FWs7nk6N4tEVa3CjT7HBApEXTC7MJ/7nvV5jr9W
fq1/ora42xbiDl5GYfUS373NijD81pSRiN2AIGokn8dTcrBJxRXtiQDdYLL7RSDx
XaCnq/cczOL1oIwVG+8RpaGDHQD66gb1nRUVWXgw85s4blhk3HH5SihYK2FRAzUK
rWrDqdKAIzHnJPs+g2OASO4u+rDMNosuJ0/YYT+W32FfXG6IQOknNLHT5yypHb/t
fCW2pTv+sO9EFJmuomaIDdRZTdHUznv/InC4YK4JWIZ3oVWvtvgWfJ/QkEeYXo8n
NVhcQaSCCSJCi7BqBg0WIKj09x0Um0K/nvTj2gdrTCJFaQ7URmo9xYJ0lhB+ttlu
gIQU+wFULfHwrDl/Q0W1eBHZ9+gAWriMtO749sBKwl7TX8lihFkb6cuwObJokPeC
15oXz9ypHcGFhshJ3xW3vQzOyuwpuTjMyPVmrSV7hWmi+W8L3C/1h25JejbBUpFY
GFmk3kZMvilfRmXQ3ALZN0HNwLOFyiWYJ//kUrvWlO1WJTwMiKHA7Eimr4FXApBC
rTyuwe8yht62yVEYw0UHKAKUrY6d7MALjLTbJdnma7O3KoByeyjc/RhHgH0JINgk
p/Aj0RJ//pylRN1k3Kl+6CcjJ5fqWg7qM+TVKeruPFQzse1mNgjjddU8+8YzriOl
2Goswh1pjVl81iCz0DBGw27xE/wD71JWmm0ej5HJ1Ex6NY5Oimvu0M9uBvsa933U
ZR0GpSC8mEQyb1uciHSZykoyoAsMaLRoifaNCj4qOrGbso8YBIka0EQJ9CufMjMn
igvFYBG0WU2BDebvIE+EOStZvPApnXgNXCQpkSEgH04YIhAcJ81P6nitRru/M/I3
1c4gWtxxhBqA1aVpaMRHR1zyQkUzIJtEmLo5cWLh3qFviw8XyVfIWfy5esm5NVca
79o+h5TGb97swEC9AjUjIwkq/fq+2oLxFCm2866W+hPbTfcvab4M593I4tdXUFeJ
6VuPJApM5hJq4grF3kAVHLGn6y46g2ZPXACEPQ3jIDh4uNHFqRsmu+OyTxyeffmq
rZfTebG//0gHRU9OOtiIYJy/zKndPRT0cTxVEedhSuZigv/aJ4YKQSALkToagBDY
CeL9cMsDXiONPm9vIlDpvGfi0p9ajCSZo1PTIRNfeLH/eGrtT79kH8B20xGaja6Z
iobVwqbjGF8p2ZOpeyKqvf+XY/0QoB0xzoXcAQDRFNeTjkGSmiJ4FT/JKJc2SKzM
S5NegIQ3ypv5bpgp6uv24yr9+nJhHOgDtVkKgtdrKrNngUcCkSj6mDaM5WqPJMOr
gaYNXhscbaTml2uzozzNiB/gnHvh3D/BJK4nWhcvmNlKCb4qwOQGjoEAsQhTRZX0
xgxBFU867nTeY2SBdVFxYE6MS8gi2EH7o0RztjUZ0MJdNhLLZimt2qK3linJM5Ga
t3cvXSuHDGF/1qk0JWwUFCQo2z6SupQzBVfhmCheH7vHkGST3vtrXgNKYlOhv2QX
gyiKMzgYqlggdSxzcQglRKPrids3NAEQJBS+wTK8NhiOMerQGRoycrpSGePQf4uv
6rXbhdHZbHhM8C4fU+2XQRcNw+0HhMiIUoVLtTsSUUkays6Bx9V7vDIw8yiJWI1T
d/GMuOTZT0C8KsPpu+WTDEHbU55vNaTN1VJRJ2dUsKe2pTBQ+H+vSIGClXp/+Jn/
l6YBh/1k+HktdGPlp+Q2td5ys4vZSMr/4GvJS2a2PNM7MYqw1dMoLqKQSC7l0yX3
EsBOqFLHcZ2ICPMBRPRgTYihX5wi6ZAK27uk3BZbMbWeVQR/iFqwTtVYVCe7Bsxk
XqmFUEcUj5jCLoL6epIYc9U4pS/aZGHNnoTCQ4Gq+D6Hz8EzuQIpp55fdA7wZEaG
oIHGhxWZ/h9DHHu/u/t1VWgYIXmymj8qV8TRWsgb2YQk6Q5TfaJIh2skdJUjJ7ed
/mmSRyPqAASAHalZt5eI87LaIbVgQBCmTx2a+C1rqXplnvlwkroR1X9aBiItzUzV
x7JmgHqvYrF26okYqX9lyaNzaMToxbKEGEsgC8kigCcgDJuYiQb4sOs1g8C5SnYw
htlyflrSdhwEGnTrF/i9Q7E0Laf2Plvj/ATGvEVUidP6f1IlBu3oz8KXuj00wyAc
omhaInu8XTSkiNxoU99plMVjReLwUOAZYSJ5eeLo7ExwHGKGJCKO4AAcHqq70ePH
HC6TYehDj9B8qbCt4ZPV3Fxjc8HGyw+rpF42xVPjCG4D/K8gnrzhd3B/4IKGT81S
LZRtCtDglhXAuo6zcdgU7Kyp4Yh+vzjemX/66gQAxRQ82qFwpooqKUi3hglmZ+hw
5czHDKni7kUpAeZQc7Zhi1UcB22IjC0ptIIrvUj+L2/ldykwo7GJdRbhBDZ1vzlJ
LWjYkMpPBlElX04298Vis2LGwNIRbbObZHEiJR3durlIT77lYbbdEB9EtvnnjbxR
yk+ui6kgH+O+D4Ecay/grf/bZv/ZIMnXMlfbC/76hSPf+L5JD67zmWo4osvJIBEJ
Fbu1lmfoW62q+17zwI3almkBpK/8jlj+DwsHgs2hY2vwbEpVYMQu3YWwT37MXz+K
KAqDVQPKtEvmzr6JMBFcenW+835N94b+6pZDHWaTv88yckM0e2nSno+Mek+r+6l1
iUzmSLKBEJto9PIGDPock/uAQcbKLolyPUILssF6x+Eo7xixbcMpAOYfhVCtIBWG
YVCsszHFiwVBCSoXs6xa4TItsY/ae1UiTblcnLA/2TaNZcjfdu5XwwyI3lRlYmnr
C8sVQR1rqf4q70OOAIvuTO8zLtCyVRa1N+1L5rrkJJ21k8187mApqwI+RHqy12F2
JsFU+FBad+aWky0rw0Wu0XmSBnV8IFNtOROY0oL06WgbtnecQakDt6cBlo2L8gkV
06VvK4jRClBMjFVcSAvAKKvZeN8yB5DxRVwjKg8mqTyjbgovYJZTtvihTqQrLuo0
ZrAiqlspPeRyHJ5sGAu4w1GxbiFy0Eu3XFzgaX6I8tPY0FxCtYhgQa16VK9epicd
sCtt1Hmwj9G+de3xOjxzTMq5lbudgnr24gIGKhA5dgt3QJXR5tLMGjq6mXXj5asP
Y+g+U+Q1RQu0kpHSI4DcjgywS5qll5kIfGFiEXe+TEflNIlGGhP2sYY6A9g/Cj+O
ER9Jn9vFilrXa8ojxHA57FJ/T0c43jPrzU9brNma3wEdLo1k1d3LZmcbB3Dbhor+
r0K7x3ovz81NSkxELCrJMkjFg25VY7Z0RAAnCeoQODn2U4FVw0A4m20XFCcW0I8r
+x30Kswa95N3QxjnD2gUOUO1ba8PpirNhDLonhY+2Q66INtVkoufN7eCM3OGQgcn
bMd+MbnxkbqbC5LZmnany2sUhP/5QgB1aGE0rP34FOIPFtJUo51usref5bRUa0Od
nPXwY0JFzc6qovEiFOAOsqQ6NwgvgG72/xBc8yxzl1BSZl4YSGKmDqRoR8J2qAtO
4iTPntEAl/goTdr2ley4PLEIB6+uSMsF9EvGVE299KaoIY2EdlnrnbH+23NKHZEb
ec1a+qaeP1qGHWY/EsfxV82tR1kYuQbJoKlFPFafsVHKO6Z+HVuQT5OXiTpHEO7h
/1yA66e6iljdt31/MdcbIzhH2NrglI1f6gt0b9uO2bkosS5m81T50Ddlkw/N6E9H
2rYIFFqNOGSenY1WIAvtMLVjMVbL84VgRoRcWBhqtAv+pxMm0SzhWne9UTsmp0ww
BG+stKVlofi9W6otn9IHhk5+npghhTO1H592BOkP5gJxo7swfYDgWnimpT4kOr6Z
6viGn6pZosKa38INvHpVRYZBedmDVVQcqGMg8rLBee2zccEzydRPbstey0HLSZ5j
Kyke/pLiO+ON5u74b2OPDTyB+CPQKv9DcNONu2aeqWEv/Y/9xgRbVWP0RgWw4HU3
noPlEqNzS6jACOCnMAF2liPgLnRrZ/W2A0nDEIfgZkCXe2ccvJ/mqgLyLHQfVWT2
E4Qoxj/0u/TzGzIa5w2ZMWoc1MoqnlAh6pwy4GxyKOWp/PLb2PIt7fLWIADevEv7
Gl/J5MdjDLedRNe8p9FiAHrLQ3ORfX+30lf3+2oDVpj9e2spIJ0XZtI2E7AlRISo
KHhsvAa0Ne4tyIE9deuhQfiCySLTdDI8J5quw03JnZFX3uqKJU/q57uwtezE2G+v
OFvStYqR1Ypg8QsI2PFwFHFiuhF3+X5uYBnGjQD5RVMuLtc/MVgTQZWnauy2YYsL
19j3m1pvkILIXB2aT03R83GOOOFuU2WiMqHoI/+UfpZJ0nTIr9naDthTqpyclPKS
rSt7orynh88At63ReIOau8ZHU2RcP3vAdzZOjyqfn/pADeROlnZ8inWzDQslvKDS
zpDR9ixYCRH/h31lrcRLP64nP+Au/wqFZdIv9HgEOLMKIhFlaybzKBRD1n/owrHg
E5P541jQy7AU1mMMPgY2bQETaE560BQcBP7MNXUcWoh39PoU1xN9xSIzUJQj9Gxc
bXMHMOfJJ9dwIpBk9RGK8qM8PTqE4SC52CGEPKbWMTEThfL8Q7lIdeBv4r6kh43E
CG++HLynaSp4TSfxxi8ApNPcItJ+2flU1hF7ujOX8qohPIhELm8e46QGat4OU6Ar
0ajJ0DSNs/+1D/5MLCSBx4Ywr2Uo8YExGOwi74eglQHQqvaDpzZsJ2iVOyvM2axU
7WXbn/7Kd5Ghu/gDjlfSi+DzNvEn9LBhvgzAfC2r0S90o068x73lbNDOhy5xv2Rq
TDw6vUTVHSYM+eq61N2LR7YqI3GlKVh//h600ifPWHUpXuUo/nVmx14FbJuNVVO0
QBKBeFvpkBAqxR+XWiUwnbbJSKKQgDEFeTfV7P9RYB49EKo/8Wqo5DHmlH7WsukL
qkdcgf9WhrAER98zplmO3rP8K7XV2uMU5I7yWo19uF75SnMS/X/ciN+gMviA3SOR
6NV5wXslWPJWs58fNXkIaLPtVxllz21KWR1KeEtiKXOb4L70hEJbX8O/O1siH1ab
ql/VB33dl/15AkhtESTXX8XQKdYVGXLdfbOFAu//kMX7gv6VEJtOZBEmkWIKQGtq
7xI6zs7uJwT68KnZHXf4KkvqKGhJ2hzG2ldMUi9SGdm51EIk13wRk6WVXzot1YvG
KkDMhbQtIXZOCxKWpxvoldMhxPuqLdkHK//NK0L7P/km1Z7cuPCrEB7yreZz3cBo
2TNGGp1KgCy5JLUGXQFhHunGiEUG7MSk9qnkBjA3+k3SXWo4cvM3eStgE8iRbrSO
v/A/w1SlP88F92v4ybkmBBlGmRo10wtEmvkUIbm16s79iFE48CORGKKGks+av0Uc
kT9VtEcASCnWdmTTkOr9ZKdfSAdkiUU2qZ1rE1AIbxPavEtaDSdMCY123NySfW+Z
gVjKoDPhBHXNyD5wOXU6dBI9iY7NkxZETFUb4wP3JtnR0kdXIneQZSs5GAdmIgaU
3nZaROH9aKgjxP6Vb4MzhGd1KgjsesE+heqAMUM4Vx1eHWxVgiJCD4r6yagSMwbC
DHMsWMEGeRcZ0L2aTfszCWZtVfFrmk115h4G3I0bZ/OoCzJVObar6TzXq2mOUbMi
gTVnXQxaTvGOquCooDRfMTrPl4PuDX2Fc2cCZ2wqfAsOvxJFXlYqxBhaGdJtewb8
LYD17kUW86JJQNKNln+iiOmu6CfL8oE2b12xiYpISHbn5lqN9mZi4ObBOZNR8lny
OrCWc+ZNu3uTYKXSht3gLOrD+8a32/0+lxbiBxcFexZdU0opJLn+/poQUt805p2x
Vh10wmII081m9dHFD5Gd3EzO7RLPwWDNqSIUTGi+b1FqiOTuU891c86TLRJJVpg0
vxitiXmkkvYe9X6YO8SczZPXwrKp94tLv3xSjj4W6y3wVjLJXXqktQSBKtDGltzu
0ZleghXhJRWU9rRFyOtEzMqKc+P0Q/uEPeowQxV6MMxxbUaYHc2PYi+l3KqFE/GF
xgaI+lSDwboJsioEeO9Y6QD/2i6STp/6kiMAx9HAk1qRWlRV6HYfahQ2bMp1CylN
r8gsHol7jAitwGltvi1iag+05EKbuiuEttYMKlZ8jVUlmdZY2iT3cUIa9vNF2Q7r
6uDXAOl14yCXHnOASscrrLm55E97hY0wcIoQwz67YaxEP7D+U4jmK72LJRL32Umq
eGsOc80wBTXpBeae6Kuhg7ez544ql+xPZ8X8A0bupaE9PggBum6WnvSBa0Srq1Rr
qhIwSoCDAZuXN0pkRFZsOESy2KUVlOKsux4oXk8nMBio9ZPSIA/02/RZmHeg8Z4I
RT0qhzk8XK6MY+p6+t3yb132+mTycWoVBRiJsSyeAnUBMC8RanU9OrURmqx6eIGf
TNlYcLJ+dM5Fn94OqwT4TdKr6GSNweBJGKciRsqsw/1lkHf792iHfeAqucly336D
JetxBSlJAqCTFqeMf7K7HQq3bHvj/mlvAyZOY2gyQ8Vv9dJIWMl5/Ltdow55VCzK
Gu1r7J9+O/WY4JdwC8aAxm84vBmpZP4DqnJa4FOsJ/8bJWZs+THme29WX2fxUa2r
DlU7MoKbda/6BAJcnKatOQwKrmnhR3CCDgxzX8yaphOeiBbqqE4zpWqW6Ls4hfD3
9oimyaitdtfOv5OFbihLE05kXdanYdGmHQw6fWCdjDnzET2Tuhq7iaya2HOeFeID
waUWkH4sDFolyMwZUP06hkNVs85duUO4eCugx3v248mKBVF3UXyWio/VTIKWn//z
Xg/da379mVF0xM2P5uZEqJSfswbrrAghOmI6H5e5+7rhIl6xswFGulppMC9o5jC5
y5PgmBfj35II2YL7KHf2tvlOSItCVfBDKpxBI+aPLBMZtyM6LbVFmeDXPLznHP+F
SRP+SU7fIX0R3bQfygscnWOWyn3VEaBIZrnOs4w/VkXcFc4C42OQ7fPMjSG20JYw
cjiIWGPqPJBE3MHhrqz5kL/G8AgEH5wBQMJHwtZY9xqnh2pE6pxnprQXhWqtbqI4
sGbBbK7kgjsSZ678mMhOX7tbbfgyym9rbG201/FmVOFu/fif8dVvOuWglGFxsnix
Bv8GqZurEEkymQm8mgOX7Br3FbXdGFPaPK09hilDzf5tt/OssjH6bGdeW5/LTfXf
fDnKgcHBm0SctjVMSCU4hLS4KfTL8kOD2RaBQxdZE8plIAtVExve3d011ciOrXR/
myY33lTrn3Sf+r+OhOeHw8NMuiM78NQy7rPT89sew9/I+2o+P5ZMLAyuf0I0f7VE
NKGkTywbbxlGcJlToEoXYiO9Say8jdpC2ZBsg72Sz6sylkPATG++UeBX5PyXZ1Xx
3DBi3XH8nGOWx3eOqBa82J2MfWoRyvzPU509HH4hHcB4pctTUG/pM45A/EhyqyDs
kh2ipbRoI40anVG84fVR3G/pJ+5YhjVrL8M8Af51M6TsiVUmpXa3Qr+qt0BmokLT
BBl9ekxibY7SL7OqqQ7mS6I5UqVNORwPB6DZL11Cg6x4qOrsYtdxEBg9bZMuzZNx
U3bOUwg6QLGhG78H9Uae5iF3pzSiRdiVSgTJCzPUcU7TZuExJWTYQ2Hs8JiC5AqI
6+3sdWrlsXLIj//D2LAOrSqS2kIKYMf9uc/5e3R6ypvlHmzvoUDKQvP1eoO4Cjfs
tv18VhAzwUX0vkpK7ao4BTuDFDWEpX6yPbu8I0eBmKVsO6UMET8m7m29Ar/ZVLG4
Dof0jKqDtlSFcHzHo74pF352dfsNEN9x3Ge4xDb9zJJ5ZFz6riGOy1HjeC7eG+ob
Gmx3xGNwrxcKte+ZWyhZARQBeknmEHiHL+DtFi1uJrGUPmdZESy82r4bRpIqhmz3
anmpUus4OyCxxUQQo0cr/Im8g82+3FlN79xQ5MxmqVHrFKgd6FqB+AIrpGgA5H57
+MhYz5C9FWaQY75n9SAQeUeTPV7IB1ytuDI6xpVfcIhVrUm5YsUa0QQOZaPN5+Dt
9IKrlaZXeR5ur9guzXp3aaUK5t3IZTKm/Z4xICkPJMen3vPT7J2aOaoUSCiWTa36
DiSMy+pxbKscwTyr+J6IEMTMj/cCKYf1HI3EsZ07kGt6c0hmCjP5ap4ey6nLIoGW
UZ9e26cEYd3MOFOvjauqO7HF37rtfmBX1so5Bo9n7VMqE2iX7+h75lgRjHJskXOg
a0y8IYHVIBisWPV28uFEyU6GKu7vvtTUkyBffrqprsNr28+WYJD6JsAW8o9v/3jt
SBW1GMz/a4zkGK8acq4zkvYsLd1cg/qtDS22gP2gMcaTRTxjIJG5dXRYAsL7JbDl
04QBZl7niH+RgvVuRAn/kPlHtArXXIiDenqcRQf/ClWFxHvqUYwJqefDTGJtxprK
Fa1xwpTIWdkwfwqn/UHhIIy02go4HGl8YHi0E/LKAfSKYLxgyf3lBFh8B/pqjaDG
47HYivsQvOqbRk38uIE47cQ1ozc8De6RpGXZ4ru/A5lqLimWVIjXqrJ2B2owz4ES
gH3aLf+2TLme2UOeOjcmJPtxUSTxfwTqDc1hkEGG4ujuetyZmelTORHmxPm4GZiD
gsCfG89BJZZcevdn0dyvdG36+wg5vXjuc7bSUvV9vbIb2sZw5+7gAr0b4Gzoq5yn
pXwvN+yYc0/VhIQWt+3fuQ/pw3SZScqEOwRddGOdCUStpCZbIjUX9qatou6YZvhR
J1uKOJpNEWSofstnodIf6TYbSPF8yY0Gc9GjMDeGMuL5yaaGw5H63DPOQTnQG0AB
SzeGbap6iy0HNOtQvu/1BXrWLjVtRHLEdOYOq1VRl4yWavOVS1GOzBWoTEXnMg4i
WfKxRBSCgrqLclk8W68oqMxEmjqIMKtME0260OC6w0e0DBCBmHfvzBK58w+0sPiD
NlyW9ak5MqyUof/gGcf0eKGSAfBQM26jLsNAtaU6DJ1omCJC1Ki99j4+3QXECQbM
EkGFrlMxlFUIPRksPLSZt9JySkDlhgjfLlsZHHnWteD2dawTd5q3GLBHfIGbNPdt
j9u1uNaYv3mY3NIQkKnM2CCW/mBFW+BM7Gs1Cfp5RRpCvYkSD8ALPb1M23YOhPOc
H2rOrfnQlGJPh9IS6/X+KZswt9Iiul+YjIAcOF+ui1MRJDezPib6UhErXbXYkd2u
N/91H0KSfGEbAKFMz9TRjren1eS1nMQCYyGwwpwpJTbBbjKzQTKCq+FZf9bTgWlz
jYSv+G6gHdTBcTkCadpHWWNYHnD6Odq+g3ioqvgfJSycna3f30ntSSFdDqo8UfDM
I625VYADNvjRVMyfQrN8AMqk/s8n4W3NaOP+2ce155aQsuxHJhaQg5VB4CDxqF0w
ot4He722Ii80/aQdqq83zK+eb5X8efu32D+ZdB2mD8wKiUZvZMHKEw0pDY9XyDMQ
DVBMYaUbQ27lY83Lw5cFMVRIwZcrXxPLx+bwN8s6NTNWGD5Xd844pohCrFINfqJe
ZCWTYqEM9sMNP0CwyK6qDfFvHSnvGm9g7fAWxy6owFbetAZO/Ls7qOMLvZehkKRQ
8rTW7oFOHyuJXRO7bvZ/3ediNcrOTlQt6BC7hCZKgcb3mqrOrgm3iSODBpGTp6BC
gijIJ4MnuS/wR7T+07ibc2bm1KE4lD3j7ZD2UE9iyYRYPYpvuOihiAFOAtDnZIYH
t5WMja8hOp6KwImZyuuYRaJ0Se/TTMU0WJv+SxVexCJC8jJqb36Q+sPrt6DvdTDf
NB6+AJPNPN9yQiZyLzvWXIIfKWrPRSIYYdsSWuukCNzkIk0+bFsr7keaJKv0W9wn
vL1Vnbi50flfAYXiJeNJ1SiCBpJ7maqWmtNkB2c3dvi93tOcA2Sz2GIvmzTvUaA7
Az930dVvT+7XQFGyGWXt+xLsX6ATNsCAS14zD5qTxqmHmJuKV7Ypv+/1HJJphCv7
8wStWbR76ACp3w3QWsG205Duzpx8pFAKOtEyNHNIgcJ3/fo/XnlkSTX7zmSwmJeS
O9oyuCulnt+h43vOn1kuCnDg45dqQHxeiEUCpmxjuMeF/k0HYSZcb4do11kHDLvz
Q/n4gs/dDLnFkijVfQ3Wwloc29aMjjZ/NXQucpAOhWnC3NlNIV31hbOt4NqeNxiB
O/+wqTze8E2DyJaoOhpZMIVOCJ7zeGr+rvDrBz7NcYYEyoGS4U+oBdKJejGzJVMz
T3RJr80/+d+/8mO3kp2pevO9lE+SZN4WMElaciEUMwzUq2qs8fAbFp0JeXf3mxT6
DaVmn7SMoltzrMbNQS/3klseaK3SFQNoPm2AAnrtEWjNxrqhC3wE/JOGqioiDAfT
8zQI+9NT9DTv6CPj2lruF1hkElAntLP2hRwjJf79HpVm1d3jb1/U/dY9eJJNIA4g
YYGRA2NJ7wBCq7oBoh086373mF0kGUrY+wOOblNAywBOA4J/e9jv9xDuWJ06nqlJ
MHLD9Av7vqPKHFS/HPCshzVIXmVY/qt4ljzQh3/Z/4R4m36W427N07X3azkpZ/Su
gbOrvG7xI1j6EWECttcsTQpARhPSk5ojSto43skfdP0H0309MD4VHEt9FevbKb74
BHH+CRLQdp9jkD5QWpbqm80CMuwAibc57EZkcb+01EojjToURDFGVrd3j7uZGVX0
HrbPx+QFvu9etRPRptjllKHqvCElps/cFlO6sYcm7zRjDrKxIELA0GHvys1CKyoV
x//AlcstUfLKuyiNz7leYF9/UfM6SYbkwqS15CdGCCREScIf8elQdid2ugQ9bnR0
R7GF+IirVQuapNrWAe4iGxwqCo8/OTHYLkG6R4pCbExzxJ6w0DvLwdDEnG/wXKWi
lbGXEyqihT5bPn4q5r5TeH3HvcsGiGAKeNIRjhM4HvpqaZodboM4bPbFEJY+7bFx
A9WP5ByF7XgufxnWUDVFhmUC9VKdtcrfwNvhEiHPjO5vkTnn9vpvURxdfi1K8zIs
SDugbUbxktLC1OT86pIEz2ghNFWL1I0gCkK2qLpy0CdoHjsSgSpvkMYO2AhBNtkN
iJzjked7T3gbmp3pSCKQRb69IgDH7e2EKRdb+JZ5YCEmBNQXG9HcVEvcRIGWx64v
+A8K1mj5g72IN0mp11foE1Eg6fyeY5PBVgM879A6cOOUVO6nW6DVh4Oxu1lcH6f4
F3YTPyu2Imiwwhy9BsYIvERcuCzeTCLxcDpx1wvtdTllpM2pfSdn/KY/mBRCWPfp
IfuXZqUPbZggTk3/ZUosnv+REyeEK/jVOd0ZRyysH9EWlHGV90iRztk2AmDmw6Qh
uAIu5tKgeoEb4/nDSKUgv+HWgTlewWzC2njTGwPp2xeucwA38VTEZSis1E224c17
gWH0P05ckhIX+jXLWh/kFyl7P7OWC6OKdmTRHETVNyqY3Q2TvVKJ9fYbHDRZqKKn
M6zNHmFxIqjb9NxVTbMxAsy8O9L/XZST0o6L8BPvFd83skNsvuCgcBOovMdAhDrH
IPt5tqD5RsOx/wmp8A0SH/nbpiW/PpXScpd6OqWND2lGgmFtn3CuB+PdJ6I6B3kq
pzqZcRkgmeONTEYsd/cb/zm/5cPHhjCtu30W1hn0h6JTuZQIbAL2I2xsc/gOVrjC
BeosH1yP9VsiZU3c5Cgo+senrW6N3JOfPwLnTOryd959TR0qrUCsCUzkD4uasWHA
bNapb2FKYaiYmxnuylWZ5h1E8NqanPDj985mbzhU2fBtieNvC63xsJjp21LqeeUM
HFHJM2SDkOEi1aP7YQc4POmz8c9XIr55vJCwRwYJkgxFHx2KsZTtSbJgKMjdAGkV
T7098rjGld47z+WEe3SfVOtfMsP20EZ8mCOIP4zdfbIoGMElo/qXFnqx3UPHUnvx
Rz/9vGA8E8NB282tRkujArapgD6/iLoma8o1SWJkLgiVQW/T/MnH1b/tvbAhzIWT
fLK8bJdZ/VTun0mz9nN7fJ4Pt3flAcEUn5KyENhoNrdIhfQoFMDnqhX1w+864Y9+
ihjYIJj/sSAcaTjx2El/tDAMoH8QdXOOWgzXuWbZdG7yYCeDhlj7JuSO5R82P10B
6yS3V5TXbsVLqNLLVrEM2RqibiuPDUHF4forts3LQkWl+8saEtJjpkSc24Ur/E8B
3o0Vj/AGRk++llQ/akdTKOufox/c8IzhYdUAtAMoi1S0O+Gz7VkUmlsJ3Z6i/yUr
ucHaXfhrFRHNmbxJmMnIBdb6mFH1br4u25+59r8e6A6gPRAS93Yl4knB+gkZeqr7
61PkI0vZCKZG2X63mI2FozreXza1PcRWH3sw9N2K8L2jksoLez0tffiWS65Twz5Q
xtFk7gpx58ExcubdFxZo2q9bvzCRhBean9rutFdsqihzQtqAz14GUtqdIwqTBqrz
9NJoPOID7iHUM2e4W4Z+YnpBT8Wepwq5G/EPgW74Nkp4WfE4Wz+QGzLYab8SIlEz
w/ZZkd0XkyOjmdVRPKeDLipFuopF1ZUQ42e6x6Hy4Pod6UdrnjOgl1WrAlvuzaWP
8WHoYhXetHODhc+ptE7sd+ySfYRaWsZVeYSesv3eKyKqnasRLSd9TbRxXbFGCNQl
gCFuXHxZJWLmCALythMcMJRWPQFlHjqiide1znGpDOOUAQPNyydzFahlWxphzp2+
BBUX1b+wq329JNaJ8v35+RGJzgwiJnhCOQmxTkREL0nlIOQBZT1v0csfQ1b4vhBT
kX8gP/l8ZU6uR7wU5SpCvKfxi0N0OvNxDBYY1GDllMWq4dAnY1MI/MlQK3hk1txV
NqubR/bX8Lh73U5CBpheCyhObIOhqXjThrPuy8lx8OAt0QuEzWVgPVAtaZOQUdII
auvF0D8o7Cc6SMtOH2WZXEQKCe3bi8LBNjSqYlRSHIwTAw/cRSSa+xQHb1uq3jUj
CUG0Y36gGyjzeKbCNr26P47X9kq3XE9yhUiYTFauica0r8fMojxxGWVv3+fd2mii
DhoZCZuEmGDD+YHDm3yPJT9zL7Ln59li5yNd5HAqvj98qU2jhSTc4OmZbvDYwDFb
gYeoMgaJLjlBsxh0+h8WcCVfOm4QW6jfvGxERQJGcDLkkmI0fWHKkeUDHf4D4KBm
idLF4lTxzuKOVSJ9+SFjaysN0W9lszyBOatLC6RBxeVwGbxT2BC/mFY+LuefsqII
rTKcvNduLJXrt+4sVdKPtdkfwi7p1b7fFOlOh7xAvM167jWQ+Lwxw/oECTLX8fts
Mo4EEgaaEpjPhT0FU4BN8OCuMwCdN2Q7KP4tRcKHe9/ggITtsje/+q97iswxtvf8
/WV+WpqcmaJMLOo9Bj4Mid9eD3ANEeSGeU6BG+zsR5xaxFroqRaE8rijutlxm9bo
slP3EpXhepv3jMfhzr1Ci8hbbKLGzWFzSt5ivlkApPW4kheqcOZHTQj7ThXXKgif
aO/V3fhoW8hPYZGHXA1Qx1Ki+LxBSO+HazyrqPyPKkb9mA+wwdI8UXhoyDxtKNuf
l7R4auejd/J/09EacBHyo616evkXWU9sFTvP5eJJld0rzeK9hrKE0HxjX4Tt+R2K
SyKKsYSALoFu2DmSgfAiJSAA9ZELsHgm3aCoeBD2Xz7NuYbrLJuP2bz8rNDoljAF
5K7P+U8q6nzQPsvi+psXyjhAPtKBE2nPUofLiOSWewZAMxGFaho1/d/pU9Vf+gaC
LVdHLcGAguiv8m1JQ8OXxe96/gU5UeW+5xE7hPcojSCiLfp43/KU9E5QoyNk7qbD
UHivIeQwqj/YmZu1ohrq9Ql5Ea9Ok18+Q00CAthUmqPtOl5mpdzdyQvMS0yU0aXi
nSGkhwMRn+uNgWuvqDRyCnp0OUOGd3MC6xlWCbOs5UxRHfNAewTkJ27B1NT2Gy57
UyOKhapGd1yHYvrNbmQ55r483/dEjFnaWAIvek8+gQDv04FreqsrNTnh6eC7bQd3
ppbjX2Zw6vDQrwPyoILSvx7TbEWa2r/Ic+CjEN+u3aUrfFuxHWU+i/+b1vBKQLL6
hQwyUYsa+DqGkOLjARcD6OFWyW2beqszez7vNILwMJqPXDjYeU59YCwQ6DQI4QB4
fFtpLlNYiDRCIiYR7RnxNPcxa2Y/BVwoTuD+p72eNnhWBjCeURZWIEr4Owwa1AL8
5CZnKNbJioHGFHe2NJ9rRnGEGAT0YOORyxVQPGDFwkV7d2ukDAqXG3dlMn/s3GhL
BdhAOh/LsVb1wsEG3BVW+z3b3vCTSXKULxemTe5qJAQj7IZnxA2elDMUdkQ9bSD8
gc/xUx1OZaJvtkWBJ57cGKxeEtlYQSexuWCuwCWlkPb4FnVfY+5+U9w8km5/yqwu
JZz/YVa9oPHB2Zqtd6O1OumvpRy/adnBB2qCsGni1tXGe032yWwqVXLdVNOD0vFA
3vN9gvUBBMUIvMC9VzQ1Qh7Q/2j0sq8eYuztScgiWMsVNk1UzLDe5he5JEXt8jV9
Vh67jrLXbx4RXNBKxqMfofxyby8TfSfcZ4Jm6cUH569mKX0pti8jxR7t2sMzv9sZ
h/iKWxO6DR9Ndt8K7qx597dqS5ilK/XCdQ9yi4FbdpaTf5t6fdqBmXQMnslghjam
sAARr8UGhh6niANMiZw12+Vwtl0jA3XOSqRTl9JH1U1pKRbdagXkL/y+KQFdYArF
LrbrRsRTSWuWmlF8FMfPj7mcbvFCmggDCWpxFOMPAxLeuZpo2G/aS1tvH+BjXfr4
bfPuuekPZfGTFkur9efYN2JhRct3jYFNsqemiAszt50LhA9PqMP3sKBSdA0mtOED
+WOvHogyxuKAH03WBxCDjmpB4k8wLWXR71OwhS2Uw5iixTsvTwBCQYtlq+K5fxBS
UzEPRuOTePeHg9UG25jxnTzjRyG/9wXmMBtyzHg5jkYDGDqguM9x8da5sG9K3d3B
0IckkR+fgb7Har88401yix6bCt/Y8PnUY8vMTdg8OZzUZ0eL3+itWMsmBoPxqBxC
/x+He7GuUZF0FBmxqz+OTNcfEmR2bbdO0Vu+dF8XAyc8A54Jkqm+WVhaSDuTc4PW
RcuGErRRpu9HiQDXgxtzdDu5ghYTgGjn3ijU+TZlcmzc3lTGBwcER6QFczdNY3so
8nOWf/jeneiooGGF20lDVom3x0c1p7sUXZVnq3foZDq5j21n8albxZz/RBMdGuoX
eY20ghvROoG0xeTS+intfnfU0zY4wTSB9z77gRF7d/B3f6bonHqFs2z4eakT853e
cSegMQGb0D/6E8KMvjF6HGjF4j7vJWIQiaHN8tdpmS9S/uv6WtjfqdQvNv2jmkxP
WgsbOQ+NsY1yYcQ2IhoaanYU0kUZ1qZlO95HYkrlvMYyALI7Xeu4gNPNn4Qc1Txs
2lbAUFFlw3ZjZ4SEHjwaNXh4tU+sZeLdPVI5QwQnsf7wD3tBc4MRr70SNUhw9rWe
ozH7xs9W3hbv38N/wDx6f9ll/7PdNYT3LocpEhZhXxIpdL/CG727rz5hfuUkA808
faignRFx0JUeok1kRARti1mHG2RZOpBJuqYXKgQsbCI2sfybKbO8zPnQIVsqtK+n
hjLM8wHEv/Mm/XZmMfSQTcF4wXGWeaTGOr6VUwyoQdASHau6gvlxb4YjULIWZcbA
GXUP5Ia7jthaNSFyn6sXGkDA4KFqaIrL5s6QHZXVl+NpB9QPeLdvlpIak4esMQQW
6LhZhKfRr9bFrXyOHu5ux8Rz8Dy1joIyJ8Af7YX/uKi9L+2FmvrdiG5xooGL+1nl
2JuQRFby9TOE3D3ZPdgVClD2eb7lOv7+juNJD5ond0yiMyLRN2voXdkK5ksjmQPF
Z+StGdVpcaQiGC2ce2C73cP3SFqOs9pTDyEwpMuFBymv1nAJFYn/R/xsQBLY7CXK
wheXTEcHt4n7ZQJ9Yd3ug9jNXBAiHyB9jIJ4JrHfh6c+2dOXOn0U2PrjbfhdsRIv
5NV8TOVoXkuezM0qSlx6QOHpQon/yoTIhT4D1iDFiqHcdkvArgJEG5sPATKNsHIH
uGQTcOApqm2eIEBVF8mkk9NZ1r+Iac7YEPkIup/w9ONXNsx3ryRiuanA9Tqaqb1U
SvfIp2Dl5DWrTx6M8raqJmRWfEXM9k7G0jHgT+FfU8YsE45FSCu8GrJbhoLPkDtc
VP9m2INLxHZ9/8XJFyda5P5SC5WpzMQ33x+sB6xeagPIpfRIUVXa5SphYepmLgKQ
7+GyfkFZb7aI6Y4HL3uadteISr5DmrMG+DsoyZka6TFQNZNoafNgkfyP5ouWw5JF
im4z9myWSnfJicpM3zoxe+OJJO256wpdy+9dEHVhi11CM/GZf8QGw/VPQ1rI2QE+
YWd0tWLcYDZ7VQiZlgaQ5H7l/tebjfi5O/6O0r8RQSP5K1DsxexjrGI/upLVHAu0
vqLU+DEGcuCsarsl93IOK7hjXMvxHe7VLGNnZ4yyVi3pmFuKyNrP1cYR36gWJB+b
wCih8LpD0js/ROQUfaHTEl6VlrvetiWxDi228sWrD5bMcaEwZ+nX+lM/nPfPO1JR
UfXTbui2Dlguzb/12sZIbs+c+Zx9GoR+/TZTHgQnaXk1N1OCT/dZ+ITdt6E3A6hH
AX/JzePrVOhfohiPJOv4897M0FTzRxRHZeVq/ocvhOLEogXbesphiQtsQAD4nGKB
BjkMrOU/+wx8LvenqyNq/r2KCUJMpMrwwKS+shEyioEjBEdGyjOc8zPyIUysJNxZ
WtpY4jfMBYcyMJ/lEGIz80bjHihas53hejdC5NX6SiLukiMVn25ecQRmBRqjVsqh
oD/z8YCVuHNCaMCMiupGMAs5HGLIzXoK/ZiqpHnbgkxOSS8JmJprj1ki4t/r5+RJ
A1QVT75IpqrFzcrgZp6DG8bTWWedZu8jmDRsuqzbuScZ0mZ7bE/BgtM6KTpWGRfL
Nc1SJfI8I43YVnqxW3koYPIbsTpn3OnwFBDqAYb/GyQEbKvai1NcRJea5dl2ZN+3
Ox+M4DTQp2Z0nj+0e1RgkjU+7K8aDKgzeENNRqTTMAjTrSqzN18rFB+Yo7cr9upY
6wEzqF+yi/FPkfM6L+a+7s7PueS2IzowEchmJK8y8ryrOBEOA7MypcvkN2Vf3Na4
X6lLRMH4H6KC7rrDM5J5RtjQ9xzFgH6kPj+urIp/lFcZKArITPUJqAxjpqXSpyii
8QFgj39AuSselW5Fe88DtVgfvY9JkBAAF/5xYQtS+orvW/sAKxZbFKrwNEoSxX2+
FNJTIopg12bJnb8bgbr72oRuMIB+Gjh79lEphkuQXBCZF5+cfogH5GxO+s+QhLpI
HonRxj7xyO7yS72IMX3L5KvpewPeufNdDXxX4qj+kf40KREt2aDFeGgdu8fKYOVo
Lkh7XsMm9kMBpjTkJv4/ESZ1V5bzViHQQvZVttBwhNcq/Ue5I82mCVbpJMlZ+Py7
NadG+2S6fBLbhCCcmjLouOyYAOat8ocBvF5BMdD2kABSxNKyPiLa8c7k9ZD+dNxs
xa9esh70qyvfew9AhkC3xiFBeDTMZ3rAooasVJ3rG4qBLd5MgN26iy96eKn3PwW3
UxqIRXmZBx2/iysSXKQesGm8lp5OSfbRwLQH0FirCT/Ndfo1sU4HSLAjwhTqMeJ3
csaftgV9S8MppwpgZi8JPhxArYl8vYEH7ixPsQQGam8IqEIuzj3XnmOYFd+C3LyP
q6JUHZlkWphgtdHRyRjaVlmXVWq/iL6s7btNSILWYpo6FjXBBgR4AVuqh1uVoSFx
GExkyKqrHJfeMlXGUXRB3XDIBncZit9CBD39mkU5Y7FKLvp0WcVCnbZa2g1H/Xch
acwRg+FfAnk/37Oc15EcLX3mnnZn/7HlPRWqcnWXqANWr3cjZcAVgi6CwQ65wWZp
EW5s9ndhaTWJ1xVGmC8W3lruyTE6xyi+rnshAlidiNKrYJTSmm1ko5hXqDiAYqYG
UnuRmIfuRoZsBXHi8f+8/lfYldnL0Vx21lD+ljXEUi/P7MkQZZh5DC2XoiGZd5oA
QUQYV9ciDKeFz3J44P4FqW8nPE5E5IevlK3BeRXzTL4wb1QlUz6tWZdlumyN2ZFV
Emy+stoFZq1oxYEfiNEFGj6sluw5zpXqtcb6TIvFFiUD7SVcpswVr/Oq+ZuSIJnx
PzPaHl4+c++X3U1QTJubgnZy7sWRUCwgyjXeD1ksd+Ntc0pJJmwawHsurBc55aYg
Pxt8QbWmf1SxuIMV5mZQ5zWXFJ8CWzrBG8/L8fKxI9BdCm3ZaNvIeN2pHeAsOxvK
8k+FdBxFO5Sl/wiMKg3BHZktoq6FYpTyexLgTP7QxFnLj7y9FrneVbK7NuKb7Xdx
skRIOyLqBjxabZvkpsCtaJIOX0wyAJPGqK6ucXG7VwH7cxNEk6gtP9900PVhqDZU
hyiHld15ScnaFWX8Yopi0U7IaItOzkji9EBYm8l3zYcbhQsXHCCuvqglYFzzw2wv
dPK1QcpqZ579sTjT9r5Ne8UypEi9FOXdj7uO+FZtAXhccR1SU3YrmNTfqWnRgZkT
VjNeeTSo2dH7HwcyWKwtignWU0J6TjjTlkBIwa/NRsSLpvk4xkyKIhTLsMb1pPuu
IGvW2XQ3gU0mF9XONDjbxQp6dBDnE9pALSAsKt10ut2tK3tFgWpEswmNt2+/aSYW
IOJsy0gUwRq7AGIxs02ancNnDfSyMAU+chskmkBOXYN9+e5iAMsjb3ZR/cKHCfgp
y/lucr1RPsSYPNu7nMPLG2sFL6SQgZ9BWCtpfAWYwygJkmahztdKPZmVAeD6vxjd
Z8MtrGDu4fMi70RikhqWSlSeNsfU1d0ELfX1hmSmLsXZccOeaQLbQnxVD9DuaUMD
SQzoUZB30sRLO5tY54gj0J0vnbqeWbeeo8Su7CmeuiVdwyGV0dgPVtA91dt++ucZ
AqJ3JDvIPTLnr2Z0JJPnp54yJ0jQbiMcKbzU3wCP8UnW4Lj3BAf9sWVsPcyRoPBR
s4L80U/XjfsrVf16WHAW2XxqH3XYABBEm2UZqNXp0CNYwDCQrDFV4958vEkkicya
JzR4iV7FiOiB8CBRIBszseYO1HHunfHWS6J1sloFdnI9CMQRadXOTyNnWmVV9h4q
tROLMSzuSoJqQbBlJzxIopO4/NEJtxyx1W4r5x4VHUfPVHHktFaJoNE1wmSUXBnc
nGWENLW9JQLB93Upj+cAu6DdfzxFAHEnS717VnPXi63kxBGNfcK+VxwCv4JASFgw
21lAhsrVD2QzK2ugjmcg39ypk0J0YoeGUyPjr7EvukLOrt82LTi0PNEiGCrFwspX
ih/egZXlTLLcbg3TnCmHNUC6k6u3Kt2v7rAPiaGBiIoBStUpnj2U9DYqrVyJ+gr2
hIBVx8CRE9ZNONcGKr/Xwc3DXnGKvKQnGPGHj8Z20uUZplIUDSrA8UYZe/kq2ozy
DlnzxWHaXYGur0QxNoX2ZlOzoET0SVsOvzhiL3Qec8h8x69y3noXiGXk35Ilq3mK
LSaLtybmsI1v+l+Vuaxe4fbfHaQYwhA9ajcAeUVOw/VJwTyKS6xL1pwxASx8Z27F
7P68s0rs3kU17pI7XmzOVsGBmSH+IUMazh5/9koQ/Cda6KNPo1yN6YM0iqi/qHAs
rLuHTFuQlYDHnrRMRYj8UndxLQjR8/R5yUX4k20hpc5Dkkp6ZKolUKTIBcqtgMFr
wShVukn/G8QAHpaqrsVa0infoQ4lh6y5gGJ+lOAtoeYi0LxC7Iex9Kr7nvh+DFO+
hys04Ge+sXPZtXF1bbia99MqYUd10RQS/duOVl8NUzRDcjXbKwOoe3y3r82E/bh5
0AGIitHTx7EgDROC4iw8eGAEL2hRc5DUP/q32sdh/4h0qSOy3lkZukXSe/2mN2/P
BbULf6ypBruaF5mLqH6bQwjSm4Wdn95xSVGKgfxw9m7A+7kr1nH0gxxCC2cRPEWB
3b9l6H7zvPqL6r0SJmHAUgYZOKcQG/YWxP03dec+IXh6K4fpHecZK3VDXKUxztU5
1iKRxNw9DeWwSGwxyiHhvod+YQK8e+YMxd/CsKMl7iTtgd+ZI0WpzyH1iGS444TR
FwxOcCIccmuUzwZ9l9Kub1a42rbAO2ykfccndPxI+iZ6bzEFGkokQuSMSlcpqIU3
ZmNhs3kfqyXULJTmql0Milh61TUCoxJSVOsSw1t8osOSgZGq0aUdOeMAC/WQFchC
dOseWlH2GTEMFrGX2pevf8NHIzDWAvG4xhxrb0TKgQLSeQDq1C3Jldxr/oc1rOFq
6WN0O6uwvSOYNU2LDBJKmjLWvECgGNT4i2CINRk1tujs54MN+bBEbtkRKU8Ns4PE
PABkXjwmwvFikUn/1WCqBumdrvOhKVYj5U1JHbVAAtjbqkIumTmXsKWYC/jJxVjj
626Hp6z2upo40LlXf+2RhOVN6iBRgDxSMfJuzmNcPuFY6gcJUKgjdPN9zl3kbUBj
EftCgRN0anekHNOBi8ylDs74B/HNqrSsUJV3+BzX/yCAClTSRSd1/YEYL5THWugo
XFyKzvYvDkkwiQI+XGoyoY8XMTIO+YvlJY0CM6OcdDzwJFSR292IDDHuWks2ybWn
nuSnRgBwSGkn1AtrvG+PmlEV1O4OnwOJeVbHZAVSV/nfDHrMWBuwCcXTRGj3OlsJ
T0liZ6JnQAJGjetIzWDqoW6YP4gViv92WzV5/1N+0iLBKx8YtsxIDJ7Kue88Kwc+
j8BicCsMOaQeu9pPp2MSWFWVr92qksLJtaBDhI2I1hWez/PcVybkXK3ZegVJiHD5
jBaKs8us1CvTyirgs+IGPL+K1415VdyyHY0CAYxnljE/rN3WleYyq3OGmwAjS8pZ
xvlPYQpAC8E+akH2XLWS4zISmXesDgw/tq0iQsorWL3YpeIgaNvC4BkGdZ84XsAv
Euhg4dMWCOJsvCw5wGiBPDfbWvJHFRvozFrjewvZ1DwsWNWvNcy+Ch8sqBuM0sDZ
ip5bJOBhdh7x/3vmokBHmP1sBS86D4lMJzQ7awCZFyGkPPe+ymy33uPyiMeeGRtk
xMAQ7v/N8TTqWU2k88n1URgovkJJD2WDKGpH6EXxEGalghUhqZa0uW/LakzqVGr0
C6B4JAT/DofGf9cG64poEuACtMCcuCOgs1GPddk7EeEXmo52j9jY8OJmhUWqctoS
s2t0SUfT78gNOL3jG6x4dgftqw+tEjMpHIXIK1zKVEwfUeQAnDI6v7aPKVQfCJ5v
JMCy/z8yzMOxJxK0mR2mbAKLUwG3e6UREyqpDxcDSWZw06vZINV+3OGCxKdNwm/3
Yfd7Vloms5hWgmtU2kHNvzdU7BjcXrngvxdrw+AleelxAo2P7rIUvSKUZksNKL9s
vj0Dua4O9BUXmr1vuzOOd9O9Jmte8H790gE/53rqq0F58MBxdzeNxJq2+8sKhsGm
nB0lQGaEzwj8CjgxMyMCYN6IRzk8E9/2ay59iVWt8Yoym2qDrckcuVkCdrQlWnch
B3n20U0zQTKe0LL7fRlKghIs3pj6nO+k9e0JPAdJufgje1Fe1YAr/qQQzlnfEmaJ
fQuLf5eMxRdJxidu0mCdDxyYS7grhfQ6g67qBW0P7gI6a/LldhOIN1ITcw5GIsOv
H50C3XoMXmuwzCv7YQxlvjrEYWCO2UHuCwICZpi1mwP/zr442lslLgWfBRwqeO+2
KDow87ShPpUK6ZI1PteZdk3aUjEP+piPaK9toRtkIWpRfECTt1LAtLgCpGkcpw70
ng7EiJD2bbRRvIuRWmfgIsfLLFPEGEOi0oAwbhsGVNOEIiuI32ypiEgmQZAbYjJ6
MczaXEDQm2w7+AldvUgLGVeivRVMnrRBC7EskhZmlnS5bSVb80xjNNR94+HuNlLB
FZFEz0rgM03uYej5xk/v/SV3P1tpMaFKLlEAP7xY0TSJ59PF13vKMUI646D1406Q
FtlF91IrMdUy8twiuB+4O3VSl30qjE3YFkSS10n9wHHwhNtE2CAqEMwXZJyNPnRd
3tWf0Qfrw29lNX2A/4uo/oG2rA/Cg5RlwG40TGISl2AHuHU2Vajcy9PSQyrkVpwn
mJxMUoFrHLUpUnrOvr0J6Sv/rM7ZrxDZpxlp0/6W/w+kzmpTuPhia/bKNttw/uCk
iESonTuehN6CTcqByRy5/YvpMoqp1TjAds1iVljERiaeXsdEKSJh5pJX4M512n6z
kKx8rZVDTjmutgtn4LYJptoVbkCSvVLRL/RS4ROmNZew51U9Z2LIk6DPI1UoS+Fq
8CWkTMHUTQfekzzn+OIEICfv26ZmzH70SEuOg7jzrnJtomsz9mOg1NEzixPjpydA
kDK9Hk9tcRWKGdIFbvyBkfuIsdwL+xXwPoGHJ7GDbBwxvGmorberLubQURpavIuO
r0eYt3K9Cxmw3APrl8KzgwEGP6Lt+NvKPlWAVzSCRPMTHKgkfpLD5/0UDC5tBASd
lLUWLVPbN0S60Vnj9Q9Dn8v/IVSu8n++nHfaoBFOzAM+i76ekjhfyF5OUa9d+HoX
XYUA1ocppdNq2ojBtYwISs6lCqDAtR2Xsc6rm3DbZ1MLAXSVJpzwpyyG0ULbFUCa
jX5sAdBhBNKCEwz6A5DxI9JtO9Eb8Ya1ZkOqSI0jxroJM1fzzWUFXPN4uMtJX86a
CK90ayFab/EDVH2be3ah5LKoKyRXvf88F+9pggL5p56nz5R38WpTNWYnYz++/Svs
nFhbLU7U03ez+mJWaFW7oWgdrdx7h7K5ehI6CivqKqXiSAjCKp+VjvSn2hQZj+UL
YENgzsnOVz1ciE+lmjuFjvZ9L2chqADKID9888/1pg1IEHCyPbHfH0fIR6GVINOm
OJm2m+4t9dQ1N3NzhKDXvjbMUENHqfXYzZ0BKceInvD/WcfskhkQdwRuCx3zJGat
HYCViwRLURQWHGTBKSNxIQsm9PpWqVaS1Ws69Z6MNDZg4Jp1vfLn3Y4KuLgnuYSf
MDzN0tRmDUtec8GSPHdz0Ilbw3mpKWLpr2bm4rSBhMI2d8q+Tw5B4oijMWBBZv9f
IC2EtIgxcnbmXvcQd8YsiGnQhe1ThGYsCkeUmca6LdlkWN3bvs0V8ISgA3DNd7LQ
/Qcpuxs9pMSzkSiECnBRS8t6L9tr0UAkexPppto+337ukPtZ7YdbG5ghEwiKy2Kr
CwRoFLCaUVpTARWF+T1VQg9RQXdWpJttJnJoJQPpuRGxAWshRgpqttqXOzYQ3rG0
8dxdKt96iCOobHnfGDRjVNSM+QSrs+071uL1uP1jjnHlYqjN21+vEizXZw/dtXQm
uCT3y5lHxIGBLyupjtTRtrBE3GxULnWJL98W4TvEY9v9gpE9W27AINJ+DrqyRbpM
xsu6t5sfem3GWXP1Fx7Wbmh6La5WcKnI9LG4eXPmxAkKH0vl/nZYX5XEWWT+oYJt
8fOG8YBGvVr3UMLaPDuJvT3iwPShTzgIritCWIvY0eMkh1HigYBCTHPjWcczraZG
7iNG4Qfk6KG0ACFJbRkpBPr66gZcYsUCAHHeybUed8PAOolVfzZYuLPkJoFetQ/o
wXoqOv1gNrAGhEiiT1JX5AXS4vjdvWy0Ue0nLngiks22hLBrspHYElE2ALt/PvNS
EreAdJtFw5tOPvf6jQm6gWxSwBiZ2GOMOCZRANR4sXoS3n9tVWdijG7KjBuGJSXE
Csp4az2IyMEMCJkUBEAWHUsPHiuV0YDfjCmO0XeEoAK80/EJIPfpuQXBu9fc+jLM
8t2Jn8tYc1iffLx/3HDJny62HksHea45favs9K70rMlowh3IDUpKIpF4NH5t8BZu
1u1BO7U2eipRUn+6rI+L9M2AnkcpWSq2ez/oI8MD9vwEJgSZ6LeqzS1cLNW0qiyU
qrCsyuJVNcwCp1FP71lR5xyiJB8h+0ri2dAqV5aB9ynpBAd2aVyzZudixIuW3qaN
58NpRIL5am9HXgqKrk5GKXuIIC9w6nW2oRbQZQsSLQ7FWn/Z0KWhk8h3lerNkzcI
vURAQhx3i5mywDiX5Qu+btQN0m7G+za0hTG4sBXC40/hLDhrXLAFkFhbeJHW4yr1
05+OHIo51KbFn7AlsP+7tHG7XfiFg5KkXn5tYYmzInhOio24CjmRPJyeIiqLBspK
olJR1GGFbP5Vk5LHc+ZeYncnRzLPUgzU+jdf72MizJbO9USiX+jMRkLtmWfYC1r1
KxljI24bQorimBjLwchnVN9anLBR/gcU+YcVr2IhN8VqaaH+rJoWdFK5ZABUExxe
D7+3bNae9xjhP5aUfBsPOApohpwgat8K+caeb/pmn3Ty4zsuYCVqYsoY2MU+gwm9
FLPlxCMt3hGG56J3bkbPZn/+XCNveaSYPj+qC8XwuJBVuh7Y75obDw+GodeInvey
Ff6sPRuuBUIN6YX1ZWDOJkLaFMJr9B0nuTwsJnRkCta0i9KT6pN0u55/eY3CF8i0
niQO2u/PRovGy5kTYVkqiwf/Zx36TtL/dvIvn1Bw72gVbn7WMiTN4SfOxaH9nDzB
D1neOxFKddOCDUTipXKf006ybBT83bs5KnUcAXRvn18lLj+sbEFA3xCLLBt4wg39
zMGH0sKIENCS7BBzk5MGnFcKcoaaZE2DkZxFQQ+TXAb6KOo4fnlgrWnrRpKPPYjh
p4UdsHK5EMjEwFvhAcVktJf3xbsp51EJKFtXgDv/Tr2AmKgnYEfUq9S7LgiHaM5J
dy/8+LEIkyjiUguVOERaah/MjeMRXhxkFhGLfGqZ68WbJQsnIdmJotcpFak9/OUN
AaYzDDY3VtMoc+Kls329gB90T7Hz3iLLXK5jSoVGdzQRGOOTxqlgRQHJrgn0gA/e
CUpsyzdXLmWcgYhuYaM/cy3gHVJoVNVrElKt6p4kqWYjKzQVHkDQ7ZPUNl28+A0Y
AliXqVW3IM3GsM78E21gU5U6kNqCn9wBl6N2G39YuDEAs802EPbgMmtMZ2jZkVnB
vOXw0ynfJJIDnrrN05VTYfPShOXbbH98k00AoXkxRqBmiLV3NubnRgvEk/4+BFTk
eeqrYF7aDR67AVHbGr5ttMyzPh39miYqy7DKqa01qxU2MsSzpTti5FoT8iVRE0dK
WcSIV/L7uDcKuszokh46cd+SjgJrk5C0e+yIniEc3+gfReim1sNeIIXw20mBSEPk
mvp1l32lVgjrR0hA+ZUOVrqQYv2Bn3bTJf8fYaNrcQ87tGusy73+PIpYrPpnQ4rT
HCNjPr/y9HU5XTWb3oykc0tJT4T7vYMVluKgxq3JS2QE4nUDuo0Rvtwui850yTH8
rQdUIuF8LRdtOPyRqnJCkAkjPS9YsrQr6FitJb2mY9fOtTcBbAbzPlrWB02/hTXH
3w4dC4rRsUQ9SluJvT4LBdVd5ImrANDHTCB/AwuMkkCoy8znTv3G/+Z4LQSxxmdf
dB8dEP5SQf5dUJWpwbDjjCmE9qlQjhk696/+tLRMmR3acubNzkW66ay60jkeVJZ1
71har+w/nqWHrKaaKlabCnwOJej39bj6rdFJ0Hx9Oze9WQ7BMSe1DR5rqg8aCEPB
peR3Cqz02cparPKSY/pzUNOhZNWiUmAoLjW6sscYzt/MrSa2MQ/iPuL2yOiJ//is
36pjJu224Q/k1G3EFDg1Fn6vFoaMtD40dOrSaNbymM2KzLEm7t8s7ZBP32CgyXdT
WVGdfBPP/Hzuqd0hbsByXFq3Pgbu+NFfWulWXBzd60HLXVSRgMLZP08gdKi8j9V2
8wWtKP+TUqxW2J8EJh4/CH8MOIcRMcCAJEZyjTP98ei4jjLl8FsmktkVd2voPFjb
snoTWFlyoRl6q1K3oy1gBC8OnDQZTanpH6LYb3BuQpRHqQ8HzpTI27slHL7fIw9k
/x3Spe2eYM8HLUHkeLX67zXnMm3tNWfEiLlWu2apEudGndTwIeODFR634eUiBrzL
j8GlJ5XoaPL6CJFfNyzCzBLn7YTDifvk8yUr1tm/1RByf71gwd76jyJVQYj0iZoR
yhWRQVxrhLY5Na+SochDRnBmHve3TAusRo7jMvgZRUMyOkYftvPEenYUsfrYAB1+
r4/gU2jXHm8nSVdYmLvpTYqj4OoE3g4lC5+g5tK3A4XJzz2Y+rdF/+bNkUdDvZ8U
+avIvvjyvu6lFPH2iP+f0e2NSAMwlGHU+aB/MJ2XPVskWYwaLs//UACUfCkWvRZa
/A0DhxUa/Mtg/ZpiruWXDylmGpVkpE+9rz8zLh7y/kwDufQCgmm44ZjwkBbg2AsW
Et/cj+ujQB7zTvxs9Wzp5jw9ZBrS90bioxtxnqAMnLnroG1W95AKDOfgZPaasbQs
cqzGrc/JqFTbaY6Y7MZxrESuY/mpV3+rx04tXmgCKKoj8kI3tA7grqe/QfAVM1FG
xuKhRUKfXhXukTUUx/NSYQb9nph9ObKYsImO+WC+XIrZF2RA8OGCPmQS9e3mu+7z
7eFdbxqhBjy+jZYjp61DjZcFqRn/aNU1xFBMD22HBPNU0YQueBZC7VMzNiKx6tSG
3Bi3xCEUwHHfYytZJmau/YlVTb70Az5TGDwk57L7OqcktNsPd7KwffG/u+wsPlDe
53EHVAJY8I9zwyQakKsSAe8hWNVQEidH3Hq81nV5I4yERyuXRZCaYL42mfKosSiG
8VJnYXqv6dLimtjdss/olYDXV6lCHKRzrfFZd068YzY/EVe3oC7cpj+MVlcxIL6l
gHziSVTMJOmW0z6q0HSh8TzBSxG39fWSiVdYOvZUPLA/wPiwxRE1y5OGHQWwaeKD
e12dxqcdcmywE6sLUxtFhUsjK77WmfX+4CADhg+UhBoumuygsoETy+DL/dVsBH1Y
jH54siTI53cuDjGx5VhEn9N1TBSv0H173Sq8AiKBaEzAppfPXLm8SQRFI1OnAGLg
yTVfo+1Dpm6NdsalAZ4aUdyr4MEtF/mzNlU9WCvf5mraUXuZQ0R7XYVs4nXn608H
2SQ9AOcUlnvIYZP/N031bFoOxQ2VN1AQMZAcxUQ/B1Q94oIFetw1rFpJn7DPfOhg
IXKvZBiYZO2+P4g5LfzLvAWk+6LNm2dqOUOpGpzlBgtneFj+4Os/rB/UYB1UyLuv
zet/GMhpVSkzN0PemSorPnYG8UQUBcZQm+nt+68jneXJUghNcMKWIUabgcxtXKIy
0ZAwOz8gaevsUCq4RP4AekM2/YGfyvP3Dw3HZ9D3YwkTpTx+KdHQaTX99i6Tn3ZQ
v3HX6nNqBL30JskVYJXW2smajca5fCyJIp0Fwgvjdq6LZn+e2iHS0ROAiPVGOR1b
xNe02KWk61dK7k+wn8qEV92vzpaFp3nWlpyTcbaFxUMtYKYhHBj2jRgGIj5x4rMy
4+isPo6IPPrjmuTQzLlf3Be7BZ5qNN51OWkkDP1F5f8OnN64ym01LdL7k+q41C0e
Wn1XopwPpSyCttH/SKN6lbul1WahsocNSxwOA57Th5qx/paDPia76v/2B9MyWjRL
zxX7Xwx+zROEEs0bBh6XfrP5PVSQnwQmfC+dUcBrU0UjSJiUVgDH6vPXmh1F7iRZ
HUAo5kJLEgcbi7+NIhsGTbntzaVsQNdpJLeVy5AdA2cp3fb64hrONioQ3MbZztVR
k9wg/6cWOq0WhFV/idN+F8X2+YzjNGCf18Rf4m95uWplr2cX0iOxFTKTnvROk+yd
iWz3MvxvqtJjteL24M6mXVBPZnDGIQx1S9XuxNRTK6RjR4mq8OnJ6GQtnyLScwMT
f3cwgLJV0rR/oa0RVr9xL3ys+sax9+oeC5nxcAbBWsTjVss8L2zlXXcBxUNdiR05
KvW/WfAjivqVrlya5/fQJiqaZE1z7itUAov2pLZpF2ItKhmI5ej0wz1JvGH/XII9
5bYSjfdC8hfcdx5pHDGJfJtTySarJOGAByYG7MNRo50moXMOaUDMh8StxNFiGxju
ZuOg7REb9TbfGDenRnThimkkKmhfsC4XLWi5lDfu89u5WGQb0gw5tKePEs6U9ybs
ogXrlarvn2pe+Oc+pDu+gsymNwUmkMss2uOMutXOR+V74xGyD8y+BUwO0X+/j/sU
Mer5aiFbBNrTHR0UR7lETWNt0abizsmKeJnU8fCwAvUZ5JyZobrbbkTbbWk6UX/c
AMAs2XIkHpym8GNn2c3yMhYMTWqJa44D+1ALTqYUh/ALAhdOz0aqjicWbAVlBTli
zQF5ItltAcJC9Bb+ohNBhjBVjzx1DEp7hheB+15EoYp90wamMS+waZ6apmxtfNUf
GQg4FYyB2oofzVc0yH3Yu9OTcn6H4HJ5J5mt6yWugr1ggNMZ8oUVYkDGqAlsjSA+
UAqm5D/TjXq/VkqzzlVkOitnzq3rp4eyK0I8SzplYLJvu6uHp95F7phlw00+3N5H
HhYqrbUneyCA72w0uGtEBA2f05QsFiRhJN1d1RA8A+yrQiulMm/6l3zyky2ccULi
v/VUKE30VxZPBMkOwijxsrFySNy/h0CbDmLyIUlc46lQpd2CDyTFnv09zq0BBvA2
9rTzuvfOUCfJwezM0bUDNSFhDpWalPcA9L/uetHb5AJ2Z24oFfRP/AN9rraSCfaX
DT9ojl5JkW4KbWrU8ApBdL9EdJcnLlZ/MDTU+uLMJpSAPRVSBQprqg6zmZp4xHvk
S2EVEgcAVUSjb7jLzY154jYisyD1I7ETfBIWVCHwjdcuOBqdbeDwlSUMF1EsujZz
HnwFC8BAMD5oDmXUT9uXtjca4dDtFKZU/0QunVJq2GYcqEOrimyxRGWRWoHYcfxN
FJ+cIkj/TqjdLZy0XF611526HXYVBY3NAsWJUqY0HfQKv/EElqMUv6yeZ9wCYSQq
8fIX2U4UOPyf/vhZAZURNMxbelTR25vQk/4gJiw5GbUycrFePL989udKDjfrHLLF
FzmbDv7y2xiogKMS+dzd61UD+fH54yVcs4Fj15Sj6guAUDwK6B6fzoymSJVEb/Of
wLy4tUaRcNrzxIHcHM34myD2xryyM/Vh1h4IGDcHcVufmZukZcVLxH9b9Z6/N6L8
OmAqYRfmE/57W04rQHxRatxpm0JBtMFF4nV/D3KD3/E3c8oRb1qEOzu4L2WJ8KoW
vH0ZtK5RtPP17P6H97/XgwXDAYi3JjFsDpWyA8NSL1uxlgCRzCwtq6yVZ3QmCY3o
oo5DNEbTeDirm+CUwsQ1i5yWjtkCImjidflOeemTh9DqYvcaAtE6UF1YbDUHjIo8
DrlV/P2H1y3RYVWfeJs/q0+Adv80b1YB+W/UwjuPXKOvnBOcpbt0XATCjp1uyDNo
Cbk72htBSzLyi2juDWuLXE6nBT4kJo1qDnp48urG2CRTy5hFv539AK+Du/pb94la
NDWRRq3bLV/YuxR3lrJhfpxTG9rPspH9vskVfm/88CQfU/XFluSDMx+npY6PXiQg
Vje4tfZ4yuKqAqIldq+VSAKK1RnzJEctZHQPmG4bdoVQP+Ju4kzEAI+nspo4mIpB
VlPgldvgiK4SzqMXUg9r9Vu7P4Dl420/17/SnvwQ/j0JUiXwgdC5tblYDpXFcA04
+LO7ieYHtqwdJ8TDk6wrv4asnTSrRTEc4NcDN9ha4jXLoYIFvvE4xY41DHUKiY/y
82LR2UL2K8IdoUtOxF4PFHZMRdQ+6L3M6IEE/PBds6WS5d8ynLrxIR3ZAtDJYSID
P13/H/MN2RDYcuX0+RUQEdIzKZit/3AhF4vJw6cGPdeEfVwBWN/XGuJZQ6EQMJdC
7WFUQwd+RqGWRQWomK5j1fWP0yFYn2tb/oIBGoMqNkNXuTY3X1LgFSqZHk+6n+b+
HHtGnYs96QPJpn+fkWay2j+oyCkiHAQlMZqdk/gcqwGjH/g8t++Be+wM9BZ67O4B
h9KtDjoGmj+Ag4rTomSVETLJuYhu67CR6Dc6Q9jGw8nUQbL3O3JNP9OgeEiUlzNj
a2mO75ZslJhrZiWiEFk6dOraiBenrHMq6meKZOo0Byg+rs3WHJl2azYT0ZASUJ8z
Vvc71ZFjrLzsSTP2P+F0BHCczEBRNfmuB0q6Mna469/gfwdSJD7g/KlKqiGomI9v
oPjcxe23RCtsw62NP917BIFF0j0R1T8cUXqqXCu0kE3EUa0lIeBRU8XkeGaveJou
bQAi1+dEGRSzvaY4s0aj9QCuTz5iQJ0c8/hKi2WF/pbSgGACtkXbuQ8GAa8ryFcf
UlP70B4nPFqWUlO91P5A4MyGQLLkVME2vYduh4zvsfXb6iQkZb7ccfQsG05QsOI8
4zeaVJXuT+6kVODP+/a5LlKBFT6dyiA3hsXqGH6Bhw9d8ml59vfBalmt6efZDU+8
35vHzMQi6g3x9HTCWAhSbbun8G39UtBAi26fbW2HTNiaxWEWCZMdBP1GYZCDQPrF
w2QW9HaRx63rmGMurTjxHrBdA33BnB6o1eIzPYTbylSRIAeUH0/QXdTwa3piNOyl
/hy/54CuSm0Qq0aQt7P4OQLeqPbaPTBlVNtPeQXg+P9/grH1LRX/qm/9CKQ69wwQ
Tc/vc3jcbIyALvbYyYcZOjnsUnqXZhlJ9xwzh8yuLOX0bhSiLgeaWXmjscSadCxn
NdsIKjX8rCDKpMgKIN0ixMymmptdo04DuWLcwcmlkb/f45d0YZzoEZr0OuyNOyzS
POH9CYwCU9VC+Iue2hCX9PP5qsbQlSHiPEdbNMWFC2rKS/Owy8IMSnaLsNHLPycN
+d7XqXWp7H9+M2g0sEkHB9lZvYazYXRpmxTTW7ap29HKGAfx5FOWhxmXvDL1s8ta
FKrkUnQzTz40g7QkGHGMcAiSx4f5wxFw3gVXLWotTV2xGhVH/+qsMXr4ManJBw15
OeqJ2a60sGZLYzopjHpu8QdGOiIlX45naKGcu1eTcmoYyGli+LA+X9qtjaP9RP7I
U9eMvQsftnzJLXajVtfTRhFUpznARbvhaw6w4hE699Zsq2ijOprVkKb7u6N4t82d
9e4Ifeqnkd02x5QIqaJ9zsApoVJNxOODFVXXUrvx1p/9knToB2sECBrWc2zmFZHg
q0DPnxeVmEq9tQcUtqAbWHilnFNDsFWWiHNjEHu1IZ2O5Y4DM7qHQxkKv2wlj9sQ
xWpE2UcB+lq98x78LeOnlj+f3RL77PGyO7/SwZBDmijMp6ovwIXx4VJOvMe7pCFs
RN30O4qCcUebxu3tr/sCM9gZ0KB5uXgb/4UZuIm1jTzHbBvVKSxIU4ypGZaAmjeq
68tt2tW6YgRexKeANQQDwyA99yTqwjR5tOGjDgECOxREnfylj5k8ELAEYT2LqxIs
x6A8mwMhMArm/b5JwOZ91Nglc2p48jwjV0de2l36e0VSY1VpUwvNdiWjCzFL+V+5
+/ZnIxcJL5Fx9/uycBm+1059T7t2MNp3UybQP5dTgx3ZVfe+HSrLqtZl12T2B/EA
pQlotmsHV+Q19FYp3sqNEax4JOo+ritnUPClXmwNhUxH++z7eD04CkuQjnPZr6Rg
6/8QnzWAY7G2yRaK3yW2FYfJkiGT+XTzhDIWdlAqDPaXaCIDaBodlrvLpB2qJu6F
uVvJr03xw/rZ8faCztON7LF7rePsYjjCTatdPYnlW6llKa8c4VusaE4y/nVfd4Mf
QZHxWxr9g8qFW80r3ZD+sx35dr+k/HD41ora2OSZ//Xib7ycy14uJMy8GFovB/po
akzvsJAcwGLpn72iNJKduH5yfRgenJrKemP7eJmaSFa1CdAGH0uISswEOTSmlDV+
zXGLc4tXiNePOLv9yqFu6RlrBglhhZTnyiNsJfRCtxajeHaPCFeuyBIZgCD0N3Pk
ZyhjhCy6XcHS2EnnpSjw+/WbA2KYwxsHFWU+9NjHLvC+qbiO3qRUTOIy+Z1syWPg
2nxGRyIZXpmgGi8mlwrAAttdXE4z7o+MqP+1PW6Bczrt8c+Zmn5z2hw3quJWTmXL
N9e745ap3faz2t9rJqnjQvYsCfKQlKvAz3u9nGOsN5UlOYqtkiZ+an/B60FcPDS9
r1cUrnetWruLV6H2VVAPH6/KhwHq8NUFpjm+SjAxXhhsfexngrZt3OY4l0i1hQXq
ja/IAFV9AbY5Br02k9F1eBBYQXjnrFmvD1LI2OyFsxZr1PaJoeoHWSWr31JasJof
EoGrCWdeMKPeiyROlBtj4RjyNYG3oDSQgK6F2yv+9LCb3XaDL4JInS+1UVa562xt
NPkM3uVVoorE61BAL6Pg4XM/PF7IF2vUUhZ3qZQD+aBzOG7qk1c5/zBj9WjzZytm
drUznfYnDyjBqi/1IV8W+JfCT9W89P60DmIn6WkBe6t1xcvM9r6GdqnTnwFWfGLG
mfvlY717ltmNth3w/2KrfegONu7ujtvFQK94Hcv+Js5DvZGHYifyvErlzcYR6rxY
VoMO/0HU9lJqC474XLBfJKXHIUocPPQJApfMqOlp9xeTi0jfxaxrl6Q4QRTkzdqy
krJm6gn+Avxju8najP7L+94f5TYqPycbjy2bILvm+xtAi9lttsUWwAm3YjUlbCf0
LvW+wNlZIGZF9V54L9/AxUKvjs2CtNeLcbE1a38GgqZXJk2mcwa2lE/U/Fz/H2zF
bA88khx6JSRW0wytf1JmK9+DOFTC/0kGdMGGOGH85l/7Sye30xH02mq4RlWXiDSt
4H0NC6pS6XbvZGxH/t5MkhDfWP00lVNde1yXL9+OUfuNnCczjOzS2/9aWaHJ2sAQ
tKIuj7q438ptaJhDvM+CO5pi3cyvgQDZgPu9AHTucmSvOZHp95k3itc0oAHSvKnR
DmyohRy9rNMaXPKkKCtAT1uQfq0hH0hDoRgiDgVm+fKfj8mfVvvg/oHDBG4JJUcM
shT9HCWPf9ub0rcLFBDTwxRq7Ajhz4TBxUjLwXaf/DjILf9ZbZ7oUx+aqGMwJ+NU
hEliK2+OgntoO/4VL5EQq6a98nk0UzV9L1grRso8K+BGmVOZjh9UcBjminMQgcWw
dHYvuDA91NHPit5zPv00O+P/XXuHvpNkgMPKMjPUE8YK1TS/hAUG0H8DsERgz7ub
ZJG6XY/Zl560hA7Tac4hrvxQH13TZEhk74oplGo/AVhlV8ii6ZVhMks9nmTxjR6R
5FZrltQt0f9WvYgM+rwFcs37L5nC+/1evIIelRM25XjtJ3RICtrJmhxBmr2nU+w0
lwg1MT0biLx/J9OQpqPhD512PXa6xPrE3XbtZWkXEEK80osx7zvYCwwZt/WPT1TV
EQOsdz5fxo9V09VWnIS0mdIXe2v4f3Kmm0Q5LZ99Yhj/Bf808ZMOIoCtwBXjrh5v
6QfFYiOa7a6pAQRrzGAN/q9Sx4SoRA3S+V26eLm8du83mCLpADOUdbi7nrerk8uk
/ETmQK18Qd/uerSZeX4PWq/PoXkag+z7ieQN615wXTEC5O1qYTWCZRaioF5B+scE
LUrEfWY0rWuZWPvhtq6dV72jBuX/J+aBRcn04WBkh0ryGPv62jtvSWmlv0sNGhXY
ZNeOj3fiVZCb8hcVaTMq5VYoNSOXpydiwPvWncmIemIxBjs5QSwh0LTnrBc7AvZt
u1Dw/ff/OJBBvFx6hm0sjPOEyanKKHOu+zjuQzLTGsd+Ea77OuCm7MqmwCCZQM4k
DYLB9TiqTcmxJ0q5siGdyoSxSm1iO4RIeQgtzPPscZlGYTRCKe+pVkqiovBuc+F9
NJh4Stgeqzjx7yOvAZAyO9HBjAlNuy6t3RlBQGFyjN7b/HPtFm9G44cPB3kzVjJ8
yunetrnZ5Oxzt26jYp9/3pBESpCqzJe7l4Uf9xZ259xFSVNGKUU8bhs9AQkZGPyg
Ca2VKtcbvdPuhyAFPdTvvjTQPVZ1d4nos3jzCzFZ5x0D+zcppCeM0ZvmPB0Hb0oB
FPuMQCNqvXLpzK1MZH+sLfRG5IaKe0VaTTtI8PCNcQ2OafB07no2KOWgwkfx49w2
6eaMxwxX6ixbk3RyCz5YwPCQut2o5q4CwxHibz86c6G6/NwTikZbOhNRhqfuYRaL
C8/VP94tVCDiKMgQj1+wF/aJoS1A/YdTLtdmJ1o7U1GOiaTjZAA5l+U1Uel3n7vw
EjpAz7KnJjxGOANv6LDPk+HRsuX0FPWuyytRR8GlaohI0YQHDCtv6hAzInq6I9wR
vghIJvUyV1DwrkSkRoQpafW5lDRSzZOxHtXjSJP1Nhcjt1dDfPZiAcu/0Zgzkzq9
fWpF1OId4HmTAPdRYLWoFp+fWuIfsYww1fsZ8M4/Lx5m3v/x6C9X1LnpuqLsJr2Q
JQhD1ybTmVNtCxqRtExd7V3/vgMEjON+9vJvCGpzf+qmA5MjV+HhYkfcrGUpRCg4
Nglwi3t4aOVCvbFLlqVyvHczBeaUrQTJ7F/sENOc793DEOOhwSoa3aKdK4iFZZBz
LTz8FP+5sLumBeZMvSfnvPztqlmZC0F4vQbVhuXFtL0vhSU1BJTGon7qsCxOrzBv
b39w2A2oi4s9TykNfo/miuoWAfNHmaJQtqnL+r496VsYfLAHugdHc7Qa9EPVngFz
S4otju2f4eYWmAfI4VeKImryDBq1q+jLk73QlfYpfhzJ8mMX/kpLVUxyVw5OX3Pe
peHOoyYbobq6xpPDMEfPdZddhSGOE3wmIIR3ypAiSi2GOxbKkT2Z+GlilTXN9i7I
uiF/Vsoaf7uV5c1gEXcjupZp3KoAxend1/6xJOiESFgOnt0DUshpXucaMFKR070Q
MdR1zD3Lil2xcbLUqaoo1Y963o5+wkGAw4UxE9dCDofc4nQCmTjqKukeBWSVkG4Q
WwtH0exFca0dw1R20C5qvoR+zxY5LkNKAPrYNy+ihu62kWXhqi0r9DI0Hvut9XAS
KJiuOd2PH7S2ZlaWOd5I9fmjv0SYJxjoXC/owC50ipbkQmn47+Lzml6HQSqnzYAf
uTs4oKgTHQXfmVifg14+2Qc5yIuhqlejgpsFsIOYppjEB7OYF2c+WoMczZiPYSPo
a/P6j3OkVRwC3RB8w9Q/GOBc808ZsxJHUl//5zSYoj3iuCKKDpBdUqX9F9h/SuAs
tHphRPh0oKtn+/65X48dMzT+uhBQfbEbYsGol97LxrjZpbib3ZEjbDnO4CqPeOk7
o+ANkWD+tdO43kjiSni6HajHtL3BXCqzKDcnrCvGE9iqiuTXwItoZii3GXp0oqP/
b412vGwGq0eJBlL3q5Bir3Iv/CsV7XlbflZoUCF52lFuYEsnhjOB/yZNZ275p+l6
h6BSkYMf5JtuJaA7IS2Df278gFo7fkPwoM/2wGMj6/GH6hHn+S8fxkhhLF0CyVpX
1mrSH4gs2tywQSNG2mxNvLKVgZsRf6rx1zbuwAC+31p9Xi3XOqjT1Avk6X7igjxj
zwDd+qw425bbSMTixglAMyHwZ3e79hfaVou0haA+maevu4XyTcwVGUIko6gIBIMn
8zrwo3PdffFnG/4U5JeO3aYIOi+t97SEV32GB0wPt2LTfolBEbdB/uFUVp7NFtvK
N0MNodfCGoOZF0RjrDZPeEqHjD2TnWQVvubr9Kkv2S9ek1BEC7yzBign/aco65Ip
327Cqe8WutikGECA45fn2bX+6gb5N0ohX6LbJGJXzI0VH5vVkC2gZFcg5mmFXjnR
aUQT8Dx81hsdAm6a6Cytt3YNAWd5cytFI9nqVaVaQp46pOkK9lCb9V+hmiquIkvr
guxlTzLLeLmegCWPEazznitMN+ac0c7xer4Vr8fWeJ+ix7FUutTEhDLAnFxv3Nap
i/Jr4bXUa6NzBrrdh3Lvtftf75mXigO6mjy2DbH0YQMFQ0i1z9XWW/Y+SIstELz8
J0QQpBjHzcCwhv3dU2ZXW0BxXOB0dwLL9LWWG9sXE9CEszKgZ/q52un+ejaRLEIw
IeAgKrRgAtTy6H0m0T1IoH9gg+30t+Tlf+g5mRqmNLWYP4dVf6EpBYiTjwl6dCwR
qu97kpjXUXsdvZLjqaSgoViM6v46tlpFs1eb8ntEzkUlCKGStln+AGhQL4eNfDo4
DlHNaZEunEeOqqRhWlshSgqlzWkN6EBji/9dH7GptQpG/2NfUIizV6KdSvKWMud9
K9kbbGCeRMPoOtJwsGdGZA+QlmJpiNmz4c3tVY1gtc4vMsMkQJ91Z72QjzPnmJkX
CD/zO4DAyC8I0d+nvrhu9VRfuGCGvJMVp2A8PRi6SmpE+XyXzwp3PCpoy7L9rwtV
cKKmGzROIG+u8leYkXhucsfKT2BFzLZciSbrLFUTZJYyKIBRwItRJSxhB/nZlmTG
nItUK1tNcyUOaNiewPR8WCkhaiNuDnyeky6EbeUukFQlP1fbdU6JyLXqItIGoqWg
4QnQ6bhJ4EpBDRRnNl5yFOoK/xiCyzg5giWXiulNGKx6/Ppx4rn8GDxOsG5k+RXo
fWejJpi+uoeI/IOrnZazVGK4KTIPlbuLj+4vuMHHWRa93B5Pus1+MNgVqihaftZ4
oVXI7VyJCnPgyLYngynHbF5xm2qtAeojOOu3sSt4KX6uA7Vjxwy8p4H3zv29h85w
P91UMjPV2JPlSzOSI+0J35EoKXKHMn/6dHkTzxl+g99y4owT2QggjqWUSHUrzwox
VBtaexalJ3HryiLcFcHc5zCHYXOuyu1GBrxFcmQm+UO1XFx2n7kVrwSPtXYEm335
CfwmycCvHunvUFtI5MT1p9gl7e8iHAQLSooANny3ASr8C0fWBB42Sbp3+qOdt+wN
BJRYXX6v2zXfVrj9CAsu7jROUJGeVRVpveeqW+QuXcwCFNYpPQvo75YvZaajODf2
sBBMvwW8nKDaMDG2+2Nzu6oLhkbZeuMEzd4sdqnICh4JUPddjASq56DQHT84Xpno
op11VZfm31NBj4rvqolpt9IUXBCZV2ftL1SSnYpBUcjTuzC4rXKmX5qN5lj5Fd6z
jt/p9yqBUYVXQqVcYYbMS4StWCUqNKSnc6ClTDyAkvhJ9OhAJt4aNDEsZYUmFtPC
QdN8KIax41CkJ4X3ZHv5zncH5AJvJgQjBh6Th4e2ZydytUYk7UxqWH2pII/A2iuJ
AqXChuj3O03f5hcoEMjQqqfk/SZCNezNvs81wEfiLQEzXASaTPKJuu84xGuCiG5R
bAGVV3VH5hGcCm7miJn3G8IN9XD2U4H/bKw4FlVo8q2TnuYY7uWK4eB7ixGjND7o
GzdQyBO+byud2k+haSiLk3Id23meM/HuSNCmluOICeyXjcn6HpmSQOkCIvvesN83
PfKZKx2AeMh1JpuLdf041/rulgt+scW36xvRahKCM4VAYofjMycfOXlusLpPJAW1
h/+5qjSOI2VH1T7XPUh3968lIPLwLo9fIBonzM+Aiuai+l88ikk327a/bfF0nUjO
XacIuOPKZq6jsy+l4DRZhsWw2+LrsJFY1AlPGO17zesKp496i69sBDDOm41DJ7v1
ELQsISajmHma2SQzZfNzY4NYffjCTzEzXcQPeIcKfLeSs/3OdgSE/4IVIQRJjNjM
09tARRzE7aEH00RXkX921/EPIoF9m+LL8issyYGCVYuGcCf64Dp4vTiXUv/G34+m
SnSaHIJErJGCRNz1Q73DAztL909lsOfisdiqPAMnCatS+kXM5fTLK4Cr6xxzHLzL
7IDVgKtHJCgqXzxAkcPoE6x3JUQ3cDiLYT1cRprzjTkI5JowAf1Bbf1hH9pe8OOU
/WvE7PPPwxCYcvLnNe9W3eqTGez6c60SC3P0zM4kRFhrODiSGnJP3V7putiJeciM
Ce/V8OqMk/BBAjD+7hMKXEmv7uP3/fHeXnKpL1BfnerWwDr1vcdQqP+Zl47eBJ7w
nQmeKY8qJ6VEFVRhNn3YFWJT4mDvQd7+ZIKXfJ2KvpRcXn4zPU5a+CuZLAdojeWk
H7BgYeF5ZdCLhtwrDlGbR01U0hvZFlvDc7N1BDGlSLDJCR+8HwLLQxVe0yhx3ngA
p2ARnK/a9qoP6xMPusQNt2gv3in5qIxt4WQlnS+n1LJW4IfAYgkDeBQmHF5gl+7Q
0+O1VBXwvRRwO/slhMmViDtEPkpB56pmVlgyC/AYJMFYvuAcKdhzHca4iRZ68eLk
8w2QCb0U4Xl3Ct8QfgbR2f1tmdxkHvRFZgIlEnkZQ45TeFwGI3oHJRG3P66/RjnB
GHlQBueaNCdXzwfaQNSqqTxH0l0RmYC3krn7/02vMozIQEYABsJfJpxeqclen1XO
dKS9G1M+VkFlVzTt7+QDtPKPbV1hVLBd9uvoJEr9Y941GKTkICmOi2ygcC1xdfqb
NVU9VvhHQdXxQv4lR4UH5EqbhhOltpHkbqRqSGYQdKH8KgChhZcBCHPKji/3vs5p
aBNdbS4rv8PkE+WaBePMcAK3cBdXXtBR3cEulQ0XKhyZeH62SUrmtZYQGmTTfwZJ
12xiuWDulRAWS0rsC9HLc3bXlTW820r8RKzJoDo9Ju/UMzljFY0S4ndnU0DjcYeP
pLmenDk+Rfa6jTN8Y8ulH2j5zavKxhFTCSjaAKi9HXj60AG+7PI438Db+oPtxu54
CZ6YKkXWuzo/TYH8+s2ffsnsUgbL8TPwCWIvVn3Jq/UaoRGbXZgJmS2bQWscqyFL
gbQ69h39gkNG4n+ZRGORhTwULncbm9V4Dd9ESzUVYdPfFTlB65Fk/qYSlLFf5l/m
Qb9u6Mr9II+8lMVdk4wn5disIkOygK6qlRHShm/ncUygLWuGA13KgJCjLH0yBonB
MfdBZu0jxxpTDriNlfQwWFVPheg3DRhT3JQhyR0eytxNTiZcugKT35RrsSGxwmvd
tyvMwrEWZ4cDJNlpbYsDibdou3u8M/TTWnsizJ6CHYY01AsZcHv5EVSjrk4LKL17
5+xTCE/Ev5TKoKch4k7BvZ5SU1XH8q1Lk7L0rYqHKNnEockmy9VR45uIViQ+Y0BD
ROy9SyK9o51V/tP106zPlP3NzCy/IhK6sKgieshgGSyiJGoTHz8Ylu5ETQDtJAB/
hWn3iruqI9FiVKXXXisFMwQVs3ENWw1LUi46oTH+/D2P/JTi9X/SGIYKE+LF6VeO
mHKHneLcNVu14NCSPNvv91wAXTSkOHs3M8zZ262UztinA/uZRYLAiwer2Ha1Mohj
Hbjv/H0cp9cvbfIWBjDcYoIROebiKwFC8PzMf9agaTJO3AiIRue2JuMB6yQ3dHby
kGmPUN32sH36cv4/nhf21Y5ykZo7KKmru75QB/8ypB8CztMSlS/UPXqQ3B7aUMYF
dMiuDdIKvJOB9zMpzGiXjP42/OqhIQIlplhkw2H7M9L+URrG6eQ/seDRCHs/LXLI
SsQ81YD4TK/r28GF28fgBzEArsz7GYUO66cmAV9smd8tkGDnaKlAvYApwkUY1zWG
0058GXWsYzhEiWI/mWQ2n4VQmVHMIKrnRR++cO4WSTEztkSk/i2xfkzvFpBEAPti
qoPaFTsQzC8qUClnwQjZdAJxCE2CfNZPlpspq6lqv9CxrEKjUvcUABuzAanCem6l
cUSI760DnTNgak+iRScQuuY1xkB9gq0fIGil1W3a5mQk6+obxsT4Qar7xTq8CUbw
iaXzy0gkpbPU9sEH2eMoaHtNCc64vjPxNTPBywekkF76K+Fyk18QidqD7uegm0+v
Gp2WLNhs5+Z9CBKWNvim3VZaIRjwrbKkephOgWcPzmfE7wUDcH12tDIEGLPcIIP0
Zoi5Hp0cXO5FH/Gu1JvtfBBKdHDajJ4cxwNOaF5SAb9l1Kvt3uJfXVdmZy/HeBIQ
ywI7ia8DtXyRNTJdYSlLQmaytX63oVbq/rIF2ULSM9urZiv37FVsWEBb9ZNeYz1w
Tu+/Cz1Z5tx+bhSYtJWxtPfu+vBvTrrjp+wV2A9CVdvgGRokXQ3hitGq7EPFI2H4
CY1VwRjjY7rJ68mGxwopQjgeynB3n9d8w+NiWSohzzwmTN66fEq//qrHhWjD0RFm
0wnd3QyY72xvVhuNQ0cdlulu00UrdQ/5TT9mHCZh+M5v69xjnCarM+BW7HLGGlXW
OMoYXIb7zKRAhZsOxvTI4OPyGPkMH926zkb1HAXSRmuCln3N6h2KmgYwXkAVAcIQ
vBTOvyd7qB6trQve7T0yiAbU0O4/Pv3u2tsGyBT89Z/5va51Y6GGfRxH3QIyHlTG
0tgH/ki33spZ7odLIW2V0OJBLvoTtaE7yhEAby7A2p/loKqRMz9Ntia554lLk4T5
gDlQ/mLod00rWRBf+Qn8NdSq+b9zRXB4aL7WcYBcGL0trfDMm+C3HnhA5BHcdc1/
Ul8QUM9XThml6J+ywqdGgKsDmok0+NUUCiHOl72yVTepV4YV+ZiPex/WF8+9aObE
sdVPKQmaTtHoTfRGTlYHgrwpQJWpGK4w/DVUsyMz5/S05u8yPnixq8rJv3aJhwrH
G46B6dAFAhoj0cHsgYKjTPcYis1VHRyn/PoY1jP67MLNPrU48K5dgOjiB59Q3WzE
w5Hb5AA8ak9aVlCip6OWbJEj/x43nrcjNP92y+9sOstwYuFV0Z5hbaoyFl9MnqMb
ru61w4FdmmYlqDC9Wg4jFw/XKMZoBr6z2jz88sVoj/z7b5tCPMwXy3aaaUBWnIk7
ccK/rv//RdZyXhRIMqgOn40wKF+emK62yEv54bMz8EURpr9LdRWoVG5N9ph4JZ/O
/Y+3h3CHYu9+X/j8nUUxfhAgbbLYjhSpXNdLilLKBDgre2vZnAzfk9GTaMQc3Gmd
+i3bh7dsychjbcP6rlygEij4ziaEyo2ZBNh+9yfN+zOQ/vOApSfi93xaG7OeTrGI
3Nz4x7CMTCejzop5mOco6EJq3nbLJKYdNpmpun34ftbIP+lxoTvM6GmAOfbGgl72
s83FDp0gxhR6q8tQesR25yLT7fV3/0gqJnjZ+t2iIMNjlRGvLS7FIvJ1J7tFE1qp
yAhPfvOHRHxn/SaVgbtLH3gEQ2DcdT7zBzOynMBEIOP3huhG+BLp6DM7/smZqXsy
8YFNo6Im95zhu+ICi1A2RPzrJGDjJdd0Lv7pgLsM8p8oKLivYGEqRyGDMKPIXylB
rwHCO/Hnboqhk2U4w9FuiAaIjNCNlqtVsBN4lXeTIQpQHNv9TBcZlwL0e6KONVWu
h0P/32lueWSd4IbCZAKVR5o/6GMU75GXJ+Ucub4vH9z8zNHGUAYdlQ+e0Z1HOiI2
ElWUWwLUHvPh4X0aoO2j7pCBZ4pvGWhpY8LOKCFcrN+elDvRJ3l5g63hO1TCm9N9
AQWMpkPXuk8S7tLFlvQYuiH1F7TzHvkqR1jmsOF6ENn+28LJJw/uQQ/OU/te+13J
9SPZVQxa+SFK0EKYn4w79qDC1Ddz1n5JL5J7nh/bOHJgCuUMOzN4bV65V8pveSxo
6sFQdpkH0Qtg/HsvUwg9EoP/RRsyei52GOVDH327Y45qRL6ti2gOLwPgUODAGzjX
+5yjFgFaDp58KuErjPNwDfQ8s0vMZBIuHRdhbyNejZiQUQ6Tl8EKI5l9/q+QQMRS
qC+JH9tu153I2tp4ln0jwrejSWkBtbHUmujF3ZGggzboujyqthOTh6veRXZq10qg
PVXkgPW/Z050pIZDe/oleLbK+mbUVmoip7ombGOMgreKS1/WmX4p7I1Q28RNnKAQ
GALZzEgn0X2Sk2hQap8lZKrqYrm9KL7xjSq/78Xh+aFIK/qpzIora3aqC/qOosSy
NtDFoiTgB9BMBgeN8WZFgQFJiUVZAIV5Qqyb00TN3Fg9qAp/08C4ubLD25Wajdgo
kW35VYWJrDkalelNKe9XuefXZYKuZcagNPtqiUu4ofY+zdyxs8cVJjONk9OpG3UT
Pc9ZNqvs7D0QYiaUz2F2NKg7ojhppOuULii5Z/4EBGSKQfgY6wD/i9w7XzcOtzRb
wZGtO0Mqiu9NoRmiAmh0RBdPfaNp+sA9x8ulPCvrn3eu670fSqmQ9ANOLz96ZxVK
H/1zWvNtM+att+4Opc+1TYwBhjxcUuUFDca+ko88Gz9EnU1L/fI6+Cj209tUhjTf
NSa4NwxaFM4/rGzBYCq0yky9O5h833pRg07xXplcZ/yqzP8uvUeM5d5d5qaBYTBD
914E5K42A7H3wMcpf0yiEa08akO4gM6XmDbp1TiyauDD/4MybEgHabe4C9Iq/WsU
NEgE/mK+Zyi1/wA1Vp3kwoQPfarN4Gu9gdGyT+baWDZVHMAEHwQ88n2ZCIwnPx9I
pDFrM//L/1HfzsqosOqEVTHuP8MWhmkNieSJjlaYyMSTDWTLjAxsRnefPyMQ4PTH
ukHmEat2n8fvvhwdWt37+GCILMS+J0dWQv5Xt8ZBlNLtSlP2HMbsXlTRoevz/kdx
gr7zBlIpjTdYf8gdhi+bwTjxvJvDLhOmIySub2kk9rJko1hQxziEWl7Pynfx44iq
sXFxbIWPzN5jiUh9H/AUxCyyCNcfflItyPyZ+Z5WUrV8V/UrYd4EP2W74vBoBTPZ
L1CWBHFyv0rjLb/2rz1n4v8pUwC5uULJvRuvprmFPmwozwgxMF+lr8ukoVoxl8Tb
1BepFcwEsl31lYFUU475KgedequXUhhPhE0XHuOrHS1paJV0Ug937q+LgJ/yxYgN
nPk32AYifvz0++AZjMiKmjmUDoyFzgK6n8bFCfGKJCi9U2l3xy+jNRe4B98pf2t9
ZVjlMwaczwBMqRjY6qXDoAgWY0I8pA2pTbpt6vny6hF9YGxqh+5US5O9985W5z5M
8ty2xAY8sm/4j0ulTWab5dUTkmPObf1s5ICMBanRqxWH6fHlSLxdtTpTj4KES8fR
HbLeJ2vYQZYZp+KA4IpACZGnACupB/4ffFNpk9moB2Pkwznbgi1GdrAAJDAROBMc
ky6BLRbnxjpfwslV9gh9n1es/wPv0fdCZUs5F9ECmEBm44iqvu6pE9VJV4q153Yc
Ivdagb33wHjP9AUwYBB8R5rOENU01SWiMRb1isI9X6y/FAnw6NtdwasqaIWBxHUM
JG6fqT0TlprUP8u0ARWhM+BM4jKfEamnertSPhUmMx18NfEu0c+g6SrnIHlIxXNo
7BsGYez/Sag3n+HBlwpgvZNs/XlNjvc4vm2lIWFoTJDdpo/QrEGueK0fUrXKRLkE
c5ykgj9e77L2F0MoUtZLfA9wFca9jN2KTATJK7Zbq/EdVIySXNzP8xTRGGBCfIbo
76Xw0Zndo31Gqmt6gnfloqRvm30yAB47PuktQiBc3rPjzAvYf+ttOMvKAVhSLErT
A+2Fqz98ntpLvdgmR2rx+3nox1HozuG0x9lvQqiVDxUG32IIwBEvAJ77ErybdLzp
BT+lUtJfug4nXMPQDGVcZ33xRP+4AYkmLC83vvJZOWxDfY1HGLqwq6ZmcS0QIgas
3qQvcktMsQoSUiaDOUMsXQLo0cihorhwDV6NjvcKoh05mPZDpxRlH+hx7gHBzY5G
vWouya6l4qvlbTVLVl/QAqgLzV77kRMPrX1YMkiqffNoq7ZQxYP2x0/4A5jsZCYx
ddsCDobauw9XOARM06uNDyl+SJwEudI2xac9qYdoerNmNYgNW7k89Arl9IkZunW8
6OLPS3v9029aWJh+uSKTR4uAJVP1Hf+S4tBA29734yGOFP4NzLjzMAAs6l+pUzaf
Z+87pDAieQmXcu2YCA2t5bSeN5fC0n+LOGZuJzzw8a4mJ1bmUjjboGVbg8lwmyvt
+gkXWifl6tAfO3+Y5z6cKnfqllGgx+85Ro9rA4QqoWDPglHXrq2FNSC2C+tK2S5t
nY47l3fgQD5Qk5F3jD/f8f9SztwkBnRKwHszO+vJu48P3DiVMN5YfvpC8y/W7mo2
9GQ/mscs/pNWu5P+mAtwjJA9U97+KnjBPBYWCLDGpcaYzzwYU8q80Ww5+Uc8yhCS
FtmwVPSl64CdiGTN3HtAJlNXo4or3LwlsON+m7raWdBZTmq0GpANIitIJ5U6WoCM
aWO1Z6OHBhic3IRdXI3FdmCfjOvFB7/7u+PSPN2XCilbW+PXMocfqowF1ZteIzPj
r+0J3JdrMOBZVx2M5nlKtBxmChR/p4FWj1kX0wnCEU7NcfM9itb0XFKKnUMQblio
xdcy7PRxiEK2ZU2pM4/eMJ//8BGRuqZIV+NkP6HeuguFCQde+8ZO/fNH7ig+eFK5
T/ED9WOU/ZaTiFklpz2HK+cv+YYTxgiQASva05aUoqaa9nmJ35sR/8apf2LN/gwn
P5P6wn5JpYX0akzBNQZdc7pOI+4oP5XsME336rVfImXWDIDOFnjocO+RRC9fnLWs
FDKv3gxO37VkqMJO6pztkHAEiVq/TK8i7/BoqKcNarGZUwS78bIoE9FbScruLRHN
B6yW5sfh4RvucB3v6HVHXjGfDoDCfZ76wSWuYrnst2CxrCqVS2eAmoTFgQZajvej
3AGd2kSWVW6SOHSQDUwQ7sq6PGMK/XbGDIUx0k1Td2BwuUeFZ6dpvydxjVb1+FRL
jGTZuJhdAyYgZD70WlRsa/eYLbrW04pF5lIrjSh0S7Sg0/yAWP4056WhLBxI2805
PJ7MXgBB0suWHaVuPd5/LPS97m7BnOFdxU2ll6047hPLrXdOVMePFZhUG2A1hfkh
EWXTK3xu91mX2dPn1ZWkKZJy8J/pSWm+jF5AfBLdJDwgt4v2vtVRbCfulmQ0gy9l
UBSLCBBxqxNzwittUtXPeha2sn4Q5xXOIUbyok0BMbFmiYGU1VwKevdjtS1TnEff
3NqY0Y1MdBVn5lXkob6HksePs/YO+S2LedDYnI7CARXP2nfaxi1ChoYEFumzuj9N
ZH742hIJwZ3uTG0ZNi7dJ9Qsl8f4K7Lai1V96aSWVIvxwQAN8GoTZbp0ZVVhoOVI
P55AMj1J5UGPaOmR7bN9HzxIVnOKKtnH9ooLQjJfYBYJhjTQxarbZ5NJ+yJq9qmJ
yHiA/K1EIQ2Q4b/V+TsJZhnZydf6IwRu2Ab6u+AHso6SW4tDpx+SebhmNDPZIX+n
UJOWIQQKqGdnUW31Lbo/76qusdr79gMTDFPAvgU7GOJCFXMTaukrX/FdYaZduEi6
e7d5snKyKCI7ttqM4IxQlK+FZdpIWkrvPUjehMR7vO0wkbktLil9/m6CGHGxSk44
iEG/3Ur33ZcAlqq05xZVU3SDxTULnglu6bFYA63f155kdgdeYwSSvbxOawFSpx2J
aicGqdpoZ2N8pQEfkzjAaJtKFgYGx1yno97S53+OF+92NUGi4d/ASSy9Wt3WrPKr
RQXJAgNkstmc/B1C2X544JwIdWhR8b/2owHEAhxOKP0wgMcwJv6WAjCqklUZI02o
bs8jT271VGu2xF9cCk6ybmXpqcWSc6HkFhafcgFyGfMrZq9ag0vhoP9ynGNlxMfN
Yd2K6QpR59lg6Sa7qGRw0PMm4ngInTdWoWqQFAZjTMFqnyxeSrkT1FyVjO7bJX6B
tRGroVipF7TPGydWDA758uDyHffEdMuQhKSlumISbKKvBJjJvli1K+7/3F9zOA2t
rWlLV3YRw0Rskyp0v49QV5fdajjRQjB+7n9JTDn8dp7vVtnFyb2J/zMH7YZ6vZu2
fpWLHFXsUSwpRYLvJgjZNUMHNuVjk3TB+Il4nSRLcYseInCEMUqOz0GWw3M1+vk1
PPfBYXmi3MgXeUHfzKTwO+v0TUIX1HFpiu3tW/LUp02lBw/9/zgqdaikRoa+zDnU
4xS+8ROKJ7/Kw+LYao9iqWXgDq1rVOcl3NINXCkm9yPFMsGL1EMPjIp43eJyVno6
FiKwk1XQmg9JQnUByZkI16sup22GrI5fr1AsA08h5+BSl5lnfzhxtBHVIkD09WKb
tNOBSrH6AuVD9lmwljrEfc+QhOc/XFSqGV8nJEmmiypkA8h49BtRqIt/cBP7bayF
5ZDonq7enlPyqdaNWGTsK2fU5KfsVNu7N6H7D/5bBwK5j6aUjU4CoSrvP7e/5OTN
sy39x9qpgE6EUc9NmBLGYVtrg5W0NUi/IqJWNb7GsQ2LyEgBPlBF9Sl9beT1ywga
QPfvlZcypaAf9ijPt2PXnNPuiVER/iUBV3l81ucP5Uau0k/Xq9YsdcCtaz/dbJCQ
OfyEPZ7/ZMCFUPSNGRZ/v8HSM3Ye8Ej+rQ8cDwgScnVNcq/zG5ip75ZDWfF6oyk1
4QfqQovhcVyFALVK0R4NstPtQC/J8boZoRZFJWyubpeo/FNY5pDFkzVmr2MwQeY9
hQqCVNPKxTs4ValFywZquJev1k9165Ci1J7U/GROusK43nSfMdTP1JajHv1R66a+
e3TopQD8hy5Yaxedx31K1PgY0WhgCCXYfNhtvO7uGHW+wUZZC/WILpMENfGWvhUW
HS4M3Fr+iKhq2WNDqfj6oIoksNvDDUVnyBrrxA7xz52wTsdFhSLPo2Aw7zDaDqgY
R2M0lifQ2nFRlZXL9uAgjGzd/loo1go2ItI7Hc8qYA2jLHx/CSxfNqciR16M8ndT
Zmp8xX8uOcq5odABxTrzggbKVmYlQtuJDhM+ISQoQWoKU6OzEkiD/O6/oxFDACgL
JsrCNVypRWcP8/+41ssmrzCNCOsMiJk7GN3lyRJAHTE0tenNmi+lIrOYW76KFWF4
F25nkrvCvkN2idMqfTnIFIcUMoPHH8KX+WjrEJFBWwA3vTjotY4H0ZvPIm7DwLmA
bFREAHLTpBdSC+3pJWmZ2JzwWAUb6mPXniWJ/Kus70yrSsJ+dG17+Tz9TKFtzV/+
5U40kNJ4xkyBn2Er5JKpoA6nsdwN32qrBWCArkCI/DYrTUz+yTVOfc6kxVt0Zxwr
KlSRsKHynAL4b4YZY2SjsgDN/5BOSiKBOPTx0hbB8UcVyQGUHIQMadpxHg5xcnxh
Kb8xRBlj88vql8SmUIP0hfyY3Yt8RRLvZW8SD9NsPoUzPPn73JzYvesSGKr7Y0+q
lfYc6nJeuNV3fZknYemF2Y6Lp5ahXDQNyxUY3M1v5y744cpokVlpwuGXjXtAY/44
zjgVhGYfUIfLQVlSD8u5r3N2Jw3dukPhBZtpLwK1hvS53uVe5fqWwaLNI6H5hGFU
r1WrNwFGy0ab1p2+sFtuSvK8nYTdkfIPbZmSNkN6isEYrnMcNc0sVnVMmdRqu2lt
uhPfgyjFk/uJ3+IFWe9EQ5esZBlO9mStnNaa59oqjS2cMq34kU5pckUBzbWaf57L
NhCZ/4MJQ+pXZxeX521XTF3hayotD5jZ3KVLlE+E/kzf9vQ35JuviLGsvDC1U41m
KApA5Ph5/SypLgL3xVgvLIhV9rHMzbuEnQoryqOa+Hrm91a0lRLMp/DqH9sPyq6m
bMV3fqoDyWyLQzBmHvQHaS3NDcHYoGY2SjMaIetxEzxqX6gfwG1mlKXUZKMykiRN
DuS4z86jM6m6Q32z23bU1ywyJBVNBQ0Er6FioKcGIezYd/J/xpXVumObhSUAVHot
lwKsWnHJvOhBsArZN19u0R2L8/Fe0iTBzeXcvCpBUx0JcDJDJ4+0IV+3M3XRtriF
3xcRvXqQfjC6dB9VL4N0zf7O/xWgrqB2YEtbHF3WGjnPPxWTkuUsW2/wvO7e7W8H
u6UyhDGA564zj10H3HXasmyV50mHLd+w18nxF4z5kT/aSjvBoJ1p+xtgsJyVVt4J
7iyVvftux8pmtdMK3Tjl8KUp/Rgag0ubhIZgXzGiw1XhpDsLkIkk5gV5tlyqlohx
l9EWbWRY0a5QuI0WpLQNruzyONX11HGDuDze42Cd7ir21s1S2fFffCCWGvJNx7rI
GuJxcDvLj3P3WlIwtlZFnNDmvqL/EOCMIocgnwl7/U63VgNIck/KlHDPxeRmZ3fe
55QOyHqEuAqBddN9qd9lPbLALlRSxE8uWRsqlJmg9AHxD7fov4BS7qyByDYpzQpf
BmTci8Ih7G2StxWINMbNRW+P2mF7vM5Jw/vKHaBSkcki6AMhp2Kalafxlw4GFj/a
wokHBdtAKFPwU3EnZbh0h98JpX0ezU8vyiAQJgG+uwjIVB6ZTpofxrWZQnwSX+U9
m0ChOHybQUfbJmQwNXNRNHz09RQUxQ43D9O7Nd+MRay+PDsDNslsHlu3BdVyW8hg
1drLT/+y1nZ7YW11ogWUDhAKnryvS7Xv6KsppB2VoTIyVZ+cFYAhG91b4T7uq4c1
zmmqSuEEvtl9hIYXsDmKXoF6IehVEglFxUoTJlWKWEi+18EfJ7DMnOCzHuY6t8do
zmdNaasd6lxiQOzDXcF+J45SY1WVkl+M9qoAUg1RbomZl1BtzAa3DTf/iDGHPHi0
gR4NykbkN70PVlWrKAV9nno9ma/RADw1wNu2Wn5oiaxAOjgNQRqOaC20T34Uhb9Z
/3eOqEe6bE3QXAULdBxwIZfJhxz79Wb8mP485WGj37pWzfCxfAhWgCoyhhTNRNL2
LdO+Oou3ITEmSYJ6dzPFAxaliKo+yE6Tq9Qk7Bp1kf8fUZc9CXrLrzQEbab1pocz
lLiLPGvgeSNBixWGVIT/7Rn43Z9KEdNHp9DVWGoIQVZqK4tdxQ/GlhIfvjpOci/N
kYQQtqF0RiH8Eyaa8iQ8Yidx/T20UtHudi3YUkWmSXXpBwaLtZ2nOSD+48+1P9H6
LGQPLhjWGPttTL1VZyRhwc4DPawWoYEpuqssjNWcc8sDJCoIo5zGxPqrqHKHFAby
6k9FDeXEycN9WRiOt8RbiYHPFQmahAkuJsZ5lLQPsNN4ozuaHq9GibEwm+4yuA0W
zQu8HuTPJH+MB3juLJTI7nUK3iBwcjV9ntAQN2o+hB7M0rmzd6lQteRfWMsK8fiR
DMvChMLxjynjHSCjQ1KB3LBcUJQ4rmN2XQfpvahwxiirKzHM6DWrhrSo6IznSafF
SB3LguOYwoZdPlhwpttqcQSXzL7Z9jKSrru1WDG1tQCT/53m+ko4gy5zVInP3lbx
RUUtS+TSaN50nreT4r3o+wlhGd5NHPvA2xgLVNlxSWXZim5OTRVycT5BdrzxkWVS
M6rWkgQ/V853j1Z5GTrVZkSALevNofw6T0gq9POS1+yfTdXF5VyZ4+pGhvy5yA1D
g/CeuWDPItRg7e6hiZJPnmvhc9/7+49ctFXvsuczVHWlfk5kyFi4s7QoUU4Kv0kl
y6xpU5HOL1h77l37TvCpHHufjmRGCd/lj/zKibK1BB93SKqMjefihloVAfdLr1mV
8Yk21ykuUV7jSAD69rAlxz6U1XTeT/KjIV6JdaJwhrRuDykofZNfPP+fo3D51Le5
kj4wEg3Myh9Fz0dM6ifTd2z7yL/H3vmfwbRUFMOJQbPuyYEUAm8T8nu56TLPHaml
rsVNsZQSg3d9Pby2vmHI5hqIeieTxjuERgmsLNkj+4WoDAGkVUb16kN86TFRjcey
rO9dW3OZhmd/lgS7fwTrOPm5LrRbsSrkBpwwahJu+k32bp5qJ7A9Ygg2SiKy5myb
3dhIBxjkB+EepnkbdsBr4E1FCItc6RWSLjdWzoc0Zmt1whYqSOYlbYAg4xor2rE9
Ka2CyCECIXa/qPplU40KZODigzEsqmJAfrj9olMvFm9vfElqlpkgFysYfO6YNl56
H6kW/RBH1H/d8rJJCCqZ/9/yzzLIZsUS7MJAftPM8sFOya1tdiD45z7UfQxrXGcR
Xpca2j3qPIckcFDFmunLhoLVAsumGLaYUEMRYVGn9TneELBK1dUCn59G7zvOzZdR
Jbd7Zrvs3TLodwECoYpVNa6+8cE/UsuQqq1ZTStTV1+v/ihPXhumbgjP3M/WnVRO
nTnfRC7G9CjKorrij6cdMcbB/GkgkmKnX7PInrh2I2NYcY/NJ1Gkg0+W49loz6zA
TCkpNfPjWtwfx/SCxlFvAp2Trwhs1XkraFn+k8zk4cNr/Dyl4hDifv0eGWD5e4SG
s8C96dtX8HhGqHPzAG+JVBmPGStM2apIibM5G4s6fStpRCPFoBrfuMYV08aGKEZ1
OJf+sulIDCHEPwgN4d1+7vOLRrthglC/0USJsAexvhXWzEUFPFGHREvOUrjwpCum
oCoICRboUKRiMrL8uFXA6JoSyRFyCud0K/J7wX08s6X79M1dXOi+bX6vG5WT2G+H
wHImMBCSBxaNQW2JEFZM8p3v1Mm6uXF2rqJEh7m7q52QhyE8wb8EJBz2G3hj9OMV
O+nn+tM8W9O+pMtboIaxUHjBcjbKgatYrwlhiIloYhybRYeEhLcilymAIoTEtKFk
XXUWvQ2zNq61/OKqJTAIgLk2trj4EhdtU2PdGtZFdU1FkOopNwjsK34dsXdZj/D0
h2Uwzo0ntDc8VEPlYy3PBRxoETLxgjuNCH8EcwOx8AU25Fe4+YkH2ARIky32iGhB
bnCZ/J8ps31Fkv6zBvhLpl4q1tjg9kRXo7uK8l31hZS7p0eJZWKhEDTAZx4TBU/I
V2hRxg3ivrG+wLsK3zjZ3LpplXAWXDJYePXvwqF3pNMJR4mdfdM/TPIDGkNvXd3B
TMQI6tjDff+e1tDY/5TeGiFgpbN9NBAY6lkCvudKXVbXs0ImRLxGe+E/jikNaa7v
BVNYReIarPjIJdCcGo/zaAL26VQOtEE0hJieDnzYs7ocGLSdKASaAKlnkuFjfExe
L8yWCgt1IgBjhoO0FDhyw49i1YFMJyBXCsCKBqT8Xug4Rr/8De/3y+m4h4OKrVrt
bZfr4naPp1z1H/yp0npWoggA/4l86/wI/FwZqh7+UERN06m7GNDxsssAJZA+m/Gb
Wkhe4wmvw/WPsC+LQ6HqrFPgDKjdNvi2OJ989to+PZ8JpLdjXeXjknGBoyEZJNLU
//LWi4EoKPlSq/Gt8xEhlMrpp+bRJ+lc0jqp/39fF8Fq5FYcdsfgE0y4X7H7XQjX
+N8PlYNP3FkA5XDHdCpXSBqa9igkIGnxq7DW0eMsyIOdrEFOIxofnFSLDYFxHb7A
J6TNgQDFVqlmkKby9gizFd0rjJGwVbqWzE8qf/n0Qs96Qy39mlxzVQQWNEKQTWZk
tQu+5iBAb8JjE9Ri1q6Odip1VWUhv8iT7aIPEKpNsa76I1yIGoCmBIbqzToTkHmo
e6z4aPJHpRb00Y0EDdOr+Sfxdd1iNgvGIG00WtRvbe8j41qV+oCB8tJtz5YHaebB
0Hr1qxVaqyQsJIdfbN4XFV1+Ljy9He7XBcCIJD7O9fTEaadKp9Oh5OYUIk1+0qp7
Y319CywKBfR091Fqj1BxBr9jVQtiXmTAUvx3ul7WEu6f9LHlJOIHyVqSR14HYjh3
yw6PZs6yFKkFoH8ZMSRHzbT46vX8yCpsbTJL0GGTts9c6v7+fN6nv29hXYorAy6+
SkAkjO3bcIP7LA6FrL0Kugv6mr/ODPVaRwbZHb0dq85eC6HTq6XCPSWZCbT+gA9R
q45lETdEYfBDZ7LrClVMYCsHZyGLSXddtv/EwcpBBp3ctZWNaKJ0vcNiAlhlN7Ir
y3syMvSFLGTe9vvGxAkBuaghTD3n9b2Iq/okAfaafNzvP4sLYzRoPhbMHk3vd7GH
y6zhTMnlabEjNUDzDJegqktad87lSlgJ88bXan7d1dI5+YFyZASZQKi32RNPFC4Y
3iq4FlCLnCb0Byzu+yCI4kzLhAUGI5u/HD+oqhoNGDpvXoDe9Hr2DyU7sg6M1qOr
EUmOhRhwuHedxL9kPouaxCitRnvKOBGA9sWb4tHbkv+UKDvzUCsn9APMDPey3ia/
Zj5epTKTK/Dj9FOQ0hX7B3RplLRqxV01XKGdEl5JBpgSFl2DePEAz7JOxxmLl4IO
6UfQ+/XtyVsRiHpmusfGbqeeLE31PzR9sWBphxi4XGyzwgvWrfPRwrGVZoHfha5h
vzhaBYEWjnmXazRX6rqaJGDDtDAnrlB8YVATggT3O8SNI07pSAZteksRU59ZE9Xm
bm7LYL+SEtBGeNZBConaHN3F6TYMMsaers59upHHUT0hhLuvaLs7rGQrfptgrj37
VM1BhP+sp8hBUQ/8kCBUysaoS0Hv+jYlE0++3tUyeUUMJ805CNs5MRc0N2vgCSFX
+dh65WZcznzM4uNe0zNEqh6ex4eeqyUOrkCQCfBc9cs6nd+vZbu8qZOYnUkvgKnd
hyS0RJa3/OTelN2IT28ydVX1m3VPyq+gWvu0ENnaPB5pTmmNesJwiVAayk7SyQ1M
o7kMXOpDjCIsPBWLdOf+kpxUMbTFAeht/xIS+XL9kFs5s9DepPKrZ9kye+sd2mLV
+8k+4vB8GuV17G+RAareET4POfbZ1UojimTsIWYD0LvzQikPs7+te0HGRoWlrLT+
L/rcsNzpg216q4Bfz1KC8E5DAYNTm8J4WPerhfARmywhHl4Nqi7zea0UwfYXQY8w
vZmasrIq7ILPJ0O5pa0jd9VZ6AiU079TNKLBpfYv7SuiEFmEf0X2b71tTZXC2mjY
35uf3IPR+W3PPtmTELmnhob4zUgDR5bRFifE+kFznMwUeo01POehwa/iXdJXrcI4
cwIUHQ+imWCu5SbuHageG6JHkoJnCzO4XNLC/UeooKg3AzmFf+mmcYId7XwwpGNG
kPL6p7jKN/dIKL4QTR34HYfQG7TbpUPQDJobOcE3WkVpjEO4pWzs3UHwDLRVCxQc
/DbMDZpDF21PlTq+09nc8qnlODUj9SDm8yG+/Q88Hp16k7cXXgo+MRMSbdxzezyE
g3obR0+Bkd4EsxZ2K/fkGc3bZmRkIyUcPj+WwnKlJHVpyWxfcS/YQDZHHO70bmAd
4YTJKtLVxpDnb4YmaxZBfAylshpyqPQRYWhcjiBAJN9dZqWFduc02IkN1PBAEi8S
AKOsJCXsdDdqRh0kzl5TLuM60KBteddSD3JbsLkSiFtbVmCPsYpYgTqy8srbI5tm
JrPZXlC55fS/42UP5sOmUU/schfDKgiMqvFHb7RucolbWdKkjsmbrbcgplja1w/Y
mFdzzWxs0+PErFRYdmk0sXHhJLH3tt2+yJQnBhduYLPk7V0IQXb69pQ1yP1Wj561
Jiqy7WKnJvwE75RUXkrKRvFbDWvwvLajqD/fFd1P05C4CplBD2Al9bkJTF8yy0ew
ixhS8z1cfUB/+uwMl7szQumpRvyZQlS29wUVf1XTIbD1DQ7Bb6uzHAcEn8lR6P4s
5PZWdDEfdfNW+7BuELk1jPm0OcjTsyXwsoV9CfAw7fZI5eEeE8OD57zE6gIazNuF
Kr90YWo6tgTuJj9VdKPAl+22WGoLXZhxvblIYzIUV4wi21IgzIZpqB+o9O2ZnDhl
2QNsltyuE0Ki55kUu6ll5XOXQKtfKdq41k1Go9PUxDYVCeJHiilCmZ54/1AVidkd
Oo2IXoiGQqkzS5T0AV02174gX4hqte2OYDOLOQxGR7MGsgI98k9x1TVLaPQZgaWV
D/DXXPn5GKAs+rLyd2jLLfHRreJqyxNHM5ecBHjbTn/dbf3JRAoPXLvYm7jb3z9e
0eesaBq0jSdQkCCWBkEd3jQvgVD0C6OWRIT7+rXCZEYT6/sjE+iyueslPwrsk3Gq
9Ipu6rPrPTb61Zm/ijYxagxTa2/J895p0lUcA/+hnQOII3rdSWHRYb4Qnt+e6tpL
kq2yFzgKFveqMF5A1aXzqEm0NSui8kYNplNI7g4xkk+hlRIAdew+usUwvn+M4Qq5
HsUyBlLg6QVFlSwOsOExgXSveT5km8t1VGp1cMv42HwVFNBMvglgA9WRS3pV+fSH
zLMFQqI5MtU9Sr3IMV5b9/KdH8PKLAv0qy3HDykWF9qpIhsVwrfL+bHoABSk1lMt
wZOeW4iaWBXgQ4YjwQJZeSzwhqH39VQxzCLIroqq5jmsSwR6eazsAh+FxPhgV2fq
D9Vb1n2z5DAhaKJoL9+7Y4y87/oqDxgIZSVObtCEE6S2QzjDsY/pl0chNjTDEdCa
Fk2gjVNXlKbDU/G++1a7HUU7aPibBKw/Gdbgr68T8NoXSRC3Luxlm5cTJWyY4QMV
rpPy3OwU8MQMFrZGBNv+LkkLFMgbI9sLaaox0NdZvt5fOvXK7YcrQo1ZYSLt13/l
2s/JRf25IIFUqJGLVcVCthwWVtmhBuhod6fY794CnP3576XvfWDV7qw8RFQqni0t
cmFF8SO0f9x5SpagWP81MkxqJMEIELrWu/AYKgrKkqp94Lr/hNeQD/Wvj36a5fsL
yX4gplmfndDiGjqkBK7wFvZfDdNHes2PvbrGbikrTYz69IE3wzes9NaF/nyGe8Mn
ODDfPsZj6PZTqf54PaN4e/buYzJKXrAu96RiET+Aa0nMRFd4yApXMw4poD8HLcpx
mZ2iTfmlm8P48NAEOW4oKmwFjzS9iwlB/NEf5QODcKuMVVdc18GJSr5e0xLGhxbj
SJ+lIS1ha0Ny90dTtK1yK/CyFkK4x3ZwMsicQIx3tN/h4FbKZZZKKvom5RLmS0KH
eyHJ8XrcIP/Dbisvlj2e+a0fCFSUg/9TK4b1VrvUkNmlBmbtvijCKD9UQOc0V1Vn
bdq7krr9OoVzsce2cKppvEmYjMoNvj9Ta262r+XaPfS/fy2C6t99OTRE6b2Oxfel
OxmPGpPg5qTI75LZBa9CXLmuaz4Yx5ezCW5OOtesmMnYrrCcA/a3+MJ1s94SakIj
QSdV0JS4CTwGc9xC8T7vr6ojKyxSRx5/pOK6857mZAlSnRvvVawRkhAxYSk8nve3
dIr80T58wUkWgUSOWpuDOt79nuviylKJ960nYVU9TsZ+RQneD648aTx2DIcHCXAA
5lrysIWXWQ1klnXvT59jTgIbJfFcrmU9c75kzJtXKcD/OLluCqexSLuBh3rfUWYq
9mhEjaTPL4IE/xKTmgtzEtmS/+4SR2eYTf/aZ0GUJb6pAX4Jgn43ebPxZazao9ON
b3EyrrFSAsZ0mm/zTkjRyh+sBsZBiLEyodUIKkx0/nsNj+XyseN/qsiPQb9edMgz
H8LkJpoTG/WVQTgdo+zpUYfgSE/hTHrKQppXn6qKR+F35YeIYKkgXCKWTi0jm++T
uKHbXwRpk/4crQpK4PkwyyDyd9u2qvVk2IO/Yy+snCZFnREbN5K88cpfQ/fNAiWl
4BBPwVaQJlITtTL21XmqJ5s4G86db6UWNm5AMgtwKi8Y/jsgwoOstDGzUmL3tGyq
MQYTihIdl0ytf17kBWxHXogCLEgLAl1WMD13oqom5tBZMLHs2r0pN6E+I2xvVF1F
1LnctnjES4IF4W5WNVrW9FwlW7WDpSDMhtPGqv3qPftOfmyBwobWMInTNReyLzO8
0aNPdtKdJc97IHuEXFtwSiYKnDbN+hXJhJN6UewwoZtTIeEw3H+41Iq3kzlVcIET
T+MN+Qr3zX54TOOcvLM2te02vo0Xfzwwkb5XgCAZ1drrB+ljqvcCZCBjgsAm8a4K
3D0VUiG/ZW6IBaQAX3GXDSI/jxdCF+Nh5GxqhICpxbu2WUzAsrM0vqkWOTJqnRaX
UdpYpP/U9R6QhCA7vZX64/y7HuyBXEd0cJHZAgnkawov9UupS7U9IXFmnE32vE/P
pnsFAQctPwYCU2fkyupbtNffF2Ykn/znAC9jijRRiujemWLhMfAEI7+NLb7e8rV1
GoUN9SpvqXsatP+G+zhD5pGg4YOYzukzZZoLhjJOy3yksOcZfoGfnX/cCqtRnlQw
7RcRl4dYtxEgXsbXscgtxz0FjUvLJajDz3WHLeGEAtYWLWX/8gMlMv/r8zFlo8dq
0cHzxVANNLPsrVz9W9v8mIzUaSl3b3RiiPjZYeV75EFqRvATRdMa2TLcUnFX32+u
CDRHsHy0PRTBzJ5sh+2qVnGb1fiB1U27+M8arA9hGPUUtXt6XyLH8Mls0D3vRpc+
+WmB0Iupd1c5fyLKTu4lG2Rkv95WSSKu8No+QAyerfCRY/dXKPfsPmBvmCSP2KsE
OCkiBJuRpzpm8Blk/5m+kAx+/kao7ql9IZxiyTZp292DTL/sXNwCgtJH9Da/3NYD
Q+/H5AG7ADrjRqL5p/94LBI7A2Ys+XU90hw0jazjRhRXY3aqOCl7dlvl2REQqjL9
Pfy4AymeanClsKVLS3S8H2Ch1L2wYB+gX+x0cwxMeVyYWgAXgaSSpj7u7sX9OJar
EXOmhh9LaCZPGBcToiMMUu/XWnHS9T8rDg3KFEo+v2nLvGD3jzzhaAMPbYulMySH
BioXToPO4KML1JUXzozraOP117OUKmfwNSixysKvLe2tbeuzDa8ICwFaTAXoD4Ch
o0Esw10eYWe4tn33AwhsgO7H2cwttGSFRIjhv54e1A4T+rPkOFWziuXjOXBOkHfU
kpEgp8RwgrKu/TfdnxEN4QHBiw/n4EBfd9yMstF/3TxGIk8w+VPFeFiuhkmX/bIl
QX2ziY4+ZJlCdZH4d5Qv8wb8B/ZF9Rj1i0lClNrTQnev51xR4QoBIz4j32L/f9H1
uTd2MQ58f4G2XLYZiSqK2XgHl2kxXD6anEblrWcM1r5rUKh993v8HpBCWFl3yH9i
ExYQujCk/kcqam4WA20l+yPQ2TEQJbc+a9dto80HqrBuhwZoZ7b8HQiDizwOat8c
cmo+hVbxznuv+ViEMUoKm341Ge/PQoAAloIUUFTPrbvxVTIkKdC/H42odH7Mud4F
DYZ3RC+nyqS4QuMJ7XhrYVrtWQgwf+tfkymAsfC8ffuji4o5ebRYEt0xiYMKKrCR
MrTIC6lCS/akJ6LLNuGBDvnJEtbqrWS5CuAe0e9yNEVEtvJ1jBw5okoTh/KSCWvh
h6mtP44NqKQKjuLHXAgXhh6zSC7/nMWQNYwxNY9nzFScbPDBO4V97dLqlASeC4j9
nPTjcSd6BfZr2DvyYVpRd4P505oqfB6tCyTr7j5TRFtNBVbf/ki67mQm9LtsBF8E
7S+UgfxqliDSrMbLNJ3Hq6w45Jgs9XT0uWDAUTbfin4AL62vUkBS79s4C4siTGmr
Tirg1+dJ1aM+ypHi2hqMJYezF1mwtrt7HgX5OYiWMjU4QYH5SeqZ/4OCyenj6GxD
8tT8uHN2SuQlJ8O0biF1ulKaFeMAId/ujZ4vziKgPUqtxtpHe/4p3HlJiVBWUEJR
Dc+HFgLWCMeGNEcyyLJVect8qkdOFWJVrhRqFxIcwjVFCwKWxOX8BBIcBR3p+7ZK
QYUkURV9/72gVA4I453f4cXJVmfhIOEYHFCYTFRDaPX0KeRXAdJPvQIB64b+V164
3QhdExdG0VooWsrNhvKXxCpC97wAdzmO0KJQfakXzgH8OgaaK2DNOKMD+zmJ2unn
m7KkJw5aa2fh47J/5sxAMiLDMFxCWF8kIkvpegC4yuhnUDbmT1SgBtFMihRb75CJ
jTcW2IZ1DlTxCdBe0OGa2gFhYSsOWQod2FH77/Toi+SCh9TiaycaGUWKgXjDnkHv
I4HWbuTTOnKGZbVuxnTN0IhFY8KxEjZiSkc59gB9M6vRB59LUeW6beIqnt+kn/AI
cD5vKBGWR2VFWtVHNobe1Z6CvFuoCtisfkuUl46cjeFA/NKwl1Kg25Q0w2ZrKcdP
/u5sz4fdfUcz+fqhSENybk3PrGpoOThbvtzcjkW/pGDAOqS9+kpMNLoNXmwADTfe
lHGY7mYDVqlU+O8H4LaWluW+XjA4/lukIlbqiY4XwzfRrrztITGsJMQBaUBvwgJW
sniFE/fblsTrbsjrUKe31tGgr95qOT/UkYau2kzsowm9sFZFH2LAZnxCEDSWQVQ6
Z9yRkIIa3fgZOeF9cvAZKuUvdx5CbRjXHtg3u56X0IAyeoQENxLD7WIfgXtkp9o9
mwz8TM/2CO4epCqAEXNxbpMQ/3uzBx++x7chnswU6qUC26yy3JMaLkAhf1vIXF2z
tpOVo291ZcZOvgufKiHMkN1288ungJBSUFpYja8oIUNc/jR+jYV0J5cA/LTZyeBv
a5sZcfuXUMKPyXtsHM0lYkKYBoynNikcmS5lJIzQZnu1lBpDgA7TGa2cIiyF8rR6
J3Nzssia7+qSwJ5NjfJ8kc731Smue2ycyrL2mkAkrb5nyOVyQnqjla+zqQrGxpfV
J3dnMdO4gMm8KKQOudsad9N9OGlQoR7ZxJ79/h7uvSSv8J+cSxODgyEgj5JwSUWV
XIQyJdGitLYbYRPXdtRaaQdoYwbMrsjB/yOjKvEky07uQd/S6D0n0YSzRVVFke74
wpLvHs4CWmP+HBya0U3/CWz8zocvvHodqFbe2vn6vGK/ENK9XVbOh4k3tubz5y/a
KKoNe3oyyjcIaVKxroP99MBfWFl8m/w3uB629J/2XdBS2oxmHiNyw2fip5fgYpb4
q0i/+VrbrgcHfwNa31Z+J8GlFEpptjSTnsOJESbLUNb49dtyb+Ol8JHL/sM1io6C
+o7t4unWoXxoVBH3JdpPg41awhX9wiPhgQlgbqSdHRwB5wT27ZtwIWpZxGBBXY8v
cAfSm1BkjKOEq4bISXqCVDir5QdySfYBncFuZqq8COivvzgzje9+UGkmNywn90+n
T8c0kcHhUvkC3ylecrOW4db6cufHs3ihlzpS7r3dSjB6KWvApMhB4zOa+TK3GW2J
rhhsac1ExtgIl3XFjp3ygbGSrHyFySYmF2BskS2PVpLPpghT0I0o+VRXRhkJTCqo
IacF7gYXVTizTroQ+86PJQ+ZkZztrXrCWFnwuI5+PV7hKwS8pkW29VCLpuJaMYpN
e5lEVEssk8jNJoj8UmeyWa+HUlPTYL53dx2SiVah3MCcrInHJ3yDQ8f3M6nkuurO
2gvOKSBwrIPqYOyyf6EUU3zCYvVYUBI7ukzNpnqLUOg3w2bi+k0TMdD8HaxeTp8I
M/E1mrnuG2aOM6p7iJoZU0O7uSd4KxKI4RrAMQ+EmkrXESU31XxbRdILRYGZBh/N
qDrGCi8vK6+guceZOqWB5CTDso4VgtnNfuIqVfmjSSeEiuoSipScQyKe64l9XBt+
T47lSNBEvt7KXYz1kAtew807FcnWmfAHBubDIBuoTeXBNTuctiTaYmx5kpaFZmk4
M2DQ182oEc6tMrw+GckjXSo+KN11vvnIP/pDXQ7KHYcoK7CrakilsPPii6o4hCF5
jTTESrokWuixj2aSrGr8Zos04s5q5Yh//oDda2Q80boGkRBLN5da2Qn//af9d36e
x8RNiTMnsQ8VKrzb7nrdQgTIsm7IXMHPkDtXHbjg7Ew7TSt6NB3gjYi8v+U3E+EG
dPlVhHcj49nnuslcfGpRzJfn/adrgkLXrgdoVHlpYgOFaQUAbCPv0ldlCcg/uK/B
NAi3b2VrwCamfwiZ6gRGMpHp9o4Px3zT7qRcTsBMMvI6w5QVVRXKEZtKoqmiJEv2
wfXPnGjhj47GSuPTX/LDlyUPoWccSE3Nh2AuMfJR+Bs+5DtTzH4acweMPuEK2MhD
Kh+3hmvcaFn1+1Tgi327akWDhHRkvN9SFguhpKWRc3JO1ukKT/SI9yh7MtyuNtL+
idwIvkHea8QkaRQI83PIrWiIWA8xmUrEOkhaHFc2bs467zrdUsysEpVR5eJOxgZx
8x7/35ETdY+R9iU+xX8qmn0XiXdxco7X/W6gQWPK7bZvlWjkmw3Ja5HAPoWr6wXo
j0etG/Y4Cz+9FgHq6OMIZ7KaQhCRbPG00W+8Tyt38GBluhDDI1/uTxPzmQoY8BsK
ga/OjqQHO4eYNNdHllkz9Rt+omdO37Izzj6pitkpmdRLbhLj+Ur9hH0r1WX7q1o0
Ht1O+lHal8wpfazV5dj75POCgPH3SuX6cKMdG/PJLz6k+CbV/vbWtaYmmuUupFWc
5BLjf1rmIiLQ/Urtm3OGznRQvzS1uwjXoioz5VbMzwYLJzmwU7Bh/SW4waNm+TQR
+iDhct5NsSpwJtaYZ2zJiXjNIgWYX+nQuYOLsCWKEahYJwEVESCkwJz9ZIzuG4SQ
epmLgVXJGkFERogeur/qWTvValHruDiPEIBotH9pmH7Q9Igm7jEMSnZX5viOe9mz
9OOmX8UB2QQfpvbnZ4l7o1K9/5Mc3zcjnGqWVKzcZX66It40ySwM3u7uOn0ECDnP
PE1cTbCfVGHDjoOOXQE5rQ9WrC+/iFB4m8RPE4KUO65tk52obEHONF9uCoJw/Ody
Ga0zcW67B2w56+ujJwyG+ETetKVtS3pJkcdRFy69mgXNy0yKrMJ/i3pwnD1KlH7F
FMqdJrLoyYhnJwacrC7hslgw9PUAD1ysLCoBfKB0xkXfBgIfAvvJ1k1ZRDZG2iz2
Qo8QePdblMVXg3oe4kYFVB54ENPWl83YN8cbmucVa/c5nKaz3BiiRgUhN24SyNMH
OmWAiEJqquivLBoKQRqGdwIAzlO0qN05eJY4TfZfpvoQNL7+RCYyrdlmyhVqglgX
OfC4dUk2NI+DPZcKnWoO7jwZBBJMBrjKlFiodAOlb+QuE4raTiAv7/Wf7f0pbAsC
Uoy2B7FJPw/dD/OLRxQa+5UtWNlXffQmTkeh+817OflyZ3cQ2UFoBEe7Pa+HJdQn
+VgmYepDg9lpd2aaTMAPBFXg5z8q9VtQW0OvHmwuhqGs5kpWRXT/U7Du56lCTbaV
VnoqONSgGSDWLHcapLVN8E8zPc8Lw9ElU+O3yxFH0kaTWuebeo6Vb6tq8c/s1DEx
6NYHIMg0SvFDWmqh+uQ/EybJhr7TAnIV7ypbuXBM2d3tEV9drVQOa8BIJEPBtEME
pk8IxBVfR+qrD8gySAUxyGqWpdP7xP0Ejx+YAG3X9aXH+qj1/hhlgycIBO2izmX1
cMqHXp9kBIkz0LoBXrjW+A8FWLJcVegZdYAOLH6C8wR9IXTVZzO3YfW5o8DzDyyZ
A/KwWi4CRzBvUF19jupUruuMO0uZ9YTxwoALwgmlNeGWnpdkhd1cssEsfeMuLLAo
iLV1/oc9EqV/fEvskAi0KFimPKrFBsctWcj5vsYIf6rmsPms6LWln5kXXBKI0Cas
1yFpfUTM5VHVbSyaTMWgw32/uW6kAF5XWqp9nuezaOn1FM/mmss3alG367nsRb90
QYstY8v3i1IkzOJPpsPTceQNIelw03xerP/abKXy15VBqd37ymAD1MZWVGTDN4wq
khoBKGDXn0nrDThwmQqPOgOsXw3eeA13XWB9NcwHB3EjaYN/Ox3CiTkadDRNffXn
3q0QS07DZ0hrDXBrv7o5Gtxxcx9YyBpI/t+p+ADOLXVGgMfPdDTKpfHuRJgirhlS
aB0SjQ6XzxcmUFVhTa/79oKK/+5xbuc5075bmWB6Hw1szBEPfZapR/a323/R5Cmx
7Qn+wP3gH6Q+P1JpNlk/smjJ4gZGMnlcF6ty9tNTEOkaig7bdZuKaQEHnEOOwmJl
7tSPH+yE4+kfWbduAIQVwHGjEKeWSfU12MRQFn8F7shauYnOwOD3KWNlYiMYazLV
siHyMXtjgVWn99M68YfgD3uKrkbQzANE4Vmp/jdouCdWKfe+YDjypXHopBcYBzQC
fTMEY1BRKPDAxo8yNkq7cbRfE36dSnMyx8qWjzl366DVTZbAvdEn8D8zzqR85YJM
4xHOSySUlTOPEIZnqe8NbczBXfnHNdOho7Kxo6VotuPpuFRtwBG/wo8tcSfYX2i2
DcFUvy/aYcOAWMlPKZUs2KFk32Vv3zHhJTMUyiqVZgcWd6ZjMWcgl4zfpZnn5uTe
jES+N6jZ8EMCScAfpfNTMvmjCOajK0TOpGHTFRNLzRyzs8meQrdqfrEQz8chqWMz
d9O/gWyqbidJfDr0ogakjv48hnC0nyPkdou8wiv1B9WowR/FiNLhuyMA9vs6secV
jUUDFBsp5deNp2dkw7TQxwzDiijOrmjoGJM22L1YDEgAo0Y1MGumeY2j+VsarYAo
+kCPh9qrNW3s0WlVbQ15DSEkg6/yDyA93K8xGQn09ded6DUq/HeMzjJEXEC3miZl
6d/CltJSYMHmrxnyJXsyc7RJEu6ndBT+rW7eegQpHU/LZTDzEYJP79tMvDpf09wL
bX43LBlP3UX8YBu0JuEYjsAlx1LGlP8G7m7ww1qQgJrsdQEQn+MQtRiT5swjYqIv
nwxnhWfJjrnDptmAlVvxgEhBbbsj17Co7MYy7m9v6oUW5UVtKig9KmvrudNoyAoi
4POLcca2ZJhDrJl+RtOgSvtreXJvgWDjWmsKsO2nVgfzu6TwI6Yeyckk111OU0ea
zbQHMpl2ibCRmWErsv25gVPlDNjmasrA3oVdKAV5zh725qaK72hzrDSFcTFTE4Md
7j2UTOweg348GzenLxVXQvLvgquwbdgJ33cpxnGSqc9pdJ7slFob/S3+G5qvBL8Q
H0BiVUipScJHyzcNAVndZDv7sJnWPeBrL3R9ruJbweMn2W1QVWw0zGwyQkjMHJdL
qrrdBQyGX4AxXjdTw99tnDACY0j0axL+K0XFxvxm+mJarUwicbC+qieda3T/hybB
lBhF4IemVUjJI0jULpateAARK94qvOAQ+lRdc/Sr2H/r+EIALSpltNWN9jlwyNUX
8a2K6LeBTcC7t/FVqsArYGSjooypUUTE7k2ldyJ7KWJawqV9LU/VfJYxekDpW69R
luj2Yu2hx53E+F3CS4iAEqTqoQXCvFXlyGdDSgOSWpx28Eld76hyf1MIv2q9wmoN
F7yQ+cUPCdD5PeH56RKfRrqIKX23iVY9wnKkm7I8Ga6/bikXClswx3FPVq+uE6If
KrcDy+4oqhjc9lqgVNn0qe86OpQOOw4vGbqrR0kCwvSMAkTMtqLpOzxu7fdk2aAA
6dTqQrMe7boR3MrF2hvohaOHfOG7/xksUeSVelnXh2uFaCVfQUBHWEvMWZBQeMEV
JONAeuR4Iq/fvtXAttksW8DB91xJynN655GglvzLdGNA93wcZKbQTt3mFdwwcu3v
BP8OdnwMJmFK5oBiI+jZn8TKLgTuP6Os2Oh0KnK/8Bc4QWocudnenGIIP6r4MCyd
LJOqjiDH/WdjzqQJ+G0eub7T5nJUaYZ8hDi53FImvTulwSFePcHfSJE2/r3EO8y7
66ryTLHARkF1pAMyYz22p98cOJWhNDev6GFCKkuWqqgO+297ZVK6c3h0DyK/Na+O
YaQ35LSg/HEdxtEcvAZPUWFFNErx2xL6WQrQyREOQFS+H7YXOFEz+eeBkcAePEMK
ZYykliOuZ0ZJCvwQT0z/Y1W23AxDMJ8mtd9XBzrSt5QbzUA3B5gqEaL978KZryS/
wkZRREvdS/6xCxbtJeYRcBbn0xz4Z655ryKhBfcDXSEb2LeZHg+a/ce10uH6ASU8
FdNw3lokU2RqJ1tdEWDaEPHoSvUxPU2U7zjYTIGH0uKChm0mHAxhE8lnCWmR/lqJ
NfCx+zAADkSbhdg88r5ZHU/0vGY/3AOBjYum/Bk11ENMny7/2452k6T+x02Ec/sF
X6eab8mh3b5ZLlQtaMqLIODAdaIWfVVj6ejx1Gpe8rvWLqvNXI8nW2DniWYaNyPw
QHOP7H36FtDuE5Oj/wQMKI/zzE1+Ya5XaiVHtKpLgDVS3k+Ren/LJlmRpKyqAWPY
2OU8HeJWtyZtXN36meilDGMcSs06foSZJGnCR7TY4TXgEwwdZ3fBO+A5H7onpNWz
n0CtILIjUt1kIBzj30LmIaCUYW3nP4VIO5s8VS0H/icgce6WxnRXtRRMkbCdvgkC
NLO47/D0e59+tlvc5YnwrRKn5Vfp3hl8VqTJ5zd0QqDUu9Fahgr8Q6qqT5c52R2r
HvW9pE0xh+DWb10Gxtlt1zUBkkuHk4JIai74sTrToxq1qClejhKesZ8zVXd4Goig
r6f6W4vos6dIvh7moVCbeCU3wergZDmcVJIJf7oXfTWivdKYBxPzmem0QQxMCMCL
Zqbr+TMJi6NdcuWAYPRO9ktPpivWFd4HlrXjSbv5EtMmafV8bVlm/E0rgATf+vXZ
ok79v785YG2WzxpsASOnlwFwf+S9tKag6KB1fGSgaUyoITJRx67LF6CElAO3vvDW
KkGKUuGe/AEdfqbH1OoAsvKlkh02F2sbGdPQqY6QyDd6/xr2YkriTRTMk0Vpy79n
NZm0DtqNj4dLzyOWH/npZeOIrauNVIAkshBuV0kW77X14CaFVqXbAsA6VgA9VbX5
wJCihdKI0yR1crEoIEenhuobNmiSRBmJqEOfNUw2uoWs+vbOSdNtpvgKWQ3Oq3It
TaJCrtUHC1dMNDdDqhmS9IJLah7NgEobd4ArmIUYzQdKk8sz9F8YqmOJGe9Fjgk5
+JrPJMTBbru3IuswQy0fDzHH2SZIfCRno+3XBFicXVyr3Zjur8LkK1jIfbVBQs0e
bBUt+T438DNj7wY/+15gug69mWuTg3AbdOstNfBf23xixq3hqH8Cpg9n/UXVjk7i
OxLPTH5/b+6nT/v3qgYhalrPQ1l+kc6/c2PM6L8/S4Uf0COr+EyaqFbXbexSDA0k
XHEkEtYPhn7OsJnSqYhE9qS3M06sgaApCFALyQV0BzhMZZENqh8mcpN3Dr5cWDdk
aTakkf9vzPn6cjXeVvE7WyeUA3OojVwZ9yYAdwvqOgM7AbYvvHGDURlOuHG72Vdo
gqndfxbwYqkBq2Q846qapsvTRlTe6UMuCTtucSANxt4UqYZxeWhfg8qz+erfEiuy
EeS4QLl5JyoJyPdaziwDmbjqPkKaWMQRmvw8BOtLOsiyovjxsbb4Ez4sWr+fRti1
CHA7rDR71ZKO30k9AfE4H2tRSYCgwhfHrCepRboRkXfACgJLxAYkZHPf3gAIHbEm
4fVGngHLMXjbPpQtMxyhcQEHZSkb4r55LdcPt7nCl+3A10Ks1MdeWDKqPRJEEziz
PRcUS+DgGOF9Jiwb6O5K0DIG1WpxNj7zCOcYZlph+Q6t+O4T7ca7w38jYWHysD4s
MlP+llH06MdhCAhQ90GUpiTeMI6GdprqzsZyzDyLlGk6emfqeicoNcQtcm+NDpHb
gXKzXdytYTLI7b741sVgyyBAkc8SW2TPPX6VqeCYOjXEGgWBkxesasjpy5xxEcM4
b9KeabNP9wrTVe89ZivcrG8Gj2Y3K0/oixUM6XHyVdEt/ksqsl+4PIFsyMOtaHkR
PYfvdDYL29j8pLR6mm1gGEJ+LPT8r7xw1vpI8ZuP/MWLoGesxxhz5S6NHXrR3rnY
HXesh4NEZRP93mFqrPbJliZIkPzVwtFg25k0EgK6LQZkS6TOvlhzGJzygm0f9Qyn
+2Ags61PfP8aJZbHIqxQrfcPL/WdEyeGZ9wFWZXMYEUIS4f2cP4k8sMCx7ynMoeR
39UksmwELPo3Inf5sm3yQfvTIQXlu2CzSUXeNKF8JNdL89yKkFNUFGmeDLdm400C
q27G/TibHPwuHLAEUQiWTBSIlFMuKF3yiY6jGyFt6D5eB4vbAUf2VKrJFSojTkao
guRpsCna0YdyydSamljnQ1GaWQYzAmJPx6+YW1MhpAvu9di2rWz4vFTo/h6Il8+p
hY96X8FPs8Gd4AcsE1bPTJBEb1v4oDAothPdKpPp4jjT1nLEvxfvNUGgtGt6gO41
LpOoQNIkdYC3uNx3b96UHKi8EIAtQDGItWraEMMxMsvZRpa11xMVRfMJukRr3/mE
mrahrcgf33JsiPoaSyVZd3mEUp47n47rG0TFP7E+VDmGyqA8QKsWXTfk6bbm3qtp
hLsVYiX4NPfXDXT/uPDqT4XdHypbiOqbW5K4idTvpAJRJ6tI8NIMrdLAucEnCNJH
0x+gL2gWAP8/Hu3na8H6emhC+vzf3fP9zWCKSiFqN2YmyHu9t53BXvPkl6EbFwLx
pBhpo37vGPEyrmQRAv6XBnk46BajqQ5n57kyoF2SIWUOykpB892Fqr8jICnVtjxE
RbKgLPGDDmN1qFwpqlXjX7fRy+K6jnE5kdgOBYnrI0hNdCq5905WuN5j5QFp3ta7
PlPjQ90vJ2A37XypwH3nhXKmNlWGGUSfKyGhRvWtF8fa0F5/IbUxPIqOckzHtsO8
7HIOT5wXYtcPM7zpPHmg+Z2QFVZ8KOb9i6AugF7062mOL33diNLVVjJiej00jT0K
KA90nMJw6QvuRIJXRiAP9hHchmrnGsGxsNpJyz6fS8xdmUcFqKHWT+XUW//EJksb
d62IFbObsTQLwY+K2tGXAS1ikqtzk4IzzAX8Un23HOuE6ehzAHASQN/D/DLOABVY
nCprcWC60FQpV/4RS8aW0SPlh/MUJIV26Tl+g9YTTYz3YsGaBR3rV4rYxgihcxPh
9GC8oK1oI69QucbVEJtYWiHZsCmDmJGqWxkUsFbIshnMBY16IiJOedQiphI/4prA
Yz5VQyvZS626qf3FBfFh8QxB3RJIXvrfDWnob0LfnodwGBer9UsECAJW9Xonrvi/
lpe7CPMZp8zYv9Q21smkqWrZU+T+hveHstJIgpisoj75LtgrZJyZKoj/n+bDRZLw
Ei4eMUfXI2hC3xpwTk+k4m2liHYK2/ap7UWXEQAXPzmJgQn5Szv2lVP0IX0yunAV
5HrToRBGO++ORBsxdXRPIjlOH9nCc8xRFLkxxM1X5pPHL0lqnGjX5AoNpvmX7RB3
sF3XDk8UwgytCkFpgKUd/sDdrI0GskzdfBEVImG0Fja5nxg8maesshRC49aEzMek
v8vP9OVtw/ombVQSlqpJhDMmPAahS/Vs4iFO5u4vCe9c/uc3zkCUU09F3pPq1VHq
WZJVQWNvCl2He2GLdMp5CEFVpu7vNkQTH0SItTCs1qhk8JckK2iDkBQReGg90PkI
qGl+0BjfTORqMAjBT6qx6FKo7TP95j9FJNmy1fRaaXyxhl0iLjwGwCYb3Es7u1as
4DlTsC/ZNrsB2ZJZNiUJ632KVawneJfPvZ4loCc+dMZ02XDawEaYq6nnPBix/lLX
RjP+94dULJ3oIiAfKWp785NdH6AQ5qrGlVL/GQ/jNG+ENSQcgpg2l7BQqmWEOYYy
0UOlhz8R58Z1xma3LFdHqIBomAApZGfqZOGcUnrRtamMkO6npWRwhOKlqA1Jlq5a
TxzuHd7S7KZRhcA11SMpOgcr2coROwTuTI5Qessa4+3HSIIPiXHjBpTYUkqQXupl
QM/3Rz4b1neh3kkGs5F7G7BDN5TF9FNfaOaXr8aDVXE7WkzkAaYSVcUgjrK2iNWg
OjyB1B+Aa5EdwOVy+eCSfCpad6HnRqII/UdXz/vBXU1T9ayvKhbJNNKT8pT3cM0H
vPYS/DZymzbkkr+rC7BScxaN8huBmr6Vo3oBpzvU9RuJF15/QaAIvS0pR2/yIWJ9
lQKgSU24/aeaw7WS00/pxjC+AxkSrYCkOCmiVKmtIiEjVlDO8W3GsCuHfxQPlwFZ
mXMEO7WowbsLTdiwTldmqv6Zei3j4I4/G5rGOPMBc+NFJo0AJRYw/PcB0O4fMP96
QjTY9LAEV/SUnFOUstu0x9uEwLp9JPuYi/Jp+qxdPVCPpMFWdrf5V5grRxD6F8xB
f8YNiUtlaFQt6kN8yrzqqjQeNqjXI/l0lfZwXRswx2HMV9+0NRGmWlpGiDIQhgsJ
bd193KoUfGiBXnqhgasEYE44lGPYDRdy6CZ6cfAvm2ELjeX9SktwPlLoLwhEZwbp
WC0rTrs8r8IATCSon7NyjOHJhWla53tJFkNV6uDqdblhXhxSYLW5jGW+4EBrkp2K
rWT0hopFWI0q+6f4WeUNZE+GgwYeXAhM8loJ9itFsTs8knkNaRTsBI9r0LRHDARm
JmydPOFKmDkgXdNZaUpYeftMe7iyqMshnaDQqR62jWdnt3p9EaBRPIYa7z04pP2t
I4LmO35Q678/ri34vNrHp1/phoIgnW3/NCf7OQUnKnC6XYF9MRKpBDbDIYYwzqPI
ph8ecPJNAfv7YBMup0HtxNqfbSGBTM/ECBdXQjHSX156C6HxkY/U6HrvdU359jBz
zsjTG+QBj0yCezpL+n4x1J7qC3MJj4AYTeM7zM23o8lWK+BJWbmNsBIO2ZbCWrVv
0Fd/73hKkTNsJZBMmpkwWBEZ5E7qCd3RgVflwHj1a0fZaRK8SEoLzMDOfJR0ieuK
0N7Jrw6a+UwEgXVFUvcKI6F4ja5QbfuB+U1aKbTiiSummjLLclvNLtpK4MSPWr50
0HRzEt4T+OInMbkHjC0ztspSmwUAsFfl0gkIq3zyWkNEqmeoYqW8UyBBKAgc8EEv
nArm9mxJ5NRKF+OPdEiUacwqWX3MOVENAulwFalz55+JwR3yZFoogjxO4K4l6KSp
UN3EkAQjcisG7YMEdqrz593qUBubWFg4h2hY9PD1+kMB4KXC2m0zQi5iNMa/MgsG
1DaZ97n1Gt5M4TtB+mCPmOa4Vl9o5KUOqGzuc8JIfZSCuI/952uNUUuwaNRA9NBx
xfNZJVazd6mWhiXF/47v2cVSZMLYtTahJGCvlB6tPAHT5390dkRglOScu/DVMgE3
hlmMZuwZYc7rwInoKT2VR1VgNUktAJaSSsP+zL33tsfr6mUKnv3zxj3Ce3J3JVum
wQDOYRMApFWE4ieCpahUhJN1atgy2nHsIhjsj13WjAsN7p3vR/8KilKQMmXbIquR
zsK0HNl61UFNJMjbmfRgpISkeN739tD/yvWFDUUFn0GGa4i9suusgbmwgDeK6pM1
XFQ5Z39i9RfHUzqJPI/+Y4mfsgT7uZ1ET6Ky+DfISDyZO3aiPBo2hZiFDc+iZLqp
5tnQIr7HI/HS6n+mzLdNrxJ0y7ZXRB00K95G27TTzL5hFSkxnfDyP5f6Z7qtWZX9
so5DS7qt8MbjRf8yk922NFHYw21l7jkLHaZu0QbM3B8mdwVgW2t94gkTD2DwJBC9
ySUsPSHPO/fttJdnZaeJcU18ETW5r9eVfDTNF9p0LyIWp3CpEDCeCjIhLgiXwEzY
ldUQxVr+DcwEhgzKC24/+GWYFv1lU9nvEqGy+e5Ny8WhfsrXe5qCt6Kl2tnR4FcU
6Te5gBs7n4Q8CUUvGBtr94PIyZGj2+4h86m3Rry7LoLCEj98lBAzgLJAqMDUsi/h
8j8Jb+UgO02bFI1A4nj4gx3N9TSqpTI1sfdh/Fw7dcHbDZD69dYzbH2WT+uZpDqn
9uBlFMWpVGHMWQ25ijiANn1p/uy/RV2DjiEtXUwvDofQ3UjVVGTT+IpApywD5ZkT
G91lqtNR0GfMbZ1btDr2rSNkiPCN9xO4I5emAJEWMNKlVTibKCAAHMVZMr/9NPaX
XziorytCBO7P9+BWC2fN7qxH+3Q7VPFyxmpC+mze0p/ov5fweacjVamGkPZIjwtU
lMVZwJXic3lAl2hNXNwippROf1RmUCIGu3MBTf7M91PWOyCfxZgV15RMJje/7Dac
XA1tG1QXoB1X/jhO2SS5oIW5gay4WbQ+cspJX4i4h1MCuvBMbMvmobuf8wZ8zUzX
WptE1fuFJ+Ur+d1L/ruD5bP2tcycrnJBqG0RAvshDMQ+NYVMP6cYPhT9GmxRrawp
LTeQ7BSw9NclYN8ykx1h7IUwrWZafP6VW2llTHTiNk5RtiXxW8A4W/otzqGK6kMs
hTAp7e5DoLuhZK5cdb0Nm8kfsR9QOuM/hxNthEax/uoeTnPIb4sUQljV9jt880sd
6iBHFXTVkR8QeYHiPras8mYHMZc0UBSEP3PwvLHn3+H+6KALxpfoOlH1kctsU80A
FAU4YhaCzCmh+4NRFbjR/ceTHVKBBfaUR7oKfCpRy6RaPq4dLaU0NrF136HeOaJ1
DlZclg0mK3Dq0G68SFAxbPF3rxgSGpXmyiiUz9XIqCkc0i8gxvo2SQTpOLYcvwM5
jgxcnW0pd3JwCUzdMSiCjto1cRjW8pueLGA2MCNgPwnUmy/VhLnut+VYMw/Nrnfc
Ru/adkWtotorMk/cGvD2dSnkczX6tsX6qyQ6CB8tycqb102Eo/8hUIAQHZRuglFU
lElpDUhl+9BNS16z8AIiY3qYSL0jXOWLRWhsz7aWd4BeJGO6ks6R9iEfI/diA5Ay
Pp4g7HFA5UClfuSov3nDfIPaeWHyaO+6f+gmhrfxGtHtJOKM0nbQTqpdpByczNjV
P8jHyxYn0UAyIQ3pMv9njlTOMlZw9E2pxLywNtfLPZ1gw3A8rDwMj2rXEKz9uen3
TvIddTVDs3LpHnynwtrQli2M6fpTDyKTF3KWBTm6wEHOM53DkRTcfvNsRZlx6Tpl
q+cXRBpolyGWNmJOp2fFfOnigQcOID6v9dJeUfUe/iOaKd/KJqk/tzrNh2mBTFtH
4QKvQ6JpQnK4iaRSQ226qkDL6ewP4enZLJzIINWlS96obAPX9OMrMGE7W+ZEpj+d
net8mOkXSmRM1vWJRdt/zeK35E8HuYzwgecIcFc0kVqcliysXV+Mb8GdtX70pK7x
ymV4GwYukWNpS0jgBr/bU9Tk33Oz0CiqjeNh2wNExKB3C+Z8FEdZeqB7QXafLPwX
sWZFJ8pDUneaNvrr/NnuBpWQdMeM6BoehYeoihVZFjpBi56IZsBQHuSsqsfwuE7O
duH7DinUGgpLyYqoqzc+yB0mtKfPb7gPAwXPEzsO1oANcXFpQE3+RKtWwEXtC+gC
PGgB+RzbWKrw4eOwRHKjoei2mOH4Jpc2rzBcSDQoDAYxBuA7idmpb5ic8Os0ZhhB
uT8gbLURs6XxJhL/m3yVrMIX97ue3CdhMhv1GXCOy/c6dRpi0UqwquiF3TkESC2n
KME45AsW/Y7ZkAsZudo3pjZ212fhJlG3+mxo0b+z6cJ3EKiSpspguY2D3M34TksJ
PkqBSm9SJ40qmAF56Z97ohqA0buUMaN5UAtWA4bwo+VKNSIkfmhrZtKQEJQ13s8e
xl8VqD/p1hLQ5gvZ9vbVyk2vOes9fPKFTJCsnW1uRWdm+kPiNTkMwjoYB68u52no
iEU0Yp4Skwu2DhBUA3vIWBk8668L3YRs8cpEhMBcW1E35ftev3B/6KSHrxWtJVOb
3EgHm3C4d0IsdnixW0p7yL5zdgJWXtywsagDJ1Y7o0FzTH8xSSKO1FlBipCp098K
686yRIXEiryENZB1GU/noEobF9BCKuoqn8+ZQam04HAf/bxfANsbUznavNZohtEG
0BnMmOeQblI0+/9q0NCYpGhX2xBZ2dags8Eyp9/GLvtUsHIAC+ibzF1xABpeO23+
yzGaXBQq5Lg+JrdjcqAEVCPupKc5w9EIbXOvaSMkot8o+zEixM6Qw/oI+6s4y+pS
JVvXOmD157jT1LmMTHlCylWbMXbVvJ+TMKH0dwhL+ItvfKtf53MqQW/WJKMS30l4
ZtJC/Ss3sDf3ZyJOmOxREF5Foig3INJfxD43q8gYXJrXloy35pXEkdDoEPYqDzO+
1TMM+gyzbFtWC2nM23b50IOqdwjmnD9tkFYJ5PCnx6VQ1XZD+UlnYtGWRXR2WceA
YZ2SVIm5iLd2WKio63Ugi+Tt2szNZVXqhGAszof1HubjdawNR2RDrQs6I6ApCZkd
SMNASBuwIWPNbNY7unWthRH7lwCSCmAKI9WzLT+N7c/+n6h4VV8EzLcPlDy7DeeL
ibKhl0fi1FUz0P/OfTKfrE8zKMSqTR5xEGk/2GZZilczHEaPe3x8c4501VuQiNmK
9cR/E+/odbrPZacTmMr01nkwwCIest8YISDnUtkbi+Rr3weGLPhGlovHBCNEQvR+
n9EqnDpNIm/Fx4HxAUAtSTdgfu27IItyzmWHqn3Kh5OrNKwec4qam8ns2VzTURiX
gMBSewZckHqInnjVN3D4zOi66s6bbe/wiJUJAVGVelmm9L1/xiFJkO24M+pVIZgh
k+6TcH5bBX3IGlSuKnB2ovVtK/96+b8OBRXbr/WCiNc9IYTKIGd0vGC99eLKa4ks
5QR2KEwwkQHyfpzWGqwyi2419FiuZpHbsWyCVvqXHBzvHTRoFkvNYVGXclplqu0E
jC/biyeDL9xa6cQT8I8BSwd9247hfsMI7A8V605U9KzmsFovsLoX/lCeRQI5vwYm
hj+qDiewX3QpaQ4mI8kMcpnNy7tjahXjWMr0vLmVC7yF3tiCShrm7pdYG0r5ckmR
xyU2P7N7aQ+uoS7OPSNs24cR2cl9/PGCT9yztdZi+m59/xwOWNZwlkw5OvGiweTR
MhiWpYCQRqDU83bL0CzuZrzmMuT9EljZkY2M+tR7FxFKnQ2xCGS/TJP7FK7nM+kr
ndkbFsXpfGs1x1cLciUM0AmdDNpS1PhQP7uM8poRrAtNpPisGqR7diGqjuIMoaoL
qH3HbdZ01y8fir8ppuWR3Dd43AdFK6xi85QnlYbQ9EFsoNLwEAEGZEnlPtcK7ZM0
sKs4tLF5FviWbrcGrM9iB1SnWt9vEiJ/lqE8+J57f3aZgj3IHuGg1/ZpaT3rfFEP
Me103nNepML5z7re1U2IF92H4NYogVqH236JL/G4zYIw+crV/6pAGbf8LJFwVh8c
U0L38r/JoUSuH03beYYJIpkrdnS+sT7yuvvctBSre9QQVhpr17niT7ew53ujsuMa
PJemKW7FzzjImJsYzO9z9n7g27FLgAFHRUDMieI9Gj1NYKJmyLdA9XVwcd9mGNdQ
FRp/gI7//NmyJH7DaVn6I0KAT+iKEW7HFy5ehUsrirGapsq09D9RGaVUXqVCQLvA
JmpR6PqBaAnxIrInyImamHYdmoEY0YU9uV6X9a9kyPz5wnOYfVqAkMPoILrng7ST
jr8ABli6gbRZSDFqO2dHf/pprZmTC2Ytp2/oCsHjFGfoHeIAfEpgdjiKNOqkS1MP
lY8MXRiVj0nWLvUQ9c48Pp2HsG38IIup6mRs9G6mAJKnhNy3d1UGYc7AqYHcM1X8
ZMMBsbNFkXAOre/5TC2Hx8pNJMmPrznjWMsR9L5Zx0D1stMMSPLtRyJalPBHnbGe
9fhYnYkFvG1QFeMOdiM3UMBkG1GqxKRwsVxlLVBPedLbPMJ3VnMRImi3NQ2j8B3J
r9l8YYofaLauy3cAtl7LulISJGk3JxUQwab/wxyD53MBm5/FuxK7w+ZI2ayxYtbw
RckPHjFhKwCNEHQL2R4nlEPTeRg7DuHEh9wb3N7iPOfCQN4EYPOVZK2iK1QR/wwX
EK7/zwgpN8LA1jyFD+4PZf8g6XDUF7IUUKKoTJgLtonC3/Uq79bvNPxcMcBgt2wy
3T7o9ZKrt/66peSgzCl1kvwxsiij/fbcNIaBV7bhiZihltDyZ8tDbAsuf/B/B/cG
M8UIJla6Iy+BcKtrfMTvB1bTPNlO3qPKUK8YoANfWNoc1+GuGDNE5SMVA5gY90Bl
BCzHqfcxhG2VKv4CrzY5jXPOKaZ/qu6cbloWPnAaRN8kIVJ7Au0dVlKkaab2Qul3
/77x0ycit5RyEwVmIiDfTXqiAeMrwDCqUFtSviMeLb91EWz5ThLSDN1PhRGKfx/S
oV02FxAfn9b/ATFab923GT1bLpIpp38XeVugOlGwxxHrbePMJzhJjX2WoVYoqyEi
MtLAecmLkt7uGYU7OaNZaP4RqZoeh0rcavaDjvItdQOIZ4He8pRhrkNxyMFSFgcx
FLuntXf0F892QU26AWjziopicWUxYK0CRDKVhELWS/UjhQ8dmpce2CP3MPL5LH/N
7ZKBdfl88ZxpZHiZHaNSbnM06pmw9+lw3P7BphHiSUE0zcH++6aiKI3e/YTlAO0k
ZONBJWl29C5HzqtPSTTq4eeXTc99kM/YYUZh4tU3xqWKV7GkMaM4CBDIhoq1l8pv
5XU5KzNQ9Wbbui+1kMZJrnQk/GCiVd1rRkugiCQQRDkyLbfYe4BLuNEQypYufSDk
a9b9trkP+UnEez6LTsZwn4QPhi+T6zAvdBIOo6rR/e3T5vSqB20s2rLIaA201F3e
xtLrP5OTWWT3zx5Ey8scFW3MD29Xk+IBMpoRTnj0R0R+JiIDCwV0ysbEtgC57x77
fL7b+MLSMyx+9KttXmgbyTZKgdw5StDE06xIqiRW0AIITTbrwqioawajmVFQRGkU
jyfWa6CyS9m2mL/uUeiL25ZmtXlzEWnyFOvg4tyjFQhVP4S0+BY9yKw6XVG9AI79
kEXv9FDXoUNwfXcF3WPSNLHm3buIeA8UcXUPyGERJrqNVihQkD1gVzoqp6WFk+nr
A+ntVgzJDQGsrSKgfeKJNlDKtOJbv60b8QUM6lXotmLZY1sm757tFhH35L6IUrMW
O6ERdVIQ4eEPfGLuf0RObdPYC7C+8FsRf8h2s5JyPp7oduoHGcWLbU42Jwjw+3ar
102ZfQAIp2RXg2nXh6B/Mkv+u8p1noZkox/WOV0bQDdX5CPsqQw8YVQ2e7An+1tq
r8rl/+1v5yq4kcqSKv6HSv98OJfEq0OBREQ6oBs/duwEuIqgex3X8AJrHuE6swhC
j7ECtSHgpW2GGUJruFHj96QXaVckffRT3XJQydkJCEEGI7+J8THtaPzSTkNxxmij
L46BJghEa0w1i3jsAAWL9bBz4oL8m9Nuu5qBsYEgiKHqlFWZjeKFzdYDBkDcb2wa
UCKHco6jPeiTMPo3RV03N7Wt8FeYSByWzcZR6VVX/k3jUiyGvKnDwOln+tdqi3Rj
N5ObOInMGv8GgZVFoI6g2uSfpDzr86L8lZU4I+zoS9SUC6PJrzp+D8ikDJc6biXi
eC4dZvugsI6+XhFSXS6tjpEsQg33FdEaQURtg7/bqKBAiMTpQOFsmJ1LcFWUTtYp
0+l2Zt7K6Zv2R2s3ULv2V8fQ7hki7y8ragLiqcaFfkGdEnNpC9EHyUqVGe0l0PBb
9rN9ilEnBpZknsJOAKUA386lwZ4ZTC8CV5grctnFC/RAX7a+/IupYwZfg63vZDsN
HHNbsE2MczWyV/ZWG1gRjEmKDNb0h9SJBRgIAmG1721WgepwxoZf+38xQkXQ7jgT
1yeBgUClqziNGlp/ezoPRHDmAHvXPQyAiiVAlWrgv4XPrJtB/TsFkgfzifLeDi3h
aZFPwgMuGTw/FICV1NQB6CcR4qlOqyzuhSevsYrO4Ifq+89flkDCzqte4qUqaeuR
acdDIm81M1jYyKQRzSgNqFu2FpAxnS7lTegW8Egft9geQtMd7EgfY1SHhFzlJ8h7
4S+GNyL4DX/tbiOWbKjfBVajvEH+A8snDcoFAOe8eVxG8fog2N1ivJDhG7d/lVSJ
I//of55vOlQL4LH1HCI1MILSLW4IvxoBEQaX8bjdKIwnDVfQDi3X6biz1crFAsyI
HzzQc50zw+TJKl+XnK2wt3TWnW1RXknsu7mzemtgqqiVry+DAN8aymiqCDIAg3wj
Ajerhm0QWDD4Jgb3vDpyuq3L14Z4a4wtH2s28Xd5ydxA3W0JNdhMIAbHlX+l6fNJ
Bz7VeySS5YyIU3w5+P59CCA+pRPovl/eblcOW5Vzgfx8H+SwQ2DodTPIv0mcxsHj
dFPVwXLeXUd8F8w+ETCd7ZMBQ2HWu0N44rTHDwjZx5yumcpF0JXgh3oXp5hsIFwi
YeH8v1OsH6lTXS7w402OlefWBB4aCWh96mgX0JedLsG3mwg3DWAFx59mYBhYIrUn
6Ij7jMwInqkiTXiNQ/JQ1LargCA5sMAhzA6e6FODEV/KNGRO+NaNr+QNHRJ7fd8l
m2kCoHS16LyyU/pGUXSWxriXPiXGVIdgJjz0EL3r4hQQRFFimX9lHEOI9jExJqJH
Pmsfm81zQg5uNKZM92+w1vdl1HF+HQOSA4ZCydBJ0wiX3Mh81ja78HX4079Ixqzu
UM3E00aruBfYBtipDCyJPm8bSXP3AyvCV7tn2Nl9ZmLqaruLA1hC1yoLlgv1Ks+K
WDFRPcVOesm3ivSC5qKpeck41s9koEorkakGSJuKNwAaEnpWsHjS6EtIxd8MHwWg
1Etgs3NxwpYf+Dn30PsXvTijJX/pXn8aGrEwXdMJ1DZnux5xlRybnw2CkV+KKKxt
tBQCaN67YXnuLmv256x0MYkiPdwh9BUSdNfarRQpoyrTFSzc3VmtrGOP9/w+CITH
1yFC2e3KL8xWKjqT3u9XvW6MmjyKVLJg/fbA0P0S2crM0iNr3yJBIC/T7+IppAZe
oRAJpb+LqYLXLJy87kYPqEWuD8C7/eRLlNPVpaNwSPNg2HAQncjYeXlVRenAFfCi
CbWUt759w4wX0kxj24ZbwCIgoX38tsnlAVO3Rj5qsBdQsGo50bSaIa5u8lLcix5S
WlOItiETNMMB/e+xueO3/u25fyIIYafUFgEf6/rITjBTnsX8MSJcd0tntGwFvaRs
Jb1/rNjIU6IzFjUE4pQT1nAhtaVyjTDReVd9awAdUFNK8ypVJVcZgSWpgwqfoIXP
YQ/OcaP/wmq0WJ2pcDFL+b3+nMVnLChGZZgkW3LvtewaIAZh6ngpiU/ueb5/kR5I
NTWnK/23ZH0CIBwLmcFzzwuJJKq2sTXuc17MBIvlNYTuQ3IsjJ0bohn/RoHeMIMd
i125hAD6tCGaEmRwyHLtW16g2FxfaG0TwFgFnuRT+c8ShkKO9nnkZDM0YA23xoho
RANWZZ7H4phuUXFYBKBSzqwwYRzD3k0Rr0wDNgg77ZYFXHoazixXDwlB9t/R68Tb
0AqJ38ySEfznThrxtBVkjCtzE+4HriwU9xtBBTuuXm/hFIFbGtc4tm7MV0jYB9/6
yc0IovByhuACtau4Os6SGtSzPIPofJTKkyrWTswFWz6iEkTPRLfQZmh7FX4hGxcs
ZwlZIQ6Zhuvn0awzKEfHbUu9iTD226yxb6v7T66x8kFzSd3GC7uf3mukOFPA4iqU
unqjZ9aj4Al5YKAU5ViEayzsns8hT9j4iCIrgiEX7Ix4T+DRKcDnGxwQVp3EWngw
gT8ZxbJ/gYDTn72nwbxpqcDP85C+ejPOI+XrSEBDQRdhFuIVqO9BuAEUuNDJ/GRy
1c8Ipq3iM98JM/MVkWHXw6eBraml4ohGchrA/lB7E5b3lrWYEiPor5QyWvvLIX9I
NGOEQ4CQRAiIz16FQAcsjemvNNBp2xlWMi0/fBV21vTLUIxBGDg52xn8JbhNk7Wn
bOFmi6crrRfaE6VpbxtBPgR7O3AibH53nyVN7R3rulNHsTc42My7rMjwi1cc1nGB
f5UiF43xbPjnbRNVPFBR+p3kfs1pbLZQiKCrhEl+PEHEUxz9dV51JqS86gWOxg3h
y0xISP6y8upjfub7D9GyAZt15OQaDDF13DgfCeBsrgYjYerlJEZB7ZKVpEUmbHqr
dfwocpxclqJ95VeXPuLPflgnSLeGYJXZTyOYRe/CMOISxuYQ8w0AvKpjjHTPtQ5E
o4jke3wq28q4kj+Dgj+FGunN/qXTmZtbSIWecFwJmJRUD1NJvFgtnKQ/yl1oMGSp
moKXepXkD9djSyo8jPujOqbMRsi1w9Ay3PEX+rbiwQzVyCTKji3ua5Szj/Qboxtl
rkhW6feo/pR6HeJfZU1vMD1uiyL96ZVNvB6E1nJcGQw9D11KmDh4SBKclnVN/+kc
una4R076KYQwjPZ4E1sGAc7i7PgMf7trWRLNcQahADmUMBbhvJFX8kPSooA5MlyB
PQIjEtikAabSFOL8IIsHujG4mBqi2x/rzjyVcqS1Ardi2kagzyOeh3YqO40rBCcR
A6fzAVpuporQjpEhU0LtgOMKBu9B3V3IeYJ6iFlS7PPFy94kq8zfJHHGQTQit6Fj
oEUp01UgHBnRcmRX/M5c5ea4u6q8/mLLHqQPb/9lb7Udmlxs9a9zBoThdr2BOJhL
QrjWkz9Kxrzbi/a6LdeT6AIA2PzoJ8fM26s5ebg2EsdyrJsHAUrSUYpGuSeSLoHr
Ven2HsRaT5zyIBMWpCmOelonT5OTXibi0GUGRDwKERH9xB61I89E1tOHWJ8Y8UeP
KuhgjFSnXXbnrrz7UmBMPhE2tPtBqseRe7+Iy3OUd7KhFeUCUJFJUTGUMahVYXxS
3l6kvyAzrg8pl8Z6+3/3crPJ3IGJAP4Ew9ZrfeVqhdb1wwnFK6dnnFxpzV3xfjZd
f15BXmXhlj31OdXcHQ1fmZSEY8s3hsc88xqTfDnyCnMKlq0za/gdTr/HX3D/3+UT
oseE+eWkiAFTjK6xI1GGp0DAP/7I4WBUYLQ66xm+jthvsb3o5pMSY8wU06o36vUR
kOetM4hhoYaYRcCCAVM90Rux1XbSLfDAyRK1ZfY0emy4He+M86ix67AEooB7EIhF
vusqocANBoAv11RA4hSChW9zv+DwMitxQrR4FpmRVVxAOd8UwlRl4tJbb1Zqqa4m
sTUlQiiJSqhS7RIMUoTGiWM++DHhufFbLlm1BW/JvkgdXOOIMEwAoJToOHvznmR9
Ki0iJZ+nAPCfI6sG2K3e+1w2aCkmWhPMB1ovmSUD7yMYy+T8U5j2owmADSJQ3kUJ
KtSekvpszkF18qE+XqELa5N+aM0YlullKujZf3tsbgCcEkYe2k8+8Xerhq2fWxBm
kk+fZMm87Y9yqUQEJNoOzcqsP1A7DTMCSk6CxSFvoVxnluwdAqRM4XpE/XZK2SNx
jqhVTLkYp40KjUaIArXNLglz8+PhJogLsbrtzk7fB3slnPU7vcVQZSzQcGOMt26n
U9HIXylTtVrIbfjxbO4lTU/SgOCwAEKxhUg8/8UulFsUvx0TjQOGTdwhqU2jS/6y
VVjSnBeDWM+irYeur5aMgCI5Prao4XHUhpNYkzEUsPYPGwn3m3el+6gclA3cEhB1
g8Ut+CBXLuTEbqZOXKmV1FxaYg9dJm3DijIbyW3Tc54XlqL/8UFuTrWECEv5mxLP
iXKbVjbn24eFAyV65d9yzyGa1DbWjvEdZh69xq24SlFj+Oj06rcxHsgg51QznLWy
LvmKguZS9rw8rPiIKrnHDPFjz493Ohlj8oXX0yofiviCOUwPGLmBXsK8XPE7m8jN
fKqzPefrPiwBbTQD3O2h4wuoPYL7YQ9JUbMxQrFlCq79VtzyLU7XI099xM1BfVHG
fEnbVM9v8ycD+igbvHxxHu27WLcgHo1DPG4RCWmd31fBkGSzGO0EuRmlAnlHi+qI
FG8OBrQa4Wl5mNYhk/i0CLhGEkmJC/cN8/wiY8Mei82mT7DWH0cDXhyG7xzazPHc
mS4Xie0M73JbPH918P2tJtr8CM/G+NskoG0vcp5hLPfShzF7/S34rPq6FbuGX6R/
gGcfqIuOsPGnncxg3rL6RSOYMP/zgGnBJ0uF3wVQM5wAesqYrOvt3Ol8A3dZ8p3u
uc01mRIPfRbuZTo/7ooeZDTYvWdDNDoHiaJEptfEBNqt6ArzhVpgKzb4PWPHc0dz
Kz7ZZthWD08k312e3MVxZD4cxY2q8xFoyR/CXMTCp/5Ze+7RDUJSb86nLVPzlEVJ
GVRY4szRVm2t1J92iU4pF0udzNFRC1RQfL1WWaH8SuJHqFd1TJPhne4sGdJMuo0w
5B5v8Af/17HImn5B0ktwuI03zFKXkz+cgUUIB69HVi62VZhYQso9HW63KisekN0U
eGN5lg3WQ+Itdt0yUDkh+K+n2KCFMhJne2S+xvfTaIGBB36VcTEUBCzjKFPzMRT2
P+H9kpvkFR9Os1On0jr3cW8pzgnMmJJfvtpyOcwfNwAyuZzHNakRQ+fvVZb6Kklm
dR62Nav2jBBVcFy6rG85IAjCOmPmrMGlPhftKEFTOr0ctcauTP9V6yXJSMmwR4eb
L+P2u2Nl959F8+V2P9R6SBsJ2Wcaa7BCFwSszZSvXKwr+q0x80AEcyMWXfPtx+kp
RerOQqgSHU5FmROg8e1askxhhSg7o1gQezf459Wpcpj/P1nGiZ5MKH/+QpnnXt29
9RcYBaKe+5pwEOetfJgY+VfAaIUWkxB7vc5lOnwN8HHa5n+tXU0l2zru7x2QiiYT
FSOk8ac1TVpDWg9HdVz9J/caVMKJFEGhds0StdayLyl+2eBy+tTjR+/5X1dsRZbD
p+Bhgf6u0UiyiVjwi0GWRtrMqf1R6BCqnxz2LyAQ9X9CtI9TmIuExrBbvqAnoZaf
AZ8delejkI9+cJP9ywza6ge8aknpyzumuRmfH4J4o7J8VdvIVj50Jh02xbSPJb9f
0jHTrCR/qDsMrR98VpKg61U7G3HQou+FX7NkM44E1NakpJyvhO69CiYDns+6zAgq
R+fV9qy3EEBv7BZ0PyunZzRSi9KI9pyKVu9XP8GJIx65p7RJeTFwzltOx0s9akdj
Gt/jOn8cxNeMziTUctINGSfMkzkcz6l5npWwdELdHxnY3w5qz7LR1VbO3OzV6tVc
07QnQunOGPTXMQjWeTTfOVZesb79FHazexjKKe9dtYm/SgVRIHcr01ppDUgF4IHE
EmkUMZzqFNZvSNVDQm7fD3cMndwMeHGPnlPehxd/8c5egJPkxE9dgJ08XLwNnvL1
QHDNUrrUZj1Dtfy494LfAYg2KWbO1QZ/lJulGdwwitJdkDjCNKDnoPVi4ztP0og+
uxaPTUicaX076UI3YwR+t5j0vjAm5wM/pVXIHyltxuDYAhrDN7jHioJlsUWHBNT/
jIFiibQKmz2QYV1HMXir7we8FJR6bI/wgeV8q6FEWJ49ZdoENP/cbgWb2pGnEpWh
N/3NKORwhiSabZONOkHW9vbl2U3mrTk48pMonHoUEsPZCPVtjfATYA/rNapN/ZNz
RIJCDgfAykaYdUFa1YnpxV81TIDo3AnRBzTpSaaXkWfFCbSOYq40gG/xyaC3O0J+
ead8hsdLDfWAftMN19UpeYeRT8beUEg5brOMw64rFdB/o/5Lws+F2NiV/Ys/rU/t
oiflqdgEJHOLcyQ12+4n5JkHK7eMYo2dw9S2NkR/IHsfTs9tQgviVyY71wXbNx3M
hvhs+Gu8p+Oug3K+lP9Un2E++tCIkUGt2hKm/xz2nw6YdYhOMKnBgQM8uyH3Sw1m
IwfQ/zit/MVJoz1p0O53KWWFX8PxU9u2eHGI9usLHIk/mU0jTd38nxprA+Xs6npt
mLV9f6TUbIVHdvB6PRVBjkiPd+5eXw5sa/aSaRxfDDKypARydNBxo8VtEQwqZojQ
6aBkc0pIS32NaKZHiQGsmsV62few1LIdgZ50ykx2JlGjs3NuzA0EZRhcoWNza/J+
32RC4oz9RL9NxWdtpY4Y+ldCoFPjGuMEhzSYKQnTrARJ7llheFPXHJtCoMAUi2Uj
NarFXT6yW9N2CQTnBN/ASsOsN1F/tsAynUhvGdUOWhVf/DnQKIkeZl9Yg7DoLFhS
D1F1UvrqIcQVSI+BtDrWLucSTqgiqPdAGQ2FDkBwwJ70eqx9wsoi9RRFtlC/StJg
Jhk5mSO6QM9NVrnT1Ss6Ekcow3Z+O/D4wz2e8VXa/CfbnKqNXtvbcTJfPs8K3p9N
e/iwHn9qA2itrJbuLn+gFWRrfp/lkJv6tV6pmZdPpEWURFNvi5QMd/oBa5XxBGMf
t/R9pVzfLV5HKnw+E1feBQvTune2yLeqRSnlr9Ep21idUCaKrm4zNW9AUxRd3GKU
S3GaTztIdEk7/lNSyfUXFJgY3UceSrs0yoj6bbGoDjYv7rJYK3Ogjm/bkuM2Vd74
naSaqXE98LHOYmHEn7rb0yrTjZqycugYumh9+OURMnlcw/4sp7bONe9NYUMRshtr
ZHuAbXUlAcXj5x+RPvkeajHvw7GP6kj3oB3PtgQlkhEgdWDvg46vIWlVdH+5u7SB
8T2H+f07SkD+NoqlJ1UjdufCjblUNUV88KMbQu9S8IcNi/K+JxaqDJyuxWd8GIMj
eEzcJmOTXGDru5a5KMDgFFcPRntikJaofvgI9RpCoFpi7CVca/6k8SL/V2nvFZL8
g21tH7Exlmyb4s3vWHIcqQFdQok87PDmUTGkgNkZnFgdeO6htMJuxmr46BUAHbuU
l4qykWJQR28Lh6OsX9MrtLnPLXlgveUd0D0Sv10n89Iw1LcAfLXSGvz7tPQbYG5d
MTmKS1jGakooh3mwKY8blCSbW98+/XkwesgwLbI8jYFhNbCS9OzlxpsF8EtvO9hJ
wr5TbgFOq66+ze8y9QZ2gMcW5AaiZlJAsv2bEnx0pNn2iObL3ivavLvWfsa7Uupd
v6vl9ie3vSE8BQZJhOee2I3K0yZcmbEHVlmyeOl6eo+P7pAjmof1jw+WLIKZBtTF
czLUR0PlSU8Lt7KcFfjfZR5sCBYmmHNCDnnn1KgOB8gTvn7LKU0c8pvNParDj4ZD
rzRN1xs5nzIUFKFeoiRirwELjUuSrm0VvPQYca0Svx9UMPETj9uJy33AN0xJVMYR
LjinPZIQJzGy9FOLVbJbNI/Ja8bh7qI9Ois0M0GMUPzq1xh4p7eZGzQU3G+LQNWT
F+58tQ2sMAlAM2DlItoMmFO7EU1/kTqKvRmyen8YScrqkjxsDc+Hhe9XKtUb35HA
2CPd50OjI8ox+y0PnPLt8JbZiEymC82sWhJxfQjxiYDHNPgmvdydUMvOHAT3XeBd
VWkDUbiV1Mcw+Vd099J/Q8yp1bGHQ+K4kAAVCQuqFCUTs3Q5bg/X/bE2UkDMxZtl
KGcJrOlh8xrtPjYEQl890po2Lrzr7jv1Bzuz5mL7GGQoeskp8uxOIeu0tNTFK9G1
7rY4KZwcn4r8j0kBqd9VFToNiZZf9MnJKySC5SGscLZR4i8C5AlPTEJ/AEeaDN56
690Zrrl2r+Bxhk2U0kYe8FUc2mLGTgv1OcWFe7AvvxEiutyuwFhWBmQ7L7rJfkez
4FHoTzGV+xCsFwuEn+drBtSL78696sQUDS2amwTcF5Q5V/b3rmuNExd+564vtXV2
enXp+ALsWsILDrP5NBKjlI0af/kCvwyMTQd1yqfcFy3Ns0QDPi7kvVJ3Q626K62L
bmUrQsJlkJKZ0RWEf7AwxPIpoOhJ6ts6Sgui4wLxVB1Pth+hkeBXFtMHEHEl4b8P
wmksFvkzanWBtYjy0+YR0pvCdjIrBoktkb71bFc+R1Arxb/gC329Yz8ScrSuI3QV
ya8PvewSzDQwr9G6UuGpuUnZzsZ5HiGzKhE3l0S9uT4RpRpxQ+3BaU6pCN66RGie
T+7mrYHuJQ8xgk9CYGOC/dHP7D+E9rm9L+3bc5UVknPJz6WyGS9Nw1Pq7NV+q1K1
gwM6XU42Cda/iZVGz77gbC5X+d4O7DmUKYhazdGPkdJqLwuBJVxMZN/MN78q2F1f
foNYNnLjSj9UmCBl/IZvyfkl8LvUVUe6FiPrOJdFciYeDtRvzh7DOKVb8uzfGk5N
TUccOMBlYVpmXZE9YbZFbsb2gdPll6qmPg2UBrH+QVlQnhoCmDVF4QwPnk1msNsh
bQ3gNmnzmJjuMTQm4lIrkCqe/LckYgovzuBHQnQSv+xD2FYFimcXRCtFNF7bXtsp
HAYj7P8zHlxA3a6DsDLw/1IJzm6sHLkQNtu9kiFWmpe5cUgR1K2qabMHMLo5CQAy
24tECrP4OyK8iBdXOuYpTu4YAMZnBScaW6deQVHyc8v7RLvz/Yk/bjqg4U3ClLIn
13+TwOW/o0NF4pKyykjiGPbyynd+HyFVxGGzIL1bG+QmHPDJ7WZuRVhmPvdx+xOu
S9MoLog75H8MM1upSh66jr3gAmJ3De6H/DY1McUHWB838PXnYkPldRwB8ZQf5JLo
FJTFL21q5OYrnm6zFab3cYokUtiOkJ3rzkcXLZLb7JYaUpvTg7mBB3CLq1qHvzPj
cSWg2jow8b035Jykwb1uL8Su3HNeLS+qKXUAQIkmt3396dZc2Rgf5ivJ5HLl4olk
8AqWiO543E3UhxAYZ3Tin2fM8nMi9rTMGrYJGo0irPy3iZU9Y/gkcZIy36oeKmEQ
fCGwHuY6/7L5WcSbRKUVuSngYgg0M68eN+PCpA4bVsqYgBiW/6t3gZ1Ls0i+12lr
hkP1QPV+YPpdcFHJDnBMgDIvK+jNBN8trZEyY3Ij9sN1QcUIlZXduHKNPGY53ILF
VjZ13jb42mz1pReIuEUX6BqudVt+2eGWaC0h+afgWpY5ofpyYrMSJ1isroqQOr2U
T+LPb2PHHE87J5heyaN2ogU9lv7+XZRRPBMTibEmGxcr1InVoYVZwAPJZgI4BzNy
ROpeWi4qkRUqnXA5e/yExFKTiNFTQ2RzWATDl7GQR1egUVPqDjS1wWT2SjFXHDMB
DPWZea3uDwPvpK54sOTobGXBZwCO9XtMnG/YDewvUvrCyWh6cMZOI174xD4n56if
gotd11bAeJAt78eisW/M82eRzdlytjRWSw0JHW198Xb4EjSkFx49NlYNeGpVBLBa
atysx7j72TIw9SOL3Mfvu5P8PnNGiNxNEYXGtT5dRBw64zts8m0SGDKyGdszjKrr
5CrRxI2Mf+ddNGDJelnVgENFjDCjWw3gx4ciuTBXBWwLPiL4tdA6Nx+sc3B4CCKN
GGPdlPfalPKyX0schFFGPcnO+mDmngHG0fbdXH2ThWdxT5EMpYrjz7NMy2YRNmFX
t7TT9bEBAxjRN/2e4i00BVP7BwwllIzAOGJwXxJQZhJnI007AuKzStSJYqiMLz5+
zDSGeN+GJrW0w7EnFTIjxowudHLUr6RW4HgEM2MR0D2+c2spSv2oSPImDMaad6kB
vz+LGlNL8tTxSojdZkCA9wmzxyeWgN6ojupDSD7WB21DjtCo0KlchENU9t0q9Qc4
6K1DsWjtYnic0K+DpmkAgEYkqfYETzDrc3IPKc3p3LhnQoVXVKirHAvw9RbdUBi8
6O7BlD7klNNxHy2Mrs4Sfl5ZAIxoju9Vq6uOdlqqzMgUXyV3TGyK/xRo56990qqh
u7BZgns4G4ozjkqYk9hoxoz4PmiKtfG3noRpJKWO9Q2F+6sLHOjAxiDLP1OLEyjL
CrwQogCoSBujmThaNiFR7CRZcRp9Kqe7V6rDuQPvzKexNJ/gZEe/pr9sv3Y/kPCz
SsiJcnRejNDnOkvHB/9NQNB9ZmfhnFhc3Lf86ObP5TXHVD2BVHj5i1ajSIUl4pit
cwr2xtqtqseNdIA4sVlz4YiWys7xBdOgGpB+sqzxMOmTiiN9uhglxDfA4qnXQllK
wyNdCTkzURRivDYVZkEOBU/pBCibvHlbvCyaqbuLgss2tvSgyn3tUz6l1uD9FyPJ
HNQ/9OdGIgjmqAzKQnUadNpGRJr3mYrAttPytD0Xy/Vgi2h/4JA4vU6Y7LEWX5ds
rC7QbVgsj4q2kFF19qI1M40wuQ90pEaB/ErU2tjvNMokU686eRt6pPR+I6oqqV2u
CZOT7s77EJc55mn+Z32CWnh5/wTGoAmgvd9ovOPgJ5s4qV0wP9z0e2jHKIoXhGjh
uiImBq80QLSLgD3t2lv8Zg/rXZuhbJcMh0+3zZegTAdOiXyjEMPLv1eNq4zbY/OB
9mv9IZ6EEbAQ6IMaUSNVn66jEu4gsFxmiH0AeuyHc/Iaw52GNbD6LlH+4KfS+uIj
cMZUP0V/kdwUiRdNZJnIHGRqLQo7DyVhtEKgGm9/XyIhoi5i0OcfiR9ph//Fl7dU
AieWLhoWAhulNXbWr5KeNeja1xkmc8A+hPuqHQf9P7xx0d4bsonttClOz9QLH7tP
GMhcXvVtg6/mfSLXrOEd77Cm3/Bynw8CU+Y7EM2axxEwa0Fzzxizc+pIbO8zf46z
lSWFIJhyIJheXfbIoqf5e0qXaz80AfELNW8SoHz3tVlUZ9/cjj5tCj0jDa/femST
th+6YTUGgbEZhzu68nOYwMp00ZxlVW9OHboDfFq9ymyDiOK6Esz5G6FcR5tgKMy8
auc8aiki9onULprNphG7fBGs1uZhDPVv6PjhvYLV2OCUT8QUO/sWvKxUTcWizVvD
saQ79THgUXCyFdu90oMBl/cgLlHGz3qTaNYO/C4CPrba4mIgwoYnqaW2TTBk3SvF
ALTxWow6dZqS0B4+S9wEvE0iSAX+23qUeE7+pgIYqbkGagrMr6XYgr8BAq+RvX0I
8aoNc4i8W9hwOrSboA3TZpGQwb91J2HbYzrSRehjghr7t7USgzomm4HXxg/0mk69
4zj3fk0/YlSuE8InniJLRk5pS+W3iiFywF/fXIWIdlj3MwVivaaIrgdT9e1nTGJq
kEs0HW5nsRCYcfVq9VerIE3ITOISkZtyp1XWOtf9VQ8PkMw70haRzb8YIrYcvC3J
MsfaUTwRFBERhwUOpyLGWdFL5DUUFME6/jYXszZpuOW2bbuEuJB+1UT9qBjnAjZu
Hg0NcOAxVq2HrrI5NQzLnJvboOiF9uojO7P6JNeeWB+qz2RjM9Fg+FQNW5lHqjj7
VamRMVtFP4TufF0463+nj9mG8fiOWvisNvw97llIlFgEaVHA7Olh2pzVX4gI1ywU
J0Xk8X3sC2HKag3Pd496UdZHQTyR6IBSstchIiIjyciDEXapO3V4yAjlRj4lz5+V
5UXpY85EPI75rhmFtHBvWp/ErKln9b8kOzQ0lJZ/S8gJKXOLlE6SLIs1OMvmT09r
4IgqryMD9iRqWiwzR0NMrh6mxz9pVEE1zTiEXkzLxBxY7QSpnBnD0WJqab3Ijh0E
YsJqXqsxENLu+SD0Ae06Rs5Rk+iiE1Sn4TvL7ATZoeFaStIulUH7vKSnTLnPQDTE
xyOiixZl8su69R0F8mUgpNxz5P7hGJe7fh7GdK47dDzCeytKhACMiEeYWttuDb8C
siOpSjqOQNItMmmE1A0VidvW0zjTNMk4rO93Kgque4DWdhMU7Uw2zdqrU9qm0iDl
otM5VQP/oLSvarAKTINVhr7MprTIeL2erHlJDEe0A/7Qy3pdUVaBACleEMF5/FLe
jYgPDdBlN0hAYwZ3D27PNHkO2/haT0Tq1nMQYyNtYH3B1pO3vf0XhmwGYH+UnIWG
dlE7QhX7I2yTC/G9vQs2D26qgEk+s/sSNMibskKpJQ3ci76oaIQH+WWhx/qE7UBf
cEWA8QFEhj2aSMz3ijr0JpGKiWlnVq2LIPegHYZ6vbeEl86c2/RZXeV8o5LwHYrq
biJhfF1Tbk8zZ0kRhU9IWM7CllxKED004vvQthYZPMYanprRPLsGZJgGsG9SupSo
kXsvvNAxD14Njo/TviLAFNhW3d1yquYeNT0mmjFn3OUStGwvFVf7frwYzmhvzt2E
kMuOhJd6Vq7583JlMbwQLlPgVuvV12s3wgElxdKF1faFTeA4UZUtED5kDlbaorAM
UDsPKSlf1+RTZn+x9ZtfhD7ZgfQnkn+YMHRu5BCeXr/+Vvx34imT4j+rBc+KpvmG
EZn9dSDayuDUBN1edSg4G4LG1F0VzK6CAlibgLT8LYIpqLSUEtOclfmOGJCGUWkk
tc2n3Avqhfouty5SdX+Y6htnzeOwQHLt4Xmm5TdpNkdn09e9498E5ojIKkShveb4
yjhqtPh9wwsfbC0Qg2/clJbOD7bAluJ4MU1VXacupkAD91ajwMIFIiWyx067LDzc
iqPIteUeQkTkN/IYW/kciH0RNNRNo7B5KQhUS5vvjUTzihgJ4pXDQ5tSrFYfPxCS
MXALn9MVIfDjA98YWsOtBpnDY3eT6Pw8JpOkYwqFoMIML+ni3twDN2BvBqv40Ghu
mUYDsVjCndPKSP5zCo44NTfeRGG6M7tmnd5O2Y7ISnEP/4TpnOGfvCTPhTn0/lsN
hXuXaBOn+PwQqIxJt/iR+W5oISKsr8PJ3BzItgzWBzykVsKc9wmwA32XDyCJfQw5
0j1Aaa2D5tHS9F/wVHghpg8LOVdf5F/dpvrBq6Y2RgyLiKuQ7zXAG1x8Rof+NtH2
6NJiUKl6lVFf6sQKYRH9Udqri6AKTGw0NabQxKJo887Lu8Aq0gLES4QOR6G9tX4H
H4ljzUddi/rpEzJLeemeGOFpu42lrxF25Olg1mB0VZwxsdflKTguhXYKSDGdBeyz
x+MsiZqSzN+JWDeuJFWJ67y53fJFyi6/6AvT9MOCJa4bx8oeSIs25FpEFHOzM5cG
jPlSkVRnQui4B2yS1o1X0ei1UuQNnSpWRxmp9I9qdQ8UWCkwAU5N1uViXDwN5QiI
0Fj+CoqWlZxrqPC6YLv9umENOIP96IBkcpSs40h+LNsjul/WzomVWWt/Gv2mDUI+
Ds9dNM/3GxN4io07o7DTIWpPa2Il3PecDIpZK4txPosiKJhn/XcHCCNzo9Uoadjo
VbbfT0fS4m//3r29/diEwUqgonM249sLzsxDCk5aO1F3Rx5q80daP1RpzuD0e4d4
F3X2ncJRdd5+Gouexwszi/vUSb5FBayWHW90EIkWIPfjU8xRtrfYOiBcWAAieKZY
2k58M0mQhSO5p215Kx5BatBh7nCPBlH7Tel1L0Lxj9VfDmxzEOgcVlEMnOLdlgsb
/c0KkR9N8TrOIJvzNISu93iHDXhIYrmk5iZAlbKjXJQQbiUzYaQOu3W8uutCdqSQ
Nm2BlxXoMTu4LAO4vi//OhSAJ8uB7YB7vPepqAC8EPUcfHCaePYUc/5qvSCRoreG
it6t3vL2mu+EELRmozceUgpwyj0GOXesfmNkbXAgcZWuDCkMD42k8GrRRnNETdO5
q5OQFs7mQ/VDi+2Gfh6Ofv+lJE6p5q+EPBtKGSw/sqlq8GnvqcNVX0wmAtDNINgk
ZmtnyM0HPjcOJqzZ0cw9l2Iv/jF0yYpzCXdSPOujPySDw/VacnnY0PZGu4xaZWby
Cc48fJJigA3f/zptpUM11GzBX85MvWXIjHbq+CKHHdWDT9Ui+pIok9OFrx+2pPiv
m+S9R8hlmjfTZpO7daRcyFO2NXiDVjZez8NRuOkNAP2sl7A0VDr6j5YSHrRGa0lV
qqVhvf5MfJC4axyui468g0JT1wtgQ4C7IKN6l3p43hE+QWp72zTtdmXux71b45pi
bglNCcu1QKqIVNVCxCLeTjvrtXrgg6SjJK3M6XoCJYDlJJl2NRq+Rtl0zpWcQQmk
6gzbeMcClmZ+9u/vwbg07XBjWfbuxgmwlKRLkeAXZEWD2vpXnPOMebvEeINd5mh5
81eXbK8Z60wuGa0noSP45x6tJwA9lHuorg+5rhevEBT5hSR6DIqlm6kRT+IefRfc
AVLCL1jcuFHgUqZXKyKgeUpfCvqetfjpyvY8yNVoSz1WnLFjEnuejckGpYEP39dI
wFJHYVGC8MMPBUNYinjd/zXZ/uT2OlcahABQtAoRUsZ4HdBHuEtcHDQk4nS/jZhE
7V5/M7oZSH7TzxgEQnF4jOz7q11wQ0eNoqkjxc05+QXVuTjD+739SlzPP3LbfkCr
BL/BklXwGachpKOu66A1HktncsroQLjkhFEkn0X3hcjEq0ziPvYiauso6qfzva0V
rWTRHFqiSJLmDUZsATsvOEcEIaa/NIr0TTCUZWy36Gn53JzF3+ROU9sfiYYRdWLs
+LMYAeSLJwYNh1YWS0q7wqTlToT35iS78Ghv6V8eX79B1Vu/1Mb5vCT9gvJrqodo
h6BaoJv/Fa2rNUmB0lPKIqz2/nGHKgYK3hbb567RGcfS+yjRoOquS/C5QU7QDUcb
0RHMa2YCXD3yrFUlGcBGgdc/18FHH83QDGISXDG0usBSx7C75VC1fffV601n9JN3
BQ12JmndeZsiUaUvBB35iC1UeOgbHeb+Q4/PrpYZBqBnKcphJsaxfATWhMsdSNz8
UZJjcFs8HevmRIFEJz3tuN6PnJ9yHw2iXNixVwbFgduBKRuhKvGQgUHPGOeffMwc
HCwNZNhZNQTvjzzCpxKuGktGv+9bNjLQrEXOwc6LtajLdJA+l2oQpxJkgkdHXbEU
CUs1PAj/gzyqlvvwcS4pTSTuxH+fkqZ2jY5JbFBlDQlwoVdnSA/W7igDYTZ0KseY
UMeGlEI0yYhnIpCn5ArUM+1is5AnmikEppVr0KLIggG1Q0lkwZFhhLTrgfVJ8Vsn
n12LbSWBNYUKu3u+u1Dz4v3UAr+8/rfm3j7cBzS7aW5XBK7mBVRcOQGKT+MfJghC
L9oQBIBOs734F9oIir0eoy8ct8NT9ZsnVYLEipHqpIMULBiupYRlI/4iTbZZ8wmw
XX5xL36+23vd8qtVTrwh/LyFJba3uT2/y4LkTusAkvwcl0Y5QcF8DsiGMwGbePbI
rp0C+KrusFsoGVDcR/yNw+c0ERlYIR+zTclB5fEDwiBcg71ceMQxt6amKhgXnN/r
Q+xhzSbwpLZNk4Rksr/aJVpSwRx6n7qS3OV8zpXp5c9v+i5ydwMviKZuE7m3hAg/
g4e08q/RuOqHHetw2bnwxA28jGf5Ux1BAZm7tc0aEQBXTwWBMMzKv1RC+308kWu1
Amori5erdh1NCEAO9Xn6u64xJM/3NQNUJI1FJaOmR/JZj78VY6VI53DDnOnHALzT
fu+Ma4Jkw/LGqHIHendqjw66Q9x5+wQSS9JXq1JP20CTi7LoxXcxuSbKs5oHBpa9
5dWp8rN4JznMCc6JPjsRp9leGsFDXVqAxcggWMYK8F3s8M8NUQP9SR49jvDfE/7S
eNLwcWeA0LPYfWReHvXim893DXCq6aeElrjKXWGsNzkIihwWOevbjkV49LbmeLaH
GmiHBB78xjTROjOmSPrvWLducpltqYNwEOTGU9xYh4i1G6HbqTiPCU5j+A4Cy/DQ
9oB5o+y71VTkz+Lkco3Hy++PiFCWyoOMgiMNKX1PzmoJA1CiNvzAFccQVsTD9xeu
NQYALkI0gxJK+9upiUnROPUYSqw9UFzDR8E0vM3cYZewQwIld2QCjPOvDaFSJVFv
tAMWBeruXBDzBMOEDFFKc/Zc0ssMYscy0CqDM4U6ld+jUn3XyB0PsbbhoY8s7qa3
lt/o2YrnKC42dqdo79VPFv11y2p08399SRI+1zUMy+sZQBvzXuMF1SPjECmN1jaL
ULb3aFggTwvzzG6lfhDMseCnUu1Vl+kvUsX+cR8qeo1+xvIauZ4RurOKpcokGBxr
Ec0I4CTOwgH+wZWjcuBW2PfxSPlcINqTM20tGEX6Nj9J3b+BSsB7+MqklEAOpY9C
WK+dNIhqqAtOnTqUTuopSfqB55dcXVuFecN9BTgJzze8aKwecGO6BdXE3Pd2HrUw
S4Yt3seOH50L4P7nYESY4qK4G2h9BL431kp7HQCiXxhcY8NX77hYH/y00U4R+H12
U6W6qKIGNWVb7KP/5aJdNiiopJ3V6ZDtQUk32JC1tHbrKiDwrBB+e01Us7TvmhLE
5PxZ+zroDFxZeJ1ZIZ7cBHKWyk7QXGGCUtpo0tUypl1y8uunSProVOVBMrEfRWI5
fisKiC7R7h+KzEONdP0cgJAHGnNTa3Iaz1IPBSSyxk48qKpNv0SZgBcwbZ8fLbW4
z4rv3fGNjFdk5G+DMIo93AL7/4Ntysr1Xfshn7uzcPewYzrp9xlHFwviIPiXgi5L
0IYyikF3QbAgCmk5iz3s19v7t2ZApfz2ov8jfNdFqsieBHDmMlD7xJwoF7C/zmuz
9VBav/5TAbNeDLucen5AH1SWtRf/mC7ZQ4wD7HWUVD8C3QRvo/t67IIAkJvUtt79
5fVopiS6lDjFcTWjIXifZLbH44bpurHwWSp/mf+LtpvX+HKUJppMjIqUwXZ5MLe3
JsamQ0mTkZcWeKOPT4FRmNjVf5YWGoxVVnYkxXTgZHemlGBEJmI39NAbTBavYcdS
KfBUkLtHGohUKYRpeqoiWOKvNWqaALp4XK1rZKIJk1Li6sGdayB4iqfkiRCLafu2
J2JtJPsckkRIJoJRRerV3fDpGph5y1mO2fOKWKSrY/srR6RsfDLslDKo1NdWmv2c
LoJjEJXEZeEiz66NGk1Cha+kmUKA4jOXRsaLYNOhmRV5yfH0NsU/aSOaWp/MBlT1
TSgyQB9uwcv1TwCksEqlOZGErAVwVLahJAP5Oi3WPSNimmVTP0FU6suUd+zpxvAo
tNgLzjZHRJuxWu3aMYvmQOtwwtNjDnlZfTgYxcwncqofmz1gT2mvhvE9t4IH/u7B
xZUpstt6CW9tRSXcEOvdpxcOwNszWdp/aUcwDfRpwe5ZdE6gxK420VHuNvvz/aE+
ZhIayL4CURVEb73DGbOU083cmnQI3gtap72AofFhu15czzZ/GQ6W5IV2J9QNxYxk
8g79RdvpgUYj+wTu+dMIwPSiXJmI8GOqKGzosP6LKcpZfRQq/ixVkDd1MjeTZ5HO
zD0p0yD8Y2OIUs7aeqthpZ4XwLOSuu0uU7J76w66PcewChN5NS0gZR/QhAUUEHTQ
0XpZ4FQtgam2YPJ5GVycBsS/wXFSDfPrDfCFfEU2pkk7WfbIhlwz//nGWGTzlfqk
UREeO3cjjgYAASPhxmsVbNKm4zlLc1AnDUp3Zlw+4WIywcbd1XTMwojfAlRmN5yR
nJ3Wm4B29WpmcWK4ZD+t/EyWAUXkGWCSpHqjjHS+yZB1q5DBo1+nsvKp/G9UWVZZ
DkIFRShRUrIlT6MXQFVPwDVY33rUG095N9vqUte1Otf/2lpHDE4dUQe6zl2WoryF
WGKRy5E/rUcspG5vaSuDRsxatiuX42G7K5Yn/UpCx/MH69AIuek0NxNAZi4mZKX5
lMJmrt1pLoLW3gaFkT74PSiRK0/3Ksw1rZvwI3QeJ0iHDvBYs/+qHd78P3tZWFyU
sHg0VUQRBaHnLko16zcLCLZz6tEhPwxEXcFNpJD7CrUyK4gCIn+0aQ6kPeeQ6HHg
7zhUdxQKc70+rp1idpfrdsv0oLBnsKO5CPinSvmo8e3pfx+b6R57LcP7erSj5N49
Cw4tfHoiONrIOgvyepQGl+2PFgF1Da/tG8oQi9UBPS122wt57pWedUQPYTeoSZ2p
ERud/kxI7JWl1PF/moe48d1kyW8gkQB9cWDqcInhTb1YGvEXo6KBXSjrwTxRokot
UnboxG5SsWXDVGXP6yWNq99pMiGldOcltiCIufXac7iwObzCbIpF0MtpNfsDGr92
SgBxsp/sJIbFiqz5iJYE0MNUPms7feNgqFSQe0Urr1aXgo1ZVc39yPZk8Jkz4O8F
3eWTWskBTVYAIUedrzUI/wAAZP4xtjEbyH8vBlDcj06vEbEjQS4KOSAYmu8a5OIL
22aJsfvYFuBuM57tX+IHHddOBQ7WdP5u9U1l4A3TqE8F7qKg8u+Vp+PkluuxXkfz
+lCNOURanxxVawstZGBm2QKR/j0mb0z0RRP8wlhamXZfmzq2Mgaon1V8wlimTZ01
bQZhgQD1hyKA3NM9f5wbtZWVPgLzbf9vaQ+oxEtn87eJVHAlGPXiMdBzeFgqsi8r
94CAB3VX3gZ2up/o7yx4QUvzLCuNfAVOYpsRyCJ8thvk0FaCkPN32VjppjlFLswt
/joUKmUlXrlDiqUD3xi5lJ2l0OWMnyepmJWHPIF6SK2ByzxeWkzI9e9k3q9ejbO0
DircCYqGAHyfVcPt+qmH3624lVhPR83CHW01CGl5BQEqiOXPc9g9gvMA2O9J9Kbv
Xp87ekPIlYovCPuRUFNrMO+vjCV2ZyGycUkdJBR7V9ENhYZKl474ncRoVTGwrVCq
0NI1ecQMuZxT/VTfyztoK0IBCmzCAh5wV8rvkQ8oCotoQTy+7VP1X0Ap09sd2nO0
fRy+b+EcKBu+7lKYME/fx0TxKgQxZETZsGvRUw7alpLhOHr6hd8lHYUp6rMKHmex
xckUb+ep9IvAHIYj3weHqaMzBhoPd58jg8T+2gn5jRZUDjQcgKm4gBYGSh8QFgmW
gt7T8aipc/bO6El3Iwejrhil22qGRk8IE6raRzTn8fEke5iWidvOoB1OpPVVxQpV
RKv4KKZa5UKOhmGvso6rIE7GV0EF5AoxWk7oJA2YFircEJMB/jJP2KNjf/da6lGq
YJ3bNcwaEXD1WIsmq5chBiCVKYEAq6B5Ybf4bSDXYG6+/e7zLVis10Qik7Qs8Oox
7vkWyW83EAYpcc/gLjt+aS8PTrYgBvtkmaMpAi2nD2FOjgnd/5l0/dq8VkIlgX71
s8HxsOpL1EE5Ak14zykq8qKlLJwhvDBsrPTlldARcFretSWmnm70zTgq67JN83pr
lt23bST5vdS5WEz7FYiZqJKleCMMwG7sMFn9MYm3LsCgX5KiVHjNfTAww5W7zinK
g2e1+n0agijFknKaBbjps+I2PSwqUi69ow6gT/xQVzd8+6ESVhFx1sRK0fK5QnBx
ArqgoCaSCxe8ChthXDyagGx+7kWvDK24P63ewScp5FH2rt/deuN0q6NdONjnY46C
38j5cTNAKPFrUSGhuquwBMQiuFFulsVUfQcuCL9G7QAZl/hN681ws1u1ufn4MfHR
aSzuVEfBzdEUtELb2+am4nTPENkmdsw1tIuG6v7sUkCP/YDiZvJ7vYsNdboWbzJ/
jwUjF157KkbSlGAOCZ9NtOmF57do8IgASoeeBu5TrHZ/t14uOKEIxvZ6rESGrLI+
V7myuNFwG0T5XPadTUxCcC2BZ7TS6b8EqeFx+r83cdTcBbpokKe7TCsRAFCSA/Lw
wV/T8WzqxUdMF90Gtn40RbDzhHqS7TVTxWpl77qip/db6SnhRdKA/kZ12jrcipST
I4oemND5qwkm4RHRiXFhaEHlNbU37Tp1/qOky8WnZeBt/WzdPU/CWEashIDPmGaP
ICi7wRbul952hKTkGaQmLVs8bwXameEoWchJ8nu/7B1fSuUHkqAQckM/+Zmb4DNb
LK9Te52J8luT8wNxBHW/neyiPCOIE4d6DIyPUV7g7bd9TZAcfxUFEcqH5cvL1DGy
0INobV+LGaLnOp8Lv1P1QhlE6pkfXaCfcUbXaJNSLyTOlvIAHjuZZHQd154TDR0w
25EYR2Sb740qEw79zy2HTDLrWVedwBWkHuFgBfnD57tuLE9YrocfD27u4NS+egrT
A7e9PjcD7vUn2y0FgirOh2PiEo+OWIi6CtYzvutCTHB+b7LsXCX6xxQhdhO0awHQ
UEpp+7esPWfXljyjg8R0pE4WCVZbBv7PiqxHJFtOgEcogcuZ3Fqnd9TdAeq7nFil
K6UuS8qhWLX7IhgA8lMgBF9xHigyxy4bbbk7lZNxjCsT5Es2jsCxS3xVq3r35shB
GjOFYnmmrPCmsKyJV7u8ln87cyuBO7bJ5uRiMoB9GBIsIAcOfzZ8tpp+wxEt5zz5
sOIxo38k+lx7ekYHKJ4xD0j9AcvMahcdlVUvBiN+Ufu6aHY7pj/A46lUYWQ92Rco
4ED4KTeuQsmZzRN/Zr5GqFwYIQEvQ+I3EgMPLqyUpQj5aNLxGsdbGpcI04ob+RTi
+mLmrlkB6xU+mwVc8fytZduc07XhCPsX1LorSQESmo+WROf+yTL/uoFyNiVKUB1Z
Ez7T7SLlubMfqQSNToaXN650KiBz34L1HDwM+6otMcBS/7xR8THBhD3G+D1s/ZiT
wKK4/3KUY0S8pMQiW0ZnNi3Cjp1ZLpCGnyUJ/nPpzMzYb1S+wNB1i5d7y3Vlamn/
MnauNmu1OjzKYMojPOl0vvBzQ/YC8zTZOjNBdX3zlO50eQlKbhIFUglaL3noqV2A
cgnwsA68Qj20pVRcVD0nqki2IY9Iel9StQFjqPeCZV6WHKXtc2Le6fyIlUWh1gRn
tLXbhtxxg6PXrI+uipVVDW9k0QgOPril0Gi/rAFtR+JNZmZ4758QngtHCJncnRk9
2/iqlJVH5PNSwm5FJvLhGzEmpyrnDGg2O0J3l3Fm72/7JAuEblO00wttFj5Qa6di
mZu+jZWCcvtFprAEq4XZAsZkDG+i/F4ZtIKMOZmPADvnxUgYs4aiyA1og0ieebKL
hwvWpZixzPJGM1KdGSX8k4uylBPvzRMzfkpqy1oJjuWzpfPuFwPT6ybd9idmbXbH
dDCsEIoUYIYRc6fLLgRx1jP7fwABhLOVMeyMWPO+QPzCBTYUIBU/3eUyTBKF8aYF
l2JoPaiDKvykw/G6RXvLsaO5yYrULuCjZevnQQk3nZGEYlyAPTrCpQ0GnOv4R1qM
924xRS1r625detJJLo+4m8dqg6yJLQpXxT+Htlcc0fPU6a4odrAJMSq3YVz4uFtt
cTtOsvlvZ/1hCALujMaYioys2bOjYPL+6p8XMnvD+QnHRseLi2lJJJxBKOygM+oY
bkMlRKz1aS4G4SWXTTNIvw5801xP+KTEP/KhhnQq+PVRqiV2ZwQLXumEulPmIYSJ
/LzXVm57A0GItk6PLTfaKPObV+RKy622KwCzrU/jq34T0huqeis3t/pneB0tYhBa
2exd367nOKriwmithAnYHMR03lLs9f4tOR6oTSnBbJ4koiyGj0lcnLKqxPXp2lLm
1+T2abJVViR8OQ21rBNhNF9+srRD3lFqIfxUiAS1gRdBOYUlJb0CACbYK5kAR9Mh
olP4a63kzLQ/83RUWY+Q8v+qJ09qZ3uftZkk/Tda0Tzl4CBltVsR8TSFLLrcrTA+
VqXDSIDdGauaZ4RD2IsF7MBHnBiDFbj/08pvxqM0ekWS+HYeWTLBe6b+XvBLvRsS
2P3F8jJTsoqezhLveEgUbVLyFh9NwNZek9yvMqfjWatwodioEvAGr6+J+OX9uCm6
7NckpPMLCQNuPzJEzPJn/EBvPXGTleYIg0HxPGqyoF2QLMHMbRp2zsBAlgLxcvuY
9QUc18mYK1hvLdbqYr2ZjLfUWWynJWjX+N1uOPAT1X0Im+zWtIGdcMfnhH3RIs5M
2pY/MkNkKlY7+TTA9db2MKx15dP3jx02zm+dPPARBBRfQazy0Q88hdejWmEDagwK
T6z4T/wTLp89f6d8i9CRYxuSz1Xn2149PYQcec3KAfOHpQcCis34QUQ+R/ZwAUzA
Xz3s+ALQR86bKmuln0kEd8eHn/Ya5hRl0IRlxbxMUSzl4+bF9JN6S4eOj/A5nyVC
NmrKm6vnEShPqO9nRAO7h3PydYhlilkxnU7QNK9gDiLjk9MPHV6HoYXAK2eZ/QxI
KSA1/P36t0hIEntgiAkbnus6zVY42tTcuDKTMLuZYJ2FDtlS+ozCxmSfQ8Vvqq65
0U5uIEuo/uBJpS/5k5VWLvt7xawpy5CLd040PGSP0VX55WoBzYor3uIz5tQ+X9WW
EUwcqt8ZMCRPIf8g4oB2gegjB+6VkZCiu0d8VXkXTsmKDaAcWLZNl5DGyzdmQWIL
+/EoaFr9ZegPE1j4+bhk8D80JKRwUihgKXx5U0hsLyjx06ASkMBvuBrGTrVLhwS1
Dl9s5G2UvK9jCdyuN1skG/3/3Mf83Nk9sfg6GeekENwDgT0IRPuXysONvW+cPkrS
tKAbc1Yped9+iel8fIH0gQEN1BKRdvxPLU5DtoTPoHOSn3Tit5b5HG4hTWbeoiOZ
JACnMfKUHuYLBocxjSW2qSBH7pPiEZHD+UPAbOgjtRVh8w591wKQJxt3Th1v1uvY
fjwW72ARYtQG9gGq889iftd/71X9UJ98NztuOK9YaAaj9z+uasEsbb+2npJOEemg
d3kQmqNxvPBGE1AU+4wIWr1PSkOv57WqIy2NxNgZnZ4XLYN9cuiAOEDxNmmEPvBh
DDOknyRKgcdHFTHoX63TPrbpyk7RKptKOVOL39pROju4cKh+6Z4na3whpnKVFQzf
sOTdyOyJvtbXXx7tzOKVRyyV2d9JioeF2OlMQU+R+cKr79Mfo8WaS6eoT0uFjbCj
8HTgbS3cq15KNqNKGSdnr0Krx20T951Hpd7g8/tQ8/7oTAuCc3ux4iKhkeKd0c/+
YYdSAiYyaq0t5/u44BNVjVBk+ThhsIcB9eETmqCEnYnpulfd84gX5+WqqeX4TNA1
KjxQQWDyS6YO5lZtJecdV74tN2vnX7DTPLuUKCkHIF8OFdVVj2C3OFPSBbipWA4R
I3DO8LvTlwyI8fftwLGtlMT4cY0RbZj16TJwY3/7xk1DZQVO+0ri65ws7i2zhG9W
mskTlxIILeBOUCPPwktnMCFIOihPgaXu7grWl2AqGW+J6Hs9uGdVfy7NfpB2ab+Q
xwU7Ob2SNgcoeNA0PMuD45pXsfdd/TOWb5sxCt2+Qtj1Ys/k+76qck3PGzM6Hpt2
z5qZ4yMl0e/cVCGvXu26Binidk5Apz6/sEXHZjp1dt9QjHZ1cwXeIUE5y1o1l6W/
sarwE2qowdWi3p6cyP1BftE780oa4masrIypXhqbrMoGwIRCxZ13QZ3hJCkL54L6
tqO8DABWOmeHVjbw+cQjwS46fxcXCQo32kHuM/P14esMHd+qvWWZiEqwci7V9OXq
tNCMkXupE3wlLyHJ0b7XqVEhYoT2fYAhX7I33Lw83IGzNkb/E12hyDOynMF+Veo5
/cJmqh10yEtShD2sRwO8oN0/4sHfA77Egbhre1rXZphbPVBT2CLVOGEGIeuTXzc+
fj1aMGMGnaRFoAVme3N7z76K53ejoQ89eCgBre3L+gTfNf6Dr3MwI//4miwoPlDw
CpXWYA9Xw3ucthnaYu54OpnnNYmbwkBTtp548DvkWHeLmPWjFFt1puQhCZcsfZxn
t7EJRcYVU6DMOaJkocsYYeIxAYNOKya3m2WfPJMa9QjdhLqZNMVse6uQN77hvCwa
rlm+/ggAvJ09CirFhcwOV7rqLRNieRQLSwZ9wH33UvT/JpjmFfKj6Dm7ZcbY63OS
CXcxp0p/ObN4F8fBHIKo9oHHN4v+W/nQp7Crwt5SxDekAzbuaj2YkklhxGb84UXu
wlk75IpS2oaoio3lkmHhvPpF15zKvBlkqKr4uxaVsWOZnQhOgUdgv/HHe5oiX+Ac
xOAazpQzjZGgiz69pueNgi41yIHb83k7UxSovwMAsoVzNk7VJ8QhrlCNMKcxZwEJ
IPxRHAdHcDTIR7woDfqeY0WusC9R20wiePiqF5df92jTccBzUARzLvvg2smz0dkV
QwT/oUcWA5B3s7XeWZPQpXsGLoIM5EBNwqGvu7JyqSd13OpJlFV742Vy5NSbWS5d
qmCpH0nuWmOzrfNAY+v9ktk7MWzvxfng9hitzaeRioD+BKqK1MvFjhiwDF+dI6ie
lqFeaRBbaoGmZmx8YfyR0IJnT/sckXFzfI5hKyAcRrqXDdWScTKOlpiUuPlrO3DP
D28lAtbvulxNIYmuw2iGDnPTprENtPWaRcsjnur+Z4ob+k3G2EOfsLd7OMCg9sMF
IBHKHFhN5FdeuSTTqJfS22DezEks9VWLB63+X/11Rdk9kib4PV1sMdRRKqOO0+29
KFGB10VKgYyS7gS4CdZEJiPLbChLaurMr8H0qxC69xW2rUcqUF9uy7ySEgXZ4603
CX8yHOEgNqfPOzkc7TEfrupp5+b8drg8I1ZBAEo/N2z+1YTA1/9I2uI/LXlW6SgH
9seTbqRAWclvNgXJJqBLKZe/8FeV2m/iqQtr+b/lBIO9sSGT/JRbwvRfUMZ2m59n
Xak1983p3+Aecch4EXIR2qi0OePA37PgsWP+n2R2J+m3zQU+DIWKlFtRTjtJaMew
3EnFjR1coceDLSvAWDfBVb3lCU5FizHIq/3VZogIk1iEvP9MyVYXVJSdPGq0Fdo2
g93pJNah34C80ZRJ7XojIpfezY5wf77QhFKeqgeZpmZlGuX3cMDLsVBsIQDOgl1f
/sJ4AdOHS7TQ9dN0bFIpZ6gQDn1axlKAZru61q2TyKllqBwDPwMEFiXZWO/fOtso
vuQBXvqPC0VJtgMeFMDTJm8wByOyrkVS/6aC4zdmbWQRzCsw0T7ssqRqyWJ0PLgr
6Zu6jX4jgG6XWjCArEA52poIgGx/2jwfA1fTvSg2TmqO7OHfwM5PN295sqH7PqMy
DDoiQqHQ7OxnaiT8f12Axx26M6ToEJrvLdw4fjmf2JfEXq+YBvda4J8UbJx8vbnY
Txfnvpz8G/QlrXcYdSxZ1W9h0drDa37ZndggTCIlOI8NpMUfyIguHbayy54wD70Q
HhZmsabLXYn+0d0IVcoWxVJtQ8av3pNS4ynO+Fv7vDcaH6ToU9TuzvGvxZ3Gvj79
pTOu5kWxK7qQ9D7x8djM+ETwJLFc8qYPLQYFTSbgvUsZNPEpZSKM4IRa46ofhbCn
awlEtzM3AxfUnU1BIDgsrD5cJnGnJ2PsVhSrlDBx3170D0ENHlvNt5MKBveCaAg8
GmusfldmMnPliJYHpfkMJ4Ei2mKcxSEhswlpJRzt4lyuGw7hQf/Iu+Bh4j4+Rztw
AnL+Srz48uCX+sLvGpYEirT+eougwXQAO/yVYt9SJ/MjCUMJfZd/culNcQ+zEv46
RoBPRyucpkjfchlB4kPY0VjChpanG6lRgAY0K42Lp4XblnUpniY8Yrezeb4c0HgE
6duojr8NodwVyUv1g6bXV0LX3M3MGVbvdOWnsVuFalxEjRvqHQ36d33zdWYmNJb2
h6gtMjoXIGhhHYJEQys94mIwF87q2yBGAC1iptkkCW1cG57CCvBrtTTMXIx/Dax0
TtgFkpS0wDWh/RzpPPHqaaNs/XFQu/K/N4Kz/EYel2sR/CSjyTGwHnVsHgPb6Ss5
xdZQIZ9Synp8NhxrSaHG5ZdYctnTEXCvnNxilUgKqFZzYglt1qOrk6Llox56MH4Y
ViA9dth2GeokTXApb/QAnfx+Jvx5MK/w5IXCEsycNiKE8SAgUgZ6XxrK1GWTs109
hAvDeZB6Wq3gcR9suFpiaMH/ZaBt8qaz6V+pql5jT9nnFN2fWnQWWFW1YTgw5946
EJBrVsY7yKpJOHFdXgjfwRQSCBlPobq3TISs9Q4xlaNWQ0Y3enOhgnieHZYhwxJU
mWxQeFu2U6EnSuGDm0BWgYmdiW1HzI2eUmSEJuK2Thtx8RMdvnitsMm9qVlEW5JB
mwa0mw8xgavJcbCRafXozkYYWzdkmZ8RJEf8Hi7CBRSPOVKekttJQcovkCvN3DQF
8gUqNKXzPSydpetxg2gr7FURHKBC8Iql8kQRduNX/OM4aUIgHeagUCIQK5be41Y/
5Nq+w1NiSLqnOyCK/MecneIWToaznrvsQhLg7xt9LfcIFYe9LbCaaXsvOgoX+Df4
sDuiedW8iPiIj2qBSI8VRyvFo00l4SWS5G35trAVuMPvwD8zOgKcY/JAa/JagCea
5U5fVJFpP32vHuzPrZewK/rITBazAO23iQTMpj5K63+th6J4liFtmWtTkhN0sl36
8NME2A2jqFBV59O/dRNfsU1pDR6r8MJu/ZQ3Wnf80X2yU84U7LT9339xYyfUHaPT
+IA0gXXguaN4CUNiknY1So0/izQ6Glx3RewOSRoO8KpQr0McavgDCjCYhRdkK9MR
iUtvROdhJYIOYhcWM04RCIJ5t4G8Xwz7SE5/L5rJqQP3zlcN7vTUrR4yDwFk2rcm
k5JldZu2nFPHFeW4+7fLczW14/ypqoF3preB0EE+7Kz744h/zwLIIRRnIq4Piwhy
zRHOS8zkMLF6s3h7PTKD/tnHFu+zyRX36QspvYQRFFUuMHdEYSPbBRTbO+zD0XvI
y3Wj4s/Y4nqN59RurQrTiQDmIaGT0WgiJOfMyx/5iULTuId4WT/FSaRo7KZXA0mE
er35xKzqfNzD2yw2RWMoCQdYgwj7UHLBAFHqSz9jhM5mvjBuMztoPu4eG9+3dvAs
J/ElK6uZTWfIXX/wOR+MvzLfqfUx0H5zJuQpXDXx9aeRnz2MPYUCOfY19nKsz0zC
khAYq2SUnmnRF2M04ajs+PCFWAW6qbVs15vZOoa9hQTCK4J+T0w6zKz9o3dMDW3c
s74sFnisgfSI+MuuxtO3hyz83tqKTZ6DavQhW3iFL67HT70/X26BHuqdp2DHpUHL
y9I/Ubej+t+JQfxPvddNIHUdMja9aJ0z6kTVIarD8WFQtAaGy7ie2n3Q8TAbExBm
GbUCXjUe+nKiJLzOdrnPoN5+Hu6untx7UnxKG1ff+zBp/aNWR827hq8NxV6TjYYU
AYM5CheHDk3iYCrVm+eYT0AQY4UGHfJYDVnAVxQ3OfaLUrYHm2ArvgN2ttfuKE0L
fAX+bIEyJdKMWZEM1wAGtlFXGinPShZeFWydPTGkTyFvze9vurqmJL3pswN1w3rR
8P/9CgoQSY+3pF0YHTHa0urqOc/Ya8UMJE7TyOvDNSOli2GCEsWzQguiUMbAxDzW
slBT3E17kaAfa1Uyq/KGwzRmJHFNUwF5MYOZQZJCphY6FePyt6ODNxqmOTuP/EDL
m9V4A/Fi+FOpc5SAWQfXk2/bzUdbAk/3lWlAEemvpR1/K+x0LQCplEC3MAxZFomL
0+jG9cig8SveXXsWnHXLBH7lfilFW4t4hiMrXNzq5f0pg6g5c4emT/n5oS0vB9ce
jhd8Lmk7fS4Z8NWOg7S5bcQE+2obWbNjNrQ9dz5E7E7Y59k4lqDxXqgiu9SxbkbI
HjYzZrE7Lm9MNPLjpuMmzclNwOnfvmxp6Panh4lwAQpXXgsiwYmguB+zbbmQAvVE
j1TNXefMLiredaWuqmoGLsq1qzO9kGhslJj0rthnfJDxlH2OlJmvt0tuTR3723mm
6IJ4U0sKMdRDyiIBTJF53gbGIDkuJWTtf9q0UTUtYEZQJVS8eLn5aedsBHD3aEfp
6ALTmQ9UmhHAsvB8lWmXIRZFXXe/C5okCbSQFHsFj1DZfU+hlAaZVWVv9Hesk3bD
RmtjGHlpXCPtWebHHWuD5yIHlR/vhseuixR93T1y2Poix3MATWCuQ4uNwOQWJj7m
sz2dD65vfMAFxvN+UI1QfVphCvwVM8Uf3klFpb6NM2I/S4vXTZDOYdYAq0E/n+jv
8H7U3AsXBzRHgyYnmkWbCE74XzPy7ogeHZewkZBsoKaEuXiwi8xvvR6q63LPPGJ4
TIFOg/+MisgzVH4H1/VYE1haAALcn3aQYT/TWmAGFLzXY+tyefDluulKRJaIzint
Pe6w8KARd6RstY4lh5/g39I/iTUZD4XMFwfzx/3VYdcCBGp4cPjI4Q/1DtMtT0fw
TwoiQY2k7p9yumRmIYkLZJaXJzu3vNTgZ85Ncq+Qo1nMvDE66J8r/inS4zvHrU6D
PBFGNdBx0QG/2pK3N3Wtj1ZR1CAbQNvDSo3+1kUQm1EbJ5tWu5rmU7t5nvdsd+RO
dLV3VU252Z4LyU7OtYGpZDFnbtBH5Ev+M+I4d6o/VWcPs8Ssgq9x3KWIR/e6k9nj
c8k8BK9enn4lEBHlY/F0eQyL/yj00WG3aEKbZIlD7BBs1Jx/6S92XWcuce02QrAC
IfrPpNdPyF/whid5fIamCgwQ2ABiinmK3A82C97rVWdsajBTYaDDbguhh02m+J/t
PdDlwxxw8g5Dy5myuRE2kuwgdzxWJGR+rcsZJu0ssqHzUAKQj3XqqzxFj4++zpYk
IJ6MZlZ34leKphg23brMo4M6/DRs4TPJhDOjuphabAlFDV7PlwsTdQkK+rF9ASug
6jZ9w+6ks21oIes2y+2qrJ6OakBY3ZfykkvNUc5WurUUHYVZbJ8qmcZEoZwBejCK
zx8ekzZK7Y9ruzEW2TQpUuT5QL7ahEWbUclE9ugInbNU36inBr4RHSuG0vNQOSAP
9eua2FRIfFFKGP6uXlTBqNh47LRmlohKYKVUI6wbhq2AP5UmzX5lAqnfeqsH2GL8
96kD1czA7FkEyJz74xKTKzLed7Mju814uXtf7qSaqM1tre8yKXpDatPwSZclSk9z
FYrFMLiSSIS0CS5ZX30DTSdhUTKksN/y8S8MDrGFmfANOd/SuDTHE85a1xwaG6hT
qZv959NWpgsdFBdpahpyy52AZ9V1A5T7pF3RvNYu1f54VO0lGTT/cCi26hJcBzD0
5qp25v/Ck9qYnuySMt2u5xJAR2QXXqBEPM+/6etbgouOLfDtWF/JwAugEY6OzRAm
Y24PWoO2V8kKUJixPK4au8W1SyorAzRKilvSxrEx1NFEQtXZR+AqQ0Ip1ExMV80S
M4FMSy6kPZ/G8bVMO//7TlGEOvFb7LorDM6KkOpBycLgIUG6yA9UiDFGq7BYsxgY
dcPVugs0tLgG7f+ifFZhst6nExjNUIwzoZr52fvB54vvK0dM+5OwTfipZDvCaGty
3aijLdK1A+aXmUa+AY5U7zDHRpVQwM4ezGyeggKT/6rmhMazT2FTsSoAV0zvwNVl
01ZcDDHNzoFw6sS+zGArsYAuorThJiMYaJLtwTH9py9esX9yU/O8UgARNgaTq2y3
T3C9TIL7V5LPQi14zY365OnXHvf/ZhUn0+niLHVcnB2Akc4c5c4Wyrov4AEuZQCc
jKVo1a13Kw8f7x8RGt1n8qHP7sLL7oXWwxXXauElCAwfjTBAhFMH4rdsYYEkQMAe
TWeQYHz+IRLy1Fz9eiKKFBxhcjZ1F//84WuO9OmGifaEMftmBmDfrxGoVBwUaIkG
V+UElRmTc5qs83kKMHWntm3Dk6OOW5oiYOwCAio/YvzIuIJhLs1xY38KLDVU/KSn
pwi0TdoshcK7ZQdvOP44ryz0Mc/x14g2ffm2KK7bEaUooqXC58wXW23USOZt5c+0
QWzLPeQYwFP9JKlcvFUZ7rpjoXZUTZQrCvc8/aqa1C0DK3ebzYLZJE6VeGPtKfxD
QHSoi6q5xTSwNkiCFmV5Kvl6ZZMhSKrED4lLZIlQO4eCG45/JkKszCrKneTn9szu
BUKlRend7//DXU65/64u1u06Izu99vyD7mJmBY6qT0hy7Tmek28GIeYKampCDsPY
RqKFj5Wd1IPFldGM2i1Gx5ngt7M1di2FT2grJmH3fqnH4Z0tjz/2JuaNnNy210qg
5auDOW3cZQrAe0hEFr20QArZz8VXh6seKHp/qjvVUCw2dmppuomH9/t502/Ahvu1
BSIQMEWhz+xWrrW/TyIJe2dbl4IpuSYt4Qfnd6sWNLWmPVB/5q6hCwDtJaSWIIBD
l9B0ss4+GCkBcbMAhh3s2p5bwISXKjAo/ekO77/R9fGAuL/sBweouGEKipkAyoCJ
E6Lh6NROxmyCISPYdU3nWOsbpM9DW7zMLSeIbvIRsnulgKBdvINenRW6NZHfAAW5
OoJIKZST0JlpxffMhxa5FD9czNDRCik6wYMb/r4hnRwI4HXicnXMRrmo/CEuYTW2
3OHgAbIqjl2Z1SsBYfkM8Bm3CFDNZZMmmZVO4sHwv9fahEVSorUO+Sqvztr8iz19
ELDQ+1fqdy+/d40VZOTuiup8fk1kUUPRPdbPrBwryT10m00PH+rQgMCFYE/7Zxyn
G+cpGjsf//i6ghMm8GlIi/IlYq1etnL10VIqteL9W5aOa0QVYsuY8TlEdF0syp3y
AaGNalZYMah72rHjaovJqsrAfoaXab3gm5DbIqYlNZsv8rmYOe4ajvIhEuQmz+Za
+fDzp4AVL/EWthXlXmuKPzR4Nf3jyX+3PaRPxU7Vm8xaCKcsdypH0YxBMOih4JtC
wAan+LH3F/FrxaPAUpBHy6kDaLUTrO2se5BGzK1Xsa82uBoI7pJFiDfsIJARYHGC
FzScuuS2TT128jW7eVAKtEkOb7z/HyPQ21n/AUmJqt05rcYWl578ozAEGaX+7n5n
4gOAQS1Cx1ns1vnuZezOeoxpZo5oa/7pPZTdzUeOIV/pPobO34FNvXF1fd4jBdHh
GbK+RXnmRYu3q6UWvvED2xjBqlc+lFlUSRw/5/sAzlCdJ/TZDV349ouGjz1J7hcV
5t0pnK2/T17fmrijQZK4S2rWvToYRoEffBMevxidu1Jw40aMqQwvl9CNwht/ZqyQ
ZDL8kC2oUbGY0wzmCOEQRnhRlsc0GMR/CAOBO6ryf5YUnoId5I+LG304zP/nG40E
cwQ+jaYF+4IlcBEZdV41h0Af9pT66V6WidaWKRGAQLvdLnTdxxF5Xvt2NMuCd1Nk
2FU6Fopd1+4wFiRXnqWvz2twtc18qAdz7vcmgbtyHRSO5F6L+G4g6Ey2ctdOZFXg
5wEvVIK8ODqDWDvoMqXrAgfTYl3nAUyhWzKX1P8B4uVKa0zxWhMiZu7DKiyQgrcP
00YnNIXRjXNaxJ5QjN/xOF2H1Sxr+6d5Ulbue7pE0JovRAsqniJ1SZsavrIYD2el
A3NEzDHwhuTgeYy2UGAiGFUgZGadGiN9ROEsdPiv6GjdsDrY/Z2fZ6skWkad8/WD
3SvWQpW1isB0ICNrUhmr6nvCXfU1Vn0VGJUaRH/8dt+RHr0IEK9noDk+mbKNiJTJ
kfUEcOrB1V9BJNwW7oiCMOzDR2yzwQG1fIrfAmykuxAdhOX2sDC8ISaq3YCcgvs8
5F23n8mQNQxdgc6kEiDJnUAMqEzTZqPJeALSsvgF36SeNzcQBe8L7hEa2ZaLcNET
EY1Bqh1x4+6HnSTaPojpeE/V58FjsRGiCT/aRMhRxfOkS6cynxfK52HhJ5/pQETY
niMy5+ZRl8nOICby6jvTETeKeFKbfi5eB6/zv6WHkmXsh9k8obF5Eqv2Ib6DwowZ
Kc9pN07VJkRFBHWvbnu4X3eNid/Eu23bOvf9Flc3VkFNPj9vGDv87XJHFDgal0vi
yF1QLLVvlIAIZyqIfWyaNah8FRxacuTK74RDcPED/Ye7BeJOir4tAQKxdC/u8eIL
5DV3w+NeC/wcV7tFE7cuRk2Q0z9QQtbiTqa5GBjM/b2ImUG6fhX/s8cUrUXDtNxA
T/rJpwl7IZR/yUrIJ5QV2gJ3N+Z5ejFvcBTdoB8LlbAUI4eeQxrh7caHOBjwmsHS
c7bKtvwWM3BxRdrPwdNtz5RaOvqoxUmytlvBP1fshFR+9A930F3dKiroG9G3u2SN
MlYkgM8TZLZo4PbJKu7Qnb1XA+wRqr9xCLpuaD2kXl1giS8JWv7DEDIU0k1rYUHM
0GVXZK9+Wsx6eL0Cx+Ky12yr8hGBF5SMRqDOh47tGsvICsEIa6C18g0LIM0MDJhh
RjChnscmN+sUP7AzkFgq+pXuvX+4ijWO20VLNL6aZOolgpGjaf7PUWDISp2uLYkN
odXk+AxSu7IzZ2712sl1HNuW2id9Qll7WDyfSAu+5TGR6rpBPDhDtvh+ZIhPDYC7
SAK4aKZYUNwdd6atJPH7AzqEobkWvLgj2VI9TeuxViaJGP5AGsU5ERcxCHqvAnut
8iCQaBDI4YrQ+czyWSuhsNUZ9OeT5wQ3iybKQkcM66y/GfNmBhsuHOLX2IySCrZt
jIwQM/K6sl0/Wsknaop/ZIMwXdf59FTPVFWcDnExSCPwigJ1BA3Dk0E/PF5kB+Qt
FefUkvMnf5/vF4mu6iw2HJlcJyOXOb/DRPmFbYr3J8Dmx6IgDKA+XI6NXffK13cb
oOj5uKfDbpGHG7D+jmuhOJHJp+TNJrIZPMXU0TSHLL0IsM/eZ6Wcn7crmXqoy1jE
flQPEv8b8x1maVK2VHnVn+F1XQlmS6Zrx+hm79zd+Ch32Qa3vNy1bWJnTWWpO3e0
8EoWb0PrEfYUFKRFkPLGMTO6d+KwHoeHEjJwI2ha9N0Mst1JBhVhvZbCDpDAp7cF
7NEy4Po8mts44Rav70S8TdYyfkuG1abpgQcHFh0d6ON4P2zajI4FA1jlJEmJSkPv
27esDo2Gs3IsH3UjRqnlxrIE1x39jpeU9hfWo+mw0qfbZco+ipcsNDA6IiQxWZIZ
cEFAOJISsTd9leRGjxNInXMpBv6gWHAhk6k/qdLcCEUarSa84nF9dqyya6GdVdkF
qvtlmYypdJ2hf2C+XT9ROhL8c+7j1rei7/cI5yFnPSBFe0nyr7uz8TJeWaQIZeNS
Fk7uxiFQRAhMR0QbSJMu0PlyACqEkpCbw8hG2u6n14hslof52rrdxGjNAISI3Ity
XQ1nqY0raf2OvDR9gmL8BmuO/IXvBnvWOBNhy+dg3XTp1CiVDddFQSmd+Zam2sSZ
u7uXeOSXHk0D1IZqGGBKyrYeoi+uQBG6EjdRQhRL07k0Wh3SjYZzMaDy2XilK1/E
Mq+jPz/RNAMKtcHJGNi3WSgd5LbBgbQQ3jseaUHdKpfZHksmhOerfse4zTDfQylv
uHtBs69iLv75C8WhGZgfptdEEwx6uLZTIlswswoN7VqpRiCx93PwDFG0q07hjdgw
e74AyzdNKgEjI4EzHJBhL5QTRT8pgtwTD6w3qcA5NI8CK5lYaNXki728xD7V0Y5r
Nae4hoU7NUeMJALcr3o7pUxjHMoLvCxTUQ2AeubqvsfqSWWruQzqLpn2lf+EuFQ/
/lBuQnV467mVc/FYAMEYnqraa1K4seGIDmzfC69w1Yfui05vyCdkF0qJ61hHReJQ
YptHAbSRD0y8xPn4Tw8e2MkpD51UrM2XD6eUXzBIKSId20uu5ut0fhOEkpD30Vj1
Ga6hVTU40WMmf4k9i5NeN8veaDpbekZn02kvxzUG2XBdPT6bQYoMIsvCRVLyuUPA
4Khf288HSH1/zB+DO0z1CfOeblPJseIbxGZ6G2w/8jiG30LfjEqIRNXl2aRPb4oa
NN7FZLJ9C/poVGl51iAjG1muqKHQfgFJwMLSFOOl9Hy7vQzX3ILf6e9KnOYGGzWx
KApvWjhsGSCqnXlKA0XLozVqvwxyGabDY7NlI8e5SffmlgFdBk9uhMYRARs61Lpz
ngyVEdAzVAca0gN+GY/q9Guziewl8KAKeFahFoF7xxVXd6SExEc6M7QnwnlfjmSc
MuxNK0sW2ByFYqt3bGNmMbk6i/wyH6UBEVL8eWst13Ze2Go9izoH/zF/cusIdykB
RhT7AuQ9ztAr3/93K0WIEMm5UBEXAj8wXcOJyP7zu/7hGAjjpcYonf1I2Q46wCJI
nIV0cxEghjxrfvLwX2EgeCeRpaJ8BxZemZw546Rth91Nm9dPjrNIqDzWylZjTF2K
o/PpZaAZLGBoLWbKySdKWE7ppS/raOLFoKrPBThFRr9nZ8rQgTRZMqpjtB6iCgHC
hdmTL4T0aX3ZJxpbC6G1aR3f3AN8yT6LVX7D6LjB22VAOQEEYYki6g7TOQiiZMoJ
eAJnV8KTwfe7KjzgKuJhYCImZYWjclULDVNcGU+qzgeR82POvfVb/lBnW3uyIXcJ
XqFikxZaFKB5qzaBkOjyBuxLzawy9WgO4/81h0yJmLTmQQreyNTgLuYg4EckpRs8
5pWQpqjXN4ykwXp60EXzNENm2cNFOQCrUpp07qvUH5+Nrjn10CxrS3oKjGC98l6b
rb9qVcIMN0F7qOrMn3tVJ1iKOSP9+uleYaCmRxWn33GgX5JxIqwLOvn6Ko86gEfO
sv2EhD6sbLqLuKQZEkpRK79Ni8Po2TQs3yLW0FDVtrvXXQE8et8Idm9NW+SlhGen
4sGq/YVlZZ/2OwjgG+QOdqhASSJDKxlVSlYPo3jB6GArkeouxP3Zo5zWPeMGUY3t
iIrtfzzfNjuBSM3m7Uq85VsI12XqCUfJvkhM6KImWQxBMSg0xpNvE5JPYLOdXcSp
+/Yi9ksxGFGDpuh8JmooRNB6s6T6676PvzdTPq8xKqrHu+wTimH5N27DIopwCH0s
tsTNunwdC9QIIZBrRcprY2Y9mCr+FKyzB9tduDbxv7Hu3KrfTTPq5qu/aLX+P6i1
7jL3/rSv97sHOSWE2qMgKcYTM1SSoLX15IYCiOeX084u8slbDXPPxCR3TRCqU+wV
RcRMWZeYqWw79EZ9c07fi3Gp3nyZ5/uasDf5t+BJYA28gOqlt3iMjV1wjGrPCBLd
KvZzidw35Kio9uL4MPFuwjJZsMlXrXrPe+RX7MzVqpTGYSGH6/IJ2QFNMLIV36SB
WBjE9gxZ+95DxsjZhedV4KjrlSXLdWFmLJ2pmzswBCUCaTBHMBdKfD3QuZMmeK8d
+JGHmWDG4GBzXX3/Uo6gCm9VgZUMxqQ9Tfpj6xOEo+1615uxBxHWLJwRDM9+lIEw
8icHFtrnX3nwrCPrruWsyKC2yYVGPKgIpZjI+tDO0PDbdvhxbNQQ+AnDdq1iUAH0
VsoZJtI507DyiwiXtcVzLIx5oxOvMGDe032oBDOM4LUqEnKENRfsL2/SFFZrfwzX
1pf06rwPMqCmsh5WqmkomE2YIGIJAX0awsIlQm0aNB/lMsUCI/aGXht+/oKko2bn
LjQmMJH59n3U53xiyT9L4y9jpQWzvs6rNx1PeOTz9MbLUHBUQXJJen7OfyDu3Tfg
vopoI6rMmt89qI65mW+9Zk/yt7hkwfPUNirB1KlwL9A1fk1PZkLkdMH9a8Diqt4x
DvJ9M4tzImXY//SUPsxt2LHhlC0/YV53rQgtRtzk5+4KUUmKN7wM1E0L24yEWVhx
MZhSLTTUh+rKQFThoL6uMruYdebzcWNjAPISxLlja3/LuA1YrR5uIkppcNIcEOYg
NSEH1SQjWm0adOD2rpjm+MeUQHzJQs8sjblZqkUefclXhlhJ+SWSbeP+FVKUXH26
K8HEB8ZeQ6DSlnNXKYl0lVGJBv9wY/BFLFQoTGClU1ATrhV1oynx5MeZLm76MpNB
HwL5p7zZcZ+P9EdpiEVPeS6SuMH2DSs350d4Kxd4V4k5Y0bPK681c+WaI2Y0xh/O
T0cxoo5ds13FEbQfXbAQHa6Gr22FV2m3EufjZA/q8+4LtOlQR5f/E5sJBTjc7dsY
zBoV0JxNpxikcw30etH4wfnOg5SgvrHmpIrUMbG9/fAQUXJ3A5LzsdojGm1t95d8
q6ue8s12IJ+kVp3tX3+DO7618AbdWVrO6+QijZN3TnrwCIMUOSVpWm/NIaz77lpW
FTZJ4gDzsR22LwITNt0Xo6NBTY9BhXOzRsjSxCn9UrA78qG0wO9mPBVCwViFAnNG
Vx6PEP9nMcDUR9uyQW3up8ApYg0zdvfi85KmVvWTzlJcgbmQVNhhCagtZjxFULKL
U/9NEDMiiHa8HVDpQQyJDWsCWiFQ665cYDuUwCOCTYKdoXJTJ4PWVFWAJjR0WHvB
VllipiXBRYBQlWyoluLYPVl0z0Yy8KzZm08oDP5HhhgMzcTeB4hngOi9yNcIUxEv
ga8SvWp5X1ygi2xJnzZ/CPqLchQhJQXOGEkO/dbocrOIFQKAoGlW54AUR1bbnySp
NsbWc7xLgmb74kcRNRQ5mC/YPk5ryucVWTs5xfT9wp0qoTiis2eUriW2+K8mm7sV
gIdhex1/s8KnWo5NoJF4yxwLuBC/izz7uKDc8/8QtJZysTpd/ddY4ZQo/mEOD7X2
r6fcB3eitOFFUIin26cqMljcH3OlGO+bQ8frx/Sv8Pdkejvc7FiVI9/loEH0nHs+
dabHyq7/JS0DYj3g4MrrGdThrOKZrvEXOVcd5BmPzECwVPKAbEs9/lZPEKhz8NmB
dfoXyIJR3oYWzBFdzMuaPexl4OsPTowKxp1wT1d8zChEsJOeCEAlhlbS3ZMnHUsU
IWsQYpBQDv3g5Y/38z/FevUD0AaBLJ8ZA318TVZ/sFIOpnLHTUg1h7RxkrWvIAvp
6xVPfL0OTK8AN2T7AmDdkNo4ioKf1oXwmeey16YAHLl7OfN6RxHU/a1h4dM9p8TU
jYTNRxW9l0V8OAOjGYBOotlgkytDilXo9rCEeycY1TfvbRBTJ3MSQwwHqeiPbQhI
Avs2/SkZHkqe8g+aSLnM9LpPzaQMSCRmLBPAtPc2boRTBpe0lq9N/qUMCAMmYEk1
GepSqgaCcmNIdGtcRMZraTxeQAZNdmeyGey3eIjJQaWMEC28kcKZm4gdnLMmqe82
5geKtGxtQtPjfhx2T19kD56fgdUlxgnlLJjmoBIG4lL7rtfVCK2m1qZIMZURYtQH
Z0MwtnqD+XregzbPm0t1Q8pK9Dse/pVQ62+t1f8yN2DR+6xHvIE991OUAi/anIiW
w8Haq0Q+F27QemFSjieRerhA/YT6/qgmQ507qz0QBpTqoO7YwR0uk/NT3Q5JBdy6
TD1qQznGr1SNO2hbjnm3SdAAF2sA6C6M3c9sJ9TIJTCHx4t8VpnF//D0yBqcyiGs
gzwxtzH4Nu2yXAsuTSAYyd0VEKq7hzxsrUxfmpjK11Tf5ZP3NmE+fcHb1mUnZ0gU
wnOQsz/itLEpphfOw9XCqqKOoNQA1T8DU4xV/Fe38gKro5j6k31qMZQU/ukVYcOm
UstegfJHn9lPyGafvqX958XkAQdo6txdU5K9exy8sBp3EjlrRqlaZJoxvdZTb4to
o1U4rSKzpeO7IL0PSYj0H+rfu9IjlEO3LGz++FXdDfpzG5X/tu3/v0StTwXxRPBB
FxpRKOLCl447IZ3LKwHK5kJxN4tW8jEiSfs9DuX3MjobIXBw16JHEYVRmLz3oIJX
PXRMjMenVl6K5xcGpH96i5M7tO6lmW/0qrOrgAarxU7NqWoqzFYENnXLggYwcFjG
3+QVhhgVJiTNv8VwxGuAChsGrJPVVzFjFY2uH4LBtk9X34oBd7D/d2kTPfOX5CHG
TOjcdAKtPpRb2lElajYb4zB8YfxlNXCWiLUCX5gf+XV2c2znwqYX/SDV6UU2lpen
NZalBJb6MiRL9sqMOGubGaT/OXWzENNxIPB7lVSIIGG+qMYJDeFJhAb7urfuaAZX
okf0k4Un3bFfg+mGtAjFKypsNKcNBQgY72EFUEUGEDLkXI7WNRcMG5qWd/S2Gnuf
ezeehdSTK/JdiSb5gPUf9+XkwLM4iUM3MhCIskaP9oNF8yRGpBzg6n8lDN5kT1eF
cOPd3z2qSMmcXwy64fXA987RVvCo7ntS35Lg8s+oQ58Qx9IE/lJCJg2WZW0o5wcv
l7Dl1JOacibs5dVGMTXw/PPmWRE0GYTNHEX0Ygnq2SRzbhKmnfs5kNCpXpVnxVa2
613X4LGbQum3UHEx8jmablHxt0KYpTiT7ptt6r+Pn073B8wkycgLlG4uah7JuDPy
PycJFmqEwJr0PslX4xguMN8DxxkIV5U3QOk6hBPFX99LX8GYazzTWsGpgzMxvQfy
LqUIDFQFeAsNj8RoKHyZQYCZC3o12V9+K7ernQbQrlvBjnNLpbWSRCaDObCob35r
e75JPMeMx+PkI3IufdgjgQcgD8FRSEp3Fzv3WEhyZ0FBvfkRF6tH8vd4qq+4G6bm
D4HttmeXjGn6UoZqyfnWPH4J4jQNFEpHHlsTzq6ISOuEk5bkotyCjNkn7OG/NWOq
P+huv8pc2MNcl7InBqL2hNlA6QJ8gNUZwXSZw9m3lAXZQUOkvMdKC6Px7as+buMg
lG7x4usPG8NbWrsMt3Iv+/d/iW0M7EL2+v7vxxMpxQwS57Tbb893nJQ7a4UpR2vO
ckrebc7OU9NwAq18KCwmFkoXtKT3iQT2q36tOBvIeircKTy9AWoeAg8Bo/zDPll+
WckxjuOdFjeBHZiiIHnzlslL8wpkYSlfbJGddlM4ciaDklqlWDs5TXeuqX7ajxYa
qHdU1SHSQrTld3riknNgb1LMzahV4XZPlHdhzsoxO/uQDWRGAi8IMS4tD8SNeJ2B
ZBVMFJ7dIoN9SKgZjbOsClTggOdEL+e4PoSsJKnrb32AdEGj4BThz+F4TBv1fWWY
bEi4XnzUttF9X77SyGRJ7AVKsmBfW+wX0TENouiiHDDZhPqZVBRIEj9U05vKVf7B
13b0KdQp75LBUwdQBdZWwlYPZ/E3cnwlwAKDCSThiHpfD45GEa13Ui+EyK10dvrZ
rsOKoknhrYqY8n5jG9ilruFhov/dbD1/P8pKh9MwjE4I4+5Fdc8C9kkcyuVgpLp8
v+QI3TCxZdCl5zulVaoajljAnbXyl4CrJLeeEDgHus2JnlZdxQ22GlNfnkLdj5PJ
1LyfVaEaDAQqJIDVo7h+Jp42Xt9+O89NRwba2VARIizlARDbJ28Z3FW+yIX5Cjf2
GebBRo4/P72o7RqzWI4hzQcr7H2ZiFoR3lu+Mz0hzazlhQqaK7NR0c2ZBM0Uqj4w
eAtZOZRY6q6wqWOPxQ+Tk/29wiEjOELHKs7xb9BZbPyYvjyCNGq1gkBikZUlwihH
efZ6pWrqxHBGZQ7WBzecTdo41I4vKjfama/vOJYOpCu8fz6mISmpdrmSqzzJQf4Y
sKDJS7PFRG0xnkQHBxHbah/qMCso/Utpr+IViC4UZajBMglrxh+/vwOOQNaA6JnL
0riJ6akQKgyOvGaeHay7zGLwsCmoF9Puzq1ZbxHZuigWIyAgxbMkaiNoLNbABS3V
Nf/IK2HZeufB7I0g8YOfhJ1FCNBjwYrvz7hNWtzyCGA9IWCGGOJCSiQH1q5CD7e4
vxnCGgvWdUv+MP90t7/aIANLQWhNNzYVwpBZI2nHsWUTaHM18DCaadlc4nNZ71PT
w2IXdEW3GNjWOau7QAN2ntG32WKXZotuWYEgbw4HOP8a70g4apK22KHaUopMXKIg
pyHZLM1HPP/5tAGNCNeglKSirIDdYLuFlIrlP2nHMqQTgNa3sRToSo7YqmUvdmAA
DsYM/sxHgRdxgZ7v1M68WHE24pzkWVbVvJJBaRubdfwTKqi5wQeZMOnwwVy2xgok
OdBjVAx7A934qwSjBXCPxC46X/am5pPDmCB55HN/NWjh8e86yldrKbAKx5iPDxVo
QbcUZeEZu2sq8V2glcDjpCcUDzhvzuEev918WxZA3sdsdbuAGW9IJ8u9QgqWqDTH
d+kPQAlp2Rvw8zNVgIhgaH+Fjec0qBHa9CK6Q39uJgFCwec2K6sGirAeYIRsjNAT
cx74HS3gmgEQjMU5mBqIQ/l3nN3pmgjfqd11TwiApMiu6m7d/oafxyfm8KcmFFQR
ksEfX75HBn+KnAGuWr1UArX4AuPmMsf+8v/JQ3THMEWLaogPcJ5kKxM68OvjKEg2
nQDUnhOoRHt7tkHyy+r4fZveKtETKNK84Hrd7068ykKIwzlBrJkYJ/G/X7t8XyYk
goJaHnr9oRvgZNHtqqRqgGTfgvS7z69JiUrTFl0p8hce2BiTgUWazJSPQIQIE/6v
im3T7YM30uSeIk52mY187ilEDqCaMQnvyefdtfyeV/e3gBdRV3PFJWkOsQB8CYY+
i7WDqVmQ7asUr4OUhWF8X9OsCQElRAuolbz9Kreh68gb+RVcr9TIDX4G7xtoWcoa
rzVyzpSob1gvULHWmNVEvlPDlRPrB6hf0BrnpGKUDHlCR4rBO+TW3iwesubNIW5X
a3e9Q1colKvap1DF3t8TQHN4fmIz9+nQZCgqvGhIpL/SB0P/4FJYoyN3vo4TuOwD
DKMT71qb7d3rbW/3GC8I1H+cDj3fi/ljNNxSihfVMqEyTAI7+XTHc8xpl/0qB6LG
+XM/2hrcklxWBAJHnBndQOdHn5NgLwYmocWKtjYHVk9qrjlu3qokyywSHxbg0OD7
taoBluYBd0bv0AdRy4efKtp2f6yhgJV1bZzwxv5nA2OKAk8A389b4IJjdAVpNsY1
fQDz+evVvRlJ7k71yBi30LfC77uMzda3261CqKmtrbt4UZPMDJehnH2hvF5jI9fx
N8oAA9dlWw4YUxpD6lQZwC9agy/1H2jHVlDsv6TqlV7vChVQZEFlbJSul8ZaSKm7
y0rHAAZKjtGLO40rgFPTn2+dOGrh/j4PdzoNJbVHBc8kolArmDFNty3Uies4icKC
GL8002lndcg34lL4PN8vBer0tR8bDS5DP1oZ9wHHk692hUPBF509w65YHvYndMRX
FFAwV24B0nJEhnPMJrZYcPwAqzV3G02QZXyn+V0MdEWVuqIcxj1JjxhBrbgCxXBY
l0xO0jxB1dmNcJchg9bHbv0kkKVP8AAv9lUxL64rBDZo4MpL8/e3NicRYRnBX6Zs
8Lbju/M2OEgn4eMT9wVEk4sTlaCg5O/NeXBnwZSqf4bwk6VEeUFEHfq9BqQ1m95s
qU2VuukN5o4U3C+qDChaiW5n9EkmKuhNvZ5cWa79YhNa+YFwLr1SKO8VISnjdxi1
kLDpJxN+DLu1nlhnelCgmZRE8vWu1QkLiELbc4Aakgd0s0JXiwiq9PdzPU4UwcL8
43pHgGYm9pK35AqaSpHggr0pBpCKprTBapfe7dD6KaKF87/L1vRItqS4lkn4gUax
9MDsrbV7AgrktmNfCOBgvLyGydeTZJNq605z779e+Hp+IaH3Ou0zJ0qb0TFHoUVW
FM1+OuDIfXMt51qkSquuQ1YEDFUkpISCX/4VcBwXYhp71PxDxjS1UV7VPsLkRNeA
X7dAptEM6FXeF2c9qS9SXXZ9cUort/TwAsS+npOshXh203lpVDRnTgY4+tPj8EUN
bKDN+lW6BhpQg1VCNsMETYJQdhfJlfqBH9kZ1PoBLYgigw0Y+w5dtsGSPbKuEXqN
QnoVAC2mhXpagVCq+ef15BgxnKk3lIhdAB1whpypx3H5W0BxkR0V5gFxDYH7XkSz
EHoHGs5y+lyY/D7mqFzuuVTTXjHMjs7aqCMotN0a2PtG4ECVWP9i5UguoW03xnMw
xyeERRrVYXCAg8nST4RvDdHGay3QXhpKrhRJjMpiXiOe+hl9LvwsstpVRBhdnbUA
UGUIiZ2wjYT+fF/MJhi9JXNYbkRKXJwjeli8IsAS4nZpLQXcjvRZ0rTZjQayO9nb
ppoJsqZfOyRJpPlvNWoKy+yuA2fOMalG2jRwkcPCa65cb9riFWOJ63wP5WTDDLVs
TRONReDCfULQcXgNxQjBZlXUI2oV+WyNmSV4tb9//wVLGRAQWhQ5o7LuZ/eMi3Od
BkGYDuMIFy6H+4Y7/u2SK0cqQYBMg9s7a3sM1Yc3Amt/r0vyU4ItbifpWN8qmEz8
NqtuSIege03x18+UuwEqX03tJ19maaVjeVExDxToueHTWckDaZJomIjqatfL/6L8
tEAFEM/qB19OtRz4jvJpoOreOYjKNahcUB38ZpHlNrvXuGG7qa5TAcO+tzlfHgiC
ZR4Dz2xSvkcvl5aqqTGGWIMA+o29C0pGHcVsU61u/IJMk7wca9UAqakACj3CeZnf
We/OgNY3ts+tptXVyPZrS1yJQd8JaTdi5gZ/yptDj4+CUEMi5LrQ/xMxANHkY364
ZhOKM9HWraxZCQkiJFy49lEU5LalKUeJTYKhmp4UySRuPXtmT7QJFG0mMjnrm1dd
DWEB64BJZynjLgZKiNIIefMg1YIYDWNHUX+fGZSqDFzGVN+BVI+UXEdXn7tcGmdJ
Efp9qe0lpDZp+yOl765BqCJwnbDn9AOiBhiKRmpT2RcqFWG9wGKw3u697qUJ8coY
tLJjibeAd6ga16TUeo8Ghtkrzl49UrGJXprKqiofBqGpkt8bkJNhQx5khulzMLow
1xk1A8syTRVXN5nwdqy2CrnH3wvZWqwAkROpdVajDU8UV+0G2zcZ53kE2k0+hq8t
8tf8dm+J37Qf2SxpGKT5X2LiScdole8+XYpGhFhbHHpS1bRR6mF5GpImu04l9oUA
VFgxIo+b+w8Q3tDYsZkYoWwngwDT8EG19wg2Rb18ndMEbShH6dpfDw+qc1GPdF/v
9HONaD0KPPTj14AbgpVwA49z9plLXCFOb2s5G9h+RXSuaNFPrlSduZqFTy+Qa+HH
SlgokTnOI2dRE5024G4iGaXO0m6F/gUEq7+FjB+avHN0IYMuexaZ0olG9Y0iPB3D
PsOQU4/shQJxlXJozlWIZCU+F59G+ykGk3+C78WnwfJa2rRcQt0PUyBWI9bdNDOh
th48yv1hARonpv3Gc9jDn+LX4bymMszbzJcoB0E4UHdOgVHTBc8m/A2PISP39giz
dSxYfs2tBBIO0hHQOcmEKIHPFw4STXN3IgRQ4OIa6cFf4G6Iqj1y0VRv2DOo/B2w
s60zMVSEF2FePZJ1Kda21Rg3xjb4TGtod7HJ5CdP/Y/0F7X7EQNTifwcbZpdEQyh
Syzwg5im05mZzkcFhPCCDrqHHGFGgXDai3mVUMyuFZoV4Yguxb6XLcvZ5mro/jIQ
j3HlzIUXt9cU9CqNaTTGrF12D3YwgCgHfTQmmM4VsTPOPwxSq+b1SSrLA+lcDJay
WS5aVbUjKynWI5fEUHXD17sU4dZf3KRNyAmpbMviOmA5zA+SGmDvqUBzhFMcmRWO
MFXa7xuRXx79mTfQFQZRyj7gzRnCil0i1szSj4sKZRLTVOheD0D9J0EUWina9x15
n8ySsGCvoS3C8lBJ+8W3BSi8cGZKS3LJEQI9iGsFVOXmtoYHyjzME1R9Kq7s0kKL
crzMor//S4RzhD3EmD3kbtY5m7VOtRpyq62Q8wGGMQ0b+EA7roZr3moMTKdU5nIV
7q2rSubF/SS+N4ZYac63NgDydHtk17cXP+R/sw1k/1ty5Xnq4kWekSNN35YL89BR
5/PiThmrWaqtjefd/8t8Olpti+g5W9hEmWrWhTABHGIM05Zbj8v6c0COx1/z9dqA
kyptl6THogaEAIWuug38mHivksXHDzENPQgir4bDaXcJ8SjTZs1S15HbiJYzM5yu
3cGzzrgYDMjkW2HmjQAcEbC8nJUnYkoAaLnRFkXM1oCqe4Uts1noK0xZdQbp80mf
BKqBpFp2zAooFS+vtRKqPho9nYwGJ13f3+IFfVPIx1PpAzKGoK93DSnL+OOBpQZo
m6iC1MUFYvvr1TmWb7YVTCH4Fra1ZNIsrfRtdfkXWbStw+O1RQlzJiGklbMm5vWq
3dPawhBTkSjOdr0SK8VWyh1k76m4i2uJlF9kSsG/L0DBSHQvn3op0F0Tm/eCxj1e
s/h5jGf8rufjLT2C1xVsbC9pzHWdJw6R1igmkOCTQlgU3AfZOQWeXLZ2A6Xw81bR
me8ClYnwWvkt3I/1xka1rp8iy848OnqAtkM1vgtuwMeX68p7JAYDByH11V6d4YQh
4XiHLfguLd8rNi8bChMrIgNZnq4w3rh4x3Mj0Wp5AmGSE5CE5+4gdY2fhhpVre5N
jYaHVmG3h5/aQQqWvzQVEfpfhr6POK7Y7G8pg/ezoiusIJPQdudIjHi7TpoUA4Gp
s1lw5jktQlh6pQqvCicGP8USN9kyQO2wYvpEdXo/VT33pko/6ffog3PDy+jljkQI
YLUPN4DDaqnoCs8FToxAe5ihbyiPNL8uqMqZjlK7AUjztTwXIcexY0K2pSsZWAPx
KHoZT/GzTSv+szXpfWOmiGzRJtmHqvvbF8MNB9HrITFFpkq8k523yiVY3LI4Se68
8QN9s0BqnMoL6gn4v+c/42XdruPdmMz43ThMH+NIJ0/Zbz7Sjo2DN1Ch9DlM6ySN
T4ViQJNhdSlmuPMXnxkMiwdj8JLp3tpmax0vGiAvkvpIQHGzV2RCk2Th75S8C46a
ZCspOCKEdQohOp4jhkHe11tacMo/pC13mF7E3ey6Ownt+OCdWrKkVDU8iYvXFxSr
5NboiDwjJHbonhutJDhFi7g3PFzF9k3zv0625Ye46Q4Y7lTQ8+0kmeUk4BHx+BAb
oHG6hfaraitYplOxj48+XPZ3V80xrbz49UqyCE1XhXCOmgsdVxgrqrK5v+bu0wvX
N74i32k2zVdCUxhmEH3P672u9LyxeHdsWQpLd0EDjl88A87Btx2EHriiZAcABHUZ
rCvF5cOTb2eSa3bkgeAlffDTBnE75EZFJwCfyKC52PB8FCnZEznKvLXpwIB8enSf
EknghY32CXhevPdolseEVytywgM+qd9q3/7H43/HkJotE6zs9KTzcRjMuIkTaXuZ
KT12/j6drfCSuURcw7Ux3TvRgpXH52P+lcFKIN6M4NxW0NseN41O470Aiw4uHSff
S/D1LtvjWk5yBW6Y0cxiPg8O9sqon5etTyPHxCMShjf08Gffqm/WQvHDYx3o4Pdv
VLC8kcaN3LJztQxhIJi03wHUCup2f4NeFkBs2YWii9+JbGrFlF5ID5GBGPgXC3vR
0h9mzOD6iIeMlgq4dJeJmU1yRQjCCkuzDo2DaS0Tkd1W/svSMyNPsThkB1MDuVS7
ddKmuGuA35BTKOmgXgtz3UuVd0DZzgg/DyJ11nKgc1gYXNfcEYfpJRUCaDLYctp9
jyHOCNoHvj02u4oJ8/WMNzpClbS0CtdNiGGXjK7dSvG9rDihXnTw21gnj3NNyx1I
yhEyILm2QDrM2TzvX2cVxFmlk+dbvSM53LbPDR0WnUl76ELnwiDInSSybGJ0REeU
3aTgkNZE+/SQ/Ws984qrIaRMdWrulGmv7fFQcKHwf0VH6Iipay/ZjJYKao2PoCAg
aCehE7vJYK8PiVrzhdEoaTXBAGzmXROk1xSwLAXwX64jyEeTYp6oWQyFX99jyP2S
A4o0bzYEhRCuLIml6sx70F5Eha8sU555I1TB705TYIURf2R7cZ+FL+yfm6rmXFDx
RQK92xgUzqhFbDKK1hrOiyDr/DSSpR9D8KUMPtftsvSCVv+IWK3YxLA0UJKqQQ76
Z1yiHuU+8AQtiSAgPjjYe3yOJnnqXYPBjG4V1NEOlF1JNSFALQscy4WmLkJWdh1H
fXpV0EJbR8uci+HPMGL80qY+2v7od/WJBVuCWYvibxLxRs7LnudD2vB88HVE6Efm
sAS0OABMa+ZOlebtZ2+qW8iJ3dRs8255zxqZ9rSCKgvvEkQLDfRRPM2GMINXmadb
mN6OSmiXJQNyuZe8zL0nQcUCnefmmTE6ekarIF1ee1EUsZXBvnULXXEmTqwTxV6I
hSYfnJ/mVyZoVgmiTEW/tJPsCfdXKIn6dBfqLHQXFaFFdFxMTEcxlgX9ZduhheGb
2krzcdu9cksBFALqhs+5LiJmVRA6V/gAkewJyqeeLXykZHZTcKv05fjetSBO12Ec
Ho5zX3y7vyQR+Rs1Ag/17uVuAdijvsyaqRwOPWh7sa93GJB2aTgEwnUHgynDrsvk
/+0goiFCGHEVxpo+jywvfvSVZHWnfB5xgYEgb/twvOc7Z0+8aWN1LOwcRrgD/X65
/oBnl7ZlGpjV2cViEhpwfmJk52VbIT5MbLeuw0RXDeqaxVovx5QwPj7U/UWYkRYd
dNL71siY2uMEwzpKwwYLdxWHf7OffYd43VGjQxN3VG2SLb8bIZQRxzizty9dicen
lZLSx9A0yv03ytLLmm3tcdJ+CrmNSOv9Ok2RxNij56w9fubRdjE2Mv9D0cvaMOGT
oyhBYHJ/eT7z8g9Tq9Wpd4IXWEc42XWXrFOGH9tRLWQjxm756Q5P6DeZO+59AulL
HiFQw1C/+521lvQe1pHwSGKPhQTJtyqyBjtj5myAqYbUl9fVE9mvqIm/VCPI3d/R
mYHtCGNfpmor9IdpT0RktEuebUPSvtnkAWSx2Wo14SeHlsgaNdZnHXhROZXW4y2p
wF9OHkgtiksfNkYpmmZ1Ua1/Q8NcrEGlQ1dN1DK6m72J3FbdqkcO+cfLD9m8kulX
z3Z8ZbZHrt/CqoSjzON8swOWr2F0KJ5w+Nyf8fM5SpYe71OP4KLN4MSiHm5h4NvT
QMgY8zMXfjFVoApbwXpp/MMLsallWkzzWjLPQ+xFG1bOK4x7LhmdbtOFZ84DZK/3
EUHI576ZB0VJWVJ7eW1bw5B7czbNFQ2nOI4k5u7rXGw9zUn4tIvnr1G9CL4rsO8t
LMrJe8DujzyAvCByLfWXQYlcW2H+/1tmjwZPHM6uvDUVqU1pW3jKyPSnOOyap/eg
ANUOWyE43uhz3UlX+52qyjWRqnbn3lWOaTKUM6car5ZHWpNQYgh/Xsebuy1SH1lj
jVkjA7ldesgHnUUMtIvazp3UrmtTc9oPNtZrTTYF1u6AvHMQO7BuXHnX+cXK8TJP
ghEdNNnaNGj4ZnPlT7RfOvBumYrC1UVrjnv5SB1d2+K5MUdG7jmHX8YuNuw3dLWK
RKWu+T3b2u9w+wjJTzoJyb53g79WFWFEPYG/zN5IaAeb7JtqfAy9PhR+7RXpy/AX
W9faEh9M+AYWhlEk8rLnE7sczg8Fdg1RuUVqLnrDXfaVkc2eqA1zhEjEqHL3iZdT
Et4CTntVF3blDVmB+qxhEAZTKDvPM9YZYTyphI6yLbLUy0UU/0K8C2bIDMIXAT1k
mHFoEoUWIOXsrRy8ManzT3XYZqMA9mLHDwz94dfw6CWJYxQfHNqxrw4uLX7QU3VZ
H3kVLvqm0KAjjk24RVcc2cK/ARAi0SdEHZUuOpXvmjMIN5Kcvjod+zLi7+zUqUuQ
F1eWdzum1IZv4haTul5oOkUrdLhQnmw3uzTKXGq/n6SOpOcX9WWC+5a7Mfdc2r4U
MT7Fzr15TgKPx+Y175EIiwRvLgJ3aZph9uLCaYnRbHgGcHrcfWH2cV91VS4iStZ1
N4XQKInW6jVUplolHed+pcNHfgulJAVjSrZDkHa78HUzSgAY72BdJ/eTaaFgAmDB
e8tdouOSTYXjC+rIzp3WwxTnmVB1bIkR5R37a58l3JPAIgM3Q442n0KNyonXckzy
EFqa0EfnnBKBXOuI6t9XgtTYAJ5EP41s/8x9lRb0wCx8u+0f0UHYK4C95sZjmYnL
QB3wplacuFCXAZ8ktk0LEFn50OCdcu6KBW7CTkCxf3+wwY1/qeqJX98q738Sc/PY
ykEMROPTJJzY7+z9mY3THFwnrRFTbrokpJpwH2c82xITAc2/gmwgNyg77N0JqP/l
VWwxZ2WN7FCtFeIPAfGMHuEzA2/vl944R8QXDnn9zeAqPKRfBFBd8TKWp0RXfTh3
rZESHq8z3Vvbz/sEWY0UgbXn/XD97o8Rjp5+JsqtDZITPigWKEJ/rZqhlEGH76NV
D0lM+pjXNDGMWu3x4xopsdTnzUrkbUBcxlTYfo9TGSNgIvWGEXzUb7tYu5DgRfpt
UxIGKXFKNdWzrlcycxd26HWTXSZqaSy6tWsMUdZGletFOcM1GsrRRhv9nJYKrZzs
G5dCfTG/KjdTEQSTAvzYAYlOIl9nsG/7Bid5EqwLsMvEyzgir4Kc7XDnO2sfNG0q
rG3cbZRalV7ywZAV9Ccf3YYXdVcBBaNr4U8QiNIJk2WrUL6uvOEvBdnUnaqoNLKG
ehl3bktCNDiQCTOtV4wm44ABO2WJjHaGMxtp9mhYQuraPkAf7W4sPBWoS1t9U5do
WGBkF2JypGRJPTmdUWtImrrV2MVYFqiycVr+sMaBRJvfaNIuGFTMVtyXgDfPAmU6
nCI5AV1ztutDwgNTdZsmIh6P/BwMviBuAK7VLva9m7GJ2KYnKF3tBnlu6gcVBARx
RYKmT/TXnslTMkL4KSuLl9I8c0VDfiQWkRaKVUm6PTwxg276RHSFR34InNSWy7US
vXreqiDkjXnKBVESx7Ac2zv5uoRkdws6bk9gRB4Kbdx5typP0f8x8ObH91kOK/Ws
UzaQmi4o20w60IEYRVylv135v56ePTTSTWxyhuMUh4YmdwtFz7PKWnY9pA4XtD/F
6Xel5GkNfYj60l+mHiaOveEi5Cpk+1rG/AKs5XRqsQKR7F3oDAh4+WEZU2CSU2Fd
SsCE0j1h5ormiMpveidqHZUP0z6KYgbxyhdQrLxsDqvHhlyJLuhu5HJ9k0wE4UJ/
/Q5wGTlsUt/q6I9mqQous7WNOXjpLZuVAOwnlSdxPDqs0HKwC+c5xIx3GWxPgl5i
1dJAh9Ro9mkTpilwFHwAybpiobIay9l/3gLwy9cqKUtLlWf1LwOplNZbP9MP3nwE
ZGZIeXIQJoyC/wugp4/TCzUNlBumlER8SfHNr0EPvunW3lGm3YwynwOsdS5qfDns
ul7nsjT4nqDJYB48c6gmQP50BD82ttSUlk7HmvhQ6GNwpw3tcE7pzQv6T0+rgqm5
ifnE+vSfHikWRt/gPuPC/8+iyuB1e+iaIkdyIVIAbRlOhQS+y4a2Gp/lYSeOwGnV
FNA3buiJ5bnLVA+/1UMQhL9BUwmV5GivB+ZIcMGyAWO2eDB9WSIjPW16jgSPxA2B
mWXCkOtTceGSBsO3p9zwCFfXDQrTYtFw3oEj6GmXA71zPTqV6ntSYuXCO7dnrE80
hh1+UPOJ9Oc34T366wDPNzgyjztIhxxFuX4RqmkEh7A5qUwADGs0qbwHUdkL8yZu
o9urgwwC/7O71FIhMgNkMVaj9nVpRNsEUB3t8vF5OAwTnkHIEdGv0UCypVh/A21x
tz/g00os7ZMF1HU3rUqjy00zAckgR3uUyfDjhoRr/2WN2sAlLl2TIfzvA3mX31GE
qCDOp3E5mW5Yv951U9kA4yubs0dW2Mkt92V1ek9psd59WYPm9/gOoL3CIB1Cuxv5
PvGXKEVl5TanFAhkl5odR3OJhwY2O9myfC9LtGT7CDfFfc1ZH5qPqHrCY766n9xT
FPZJjRSiXHYuyOIDmF20oR+83fGZX+PZsz078p+GQ1a7mZQ7JuDJoHyzMhS/83n+
wa2IRD5KcphjI+MxF6xnNT6Eo7SYfFJ7dmqORAxhVOcPGoTGJUfnYY4cNPUxyT7e
y0lLCP4MbCGkgFE1kjy3YQYWld7QGDRpbzfLqnfeRBSdvWQQ0jn9+ktMZ7gi7vP2
h73aJTRzcqjCWT228CaQyUTz8oDCb0SxYxVRUia0NR8IYwTuoKUw2iuPB0QT/CDY
bfuO6C3GdBUdbBS99xKdnpLOIoxpKnpZ8B9E/kafZanOoWy/xaBfrrcU9sURvgOS
QpSXGihjwnb4r08cvKDLEwu+ghBj8L4n48vxkUr2TfDsS0GeTUhY/RS2tbI4qJtQ
nTz0MmWLkPWkCI3CdjuHUneAThoRoSixQIeTof2a47YY/kgzlgVoMYMFcRd5u3uS
z6o7Ca27MGbA9YgItDlVRVLlmxAGmEOXQXpE12eB4QGXeky1aGx9RKi8/yDPnE8l
Ra3hT1F66xx9bvufqYuhI52y81R+tpkKcyGMSKS+mJAxZwbVhriWLqeLajWte+sY
2cueX3cVCswxIjEk21JynVNmuB57mPwzXI3eOkh8OKr75Q4NtlZtvoATN0rpyBCw
QmVHzW3DwzO4g9R56hbNF4hpjdSkAqsCG9io6y2E1IZ/OpAPMA7678OAPVd5zxAM
hjgjSQGy3LynEwAXMv1pCTO5gGLw8PbzcymhODgyoDgrLNx+jSdTfAwYNqpPIrkc
RNX5HrDJxUW/O8atc9KQTu/EN727AERP2TI6HM1uNPjOO3mj5Vxus2UyQEp8KWJ4
dSWWkTbal7bDy2s43q5kQRqemWsIgReXlWFj5xb+KO8PhmlNTANlM/u5vq0cAJnG
fNzFedw6SSGvk6lcZZReHGpCKb5doVH0SbWKybO+KL8s/PTvXQca52lbPqM1vTil
ZwclsPmsSv5ZOdFM+twxdhc+wPE2B0ugW55BjpS5Qwoe/dQbkoAEGys9T8vtOzjC
ad5PymD579ZyzNWPkv9CBT0Y/BzE22kIzcqIWTIYvr0SOBNFT1C7oJeG6eJPlIOF
LjFTTFGyYz30ORqdWs10WICZAId3bCJVwNnoT61RZ2X11Z3UF8g1nLCfG8+FTJH8
9mP7nt1sCMmbY8RbEVr5QgqHDAQ5LGnoCKrDabO+Eb/Sck0SNEjuNZ/4zUzC7ugD
NZJua0b9src3NYRKGqi2WeuFOCEN5mHpJeABjTeeDQwlqEDQDFvfU3QTEWBFblI0
2AB4yrE25eM0nNELTmyqC2UA7ZHNPzHVigSloYNtRJx6bUOq7HK6jQafHi50JwMC
jbddo8mJB4EqAUb/6SFWPhBReUfxIUom12FITAVFF9r6FH3gSF3SPm6U+0fyeTf7
d4+ArlvdTJ/EOV6dnCjHPlALYjmat6ob3pTpdTNzTLue43Z5JjCkI1x2jmHmSqY/
C1qo9IgLAhgAmcm89WRracpXot7Mog7HZe3UHLIXUr8kDNX5oNxIuQ7UbRYWsb2t
Olv8lOi9y9NFvF6xUHQL6aHR6EArLX0+/DFpEM/A0iF03CNP1HJloAIVfK3xenG2
vLs91H2J+JSwq+aYqqWc9344zKIvWse/32tHxSpN8O+HS126lfx5cemYmGVDAxzP
PfErB1XL2ZBy0vqVRTPlvhF5bXr/PPEw1KyoXZ1iUtlsfV2J8YFqx8izSplSS4BF
/nWN9F8sUQEtRSkdFPURCa0PlrIatnjigyJrv2KKMMkvB6kCNQV3zH35Z35F+yCt
coNJWt1cByj/S9iFQ3ErQhc5IZ34RDFL90c9jEP8fWrtQ5xMqqZRE5UM3O2luS9u
0bN9GsJs0Y9y8DZXH5emyfArAvKP5bKi291kHM6FsdWKSCqeMRDNSvJnmulVIgZh
uy+BDeIQojHr3SDIf/qBa66ZzQjdKZ9UT0johssnLuBh+kN/sv3NxJWhjHLuI329
yfzkp3l0WJOD5nSEPZnRa/LRQd3dmI+4oGYq9u7qT4V2h30nOu0G1pthmH8gaLwr
T1MdbXiiVhVTS9j8/A5jCrJAt22QemEsJ+ujhKNq9CnW18lLoyS/oJk5YNdfKaC6
8YQSq6OeU77d2Pj51wl+NfYt8FVfwuPmx35R5OxpvT/rh9FT8qjMHcGQQZnXiTXw
+AgR3LiH1LRA9Yc46+UDa4yBZ1AYwRp8waiGuXZY65Dh7gisCL53q6O54ijiNeIv
PEk8cOvbhCneVu42Od/QjBcUoYDwEn2/cMZTHnsLw7YQmbBKOF86TtE4J3zVYojy
PfuWz0jNsxSKCLEWuaO4kFUxRQB2rra/DdNunOHo+jS0oDp5RMDlNQZVD+cw0J57
1tKze6I4IhdzFjfGnDivTxXo/CBAlQwqRZc93CpkzQDX6nXE9MSg8RXPCNXcGKhr
1CB3Py6F3eDAVkysoj0+jb3Fe3rHBgTcNBlQjYqq4deS3nUjycAqbVLWScu4a2vo
DCUgxD1iAk7g9bQ+9wTzZhrT8z4RRtOmTl20+6ZhOCemeirziWr9QyB7mrC82wE6
45bge257DKktzPdSVprCFQsAp3K4AH2/mn6uOi2rsQkp+2zYypEZX020CQWFRtq0
Varbg+yqeQ3tJj0Ny1mvcSbrJfzH5lef2OBh8u8JUH051VF2vkcsxYzkg5smlx6W
kr2DOi3GPb7M6tBZbgdFETAUboTlGvg0eLEjhIo6riQAKgVTEml2JTJmOeKIb8A4
ZQLTTG200m00ftgB77eumBd3pM8gb3SksjL7UEWElLEcBRWaC1NpCy/PGXagkqhs
jhQhkJUHFVp14nb/iWZRdhRJKoZXvaMD/3+X+jn2NI5rXyZROOCneYC5ocd8XbTR
LEkfk4E10sK2uXb9k3mlxaqEPPfZ7MQFskLihu7t2297qexKep2vdBW60npf3GmK
jTuLdUC0OyM2hCMVaQ7VumjXzSIiGpXEHvTU/LTSOEhLwxU+JxI51c2dOEnuReoY
cCNFZKvsJYvBM5F1FV4V5cwPOD6o8f36n5Ya3E+KwtA0krKuvHA6s/FG6YZCVI7H
kuIGvfnM+HQoVE/rtBbsy/zf5xnizr+XVWt4TgT9gyE65pPVZKwFZXpRfPd9hx3v
UKSjh6vgG9hKO0ie3vz+Yr8we8UusnalhMBQf4Iy+bWDqhZ1fTec5zJu/okCmqvt
p83jpaYRCMhNDwI/1cfVEmzKb0ey6Udu6dLVFHrzZLsJ7q1x2BV0HnSA3HA1DuEt
nJGO69D5ynKH/T2gEvjv+qnov6rC87r52zkJsSKmCW4FJx3KegOMHEEPxVOOtxPl
aSCAiaVH14K5h+EMbS5OkniMKEf/zgg3fRyIY55YiHJ0+aTCYRN9MMrtiHOi7tYt
6euNZDjgojAcBO02J5sHeVZCRRdZXouivIxILZnhew/QJX3D8GN5SKsrIWU5rVHr
yg8P980R/kWX2uniKEuYRNuS9QWhMIi9EoQarvKYQS+BoOuP0E8pGLD9V3WlEXoG
mugt7LsgxSZDi7Lr60C1/KxRSpkhQw+3SpLqsAHa6J2bFnNiAzEjErZTHtjPJjDT
cUE80q7B4t46RsKGzgxqwQsFLW2EhpvPx7AN2bz8qvVgY1XElvHdp4/4LLPRkZOX
OyGvbWoPIEVA38sFjQdpLWygVgaIxZyFEwAbN65Oa3OU7CZ4QbiKuW7f0MJCAUtB
f8L7ra1PFVFa36S27uq8DKsYrqB0c9GeEgPlwSloATDogoqFjRuPKsV/T+5plMWW
tirmyyNLZveTpC+52th15dvFIeaSK6L3jK84JzoUzFkJmbAtuyaEdHbtIAfxMvpG
/abV7DPAzRLhSVI4QeUvG41K3VEJzq+30pd+OgOvdCcrULTiJw2p2CkGoSrUClcF
dekJgfShrKlfiJ6ctFOSufGXTE2kE0E6Zn2JpURERhCisomVcHdHBiRPMWpFEj2B
K2lJwyxof782LHX7wiBsThmi8KlUAVYzHaZzhZkcrTzKA+AgwB9sEkO2nrZK/Yuc
h31MPogTgSotz+dgJfTvsPTiNt9BtF3JGsPjsIt6m42NF++YYt5LAh/8nuCGdICM
US4spwnqjfj5gJwxJvkIke6NdwTt35w+RoNAbN7DeE5M6AqFrnF+utH2N/QGCRLN
klzgW3gPxGhLLOnoGI9Q2GFTnQc2ZoxyBXPvqrbHY+W0wN/SkLmcE2F7H+WzOegZ
D5OTTEeiJSm8uscdUrrjmUDJweaTHV1dF6apdZwWw0NE7utUhNN0xGFkPJeYOCgN
oxuCsgSMB0o+CZsEQXFi6EvUH9BCbcwm/DEtqzIhx6LiF/jtx7zsuSC+j8N9g9lx
YZP28uLouCni4V6BCf53dvUi/RcdRKY7i9TlNVATxMOk3HmBJrFitaLtobBx2NhY
NDT0zDAx19gW+zFb8xal7oXyEEwtp3ZANU5HUC/VH9kvYMySegjRyJYhGQk0IME8
9HUsoP4oWlP9NT4jUqbAvQ52kqkTDuFmfduvp9dtWeF5VBwnQ97RVzQ50m1HBi9Q
l5/Iy+543AhwCwK+8bDESkBf+ysiTv0wUZ0EjlbRj3IlLiLs+ekmcvAo2IL0AvrR
SKMqNtmIt04gL4h48BYiC1Q32sQ0B6P2Df5PHLhTzOydkbQbZEafg95n+hPKBnKI
+ExxIR9UyZqSgj6VMPc9ZhatwaTrYpVS16CIgi0/688eEIQMBwlz73JH2WYnQ79Q
llJC/3VfUaJK3kG+7qv7px03fLpSv+/285GwaNPHXE5kWUG8RYkXq4t4KXzAwkJ7
JkfvVHqVWLv/XgFErBlnk0+FXTTsgmtrbentOVdbkHDGyBua2wIuMb9uB42ONnK9
PJRHrbGunwvXvDOonoLjVkYS1aKV06lM2RUbDbRqX7s2nU99Q6jYv5/H3n+L/VT0
tv8tOMlZCpxPEH3TbyvJDLRdGcwBUxhTq5F68JbD/BbgP6pqMA5AMHFeaFw2kNmp
mRtwSnR1/AYChdYRlvS4640ofNzHdPM+1CD2BsH+Ug4P49ZIuxuQx137Yj2FYpnk
G8Cwu/u1znBjrYEAKh+UgRZkxrOefu2q2Gye6EZNnngyO4iMsdjgq3V+oFg/oeLm
sFNQjwdPF7sdUIOAzMVqDKsAGnVV8iXEMOQCBIvDLiH7n/wNvP5luG5qkPqciv3u
3XusWcQAF9I1IvNsAvxqEmRhcUILeyjgSFUkOhBeeNJPNE8uX4dYBW0USoLAbPVC
TGJKl8nZfK/UsBLr+ddwnXV4yvKnt8paOh9Sitcurjq/8upnSzC66dj2kROmQmwY
FSIWSXZwmAo795P1NnF/f0ce1t1NEpvfvsGquDkRk26N9RNQtv+Dtrl4sb8QRDRS
kFMt9XMJYykJTjTVq/8FicEcX4fwJeocC/bfgOJqB2ID/+01pvKVNzLeevasmOhk
CSh7PYApZQ6jnEDDMfEYRcu+tS99rIn7WdX74btQI+kL5k1XYuBdsfmR97ejfbP4
C6aARq17yeNN148pd4z28VQG/A1oFlJbW2mrodzP2+MmClbvOgysHnihMGXJaNvQ
N0VIWN6zNjb3kFRN+W0wefghoF2d5Bi7Tk3uSPCDKAGUKt8SeugEj76cjvgMlxbf
8lyN2kjPrHPJM+Q3O1q+dGvscbNeJ0EoNKyCVx0hzJKqJofDpMa78HolIsoePLPx
ozDGBBdTbGvRb0b0ckVUXCsGStLXLa0w0JLEHtds6w/FL6cgcLu4VBVg80ynGMOK
QcGKdaiv4MGhK9U/yjaAr0RJTLw//gAeOup0yJurVZg16i+QIeVXBChQCoEmsM1b
0JHLmHNalP7TNJAEvTWYV8zTV7I6qOkoqtf9Auj6J+e1qyrJ7W4oGJ/SnW6y8/Qy
wGp67d6yrLLADiNYp6RRLCgQ4E3SPnapuBeF4GavDzt5lFTN59A6HEXwZtnlWGrw
DqWowo+EkPm8+fhpW4XH1AKdf109V6P4JpqlT4K1hok1ObTbiuCYKSkWnayZ0rFJ
zmgd3Hb5nCIaoJE3clHBQQySbDEqOiAUGwT0F3TP9ZQmVSrhUuSVfvKdq+7GWW3Q
jJcA0/+DuMj9Huf9N0b0XeLUEeu4fo8I272pc4cupZg/Wmx4kL98D9ojT04pVODn
jYavFsV63kzpQHv0DfkZCiZGBUzWRI8VR0X8Ka8OSrOKLsRFKPO4WLNr5m6lsCn7
kPbcQ3jQfMKjHD/CM3yTCF+u2iHItVpSy9PzFRG7G942LDXGuQHJjvstxMBnVT+A
dEO/1jOLYNKfUQj8Wqo7nHBUHwy5HuNvZY+MCfTXltQmM25ywKszvxfo/eT7dW1e
cbKBHunRRezUTD2jp1lYdDDa3bdCQfyEmHMgPYyvWxpsU13MkC7H+dzoXQdN+LZ4
YFo/kjuqNs8Bli4+LqsBzHeQQtp+89kDR7rro3RJbcwseEsuBATjFGe/kt082jAa
Pd9oLVFFKhBCaGFC81DjMVDn9T4RMX8cO+kQU1EYRIkqBdXJYa3925s927P6aBF7
BvUvY4nUUWthzcJWymwTvRgz0KtMF7D2aSl0E5XwEuTZrxRwqH1tsXcVQDzqSCnE
sYyqAgnrS/vBy1tkz5EqE7YaDP6y9Id+Dk0kou0e1/3gegpfERXJ4zSVbY10PHOZ
HeCdF6OVDhm0Q6HkgcmP5gkv87K7lXYyxcXF94rnaoDY6/kPvdhrVtBeJa5SfVNi
gCv9YbK6xrS70mwjnLOYpIcNE5P4JIC25cW1TPComea0ERcXlX6oYukkHCSG2SF3
XZ5OaGxUwxM4DQhN9MXNx6eismErPw9ogswTOFK7W1g5LR52IFvSsKFUxs6dfAnw
n0kjWw6jpFj+vS1LAqWTPgWD0ZFavT3SkzC9h6Y/N9Dzpt6J3p1BXpgvnacRcSJ2
D9TXtdNp+CfsKASEIzJ4XTRB/cSNeX6tSODjyZ/xueI+YoAN/27rx+D9bHlidnQn
VLJ+2g0vZSBAVOs3FQHfYVNQUI/3uYzvgcj3zBKwPBywP7v5IbqqeE4eekPMjbDQ
fH1PQFKLpn6raz/yXd7MJpGVZkwny9syhWp7MmSazAVknYpxHm6kPkqrspjTtL/G
uwZ68zZT6rXYhFgeTzBsLhaSr9TmaFdqdZuGRIwt18C0NAcsekSO4NTz6vy6fToF
qAxrT4MNedE+S8mrvjh/RcRTIglbVol3mOFr/LgOJHkHf86caQ36i0pKYJblhHOC
VsIh2yySkeGDkvPcL/2jTTS7np+LQJqnWTQXBlvogs7MKPlmPG8QWDwRll+x+qHR
Paehl1bOZzaMLdI/pY0TkkIyjLbqYKe0N9oANEAgkzQos3fzF524nc58r1pZIi3/
zWLBUeE1jxhZbBbe7kGEOD4Te91Jrf2qYtkkyINAH3dHEvlbr2qeygXRZu5EtMS2
qXqy63JzckEo1YnRszNfpExfPSrBH3sdCkpnmntOIsasGNezvSKlrp9y/stA4t6t
py6QojpQXA9BgE02KOKq6V+TN371seUjYJCaQoym6KKDheb+4tzq0xOdn05ifWRX
knC+VjiBwHzBVxrhVrwlZmt4a59sRJ17g1drBKBcvSL6e3nutxrVYNPpVNkwi85Y
y6JUhAr3udeSF8xvD+OvK7LHuJywz0rKuFAzcAXFAjPiovVNpl6iAENeIMo/mEpg
jIZxBJlZ8Mtr3x9f3M30ax6N1JO04PNrlWCTXwCnnBe813g2d8PPqjg4C0zqBfS0
Orw8tosGYjKgMfj9KnddUwhJAhtgCxbUmkXVgeDslUSjpW/XmdgY0UtC1qWHeD8z
YCvnvVo6002udL56xvZGDohy3eJGzSg9Wlq1SXhKZVEeDBIGrpWISuB8corVtc4M
ddMDKqPbEgmYeBDN9iznEBNTwXKYPyVEgtrsiXqeOHVwRa49RPc9JGMYuPd48gex
CFWqoApWgBfLJBx54rS/GskOxN/BFVVx9Oq9ERMOnf+UtSyWvQ+r8nTqEz8HFHMi
GEQvzPMh+AJZbyo7hjYoiryooeZs0uILu73nUCYQVL06jy1YZ4NL6sgaMue77JG9
DB6ONAfS7EBJGqlN+63quIVV53FSeVzzynCmLFX6qdJ0mHUp0GJIDTy64K4I3F9t
agLqIwkhPxbsv6X3XTPAanwjXpi8RxrZ7nD/YMId+9ZnOuCqvXS/SUP36TXVUkm0
jo9bz9LlxQ6ZE34pVu6TcDMO7WLq9ZyzT1Mpu1iqPwhTIYEeIx7Ma3JELr1Yfuxl
i9MW8zuZ0plIhoIpjpj3EbsdEygAKTi+mwJT77fPTyjuhwXUhMe95DArQ2Oj9AWA
QCfjTJ9USsjgU+7Wu6ErmUVCS1pxNX7s+d1hVpV/AU/2tKLVNybU1xUXzCscH/Cl
sGUHb4tTVZjg0f7zS+LV27Ki2sv10H27cL226EFr2yUu8M7lSv9RwS7ERf627Fef
IzKmSigusjRI2IoZfogSX8jM7mxHIPx3ZOK80xlS2YXecJUFZxtC9JG/tHPfgV6T
WGqXly3YOBDcSHFQKloN+GY4u59AnIPA+VLJojZFH6frqtqQrCVMXLjAfQi7vEnm
5QvubcccpxdtVU4rN9aFP9xKL1HKQDVhz8bzpYMX3YZsc+LAZWgITdMiMo1I+AaG
HPVjTCCO6wvxw9nr1vdkQ5c2QmRHQbQe8dV84eo0wxsnSdDazv05XHqpAVs6Spfs
sbIiIJwWGFnp1qzWIXaA2wgMsjIIIGm3u/OgwwNmDo5HtDjAK5yKxDmO91AHRlSq
cCq21mckpvZxfmlbt6gFGWTPfyYpJlPJLVYnC52/uey3niTSRWWxNvg8nIaCdaSp
wA5GgOt79kUeayk2jox4HMRPwpcVPTSYzlfPF2ZYXEN55SdZ+y9zkS9bdrfgmHiq
Yujwtkalv0aQDnfLLGBeRlT8G8DhZgG+DpbUys3s0nJPc7MboPQMO9s7+dZe1OYn
XKT94sFTHV4YYxYiNuQ/kEE97A7/3JcJqNrSd9DDYw5vYB1dhG0bAtDNKlSfgfbs
PGvGiidAYAWk3vmnBYuHAZZJeSQxtxXgzVp8m14ri3QojKcQnlFn9DBkk85emEme
NWSqmPivpE5wBBAi6jXOnjRErmldIMcFmQ9GJhOx7SItTckUHdJSS5Ed1FLImjUb
rpreuQSw8yv94EwMQPyXIB5bVx19ZiHOb7TlFzBGjUPm5ldq12KEEqWHC0hlw9Re
H97ZwImwMts3keJVEpZi4JmdDioSpTkBK2EePkniHSK+vPiDkXrovMvGhKs75Zee
GFl3sq6ZJdByjwqSSXZ1FogMmxGyHEvLERbVgv/oVszkkHBDHQ7gdfHKc38H4jC9
8r3GVbgSQHHzF/6V+SqdJcT4oW5hYFPOEqhm/36gz4OuoKndOy0s9NZsoBRET1Uw
Zuhy5238l5zafZsutjfJgN4sWF581W70AVWIoS77SmriqZEtDY7AXaofC0mi3fkO
fmkJ5ZhBl4EmZov5u6bwwjGL3gAnlyCXUKZ7iiqErPdtHXgBp5jUbLSFa7Jgs0es
6ifx0vrHoIrb4gigG62plH+U1P4JdGh4WPaeoWF3nScETTgeyeMc8b4e6pUdUb/H
9b6021VRkkMbDTwP1wBkzLjmyfdhgMuBpNj+ytLR2P4SDMBilreiUJM+O2A2+9Iu
nKGc8vHtEqLtTRIl09UgfV56RPLSXkFLTjI1GwofaLFaJO1fJ6y8Cw7Jq/u3FJhp
Ud94R8BFqSuXmGmTMwgjngupnj7A5Fvd0NviyAdyjtC/FNHdiZlfRIKMY6J3uMHA
W2+VWom0YJOpJNPg8DwtW0Dtl3HjSmvy/etpegK5wLQiUCbFz+y1nUPPwyAiteHh
EC0Lp0NIF7gYVaRl5lGYcVziiqskkniEmc5QLM2q+DXCjLQs4wrT19tGTp0wGYBa
wWRmcdROBIbl4lcPzPekW3CI2hbXsp8M1Og98qpmn2aBIqGbaCXZhxRwQA+zu5tm
qy1jczeG4vQKj4eICo1msuU01tdx5o9ACY4/oesV4ICNM9hFfUPZI46UUMj2j6Xg
/hFLwJBTAyxWmJdCDWvQhe0IwEsXMumLIRdpjWeK7pqbTv1gzV14fGnNLURT7Hbj
Juw7QSsf2/Up8vJt4Y/l8QyCH1elBKwx6X9Cwf5W0FgSBrgvaOZTgGpFVHr2h6IY
9jkGPljYSocExlg86xx3TOgjBB/8lhUJSD9/wwwX0Oie4NyvOcEneHVOF0SI8Sto
xWXp0llCHLPMxTxXAkYRKO54fiPUx8dNvLrXcclip1PnVFiqFbcgHNolTCIlc6dq
sYjHdcGASmocI+jjez99+yW0+k/eyn+F93j+7R2RwkuiMt8VvpHPyBtwPPjkscUg
0fo4RqO84XBpfpjPtyKGg9+gQ7D2sXYMWRtw/2Jja0ougALBJ9vFC1KGUIj1vm6L
cSaJcwEvcytQEiDPnI7u4d+Ij/d3CdguvoEb7wWEw5xRztUsfCCn2A1q7qeKah9Y
IhtGW5HeqvP+QinkFjoleItHLzScWV2nnPs9aoHPwwNtIk4xfhp+EHe29etyBRYd
9Y4N0S+ZDXGkX0sly6QPo/dAAE+gRyFukVXrk2X7UQEWRLRDMuwMYem4+ftIkzh6
LqjKpry+ssPKGq0FrYi/LJxZ4EPfX9XlBOqA6AlTbB80rdD4EtB76X0ECRosPzaX
dGXtl4GAKciWHmH9f0dXBtCwSnXga9gglO6lqIPxaVuUrSWrWoDhJi9RzgSrk/fv
YDTAzVP8EiMODYpmUjZcaLG8YTaSMEaal5Y4NQ5yudKGrTpxfDST+8vSQ6iP6jdI
6BzGO1jq033F0v9QfUZp7UuCiC2Rwf9VuyCxJJvZ5Pxj6hrGQKs2ict32jrLu4Kk
w9T4rrTRqUruYEGmRPt0lTJi7uh90eUOu2VYUS9EkLA6KTtVIIsP3xTT6znvhv5U
6wCICCu5le9CLwDXhM2sCTPDDLEaMIXIJtoeip/A52FuJQvuLFgCkaQEYTBV0nat
VIjs+mmIbbemrc/Vd6WNk5RivzrHZe2GXi0IfPyCC0XM8SxHpjKQrY/KoK0SBTXG
YEviMfbP6vK0gqng8udyfJMbiiuJJb6Os8067NIy8+PbOsu9VWUxO3PG/zEJNWGZ
QD7aMArVm1KO6g86xC8XcF1qe7yg+G5lcVCTRlvPPugl9QJfMWviIi77UUeWHi6t
+L8M3qtIMlQZuUaOp4qxZRRnNirmOwjDvB4vemvCX44uXW7YHj9CDBzQUeH/VMIo
S0fepARrmFsxhMHxo7yu0eStjYCg1cKQoJLDPoQiwYejkgEF9/X9cE8fe3oPu9nL
jdpdhvA2AmP/qRTyHubgc5pwKfK7WCyV8AYTA4ruXpKycO+fYB0QII1oF4MSUbq7
8LPSCEcMcC+yL4DI/5yxiYos2yajtL8jwKvl6p+xkEsYe8dETqHTH/Nv8R/rdAP+
3IG/op2A/nduEGwZknme46bT54woZ3sn3pzFWyRaI7HL4crQzTrcM5yAcOt1OUDr
aXJz6+ZXHRNB5bpTc1CdhZkvPfJmxKKg1XxLqY+2YH2QK2PfrVh1v0saRRtZJuaJ
f/N1Qf0iJ2ZHgTmC5mruOOuvKzELHOKPQz6mJ8mvigLpwXUIgVpyvz3ai5IcTa4Z
jjAVhzjDZ3v0TqrWLgm5D4Hbo9MiIM4ejJl+Oat1i8g4FIHG1/9qPmzMLZ6bqpMR
d6mwgCu7a05h+YBv9ynWNiF5kofVBRvgU4ZzoizPEZGWHACa6X4ftE+8nJBUmX4i
EbX6eviTexVpdvvAOP2Z+LhznOLHwQn6o1fRW7yN2l19X2WbB2txNRlpq/4m5L7L
eM8xn1tUccHcRiHAtZ1XHC0dUq3gVY3inFHnzDS5yP1i0FKSCcxXPNng3qxoSuP2
7iU7wgWwhvbW3VEuryhaYutzR+OnrnbaTY0vI8gqoqZwk1Rnu7cpRiYHrzoo/yJH
S4I8tbeQiXM+npfrXjWfIcFFlN/jDterJGmui9WH4g+7w2URxNFzdqlyJpZW80o0
juuMLWwYf9BsLpq7Bv4xh3gYjKM5U/xLXIXwA1FwhjIh9Dehn8UopqOAGVk06Fhr
w/44VWVEbr6WF5c4OkYK6b5jGeO8orzVy7cvsW3g7vd1ytSuaShi3hWmuRjaKnq2
xU3/HAUlHeWt+tidXsal884CyEGk7OWEKe0DUTjppuJ0sJB97O/uMNH00dIDuy+2
I19+UzvSG5SwEo8SYfyawB/Ll/+pFcFOtpHQMneyJYbpT8jeWOHWH8Pfwan15aq0
G0pJ+VSHm66IHFNA8jkXqRnHxFmOZxdLMcaHohF+SbwZIGkoWfQXsLOjuMfvfdd/
pE5AJ99TnzcgmUH5/mU80Yxm58QfPtStoTmduz1QTur/v4CIq4OTmnSJ5EaxSbse
2dVTBIEMzB315568BBk9xaY5uusD+a3nvsQzeoNT+V5XwbquCHTrf11W6Pj1rM4I
EYMpxZFesHRRVz+EXyIsmWmn7EHi4ywY8SCKTi1zfqJdf5rn1BxyWKkxuMKWZbpG
VG0vshlnEILaX2HiwEairQEAfxqASMr60F14figA8curlzAh3DefqUymjgDuWWw3
NyT0iyWFn4UAE6WSWEVw2mkbnbjcvAl88oKpjVJC+yM6JdvbgxPl54FbU4+DPbeA
LSaIIrkqvl09/jPyIToRDR6McC32xh3/XdB9w9/Jrn+Ewx7BvtkDYt7OZnbZKp+M
ty6qd33AeELzMpYyt4TajRlhkElxIHaaMK+dXgtR8YQj/7k3JoIkALMWUCkI4Vf3
esATCo7Gm/Gvyuu+RL1KjTvJa+vCGunz4iLXpB6UQ1LE3dq/1DDlfr1/L1SOOJjt
KlcHJ5STltOyvgmzDr55lmCmA41gKTc9yGIBu9Et50XF1v8dY5ajIFRfXd9UldOu
oWsvfHGVUqqTZrLUZvVkzfor9Q4TfP76NdT0HhYzateIXPkggOrveQAWQAtMIlnj
QftAGmVsEri0vD7b/vw8fBX09A1B35E0IHFQ6gyiM9/oQ9MmeAqer5GHPRMfwgDt
P5F+vbw7bP3u2iB2nJlBkqoE7Bp8al/Wid3+bH081FMlDOrOTQ7CMnB9b7ZD2OgC
zJCxwX+jLMb1F+OxWDG/EJCUdHrPal0aN5MW0eGTbUz/DI5W6nEpLxSkeHF9vxYW
hAxlYy47T0zhwQjyi0bfYIgeyKdJDC0eo/l/rHHLps4BqeTPB0aeMq8015BKFJcX
eVkFS9fIjxW8vYsHcvE1veRs+CFB0KnO/tiWl9naFkTcq0dzacxbgv4vjBiPMUFp
yMfFBv0aYylF+4cFZLEa5c0RA/VYWH3SL+yiq2VkUKbFjSHy3o53kzc+Ai562Um9
jIQcSpc3gOLUOkNv8P14HId+dwOLI4+/ub4kFvcu7OrjytMtMadFULKisCnj74Rr
S6IjGGbJQoXj5nr5xTgTC7l2JbQF071Ps/VozVLyi1/kaRqoS5JgLwN7X1CGHFI9
gQ3iEDhWq7Z3/M+hs4hQyaPQdB+leX4b2gNwuij+4O/tKfx+25HK+vTzcHCY7756
Pq0BqYaqXf48hGdyAPRrsEpT12O6vf6NfM5zHmp68mDR47iJbrQdH4iepoMz5Pvd
5iinlHSj97adh7taAkVDE9tFFKVwPRzdVzZd71fUE3tictctjzmM85fdMwIGDcF9
IFGfN8xKK3sSuzSvHhE7ORtQq2q4tg07FV0IN1Q7mLODVu44DtX2NQxJ3ZdZIdjL
jrKqj+gGks4WacljotoMc9aiY740GJ1r6NPoPYW6sIEhmeUrKo/bqvWN4vIMnHjp
pOQUeYyIaQIDOyWj/jDnJXiA4Ts5AqKl07Vez2LgFhU7prV2sPJ6WXJVdMBnsxn/
oHoFgHT5KS5Df9gMRInXI9UIsKAUux5hRySg+IvsrlNfrP0ARG0OcvEoJvMiI1jE
qpMefudd6AmteF3xeZExek9xF62Iw2lJy3Qsb+tXdTJISkhTfBS7zRJ64zdpJrO/
rwOsAIAGNEXzTtBwxYgQ2X7pObfT7aaPNkcL6zraTU9UMSjGlQzx1Wp4IaHRg9dX
RD+gwPvHifdlLoz4n7BtaML64OxcJ7olcrR1NxiEN6GYCqCAtSkJPXviCAt61Bfb
BsNFY4umR6O23FUgVLHdGHZrt+m3R68XjocIk6677yKB5j8Gcjsu6fQq8BkSB5BH
7WQ33/ECNyoEA5LbcbTIf/Qe4qzTB220h+YZugaQsIjip4U0vq36of9OK7BV0Ye5
dvX28fBt1AHKzhvizZbBBpTXt86Hy6yMnu7fnX5cwOYQ7TGDi8bb/yAAnr3g65eK
DSRhIo7BWHV34FQF6msPYPPogqgbsKiwgcpYQS8A65JPMUNkgB/foqyjgRSvEjds
dlAXWS3YxrZPj1M7bxXRqZS9Yl122hWngKlty0RxJvcIH2VTUFU1hF1ZpNzyn8LX
G2wszlpRh/CXS4fV7Eq5gGHmyJNLJNlBVbl4zf2fFJ3j+0R+audIvKtr+K2yqcnb
ht1j7+QZHjDG5IJ7R0aP5wXDmIUWd/5WiwgttjpgkdP19Cy/zKr3ny6S/T2uvuyl
D4qPbnZyMt2RCO/EA9krRD7lf54smkufFapqGHQKU/NHgWGTPS0Lg/8lY8KA3T6A
J7Xm03n95ecPis1UwWXlF83YEIN53I7SjDWW2pP3TvUjIE5Fsm0S1OFSJLy0iR6y
7FHEbHSdYaVlQRp4CAYHYdxHQAVulbnDONxkZY/miMCqBKaHdFFP+0W3KAh1goUl
5Cp0dlQbVS4p+q4ImBazOrR3B1emOTK8mwha3FqGKTifgSbcWobIvFQFDh1KcV4T
kBJS/VAIJcxuu3RB88+2Q4F4oz0stj9zMmECSyreNoY6RnaAkboJM9z3aUe0QIRW
95HWBS0PTadOZ5NK0QMTXdfNhkcUu0u04diRk1/K40sHtF3lIDI2xBbt9P6yCtEs
y1R/Ap96rPs56MH21Xq/RydyXN8e8/kxBK+LGvDugHuLPspE2X0iL836Ir1uN+0q
EzaXus5aObCjh70WVfMEZd8KeLI2sgV0f3/PvSS8L+imHWgP3XnmaweTuq7nXbzb
rvJbva2ZGZ7LyDhrMeKDzqS7jPNIhqmABNk1oLszeVCnObcwBekTMuhpzFz1lBzF
5zLwQSDvJ98VkdGnOQQ7nTQFc2mrX1KSiOmcuC1Dlw+XpChwbcrmtpKHPvi8eXHB
dS5NCZGiYHapH7lLLhws1ip/iWb7VejepJYVEpLBql5gFsJoELZeidBp6T/PrHJ5
4OZHbWxQa3CixHz/utWDlub4KC2jDQfYgDoQylmDnLt02ir6RjyiCv4a7dea8zjd
RwSxqCa/qTar25nccYMisJNVo8+J7HHXp28dre5g9DutWU8b543pMf5q498OWRDJ
qGclxqxCTypAhciP4UO7xAcPJcobD6WH7363p6rENN1f3BBAfk9AVIXMQ0PsAmyq
GiCwugeR16/bsPKx5z6I6nqa3oMfy++g3JV0ns9XxmhTWJBqoiZDpkGwoxqztzu8
DhqYJnBqT4Ruenaq+imOxo3MB0Cropy/OP9rSe3mgbm5UZnxQ7Hi6qtWWDd77I5u
7Nmg0L4ZzJaY+dudbeEbahwzzx+FYwPH4Me5csiyOMhR6gWca95cikbqyvjRwePS
zA09sp3zLRTz0eBIhbRMLkLGQmiPn2VQXHOzmNrValeW3dMzLyXGVtlaLvJC2rRX
Ii+XX6VeSyHnMffRDPlIibbXTjp+M+XUHCe2l+ch9oZLFX5vuyN3lMTnMOcahEG0
zTpvKz9qlZ7rgfP3xPS5CufDc6YtxH4QgP3CMabvnYbOeWYr/xGiRBKzKPI1xf6d
slK99w3vrpe9rGf+T0wQV0hFu+Q5IIdzFNsLeZ1WrycnWnCxlveWeSbiLsw3c5rH
htlrnAj9SWeXE6/kWfOVCDu9XkPl4t+7iOuUOMbRmCGzR/z5IgtPuz8KDnfxERKu
9LW6cyNgOBFneTj2WO88/3k+WqxkMTEWhoccMVcIdvLZMFWgb9XX8eXc2l+9Ppzf
NYWkpKYhAMl00nBn18WEyceHF8FkFGDCbID/F0c5NqcRNOsAJDzLDw7JczZZb8t1
rBY2uAh19L6PSrR62CpThg6OlnseUSxXLWclXjq490ZiREdgUnh7Ip6V3xRnJUSs
fNF02ar+X+UbeH6JskCXHLCTsyuxYRuxUHFs1NetqZyuLdpojNGr62/XClz/Cxvo
cNyV+U6UFH8mmvhhZDUtWQyu0zIU99NOvmr1zhYMlKdHmbze4or1hn96k5WHNGTn
jHlBSARzhcA5ux0p4+28sW0Iq7zLaw6K8DysmKWoypWtS1D8WrvEEKdsfWJWFVH8
oBtOD3VVF1AsG+fNEcAqJwSER4AtN1/DQzDTLWuP2HbAVHk5OBy97Ljx41bTmaCS
OOI0Bk2eAxCWDQgdELR9S0odoYkFXeX7E4cwBDyXp5c2RGEWYA2mex4VVM5N/4Bq
j5JttyxRYs/QxZ53W3ShWqueXKjcu3VCdVeFM5LvBTtJij5IWd7/kE+h16n1BaMG
PqWOoJK7Vnry78cI/PVD9uJodqL85svlV3xfynKzIclP5oQSmpkMujAqlIPfIg9X
r4JnKSuKCW6LorDmL0JKYaauaCXhLnnMB1giMDa3KtNuXcY21pWD1gZgfXHck5vT
4i8mnIykh3TcYX9HJmHs2YThwi2zfSVgzUPMc9u2JjKi75GaU+dRmBRv6ITboThR
VR2JEcFwvHmvn2BV1au55d1GR1gBHCB6lkCcf71Rw6Izqd0MKbbp7E4SWo5pJk4W
tsnT7SxceEWCFVRrRPh0aiTcEY5I8whdv7LYWybdBXXv66m/HNMwb8PjmmT6Z3Md
tZEY2coDAlEyja0xYAulDvc9TCND99koK0nLHb8Z2+7LwCBiuCuuhhDlcIGyJYqM
sgV3b3OMPqDVCSd21rFa6WTt4QBpRTBYEAe6/kM0bMiD0Qng05EAC/PdL2CFFpRP
XVVDDqVWN0iZULt61JnRvmVG9pqo0ssQ3uxGr/2tOTQx6gMrcQYAjEsoU77rgY4x
C69wR4a0yHMkks5Wi5/55CSsVL1wRDZ0fmUAPlrN982zsEgR3pveH3eLNLmvj7cG
v8Pm6zIarX6KGVC1hwVQeF1CYOVMbbX7Qehw3XrRGlQQL5XC4weOQyRzjjXfe47U
KW1e0trr0wRKW0nJyvPKKnsPjGuw+ao6WvIhHUUQ6iUxJFKGFc2hVsRxK2Tsv1Cr
92C2MMCiMBQMeHQpaVLwA/vJ9nh/kSVsLczi25Ld/YI2Npa2ScWCbT+tBQX6ZMp1
b+rQZuYa/TRbyTmdldZZzTdegiVHCM8qTa/mxN86CVRk/UbMJ2qmtgqcmisLMGWi
brejuOSuikjrajtiMJ8nM6JnUfdAHjiqNZAecO2yXeaEcYN4DoneBdlXVf3SQhoJ
LmtEA3NL2MUtZxFGaIKw5c6AshwxXkVRF/oCaM1SjEnuLGt76QmKjauN9EDuePe6
fU4sg6HkOCW9fbkrEP3dbWmXWmaxy40orPDmqEcmAv7s9jsU555Q97j2OFqNG+03
Ddzc8+16wzvDiNt0X+5udU1awgb1WoNJPgg29adeONjcFILqSjkq9K2iRy619YO/
t29upmIzKwuO/sv1c8WUjSlIz/GOB6lDq5Pwq5Rhr/kZUbCJoHhqDkb29Zgs2RIl
HevL2cVzN7JrCPqFI3a4EOef1BfQnt6TUvmLiGW8eimy0WsbR7DQ0wgXwOAzzmS1
JN1n1AT/lBHTMq3y/QygmX8KHtlRRXSBg7qAHKZKU5eB65Qb5d+VxUIKJGaoFdT4
m6fhtr6j3KDrREF6YV+XurtaGW8sGn1VpCQT/cNmVQdgVBo1GmaWx+t34TMMXwwm
SzkIhU7FtshGjHKF8XjIDGD/jo0HEKLygxayStvr2hV40usnROAAjJHUm4yDPNcn
Bh5bqKHGCmUMcBejXrWJGpB1Ip1x8es3wI8AiMwPEDW/gRqnqDfY3szuel8Kl1t4
3++JatzeZE4CG80q24oXNI1v1dFwS4c0XFJY+tNEubX0RrYlvICrmz00ySsQtxi3
jKkHJF/U76pO+8FBrJSIOA7Yc7zt9O1hI+y111Lq1AtYNp8pIxAaLzmtR4knKLlW
xdNsyVbQc/PJVuzLMqTnBai9UhboXqDQgOm/WyNnqSBhV+vnn++OXr8UH+E2xelO
JbNhLY7kkz2P775b6LjS5aboLswGaLkci1MrUSbmH8MX/9xk7YOexITd4RYtmZdC
/7bJDGcg6+2mqnLcmM+SneJilqpyr3mPy8H6flfTn5zdZraEb9JtFSTM6MbLQZj8
gaJwRtFUa5wC6Uu2sU9NVK4LIthWOUAT7aViFlPeS8nXQwBFFXLYmK9ggXZg/GnY
pblNG2+uYpjbWWJcZzONAcO91YZjwesey7nT7DiYZwGAHE+T4/h6OtK2MVoSOBA+
/kpK8uoaKjvN+Xd4NiO686NNLAXOP23BZChpWphcCeS5N7uWzAke8xoHtEgmEmOp
9wMaCY2N9+dhvhtyJRz5b56/IOdQ4IWnSVnlSwSFloN8BraFyCDtHx9TA63O9Kf3
xIqIZz211F+5NlHwRS1q2xN1f2hOFL7vKOOQXtwQ/X3zS6DWxrYMd9A+V36duu5T
zgAXeQ9U0/aeQt+xdnFDJ5Ecq93F7FeyLnUW5kKM4rNNiLSRO7O7WiS9drfGSAcy
FG1H/3bKODdyd5OuN6UM9MdbWURrw2/vUZBl5Mq29z8B9wSVy9oUZ2TzG1NzqxVp
O3uQM8n/WDz+0QXlyQtsDP2yh4lOBqZUqwGK3IBetQ6OcRVMFav4x2vCOl5Vu7cq
L3cDbU40zqCY2T4Te6e9m/kTwM9wBcgGqxvsJJef0gYZc4/2Emu520WSotravkHb
ALOF1T3aJRP21eoPdyPbrUAe7r42THy6SWkeuq6r529L/p6QtaBlBd5eBecfJPuG
xsisSRLfsA1N9dQtVVgwcla0f9LhcfcTzEHzGhK1dyUsmqHDcuoOidRilA6tdT1c
ItNlUPQ/7vP/dvYNhjVaTeuAfeLL2WEa4Z5VnDJxlOT7t00aWfgkIJacbQd+mnng
bPyJ/8c0E5eWI07fBLRnRWA1nSAeA7fzaKlgKQBu63pQ75YtDKfVWztFpefP07RC
Hd8+LLR0UDxUfucPE1gz6QRV3ZdE5yYcxezAzJS7+NZGkdV9wDCRjtqRIHgBBhSf
sOXYg+7gi9wrgHX89aCMAaMdo7a8w0D/ClMN0zV1UM79hiL+EUGJNP2rDMgrVOLI
uZqUk6vGiH0LTCOlO95ceRtGmxcrKbtjRrtcGpo7OvpbA214KMKKA5hD5++1aRIJ
Fw8lnQkIw5YNdQhHvnAdbP/QQ0/d8/P9l9g0NtLXwRBAfk6HO/THE1frekjFPo6h
FUuqo6Mrn8oucb8cAKvnaDv3I8aGHDFcN3PW7rx3zFrbuXr7fkv3ZJ76FV3NdYP7
kRhdMO6oeKV8qIyjjFmQv+OFTa7VHGlx9R5L/rIdDeuzAwpy8/4Ho9C/8zkwVOkh
0D+0TmFSpiaiCzQtjN0UgSlfUf5rkIpLVYNh1u+XXpyL6GBLrL1ww8mVPGcpRZaW
AHUjaHDTvjiw62SPevdberoFgQfo6/YWSNP2MhEg7Mt8WqoaNNiiO8KZGXCzXmwD
guarWGxN6ehFAU63D7Z6/Hi68480G+4XJdUMnxBIvH1Rp9wvJjZlr1lnPOyyYY05
lhOhp+vVdOSa6PycUzzwOq79jA4BpJ6H0S5+osNRPzI8ZwoZO9Iv2ERiVEV9w5Pm
NbMmQmfygTaQ7fhtkIEZSIFr2lv++ifMHLPp6I58QFHZq7mZq02Qxpcpr6CUO6Mz
H78XUJlGn4DTlHRhcJ2uc69RUPphAQXcdRqa6jCyEyPkfl2oJkrvstPYEmh7wQTB
CbYnpaVs0fwUjgExtfvj63ChAYecFYspuD6w03RLYFn4L6CZBmFhx311bsRnY+r+
ptOl+niXyOHYp6MfEmDBA6+hx5TpnumgjI+N8BI3hoc+bOsN5oZ1PwbWQfcLP9GV
hq//j/NooIyxwC51yn2CAWrL1c5xfBpLR5hXlEmX7W+CpwLuhYUgwhYBsGcWFKWM
lJenY6mwZhiVRZAfd+W1gucnlHnAnnm+FLnrbjV03ExK9x+PZRQvtMWJXI1knqJx
KHub461blMacsbMTugE+ON6Z1T7byWI3dFjvdW1apD7uPNZIiKqktAnz6QSVrt+r
Di42uMynpkgJ3yzg5YT/dXlH0cKEywk7cl7hAkuoWhsKUchexv9ld74AFZMr6gGg
dvzPwIefRUAah36ehJekW70cuGIbr+aiFYVI4Te5XutD62W65XriWsYpWicjV7KT
Bp6irArrksRDS8Y54e21GMUF0ephvUfsBfAswQjvsfaeAgS7Qn8l+iApdAfojRNB
9wFTtHeEQR92Nnpq+4xunJqmXeM7AxPXN9kh1BovnZuE7r3OvFgHDgCucqw0ImcV
Ku3lKaQbz16JfRNQ1a+hgB1Mn7tBWL3xQfcfQKWEvRS5JUagO5s9NdsvEnXIHaJO
n5M3rz0YR05gPPJ5NJHppEISfPMSWupR12gQxKDssIx6eJzBvOSXg2QsfFRGsVoo
DckEI25KpXQWYIx0O5e288l2O40z4D/sisoqvArIs+B2/6glklprDMln6tr0te5Z
ix2o+QRGNLqveh89eZaEUb9EtvsXEgUdR0PAD5D08wsJ3QPPxn5IaDxbAn9L2qqP
zPGGZ3zTQB7anR5qpMqxI+zxZMu1KNPsGtCrXRmYzcOpVBv1i62UH/6UaH2M1qJA
VpN3vv/arArBPn3pP2bVI7p3QZoZefRluh37Lmvwgpfr0sDBHWUoeLWAZuajx+2x
6CT13isJJhH7XCvmbl/v4pbU8Zdhelp7b4CIG/BAkPHP71+G4rRFH3R0WywS7QIa
UuoW5TrnTi7yVqL4fCjw7Qt2+z+hCeVTBhUttLORWrawgdpA0rLUa0kpCv3AZN8h
2Rqh4HUH/Z/9n5H+ls+Y4wJrVaZkANbrRpODzl+c2H6zcootSmRpo2wEed1Q09kc
zHgvXlpsOYADU0Ccli1mcCPq5balX9NF89Ggc+yUgWO9lQBtUXIyV7GEmR8Ysrdy
xRHcO7BW1T+cpf0MtX3Itn+h061HgeIPTqB7eMKRBsZSghIMKqukwFzapmkT1nT0
lr4WPwTC1JdKIi6iaHA2AlGzn4teqtly3lywZBSP7KBXV3YKyeOhm7I3LoLPTd2M
UwsDy4/rr7Ecvs2aH4D7QDTaSrzXZ7Zd6GrW5Tdt5OE7j/sh/x0ZvqWp9UnZ1cuR
Ph3nosCF4pxn6wshi8u4AnaTaOz2aYkFDdv+Dpc3axwyRx3kQRY9shAkQ2l9KiD9
U+NJdwgeg2bBWD94+f4cYBCsV7Np77ouavqO+9knxGr92hRtj9YQ/i+e5Uyc7ZyE
DUe3osi3xtr6wObAqLyfS//L+DPSjq5AzFiQ22TtNewOCLQFeO6D0ojPNfxmsC5f
UJ1RkuhW6CYZ86PeqhlTdmk11umwJvqOb1Zqgdg6bcCR5M/DTqGxeZknTV4uWUd/
MIciTJPBnd00yD3zZq6nEDHEEbzQIEjwtje5DtIcILXa8TjlNgDg/2Z6x/Y+OBso
e2iaaJfTrAPetC0coCEqdG5G6JvBPJt7x+rlekpoJfWHjLpxkCjV8othjkqL/CKn
xpCpkB6mb/ZJgsGU1sG/jZw7AlcjrVMf0mqc/q8cO5Xn/qpBXC41GxaqbT/ECZIk
8riCf14efraMg4VZ9wUNpdlO+UrQE1aDn6Bg18QSnej/Jl6i5IqD7dQ4IUyaFjMT
cyAbFmAnKNfYkIf1uA9m03KGon6DykccFdxV0VwIv5TKUzub1HJkSoke4wkwugDK
9Y1tOcce9Ox/mYIOM8kSfl4SjJyCbgSR3BdDokpyeJpsn3KhzQsEQ1r6SZWgHizg
8nYl0ifH+AMgUS70ihF5+bHGRoEpTb3kf/VLhUjIcMBs5muIctwDXADnbCRUgOg8
AvVi3aKHJVK3O7k5LUl7mtFhOscZ+Atrp7SntmpgIOU2p/gztZ1ndWHYHKuRC+Em
ajpVUz8wKDFb5o71RD4rCCp34Zv6G6E+gw3YUUSpRmcv+jBEWhg6FVWbFZAdOEw5
fyskLP1rxuAtZrx6v9sik05QRFTCuJ7kIhcI/6q3pycV+6ZNlO4lwswwY9KyGBOV
M3X7w5OwZY6g/TjWky6THAu9AeDyttrf81xIOF6ttPzKu+yX0gFyBOlsS6TxQ33x
OkoCPRg2+EkYPgG7wv+pY4E3sBq/5nZpi6C37sJfM2rk9PKX+4xXkJLsQNjq3u30
+ya5r/d87/rLGAcinGlBbTtSdmaL7XK5zdFBbVuKAYRIkmgL6kO0hE1o8zcubgnQ
OiNCC685pKkZfwdEi8cLkrBFp9cyAxxIwL7ieT3wkRtpqn/FOStFjsmwScEX4nz3
3gdyaBmGjjapDCzrB/+MlgdMp8QcD35XGhtZ1kCVYXhaF74+Nl1+IEkthgBiuB9r
x+H86HJOCCQLS05eBZhS7yZP889Z88nsVwRdji+ozpkfQZ1rAGmbtna8kAaxVfd3
aMhLrCM01dZTVHibnY+Ux6emPgpNcI5PibZgcMrktW25naz82qnnsVdmDje0QaTS
+1R3h7PMpwKc8D+wUq5uCKSleStQq7ZX7Qu/nivbv3Ke5SvnTYXFTtAYVATIvxiq
lsWrBIKb/U318yT74YA72tI2teg42KvatQwps6iFu4KMzLsksVenQwMT6MsmN0sY
O3UjqHCzwm0dPzGsBzGtzLbvqTQyP/6mfeWXOjtnKLQVuVUxJnP/Y5LLcP4QBtNa
/PT6frCKkp5da9u1qvIrpPapk6ncF+t+t33PatVL6mYrAsYeMkwRALvei2JSoIDC
EZt+/IO4COWlmQaCP+qNPH7TEO3yIsf5tRiWCx+XZaQ4xcz3rWvvdjXHeEtw+cD2
Ul+fcK5BDg+j2rKC/4yjRV/Ln4f+rhSl2rv4SXeh9KTIN5nzwOGjGMW1KUKsnvJM
eUrxXg49PaYK/wu/NM13jLwYZWbj8f2HM7OpH3UmdwKbRBmUBCkpnkBEww2FG5Zy
E46FiMQK3sPiiEsQoWtSb7IF9uipiPCfAhZKMCemoqSwrM8MSGjSfgpWr7VfFdYH
rUIgt04MmuY4dC6WjRgWfMFe2cnjRhr52m2/o3nE6sTfLMoCb2DfMvJH40t8B0CW
xrxaoI83HYZ8Qi3h1ujpWwNVLDTQtsb255L+n7pJSjP84LMjVBzlKriESyJ87zws
baDsoMiUqc5OCvRwTYKAdT25N9bZDmv6Fkuz3hZw+G7jDNi8NF6GPpxuNNrKWNcj
noPf2KIwkHe5gEQtamSVlWf7F4U/eOeOBl20Re41m08lcGbQiUGW4M3Hb/ZfUkF2
dbucw1i9Yo2tLlb1jdkYav1s04lKlj2jz2CGRQ6vmd814caYTHep4HhDH0Hjrc6N
Ke2TJwB3p9C01x50Xl28+ztOYQQnUDbeKRBhpCq1jNWt0gc+7brYe526Kc1Pdosq
575jgTryQVRTJ+wM4TELAhIB7cnpv15VJoIn0jWNWRVqBlHJRDUTvbxKMLGQOqJ2
B3iDeXSDRX5NYNUZKBeSNNJW9LHzFfXzznLaoxl7+lSKuu1X4OQpqLA+ga3TTrwy
naO0AxoaUAm4jfBw1Y4VMi9V5gQ5gGl4gWs49vji+nQmzRFf6LR2QiKpTkNVa08r
2gQ/r7D7CtX7NWNirCASRy6BaflqQEP/LpgAWDeRZnPxrbZEQGO7/dHcv0Wj6pbg
HUaKXBRGc9bod7icjlxuoxqH1h5ramy6Tq1OS+pG0UtU3hYMmfOgL+U03fau72UJ
jPZwJxZOzQjcpNSGHf+jGr8gb1r900bPTSlYaYiPmHhr+HD7fdHeGc/NukzVhpLN
H6NUOEMP6G0EwXXRmkNdqJHRg8KzNnIeW6gtqISFiAME2QWC5nf457Cvai8AW+yM
LQiXrLrAYpZa5B17MIAn2UbBtFajEsiSyUYS5F+KxnugjTHdhywKAaUGP3UqOty2
Jem+AlPzC1tdM0eVmOpeVEkgvEEYJsqtFxRm7Mzc1t5OKybsdtxUY4LR+p0WvXE9
FSCiNxH5KItkVhclLoiJgOUxBYbxbIeJVXgGvxyvYvxObojVoExzIRHOyZexQebQ
knU/1bKDsT65bwYuLYZg7CADcSIUD9luM265xcDxPKgbHIwkGxJZmyQhA5AnwFn6
vIQNNY1AM/H8G10UU+1QWD2Rc6hRfnsC8HGTmzv6Ruhb3uZFoY8qzUKNZUW4fO4M
cCCZuvdWX4L+RS+/pRNfjPpO/ZvXWkXz4S6qM38xH/aXjdpEaNaM+dVocp5KMob0
omvKgIn6QlHTofs7P16nIIh1N5NfjfejF3yZLv5W0/O5YkkijHmUOYOuxKBglPGU
QVXl6sLOhCjhf4BMjSmStv5mIp39AJ6FDFbRNd1o9PzCB8GJnbn5aVY/8Te+J8yq
OP5QueRI+RC7P81knEos2PZrin5B+N0PPdDES52l9CAwjUDCMSVlm2zokls9ga7G
RDqMMNDdwGSGFGlQw/6OxzzA7aeDT/F7vDikwMeZb7bc9PDzM4K5p4WHiEjU8XZ3
g9Rv4nVTQ1pALD0w7w8FD3Fx6gxThTnn8lQ+mwbBnwkGk2U2N3iGZOf6+7PVE0rR
PqWCiCRgWTLF5fa0NZ6JDTQBBo+mXqDljglhI+WZc4FWzWDGutJ5ceAKidUXHx3F
qrvzJjTM/NCpYbWMTLXKZRJfKe8Sm3dfwZb1Cx7h599keCIL4p5tS0N2y6/CH34I
Ld6Q7cnx+ga+FoaaZtruKMgr8cg2Ko6/xT3pz5DO70xDKzi4Vr+wE4Hev9Mp0Tb2
YatvjfwO2GxYV5t/YalJCnr/OLDI1S7I95P+06tsraH7OrT3/PVgfrnXdl5MG5pg
kl7ITlpTHomeu2tmwyeV7tDSEh7V4KR3hDwKO9xB3ExqIFw3Zp3dNHS/cWYziJmb
PjYCblrcPz4iyg3tlxCTuG5j9uOKVCVm3y7Tl7i9amGNHYRC6iDpH3KBppMsKQDY
rp3pAFRmsLWmAAKEzZkLGWWs3nQgHau+QfvzWppiGMgChjZQbQFd9q48GfAm9x9b
SJwhIzSP/39eQF8h2jDXAwFdTK4z3B6MBnU/UixgRCQ7g0p19iiYSnZUijwNgx+B
QxfdxbqyoKihZ9vbBCNZ5xGDlK8E2GZP2INgK2ZUWViBXxM2y9NR+ChFiirV+qW7
yH2OfVbVFgSIEyTVGCD8Trmyg0O54T5NvWlwOtlf7jPOxNRZcIOQhmdVF1Wk97kp
AyJXxk4ENhJERB8zVOMQ0WsNJd9jyyWbgooDW4fhTLFouhJou9WSwmn3w10Pk4Sh
vyjouFEMJ+go4vYRb2mZDFoL+u6fejqSIStUZWTuEtls7O8QtiNoj1aRuOB5wI6e
71PZF6NDk3T0n4YCLfo7kJQZkpzQXf/0318FQSnoVwlmAZrYmcmQCESFcvB0Myez
FDRZ4u4PmF6oiYE4+MYIxypZ3KZYoVGVzNLZVpk/QG/O0cbCE0Nuroag5TwyeT9K
xqLDVFviW+KtySt3LVP11Lh1ySnircRG94dP1A0i6VeITh39l9EdRFfWWsi6lpax
7SAiHqQEw8StNkrVyFXv51UQeOdQbfZsoyNKZX8ovU1pvh01O0p3jgKgaDpYoNwy
S0l1eKtfoe+G53OCwqrmPV0+bRFP9Q4D9IrfXe6heBsmRBBu7W3aGB/7oLz6vZiI
cSQp3IXsyy8ZOYhw3t7GGbjdyIrRaHP780fv6kWEtChyhefCAb/rdPzgI08XJexQ
f8JKRGt/fwb2vw+58/5SOp4fJO6r9pglW6h1u8JwjaMwj/ICGfy/OLsMagNdequc
5gagujmOWvQp+igY2qX2xcr54yT/JVOLVWYfQmjSlTzwf0WyLybeep9/hcEnOQNe
YDM6RbsqcqXbboiAFjYpQEdnc28eUJ/L+AWCuEaBDH3Wxc/sXC0rJWBiow9G/Wm3
7SRVaCJB5OgxAWHRKA0zigIb7nmgw40nRz16bBM/8qKpt+6sfXo77TzrSeo+liyQ
NwD5/EA3jpxSeUU6+V1iImuh5DdgzXIWgFLbLEqQonkQ+Z3+vrww746nskAADfE2
epfDfNVWL5je2VWJD0EOqd1UV6LQge9w+hjozHNGKtpcieDxnnAUG1ovEjdIgNC5
y6Qjs24QNr7cD867Uo3igB3uin/ehcs2ielMjsiir/9Cok4hm7tuLjImYli4HzaT
ArWkaIoyQQeLXAkrOlJWk6nchnz4nEcrmNjJw76P3p6l95YSQS7KCIlj35YoX1vk
uqnCeXMTBSv/cmMWjpt2wyQevXYJ2YHrLWGJlY3TjYXuI7GsgGqzw7GQBb7MPjC7
+BrHnVy0T+2A9fj+K3gKwU9bmokWbCrLU+4+tmgOJbWYIBQ73LkpBPFGgbQYLxf1
/lSyy4/TlSZEBrhVYLns4fNr0Hfo5CsRfkC5cfE9lhDpKhaTTPH+hgBB6NIDZ0og
M7F/1UtkFseV8K262aga+FrUL58n91vA51Oua56murfd4/tpjnPa1CNj0Po30vbu
hxg2Fonm+spAdrc2sQ1cg1ZKwiqMMchJGocX70czHbrpg7clOQ/uZmL0D4rbObZ+
sHmspFrgIaX3i2HW0buqQx0Z1RY0gblMekjqcZDQX6vTC5Qqu52iXE5tvSMlPlk/
gjoJpI8hy+m4zmF1ODEG6ZWDK4sEinscP7vii/LSlKG0fa4/NHf02cHQ08ASvsDQ
howTYMCjd2RPQJ3pO77jCQnD31w3KCGSwcCTHj8bGy9ObRBpfxzJcK0VYX1DxRgk
drvPyw5K6ftLDTkPYjgHEaFifoVL3UVOOUaniaaozEAIpK3jbFi2dmiOG7zXi5rf
jPABaDw7Y54Cr/Qfw6/spdktBNuCM/T4xMWsxK+G0l32VpAQvsViyA18ku80T8e1
LrDWFjqsPkc2SWbIq4seWNQvMYGRqY8E/6+zZkjYcQe/8bnUxEjRw2EbDxUCUxIP
l2G1bAZnpQAI0M0zGLaRlh+E0g6+B28nJZKrtLvF87+8VytHDgc+TRd74z5F8+C3
GDZHViEvJB74Tq7+h6f+rYuIt4JpuVhjZpRZHspYlWuYwO/n9f7Hho334CzTo5QL
GvrWChUzCRuctGSQHHYWHER2b48Hcnmpm5SXID4a8ZCngtLg0wwKx4eEPYKWAzXm
IMqhI6tEpVcpb5zprUk5m9X0r8PSHf0aHby2XGGTWY+OkkdNR6MWkUvgXCJLFSzC
EY9jnaIrdQ+RynfqwzJUXOk8yKRgy24pK3ScQbc5xegxlMOUD7lZptfl8/nhO2jO
o2brfYIEt+ywARAh647ho/uevLlalxOyCo4qRlFdoOua7khNdHswD8S6lQf9x+bW
Qc5L70/PYBRq3n4pX02vbwXv42bUTbTbOIxg/z8Eq4q9l6Vw4OqBV4Pil4SPGbH1
Xu77gtmJZVZ6Swtd4tUPgXZqXP5W7p9Nj8CjRPEDmelu2lfd6cAxAonVFOzLlFEF
lnYmWYqnjeQc7HiJtnuVHUNOyUyHKj4ZAQVMhaMzj5YiBLSZwqbrT0TZH7BLaslm
wAxK/bOvfh3zZ+q3Ef5wfCdzQH1Yg/1YkQ3xQzUlCrewid+utztjwLGAEVP+a2c9
spYR0eNz5Rd9GnM3fU1/X7C8Kk9SHqvC7sEZy5rRNui5lJk/XFv5i4lLZNKjE6hH
NSqKkuzg8HW9oS9ZzHAwge2Lw+ZmgwZJkMyHQF3PokkZB7nKklmrQKJyqgEuAXoR
+MfnQE72t25vgRVlAh53vlUOEugxt8dcF+HgvVFboNml4LhyGIa/Nj2hIqKzXtXM
Xic0pTg+RMPf9BeeAK7MmAdatm4oyXFaJtZl3PjEcRp+Y9Yhdjoywq2ZxdHMlDLU
D6bmOoOVKLPnDGs3/ZY3EYuRoRkzIrVeuddMysrWYqDVNJdYhhHM9qo5tEKvA3BC
8aPIkhNEUCBuQgKIiwcSBilFTztM3WstNCPE2YrW7yUhSvGL/pkx+5loPTt987zR
Y1CmM8ZaGZIjoLQS3IqJQxJl1E5N/54ZyuxJdmQNyrEIPGAXrwxVjfquOcb7A5lU
2Bp3GSh1zeA7Q3XaXG7YbSqxbmUjOaJmALqUFMd0EllGfM4WbEciF0Rjq5TEZJme
Q7fa+AzysJ6J/hStK5tWF70ZQXvo8mm3DkX1Mj8cu3+Xt8fzaj98coIDmrP27z2W
pmneTuMqlGJyYJUZzlzeZm2tailVww7jRFi1DKI6T/E3RCLBkKn6ntZ3BFusAMtO
Vh5M5/afZ+zDnAbPg8eN9Z4VMEgrBLcpBqnycYfi064dOWmSSvh/9aNCxElx1pVP
wam1BdPj60txOgCBrAH9XYsMRnxObJcqo3xlg3rDmo282d5XGZJbEQ9K2eRaOhCR
PiNzmMTOb9biKFf2fWw4ItnJPai0UnzXAdBtCkFcPDEmH+pa0lnCwmD8enyQOdzg
i6Z15mLqrJVE1Nuy0eavg0Mamzeo9Hym/or1RKLrpXWw+HZxtY21WSxBGm+yV79z
u2B/Vx/RLmnpBVIIyFZLc/avNQIK4DUNAQfhLPQ31KOQ3aKx1br1jYvOfpiQkEgV
E3tdCvmEaih9HQvkZOqu5GmnYNm3NOnpj8/pnIINdKnkWt/6YeKUc1+utm/aeCsv
V0/KXXSN4j+MvyPh4lPiVPc26sQklrSPkTntQ/yctpz+KujueBm6z/1wEhkm1QFk
hw0B16+/vmhFJfM7uhzhrBDouRnyBDHJG7DIhxvdbdo+yqAQMpUe+cWru4PX/n4X
iNII+OnR7ofv8FIX6Hbe5kztUPc/nxkhCYz2IDeCYv++y5QwgH66gOrlhYI26Afx
wcz4SqWD4J7hyXMmGDfDc1Yoal1M+OHKnlCoKE0YdManTiwT23+nMc3ANV402TqN
gb1W+q6K6capLf05sFfnjLc7FIcIvaaoRXzLeaPL5PYBRuOa6Ee/RZ6T6zqSB8zH
CNnms1hZhpyaCi8Eq3k9Gwtu9LGiPuJCtQ+6Qi/YA6bh6ZtOfs0gN4J0zJDQtUaQ
OLs5MMrxkESZJTEzpKdc2rEvc8tq+OUJdlFIfHaQHy5rpSD63+Z6/HDdDRK+EUWO
/sShqW76pG8BMb1Uzjeeh/2wKwXsXmyBz+YY6FUCxil4vkOgGMrJywITqdKHHPU+
N0GDxh9h+kr0IcgEO9n3UWq+OBvA/qXTdxn2/0IMV6emOlJ8bivbeSYVg00ctJ6m
Mm/3xXUsh2tSeC0YDMyvAipocLLX9Ya9OpTw76xAVDaIcmny3hiFrBIcuimGr6Ld
6ft4WhuAbdzEagid73H+I3joHGODYoLKORuJUfHW7zjRpasNwF96TmiJ3fTe1dFT
MbWnKc64WWlKNC6paJnDZcqZOveqTcl2Ep6u3zTK5nz6LnJssSzrYJ6AINpxSWab
+9DU2dPsnFoOrKlktWINxs4eRjHSX4jt/SC6/TrJHqrbhW0XfgAeKe7QY5d3A+py
ZX538wjs6EoeyiMNJhPT1/wQuleoOqjomqFjbkllGci3IdHjwmHH0BnMVjbkFibU
41F66+5QYA2orAh4ZzmQDW0k8ZD+VAv2LNNa7/Hz+sQcwOelMl4ji7KtUIHWF3IF
qF7Rrst/WQSas31IuFQ4oYiw86iUFGAyp4gvHAEdYrEk4MV6BSRDkf4jHHo3+6s0
WftrcImO+SQRBH6IKJJlK0eP0rFSx8XyLHcBi85xiP+zdQ/20lu8ixIHSCF+4Mu9
1Va+c8XRb3VJRftpwYtGVL1kOg8ocmbyHcasu2spCI8Thm33SQqh6SVTan5El6Ah
Zq3xiytFxcBzGoLRnoBCTAWt91zGiDtHc/aRgPMvfCJDbuLQ0GhAwCk7r3uT+MnX
Y2WXTBCxjRJR8b3rumnxvRXClE71Su7Zo2FExio9TY0uoX8JxOTHzuQwMggiGhH2
hwv4pmNP4YRQDIwmZiIBxJfKOkWXTJ2T32vcbemu/7KuVVOf7blv1syNzREb2oPR
e5jPxX+uCt9HE2XELqt6pxEY1FlrT0xiaNuZ54+l3LguhLsHg4Ih/xNlg1StSpmD
9guetEokvZHC6qXCFy/cgNGJ55fXDee0+iD7oIC+VT466vietAEKsZvYpl1cC5jL
ch5umqS8CHsleApw4h+8UFzM0RCHZG7HpKBWRc1ZtHD1/8w3qdIaIklBpjW9Qmdx
UID87MLjn+R3BbSXSfFQoaSi/APE79EHMrpx3/oUcQrpfRtWTzzG/JQAumcqt7cp
6JNSDEJ2lv93gpsLQckai5dQmk3/Kh8dSfG/GUmbQ2F0k2ZFISnk7e06a7V1VZBA
61Icfcf4HWQSMirImcD5OkGx3Rrz+zm/Q1xP2zl5gY8gIIHS+37ZZq2GANfyiyuy
87gMz/ICxwKuShjYEA1/eo8Oxe2FEoMMugu7bO953gkEwKEd2gXYvgNCRL1+CN73
ypKcIDhDFxBlH8BsH+kQFbruibsBkFdg3GsnAsRyN8brgtK2wqi1gFvRQCSDPn4X
qXaF/FBXXdQuCLExUGp3mru9rVRhKSHN7TCiQ5CswR5dhM67R8LJqKsEaGyBGCpX
OKmZgW57GILM451C8YIdlHAbmubtsvxZ0QiWe5j+zyKHd5hzPNocRw5nybOJ2vrz
HJ/n8RzIx560GlDzVq0JjuCKXRtal72ui1nPV0HEIXLH0li5AFP9g/YhqcP0ve1V
QZQCuHtdcw1XabFqvFJoWHhhY6SsIe6fzr/rxbZLaqAZm/8VKRWmNJkwC8xbxl/a
OJ0TEs/5DF4e+yglak9qv1biqub9iN1RglS+1Go9KprGpeoHBz9yExvDOrByW/zu
YZKM5K3Gx5wxpkqg8uVJE+5KY/8qZ8hpZEUo/scUhYU3a/X05rXM+FrPM4SAkq9s
RmmShVYKBuSaXs/Q1rGq9VkPvmN11K+JhXTRtbXfH2oPn2dfn8J/r4n55WtWjvIX
mb/wYH4oQw2Yue/lB6GW4ZYLTtJSUuBsgEYF6svg7FVeXgGlPbfsYw3wyPE5geOo
yJZRGfmZp0XpKdo9vwVRV0zNJfW9xrD/+zrO72YL/Dnp10rNPuybssjzeAEuWF9b
ZgiLb1rhrJ0qH0m+nluCLd4sVwqQ32L+WneyyacErKUpdkAa+kT4EknBuixH+XFt
fnF3w/HQ9WtwIoKe902JpFIZ7l8pGHM0gyLX6b+ME68HlfPNBDH12tqDutrzVj0N
F929YVMtMw2N+b6rpYB2vCHH5/gVTC8KLUJm0iiT/o5fgMSM2DmdI/ZGNiZewloc
7dFw9xBEc/MvMzbctt2f6kcje7T6qI4xHuNKTZ7gxouqb2oqZG7sCuBMRv4zImQc
V/9atYAeJkKFRmq532AVSezL0FQ6LHxA568GKY2jgF4zCjctHd/btusnPlq2pehj
Wup1lteyD0zivYR7mD1iJPqZ8LeHfeXqLVFrJu6H5IRTh9YmhpZKaE9JcPsKgFHL
3BBc4lWJAJrHFNRyQPMrFuAc9yAVYTFW4Jtl6OFEADEBQxBR5N9TfZTgbvnHe9+N
xyYs8+VWiuQEW9+eyWACm0NgjWs9AKC/g3tjYsYz967M8DyIYJRw/lD+Iu7Q0fqG
g4h7qvIvB8louaZpzK/d2XDzYndJrd9ZDR/lFje1YV1b8ygC0Rk57vpKM/LcFSCO
kGlCbj29Tf95st1P0fbkiXEKcpkQHw8kBB04gPxbnQA5I5rdxzbwjhpwB8LQ3bUG
tJASwC307O7ddl/zwBWbcu3vKVSkuYMlDSHuEvKVTHwmoQajs/Jmombs/spbPPhS
PQt5SVE8vJzTfF6cMWmqG8NAfRhYjpXwgQXRc8tyNFstTGRIt+gQEky8heLJNSLl
KN7zRqjY+ygcRcwnEwvMr36Iunjwjhvmfqz5Sd/f5rPwePRu+eolqfvaHEhS58Dx
e9/i0WcLj4edbMJ6ymc6oRUszXkuk80Vlqr75YTmfAWdGp+OIVNPP9Ph+fO42DH+
Yr3pArGW50CPY7fp6uvTVcIMKrsTFajXBgRfhz5o8J5a1TqqjMHTtFZpMt9uaXvw
kMVONjj5MT4GiHt/kFNGMdPQ3kx/Qiamix0TDRlZICfM8usYRwCHEuLcvazQW+DW
D1no/w9Ar9ZosALC86QT6nBbtXid8fJrb7hdbTW99JJn2ClOQwNbm5U3ZGDs/3Yh
BozTHNYqz/CeDIPqabN80Kb9i+Sz04lXiqn4zi4FBQ5otgBj7wrPo+u9IFVVKsFW
vWju4b1GFITvggk9+dBvQnfwE7CsyixeqhzO/JDMELvAr3AMTVZeuiWyIqv0tLNr
AIv0JkxR3jP72fAuy841CAN1nAAVRO0GjjTPgxQiicYfMBI+6jVaR8dGi2m0XiCj
Fyyx9UNi2Zbiaiu7+AXxsxOd3atfYxakNGDWatIG5u1J0WedwJuZEANI4B9D1KWT
/E0xocH9sxtI+qxDra/C8MVTEYPHvK01VXFlYJLsoEPdUub2TjE/G80aEK/6Dh/j
wZAX05VBH0Yy0HEs3HylDOZyZ2EsVArHNCkFwjxgcr7tqM8Em30bjWG3oHzhZyWZ
dbiV/K3RQZ1ag50wo7QvzHkaOcanXocH3o3IUML+L/nkiAaZ0NEOXtH/lNcbh24p
pbDY692RQ8FDbp3DuxPyZgk+Hhmz1qNGuTHOa6NSygPw0ZV8AqlTAak49Zn9lljy
RlJr+gyWpQKXCDmWQZs9I8ZVejOk2ow2GuTyY+7ITufYAsfd/W6JNZ4wKHWGlxxL
GTbKTkqoQdsk36oikJhDx1By8hT5n3LCEaZEZcnA3We6wjrrtZDlsu/5QdFyv/3/
DXYsMakidvMtmfgSZ1Ww+3wlYfF3pFdmumrbK3v1Qb4yOz4Z08lUnS6G0GE4baxq
fc53jn+LJPlnmBPCjDe/FykMXlohaigXDVH8dTqAjLiR180CdaWxFe2nUKDIgJVo
Ak4qT6wCd2x3amCXHrCIJ3jsdixW0AxWZBOI/fg9OznweomRl0096iDY8o8S+EXq
oYhOdia4cnA0NSMSsWMh9t0gxnEHGKm5x1G3P9pCJDr9tY+TSqidhj8XvAqfEMX3
um4Yk68rtIVAHGy4IM+Xd26HypNx67sb8QUF38yw3RvEWLK+uJwps3Nh8ARParRL
5e0rPLQ0AUXIm/UcnXRabs1/TpTYSIfGfPF5nqiOY06oIFZRLo4xRMgC51k1peB5
+itLOmFqN7LYHxC4V/HcBTla760ZiVQF1a+wSd48lm7n24x/W+gdDHn324/mtKf+
d7RktiGDM+uM8xPxyI16TFGxBFg+enLhuXpjDUjSZtHwmWkHu6icl6WHrlNwKlmn
qVuufGPMBtPlC7BRipk0Hzj8n5Cwa3TxjzUF8ALDEdewKGzxK8a0frOp1XCGLx5y
gVL8/ZPiZM/s789HDNSNChGzGYUl92lZ0i5X7b5rgXcsGPzcSmZ1P8UoAAwDCa9R
IJWfOHT9j1GJpf35mOobu9YmjWZAKImPy7eurFzY02bnD6SOIOiCe0RAM+UQfDOW
RQ61Q5evM9tuiLEMWCEVSl6Jjb4+21V9oSBPPyDlzzryHwHAL52PkJhA92PoyRw/
exdi/yoBLZe7kS83UwTybyGO4xpeYfEj0+SFRDXGCAg6gEmM61KdSHf/7/hawJd8
0uQwPvMTS3qm4kK31zj7PNOxa9dTVYeSs+768MIlC9JkaoMgMRtJczJH2e87aPBA
xSgrkaa5mkrr4ifwbjlGRA4NJ/SmIg9Fjst/+gIoGhFzLmHdhubZwKVfa8jVSuTF
iu7Ta7h5f4fAENslwkeQEWIRkdr+ufBb0FAMf4kwVdZN5gDi7Qi+wWu8h5bg6GVd
zecwHBzlV40nQYSZ3CPnEZ6QT+ju+f3eKXxOqEZcAiEd9o/lkFpwXnd6PCqkNkAj
nudjPBrkpcifRgfexCZwKSyc4TQKfsLsdhhIq56gjqUBjfbvAQmTDWlFnhvFbe8Y
cZ9LpeyuzBTINuriyEUumDf+7bUV14nezafJtQ2S6aKI3548aIWq0qJeASXPO6t9
ZX15dHDCTG128BhO8PuhMkyHi/D1o5PIqICQuwZCp/hKHArxfA5tM5CmXLZlmGaO
iZHltSrqzT8Iyt3hYcV8njz1+0UzoOF628H0XSYGW4fgzGFCYLbgfVsJTA3gTkWv
26bz2CWtHBQ1iXOtJ4Eeor/dncdl52lW9KQVJcmSJ4FVyu8klX16GxvrIhwpOMya
jhLDGSDrylwFwVH/WwgCRxb6eUGKWABOWZkmNeIU0O8s4l86UbeeAXH+L8ay1Ai+
pbXCyFdbOw0a/qbgh+5SgxO70I9004xXxP+rGtPQhOYD6c6f5hJNhEE0YGZNWPaN
vrxXGUZdiYkqz/cqaOh0nHFATi3cCo5Ttc9VOnPfMrT5lDL4rHB72bBqYRNe07Wz
kZurtpQ/uQWPiPhEF88jXfuf7C3Xil97fDafVNvSuBIzhtrnhpYX9iEJSN6TS9aG
6umIWnT3w31/DDpUdkfmJ7hOxmSRsbAhvSXRGROzmnSR9iKklvHcjD0HITjn6HgF
tjSI21ejGOKbQ2OOC9fPKKgxTDHkqGHR4Xi/QlFHNqIbrM5uXFtzf5FqIezsPX+2
Lkea67THPI4mttgtbz4hJtBi+Ur0JvViSeNxvHBeES0oQvNZxU7UVHSsv4QS2iLd
lz3aO7sJ1dmkZ2CVbXLUPRqIoguEB4r4Cj2i5xFbBQpeWpeFQE4AfmoIFYHMxoRD
sH1IGS3PVuogHHiYiTQz5p2GMWNhnFzzwygjUIB4SM0uFz5yZHTu576QBawHgmhp
Cwt37LShv+xnF4kBtzCAVkXtrGgPdSLsj8YgsxCer5+dD/MG4mxbIlxKJxiRde/l
PaI77vOIaPCeTnvO7jYU+xRB1AXdotGWKuhsi36ieM2eUV9z2HbrPfxyg1Z0sbve
kJd9PPiar4KX3/oGQ7RR4VS/tRtR4oGYhvhTtLSMAP37NrG+rOSIMfNXFnl4m6WQ
8kWWxBNmdhWaUCs9pBNAoO6Ekt/bbcJ6j9J6yoHD1YcMhBYxK2P5lXw3H700FZCe
obIBn0oKBXh31AVB03FNpLt6Mr7W4ek1X1ptk2mtCSuUAhpOy61rLK1XiqVeEfJU
2ZTIpKjEGUj3RrBoNTQ+w/a0PCSYaRFrSJ0F3+OlSBOico7QHAz6PEjveiv5Pd3N
kRH/lsySWZhi2pxJtyOMmEO5w1vkozUt/w61ZbXdH9v80bxcOE/JB1e0PEo1RCal
6XiMNb+8q/G94/h5SrQt4CeIIiywRtuhHhw/V4lEqcbdHmEPnyyZW0BCi0MU0xe+
RNfIKPGgKTpG6NjKOTj8KZPD0ICX2CWt/kUG+lmOVFWvbsHuBOcxUGAbgOFSJ8Sp
K1R7tirD/gsoWxSY9aemlS7gzrPbepCb+3AcOLRYn6zTjX3wAy2OWVZMFtrW7Mlw
s6iROKPOyT36aN7YRA5gGsckq18cDQYdlwthpSmC7CxN0G7nGt7uiVdKSe8N6gMP
SX+QrCjq2cD2j9MoYLDBkWrXdExJCSG1HvAy/HbYMj47QK4iEOljYh83xAXQiSXC
cn7+9hnZXn7MSbDJ5YoGsAcj2pyjNGrSrJ9rIXAouHp8AND3shcS6F8gZSd7QeJ1
iPhlTU2rztrQU6R6Q8ycFh7BtpHaD6SrlITSPeBREVyzOoAycKjwBq8mTmSh/YHY
VVNoF7My9Pc8H0LBF/RxJnQI4cQRYvuoeNc8orGVHa5o4no6Mj8qEMHYsJXUxuTu
KsN7wqB/sdkSrN6tkxKCmo4TWEJpAaKFGNe0RuVeAPaZW9Td6pDzRK6MeY0mPbk6
bsYL3U7MTPyYJw26sgjfNvlvIRbHcClzjbvzocaRdiKuvSiZSPn8pCqq09g4uHe+
Y0qqi77Q8J+SwGi8QVmv6QbisxLYw1wfgahjpiV8N7BGHVtP2a0w871T/+1KOlT+
yX+LRkhYXBrRY7WFX+SIsHqvRIxgdnxiHdSrcUqJ6cmiagqT9yg51Xo59PBnC2Bu
+V7OOhGie4Le6B2vyyY3Ur/KxD6hO5OrwXnGW61tgg04NfmkoL7RrROX1I1xMjsj
kY2x6Jc4rDJnHrZhp5h6+nX04HXV4icF6YEndP43r6o5ZS86gdtU7owKdVz9NFUe
nDitSxTMJKutotovL9S05tpZRvxBxsz5eATafGn+2W2pEViLqGriHbQKvdZb/cM7
E0ENau+SqXPmmhkqsy0ZSaxsHbYWAqHyrJFUUn4nQawezhMt969sQBth5KzdF90Y
2GeJlWzUYHWRe80eSapPba5+DIYlC9QcX5daEvYFuxjYiu2kIQJCWxOhcWebLSlx
XYDrPAKtrUd5Wzal9b/AS0dmc+/N8+jqPD/MN7hSwmYQFfeY0XPbDq4U0Vd+k5u9
e3pGqfj/fLl2XjXa3gE96R1oBWoMUa03tUbIBPI9vO/pmlpjB2LVAveRwrV02/2Y
INdmqhD7jNYnkDQGTFy5Vf3yCyemlBPifkmnpb6yNwt7GhMLjln4B8DoRwSpzmMl
aL7Hp/eOcMNEMsjHDoR5YENwPW6EhEh1Kxb22bQ8f9R0eq9FqISYNkTVZqbhRRKa
KnTQ9JYN+BM5fM0340Ri5oViH2ji0fHtjZKvFk38fiBlqWdFrIPPg9S4I/GXqnzz
89BP8wWiMF5EaaqETkYB1IUFH3JlgPx/15EPalO4UzydvaDN7Ja6kEpThn7kqX9w
daP8aWnYWXC1rGwCqlK40ZWGuy8Uh3C7nlxiXJ1QvJxJmjMGsRtyyLYFZfjP1Zrv
TjXN9pNRTTArFN8BXnjtD4O4xw8mhzkO8UsCTizSl9TV2gumgwEIMz8OrmfNL9At
70Tfoer7bxa6uTI1ByV7WPBTWRm7XTtSj6plRd/V1LW2cy2xHvBWZ72aLz1lvAoJ
n+PK7O3Rdgv3Gdf6QzcwthTctfge9r6AweoquzSJBZUKbGZgVKUEsa9KMMVCew/O
cXc/xvb5kUHvb3jIqz2vbshx21aSW56H15OHlOWtHP7XvtdkEc9BaNRBRTr0ROkZ
ubMVweG1K1gwC7JJipUK7m6kWVqHlRHpbwiD2ruPHUIUWw9DMU3RQoSHxuEk19hI
kj+ntCgfzSoxXOOuxjqjDAUSGsyetKeCudnRRdB2uh8fJjf4Ir0LwrhMSgn2nDES
jJvFPmXg1BcjrWmqQdbe5liTNQDwvYwwYh6oWqVg6hks4oc9OxJIw/I7fCfm2Cog
9DXgG4nKJ14sGbwZn4C2hmA/jcWle5dgYoqD4q4nhn08qK11zfW3onJ/vyOG7jmM
/VT6HyvJm0ADmP9r7+aQxp37bHwI5BMYnNb61k5j4WsPpMocVnGdD2JmSdtvwCCZ
lb5VsK3kG/5pkcSVIQiMBRpx35PUmWH579Hh+6JqqaOinpWni+HAHJujRll+wZvw
aVzzEvkSopIANtkgQ17EyO2Roj6DRkYCSrO+xnPIcoKJX8HfWTD4WLur+aZdGLaj
fws1KpMTAX3i8Sd4S/mxuFbM/ZFSeK34TllU64t2N63MXBY4zmkv9c2yd/czRpmh
MMFlW9afB3VKC2OksU50ZHWlILM93QUEoqdDSb43o2MUhJQ3LqeiNd2SESTgPaSg
cD4TMqojhxGyMDriICIiRaxadlAa1ehuOX5PINVH4cYQZUqblyGaoyi727lGHX0a
fCzGTkOWVa4ESTbnth+T7nfA3xZmKSjQVbmKllIUgjkj9WYegZiTWAla17b468iz
uc300ry2oZacDstaJZuY2Pm8gwhYR1v0GNPqj8S3xWh6/GtBKaBLjp25PwePDpdx
QaMoupf/s3RldZ8GGE1uSl84bmy4i4AykgO+aqzH5BUK0peDFhhnSGQbuV9BbddV
xlFH9poN/GUCAL+gI8d9PqW9CcwDskB4H/f6YF4X85XyjoND2bFMWeaSD6mgZMnD
MJxybpU+3k/2zKOuC4gUrIJ1SCOdQyKPIjOFycPx40rJ0KVFpO/lETwhMzZVSm8G
8TYfj7QYUebzxKbbTWLihbx+zW7z3KNUq/N5M2iPMApebiVvFmb53eYaudb5uhda
RpX59LwVn69nxb4fT1L/OoXHM+6UYMtZcKcKoFbNkEfMqP9r4kz2effvC+KAPqHs
o7ygJy/XdtKmxV4ksCzERdFqJNUNQCLNJQOv1XsQ6efh7rWGa7Wj1bef3XcQizGU
trHxlsTzp9sRmNvJPjE3lvz9SqFIzXKbK/Ipmj/yd9p1py2CzK2mYHxEIe6HNDJc
ZzQLYy5itvv9TKMg/dNsOjP/jHGrF6VHINOL7Ep83Q9cZEMG28SrIlJuR0Z8HdNn
FqNk89OCvlbvtgLZ78pp/USI4SdU+pqtpbLI3HN2/2pTdajwNlHbhBVtybJUolq0
MsTPpBledy7+2Bd9IxlX9QVVmrDcDJRVxiI7fHflVW0j8O1RefsyAmiENZc17IdH
KcIsIbXtk7m7w42OCHwy/mUzKuQzgTzR0A+V4kI6K/SJ7Q/WQNQDB7H/pEcrY/T6
uO9YrIo/8XG80F3jpu0FHMw5gdI4efvX3Ccd6brEncfPbFeKfetUUr2q18HFHO5T
W76FjyJnen2KCTDC0bZNl7nu8L/iGFZkJ3Gi0hh35GM6qRzM0wFEp93Ur65odW8w
XllgCky8Gk5xh+q4xkRtWFUjps9ETE7a2RsNg9Ng/Y3dLC5O7Ia4Spj6eWoOYDy4
nRTfywVyCRAKGMMQo3Hw6ncVnoR73ibtjnFT6yknLEa7N+YVDxZELhcr/PgDoamy
mp2GLnKixgewuuuOUPREu0Tmr2I4eMqjN4lpLZywsoCak5qW2TZSFD+W/D0QYrkV
S1j/KGMST0SzNstJWt7unq0YHZ83w/SDJJkUveeh+3umvSnF0bqTAzH4qp6xlTen
kL16UxbOggNY9EGPcYfGNpe+kiZkUQGeVl2e/MTj+wwi40R3gIxNKLr38k2wLkQm
CEFfAcZjzVddE3B5nzKxYFGZuO3jYPRkchWlyh7xwzzXV/DRXrqoU37atpkSxySU
q0kMZQKxaLmnmeGuUCJTqujNrsdRSZF760MDPIrUY2yGM9xhKhtXCr83j+ZONyCr
oZ8sAreKkKjsUKcSk5EZqoLXrlU16r4YhuY1njL6l9tPGTsHgAf9+SPMr1RU1yL8
1eCXwuA3TtPsFBLc0n6wXwVyfL7sA7zW9VdxbQJyTOu/hVxMroGL84ykJMGwVgDI
EW2tDPkme5KwpOFKWQQewCJFw9252ngCpeigYkkPq/Jsp6Ia8SB2SHid5Ucq//Mj
jW1/u/ymzCO6qAXbgoOhLAIAjCCk26Dzh6onW62yZ2xmqrU6YJuKqQFK3J0sKrSo
3N6qy182q1A7i/9UlJSi+VtpxZYyE2A8IEsyPlLdLuwzt5n7gD6RBrVhqR8CtQol
odBqfwZxuimSCS9ZdLGavkU+oPgIgp63FMldjCe9gUJ1LNFC1bxGxWBtx5jmS9Yg
6ICQx/nCtx62+MOMc7NnNQ+Ga6dwBDy44OP4sVktIscmPh0WjtHGBNej6UUOOtEl
3JSGFQA3i6V3rbEnZkf1iU0a/BQXVfzr6Aq8AzMlIpNMk1KSEwFl27KUW1sVTp+8
s1lWkf2Z3LBQaMsY6Jn12N1PvKEk/emNmvj3VLHjwJBtUTWOGGhKtdk1cdNyG5Ie
CTLId4Yi55aYDnwoKZHaR+zRbWdNVv9/g0aBnGXbKNqPqihbK/i+XhnyfnZ1BK/u
WlLmqb3FJQ/xqk0fjf+0vHJpfR8J9BjTDUhtK0jmVdAG3Hfq9K7UHvty8RZUD+im
cSEO/74Qt4J9rJsGW430J/7p9t4B67UdsEEmxihlRyWDohkbvle9ULY0kAGZd6RR
fPm52FRhCSup3nNm4pBd824iwkt/H71EAnz04KvmTggN63dGjPPW9PmfpyO7h65R
8rGgLkjnoNh0gzuQmtmqfNo4/Ec6kiu2IlogDRp3whCgMSmydeu19De2LlbGi0O/
ONLR7T01evhH8PnqZAxRNdXctNIA+eYl8hgc7IdOZTjvoJ/cQDFkNiwlrwJwPamZ
Mlf9mIjrP+iejBg2pLDof/KbS2ya0zDvRFkVH8FvWFhZot8Tztmbri5gdDqEswfq
3YrpnAHWzBc1yd+dpwt65+0pDVYHfN/0nGcNhz6VmwlqJo6bK1svruY8N9tggG6U
OpgB3rV8o016Np2+olRKX76mK/arVrqktGAB0+DVVi2hAvAfAx+9+vnHl0QM3F8i
4elLoI35ljD+/3W+bvR+COkJ0w8KU96BEMNHDwv3gFsW/EpEZ3sF0w6qwlMOv8q9
kLmCYn2ATHfCMzs4KQBVv1NsrKX048VOHlFPBuDAffql4T6ySst0bW3g5pP9Aqos
fBiB/e6A/kBhHdnP+P4MtNe0ywt572AJYdKhRDIZcSrMxT7LG1NofbnTSZMOnPHs
wnV4+X+LJRNzoXz+pa2DDv/xDAGNI6BFZM8w38P605NkIHXgvGi/gZQx/572SJds
oiuOyfmEm7iFCqTmGOTJaE+Xh6JQzmGkeak+P8Wh5GO4UnaPuNH5X8VmrojbRRWV
1uhZe7fOLc8bFtVr55tFImfXC9tQSqvkN7HhXiWMyc3aBfeCsbrfwvjaIDNyQ4Lm
c96ckALcQpRVxhLKCaOYFMpV4u1u0sNB5SZFQkbbNUeDN1yRNY4XRs75sqfo63mS
s7DfXX+ZJXMzblXDONDm7uGAArqWOIpnfqWf2IZentC0QnJfpT2Yk+eIa1nHYBJP
oGB1q/VqiuMaJgEpWly+PhLXH3DMTHQ7lcYYBlJBI06e1D8kpftnZ7aDCeGsEJsd
tVC6gDivoXI9Rtubu7aCMmAY/euYXUV8EozPlFEd3gqjKNle1D4XeHKCvV/eUfbD
0gMxfwPXqqQWUGMSXknWg/wo0ZMPkrhE4qxibKiy5on4qy4hvLCvFGawJ+8JBNnU
8zyNiATJQ6kGJxnUaP71fZOS1NdZqCRV0o2itEj7ya5iUAP8sk3QQDSgOKguHfUt
ucuKP1a5Mo6pi0IbamT7D27b8lP2cCw3wcK2GaF0C9/yocaWuPaRseFTNxjdm/on
/E20TXQgW9CVbyP/uGnZhEI2y3HbFkTvnt9jGwB9STI+jE6DZL5nn+NNZdSdUd72
eugqh9dQWentno/mK4en8LwUycU3RMw0RAbt3H9EEPnV1JVH6a7TWwKX+f0e9j2H
vNvc8hh0/ZKEsxykuKRoYfSA3IFuj6zM1b8P6l5sdAfI9Dwd52kkav6y1ekW0tA0
C1F+5DU5PWC66gFPgiL+2nxMrujVkfHyQ8/pA4dgAjXWqptDAR4WPYxH9NP2Dk88
VGwuq0/GxZEEVNBcFWi1N1ntyKF/VS4ppJlDx88j0slx8UrR03KbuEJrUTCnboIC
aiUc33BNp9Gujf05+eVcDBqMXnmGqEpXmuZFTwt9Gynh1Em6QeOA8K2X7onD/1cM
y0QpTL6AOPOidUFIC3L0Ac4Z9ILBlHM7j2/2Bq/XOgBUwD5oGyiiovz6VtUigBbp
hIvaPuD6xFUkcydWXseU2Mof7PjZdj/wnS1HYhvUj5mjub7NlL2YyJD7urghmmfM
x591yf82AQtesuCOAI94/w3+dAx8NcI3zYO0c2seLaeFvuIlRyXognuaGMZWFyOg
N5Gmdoc3IpuYnlvALMgo+dksMQU6P4RRcmDYypXaD7StcAftU1lE9/FbITgJ5azX
xJpTKHKOAP9R4AhLQuy2jpecjYZOgOwH1i6jB3iLUVPZZbIeG2GkulC/psvLBsVD
lcBaIPRzMdbtdtoA/dQ/sogQqSXzA9uvMm82B9DXEWblcAJis4uUj+k2Ezb8jKX6
q9F5g48sHkPnmsqyejK619eeJfBS0ZcvXzT3f2kcMRJPz4TSbj7kU3hD8ujkj5og
CoDcIra1wTS+VX4lEatgBXuxca0tIQ0w1XZvCLdbLJNfsOp1Szwq3b+UivowPaGX
D9LHII6FsUKj7NXY6oD7FLeKR7ghH4XVLIztWPLDQm2aOB2B+HlOStRZlH4K45Af
vGtzCwbIEQakhOWh3sXWpOKQbQjcT5N7DFqEj3pn7piPo7qi4soQrUFDbyLMgB7l
tAeypulgY9At3CLFmnAiEOHymCpAKAZDePill7t5Z24x6LzdFKJnRQo++8flCFFv
6OC8DKWZqhuZlyuhzgkEPBDvgjaLu6tiXcVR3m6yWRlK9Tc4Qc0C/xcownkGV3W4
BGKr9QC/xijnw1EOGOpze6bUPKaf38huyQkd6yoais3QXvqYPniPJrYiNuQ3veVy
n5eetdVgBX7oZbYH7WRB+RKMVc7aVZcrSOeLlo34rbT/Qkfv5Y2fThTWQWTYuWfg
1lUA2FF6KGe9yP26IZI2LBdAkLn8jgL1uJG7a+/+1P8gQMQIKn2eCDZ3JvX4Dh7i
0NnDRYT/dOYU0b3vVSkxGAx6X+KlMFv//l+K+kJ98vjZulcjXNByYP8c9g4Pkm26
fqPVabfxJnVfz3zyMHlgzD9FDfeICXy2VAD7wuci8b6MQxUF0SGyhjb8oJp7TBuv
VTf2yGlPULuh/A8UF8cLA+KwZL6kmh4XE5bscysYTVxxYXHPzmUq6Ia2xJ+7UoD7
JcF5I3/UEKwcygGOTQqRP3m8/0wgAT/U3FP+buLJkTd69HmYDyi6xfuIRBoX9GtW
aSfnMmkeTuugsbwD2C0PEGXlfx1NT+ZRYj3QBaq5QQlKvo9ZSXSIyAhf0iPdBct4
kTPU6W+le+24wHLbyjEFuVjYZmzGQ0G6i8xiYhPwMqhGWBUhyw5/cvK3iNobQPQA
144EKznJK6k1L3A8rhZX4YqfMAVYFO2R3/PXXf7bfzyDQsjZ6HPYIC6ISq6Csl6E
Ce466wydcjMwRKnDmvKfNkBQvdlgfJdjU15RQNiDLah+mW5P1KK7X31j/N32mgb7
+ZP4x4t8DVHEgMlIesDrWx7qWp2D6K2Ei7ZfjDpUxy8WcCf6Ie6zVOmpSONVj16c
4pYY2D2SAd5x1hE6+TdzSHRO15PGbJPO6Ouah4dugAZxg8TmsbIWk/eLX+HoF4WF
eivgdBfaGcPfkHpHY+J3jkd1NHScGgAflpWvajqihHMsAkgcIJuN8+EVTUdh1bsO
/jEA6N6nCVw2Go5wbzjfDKG8/evDIDVK4ut7tnNHt9khj8M1Lj4h4V736SeNhHWM
bx/83Ley+kCzLcCXyfNQl3fDkEjKG1SnqbF2xtlKmY+zM+YyITOoBxbUXQG9mQbu
EKTP6u20OfgCylJTHfO+ZodBIkI6Ap1A4hBWkNfvDgoHY3kFSe1RgoNgeOLG2phZ
JwW3d/+h8e5CAfDdR8yEIOUXTggo7O8aZg5jDfbL3Yfjqiy+ddux3y0LtvvT+FjT
mvKOBk7rxf+L66nOhSP4qcgel/dD/qDGn/nYmHA9XkLqnhXrJcwkz1n/6SdTgiX3
xjjOkvH1ghBy9CzoTZLTaV076UTEAhsmSawWhlD4FBzYo3cpCH6Et3AW3vctkgX0
Y7p4HUqudPlFflsan/s2DXDcuFmoecetQtkTVVE47EV5GNIpGZo5WGIbmRe4heli
BjOJaFk+otvjPHWB8VDmYp6pD3zqbMbrneBvPJrFuu3biGEquzjyQjZwPuBqPF6M
VUPFJIHhRG0N7aY9ARV+/yk1Sk0/MgzRJonE8QtqRPpdxLFf1VKoOhGb3kOQD6YU
SsV1q0R67+dckOlS7hENCMxJN+XsceDzleJJAOzQCFKWCAa/qTTnQ8uVIoQnM1lD
3fpaQzewCkXGYENDIA2FVqLhrB7t8wEog/vV9KZmrvMCw+fjDPUAih0MleqKOgWJ
ZIs70a69qyVQXJy1goabIupR2TGzRUBPp4Y6Sj6C9O3wM+SQwDn15ksDuGdIVmbH
ipx2GsOqSKEA76mG3xdQoc0eeOaAzrnapKiIu+fCY2h6uhxpn6A1ok7oyeV2XLQL
hanamjblzIz1y82VyryYfmaNFIy7KgjFFEX79YaK4XFf2/UebxqC5PWm5Nx/ogYX
+iY9LM41ocSCaRK+6BmiiG8ds6e1qhuV5hV+fBv+185Y9nqVAsenwFpxDyf5ghLI
ryInfaZTzd2EGMBHe4CXlwuPxBqIgzyvlg9+QzmeUqochid+Rl+PgagulHHDp51i
5LwhAgyVjXLHN0lcOkiWNdadmmeJqQZWY/aRDRRXf+SrSYhNNZJ1KedrBpaOLch8
ofFp2X0T/sJjMpIJPxMBo0L+gXJ1tFubeseOjwc3kovBch9ldhDDD99fbnqYF8me
CshgE42/r17jZ+TsILzxqcn1WKu71PXRWV3/lUDBOCyBqsZ7L0vUTsN1Dy8MN9iR
DKsd+o+nJEAMgZlOiLLIEQpVV+GfwhUi8gphSc9hcemzb9IQUKtOXmkcljaFRKcF
OYfvoqA/+4BfDK8ht98e+H49HHBFU9kEdL5rMcTA1Dd9V4lLb3zaf3+Od6eT9xJM
x7nPIJaeNtHz5ltxaUI5sPIQlFG5Me5tNKE95h2B2nxPZSuDcKyf8fVv1SYxqYyW
IwnodI7qruStZ4Vghf+YKSprYhRMphdi7jaoXIiBVrUCB14w+RVdYyxdQO1Jhyhv
3dMx8VVx2cpyiSXM628fuBi9GAkK8u3Jjv3nEJakhYVMCe3dI9TQ4dXCKmLQhvXu
j5+CZ+BNyzA/K42YhF0o8p9y6UMu0oWz1Qn0v88n/jFW2RLPnrJ45zrN/E8n87sm
f9YgWKyb8c7wCnYDdmsA/uD3nXVODQR0SM6ZRm8ehPFmfFpsq76NfxBS7qQGrcYf
+v6gT0RtcHtsj0Y4P1CbXrZYV9SocT6ndfyKGB1KrBVcWni2Hp5uNVLJ2nk8X6zz
8qBiVrWG4i9CWzGGjTw723lJo/4ICXmD7eVew4rIAhreHyDy526WDuffAGKA6Nl2
ZHlXA3gUVa8I5sMWUaioGK8hEqDuMR82BX2nVltI+Dky5w3qKev7MY5D3mbpYboq
BtLpDFmoJkx8AcKTfCeh0DViz5eDfbE6dopnn51GWQ4csg0kEHh0P2baqBbcKcNE
nFNWjGsOpQvhh5ZEeWO5rnk2vcnu2cTBNVdE+JF8RrB+GBX2eWvtaD7N+NBDSFas
Rvvn4aS3HK0DJt94I8INphd1+JfsEnkkGqIlg+K0gkumsEyWsYj0qcFUcKm+Si5J
6FRQjr2Xd93zlhrEM+lBfLApazrKOjGqJq46IXvFMxWMD6hKwzpNtpS7PU9r+hNx
N8c71n86uLFKdyMnv/lYdn5P823yyV7iDZCND1VAcG/JK0AsTspp6b9O9JMPilJl
7+9H7Xjhm29pNy8W4SpDjOYVn/dLMFc+eXRbdaYKbAVJ5wncwaFlIqwv5cw+/AEj
0EFcDhQv7Hvb1xHnXB1YCQ/L5Ni+DDtdthHT4LJuBlbOh1BZN/u5R3xE0ujR3ATZ
tpLdFNoKIddoOOxEd7+gVnNdnT/ZXT8Efjecxv8QHHNR56Tx9GkkQ582ZA/oHzVj
G1dNRkD7svk8vJdlVD2RAePQp7Dg6UCiyqCbWZDgTjczzTRNa6hDqSwtlgnm4KXs
7WCventoXPHvMTqDi04vUBTGCtvAxMNkuebvOSNJTP9ecR4SkVrML9u4KYCvhMCc
D9QC85HK4A5YtVZLwosfamoKR6u4fM0jCM6NewWC1W/erTXSApNc9UwO8WrblRck
1cONkehmmWvPZczhKR2vpG0r+lSPXA6eFjmx3XfnTWFVNCPPH1uN8rxh0Rl3jD5x
jsSjwxOaxrQKUBypqdwGvgab81X2o32GgEdS++5TztdYbgpsxUsk2hTtcufaG/tp
D/PDT2jQOJ+7NoCQbTRNZ3JuhLEOIPaMUBQuZw2vI6k5GqjTYBJeA53gWg6xfFCL
JcGLYiijjIXsKsDhwyAI2WUiSV5IY2IRxyKyqs307bwDToahydnQ3F/d34QQWbyo
rjFLwUrNY8ygwEBTL48IBKTiL+iGgJ+d0/sPc3SaF/kQZHImbmb/n6rfL1EXI1DV
2fS3kdGuL6OzyW/EtGPOXUUmoHKZpUITe8K2e5y/IIVg9AVFFmLOjxTOcwq9v0UW
/9NVh6Ev5nD/qkwK0/ti7RsJc+8cO218+txNaOG4Xd3Zu17HGK5N8hLDCKk626zV
IJ6VahnEaNka8aNBFmSykbv2dI8/F8d59/22iUKTnxt/TQZGDktyLTGtFn6M9LTQ
bvQECzc4udw5UWrXPi1mxYDYuMo43Fxl8YqMmRLbDgm8iEIEGMnc2TiEmOx3oM2R
OmGk+8I1BORg9KvLdts2XO6SWIwfyINmRg741c/xOgioh5GK78iQFVlIBNooo/2v
xrMUjVWjxdVkdSomhPeXfuLBdHvV/OF2tmYSls4C7E6sLGHAj9qG2hANZp4e3mhq
1eCDcz3suE0SDgdTN2uowWvDsBBcCFXqmb7XNCQt6YNeomDKBwZCM1aX7g4T7oLm
YFmx1TFJH52iV+Rbl8UtlZHOPHG2KTbPuc3cdZOih/RoHVZNyCgavjvZTbKIfQAX
+piLHaOPo8G7FR30wP9kG8zT7TXhX0Oa+oI4MXjTHeyAZ0hHrYF0anHEuX96ukn0
s2G6qDNSwoBmndvaV4PvHatsd+trceh+QGJL93CHrMgYQnNDU7h966+78tPFVsOQ
XkEnwB+UukxtZyKTG4p59/apXb6WNKQJWuHVcBHIPp4Jk1PLGSYt0OTjhVM/VRHj
zhwbxFnZv3CyE5zqcOCMjsu8laJXGn+kl+vR7GF5BcXUKBPprcPS9WklEYZA3tDl
AuduDVhyXJf17X28YLkMddwPY3Db+06CJbe/NqS8GjIivNKZJa7JHQoV7z/H5UJV
ewTN1JTXU3pTGyOptOd1j6UVqmErKrrlsAPzYTleMQNdVYgYUt22HjmkEvfV8EAY
NdN84W+WLe7Lt4TfrjzPHBJNuC7/Sl/cV/V2sr0VvE3yfqQAImYApCaOGKWo7M43
3IEUVYik4fLcm/SssGpFIGBMagKhq475eDpJhYA6ocezEBRa6EMMjwTrTYwBg/kG
q9Mm3yDtCRIgKxEJM730OglvNkYt6th6Pl+3LOcndQ4kcdYOVtct6oOdGDdKemAU
mHSPoegHVsh/DqaCOQk3mctJjCGaMK1iZL2LHrnMOHZ8maOqSqjQ2I9IXK9DUnJS
kJM4ShB7cVgWcxBymLDi39QV0/EP94U9Z/njG0XerDcgz8+/QIhdFRsIN0MNGyjF
DKj9aNae0TEhMUHyY5tdUT4KGSPvbEFRseZw7/UjT7/hSky199rO9cvjwEesVN9R
80FFe1sDH79I7Q93S6LewEYveRdagem5K6hleD1M+MOKrKdjcxWtB9TF7S29C3LV
x4Xh7lIKT1+hWCZNzSrUCEM08xG/ke7q4dobKSyVctgSUonR66n1bAzwrCvRcW3p
QjwGNtM4Y/U7XoFGgEeO333tLyHqGraEwXI8pkBmOVMjoU/V3OfZOjeQP/c/ut2f
l5f2chqD+Eo309VzK3By5CyG3E1ZGxtG6tXGHfwyHa5fY/g1tOscWMQZ/bxrr6V/
8FCG3yf4j7J1qISgv4Tyl5LelWkKB/9XZuVoi7ruDkqmPzEN3U52p5TYX8yIO/Pz
mdm4ffScWTD3Dp4dz6+xIiURf7FSMuHvVTNlSNejomoYNE/nXo+226Pe6qoX4+tg
dYLlopDxQEb+TqnqpRRm/bXhG9MHskfs40roNuvD07jkxsA1vUR6yuF7LautWyMj
N7skJa6yI36XRNkodwm9cdw9uD734Eq0ulfF7VtqLwTPvCL1LXatZ4txKE/q+ion
yzWW9qvwUA/rk2YmCfMkBUkrOOHL11eDb3/krwRvTrAUdxon32TVXF32Jn58hZ9q
3ScxNm18dxbYRf2rbHp1ojoiCtQA86jidDSis0wwVfyP/t88fukfiEWbEy/QqPDm
otHj9DPywbwvVDTt9WhrWSH4NhdZZaTGV0fU1sXrojyB+avyFVxSc/2rmXzrjLhR
TIvXnLiK0Tvw+3Zqq7hWNayjwd2Weyj1u/wVZzaB7NxilKunaeyQzSSgkJHi4fke
2B5SvnwuRnuZELyXtx0g9zjuE7ImtAyhXvjKXujGIxccs844VHBzhVaRQsht2PVt
lXcSahuUbhqAiEtAlUvGlee1yFQVdep2iDbJtkRiNy4P0rgtPJUC9OJnHd+bxCty
86I9EffIEOTv1+vGCMEWX/pvD/rJ/lLXnFZ7vtJm5pemgIkPNSw2f/RNDUiqfWmX
U0wqfNZioJM6i5y5hy3Snj0CMbckAsoNUS7CiXR9J1W24Q3An9I0LDP8P96jwagO
kYImZ9l8caZ8EzvCIM0tJAckBvghYOFHzrzE33veDO6UYNHsLoxmppUJ7/7KXIIx
Id29+1P480p0PCDYwiEui+dkqEdVBp2/E9wr2vxhg6OYsPQu4xRztO6ODqEkFb7i
QusM+Fn1YBLbQ7pP/LAqA0Hofssm78/qvm9VG22l5UR+DBwYijFRMy/+6uKy1qpn
RDUadsclG5/1NoUoQLQ8VPSkiDGXkliWA/JR/km1ChbTRB9Pjl+IuMa5e2AatuWl
9aq3mnlBXkyU9ybL5aIOgzarpxcYDK/auwyyZMYDPtuaCg/WQktjZ8EQL31dcNdw
AxMJ9JAzH5XB1dnaet+vW6t1YSMrxR+Aec44OcCpc8J1b7HBlDtmDjGTPIz7D6/u
UDsMITmslWCAQ5f4rR3snz8hFRQgMXyW1eLTZAXmeb68j5KCE5BeyowNUGrhBAcP
PA5QUZAdp13aSQYel9lP7lftik40uz4Rl7Uq3W2YDo3bgCd8NcupizHnKYeOS6C9
AqIGyVe45VI2DN8VEdwkR+MaapJWbVA9BoXPflhYJvA5qQImLFyEhHuaw6L8bDHR
vil9uUfy/3V7UlL5pN39orxlAYphFgKKS7x52NFMr5bt4oCQBZOyyJNjLJtCY8HX
DXidY2SFbOlJMS6tYmFyV6oonQWkkMVyLtwxxkUmxYQKXd6NubdhHnPGfB+9LNXY
GxoBIlgwWzPKSvWRK8g5xy8OAgRMbkb09z7rmfIeNKuTagef9YonnDOye5qJuGxA
0uAU6dYIgHydPCQLCNWglP1yHuuVSIEi9KwUNsW3LQOOkb4ARTgZlQwlCXwB1WnW
l7ZcvpnG1NHZaEtiUJbnx0dT6lP8VNXcU6H0qHoiiQ0kuSfD3AWVmjIsxTsRJXEJ
ysjMjFlxafKAC8uQ0QzIeyPIufPz55zsydfzvlfIrra3f+kdifVFxvFmwnQJ+UHf
9zyqYZSz2Xn1dCNqO2fydSffpxCBaruldV378hKlsN4MFXGfDSclSP5cWWOtkvhG
62RYP5NbJoZyxu9PzgxvUp6PqcHp4aeL/e4bS9ECcUXiHP9n/h1bRz8paRV4yZsa
gO3RgrqGop6C2cbXvUoTXq0qVMSzDALclp6bQ+Fq1ZEdlyj/DFKKAiypV3rkK8I/
ywasETjfe1p8p6LmMfMCiL01B8G3h0oPJDyH+3y2BhIhKZOBm7CcBm4Tkmj59z4B
r7c5RjL23QkPqs+89Zek02yKOJ4lRyHgbVfuP8K81Qk1/UxpIQw557PnTGnpln0H
IjNL+Db8mX5+PmjzzwN+nX6feyt0DVol9g2YCmUOu4+U+vroAiYAmWRTnFKqUn6w
xAoPuYZ4n9yRUvNGoqqTidLanRa2S05pFuRhr/Z2OFaY4ZFUgBzzE0EvrLGAbALu
FmoVOXjHTb7pkEJtDqqzd9Mq+AKUHm/gzbJlCPL+yV+progoGDuLF6PXUDBa3CJN
VkmjorNP2jHhoGUt3xyCZK+ynuOyizZSD52ZXZ6Ccf2JHINtmjKnPf7R//qqa4Xh
qmEVnVdPaXhoTuN3wYZFctC3X3FLYl8xt1U+j5NM4xhrS+MiJLJexcu3fAC7ojBr
gcuRvtg3fI/idMa7p7a8FlrLvZ1dFWyPyjqpaZXwSb8GuKKL/vCsi91mGAE5C+7p
PT4bpsqjSc4hFDkRyt+EyGLV7fl1wOigK+giU2GCru/cYRW7CbrYcXsbMwqs2n1H
CM+lDQsW0AWZvgqZdc4Q1UmyL3pZJWaCgOJJo5Htf/byjJJiIbu4cWx/VPJq+lUL
f38znKJI8t8pNgXzERMF25LUrkdhTMzaGaErf2yD0wvmvrZL0PHg90uupUH3RIRo
udXRNPoyUj88j5S0ws2GWrXG3aMCHuR4GPuevXhVSfM6G7yQnWv4OfKNuWwRSMII
7gsrqlxW6PUSRFUD+cnOEnq+OQDFQM4/5ZNSf9KowDKS1E3NqJ94303S95gaymkW
Bd0CnwVABSNdk/Sl1fxqxO4eS6zH7uFVmZwfdNrt5MWjhgON8X5IUzYd0kjoRBUI
kstNMIvHWhdNNaoO8drX64a3BKOgkIaf7KFtbXOC5HEELq89jFulumgZ0MOcZQqm
F2nfjWd7kzFYRWHEw+zMnrWE6CaIpdXtMKnDnIky9X9wDlMmgpCLs3atGYR0dTHO
9+bOtnsXft5T4aNppK9snaj/Hn0+DdG8G8DnRFN2ShiCBXEDFMiH/k/W/lHBkiuM
PSg3MsIbS1qe0RHR6sm3EXNeDgsUKbLMkKOjNvzWJuKAaAsOVeOrukbsLECfNI3q
wkLFD4e8OZqQ2+4m2XNlTEyWDDuD/pWiUXQNXnFxaYXeBldq5KRj9mz+ewsDGKkF
m0OfUgDYbM/zHNoUlCDIFm41gWvWPFpbMdL+/eUE6oG2pOr5REDWA9i++egmOBeh
muOdJpOWCdjFPX87mg5IETzoEbM4Xzn/iOChA+Ne+Gda446pAB+nY38Z8Wx5QYx4
LPCaN/iL91LBZ/5M7ay1lfydKSrpniCEFMD3GdQqvU9p82hLgDKWtH/N/QMMXUPM
+2+sgoath8m5BHrKa7TvtM7Q7Mhm4iEDBybHOFZuTgIjewTwS7rfKmAmsLGwm8nH
x0g2cQkTbFAnper3ZmLXw3Ns1YvTTJji6JLdw9nHW3YVtqsICacT7KyeNzcLwwUX
vwDZ+jBweG4um85/capxQr2DoS97ZsCl9DFpfKQaj2RazT9lZ0UiNtF7Dvo+bmjV
zInEx+2fcCAUak+oaQl5ZiJ/tCYMNP24HEy/Ue2l+NiWaD4cXNqBbjwUJ9Rh9Dnt
vOrY27GN843O0RWQ4v6ayHiWFYwYe9VlXHlwSCp7SPzBqrRuTvcb/hlexycwRYeo
HBCo93gLa1XmYY1Qm9ZhEvNZxYhOTJbViZfKghh66sBMTxe0fyRI4qimNSaEkWK6
VpTNTZNTQVuLp35I5210Kw6nSQXMT27pRGciF5Q1QqBw0/0DAZwDqeVRD4D33zYs
5Wlt1nSSOKauESzGgNbv0xfOEgOD7kSX+b4rbyTfGy3uXGEK2Iym63EebR79+bUB
N1ozgtAjh07RZcv87a7Eou1Z9PzRhkG7UmNJ7yyFMKr8EWq+xs5Q6IYQGYetuc6U
qMCDYriczNhtYcwx80wlEt/WonQQGGH5fJmMv6LC35qCt5pXsMOcBGhyLY804x2Z
+sJLcOU6jnaj3YlxLeZ7VQkrljor73+S1jU3A+0I22rZxlV6kV+Jpdr2JMwrQx7C
AOVXY+VlJDGYV3p950E9v2CLr/7542Z1X4FrVjyhTbA0tHPP84o/PE3Nmmj//142
4MUr2ULnR8w3yOs133kEdvcGKtCBnstAMtnuuspfHQXOff8vs3LTSklbQQriJDau
9uexzUthwyUQbjbDIuE8+q1HgMcW6OhsEZSNOkZaq7li1jAo+XLfBCENBdTwuFxG
cqINFcNjKGKK2FUo2XZQBkpxCa1d90hBbbwObd1QtasNcNvqPcL+py2OwyJblDYP
6xlakQKbQODIYSTyr3tRsQMw+2j2Cgs5EROrF7XohUWr+WGSjmL9xr2Bft/tuHiy
T0LDIQAs1atPGEGsGTYY4W6aKFQ55UwoJQ4te0b/lPkvqoTIr7GEW/5mgiRjiB5U
vDWc77iAXpBQi3MRe3YgUhZlyU4SCLj+UfPq+jGng2D3ezqqeYh5kpgnPMwLYuSZ
iIHIHNM8eUcc1gK2YhpHk68M/EjRBhCMax7nPe1vScCP3L+k+UIZNbeqYJFHbglK
b4u5Eb56kJ2O975fCfYyO9iTl02IByZXX885WqDPFSszHjdR7DVPmJl4cUmpZS2x
rB5pJ3qiULcdHZTf1pWARyuodxFZtQISY6eOENnOCJ6aCpFDKjdJosVzHMIUcvdH
o8eKLshkjs+POinV2Sr7Krcl5Py132MBwpHuRvzmkqKjpS9McnBs7mE8CLQb8z0Z
kHbD+/seiQMvCeAATlctN3NSVUdymGA33xgMOS+VWSMDZnMhi/MTnOX0LxRGGt18
AAoXH4W73CyuKGQsgn7x29FjxBCore/+eIpsETYVI7H3t4Maxt8BGS8ynQGKUeGX
GQwan1kx3mbcYw2t9GaVN/Ihn5jSEhn3JyYI5z5t3CxypuEbu7T7fcgh6bXQksrv
apTi/mGCj+QirphPRLcOSy+QzMunEkx9n5XSZ/JrcaM85x/gAxvPMm7HaQBezpjY
ejq1cWUiJgw4C2s1SY5Bb0g6TZs3APhrjnMgiOjf2A/KwfuWDXMXnHMk0yV2HpBb
cc2hFOTFkRJfK8pwIBEoiinJF44KILXHD/VSTfvSe1rOAxtgmGjCJb9lqLulDptJ
yW4fxlNFDJZFPfd1NcPHjgEr0WaPhYbk12Ztqj9tZjjUabbTlPChIGWDMPRtZUAs
HxUnwhzRZ3p7HMByIZVQl22mmCaQQ7ugkG1aG7dpj+pgTPNPbOYjzmv9sa41Kg0e
di0p4E7c8OnBnIJDLQbXm2XhjIG4b7KvTh1cHqPA3F8yumfoOFhARMXMrpj4y9X2
0EliSYGHzDkuJpT/X/tnm0mQ/pJJ6/YE3fEs62vsJJbsHQf8R10/vto704q/O0CG
L4zUGGvBIzh+II1z9Pywe5JnZbqYnHtS08AwTScAuUfLmQN29ZU9GqWSozknVmgA
JA8A1djZJ+LiLAsbAIU8h9V2b8WkRdWdY+LVdKk+4QhpwAcV9bNJqOAawFd3ypwd
AedWUws6ATecQBdsgAe5WbHPLeo/1m7OgtVYr8JppcrlC/CWJP93b6GeV/ipwp4l
6gUfd4UGVGTEBmZeunpafq1Jtk96BrgII82YdHiRsZxS1C55SbbG2dHmHn3ezALg
UnUxh0BWhb5Ed8rgDnK9RxwCrwXkD6g5PfBgTc1TVc6/N07f+hThgFhFHrkOTfMu
OyGwvIvp0sc0bmzUA4XZY/8udaSJb0UGvno7vgLcivEyoE9T7mVWdtuksK5iB7dg
Hhakne+JHjpAxJyocqOI85Z31GlgLFO59QjOHRBoZkSUptlsRdSCSleY9zALK9ve
r01pR7wxlZv7rUa/J4gcaVQvEh7KUrbIcN3slqvt/ikLoshi4Y3byN2aaa79FVKG
8f8gRuba0LcZafk9BZCVfztb+xfOdMMfQttCVlLDJrqTtXWT3piEJIHjYUO9qSNN
8EObWJo6yVOVt3GLTF9FHR6rWofcbw8OmdmGk3As3qZe1ZpUQGMisy7vGeoRv96K
LCw/Dx0otj77Gr9YHItnsoxgODeGK+TVAKWB5x/TWBOlIrPXw0zy8vIkb8Snz0TM
X0bEtWgaIGWQasuk/ONCVqxO0gr7QJ8pkQcA1sxWFrQYsBfeCL/yon5V0R6OgI+b
2cq80HFYToY9UPyRtsHTn6AE9ZTLNpHiN2NPX/TIPowEtXn7Ibk419CkjnsYhKIC
IiUc7GXNt+tvMAABVjq06QxLFvIK5fMdm5hlyCKYOvI2rO6gtrln+nNQBnFgslrI
j3G7QYMnPt53WoHAXsmCrcvy/80TJBSXxIwyEoFhgr3sAe0QlCsCETETCF9dEGnX
VbodZQGhC7cRn30qfwW7s4DbdWE6nt9nEzEMzt7Q3Hqf3fv47ACGEspo+CIe6bV0
fMjXGCCByAvcfpBTLaqCpCAzndmJaQn8ERZdAySUYeli2Ocu03g5T2IKsFdS/t5p
ywf7CYlNefel792AUHsL7gfqMXmrOPteiKJMr3b1/kyhFqkNx9x3CsK9dvXv/oUX
LoSME/dSKjTo3e185DZKcijqTAv71YDmisLZhiLTP1ntgcpZ4X6Y6k1729fHX10H
uuvjWlQDokuGoUwzwoHc3o8rZJruBBnh7VJ8sCd5luN++9oEC/P0O857TymIyldV
z6exRBUSJRAZpfXrWVGPIjSmYTS0mXxJb0ca6XX2sGgx/th58Pr4RkjkDN7KC1cG
vbHbMyCgwqoDIZ77kGArVNWWQ8yrJv/1hJb7BYtvvweHpMCNu3vt8okxtdz6ydDY
qGj5qen3vePsRJEGUa+tHKxbGv4lLu921ONmYvmxQc7R7oZQVz82gUNMvoaa9I/w
OjKoZ3SVcmkKxv3gYF5yKn00aBq8SfvLU9CO4+Xnj69xRYPzUWJlOeT6/vB3/qt+
2M7OZapNiuoIXdVHuCcM3Gc7WnLuUtWkg307dTaCYXkLq1x0b98QVWTRl8cllI85
39qwND8/JmWTLJPtPzoySxQ4XH3UlD0EDye1f6UhvJ4shbcUaX65qaSlzbRBWMGf
bWtYMLP7nqkM/FEDeJQg3s1JBsABuFWNMXjWhVHxrTKnXqN9V4VCy7XJ59Jgk0o2
rpaOAn88//8CtQU3YYP3/PBo0pp9YvJjKyVqMG0PFQc1Av3ouHYLDug2rzMKhbVk
kC0GCcXf8C/BkxX8cxMMCaIg1gFCb99XD6KKMLB0bJnvtmXdu0POCs2ecvsVVIxr
Bx98tTR7ehZVs3mpfieEC4wpM7RhUqP7ud4Ls91WqUQyE86XCPI1pqmidvMCTQnE
3q7x48pvyNGip3Y/bXwKWgdSI+WPWv4nzNnulHwrrpGVi8gLw7mKKAEhD0vNYo6S
GQX/cFnmAtZQwKmnfmdzbchmDL+cM9zyvndhbMlqAHf9WI9wg5LqXAYVNSmZcgwV
zTgj6AkX1iLTLrI/28KRZ+4Wsvrfe83A5MjiwHJMzZRLMuKl4rqe1lgUQLzBzjYA
n1Ph+23T0e/2/UXQYWU6wkpZlxpa1+0Y9FKnx/IBJtBMBPdQ5SMDZqvsntviGazE
PUb5Gpzcq3d0jJdHtunD7BUfg/FrAlXD8JfS7Sq0uA64HLwzuDEP4ZC/VFz8OWuA
AqjJSqcBtYcoXEDRmjY6k7MtZYXs00bIjp7cZRT83Swyr1AwumLKdg4Np17egh30
bqg6dA8QnqwzcW6FtlUufPsLiXiqfW8jMdrP473bUblFQ3Xmp95SzQiBPHUKFYMX
8C0wpLZQanSYMxoXYhaCeW7ESnkdKWxOhciGTALwkEm9xj5kVvOXrDfZXnW/tl1m
JnYzTOHn3VkgQHZvYISpwE4kxQfRtSUf0jASSN1MwJVP95xoiIT43Z4/7ASSQc6Q
IupRNOng4QL7B0w3D+9gLu4YjMSqvNXotE3FeOluMrDI4XefQuN7v6JURZHZeJpE
9uuLNYs2XnqYmSVZO3fJxIxUTZzj3a4whoMKmc/198M377hxm8KFyTpiVjIUzKnq
nsTbUj3tcvZ+dzOBx2mhqlhnPJOKntvXuB1kbzl1u7G8wR3BBuqcgyl6huVDxiXN
sufvcvGax4/Qy3XWF7FYfDUbNiIH2dO8sJ39T9Ziqd9nqbzE1PqW46hpFyj4qxcO
UNE136pChVVtzBfbNFQgYAiCpp8bSh6FKh1ZRxb27ixjn6HG6SHXtzZAKBnU11EH
+778bO53+z+6E5A4FG6mLqMuFrlm8uvhJbJ7ktOTeNi2n2sowPQG9XNoxJ//GRdY
ROWIP2ywnYpfDiShwd6eP4aXo4nHr/E0KnbgoW41JaP/s9qACyxcw0Jd3IMzOFcS
haJpXg+6WCoYHdAjskEgLCGio8RTIZzc8IC0ov8vI4oCDBFkLTz/Qt7eDvUoGRZ/
yDHt8HKp1/rrtqvT8yY1vMInnr+qbcb259z2HNYQxsDoro03hMKSOUy0I6Ku24Gq
LEJT+4AUNr4xYsrBTZcjR9cbJgN4fR18cqRn1+kexwfXO8H0xC5+9NAW2RbxcW+e
vZSxEl5Mnob+nxI2rF50WaeBDGAmIYAsNVAUdOLxX2AYDVeIt+n2DGexoNRpmIZb
RD8Y5v7dkz4+QAVs/qhablU8vRV/80ohZLCeGjz22HXRDfD5u6iaCdkmjW5DHVf1
TLo3cnGmNPBQWvjZkWX2Enpe9IlyEfhwbDTmv1cubwBPxNwucqxCRw3h6Xd70Y0s
g0L/4cmDzRciZv2Koll+xPU+wqndRxvlRsMIw0zco/Ds4oYbpgiIj+L/fb2EQRcR
a8B9Gl584Tnxs0XDfE7THOrvtAm2o/SEB9rXvox1RLDYRfoshtjiLb0xewWnmuOh
9SR7hrYRHCUIIyAXYBeDGv1HDg0QVt4Nk6b+7h53q3UP3/GKgirM38aNmx/6O+sB
sJZ1u4TfZXztSGtA4bg1WXj9gXob8AI1d2O1LbVD8hLCMlzd5+6YMd/4nUNVH2ZT
PbbTSLsY7h+UclkZtGeMrb1RO4bGqqmg6+LmA2000U6MbSjW8wOeQseEnqJtb7B5
cV+2s+g4PdWDPfV2r2cpOUvVcp39q/9HJXkJJs0zkBDKM/iDV5CPVEuyFZVVvUJa
DgzKJQReMbZk7MpFLzUxBY99j1sQMYjlR+MH+5F6KL96KQn4et7PbjD0Pco8J8sR
lzAkOwglFRsFIy6BkVXog8ksefLiCAkDT60hyI5L7XQex0yv6kOArWK44Z0MQIXl
vWnOYX7Sp3DYcPG/95H95gX1PpEcRaNNoSh/ImXyPLc/btxpRSBSuKz0sSTt1VbM
lDdaTRgeeeAN0F8qTwNsAmrw7ZchMDDnNJdgz8jhv1gOKWos/zccisdEJBfzllPc
GxdXN39DE4sxWf+7Fxj7/N/6vTeFjQhIgNe3z50TVKcmJqpOSsPulOvxZ0YEY0KY
+zz7pVvwZ2eQ+yMtgL5H7eeHYE9um8v9+EuN06KYVeD7WlIGfWDjq6d/dTU8h7QT
U6+blutCU3XS6tkqg7TQxeUmDZ3kcNBCU0eoEOFnCp0SP1BJOAI5Dcf8YOXNXGcq
vmp0Ol5hqZ8qVAeSvc71uapyRBe3hLNM0lQBl8pyLUW4tLG/gOUkWUMmylpDD1nt
/XXpSzvX2RudcNy/5g4N4t2lQSAGjvAJIZTBkOahDiaoiks2yVcloCxymIJAVyY7
WL6PuMzGrWQMIWS0tJLX8sWrf6C2IeHyVrQGj+SSDt/ESQMOkPOQDdrlsN2xfNOL
2WqUGpAhndvsm31/QHKqJ4RiF7n7dVjQPeu7QyFhVi1JkUWF6OYUu19HGfhdFhwr
e6U04vrVEigw28as+WpSgBeBImbCEkRks7JdohkvBZ1jrtIRh2VB0bFd7LpTgS3d
Htq4f4YCucT1EAYcfBg2LqlBaTTWhAtfmEo5833a6tcIx4lplHtNtlicRIUNn0cn
6ja6PGkkghsT0IV3ADHoIH5SjXijbJcUTMiRJHXUXD78PQ2oYgmP5XPre5byvSH5
BskzcxU83qEwRYqrbhsprMjWBQ+XSi8uU81BtIHBry2v2VsfgrcWFXYmonFiJPWr
UwGRfN+VMuziM2hSL1rd0Woy2jduOKH12dpPXGn4kzaQ3IMmdj+CmJM2PrwSGZge
Mjn8Si58Q4rb+slCVBKWsPxzN3O4Rd/IvXCrkLkQNtt/6f+IMBwUqT+QWpPgACsZ
6CIs6lGWNXrLWeOhTGgnz/2KAjIMKro7YGjRGMLBmOWLBdGXxg8ZfYYuETFRvZgS
xUmAZgE3onbgTW2oQjrzxtsTTassq24NAGEjoFi1uedkogDEDdE8KYI6RktTynOx
zw7Law7Hq8tPQapbT1xUWdTB7E7nvvKRynn6/h8y3sAcjjCfJMtf7ta4WBpF1C3n
0tqmssU2sfwotRm3iizzfx9LD2d55vHEViC0l2enyZXZ2N3dKqyBh3QOn1L5ujWZ
yes74bbJCMhS8B6R3hUbQqkxxFqYLRFzAbyBguI+URvauvuk7iVmXpYm370Ib8Mf
Q1oojYMlIOB31oBFfUbaK7a9pB5tD1GzpyXpQU0DQrMhIYhfC2SFM5E2eiu7bqJu
Yd4vZnfjYtbWgi+vn11HRH7VRERcYMZUyIkHzYlhvuCuekf2+IN4GxYHl9gpBiBz
P08qlMDW3oD5Y3u71b7EFmk0VbIpW214UmM4e7IkIcRgO9uNxRhIiwfZm6pWf/b3
ADc9NztkVX7JCSDv/5vCY66NwiTMx7lZeVqNJe8ZqsZtfDD+CpFHgZ+1FCP7+mHo
3fr0rWNB32wYVD/lAMyeG4viqd3RUg1czJOsEyrG/MPPCb+uz1E+jI1qiDBRkvff
Nl+LB2Ot/9IUOlPoxFmLoJUT/Oc/6QNlAr+fAV8rRu1FA+jJzIKeLKtfupohaRNj
bufGDQHm5lDvH30UsdDozR5ozHe2nl0h0SbmuBNWn1MY3aq++e5kIwDGG6XBo0e1
Zsfe5Noa1kj4P+Zl9VTa9LXMqbuneUQd5CAuEnHKfaQilXg/QNobfwvE6qB5Z1s2
RjCw3L9QeWrqYelFxxQZXX1FaAPtvdi2M7tJ1OlnlWqkCqeDYa2oiRW+9O0DmdHr
nnAI6ym+baAcjsPFHDe9f6I3c1YWUgG1jxwO7Y5h9vuNQq7iwNZOzdUs4aBHKf9p
HzqfEUUoFuuJxt0Tf+HPLfG3DF924N3UdJDCybmlcaUhYq8oZg/H+FlJGeVdlp1f
9Ztt7hh36zXaiOx8CwkNb5WEPAk4DM1Cvm7XB3M1iAr1Q00MHCemoIg+hTNpKfwk
b9jstM8caCy647w9BRyp8/BXfWUM985nNvttx55b0Dq5XuCwIp40KsLYYaAh5NG6
TUVFs6fr/2Ssm2Tt9KTXHXcmYC9AES+F4StKYZSO6sVjQjSw9vd9oKTtqf0g5H/0
LE2yrMOXsYSzo4yxJ4GQsK1iS6vEM/5h26eVy7wyVs2ooclH9zSMYmEzcUCu+qOb
cbs1XBpUoejdC0CMXzwsALUI3g9ZfMcsvS4Yu+bF2oOW0CFh5+P/yEO8b6+rm7ET
ec1kPXemsjJdP2oiEPG5l/X7VGvLYDuVLgCxNJJBy2Ql+vnKuieiYOLAuzPqchTt
jzENlDns4IKyxiy6+UKbOqE1DrLgVH98fq6rBMG+vnvualRVSb6HtKSM+eZBRJAC
0L+X5AWkNV3pvFpeFWyeM2AhyXrhcESXnFi8++D5DGPahLOFL3xsMiRymXkg5jBG
v4jsku+JEQBa8TVPUSfqUuEyeq+7v5JZeLdYDUbC6xZIEGlwyqV0RFRNLlZS82bu
u+hCEEB99klnDc+pYZgX89n7sFY4DldHyMK5JRBeDfpTP6qjgD68nh2O0n8vz8zY
X4pvZ28L/Xb1IUuDicF/6p4LwUnW35GoNWE3j0iipe2tknx2uF5VADA2QsjKABwQ
bNhLUtdDsa7/qD+1PJV8YBVHlcHd9tg/ZyJOjjXEpCdVklz2EN81Qcm+D1lOrArN
61lBaiyVrbES40DUhiKOLbl+inbuDa/oCpY0yTZs8ZAWmdiXPOCsEvfAZ+kZJ6N+
cPS1tONvjp6yE7IE3jaTvtmKayogULEKyCREVZfmA1vPVs1WOpwK1+A+6am003nt
kZBfe4FdApNg8Cjm6WtlJBZQpwD9/6rVxVIMIkOvgt2ooLWq3YkEqeBnknU7ZISx
2PPuTOVvCwSniU28IasGg+2SEZu7qGN74Ij4uLhqROeyxwmLQkiBJfrtrvCa3MaD
I0+OuZBYioRFwQRN3QaE2yZRF17ii9Cc/auvqlJYHnGiwx+amtLWa5UlyZKnnb7/
TjMKNhs0ON4YrH9mzGV4JOQn/H5L0608NWwuTyQpAn3UfSLVDwneEG26Ywvm7qgl
Qg9Tk8jZ9IzzCxE3H8t5nb8gYWNEjwu+mKP6nsmoFVzQLDgKaW/ItnATilOYuPGU
16QcjUW6cqJs91d2OjkCFVOeeW4+dIJ7WDesI4BhAZ82qzmIhV2+mRBeXhE3hfAT
2GGKe6hcuQ9eL5fOqYe0B+9RBEqO43aFeFhDbtsJ1mf/m8lKypi3TrjBqT2YVqFP
ob6aY4nLkB4X7sxTAfEVooagpqCjeWvo72knn3kCPeQqmnuQ4aycwKPfTJSK1DJ2
Ppj97ytNjmMJ0mGISkj4pNqZUJ+ucIlCTErtMdAO/tmXUhWmwLNe2NsyotXPJ2f4
DNB/xnnpCe62JbGx9vJ5fn0a7jf8w4s8EH6P3gicFzw2r3ecR9w6R9K+chg66KvG
8DwDsXzt3qXkb4LJP/LAK8cYmfdUPqQpX0iXe1GLeVoTgpM2fhtoiMrSB+pA4Qj4
vZrYOfv0rBvfiZQle/LWbK+STmIoyXu+Ro2krPoc3NL+dqyngabUJ67HmbrizRyu
MFXFX9IMs1irP9XKa/eS4l6Mas0TEZqaIuL7rBxEPO6jZx4P5rM27jZR2h//Vv1m
IVtS1tUBhw+BNiNfurF0uCQd4SGiy7a/J3h/5WOmB+XjuSyTt1TqVgQLXwxa6PXq
Dz+ohNoW2t3BiJKnGrSQZMbjA4B6HTXkv1basrBxCfY7uHJIoSt5wOFoP1NSOC7N
9I6SSydLmd3ilFbNFqApgLFXoMvKNXQX/8OxLlX3JHL2s1zycW0DMNyCTsed4Yr2
PNKlND4nEVX3pkPv4I5ouMa+vyvUBtIZhLnHXDK3j+RTvuBXGTkT4pmww87JtNar
d91K49+PqhtEHrtgls3JzlwaUcN1tAwyDqb3wurTFq3sJYSqcQqFOYviEinbMPPH
GpIrQvWmF5Y19oBYi6V14+hP7uPU6gZM29rVALwHZiLheuH87qIwF+LKLHwKIgSF
IBVU25gqhFmJlaVB6y4Lla64bDfc3iuD5uMBHeGUSQb/ICzCmMX+2ebwy50BhpSK
MH4SnCFosVGaiZt4ZR4JPTpu3M5Ht2j6i0g54BH13/b1ZWK5J5K8K7IvEhmAD2Yp
s1XT7/ar4Fk4RTOmyKL6trExIuVLnat9xQ+J474MC7pBYtqyny+cAwvmUcgYi5eE
YGM1XNDPdX/45XZD7wBML8dgY3xWidlU/mhI4bzhq9iCa2k8lcEdzLgFel0c2Iij
G7kTW8C+mhNGLyw9L/iZbTkF72aUZRlIxtAvZC6nJ8/TJQLp9C0FPl6RzgDCf95F
VzfPzxT/EhMa42RibWm7KW0zq6s8T7gRv53TPPkDXaLPhA4p+xALtfFFgYCHGfiy
6UPYs+DR/RUdoSMVZSmFHSHPUgz1l3+6Xu95ASL5lg5+DFG1rFyivH+XtWPj4phk
y6x3nymqfRi92m6SImu4j/h7Y6Mx2QTE4/sr+DMSUVFePF9mx/izR+Ve/+nz4wTm
PLPMfXwRrPKJ49F9hHpHSOlioBie37oTI3ViosWoLagHVqIofZ449AtrXPdpmJ2k
X9A5AY+zg7Sgrkhp+vB8BpdXpyio5msLftnpkvKsUYucmtcbWh1dhShgnL2lhTbg
CQwVKXQyotL+eOnnjSai0zom8934ZEXSeX3s87QIZkutAy1JdhUy53PK2pJc4IW9
ywq2YgQmiInZ4J1osnEsMKXKRXWKOYCHSmP6v9YuBiZyGrvwPFwQjwG2wBWAg8o3
dPrafo0Tw0Y6O8g+PPcJaTKPHgVJwV1I2BIGxq2Zs20PUT+RhselwdHqG6Ih6ulI
ZOJQa7tUVtXYBv4WI6Gu1Yhj6Advi496vGtnBJ6Ln5f3WdNH2Nvz1isO/XcqUQlu
8ZWCZjRxOSR9XA5duarLJoBmiRfRi5k4Ficx6bi2ckiUeqkHbq+xAlc9Cd9lC24v
qwSEVmJs4gn+Uv3n1pvAiN9n6AyPSkekxMhuBO/6V3NWTFWZvpmhtfg/9xiKeZ1H
LRnwUfLsAa17oCevegRnqdNrpLv8+zaTRuBoRamooHor9qhTDPm4ct8OrocYjDcX
UjXRraz2b/p7XNhVkWWG3Tcf3S0pTDA2r+wdCpmhVH6799ca9hrSqnefN2NlVqqA
TXgsbV32r5lAFH/eBAatgp6sOYESdxLFI9I0HI/96TFcv4njrbmaMEoop9DqKz1/
/O/vZG9Cb8Wa95Bcp7vaCJz0HIxFA4+8gpP1MpkaXQGyMP7tNXHlSD4dVOV4SOsm
LT5ylsWfGPckGWpgyPvAbx+Qbx+7zw+dMfRxhIck2sBwExccZgw6pXfKCv1AWFgB
OnsdLUJ5G2yyFYpUaEKMgt9U/FwDJaRIuHtk5aZ56pK5sNfJO5EnaWKS0yG2TNdy
aXpYLeC7tQnV6Yi2ljQUps7/RTa+8+REKD81UzVVab63elJNKjzqGSsOVq9UqfEw
r5EveQl2Pzk8t7HVcddUTX/Qbm8JskY+kblobEDi1PU19BcfcyXVRuzqJZXcLdqr
6Pee6jsSf1vSRxH/jV2OACbXMBF71yHQ6d+LiI12PB1l6OMof3MYDqODMZVsZcYi
fUZ4VvFk+8VVwiyR7hg2TJm8ypN5ApdeMer/5vVmNFW4nCnyYMLEaCNY4pgnT/ww
oThfPBxwZzSLpUtuCks+feo1rp6bsOggUbVePRDVT8XjFrtYSZmXPpW3XIPKqzRM
E2vfTTXufA4oRhxbflbIa+Mwou7Qpi0KBVgB5GzITr1PxxwXfjDvuQ0v2rFo8sJw
Eh5+hgdatNxAI+q3o9m4QM2j1ArMDDlrUa53yM0TuZmMkfufhdS7MDkQwT/p9Zlc
RSJUm5LssDmyPM/u8h1mx4fgKGcJGCsaot9H/MS19SQL0Na/HxJPMqdjqNEWm8yR
6naj4p/oibRzfswsW4RCVNnN00kUf0c+JpV4j/jSBFZnPs4ztSs1IyYe0BtBYkk7
K+7fF9L4Nn1jYWgjApirwlExWqkjRXkLnBp2kHDeQrnosGBl4esgPFUfkaKPp6M1
RAOeZgLVnW1KwYdXpKd4rED90oNbswEwYDzxDucaIIRgu0mYMXL/hpBcMvzKFgjs
XGQALjYgLVO3CgLiQVAktpoA62Qy5jDTyU3qS7NiqrXOFIrNcwO9km0FmyoEtkXo
6MQGMjgJVKc/b/JyRBjZKu9JY9SrTWCNAVg/VlsWOjCWyF5gGBDnZ3O6ILKPY9IY
y1dQBB/S5zUnfl5cq9/C0XKZVrkq0cskWmcYV3gJQNHqBh3PfFbMOYpemKRUp9il
u/Zmn40fNjUWRO7o5mNGljtiJqa/lS9imVjGR+V694EdlnycK6qtGyS811HE+tTw
tdd+xzNYAL7b2FniiJGCYwjH+Z6Ed+Ryb5jD7jlhKTlddrx2UESQ4YXPCrEHRvnI
z9FP++WJJsWPzRSwUSMieMqq7YXTuArgYe0zH4cb26wiho4AKv+KsvVjwhZ3fh03
BoKeoc2oo0krwquZ2WiQyweDdbqVa3WmZQJleI5oJo0aTzp0ehCOCO9Q29c4sahL
dRwWKxzAzyIJfiMzv5ATAfhA1nEhWlNeb6rZAGb7+bsu+M3vMWgiQcPS3J4riUbY
PeSP6Qtr80laUAoqDJZEgFIwhL4wQBvl/Qt73W0B+SixK87/nkQC7C3PCqm5tg7j
Lg+987weNbx8mNJdDB3P3tbWmhXvgWJTVVHx1ODyzkBTDBLlkJAFgMbJNiZDqHgS
5hB3hEb5VpZzHwZuloUsNY9oFdyOrWYBEGh1X4jbqkQwO6Dy90B/p53tzkvcfkoR
OpnJVdwkWeqZlG2+Fv+QipGlBvz1pk+L+MAulh/91rx2BefvSDUR0YTxExdIx7JN
HOHTHjgRz0hkH4SXRjYL9O41HQLUEH37UfCu7qJZUVIhNp1OON9wUfOVj/du8rIt
AzQyBt95WCn9vMyo61ddUtnfPe+DiKEXhWpDClP8Vp+XnLDhqhF0P1gEob5sGH52
Jbqd935o7tTi1D/TAEhR9dAXcqifskwovedZOaXkaKXuGfyemgW8MOtrxUprQxyT
j0sJFsZRvePcl1Du78OUuFVqE+jKodf5j3AggQrXf9K9uESAIKtzB/IFrpygd5Dr
6Zm8uQhc+n88xLu851Fb7cmKGIoRvZ6mTY7EolHqjLXo1TDUAxahYF711LZrs0vc
ScE1Hr7VISmBY62Z507cuYYju+48/ktb7tNYG4UcwSSgH59QE3qefjfjNRmGD5Go
RDDZ1DRDC86R4qWAyqhNbrLQb9do5+ifKiua8OrKicG+vTa6VfIRhQsJVhQf/30B
t8Q9PGkYPLRA9OYiRpMSign6uSHlt2XAbcbKgQnbkCPfuoVh9gKXuNvFpwiwyIKF
uODHmAO3qTwIITJo2BbyZNkthLs4DOqOs2GP1pkbKFv0E0dih8id/99leR8aYNAB
PMN3IkPBC2KvBgsKn/N92x1FWkrwysvIxe1S/n5pRqiR7WymSVFTCBkKjAk6N8mI
vzqp+J+llJVTeMmii7S4VYAldasnihIodib8wk/RS81k7dBclAuM7M2se1aZSgEf
F8d3NnYzyjsOh3tTvLC7cv8LeBenei+Rif4Ns9J8T86ley+3d749pv3M2hvgZXy6
MqPbsq0wh7Vs2JP5kT4BCUwV2KBPRmlt61XZNSRZTTvBgmZN3NV+2xa/ADWc9LQA
7+s8MGIyu66mvAWUyXwUxpLgCmyv33gTi2cp/RifH8y/Sh7SWZ2F/y5iYDRqQPmW
hE0qoMz+bFut9qkTM/Qp0chL2Ip9KZAXVE48ald2u2jNRzvRdlVKnKpCB59Q9+m8
Dy2KNHyQCPEj6hyTCluLKZf5OT9hgOazEZxjPORNBXA7nAmXWCaj2VHRNLixTK8m
BYYD0M6JASLnIJp0Tm9+AeKOFSFG+yCu5YwOtiuHq0Im4bzSiEbKudaFwncN8tqb
1KZVC/s1Q4IS8iHK7QCgjXmi09+hngNxEwq6T0gTcELjhEDe0ktR0HHjYDYZOGN9
vD9nHAXuIlgzJUR42crvDCpvc8oRXYAA2YlehKD4TnsI6BBugdWi437woLtZRLHu
dcBcGvznhl2U+5s7E4eLoCKhtbzWoGj+Hut6dQ0/Nm/vTpTeZLLHIHaaSAngKZ8O
KtZ0m5r/Q/8ojS6+ABEIT8rJBH6B77kmjm4g5nEub293ce7GWYpMYqV9POY/lCMj
k58aKVj9WliPcRK57sAkGUYfeAaiA8YYxAsArN5NPreTLueHE1KFXupFMonMSti5
8LJGdIaQ4vBepxNrdw//g645w+KbR+Fq6pQbd8jTh66XHNJBJ3LtC+3njKzlrjxB
C6ob0clQqw0P90Z+uYVACvOxfLoa/42uL7uRhuaseH8QubiWW6Wf91fCoTc5PL5V
CYXZPaY7cKPDNzCZFmMi8WCc/mbg0kue0gGt5VmM9tVjSLTZ8ZoRWx8a0sFTI7e9
Zho4eWWZ1bWSGkT6cOExXSPuR2nq4f8JKlFhgfWjKHdGQQEhkcBc7N9FInFAC3jJ
e3s6vJBJFlt0YNUEEmox+SYc3qR1MBMifjTJwIVex9d9UcLLJ5C2SVDxPnwvWVG8
+x2WSxzMYYG4tvPtXD02aQez6hounF7HsB3zIN18ZYPe5TRz2VVfmWIanUzXdKOl
LYbsR9eed0wtjcaIL7YIn7U1lPjQLpU2/yECmCYnbz4il53oQdgbICSK4bZlWi3i
cX+y81E1CKb6eTEZiXzkI7ptoGmJn18L/Z6op0RaPhSFD1JiP+xtRsFig8qqizfR
FL/LVpCLBbRr+bkAfNW+xZlSwzm7dADMIxN6RlI1zDHvXXIHTKUdc1UHMTeus0dD
GfdyAQPtmVir3g5a8jV29c+SiwyhQdrCXlXTFE2IsNjsXEnVkdUWWqXPmf9suN/v
eUFIZzHAeMa2zYd+pHt3RdGPLKRKFDcnvD1cuWZKyVoGJh7ObVI9iDjOhtbXlYdf
YNpBAoTUXUuy36DjAiB7MxzXYA8oo4xq5NVquz27BGb6sGthSEM/JMz0vBfQX13X
5B/V0kRH8HbG6M+QxaXNwp0Hr5mNJDFGJmNdo7J80hH3fOMPFzRrj5uh9KyQnFl/
Nm4dZiIRggC0oU+AmjTKkek5tn0Jq7nE8VasTAgRYrUb7YyTHi/CAiJ120IgfwWk
ynQoGmYG9r7ufNMf9BG/tgyLagfapHi0h/0jxYWK17iABdBwu5LbpThmJj1km7bk
UYwdYM78lP2PCbe8k5+jFNcyoSsv63Sfkzx7iZWWNeOvRbmYFd5FGiGGq+NKsiby
ZVtgRp44kjQKHMVLia8bvJ4MEXqBUcM6I6MhEARCDSKIs68l5jT6tSHto40iAnwd
TOIVlp0HGdC0RTKNrXO3kxtAlHevdGilI3q4mVW6jIwETR8mm7RH85YUg6RJAoF5
8XRxCSDXkkZBgTvtANFTIq8ImRdUHoTUkNznYLirfeHq54AlSVNKq/uF/qG4mCYL
/y2m9q/Vji42Cz3x8erdV4VwwoiGtbV0IsvOX9IrkYOPh+GLscxOxQ/EgqvI1Lhd
hwsbxlzFrLDDXfg0MuyYsm2Pf61EOxugOnNIUO7slYX4J1xWWzXbYzCC95hBJw2A
VqmkbVuPWovh1j7ngvLwQC4kBs7WlFt6Tk8Jn6ohMOUEj+2yJGhei+zonP0yfhQd
HS3IBT7UFAcbijImJ5W/+sI57pasYpzWgPnWDhk7g9H+2KNNQeRo3+70CnFqZ3Zm
yu3dfGjzL197b2hiIN+FxP7ioLzGVRntYh9FYF6HNazFE2ajYFlSS9KVcVdy4K1e
jNskCCQNXz3QFfhBaYj9VLge0J2+R6wa6pJjXUltQSmLzXfWFE8HEoBVLDXj0mLJ
Bxah3Gil9D7J4hUu/H3tnNFmUZps8RjiqOyNYMKYaFncp+NLOUl312tJl+j5gdlG
f7xupFOrRuMudO1u5kEpnvPLqecPm0ZxSgzFSO1NiXZfcMzBtVWpQsdrigSe7k4r
VlvYGpYcqsjSB7scIQJ0ExSps74Krd8og8cJ3iqrdlsFwmhuVZW191lJKhGVJj82
x7viRxZRKH+IZUc22JNWDSgWUJjw61tHd6AjGkSTEz8qF8OHCH92J5Bdi4aydKsZ
YBAXU90hsQJLvYhZEIWBq7+wNnll9J8gEi1vE82eaS0qdtMkVOweLjP3n85LTIsR
W4AEC2pCz6rnPrxH8IKKZUerEl3Zg6s9e/lP+ORY8o8BLh+YtVpXxq84rItREQep
O5JNcX8O7XjZ7dBJCyH8xihgBmnwHsuJBPMM1Gi6N7+DqdX+a+2VbIDWjsrVSMvS
YahlpeHVHNVwztHJxdBdtyFJ1LZ57vWhBzJpwVPeIA50ggYwItm1lGpWcDandKuB
EKS8W5EJDG4okLjF+kGQZ68Ri0tc6LgXZaAoqeZWJfpd4X941rT32ZUZJeyZ/CwA
lVeEWqgeRLvNgTyI/X+MUcHs2391gsXW9dEAjgRmoB7gyaEBFaINLN1BJ/mpd/Od
ERtMHn9XJzU7mxBu2rnV1VoCxhUQA3y65+MYnL8ca1+bsaFGhj6J/NECuR92xOR8
o03+3cSow3pn/YmWlTfj3/4WG40t99L/ZbGirw9YhmAd/0BiMWursACnGc36jvSS
R7ZNxUzCUynEq0CqfiSHFqwlwreKVor1rZwnkvRolR8PlBfRePFrFchOpJkhUNui
+E6LY2rKlZGrb+18HVT6GU2M2oCSRWCWRTPNrUQvX48qqL5q4WwA6720+QMw58AU
1D+HuVMPX5Cpq8p8db7F710ZjeeAqW9vvS+VeMfVtwzwvUUzc/8MlhJkl+s/DJ8t
ij74qmGa+0KnB7k/0qNmr5cekbafcwxzYsxvOd5AhIabv0WKrO7eXPzkRJORHrd1
V1wfA1xUE5tBxMfBYwyaTYH+nn6/2oud4nYs5iT7+RpnPXgCoGlRM4u80+X5JWo9
OVtbWv2ErsONhUGSWMvN2vhTmBZGo+9bz4NXWJDWMnpT4lhvjdLZxlAjFNlb5bEu
RUYe0Ly1nNBB3Bs3+nnhWFIvB+oEGacE7V3IwWIg7i8br4SLAmGzIcChQ/ZPN9Tw
Vbx98fJspN5uORVmzsSKhhmlQyx9r8hVdB3TMwJc1g7xy7P/25/MW+J19Crxe0kI
jIyhtl7tla7XNNlPyOi6YMt7bbapnFO9e3ePXgTiMZbFVrjFoUPeevuzCZ9kBu1H
keQeLDrixx9P14/cizmzijzCeSWlpI7XN/+Ae36pIwOy9GPGHK/ZEvzJD7PbHyBC
b2kw8IpV7/jt2gQTxo2N0UUoYTpblwjIMPasH1BIlNd6EwlcmI3CQecAq/3ZmMJ5
qZky9jdBKh9lFsQ6C2e3vdwfYtXCsEFbLs9iQfhYPPD2UzkH+qgyCyAVMQBzkyue
ROLDNG9EmXNE/BTSnCqUSMVrjF6wy531z304pPxeGZ2zc/Crq5Tsf284V+eDXJxJ
Tk76XMK5snTHFDBlnzocndV1pZ+CbFInOK5xS+VIHGoPH5QwDI+ak4A0IMvaZ0y6
7pa2D7CmTXRpDCL41X+hMAhFlnyXzJrlGsMEr1VfdotP2iGwF7O5fdEFogABzRjM
v3AbS8psbpMNeQCAeeVjojutH7GhSf73gwBS8B03P/DoGV2LLVaLzaJ6LEdtkIPo
PfkXK1hxzdf0miulFDCAFHze6OqGZPYV/MX18lfADuk109JHZOIw02LI/9MuUcvW
X0KWpF6OkI/YNk98c6Yj02pfFXH5AYLpioU5U4nJIINRQWej9EiisL2Hyz2LK7Pe
iDPPq4BwMCCO0YA/jOF7MMR20CEQTBDJtkhsZpSu065JeZ5CiLRGd6JralBH3p3G
bQ9P94lju82eY/qbO0OEqDOKNJ+uYm1x1XIjrOKmbG6PicbQVImhh3JDEEmXvlhr
owEsC9nTrTFdUvNSzDc94qpi/vKzaOZobNp1TttLkGGU6d3+1PNX2VvrE8+x8u6l
kKvHJ3Db5I5425oUXIaCVI+ACETwnWj8mXQ6k9QnmO5FFTNrJOhuc8b+pgThSb76
KUpc/8O1vJYDT4ifySRSEYC7E+63lI1+NNfvZMT9rIuK+CLd5MZ4TEKBp5clOmeo
UiiDq50LPqrUa+Ogo9kC6nABsWugOK6JsvRBvXjRAoibPCaZ3b0bl2FgO8fOacbW
Ogp93MGhmPQ/TpHVswl91T6ZanPB1fZRrvZN7z7MEzc9TylYHxDvWj7063VV/ti/
vRXktnHaMjVQBcaLWeMZlx3jVHpAv9N1xYrNEz48RHwumbY93J06XWeQOOwxSP6s
gGYflQAO90P+SuP4LzEmrsqQHfs4NyLHpZ93iP33chguUaXvlPU/tlb8D13BaHox
LpDXAhXXUDNF33e6q6aHo1re3WvLvpxzxkpJioQJqRGKXEffh2sazpcPOaQOVvAZ
q7wvlmAZVs3+YxPHhCZJ4Wl4zLEuseAzQATt9AcwMwGoa8fFcqaV2r4CsnDcZZEg
RskiU4JaBhODpB7JPDjbmjNi/jZjmfnVWjWqMWksg4gn32guuQ5j+9i7VuYZy3mx
FcFMEhvs3UOzkSg9PTbraM3YpMgwWBIQDPKBrib4SGT8PcZm1099Z8B7WFAfPPi5
DWo2fopbo4n9g6SjJixkLTUn5bZGhLPm4K/SLkC09sTtJpHVwAPM2K3IXBcC303w
rbqfmfzYbkYdfWtqCPdDrpnHEyguvh80IZNFmsZSUb2rneJSQOf8xBm4j9EUns42
cVBzqKFBXPY7pX2zl6btiW7R0hu8YDj30h9MJCCDNB8cJVDCzYmHj+MB6S6LID5S
dCTipWYx1en/yoEvGH8/JEoOveD+DBBmXZ2YBv7ZGbMfnQtq3zb38Y2ixmJO8sPs
6pQbaUkPjdYk/5457DPyZnk4Y3m31cj1QjTX1eiYOY7xP5JywOaLN8Am7mvHNu5e
+XQomtv4BQDcKwOT+DtXeGJBQ0ww3Yzus800Ly8MLlrWzVih5gvvblMuH7jXBhEJ
lzIiCxufIdBH/RVHcVcmAzotmfjEbE4NbVeTqjQ8e42SuIMq8LxEyRuK1y5r5wVW
FFd3FDKIVABVry53LYL1VXyJ/xCXtcFTA4vFp6JPjYm/AalAWCco3VJnOmhHgg8G
+wCwT4iUWFjOWLVTGg6L6gubzuHc1F2/UMSrn5/2qKdWTsWUEbGnPC9jLKis9yDL
/ZzNI+53wza+uIBv/IGo+q2AfAK60zq5GHwS8czCKMGUcqf1o/honlECunqpEbY2
wCCBOVeC1O3cqLCXm4GJngv0KzLVQGYItHIbiv0/gUIBb0r55HHRtPdHhf6FPeZZ
mJbh80UZA0jG3NYs9LYK+OIWERnBEpJN6tH2gO0QQbRhhke/VI9oxyY/7+9JIueT
IO9IFsktW0VIXXFqjc1U39Gtt4/es0oOJr7uclrKDcfnqYLoVSzPx6ge/8G6dfKn
+dIQ+vi3xy2urCOBu7AOvL9NQ8rPlEDXnvl1kr8ByteX0WnDzAJXC8+PSGmagrLr
weAt5ZJ+SyCCTmN/uCan48IHxNiWIymZ1BfhZC792JlcakOHHvLg4girVdOOg/sD
oabp02C9wYHUoWBPvGfMcXEmo7oYPH/8tn8Y65kxLL8Uthjyi5X43cz2pcL3IuQL
KRNV8pSCQfwy9riofhHGIXrtFvkV4xDflHxP1cv8IJNTP41r/+EaCVJVOWEt8qDV
UOzBys4KqLku5PBb7naUA/HdWzBIbxRR4TdY0vAnh7nhgPCqHgchNFQ+aRUKRpY+
D/4rlNHID+nCPbtm5iCyVQ6+b4U40Bp8hNEPivcz0e+Nt7bj+uRGG2DEg30io7iO
cHK8EVb5fNKQgtBh2zRBSduQ78UU9WEaE9asEo8/cu/m7FTlb+47851Q5SUAzCE/
yL+cvM7Gx7V1cY0roiGnGycZ4htnXo6yh74o42h321Wt0jD3VJXY3Cmm4bLmhZMY
+67eMAxEwADzte9B1VlWQwPTXythIwyV6rx3DdlpunjOJNwDqYIQaZi9KuL6fC9w
kH+GzIWFDPNAELUx3Qg79RRDkLtw/1j2Q8ZNn8E1KuWOx+CN9WGeEPmtK/T/zH+a
LNhNaN5+gZ1GHFMV9ZJYlwaYPntWs6Ll9wFkHNmVL7jjZBLS9WKE2ZJvqQU28D4F
rpc69OV00V8UftFR5g5zQBNxCzVhEYg3WZizGEf4gSH9E+bIROtNyPk3CphnCQDx
//lYsFAwihA9L7KIfXWBTLCYGpqtLZ+clugkOqjw6i55GEP7jgxB/XrWzcxPHeS2
xRM9bLa3+OiiwSuT0Yh4yKP7q7Vo0IAxRVbUkJHJ9LALMnAOMRV3X060xL+3Gj07
FNmxOfasOFEW80ANGyTCLvZMVjH53wdGRci0wZs6a+SXNwOvWCzfKcxAvAXK52xZ
vJQ2mMPGae1KI+4LB5HVBjmzD6CbtSAwPw6FxpjKBIVtXD9pFEeaAMpCxr/tEfx2
MOwXUStUI/Tna3kUFM9j9ke3iNIgfMzKxXO5Gj4vCvI2dsR8eo8W3tF66r1/a/RT
dqUOucoPhmNvf4X7PePyJX9PJIikGOs5B24BZmCKed2Oe1qMq2LIXyo1Fn3UTnpm
ihHp0e13qjyf2KpyYaEKHJAzTveVZNhYwriYcBGGeD9laa55vbiKGj7nKPE8mqGJ
SZ08vKiau6TpEu9sEcevDBherf2CkDGel1j27f1mLDOcLmJnJ2OGF41Fsir8fWoK
p7hpvXF5ZDBE/OGSgVBetVozQyirY31Po0wnhQsbiNwALIcsYLZlzwlCXC3AxKFb
ZeH5VCPYrEKuS8XWSnr4xRkAEpiiLorC12MLAIKMIdTNI7WqVPDq0ZyUVDaMBOiI
+PoqPftimvKoIQoEompruq5adWu+BmhSND1/tt36jS+W50WM/sumxpGLM7ZMfWXU
URuOZ7WhZU7+oqbhaqm8OngTeY9571rDjyLVwAPEBooIRChRCm7/dQfDjA+dbZn1
noxcPIr+69BIMXuQUFtIGPq9yz24Nbz5XEDWLUBBJ27ql8ZKkxHdj6jja3EnPHU5
mLhZamHUIIapePdimwX5dG20DmuZRqHZm/4skjo/9Bsn4frC/Uu5JAtwknuFphIg
qakZWXUa71zI00BCGnNh4/1oNnKq5mGVWqPe42Mkux5Ey/2rv1tmhHzJYeMPDBcT
Mt/+x6uaTCf14Ts5Hj/E1sD6VG6TCtfspPlzdDzeV50x0Rscj5Y1QJ/dX975Zc4a
15wqbF2KpTNMobC8LNXVM6854U+yqpdwVsZmJHZ2xPalV6ORL33zCQVLWORvHrz6
u4rh4UL9aQqmetma+3NgINo3whHdJO6ZE6nBg4xvvKhfUDRAIZ2uZbM8SK+Ie9Ns
3HXWpNzPbaaZCRmDhmJ5qFxRLHhFmXYRl5H4kC5nBnJ2oVZRdkKR4J4NvoBDoHbu
53UNYlvuu4TFUMIwyh5O2eYu/TKHQratfEM93O+hQyKS9v4PSnzyGoskes0fDN9k
wbV+A1+3oWXmRi5xxXuDwll060IWbYNvp+hE3QZz3SCt9uT7FbFFokcCk1gEHVmo
eHwk8AlXaMAvI3zukSRBtDqL1PWvGnlahMlcq/q4WXuw/IzFil05RCX5wgB00/i1
xJsgusmxwcBVFDE4o7w5yEp/ScYxWmhd/za6L0qOdofOxVxziyB1G89IHRY2Syq5
5VSFG0krswflV4WpBZ4xjfABlzIUMXwsVRdq4GL16+ike5+mQquqx9/mDm4gC4TL
rqJpJZdpCaniSndkWYsDXtnPFhjfpBkaMO7jv2WogMUN1Hlp7onkrCxsjcmPme8s
7iWhSuAwcQoaPp6hJcZ9bdGbVlVHcqJog2EZ6hgfNMBAvnWvAbKy6dbahHMBBvI6
7o1YO/EU+lM5a0eeDte5l6ajF9lMWCfrcjo/EkC4bwh3IMHmoWugMQU5WVbrpCvF
KLUSFxL7tISIFVFjDlClkLMH1Ao4lGPHoZ6p7lxDLpImkVLsUvbvu2XgvTKXNsth
yrnW7zrl8QCdQEf1d9AoOI5e7A3WQJR9cKXcAufW+tJd2BJdgDwPqBT4jtFYlEyF
qVEXhrzSXDOGB5HG1ajPoE7BhWxo9V7tAriyZKJaz1K+T81PqIp/R1d8jDZCxpxZ
OuD8Mv9PIeFaPmXfVRUHWv7uolkgVUnbKWwi9h76zttVzudpTpDx9WBwUPJCGyF2
aT8BjCBVSXCnWcsL4NmAhTpkI9Ifktupu1sW/lUp3xFgKYj3fncdVMdgcCsMoKzm
psIdcNGjlGPEQrKPCnJFFcugUwBXqbi6LK3CDJNaXcOhAFykGyMvj24HXpr4oY/j
oaasmj7OdjCHDcnAVD6ymP22rCV5nzjtMxgZ6Wdj3CivmX1rpm1K9j93JVWz+uQv
oWRP3LdghxfemtSDCQyvFmcsW+iQy4SQDmxCSw5ujyWb700stR4X3jbgPNsg1p19
0ipTPCy0kLtfICdrPKV1XqtZ3u/7FlttNawzBoalK9t8+xfmXtiy46foDrlg8F7Q
RgCg6b3nMZmhCJ4PEkJybwW1SpDUfuwu3QrJ3pdO1eFA8kES5L69207wLEKYvKKo
7Vao/X5pID8wBgohBHSGLVm/MOmV79fjNlAxGHNn6mmkAvVIZm6EM+DuNgNiL+Xu
f8j+KRGiCJtsshpGWsvGPS7QraKHei3FfpNpLUtHY6GpzX2MhXkSfKBz2Dy+44zq
hpT8XEdL8h3c5kx28B4llIGFdnlS/uy5GEBGHXzDuIxdWSvLYxHr3qGzu6z7w6Kv
53iiHOsiPWefE23kBCI0mFizM8yJRMrpyFnFDflslA2/qyVdJk7IaJlbby5jN8AZ
5RbFwCHUMdO1xTHVCCrWQ95ykhhBSP5BPWeHc/ZwsoYFtnGHFf+UfQGnZa6hYy8/
xSgryr3MmjLZSSUcuNWyKo586OyyPxK8RObSur9BCFtC597gQEEqZGzSLcUPo5dn
B/OMyB4tn+XgIzndxnwOqj0+Oj3lbjLkUUyScfUm/H/u0b0QIwTHPSj/lt52/bJY
Q2fpMtGd92ACAZ19BaYNPdUXM5jsNMQNMbe0H4D6bgXsi2EYFluaxpJ8jTL+NrIr
RqnfkXPaEjnpYFOCFNbC6k31w+29K3OT5urYpyni89yfr7StycpxKa3J46fOQ8/S
P05IGjqwhg6IqGqNNHKKL2AZPpjGJ/Y7z3eQupHcs8ovf5QNyZpEx2RbNNqhThkl
3sjHaa2NxSZBbQPUjcy/FkI25v7i8PBeQHToA/PYefVi++Sht0Zx29EUfSpalFx6
vCP5t8gb7i8tKQhRbA8+1WvUba6yay4hs3dwXK+85caMoBizMQ1GJwv6sfEvgJ8N
Zx3lg/BRqnN4wnpxge6O+OopwVU94JkT33rWr5wEzIaL0bmYHO5QgAeGUvvYVmDV
/225Zb77kUaLGRqwDk1p1t8VMkOS+sO6wBw0EHJFcOAtiCyWOTJz9Hzht8R1R3pl
ffEscBfTC+HF41LMHI17WjwvhqXXUJXSxKzWFzwtkHQoDhpw/umeToHQAKd4aQ2L
v8NOsuhm7KkAqLRXac4NrRk3Y5zGIehmgjJtFwvFU0VUgO2ItFVdUkpZgXsMxBwP
eNoCJNfWNyfPk9ImNPuPExI4sMXsj5jJbpUe+E19t47FecYXupRNTa/b2jiX2ofM
o9iXZ2IWGHnoKBTEu7RAMWk0mpVlFMm/psO/PNYCUBmwfHElXG1zURxTyEquOqpD
zxzEVLpbaD8u4CE7j0zCgra5spg2o3im5NfHvoqjyCwttnygdbhrGVUwbQYC0drG
4Q7CdQlb0I/SXaUi0UBtnj6wBmxFqv62viZY0JvaiULTlrJ910O/pZ2ibPM7v0qE
JJiypw9kZdnlgdQLrcC+e97uH4bXY7NeKNCbLbY6rafk2PhQwQYT/Ku3WQM6XMHy
g3kJL9vZDdqKhXe8BDgy/xlYH31+gDTa94PQuTg/nFNrulpNjxfOheUEsUxvpWxz
Nkol9oV9B5aqGOzcNHhkmaDrDOy/4Q0oYVWonz0VphrU3hjZ7IwxvFKdC8/cZBgo
Q/IEvUrvETgS9YNBTvl1A11oBq+qyU3Wm7WT4nWMrKKWemBllLFJ3wiEf9ieNfNx
CTZVUkoMF5vN9eUDDhuW1qqeKUQBfqKBXXZAn058/EhWF9WuZ5B3CdiZH9M7WKi5
beHBzQIzD1ti9KUDH4i91vEWBU1i0bDriD/ypxyN4agT6Z3isQ6S+LDVb2AMyjBP
B23wxAZmsM3XcnDHNTIWqe3alroJ+O26DKii1PQ1Ta+9dRQ8Ru8cVatGAZqljYpN
b64jxNRPK4wL2GADmbC6YarpDDo6DhDa5XQZFYif+pn43GVWAz9jT9RXfcqMYpd7
ynIS9N5/6Km6K+QvuUrDBZgThFFHCwF03QjnP0aM9l/Pex3f5uldimhhAbpZb05P
Cjr7ZCD7qjzcvUWOeBpclicGAPliL3R4tXJ3ZM/KFmuIOMa+7NOk1habW0Fv2Ie/
v569I67GWTbl9p7BSdMLeRRusduPCIo3oQUdV2DpaKZhSYt3lfa9S3PaeszRpSpr
LVxwb5BOVwea10PvSAm8G5/Bf6U1DcqzeEayQ/OHMPyDWRtH9vfeeCe2jYBHUwUH
dm3NlhcrnxlrHEFYpwZ9McKVdXkhvP/kE6t2wNxyGzEufMBgd374CoWbkGekdT4/
ZlaucPciswD+uZdfkrxaIpQdvzBIXtf9DHQEfTIL/yqO66jL6xGbL4j9CDVfoBZ6
h81M9WpciOG/b9dpMYhGtZf0S6OZTxdjqsekrSA9yQS24h7K7VChnNyeJm3zDqln
Cmjxnofrurwm+AgAWTJgnr1S7ynQto45ykmks5go986AkssVw4e+C0jEZSDEjIRJ
CPshzH+yCQKaDB5r96gJdLr3S8rla4wN+b9GrrT9acno++DeQ1l+7eLrcJN2JDZe
F1L8DYFhH6MiC2olwAA1nGq6dJx37RuKo7iiYL/q16SPyeK8oWVx/+o7tZS5cUUe
rXs/NUuFKkuzwpKdjCYqSGaURVqCW8NRjDKYmCq6+JuX53kLwcvexDTNDTkuNFuA
elXD4yIGz+OSKaxLOU6cZKsfwxkCjPKGvdge4WviG3Cde3k4n9/aJyXCM9EeZ+3z
WOq7pJMtoa+3+tSKGr6xyJoW4mHb89T0FYX6JgeOmSyjMAHc8CCqLoiIGACIMpqh
xCfKM7/9R6MqcCCJtXLlQb/wpdlSijnyvtQvtZNxvPx1iEYQnkZNWaW6Bt8NnoCB
N0WuXAVNJSqhIzJhQFrON9de62Piam0fTI4uK1zcycZueIXasZPuLzZWSgERBNOV
55ew2Pce3S5MVakaEoc/AxYmeONvYKGInS0YuT3C2Vh0VQmHWztfiomnMwdQaLmh
GRfX4TJcwddsL2piVVI8944k5rvW+vpreZp4bArKj5vxeP7nsb6qyXecmZ4I7Aoo
YqHjiRr2WM7+E9fLJhy0HIT7FBcD8haTgsGlP9iE5Tr++8Q/UmcnDFEAyVWgn28d
2UHJjt+wh+SwdBxdZoz6LH/orsrOSu5ARUbc9CdXQJ0Y0WIKegOkTyNpeN8OY8gy
8SUIwPc19cpja1NJkA//b2X1YWRdxdjptUDFUq4pi0oHcJ4qNM+abY+x5YoLe190
nLy8VMUCgSeKO+E7uNMfCLxyFPHztSnN0bXinO/hnx90SmTOC+tH0GUFrE0nOsqG
1nnJt91lrV2FedN8aYi87LOE3ud+t9OB8BDDq32hPixOKsF+phtIRi1gQKPplxR6
pAHHXXz6pvJ8SMG5Vdi1viXVM13pdgMB3nXqSNokuIxZwSlBqs/Pwqp8VqdLxagB
PHkL9pESh5os+G3gTyk+7QN1Kdrj/8eGoVzo6iHq4VfMv16EKqBE+Q6puwde5H3O
WVsrqbVwbxpkgIVhJT7BPLWjN8kf+GrHJFPXXyANc3EcaLT46kSSglFc4tl2E6Bc
p3bwarVc/12cq8fbZpr+bWducEKHueH8twbsFBA1lkQ001ajxHKRvsooIivkziNu
mslt3a0u/s9WZYi5BnJ8BSCa7AWBu87eSxsfQBSAXivDCE6uVcEaLuABReDTNilT
+8w2lLSE6L0mpxdf/c2+x1GRiJGfPbkqbDucKasrC3Y4cByn+yFj8/D9pUEC6fNC
340zJeY3eYyDXSy6Ngfsc8F0X/qbf9bRR8EA3Jg2AelDAOUwjLgiLm3F2aKxG5Vy
JbM8futNGl/yOkQqbrqYHxydvKw40DWgwWRc6seMRml4FkNpzlwaH7A3u1wGPl9j
zB8k7/h8t+dqFzrEET1HHZqcAj773r73Zys4VhpDAaBuSvEJuQ3O2nZNpJMRKLJA
hz24/JWa+WWgDpdRksupLpaISx2oRBnEYHes/I0BIHaMAwSoWR9LreeL2t9OmzKo
40e5rmxaiH1fiD+0KjuXiAhv87uZJm+FgM7xNkbSPncSKLPNNPxKG+GqSdnYLVhm
6m10ndJHLm9HQdKn9xAB3We0OZboDsoG6Ql8jYReLLKRqmkIeH+xrnVjC9ieaQ8L
PBEZtnkG3JfQMbNsv1osVbs/aN9Sof59L5dHjBkSF/5vsEQcfPo6I3LSC12WEugZ
FYHbQypH/qel2RTMiO8puBRlN+fu4qdTldypeo3TJ3CMAdXd1cz8iqcrf2wBkLbK
qRxetxDNjnLZ8WOR9dqCtqtah9UZQfKo36SwMU31bBNzDQg6gD5Imjnaie/xOg50
36HhyCTtXWIzttnlLYICGJNZq2S7RiPhlGi5josfE3EEWDgEB4qYtP4/Sm8oA+U+
po04jj+yKzwVdavuj/puF4Y94xNmo5iHYICSRFf9yE6y+w9sLvu7SMtmx9CBQIJT
gR+X+um8xJ1JTUk2hX7c6goPypcb5Dg6TXAGgZEd2k2IGZtn/74qqw1m8xXRpsm8
dMGXk19qXldXMWyBY+mNMNv/Gq7rB8MfMMR+QAj9Z8kM2+1VJLPlbcs1+C85g/xc
boExRij0hmXmhmnuSI90eo5fLW7YMQCm16kQPQ9in1JzTOaED+tKURnnmKtJ4xhc
8K3739ybMx+wasy3+I9/2L+AvaE3s4JRUEpsPQznpht8+JP9e4zAHYozDroxsOjg
CfjAPDBFApXOk68AhAuP989OJUH/cC7BISCos+OTmqTsP69r1HLAgL+mAK0XcXCJ
9EJYyqhbuTaxILYA5L0qjSnJZ6ihgleOugpSvFXE3sKfM8k9jeJa2ec3xZ8FA0ON
VaBI7KERAZqfBzYnnBcChgD/CXKEyvexLbWMzWJeITZqoDasvOkCZakLuvR0XLjs
ozso0SHF+LQUSuShlmjnmQM7dWNFK38FGpUdHyVX5Zxe74jHQBd1JrgsAKfK0l0A
LeED2kuzH7hrfeJoqDc/UbrB/C20iRP7q/LddYcIRfB+0vZXknlF33FSfa8h6t7z
eMMt/8oEiJt4PMutg1kKyU2cb0S9PwEBpp5+D8BLnNnZbp7D4i4Ico7qP6eYGbjn
L4SbOCmVUFj8h06xM4UV4LZ/PCkXZ5i+JxUB2w9zhunPXJ1J8Ff/Vl1wAEATrxe7
UrSkJC1EgZMNUAVgTmzMh/bltRkI+INBzaVrttcQJgeiM6IpUOOXOzdNpeiez9yl
3hD1D88EKWIlap3gArixA6y/kdAuwc/tdd25NkR3k0tvPx42IjlmqdDtnAXVPada
GUUdS2rW/BxGYh1Vx0YQaQoGpbUuRH1Oyg5MG6Yqhsgof9W6I9QBDnVbzE6UKg1B
CpBLCJEClVWx085gYGsq/amx8BLWtmw+Olalkf2xtN2KVhGs4uOmZ/DLbuigp9J5
z5U8GpFodsIu1lbdiicRNCGsibryBjAUqdB1XZGTpQbDHQ3wrp4TOprEEADGr5Hj
stcyvjw0EMunV/TTFpxjaZbYxmBjkaxEY6zE0Rw4/+cAZ23zXDnJ7aaqpTaey0xd
4r2XDDRPnxJ8J4ITPxUj3y0OrBgWkHEIdcq68YVHqFZAQ4vKs1qxPeJPdfrjff6n
ykPQ+o43jZ6jMvXoWvU/1OAedFARcBMXo99Kv09NLDr3AQ03zaw3SJT2nlhZTf7a
n9fi4MNTMaeRKXE/92h1xRnTDv2QxQ4mCnDeyfQhKXUnU5bFSk2JI3SX3ud9wf0l
7aXENVXVY+N0zijE0YfYIaqEy78zD7uTYFQmVcR6K+rzV4P4pJK0WTCd9FPNzAfV
vtalKDrPNq5xJZlgFfl+xn8WSeE6zE+HbsHA+VnTM/fSzn7KbrDiAdJDiroqN+o+
JgB2oO/isdUACLqshoMF13zC6tPRbyfx4W+5XJgt+abkPPGaQ+KWb54Tjbz+LQSK
B3Kc6Cg7EjY73NQqzsuWxU/HhWiF3buHj9RsjtFivrQWijoN8CVdwIxNma8D80lc
m5MxbPjFmSxxEmGUFNu+l9uxt8AfC8C/4u0dCh9Dz8HuV8ICSaYQ97GSPiI1jLyR
/6jO6lW0S/yWyyXA6epguWk5XGUxoUrTjpqIGj4K6l5kPcxTbuE0MHDCK5jHkgw7
5Vb3lRFHpGWrlC+nCqhuWTH97l3AcwjJd3gtf7r/b6xS5Mt6DATK+aXLSi4g0BD9
uwmEcXwnaTXHU6jfW1vKLVeccmMBu46b1+fLW9XZaLlHJNvhThGEBdrVoGhapfCj
paOXa9K6OUVgFo9ULVqLv9yZVnFSWWmul4112s2a+as3klSv7jknSPOnbIrii19O
yJt+07HOfkCI0bxxB3odXd+1QLxTU+FvQoNXg6hM5UC0MA9vrcZPeny1TQrapTwQ
RpyDmnKmxhQuE6MxBZiUphK/WLm0NoFrPza7PuS/ozbT1n1BRlysbJ1RFFrRTX1g
OW/aaAwa+YtjLsyt+/LKq1R97AAmvRZLfd+lWcXEbfJMPawqILdnZHBRH2vm+u91
S+5mhurMUxgS5JlSjGteNKFMmmm8etXBIhTrGF+F3GsMcxwIKUOpJHxy85hde2CZ
YKpYNTBpO5KGRn0Fwmj5F8huer7AGHrboG7y7L3S9VgVv6lSu+yAUg69gcXRRxQz
pmjGryTqud9PEE4ACRS0nLrDrz9nI3b18rPJhlN5jboklOA0kZdiSWUZHxIg11nt
bw8wgl6XZa9UDBHGtj4/jp4Gl7xjP3HT66kB1jx/d2xwTnc2QK9i7dNfQHZDjjop
xQ078mdPZ7BlTBozAfvgAQr9OgMiJ9zXTLtKoqfeO2BP6/fypUBBsvETFLp10nt3
K8Jmru+sRURodEkSIe5VYinZRF0gJBPc0772hH1xHcfsohdSGSm0u8OatIgi3r4m
MJO8wSfERX0nya26IIOjE2yyAwoci/yPm3AfjMgtFP9OJBKpCW7meOUaEmFAWq/y
lmRkzaXsByHBIrSOzKcRLLN4h/j8Qx48Y5KHDFhoiu80LJBohaopXuHFNyxlFEyy
uIsvdwzH6bwP0/tAwCMFg3fL2OYzbhx3ZrN+v7yF83UxZVm8yn0Fk5DDfPvGL6ky
RzCPjqoZX37cON7PYI0fdf1BREwINZZ9P8vdPqVCJmTiCrdyQqNmaytqYB87VtXp
dAwTwCdT+funs4K+jj7Fy4W6kFUNZpm00slfdQ862SfUD9G6WvqGOshp50Wm92KA
tmL4cezNG/ptEByPN3kc4UarR36PgwOG8HUkTWtFfOTBCXJO/zlNZIOZdmpR5MGF
xfFdtDGYRBaLYSSjz5sP4AWKVFvmkWDjkNzjHdUSKcKtZX7gp8yqiA8ijF2TtnWV
n2ITzUk1sHZuGVd8eLHODb7vNqTpTNKue8GTeXAbACZuK7f2LiNt/OJPnFB5Pwkn
QYNJor3DMBsABvqZkKvyYM6no5rYCHNyNxXbFoCztDI8uyiXvPLH1cZ47adgN8BU
tw4HJG9QMxkHtC1aVZyBPyn3WXxP0F3WLM079N+Xc0vGRnma2v6daGWonjRjlM3v
Bz5Z+EJxUfIaKa5LZ8yFXgYjDOmQNADprChhykZ2U3HAvjYYRThvU9xCYpdP9akF
kTHDUsEcTu5J2JRnYvqKVtglZlsH4tzoTgQBVdRvSzrbtkLHwC9M0OP4T8MUeYrT
u9qgYRSoKx5CIbpdSPk52k7W/Y+ZOVSkOOkRr/b1jho5vE3TbdwGHovsY3BWSW0y
nmIHR7tpFOIcnsYLRF0amu8CB1Wz7jw4212JNMekF2egLrD0OY0tDtkpAKkl05Zo
hFMdDf2bDbZQ7UCGA3MV5K/dqYPoyGZ+4UMa1bqzhJxPE6XVYxgshu0vnUTKft6G
daOs+b23uIk+glo5Ast7flyo9rdh7AuRIwiOAqafdfdOOoahxIlue5P0RC0zkipo
0LiBIIpSvMexIBX8xC896kfEk9+3/oA3GgSJIx+ZVxs/HqgS4Iz0IRoNtnPePfY3
ICrAs/fJJIIckPRo1wFf1k16A9gO8U5bUo1iN30gfdOxydc+lraHLJksH2dFQ2Sp
8qM9CuRTg5PDBbayQtz0tq4besiSFnUYOBPECUkfI+l2A/1zv9iIvbJdZUml8PZR
MdpFOwGX85W58jJPVO2dlrqI0ufJMEPbuZ/WW/3wyKybhSLOxHMP9cNU8spqLZTG
acOnZOPCTYL94uDsEXPUKB4i10YjQ2oEpsfZ86rLHlc7upkZVuZT33X8Vtgdcz4L
S663kcsrBw6TimwZO9RW9NI7WYx+kvbN8UYrUvqsClqVQ1au1gcZDi1MjqeWLa+P
5we2Zs80NtrOlGWWkMv7KcBgSbSocMZkQgNp7ScCnzgPEfjlNUCvQiP+9rHFcc2h
aWy8UXl/3WMYLvM+igcYMKNzLGxfS6BeSfLi1rDdzqI9hwq+40c3/6hosuatoD/T
Sdm9z2Ppgw6rJYItUElFJtQ2t+lHdC1cCnptQLraqSfVcLcOVarBSobgx7qLJQd/
EoLZbkEFd34/xFbnp3P22lRdUwjPnhofFv5nS1rG7HxBlJE32nqkeXTcNdBe8Fp9
XAs/jJ6he8r7d48afxdUCthGNMYYlZ9385TGB2pOn2seWcTaj4cUjkVlN54HiirE
J9Gna29k12T8rnygxR7zZvq6CwlyNUFFXtsGiRF9k9MbVAZ34miO9a0kwqkVFZ78
PESZdtRAdbhANpMiBU+9/mc2wsZryBSyJMNMmGAodRrZL4UhpD64RDheJtTcCO0Y
8KFkRRDSBfemLQB2/Qps2LPXr4RbRYA/xw5RKrgN1Aach17TLON8iGQXJS1B0Jet
5RoxAwHfmtkkGWz2/artBWhUipOlo7AZwv9oExghJxUcwaO6giIXEBq6ml/U0C1h
FU4CGtOFFis75BYEA6mSz9wCxmiKK0Z8fY97T6NfY6ua1WAlcp+tzTZFtyALKtEC
VOB7phPdGrY75dxUtYo287htvWlov3u6DT0416ps50fwj9TXwQ4HO0lQp21iPR6s
760/JXNW/VcDFU2s4bq09hWfTG3IJx0G1uzkVB+tLKG99+WCmseqKlH/+mNTbW69
3NrLuFbsQD8xaZVnjTn6O8NXUJ1UwQtGzz/rZ43AP6MncXavr0DiGILvyzB01xBo
hHDiP70PEDs94bCgrx62tnzYcBgO6JRWEb1KcG9OhP3clMtS3/Mz++uy9vwnlEmL
rLz1dZ2JBSdJ9X1ZcyNzRrbYOQEeZy8ZWT3ijf80MD016Zms2CyKf+rtsgynt9Hf
xn3ePJXmzbGgAz94YPzpqEUr88hl/NPbGHaKp6+gQlBpjtkmyJyavtsitdbPWSBy
D++Mt3SKyWmkxu/FhK2AoFnjVumCqK9p+WdpxA9YyPkzHorD1jmv7VeLEtgGJvQz
t7X3XCLC3BevCCjIEMOMOvsjg4LPWDSntcb1FrR3USNHgfUFK9EVAMRkDzFU4TZo
0qsvztcQb7kKmAC264sUODbvU7/AId2oU+QF5nW7z1y5geNkUKOX50purCT0IUCm
Oft0FleSYl3o66gci7gssWVQV0sSExDSzd53ilEIrD1B7tVs21WCD76sgtCif6fB
x18gKd0HeGqg7YNWxG5VmlxN+2MJr5t7GjkoB8kjPEf7lYU/VB814s62kfYDhKwQ
+QJ583+Evd0qq9WeEfVDuvw+8so3ijpSNcUuvxIyD1x1x1ueAs99CDmrlomgClV3
QZ0IW1tNOHMY00erromsUVDIKDNAXJW8x7pVE4wUfcAlVxO9R4JyaCB/uKh7pmIx
/n4jZaY0wPZlskq9G1Z5VMD5YcaEBYyotTV7QsVRkrkRWBlspm214JEgRVZBjJJh
SgypSmOk+5jcRvN0YPW2GytWXmw981J3zc3zE3PB6Cyr/oLYoFuwG/I+Ke0pysTJ
4lDH7WYq15M6QgnKeLtRpp8zf9lXbP5+z3oqfkRo77M9r5Nq6mdLiLYFNZONek7v
mCwNXQY+0mCppRQcXBIlCCuXFLQKkZAxOay1yauaC/c1g8YgHa2O4recA3m97GKJ
+NP1wuBcNOFhF2gkLx+HZ1Mi6KVC5YOOyvVrm4+zuPo4AgVzoN79cjnHGcP8HfNc
9XkmqLb2iIpAMUVtCEQX89wT8EFuJZWrApLlDUPXVc4JSqOGUTeIcjLqywCFS3l3
ueDvmIlFSLkAdGZuaU+s9VjvKiQVsF8hAYLv9AFqg37fidZJLY0C3ku4djP5yJEc
5UvstcxUV2STTIpvqjSqgLEnBM7/yyhrsETqnBA6Sb5cXMmHRsWo/E7xIn+gGWQn
OCSNPu/O64k8rLj3xCZX1wEU2mio1UW157GKvi21BIbIr60J9xB213B/im2bAqHL
eh51wuqQbjz4s3UrUigVViXDTk+t9DHIvfopfpOyXQy347JzTo6CTYR8bU7pufCd
T8/qysp3A9ERbYeFf4TwNO3qmTBVVjI6poJU+AJsJ6lviCu9EO+K6mujMDBZHvQp
KYdAjE05+FV3k+lPa89ljqUKn16aaM0KkidvDZO2ZZ1otoM/B5K2QtMmzTxHkCgj
DyJ3gL8baTnqvSyj/iFB4BRwOVQiwhwu0CqkYcja9nDe4i49m8goq8pS/1DWvK4E
wxRIxI5ucaEOZY/n6R1MaSVGKEfLlEIlXZibgJCyX/7SVBtnrI+tMczuNTRZ2RXE
L6R4uZ3mJCaIbXnbHr8wyplWs9NbeFpAFEFjmdVT5WcGg2SYgtPM0/JNavhVQQJb
h49YS9vTGfpDstv6bxS85os1McQfQy3Wy28Adzu1daT8Bmmdo3EuFR8msm2ceWtZ
WNgy7b6TNZUCfvUF35c+dgjR/sn1bEqb0wCTsi1baWsSiTFRe/kdzF5Iuk025dKP
V0OrTeX0jaY2ECV9CUT4RrlGnMzyeYaaxT3A1EfKSgCkWgmiyuinHI3QJBMhnohJ
X43qgEeUmQlMVPwCqvFlaaHLW8yWLB44L28+uiTSMDkaUCsv8WHZYQf+XcozLyTa
3OFWHqpLZtwn0H5JY7JDTs2mJY7GDy4wlDvAc8RXgffpbR/KzIjSJMsObfJ81Nb1
5TV7zcP0zoV3oA4Qkwm7irfyVFo5fasofJRiyDa6PW/fKzv7yy3B+a+ms+coH4EP
FQMB3EjlgFRJDabMg3yMqb9XJ8JwuQhkBO3AYzU9w1vKgXEKo6CJa40G+wwqOpMV
QzG2nggt+BdWTE7cBXKgjO6varDOpkQFxXJpYZYTz7UaTAgbPfxXZEhN3G4GIBwQ
J/yr7fV8tRYHpXYzsRaEaynsnVwgnAdRIZK9lfuK/d/Dpz3vuVn2EPaoW45Wztb+
exzH1t+545pzIVLTU7lXae6Ki/Z8I5wwPTUyXdmP1MI3sJoKINAHUTtViRAOO+eF
VJAxlbCh1FYnTi5BaONzkyFrK001/BSF6a6+WGAWZ+IvvVbe117gSG6YuTJJ/96L
zd36rlmAH4cIZ7v0lTCFmd4tf4hpcNV3kfnQb4XmQc4N61YAmX6hK8DkmIYfW689
K9Zq2OcyVXXMDFnRp+dxROwhuQzcGROBuSCMm0pbZqZulgK2Q/dQdXe4WXGSOMIG
ZSFlluQh66fZ+XYR6dxp5ByTpjlh4tHbaZiaSUpdQtEoyF5nBiwPrm6mRUnulHv2
Iq+9DQkaUdCyUh2ih6tHRWCp/gcGyTusOWrWdvCexwr5CxP4MWeCwqudAt2xF4om
vx/vY9dNwiYHafZ5pCR+6R3ari+GrVECwz4srUEqFKEk7EyBLg6LRbWWe/N2sqCp
rRnAxEEiPkNzwY/dbPR2b6PICCOizZQOB92ms2e8FL6jWhPlCXbaLDvaxLz4lN2a
ks0l/iKu9XIM/3jcFoniAVw6Hznkek6T32FMWBQZkeTXEONcxGh9wAF7pO+nVRXq
wNtajSKuDQ+4X8KAgEB2kceYaltsXhvk23k/2AsToIKeqOXAr5M8PXTilvYRSOMo
ILz7KHWhQuf3LcbXYT13LTiwFmzjJJ0v1kJlmOXKH8FG1ePxnzNpbFxwCgh4lUqP
SZhMPY0NRqKhwT3DvAH+SjE/gd+cEFFmlRBWBaQk92Kzw2cmVz3x78fmlTN/c3rS
O4U8lcCL2ViTbwJzE2Dk7rz0jR9IDrsBCR8fphyzXw0rGW4aSo5UzNSCFclntivq
LUkYfa7tj+FZ52BDqIQK2uDrVMsKhgZcM8xsvkj2Rwf3SSwbVoXF0w/1TXeSKtUh
W/u/vH3RH6rb+1Z/6ZYjM+Gj5SUJ5g+LtC5ndW9Gn8z0yoL+O6BlzTefHSBxMIuw
B0BrYvT+lVOEG1PQwCzzB5Sqt5HVZnAedcNVhhkjfh4EcTaKZZkLwcad4tcXStJ6
jdCxIigO+5J57+PZoVockUMfK7vPpNaH+qeS7ij1+MUt5CVSXzNyktJM7iCnpYDX
ggaK8Q7Ii67wfE6n+imxUC4lrtfvn3Qw8/QtR7VGsCcBZLkehOjBg/V0HlcbzXEC
hIhpo7uURNIeatHHec6Zkv2Q/otA92qGiwG8b2PIYrpyJBFuXg+vM8VltiKuvvHV
zEoO+quYbnHTLocyI0pZc1yl8WQZvCke89J9shJK8CQu8cSpJe4qiuuxP6MJ0bMC
D4GcJuqQgO5ioJx7rC9jsRnKLsCmchib/2OB2iTwAyzdEgm7SrrL+KfEvBNp3Z+1
N5PTdqrY/3AnE7ZKWvOPGcYv7A+yz2jXM/lu4i6z/fMGyMkW0nNZGdWUWAPdz9YO
BsX4TZpEgVmO4fstoYlZvj3D7EYnFba77X3Oa8uy7Dpaei1FoW4NRAtxCTPgrge1
CI9V4Ixc0AiIskrBWBjNXE8KoZ5QO2c/wZA6AWsJsmjZnXqZo7eWXyANicIVGsmB
InrZ0NG5LBq8yRFIoDDEGzramBuUSHP7qGR0ZAYCUg5AnhqEVfhZCJNTmNB72Rzd
BpI7HkoKeS+XENhtpaa66iOno2ue8sOU2GciPGxjotSdmKqGJUHzYmdvFIlYcoCI
ig+7BDqL/8w7h6jb6hWhYCXGEbc0eWAVGZZJsb7KB6i1tjT4jZX4SF9cxxdGvklG
XWFEwGh6hmWUbjhuouXALZcHgZ8dMBezmje15EksXPc/ShgLV5Aq8Ixl5JjaK6y8
pJWXrR1BlkH8LICdp+WTwkQzrTjJsdp/cIgEBd/qyLrs8bpROFWnbCAZduTzKWaQ
NhmeeoPKOBP1XDLQYnl2zL5a/eXxbg87vjmUjRxikeW98ONB2BOalIPQ1LRweSBV
bWP6JAUU9t4rxbTt5vRgo+9Aru/GCrHujvTJACxbAl/BwRZJPZ6p5bB9O1MbFzGz
RoPYDx3liTdE+wP1PTAsH0MjWOwmu5Xns9LJJ0UAnvS8c5EUSJkf4lcDasmKkPTS
11NlCPAGFn7sXqK/MpsZ0uqAQKybXCCE8MKsVeax6vMkOOeWtEKBL7Pe/ptLCDGr
KwoyTWlPGXerKAr5vhfvHKFQDxp9s+SG05bsuawjdHxs4AZWwaa3iVEkNho+yyYp
Z6hK+1eNmqjpXEu2L2MdePPriyDMDDogrXWNkX1zf/evnwhrV5ipCvI5XQ57qC3i
0AG0ONg3VxOquiAR02GSrMXDj4TVOuTYyfVQEvsRJjOM1/Mr++V6Cz5iUrczeBj9
hPrGoCCcLR7oMixO0bk+4SELlhP85bke1fdOYtSAd636+zCAHprIjWepGE9NxkFx
qtf3db4paRn5giqQxnGEEeH1aYoEuD5S8GZzuaNfp+p0OGN9OgjhcQWnl39UYGaQ
QbM/Cytlgyc2BFvTwdGkPtY3w1FTQSNTNMaG7mefjzemKPokrkE6QFSWz8Vu78Kt
Cl3Svg7YIAhZiUA2TcEVifTn8lyRJYhGlzfIqZt/4L2qCvTwxgrnNma8zLR2YPpC
zSAwqJkAl+liCdv9drx80yvc6SDRxsMVF83qgoKdv18tHPbIQDf2GJoMflVGqgyy
pu93ds0ahG45QL61agk6QdHWih8EyE1SGM3VaKc62EKWu9E674tCtJCiVAgjl1Zp
KQsbi0xEnfY+ADj8OJuvZFSV3tSOzjQvgaQ0DliX/ZVoYe/H0kXK3qQT5MsWPQh2
t+Y0PZ7N4GDeRwUME0qXlJjjtZ1Ab/YgGsibNcbgX+FhwRlqVZE9cLxwP2+fttd/
VGxfHS4XDIGsY/TcezH/Q3NtXu/QvTO/z50I15qLbydEJjqijMQv5fU0/kLMmYdw
oI4OWm3z98dijNm1gkEF5+6Ae12AnFPuBTA6mNldYcdbNy2CvTUK64gmd+0waxp2
6vehNAdHi90eshDwvTZ8lO74asI16tzUCrT7XY213YSGDQZgpEarcyZCwkD33ivO
ufYgzkskuvPSMYD2yKJe89ehiCRg59hLM8SeVJeowHwhrG+wpu4unQp9PqqSY7O6
LWSFeJ/rqB64GXZqWSCQZ9k6eSes46zN/Eidl7T3Ju1lSR/JJwOCXdWG7L1XOyCa
FkWwMt6MTXEROsr2Wl/sclXRiObDkbaa3FU8rDjnwWBYDAu+prtvQDauU/P/KvPY
EIPNijxboQoFvyG5KTeRvwQRKdY5j/lMVAsuHyJeAPVrxdmbl8o4eNcK4JsHbRnV
nlShTdIq+fOaIN4v89sgsmqLcFgL9+whLiYw5H8sJazVcB+tAe/WDO5KcIg81Ydf
jDw9XGK20yCKtDfH8q6cmIZSmp5zq2b3yv8W/wjyjEQ3yVcyP6BU/XYH3aSUr+Oe
ZVYu1F9jxoVOBPLilcUwtMjo5kwLl9aJtAk7H9IViw7TiS/u3TsHM2Vmu4CDxaXE
icHzjgJEVFKm2ladIZHAq1cB+GEMgyYJBihvjwjqA2s8lVWoPovXHMRGhg8c4ClT
zjXQZixuTpyoJSKDoY+3EOwZ1Ya+3XG8onM04IM73+F0AKhn4SBucQo70P5FmbwR
BEq7m+dmH5cMcFirgxFywQ5+RE4UCRlTyooFGP23kCiFFA4Bnr9OSsDJpUG0evRI
hp7PPMml8H/t6SVw+vaMG6mDuj/HORwVhRs5z0LXJctRZU6FXu9uEOHNEsauhML5
c5zYIhae/eNwrrziZWfmNr0p+OLDPi0VZvilfS249bKvZxXjgvzEaYRlkuk7Ss0X
Cvmi+tJUmu/qXjJkY/zFNQdnFZp8xqBL8rMTpiBEAWoDzfHG6SNWP/Cqsu4uEeKt
/EjXsbDw40KKqJ6C7c9akw+DWVxovQZSHMaju/MoV4GoHl+S1axQJRrbU7y/wEtn
LRqeciCgr2NzZ9pM4MMD+1hiqQQyRsgQ/3QmejSXXTbiwHQI4IstiuuIwU8xkXKz
v3MCyO3qJj/np+/IoXIeU/aRfeIqvCTeR++9Q5J/MTn/iZ1wJCTq0P/thOWwH65s
iHzr7VVsA96Z9pCmoId7j91NjRA8p4KLlrALEuMkkHl6OkOozEmgg/vI/a2r995u
n9KLHN/iCjYBDz5kvYscYio9OUokMRIRNMImgECm/HXbMF3+29+rkcP2/TH4L1LB
O1VyhgHf9gDh7WMNVZVQD/0T0Q2GiCN+bvWuAfRnY4iEPWmQR9Z3oS5dQrTJ4GXN
YmnQKFU350Zn76FEZWT4GIuFCCGIQ+pt1ndpG7fm4wDv6y7B+3Ncz3/dS4+8mP2d
MGtcqoZ4Q4dIbSfyZtDENkMCs9RoVdw7IRq6O9a1pl08sg5y7xcyc+33Dw6YGEwb
m0OyFf8l4y2Bz+Eht4+P/l0IdFBiGgSCVJP/DCqVVV9TYldvYJczJ+sE4Cc0OpOn
wqCS9C9umDD1zqkQ1/bK/RLHH5K501cyAG9L41ViwQ19KV+sVvPEBuEPI+7oyHDG
06v752oNVNZm1ID2ym5+5D2gW9XFffZ08hs5MPXHhd260d2tt3zpWKWg9V7+Mb6J
ozHyeSa2MOcS4BH+PvKDGL9l86kj9cs8divfSWE67P7Gsfk1MqrrTo0ACQ5JSnNZ
cxWtZSD6RqIpTQ0u3xr/hMuxB5b1eLkYvACFnVbTCxwfOG1Db+BICr8sRLv1Wcof
hHu66LuHuRecFrZtaEbU3XNjdP1/DGi218o5twDyUugl/K7aTyi3LyoQFuhAV6BQ
M2mThV8/XjTUJPZsHcSXK+9ZOz+hXsLGEblnosemXWjdMwZ6u/CQF5sNYlPNS0TZ
AQcl8KhD5azLPcGcvH5Os7GWEp22w1kpofDkh0lxhBN5UDa1wTiCmV7uQ22Gp1K+
xqGjNwXNNQF+Xqgi0xbtOHEjyHMsQ20S8eu/5gE9mIEgcvskSNW+uFWWI3wmVOSr
ssTcODDWhftihPX72glVc57Kt361s9Oin/T+/0u6wQrOmuykG9jsTcL5Usi2ea8S
Sosro0JlSnXnu2Xdo9PgDSKcR+oVNWfG0qKrklHxxngtt6R1M+Fx++Kb51TFrHyx
c6X4d+G/+6244Uag1K3dDCCtJd1m+dxNX8bxJk6X+ql7HvDMj68tBzRGWkLtPzJR
M2bojqlZE7Os6mPvFhoYeI7cd4B1UFzx0qdsdL6ng0ZedJFKEhVC/e9Wgit3iZI8
DESYAhQuonVMB8LLPNJ4Sh7QBaqMmLf1k1HyBr6zKoyPBi+v7QHLeW4P7P8AljMa
eSlWooRYoHEVApqCg2JSVipz+n7MS/3CFMU08EB5/TJZ+LwmfbwkKPfkjvltAKY2
xWsmadYfIgLXKu9yBBiSiW43kgYinF8XGLQ8qgYcgshMveCJGNxUgSffjbAChHRu
zoOVqaLz7rEeh8o0/Ea4yo8aPirg3xKsd0PpXwxmLPCnPPDBGrXxaa0+5rD/6yRM
5pneIkSi5VxgKUVflWOQjDL58H5Wx0G5LXgyzxI0CuT1XGxJuRcFf2xWtoOnvWEI
UFOqGMy332sgKjsPXuk+mC6JUL+Dbfwv/oHt2We8IsFltmzGv+VMM3v1JqfTMO+h
/8K6j/4+nDS7RzMuld9TQtaAFQ+JH108cbeQU7uoTajYbPLf4+SSvI8irTlZIx/D
mlj7vZvByayP0Ht+E8fC/IC04ch5acBv+EwNUx2FjyZcQI7yOWyLkuz0j0nyecPI
vuKz/IESqLF8aAUWSVB2nzpNG19HPGh2lUckjJM0H3iC5rjMKwDpmCElQjRIc0KQ
3rgmIzAiz0JfHadrKISjZepZgZgU9IJyDq/Eqlk4Zr3gfhLgnCnXfYkbvFYYuCva
Wyf3EvQj77PoY+ETxS2YS08t4LRoQF5QAUYWu/DQHQzjs2lQ1WqV770ZL/S2MLPF
iUyTxB4j693My+mcdogXJ9INReGgPzqREU07bm6Z39WO7da8FrmYuliUMAof8XcP
iGB/Jr9o7yukX9kyEyZvKpj77IE7xgjpg+T49LX5jXwHcx7IawwYECVS6Ck1IeZX
mEddlW98+cgikqOGY0aoFrjsfkdn3gtMDjAz1gyGj3N+KfEdKd2cTeH2T773ETfb
gCRP4INAOc6sbr3udpUPtzRkrPiMjHD+agk72yETpDWtcGE59MHZJzsRv8tCfihy
V5i+09NbS4/YlbmLS07EnYGox/vefTQcImKu/T1DVp665cF1SGe6YfhWrtY+r4QP
R5BAehN4d/Uo2EtkhVCqtzuZFBWeFTelSyGQIBbFChLQJfJnz2MqIiH3KGzrPeQt
qnNPgs1257j6z7Qsgi936nYoL8BTjDOlKwibpWzyeRDCkmGwWqC0suFHJI/sBegZ
W80U3hIP5i5dVbaiZsiUYC37tIB/TuMXZMi597AUM518EOpoewKp0LW3LuzodbnO
h8VUGYyVtFG2INV6qS1jK5VMWklkleXse+NQKIERdWtD46r0WoPQrEJB8JWAwwg7
ibTJIVxq2hJGtDUAy1UxZQZIjnQEv0FsJ3vWonmRvEkytPM90X2AVcOCjtw0qyFH
uy5WFMneLiJh2LqaISHgNdp8LFulzar/xtM4R9bMXS7tcIHO9Ea0VFumFTXTenCN
QZbYw1KK4iA1Nz9N9dXgv8jaOlpLFgOhyZxKlW5SygsK4BdlLE6fBjY1qdaCMlmI
Pp1ZpkBb7wsWdKxcTTKBMp/MaZo4d9FPFfLfMLbcucqlwC1JmityWRzeOo1MLGjj
FHYCyKzFwFilbbS5jokPMeHbB8CmN80R0kR3NVSJqF25Ir4CZNgfBDO9ho3wup5G
dsFkmM4zfoMjscPKMtb1zaTmdW9OXlNY3VOspK4lalzRiCEv3RNjzWfVxroT6X15
ULWBsRKuEJEuV3XlGylQtsfsewYQR4WNkTz31El91cbJGaGD7M3kHumXfzyNXPEU
Ix/OxZldq2vz9B8HH4IaB2BBCLkAItl8HrPQSnQ4cqv7F3EGZwFhD4ouIUY+oGhP
Zx998FaFZNLpBl4bsP3lPxqJESuv6dIHKpYsBM2Y8lAQiuG9n/lwnz/KcBeKCiMa
A2YEPoJ8hQEQh2YoGJh/isjYA8QO1vjcAvmxa2aYDIFrd0+R8hltAcRlZgRoqSs1
5KgIR7ymc1lOdEGq17THqnuSeS5/Pm1QPm97PYNseOtNaA0jtPTEmLwjRsj4qqqP
ngJmmeH4QtpU3c6FWx3XpQqhn/kfHVbCLbdjUieHNK0A+W4s9hrZyupXrYDkYVaj
OGRoNdW0Wfc5vCsKwhvrHgQ0mHK7lhBmzedgkseWrEHZWguRiHiwC35XFf9LMXI2
emsIatt+tKwZWCal/HRljyP7QbhNTGhGXOjqEc2xjj0xlypx66gdadNQHpN7N2f3
tdFz2X+ywrLdaWqr4zZ0sOU/TrKmkGEcaDEX+fivU5X7+0NhDALRBqPfg/NP/Unz
onJXx8tN3W24HsbAV2qSHTMz5OV03ql6IQw7M/JAnMWLlsw61hDw+JTGih+4R4Lk
mpaYCKa+SWirIT0goJqsTcwZYWr8PKW4fxo4y0d1icwunszvOSMPyw+Ttbbrzw3h
SLspEJB6tcyCMQ9rCuln7zeTs5F0OJ2TS7sLKuA5uf8hsusDEU5CYfy7IXQnhcdq
dq+VfldtthTHhgxJ2bCGECnWpcSeVwWlCwK/qPnafYGsfK4RyWCMC5cjNgu/JS4f
zNXCVM/F4iHwEk+NL8XFQYzlg3qIw/hg35djRllgw+6yJIevXwVJxK2p43KkzC1r
VZ0c8+H+XttaZbe4cXpzw56m/OWtnfk0P2qK5YH5FJHSkXTgyqTrGeKLNJDe3E9b
CZkZr5K4yrJHyuRYIncn/qDFUuIe0m5+STqaYzPyqSDSjadgydzw7HE9MI4rJJjH
F8x7ynosFBkw+oKTuvSBVfbdYsaHITbkbW/bPEbQC3oWj/4DnmVNgqgXQX/Ae0FO
aLYSrjtHElJIIiZSWxVn7K5RZlRZvMblQK/oRKJ6GplY3eCVb+zDNNj4MeuVwX+4
S5YKhwiRQ6/JbFcHRVvp1b5R83/FuOqIQ9D9Hn9j2sw/ZFJyhUKcIxa/ZbcemxpG
qf6pocdkW/tmpLXIivRlCUyFe2PxqubuLrBLR74SEktKLUY3fW1WMs1+RlSMYVAc
1vYlUjsVk1J6ZFxNo9kc+ijfDP/A7d/t6u5gOQcPSfLTEWWrYKoxhgYXRUrqmrmo
mUGJBeJwHU+rMKXIBY4gyt3vNnTNjDRlC7RXRXx5687eGUvwf0Ddvf/jVFR4ejEA
8KmwLm1agEczRp/Vt5CxPybpSgvX5iMIvLPkY49cbh2jfGWM4VB5hF/vLiPsyoRY
BMLfBZ+UIMjjV7JYKC+Xub/QzC6FAl1pvnKJbUrBXH2tnG2YddmHyuVmFYjiWLO9
V01SfOG0VHgVYA02C7pu5bzw0HE6wSh4Rxapyu+EutN4cuAibSNbKup1Tn01dWfK
b1d5WVZaZSbouzApzKWVHhhmwmeS9rCu3jLyJg1r34+y7fRuqblBFaYnpJLhxFth
sYKL2ZqLEUJGHhRbZw1A1eFVrDJLzaO6ynyxHtm+cEaLGdYAbU9PE0wMQZcGQedI
MRiZgeNasQm+vbRShs3jvMW8sMl9a6AXhTDx1OepOxSQpMlET7OUhOF93PzWIG3e
XRycP98TtmyoYjik6p5xcEvbzFlpSysQVDWBdAGK8B1uazQ4mOSet8wMXiuofqjG
NVU2WJHG1ofh4eVPId4TgDn8N3gVzMUCoJ3sybnTHiV2G525tTVZGxWdxQv+Es9l
PWQX+uDJq8S+EtaGd+FkXfD9me5IxRhVHTTLhJF4tN/8aUTsDv3FRAle/GfGpCAV
T35JrFDlkmS4mjnRWtbOiG5e/QQl9/n/tjYCzGzFcWxdSI3xJ48uuKzYV1BQ522K
V/49yC+GWZT3wIceUJdRZr7LJteCzpUNuu2jw0WSrTP5oE3W5W+IUR3CReZMRJqe
7MzRb6FcXmdKBs3SYch1Rs0Rj6pWg5TfNRuEwsVDo5EaHvTL6trBttitBp/+3M8S
DFz6qjswe/gMWOu8RXF9iddQjGae6AmZY9OPVFxJ4vcIZ4cduwCbV9ZjbCKwYu9N
sl4ayDvHx0lU+b3xIvxCofRhtNwT80m1WKJMaK7mQPa04fLctxXfsDMkPaS7GEgf
OSLZC8aIGstQ3c4JvQVmB+rhaYAGAeRJRe4TV+5hT9Meo+ZTRLOyNarTJoLAgGt2
g5ofj8C/rWnPI3FmwVri8rH0glbbVKDsUyEEHtfzurHq2wb//Fs5EyFSMYe+F/ip
OGpytmYCoyF/5MybBLuagmRknb++60fvWWmIXTt/PdB3fw3xIXMPyJsSnaUpLNmk
tRPTP2418aiRIoda2bbm7n8/QqSGgBT0yxhf5ARuUrOp9vybqnqID1q3vbkDjZZx
e2oANpjyTWECcyJx667F0mdQ43gEAHGXoaRdqEHUN06R1H/gH6RuiwSN98D41k+0
gQ8xlqgd+Drho/9257tkGarP23zeEGvavSdv0FKfXwwoBYgtj4qhWmk9TdqLnP/5
C8IC3z7BhMysD1Mwy8GO1HtB3+qeatH1Xr9W4opoHb20D63ehjbyvkUEhyc/UNi6
b0XupkoM0Z2sYYVcdyG5Ye7DKlRYp/nAjFpJbH94hhKYG+QLHFq3rVSSKCBKfZH4
8uzKrL1ERNz42HCObRkhncu5kjQKdbmXIoRGvM//RQkgY687TDqymYvPDgEGOk60
NYyXOIldxiZe5i9FRCoKRr4hYV31xOftKIbT3uqsSb82LMrJ7thPwxYyiIoK4rFC
jV4WFJIfiuke3s5JWDd3VAb6beC52LnUazDYkMzsP41NQfIVfaFozHO0UpJcPEpt
MYh8cbewspdsMpxhWLt6tPgwKSd6Rnmzv37fSz+sHgDWepbdgGCWqW5rPh4oaJ+2
jHSQz3gptwoWM5+5AwRnB0n8pTWi23C2Xeeph+0VwEUOxuq8oD+QfNGa4xQ7tFbS
JnYAVylAQPVD/avVWTPCgRlZpKmj5DosyhJ2RuPh40+KtkuyJSUIRikPqzxXyOKZ
73mJwpWDamO34E7/sWNdh2YcLwA/Z2gSqtTA6/MYBcWriCSX/RgjZzrFcALNK63a
4zFrHejOcnn/Qgv8Y4Twz827S9XKv54lSWpBoBm//6sS/ae8WAesm10Jf4kJYtT3
eGr+j9L50Z92liBv0VfQAqKihOzGgiWNIPRcPIupuGe8zz/FDCieFhiBKxXqVEjP
Bo/a6piXmp07jXyYtn2ZhF/cAo8rGDoZwgZ0mZaooMBtuJ02j8ESwbvaBUfp32Dt
qEdfQTlt9+N622MDInGXMz3wdMNINHTYLdFf0LN5rA1cbzz564as0XFLP4Ni5D1A
KuIbCsLSjxkC1TAkIbLfUN/j/wwcDH6RG0iVB/Ft+Yd6SdikvjIeb64yB5pVqOSw
rOISX3KvCW6yzSU4NTJQot4mIpwzWd6SHQCMPsfJFNcQDNg6jwSAyTYO4YyZeiCR
aJOEb+KMHCB57i1bBwBpTf5ZVaxFBSJ65bfqwEdE5tHB1BQOWKHQTJF5CNNVh06U
5nZ7ehsapWUE7N0atftIxd9rCDt7Stnzya2q/ilJIw43KVC7ETbrHCZfkkK+Er/R
Al2uNVicE6iIQ4hHVSrlUHB2+ypzz6wC/Kbcnuq3/AQFNisoBcc5/bykAPOqMUMF
xpX2WaL3ZfqD8fvuMbwJqs+MoCsb/1YzZQa8NiXM6cyzFXsIXObQJaoRLTNUF0Ez
M0kpPO5yJlriZWH1Oui8xE+KcU/7jMUr3dscMISFiDl70z+yeTJjNRNHK/ijbvDb
wbt2fHph6gt47jcROT9ELBgcVk2+IAOZMRor2Wu8cgy3vRF67UOrNDrjZuSCfu9R
Nq8PCUiYlGj7e4MmI5CDffmQ0nU2wEo4gzLdbpLvGf2VUDb2V6+xHwn+IlfuWsRN
wlFevnzHZ8unx3ekN8yZ545hFNhGVJ3hKlM1pabn9mMoDjOkaGjeWm1roXTfKm4F
lP6SsWLs/L1ADKjHm6IZtYzOYdKR0jPOtu/DF6AbUFTt5BCzAc9zVhJDjIS0SMxP
Oen/SG8gZMRUGVBb3v43s/mgiLilsAXBaDVc2fjuyYtMqcVaK36W5uvqWs498GHF
oIMrdsghXBWGfmSEyxmtr/60Q5e7SExC9biLgvFXYX3VdGz7y1VUjzN0nMCA6+23
ZO61NiOlP0P0jXOaW0+HMK3PXjq6GCDPK/xQsitu77ufJVeq0g+DBpXawKr1Kh1j
pYxV4tdnr/Yw4gQum8tv4u9hp1C7Fdbop8rnqXaMxsFyrSamMDiRC7QKefG3NwEP
izZLpKX+8hQBM3efdnkHtXHZy2iGuMjWnBYIH5M5Lmcb6VMtiFBIOvTOyxEuV6Jc
VPCM0ldiP2z3EQKSOytr2l57W6xa+itGCaQ3W15xl7xSlV/N8legu5CKP/MyigKR
OKkN1XU+PS+mcrLg9v7JK+OT/MS6O7GVkZJCjw6tFixbidA0DW6accZ16RO8WnCK
oTaL37yz5UrRokHXkhV+GL5p1zhIQTp2mKHWTw6JCVfGoyUpZaYB6z8+abXRsV1n
NkNA7jTbUlYso7Z7Nb9Z1/E9xTmZ/kOznqlD0bn7aAoaMwvRztCmWAUxVs6F/KS/
URdZ9n0/HAN+EuFiyduR7hCgkqr6iMn72QKVB1+pXG9tgL3QoKwXD3IMk0/L/KgP
K1rScG7Ed2WKdsgZMreF/34de3Xl5CkwtFEOfYsy99HAdyxH/ZxM5QIgakWc0fiU
V4SBnR20I9BOfD3eMLRY0t1JQwHvPD3ENhbb96D/6kMLzqpUPDv7E3U+TCUk6WpD
EeJ1zuQ9gJsuC/v3Npj13x7RD7cuA7PA/TsyOWXTOt6Ju91albiRoDOBDEV5/jzn
cVT8bB5Uaxuo8gsTD4miFTgycnr1txhcUm+Zv15Z+ZFTLv34H26kqyIP7t4/29zD
4z+NgkOJ1C84WoYFywjJVx35dtDo7tFYa7aovCmrtyWGDrwiHsEHf0yE5XVoQ6OW
i97fVLC5FLQdbnGGucy/DEJQPNWhVFw35gEPDeHLDyLhavAtzP+gc3MqrdumB3A7
0VHuJyR8Z+VHANxXz3tPiWNouOAkfaooCyEQn6AsYWN97JLk/zYpTMlc7LHWFZ2j
48ESIm2z1hMwA9lG38OCNXq5vlpH+1dzCoYvus6VX0dQFV9suZZSeA4aV1WiSklP
4MAmSnUN0VUcEUoi8MQIocN9cd91f/JN0xQPSwjAnqbZfscpZAgxv2N1bOKBdqjG
5JLJ9G8RgGKa9dM/qrOETIDTnZOf3nmmhNIbjvIuz7BvLB9yjWDWcXPibvr14HMR
vW6VKKd5++qVclFNPn8UoNlfFL8Gyr3RvcSMKAdVrR+kpcX7ccx4wisE54Zdbynp
AeK64q0OP9xLh59GF8E8OJXQag855xUNJ7NljjQabHhUeDj/gqg0DbASDauBKn0n
4wFHFq0T0c6wIuLaJ9OlaMe/E9EL4bcNM9wtbt6mvO4sLAphJnETw5gCEcazQBbm
fF+lVy6yXH7js8vggbreC/9r0Mp3Rq/NqbQKp8RqWv1hooKukbwNgYAYU/Ddqeig
8hRl2HeGD3wcqBVvP5+zFcqD2IYXcCMsOOijjwyLcI0pgpKPHWnvgRAgsB8+FGYo
5q0JDurblOg+mkLLX2z21xhaLxHcYUhaytXHwOr3NDOTcYpi7deSNaRJHolZeDfu
wUwGZVtpR1hjkpaz6fr5EfHjXHFwq//gPZChSlNwWWZ6wwSYEERrUME12TNTWh3t
QMvfRU2P+F+CZZK8fc07/uyoENe1530A4DQfKeGOkEMSPGenF8Sd1BYOhRkmVChH
boQGVvFVNz8FAA4AakVGPLqTNQmMtN4k7bfbseEzjnF7mIt4la6P/Vx6HMTjXN3Z
k5mJlBg9ctoq9PuUleouiYZXVmyGOosusRgDh2o5mOAFJLwsvkM5sOYvT8wg/i07
m1GShW5J00c9ZQbKRGHO1NDPMdGW6XjRNlLRAzmBONF76HmENwHyNpW3RZmAk0iw
g9wDEqvO45Mq8ROk74cnaJCfLvEc+AvGzqBvrOx+0qN88EZmFCWj7PIsust2r5j0
1SKVbCM+GdsYiVaRT3ByJBK9ZvkYiOMF7o/pDPi1PSM6FJoobfDT5k98Pax8uIaP
gnUkLtRc4T9xoFNRlLnBw+Qa2iQhWpgeVPxLIClLPF0AuCwR1obbQPjsa20avoMG
ER+vtCYyrJOSxlIOX7iqYJHYrlWrfNN3G7l40X+sy9emlUPVMfixNtZdynDBF9zZ
k+s+x812dk8CTvn3H32GkpsurgPPcFI0zRCUadMbAmH91bLJ9f70KUIzOk4VwgK+
PmFfWBvzrPJYHcvqPE+O2wOCwdF7AGa5IGzPfQID652i/d1bVxf+vAxSMo3RyymT
yEbB8Jw0hgiAAdth+aQX2DX45ykrDPdIs3RHgTGnU3cb6d4l8I+jI1P1vsTafE3k
igm8qo5an6HDowd0/0frtRhNZpAB4OcOwFJmdV3NPS5lQrbTS/HWA5VqRmRNsaHV
ftQ4kgbN0DznG1l7x8zW6oSnNjollcYMwZZvp3TqCbcISsAxQygWdNw6QvN5AbM3
zAuk3aHaa+nrKoj1ifYdERUVOpgsZq0lUBscN87lZtvkB7dndXqgIVM4SZg+NjiT
nIk6rRXcTEYd2f1CAgJAmmbsggO1Jtb66bT7n0Xdz9JaU0jxjjmIp3mueZoDuSsE
fO72eLUq33CZmXDfTVfxCVIMYOIDsf7+DvuyuSpbLt8i0xTEs2x+UIXPKnUaONr0
g9EV7lbcqnxPRmHjjyR9OLBkVCrozUnHEMaSfyau+tBEnVXoDjMNnfj/tRlhWiid
cQfgPSSVPY9Va+rLOihtbgRD3CsAy73/Tp0UF9U20S7SIh0P+bb8rGCYMjdjU4VK
LOnsEG5kIz6UiAfRwRyYbM93gEdCf2DezqHnQ//70CvNkJ5WW0U10lZZReMB4xb9
lMEjIHpGgw4mAf6CD5vsDYkg+fv6nl/vfsnScRni+zn3Scv5R714UekOw/Famekm
SYXsGV5pkj7g8BN/MhoqBP7J6i9LqAW/+/9AnTL7XghVB3FocaPwOy1VF/6eJjXX
OUpy59wfBupsZh2B+iaLBsb1HZKRodwA7NmaPAWWXQX2nMYFI/+HcHao15uK1y1D
hLYmbJqw4Hj+Esl2I2Tk9tOUL4y77YN8AeUvn5DV3C/0am4xKb15wZ/iNUQoa0Lw
zl7Od1oLBWkTgKTrIuvfYN/4MtFnZ1QszCOA/cC/kVsaEW53WUZH1GShVzH4ukkM
G2lcmCbkVDWAZS242jYEF64uHOiEk0DRokp67A+OIPU/lyydVlN3czSd3IsIN0AS
oI1TrgTHucZ0lcOltAdoNR2yBSlgrjcgRJaA83YpeaWIH4awi2eIEpXliLbZ2cQV
IvZi9AOeg2+7+lMWqdtso74vHW2Ztnctm7i7Y7wxWkdyRVT31bABxd5RWJ8hLx8i
4MzZ3uotClCVYqMCF1NB/LG32rp9z5laTyO71l6krrIk3AQWjZ6nNji6H5/EMWe9
67LBdyCZpAGY4F2GCO6dU7w+G/1yZuHPS8A8NVuAZPIFTuHTh3JCnpdYoiPWORTm
cyvV+YhxWbReI0HAvmO+BB/yQx4nY5COIFfGHXiV47ZTTbNHptaFNP5rBNDJTp5a
FAX6IAronqJ1d7vXpnMQ1Ekqpg45YBLgZ7n3NpggnjcZsSs5DCJfumlkKG1zVpm4
GR3E9bzySYj7DrjM3+cP+OYECQUY/DGsspWPE9oMjJsmtnsDoviB2dU4Zfx7261U
pQUrzv8MdkvdYGeefZ5uixU3Gjph4tszFHY8zn+X19Jw6sM+ns1cOmmJ2Yk9YyF+
ArWvxRR+t3Io5nRJHw5JjjciwSBaXRtRSSXBQmdirYFaIyhnXmToLOhCNDN1qaVE
bTJpF91GVclfP7aYTM+POInyBbaLhooxvwIauBX127TVEGAOOEjbo+r3F/D7LqmZ
Nxv9ehXKqN9MugI2y1X11sEoMDuq+i9T5GhWivqCi5bv8X9PwFfqKL7DK15Bf8Nh
uPEp+0iakfM42PKstdrAY45yMtF+J3h9orheVG2T/PTRUKypix6wcOtrmwrSgrdG
E1fy83uiePB9Jpqk0Np236A8RH5aK56w2pHqMTXpWDCNojxIOahx8Aj6Nx3vKml1
uAIylcMZHxOtyj7v14m3XmPlJwKza97daIZVIWnYmID56bed/UqTZfdKo0C1JkVN
f5V265XcVzl8nrici0C8vjSeb+CGJVwPZOM0RhMJU72z8ik6aJaxF8B8rQ8smTos
0NhsIdjym770QNupmR/GdN7r1EFuAeLSg31MWROfw909ND9BQW5Ltykq6kyLeErI
eXkbX2DsCKEaaJO0I49Ds5Qx0H2sfTqxE4SPStCy3X2D60hHzMP2xfw1TmvTwluH
7vXd9Fh3ewdV4nkjJnZsVA0FPn6vLHRcCEs5MiCBGjttM7eyjOc54fyVwoMWQxbw
n2qQHB95eVmuKxhqO+5TGS9nNlidJTX0UEKXEJKKrkBLuqe37IQzZVpEgzCOPBP1
UsEGh6ZE0NG5wYr/w0jUGmVwHGEcILmWMWGdQSzKEjKf9Og5EGQGOE5zFgGCggA4
zjpc4QBpVyEp4iQRah6obzg+416I7s+SbccedhF6B9/8dAWJQ8UWi8gs+vak5024
buVRK1KLhBWjj9tF0OLvyucWTZ16l7nTIT3UNcPJF/edk8jMIgPm/BNkSYo71wJv
Y0iGOvTfpQNnauKsFVMY5G/u8JeOCdk/ft2LjnjPmBok3DjQr6dxpUNaE5I5kIE2
fMTsQ/daTEZxXbX89x0aXgPuvnfqalHsjLE30h7OMTYQHKJu219L3e9Nm2PEv7LL
8bMD+eBxSJcFlD0KgNIpB91tFNnOHPxAvSg1ONZjphuYuov4Oanw5titxLgtW9pS
gYb150OTLZzPqL6FSUmKJDgpLo1KU1braicKyFbZNMNdYddpgtsnPiQAd87rOIwT
mGl07seDCIOoaNs8Te9SjpmBUiVt7lEKduUyIu/zyU/Z8GcqHt0NZU/g+iH1XYIq
B1EZ2F7L/UlqMScDnEnlyeHcWgVjJsG6jZFLSdTPtGGGdfkK+Z9zpTK1bb0tFnrz
LW2VrObD1reA8IRCWrVGW0jlHlJjsgY0JxZl5U2v48WeOJW70YIkCqMX7qRIrTdg
Oppt/MQPigBMekozHQOcKYozjkJYaSnnTgK1uOKKnL48HKTrmhNSBOBT5yZscBWJ
wI4zNtxz3GeZKIqbY6MFME5TJkuOoZBUvPxLJfUbwkxiE6QpFk2TsxtrRN7hxSrs
el9h6Q/RSoyoQI6BFKwPZkZ3bguUP9borNbPVUjC1VatAxDHlclJsIXIQzoaNZ7v
XgpHs/dIA8DjXI/KG3Kz+4o0/+YFyYwMO/SL8Y9L6dPJ+/pO0lOlY4Ra20SxbWST
D9/+VgKl4bH0gRkf1p6wzFIalkNRzGwprTfpeR57/Xb7lrh8eMT5iI13XKMRRYdg
+x5mN4BGDuAOFglqUeHtmkNa9o1oLCgFR3Usy1S6xzPIEsyX8bn/yLi12Mb+oi2C
lBokAJ4bH+1Y0o6syQVDZGSuxrjIR4Yl18F+b8g3qgtmaTivrlgvnGMkV0u5v3t8
eNC9fPbE1HErBkkFV+ju/tKu9Ps99pyY0dPge8jqr/+rzzzDJe8g5nQLtYQLsRdT
wgR+XQ1E9kRKUw7RauX5u3eiBOVJxTAHY3+apAomEI8jUH847R4XuPNXRAAttfaL
369zbc452XHIh0LX1RhBS3A/lUazF9vuoCqP5BS6PnT/A4fcDOZEsN3yl0GyERni
C7R4Vyl4yMA0ZcsSOkqDB1M/q6nWbgF3lvBqCii//AhQYrcFHwf2VvkLNcWcR50D
Q7q9ifMBBvScAoq81sLP2aGHt9a0qo/EzFL8LMHKcJks7JT17mOL+dfBFENHffF3
Ge6uyXAnCFqv3cGjTUMOD7M8Dc91CBIAOcGLvE96gV9UEWhmEs1zR6XVhB+ZhMGM
hHENk4elzEERw0WND753uTUxUqMXifT5q5SgNWlPZFJ4J31/KcVsJl++3kLIvEAc
nnIeAJBj1+6Cm5au/rv5HhOsyBbBl56xUgbU9lD8ythvcv3EsNFG7C3IZvvxObbW
teY/Y5EVauYkGOiMihKbFsVQuUYlmcr2oQOBqKLoB94BqQPFw28O4JBQ4D8/7wZ9
JbHB8lbKBH+y8AiQ88wzwpRAqCyRg3opcYWwcuGggiwgO+F2kkt6F4TurOZB4+UM
b0iQyztaOESBKNyVpoe7EePqWpl6kDD87BgNDNbU/Dp4uX4OiQKhXnulJhJ9mXqy
nczk3E/bMNOZB9UijXvdpKj62UX4oUFqESPbXx+eNtLWAoS+SczGpdbTXYQUny7F
8nH9ev1uuuvBs0ORjeFgTBDFE3v6b3DKwnFHICadhMgd3jT/2ZKrsPnlxRWEPhMd
dPpulQSfPnxlREq1UJkGIiZA+/3cZCzok/WfXrXqnKYRN6n54m6hsCUBvZ/XiSp/
+nl7VfsFsyEj2ovBNpNeDzi8Ah7I+YhqJEU+8nyeRKvQpbrpZ9sVZgUwiJFDzko7
DgScVs+1djASOX4rxqSGIQyT6ER8sEr1nyr9Glm1hBOpzFJKz1pyif8QBMx1eCAd
68kCcRYhbDj0UzGWpyw7WS68s1oXVfbr3kQ1p9aNVacMZ1mK8C2hwUQGsFHUKBZA
/ZasNWop9EuPXGswQoUsPBG9M0r1IZ1N5vAfU1pbYkWGcrK030wrXQrcIHSuJFVj
OmINm6NI2xNPr7AtORybV+FznDCsCHrTyR4161xBEYQfZUtpJURXWPgqgXrpQe4J
KlXJOpA9f9PP1xRzFKXVo/mHqJ4i/Hl9rmVE3SDyEx/G13Yo9O5/JWJGppwY5gNq
IfGEaXaBU8pfUCb9C5T7BaFfXVG6s7UtPADwIU//xM6TR1iUJvIQq3BX1YIqbJ0g
LuXXBnwkRShSQlH2ZgeJyQKVNXOcnKxr3IwxeLs3SaLJAA56FYP9BYLq3G6zjU9X
TyFf8rlFLcOSJm1wVANWaa3zhI/nHYTXcvPajYIkOJCMfg0vlH2kBlQkBCSet6aO
hg5w4Cr8haoKZ8l0EJVvu8G+qxSFMG/fhUACkoPVYK+pJb2XEsRUKR9evMtTZ7Cn
o5MElxWjwBKFU2FSIIj68qNaVzgKrI9eCvKcX1e6fHsrOe72VNcplhbPP5LvNBth
TkYd/DvaXiAKq1cLlxhmaPogjIR1xg7a/EoyJQx0+I0gsXsxiEFKxLpfn/aG5M/o
D0TyD3VXH5i1vRx6BYDRGK3tHbzk3oohriuOLw18vhLkTHxt8cy1K//bRw9KRAtF
7Q6I0FCPI6Tr4Mi+XgE7RBe9Kxx0y7fCsjHDoHbNnp10bd5UKpfHHDfc0zlCfqhk
7fo4xWKfPMAqURODIG2Gd39/Powj+N/za24aKcC7AHetvYm6eVpQon1iBxIIXYyT
upEfJted88N1vgQ/YlWqSYHCf9MXisg+8HSWozojvOaQr6jNPf7Bes1oJF8OxAub
MhD2ixcf2sQZXzh5Kjh0ffmzi+XruhgB2L+QI2I/MLsnxxSlNMELsq1ohcn7+5oG
vYzcgW0c4vZZfxymRQYca6ui6Inbrnjg8yCVaxkqU09X7JbeL1v62VOFAfk83mTb
2HHoUlz9G83io3hU7pdNVE0bewTk7srpxPfGAO6ohd6s5LEOeOBGuFzVXQADWwi3
9Mm4WQtsHrBnnhk0v+RvWBH9168j1DKpg8RZbh3RT98LEGDaC5PhyiMz1vtoF8xc
+KuM4k3INabKiMAQyy0PMsA8EYD+fla3RxyNzdfm1ffooC0Hzt+n0mI5tOota0pi
PY8J865KclO5dccqLyTyMrkY0s86n5J+jrLEWz9WedcNYmswf0omwRUO0XkzDman
7b4x0gb3swwbIt2w1PVU6+PbmtvQ0M2dsUvIn8Jt8m1aOFAiAikw9N1e0TVh/nX9
K05HTatCFbtPEKeQUIb9z7epVCdLMBJHrMlINaWLXw34KL80EKAE/U4lvVsi4E/n
loR2xw3YaS/2uDswfKgTI5tSv8xSgj68LTpK73b0/tyioUvp6c6dgoE+byu2/I0H
QArUIz6nB2J0h5Z0UFFgDQf2LCk8ctdxFS1Q3w3XOXWi76mKIO1i/pTU6wjjrpcZ
EE9B+5dAFstMmBOSXWMMF7FGwJYuFenY+CxhaZl+tj8uPVh32UAe9Xmvegzt2h2v
qDF5WBFlgpY7EL3TWQLfFdcHzb/xj2NJYWB4TBtcTyaUeJmKYefa5VBjrihdIvWM
22gkvbPlxrilJC1jsJZUUlgwpvUH0Hwx1b4rKyj7F9+ErfIYVfRaDqpX55BWXtUm
RR/5WZrH13D/syUytg+pyFF2zAiuXiu57PbjcisF9mFxHkKXz+vN+U/NGiSCro9q
4qfD+Is09InCM/Taf1uhV56zuJKkfSG6zJnOVnuxkbe8+VvbUJ1fwGS8Es2IEbHb
h9URRlHVDUB9xvoZY5IenuRs6wCOdmSHLgW3ooDjfkNyHdCD/ZOyrTPS7dg7CUSp
uzpjIUow1jUJ6KvAbFANQ301e4mRNgwjbmHoyg1qqB7tzaZWlcnVsRWEY+MRQjRP
Zm1bjLM5JEaB+VgBrhFnzoWsgQVj2yAcBkN7JDxGAepZULRfLs7reTxLBrZ5VTaY
zpSk7GqEW2VNIxeltHsdTrLzOSCWg3CQZNbrC4R7kfyV8ORZ29Wp+kD0sOulEbke
ZpYDdggjU1QuLEbiMo5vD/HOKrv/pxfyGbANYqe+pI1LhAbO96B9tTeQkSZSxjD5
o3SNnduZ2ujPriBA7q55YIsAW7Nj5swobEeKuha6JJIXK+FhY+6N9Y3OCUQbBQdi
ePBTnutzuj6p3n3a4YTaOP1dXRu9g/S09xyeaWk+gEhojB5Jf/uuMUfpFjxLKNQS
zsLn7e1eY9rfiPmv45yzpmSQZuYwcYNSEdm6JY3LyUwR3ccNbbZSISdbijkpoPmd
2nwOz5Eyn9oNKHVT/DRqGVn0F+vCeh/fQTG+SA0UbHuM27cUBTpItbAZrRTtxr+q
Qxlx/3I81x3q5eYjGp1pDjnmsjiBZryXi6vZeZ/sGbOP6sF1YemsuTpwNYRBpnxf
IqgFk+t5zd25ESgRZI9HcS2vxqORedlotEsOs3913mlVEspUnrW09AHq6+U67KM+
TLCpfytouVg4/TeY1NHFLCc37V8V9X5iN9VjWVG0ZmpEPb+YvO2m/jWfA0jXqBW0
FXiIfPX1Bk6X9Pc7msgS1lsZEKLEWRY63DKjzCJ3cKGxcAjC3lMiAb9ToEHMT6SO
0THrR4/wFC1BjgxoGONO4zn8OsXeis0O+vSsDgDRJqtUjFm6w+yt3mq9Six6fcUb
nDh17nix3AwNEpAtZQF1tABrak9WVpNvtyGlambFa8STyZI4Ke3BtEjQzG5ahOqT
w8xcnNRolMPmp2JZLAB5N97OoLcbIq+tq/2tvOgHLmZ6m06Tz3S6z+ZGTB/wHFXw
rzarpoKsotJFpE2gdrIqJyWT+FShP4M2tvVdNcCua8MMVR3WzqKUG07i3zFqBowt
dZbkdF5btLIpptw/Vgbf13CALoe5cKEN0JBYS0EzRAFYhTyaamyyMdMsVOQCTTcp
ZhWIHliA6Bi8VBr48XV/tsoqKGZvFTf4G45aSNk9Zw3IfMws5LjUXvpi4TbRff84
qgzvMc/7MlmV/uaLH2j0roIMbeHOAVSrGFxDb1a3/rVL8PBSEfFiI2SJBPOPdrwi
TPW3yXSJgvl/645zp+tnxtGksmE6YT1fLW4zkWqgVIoDaOP4YTmAtZvEZJGLuS+J
SUg9TMVl8FMhuZZn93anccbZ3cT2/uYIMHQXU45nsDWjwpdpFHZs2opWVUQxxm0x
cCO5V1JKVfV55BKHdgfxd4ahNw6MY0MUijeIqj1w5HImgvMqDx0K+x95fg4ZtyXf
OR4JXhloucTwLxom2kukQDxH4iUQPP/DrKqyaEn17XSuHzQc9wdU6qfbEFpwd8mb
QJIQ5IDAcQPbV6VVmISnXuVYN30NkobGj3TtkGDreIe1QZ5XBwUpgn5H4Af/hmbm
vrvlsu+OEx3nQWM69KW8kWwq9Cy6uShzlx8czIgBtBmnKzkRAt7IgnSIo/GpzqX1
CNTskqYs2M/OxPKnnqMb9Zmsy4+9ECgHA4UrsuGKbi4e0PCI2YA4mmllAiIqsd9z
7e9EgExtwprpkMFjkvkr3HGz0x6sa8a/6QLfG0ok6p2Q4tJ/5ttrtUyYT+rrrlJS
PIcl+1RaBYVcuvF1hmAYPnN0BiQd0ZtRVkHbqdO3ygVl28+lDuQ/THQSAbZ3fiVC
ivPengjApPmjcjOmy9ixyCrwxJyUv2kMykwyj2NQ/CXtFQE97H9NUlTL3GMl3G8d
35SnVBKKeIXTYuRtaZTAA5L6b+v5DaqP3hxHNdRoF+tB8Pq27FJJHWdPiti7ube/
THda/AP1qUY1HTYnt7slQ/80ac6O3QfI8UdiGWs4lsz/Ev7vFEGMaVUMXI3272/n
ip1EH7kaTr8iVcS13qWpzKcC8qH1ahKOD+FJEYE13Ld1MPxHO1UJi6WBq2kBD77Q
ljAqw19/xIHuODRrys/Ul/cMAwYdjPWenBGdFcFgXrmeC4765EAFn5aqVtpdmNg3
hTHA2Ok1sO7JrvLFPFH87ogTbV/xcZZU35WFNm3+IHl9CCzwDcli+uQQ0paaPD0X
V1amldYPHeL01QErITZsPzfPW0oLwxXoNSpPMumlLUSJTLkaYLBKv+9RWYG5+KP4
LBc5z7McrCBDkuiyAQvP25hNQ+vY3iX19xs746xRKOTBqOPlen2ZVGVC7SKBJiG7
0kRi7SDgo4AL/YKn8ntWiBlbtMm/74X67YGBcXXxoot+U5mt7QhPUW7ZYohetEdv
GbfR+l1xo8HFUEhgk28eNZOLs+83aj1j9HRFK4TELG0x1S/0TE8oBcClh8lW5clz
iVGkV7gHOe4LuY0SnlBAXyVa5BqfjM589M05TkK8vYyhCR1RebC0hVrTeV9LAv+3
guK5Na83l0HuEvvmYlP77ZFsRJC1Rh8+XFftCa5/UN6xkfi24fFRa4S6d2bpjDx7
HOHpHk4nKJrZo2bcxp0WnYqDGYL3dBaMb1Hjug2jE8C9Ir3D5PkcDHMsMfD4ogU/
uywXNg+C6jZ92VxLWCAAmJRe+SykbSdcJhcCK1L8MsuuSIK0qviu6+rb1cX7kxxW
RDZe2Lqlt6c5dGzdeqgTOkdWQilr3DakG0yduaw7oMIKEwjpuGZRDANOXwILigme
/+xUVpi8o3T1HomIAgh4zrHsYmi9BhaKLpQ+9fQge2mxepDHKLFOihuPTNpruLrg
sXpKYxakWBygZeCzzTWgKyY3b6uFg/6Nkl+Q1zrrUjvmMffADVIKz9vM59I0qYet
bkQhJBxgKcSo/o3GYxV429A7xl6pLumuzsL/VLMRy6ShANR3Kubl/GGYS6qyAqad
QmY7IALjwwp0PCZdPy/v8b4SFshUURW1ud2/Brwq0b3y8wv8n6bWlyEr8QoDSgQ6
MXG53r8eVOaxJAqQT0iAlgqOSALWTWaQAuN5Jkmc5Y8VkJ5akS69401IM+y6ufSx
kCsBYW05Wh9TP+7FKTTT0ClNFxWhUfzXhLdwTgKf3LmOj7j9+YaCh/OtC5lEBSeg
jOwXGjUeQEwlKhSTvH8B/b2jMCjC3Y2xnO0b8amSrTY7oIBhbAKDtztlFpo4lQEP
kjbLg+MMuuMAE+91mjmc7LErCeCO3Bjw859MJglxpjQrg9sUj375BnDfoyLF6OP6
wBFvD+8au2YuIuq4JgTLxSh2yJNoZXn4UuB6UeDEkWLlTFiZ9oCeAyXjjWM6O6Tf
RyGD0rT3jG+z1o9OF5lKuB3xDo3AVX+chsnQaxfipgFA+PYfI5V8zpvNwq+GW7a9
hsJbqI8FeqgJuJ+PqEvCPJHVP93WHxL0kUfnXimKs2TNvtxDKQ1He05QtPsC0bkQ
6s/qQoEYfVsfkbeVzT3Rs5zGZd2x3VThH2OnOF6jYuU5iVpHK2zXNyI2aNAMSOpP
jScxl/VPNCdxbVSV9CxcF+0gIpR0G3/meRQAgZLGIsUuVXoMbAnB3JhXuSXCnXju
b0n1EqY4m8Mjz9s5OztSQWs7aX2/Ik1p9Chm3QSKWOEzY4XnH237RO+I6SAZ9ftl
Oy9XG0lJxREaVv9Ww/OugYUx+hVENMQLyvydA1cSxLilhUF8GAVWMC1Xc90Cnb40
tKMx1p0iHjQNjaWDUohLMRdOMIMpco/3HK9+bJBv9bfkhEk44ZoOs/617PY3+Zqg
OvZalrZfOtiiqqyFHRzXefwmWQL39MqiCmjerwy1C6MI7cU/tI6qtWueGqzaOMK7
2u7iga3Dr5h7gmlhaIk4x7UPM6855OCS8volnz4NHm2avIq+7pS3Be2xl6h2F7o8
RUF4hGbDuyGxeQUlYBNaedXwMxC4WuIPWfw047GcJapn+iWo2yAmYLbMTDSikX2P
w8MsT6CqTFPAAicPpv+86zuP92iWcz/bBtPyslCoMF/0pMWeRZ24oApsDsgPsphc
c2AOAvCBF/E3i0aFCE4XPJsQX8QsREQ2uc0OeFkk9cSrcDe3U09ZsVYHg06XO/qO
ew84m9zQYV0pdOq3uyMJV0jyxEP+6kW+nUP7qUYAOgn99twnhGJoifCNDbg0DPPv
ViglseF6tNskbCO5mdyH3Y7Mc6l3dmbpbCuXD44D0Wxj3r5ktcPuDm7Yt/6mx4H2
vqdY74MNcYEnDEoFWjXTDR0p4P3NJOCDzI1bO6sLR2hBXU/bq/11rFB/OlRYAUHa
DWqCja36hrufx165SmncjFLFkpYh3BJovS4bt7JCy2HIv0weBmYsQB2Wna9GcbBB
Eud4fo2WvWJ7hB67XJljramBuXPMExtDSUMQqpxd06k40O36QmVqHvc4WlEf+esS
eTO9v8EgXxqdtDvk8NXWhJ5MsPnnsBligEiNF01RX0qhggk05ycx2e7lFzOhtgTs
MzhA1OTMpjgQl4O7JbcDysMbEGp5xGAZfmif1NrB3FbkCkLMLqdeYRRJHOL6Dy0s
2ZvZY5DCO9d4IkgHtvZS9GkSqfsmVQJM4I961VZWBTUK/O718u/CQCY351bLbMdq
f9YMGhYABCSHBKf6jc4hEuOHaJJ3sKE4pDzWPmKUUgo6o2jEgN1soBTASGQqj8gV
Epy2WEKeWeJDfvWm363KNcLjfLyE++Y6lI8/tbwW4lgMGSnar+a5VDZC8pcLdJiD
RW6U54coY+U6R3X8dT+3LK9FpFQTKvlzURhe/BnfRaNPvtp2QvnC2fVpMi026muB
Oa3wb4ZHUMcuPnDqePPAVvwXksIn/xJX07/FOMjnOI0sB+pFYbu3iW0jpq5RcZ1s
4FJSqDs86SNilovPyj4wJOkvnPb66rsTDxyPElzs7/mirgDDPhqopKmhNS/Et18a
qroNNP5E15QB9GrQ1lsm+RqPnXZVyIqFsl6uLsG2B3AqFyRNuSbaFEVFuL1xLIpI
IpnHMXW+Bw822EVx+SnoJL1tzReK6uooF5TGrGma7atZqe1qg3ArI/FV2Jji0JLW
wvpIFPu4MlFicsXgYBw7uVh0id6BenY5wiCWZ3xiz2hT67Fc1jSkk9GJJjlJoH/l
oKwNegiVPGEGP6wvVNdvPCh1iTghd2SGbQ8Aol6PEq0EnP3AQMvzTxRJMZATuNP+
tZYviKbnny3ar5Re0tfaD0DoXJuV0etxp/SvXvuc//g8g/UE4EVBHcU5xNiZ4yS4
Tb3tCeDp8DNUQ/HmapUiOqS9d25QtSewlW/V4Sv1vCHbRPqsmcurgujWTR6p02J5
gfa9O4sVZDUykWp5bivyMDypAzlHaqv/uW5aLYf20m5A3xyCKhS6MfsT4AzMGoVZ
eTFlv7yLSUlyRCFR5L0Iqo8xGzdJIj9P1JbTnPW4iRK1PY1ntgBqANTD1IE/dJaI
dlDeucXB7qKeheuLbHWASeufabtQ7My39BMmZp0ZB7BdaTPVMzplPqm5iI7e/0G9
9zVtpcQJqU126s6onN+92wl06KxrYsN/VmtU6Rqv6ubQ3kKzJcrIQNRAl/MOuXqY
G19rY6mP8rAOl0RQvw/+SjDz7ReK3T/5WGspm0EImMgn++LRQASvoTsc4oRjrmB3
gB7SFm8BVCPyi6vlD/IOy94eX+KvltJ+jefwI51z1nw4TTlVspkJh+sDVC/taGaR
yAgYsN9zeXKMKKaXbb6eUaxiP+bpDX/PmvO1JCXffpTtJjv4r1+QPQLN51GasdcK
svgrt+FdZuHQBdDCVHMX2ZX2s8eXWD4Jh5lkJzLwYoNZQhhLbCboYo91cWoJ4P9N
I9hJalpXkC9rGAYpu7Jw3gbgXM2SwIPpx30WG0x/gursckMteNZsbl/KLiKh2UWm
TXy21s1HMcaXqYMfp2wUysVcnTNYYsDx85fYaLeDedkIKFL26bLbZa9iGHupwjM6
EA2LkwaiqQsplKfSDm0UmTTIePF5rbO/88zQmYDdOzBlLQsdlSBcGO7CrhXbBuBL
wY1lf6mC2UY6cAsvSTlVx/cJ1SmZFg/MHcaKrIlCRCJbxwaQ3tm+aZxNygR6CwgF
ZIDcnt4pp92WXatWoqRVnyGTyYu3nRSohYhifqU2OS27/QR0068poJ6kat2xh2CA
d6FDonqiGdo+Buk5Pj3k30DB7rHVt8MLP33MgWCklgZvbyC1iag6jHRHn9D+Ov3O
02HSrWuIwtuZb1V9NXrQwonSFT0elV75xCQts/Z3k0RdeYnOZq33TvSOCa2q10ZF
D26nqq4+7BdSuq6NwXn6javh6Vyvz5nUxAvAYeAY3+DQQDiCjLVoAQlkUVRKP/lr
PxiDRSuk4vNKNksXcfjhHgDTgHKGmtbj8pTTpO0P1Wjntb6Pa5qPPUlO2RVsTRtN
Qj4JfLva//Q9k/y/isCBvri/kIWkeoRMmNOAb2xIfnCzyYcRWFfQ7njWUuGgfS30
oFqTil6FtAwNHeMnB0wilDX0hlIzDKYrLADU1zkrOIW+n1N7NlfnFJ/0hoDjSQN+
4TwyGxP2BRsoqA7rrl+qj23e5OTK3gRotawOopeBX0nfHH1s/3qzUVThmcHpJ9xN
XcUDP+ISpxr5CZgHTo61yNwZwr3vWclu/XcpXdKZWGOgp95XtxgpU7jZUD8qYAf0
kUxwQLozm/YJvBlZxIE9xroNWs7XpmMXRhkZDEBAQcQzPDXZVHKC/cRk/fB7f40s
tG5vio/67ZISUrdlHCwcV+4+/HJX1fPluXXPmupiau0jooKCW8J0dnwuuvxHYudy
+iG6rRRM9oYtDsDfuxw9cw4A/PFxGDwfV5cD0PE4emw05wZ4Vy0XJPB/jEvs2iJm
KGtdAwITt0F7rhaZt5xg4YllmFa8mwfKzzlZfQW8LYlRYgUfipO3kjWNrT2UHmxi
YwOFRoMMCU4mh3HouOGfzfXMja3uQ4REON89H2j5BKcj/7kuWT8em3bDn+QtNLrD
Xru5QUIJlrx1HBz5245w8ws5igE00m0o4rxvHiOm9GMwlz5VKKp5DA2x9h7gWOZT
YKDzHCHHuhOLAr9WhrTLzTPzRgd3db/VTtp3J6GVN58x4sp1xs05H5mJBgbjPHzE
83tY0GgU+tUhzJwkbIYQs1OSKowgD/52GbPktbkjVxa9L7hPRUMtQqOpgWgvoqaY
O4aQ4HsY4NKJl242vG+RVlkTbefkR978rMPCi97aWUtvI3PNLDj736ts10q0lwHB
fJBzL20uR/t2T9GsOIWRhCffK5fuVO/+CBEXmc4wtdf7slpsF7ZV+A5cq7uCHxmm
Ybg5non2CW07He5WyqKn267ZkXKYYrjvsazN8AkDRtl0LGx9bOWX2yvt6cjoudtF
VWut5A/ZsMhEG0vJqUzfuybJZpHvFXSCUe6gWe7cGf/HemZAKbnKFX3fHx2tnMmu
eMj+0haXj8onyya8KmOf2wy+pNWhE2jTS2khkrfU/smAeK13jbZbGTJhy4BO4XI/
qkz8TyNCjE4WunsUxKHPc0w/BN/i7AR/wHwW2UcRzX+sjrrm7tqpeFRc7Xm78Owk
44olL+mHv2WUk6lmDKJqsET+ge52kQLgapzRnXAc+e+puKjqoS1yNBbP4et2ppGb
aZwHWGQXaj43s/CksZnyWaK1DGV+lRc4Jd5BJXR1nePmj4I19R+bxODAYo3aw736
RtpzRKnHaaxMXZyyNdl3P4quygVc+w0OUbdhh6deysbsT5pD3urvbSAO/acn2mRq
Ed3Xtpyc0Pm9I0xlQgbWsQ+7Vr/qiuyCee16mqvdjII4fFWUbB3rk+l0bVdu5Yfb
Vsreggb6uVntGfhT4QS+DlkSfkbkT0WvtSiqGIxzEdc466iPddJ0/nfn9ieKGeri
fwRZl5YOoQlhwylLQ0+OE/jF7CMfCfrF+1EUlX1s4xvQCDkC7ssILZR0AjQUCjaS
vjilIQUyifkGqM0emHMRnaDoer977LlBRa2RY4OhgvW7r69AM5wzJECTU5Ub28sS
zFWSN124HB+ww/8ZYS2F2QANHT80Xz7rrO7GFFAAbygtpPbyJpHutQFBgfj9BSow
hFytcck5H5WCtMb0oZ77O9NfRzr5/Rx2aPq288k1Fh96nMk4Aw8Lj1Jz8Zldjne5
fT3EzuhZCQgDBnLXE6FyhRkYAzRVZYM1MtgQKd8Cn08xuXEVBzSECKWKDZeNLvwl
ib6LiNFKmEKwi85gyy1rJqDYhA3evhUSg4D8ylIcJZ+wtH4rd87eASGMlIb7bT4x
8nnj28HOCVOE//fpaYx44Xd7imbUsK+Qlh8wC8nP/azrkCx9ouGdLGTRVg2Xcr4k
9TAbR8RWVrEN5ZOa4YZPx2IATg8hupt84wUMTv8Vin7Y/Sysle+XOKjARSDaTmn3
nf9iFuwkhb4NAGzvoP6mUy1A3ROLo13+82AAF/jeIXjA89t8Ivn3Nv18ZUd0G1wI
zSMnIeQmEobdeVofxjk1np6sx2kMG6OZu+2kGEzZOphyPzOf+ucbr92spqeiqmh0
q9u04+jFM21JQhoDwt5Nat/w0xz2AhtoM1AKVvUdZN1X8QhETa37JDTyRTLz3r63
f2oQfMjqyzY5/lylSk2rrSr5W2votu4gNRIl1CtTjQj2ykM9PrRn6nwvh2Ap0OGS
BWKIP1AZUnKzz77VaVq6f1UJ+emG5JsHYmHfwi8FGYSTEfZNJ8pugNlgrye7YY/q
MwoFWl3wF21DAiIET4/fC93ZcLSf3hQwkRDRQ3EBdIXQ6gaRqgHozMvbOKWcCG5l
E1inthbieXEHdqu2fQNRZyg8pebgolSgHS1/lUBUWf/oFBhirnpFk3iwMFVEQJof
Ly/pIXC2/FMe9fW97QTA8RLiYRGV3pg3NZHGCM/6ImLVMYwlIqf2UQLIrSfVzA0Z
S/G1RBajcNTmCkDcaYPCubuLErbOqe9Gw+qpAPhPGBw1PRjHq4rMnvAew/rZFaSi
wXTqS1lbQQwyNXZ1npWOVjuekzsKEHAnQB7h0xmdb0Ok1VKJP2V9CbSVFfeixKxe
iBwFNnpAzVIm77Y12/cLAKt5FF84Uz7tIOZSw6FhvFh2YnM9iperj70EhoVlPw39
8QyjzlaY28DLE0HErDbZMXqMUzS2BVHz9cDMqk3kOr3bNXxAOWysFoKSjNYcF1Ut
9ovJXmXwS+oBzn14me9ofqibgPPFvWz6qQ1zrBm2PwX9WJHhgYBl8LLAb1Z2/Iwq
hszb9Un42JVUsVKEydNZFY0s7vYcQku5xNqFMdryEJnsaFmMgfLiQ2wOrPE0w2xF
ytosqXIKSeIn0jdN/D+YtFyJtpZet5b4XZ51aD8wpq75j2AB0T2x8A3nH94E9EgS
gRpwUTpRXuVJNFa89Xs/UEdeTvwBuhekDeCo6coxcXvrtLkfxbrWVFfnJGsRKnSZ
kh+K5YqrdfXRhrjVewPNO69ZBHOiSWFk2J5ZjzmAvJhDhj0Dp3URDnm269OBJbRm
DjoTr8omBEI9r9DisbAiyY/7YpyZ7lMvjkoSdhL22Zf3IOZdc4ZKMOOOzJo5IwwZ
J7xUOGW+GNGVgxanTB3lkd9hqiCBTw9BLXXKKvAu3vvtwJvatXnnbIuaqzv0+x9W
c/IU4il2UBVZQkNe9ym5lHExNxwjlQ1gTW6vn3e+MzibfQnJDQfwPCtJqKG+1gOR
iC3m4F0D7SBgL45T+MRD5eAt4RuMn4RXYqaaAcuiamjp5dW2WPb9LhnzQui5vics
1B+/lio1ldS8NobevZTqAt9izV0d5X7tUrjUR4cEm052o2p8LxIMafBeAyVD355o
GqedR7vGI8M7cSgB5iAbu9p60jQG0oYXHdIsVbDJE/CHiVqsXTSquye4Aujr33l8
JhiN2DNCY+++SFx1nKvlS16QDr4PgIsbLipXI+IKndJP4aYuKaQU8dTo4+bdpkpp
51toM5xCM0KyzSB+xNV/pDXFR/izvnGV1DxRbfGFvCRAeZtZKyO868iHVdMFUeBQ
8QN11HMaveC+nawmV2lt+iZ61gTC3larstNfpnuUYTKBFpnlQNU7ONMPMrunEOci
BXhc3ZmjlRn48epFkvdB9vRf5qvQyUW0tEW8Trl863RaMGW4HNU2rpbrB0EvJauV
6v9HLuTsaHWG62YQw0zjeXoxAk4znjjiwvsOuhJdUKoyLFbKBWb8mZPy5ByFp180
ebfjZFMA7JM2tBUzzBsbvs8X/FWaFAq2NWPfQrWE4uTWMmsKxTTEzjoLueVLx9ei
e/FBZHJe03O9lG4Jhe3LryUttI6yt8CLJVHkn/6/fX6kVaOXp7Rb/9Q/fTisXhyL
wn/kpN3aJlyQg36tbdAS+EegHXBbgBb+bDCwG49RfPyQlgMiUCM/WlY/uQFAhJJO
zV0FgB2WdSLlq03pu4rS5LckXMhFn3HC6Jjz5EuI/Ry82K4KXPhUnVJRptT9qudt
fodGZhBTOlAb8GkSX874z96YXTkw4D34FLbM+xaz8IjCZOOrEs7vG3nFuLumgqMh
f8bPnIQcvar476wpC3ojEt2m5yk/+2EFNkeML7Q+7R3Uk4BZdICA0yaA3o9Rmc8r
6t+Mrsl4AQ8Pc/NFVC8JZXI40SyT2E4R7yhtG1fc9bCGecaF3rCfteXfqXZ7MfJ+
8BI3SxraNiUdZ7rNN+qpTCRjyQ7Dt78mwRM80oKmUyaHNaZ0vuGj7HtGnCeCGGO5
m1rc2XRJEUiqV5DVX/ZboIPG4TUN/5BZCJAgDzpt29MQ/4mtz/+2/FBZrWOI7emA
BDVoiDesBOCmYBpCk1g3ZaD5wr9KTWPLLM4tIUsNeT9+U4R6oljIs2VOP6ASqAUT
3nC8n4y3U231hZ+DvDiosOimalC+JK5QAXMVja+YiviI51C+aAVlGC2AqlM4siBF
UZK3XXdTdVogN6mKPj1x8w9vKJrZGzSxi0AyfRuSdpwcQeqPcjuVGVGvqLCy4iro
qRGU9n4cFWclm8NAfR34h6+JrQ8yoshDtZX4DmqlIDsEG4ywwSBJKpij596MdKx1
OWkgHxBpmN6lKfaY53AqXBFENwknROYfJcvEOP+9ZGKjnHO/GULmidMrVtzxPnQ7
ZmGvVUEQ44UJcorK84o82CllR0lZnHOS6npQs/itxrij/bsfDLcI+amq2QUDAqHT
j4/d5x76yofJBkld2iPMudEfqUb3w6SIvFqsv7bfzvOkLCFTVuUCN4106nDnSfMW
TZ/MRRkNZiTqPRp/6B87dQyukyUxnnC1GtuOiSJbojG398wAN7IegckBwG2CEpL5
Qc/PES/0/mZ2iZILYJpKnsBc6JgYzGF9XZ9XzKmkrJCzOy1e85ztr0EEzvQcq6Iu
DV4P6BMf/5mE9iokbCu89Nec5lQD3x3p73WKrkWy0AWN0yDwrS6bhZNUqZPuR+gC
UOtU2CFc+nld+p9EugkVDoHersV11Exp2XJrxozh8/Ezh81v7fn0o1wK/Bq0Ooq4
hyl6bIOhKO5SSCiQenRTQx1nCWteUUI/85RvA4whe74n/nGUQw1GVx6SLqkAHbx3
1K0t/EP9rLg5b+xLdqOUir8JOwZTjm+t/MDGdLTAJLFAOECb+9ibyiz/p7EUbUxn
lC69bAVwm2ZpUeF/F3ybq+FnF3S2EiyceXAOMbc+Wb2X46HHa/eAmesvG0DyRudU
SWFPdwSynCpqarYCxlhylXYTYfEJL713EOjmMCbO91Hp38jKto8nqLlrK1nXHAGf
rGJYv2L8cJmzE07F/I9AolZixg2erfU3pR1xgyZh/Dc8uQXu1By5lkSMxSAKRkCJ
2uN8d4+UiLLql+lAiCBJeEov83OlxzD3ZaEYx1DZH27v3T5CJVcraacg/GHr252m
iPLepxtKMY3cRFR5fuE2H5W2MC/PfxZ1gRqvP9XrBTNRcFdbbppJOmiqCatnY3Yi
7InXUHfDPTfCMRsYkiy77+uViJkWOl1TAuaRkyJ0ysn7QHpIe/uiwvfKzWDHrowb
xoQ5v96xrOn0Jwf69vliNAmSj/DO1gQn2EMgEPMv503zY+Uz4ExQx1yfVY6JQRTB
5driVCU2FWSun/34y9o9tSKdWgndjXGR5Txux2K2osFoKtMn1cnj8EzvaC7pts1V
cvaGihesS1r+QRrQv0Scy5Y7iKg0Rag7ESsWeJJqFCVzciY9Cw3TooUjYMMFkZHi
FqFkSSkBXsV/Rfx8uzxfQML2I+FFsWlOttjMetRK8Ern4s4QUivaif3CJdAKOYYf
y7u+HTxbGmf8ESzSL+bXnJHeWjW2Cnq8SxC9eiQIOOokEsm/hh4E396RmgGwQCJz
lu3Eas6ozc3lmz4bMOfOIwySJh/tpg1BvjiTgGw2z/B8q3kMadpG33b5i4tmmnzu
TM6tfYused8lj8hFfhR85oQV75gYJB0X1g4Gh336sCIJ/aGpu7e8l0LrBl8izj3O
XwuAbnLglSfVLHu1qRBKqhI61wpq/anA+k388hQrrx78eHYO3SSfU0ar0gf8dqAC
MU6btW2nO69dTlRpklRauEfC0/IFYAQsZvJmCQjveX0iM/S+F2jS/YXHv4/j09kH
74QwzJ89yt2K16+beJZDLz1jIBVvU9fxGWRqLVHSPJpmaXpe0xrkmdOCNSL8w/z9
gwmYQB3TyfRYzKKt0n0ICjN7TW9nMGRH2vdOPJK21s8/ULVzqFxknCR0A5hpaR54
qvU6WBtsyE3+fI0uvWegT4gPJwXJzRXofxE8xoV/vg6znKC2l0VLb9DF0o3eIJ7Y
NebdVzADHMT3eyvLV549TjZRUIJ+oKJsDkUTNGBgvMfa7VmWsFZXyimLMtOk61UZ
xuWl0bAZZlgvR9fTpvx0EyC3Zf0ox1OnZBo3ZR6VX8eii0mcigfWBCJMFkI8J4lb
B1PVqAvEGrXUOwDfnztRKmLyhmYZkOQnU2EOEEsLKk/CitosvsxJOBqs+MPyJ+UW
wMciyC6jrNXxVa8UOhEWP5nzkWKBPh2tohGcRNBWpzGtFLlwjx+vJHRz3N013mI+
8n3l8ccdyet7whOYyayRVGF+lRFxj2kukn0UP+TSi9sg59dQf5FS28S2gb90alUw
bI9uuA5mlXPTZtNplLKdi3HI15IT9gblJfRN2lOlb2B9JQt++OoxhrIPk3S4DBXz
Ij/uIXp6CU/8iAOD+ojzJKOlALfHbpxo4owMxSoPn9U1xzsmAxOVNO+wyoTr9NOv
r07nqar8OjQeMhTTPMCp0gCIqJnzPJKxb6FdILscSuV8hFGFZyWJvJ7noZh6BZar
73iPk5NgPko0R/4zTvmof7qYHho+XHoQBFqZ7alMqCUr42whXDkOgRKpW8Wh28lr
rDIrIor04jwyb8/2slFjbxxwhjx005Se7piIAyeAccFFZq/8ZJ520s6aDgddKdNi
vXaKBnaFO0/LU8tfXU+5JGAHXC963bIcBqYwlQCOJCe+ZpcRRzB3pzqTbDAIhUC+
Sfc6HqxcSZbk/jAXMUrHRog0O8W4rMdKoEpYwtWtNrZcVQqb52CPD36FdiiRYkfv
bPqoW8wfHQH1KqxQvNFQvpLVJyMUPAb6JHvD2myrjbZ1TtsqucaZlRDMbOZvWOlk
kWO6FK5TVt9eiG6NSKeu2tI2l49yjk9Q8+DzJHdQoYN4mCPIkyIKHZWTMJPWQNxF
d4/nLqwHrt6L07NeabqlIfgH/XHS6s1VUh86NxyQfw94GmBjPNvoLC4V80XEAKWC
18KgUZ3qCPpJ7JY0Fwrf6SWUugYocn0xhweF0/cbQHan/MDK4crjUP9inWH2hNnr
DqW4G3iwRL5Vr7xffQ8y8D5ndg75o+x6hu6D/hlkCWFJTltvJZpPMBVBcy3hCaRk
UxadN3QY2PprxAJZuuKGaDqVjW1QRgWaoCFc/GrerFsOR5VlRhR/Y/7qBXyH4KSf
tjzG4qRd4bZLE91/RXeIWCbdmcIHW17JY/dwVTISwPtirJ25OVCnc3JRs3ELzzbi
yZCiQ1vS4tW1JhT2O4HtWWtfDmO53qd7G8TwBKCug8D0aUpklCW/LiyA3BF2BjeS
B1Kob9CNIfvvsQCkBnoQkUihOPAL6rK4RRG271y2EQMb8dU8fPHSRAxlgd6Qiivj
3kXRQ1mPoPk99foh1UZLSrFnUZWQ6Pw1P2gsZIW5UG53nCxoZin0XqYOtcj8Nh+i
3PDAnZspJsEtjJh3HSJgW68wfXrDyQH9fi7sHsQoM8GlXKe1ErVqK9P6wssVu96H
eomsYDEuXtZ9uLf3hak3Y/b9uNoEDGhbgkPao77sq+s0UanPWKMrg2WhvGrvRM2R
PgklG8BDcS2j/Ow/37BK46loBmWY0jrTQMaFmdRzQUG/w66+5xgJ+g3ctzx5wVKF
20x0UVFs6GmpLYYUnm0xdwwfGfceec2N+W/rnVP4nBEan5lKIOmFPyZH6HSa01Dx
QW2V+imxDST+Vuvz+gwwTabLSfxSffZ7Cqbx/dxZvLbiQ+91Vi9Poy91uumCdB49
0Zdt76P1EH8INW9eC18NJD4V3rEJyPqWyVdrL5dGP0llBNLpx6JdftMS2Jtci7ZO
7JzkFJdKMuyx/oG+fPNTLCruGgxfjkmycCrIY4KMDUFi/tiABPUShOfmKtCPlvK1
GJJ9qVokOSQwr+QoCA0La4HlQpfv4hVVi4kyynP9D+rFsLsZeR36sJBczc5BnI5E
73Q13ipRGgEd0jyYpFoCh01QZLuap5P/K1DRcpkdyuMlEq/pO/moSZd3gXoDEtS5
WH8Eqv0OIBlR4ejrau5T0tQEs0/Z0G9R4QwOw8yCyk+GzA1zAL7lKr732L0z4M26
UkHOT4PaAymjNi89kTqUlRrzXjwkDYFATwRreJlFwPxeNGX4ZM/QvBE+z73bMsrs
gmd4obLXN5fmHdFDWy6twrQBQN61w8Al5iKxPueqS7WlGoxncqFoHysC2h/gVRle
IS+I7mjl3IAOrQAAjYNhbz33YJ37p6zZLnmACuVc8C4Fc14L7jzhWVA/x/7a48H2
BuY5GTgh+GOLsZ1kfbBQH1D2ivQKce3Qv+qRzp4LkMVenNz7eon+0wPaZ3IfE5f2
wuRdxKu/ogJ1DcDvp2niEpTJyolqLaFtyaut8ziSyC3/3EUYD5LSuo3dJ0WsrMWf
8jHGMIHBRy5B21kCoLMRQy+B7CE0jco+HLZ5WKYQVsMOjli5Z2bLViemN5RMzqWc
el+RrkzPYwvPuFyEPf5knOwyybF0mSIX016BKF0lJTU2cs5GdUqDUGXYcW+lw1H/
as3EwyPjX7AtJ3BFmI/BwqGTiU++RwrdsIXBgxY+de9YlVHeXZ2wPX4ge7rWRGCx
We2KcprkZHg7QNpM3svC8Vo8GifTTdT6NIpX58VH7pEFqsYt2yjp0kzz7rTRLyqs
PwknoGFER0ETuSSkj75BRurcIx348Yxbu80ZWFPSI73AHQl07tlHJW54ancArren
S7N0W+neU+Y2T0URAP2SZW8QI1YUxKGkmh/5oJVBuKla/hHrQ8S1wS98iHAZ0V+Y
vzLOLWCQQ0g+O2ZbbVIACU/h1Xz2a9cScn41Qk5E57BWB/xXbXR6DulzYJVt2UAY
vVXUn5noyTIgAr26gWxtRhuzRETorCoeBaOO6F1ryiHxTjEFEy5k9Nw5Ad0pBCnH
Qd18A9UPAVxX9DxIEtCX4xojDq95wtAo4eTr0BxftDPpRrVFPZzTp9Iux46TloRV
DPwr5ANp6HJY0GpwsyfwFBUOXWQQ8xscdZ0LRDvBO1ZSbrLqZsbfBqam7tp/d4db
SYpeHNY9mZMUltoZAeX0k5Y1kUkmB0ZRLYmy9KA88b9LbX1g3YSW1uugPb273Kro
Y497Y6IZia43J94uM2JfkhC/L69UHLLtUdq7xeltxZAZxBIYaryDGvuUeSTtau+t
wq2xRE49sM7fXKYYv8Ywm8Cp6oUN+IQq/KrQGq272qSB/8h4F7ayG87JNS+gddst
I/WOsydOeffjzDj4F68J+KHwYzDAaYxshM1tYTRW6IUhF6fR4j+B3sEd8PveRbzZ
UfLUr2UxBJSwZPCINL2f6c+wdseO4IEFsDB8U00A/6TdMVae2+oT7YvO+Sr3maYH
5L+0WQXzCHQMRt8MFfPKCFRaQkqCZ5ytk++hXFNf5moiu52pmIs6zN/+6HZV6v9I
M7tqhmPn7JEfQBEU0kufqJApKcAw5ASlGTsfCLt1XOEg4QL9A6f4+gdd+LeE5FtV
Qg4/YDQo5p1ROoqjLYohoD7F7C+NDYeNHDoBxcS72XI4kkJvoyjIEyZOR32hupYY
ZCkwKb7tmRhYo3AyQUpcW4cjNm0ZghJAOs5arXs8R/RYTUg1i2gKRYfTx7LPAo3O
jJShyoONrPnnZ+hdtClLS6Uz3X1MmkxfCnoGNOE/wBqcTYWhnMlc2KjpCfVW3nPL
4TY6IJjNBuLqHpx5vHzrMUNaSS+v3RzRKBcVK8F6VZqee3Vs+/UlmmGxB6Tr8hf6
6qGvAjawbfDmzkO2bSVuZM+WKhkfLUugqPsSdGw+SkCQO6DUWEUcydM4jtm+oEyy
bh0u74lU5y0Yw9j8abdCneIOhWhBxsXNqSObEHkx1kAS/KTiDaC2zm6NMSfCQvqB
MgCgSHuQH1ajSpv4+wfIjpG4QbiReUS57RDZV4X10v+ASY5DGvNfmhAPS3e6fI9Z
UkzWB7mgmM3bbewhegYeCpx5lzQtsbU5e/BCriqT639xZktAfHTyPkusGUI7NUmr
icA4uicO0JyHnh+WQlqDxIeK0oLkIynBBFIsOyKTVqsXvlvNEcYwBh7TdQLE41cj
xhlHElecpk2lPcCUdSYIADE4OPWQo5LaByCdBEDX+Bph/KdUvYKPPZs4zp6STt9S
mHoQTFa59JVGLb9dgsEpKrik/wGmXfejXRkpksRFOi4WwCFnDQoLX1eGd3rZigbT
3d4TLX1LQExJLbMNYcRTI3jkheOeYJh77sd0wWM9Oo/TJ6lyhGE9qJ1fULY3KJdh
IMleiToS0xK6Xl6asun/qekY7q+xa7HDCZewJ+digVuEVoLHVNAKt/iWn7mh3/J7
Q3vLzxjKtX8ZK/mvHungv++l81pzKyL34Xa3cvBU1ab60sDNv4AuFGti2aOmuNkS
YcRtQF3/n9/c66KJki8daHhlSVe4AYTD6n2H8K7mHp9lvnvF29gNanRj9I7SmUmr
Yq3A9mG2PYJLkQpdg6TlaWKn+WIFAuCJfyZt8G+QSkPAEeQSblHaxPQIkUaoHXIJ
DbpwOTpXVYF0q36S1EdE2RX0eCjYfg//ez6If84rVmVblbtkV2oOyAIfcJL3l1wH
ZaQHBCy4y0FwoI5XKA48pcyPVwj6/FZgtkSKHupXx2Ge6XLdHuyELAdk3P6S1HTo
Rp1rmY/Udc5ppHeEGKIHHrX/1nwkUyFPgn02SryfO6EwIIZC2Z3xCRaqANSQckDB
Wg33D2WNUAgKeovfpdSObZZSS455ZEb8SKCkoNfwg1r4c+OXuL930MwKrnWk4G8a
fgQPkFXhSfegEVsyuV6wEZKfTg96CzNpszRqY8xuN8hsXLaTsL8ZWvNqPIho7W8K
6LPmM3Ofn17XpVqC4tKRZvyadCKYYdMxJ7AUZNnahOE4BkdCZhBuxBYmVJ6T9oMh
sAvtsWKNw0X8gtDJBcyM4M6bdfjoeRC0onPgWVQM7XkYPLpGJC+1tGijKuVFpqeT
+Mc8H2zzt6/OOFmPZQ5StyxvBFTz2FFuVAYKMk8DbJl8ocIGFLqtVT4dTBRqzISb
jM5HjF3Zvxro6p/GjdyeX24SUTYF6/G0NQmVJZazl90s7ROiiXB8UrARiwGNJfYZ
oO8ZmdgXhYn9yULLAsJmEjMIYjVlRUP1vlWJ120GRK0gCKmrySbjnPuVWhv/8+np
TomTEYB53crflMXxypmbUUgqBqNcTFUNch53P++a+jFk96q6mg0qqYZvhRsQBNHp
aIM+zvcqXi4tAknp1xR/9UqOwrkb4IADRl6yCv+bAQClwNHSQayjYYZz1OFbH0Tq
NG7N+F2ELzDHcVK3c/oFccHOJ6SDjfJIxLpEz5baRlr8THIeI7j6GXs7YwzNnacz
4CbPIv1kPW/i9qG9wkn2QVyeMFpgUX7mfZMnasufX9xnftVydQY60tWIXhxtLU5L
XVVtWyUgtbOHigru1Xs+ihPFA2vWuOq5aYxHCg64tkTl0KJ4H/sKL9c8HzJlla06
b7P0YuRSVbgPIIcXe/uwd21SYQ0gwjpSkkZk/Poi3yZ3wrKNqVRtUchVoEGAEhXH
YfMX3JfbelCVJ/CpD0hNAdFQbDJwf+hJHmjEMPI43I7XilK6n0RMCp++I1J2FaoQ
s0ttZj62QO5Icqnrudh+Z+lz8ZDb027b25eP3hjZHNC4If1mfADE0EBCieuqx2C5
9DShMIlHKW5Mu9bx3a5+r/eluWDStF/ll73eyXxcXoqPDremAWN3kO80cw9B+5Ry
d10RIgxG5M2rNCURv97lWqefC+iKClkVFU2Ij+H/q6H7GORc4gMIFUpkgD6f2HuQ
GRJqncQKsC4CLrnLcQH1n7qxFhFJRC6wQoGBxnnaMAtprpJ3TmBigczVg8GeUNLm
9spY1V3UQOkGFn3BRBH+q6PBdk78iNjhLRWrdJCGckONClrILM4Z6DcOXc/+Ej1e
uqXrbHO75mU8bb48mcUYxdaduh0E/89NyBXnL1Qm1A1VXIQejowHvT0TAOeLDqdr
SKJfX6wFJ0F8V2NMEh/0RbnmFXUHDTtHlQSchzwctTknZIUvWieIzXXpsjV/kOoU
BxwtBa1fQTKcfGRnUKlweMKuR4WZMvtnyAcQibiewrcQyGoUXvtI7NVf0pYMLD8e
tnX3zMdU3OsKFrs/hyR4ECRKR9QjiwfbV44bhJalwzOvezINzkhfAx6afc4VAMPc
O3Mi6ffAgPEzmk94nwA7iuVvuKDqHNo+vfo6CJKHEtTRb3Uem84oHdW2/MFesKFs
ve8q+nNjQW3pmu6WDYlOUfRpUKl9bToDfu7aVeJVOGrT5xRnrPSfty4qKwaticFg
fwGdVlsLRWRXWbzMEA+n+0igcLPoWKWfDDRzssHhfWSEy+2QFy+hQA4vXD+pT3Kw
yr0fnfvqio+LZf/jl+k5taT08i2VByLvJJFAI5AAIWEVXVZ4VGo+dURW1hMpMOoh
VIyxTCdaw5c++VkP38kWey72qeyU4kln541R2PWyZdKwE2BXfGXA9TI2qNRV5kLE
7BtHC2maulGV2I3Z2UDp6P++EbWgpVM30W+tOBZgKiKbOfpr+dQqP+a5wQuOKJn4
zP282EZ1iYgd/W621YL4rEMqXXO6bj8RC8DxoYk6YOuYGDdD+FJSGZgsc3sizd0O
6VWb5mHC5xMGBcxmnwoIvq3nTusPlGm2MNymhnXrx7/SdkDZqJlVLKv0bYC43zS0
3tmFoQwxZ0UYboM8qgmftYetOME6HcPOWXaL1sGaG1LUHoTeeEkePxe3rdEtkxOI
akc2+49V2759haq+8NoUC2v8k/rlTleg6VjRX8EaYGrKHV+S0ZZGGGwdcmoQqVA9
CuAPJ2rawN2ji+8uqic8sIWnq+JDElGipRQB7EiGWpG/xM9VFQwJGKtMnm3QNvlI
gsIac5OyUq/N9wiynSWBMrnQKTDkijIfQh+YCzLjmrM9DgZaXn3afrKYlhwnVhV+
PFrch5PvUgY9kcYpK9KDS5eUim6cwlQI5ahU9rxv4oyefAQt3v0+sGDxZFxu6Nmn
FJu2RrYGiopxMsX+qvzOVCtD+gUoIVhpIBlcbkRrEtiHjylFFNCBMCNkpKmYrFvx
CGrPySPEWlGJn7tM3R5FDByBYjvSWKOGu/EZE5V9GwWfet4c//kFkl9m5mCVFM3l
l0lqJ5vqQN50Cm8KO3ATsnXMLqyDDZpCIQKrVEdVO6HDzFT0Btp2XGf+IIkcNMOX
UNMJLMaao0UtEWY6Txx/j/oVioiFffy4I8EtcHNhjWrgN0dl9jTUIoNp+MMjYOv2
C1Vd1ZDZyGsXu8FmxwraXwuEBK14mPR+rENc5Ix1nj4Y4ER5C8WDgLdvcmNC1W0n
cqdLB4w+JZ/x3z3VvVuvueladoybX4l6azWaGN97+5hblkuqN/Pym8rr0DnqIJ7d
esw3+r8oIWaXt9n1R/jIdAmzjGGQeTTdeKEseqZkMWZRxVZ9pommS2NurNIRAF37
y3QRFKQtF7wNB119xMD99zGvl14kFkHuqF7QvU2FgQb5LbnG3ZRTTNivjK3JCy01
rMwgRqeD8zwnsM9skDzbgs3xtcp7IBBLD643T8+NRkWri86abyC91wt1v9Lg+ehV
wxu4HEqVYeYKfBoHUaV6sb6QReA4qVMr7cq6zDpsKK4YWbMObkKRCNF8yWaxYR6w
fCvUfbTJ/+rFXyG6cgIh2SLOKA0zBYNUQbmyuy7zbTaxEoouLtOSZyeDznJzvNL4
JaXS+dagOSV3O8RbjUYkrFt9e2hMid7J/62+4KAmxhDeW9a6lmB+qFbilh58AerR
ARoS7vDKlZE8cau2n80LdnFNKiu0UimguWg4Rg/qwvZDnILfY+KmXN8y/0hZXN9f
L3rZQTdt5n7QCAUTaihzhQ02p0jHKnYTZQoUytWkrkLg6NRC0qQO/znFqYlZQzSd
5pO36TtFdxio8Lb3lePw9ATUIk2/B3ZCuU79WDBFegDSJgwu10Ig/wgaRViY25e0
062DW3zmnqMv+mpw61xJL/qrRl2FL6ITM0XRxDqsKHs+k7uybzV775g5xaXji9vS
qUZn0DKsr13zEaNq3vDQuXHHJkOiz4+jTV5cjvyyOqgNZfZLYsFxjZQsB8oyhG6+
pKOzKbY/ymqilwiB0Y+QPIV1Kx4Vua651GBIMoqvcYhB0mO04417QMmD3gG5HIpZ
oegTDf+ufAKXOk+BO47QVY3aU7r57D+gyp0l9NV3USOV5QpIWOhHZRvWmmtC/wZ3
Lw/eI8muX2eUHigohn0kvL+auRQpvOWtWeXwl83ZssrZmHFmrvz32Plh1AuHiLmy
SSRP66iYQAz3/UXrPFC9OQ6FJso5gaOmL8KTNfbxhW0JOTpc0kE1j4D0aduptaxu
yXR9DEeEpb+/Z5wSa8/2VpU7REDk/nzS7v0OVH1ZtUGdU3/K6bmrf0CFXPe8TJ+g
E2vNr0hqN5xnjATE2cKraIhHYxLH+d8ehkeYeESf1mjJQ8jzDK8iBhD/ZPWYPDq5
8VpHb6lBY6M8VEYY/gU71e3w+b2NZspTVPQN8kw/1fA/8KoDSkNaYoVW/ELWF6kC
3Z0QsZ3b9XLawfHMYUHT8Vu6wvPeOWX97/WfBW4n++0H9lVsva9F0+lBn1iliqyi
bCFrttsuEOvhv8GM9gP7sUDuF4YQyrpISOVQftJsqYG7CpR/5d1fiWMtbvEKThM1
Ge8viWKuzfDZ+ma0fMGS7m8aJj0gFUC/Tw+00Gjk+o1yV8/Fwhjg3VHfFicqIwCF
ARapSydkbczyTSKS+hJ+a3onHWlwzw7UwVo5K2STS0DpkkPTc1Tlmmfl2ls/v1HW
6mBYYaH722rtjMY4qrrn33qpgiH2z4DScwGdtkOk1R5xT3iw3b4VAgVpFVxYFw0x
FXOeoWNbJcNVmOm93u70TUuzZPZVj1vD7MQp5i4hiE/49qfsxe8YnsmGRIHNMMGp
FInFnea7/eapz6Gc7Hhq3bm0hhg/fTa+A0aMnTywADAxqCG/x7yJqPQf1FnadHvJ
BiE2QShmwP0BbNR6PyTp/BToeYzFCaC/weWcpOeu3OuJFFVDL8EHiMDEePSWM8Ln
3i9h4JtYTUxyb1Szx3kSGfTJ5euw4E1Yr91DODx8xVxxi53Yr0TAVhJ0mlW3eE8A
Akgi7knK3rQy5KQ0QrzrQ1QV6V2mn5kKnl5sQMMaUh8yQTVid2WjReqoXq0dHhN/
B7OeBpOAWLugA6Q/G8SpirfElOzIzeSh5DaAM6RCIheg5rlnIOww5ApbLp0rxBKO
ukP9YMeR7Y7T/3Jk3Qy3bL9YZT/pOv7tX4cpQLIFhIxuWQeGTOb986ec7aa7QMpW
+El/huilE07doQdbWpkXV+c2vxDUPO8alrXke+VTnCoP0jX0rYOWtCNomnAYUBBu
OrxOjoq1QeugDcfrWuQA5EWAp9xFGOaJ1DTWvgLSJdL2Al9FIF5GI9MdEkVbL+H7
q8H3eo9jS2LihcZTLmGwdCtFcyalNSXU3LOuCUbup9VOErnqdorvVbthCoBqCm9E
WJhsdloLiYzMbbTn5388OxkoiKmGsaqKozzwxuovYJ00qdqCSs1HUWsRmv89Cx8B
6Z40Hs1K+siWVwDhrRSdwZQLV6QE2bgRrjI+Qvdeh3Dlm2B8TltkSpRSFQ11OjvW
b9cdV/gswSCWLG1Ya52/kuvA19lmnj905YWWhzpMCuhnqKyhv/zBUEmEcZQGwF6i
VpfitIeKkI6e7WL3+VQ8LsbQ9W1GXTLDDrO7RebWKErVI29paiSE6cMhRbN/qBcx
jzWkucsYvYA2tX1ZWBNpy3XMYvxbtw63L3lTWPgFMNKU3OXRoCUuBJzxMlzDw0L9
HsFs1sol/pC0mYWl/xyooAMja0Tyr6vaJU2AKuOIUnu9lVF/nB9AJXntgdZQ92el
J39nu08nkIAmTS81vKxefUKUheCmcek6/6FRgzjgevhyLTnhmynbwaiLQYAtuCfX
ANd6GCGhz7sIbGcANfbJYh47QivFra3Bqb4VH8Y4wkegd/U8B8JVn3Es8Fs2njL0
OgXfHGjx1IEy41MEPE4wcaCOF9TquNU1vCWAoAaHxroMC7IDYPtEfrmMs0ErrDDE
ffecpQ8xIOGNKDSW8WqE1rURXSqRulAfv+PLpEusqkPKcFN3On9/o79NdPzBd10M
bvueG+TMFcF+awG3GCfPLuM7p3zD27qMBdxrA/eUvLlCOeucF6f6WJfVYLWLRV0m
SStLNaLCmD1ag63TKe/+eygZxe2RKRS4oRSXnFlbx8Du0gFpHIDlTQT5HOIlSZ+L
kKqh0Jf1ioYQgkG7ZbH53HN4e9Kg3oS/cFGp8G+XbVW/vuqjr40YvOaShTuptpiS
56DYrCGCyZjLno5nGlMThAcR2J0MSwhWnkNqSPRXgJYEypkx47sMFB9pLTfD49nA
rEUqOn5Mf+QGTFGsKivUBSH9tBjqZ+AsjkKBPBtqP989YV/e61Sa0coz48/jNNHw
BgZzu/793JV6Vxg6TQzQ0kTgkX6Q29wHiyEHYIAnZWiJcUco1jMyJvUOc6gwFcUr
I/xDigAC7dpB5EmW24fHwQUnsi8fz+qN6eEWrIo9iaZ4UD0xMfR3nU0pH9U3H/ue
Kc0GcA3HswCrNdbY9ef7LXpzlixSF39FOmraTpmXMqkEuwqVFJUR3ign2SiiDgGY
N3FvN7N1m0jeNJCrvJvYbYrTaEak/ixTbLl9GqSCKssltsMBoqDIMijTDNcwRkP8
YHQqSK4UzYHrs4iery5ixs9AvKOOC+v4xlhuW+p+23HsBD6bs9Z1GU2OKDZHwzBt
tj4J+qKKwgPQlmkPRUAWMKRQFyJD8eDnPM/bwmaNr8ZmpxbIS5httQXwoFDpPKd8
NOaTjuOgiV9p24Xn1Zgt80HaEt5ZqgmSkX+knzsvl6/vnmfuVrn5b3f0ENnn8IHi
8DBBKNR6ivtNu5v+HK/FlTYaUQ+OS3dQHt8m3xZJRF9DwHP2Jexr7HYvKBqN3WS6
vdo30Qvubkffd+lHH1TN9Bze3OmXBPYUCoQVwW9DBds985F54l2+M2T+Lv8CkJHS
/7dFtR5ZgDAAsKi9ucANekieKIxryeEReDtboc4iKQ2JDP4XaNfwUG0WqOaGCUMI
+P6GOkvsWad6lzlBDU0A2k6JwDJBX6mz5cuhH0RKEEcblEyoIsaA6VDDyNQp1hmx
SpPsPpAGqvCBtVuZBWQ71PU4rgJterIcQa40Gg+9UH2D4rP4fMZz+KgbblsSjbqP
ATw+2BXXAlgHh5zyjaMlOBZN6Wa6j0+d+sPbgmElPEpSHdSZj0Oe8pRP8cVM9/Bc
SiANTl0oRtq3TPYIewBk+nmyFoZBDb9/FZuF+CBpv19eQcjzdqt6S0tc9pEojiS6
sKYwiaAn/7HZzGxMmt9ZSWuxfLPChS8Zvn8mqKyeQaQScpw3yVmuCqZuI1G0AFNB
I+WVKA3CEX4n9CXW3oLL+UegHEcT5i9/NFzyfrG5EcAjCYi4sBRkKMjY4OTdZaJD
PpyqEEUm0+ziovFMtIFAo3RPrNkxWPOLvlp7Zhn6LDXf/bO9xRPDmPjcQ0L0ZrUY
ETxZRjiHfNYszFBgpiqUQPsZqeUt/dxokkjSXWUh6DvqUNfRwEU6MQ1RAgS7BhHR
32JHQ9bhua2UftM4W/keO4+1DT4FDnixkNR6vFqalvUXW3eErOVnpYrDRr0gq0dx
dCQr+uab2r2ZfTPqmpcSko8DWOr7w5SXL1/cv+l+yzy8A6JK0NghHY5AwZfCM8Ao
q3Rj5lz2Ec2xuREoYZQOdPAGf4BP8bpTeVwBlk6ILz2ANcPtffI1DbVa8v3P+yyc
PRjup0hHxTJfKXHoCm86b4WvNc29dCNPMhGBYxcOUdaQ48B/QGNHsJl3yjGOtAWt
g8FU0GXRB+tP+9Q3eSoQ6XpcaRRA+wiB9nLQfTuoLn8bBmyYeM6PPb6AHtIssx5Z
gDKDlwl4nySF7ISuQYHzGJeYCpDN14BCwY9GO0xGGoY6UWdXtwfF5HNGXx+GLg24
fZAn2yckEsvlAYuDcs4BlLJwQmw7wNnz8cLNWGL92kwGjzGzV1/TybBMxiQPtAcv
LhYUvP9zbGVmXofUPDNdvuozTdG+dXaBvIhL0B8rvpOwt93wjyCGbo27jDzVT0x+
0wOb5Wf4dLfc3iyQRq+jbeTRSI/Y86RgQbFWiWZtAioTyN+9waEU8b5jXwCoAobb
ZCucHF8/XkRowUw/5D3VqrkXmEqF8/R2lBt4H21AU0iV9hdfNDxsSMnWSYUtqSoy
slZ/DFEqL0NRoB5QPeCQC13b/EdWOj+bmzfNQfNeEWSOYlrbJwLWYtsmWzt+MCii
+Elzp2Jp3sUdV6gpVHQ+gWbxSIIPtzODDpTN/q8f4JFW79IDWREHnVWWqmhTpR3y
c8ScjSD9xvg84VBNE610P1FyOkfpJJ6R1M0Dl/XriixAN2MzptzZCarWvx2o5HWe
isN2BU95ObEmEEr0JfsXT6WAlSPYMzdrV3ibRj4MSjqyrXJKku7w853YFojebVw1
i9WtoeyxvKMopFpKWbhFb2QfG/ED3JMg7ivK7BkNI5exktu1oRMBi0ZmnVMGbJBn
lFGmXerQCMqVv4jE/PT6BNzrAgP7mF8Gx5tQb6Nng7AfuAhxaiTtf4+T2tYgucuR
Wr0PQh2nQXuN7uLxos3MaDeZIzI5IsEFT6Y5CXdOLlcriz1+bflCkBBdINuEF/iZ
PfUTh/vH0xPY/YN3Jn/6RxELlwINfLAPBmr7Ejr2X9cb3BgaRA0MsE/fb9QiRz6f
2jQJQ6DeoewuY/8Y8XL0GqTXx8JstE9IlhLspBi46DUvEn4eqlMXWWuDyGcukEmZ
fCJyXOT52vehUKD1Am0Csg3qugwhXokKQy6W/ifBOqkcJVJz1vau5gR9y8dmewRu
5vftAQgwSTvh0ALl8323wmVLlOFdajm2cjGPIA0apjao5oEhykK4H45B5pC8wcUM
Tjnqmc7hOkpHBDwTFEE7iGuO4aTamiBdED4mz93Q5g+dXVVbq6XlqpDx1E6kjLp3
XSF0ob9haDqSkvR77MRMxSgRCm1PloMfHPJXEwx8rtZrucMwb2dGnJxpRxaH+gfa
gQKpTbQ2kwgx0BZt7loX6AD8oAoaC98W9g6lHRuGzrNlMZDUU12Apa+lOGg8AXXx
L+XvT6OZqkzaBgMF7S99leFTEiSuvu+B1118zQcMyxVKL9aPVe2pv8rLNgi2q/GZ
hcON+1Woj96gI4X7cvQgYyTxatzu1QNXME9HUT1DwEF+sb9RdgMstiNeUUDH22PJ
l0ckgTsOtUbzF+lmPgdA8iKmE1IvsVqywetNqdd3V0efEPRUTHb30M9qUMfPIqjl
D6Vuwyg5g4JAO+w6SjSTadLurclFE3d6qCL0AkHRsRXba4BQuk9uCBOWVnH8Avkw
L3pU3KY9EH1eyRUCOITW3d+Iu3F/e1fYrbhaQW8VdE+ouw7m8mujwDpYD2JmIN3H
aEoX2Ug2CTC5rxG2quKgUIYGYV9yKpJS8JtB6ZJT3NV6eW42KRNvscs4mROzRHau
7tmErhB7RQBK6oTi8O6eFMo4Nd/crRQRePlnibnd/btreloDPKzIRKmockcBiVty
chfmsFxSr/G5AYJec2Dwt0GJMh8r2Boy3n6p7ekoiaEE3V9oWSG+W5Bcg0HRc0gW
I2ibUBOEvozEtXWBvFdnELUhxPwL1uMi7BCgXd0Sytwp02p8cm0/E+sLCyowV1Cs
q144Y3TRDXIgBURzSlz4dU0CW9gM26G8NhwtDz/GiK7lxF5pV/8ETP/1zH/t6b3/
HzStUgc2jEbmTHGo1enVzDLOGoJb41fekjcERuEYdRN+d8ju1FJy0zckXDcRucuc
OnDIJrbESQerfOew0yK+c5twPKz2Q8zHsop5sK7FarlKGmAf8s22ERziAdWGpodF
D6SKyMgXToDwDa+wUq6XroG1CG+flj5wS4S0iEnopYeXZJd+O/OMacB1Hm1fxVKU
AfU8zszmjJxnfAOOIogNrtUeZoU9HtF4jnaEXB4IYrGRG8cDWZB5NtlsiW0XOEXH
1C+tV2DhY2O3aOWNZjC5MHF/RibMjLtCvZ4Csxu3a5i/1cJVHx6QAyfk2J9xZ0j0
ds1lHjGaBxDP4sOn2md6BoOI22/s89hxxNhOnvsR/Zx6hQ/HubkW0Mlm75N+43SS
wjo71xITk9Rkq4A/saGbsYUwLEsP6lNqFeGkADVEl3V5oQEKqSf8820zbpz2PZZi
l78IRzKtrC8igGFJtN1ML+O9OSuu1Iw1bk2rDZFCybcUkg2czmDJaEw7m/EZibPz
XcSLxTkHlNG1dZcuNrRtobam+w34G+jmNaM89TLEQU697s0XsWochxufwRFD61u4
d6SR1sCeaPL4kIv5LGJgZQK4WgGJ0mzsxsg+jL1yzTORfhURK8yXlVhlAt1p03mQ
AQ56QHt+APxwdffTdDOYayHmiBU6BfFqVXwhasRGYfcB5Y82qGO4SBxStMrkKQUV
ziBHbhekNEZUOGvq0gc8XLoIPVfp0ZeN0nE0EzQuvnptitygYwGqRuvhGau1VqsT
N83MHfGM5btukFAOmd17H2QOKr5npXj2WTA1ZiKDhLddW3bRtFPJJUEc6XouPO6u
T2ByVT/xXNll7sYzVLewnIosDQeBu3VgAh/kCbd1zDYYdsiEsvGTAnWKj0sjoie+
pf6MDGl6k0IGXJFGDMYklk8+S1lCFyGTOiEMwB2Z9aqfTu5+1sREzZzKTiYkfW5q
is/PYhSDMkYYx0akys3UgC2LwPo2Kez/UlymtvHsz3ovvaVf2A69CJC947bMhob4
RisvfgWUIucB60XGc7D1xM4jO0jdhalbDXma+ppnbKE7T/TXzWOARsEvju2Bw7Mw
1rI5ESvzSFLCpdKRJoO9YvW/G1yfdb08Fpa46QAOnBeWNXOilSxwh0jiEstu8mr3
OwLMVZr0imKOW+Ms2SrroVJHPV7P64+jb9CfqRWL7Iepu3DTH+VZHfIwSMvMPl8y
hpGZBKvYgR2EiYBFHASdeNnGcRyheVyWdAifs4apWp4eSZbUrlXICGsN2NNGI2a3
s5hoXnsM5n/9nBYAiC2AYafKzGv1e9IxyKBPggDE3Gidk+D4jNnmfCyqOGLDPTzY
dkPqRSz/8Yv+fTEWEnZlKpbMndDOZaSWEg3sOCz/KlE/qxad4V/K4/njBch4UPHj
SyfJuXSqeBMyRvd5jmOnXLpJ/JFtmkxz8JBzTvuvIs1wUbGB9NOyq89S0TFQgHsg
wgcFD51I/XAE/Izc4T3QO9L6omGISoA0CEzkoVigQoyB4ndU8OzAFQxsJiM7mASt
kXVFYXu/djLf6X7njumkJFtPUYV78H4PfcQ+G+H6eZglO85PbzS05djqoCzPJV5M
iS80VDe25NQNCBIEkp47SZrKqffNtZs3uXCboQz4w6Jqs0WhScJryYgvb5KugVoK
jt/jhZbENGCkyJ+bpi9PSj5Z90oHYwZ7GHmfHmrLPkY3cnxOFSugsL8ddcDz2Hu1
ei9OP1Lzo5F231xhuP2vLvz5aBcfritretDtDxXAJJqkZ6xZ/QVc6/ah5tXsZwbb
u7Azs6VfYA3EywpjbFYZ0q9ZyR8suNVE7AjJMEqZ5ikMGZcNSe2yLwY1xTMssb6o
EeyumOLSuiiZj4XhgljsG0X5JvMRLL2I6+LwWSTHkTSNcY5u/IG16yxFAZDFhzXi
OTROiPWsPASweYtzi94T80TSrnPl7rS9hWfL0J89ZsraGrIgDPfQsXpRvmzU/QKy
wloLDLo5EReCs/4AkNSopMz1fVeRJkO/EHFBsUOVLVP/D3m1JADjAOshYlhmHT3h
JGYNO2jGeOEIDE6MZiJ6GD35HAgWC5b+fAYdVKL/bpqMhYMzbgAfRT4gjC8Cgu5j
izlqT97hO9sXwjCBHAp3L0Uh02jd45aEypo4FzNh6+8zvK9kd160oY1C8Htx6+hP
VWhlHx5lIuwmIY3Zs2R4raYhZJ7oLx36HEL3YC3UIyk/m2qMM2WvCr5Hfp8dXQQ0
IlffJGOQLu3Jmn6ZgT+5fX8Er57d0Ln/Gfjvy0AA5o2zPf6nfIrr9fjIMoqsQqRM
mr3LrC3zwiqrZCI0MWRThP/CJ0c6sHOwD6E9fd01Z4WB9BCZqeZpYVub5TVOuPgG
CgFEsfRslQAxbZN6IDsnHWMfUVt5yQQ+c41vrJzwm2VE8v3ygj6cKd764UFr60CJ
BHRxuxUrk5XVqHDXTWxYXMcRsa2TY2hTPqRy865T6TuUnS0nYtwP73+OR8AFpBPw
NZTFE0xcERAxXlsQOjxDB54xaIAPvEJNp55Jt+8AWmaON2/A9llupfaOqO7MUG4j
KK5InzQlXEsRy38Zi4Xzz7leCIUEy8qhJR3YwgFS5JwqAHu1HNH1DPL8nS+p9+KJ
wGGWhTPX6+S+bFsezc5VSWLUP092yXVq+lpzqF3nvH70qPJLA1rtGuz2cxkIseQJ
LK4e77QixX5wQpsGprHqriY9ZGR90mmK8LSVWZQlImwtda/U1yqZrN9hp6Gau0d4
na4onQ19A4+9DYfD30msqjxrivhehvReQV92F+46YHg4qdLODbMBolDQQzcsy8T1
vNJ93X1EXRQhLYVVuTfOmCi0yZFHA9zOfWShL7YCkWSLQwNNtTSczogNc1JDrCLP
o1cP77tIfL5QjSsJgSMRE0kG14BZ6t3mpsnP2Knglxlr8Cg7M1LPL4edcKtKlFnn
9R/omHlDJS96HwZT6M1pohDEnfsRsgcGvMUtdmL7+X3ZaBUQEFryhLwqTpGia0kq
cgralSC7c8r5weGzPHfmlgNKXQ3oDXek7W63IKSZYTtkyZFloByp1T52274Yzkai
O5wStU21P8D3Tp9vkJR7Gh8wRAmznd6ThrGtyhE6yIx4NJc35jl0s39aBJenob6g
hPeFT2RI5hcP4uBasrtWZR97tmTwNS6kzUeB/lxvG/AasUphz7MfGCzc6GuV0YX2
PSmY87+BrJV7WcgpcAPZHJyFy3M0uR7I+ZzxptaOUWA/Ao9u1BIy/4n5dRJH+l1E
kRn7ypAS77heBs/9yehl3SqgWzdvBuuXW6jnpZZjUJenuZx9mIxuPl0k2dqcWU+i
ADtE2pJ9JLrR1OW+8akSkqnrlYC5dNR6J3uSOnU1qnlqR+/I6FzRCeVogowXo3ze
NrjHutG80ueE/PaAo4W6jUvOEjerKLLCUiyQMfhhHXlIv7WFgOhhogHn83DBbkaz
Lf2mPj8kO7ghVjwz0AyRUKnLpEt8yKO7jHlVwWuoMeuhWXvLBvgWigUcIhvqqLx3
p+Ft9tNHibNfKwCdxVhLAbDzGh03S9NfVxUVz16My1154fXBLwvCetS/5Fb8k8fm
bDBs1vAvBp44QM1clmx0Zab0/Av3LCBj/5qQeeQuMFVsGoxrl7KYKrCoXagehFpD
mih03dr75sFZsLtUPlESR7vu4lUDC4+87eR7Mcynt4yDTh/GibJRhrFpBN0+OpUk
7V2unlnwap40TJSuy0kgQXx4K4D7TxMTcd+4vktNMz2uI1yOK7fM64S1KB6CpSgX
Q36iYXdlVLFvvpiLDUi9Cv1VGAbgJiikYcHaE69S7qRd/yVHAgpyb0nFrniMad6T
SNWuHjCHid14ESJ44mM4TQIO0IXqtLPhHt963IIlTmvQBOMTJoeJIusDIEcx6kE0
jjzkydYbr43cLbi0KoZAD6WxupFCDn6xaXFG+uvi6z534UlZP529fni+5aSHyANx
AwUrWybW74n1iPRV7TWFFAtVCVmG00KLEct5qsOEeg/PQDxiXg5IRjAK8ybtvm2s
gj5Kq0p1LXXGndi2unzDNBE5Yxi0kEEnQXbUI/YPO2Rl9Xu+V1dGBS1dq/gXqAvZ
48O8/MrIpgtgU/U9aXxJBSI+wwWSYBd6LnRilW8jtx0qbHItYguKVYJU6aejh/Bk
C35IPjoys4+s++4Vp3L4pAMCwvMoX656coEd+jnVcPmb7mP3LAAM6Vj8WZu1Xo/G
baGsnm43nqzjCSwVph/7ydrvEaSBAh8DZn1RTnpD/ShFdO4ubUJwENHD7YS9d3AK
i4nnavF5+kM/2ICuW77Ibg/P0Zq2G8UM3Xs55hJ26Ck/ix8GXFzdbj8VaWlJUwxJ
4Bm1QHDp4o+00oHunWH5IDMT4AAdyLQNBOuqUKEJMZtIJTfx/SwHfkRV0Li6oLbf
Mn6gSLIj9dzXC5UnFQOdck/4HtFBQLDvXG7kCp6yceiDNrG2Mag6JLk+yfk6g9Gx
IqcDP6O9gDfmkVaPFVdixNNUu7RvRTJ63gWlz1N1neye5wkQc+0xoP9kTij4azy7
SZJMTJyFbxsKlQ41pQR8r5evueH8P3BsipCje+rfZUbGTk4ptLZTnNkIwtrTUSVn
fJAkPULlRws6L3UnMQcQjFK7bT/bwtsLsrUfWJM2dm8vl0dhBDCUbzPc4/q6R2zw
9480fgtfmEZhVWGcHucdtzoCyM9wp0Ch93PvsfOEvdWUoj8lQOpCoSo8XX7VdErt
7IjPHHDkTsKJnMBz+7ZVn873gpKCHjtL0fBVz4Wd7xfnAmVSHtzHtkjyDjkwbzYj
aBvHJr1o1Mv3R/AYPSCR8QgORQTogR2bfh73+atHFx1LH7wGn83ZMLANgsEvaHtV
cvWwYrxldoSRyRZHV7HbeZJueTJ/EcJ4XSkPQnZCcHpVgUbRJ3+1h2caoYDun2PA
6INdQFJEoKyb9RwDfLbVcDyRQcLcqmjoNBT3kd1DwjLchhgtPTr5rJwAX6R2QTRi
Dt4lbZrgma1fHsAsDCC6YJpuYroZmrxhjXrwxMX8wDIHaXP2kdW+X4rjb7+w4UE3
+7eRHTzyjk5oHW5405hoObYpnwrczK7vhcwwJjrsgcgGRcNInOf83TIrKA/jWpGI
VuE6qAOaXEI+UBlNDs6cKIfqe0jfyqd1Z3h43QJhDbSEDHyiUVKG8F5/tMDCeU0h
KwHpRx9eUHCauVEfmOn/fFke1Mx1/pRtlefHPlq6hugfrrW0CjqHEs5diQV3gVws
TMRotKARyT6YV/K38BXVP4h/yVUvuO5fmwzIS9htZUxBkTAdnZplL1ccIEC5wbQD
sQ7+5wA/Qwy1oWqHUzf3ikgMfKRDfOmDasBq8Utj94+cXIaSEW1bOEJch/PqfFxE
l8lvC7kGd40xw8hZtbeM83IoaEXDdEIdQAo9A04uBD5+gMgmrLHPkzzSkv/OL+fC
znPZ8OGgrdvDxMmHbxBHSxpeFgN1SVBkEKnTDtMgLw5bzHjlthAnY3q1coe4BT6N
myxL1UqpEbPhAoQnHppCIRlQgc0kDjKAwlaiwvTTNNwvM25N/OJoIyXv3PdOwdgI
D0UWHhvsPs13ohoUrSaqctO9eDYDtyY5Ig56Rlf1A+4YpPZMYaOKM3TtQnoLSqso
ijl3SqULu4Vfuy95A/1AlcLYErV5S8m2OkdSJABf/IMSmWXyToYDsHUGjdVX8Mdo
5TeWm9TcZ7ViOYTHT4BFmWLE1p+acLgTgptVAY1Mwa3ubA8NsPPxQoAaNFYgO5QK
zC4xKZjoCvhq1/tIkgVTfdUBMyWG44dal4rPIz92Zq+LNHOOax++/8ZfDyFp9GQX
qQBB3jqNFpD9i+L+FPZYY1I201rA99JHeRlODEMXvE2NgkE44JC00V+XHNXaiZ2C
Fbigq7pW43WIa5hNwxEYX+DaMNBscK55+FQ4sJnw5WPpOMwIugWraHgaa9airSNy
Mz14YgMOTWyqzB2Zqk/vwpBvxwFs+phMjrOOjsob6OoI8k8FUPbq8GeLYi37X6Yl
TM+P/IyuLf1Zh8Rj98fEHg5hw0HlU5vAqQg504J94vZGsik3p5CfKik0oFT0JZe2
KL6t1MNBs03aMHRucOWgy6T4pb7Af3kv7mnMrFlUThcSciO3gK8lyjGoDPhvsXIv
BEEAmJecZC0VaSK+8/Orpd2bcfUU1zmnKKMxLpdG7S0oRy13Xg5nEYMkI5XYcVNx
CbKP0EMZt8HqvNOcqwkqCrGSa6cdPWRuiA/keZn6CDd2SMSPraE0eBuq7LejrrpE
ugPAzMV12JIzvmFVSE84c0cnhka6d1Zz3ZudmTQ7ekv47s6xzDPm90qz6/16JAB6
o/gnk5lBk3zC9f1Wnra/DCGYl0RR6zVLBXgFJA8/5v//pUOVLDsnvQ/YMKpB2XTr
qsIJL5hcQdqCusj38tOC8NNUl6SINoKu7xzqUpCtfjsGTreFnIrdmTIzoArzFfX0
UisMmRZ0DxSVjSok0KI207Zfau4Ue9vOuod1aNuxlcD+fk+ESrPubDjPKlsxgUeP
78nU8JjgkonkZOjSlF3NkzEy3z0jbMnSCkeSgD6mUUbYY7JjUfgFeaVSLnAkLWBE
CZmYocFMjeiTbjU0prBLgOL3vCSmIypzB4Yh1mEnd4v7g9mPvkDDuxFJJPhnEyLJ
VdicJXN15hw1Zsf9LoO+MgG37xjyTQo6iIW4a6uJwhZsly73VB5p94p3gwJ2wxvK
sZk8X2h/OcsakGBocZBko26UxdGz8Yhkdw8fIfJyd28OuGCD96E3SXd6fMuI5hjo
ehvIFsdimEr01RkykJq5qWfTAcdv+9y1uRe04qOh1YokwXl8s0hFbwDiqIhRTUYx
sbz6Prl3EZF39dXUl1FyDH9t8bT+tx3DvmsPJ2apg+dPWuhcQNen4zwZdcyx0NDl
H5KHVUw28b7dWxjf7Aq35J8Cwmyuj+czUEIGNanntygvd0EsY7Hj/sBKfBvmCrHS
or8K28kH1RJrGvKMhRL6xNX67FinF2S/9bbK1l6qZpEKKUUguCQBiKme8GJ2zSRs
nltN0Xlal/FyaoDmII1ppFeod/ZtkZWJ1z/qH/ABcpapJKQSZInz2Qi8nY44cj4U
pgKhHwL5dwkEPiDoPTF+Lzxyh5L7v9c4toq8RQ2YPI4syrrTy6Q3VkBNdoHIlRLV
1jM1pVgUd4oR+L3g91jQ5Jxhmkju+nitmT0t3pM2CAr4cqHi2J0fhIlzkSobQKro
yCxoF3fn9Dcj0UBjeiVkOHu5Z5I29loo+PuCyQGyXUGqz5vyzV9AW8YEhVL2ozyj
lOdHMjS9ifJqFVPHf7ojeN4L1h345bNJ6MRw5x0DkzZeDLm7YXGt/Xghr9fWFGNh
2GU9kAlcYQeg52f5hRJYBGUwySw1mMvJ3AXdDNG0bmjz24clLf7Id12e56c65cMc
nlVOm3wObddgBI4on2RLqMFhXYY90RUf7a4AhUK5MK7/MttxUKWvJde1qBAZTUk2
YzAv1StyxEDiv9ZA6WXPhBJq8KiZxFJNCh0y0EL+LrjtovgTAW+So00/FRNwzIMX
wfNo8PkBwrO+9gpE/zuoZJcOvaQl05tUDlZzz1miul+ZZDM7+BjPfYHtBzIjL5TX
DuCNVSLZG/2qZ30TOClLUJ/9r7ptaIX6yIRszirtOdeF+X1okYu//3caadO6jg//
F+6/EfXn/3KXLMUODZ7Lbc5ETw8nW5lLd0qgHB+93YDG4XFZOOVCSU1SSR+8h7p6
2A9cZtIHxqHimDNoOXIgC3rGm9dZO7gFedq3L9Emny7+cYQDodneImdna6WM03SJ
5s8vQX7Bx2vjTwmjN3YLBBbP6j0wUyDcHT9RkCiY+MBwbt7bdpRQReDKOu4jLrvq
14DqtWW2+jfC+IJBpHlrDffG+0sRsGkFsCV9uiZMadwQb5VJp5VC/npqe2mjzIgl
5VEkSnO+2JlprPeuI4Hzm9KlndEX1T3utYI1Lz1ceDQGkWJbfhfyn2LcG3yU1j0z
6P5D5cDEsgTsTzVZ/Wp+7duIUY1ygcSLKZumY7WnqFoBsdwo26Yb5JBpkTpSNBld
OwkKHBfcvQ/k+q2RJ2+DJZFm7TyuFSRzqYsBFmBbVvOYOz96UhVXTPLwQwEF51GN
RLBAGzdKDEZCC7dEPZS1aqo7vxNO2kG9amR4TVWfUT8C9U3Xu46ShCafqYwKXd/c
xMeYLYC/OBsg2z2crMf1j9gDM5F+nxv16HWeZ+LqTnahR3Guz7yTTfuSrqJSvZmo
kyqVCCoKUXpNHABNwQ/R2kFFrdvCDF650J63z9KYPLi0b3doyO9uMUFHCOrfwvOa
ZxFsGoc8ArPjwyYA84LlcS8JcTpZnCdttOQYUqFG7v3i6wV23whI3j3tIMRa2lUU
xep/JWzlGsArC98gqGSQGWH+3iu1eKAqHij7LzVoH0NVJACaxEUhG1mZ/jzBLJXi
sXWhKjTsP3k1uKI8cKa4tb6T0AhaxZbSyU6upT57u1sOrBT8yczg2YGbvt96rWmn
m+x+jas964Rn3RD+sRzUvdrLth4y2m+rrYFS8/cHCwrTBPypb4TETQ939ps3iUhM
k2VQvAhakiH5vt9h9XFL5P/rc7hFqKCtp8XIikbRNv6Ob7OHMQEttAMYAG5PgYb2
Uf5ntf/oVbP4YRksXBl8MzXnntZva574qbxQIFAbVt6MQ7/UM6EcunAH/o/fVpwO
TDivCSqhwVC7ubmfD2gScyJUBiZXZthYIFnUGfcOMhR7YuSKJBHgVX9YDzLboLJG
c0rlvmGi5EuK235jd7dNwFZhm8v1AaU1u7AQnELqMsh2+bJrs/al8z5GvJ0UytAf
Lz43LdRiTyYz1WtdgOWx/QT0EvLhs1QV4SCU/6mFiayfaMSh5/C1X43FVKI7+FQy
s+l9xuza0EvAf5gkdLHjUdmUoNN1nOkyZ+b3ypchqBOJ/cZPa56lUzn0SXnY/Evp
9fHVFKHe7zbVggUMdsDSdhDQvJaiE7o8rRLX6uR4XklwHsmK0UY+YYU5gyYx8yUG
DCAtijlfOkQSfNcNiGUH0IzUA+vE9e0InkhLwupjMHmi3gW5VFTWNaeltX9OTxND
95FIxTCLYvU5GRN4XVyLLR4ZpPn8X3gMw3LWHBpFwy98oNP3Aqb7DY120YIISSC9
XJ1z8DMA15q4G6PrLM0zrzaZ9QyFqKDrXSVCLos9BL0d0pr7wX2VHKWZQWruFFOy
LslwDCSSZxHLi1xLi0oUBL5Q/F32zkYi2Ea9kWt4tPzzYsJ7RbxO3nGicU8UsSo/
9Or7Kxd3823iygucds7hY6t92KrZ4tX2SA3Q6otxy6SDUh+TYPWVENbeg+oFFhwe
VX+mkqEJFoZg4ddeFSEuzZcRfxAEzPMG9Bg0Ypfoc0DnvJpXNM5h+iOhrw55gJFc
0ewWI4YA97suSkH325bJIGTonUKJ9DfZSn89wrCmMnajLEDqKRl6HkuIdJPbTs+h
CQI2z2Lbh0LSV2vD9huwN+C4NAemqZ+aWMlC39iM2YyxF7zkRhQrT0yiKtWiYHE4
+zcLTO41W2bB5WR46T7jI0Iv1PmJBpnotPDs4YzQflDcQOClkqlH1qZ31alV4bxT
2tJB/Mm4I+xvj25FYvbef4KCZ4JLc41LaI9obLdRM9whwVsDYWeM6oZiL9LEJsVD
2q2ltnsU7mSqTGUUcmmnZhj4fOsDAKbe7hYXCeSU1oAX3nB/8i/qdhLta+leAmY8
cXMkn0jFiz2KJkRWQqaWNLq/q5ry22ND7DKQGCT1UI/lv1M1JjpOYewZ0NNZXBSI
/XnliOk7jaesUplK9GPecVRMitZKcTDRohiefS5FWQgQgGcBLZOiSeRu18w3q59s
4R3B/Bm8jnC5X1Xb4kKGYfFdNwOgACWXG2i+MxCj9icR9huuCk4p92kFPO+VGqCQ
S2njTddq6mdw5Sgl6Xu/XN1uNrSArPcb552xzpdxLtJsUecc9MFQOe4U5lj6u7KW
t1p78qWkZQz5tx+9rkA+/1SetNlE1AM3JaLKjmlMNZfEKfkQwNw9Si9//LfVkQpM
X9v0VwIGvN+CfX1XJOov1eZZTDSPF9ZCuqdqmYaVBa95SbRcIa3I4RFH40Tdk4pm
ONnSDL7zq8Kkox59UgRWOU3hLIN90qZpa0ObXUrURGFstZbpbBGdMNwKvFAbFaGO
UjGAPEjjk0EGNtWN28QtzZf6LCNNdRhFvQyqRBrY5J20mSbtR08Vg2wVlztGmm8F
0OlzyJuyNcCk2Auf8nJrIyVv18gWIxlOfzuTjToQ1AzbG+qQPwhjlJKL4VW42aH/
N8j9BATWkZV+2IcWiCE0uHGzgOa62Hb0UZ4n1DjFUimTtzRMKUmSxgc4jMSly3HD
xDIF6j2v1cAg0yklUHeYW1G6+/A0ut01ITVBiFQSrLl/xcZUGUf2XquiuqcIaQwm
M7BeI4dCCGV4uSl/CBbVOdI4KvUlDKuM7lcE5VBvDp9lMFEt259gnS5x+Y1V4twc
kFUu0MxD1lDmvm2dFiuLL4JLEWD2pY4VaUxomlXAHf6flSW4b83Vpsmd0etaF6H7
BQwQCIX9/p/NvHKgu+iggTcB8YBRxHSOzVC/698KEYKh/+q9F7g3vu92OQICmGCZ
t2BaclEhpllAH6NYUbq/r+moYZq2PEZCKfC55bP2liqI4mSYucsL+uWA5TKaLg04
t4iVjqXXkAst81EVEZyZ/MvjfYu8tBNrFEPS7dOCtWw/E3dbePgZDsrk0yI7L20n
CYf8PtWNZTD75IttI1y4/DKsGTM8CiObRtvGXcz6KxFZRoAnmLqRuv7LSbgDx9c7
i97gs8gdwCGCnVsLPIJ0ITzhoFph+Ryfgg/eIL08irLdRZkohCsuIUmVlxeqz8nS
AWjB1bggigSI0dt7dWZkL6WK1SzIxGDzkZeMdFECgxtF3I40iIvc9jcTLJDFn8az
ROI5HQ/F4OF7Cto8QxHU0xjwsBugi/vSjVwg1Snwko7UloiP32nH4xbeh+tvUzKO
ImAkNypg5DNcNeUqujFathrVTKy4s06M8bH8PLZ92k64vcgRlEE0USatbLpAiYlJ
PDaAiN2Az5QvfP/xAjk/8S3RRarhGlj/sis1UEr6XK7UGjNPnxYzNrjupiqlZHnP
DJhK7EOa4j4ZruEskUHj0x8y0RbBbSe7pb8ZKCoMOdWvWf3DaP1aHqBKCrp1GdSv
FJ3bwrb/kz/Lr8G/5yNreErkw+g0dPhfcgwwnd2YbpE6rOBjePnR3jsx9Delte1C
y/OewhQ9uzWOkVsC5q3zKBFcv5YSuJ7XjJoW5DlCzsSdTy3c6VRQ+iQ8h6RcPSx1
elNgNsAEyedz1p4wHkQHyOUWBj+SYQwsPbvBBChrPiykuLJYvT9Gc3uNzybBN2NQ
adGrulGWaRiAcYTsfhSr3uv3MpDV4jv4GXBDE5ykjtoioMTAfyM79x6v5UeMXs4J
Xdl0nzV7bRrwNCp7gtEYNEmQgZQV/nDsyCHt1tNhELXJGoNmZCUdqUfwvZfq2Czm
/Orf83erokQRHAhv5S9U5xAIOhzy9lFDtHxg4sx0XrsWYji+4hBXpu8c+PcUqlrM
FVP9CpLtmraPWMl2EWdAiqkGcpmn1iyQVV0zmjnQDaK9XS/ngcizsB1yYcVA07UA
sFS8DweSmZrM3Go9ELj+VqKrJySd4et1jR917LHvG+q4JaS/d1JjIrAqy5SK/yG5
fsijYADbGDGVRYFKWJBIfOMiiYEZq0lPgkF1lEH5UErWGnGDAvFtiTZvSurs6lgj
mI2mKPxF2z3pvw3OTsQtWoaYVIpodmnQbA7CGjlEcyawJA70/HbEf+u2tDJxECnR
lcmSsdUR0j6p+IuI8GY0IASIg3GodwYQr++DTvzO1ppvwgGQvFA+WMh3eh31S9xR
VoE+E4X1By9YB5d0ge9NRWttI5nNk3svm3ygRjk6nmAIUIzKcExKqNh/eXAQ7kNa
nfBCzTkHr4rMcfyTX2jKEKI/GbbrMMyFyAfcOt1e+wlxRyuBNnmWUwEqN632odre
V+pM751zVlqEC26SK93zJcx3IQz3V/WXd6fiojBXYFTikPGA21iTw9YGoWRSofn/
oVMmtlaGiu/tVt8EfO3slzQg3dJIWc8GvodyXvrQmOuVVoMVCj/h5M5dN8xEvcZ2
izI/M0ozZRuOU+0rfpgn+EoFpYXUApM4VXxuVs/q/T3PHnROaKF0lxxiqMCsDZPT
MTdOA/KeS/6M2OTGCzE7e4Lpv38USM+78yw3mNBO9BvT8AUnHg3GoqMNY6IYMC81
g8K/ReL0XDBNgLNzH/K9DkkJ5WyNBGIohd22WwHYVXXBKSZ7JcbcoMgoMCgGalbN
c0k3WZIBdaULyivrthRp8nDR2ZHu5dE6aoCOrG9Q89AA8xafBUNhiRZ1Jsh1gSpq
J/iODbPwTrboGGe1FlQrCaWLPAcsdi52vWRzje419v4k6ORtkztQJojgBlPFU7LL
fnQH9Akv6ADxkjkFrGKI+nsW+R1lUsZp+/xBauXf7mVRGxnAhBc2MJspqTQaUo+n
DCkpiYrxzz8anWMy2wHi//XlwD/+E9ks0coDMiIaU21C/jVr/EwVChU0tsnH9Rg0
8AGU7F3LN2Trxhz1VzfR83xqIMC0+z4EFS6vIRZlgcpI00YIqkQ/oZdUJKokjsl2
cvSbT8aBbfVmZlEJRZswM4bsX6vkd62VegtFqqUbJPXu70Bqrc12BCYVDqIlbFbf
VtV46J9ahMiQtscVctl3I/UN0kD+JXC7AX0Q27+9OxFKsHo/fV2ghgcWhdrpCMiX
GPO0gUTeU3VhANTcy+NS6nmxO4UKG02FIMTOO1dPtwtBzk/q0X89SbykfbYCX3YB
8gT0k6VGSIrZcipS+GkmW19dREWCv/OBZ91Jk5HKmDi1WxLFCP8R1RAdlRotnGsG
URIcUe/DSkCZyMhMcRaqkxkxau4XCr4z2DYWT6iLKC9Kj+1SoLsqGgHFP3KBpG4E
b4X60qXxssVsgIi5lWM+0sseUgp8ScAeu4hTfj3v2gFmsBvMk5yeT9E+up75BnqM
a7jKyVvEwzqqW0hcbjMkcm0rAsoC+KDHPxumlMK75xjDRpDnsXgOnPW1n03TAsBv
xcDvbpRtKV2kAP3A6rOJR3XMx4l0F+ZP6+EQ5vCM7M5ZXxgZoiTwe/L5lGFEZa1W
DFStbGaFR1SuzScIQUf4KZjPlnbnLSuwfaVneiUSRH00oEn1AFMbMi4fuDfVV+bP
5cER49VgdhyAia2/XLxhrH9sGl6qy9PDu76qlEqfqlq5eaLvD+Op+4OzwXbZ0bz6
oTe9qgGPDUZLXO6B3QZ5WkWBPUUGu5Ic0BSzU+z8uYszARTfdfDdhL0pAwLkpU6i
1v6UXCuIBlo/vMUuYFsh1QDMN0/EZ+gsEJztG/XGaHM8NUDTNbTjn5rQkB4iLdZZ
potzTvHMAtM5X144GL3aueduDHLSlRUJ5PPVCMFRe2sY9DGCnVFA4jSfuKpXz6tz
rI/hxGeZ8KtCtp1Ul/EkVwkr1paupRsb6z1S6+2hvuyXVHcVvMBPJ+Ki4m68xIHh
bfzjENj+Y37yXa/21A5EXRetjq1r7/kXNbcsxHT+NIyifCXcutkMFBtUd53w+dx6
dKFXPKL+RiCsbQWE/HvrPwA+LxMM9wjuwIF8REhT6RDCHfwuriRrSVe58IyJS8kF
tYatrwfw5dqOm68uYnLlOjtP6YMQ6zCEiVnWf+tlmNo0Zro+bWwOxblNid+dFcMY
VUq5E0d/sspsU4CB2Ue5Ej4OShddAUngvwos3n0jSGlo2TD3mAYeRZucZlMdMApD
QM6vcdlcx4hotrC3NBm7SiK8dSmiUJd8vbpG+lu68phaF5Sn4GEE5qqD7XLLjiaQ
MoRqb9wGMzwiPwabA+T/xUG6MYm6Nw+XLa249HpkTkewbw4l9Gl1HPrY3oaIwInA
C5wEmIC5hA4W6ddlzxgZeYjirW2vCJxcWqEH8w6kCDlyne4ZG1FbqDBK/zAdgsT2
8J/jXqAKNv/Jt+h+p1H7cKrdlSnj+KqvUTc0wdbWLsAFlaOXNISSn+TzRlKPGzZP
GrsSMGaRY2Yu02ED9SXrsYAVdDFZF4Oqd4b1DfgYSIzZ/uiwCqPVv8Y4R3J4xHjY
Uj58WVDRnrcHUk+IMCy2vexmeRh/WoLdQ2q9kdTHzk4LdPmZSF2X+9zl+53D5l3A
gc4ux2BiYHpRksvs3pE63agxdjUtu1fTXTI4SxWpGXx5tbGI0045/Ws/zfbJpz6Z
2OccJet0F2qplkiKmYHsjiJmK9O0W6TVYNTCZlWW5vkb9UaP+LqhmuL0wZmpDqHp
FkzG6k9r3JwN5xJSByT524h+p2ol+APVyErDGFDNGF8abMG3pLTBV8sMYbZl/M7e
vHWT41/ZSOiMvQ6lBHPJsVBhq6FvFsS84rihsUAQZrSZ/mpT0Dg/pv1Yqx5V0Wgu
jRkOJdoFaOdohXAGbewbcmtL9Be8e1li83gDcQf+X8lRdbzsszMn4dvAUAwn0Lyx
vIwfCV6Gzk/dydNRClrKWRte2AOy3C9yDohl+POHv6NdAP/4qBjPkhHSaLlCW9gB
ZEkeOTrVys5yqYtfU9dEgL1QBaC2OTXpCyeDkaZdJvMK9Hf06ttIq5T9AuZw90Rs
TdAREaXVvemMvs7/3LPum/S+jn49c0S41TXBT82tHmL8wqaD93kd6/xJ/M+dqeOM
p/nPjgrTRr9M711jbcdBlX889KCoVs/hBwDIP/KkCAtXq8HIuuKeC4RZqm7r8Kna
GepBk5BvXztRSbKeYmFblnwWyzbV3pmWZ4BIT9F5lCPKqFQ3sVyZifouIFWQcWSe
WnbW67aqny5nMjrEfy8FlMkRvpxaOAFZCilwT2tt8oSqIx5kAVzQr7mJJveE8qUO
e1w0TMTIeZnUsrZzmZt7eJgjr+7sPW+bsmjWnKYhbXrn/WPZzD/dX73wyndTtB/K
/fQBpGRgqJQSiixWmS8E7hZ2K9m6+G8HumabG0D3J0Sx7/10igBEe9KVr2AzFiJh
K0W5pYbXUHAc8y2tEs7Icryb0qQWsqoxkFd5SaFmN9fws1AuY/uQBPNoU3dRebyW
wjNttl4CSo9Y+OYZORNW/Ye3py7s/lR/wwePjeGccBsO+ph8RalWaARVhkX+bdcw
5IVCsUYBYwQuR2AsmP64dR9hutfO4EDcwXb7gx+YJtCzIMtX/dFjYcxzuBwlxyzv
vGRf1WDbjxiOVUi+tI0jMNw9uu9BLc4fTTGfUI6tO96B9vE+CjMjqW3SduaZm1KU
5gSVqlkGVmzsfdkXh+npwOX7RRKvlSnD70uSFJUeRWubWn0bdeP+0t3P889IRvRN
lNwfGLgv/jeo0fkhl8XLzqjJIDpVDsBZhx8LOa/BLCuXL8NEl4IW6s4idG0BVmy3
g8ESy1y755LaDt8q5u+8DedcUHqESSUwbs6V45yEtgnQEkhImLmNHXPRTLauvMvy
IwMaqeWVFS9JI3Cd2H9HjzcgNNV+7t6f5TtBq9z8aUt1061YxCshd2LIAkWdJ1Qb
V3nhA8+rcpDGGK2p+Lg6whCgQo0dZ/06NyZrC0lZtew0cgxKzH5JPxZP/TqfLxKe
CKyM5m4ZF0ECN57dXweA3JA6pu5njY8uHx2g7DEwuUT51yWvzBcBN/605WYoZ8Mt
0ir1QdcIV71WkcEdc0nxuNEEy3TSNFnzT1B20bzPwYyepd39cPaZaimJA/ZJcKlv
Cakp09tWihDBRvyZ7veYHFAlczfRDOrDA5AGlrmtBbmiSwG3pnjmJtHcl22OPZ1z
OoqaUZ05GYEFVK/WR/8F5GWNgh/ykOG6ZJR5AJaCOQEX48bl3z5kqPMDC0sRxz+x
H56EkkUvErOxOKhOkxiTHRIXG+bcshDEHlCw8OpHqUkVFRE0NTiW2h+/F4iHYqWB
PEcU7rtW3t/uKccp00kViPulw2EK9LwSlllFUzzm10dOjdpdGioFZIXprgDMDq0H
m41Xs6+vS5cYueTDmJKEBwhR6l7RXb74fpGVr3pYySgn8oOq2OOzZp/EGxaV+kuI
POhwmL+XQvcokQ4qnaEgu0Y9yBYX/ZLOeRtEawOQ6mAHwKPx8nMnuxe6PNCLAhed
Fz0I9k6UPpaw2RJ9gDUha6F/d27RzIxekG/hMD/plBUyfe3yLjcRdcMWywFzmAnY
y0UfrboDuFRqLYG5xFhei4Hp32cxOBHUn/tdNl8AwwkzsAtPEGBcrCYNDtLOqvhM
ppJ28rQBh7w6eMnRHtj4O1g7SK+gYbKC9MPntKEvXRCLMJjYJrvp93AEpvCGx74p
PPMhEEbGtVwtXNk0sext/oeX9B8bZvZMi5HV2p4UmxISbQqPwZ3pNkt+jJw0ZbyN
ZP8ldKtlvxhWmj1C86DXF7BCU3g6ixyb/QkxvYIz3MYcjQGphQkzAzZifaCtgak3
Tpup/h2La3nBOnUjzCPbXg+7I5XNdNQevne9HzBRRokaSRaW39HMFzP7xNrYiepV
9/MS9LxPWiqH4GpZ3jeL0Ll87qUqP4RkVOhiUy4nLMhmTzuIU8VywmX1YWwNqdpU
+zYsbIGnD08jQe1UhyAPy4dP8bxyKNuTajnriBFurEaGEIKeFb/7jox3yqal+/4P
9/ljh6md6JbX2q3ION0tAHhEmK+UDb9mWEA36O8TwZRYNmxz6TJ1Cygj+DoaseT7
5CRt1tYl7RV9Wi3ypsNCUHRI9tW7u82XuX7frYLhJhl7cFeAg3XPm9RRfMTE6Ufb
k22x/en0+yJqL496fljlLeg35SmuKgnAbFyV7ynizjNVWgmhHFxDnZLBuN7hKjtr
DRjhFe4dvEWa69G5U5zn5EZsfWAmcgBcBsfdqMCuosOqrXlrZz4qTZ8yG1bbxXbR
/gOAGoq5aloOT92y1iDqF4julYFF7r3GzWVaOt6c+xTViLTnIjxvZexGn9DBZfah
05S3gDbMokFtCWVmA7y3E6JjYoibo7+K6nFY+JFecYFJHtJVMxUlHO+/8DFgCJA+
mWbm1CFzarhTjZ6rpZSSmxo86+g8lA44fZfCNjOi5qiA/Bw7K1Uv3frAcaYKGIHM
M92hHRwy3phVsLASQXJGBr2slQSk3oFUzupCCrjf5eb+pfso3/VYJP5u713nVJN+
tQKhfhURFKJrCqbDDIsfrEoiIPEnbR1La495QgHPakwE1UgCaRPud0dtIBfMgDsa
g/uSrE8RZK2FSjKgESdY8T4xqd0TxwWRbWYJHL8H01n2GxdA6EAUZRQzl6B1E1p2
KYw8Z3VzdpyC3qVQzndakPEzX4uC+ULFGLjBR5ID4dcdM3TEV9IK+xwR9xc/OYXc
9SAK9V/o2NCmbmgWLWDJPCTnfLsciNvMdHMBSnUSbbxtaKM4TH6hLeBBvQFW4H/4
AQ22pspXx34s+NZAAvEIRvPMDDJWVmiYXcnaxphc0VHXS3CMHcolTqFsjvST0dfs
CNVxaL+GNecaUSGYc2ST3bG/HFuAuAAWUqWSi3Gx/fmN9MpPMfXxsSHZBLp30SQs
+jzfiVzRDXxmoS4TgO+KqTUmYHUS6szkOkvAGZ817H6ZGNmc7HvW4lPcvYaUWtg4
VxpbNT7Uo2kTRYQIEWSdFJovPZfvWuV/C7GMkOk4kZB3ysskZn4V2PuZoVl6knVz
/YlFCUMNCCnUdta7ZvxOgHqV6flsgG7CLsM4DcxEq91unZogO42KEs5hFWEgoPSS
cHrBNidwETZ12Hd6Ez58Z7GeOFMZGAReui6SsKZu1EpOGlNp9ILcdhDbcGJj3z8l
UG0KFEOxj714WM+UxsWD8QgDelbYO2e+OIAQVbLzduz4NKTdUkYjJFdnLu7A4wBP
GTj/l0Ww4duOnPmbzJf3gcHtjIhasVHET++79BwbUMDXLD1VVqGWrRwPVRhXOIHa
bQ7dhA+9bdNzEbSDJqTwilfl+iyq8TbSI1f44/V425TiwTSw4vMp8SPvK2eGyMZ1
xlog/C+4X6atQuDSDXLI6bVn9LOje9kJ2IjvI6hTjOcUfWaoNbk2Awj3OjBaBqS1
AITyxE6V33gUJwLdCDLewa2nqGrLuv7QkYh15SACZh3CVBHyYYcOGKTCqmuYkrG8
FueAF3h9sZDzXaNW5K3Kx9a1kX/ZfQj8uOvVUF5QYab+mDqzWZO0E8ih0OkD6aBU
L4r245zxEzlieLZEkSb6Q+ZMY9WtN+caIZRQIciRrHtIC4mXHe0N8E3b/QltbjgP
KLU4JkLe53O0981iVWU2UtN7VTr8il+j0iEdzuDtC6cJuLSaM+KM4Ep/44OvU4An
KHYgLm/JuXv02j7/Ul/nV0E8NdLXVHKBXucbqCokpi0nGt4sLcYy2zh59iJfIBha
gfcNQK/pkaaPp9qjq0oJi9XFw6c03rcJUkbgZJJDlS1Tda2RgFRfsiN9nsopHidS
cVYgywiQuDnpdkLF36ptes15HntEh4BShdALzRHpl4ft9tLFqYVejnL14p/Wns4k
WSYKx8xOOLDXonmS7/tgxltsYHf2BxVUy6wY2qnWKzwOJACbv5HBKx8OJVIxco6x
tTNRkH8ZL08pxBCzaBxmgXi9vunbmWFApgTc4rNsGqwsBZH9glGHZOtmts30rJ7t
RhpPtPH0T/5hlHih7EHswXHbt6A6j8bVGPnV3JUkUKoH5UVie6O08zmU/LfZCwhX
v1pCQByoQm/d27o2ndjsEWtzuX2HY4LbrB4Tr1HsfkYfo6rbu1einyI9eCnVHvNU
jFTEUXk5beBsoLgtp4tu5pZH8TPbmsvkLQil8UJfJXn4lqEx+N5xIAhulyv4dvst
YUbcsyrvHfp1eShQfkdyHKBP8GqweukOblymDOjQH+CrNjqE9aP7D535C59quTiu
FY2LJcoIvBhScq0bk9H0Z4usJjuUwJRUfBz7D0bDtI/j23Usy6xsHk3mTj4MBNMn
WubGgFA2+zvf294d6RV1olAtBlmsqI6S/eVftQmJOMsmlpnw3YdgnJBQ/t6nS06S
JzkBC0ikNYrb+DBePzPPQt4MQB4loOk5WoKjhdmuSHEtJGRrEbtYcWARkAIEfPoo
x0vIQiKG9NwvfVhO4fD+DbxbRJGwjq/FzLvTP60LpKPJ2/pJ8n633GmBUnIxH47P
dEGHVL/A/hgXkyv8p8tDy4SFTdZs4ADUNNyRmfpc+xMEhWBYSQj4Eweun20ANBW3
yxAphWF02t2JRwpy+G6nfOoZosUGRD1duJ5+U+uoAXXaxwVSfS8ubw5zh1GYEsvT
EIAfWbEwowgk32jmmpmgtUpgosQ2KiA5OxKFpVzwuvAv0iZ8PgmK9On4pKspFPRg
z2E13vqC2aAGdcfID6b26HJh10L9rDjr9RVvk8bw8gxPNWG2q7EYdqh3k90pHkh2
Wnmm/F2OoNIcUlkunNWQBDzdepjMVXjp41+sB/W4Fij8hgWNMCOYaIhD+A7+Dsmj
oXNgaYdQ3Jg9qSmLWI8FOkN/deVjXtRU35xvb7wTJLNE3NA6zzGkTQXhmgAraIDm
YmDNFD+KN4z3LIlHK7HSKwQGzL+IsOp1yq2Y/xCa+SKtTwHCMYbUAdV6147KaE0f
VuhZcPnBtHzJDdHiMPkRVODepP5i3WeeC0D8soXzwU8zDJVdBGIJT6uYVCYmUgj7
3e6B1kUNXJ3C3d7oEV+fEGzMRHTzxtfmgzJvYXV/XJGtoaS0EZN0NTUNaA8vTqEH
YYyez2pgWSkzTB9vZMApH3t6fZIV9ngtoNIdYXRiTPSeKajRFHF+/EHIrnLSHS9O
BmXn/A4oRUVcLtUs4Ej9dmaGg7w4NnGcsVrsiwdCIvkEoh+DAcLGF5EvfGFUo80l
TtclP/3tkFyYarS1BdC8OzcasGM6+Ke+djWO3fzZ1bzwAI9LCJQVmYhZ35kB3Es/
UbtAkPIZrjmNWkv35TkgkaWou95bF/YGIihqc+nbQ+LCNEahmektjRt2SBz+lQZu
uu8ytPv+69YPJnA6SDJkxw2BjbO9iWM33NTyvJxxwgHPlERmcaos5QAI6Pr8FjJu
mWSJK+KYYQWY7twhyFNcUpqWlQXbvAUUEfn29yKQPLRE7C7MoYlWmaBRgHMbiWWg
pjTt51Q0ZLspaoTKBYsTOTnKvr4Wo7gpib1dKn1Lx5rK3nHjfYiDGTGc0619wW3L
X3v0cybj4yQBIfuhYIcQGg+M4bWo2L3FZ7mqvaZWSGH4o0XHlBz9/jVRvR5/3X3G
YHxN+y9P5hs0sh/dM7nCS1ATMclR6GWuFCJJwcu8XfzsQupgfPf+ZkfTaaqIUAEb
9dVkKSlDb2HAvoOZ4apyY2/KPlBgK9XDhdtF6CW5qFt14ZOdM3eiIy1wl0RiNaAZ
nxpCgAMV1OKy+A1VSlJbmq1MBH91wn6vhAtLet4As6hdtRP8iMwMg2aRGLoB6JQZ
ryrpqZ1NDx8HzggdKiTVxmBjpylXnPvJMwL8GeITy7soe9//1C8GgnJRNH6TqahM
/sQHxZMmcfbU6Xb3ouazTDQY4cv2+nkpBipzTFjjs5eP1J9IPYZaYfppkvDgddiO
/ZCPtZRV+Ie1N1w+1ukVN3l62pqLOos2lQdq833Q/8lFNFB2YLcnDt5cVT2iqKV3
goctzjAt0tbVKxVOVLHbvEst7blEYqzhRequUW1OnHybhWu4PZlFsGTQc0tRvg57
rmErdYMKDXy9bz2h/hatq52VeyF+hHrszJQIv34MVDcsEonJfRVws4i3j24lxFXC
kdRKdjQKmU6ta8fKKDqmfg+xDux72bn7H+e1+w7Q5F7UnSLZo6MIK0F/f6l0ZJkz
EFJr10ZdAJrXjfK7b2hX1X6posBhWmbUm6IAd/myOo1p4FT/XpMGU/AijHHksUwg
bq6YU0pe5WNuQgiTypDgAN/m8Tck7n8+Tab9ekO/i/1Lm7qCy6d3TEbX6NmVbcMt
eO/YJ5YlqY2TKPSRlhJPwDRHthkIY94NpYf6HyLyIcKmBVwkfi+ERBQb9ICSl6Pd
YDpM7cJwsFmF6QhwAmyvKXrtoZtN3h0+AtIaxm8q0n/rHRh5Yp3IUuFXXaxnJ2sC
59lWjZcVOZFDhKimqgStezB7Lpjt2AkMnLwdf7ZvYbG4K0ZvYfi7z6ruDCCvcFof
ps447X7KNcuvtYJP6jWujFRWzWb3zQQjE0zeKW3NmdaWmqC/sCEbXxpEE3W+WyPZ
tIges+Z0HYDou1XwjnzMEU/dVQRouQrwLAMcsbRBPBp95p3ArBTaSIF8Z/1R/g9+
6odZ/DSxnoRQ37s2751FuQwMRgAG+0g3enIkxQb21nrSnbbgSwSpDzbKE02ba4Sj
c0qIaYifmtr2BpXUtyK4WLwmouGuglW6HEzo+dAyE7bkv6/Hw0j1N75fsBatRd9l
Wtes+MHltRLPgN+dFw7I8qU/Ph4TQQp3seJITBlPKy0t/bGbArUS+KT9n/0fCoVn
o8pT4jr9d6yBZyRrimo7bFg4BBIz8S1u8aX4+at7yGcRLSnC2W60nLieaFs6gisN
jkUz5oqeXl/4GURNDYLhBJ9bczNgioCp78j1AwqqVW2MZCbcMMBUwZJ5s7jJ6Lii
HqJTRD8KEmPo8Buu6Z5y1EY+Yi6Y4AcN2VevgKP58rMRs/1ZY9gKB2MOgo+Hz8zR
PXzOd5jOaKi+gwDzaUzhEYROrY/6u66dLSUkA7pKL5AilA+eIS1Fk4EVfNIuaDYM
ikKYIxN1p7kwVr6ilqmi5SE4yxHqFH8CL+GIigLYoWcK6fQzbEve0GNB7cWqx/1V
RUyoJVPlQW17unyG+WSZS5q1EKf05VLteAnl07zXeE2Sb9q8i2MZQEr+UWVXCxAD
erNCbRat/4of3MZpxJTHrjwcVRzvfJXuay6yYzAOePLfw8TSDUrePKIgeShuTuaI
ntr8CzV+5FU9SqaLMbwigIWhMNIjiOXs0o59Lhi0uXv3/sZ6VdEw+MszYI/y0uJh
rLlxwZVGhGyLACidZic7LK09jQhM+VPcSHS+gjYgZRJWctiAQhwNYjKXEJM4jutL
gnHFYTJHgbH6CkUNJHVhs10RrPaNdih00LpWUuHLS/dDxhg4gEv0wesDB07Qhf1/
/WsUvrWi5Nh/T9TgeckPS3T0WzXSBD+LXnWwslRKPzTW4eDJrU71v5WmLDRbaCCF
qQaowucJUHDyRweceKs8kWbZ/zR1tF1s0irjHIkHLp988k8AWN0iTnYxNkRTbzkM
IS83H/LK08DRHdHQ8lt29rCfPbfNa07u4unstkSQWgfL8oHPl+YAEujL7U44x5xa
zEh67JCT+yLQVcT98/efg5YhC1GQ/f3hgmcawerdXtV4mGIv9KxTt9qEAfcQiCn4
fUwYYrGyp6R+p2J9wfMtD4wSXjaPHKDJfXR9TBR6dORVJ4SNbrGoa3jviVkTVDJJ
OPDQbcg50hnjg20rNLPv3f0YLzlUCUYdvGQisCbLPhVP8pHcaGoHlIob5YAqJxnU
r224m3o29Qm6KsnjoGI0r4MuTspc7JBm+v4eVKzDzd+d6ETOGKEfixT6g8Vh+kuv
OJR8Tzf62vyoE6oX0W0h7xmN9mosmDNnp1dofOmsqnM1BrUqKRtVfWz2Tlxq6yd4
5AKRso0vXog2jFNbtzDKDo/A3EE/9hjV4E/jtZLv7DxFwXj+JJHuMpAN5sdRbxOW
Eww+7ZO1H9OM0HNpz/OcItoeFYPlu2v/N0y6KdD6Es2OSRMAiS5Buo9c3sEoyPJJ
N+bM3kafMHJOHhMyIFwPgw/uedTrz0jUU+zrNNSJSciNvcAmVtCzrOK95r9DH5AS
CzUP77tBrOFHg/4P6s32uq2YMRQJJUoEHWluH83vZx7nfvF91/qlttlIrvoJeDYz
dZkCWZBmDHQRf8bQ7GpWs7jU2ItcZwK9ILC3s9sn1PAQYd8sCnbrquJ8ZH9GYxW8
4Itf1cdRfFcQMyCq5R8pV9tCuEd2Qbj53GG8xGnRffSfgfrXlHfOe696hJJJErZM
Ka0Qk+FKDV6JX3nLAtXAHDJzYZMIh5RX2YumE7JTJ62J0qoSKD6A/cViPDvb7eaj
wz+kmXrUGor6LwBxWIJ5u3o4yB1NOi7+MdGYK0VZ9EuolZucI3AysUKdcslanZKx
7LNT4edL9JpnVSv5/k5hRIWnmVp3Rk8Tk8/8jEsbLUMQnQTBxVVoMc0xHWdNMiiO
F7PHU88rP7jzNPFQqR5PyVProFE3PEHoTLDS4keKWIto4VW+d1DCQjoi59S3Iq7c
TXXe5sSa4WB3PPz1qHHnoYCTHFmgaBv2ukhzrp3boNUWfy1qElA2aiVHTpnHygnl
eNTCG6evtXW8mvmFhUGHSG4IKV/ey+KeDX23OS2G7zFLB3eEYpyjCPRTGGm/stFe
JAvA+rU8Nxhf7lM9A9LemcChAr35rTfDwMG5AYW3f4xV93oDjBKStF3hDyN9JHmt
cy2GlucVX5uGq0DJ2vL79PcDpl4+IQx/CUkzy7lLG/0YaDgm7a2CTmucNxekfYx/
jtOCiIvmtCh5vNzXBVbhcDcbQtkVeCtw0Cd8M5eGo+gF4o6s4f/uOIyBStoAQi+Y
tbnzVtY2BRUzaC7bewfDumRxhzN3WaLZVHX1NATe/jpgXBAM6pL89YmN3GGCYZrn
HLpHZMRb5la1YbudkXmVMSskLEcQz0WDaVccvAVWGVToxWl5EGtUAV66G2WA9fzH
rc/G3zjMyTNlhOsHsrQaUB0U50Vszgc0zujfl9Pdj/7Yn5cz36jWmyqC2ikJjOFK
r2N5bBqjy1FqUVuxBwKMjfSsqCNyNW0lN94osr7/dNBo5EkTXEyJy50uW9Doq36T
6xaDq09EX1BFM2ELMMZPqUAZGpn4P4IpJ/IDp4AHyqRJXncduZA+jkwvKC+ie8YW
3Rblt7e3PdvsJ0UG6nX8I4VOkh0037+xO4dV6iTYqVZpAJil0AuUTLgq1E5WyR97
AYrrOJx+SKd52uQqnkwUFvEEO7Y33x7jUbK/WcES5dptAYgXKoKoQwZCZnRnzfen
wbgSoFStE0k0lUpcXFiX1EwL/FYSLB/Mysj1WDaptlCqJQa5z0QEzQrOUylPQ77S
OzW7DdBD0gWi11Dls6+G2HUy8UgVgvLJhqt6QKtSuVyuQpFZs6zmWiLe3fqRVxt0
dfAAh1f1TBXC9YS+v69R4dsf/K9AuTa/5yAG2Ri8s7Xcl+apWUtX74NfjNLEunJ1
6YwtpiWE73N60LoO/FpBPQk/Rdoa3Je0fx+xZbdfIhq5c53+GLivic7G0txSOi0W
A5aa9DRn2vt36FJZ3gZM54poiU127ype5W9m/A0ccI6Uy0t+3vVNThn8pLO5oU0k
WxEgyQTOdm1Y8g98Z3Q3qzdhjSobHBW0NapAZSqHyV2BRH6eO8GMEeMIHMe+yrjS
bdfxdMv5vsXtv4QGL8NQPySYx8tHYR+OMV9E3P2UYvMqJpsfvJix1hnOaSC1HDSJ
8OfjD6NwUCk60QCBwq38MQeWItRzztOH7gaMxAbV0TCKUrqpf+p/z8tGmDgzE6CC
/VfKR/4hGavGB/9RpZGkz1vqCleL4NYR5JlOLWG+NGfikgas9EJToBR0z8lE235S
skyLtB6erKvBkLG/0Occ4fqR1JFnmWS8rMG+t6wZ1JZwmaFW/Dr0uRTy3GI23wW2
MVei0KFMRM2p99rx1RQgCzzPLrt2Zabe5BaTuVH4Wq9E71R9m5nDiFd9UkFTJudK
H97ohLW8udR8BWBis5rJ4hZuNOvfeRCrv+HBzhtV+HbYWWXKWO8M04hYIVbSaewG
xhuyh4YyttssXrJt3wKCGzfJU8UKNg/T+tpyGbPBnPo1c0TLB1MJH+67IvBL2oXr
NLg+Isw1c+KTkX0fiCrF8Jsogt3qak9E8NCDmZM9i6fh676QT4L32gRtZuKOfILB
9/mrQCkU0mCtcdhbRM6RM856bl2URvtULPTxWqp1jquMa3WBCiKtAF2ymwE3S+EJ
WpWFvizVPVUehPiZbLYMOdlcVsOLlPF3Sq9JAWDWzQYqErAgRKzKqEAbYUIMCLUG
gpStQPM1M9boZPVEzmeO4Y5d2rYPgBOzPxMuZWnp8LI25ys3fZxro3qf39Mleixq
Z8Jcb8p6Coz1zb5QrrxWw/gmN6Vmarvj4UBIiu4efdrrxFrgIID17KaPqUzHERxm
xpkIGnaGPxkXUdBtgdlx3EXR5UR1OC2kuCnnYp9n9W2puOQaseqLkBIEyPyaXKCS
U+oqvbKPleocyVR3IM6MmuVFQu99KHVbbBXclGA1LLiC+ftdShfDIXnKitxJs6m5
OrcRO9tpkpQFgkVOhDGzkEY/LtQv/kqWPbMwb5Q/f7m6NA9tVzAXU5HndxIW3Gaw
T0QbB5Owyt0JMYmQLwdSMpo+XheJMR49HFNf6ruQ1X3JtUN0vBEZOb1w/IaTUgWK
jhaMV33S92rFmmP6ZYnueX2hesrPT0CZP7l+fArugx4aoF9N9DznGTnfOC+KJh9B
bDLyGzkbrrn1Fluvp1K4d00/MBP4wnHn357I9/3xZUsWinL4q4FLiLxzsJ2ql9BD
5RmuCapDKL68BkzEvO0ELnsxQv3QTKaf7v/bWp7gQhYq61aFYHJPItnCBP4xecYF
+pw3M2T6+2NyyIGJJ1aVFCU+dQvysZzzGstG4xeNoyPbgI75lVQrocDDTvxHFf5t
XNQR3uj17mTPSx9m+tAZjLW9XiUB8dLd+xGL4p9NdzbREGinVa4sRKDmHZaYcEYK
nnrr7pwzJ62TlphP3fZYCvypUAUSpdmRecf4pKD9wAWfJvcQhVlWahpBA6IggWuN
bk6eKZFffsc0Jr1nqNdpQv9WU7YEnuTof315JiL8AUpQEKwuK7Tk8niDdBEIakrY
AX3KKEJSMDd42hNYhJCA4qUACXgRreViiYOy8ZCvG+92e8YrAXo+8TpnAHACN0xp
qgcUpTyej5rtvrJrVkbfFtJp4DqxXlXaRf2TbDtTpnvIbzKL5EKlTExTy0XfPgDf
my+EadTNXCn5OlBG242D7QjdoBedawHCUdHTblQi9cVlFnQPkhTEZ+DU3/5f5lqu
FREscOLlyDiMeBqDrdNBYJbVdFzjBom7jEGQduIQ7jtdjUFuDX9wGqCGpSBQHUNo
+FXcwRH/oWFRdgAcFmV5tiD1Zrt28hJaiRa+jnf6Ut09Eu17B/sKOy5A0v5vIy2C
RltAXvFP/bBwPVGU5MoELbWgOK7zowWsSvCHdPKq40qRjs7h1InZx8oA/SlUvLkM
kU5OkmbM2xSA07zK3qsHvF3HAdrK7BxLYJJkx0lAESocctxqlLTmH5kjekLIsv9W
0iLk/21eKYRMdwKGEeHKj9F9rlsB0520fIAP8sQP8JigEcyE37Dm3QZ2iRx6Qlbn
u/y3075GneQkvIE06ySnBblvd1ParJS8L6fLMA3I/fISXw3fms4FgGO2UOv2DOCT
pFo5po6RXmskzSAicTBCGDE9Zy8XOcrJNt9PkbpEmRQrfoql/5JgIrNvYwZS3jmA
d1EnuYrwj3xkJyVR2TW7xd234V4l8aW1taUdH4f0CbG5txtUNHJeoqmTdBYpx6qk
IkGROUaEVGa9huUCiWUCcGEpvvqMq/l1Ekawu2FVBpsnypSVm6fKG9nkiT3ibVGU
BgjaTbJtFuatdTFuvG9aT5n8vW6smC3u5Dw0DH1O9PXKEqSqRBDvbeshxHCAVQxw
kzv+0b8Nmsu+BjnblDQIwWvd/gosA2k4y0AXbElQy+FydiBeP9+MXi5IafluOj7Z
lpMXgBZYm6Nft471ZSkzWQzCfS1c+wB/OOOKXtRFq5DIT8DKsE2HMTvufOHKsDfL
ZYTxkfsNoe8CFR0vYV/mYam4pzc8w5iqAWO3tBgiwV5DiPDOWAxmIAb2vAE+SbRI
Ep3ScSSSIaH2ZcPMDAXq7+E6nsbbXPoFR+u7CtRl8p2wi8TVyVVsL5E9yxmH1+nD
KA66kbiXLb/1MpwbBMAYZLwxQIl4G3Dabee/yRXD74U0J3iXmU5qVqFvs5F2ff7H
QXJABHmKJ94EtIC8XHHkxj2gNX88+DXjhMOfqPnd8+yoF+zMn44XTxudIUwWeUQN
8T/devs+M9JmXx0QZwCcrg4pdCyMXqikk/1sSwELYJbO0lXJDVqoh0R7eYvo6x87
AwHv0QkLC5E8MUxjk2aId3QBBwXU75O2bBXIUCvI9xv5tE+LhuT9+zv4IoON0i4n
wpd/j4vjlqlzIBwcr9sAZtMGUcYMqSTelEmufi3Dievb0ygo11wAFQdQDfKSq74D
HdKAHqTXm/HWylKzdER/iwX5u5kE2vo0H6gr6Dc0tpCYoteDvTOCigDUhTmZZHTi
7RnHQCS/qXh4FQybpFty/94Wld5c3X5xkFZLbLRaHo0iRHC1MbZdNK0tFpkgUMHg
+ijWJ/0VdnMTkB8K0EWibRotY2UVipW51YM2AUeBdBff1AqpOgJ5e+qQYaNbbBoE
F19b7HdNqF8FNE/Qtj/EMW7OkP+FHngnjN7M/3HZZdkfBaODpwHR9re6koHfu2bO
mQHmQaIAYwcjGq9j3DD/ZFY0JfH2Z4cE3mAoSXpQuAh+EA80SmsAR+UAv7FDhJ4x
c6Tj7wrV9cyx2QU0pvPSEp2vMa+CLNCFRZAG8sOMchCOnhTDSu+ZkecGpQyWWss6
vCiANZ6hrnZwiXpbpKM7T1Ab/VR1868rWxFrSRfv+DwOVNriLdGORVu7eY/8by6M
sVh53Fj7/6PAv4BgiOR77C6JY/fjqMKnsKsRvEaDci1dvcVq+XwRyHd2diVh/ob1
j4b7Hlr3rYYlb5V35wJYINLelPgXBwEFyLvSbHPn2om8q1DSD6MCQoFAR8DW5Nhv
q3j0rr7ac10Ml/Ireh32XDpbT8kSuaWa7JJM3nzg+Rkd0MfsgiU6Y5YvXogFuPQB
N7MXbkC7UX5pZIp9vqIofNLweUnCWSs1xjNFqSqySqg8oW3Q9bvZbwUMkkw2lATc
WQmHPkdJAMkLnINJlsk4jEvlSgymUXDum20kclOTYz0acq5/fLRweSfQrezqo4Vv
UUlrTARET90jQGy/MYXy1Ttq0qnGSq0ISLqEHuyZssTK/2m7DckjNAZ7kHgtQyxW
TP5fygf2BugmIjkaHEblFZyNcYyCuCV/qriWLxww+0GzEb7gPgPWQZzHsUvXsH9b
8stBW2Ay2xyAqXQBZrxJq19x8bWvj95nRMjXhWL9rSzVDwI8v625tnBCUsaHLdeq
dT03cnIX8BcHPJR+6EJBjsLV1fAgUgmSKJFLy2sHC9DC1vUesDGlzVexNbGYw0BB
A7Uk4ykzuKtViTqI2yWzMcWRYVOKd6248xYRFirffmRFKRNYTRiBhEwnj1h5GiOf
P2l0DJ7Emvl1BafIgW17dlP02vbiJ7nrGf1BNrefyhLNn3BMXCDmRersQhEqQVG8
HxRpHgOuf9qLUlI2sNgVTtigxVgj21HMtCqz8ouyVm6SbvhN2cg9py44bp0OZSLT
wYdgxbf8sQG/8dVqJzmAtJ95N8NB3r+Lg1tWGAzOeHmAjig8GYu4qTF6iJA9HH7t
0s/WqH1PPdwfRCQoWjyzi1d0gy+TZJTbhKGi3LeMzcVnlCkNjvBlXoV9hlXw399m
2eMnf/DKuBQMzCDXZBKmRhTvMXIEiV5YrCwfPgZC0JVZ2Fj7PRzLf4wqwd6rUdFR
x2FkjV4z6rx/11RU7Q1t76tVnZSk8nXamFK/S3yN6Juzo2yzndVGHcWP3vgBAQHT
d0CPDnkOHIpMSPjNniHJGJfabnOA2aGx7+CxpBfzei32pwSJ9a0TkFfKAZDe2iwC
YvlAMmWjw+QupLGUdURSIa4EkDUMIAyPCORMPoDovQ7CwJ0SWYwvT8gBpzl5nmaZ
Dm47m8KCiKfTm9hpX48V9KAZ6icfirbPz9cxRNzsDJ1UgCA+INMlUqqtnybUJtsT
FnvFASP4TDOlwZ7BL/MxGNM8uTVk9filZCEYw09BYQc2jwICNCAxNYY2TurceztN
gDwZa57PWab5+tZfuo7rdy+0IPNPaK9FiaCnZe+KN640QCSUZt7l89Bil3HHq1Em
+Hh+jrpOs9R1xiM9vT3cvLl2fvC0lXOKhZTjCSCGJff22QRazvXsHypya2XBqM4G
ajgKdkx17HQxQ3G4AOkfdjWrtukHSeYD54elu/voiJamHWieca5+0rrXnr8Eodbm
aQvfwtMY9HQXEmLs+gJeGIbFlVgD6bqqfGVHKqnSQWinph6PnM6GDdRTTBnRsrSp
5f1nMtc22D39hYnWRG94V0U1givD+cDUKoaVhXsBj0YaW0+HECJT7cn0QzNJplad
8lMgWZhvxtKCwcE0KKHOvDHokb2JCjjiVhqFPy/LYLbN/Dvx4yIpecpYIEHwWXpP
VcMrygomzhxF7QELqhOQ6RmSWg/FE+/fTENrv5q6Qu/oJKy2Sy41t/phSoSjQ4/H
+KHzcQA9pjSyzoKsW9sH+jgRjyhxs+WfTctwYxSHOWjcLSutqlI9JHKJXt1xyDEJ
dVc4eNZk8851CBXZ3eQB7poK5WYf1dPyWdKFPR4dqTVkZv0aRjDcDWAz+O9qC1SA
cC3s0pkZgT7ygI36Nelbg8wCi8ALXgn1RQFzA8ikh4dY7lDKUZiR6YMkjqBVDu7x
CBslXbX4Iy9KvKF7FuSMi4TjR4xseAfEt1s9EO8cdK81d04fsmdVpHG5ioTzrApc
qEz0q8FQlNpLDDtsY9jZW1uvIAxxOdbKIZkGDRu7az5JYJzlCAkKrXu/KJtZ2uKb
GREyo5geau/S6c7J2XokR4AXfqmKkIwnczcJAeuITuJnLoVePQcVZ4dssIYAB3y1
ugsbu+eOxHk4toLb70OuaXHI6G+ItsI/efoSgWaaVIgffxRe71LWvFDwkj/MZpzF
yXxELUQxvWHZr34zeFTTLABKT32FofE/cTP9xcy6SfILDWosFG3wbd5Cn1zKKUIa
ReJcuK27PkhZBzQQBAf2aLZFma1to87/UerLErelvlU00i5GiyfdWZ4MwRaKlavG
YnzyXTxmY1rlBchknz56MtdPgQTND8kJMUABqyu0weXtQ7ZaBPrvpnxJatQeo4PV
ZrlMgIzVW8RPvX+hGrinckF21a7JjpFyNjrQhVM17ZRGgIPDqd8TYw/TZBA31Fnr
BQy6jiERLbWwoBAqCCSMka2YVmtsLTv7+ggn1ClaTxAnNfm5l+15R9t8P0NXOREb
W/91KbXxgAikz9YG5EGHX66xf3VB/hiinkd3QIzxfMsaAG6S23DfY/EZgS7KVHBR
/lSvGhOpl9UH+DvtBFedaV/3Uxr8d/VMilY3WJ157PDBqAnJVw4AIOqk36878VKR
YwyA2CVBw/sD4OHvV/HoAXNh2NcPbch+NVYQXC1/yw5F5XPEgCPoY+lwQJeB9AN+
sQFtI4OZBZ7km7NfYdZlgYYO4xW1qwzn+1F7NNSKHsrYiLTvvE56EbmCU/ln72dg
hGndZML0gtkRlrE+fJlC/PLhSKVh20VPeRgjgFmx7mOembqO/Y3kS65Z9X3CqTCW
03tYopuH9O1xp/KKB8tJo/4fpJvXy3AErIIz9s0KqbpBIEEay7qt8sOUBPppwxDY
RgssoGrvQRbYPF9+LE15gwITjXf2F0Nly5o6ZavU1gHdJ/Y5PGmndJIPPl9sJPYT
6f3VNI6W+Bxy9OLhpy13QrgOw4fcBnXUZ9MhS5Xo6iE9TALaS9tDwQ5lrcgjOEvp
/ENely7fQ/nkGa4OVJdj3uE7TAxQIpt3RFQsIfxyl9Diflm6ClRDfy430JYzWGR/
wfCzlOVj2tK3o29a8NfWYY1UBghvcBvPWUwA3MTrJPfuIcAtS3M7InPWGchQzuC1
ypc/8cIhSiIW8+5hepFUm/4ZhWkgN2SSJDRIT4kgtOz8nSOSHJqGLFNgr0CGPkmp
ZkSPHF0Qyl+zRoQLiyXRt6W38JQdaVsZIZoZpIn7+xj9NU6H9yuFUvFT5Lf99EYr
dG8wSlB+Zodxxn6GUqQ3dNylwNx4SoKVU1u3rKoNNqTH3HW+u+zB/hqUF7YAoTXb
ZgkdS9u7wQKCg/huUwwuokWWgzBKKIUT8c3Wsy2D4g14kroDVAqP4tnFUgDlzxI5
Usc6PO575LmFjF4vYqROy10IqgylqkHVe7/hJmX99Q97WUx7UMGqtDzlWBmCE8qC
PJw6NRM2VX8VV2RUMJEtDe3egMS0MzyggB8zlG9G9gE/gsd1DP2qe16mZm5UyIY5
ErcecjWILqAYtgiTTWcfaoFJbnpzFmYzSWBh2oBknszgVUFiX6cMehCWLdgN1GwB
UTLGnVcatCn3wzsVMiqJctEi3b46J6BQN9T/lRP3ykRqTBCsKdGsFiX1NiEZ0it7
jdvHIMojvBD/cD9uSFB9KWHAF+n8hSt0YG62Xa1UqK4snSrW5HxL941M18VHFRPy
30FJiwwIBq9ekx9ri2NmcJPdeT4czKaGhyOdHGUwDtQcqvnoO74tubsFGInXdPvM
oNa8ovPwHzN3NM1h8pxRC8rHPWtrNi6/rid/IG+kvVhNi1nBtt8/KBrVs3Nxrb56
2Z5dvFvzhALE7TMQPXg/ejUG1ZyqZrzzV04efeT+VukdYS6b9+FDmdA/OBc72wbh
IGp9xL/hdDqYH5cTeJCTfbs9Z8lQq6xC/MWQNA0d/+fSBV4F30cwWv80TfFyxM5a
yT3OHEKDFvF040aS5ZK42fVuyR6TFS5JqSBlo7UbMLpAsE+8v1EFQ2Ukv0H5pg0Q
EhoKq76Gues+6VzZYcNQj8AI31rkBM5TFXuYmkI5O1T/Kbha2BvpDlVwP4tr5WHH
q6cfPsjWirl0X982KJ3U1BmlGACian6ISmHF25oL3kBuqNmk2L+PuQUaxIz3D7W4
3cWnrkzXrldST+X13uS8L6S9cdbhCY5Kx41taGOLTO5wZFUXDEbOFx09WCb+DpVW
8ldXKW1i5j3KhsApzjHJtIddbOl9JKz21jcsLDFzguwg64gC+4exWjni6Pbw48pw
0fZiJcQXIpPa8IRWGevtc4zPXsSqyCIZS3hZfXh0U91Y0exJJG+Utmk4P5Z2Yqfd
y/4kWRg/iGlMYA25f/SxLDAjlS7Xy10wECxX+hSBksKd5eO8qyyrOcRLjXKv3Nds
IOB1FyEvTMH8Qm8DBLTquRUaTf6Z0xfGT1RdVgbiMO4MjwklxCVw8rz72g7ewJq7
kvF2E1GWr6rgt36CfL06ZnznsY9vgykjgocRfmuXiRcKgNX8tSrNb3e7vE5H1J3+
DiYRoKjvR9qrcwzJwIAUzoT+al5HhGzGIANDBvspir6rZyR1jNbKF05rmJoWzR2R
R1ttlfT/g3W9tZlJ1QSPJZfz9dBDFIIIYWQXiBXsifi7mANYGnu4AU9HUTl9ntxP
56zrZptrXmrj3ApB0fIkKchx0v3mb93r2xBVdlFkw3Ft0rf7bZcryjxK6JoII1tg
OQWi2o7euDamWLao/cbZXbnJH/gkXNhVMRrXZ6+GJ9NC8/koIRgA6+wAh1QnjMpg
esetQPnQ2mVUoNFUE//PLrbSF27KpU38MGGC1eInlN1kakyoF+w8kgXGkJe1+MxL
WpaGZ0sFA1jBvdTYLkQg5uYTrDSIaSr5EjH7NJHR4xXHgdP+pnUfpBNCcQqupESW
Psr2QNcCuCtfTOttkZIrEy9K7GPi9zn17hunZg4ezEuKNrPMoC9SouFTkP07UnQ/
2Qj4xdq1eYDh59U10LngIm0NMZ3m3IMPSI+9ngKN0WIG0pQiZ1qNoCU8OJyFnazF
8D3uJNC92q/WnhOicmzr5DQDyqmvqw0J8Qd9z/OQrR0jZ5UD1TWG1SdjQdev7zno
lZj/DndT2jQ0cfj/bnM4T5TImWJZhoY5uYwthBSePamK3c7a4zPGcpDkB8YWZLlu
dQibJlcRJ/j3PStcTcwVroFXgTZaZP7a7pKd11l3yeSN4wRt3JWftoAR5UDvcKBj
vdmBKF2qP5DjeiEa0NHhRnvu6tCwAENACrLUBW8SNEBwFC1F3EMzr8EXETOXF32H
fgnnl0RmWNU5BDCscvKbeiEDTOEjQqQcjWz6RfKOwJXp24tIAaBtTDa+bRLsdXUE
gqLEw62DuNitYtDUGC0usS9S6MmyKNNXig9tm7kgrQ0vjse00rjYYpLcLek384Du
NH621cCqnMNJ6ff65fpIWseHCsVW0ByPyM48UNpPf5skpph3KL2zXL2V/eSkFugA
1KaZv55IdGErN5ccHONRYE+ymo/v7y2aIP1wArpSALzynnIbKYzrvc7yd6cjucrj
1ggm2Fh/ktaoA9WvivXF8LU4feuVWY9dVDwD5/8AcoMjgwsOLW+Po+e4My63IqRa
i6GBMhvXHXlkd3864uaffp8f3TPU8rCQzei9f7xMZeDSALZ4XrkUyY6CpfHcQKC6
1hTX+2l1IkVLLknzfDb0UHpnLK7JXLp2bsZ4iTyHGsmuvBnb5iD/rQ4rZgVjJo4n
njvLrXp7/HYFR+vcxn75kiEEWXR55+Octn/XZv/1cFPR8Tlyao+3O9z6U2u1H1IL
UqFm0Q/jACowhoUihuAxwloB6ILwGa4ig6J36kJWOWcjMd9lX3QdaKFdG6BU6B3t
Ktb0xeYvBCJU32gv4+wZmBkgmvThc5AmJ9+iDpV8l08FPs4wshRGw8a0A3ReExyd
4QX10SyilOCPS/XS/HW5ulMzohPbmTa/vCeVL7fRZXj1Zls4w9iNVXQaYjAtxr7X
AirTiA3oQFfPuy5+PYmlgmLtonnpM/LNEzoRpibVZhVv1JeIYg3R2D7wjFeYVL7o
HDxOzpll1zVmnW7/Oq801ESqPklyabrMr3GJ4V/z4rzWLlovbIBDc0gNmvmpXWiD
5DUp28/i7tY6tpTt4cltF9i0Ey9FaPg9b7q8jioQEBc2vRJd7lCWcaOS6Ht2AJ0a
DqaMELDGiJjiHx1rT7htwHiekoAGYzdGWJPRaEysXgzcaSvq9PSyjk+IrSftPT9z
Tqchxq9DvtnFjltFX3X60JA86Ghw2RYDjwI1KI1FKgBK5j4//uAXia1PJCfAh2qL
yrOAILrlv+hXDIgXkwb0CBfRpln/x+GDJQcN3ANJAR/vjw9Sa2CB0Qo098QSrfbP
aygwTcSJAhN/4czP4L5LJBx2vHCybZ4vrIUan1tGPnq5vNlAeq2U8rbls1xx3IqM
HJFnCthhQ/cm8+2hzaU5+zsle6c6Bdl0r7Swd37246Ee42KaXpQuIseA8lJRgebh
CukbQpcIBmg1mPxmvE9CV5Jz+c4S4RaAAeffuvm8ZafgrFX6Iz23ogIkdBh75rNY
xoCjxPO0ecBoOM2KdzFOnoQjNFP0txTtsUDBwQgWM8d69Vc3Vz/5y1rSLbOL6PMR
zW/77M0Ks5IbGK4PdQ6Yzzhwwg8/IpPCnq1BxtCPcPbfPoq755VreRczqfirMR9r
XyJpIi6LJmaYLsvM8jIBqNKJ6j+1WeHCwg/4JV11JohN9u5/+6mZFdYmwWcIoAlt
32oTQaU+fn3E3eRaEKk9OKlGYKfmb+Zva8vx6Q/avfczwY9gcEuE43pgRXjaxsMj
GPpsLSgEwobFmx3eOpirl2X2M/F7ChfKwdsRc3ydwIrT0IHHHrD46uhtVeCWLh3d
NO9xIGlGF6Sd9CXuNYjVd6KtLh8iZ4Gt+IdOOxYwoFrvRqRJpFle5NBNBklD5Z0k
eywM9t16WdWjyJsryYwQPtasOcB4aIvbzbNwutl22YZaTG7T/62n54oZ1QeM9/wA
lVS82XFLm1ujjzYQJIjQQJB2eYw0EUj81jk8a1Dgfcwn/52T0TS0pcgjDufBr35B
b0BYIjsW7WS2z3UmMKrDS8HR8aTN43varAqlLTmQ19pMnQZyZLb0KfJ7ZwDNrS8T
+aaKzYEzmqzHMdBkqS5KzPd5rqbJSmlmDz4j2j5BgLhQv7YlLloKF9A62jgOH4jY
TKP+0E/FtAK135ECVuqa7EnCNYA48lztX8b0jZHSGgE83yh6Y4NAs8CzUDPYhdlt
o4pbJnbepxmbK4WG34L7BGJXzBF5JCVpvvv9UzJJ23pXi9x+T0EPm390df3Ajatv
zPwLgvgce9358mloPoBQioNQPgn+vHQbdaD66jtUG02fJpEJPZAGgOFHVi8+7THI
yaTpewGdsmjHp+rIYZsWDcWn90lvFlOWdzrxRzTZlh3+pPYqsc9R6Z6fisF1BrpL
saq/Ssa1BYuPIK2bFniSWdXlAFWHoyg/sTzGf0iH8dp6xne6GjIka2cm05791lx2
5r25PXzCcSKnMDeivhCLDzqfkspJWjUiBaHS95IZ/mmAWReGHksoGdMQ9yW7QcIJ
N0aJQNYWZlKc60uXRRb9y4XS7ZFSuNSFRJKj4kT73TDxEAR2Lqu44VjKz8coIdLL
1s9+7WiK+Zcd5Nks1gaNFIuP8MnQ085LJ4GIXlhdWPmrceE0LOgUa3gpcZSRVKgK
MiMY0Ezqbni/xig82DQ4AXctIuyAtvMvlW7Z4nX05oAY/0zipeB+KIsqEfFuTTCh
N3tzCjtVQb+hTvkwll85742aqxGLVFigzV2lavINQRkDiL5vKZQMIIQuvVZ3gbuj
HK0IN0nWEf+tAlE2LAOhRELyOLpdXN+gHcpq0EY3Vlq2R5XhzrmGHsF6AZMtM7br
6sDK3pBqlBg9PAIMAWS7XpxmdcQOJJro8y1H1kV+iHFvGmyd7ZabSWIWvHtnaITC
Ny16rj32EZykCt/v9DM3vOs+yGwdgjxMcaLcwwNn2kcOgwnfPA4xeQJ0E76WKEK1
Fr/kbgwwb2Cv++3bWLctiRL3K/iNubC49wMNRmqCuRay4YyJ7ezhxSWFHhLtbPzR
ZeJl4TAa7s6uERPBLrJWidHy/TKZ2mx+EPoihexKdsA/PeobmZ9TYopjIxtXQNqZ
JKxzaUCaWpYIuIxcxEoF4qiZ8rvHkHeB4b465IgTtkJofIAcdguPq8GVcOlvitjB
Gje5ecFWhhWGwnOSOpzJKhmws62GxQW8ATIZpbkzoeZo9GnGxZeSLYWC4f97RsJW
gx/wiCVgb/L1zt8MztZBZ2F9mwzpuhS92bzQEsryrIyxf7n5FuY1sOf9q5AkfUhe
9kKZTycLpJEiiOXEgqZfeFArqXuJsnKFkpLTRGm9Bx8N7NXh+85vmaXPqNIWNtMr
r3wj+9JiUQhSE9Aj7E3cEowUism122NrLFej23mh+QK7oqZLuZOvirkBTqp1nbzH
FJKYGmLDFPCaO4b41z0j1NMX1H9xbVztCOMGn7eLgqp3woAor26RFkL00U0/slKl
BF3YmXTrhaSHSAu7z1h0G7phP021n8L8zJB1tXhZQM87HEfpXx0dh+OyY5pcMCdT
GjhlNSOoD0s4EVZ1WI5tWMDQdFj+k/Q5+Cfc5owNOOXNNooQCDAYeKqPZRFoG/Ds
Xr8nYfXuGol6KE10yxKBGCDZ1YMFuw2n7cKWWwCEfp+mqJgBHOKWn6BKhfyiwa5N
f979K1GOKUJOE+L62ep2BTLiw12G2Cmo09y3ckC4DjNT33uODQPS9jDD07lrOdH8
il/j66KzK7sHz2Ui66X8pOQ4EBp7Q/kSS6EhSsp3IZaZBEQs/pgWSr3G1Nt3Y1gZ
CVuBgSsWKn8s08w2kRpmSqs95b0HLgFlYlPT1hCqLBVh65SxMUBuQe2Hcv/5r5wD
3Tj1p2/JoajYNQeWVa5pwWWoCgW8aJHhldJ9Wbxyv+I+H/X+ExJQkt+j8R1SJzGZ
kYzGlBK7cBUaXgHq8SkOhlKdpZ2ypGZr/DxoXiKsmB8JcxTDZxmNhCL5ZLc2fKSR
UWkWEuUvZxkZVEnLpt+YRTE20LEc9y+yt0moGa/31nT6dRTUnnwjGOSQLCDg+BxO
jKqImMWin/iuNu/8M5Wn45mh7kgF6klwOciMbYlGMl4q/g+enPDJ5y41AfwDH1Dt
hAAUVopljYjAA2adXKF/4kLc4opjCL/lsE49/709m12vguIAkkYIKN2rAMyiv4TV
+ik5MZ9I+hiJ57tGuCaI7fnLc1iJX5DwRrbg98EGyJp8bk8mK31OMnhCfxPRvK6n
rwzUTDjhpAsWuFgw0r2vTaPD57JEK5tMVqOlVXlzfIb5mSa0NXqKVN4cpde7OKbi
LQgKIAZaf5eKsc2B9aGyuNttF/az2KGMGIEAhnMBINeMZfv3tueQyK87kSRehL62
lV2+guYpeC0wZahkUxrFtFv31MJEi13hOmfxWSl2W+CiwGRCkSi/S31xQ4EDHwJa
daCrl9i6SgUOXjC3bFYQJ+pcZKfvrk7xDCx7zaqpNFt+NLMoNlUrw2pZuFd+zOa4
19g4cuf6fLYVKfgRCkyw0OhoQCM7zFZLARsbh0cOpHSMqpzKPQVluqT1i84WZYTf
MrS3bYX+l49LAV7n5q+FA7K9fE2J2jAc1qrvhaqnzMc25Wq5eUY1WYSYhbogAttO
jw8VhFqClYGyYr9kCWJyGYQgX9tTP4MOtvzG8Kisa1aHHuwbvu+KOsVCsvs/ZcV+
lg8jhLeMeuuacpfa945gjuBkeAU/xFWVdWbT1iDqtDsPU7az7OVeSmybJV8Bs5b4
0TQ/ura79sHqfTkqeHAVJT6SzSm9oi0Q0/m/LZIZrzuE+VEpJZrbQDfhQFAY1RF7
dL1LBQi64F0Gp+Do6GepROKZtxDWA20Yty6zK79k0GUqYrrBzIXJCEceN8Ea2fps
uwK9NWZv/wn4hJgQ0Tncfv4CM0YZfOL6fWu74crqUHUtn6wTcvTwWiqgKrXkls6T
B6LX456yhovYIqyvSm5jlqcf8ce/U0Mg0ddEoqX0b3HWz1KlygVlZzXmSuoqk6n9
E4XFPa8ssbwnrJcRB7KsO0S+qoQa3Tue+rmGDgRSO7/4YeXFBL7hnkmiMil9cqOZ
YentpzgqZUnWpW5SKsD/aMNwripjDTf9xa9PVPSKwU8IMiq+/ewMXJ1B2Z+JXEgt
3huSwFA+LST0INXBIHIKc7XWL7LO2fkfq2MAiXjs/BBqwHT35vbk2PX82EMR1tui
Ul3cVspWXFB3GnA1KHo/cy8uKdWdQ6vN54yWmSjCUkcdTPBkmsOlaW8PethQ8bjk
lR7PnDpaBEDSOprqbqW/gf6SSuBUun4v2MaaJRUu8iybDe8MC/rM8SjoOUQYmDjM
2U/InZzy801qK8YgpKuciN9fhNbP7LgJbpOb/+bMLWbdBRN+HSTUZmGQ4Lh75Fw/
1Jqurpj9DftteGpPK8O9/faGYTcXiHYsAaS0hSAXpgg5cagWTJOOmSPII818pgKj
EYzSZWmUMUsokV7+lx1/waprcaVSvAHhRMcLL8rCE9KLJ6U6gj7FTaWeifP/WO6F
gjgY1IfhwcJXOXZeoaT/7tyYXtmM3b/3eTUdl3Uzm7qEIxg0zrpW1xgEM4mnxJgr
Ajhjcxi8jIIRTJ/IxvyRZ+SKpXN85fOs7+cXQkeZL7qX++X52KohMMbyWj/qxvMQ
s5Tjw5J1Y5xCXD4tdwh6qS/URzAQi7RCPHYeAmKTPQLuELDa9+Hvaimles0yWMBF
uw1mwTKbD65giAPMJXBmURa/8DRCbpVbcRhimMEP5FZaMloi0/v+XdT9a+/s+99E
XFucKHvvxxH95pEZTOHWlXLj4TlVRySCltfmRBnrgjk3bRQk82CTaGcB0yh7AwSp
AlEA7fK+9uo/qb1FBjTXcVwV4iCyKrfnqtLOnMuRfNJSqNmbTFDyNFBcbWw4Zn6L
gBnSIbV9qcYDlwimv5dfHih7oXiPZwLIRiJgRxQ8mJ7MxlIfzzmtNeArbJYBF/MH
C7S/e1geKlDYF5dpGGdUyAttsl44XxAcK4eeU1L8B3qzGthVayKLiKsSkHvP+SUS
eudlFdegEIdBTwV5JdsB1Kr0Tcr49mYZPU2YejOQjEWQxfH3fVHuB/s1FIyzwya+
NUfzDzTNv8SmkC9WG51Kd67rUiEwhIUR2tFh2MK8FeplyW44PsmWDamWeOdrmNEa
vY9gkWrC7ZkI2nIasMHHU14UF0c3qIXH1f/PeNZi2YWEm31CFa/jtguGt2grtc8F
iaxLlUSjQeFkp6Zzkh5mR7aPCwFsRbTKZ197c+RAO+ixmiIc+d+09xjBMUrgJICx
OO79dxoIwbzhJ+dehsaU1L+jVB4/DFw+F2R8oB3GneEm31IGra30TwNAEnKFZrdF
PRiwLac4GBKv7phCUJ7NPZGvdF5kJFQkUz9iQHR+3gesi81jDWZRkZAm9yudbTar
wjl8L8PQrqHDcpuRuYmk1PRotZxCmHCU6zO30E+bP6WopMHHinbmwmPF7w734KHp
h7tykjN8fcXjA8LEHd+GsAW6tRZgKYEQQv3y8fNw7wavAdl5v8NQltewW5GDKEH0
DU4OIqwv7cZp9rdVrXc+W4CNxCIoKn08uS8wALsCemp612gzFwmCK+FJ5ArtElSk
toic3H/6vsCGHzdakOuiG9e1Mma6g9ioEozCpIiNzERNT9wK+apQDD/YvYcC6FIW
vh3s6oC4AHHX00wF3k6rWoap2pr5fVkCaQfWvRsAMx9w24s9pUZOSPjzrWkVvFQT
BjPpu0powt8e4eDq7SmF6jUYiHyfiBhj3Ki9fsF3t061KvUnEgIt1yVRZx+pjTy8
u6M2f08beCJ8iz36LHNwik/waxgCWRiIQDmrbjn8MIDrOvJCA2mrS33zX3+V1j1U
/GrthrVA05qV3lybrMsbKP3wjgyT732pD8yH6P85a2mP3/hl9jghiTsa2OUYfh3J
pXhTOKFPTdadUW0ojCPo7hR5NPquTI7iMfDFYSfl8FYXIskH+oyGWcrRmgBp67TK
IcU28sIjvYpILR7Xvukb2gckS/R1AhV2G8xli2Ysa1BO7BH0L6QKcXHmfaGZxcZJ
t0e+xwZhLuLWmgKHKw2RRU2l0oJrgHVMZw8+rJ8IRJvUI07gRLNLYl57P3689j5P
4XN+bivkWPr52YIcsZjECRWClfY+skVug+229Vuof84aQAgHF2uwcpKZ/fzqgBHE
jFlQuN/z/l9/3W2Wp6dc+dcDJqt3e+dnL6wThujZ6ITgbxSPkZErG9CL6U5YEkPt
b6pcOcgS7SJtBC4RZP/V4W+i+8SK7jRwDqtdp+Oxvsqj7l2r/8h+Y5etcS3xX3mX
W90UgLLwugYrbgZjQKl99yalelQeHq51NaXCQ8NBgU8UsG68KsrpFoRt/CizqUnI
MafqJ3Eq03Q8bGBbI/YokiURZynIs8VUf1gyjV00OA8DPSZJDZ8fWdIVctZut1ht
dbvHqlEWSBaRst0/mFurlqfWlUgdnWYVRY76XCnGZT7oWMLOt/G7z5Zza+HgydV5
c1zW9sMivMJ7yf4p5zHMEz6zLUdjf1DSuo9AcGTTUnqpzZznRTSQ3qEcWOhrktlJ
Pw8vM8MjU6raX5+7hP5R46TUZOnhvrOreZupzA/tEirAuvoxw0BN+IGzPCqu5ngk
NffV9S7fN1780PaHVGOm8nLslcBuQ+HR7FQWbqnrdaZ42SojdhCjFFfdSwHRE9j8
XopdkbPc8xtezdQ5LwZqRLltoLafjMz2BgTYJX5YFVsTtB6R7dhe17e7fe1jl4DY
clFFjaF37zRzAJb5aQczujAqqlPKIW9MfmxlNqNIXoKLK3tck79x7OR0cB7NpmVr
XLDMrDnTwm0FIY9SJsCj1evBcw5JRe9xekdwFpefZ6OyqMWFspeDAjD2yrpj4YgV
qRMu61/wsiszjR+x4Qw/MwESSJ1yrg5FUAJdXg8hsWEHBQIw40fCo4te5FFAgcw7
qJfzJFQZvbVqahHZxDYduOQVAkwQMGNz0txa9zF5HRcFqyGIptsMiGwhrmya5OFm
VcsFSekckEvcMSa0LxT7LAd1JgkRsBsvvpm3sLrAZ4YZCeCFhBUhnRuG2zE9V2AR
eMjmmc7l9XAgJUtjGsE2SinzdiiOMVeTlj4ijD8s8W9lMo5q5O7e3nyNiK2iGL06
8vIg3dh0zfzpLktkP2KK4d3up+rdEg+u1L+mhFC6y9anU7OUNzRW/qvFPp+Dijqz
GUslpWNY64f01tidQD9M/+iRc96rKAmXPqJhG0WvlrknPm0Kme7aA9/SEJfAuOzH
u4wWy3g3ffMoR/Y7NqWRbupPhXZTvGxHSWaQD4XRJc/sbcNwH2vxqPtbjab3kHxC
R/FzefYHb86b64vkCefpLAAwyTXGMyVRC7OcAp8E8YqVdYPEMJoDf8ksj/bRC4rL
/Me/wZneTKEPBNtmMXIPXTeYAtKrOg6tTW6kzaEIne1s5eSsQ/iQDbOznrfwPUfC
dHCCQCpw9Df/URBZAI4arr4cbFaAZumVs5bqo02pW8QSZLXSRs2dQ7wURvvafNbF
Wx1oEOpuQNmmhxDnKGqTK1sv2ZVO8+8pgJMkpaBmBVW6ckvcW3pHxLReftPVfCa0
CpEVQZ0TdIRED9VPd9TIr7YnGVxYiCudljB6HRcG+7btdH9hAkWGcitz0sEBtr55
BHS+iwxKIRx8FDbgLjBN4MHkvQk2KTEKjWYfQGFL+zfqwfSdtL33hdDO2NCB/O+1
LTtcDsV6fi9DxMT4U/dYyFZFlprzgCKHHr1CQU40wREGhzkSfZWXjqs2St18gABO
sylCDcAZaTYT0yWeb3t/65ZD7EVLerpqRYxDv8oOwCToZqN+QInTSpPkEwyEvSWQ
7Y61DkxXeLWuknqvJI9PV4YPaAM1N2jzEhtwBZLtq9IHQRclxSLlHDJxDIyfIkGp
EDp0H/3v0U2aG3VIdX0yxt/yGXfJSiwiV9iGmyK32GuTaiJ8mvRzfPxbKk9gNbXF
IIhFbH4CO/E+3xYmZcmZ/XEQbmUcrBiy90aKnu5L6bukVZrqh6vwZF5iy+7YY1rk
8tHjbqdpIDp17Hjnm9GAkH52H/S6pw/2xEMqMZQpgtq6Wl1PnOr+6WkuT/igZyx4
1xqdp+UzNDOD1tK+X1PNvAZXWwNgBuZjaw+Gz3aHpa1UQyJ149eB7GHAty6W40c1
Iy43ZvhjffPVRawSbIeCfwOnJilHhtusacErDhHS93Y90OSU6MeWt8taQzGaJbL1
cl3jEfyPBxw2ilkehUpaaiaQg9RySgvLhC4kvOha0cNFqnAhuUWGUdeN4XVv6rmL
McFJ3sVPg3WKN3WCqKDoAdGKX9rwAId0L305pFT5jS7yfPjL7uwJ8fmXv0LvSgAz
4urn+wkLoZRCzoNUKgAkqzyAKsnZWODiOQRnpCDMoNdZn+XL8xKwVjePyVne40Eu
LFu2PRLg6Gs4jqA6Dul5fNw4QsDkFL6uTs5DBfhco7q3LXVsHIgMzK3i4OoWlMES
7q+bRZD4fMPgKXS+XUtsVZT1w+g4FJnlfdieXmhheYw7AiLrPi+2svNdYG+NMqqx
GIFI1OztPK8cMy55j6D/TDkIAhsxUvo7WgxIi8tPOUqd+mx3EcghNV+yU9EInOef
WaXLWYLwRXtXbwr+IomQahjrthut7wzRMOPr4yTew5lYDwLnlPVfZFHkDsCQZt/Y
TpshzRXlkIJvd9BdkEe/A84BOTFbjbS7+ammYFYzNF5LSbbPbSgnFxMlWc+oq5ts
9j59ZisuvZ/KKF50oF+tG4Ks54uB6mvWwSV0LnT/ijb/Mw+P+8vfNksbxZ66+vN+
5niw7beGPejShNsUzrz2fW3vMVIDoe/QYOMNMskpssUHkQYJg8vjTKTNwEZh5Kq0
iFVfOMBcjS1wYthutB2EtFupJVubd73ZqgjvylvqXpIMfwt7vvVqhHWb0rW6mkFG
iiwzXIuC+/MEPiOwk0vJzfT+h6qw9JsXx0K38JRzBKdro4yLi0LSU2/Oz+W8cexZ
lTsLBll/v9LywAeN2LTwCKGFu5K+ZYouvTG0DzJvIwNmg0T3KE5YLvWyVPBSRMNM
n8oNOO/TVB0X+zMcTddY+mPFQqE+HHyssodWHmaQHhuKSlEZGvb53nHnyev8WtTB
hnLdQitVTgXGejJ10khkT54m4l8hHbsn+YSYCm8I3NRs5ZR5nYg+jlNpsoQe4vDB
RfbybnVtDgkC89j/cTucNgIdSi5b2XYy8hMRhD/BmPm/pxWrywCAZGEyxWntRvxw
JC2/om0tBbvFu4eaHohszjDNfHR+XHS2Bd6V98IF9z4JFmhIr4DqUrR1AZSCUWrB
jhnoAA5l16LADzoiIuDmc1FrQB3+lEul+f//N40xpDl7TPeFh7YiYDpsRdXwoxCf
55shLHC+FuZUs8Gh76tXW6o4hGAsJmmUQ8HHd8Yz4ZDxKymbWyVXbDvqkhmsWZaY
SjbdW6p5GRtIEMlL58no3s03Tg5kCAO8rcrt67nwulc2D/a/Bn5CtYvMFDGeX6t0
B0tnAB64eAKqwfQ/B0IuGo21N8Q83zLsTNHuIeXCoNDXX62rycG6o2Pc8gelIGVR
TgQXQ42UsNB2epzHbyAjy9UCjm9Ezq0tilu5slGyOGX8T2Ap5udQw/lz2lbE7EZr
yRihx6fV2LBl0ccSw1vmMY6M7dfUt42iea7Me3Bnwrsi8bprcLvrBDN3YjPnU0dx
GImNsrKBWU4dytzoWMvtKG59oECWGZ2OPpgCMf4w0D56c6aIqxzH/XpEuWEdPc2s
rTXRpiD3nhgqTihuhpyJlCzE8EBYVhXqxnyH1mPD0NifPM65q9/bY4KOHFydfRV4
UFetREj3RUFv5/y+cHBBfzuqwKXJna1KT/kl+2WE3Kvqi630grvSd4T83CXgNqqQ
Sw2K8alYIIsicl8+W7c+HRpCQd8O7ES4EDh8EZQ1eDIjRSMhsJ+6nFHtOR3yNw8x
1976ZlVTWRIFsNNObpEB9PO0GI2ZEjKIi++PlMB8xuTqrA9+wNwdqhdsVJHATfTw
3yEJsRYKjHz/tJwfNhsz0B7pet76NZtcasXEElFJF+V70COEibWQVFdkYsVdv2s5
zhOA00uNFpfnrjn8Zepimejtrp6/wpSxJ+Dk/5HMoX/r68UQrTnjZcVH95JfQpnX
JPkxV+zQVpDjdSq38XBDeJmrMJXBc5qonwguXfrsYVJbL3sKXyYcy2iNE6vp/Orv
92wBd0bORktbD4dgnfjLC/CNRpMZvFe3pbuzjdQqxsKJUee3TDDFILvta/ff609I
aMhuN1lscFpaI0J7wkJMlIiVCdZhlSwBE119Uyx11Q6QEOhINPLlJWxt5dGAeDCl
HcGxoEv933on3Tw1zw/gjkNMhq9Y/BrFp20owK5jQ9ug0ljt0hTpivd5jZeAsjF+
Ede2n94BGHkGxy+3jESBJPbHB/7XV8GXt19pYnxmZ8SGmC+cKbUAonubPzVKHz5+
pFILU5B72iU+1iMBAj27mv+o99Rs5+9zxV7Pz38zbTNZITfRmRpmc5kZu5iWN+Kt
9c7C16diN3e4DBz+fQHu1RpLg/6mIHiyqLJnva1VRHnjK+ooXZU9Tly9Aws2XNoY
x2NMMxYtv7AeuES/wjNqtYA5SGJS5zyLOvaAic9m850iXzqJcdqiJagKaaPf9/dN
jPo5vgvhQUVoBU/LFP2/Exjp72Rlobfnjc0Zi76oHXPcfXo5npBdR0mjTqtHXgFn
zMnJFVWYPGSwGNVvwVk84C7+UOfiGkECSQs3l7EUyEPNe5AYTn1OS4XFV0AVVpPl
00xLNrBFZ05eMgrzcGlIQzgIB0BCuI6S/wMljCH0MC5twm4r3YiOfXYaBh53yIKT
75liOKhVmG7XrNcATv1Zvufm0JO1sxFilH9q2HiryhyXml1X43F4g9vtqq3v7JQr
/It6ATUjVZvqz1kn4jMhwhFSec8EyOOQ48Q5F+1pp/H3jgXRZ3gL4jSNx5zmrOj8
A9CrLM4HbIDfEUDCneFqvhM6keE7L/wIwaWv9WavNL9EVT8JhuRboLqLbDGkNwjK
pxYUmQSHpqHjTDNG6U4Am0HKKtuOfUG8OSnz4hLTLdwF6W0dq2CxjSl+SmEbIsU5
JdOdmgwhkzDfqGImcxygcvMpTmhFtIkyDsztEIRzi2oXZ0XkWKltP09/f7ZyUE/6
4d2qbXYEI0kC3fB5WLeVmBoVTd8L8RIiyoAKvP+TxtpBE86yxcLuzZs+RWdkbjPL
v1XmxVWrjZzb4P8K6r9UHq9UYqeA0/TdqPiT2evjZ+oj+t42x8cCASnXd/5TN+nu
B3c9lBn7yqnqAWoGsTj/THLfhingA7R8XCFEjLig//PFFhA1tJA0Rt0xRZau+F+A
U7uVvokOi6QSuiNI8i3YY3PjNtTSsJ8OND9QVFwyzsGnM79AXowW0fQSSVm5jpXp
lCdG/yL4V7iLuLMTSvaTnxWHSMF4iqguppHWCJ8mUOdcT+q7IY7i/x7WgXfPwD/+
GRpuzHZzn7SkRYatSb7MmVoMPzsU+rP3c4kSm93W3HglfqsUhOhzaxa6zoXyh0ch
NY6juTRGkMdUX8cmCn4z7z1DPBYY87hGwLqUWB3cvjWTJC5Dm1r1m73t7vCYj9gE
auYB4i08WllpOhJvzLUmag/aUPH7FyvCY9dlNX1DE3VSgIAtetpT/1xsNK/pRPzt
RHgGCOrX9D6p60u9N36uM1mGDMUFliL8mQacvIFdqNxtq8jFz/XSB+7ut0aWMrhb
J39ztG+x0sP+pviaLajMO9RZOwuK6UbeHDf09XurwpmJwO7Lh1AqwQiBNqVmWv2e
oScfOO2nsk2YCPzEMyN8BSgB3so+IUYIIKQD7sst9I8nKcwSj0UBdf5JYIp69KuO
jvRRp8zHUm7hyxpUOU065d3aHOxvZpcJ8gt9MxhfSa2xfWScnroIBSQPwjlVnywV
kR/T6TpoAhAUk+7BgnwTNXixU1TlP6iobpxfKf9pa0v/GeH6Cee3axMvJbq4uL/Y
fbIu/4fqYI7YnWX3M42lqtp0jrz7sgDaEd1g0h9LT77S0aal+cQOIYo3jAPyG/u+
umBG6OCp/Ncbo3TtVrc7eCSluCXj2JaLfzM5Qvr2paKRnL6n+4okX88yjv8bDnZd
piSup0nhbVcLWgoPPF+rViwKBZsW14GEVGOu7Zoq032fLHhdMxwBzQ6sd/kcO2iI
pTxvTQG7bW4GLoOBbT2AHVxEc4CFk2czbtQoY5RH9RzJ40b0s2HZc0Y/q3dMlMUu
+YiJ7GNl9yp0N/jr1uIPrPVKBTTCIoTaNOps7ES7UrJPPvYJr+AILkkC33HNclv/
mtsOfe6QThLWb8CPGeZBBcaAZtbby1Kazk1+Hm8qvHeqLUSM4StKzPPnhgbKqEbb
Kr/51A/Sv2QzBXHgji7yKRRDBwjtod5OH2R4RpfPXzWvYuUDND1cgopS+NmdMtlv
4U4VWZuutunfw4R+AFrBhmtNK0Sn9kUbfKI1vx6GAE2p4ez6MnfwT87Mqx6wD34H
rCTdC4//ey5cdqHWx19I06j36yKgIhsoMki11VvIEXNnWVQ5nll2sEm6aUwe3mtV
NGsG8/Qy7EdPFU8Uz19I05kDooDtUQDux/S/Y/IgMECmWC66httKeR9hinvB07OS
WrynRRhWDFGR9h+Wiaz4EASafSPgz3U9SJj5VeRa/z7VopzxDRtp+wOEjHAOU31s
vXDCevCIJf4O6iRiGjYjF8fu/iavezwOWmssXyKW9z9B2Qs1MQZoDZR/mpTJhPH6
0iV6FxpgLtv/iCEemp8r17LUeauEvoz2eVOsFoTO9K6Sp9vhDi0Pc8FWdr674hNo
Psf43MBjVTb5Mk1zXfsAsbfqI3MONudZIhiD5oehqOzkgpOfMXL4piaNsRaLuNZB
11aBTyWoNnlMXavb0mE4kWZkAcp3+j8vuXY8FNN11nfvo8EqtVf+L0aTDhC9HGVG
ENsiTA/XNQxJUyyU6qC2OJpxfBHkUWi038AafgEynb4kh25m4qheCygGsJSfQKFt
pOUx6cyOTb+J+DmotWJFFBF2/iB3226H/2+IhkG2cCcJpn/sZ+U+m5Gda548bKHC
xTiEYBesCKS9HEW1j7emLKY0p9u7PBlT9PUhzRt9n95t5PmxYe0o7AXpyP9BYKaT
ZIFpf5oWXAEcNNGodfU4hym0SZ+MsunIl5Ak9cqlkNAg908kf5VtuK/VeXtH0L76
Gcsme+TYSRLbWg7n2iYywd7aI03f3LAX9rfGAsQjvmyMIBdfIbtAgDusCNZbeVEX
sujdJrO04BKRPt66xMQQXyiZ5mgO7lKaaz7vkcDE8r9X6376AenXF6HrRPthfOu7
HIH1wJ8/dgOUp80gvCqfqMxZe9cQttOcD55hqTSISgbOlrVIbxkXpOQa7mYr1SqG
XQpXt6KGoi/nRxCT1xmxAOjLmGD9HDLz5+ipxbtGGpdIxwe33IxCjGkrHzPaY2M7
A9/gVeUvXCHAN0QGWY5BSJtNfMM6DtT2t13zSEDFzd6Swt5dNUPBTMLDbBO0+TKM
8ZOb8loQahOtG2ZeS6fWmB09p1yJTwjqYQjRpH17y6OIgxY4t0zf6mDLQg5oB1Xn
7Qz3B+gAffKdLUsiXtDxMHL1YO1nrLY6MqL/ZEIOBlggoBYCfkRfAPR/iDiE8mzv
8uHd4r9HfTJ9O8xyHD0hJixl8h55qB6OeWqKnSoC4R1g60dnd7DvDosBQjeuXBBg
+uD1EXSc05PB+EvP9V4NLOSDi9Y/5QBEVZA+MbBVZtKSVIrZnveNqfss3diWFpbb
dKxdWrpUxmObJgthS6/+tECsviW/SxAZxoHNiU3KpltikmfhWKNUjtRHMifqr1Ao
/8o4zOc/LjLPHMbaRYH9Y0ho0smz4dFecDtAXyDJkMKFW177GDfZvQhrwboAa5Ra
PVdwJtdzMnCabSZ0nnZ4j8A3AbHxN6rW4lv+ncBBpQsD+N7NoYcSvAn3W7uz3Lfw
/ebbIflkWKdoo3Y66dp2vYNYUsOV+irskejs5LcygNuxQKvvJbSZtQqHkMZ2f9FZ
DMMUTc7kAnLAy9y14qASH33Si2YgcJPida/H+C6jmh1oVYqdyDX8x2nhw0x3g5gD
wLFODcA9/EPMWKKUfZG6YJO0ZYP7/Yl5tYnW61BuBWZSf0LZuqeae1FSmjcl+tRI
LDkSKnwLhF3pOfLOIIksI1R2qYRmqorrlnOl4qaBpar8xoMcTQTvW7oSnfXnO/Uy
+mtRTThORsVqcEadxMH4mQFvWfBTCmK4VOCZ6KdZtWTQPjC2aftrvAsA35pya3OY
Ak6GuQIRDi8gb8nOnaThWlMgvVJBA1KEOf8oiPE/0XxPmeypV/QHjsgLyYDscK0h
AEm4fPktxdlT5h7qIgxX93MN/wejuHpRxubEhCMn7SU4/5W/0v4phaydVVxta0vW
4Jydwf2NbsfvLbdXZVwdc4Rv/Q4W1Vc3qY4ZJg4+o0k2xDmB8aExV5ermYItPC9Z
1l742pRgxVzOPRaRj/lB/qtVMIIQFtH/HodeC12CRHLbf5vtiebk744/kB7qGY48
tepjZK0z51TpYLK6MpVAqi4RGRC/ZNS+bcObl9dNE6l64SO47OSxMON0eMm8J1Vy
3fBsIycjRqJoXSFN0lS/psC/ukUt8uOYVaaPtT0bZoQ9uaplU22z+7kXqwtKXsgK
5WP+aiPoQsr28aJ/HAxxr3K2bbHV5LsBC+RdwBvhtbVt1nNj+IIPJ6Afi44+7Irp
F0v1FPIMnttySc2gazsQZERK3ZqQNcesNNxYOyEB6WNMxKT4hlTDYYjzSmLfGzlz
A2kr09aDNcYY0PhsIZCjk7qWHURFi6Nl1IVKSokl3AeCk0dQbXITtpcdIty9x4+v
+Rlsss8FgoZORDGIqrbQBaBf1CkIeQd9C0XMJyg8BXqDkQWQsQqgWZXFrUXVAnL4
bipHVsMfV2RxI9lhmEM6es9PpW0YLfOH4uUxhXOBU7IZPAFnLgEhMqzsYyQgq5Lf
HaYJWKYXy64Bc6dwoUz30DudyCUyBr6CVMsCkvYVcI3UUy65WWEampplhLIDqe7g
DqvQ7igbVtQSMqaH/51a4RmgTl7jk/YlVI3wvZpb+CFZYlh/LILglYdKhfO+O6EF
To4+Ds2hExXtmA2utuzRUm4rIt1TlJ3Xb07/GsKZJH0ZAN5oHd3Xbe6tsxMaUarz
UD8KvPYvsZSxNpyYUGl1yj5Hnoj+GqwIY+jBXUXvuhZ+7a3yWcRiCQOjK07y83A2
mUJJBSoiDF+PAqjZH6d4t6FMvsQuxmKQAsrzBTzGQDYMuxVaGYimTPfob9KHglMn
D1iZlBGU+F/EXKXDjyHC8fxyLPFPDR3zS5VcXUe0pll1TK3FZg2VHi9hGyXKt28D
PszTW06OnknK87ri6ZGuej07W/mpflLwhw8iZq4IYOoKbrwWMYRzlsJGKLlS8m0j
SlqppcIZ0cxFS646fPkMxJNh/2L2/AunQ3OWENuV7FKVtUoH9PvasLGxoOxqpY+o
HTdTmtDIlQV0iRyk4gfqDplV4YsvwVTXg+uQs+hquQDVoVKXIEd3Gj4Bdi9xFHre
26woNXlCdUZRGIxnY4Ilv/KXBjo3tvKw+ZNLWPH5CGZ3+cpK2Z/QkxfjRBpmejYm
ABIsCxWM5l2X4rfaaD7xq/Wv9QgyGkT98I0I8Bho3LJs8Bzsl3peB73NAB3kRRhf
otRyrg79Sc4+pMKevJGMA/Vtbsxur1c7cX0oEvmABzi1kC8muwDlzcRHPsixZVU+
iiZzFQxa2lgdet37STL0J4w2sqncndYmLIxTYp6ygJM12jEf0ss6Y9LjlVRCOC9E
C5zz872GDE+K8LNNVXVfrxt/CAq8Stj8iReJsh7FKfQgLJKbOZuyHo+W5p3z/8QD
FMdhXPNbR+wOg+tai5+KjNe4pl1b/rtwa0U4fCNs7TnHJBiD7KPO3cXV6gkLmNjd
1EW8T2i77kejReRCvQ5v7pRak8cEAbfBTzvf77hsB5LJkrrIMUtjnJ0vara3d7nJ
b1eN/oUK2qcX39JHV0FXtC4ZIOZwD+PLrotknbixivj8wbstx8AoH/g7j/n/4pR1
/OTqFiLlB2t/e59UCEoMDikNk4kaWU/kL724Pp9UI/X+5iYTDiyJ5+AvwyaP2ZC6
F639MeVm2YYe7MWaDfsDKceWzBbdsXNSQp49AbGX/VVCtjlgsAPp/SO+eAIXURP2
EctFCWE14+arYYNLtghAh8f13mhSLfscqQAvEbnZ8BZs3Kvf5OI4U4O0L4RtetC4
kkO39FAiohXrrL203mnM+66WuUcj3ML4vOicsX0Y8bk1pIge4gsAO21aHg9xZCbl
2rt3uzhnVbDXqcyZCgXBkjXvgZmd1L5CtTd4AaV7WrRIFf0w/oQlmrDlLrMPpLGE
cXTOSrasjmtP4MHAcnXx+UrS8evpWDnAeHpaz86YyfDc6fNnIRyspnXUrPUy5D01
CIuhdYz8PLsmn/2d/7MeTA6Frjwy5e3QTzvI8rXBET8BMbSCIYUVMBj/WgvBJcEC
eUJ2r8zqIUHruOjPodRy0hBUpK2+CJeTpeOYpC+ikOTVYMC+kCCUhlAsI3cwX7p/
5w0Zp05Dz0gITyMJNYnpcpKAeXmqHYR0Ac3ALqxpAnidyc5LKdN5mrnsFZUQjemB
cbgUJz0i69VmjjSH3V8tWGHUrjZVzPSc7GAAoWyEB99a7LGogyzX8j094Z/XZQ2w
w9JDlkSHcAoQcQWfWqZ2hjKCknXSaYgrl4iqNjJwtrfF7b3tiEqFfRV3Bq1mv7Ck
AWJ4Rft9kC//+L/5lbpeU3NilSoSOl7bc2yJ/6KyujsJkI/1+eBpiJ3ibRLbvqYp
a9RG+T0S8pFzbsHsqCsekMGcNdqesOr8B4ODbMwlz4e85CSS5zFhNS4IWTiNZupp
qiL+6DzDcMgxMB2XENVcybLHXuVwqB+sc9XtnVbdqGsiwOM5+r2EzhRoyfE9piZU
Yvm4MARB4rKIfhFbvgdICAk+8yxtoJkL7IRIBwAIUkEo/NMNSVb2JqaBhQ1kEfOx
ZGLqC3E9PeZi2wWaozDKIxORejAEP5Tviwjt1e3DORiLW//yq08AxoDLPI/nYvqt
lSYfzvUvUQeBym/SweiQpjY1Gaz2Epa5VOvEPWOv3sSt+pSD8iFLaVdCL6ESkwlY
dwIoA+5gnIpqALl+eyD8cUkn5WiujKqgPM9CGMpBd3hIyhRG8PFZKP4VuWkWXe84
etsfo8aajhp5XVRsoTp/BBHfux3Q1c+0aA7H+0CY8nu7b88B9Xg2ie0KRLozXiqR
yy+0EA25O0L+M1+NiNDYmSwK5e9nPKKJAq6mtvynrgvvbBOMCbQMnEIMqFEybMs5
dF+27FThyNDXdRx4DAxpNxwaPEDn2TmXpVVJb3iBXNX1Udgzj1RSMGjTLHkHcpV4
Qi9BnYvfwDRN8o5rmqqBLC0pyIBoMwQGpthN4ynWa+Kymiv69ubQXpBRUJlRIZCy
fiPtbuH4ggenWb1VnLbNCsfL8DqgYuNhzIRToA+6xh+rsBgaMiWGV2ZdfmcRlfz5
ikF7tZ/sxqqKDOieEqIf+sJylQsV8MjBN7JTTT893KD9psCzcqBgiQ6t7ippZxRd
Uk1y+YGN1kHLmx4X5SejmyTW6DuVVuQIBp/bDySdQ7xCBS8dOWjmp9VKR3hrZ8nu
G4Vb7kxKDA+7BoJbJWknQIkhg4jYcef9jUOEynIbsQjVzy5gDZ67cMlvhLvOixS/
ZGc24c+rAXMzUNdkIRm0bEO4zHjQymln75GOFY1UN74yV5JG5oFyzQPwcTKavVjX
oLnH4rvglhul70H+Mqu5q5DgWvK+M2tfoZcfNyESzjnoTZo6zZtNsfgg7p5pSpZv
ZYIYFfWE0AhVL6qS7FgKJqmGZz+Um/22D8iY2xSNobzrpyvIl8073uOIn0hMB4iB
wyg/pnxBFjBPqeshjKiBx8YG/20zzWApqaqiJONz5V9uDu2c9rq7sd3QTvp3NdMB
BgHda8sf5huY1ZigUWu7hdDyflqBMn5D9qTWH27PnBLRDPu+q293hBu3rzyXmlP/
QtQvT3kFh/lJ8wWatvKcOOQmmUxG3ICIrvGbEqAt3MTpImI+pf242iyVig5JBer4
+eJBLSEFl5R4mTWmJ5spk2DnriT4Kexu48kgXKQSwwu5vZwSop1OabljYQxgqCah
5ZoWjs/hgvb0v9Yr8DIEkIeinhf2qUQvth6AhIZh2PoQaMHuq1zi0aXtuA5RuZD3
wHijJgRzPNyjLxABgmpQl5qOMiLqEtiJwn7OQjXQDKHE/IkwxyfvcxQ8Zorb0rAp
T2D8ZX5p877+kOojJ1IXtPK0ulSMf4Cv04uuAE8zuL/rlL3MOGZh8oko6v0UrKt6
1aan0gHy8nkP3kRcApcJq9113Fke69+5C6UPqw8gcEagjwKXrY0qNGdKw8RulrZf
nuSPeMHwfDc2BJ8o2gYjkwiaW/pA9ZlxbQnc9s0zOGrgAH7rUMUHGL6UggIgG0qv
aEyinn2mVPKUBywjTP0pg3+U7PyAA7aRNGmQkaz92/IXG9QCSGgxeSZYRFPZDuY9
QM1M7X6TP6BcSxYF7ZeXBQIRpL3YqJVbVPCnAMzCja5JpL2U1bZOh0qjBKEcHUGg
/BrPHEassOe4gyAB1zbiggM2e89dpbDf+w3uTF4Pfk1/jT/DrYJnDvh/3UYrrmcS
tdFEDxftiqVBNkvDP4m0nLntUeCucYQgs+5h+o0S5ecQNj/iL0CNhAs7aBCU+US5
Uf2eKr1i9ppa8cOAiyiS/jwvodeka7i2V5MYqq5ZEK8XqKvRxwDEMQtR6VbtvgFD
AR6WJHh7bXynMnS+0lsKDO00njY4Inwk2Y4NTYcj7nJQupuAZjgQtqZ3LspoPnvG
tv7EUYHYAvQYcSBmMU8ily3+QGN++zGeGwklAew3ip8Ip/5U9c6/NDOy8PUR4N+O
pg5msy3UIPhbcjv5t+Ffmv/rlUd7oVHEEyDSzm7jYbNIji7my8QkNvV6DDQSPfkN
Dcv8E7jTrM3ekPHu6+yyMMo3HqQyVJg8DiYtaK5pDONIJoHa3zRtYRxNhxcBgRl4
Cb29+5v83S8BP+laCfrPH7t3NQwwMufmvAMnLD3EgvZ1bECpXmPsWYKCfRCexuld
KSSHJdbLcK+aSUqYs/jPpvlUiVMiv+K2kExaukuze8Q+hSPGqbVHFwKxB+dyX2ee
rsQdK4D/kEaMkNIjxhn3ct3GqKfuV9kvHcTgZo4QY/SQLq/Fi8D4wbMECREQV9fH
+cLG0Y8Q7pv5cVHZEXidTQfK9Mfmq/wKXk/fjOE5al0MOpbgduCyMp5ug4XKubNk
FwFa3M5X3hohUdgoq/3JFrtXSav8HvffAJO5a79pxPkXgUpyY1XW9P6/4llgXvhf
LVT/qCtAu3fbInCmW4jari2Ium/+Ngt98B17HD6hU/FaYRulUGKJBpm1HEHG2oha
ra9ttmROB00ZaPt1WQJw1uNdHDcwyh72LNtV58ZO/k5gNEiJc9nm4qkMPuWWNGeC
J2G7MK97jPn+1Q7Xz3OItxN70vDO3FfFqP9RxIm05vjXR05nJSmTP1wT8KAY4uE9
uNiLl0d6HnXKJeXTzkCEPNpduL4BWo6+daBm8Je0RQOSMovgnwtKaormLo5nSJ8/
k9fiegzrMG80Lt4RsEagCA7n9BhgKyUcXjtWwtZg7BM3J3fiFfsOsaDi24p2e4bt
qmK75WrNrZa7KnIy9rQT5BTg/Te7m2bizxEnm6hCIWr0UTHr4lryd71Jqe0QNXIG
hK56CjqiJCLsMXDIdN1foEpUVxAmlkn2V8MV6ZSTjKuf8GOtcqWSHGA5cEZbYYX0
iQfHeQjeik3LW128qG2ZYvTPsBb7oL2uLZw3zEl1xO/BYxMzRWHqAFMGrMrKxVBm
ic7jpNkEo1DlyKLgvet0iVVrnfRqlBJCzC3H5nQivaCJVtBJNwF4WezNYEhwedWH
a6wSVax7+KKgjmMoLZsZMu7H22qlTs+AS7v36WomCAlC3QJ6m3gc9zHwhPbuuJVU
UmlQkX9PKegYkd/YWOcn480WuwLXMeMzlIdswmDsni3RCsr5P+IBRw+xKHgu6VxZ
W576czbG5H0BFUYgRWzzI63uwdM0yQBbUhRk+WxZCkDsIC2zhpV6yMMnQ0caUBdk
bCmWOnbpS9xoHiqx8bO7OJqRwRWjO2zGOziU6QDmL37p46OhQXggZ2WdY5EZEuU+
/qwv/9bauc8+FluRM1DY2j8OM/6FAX/NcQ9yljIAqcoOFddoj6NL3d1AnOWLbtHM
aqlpRGiGuEkxgFOaRidK9WD0te8VYi39iW5g4rPExUnHJg0HDY9oLyfF/jBYAvL4
Wp9+Hz9id59t5B+kRuHzII5Ykj6ZwrHrbVpJRFrapUVmpcJVGrbfvxTwm2gOU0SK
u+o0mUcF/YK57cAWv32QRjul+Fq0y6q1PoFLARRAtbHaaRSvdBJGinaBKPv2Ihuf
lBiYTa6/EvRgzRjWwlIhzn0AQsM38G9AfGGsmAekwxvNw+g/QNdyzx/Kwz5jaJaN
vU/PD8HGbS1G4++sdLrIjFuZhnQup5VJR9cwTsAXiMXv9m/pQ6z35rd53qOlj5Rv
bQpgJ6AEmJXxiOxBeIHMLXxfpsChrhC8xK7Vby/LvwW11naDBZhlClU7AqH19hiv
KvTzb9yYuXw/H9qrxXzuXk2ZWQfHPVuSeGg+ovY5JtIorDZQQENBh4+95LXPFE9z
1CEiAMINCE0VlELD2Tud+6bvx3HWg58qXzMrUwwRa8Z6C1KHvA4oDq06TLZV4GPJ
vMG3qj7/d6zFXk4ir7nO/K6GoHhyZ2MWVrs3qb1XtPVBECAjBDUf4c67gTYV6JpG
UaGwadWoGH8Kkl/SeIpGv3WmVtz7XL4tqmL8tCCd/GzdGjeE+7M+U34WH+CGFZgC
gGluEmIInO9qbInhWf1eiiwQFO2nMO+GMMHoYl+tuCKN2i0ny3teBvso2B3iUKtT
1Tw6zpbEgEZ+tYMan8YvDaA+hmjgwkHVWjE8kFQcjfnxi1dZj2628p64xpoMvhbm
4r333dtMGR8lc+ubu3tZWGc3LFPHTA9Fu/8A/KdwwTjF6mPdBMVN9L5KyuhNL3Is
oFPmXvQuvNJeuPWuD8SDDdLa5cQufrHxwhsxCDgvesWbHjWLPoacscmboBY2EB24
2PYCtAyODmnhdTvsfIQMuwB2v9X1f7ixUKvp/prr7EhEhbBa6UE+6ydpGpOHLvRK
01bMKQXR/JG84KvllYGrJ4NqzTe0dqaInGDIAS6ybwRlzbtFDr2QHIuHHE9+6WMJ
bVRP3hBQNK8cHLq8ojyA77fgU25+9SSOMyYiCnR0geQMPLMXVralJ7BvwYFORweU
FyoeXW/EhM7RUrTg3YKClrvIE2D+5Nntpvb3sjSbdJ8Yf9IecJrGD5YSDTwYu5tx
RMoOVg4vMbW8TfHVncRzg0dayCLuYGQW3hCVIzcelbqAuJXqY1XFagKbUe1Z2XaJ
ck9s2p0xyb0yzoPG2OVtJ6YuoH3JjV4Fwj6/mY3mchXcsIRx9R1eZ/yYkxGd+Q8q
RHoM4TLVKmlMOAnbjKmj4mqYdvkkN11hAC57iGm/Alq6Tlu7AgXGjiX3i+hRlrQI
pDqm+wWJm0KCmXb2+0dPKpHuKHMD9oCtl6pN3gn+pwAOOBvyy/Tb4ka7U4Q6oHWx
mQ+HLzyeJ/n7D4oCAGQyU5Max7pjrgKGg0Y98qmPJVAWb8CAnCsHNYn31yEDTNIs
cFpZYMiLmZvEAYE4/nMP1rPwT0Z116MPQHOGI2ZuIPlM9ry2vd2tgUvlEwO83sTE
3Jlz1xuo867uENAS59j3ZgslFwC+JVzHaWrFV2b0uy2Go9v2of0v/IMS7rLMES3m
icLPY36gnWfLvHuQgnmLg8OAfeJnQ97p9XemJDkpUeEP5+qhMwZesuTlG55HQDKY
9LPwJcRxLadyieYsgNrfshbjfmVl+FvUEfnuN5qyxp6yX1cTncIffAJfi49+bgl5
yfQfcfKNv2kGIOk6UOr7HihOUhhosC1bdmEO/hTtEQ4svte3aiZJrqP+9wymflga
JykX2NmPNz1UVSAGSoAHpU/LjygMPCbykistXDuhGE8WKnLyN7EZTk5xUszZRbQz
3I9ZCGBwnJOn9LWI+yHpDdzZUzUlevgumHDmNyVTBxoOIvBXM0n9dmiKmUEN1t8h
iKXp+oPqfRhtyvAOZHmF0flsiKa1rxLi5ZAJgoaJVq6TT748amYhtf9gPRhQcU9u
naE7xOacxsWG3vSaPZh5UM997zvrlcEHc0/Gy9hgbHD/98xd2QiT87NDprihOcVF
w06FYn2qjzAWF8zUJw/d/06lnuszXlihs7rdx6kPGB0O42H2uLn/PNgn62rtS+Dn
S0kQy9CsnwmSnczI2YlL71/uXgKtKu6MJnryv9Dm6heI3bhL8XYDQ7xFxnBkLZl1
id+GNE8BZveIXXUvCwDGHu83IXdcVKSmRa0dGh19XIvGRkOdpUbCHqIL3jzmyRzK
NqlExiRnaSgAHEl3UWqjoUAr1EUV2aspZ3X0zOyitJD2gyXNP1d/TDl27kE2wY/4
vwb1ZH43R0AtCzLASrRsuKvcuLDtDaE8zi7NK+zC+gx5XZDuQAoAnTTFD3cdb6kT
hWykW9TvHR6oy5Oi/ZgZlC0C36zZ9QvIE1xqC1YPAtdwYTtOYXq93LMAqQQqGqwH
ZZjlXt/pbhZXu4jYD5O8vahej9dpV55gJQunYXo3bILlYgsKJftK6t5aQU9keQLx
KtWZy7g8WtzEKonWOeVPzpprEwxeSIsXAnnzL5gDPOkcUT1q76PvMni2WtHgsk7H
KGUwLMaR56FkNoulRj+9s/1mGzyzteyP6OsGwUx6JMpQIohIKP7plfykF4eaigtJ
v/GMzsDAF4/zQajwVhZ1u0bPCTl+J8JiqimFn3fA5VDEzPD92gD7e5SrLi1ziK4X
FnRc+b0GO1VLc0GFnIc9B/CfMZ1HYR+fBpKb0KoEVxIVulq6hl0HbwNOwXG3dz7+
RWv3toyK6+QGfDYCvGpewucqs40xG7Xn0dWtnf+CTR7RikIgewHYbE4z0WPIWDjj
wH93p/tCWrURbs9vkpsqN88jcar1/iKQjCgEdYWBItahwj75dkAqK3z4rQXIp/wW
1HtA/mFDXHdAhiL6jYXQ9rn2T2IZLtkg94jURUm9gkcqtcXAzHpz86dqousSlCc0
YomqcmxdRGcH6RvGxDrcXpjUjJiga5G/R/Hi5cFQDOZ8XyB6JgPoJPrZ06JVjUnO
ozCxPJhdj5kdcsnoo9vvd6yaT6BQt+kSiIRwYHAeS1Fe+huv+iYfRC5ok2CJbNG6
1w/C1fq0sVY5XYX9bUIMe8fp53/DzKsxpMnBYPthRhVgQcOFh+Ks0p6OYQ3FlGtb
T0l3vJ/Cbc0o1B+z9rRQ54nhxt/xkHlg5KJKMLNPS+cM0oLMvXe6RDv5DikOLqGh
jAiWntWHrbVcRK4yJ3cVsoyRF0L2shW6SZ9d8RcNMYVs06wn19iGt7qF2zyI/HIN
HwLIeVNHxfVAD66ev41soifkxwxTBj5ftZt9GMAhFwlcr6w7wN6a0KJK/JsFD2Nx
ofppOco3m5RAnbh+bdmix5XaciDuc5SHcGJiuQ4h0YTrsiVk5rK72n1hs7g3U//I
KtN8C86G0NJKE9/u9aZnTV7u7Rl5XV1tAPNejO3CbnweGGKH2pLqu4J6FcdvISNT
VZt6TAVy9cCh1Xw5sfJSk4js8p4Nf0SSrjSiSGO/769BaSkk9pSaSSlDFeTfqtV+
yogvnith+ch/JtX+IITctPOUvWSHMDRaVo4jXTKgVNWIcbRV6IsW/6NdkIqLYu3t
Yt5cSACf/siiG26MKQNxUAtCY8veDg14pxUU3N7MxZauVcUkdPjp/eoHXpRLjgtP
PFu051Q21OxKbXRuX0fo4XVxuamj8QUvrzLrAKtneoRcvQwxWZqoPWeZb6r70Fry
oLld5rrwU7f8fATOFjkkMAxt1enfF+eRwDJ0y8Cj23aCrjGopItshLb1YtV+OObv
AZ95scxxQgWARoAvZLAGMdfHCUpDROrxZ0GOv2o99N4V688l4mkJD2WhMOmC7lkL
bNiWyGbEMp9r2t+EPecAj0sWCT7vYwFpn0rlrfYUOETpy0sHTnn0lS7Is/rt/HlH
lnVc/KZ5Vq8kLjtyrT/cnqkrZr08z1oZ3fItn0lzTFtNvMqSC4P8wXSBLk1VvYow
vY8YnfdOci1+GNLS28EJ5Fjn9b4t+SOxSnyKfKWmZwDzuDYkiYyxz8GQ0EkqJtLa
yLPbfzF7OU1yqcTGbQQNKm35myUyGQ867Mf4kgvuQ2ynFmug48MzVQPKaT8XsNBB
PcqYfqKITQ/QcMhUEnBekAlFVJtQ8kmWm8L7VqcrnCgHWw+1TktHpWZ+eQpQoxLr
wPdXIVh1Pw91HTOk8QnZlKaQhNP2Kp0851VmSYwQZXa9PMP1KhAG+FwxPl6tg11h
2oxwXtc4Mu8qVefAztCVEXRKTyOSeAMwOK/yLsw4tcNTsJHvgacdUAW+406Tywfj
JJdDWJrMTVxbROWB2Wn1ubc93yffehFL9Y9r20gXimtaRRy5N3zbun6lXcJjOUC3
ywCuHPtj3MycvUoAfakjliWcqZNtz/W7eTmA0LJqR1YVK/CMc5Qw0t0xNuTar4CU
YxGgK/PBmQ7S+iMd86svnD1rhjvhe5OB/lAwiQ27wtrxeIvFffEPanWzR8ShWzkS
89mYfLbSIRdh89n5y1cTJz9hYsLd8JA60Ts9XbB9rmx19H5ExUUkYHYB9RY7Qy/d
QefzI5Ef9fBrHMHdKaQOnbnwq0wZJQVXRsKihriz5cMdy3K1dmHPS6Une/KdB15P
boyLSHzU7ovINMJUFKANMKywHaU6t+s9lXA6dW75Fk4Is0PDQV5mT3oKqDr1GVsm
dn3uiNP+VSLVlrwPH11mhyJpAu678MkIquk6YQKA9tyK9GYfgMEAZQkRXJWPIDx2
qECzOGf5niybTaqRvOA2GgFCJW/hzneYSsm0/gkT7wm3SUhuv97vWxjqgQVrSUL/
lUnLWdFC5T9jPemM8449MeGFqcdS9jL4UJjlfxfMRKsyl3VyhPlimBOfR5cF8aGy
jMEoMFqBYKn8KX4MIuLhZf7er+pPesPR+5uKjssHetSitsmao03dAJOYH8bgQWJO
kr3UEoNIIEoPKL2MWAeVUN5+LBrPNnk6klvqxOT2hdeKLnpcZDRLaAcaLwHHGeFc
XeAcbPRfU9Fqpcqg/5O65xDNkzzey3UESnWJgpZRUvpOYW8Ki7XwBzHrH2cppwPj
XUrHx2GkkiJkoTPDlMUzgKDh8Y+ya+N2MCj3zSHGaKg8N66I7h8GmkvcyQgz6IxN
5b3aYZPJih4wLi8FQ0VdhY6QTKvmjVfMd6zjB5ymivME5zdfHkIqRYsbgI7t7JTo
K2NywiQb062ikU32fZJ3egi7M9Ww4vKtRtrbVE+uvxVMInl8bqEa7DknGaEQJ4d/
rJjEsJgdcPyohios0sn+G+ziYJCp/jLRHHm0tltmCmb20ygw9MIZhE6G8Y+G6rt7
1Hx4XnrwYw7Ds3vgt7J5YVcNmNOlQrkXLApFpm3jw3JBW9i+C0aIt4x595ZckgKU
rEKDYMAhnLuoN3SvjvFpPxP7A77Xef9XCcLUEGHxITN8Aq2sZuGBGgl3Qtv6rKK0
QO82AS4ClbJsF2zig+u8+VKWA5oBgc6CqymRkeLjPV2I/8LgC4YdOTWU/TH59hR8
CcTIIk535WLpp/0BWLqFQxxlKnWOMu3VzZXIb+tKlbLag8e5GsRQCVNlQ9CFGvRh
xXZLK9syNRHYSKdLa8xsgoq8Zd09a96zAOtEi3jEDFRpANGsrjxTggReQURKrOHD
462ueebu6RkHNN4majFx8kpyfQ8WC8Sdnd59+52MKEkF9+NlQRqxifpk8oIfzxij
leua2DI8ftAP8DfAnfR+x60n0WYmWZMYPc9E4ApxtQPMSmC5hrsJtIAcjK9VfD47
QdyPj+IADxQCOsEwDWFrnJun3vW0SljzfLlSdJ7dTLkAqNWXcDlYEvoNBAeYx6O1
r+bIa5L6GLk0B5VgK0YsFOPp58AifTCYbpnKPhxCeP8ApxUNuSpPObjAkBa+58kn
gL9tf2OyTKa/WAcx/Je9Aya0y7oZAglyR+S1+ScqaxweRiBg9+Ez3cziBSGqBwy/
78YLzBZ069MgAIeXNagc2Dv5WyoNc6LwF02+l1r1ZId3tDqLYYjiXXJvN1+/PFS+
frMD8nmlJNw8FNTaT/i27ceZFqBwNG0Aas+F8kSbz49lJRFZd/gzrgvE61A9B0qg
8QEtuRY614Ni+f3TuZLR9CyhEunnvnLdmMiUAv5jrEWizDfrPdDxaF0BpaxcfRI9
S7XKc2WORki6sDno6c/1BFQuL62EBkZOyt8jaDGbBp7xCbJE2V+S5JxXJYzviQ+M
ueGiIrstnfj0G5cGqZPX2GRYbOdqhqhF+aHsZg69mmFpOvu7I6Fmb1A4hQ2J64D+
oxVZJXY2F8MHbAtD/q827XRo95/6U8LfubjjSz9TasnPW8bNVqdUMHa3kEB0CA9+
Jy7XdZy0LRpirzolR0fadMbJfJkQqKSy2P5eqtBWSQ1aoj1s62wpe4JFsFFRFT9A
pNPFeqENlQeXcHxdxtmgMbw1BTwO72FOAW7yT5sg6YRHZVSeK1xc6i1VKHgDurZk
RP1Dc4vriXTZKcUN84JxfrQaw0Iru4q2m2JrAO5I7OEqZLvSX3N079OekMp+1lPX
1Rizeo0n+5CDidhTPL0V/M9zfu/6QQMFW/KSmy+uH15b15/La40iOasUbwAuLpA8
1Zp26M8RqrIwtluV1Pa82hkBLPBcuodcZ1bOQP/HKIVxsNKdyecD2oAqsa4QNLnJ
ZezZM3Fnre7ksOo4hgilepe/8WPL3yMd4WFqJKURMrhXF/tTE5q3KbvVyhNshyBn
AIo4+ihf8tDgfo3I3AP2mS5ILFwuPgN4/aAuW313L5LH2uhA0L9uE3Lj/0zKVwcL
sj1iRysBRgUJbz7VaJLzRtHzksEDoFYCEg2NF4C7rad7nUtpefXoAQqhoesWua4m
W2YoEsayaOy4p6ypTjE5NHa9W9VGWeKBOW7KXpqTVFBCQUVm8vCr3OkGaSA2WUsQ
G4ABTMsPJM7Zp8RHYk5IlxFpFy99OvdmkSCLBfX19+e6PslHPFlbZ4GKff7E0y5L
LMYZhehfdd1fDH94b3nSfrjtfIfbXMvE8PfGyUgXm7IADBfy++FmVZohQcCS4Mox
6EXF1Q5ciB4Xffquzx9+2gw9jRBLtymN2HDVKFkuXnwaMevToh8WudMzYewR5ZFa
FRVXBq/vkaH9QFskqWHy39eEFrpmBAfA/UGV5uipYSpVDOxKaDZYD5Wf/bieD0Qt
KKFlbj8v+rUR85hXacha/R4pOJ1SjSWHLziCH6jGjURNYwPL2EgQb06TztllhrLK
SFOFt9G4IGfvuFJugDu6h9L7IQDgqUKxSdnKL+CHOhGnDnA9JbtV6nu8pfPDqfkX
Nf9x6srbmxKq1dfdpbc9wdJpQv03b+McX7a6p1lCBBr2vQvX072rgV4vlftOQJXp
wTutdrL5CdQdcJmoirGWum0vOVtFH5CIIiBWJDT9A2QQKBwjr6E5YyOy98L8ZAH1
CM7KGFZS4IIcpH318y4pV3PtydeKcOHV7tfNP9F6uOhkgMOqMBjJZ+/v4vsZTfGi
RTifBOC4YOsf2fhQCP1w5hefwHJr9UjlYBXZA+MU3N+5FO8jONJPO9xr4jVM2GFR
VuK9LN3LF1nLAadZH2X4glZb9E45Pgd6Z5H1twkMjnrQmsgVdUbEulWZHxsTMwnd
dtoU/HfTNNwUYHLI9VUbiWbHQ2dyPfjHs3slxeAkxd/A5d7m3EIXAL7GT15HDn3Q
1FStZWJ81N0X67a/JuGrW73QvV0VznKbIVgyVchBEPyIKcfch4BaaZ71moz90wVg
1LLTLnpdZEgX7/gvZE0w6RE6bh2AnK9HoTabF/WI3jon1Oyd+bHKmNJb2VMzphfF
qkYSOuBbXrb3+2PN9YV/Bzh66C81f5aomg5g1wPRaVmM8VH5x1/9V9+pBAbKfRLk
WJySBMM0sw0HxZY9O7xEybIMC6JxplaTVfL+u7J3Y8prlhOh9KoxV58rtgKrm4T4
QCxHby6hoZcBXviyOcniiRPOFXXfUNowtx1izn4oSDid5C79ANr8Uv9d4yTF9n64
rUKguvmJRd5pI5ebdWizLfBdQnGRxiwXyLaALYH/28FzeyhoTw13AWW6swxkyEGn
NU17/vY15WjvlhOr7KkLig0VbXVs/t+CuHczDMWjF3CLo84ITVIYN62zo1SGjqj5
nW1sbs52lsfDIMssH4qnpazY+pp8+mCTiu1+Kb4Lsb4AoFtlpc2VJ37Dww6o9SK6
uD4E9MIps0v20WAj0KWksifNdd2y/v+4I46/22AK3Q6j7TOFwj41bhIOGDHtrZBW
rLmbCjtSsXyOuvC5ucnyb1KNhuG1Be3PUaLMvyn6BUiartCmfHHxwzlAPJLTX/kq
XyksaDvIFpiInfNRaer7eI2TA45qdYqftbxbYpl6u9UDaOBDwpIghsxEFZbkVTMV
lBu782e1BVWKsUGXdiBDZ0WJSaDXUZE8jc5R8L4drHVmJZ2Vr94fFZwPDNzUr7YO
KwMXbyohCLKCTWrZDw5PNfazqtDYo76Yyop1l7TXGlXfb0Gh5w/IN7k59BceHJ39
iKeIu3zplgeGC/13nmrajHNZQGkOESKeAzFzu933twiLi8AZTvf2GWBq7LQ2RWYI
TF8AA49Dyhmk609aTbWCFpK/8qhvDNJH+tNSnBev6qXKwGKELuCuTpDBYGcJ8Z33
r9/RHCruNTf0KgBK7ebms66zuPgp/lYo9Hbul5NQQaZ2ZkEoTfBJ0MrEkmTsII31
WDLADokz9SzzI82TgW+C4CNgr6i9iLrYNi5IZpiCZrX6MNvet9prPFLONE2bsviZ
yejwcTgF81yo0KTQlogrnXVFbAlLquIaDCpClcy+qYkasDcK3RwOBoQF9EqAtH0j
jtxfbup4Vzdbge7Hi0ToB6JvihPZ8JZs8jUSxQnrfd2SijYc9NACj15Q31hz9zX6
uXQ/JToKWPiVxVpwn/fS9H81AzOlvyq61A4OHOR70+MjPB93gTtuwZTPX6XFTjBI
2r0+2OgJBMozJ4Txvo5wwWd0gKo7BJAJX49OEC/XsHc/FlTCRllIr+VsKzq/EjlU
ZbfEAM5yMzvS6qr9j0gwY3MVAqKgxfEhQMmLf9ZXVpTZBlaSKYm+1zwYJR+EZmdr
oLWAMgKDt6FgUe77YqzYAMheZNTW2t0Vt+W95c+eloVX02ymT7nGm/GZ+WFGzlcV
rP8y+2zy4/uaEA0QqF/zblF9Qx0jOzrLMGwaC7Mj9O8YqtlUfBwyM2mchwYyCxgn
vd1rT7ZRq3I9/Z5LKK/xaEt1vby0SOLeX2ANW49YKLng9rOZYbLfDG5jcTQPci0G
z2BBynv5NPuY2HaYSIJiPYOXQGnbztf2Kl2lttaicDyWv5YJ6CSUxAVIWyQhkQet
4MkcrYGExgxL1ydKXgbqGwaHhTTUit1s0coaIpwY7oyH0TKlsP6EEzV0oVgaYoWd
V2p1en8YqwuaKNA61/DQT6b/jpODaKADC2+laSx9oT5/9Jgbgpe9hfVVzxU5cTcB
FuxeEjd1+KFG8I/j/4Aykwnll8rA8XAKf3Z06pg7DHIl70PXtxi4oBiG+UbAKNsx
py6KoCuXiZMuynljQJF5jbSCipyZXCxnUsrm/4W39pRyHvHjMI5Lec6QS/DBg3rR
vv5vIaSSceIBnTkdyWLp4cTYAtOYgzma7W7Ic6kQU6br4oHKz7pvTe8dLJElstoN
YNGjbIWZ/c4S0HRtUwhA07a8rk/tkI7efpaEw1ya9L+QnCbqicDFfd8HxNg3Xc/0
aefKAtw+rQ/zcZFQNje0Xu6bXf7g3YGURdOrxrBvpUctXa0fu2OIEVFSewQLtBIB
LWTJdMHGoHg97ijnh/7v3uD0s2NUve5xbBozjvaxACPvgsVbcZbaVz5S3p/IM0C7
Y4deW2WFCVJ4AS7dBgl6tH6oN4jOL5wJeKnv9PxMZYkyKzyaHgqyB3toLvp5pgrt
f8Vrzn/8vsfYp24z+uJhO6tcSEIWNXfSlM2eygW65lgA7SiYfYLanukrhwNAiwSk
27S9+asDzYt+J1T7iYTa3mn7o9Ft4mnMfyTvQOcvv9M6zwBKpqQg0AOdyMenh0kd
ZmFaTzMhcNOgNOzIbbvKg6tJm4ddv9MvmSmjsq52Um2sgNbdCl1bpvrNbujcw8hi
NCaSH4phGUMjXIgpQtGUHrPPfSa6ban7TLUB8car/jNCCrUJaVuPTVJKgOuWs/jL
8bLt3X/D6umPpfiPLYY96ExekdCT/CGvWNVBtPkd4qOT0NDL1LUVmcBruZRE4atc
3wH+RCcC6dd+5EGyj8iDIfzvnWjLduMy/FRNmUIs47/J1cS1RtqgLklVxhS5YqtM
WfPj6Wez334y4fqe1KvV/wFHF7LMzDNZKeH1Wawc3mS8qoPfyfo4kPIAz6Y4Y5JV
f9+B1l1LXA0guePzs1lHK1tQ3+72/JAK6VWXlsXr/0ZrljL328gCg0RRXGAYNRo+
/2xLEQSnyrVd2fDbuwusXkUY1qdiixLVBUFycEfw50WWdB7PG6iAh+uBHSkYVa30
EMt8Jpt3i55vNwnvLzK9Kjh0ieeqJzdSRENbXeviCoXcaHpNRlfnk0aEUB9U1CeP
h+y5+EFkTXj6rnX7VrELqF6jxFD8A5tKsSCunDHOq1iYwSkru4kr4cOOZvLbFKRb
ikei3AfvYa/oL/HGdVHO5n99QiAZEUEP3wouY+sWhk49iQYiPHfYRfii1KWpJYJo
u7ce6wlYVRPvga/q/rfacEn5WgZ+8vyjwyTG8VxgMb2jj7txY+RZCnEJxTHrjFLd
PhIDnz4UWyzhVSKME8beJxYw5Ta+dZkMG+dX/y5TqTVXTARMTpxHaPr98UAJEuMT
p9JGUCjUx59DC/+lHkUAkiHS6dNdsYmbMgJOY6GakKMfZohBYW9fPKFZcx8tGNuH
9SPi6XB5Xau9vW4fA0vdVPQHDVwroL+KIjGGrDvPs2hlyyWTjSp+jXK0CAPx10oC
EZFs18cqOdxSobbzWxTci6B/sER71Uu/Im6B96/9SzoSSI0R+jwkMx1YyQIrTEnD
4xr5UZxadbPQGO3dsp623XX5V6sD87MnOfLDyH/2GwQYH7Lwo7fQ5xQX3t8lawjW
JINyTQOsBG1T8ZAd1h298mKB6eU846UKy3rHMAleHq9fuPpX5UClxgyWNh3rmJhq
UzluOOed90D4ZD2+rjLoqfSDkuYc0bB7UlLQYzkbz/jMw17jCkM/L9EMshVC8fkE
CCx4Ovi8HktRmp7dFkwRj9xdlWP0Wswr/eZe9/erffMaboMSLnLH+aU1RYPf+W+3
TbyMJJ189tKjPgo5eN5rY0Az/YRhInROfNfddiJBWpTjFrlDoNI0QhFQ5vjb2P4D
5VKQtRgKz8mhNh7kwKAmYiwrEYHhFwdm/f8GE2n2O0sWYd3318QPFMYp2xOmxhOs
TpweGqG9+wFoH4ekJ5mDtZpd4VihH1/0DrUsBQufIVu+VOxZCxxxv29R2lVpjuIU
WKuaaMDs5oJqJvgZiexbbJZFz83gqsviCrGNDd9J59wYCHBZ+B7geGIlwfmwiXDU
fDeacBA9nZIx4lhres4ZV0XgAimAgIhk02VCMnXAsaIg/dEDAmzE3QynOlPTKc47
iarALx7B3EVFFd0Ix5xaLjSr2b96Du43b213vqU7xghrSa0+A3v9gfn1PFDeF+C7
GwGjrV6NYxnkxB8y7ndKR/GzWzT4g8PluG47SgbeiYslUKKvniD/yevEKla4SJWV
pZJ1pQdF4m4BbKl9GWN1VXfCoMbj+VzkkxRZBci4PL9Y0SpyIHo6QjvFlbZI5sLe
TVw09xDqhZcb/WOzHoBodliaPpjQmDMedyhl6EB40cQFxVSIe2EM04kc2BZHhXpX
WGRDXPhrpkW9gUs23l/fqqiRwAEfEQfhQnzjsA9QDlvR1a0k2xlZxlKTKurQFBJX
NzTOy2x2aBnZW/afQNe5IvzIa/YgpDpTwPaBK2QwI1ikhlxd8u0EiL1Mxjahw/fx
WQN6RUW1SnHu/oJoDzOa/ww35foBIQr2YYPXgk1ltLbStMYURbl8Th0fCV+5X4v2
HdW1ywAbqFhXADwn8QDy7LnTC9/TZVUwuMZ/5265S18I99qyG7QpXh1nGjh9f8aO
W04DKcFUERa/05la1cG1/nQFKRbTjXBk4aJyROx1CL3+nJ6T5v+vFdMqrdcrxR1w
M7LUVYoB2UPKr8h/qfnsN1BoSCly38myNCP7Us/znFLU96/2O6qc0pUGntEWx5AH
bGfRWObMHXlQgmMlo4CawVbHxnSTRcdIOlOlJDfhuUoUQaR3oiPEZE87vsiwfV2J
MM5vWCQUKG73k+NMeKLGFOe9sa6COpJLFauf8ImpPZJpq0KEBc69zWvMbqemevL5
wZ1rJLeE/nlXyPwnR7/3O2qcipX4qxI2MObDmnxA84otRFJ3Gda7i8Fq1bJtB2sm
2bgtSAgJokGtR/DijHA7dgbe3ZpkV1tia1llvaecauatae9y0AO8p3Bxz4fLMnKU
FXT5jF/Ov+ssddswrFLOQ+1enMcuKmw5Mi3FCf2fj5HPgDJWphz/5weGrE6H5ARz
kJ0LPQa9E5GcfRujzM/N65Ss2Bv+tfV7ALgSiz9ytPJAn/LI0uBrqRR7K76COQ2g
FkFPzFU7x0O8vTEHapfYU7TfECMQKEuZbknkKwG/H+oI7fWhSuQgV1MRntamFB0X
DggNwn9+h590EmE/sBr5pRNHRsvi10vagvEFtrTaRmiHl9cOFNign1gqgYLaObzi
FbflC0VwMdE0U0BYpn3XBrlZl/xz9Kx0JFhkBwp2vwrfU+ZFNpjPsNZrwWSaSfsC
ap0aCKMUfdYgiTEMVYbvn9cByNlCJxJbI71IXQisHcQARFgUSzbPnzhr/ya4v6jd
+oeRlxqNJDopwX4+8hN/DbO+Yx69F0JBAmoj1rl65aOSBu8HncsFdEt4EJp6fP+E
UyggqlcxWefSC2bYtZxmUUntLQ1/neTP2cTK00hB9C31ab/QOtGtcbkVw6Fp7AXS
TwEcappNM4bY41ucYimJ3BbbkTBeacLgVlJ/vMztSOyJJf4ILySJV7bHH4mdK2Vp
2DWsyNXhFkUfvPTCELYEflBDShOI0lOpGnl7C8GGdCWJ16bid1WN1MtVo661XA59
N8sPWFm7vsZahwSc42LZ7ef64MryFGm/pHkK7QmuGVmRWdAs2I1EDY4DUQPdXCf+
xybolRa/PXwyT5T8ef0TV2cJ6UooWrpfDT6QR9u8mS3UIGwNOTNEA8HFFnFQQljt
FlnbM/1/nj9ZFSKdEruOjtEcoXg5bzh0BwA/24SIqwsG6MrCm1utCV7Jy3CSPzmS
esl1bclv8BUqvxGVaweTBnThXfLbvxBytobiogvxlokhAIJsqcZ0adwAO0GYtixu
MlCg+M66lkR2Mhqfz+K3pPLyqub4eLi3bCfkzZBneajDcDBoBNKzRZwdUwUvZCbs
9ATdde3Nkpgwl74a1pGG+c2NqJS4pxZQaVLuklJ7By5TY4FTL8lfHEoW2CYL64pL
CFS/LBvX+tRY/+pEqrZCiyh7e2IwDm755MHb2TXwdWElx3DtvVXOuCMF7VuS2u74
vZGMrtSxWGV7+DTmMAMcNqvL9sG5v6OqCUNkBgxkxTn84emwK5cCPUFeduG1pKaf
H9EOUD96VIHQPmjsw7Z0KYOV0u0XRewQ/1yzjuRsIxTqdgosIvo8a0rfhQzjVLr9
sfwHSqmbXKEJMni4RLdoIBbrv11JEkBX8H6qRe0bpLqGMWgNhXxV3S/FZZgqZwoC
JcOLmp4YYBa739ezI2MFKuhUh5dtyfL8pyX8tj0MxWb6lQ0pn+6IMfhEOY40V0l9
mDu399klVx9FPy3im877hSXEgLyYeH7EuyQWYrI8hsTXfxlOXqIPwb+cSvHsbWk8
flge/Dw3jphcA1aYkRyyT/Fp9SWmAsFPO0S5pT03GxdmWhE7GM3VqKcuxWIuEW38
cR69XcPK1nmHTh4N3qfpuasfiYEwpfwTP9ioQqTzBGPqnABw5SmXc5CFTUZzoDEN
HOy4g5quo0lnaucNXNFxKJl3+v8INAx5G3fx/48ddZ1WhtkrK3Unp8HTh011DeGB
JO1wamd7qWLYLl7bE7vaKiZvRQDbTBmemBshvNrrBO4oWQccfKsmM8Z86qUsCQig
h7vp3WVFXU+aYNjqlTHQTeHLOkpW83JoZuBK2HbLrvD4dcZu+DKv1gghz9O76MbW
bQqJjzqbTsrMixiNbXs44IHAhMBj0F4s7ffNpARzpabxBbfOCmivjwzzdfPCfTk4
hwGf4ytnqotqvzJdwm1WfpCSWt1+NMLU7rdSak2IqFKsaFOUkTj1VuJIgwFmPKot
rnUtjBH/iC7W8SdkgZUGoefWBFTX2jj/EQ77BapzvCkxjInJOK1mdniLMBcGgfVL
+alP+rILvel9gefO9SSvCUHSySx+ILO+5DxYHG6kZpgj4x2r63uwysKzl+J8Sxx6
EGaOb8iv131zKyQfThjIqhBVDytcOo8JVvCQzMKH74xhcbHtZYg1kqqV5/IZK9Rs
CyxbAJNHawHDbpp/30UKR64o9gUI7OdjXPL+WMbfO1hTULRw/Jxu1GbX6bsZRQqR
GSvvIfqhAie3/1IDI6+zpIeoXKNmCsIy5wIEojxuS1tMgDPe1oi8eqZSguVLI/D1
72beowRJaFWCfqaD4phQKsRToryB5p3rBe7/fhl+m4MkI/BhcX0fG47/K4TCVxss
e9RfzLptNOPGJR8UQsGBvoN8IEoFZTWYVHjCbPxVwTf1uBh22Bb+BthhVcPiaSBc
zL74C6bmt4SZ/dUls1OYxTtKOCX38QyhtenBk3gqM503Jw93jpcjYLpyZPikIRl0
0TW8NSUjxEQxh4q9xbWamkjJAT6Izel2BWCnEkvNRp/frN/tXz7fUyZAP6WiamXS
1sEl0PG8IlnlIdDp7hSd54NxFEQNrOkcxo7R6eyv+uHSig+sUHNlhED2ddlaRzyl
9hbya1pYneUd15JFtuNy1MwhJLFY6kM2WiE9SWew2+TzlblNgCBotaKQGAcX8wfo
OcCv7ecOg/B9x3xZ/7Rn4P89s3Qelzgx52E5XqQEFrF/67v3YAM48x0wBaJc0+rA
Us2XwovwPwL5yamDlu//nAGA2QBNW/Qicxq+Sxm3DY7W9zb3x6oULOd5pgI8PpuA
hzMewhpVD0xDSjrCt7en0wZVjR2swyfxjEVGvdFAO0HzgjisMJm3fzpmJ4eFY6Y+
9UaJMgkyoy6eFg41HC5eMKDSkIJohTUViFPNy90BG+FgBwfE/G92kDPvu/1+CRgd
l12jqbLRR2zAZVSIRAwKzlo81/PJQb31dKssOZXOsMjvuSS/4p4saE2Rlac5wRc5
dJIU8jVM/8vfsETdzNv4bfKHjmrORp5/y5a5Law7YA842wW56Vtr4nBp6N/E2KhF
VUj9SkxFpJhcA68QWTGw+acQp5HNGvFrz0d1cidux8V6lZCvdqecKEfoKoyHvJ9m
KTULpVKsT1UOh3nhNlK0+JoVNkwe+//2Xgms4vR1/vjR9ECN7z53pU/sSMW69F5+
XFb/OyaBgE6EqavHdOCCvFBlvacNNoTxMFiGGwU3gY/IDQpIjE0mzbTrzHBo/JAP
Epj/SIOfCMRRUCmvH5cafW9Zo9is1diYODaj/tD2HO3QJAhen2Na3HLELVu7H3Ia
xySPnXBz+HpKPJeQVPJhOvccpq+yUZfODmXcwbwLgADkQDTZK2fziXjq7Em540Ul
Qg9zqYiLPXfuwOVUEiszxWcUWxtXOu4uOKMogaRW5tXBFldMBlHFbternxVfu3pB
S3tUXWuoZQgnL5SxheL+sWjWrIELWHUTsbeBjRsxXP+AeMQJCnGn79chlS9tSvgu
rOMxwkppT3nZPcoiOOb1P2uXIFCe2s3zCIdTktnMw9WwhuugDsON2lgw1PAzOfpX
ayAATKkKsmT4lh8lSuSVbwgpqQY6gJZfvNJPRJjjGjY7lW1eX0OZyL5xWqqkv6Nr
blFGDzjlrlVe0k1o0qyzBiL4NbNikBiFtmiH7knxj49XkBwfN64Aj+f1IiTcxSEn
1OKf53SbC9IJMjtnsxa3zOjD0xpQQ0BaxbCf8ILhW/rh/Bd8JYg4vP+3slBMq4Uv
eQJ0yTGrlWMRQk6gq5spVCkKrZwb1HIFFzxUeXsvrQJBy2vacbxyHMfhZNVw777/
iIKZwwAE2Mqev3VS5H3b/F6FP0tTbPaN0QhYgUmGLByx1UF1IDce0JIis1r5vmLY
4OeO0qLGzjM3SYqk6+6yu/gN1/iYoCKKGQbJU+8lcsiJxXqPaTIyU3+sDy9h2BRo
VUJCywrLfokuZGzTIQHLzr8UMxCMjPaMGTEdsbpOm1xD/JRvJyVimPIlSmehd6Iq
wEudhnaxPV7Ul57lxxvWrmDdeTfGRAH8jEV8BN4Z+9XP/8vP25BDku4wYdvkiWK2
KAkfTFHYXjNNWE7PD5sXmNjcHOVCINgdoBvMV+5Z3BI3JQtY9+JDl6+mELxyUJ+K
y/PFz5D8YUuGxRf380Idr0ikHm+bZlZxMsCyjZk6QQ7Cz9lXf5n7z+eAw+5wd1MX
cBBu3tSzHeekr10gfMHGGW/9PCdIPCl9mVW6ylml3Vwy8R2zZUjBWJBEpkqnmpZ1
qFbUkjyEtJ0Qh9I3klgDod37k4d8BA210QN+BPnq3U4tm2c/rjEkXXiJrfCZC7bU
K/4TruQKGluQkaioOVrYCHLgxCNLmBbYumbU0DEm9QTXcs2x+iLFbKh8kmZEQlRD
5LjSoF0XpW8QsPFoJXilb6i/hZ9JozyTTonrsaQuC0n7avLpH1a7FP+hhdmFGiFT
CHzd7Ftc9IE1AxKgJtRuw51D+HsDLS3+/6laTiydYVvOR8T/pMvJ3ZVPiTQeQxBh
3yLk7doIkq6st3IqXgqvdVuuHkd4qfF5sLUwZ3PofqhNvQ9bepk2SMNB/WVdGU2L
dNr6jHoZzkDmLoo+Sep8E+9B7BGZXB9QJb4mQooklqLnLGdNrzrfaS5JWHk15uuF
8p6YwSa1AIYOmdv8He71JrdXkQETuOetEJRxayAEx70TDgWa5ONQjiPB3aaK5laq
0Yk9uG2/kOfdg9fwWni53DavWV2Qm4adJxjIO7hLN7OTu9ZspvlFishIj26B/GIh
5EBh7N9RgYgLs1VUVKUCL4BFxYzo8ma7QhZRBIfvFG0c9q3aiwLup6C9wPktY1xP
W5KZa/v+5I2kfVZRZhg+1ozif0bmeYM2YhkillmztVh0ilZuoJwMauNwFQgq0PSi
WWa5AOooQVvBpdgrsJWJWugH/JYPineI8NlmTNAl3pvdR0en2TQcz8MQlrgsW3WA
lEMGS9ojSa6gCksfEILsaNXehCherbxGHdswGlLXPp6CeulNMyyNXu+zplUZp6CE
WKYBgx7fJgNBcYGC/aAe6vemJQ2WqRzuo5nYJAVJNNGm1/Hmkpw+nkgMfaqYdRuY
n7cMUonJQZHnRyl6pQocEhxfSPqAZeVFk58K8cDZIq7E+01364D9l2e4MPXx0glu
OpUKyzgGljQ9wJZxhsrUFkvf16Id1niYwxDxRXCtPbJGt4KeHunB7mV+7mWT2a3t
63F/UByKAKaL9PP448tf9qx0itPNVzJumXYgjd0alnBeKVk1C8G1CFufVRH11iSZ
cJ6azNj7fxEtJ7+rfXJekvOp5UpVUQesNhXAhumqnH3j+L1j8aT/nDvH8EIgC1DV
fnyfpweIgQW5Xi6pDvmoKOkdvEZPF48jvRFNIlsyXjJskZdbCxWxAp+kvmOIzx6o
1LZa6ORnYy12v2eBKLu9NFE0Qw6UNcEaY2B9bfJ0osF9e+acTCiQCyoZW+zFmLoy
qaYiiwHsFPQuyf7DU+cm4ynsvlitD3bu9YYJdYXmwCwWiv7MAeb/J/tcEFrxJJyQ
1G5B/4cR1B33NJXGiAIo7uQMuFfjnwGHgl/lSYwFubrfs1204XTfC7vPzubWTgYu
KO9PvHKye0LVoTryVoXzc8UCn1ZuoAaeSgSp4j6QboOvvF27gQMqc81J9o4JrI0J
k3ONHkEZ1PNE0SOvg2yNI28aQN0s9SRpsHNFSZ06b83eJWhjWVaLtuxISqBjKeaT
hWrSlYbClFypwaiqynrlJ3DcyvGjIzEWSI5eTHl4rqPPdIPCzIwtoH+fRyurkhF9
s8107cg8BH8diA3c9KKYHOhOICBl/etxyKGwCk5kfeJ/5L5yJ6IlATShGSP41XEB
UzX4ORXdeGtivZvHadHRN0h2794ULvh/eichdXHeZPWyz3iP+1B3mYNbMeOFfFLO
x5p/R4C2tI4Rd+qpXlPZZ96PIjTCVaJM9nXSm2VhqKEcPU+CsWr3rhnr9aCFGyW2
pKpHJLDkuGKrW6TVhZzjpRUwx7wlP4vjFi0fx1z//s+1AJ3R5pyD31OckI4eBK6Y
oOSniE8lZAs+IxIFDtxbkDoeKGzijTkS9gctkVO5vZV+D2SkEedtFhcbAXsQvQPm
Tn71sRSa5UOXSOE/+xVwPwRTGv66vBrbASPJbEhqDvECgOPM76tYJx4tvDmPibBG
QP7WzpbE7Y42DUn09TkX8yktF9xW/vwOOvCQadXCifPROgMYShyFbalB+3P6gjcK
aFtLLfefQY50nlqCZDUX955vZdiJY4E+hhXKal3paa00ZuosNv13GWwrz0Ik79QW
ffvk+QUu4g9245fc9ni+XrlM2kpjfODQoaJQ/OlChriK6SIWLOxrIrcm3vQdhKeN
q/SNHRpUodkWmwKeZqDQCwS/7Zzz7U6VHVRANQuOlEeC3E+KEehllnBQlvWy2xCB
rsOvQqSV33BaUyejtsFZ6SnWbUH9nvXHumfR3bTFihuOOZW7NURG96IR3srQsr8X
VEZCZypQCNvD6GmkGL6QsKu+chUV353HphZ/A7H2LD8MmjpQm75av9v/TvJSpxPt
qjG+T1nwMIgdkXB+s1JsHIMOjZHIbQRp66I9yCALbCZHqEeL3TMjkoNBhx7k5EMS
Oo/3cg52f8ryL7MqecvwS05oc4Ex9jH4wTZ2ENLwteQFW2aaR7LuRRcGEVwMwn/4
Z/amKfFMXAzzrp7oWIwEwt58JrQlP6xDtwzJ6HdaFNAnO3Xcc0cvDqowjZ/2U1ya
qgLNKq2xr2WDUQmaBVxl1alUfnM8tYtE7FblW7IERi9fO3XxyXrh8xpO5J8o1rP7
7VrlgppBeai0dMgqb1+pkYiB6jJiFke/LKTvsXSqdmBWwLaqURCDVkeo61fnx9U8
MG1TLLFtSNorMzE3FDI+5p4xT4JCv5LreTHJHlzFwDSZWkY4g1Pm9uu3oFF1sDZw
Pn1qiQb+mSWpVPzpK1fqB9OTesIp0A/pGexuuJWT6Yju0oow4FSQow9goonM+W40
Pri+Wq+I+VPRu6hWFR8j4J82TFpQ8uy5N4G2MkrgaSBancgX+jTibZ6EblYmYbOQ
S4GU7dWLMTchE1Eyv8K0rKVthkGHOwZ4x6eB2fccwibUc+Rn+AGJbpI/Vaz7vVxj
Mc1ARByS2kh3DyT8g9J+0TusWu6ByZEkb6wQ3JfFSzxgusAxB9qPjO3mvmsJxetH
uX9io32ZHIc4Gv7h/enIWtAH8+e73z06RpzJ2OBYYhOiRgD2d3O9V3qsVUWc3Um0
+Wi0m+BDHjv9MuQueCctJEfT1Tv/uKK8obNhmsB/sQ5M60EnkXeeEC1KCBqcY6C2
l87p+ZuwK2wIaZ/iZ+neis4ibF5D8XEtICwGtrSlDCjacFVxb2MDzpKEL56r9cRM
deKXooacgnNh18S+BPeBNdr7hX+6/ICDrSgOD45pDbrA4q0IIewLn6A8xBZWnnOT
pSflaUJAZr+5nSsG2bPIrWGfnMFuZwHGKhzFOyXK3SjlGtJKVe81Gj/d+f816jtO
eSQ78G+x51QEwe0AfweQKexUSgxgPEla8MAsIdAtLZOog4f0iyJv5eHSwNoCdnKU
jEC2YA1/acLzDPPxbdCzGR1J/r2YZxdiDc9rzAd/CeDq4gDkY7d/AV2w+AkwbEBm
5q9CSBxd80Dho57Sb5HCY8ndFKkL086Rw/vAEBcBwkZ1pfxEIaVc7gMQW7Kap7/d
f5d9oeNA0sCcf/ButID+jHocRxGuuLTAXdUpKyG0z0Gz4Ri9yt9QfXsk248uoKXM
vZtt7T9k0Q7HQ3nwlAmAk1LZ4sigFsfMhocq0iDK3VE5408ZjVWwsM9OvaIKYZJI
lD2OcXBNhEJbYKkp6bp1fA97/vgB/DFC11csO4aud3atsZ9W3Kp40WSQ2YY8prQ7
iefmomRL0WZH6sqG3C1mCQZODOyePhs2mlpSSfIDn3pEHfm78PBOg9337Gesm+oG
T+5yPXrRknTRS5PGu4IoPOF8gl3emfLDO44kKASSOdqa0j+xNBsoWnFoWgdgTcT7
ImXZLPcue/BgdDZRNRicZTvvaEVB/fs1N8iaSCyCeoTMQ0i0MBG8q8bltHosLKgT
/zadVnjkLXSTk1ClSb0Dn07HZuSeio1PWTNIKt967iauUrC+7VoeH5THlvFeAONV
zpruynnJebuXSjyAZ8/i5xJCFFacmooZUJcxCvjii/kg4xPZCgsqdDWRWBPjxWsY
4xsoPqAj8/cg5tjjRCRRGnicz0OsKC07j6rauhdyVwBd90te1zGMJMmqi3X/Q9qe
RA/QJR3kWtS2Zit9KuootBim3Gmv/TpIcPAbmoMWzrjYFKA6pE25f2t8QCq7SK6M
6UamAzfe6e/EUgP3u8NNIm8RgBnJMzIeYp07YsHiofDAyTyuoshaS0E3xLdumYD3
HT0cvkE2j3c0saqTbdnpM+k5EK0QJG4na4d30buppF1+Kh/Dop6Yh6h89pmQmn48
VUN5bfQXE+mTsD4Q45cY2aeNc6bfAQzCjwJeGJfNH/ZJ2ldOnHo9iYc+TgTvrqdl
Zr/Wz1WcdDZdxSHwU/vlamGssGKC+PO7lo793szyVpzxAPH1MyNCaJpD+OHVBL47
rxPfEq0mSUiqZxzpYkyQm/9QMo5lDO4FiwBxZFIswBKeS+jVGaD4GYkCmvjYTaan
b1gXb6h00RMIeibjlc3ZvtOb28NJYEwF3o8rED0ePAfGLsmdchlQvrGWKnlcnBjM
vZMQbS4UGiV87CbehbTBIwoYqPSQ1zuoqr2xhdofY715n9bmRRMY66Rx3FKgs3Ur
NHSbqdmW9fXrJlJEx52melhfa2Mrj3mZfOy9PrGHp5SHFgtP3cYjeOZP+aYFwX8y
62yEc/dFw2RQWw8u9jFbEqOX0g0wlWAOJYRYcvJqFVMP6EQ14Lr/FN8S1eV2vhRf
eiAjRVq52Kfmuj2eOyr4tifj4VEy3DburV5o3J/czRCW9SYWBtbTQqgTVHNEhUwb
IW5y2JQpAvwCFaMUbcptvf3QSr+aB//pbT+9gUvO5O3eGIUfJLTGzTkwPS7x4wnk
T76G7gg0TZQ0y3MTeigIiGRQCMk5KB1ZOL+GvzNu434fbbdnA9aqjxttM3pFPI5d
FJPLRhz6srMFDFtj+y2rzc9UIa22pC1S9xXFbNYZZP2lgJKPRq9k/oYzral13s8G
LYeAebZlfrkFpunfoiUeG8uRcnNwr+ig1MSwmDU0leirG9H5akgZMB3LsK/RwsAG
BDXS1nA1DNQ4mYcHkGh3Il8gYOhEtifLUdS436lIxz6+W07malRODo3NlD5JzPZG
s0Vz8NqF3b6TAW+0/eS5EdoKnHiT/jo7oMvVpBCohGfxqukB0ko892MeJDiM81bo
9Srl6H5RZQ+X936B1qnaLTOsI0cMrhxVXCGL2Q/40JPbTn32Jpwhjwv63cjQ58D6
T7tSX9PBBGEfTQR2NHHwvzRgOOSF+jJguPA7KBil1sYdYjf+99WimZE+W7FQfpqM
Kl4+ffMkqqLV/OBOOhaEZ/wdGmWRSVOB8xvtRqgD0ic6cE5yuXX+t+xRLOYTiJxd
StjY6O3aKprJNYiy7oe7USQnwVaWry5YcajBDaldMWb/I4qinc4nECnGbc2X66ua
hCC/pxKYUmHHcgZ/0oYNq0x9RoM8qyA3sgFcw/BVeYKamuYjGfUnwG/vqzxljYFM
kplMVpvI0Q0UXLwTWAuUb95p3+mQkH1Ds80i4tj8vxpI67w3Hcf0IF9A0ztWfumx
cFNSnVk+KAneCosobGe3hpbBUMMJm8PtktmCpKZwQYAMX6BWLwVjrYJV8zo9TQeB
DXcy+5Z8vjwOM7p6hfVZmNa60mdqtKFsegBEtfCXQZ/3DYESQlY22An+VrPrp99B
goxZuvSx2heoGAcrjrONJ+Tfl52Hre85eiS2mixiDMTuJb/2JquU8UsmWuJ4kGMX
NkJaPSnvixyd3z0E+GHWFfXJB3HNsVFQyO5S+u6FSsttQm+/izxSX65h1iy3Q035
Gf6jEtGMM42ToCtTcdFbGzUHWJyRcNQADQNNuplUgIHMR+6VQx1M+Wyd4fJEjIGY
lgwbAxKFvinbks93xsQsZ5KWnObZk0pW2UuN4zkrzgEoB05UX30Z0bPmfDkQt/fs
RMB7zUWNcxWuWG+aJ8nn3iSHAJXsat+/W9vj9MG8SCxEpOUJkzwU35LcWlW4SzbH
JXxxtl9kMloEWLEhF2ceLpmeWcEUF1CRRtGNYGQim7rKwwWF7ySiLZ/fCcG9Ozjb
6wn3T2UshnDI1KMELqjE2DRxuenCSj2109zbUluUtwQiFnNFFeI9QC+F0ZJohMSe
hl7Cv85uK5boMqd46TCxAXN0BY14V3Arb6guwEzMP/OcT+vycArwYBZu8vSPUxrl
jZjwfB5Zf1hgTV8JFjbIIl/KCZf06WUMlMKBQpwa8Kc/0B6my9TmB94Z5M4N06bM
jeopCM2//YYtXIufb4J6Wlu6W6um03tW+NUWmGN9qOKfyWqQTVouW5u1mePI7uQi
wFm83ATf+DR13AVCR+GStcGfuyIbb0L24SbI0mX3V+UuINPZ3uf89Yjjpm502VsJ
5DyAwphRioryh1pMic5h6V8EJjUBqYH3WW8Tm5lw9eRTSAR5KPGQgyN6EeY59n+H
7LF1/HKDAdpgE4tt/eP9OrY6pdzxZeIouI4qpsogtdAk+5208jJP+UgcXoTp/gLb
l2we0NMaz5X7LoLYO9P5j+rCzSPF02cXoUGcfD//TOVYgoIx+vu3A2dpaLq8nzw5
Fzko5XCiz4xzSM6jz5JnKv42lLuBUgv4R3TiGPDgDbrm8EydN40hpBM3k0OkWa7d
NbLpFMxy+ZR+shk0Y3jS+TTYlQcF+7RzUs/GaFk6G0ipQjPHnF+6nS/WSlHJJNT+
sH+pKIvvcs+P9WwTXuo3WBbbx0HjV65nwltuQDR3IXoUiRGEqjDJbytqTolcPRxh
WlqZNZnyyjqXLQF8PG9jqYHuHtH0yirlRffqWdnR+Lm0izaYG/IzV7lT8O6lrfBb
IZW/JTprP4LRSKxPTv5NUGwshA1OrJUMOrNNVKWeUp6LlITpsP+xEJSRWbLUbtsA
BUCFQqOJQBc3rByg2gAAV42iy+skpBp36ourGOPZHNpE0g7TEn8Xcbjo59zxOfJw
kcM0e/NsDakOODXwI55ZYn6KUCe15Ot++BbUXVAfqTEz2q+KtW7gsVKdPtyj8cgb
hjTj4gI0bff6KNPUEiRQi56vEedRCsH3ScxowwxnUHUc1Aw2u/HAHHG3fXI5JrNd
4YtyFC4OkaAl3BKLdVUEIvEKfouVUY6+VCp6HJEC/ms5uRISmvO77xNVbfgcHLGl
CaRIYBwD6qn3Co3ZI0ufdaIVKNLzLWZYWANpIdcF4UJIKFqgzmGpS/VnwsfyOXVK
aqeuDRCpbv27nJOl6iGB5uLjIuUvdxS2dfeaOMlD41aq2xFXeWI/nbq9I5UflOyW
fxL/CzZsQDSOJ9OZhKX5DnKLNj/2Jz7raYCjvjavqJ4EIWL1pMwnMkXUrPNcX7cc
nZJtGaoLV6gmheQ3wUCRNdHUN73FrUTJTU3BigYXQ+VY9kZ767LoMLyzEFnxnfGX
MgTWuxvvLj3PHbSfuro0+LXagzo1Z8/45zTd67DHJWgA3dI5kJaV4MMBzmozHXlT
UsKCLMuO8W/bN/WPlDXenBylqVUi8jykUw9K3+PEgmcvYYpqvXXeMk/l5zy6eIZp
e9yN8VvwwqzaHei3q4oe/8aNYiDUQuxmzUZFaRZahvL7LAB8R4RNbFrrw38DWGgK
XKV/0f9YpU9WSFBbEr33lqi/ZyFqRKIk+nhQ9grlajs47SxpbQ0JBHdPug/Mx+Vx
sxf3FPjjOqx5z9zCOHpdQOiUG6ebyEHgx0JsO6EcKxtuqhPggkj/bhb8waa2vwpV
iLgosefg2Y7SZVfcCyEA91ZBNWPVnyvdJBtBOgc6o0F7vQoE2jnFNmDmaHd5vrft
3SCThYK3QOMCuZRb0oUVDGs+ejWwRnNXTnlUWbNDozWYbCSSyi1LytTW26vkgb5L
o6q3BaI+dgtYBPjJJes1xF458jnqo/FZGKp0cNsk+NlKovsp619ZjeC+BS5hR2eR
ksmXB3SAkkHx792JBjhMD5WDoMugQQQxwijBNSM2H711KIV6P5k52Png5jFJ8WxR
6H4LEDradH8L1b8AJwytPNRaBDAEO95bmDqDAIk0guxLTFP+lJrEXIY3jsxZHaa/
iwhI0SJRFuwVFn7LsNi/Ar6IPN99MUeJIoI7oBQbMWkWL4Do7/ys14gSbMNHZlOq
S4q6U3aXIDyxRMh3c0qGGGUsEP/8zv+EhDyhzlFmyESp+NK/Kg32aOlUmc2ftmGG
/Tqmshcbufs6XMPkY/kgY0TERwgsA2TcRtqzOmOpCvS1KKtCQQ89jS5FLtauWsDB
aehm+4yvysFGVRwC8K5k75dwYCcl5qOFzhrokvcmiOhIg56QgPhor2fcyylhZtAt
YZaTfWGyhv+yb2G+kHz6DRRzNJlz0kz1vMMxYYoJTf6+Cu464bax3gwy9vzxB7jV
TlC2+sX7UuL4XIZ+d0gU+fbWYRFKI0Rxy/Bl+7lbP+9BQ/d2nRz/l2vtk7bCpZqJ
68CWPekZ8T7pqAiHi2he0douyEbcrOgKTzoQToO74YM+2lRxwAz4heysGQ0r2gGX
08rQ+fhbJGUGP0l5G8mHgjLHkxZJdHoeZeyHifOxKDBN0Tq9iapfpXQP3BVTeutF
iqsAgzk5hOd+REm/KQfhfNW2cWpCx9vMvFfavtdaNpd4Z9VGRX7NTkhGmP32d/C9
cRzYn+m6TWQtaasA9mtNkROPYMuSFmELyLKrB1V/C6C+PPkz77+bQdw3YdSbmKrI
4OADQtk/7EA9Umq7RaXFFCN7CFfeeLKz2tb8JOx74L0LCzVrynNminguoy82DBJ+
Ma2FLqJkCIfolCaF6W5jfTvdCS9ibDCHm38o0excMlKs7YdFdVgBBT8qB2J+TeUa
MSp9KbABkb9Kq30nU6YptUmP65Ditf8/Bwi1dpSbpWnSyx7n8COUAAxzsd7HBas6
6OoTfa6uA18c6fzgvRSMnYZUA4hnCQ9uSt/TJrfxN4fck3rWF1SgDrI8Vw+ekgN3
bT8LeoCPksMycjNUhn0ebJti0xXY3Z5qLo4KlAHgoEkUaLEBjM7gPHXS1lTOVI7r
N7QBejHVs2jlesPZuGzW+nNS7n1otMcsHEzoifUEhNyqkR4z7gzq85N+FOyjiPb+
zavDIDT9qpuoOrENEJsD/qT1ShQyzksb4ZHSr57QnvhzD0RimXtnHg77/iltGVxX
S0zA8by/idLqJuM9HAhyAdRNptUcIHtJItzvIuQTfFHS9aWfGq/SSuB1WoymQh4y
8FN7I71ATq20I6MgQ8v3CVYodxCOV6po6epInC9osamlm5bw+58URhgcfomry9gw
bciMF/Kep28MiLlgW6h+rjgCoCHx4IXQ2LCUsEAg+Ieemm/5tmI8PPqb4PkvQ4PY
OiqNlFspONnLqNDHhb+fVDgUUk4MmDWKW/Pd7vAHs0CNemG+Bj9x4EZStl8BQsaZ
nFKp7plGulPUdf+Nf7/WlddbdFwtByCPp+Fi8UBU47ZTBr6RpjCLGyDb1PAOw+aZ
l8p8z/lxNgCE8bu6HYbw6jlxxe/hKG77hveq3w49ZD5AwaOcTF9dRk5SISQ2FdCt
Ty9+MdGy8pG+k53V8XLxxai1r2MLHOD/H609BjBBFy5wJq6/b/Thu2AgWrkRXg7F
Mi1NeN4tVkwhTZ9DqOWZ+y1zZ6naSNn2P95YgwgKOD0cYpW2Ey15bvDr12+87oix
TbfrcVl5CWB6PX8XQplbrys4oj3/qEXsUlx1yHpddcMS5jkLYwhVvyCDd7cNv3df
aNMATYtxtJCWMKOVm8pZgHWeKIKVWUxBqq5hyNnUqWj1qeWsRPBKASLDhLMr5e0D
Ba7pNYBSTmhzzWosPgtHRzGjOFNH6Kai0hnh1foOOXEwVH3TkmfYWULU6AgWe3hp
QXGAbQH8z5nPvMLLkQvypP+SvKpM4woEMUhZxwYrgV/CBPNFk6tRulhrm5Ujp50p
Xrux2i44V7iOgNe8W7DRRCuJAa+8rmNB9qDhPOMQqG5OCF198wlNkrGnDsdW5lQw
mvMcjSOhMsJ4zFO92Y1VpOd+PXNeYhsUOX/j0Jf9paksLxkwSt1Nt41X444Wdbcm
j6yVei8JG39XwOzH79mxrnjXYcXwX6wo2g7mxStO8fpABK0i/5A2urUBCZwOQLAM
15aos8ujT037RaaT8lO/PhayPcYC2cekKaDgczJ4N2/7uGWTqwLMEtQzjf/PbAcA
OVmh8TseIilFV0F1kA0ntXfKl8b8RCY4zV31Z2tW6dYfkn33ZFrw0ufBGZwDh8at
Tf6Q5O3P4IAPK/vaGIK2RwBB2LoL7PB56GfgLNuf9OsEl9x8d30nsXM2utbdPweX
HIXbXfxG9chtGbvHJiMroD5TeElectWgR81EHBkI+j8BFb56i0XlFug2IkB62y+r
Ui5Tc41lKCbUHpdcofUmkZLljUA8tHlp3M7r3T9TL+o3+Y6/JtHbWXLg4yB9VbvZ
mo786htDSxLRWMEQK+7vqmD/CruEdSipY8xRDj6PBQSQD3cm5o784v4FT56IFl8u
k4J43sfJcYi9B1D9Qovfl/vsstJXkGpMGs8t9EML+mWvZ2ZfhiDKBzMkQvQwXYDY
VE5NcWhu6db4w2tvKaXA+cOitnL3ogtd8hsOlrmPAESIB30bwCQAwGorwqbapqDl
lgp2Ikuk1Aw0vROM7Jt1PjmOUB9BZ5VVNA5Erdm95o66GTtMcga2pup4bjaCl7TS
g6WuWNwCUcqFbMS7CeSAxGofkcW7xfa6lHUGP9yu5gtMze8pJEJ7RY6wsuzGAxDj
GGuI32bPDFXIUMAAFe7MYbMvhsMEMP2Pz8X+EKAEs4HIkWS4xl0tKPv0f8G6P2Bk
10GMwGMlw8cZqeZjj8ThgvXU4T4lPJq19y6ens/ZtMnounBFl/3upzQLQzo/FOgk
eTmIc0IFPlokkL/LXetKx/ZXvq4bup8t4oQzhngjxVHfNqDNuNFyXbAmFbABbWmn
U1RozzAXDqCOOsNvadGYe6qmrS2iGyTAQu9n28SE6ldlZhJtKGbyRB0B/9NkJPD2
S+bD9J/HSFl9F0JY9OBpuL3hBOcni5ZGXsYBweD44kGkFbnK+1Cq4w8KLN1inrq2
g4TGOlnkvWgg4d8EfeQspq1LctX/IaFBxlofxXxaeN3mACOyYHEnPAoOADdczE7d
8tDgBqddSRPjJGHLV7u/NQMobM/wfyQ/rOt1ixhLDJ6Uh4GVs2LJyO6nin12xVqO
KA7ob2tlL/qa08FtGfS5UTI8tmixv1RGL6j4Z2RMpOTmZVmlmuqKA4ldOQ/KHHNu
QMsGKVSc1kdEaH5gcejV8EpXrUZgtGgfBzzfK+UjLYcYb4LKlxDFN2gsCbqZ1INe
GkQIZwj8xrHcd0cYv5nK81gDHSOs2PbaLYFlUwXtc434T0P7KX94sIu0HT0WAVan
C45zB++/PqXgaXStNugAsTVT8MFXhiu+wzipJL8fB/EEwqvDYaQGlmrWOb6Gbuj4
EMTDUAccoaknmD9hno2WEmXsHI7SMgz+GYwzPu0KCAc3q1/GyVdbemUFz4c4xMUS
ku3McVulZdisbOcy+9LtUOxjW5jJuFMW8A9jqWkqGj8M+OeIP/uusgQ3n/DMgd1q
gqXzVCOmOBY4Zyf+hhJrDPTyu2Q9FQDfgPV3a5t2z2NCI1DLvzpQJAOGCHoaY5yi
m4em/TL1oy1ET1X+cKbq6Ve+tttHkUJvm6XrDkOzgLyjCxv+/2f0ZLY/L08Riq7z
848aMdRYx7gan9VpV2sLS3LUJBHLDl5XYjj9bmT22upCBJM8drP/mj6d7FBRJfOz
Svh4D7T33w2Yqx+7eTeQ9RuA8GVGG6tUhLXNDbbFPBaddYQh1nTGgG8gQ3UrTsNs
GeJe6qSbh2hsvmPvvH+xSrQZBAuqBdwNvsZY7pmKKPAZhzR88HdFKdO5bi2+WC+j
ZGLrR41k0exomRqoRCP5IoC7XEt9zjinCM22TdgnDkRg6EPUD19cUtiwwWJeXlxl
glQ0cej5luTkyWmS5xjH7Md4bBqQLusOlmG+nl6WvzO/I++3LJuu/nNYoRVOB/nS
+ZKjCf6+yw/lNRZTqLDjRiseALQXKLLQfq5XmxZU+xlPZHaEXS7RDiXr4tkB+IoQ
OEZnM9OItrk8doyQ5l4I39ByS6Q86GhL/DoPpxyGrdiL/Qe/KljcrSQLu6AuDXo1
0BCvQARKEvjIowfOJTgO8sg6EWqdQp+O2ZrGLfd+l1+ROuuJbj7gMM4KLI4RwVKM
WwO+ZQhg89Abda7roXCaX3Eqbbc37Gu7ghvLkEpt14h4yRiYlYSZWPC3dA2LAgqS
rypZmHc/ER/fvbpqCCbAvI1S5vOWYv870brpcoeCFg8r6U7a8/tWqlS2BNDN8A8y
vtdKKGqHvX76H//ik0NnfHN3C9RwfKYyQShDiwffGJhHKxeLxEfI0JFnV/Y0osxD
hTVSneU+wIWXEaxE208/x46IpMra8DrIBiLA6GalV64vBUj44ifFMGcUuwSWRc6n
qsDnYwA3iNjdB0aB06d1Ydz/ol4BnLu8TOvbt9xVuNeb+UmCwksmK9KMeMXs/kAb
kAhHC9tW+kN8/ZdmVNP9VEW1Z1LZq6pNfRo1De6qrC7C3KoKFJ+DmGYcCO0URjSx
Q8pOU3Nf9fFb4p8Svd7eh/xlHdXSX9Tb9iQtna75uPvt8HVj0b2mmjblOOsR56OI
rHyFTG7J/SJFO9Imfnoz/JLS2jCpoc23olhINbol6HBSQnT6Nvho5458l/cVjjgS
ZUe1OWQsRP3GPfVb1vzi0Rn9oUlZPA6Zq2bLnStQ2pvEGMS3chm0ZhYL5yfF6E9G
sdSQ/JoHCHn3ouM59SfOHN1f27KCIZI1yrvdf0+WY17F3Bsl1mk1k0wR2qmfCUoI
xkRoxBzvZq4j7/X+FrZyRVn2r7xFlQyTp/0nURWBVSGDaVdrZGnoW7xCX1xGB80z
8VWOXV8wiopuDsJTNhPm6OxppRL72U3YsHoup2TlgjHwmESNcioBJJ06Nn79V6Gw
+KKKCR+hc1EQbUEm9IXjjxtcVomkY/ymCdoqhZBcvOOtQTu2Begm2iTCs01QZ3ek
oiMU+7L6yYNqfdmMZtOcb8eVMaVjxt6oz8ZZthwTcZt8SwahWhMDGncOtd5/84B1
w2z+fmj2ILBkh4mUxtIIf+UEn8UnEr7k65kiNLnTXxlCKyIdFVqgDD88izkNVdwG
TPtz40vj2eLytZ22k4uwg3/SR+ZSHP5x0rCIV9i3nJv0vBIgK62WksKN5Dpf9Iwc
2gxSbKrngzd/18TJhsYc4JCHrSMFeXQHCzx6iilgnQXNJkqfVYioiqorKK7YBRHL
hTcZ/agUcYWijvdfJhu7jXWAyjeop0I8EHbUrctMVTplM4HGffia5JJXy8iJlpxR
j9JoX4aZxolTsaJ7CAfsRFbBzL+wGBwZj1pomFhkF5LCNveMSk79Kg5xwvKXhe1a
7OQ1dW8bmYkum/gr9MDy3o/f4CcmleMmJMVN77KCdSL5MSP2TZNUBt7VOq5KUhV3
i+gvZY0JRCgxJtBc0nF6dZH7Dv1+7N7933E28Kz87o4YtbApkGr6tZgUkpEQ+rad
EiiEmu7dwSau5+ZAOgWHmY6VAufXKBVPjRSZtWt9L77QHtYSq96CeScpeex19X1Z
O5MXrk0AumxJ+ry/T5E4cRsrStf50/nHYm4GZLqmJ2KRUtMomYotTTk5i6bFAqks
4pqqF2LFUlBvnBhgQUlSgXiqO4w6VACj4qpntWJmlcqR/kFX1za1MvmIwqrzpTM3
fKxOc+PBR9826JdCRI2gQ2p6FLe99+/0qgngV9xJkQCdetCgBN+8o4xwgtiF8OmV
ZKhF1ujTbSnsojz4mRmKqzasTt4vPd4jepu/IzXm0oKbzDVDDuI3PC6IxR7BX8sf
Ui2+7mQP+U3D9ceI2bgN3WZ70dt9JxWV4xCgZpCIjEl0XKtGLGwAJcGw0Fz6IEl6
LF9jOaAtCZuH++ZAzilJMmObAnCaCPcYFcHpIaY5IdTSdsEKkGKZDNSyOMlHOeM8
WO9AaI49Tdn4qBb6xv2Nl5qqttMZGlgxCrW9/uy2UD9TXYMWbcWv0UaQL9vyH48/
q/Nv7B08VzcLm0x3jQ5sJOzlSH3RCBIWzHKFe918wlCl3KifB4zDxZTB3YwGBGNb
VXIImusjBqPZfdvs0FWOiX4xztUwyPgn0GPxgMFf89m7aVjc2XZKp3BDlZqAtjv4
z+csjVlYOAWV8Fp0zZEh0xUiAfjH6niDEtHB5qa4A7axM0r9mHOdVm9Pd8E03PIF
1XTP4hXuZLr5nE/eu3PVJp9OeUkNFf3z0QtcZ2fgTznhMaqh/AJSzw+kGD2UWN1B
csPJrifj4vsHDDyAKlnTm61aEf413HTUVUlwnEbZTFm41XSq5gP2wAr1NsyJsqaM
u7jujmVq103ik0I1l/n8B6EfbRW6TNvAK9ICWRs3p528Szsu1F8mG/ha0+WWnoDK
PfAy4hk6WFfosvrX230bZ9nigumzj93VB7efhR3tJsWtG3AWLnrMZRwLKuEq8Qmr
17etq5hFV0lBpl5JK2txWkGzpUUaw1vF11X28ZOGe9anLbXf9KGaH7RjcGwhfgE2
HHPcjcB+u0V1NW4uMiHnFISaw+sdgbFZZmt03yM3Ux/jN7q9CrisZxAnQ/CFHQo6
SkUlr6j1nlos+46OjH5XH0imv4ROcWluD+1C4tVOJsEZmYID12njqVLvVzf574BF
1RQlr6yGVoOcypj6LvMH/DYu46rUHcbwzfpMhGfb5t/UvLgtJVILk0HTRdRoQLU7
/gpxw5UspOmE59PeT5uv3s7aWat6YvJmVUBkBEwKuB8tjJkWOpJq64tlW16csUKo
hVsgF0d5+hi8JezJxWL/tVCrfSF6FL1CUNS5U9qfCvUNS0eZiSKfeNGhmgJzsF4w
mOBlFFMN/2PDs57qLsV7VFMJUn6ugybHdj3SRGsr2iuZdCJDTSYdGM83e5AiR20O
UNy8drAxskHNTHFyu4Od06n4XE8Vd45NMFHBMzIyWhR7lqe4GwQ/uKJFSpxEzIMg
cSda1Bmeao/YHJ6EB5pZPQl3d5bq21sQL9NnMk61D9p50bJkPEsYedxpciiDEFmE
M8zFJZW0H+2g3oGysGbQ60jB6GdSagRjWywJbIAwIuBGJab6p325qS0zLWJNsLS3
9KILNGbp8gIaoeUlO8n3YlTG5lXaIcNlSaAwWC3v8AyOZeN8vR4BrRJskB83o+9O
usWjm8HVHltrSNBcR0M0a9Y6D0TeKhMjTT99GUDHr3aGLggjVtTkFUi7kvuvQd9m
xqy8Wdu1Sy1+FXI00YBzrMOpIns4um/+nZyUet78Oq1NJhKJTXmpFea2d3nbb8nN
JcLHHXQM92Pu6pHozcfUxhrn5VwnhEHviTFc/YUcmbn1VO+rg+lj3IPRBXnYRfhP
NqFNz/xHs3mD6vjc6SgPJq6mAN9DQ/T1xa3wYCosNM1hikNSYa90hWlsVm14obcs
on89UxvjrPE1N1xZrW/o8Jrq4oL2B9IQP6hc9EbldEgZTEoTmVgsnZ7KlaXI1L6z
khOL4QUXSgT8ZZdBOWc0M+6xYg0/GW+Q/D1DQrDZ5k4j6VlMY/AjdbTea9Kmu1In
GFFsosb+nW2IYKlNmxS9QSTrSv9VWtyHHHV76LVBBNJW1w/btbeyGi4w+6CG0N/A
sTD439HC0a645zvok4YRRw37hS0J/HHnULEmbQYi1CxK4em5o12doKtyA+9oPupZ
6MKXjp3unZeRObSZvSvsIbKinb5GHf0cF5bMFGlMBPcZ6V7tXH2r0do2qG45KPWI
pHvPJw58Kpnz7JVhWlUCcCsvR5YBwuA8Rfzv9a1QnQ8edPsC7KIEqF4w0Vv3ioxQ
f8jeXiT66KxX6+S8dseMptdJBuMoAEqHY8uV2wryczYims2Q9hP2uVfY9e1vCyHl
zMt7YQuvTvWZBlj2f+7o3ZHIej44hqjgwKo4OoAL6F58m93HvRh8rPONpwATQHx/
o5DLhsoT45E2lFT/O+pI0yjrIEG9i7NM5vjwrrMixRFCS+mv6pLwftm+Zfre8Vll
fSDKU9ScNzFvXU+nESFvEWfgxqa/ox3Ymh1FHXAeFUJLBIY+R0HD0Rr0p6+5p009
frAttCvq5jvl8uuDcuT6GLPtls9RhgSAJqjtf1uFghjZHh2gDIjgAq4W+E1uaXcM
rIBvhOcfkH2ebPNdAXQCw3f7XyUCgkGAxlsOH/L04o3/+9JcIIU7rjpHg9CD2eQi
VEDxTYIO9aORe1ZhRjQzJKb2dNwX3lj2BmOsegQPecB9oAa/92Xt/oN9WOmyVFow
HDra23C3ZNjnUQJPVdilnqlnmb1iGumess6FDJXDiq8deWSObnbc0h3r/uULwxSd
AsYmCETN+Q/kbUh8APvhzQtS2pjlmVK4xNtGzAk/FZQ+GDZ6DjVPJ5jWClWFvjoa
WUiCUbStBHC5yLTSwzkWZowDl80LVbitjMUU2At9v5Osa6datElqr45Vf+s5YmKc
dO0+aqaQ1cNexVJd4Qz4jPKTDuw5WE8IwVLZKiX9CnYg5Tn6hKkEPcrNjEfeU/j9
fJ1t5tWQkZbkEJuVP74xDeY2WznNugLdEVmC1zpHuJUaw9+kzdjd4Rw9B2ya63to
JZBEc8Z961wMkk8XPHC1t9haZMCHKcNJac15Uda+slJgGNscHWPlHua5MV4tATN7
ORHHZxtM4DZvVPWEQ2G+FjPbILjBja2XNvBzHuhMOs4wLHvSeLieV+JcLTXL7XPI
izlIT3d5+fkm8ubRDXJPPXIckl1cuuvYFS4EB+HHKgGStWKYMtlaZKNbBt6G4Ql9
kaNeXgTgoa6BpXqRUWCJwSxGCBH+ASJzxyz6vGazMg0KBAfEHAU5HY9ccrc/G6xh
KlBC95WtZCfpp35QIX/e20E7uLHUv8sm/6JvrAqueeCWbQf+Qt3v0/lsXsSuaPsG
utM486hbb7IUtsdWXUr2i89Do/W/V9BnohnT5XYPyWOLs1h9mqQsqFRSnv5wE0Jg
+MEQ4WXRPdHjvNS86ir7ErbOBsdF6l2c6TfFSc6v6V0+ziLfnGm0/nAEo+2x5iaP
MK9JePVVBtz0U73Bqo5lyqZwyC79va9+3fF5PvfbgEUM7dHJg14D8KbT0DyXw6vI
BamgivpoRlUoXD2Xe4qyf/hEQQjZsexcC79m4alGUJ6UnZm2spNj2kGhD3+KkMvv
L+12c0UlU8YoExQN6hRgVwkQRlDCiCCmhkEKh8cPJVG/mo2AAG5f5UHY7E3nReht
4Cly6N8Fmsc2rG/B1Dh+BA7+1XUR4N3mbnYyR6/rjBK3oIDocUAHv1zwIlcK7otM
glLXu9fkuf6YvLTYd3xNc2Jw2TDR/w6yoYDoFJHBoXQDKc/iIyEpZBlDnGsD8y9Q
I/vAcAYTg9sQOU4c8tHtmyrgci91bB+lSFh4Ed5bcFa3558K/VgQXdrWOFvFkB9N
GHZk/CL1z/OauiQ9idRKYkpQ/4LUUEatA1TXD4ZagDlBBKLEAsGxtWPFQikyMRyG
n+XOfgATr3FOSQmoXmmJTu0wn9PHdg6YVvjJ8cB1pSzQdpFhs4wLty7JKLWlj1ip
PLFwhH+Fy/uHp3BU2+yzgGyYityzUUpdRxJtWz8RP2oUBUCWp90o/WHjRNLEG4Rb
Rgw3gJEU9yO/dp+DfTN5QndLvySPoYQ+xtyFVQveQcAAvz6TUngm49xKvNiJCvuB
3GFzvYpQgyGiapvjjqNvF0R98iPtLbNDS9un9lHywJiKDfY5S6VlrKuhtmHBEZ8d
pzXQt9WeDqKy+GzE7GD42cVk5DLUNz2PCiattvjczaK02nGM/7940ulhhv3/DySF
GVIZcc5fSditKK6RANrbG0MP2UwXDOIQLmggRpdDpM9rSem4HcV9pVj5xW2Qkk3z
AHFcyw7mQsCQumJ5PswKb9NMTeVzdqEgsm2JzQrDbVO531of+0q3TrZZs4YOMPWv
siLq1JD7A8O0jGDncd9eErXqJ/Xu2ic6/vh8RtrmcK8VOZq3dSakdJC1PGRzlEWz
1typu32ILsLG3u5ji6+eCyRjAz1OY1xenSdYEmDp6FjC+zmYLQ8+ogG+9uQiDdbf
9wiCyjvtYkr9TzhrCvfBtRK6GLfFnROXOzSrPD5CKGMMHlFQnDR3s8/hXp6KLqtw
4FuSS7y69x3s9pZo5W+ZLvABN9h7pzQAD5br7IyRAip7fSXIzbzzLwlizbzRv8Fk
yAURlXSF1kaoB+EL+mrsi9WTimoE6y6tzkIf0p7h2HOmtTnV/XvrWFlI/XGfp1tE
fabr96eAHDEpGsKo5gdSQgTFPLkbzhHmDr4jps0o3b2BsSTtpnLtoyDk2IZj5AKd
QUpRDA76qFm6tvvL5kHIIyALvllGAWgVk/vnH0wN6Yd69Tb+8IgB/ZF+8aNb5j3b
Q4X1VBJVeRLJGD7uS9Xrw6JkunqatGbSLLGVz9QOEqaDbf7++M0yHkwp7wsRLJMF
HmunTmuGuwaMY1Aj/D7OAZ8UFkpPuS0cX2NP5qtMmmHjRs8zqhDH19WBqKrFfUD9
saSoODlAkPJ37Hlu8TW4Mh5fntKKHu8ai5SgNA5bvJUoPzkf4JUPuaeFHjq/Z5XL
AcPMxqmElPQc4F4P+74K9cv9JiKSiTnU8xltu7+qdVoriJeL74U9V13iANuOX8p5
LohnHbU8cHOYrGUhh6Feciss/jyjqIFFzy8qGw5iya+9IyEOT3TGxj8myfhGYHqw
52kpxXw7Rx3hHpTumH1Re/tBeT7UpzmTn00o12KSscGrhZ+qHvYP7AHarxbx2fIF
IDIDBUOyWTqUwxWMTodzg5YjNotOQC1pMC3glFUWGWJydq7zCnOquS7PiqIom10S
nQBNJHHy0AnyUxFu0yOmUKbOM+alB9yuWhQAOpaEMK5WKL56kJrY1+Vbb1Zuz4Fk
NKOuj7q++ZzKt08OnDLEdRk6D+4u8FNydqxv6UGGLQzb2W7X0PXDIEtLrjkTjeTC
hmpUm8cHI6YNe5jqpc4xtG7yqMFtDlbY2M7CJJY0VvEaPVyheWQv/ufDZhqaHJgp
+5naJpFSPvjLdG+NHFWM223oLmARDiJ9NrA+miruaKYfK4UcbXz4E1z5WlLgO1h1
+8KbQKLohlBLJYoZJxafa/JClkK/BxF5UZkz5/gsbvg7fIHEN44D4tEo6D0G/Hd+
Uj4QG4bkUNtVEBdGfGmQUQ0+LJ6Peb97TDdTxUXFGM6J2MkfmFO7V/vUQZWCG7lY
+jGg0QxXQvev/b5g1jr8mvHDOIFqfO3MS28kY4hmTrRw/nFe12G63CHE1HhBEkTC
rt0VEz2nEs2Y85Bh8S4tLPJ7l3k+Dyv7Z/FeT1FC8TSRdkEsMpVl/BL6rVoSMqp4
nEQ1qCzu5D/n7q0Gnyngu7mOVPJEZDqNK4dZrwCAiLJtuGhmkMaCZJwQK5UDTPs7
ClwnmoSIMJqOPJLU0EzLBENcOOnDoCMNYMyfrzc+7ig04QhS2LMa6dlKswuu13Rv
k+QnK/bRos45RexRg6sYh12iVVbSpC5SdejjQ5Vupjkk/juGDCDtNnpXlRvuMtiN
PYnUPfS7kTgeO3Tn6ij7qXVggU9CbdsxnvnLaX/CHqeYIm465tihnm12wl1jpzJn
fVxAQicc+PLVLFt8QBTt1/o7L1vQhDwSQvHjjafr6rEZDSjw+/vCEcl9NhmVnFeG
qW5rqDZ+2TB5XgCg61Kbd6fVldAemOOe27kjRtOJj9UuzoQNFucOLtB8qjHYZaxp
KvPiIRc4w6sDoMPa9avXn8aoe31FSnqwfDuWGG57Ogvz8cJBVxuvXIlb+LZvWZTa
IByeuGc4diKrnFtHgIp9TrCl7OQjp9qMcZmNrCHtM9hA7n9XEgswgMcxYnyUiWo6
ZFsI76NHo5XG+6GLPnR67v3CoVenYGP9oQSBJ4ASZgEkFmDxbPCIKdJGbtlyeXAY
N39kvPQGZj35vhj32Z7HSLGaDmO21LtpdVy6G9nUQQtCKg0BUm69MqQ/GKNrVEmO
Yc1aJlRfRimFDr5JQaoqZOPzTawQ8dXRKq2K1BKh4+G38pGKSO+4KGBOGBzY0xc/
wUPMi9F2lb1451nkQndzvqd2b/TLOVqdKXezwB06ZWYL8qehoiAmLhcdGN5eVuOl
no0goV3CVn1KkDY6MqyG8IxftNQSJViDDqkfFJLVbc+qEH+swauQGJebrzH1Lxlh
DGh0f0Vlsz1JGU+PwJPr4Vhqgxl3qwHkdS6xsjgb443IN9njZslLJ/jo0wUNASva
fPMyE8iSvrNAUxZ9aPwEFTyP4VsTxxltf6uPKAwteIrMvzUOiVKxUztYOS/Eyw7g
SuKco7I5RrCI4jmw5BAtGiyilF5Um7ttw/l5LAWxk41SRL7LoN9liWuaqsIWK4Tg
+admYKBYiJ8QPWsXdX5rdq30Vo2GexXpVFhv8Px2liTAmZ25+uiWXjcuk29xLKpV
RoAl1XxgKeu/lACpo4GR2huWInMvGy0IA+95grav7CRbLJdIGsXR16SIrmssj3qt
7IjuROfDpk4TNVTlm+pVKV21bFBACcSMyc5VgD0an2Jn5+YeXuZWFSfLnz9pWgId
ihLIFKVmYOtZvBaLt7G0D6A9AGcL1Ur4kTZPbWmS3cJXtr9OV4BwDOBrziN9F/od
lcgeAFhgCgiarLrHLmqIXRe//CCD9exsaHWsYqFPM9YDm5w4lSfwBBHXtFm9c8eW
Vz1adVgICHxKv+BpUxKh80U7B0UOday59GqKUZeA/ha/hSXXsHZN5EPzWK7vorgv
MSSgnd9NqveBVx6iQXm0Zpj/ZNcxCxeEMvaRwSlf4BBxXH8VlZWeb7+K7r/3H/r5
713nfQvCCe7n7amvidhLJY4Q8fcRYNlb1pglLXJZeOlAJiazvCamO1YJFdNZv+hp
aMGTiHXHFguEaIIoyPspXOfXVuX9V//kYIzXdnhevy6sSvQtRs5/GdOiod2Gxv2d
4RSFxGaoFzc9WuDk5cG6pW9VCEulqtr0ZE6oCW37ShWi93k3YstmzN2SJBgCdyMQ
yQbW3EQnQKq9KRuszGqsFXAryILiw1ODaOtHG7U8kxoaGhgFkbfjqG+xUZ52fg2/
Im12DBH6twwt6viBQkK/RCnFXg9LPr/HhWECZZdDqH727mcyK/IWpkZ9IUfW4Hzw
JpXZzt5fmSjL7w/npuVg/AgD22BHMEprcT8NdIZ0w1cJ505oQ3ufbYbz1/4nrqfV
UOQPTI97wO4/zItRXmSjCKYM3+Poh6qZAnUx8lZIm7vACCdKLSaKwg+yRTUmDG+4
Z3sEJA3//vrTS2n8SiFt/Xc5+r8FuZWgFJtLG2d3ydCNGDrOgTztF3wJ8+hNEp7r
aXNrA5GzQrmRC3v93mwYpt438Xzjec3cW5djfuk0UyLPSvHfrE6i80jX9edOoGBy
Xm+JSuX33RNyIXi9PVo4elYRvJZgzikO53xaEiLvLegTDyQIMTzlYMbrDsy6cGKy
mKrEdlZ4UVSEh4b16sQ04Ec9FtBr5euVX2Teq82oViY3e+Ow3JrUoPoeFzh6W9MG
/wkbpFEpXW2JJk23i5clL/TBDeJ3zD9LfOeeG0UgusM69Ap4YhO3QXKm8L5nycV9
fEFoVmlAUlhsDulJ25kTVJ9I2lfx1qLkBdA5SLixHLTBQrztGEJQO/XQuCq9rA6m
yxPJJJGPfY1XTRcUW4bmBKN1TC2WSt/2lZJj7s1FbwIbTyDoEFpdZOL18zZB5b/T
iFfSc3u3D0Yat+m1HQBw4vgV/pAtVJRwzGqtZ3cB4xFQ2FCBYwnALi2kLKKhqK/g
BvpwuGlB9f+AzwG0bW8ixb3Sk0jwtYDXuwDiIUyiaXg2abJES8seAySXwIm2bm19
y+L8JZj32mDiVPlR+Bv/gvSOXoynqVdG/12tTemSK+lH12XL8jBeikTxdthddflO
QejTQ9ps84Yosxlg8GEAXfT9rtr1KX7nt6lKdcrWOWD1ufYAt5ow/MTl5TtbGCDk
XMIxDpesjfrMz79WGdAuzE46IhzJLIAOGdwobAJK1gSh3gatxNmdrQxzL1N0j9dP
s07avD48ZDrzZMtvg6wkb0F0asas2LgLQ1c+LvGE86y0XNJ+6UpBEmoHqjBKYrhF
7KD+QYfXiTToU2gvczNxhIkn5E+YMqXkB9cx1IwvkqQl9vOetdH+5k+O0duHbIGI
BZMSHr5cvI6UoawPA3vMnr6Ay2Y2NQmDN+tLQ2WzrlqUc+F6Ak7NdXGe5G1LYIUt
4m6TfryW423e+yiTBL2Ai2Ozb3UZFNV/RGDBUgHNc37cvXLLRI/QKGSQvYtaMMWF
fwqMAO/3bp21I+BaCaHjDYCm53ctc1WgEF89Sc3A79Wgz2coEK8M+8SSjR2P4Saj
x7weMIIrwASSvbF6OC5rGqAjimXc+bZfSL2oH0yq3YerzOB+5n9LiDX4K1+hS2bx
va1qRObq0VDt81M/BOuuc1khmV6CdMKlrzy2iiyw3EnhCI/N5zhyT+UmSxDHViOt
lerMqqSR4i0amYOIlBQVHkBaPDSiEQItVoYLbAFWNIQ9Tr41SY/w+F/41BvXI7Y9
3Ab24lRlU+JHkbAOLlo1trgVxBKxfeOfIXmvEZvnuoyEra16rVvobWOn2Ry8XOJX
or55X6Inw5QVqt4IpZ17bSgBvtbs6UvHhzzDEpTcRcK6NiHbe8zbGZn6sikcQpnB
xT8GK9GhlBvNyqYjKjcOO/QcOUv9ohnhWF5X8BB08S8idb0RJuU+USmIT2je4FuK
AnJRqrpDbJbLCWQ1WIYAIthAJFSx8D2kw0UY+87AAAdNkV/7GGdHm7f1BjnGje6g
LJKPjmZDWxLkhS9+7Vp/OzoI5FbsdHIDv/5E+VO1/sT5zPLRTqd6s3XPmjSxNt1O
Xa+ihI3M1oPV1/loevUbtsGukpj6sXQEJN2pNmgAZiKKzV8ysFOsbFNrgtMTON4g
RiejD4Cah/+eLJSfmVqQrGmHgdubGoz/Wsc5KW9mxWNSwNxjhp7Xy0WPhWVibzV1
HpdgYEMZWfiermBxm13BFoSWmwFfgrTTcRvBAf7B9WyAcLTp0nhDJEmMQ3s/yfwG
2qf/gFs44GX7a7s38MkIbu73rslqikPGEygY9xlTaNxY3Yhq0xffAqCz4HLQmcJx
EBWv86LTNuO/uAhS/iLxs3BuREG9Hq2p9Fun/kZo2ZzZUXpUMF3xjHJ4CWuC8A2J
SCD+e2c4rJ5YgXfSwz7gD7MFHDQRiaYJwFIOCjQ9Y3GJu6YpxxmlqAc2c+fdI+1N
WKEKPgKfwIqQdFCYoa6XPV+R64PK4uhvw8jIukj7S2zMcF+Sqp1KqfrisS1/J2aQ
HeRagYrOVDvFjj+T2ryXYvEGTmzLlj6nd3mx3r17/l9tGtJGy3fBiWL2cT1afDIT
6FZFrOPFYSlTFAuIrzu1b6k7CejlSeI+qFyBGqilg23C5uQHUTQbVIfaSRtUhWz2
NIcmyys5ty/g1btgELlod2alYelebLSyXnn6S4F3EsK1WvsTim20j3tcR2JmEfiw
TINHRakVra0PKv8YnRlYp2vwglqH5RwsQaMXu0kp7GrzBbSyZFpmNxh30kMM/99O
Caov3i0/Y1/JdWkIXAGgBym7Xmqb+9CKT96i7gaTbXr6mZQBvxE2A7uzzlkOnxWr
TzQ9CUGmuuLLBcziQxTT7UElCwFgAOC779CqVvbZ9AAL+B7GveP5DHU07hdcoe6V
409cMdRaTkZRNncPmbdBK2kQAgHPBhpc+6FQ/XHrfdqi53omV+AsT0yYY2RAWVNf
95pJi6i+vodb7zNKTtgHegLb0QNSYHcgY1n8iHyJgfS7MA5CWub6yDed6cgj7Eeh
QgV3yU5ccmATC01rnI6TUmMGs2T7YDHVV/AR+o6U40iXrO3hT2A2ZFJUU0tkEZj3
7X6LFq3Ckf2LsoKmz3np7Y3fyEQjp4Tq+1kfoNIm3cO8Iq+jVwwZzX2vniEHuDlE
gZYsgXbCGUjEnI2MsV1iays6+9YHL/bq3SOWb3fJQGj4XfL6iU/u7IOrx3G+DoTZ
zkS9On1s1A+/SWLv2XdT0+xSFccxdLUyQeEDdILESamb22xc/MPfzf/5Uig/yyv1
mb+z/enH9uXB0byUhkh+hG8Y5882NYVjEq2ZpD9EvQoKJfwOU7rNPDnw++mC3pp9
4AJz3as9+CoEdPt00/06VUTRKVCztWdSKK1trIUfOJdARijI33JqXlPN+UznAGac
H3vFUzZqNsfBy+skYkTf88420kMppFylWrbmgngzTRfhf5RAWc52znxkv4/PKMdh
ykDyvzO+RFYVVW/3nBucFFpsS39/xd7pi4pVuzl5w7ROIXn/mnGv6d6LIGMXgsQn
C4gdKreJjMB9JjFM097evF4qyYPfxjMa/ngWqXY9JqOia1wPNQO3ea0Q32sR9XIs
hxHfclTTOfjMxCmz2R0gPuPixMSNPy+wK4Mtl45/MhU2GCeJlVxiBirpj6N7PBpB
YT9O7rVtghkuqGIJKn2TwrgJ/gnYX7W/iJLPuE7x7bbmQct3hxMhszKpZP+EtoDg
lIjwJ7eyZr24c5AyyvsnXoVpjjQsWwBzsVUl5yRPULaRi6u8CzaafCtFkJ5XItVO
HEKloDtwGFqFll2j/xe+Hexh8t9xzrtQgf1jQrvyKPkHpUiDQbrZtbpd8STRdwvj
jTcMcPBsISHZmdpRJay9f+by6g/IzYrUu3goHbkLm5u9kAr/mZwy0JsmcDsnQAQR
/fR1by8VFq1KS/DpGQKXrvhwIbum1pkVypx3X4RPB5yuPck5Ihz6AbOx9/9LcH8k
6sqWvalGxFnbh4uv73j3wZ1rJxctHVenIEsn7pcFaivxkYi6/h4n/VLcECCxl8bn
8K6MDYp9Zlb+sNUcIsYUze5ow0x/2E8qkyO8Y+etJG7Sdf8fwFogVB56/sxX4ChU
/NPsgvEWmJv2ijbG/HTQ9+PwCi0015Q0Aq0x9wdP8MaoBMrbVKJyvGZ4BlBpk9vI
g2XFQj/+FENnzB1KA71ywHahYwgUUhUzCrGhaeQv/cao2q6ZDLbfFh1zA61JIZwu
1EAmMX9fIH494Oegf8JNZK+TjBA3GxjHmrbHLXMkb1FF/L7fnwmmdr/zbzN4+m9e
vhkk0hcTJtVUoHl0WR84EHVtSybyezkcHwyORQ/kV8J2YmFCjTI86/mNHRP3TdSC
C/ubDEyqY/lI7madPPRuR0PWsSRIaHL2kK1bKllrwk5A3rUmizb2g8F3C33GaZaO
r8Eb5J+bsDpSISeYG4np75ExYO3Ikh9wdJHaDB0m3M5XsDu1/NRaFf3CNh8C7Xz1
ekH8Qj0rY8z5BZz+v2UX32TK46LTTXpStftgs9EjjbPG5dzOC+Uet8be7NDli6EQ
vrfnbQqrawHD0AVKCI+ehN+hQfRhFqb3R3Yo2ygOogmUXpulF/wzMD5VWH7g44CJ
JDrehgDJh1xss08JBVWys36SdNJoIdR/6krUqPkNlr5dG6lvRE4bm6T5leXb5J5W
yHGJxZrN198IQwQKAzO+BPwdxaEEzwppibCHKrKUVD+eHm7iDhiyuLoPZGpLaSLK
TfEII+m5IEgJDdn45hpheTEYEGq1dyjWST5mGaH8WtuZuWRUZcbYnTEGbaom3MGr
t9S519llribmsuMLV3k8+rfBtWcmwRiGQxKKpjL/mleLCDRgsw8WbeAO9hBmB0h/
621hhieYt+u1cGn93jciuV0tV1by6XKuvuffmMPGy393l9mcI2dyIft5newo2glS
muLtZNyudd6pgVxPd0+BFok1r0EP+HA9EESJPxDi+eAK1ZvdY0WFRXy1B9/Opl5N
ygYI4PQFEJnxbIUIaLvFnO47eKo10uLSEzLh9Lvf3EsnhRq/+ufJFid35c9j71SY
pfwCyy4DQAlVhwB7On2VIsBSXJ239m2NTkv0C3nwjcvi+8hx7XvHi8wI9sb6TeNj
HZl4Cboo2S6aKth/zTFiWMfoLRS67tiuK6QLZRymnBpRpDh3/eV9u8vv2HH2GzeZ
SUO+o5xGzkEgUgxtSb6VkBelw0KMAYxbP4UMzhnzdjMysWJ9yyeEhKrdYDqTxfOn
NRT4hqUeg2DWjFOyyXdXj8oB9mExGwd2x3CFSMXBYHamXBeuxHOnrBnXTFaImbBW
jeFDnL5J0c1iqN7wpykgh0OFNnAbmPYwKEI9Fgh+hqTW947lmkF+GroTizAEEMpF
O/0qNJJe/zsTj7Ig3LBmzUpI11iWYTtr835p4LUS8jVnvvN3rgAW+iVAXNpOpzM0
04msssvu5hsSYa0eoUbMmxIaLSEPk89Mj1JaKoe8lxeYB7sIQ3YwbSZH5YCg1F54
RqLTM/fiRWstsW668MbIkj/YBsjsjX2eCW7oftLodfjfp4pPcybGVwFe8Pgjb1CQ
8Q0hGdwR2exWLg715RT8wuR25779rlfmJSqJebNLpgCWIGu77TFjHqfoZprAtsRQ
Mi4LxuXNrAxlsNmAytjlAukZSKX1Zk7KMR4fkE6kt8G+TQMPaDoXMZAJBwLvMO9+
8BDCLVlcEzZFFMrstN/R8J4Ytitb1CdlyNtT9Ky1afoJ1xrKoFZwfuh+ZzRW8cpD
LpvcPCqF43Z5tlv4bjI6Lh4/xDpckP98yKq539p2wIUNcvlsqjf6yxp8vmeejxnu
W30ZX4LJaa3ny5vJVvxyoZrkStl3Hvi56vAeah5LEaWviXF2Il00fXIfZgloNsb/
HC5cSMI5HWxWxLBndmfV222UEmuV6c8XleC4vZL7P3GuLh05edzEmXQoCNnsAc51
jnu5Zpdh3DAKk3OSh/YbGW2Gy5bLrGCZl5u/CeFdF+QFeZRoydoQZq5EhMSZ6auP
Vtq46OUYDu2PkTASvuKJdvM2wRn9Z5iperWpJtzF6z7YUfTQDcq0Q1ahphmMHAyF
vMXYuIDbQyrzq4OAzMWyyH44KRSTcs8cybEZFceRPOrc35dRN1SrRSLGJrPr3hBY
L01fU51U7ol5nQEF3NQBdkHYdEN5mfpXP/bhegQGN45uefAg0Ik/5OGSrMAe0/R+
YqBbtye92SaVdnPLxcURy34q2O70rMrmeHXuZnHgXw6c0GVxSd9ePtCP+m3nwyW5
0FymcAocdG2MhUKl6vhxlTpwPMYc760XGDDRWCVNaUxdEkZUx/xBDsoqVviauPdc
UZCmLB9vp+iIUC3CVsHVICqH1h+dcnUzFZ/0iOuZ441emOtCSxyX0lL2v8oBOwB7
NCUcd9k+2SRpJmhn2SBmviO8n+jfUSvmc0No17rGdy1RYNsOYWQ89nAPwuPiszUl
Coy8YEvDlBKS6DgN4w+4MHD/CePPih21f8sIgS/CZ+KDJy+PkAE1X/4IJnnW18jy
32Sb+5q3kchLUsbS2Xn0meFc6YlHQwuyxNWxt/Ze8ZuObWCttXiUJh0AamAXvLmR
DM8rCn70y9qdsLZX1h2zVAltKzGsBHViZ7Yr+CSmZtoxKofXX3bVCyqLqHtxe22/
2InTE5++XzpYTjDsp+MLT5eqIN7MS0WwQws3MSSSkdB/vlJYyZesCM+vpqmz2TD3
/suLTI+83UqALtvPueqbJ1OAcsZ1eyCzsHxhe0YMnEnY955UcpOFYjjAD05zArMV
N3D5eEKeTlV9HO8zuvV/r/XKtYdDbkxyrAH94nxhDn8HWPvWE9i/REBr/g6JTTXW
mplgVaUNbnFBwC3+su8x7PatCY9bdRmYngn/CGJHoEJwVRRVxK9gQQ9HgOC+vwn1
VkVQFweGymGyNJCJ/+ikQD9wcgVuDAbdno91YSqvryLP8O++3Gj5y+CAFnMQFDe7
6rVvpA+vlISy3kEzdA2XDrss0ZxjW+225/Ui9SwM6gEg3Lq9FUCFuWE+EfxlhCBG
VrRUHPyTVBlqPbO39CShSUFK3G5pe1Ab34KRZOEw6xSX2qb+DGebMqXPhLt3Wy9o
a9GQuxTTBK3YU9ILRc08iBSgG2HM7PdL3zac/BW1NoUBIRi+b/kAap4LjkHvs4z5
nRCHa0f/cuQa2640mzj7kB8SOe+vAv8S/0zGevkRcEZxzOgHf/+ikn9kpvz2K6yr
jZpdwT0V+Zd9ydklizcwAsg3+/dSw2EU5HX1zgy+EaSgwRedL9VgvrlAvj8yXpj2
fBzdeMgLg0RMu+8OgyhRfJYMOxdaas8cM4iHqZAWTtqHrayKGh3Vi4y7M/V1Cly9
rGmrLdCKDz3p9AEC/9OtHzW/rO6u6hF+4CTUDqXfYbpBe05A05lHjjofNOq6SnxN
U2O1zTB/H2CYIFprtSm0WpcSGPOAFZfdZYo7ZKREwHunjG2n+0D4dG/Fl6UCbwTA
NH9pfgIsiH2KX/VUZ01qwaHrcGu0kGzG66pUWcLqSteqHNeoju8bgdFQwRIi8w7+
DXPjW6DJWiwqSFf1HaMHDBpOQmXd3fcRJBGvnzY9H63WyrBpCtcKLU8HOnOlm//d
LCpxfC7kKT2VAKu3hr5NaRJnF9srKD02mQlk6E8CwIQLuT7mTpMCiHHdyJHJFZfD
bHiiR01vR4Nz+740tiQziTiiCbZLwhGSlkIBU8Cn50dPcKhbBgH0/BXv1s9zDv7j
OenqZfUNQ/mt6t188nMF5N1FC+ajsnEwKvJ7Dpo2g5KPppBe1R8rC9A+8qBmJgiP
QhBILTRgY+Pild2+HB7pl9cJBkb3T7t9dntW/0gaTJgUnpLZP9W6JIq+PqNkBuxZ
GDSP9z1pz/A/Ow88rSP3Yj3HjCRsP2OGBG6DBhvfOx2veRqmMvF97jgNyVoxbTlY
zkrjl9/kGr3YWkdyPouMQsvUnK2Gru1/DtF5mAovZkAhvoTdQ5OM9HbwOYe5M39E
6iyUpSvcal9HB/pfShc+VtO1qz4DkD92LSIQL4SHka4YRDYkEN4TzQ+UyCpT//rM
yco94FfaDn8I9UUmpW4hE/zv0xQjfUe+FNhuo56OKOVomfWtSAJZ/9E/wAaTZIuf
Q67lEXR/ggRITyksGvxiF23uGiOjkyMXH0CZXxF8AZuk9v19yraAA4FDXSTbVCAr
ZHglnXHJFObtekdez1yfs57PO7Jyd4ywfVg5WI/oNYmV1IXsF2NbeATIB+2KGKme
eWX7u5UyNKB3Nqx+LFoY7Z1vKxewgNgFSzLUO5cZ/vqBSOFUUUjujoKrYHx3akZJ
M7k6vR732dFE+7WqnfQHwlIroLY4GVqy3iHQ7SDjAiTR+tqfUFAJTF2iTVbupwnI
6huIeRVTQ5ThQXZpqfTK0tjJhESvMLJeoPp1NkzMGpwUIMjiUU4H88XcpLNleiH7
e9lf/Xg8NDrH1N+ZXWqfJfp9nGQMb11O8X1/ae/hBxrmLisWNhXCArYqTUJvbMta
7DmH/6Jq+Lr2H/TzOX+X1XXwmmtWuarZHw7X9iENGbGin0trT3quzpT5vR6PDO7+
O5K4H6wy867DH9opELCWnBcG/tzmfB15GVAuQL0nsUhVrDPwSK1gxzvE1ylHGkZ+
oYox/trtGS+tl4pRDMTEv52ggLssdCbSMcE85f6HkyF999RmJ2FjbGO6om280inT
ZrVdtXc9zN4R0rKKpAEcwp0hgVj6p52eNvdFCCh/OQMHHLKxcVsIAti730x6ELkN
pYPS+mFGEj6U9qtSE5c9mXkriBcmFjpcHBANzFbNvFXYywrgWCikjxwWLV4inRdo
oVvhhGGcIbf1ju6GqZGy9WegPsGVys618OYN7G4uNwDvDTcsWxXVTicTnyU0PzZ6
I1Sh0YuNIx9nu4ibggFC9bPWd1XFcKnv8wBgx/SET3gdsMMhwcsMaaKl7ej5dPLw
YcWIWhXfynzKX6MnZKHDcb6CEhWLJBJrTom/12HZtISBQ5EdGYj6YfCHtjtlsbRl
VZaM1LCUn60hBFBL8fZ1p5QPUcahtAekdeblj6I/s/vGLwX10QSeAuBk7K1uerxJ
55OwBc1WYAxyLChPH1hIT0DOrnnZzkRpJed/CFp+iqOWtUqYtk91X+4ufwfyOs54
mxj/gJAGL8GDThesz/7/LlMBH6+FtCvqZM4WkSARGrw61ziIxOTK9AfjaKXGVjR1
D9fVvSeQo9uOOWOmWVTic2KKEQsTn8sN8RLTxc3tSDxLMoxqst8gkja02zth+iDg
1JZJAoHylWj7AvvWhie/ERUGisNTHf/WeNk2NUjHo76biovljQWW0wQvQz4NIJiX
fyIdGfTD6tSczjQUW7TOuiF8NsaXKnqk/BK1Mq6UUfsg6399V0ieCDnHr+ELrjA8
umvbJ4wawRorIG87U4mfQrTN05x5o8vd2LGoC29Ru0eFKQDKDUDHCl3rsLbPeBW0
XLL5t5s2ZsiKFZWEQeJUQivSrMkevbcgl59a8CFjJ8tymEzr5TPN569VHAhiIfhy
6tgmvbgKWY7b5LC6vKz+DkQTpKdPx2IlJtKyC+F1/jlbZP/dZxphDc6K4+n8OmKt
AShJfrBrAWDY38TtDtPos37D1LtIjImjJUQ6xPVunuDCFObb6Oa5y85MIK3pWDkB
KjvlSs0wNaySQasdf70RIewVNnQ/y+B5LlV3g+17h6muF8kvwlN8aPRq5FLYuKMM
g18W8/0AJnctCdOXVGKHUhD9WZsSoNwI6U/sN27KPVv7tUln2gduuPHFOsHMCPde
+cUXNG6PuLhS919HJQlaKIMPKW5kCjlal0eK/csBwUEeIXAJWDNHf7fgRj4zLW29
Je6SD7mNgXFogOd2ag1BgEf9LJqYnYFNPOzWHahqtPQl+x1uP+dAC3tP2GEC2oIa
KCgCGjpoGeGk+yquXAM8BGkzRFywSNDsQttTeHVeSChfyahZwMl6EBNBcPcemCtM
Mt8bSRrTRzRMKweafJOsB7bdRIFdi3j1v50ogQdlwHhdVDUnSOyR3BtAi3PSxaBK
nfWMtKVzLJ//8UOiL2Bd554wZbndgRw5wvgNKlXRnewOCl1YbVATInVfu88yyax7
PtIeXpBYTgholWq3dnrVruJSgCbgYZajN2SKTfr2BZArc1noJNNF6R/sPp8A5Wkr
Qj7b8hHzafK+MkXkNzjRZ4151yjQ2VjLw2bTKmJToHjGdMVFpDGkv5XEA1h6pclQ
pwx1zSkAptA/iiJs2kpQKyWvn95GBvS2M1OppnDlKCOhRKDe2jMQ7pEVoxQnMq0t
mu+w9tbr0kvb/ife0f7zDrDPYwah0QKP/lszPpQ39iBPM/tDNZ393jJo6eZanBoi
uCUz0JW6eZtCF4gNaJN1UiHUQiPpnJUxBS4p0Cudzuzr6uFYY6jT8lE0EZrxwHMn
wIcDnhmhwKVVlgHfSmkC7iYMIqrbS2aKkRGSYjID8CSMaoJZGK/K6EedZ/GRDAwM
FbbH8bKZA9Wt0xFFcd0Pg2KCdNktFOYWo7pcMVYyWQ9ScvYEOBIQorSTm3TMXalf
2ZZl0FyXY4ljJEAEx7OnMTzRn4ueeWjXUc2iXDLGi0skuBoc95q6KW2iJxphFj59
OBsA2oJzG+W7TiUyTp8dio9rXnv6ktJTZSfxjI+L/eocjSB7AE/c/dyyKAplrzpt
oovpcoZ6JGHjHZ7RRHeK3OPV6P6M8f8BfhZ6i28HJ/5JNjsaKixo6Z08ucle9RZ2
rpAPb1UuEnEUPJrrm68UPdWjlVnFTveOx1yrhh51eY+2DvmhfsMFWFVod4WOwi8m
dq6kPLmqirrz755sYIB3yD69xG/OM01JAy1jsMueu4vvsKuyKXYKPq4QxjRo/fT+
JHyZq9gkmhUJvgwvlFYMQitDcrgYfZCyNLFjf6uYECux/mZkZQ2DUUaona/4+KHn
3e4EFcw5KtjChVl/O6RGNixjYwHyhY/vwlpGR4BIVMtI6d+DbBDttrUZoJJxAWoz
XCeNr8QKs6R0d60Z/ZnkvQ5IYx22VP/iLoovpGWbHEW1ISg6YUzm/VSLMtxEdsM+
ALZ63UhQp4fZQrSwg3AarlVjVuYCZiwOh6laHussmAXgcnynZ4BHoJhidPC24W9E
m8HRJ7pNDplwdmM3RsHdeKANxM0YZ7E8W9Zp0E9QnHf3voyYGGKG/ZbgNdBH5mzF
0i0AwcuQQ5ee6hUd5+/1pZqjjUj/qZqp6dHr8vHsAm1FiKvkob7sOehJTRSXDAkR
toxuHeiEY8e333EZnpDNYxrYaSboOcDwDhiHf1NcYDGzjqQSLXpDLGNQJh07yzNC
Py/G6qg75XzJicpVNLBngEPFmo9+W7GAI85tIBgKTmvpc+uN27GXcMXkeCyiPLdh
gOZr1bANtaSf3l3gru+uQtIoGuUriXgo+338ExvSfu3br8za6GEX7vnFfpWz6qQ2
75YopFjsvsji7x47ilv+ITQP8B6JrZpFuA0brnrU7kGbOwORpLwz+r7W07PvjL6I
PsYyxZfeQlH8iADeih0oX/1BxJ0yRA//anqG3mRpHM3j2n4ypSAgnh0jtXemuP7D
Pnchk0dMDlImZHk0JDtgid14TwUdAkQ1PnPlAnhFvpsiS4Kpib7hLsSXkH8N98L6
SglJLsSweIRCae4tAdOVekqpIMFF7cxstVfqv97UpnK6ky/geHMmY4FeyKHe9iJ8
Warz/UlHrIh0nBy8Got5WSMKdUGf6r7gNcX4FSDid5KkmiHRRB9KYCAKujRipTiE
qqD3a/BHOmGASH2DI/PHvFi0D08GCdUMjAntTrnzPP6JX4Tk1DoKSX5e4XL8MT9l
2N99wEFZ+zJeZXa44sG7k94/N6SezD/i7pOdVP/h3F7YlO6c/Ov6C37eQIaubnD0
8tIfSm8IGa+jTMW6t9Pr/P8iZAAtY0OEXMle5bBTkd6TaFpu/zceTfqriHtTQF5c
0J5y+KV+jgk0WixKtTmE8NcjpFXu6T2D/zhOcFEYKjqXQEX7uoPSdjjzpkszo8TP
jK23PiEGMyqxUBtTxr1P5dZsU8tzJZw3mSpyju7DJnh2AwljegGx3T+KMSWeLTsR
MJQct8eDdCo4uhoCJvKkz8Aq0NQFc5jKcMuVjx+gY6YxJncoz1WH/3rjPTpQuxfp
vvwrMe/vC3JrE1HEVU2BQINo4+XHYl+MZ/mY5XxOKKeni4pGAsxt04/I5nwneVfT
eJdIlSUGN3JM55AO5IhsJ8f3UJURHuXfCWtF+xS2jspWTP6/S39AoW8p3O6k0OlI
+jfkPlWgwTYgbLgSbFRNGVsuRErFvL0EvOxjc9FE2wYMurJbR2RbWnMnkSPrxtcg
QbZbz6X5f5+fThclNkBQZbU/Tq43u/anK8II5SqEtI+YqcgbVFSJnr2Pd2fpECHm
fqcDEqb0nlV+Ep9Bi7jQRVggqfztpAC5TPHNILiW5dnRZs+BIXwmMWcpDhgXHUvp
tyUaNuYlG7kOLbXa3PyfN42woxE0eHvDl8Ca9I6wo2XDZl68H2jHOEnV1Ov5zw8G
sW9mBq8Vho7iIcCUicneozW4uvd/RJYlPKuzELvrCBE9vfR9x07tQy8mLR7QdRNM
BvuGAE/6ZF0oWDiK+xKUL2PNm+F6hGBXUa0cl2/MlWyK0C5OYZlElELH69+v7/O1
WgvP4C3jjGn/m+F7vhDoA4JEWG8d7cwkq+d3u6JFU67L65MGC25O6ZXYC9nYt0H4
luiOKVNPrGqdsQDxxxh4F8akTA9k2f/E3yeqinPYyGQT68xIYb39qmV6F10J6cM3
BEnefopMhugq7DxmhAqPeNjwdiy9+hHyjRcaj+WittiJKYt/LTI9d72zH7V8EnU4
WL5WdxFlzgw/CXMD6G4sBVgKwb8uRhUDr7RhWP/vSagwxa+5sW4+xycHa2DWUuMS
BfcVXc12n2UlxjJylGQt6G2uc3ZX0ZAr6PN4MQYlcKgj5uMBhVMUOSGg+dy/BIX1
Bwa2sPO1c4UDwLA423Zi6AUa9D/zKE79u8wolFVCmbP8qywkTDd6V4+sj5nN+OJa
p+txNHRNJ/IFQj6NWpcVux2EE8vloAumr+uZuy9PSY82rodwys7mZHwH4kUqwOgt
zXQ5jqpuB+AvgV0r2FxOZXF6P7cuPnesCdJGkuCwXmg76z8oc6aEEbN6y3zYlWTF
UO8hEpMS5pdTh7GJeBviqhUtjOaNq5yeewAp/QCIAOePzt87fX+0NgSXcmzvMEki
RZv2a5yVtFHeKxklZMESHtkfM8ZJS3gorTwYnfdhHDmwxSa1TDN6I8KVwy2Wrolw
NwIld7Ga2/oiPGq7t+/sN6Z59mFMbSybUtrkUCmMIQxa+jFqYwC4O/svj1zlys4e
xv26RL3YXUGUxWY8kAzo0u3emAvM9Q17ThIKNb9HM+QJqSasPg8p1/6d30EQemy8
4Vhv1PYSSB8vuHohLXSR1piu5pvF2BS5lGvUcs6h+8VH8uVgntJdXfCCFMvDe2PF
CoER+ORfNE8384uCYWuWdI4toftHaqNfYbr1doggGyGepGCp3ALSY/Uuf9OZecIS
KHFnhlFdz1/Q+OAh6oudifUOJ5ntDHULrWts1xiviwi0ktO19exh3k6ijkAkBkga
Bm0QpE71Dff+68wCo9y5u/TqXOgoamXRxEhzeueBcSnUpoTf8A9jnq9sr2ueeQ3e
dsJml35dhTxitMirKBTijLG7b9QtBxlqNgn2kD395aGlwJqG9RMcnVpXzSWWj0vc
A+/2DFZ9mEcsiBFCA7Cggb1u04pTwB9TJzKrvZ1/OHmsXsOWZtzrljyc/WFNLrhN
LVVCgpKFFsqc6I5Cvv6V4jX8IzEdXEx3Wek8hH3jzCkR+TeR3YIxryJ9otQwypJu
7+IgLJrVPr/euF1jzltlfJVsxe/m9krwy5WT9yOTbKhMSpf29FEUTnaEQmP+A1ws
VpFguee7RC6ic1nYuGUwSzoxteStJhDkVpTDO65o8eMLIgGje6ciWA9fqifYOQP0
G3IbFyjjGqaP5Ukb3G7khYnmVMzrXvnkvZfcKsB+18XCGcQvubTuALFZzQbiNN9X
zXTGzDYhbOa2C06hPmhP+jhHY6nZ69DUA8hWG05xtusVn0kg+Kn0+EmiWXrCNjP2
XT6hMRPM/fjPuuXerapqwRDZudDL8NQ5PqbNiNzUjiWDjNO9gmpyiX00k5ZfbnIW
UpSlAgwy6hfU5nn7yTuLTU8t+tgjYEA3npC5SwYgIobjp2NnSft6usM1TJfVvYnf
Fu1ugnAt2ChF4kYffGSje/ADMN4LuO7gYntX3LBavq1lnjf4aPIW48s3P7UuBw/d
8qDDkCBOMX867k0t4M0RAAZ10oHsCfnIrCuFPXC2o0Nf1jUQIC07jv02q8EewAPZ
vra3R/q49lObZLnJ4aJ8gQboBV+hLkq9GWdiG0J9b13YEwcDWNH0bg3X+MaisIP0
KgZTnCDKLGovVqE5JQlvEFM04oEQt3SDyMajh0kBT1TaTqfyHXFb09SjH1vhISWF
GOFVknqD/Yh6g6lLAssy9yTsOVjHOXpnQQTPAdwWLWRa/2N2LDlcLd7OVVlXuTRF
5B7b3AqOMypi8BEVs1PIJrxfqkXUp2mDo12Qr0fvIntk8N0N8vFJeinsL/lnQ8MW
HHSAH+VF4YPJHBsXToSHo2z9hnY5z75VlGaTCriGQBrxDrVxN3mVjLDdyng41rVJ
3O0wwWl7v/PmE6celQ2mW8uNNrkKM/2GQEYT1bknMSdSLN9Z0CeaPRKPVjCu4gaU
Ky0h3woZxA17U+MdCtXoPKpx+3KyO8VnxpOJSQVjujyb3Ff3d5wpYOBkki5b1pm9
fp4h2gQ3wLfWrYJCAez1yoxMc3AmbuHY57eRmm+rx50QAa+49fciLx3W4PSXGxhw
9aG01CIeVtb4B3gsXycV4oP9TFzW9WfTCB1zWXJUklYvVfi+MLZDAkFzSKykvZxF
Dj94tMWIjqIeJmznL0KILE0xqSS4LCbCEVUErQthKTO0FkeoNC6JkYlul49f4S4z
KdkBDQB7a1kn5HUEN6wdPpbmhOKGBgF1YCl/26weJoij8+5uzzFMt7NmPtJPJqHY
FVaCA1NJq26DG4xBvYKgssfA4lbXBTdkr2wQ8Pke7D6Rcw7XdQCi5DYMjIcdbFNE
65pju2HVwLaOjY72W6KVSVvNiZkYAe7TVQhun0qMjXN3Yu6imra9COTXAjw/okv3
00rZNWyppAZ197s9FcqNyex3pD90zUjJKnKXzbs+jjufKXlf/Hz4NKKgQyxXe+Qy
irA6lJL0JSPQQ2C5DaVk81FHK5gyTJJuhih3b227bIRTCSTLZGNu4fjECMolQ2f8
4iwocs5A2/JN49aCgcuHZdCCj1wrYrxBnWCFGQ0HiYd/Q7h2VX6q1JQK5MQeqCMm
vSjtiyWD73mXDgX3rDQAYvYtfk96lDSRKnHq17F6ZIUYiUR1iQcIdVGrogW1sMgO
MZQCEE+T+US0GjQplXvz3u8YkUEsNN3oj36YmwilAqgyVuxZ/2kc4/w4XaHN/Ajd
5amZ7yvh+d4RLGZx8gd8qMYGiUKKyBDQB5j3mN9kI6vYQ+pUQxKTQBJ+HnbM1ynJ
N6ko/tKxjSWWaH0JePpSEhD3S81C+EUeWawDJ+inirMifRXerQtuoKR93MXtMPZ6
ND5Z0fntl5/nfOJzxZ29vFt8WgH12lXR9GhJi3pcvpE+Anc0VrRhP9SarrHBbQqp
4coDWV4MGXNvuCj4F++optGT0qtYxceBmxmyvQ9KgZgXZegt5Kl9HxqqBy6NTeFs
C6Ctv9D4vXxpcIWxmEOsJT/N9Mey+tc8QqgWjH021ty/mrqYtjeoNsMQzqkeHrTG
FSDOeODd3VVyHSBxLJWQOc4/er7lJ68UnVv+wMQXtX3U5LPv6XQwPuiz6hwtbZzq
XCL1W10f6iyleTLTDmhVUudBh6SYw6jWRFpAGtS5PMN7a6sn6yfScDQiZ8hcUhqs
1TObc+keu0774M1dqqfW2kwpgY2AdM1LB3bh7MswxP3bDjtb+kwGYVLoU5YBZ7co
4rSHiZ+24IXe+JBY4HovSDOXTo1+7PALTwylST/lDGvGUgUNiWUAEge8W8pmxr+o
m0spcYubi3QMa0IVECEJFIMMyVn+hl4hYBJQvtNbyr4+OGZs2J/oGrYxPLLtV3IZ
jNCiFBSxGCEo4ysRVOGBhCnUv0xirqyCq6msvbPjinoZPQLyafM4Vw7G/oDIyc8G
iGlZIRWlHvyL5/UqXgBUolxZXLK+GpT4pvIKb5FTRONek55hixhAlTAxYKCyIT4l
riQilicvdMnFMBpTncxdvntNlLDd8iMfLSd2F27fIp2oXvuEtdBU9jtsndiwxZKv
XAgBasVm/S6FGv0x+YO2a/OuxUwDzgvUpC2fSWAd8CEG1rmcJPwhsfnrQj2Iumec
d7/cPzJwNkgL/UYeyMj5kYkSnOtZfcvKnFmBiAUSi99nWUtHVllzSv6fLvtPvSAq
vdjS6XtF9bNKMWS0GEE2Oslbbg4Cd4Pu8giIO/LPeGTLmr9aVDWhpoZ3cy7Kjd2M
yCWAsJpAGMrJjX6THrLtNca3p/8UEMlp1zcl3qLEsBxFqOYtVkt2Fv6e6oNxShvd
bfX7yJcs2VE2H5TXDYE+eyxuBZgHeSZOjtPWOpbNp5TqJ5T9NWrCSUbZu4uSEpdx
BEkhIWmCDb1yL/dA+Pi/pQ5rp+4PpFk6mrXKzCHKe4MuNv+79iwT0xrxpbuVKTwD
NiJI/yzicFyzN94vGZy8+PtPOaYJ0msnBfwLeyMVJJCHvPAIWmiyndL8yrXUXvtZ
1pW0N574xdQdxTJOkz+bM6QpG1T7x1SxFmXkXrb/sR1GVm9eyeVPNMQ2bbC8IR4P
YUXXo6BH8Sqc0Jgr9aFdF9+7thJMoX8C3UujyJql1kIfQ+aDluBRwclXzTpydQHh
TOqlR07w++KOiF73s3aeh/qoJPRy/vz1O5oFn9MA/S0pltEWtYEUpDbjgYvN5DNC
jg4aYC0k6yIyG9VA7Mzoo0MYC2NZjq8rXu3cVs555VQEOG4czzAe+lp2aYTulSM2
VyRCDvALtcfT3BJx0YW3RuUa1a9zTOQQJVr96qNnguCFjjSvvYNp+TxBnMYzdsle
i6mpvtMpP+G2ZOCqrZoYWohRfM5/NGirVTyUypHwR/deEk6PB/SOHd5TYG8+lS8F
a4uQ1TT5TRhtmBqAkaUNewnlC2Z0pIhnKkPq7khMC3c9sQGPE/UMhdNYqJi06COr
vh7edpMdlh4BX7XATXmo7zQpvRObMs2EHkTnyZt9G7i/0313iZqcSTaD+9xsmj/i
nFC9CRRNW5I1pc3Rl69Vc8k2hX8JGfwh7P2D1bqvwBDxsyF7lWoU89CByCYiaukW
fLL7B4t0n01AB3tb4X5+d/dow4SFkcOcWq0tslYJE46LoP7KDosq84hdU4cWg/A6
vt7vOJnS0TZ0oLY2sdUPDXQogxVvdcGRvIGejjHQW91/KxyWbDBg5kQd1IqjjlzK
fRS1+AbU7bGT9t5xDuiFD6RFWBx5q1MVCSgQCPZiTlnrQAIrokEuHHOHyswy1Ehe
saxx45Aw3207YMZKmgbIfM2SIxO0dZ11238jYlVqChf5dLoUKOtPrijEvD3VllAF
ACeWcAc0h9dZ1gBGdM9bqBKIfkPFJJzTlDjO0a83e+TRVjAuY4npagPPOhyVSGPF
ajbEgttfLf1zku6/5RLT5dEdnQ4ioa8t/JFnK5uCTVDkbrqCXyiGK4DgkNmyBSyd
VxgeO0g9DA2HKzedpCNhLRzplNgIJ5YZXrJ0t5YMgdzrDEWJx2PpCGbq5Db23L3v
ce68ZDyVGjF6UoJrThODybxvc81kpCxzYe8oarKVpCVId7ph/KiJNL4O7Fo4e0Yg
UBgkUb0aD5ZRvVYavzE+iFL4yUrsboPo47nvrmhpJj2fC7nj1kHEWHSAM2IAjwfR
31EztdVIzMWEhzia9mAeYhH8I3b5SSa7ElTqDSNHUgbYg3ZpYYzuq699VAIJnKZQ
PfK7F6jzEsgJYRTMzu/rp7Wso+X66A5EV47kCQlv/e307BCokmizedVCcWhvhIQr
L7/n7HPLy0QT1MdJXceojKCUjPnEWdStvg1f9eGyvinpK5NnQwcbMNeDNQ68iYu+
vHyG69dxBpqxNnk0auVfYK2qtdV1l6q/CGoMpy5hePaJx8FqXPotR5fIo3nLxQWU
cPcReKefKTZRRQZBX2vNtTOCVPCFMpgXEgiNkiAupiY7t1yWqKueHAs5hD6X3N/w
LShk0aK5gCRao2gy8wgpFK5we3M7OZUN2AcYhHBoButoO5rWxhe0JqFXBei1QTDf
IJP6qFhrj+6AThpdup7TWS+oLWdIA1YGiS85UJ59rl2u5NdSjodBKtCUl39QypVW
wpmw1LmssDZOkkSHYbH+eChuVwtJA2WRmMC+K2E6GKC6V0vn/3GuH98x7Uvd6f0p
New1DEbo4ouaMk8k5GQUH+KVH05RDE9Ay6U/L920/fQuVF4/STpQmghQKl2RkSFX
UGr993QdJrGPnnfr5rVsSRRAu3VFypZtKeZhn/4s0e0XwMKQJbvOETcYWBuwx2q/
POM4Cy/Ha4stWOjrar9JvktyZbwiswM0L+I9LcQeqhmUvKyxDhgJjdboPOOS3oV9
Ed5b+ML/Z6H2t6Vxv3EJWimTcRvJkjdR2iesV2J9sVSeQbvH2Ka/mmlYTuVTXKfI
cGRozqF+4t0cZQPqPzpEgBWpqjJimflDC757cXG+TBo9fhUKx+gGDLzffC+PxtkP
8gRhyf8JIeZVcHfOWrQP/Tasa3n6ltZggqwFGFA2X6G3bU8aET3Wfjv6OTbojie/
sKnoaHvoRHVXKO9/Ub6BccgFXGLDx3Dyk3SJdvwP1yfO6RT/fj4P+FxudQZGg2VN
ZXuA1reXAGviXq+8mYNUfwQDwJXwa7Liw24+4ve5Gfm+lbWC+syp/CCkb38wlqGT
CAEiWsprQqgIeazygGoZ1HA0KKqvRV1UBQk5QpbswZv9L7j9RQWe/YOq3Xj2mmS7
srgc5yfbamuYPWiXnW3wHcLsXmUg7qL/NrRRp6OfFK/RG8MqVJMkdfx/T/ibf7zA
m8ywk2jDjzP+RPcck/+roULwRmxdyb2We+t5nQawUtvQ8TNUfD1XwZn1+Lpmd6Ip
VHRyPcnud5ZnE2fZfv3+/hDUDR/QquyVa3Nix5t7w/+K6mtBsuyTx9kaSKupK5na
I4GOJawY2nZ/hc+3GQztIsWyxpGQ5Qu8yvm8JVLHxDz/lvt4MXeoUzSu+HQJZkli
o5xXc8cb9y3pFnaPJQ++E/lF31A370tHD8uk2re2ToTSYxsQZkwkHgh/TQb0ur1D
ElVYeTjRT5ALTNuK7Yef0bVuWKFZLz9NP05+qI5M5pNJJuQwIEft5JkuhO/OKgfR
afi19Eacr0ojmthfAX+w+oQqqCYsqhAR70jB3DVLhoK4dDOy8BYbwCIX9nS3Bvj6
EjmnPRz09wqePdpIWB2/wDTIxHHYtyc64YjF0d3jlhux7jVHEza98TDSrOoVoveY
A8GjOSPCVm/WsXHXG++iEYLpNz/1IBOwHb1L8xlw6e5Qi1wCp8htYUY9V3HEGzKx
9VOJ4KukfPWyL2WqhgOoj1bv8xNv5ouWXumGCjw7Vuouo0tPmpZDdsroMoeYVyRS
2YM/UBG4K6TMZlvxbfwFPVAHEcjkTINco2r7+rUHLCHAS0w3XD0H1ZclYqS0k3jR
1uBvDVfLWeOs8aydTHSF/hAULUA/W7T0aZE2jTiLc9+Jp8N8sIGlDYPfr1TYjgYT
IZHXnNn1ViHNaDOpwBReBgHT8HweOO12iRv2yjk7SIVPWYzdl+7uP0JfUurCK8vf
x9VR4gFKmzY3acBZQw4Xov/Ne8cZ2Pu4sXAfPYDHoSBGn4CbmiSF6Vk37YAF2nY6
t/Y9x19P5P/J56mSeDHbbfteqe2x6tGgGET45Ltdl2Gr/qVN3Fw75bu8JUvgCO/d
QR3L+Fb69jYAbsNkMxNxGY0lJ3SfHMfOG+QS9SSEw/GRouKVHb3Smt0qh1zfRDqT
AvgozQegdD9iZCruyWioHiiYFBdrUSLhCkNmsIWJcpQ/Ympp574IKzIqHgUCxye4
j04h1UDFBkTgth6T2joOFv4pE86/tvDCXZ8W5CP0dZlJqYywXGcCgdVjUsm86J/b
rhYYOnDAkUORksB084I0H6nB1H2lKcuDomPGAkiRIwMHtkIAMgAR2LOD+LNFyiI8
fcwRKD969XIw6cFGLfKJnQDIm8uuwgjjVpKmvI3wT5lHPymUj/9dOHr4fT4hOAAi
chKpz6gUWa/w2WSuO/nEdBwSYierJjkgetZS2H65PDABCGXv6K+CbP/6CmFL6PPn
Yx7NGfblyDUQh1MQUFUjR7LZCLDapZ55rSBhMQk8fkxK74Q0bc40sH32OdjRw14r
TqC70+vqV3xpzfVo8WzE+S9qntWp49JcXvOcBdMCRFIU5+Q66aYcYY3ftUns6s3T
cuWOFqjnlWhY68M67cNKM7zhWJipPsto1eLtBKvVtiMDkIpTiAVDMuMv7wv4pFB1
Bw9xTd29L2f4tuJ+yp9+cVpRTrNxyD3BM93kH4uK4ZgAS5f425JAWJ3itzkMwy/u
qQ3hjSPHffc4KKT/qMTAyjz6rfl0y6cJWqa7A6qduAlEH9o00IOduZS4eqwqC0U7
hGuIl1J18nIyxY+Tdtk/JmXJ/ZD8994O7pUHHGxbongY9IqhyyJuZdWcdTqfHJD5
1NqlHFJ0FrBEwY/fqrWaR9inNso+FyGFsp3LVAYUewVL9MmAN2gGB8YR7Rn2SC+J
Qfq7M9NfLj4AgqxrPt+ZKiDwUy618MFx6qnPBH6/jPBXrLzvZHPBVYc9vSyJagbU
6n/DRKGqa2ImTCx6UDDTqoZ3q1wUI1ML/LzuMs3Nbwujm8oCqHO2Ap+qU2E1Mq25
JFp60k9s9QAiVG5J4gjxKkg0gX8Zfe5rEVGEARTCbSfcT4rM0/XtOhpb8NFoP/tH
2mn9pylJmw+49Dqm2G/US9RlplryVh/O/b9h+zsVTOBPcGGTs8FB3lSr8PimVihY
/fDTKTrsdFvDpuJfgJqvKGyBu4WdyQ8hruXABhH4kZSxMCAilxoaMzwNf1d9SmgB
2duiF0Cb6KSxA1S7YiQilTIL2j0VxxatINGljxWS4aU+lQGU41BAPycNOocpGWvI
sL8nnizBE8M1LqXRf+41uB2x/QASVmsm8dGhZOaPyRahoRvsPz+iTvieraEy4nXI
cQZIG/5I4E/nYHL8riQRBzcQRic1DomGRt+qA/4SvlFQfCH9GehwAA+IJ9PsOP2r
P8OhkRORbA6kuZoL4lTyLeqQrKgVQG/vC5Mx9rzqnLH2UmKZZdC3hAdxo2BPPrUF
2EWtEPUssLqZb9IMfCo4LzTscVKSS3DxlumAA6781mcbr+8IrIhmQdYF0MdiiM3S
JnBgBqNyvBQfGGx/O291DxWUsOfA1dSZzvvLgCvZO/4m9QH/4KH2Qo6NGQyK5z2x
jfFfCVAopHwRUWAJtcmZAuthFcWq1IVI9Td4/Cu9SipmqqVj+ZVLfrAhDfBmEl97
fXUSkJPBJn3nPO3kWgMxcCf3wGdL3UKT4Y5Tn+dG4zMHrY4fWRlUc+XzcAf9m4qj
X1AEZ8tOIGEQY+30wQQ1LkvksSd31MNXURMMeDV0vm+CxuNw3awKW3V7AlHyXAR3
Xc6kDQlHYRnAhf7Nn8UiIHhpv3UAtbJ/6Om8u+KpWEnu3gc4F3JoO5BKWCUTA/Mw
0VXQYCFCipUA+pTu1di7kGzBl5kA30npC7uDGAqovZ8f7h87qVNt6Kk8zwDpqWf2
Wl3G97nSE+cCbyy8WhhxVGjl7JwRL8innkTLT57hd/gyZraCvBt13aBkGwRnhjpj
TEar/CfpKp47u5eKbp7xCxpbGODu53bxVy44DfzUz81a/grW6itpORB3cUCwjZoY
Tc2+JsF1VvKVzXOd2aLCb6n+I3DqctVsxH5Rg7vFLqGtqdkS7WSm+ZlOgt1dL5Qm
6lTA5yIrYs9AQSt4jCdyRCojuEFbd/LDYuXZ1G4iXcq6A033Kb7MH7uPfad3dvL7
sfa6ffhLN4LsXuteHP8SLbRDXztT1L+ckue23M6w0BBnK6EugPCG0HRAMNQp9AUR
xpRm55mhXmijPoHe8NqXyGWwZJ7h8Oqhtc00PLr+ayLSXWS3msk3NoxQncMojq6B
sGusfNeLjPUadxSa0IlFoJJ4mxn6f36F4gL1LrlSMKm/iXWMQxAY3kN+G2Vg8UEm
hCFNHYKYSXlSYc7/E/UkyEM0v0UzvBPXtw/QPTTvcYvbr5PREmsCC2UQFVQ7j7Ie
AWWCJtZzZfFXdKybqOwYkRj9eHXQCbrgS0I6eC2aBFrhnySJ1MUODsdzu0GnZznz
7yqGivshx3jfv7G9OO7L0fsvu/2y1tYWyZdaTiUEFQtvv+OKPrRX5a9FhO/URUpU
Hm9XcVRHD3A21UPj5CvlptQU5FPEEGpAscEj6ZlPolrfqplsp0geYlnYcrwDRXCj
co6i93T8syzdhEdJFHUvKtOWmYJ3/1/JxpDQkdv/WjXPKK/iCramTRVQtP9Ta4xI
zbwK+7L56qMO8AnyC2ORwONQzocChvVRuyG4o7jf5/rIAoUIwTHaCIOtGdkO7FIQ
TtyELKirtmi3ynp0tqOC88iJT2vNmDJsRyHDxJ3qgLZx3DTMHlkcV0cEEwLWANvs
Gu5cs5ZLQQ3RRjvIrwhmDwMgbbk+3K6cGMUXoUKYm4pgKa4yBMeB/QAqbjyLlk5m
5WQbuQrxrUUhrYcBBFzuqzpG1bqTSBMQ1jrnT+g9XvhXnUXx81GZT0mrYy/wIMos
yQAQTv16b/cAX3GwnDBb6FkncIykK4v0qxF6YA3+b4w1VU4fj2rFUCpz4BSKVV2X
UG6Xd/bopkr4U1L1IcBYfUqxCkNZFl77dvjHXN5Yb2JL7eeDLcy7xUWQVM4CMPbb
8awbc0gphK6dOzrsfm9nbSGRHTzjSkqJonqgJ3uynQzgI0vXxvJiUnQFCmcj+plG
xE+GNeVpjd2ePM0a+ZXRoCxgvrZcJAO8WWc9DwizIcnNB/KsfyLpsFo+S6P+mDgR
YpWCft1Xxjwyq/zNLX2Kn2cmbj3uYV/KDxOKIU+DLyWRGEE8SRm4u8iuglcUIK+d
O1rarlN4BIOPxop2cyxZ+2huwkHCKgGJdc3k/ArIXizq0a+LQV9Vku6HkF/JSnNh
BRFc60q2Q0vBZif97gH+pxSDtg1JsOVP7eXD/+EgUEMmIU4by5Ne+IeED0kRUq2L
BB3aSUht3U3dBAaBf/A9uFANpl/kiz89Rzk174fyAggYE91VrxsGkWCJDtfmfSHZ
46yarBbaUWHo9sqWQWJ/lfDrwUr71MFa0jixF097IgESX8TyN43pJQqCFBJb2hzO
FqH8/t41KvA2kCiJ1qfJV/CwDcvt2mHnzXSxMj5UeZ6U1Is2rpubeDHIC0VafnTa
nqRZ1fDfK0Ky1Vfr7aI9o2w/+vJZvYNaBq3evwv7BfJZERy2oTH/kQZLRrdlJolv
kdi7ueNkzDT4w8VJBy5H5KFo8rZ/wGrZcCif3XRHoIf+PYYENoNLSmVXPj35h+Uc
lCWu2jFS6ykw/83AaXOz7pXGMJEC5B3ooiBgF3oTVqayyrr/lU6FJC5/9QbW0H+4
Ver3N+AkQ7JuPoiNU71HIxfI3V6P0iIdUbnk+ArezrPt6zN4/HTCQUaXw5EVw35V
uKj2IfMD3MWz5CW39j0B7+jjrQLy2kqrr2/z9JxXxKGNxSwt/rBFufO3RGjK+WS8
hARfGPkTam1zbH0g+dbi1PQvyAdyErPkEXgPeIHn8oSOLIt74nRApBWRVOJq4hto
YT56IYRImm2gyfnHE1034VhkjlCv5xQBoO6GFnu01iKxXiSpBdDkP7bmpH9y/9Dm
qKALVWGyKUHkRQnmBC3vMo0W0MtY8TuTDfQLNswfAHS85qEE7z1nsLoasezbAvBZ
LTezPv5iV/Q/q+Ve15vLkxFN3x8uLARDq4Rv9nYLr2xRrnQo5vj9CJtAITJ+Kf29
15JWbApgWsG3KAy5FPvotW8NjlPuM7cTr6Z2nkGa7VdSjAvhTEzm+G2+lnC/oNRC
nfmN84IfG/5m0MQHNPu/i0PYg998AyZbJTBOSPfiY/SAtym22zn28NpclASiaa29
PY14xc6Oo1SAJAbJdOZ+MkK9WxPGsCGfbndqBue41CiF1cA0l8d6F78zdp1kCc5Q
KIQ/k6A71DV0tL3GfuTzUFTXQHuj98tHViK3AqkrUsPS7qi1gyPBZGTdaPKlg0mq
lVyw2vEWdTH3Cr5AWbXl5GMoybrextZyuJH4Du3K+cD/O/3sCqhqPl+vYc8YakGS
+h1zIyvPyB5S5iYTJTrUNm+hFGpHUZpJLqA9x6boBLuRLC4d3BHF+qU7HtjiaR3p
typMJI/5mk4OCDiGdTQg4k7+qLFl1jYZAtL8FPktYlZfRMK6L4zBrri5TlPkopFc
w7MmI6AqSC66qNLZqqurYtIo73DxFA6zbAQSGtvSK9P5TqjjIvvc5wiSgz8Ze0Hm
aTj95l4ElQ7wOTrHQmJHpsK9JkCMns9hCS6E45BomaqOYAcppzWTiINzpAC7MneE
2PSHIwnRzUKvpxBDTNPHLBEsXk3qoI0/cryQCA4yk4ohdqbEI/s7ZOnBIGvtULxV
SiZQDjASnpF7l2GsWN42nc4KAnilDU/mxZ0JWGf5d3q5GACeE4imlZG7yUxIa/2P
iUqA/OQvOte1NbIoi54PWrkfKQNcBFVSb9Cj5VDu1iybe+3SSmnobAZeRt75bI0Z
icbaZv+T1rSreVkMVD86nhvuzgfMmLnVREPDekkCyibZTOcO6Gu6nd/TaI++eLIQ
mmBvL8olH+BZMlkgiubn7o7Mw+Ab5FBiWcU1utGKW7WepFtU5IUK5KrPeARn6XWC
N/p8l10FqHqjA/7w/FGgNS2O9YJdPFctaym0ohXaNNGSxemJV1t6/Si/gCC/kWO9
FExKMeYG1KxFb02QldJrRdyO/mr/WgczmsfWlFmmZxmNutsmHfpto9lY5VoSJ/JJ
01yVDj/a05LLRWX3/V2liNJcqMZToAOVlVNZo+GLx2F1/FqERZijJI6gtnD7MPrf
vxknF+saOe2DFU3KQAALH2JG7ToaD0ZWSAc/TY5ltyI+lmgmaAQuDm/cx7HKdrSh
XeNtv6SbmoKO6c7uE1LsNhND/ZAdRCKMAJwxTD5RGjRGbvVPxu85fiz31o1I+4si
x/HNzhrXJbzJxxtQ0sD7F0gPgeRm4lUJ+VtlMErQ+e13Lyz6JoNCb38iDN6WiCP9
hEgMIipM4BBVHMb5OANVaxvx839sMdcUuEpq7HOadXNh7nZ3Ws5tSTBhwb8gXv0N
PSRQPygGpqjGVMl+tRJKOBkHFTWLvbo5Fi3xidfO/E23ELZ9SSeEAe6VhH6bvoH0
q59brupnjgFpraseWoO0RcOXfEOq6eizgAFJOE/7xvDJTHIJoUNuIHm5/HX5cO02
86A0v/lVzb0ob+riGhZtNOMJJ9V78lsG9xIv8MvVWu0QOT7WoScwxf/KjN55SMnC
yoJDyu6nu+wDeAbeo9zFCDZJKkWxS3GYgWds8Byu2Ha4PQm8DQYK+0sIa9x6MR3z
BNUHTcS+5NDGyMIS3JRzx5Et4K5DmA7L+OlhW0+gJSUR6CioRulIvVd+QFueiY7t
/BT9zKVg0RbpTSWY3cPHNg6Wm9KTIwrOgbrrPaHpG6e8vkigDRaT38UJIyVad0zy
7vY82K6idaWAgVEOv+9fUhBKFy6EKA/e5aS486llQzmvfBEdweUfmUsODatN+MAY
i9mG9zT5Qo1y3vz0mbSEnp2e/g2b1n+MAUdX+hmeqEeYO0+0yB+lq9UOaaYK52v/
8T0uzrRO2L5EBfzAt5osaGLN+fiO9eQWcFmCejxkx+MYebwq5sbQT9E5YmDe8l8M
3zeZWeERkQes6lC/hYMCPMvPBH6yW1cBxHSudgYPKaxqpJ2F9N3Er5BAbEOYXMAZ
HQAIYTjghviXQhiRPJXVHrKFQfNmP/C2WCRDGpMdx/9vTY8RD7/Fd/48T/93lZc1
1GEek/JDZDHmGiV0GRDpO62a6GQAy9Jn6MAzAiJcLwf/4YQsGla6AnpPdtc0gxL/
XPDu3hAaSMx31l7H1lmafB9/+Otff3VA+DcQBWH0h+2iHNBYUvk7H5tCENKTFPXq
UMDYAGx+BFbr/e5v3vicrAG5LS3pFgjt6s4mQU9PyOt5YkyEGnkaNbx9ABg8s8JA
DGtQ5VmSlH7dGGS7V6Dwj9zOyhOMrS5LnYAUc8Hg2j22pYjd3F8Qv5GNlgYgfEJp
EnTMaWw2r4JiCI8UFy9epapk16YP4gLWQgGLcFq4q8vGk0uZ+Mr+YTU5RDLwdRwE
SWUL2iWEjVtuNP0l9MAEIfLN/lDTqxHsPQzlb/GRYtrWaBuoyLlEYcOwA8HNTuIB
ROOVwTlhGi2SgkTFD8SxVecKN/A7IgHQKKk9h+zqRvyXFS8viEd9xDib3GFZD/Mo
boFa2jdykjLhNj/AW9EqQsv7z4PXU8CHJZ55OUbvnMq93kQoW6/TC+xG657JVONz
GnxkCTyUVP089oG4bQyQWa4AFxhrbXdv99VBFt1u8QadNKNO6CkoqNNUIyWulAH1
PS77bpomctYi43ZNffIsqgM4tzLTA20ZRiEJqp9W+bzKuBM1sYqWkOBCIW5Lyuw0
9MaAJJn2qt0i4qk/ZQSuRDerzmbmwhbUmUJd4QHDO9AmeiUVCwH3SHQuRC7NYnW1
OIMXGW4yE3sjr3TSccgRl+E7Wb6gD9SHR7pOsZc2y9rp6zDzqRioqiR2fcIZU8d6
4TlL4tGqETKRKNTLVcRHZPSa7Rx8uQgOexs0xMnCzteLG0dP5VBewXvmW6oAOl6i
o6/9E1etIBlPvDBhNrja5DbbI0H4utOqIdhdMF/7xO3LxJ1Y+NUepQes+DZvwgg1
q+WXdnDtbLtTLrUvZmUPeab99BNMJoihB6t+kbY5dBe/u5essL9WGQ7K58zKTSM6
GmuoMd5KnkObPgSTRAPWdIIQPxMAMiE+jX6alusnpa7c1eWwEEKVM6wLFm9SKwoG
iy4VwlFn0XUvDmlvnXQdTftpOoQSQbPsScB1DBO7guvth2tkyVjw7uRD7Sc+12ld
hNX0urION9MF3MawFQyb4pNRf68EjWupvRFtaJu4khrWGorNNCV41ck13Fflm0re
oHpW+Fy+xnuqGvmFdfKSCk2CTTIId59bLuBLAolWqVm21gXCf4UoEPtl5g1Z+HKx
+AKmTGv4Jeuktx1qPP180lB8/4Rw+yobUb3E6FKxd56wRl0bHVtIrzCS9dBkA+v6
jJZsHe9v2DWiFZd/fVQ0GciZSZeM/akf0O6UZABmmjlBHIDshXSu+NxMG3tg5IId
2wIGusec8SiHPPjGncRxKL1sHem1UDCpjuefFwaRDgDbh3fWjWFmBpry29zM3vsW
ZewJC5EAfvNTCqNhnA39g+2Ps18zfL4b1VR9HiLOAaz5PSzABmNfwF62wAMVOmXP
0MHWq+2JJcItn9hn7SN+STML9HZxQR2X5vv4xDXJWzJcy2X0hiMhsmt566ptMp4l
yjl0znyhHqAw4O1QBQMw1XpRGlH3uSrIXGqXOQKdUkZdBwgOFydnrlERue6AZfpy
OejiIg4kN1WKm1FQoYnLYfkaDmdf8wVYtSyDalOeZdo9Hzz4T8eCY0zaVaIvFiS6
uppefBO7dsx8eIkCjDtdJ8HjxmgPhRdpZDDSmUOJqmDvi5/Isezk9sQPOaxQW4DK
NgwdKRDly55UW8xyQp1OcmrlgcpqI2FwN4h/yHPS1t58oORi0rIMghS+OdWJCPYN
qIP0J409F7bo9wJshE/OHvr5Y359Y4OT7JJw3gGDZPxklXDY74xXxoJLjTs+oAMr
71lR5e2qoA1j1GLoIFusHERRTOqaxYcfJV2wUc4lmRnvgm4ZcjBsL9BgwRVk1Pm4
VIiOopa9oEQmWUqLRQF4xnqUTR5r+DOEq9elF8JIZRJhf9Wf4GO47J1a7xsHXdlJ
x2HDHQA6qzrne6h0XkvPLlYLdQ4y5gkeu74G72OZiY0hpEeuhk3lsL5MR0KSWEBQ
VRQiJt0RMKA8t2At6hjsLj37GbR7KvMwqwtZd6iTmAlAp4CDYLeoJKQcUhKTgQ8b
XNckBkBg9zyd1wd+/zpjJmViK5qlRYH5TObxIUuumQpIPcly4+DhFlzpHvCKIFPc
P5fhR0zM3rg5wjFNxMozT1psjSdiCNeoIVdp7bMuk6fSpF7448ng/YspW0o+dahl
5mnmFd/IFVu22pTxAXSFf/p7qLhIaO6XL/QGv2w8GMTAUIjL0pijTsnF5lmc7x8Q
3QMcBpH++x67gQy3KWNMhQXk7vH2ZVzHUWhYOmruzJoxpcKBe+XfoJXgyuWskjIJ
yGsz658Va8S+1hAf5h0GBkC+oUTD7FVSCUWZqvlYwpVqulCLYOYJTI0I2jLHoAzX
FIf436Pd5ZfYC3ytPVdjCHI0x9w8Tf25hc5Dg1pwb7srP+5kwChBvai/RmRVKpzn
uheSUWR6+OtqfV0BZWdcfWb6F1L1zieCKgar3h9//TH8NlfIz6+/W5QzAiUgcI6C
68RiPbx8T5Irj12DpmN82JEULIeKsiDMyaS6gZf470VxWWOwlMece4PTOmGhzVKO
uAy4i2rmcaonGcNtq7NVuwS3xj2ZMRhtbt6cKj41DWtGid16FoUw/QliNZCrL2mq
+tzv+jlgr9lcozVsrbdn9WEXan6bIK9RSS+DNDxVihqNRXnacWQ8OgcpO22MhvGu
g/eVJGnmO8ZVRLaQ++ZV1y2yVdzn4Biw6C1+yN51mGzBiQQak/64a4kAIIRtTXr8
Xw2TRZyY2YxUMAMu8nkX8Gyi4pLEf/xnxY/hdp/4j6MYQ7d8s1ktbhO9UJLJxAVy
Ngg11PPwMvNQokrzH+j6badZnlX//vN71Qgn+TJnymvsfbQMym/VtVPZc/Tz46Er
PBmyvy6lMP+0vubXOba8tsMBZ/K5dVD6XaMsruP98Belun5lZsrOVyLATamk9EoT
fWvN7WI7TP91P1cTw4+u8tNNLPqDYeatxpaW1ZkTK1oTgwnP+TN35H3VKG/QvKGh
cmjjP+K5OVDKupwX/b3MJ4aUa63DsXyphmw8kLWtsngOLgryoUuZMGj5vVTf/2Sf
zkCfnJcPGtyQSoIlwWa/Afa8+GdbI0sGIE/58OqL1dKFPYvmqKFbvq3TKPVZuP5a
G8HEryk5gj51vBTue3l8jgSR0sN3NLoe/BynZ6uTQx1vlgPWPZdH0qs/y5UDndm2
P0h7ZPfGHx9yOmuuRfWL/93DwYw+77hK3PIlmUkOayEGguf2yNc/bM221D+XbBag
z/afS/awpNtdiZUpuMPNEPdhs/o1TqDwyrn0vtWojoNFXW7FLkbDwzL6cF4jYS8B
ELCCha5XiJFUabki7a6w8HO2iu6TFYZFn2X/qTz94T1zHMxz36NSvQd1MOuAm49d
d3C7Fg5hWNF8y3MorOI9NrUsizxYvfxDd0psID+5CfC2rNEAJ0k4FYGQWUWpwD2S
9HzCXTDpuWHwpEa9Xl1QD/1Kqbfcqttln+ekTA7EEY8q7RKdrhAwGeSmjimISR13
wMyPtFRKjJAghCx204T9Xn1bt8yzDpcbEdlAkIXeSqiHsoHUJy4z/qajafT4/DP8
IQPQNJjUl/JyTIF6BwGjSuKykFFINrK4uqxLlGsu/1OOpIra/n5lyVNt3vzZFnyO
ukzYbJeO0QG7RafO/6fe7229knKKoS0O7suivykNkD86s8B8h1ka5L6JHCgKSCba
QiGaS0gSagKygZNHG+A314lVy68OucVYVh7iNSMLlZmeVg+yafAQ9vXB9L/zJBiP
2T5MjOJfTvMrIf7Ghqpj0hNoxzesYtfQwkowbXrfz1Z/keohyTScYyA5gnaBA+WC
z7qpa30TgP3fIT27VTsSVBkcd/zyBotB5YLYRoIIi/eb5P2e/TG9hd+XTDCh4Nc2
SvFTjZAuaWxtiCqcvGdkF4/BcgK7r36PP8hScT0iN5q5ZkI5KOy2OBgJPXskrY1k
ygc2wcj5fn1MIioO2O1Ha1QptE3bi5QjHJ0gj8JkFZBlnlO15GYvsxgxXrNHLVVf
2a0/lDuU0ZRyfpXH6+GCr9wzbmIEvXFazvytdiHf/Jye2r26FgJDYYQWVHoL12hB
1BXjtJbaNuuFN1tsyWqM8lFv4EnNclTJ8VZck814MII5QIjV8691rBTDqi0+L3Fm
vsiE57eYd9R8vCxHWHMV98oK9XhZp37yhBiQSJEmqTnW/Rkj3qmUqOgsyi2Wncwe
Rln43Tz/JXak88nac0R2ls349askOaM2s7Q6xgtdFG6H+jev9lEl8d22Ct/js7Q0
buyRR5A6DBbM5wFV0U6gHU1kiS5eIrQG9Uv8p4bwDL5ITigKynHyE1W4wvkd8GDV
4mm8yAI8HR+oieg2vfFK63PtCWwcvW14Q6alT182vGJD2qGlYcvQBK6fnwnyZEVz
OLdIhvUEjvM4bEa/sIXlKp5MlWr/rZjYwTQPOaE4EVEUeEuybQ6aW9J/CeVJsKD0
687WLXHiE911vrMR0pyDq1qhAJGF2v/wBaLou8osIb4CnDy+uN1z702eipU57PKA
pDGCbtFUAY1D0bCZu6VtA7e13m2CfFmyQO8/V75OyNySoTuC2SSBy9V48Jpen54l
GC1ybiwhtebIOCWqGD1SIlxJWVvuqbcvGvDoyGpRD4vgLk7EyDWTAmDm1ryLuvMj
ayVdXQuEuzEHwlTVrZN55/ULgQHnR223P/K/+xqY+578IsWjEgHi9wKcjP/7IYTo
20QiGy0wcdk9ekA9sKTKPKfo12x2HgI0tc/U4g2ZO20dX9IwCZpn0sQWdmfN1FGU
hMl4kR6GmAsHKMEzpIND5GJmMEH3dJRZaPo5+iCQ1PZ1lMTktGnobJz0mHIFXaii
+fW/G2FoqKsDiEBf+CEEjkMWuTiopdUlxa7Cusfd0V299yPzyFB59ifykWVmpCem
18KOswLFUhLe0kUlf3cuz/GV3hz8bLFI9wv+RHqhCeFbYJY0R2NXQL2WccDrE467
dqeg+0j25EYc/Stp+qeo9mTN/ay0EwGTU78Mb78cGdjbK/ZDnINAQkJ4njZHB5dd
O0vDx2IWzxREX8Y+m09URoq7dGQf4jmm/MqlZ+y2HBnkB0iTUJ+WUouUFFgt2fhn
FT7K8H/1rkgEyh8hhzjhDWztiWkFswZT6iIxCVOU0MoVOgnYlUGbXbYQ3nqFp+Fa
rBqBJhXlv3Inqz/SDdG8Fva6DPo65ix7mcf6U6DP1IN3vhQzQw71ijZOmcrrISCe
Lfxu2An9yST6tSQtMA/IMGRoaLbvfj6OziswAZ2ImPxCIPSByS/1/vdFsrpFFxe4
0PGEgwTm8BjW+QhCdj9nReTaZgW/8n5lQjedqbRaUm3oNCXRt1Yw37gNQh5WrMMF
F/cq/gelbs/6AK7pcPMOPlA40NBW5XQoIf9UgJeVHVPpfqAy24U8aNDWSHE1gNR6
+lY7ps5KAswLldArsC/AGUZMMYpnfFKBsD9raNTyfV1EUOKdQ6VYuh+Nzx/gdJws
n7K7m6j2WPfvtKHEvaw7HllPR3IvVCsQnRyHGVzUo91vGWYEcYAvVK5Z37BYtaIi
fCEu5xuinnwOvri4mAp+fUZm+7ecZ7NG2Gtsk9lHJZqqLZommhW7vpXgvmEdqFbH
7zLo85T5uFUgsegdLvIreoNBRl8bJiMZkqlEWHdKXAhQwhO7PZqW3a8UudDupbTK
ZmHhrX3uzRLnq/epQiBoqd41R9luiwQk7q2xFs3fUb2FpepXSJyZcWrotf13vOqt
9fmqE6YA0hQvXoeYFSUIwFR5OLsRsxB0j+DjkrDz0e5JTQ1G1XjhlIM9vx2wxs77
1Fa+8CAxj5Rn6a4hQ0dSnq3w7K0R6trNAqHqji/DEPf1m+AHZx9907KD2U6bITrx
D0RwdQrRYwk1Z2EFFrPVubfy+9oNV/+3e4w/vtadZXtjjThsu0G9cteIuAmobKhR
dhSvn3QEdMPyXiY70SbfO1TX5mGq1tLV0SEaLVlVIRD1wKYbM4JLSl5GoKQdI9E1
jyBkPFUMC9MXDYbvF6AOXbEPRWOd8PjpGcmfLbWA+08JvhlASsHWGxUpONyCReiS
gavlV7FOgYhaT+Ii94r+9sYzVXB12Fm0S1hMF6HyC8OQTp3dEekH//YgeCLYdq6F
44MWxro3dCQovXxpqqUmv530SEd60C9Nt3e83/iAF8O/yfuHzUUZKXTli9+/4u2L
ySyh/p/Plsmfwd3RrzEN7SSGRpouYDwnaRbh1x/04Ia+dNyaxMtnqQmQEgNTRakH
DI9HMcDI67ZQgQjE6r9nfbo6j5z9MoYBnm0skCD57BhiB/C9VYcd0JV3YjgCvh3x
5PvChVJHBP/Fkic6TTckiW2v6IQBFYPZoZ+isB/NMXJC4+Q1n7DX25rN5ROeFNn3
CBpBm2AuWWpmx7aPj90/uHw6Nbmi/Wp7dzq06I+TyDcNWLKc2CcishYOf2Vq9Aim
qcdpi7/XvWEw1TOvX25yVsW60sePvCbl2/TLPvNlSIfyN+iZbQunmAoHptstXift
+E4RwAJVnVojiNw3TWmbfNdkn9jClshIKkUc/kWPARBcByeHUp0xV163FZJXFjrl
469umhI3GGwx4XEFFakrrKmvtTQ+HbuFfhcDpXIFZquWpz+5euXM4BOhfoQeBo0q
KTGlVPp9DQ0t1vgDSKdXrivD6nZmfpVHSXBvYJwHX/y0BiLdiauZQpeJkFetZIi5
9kaFcQ9tU+OI3B6Z3i+DteY/9pP5eh4di3vQiCkQ1miCG36PotyTqM4T79OgeT5D
aWxw4rG4llBdrbwa9D7gZpgSlB+4ywSvWefmiFPz73ts+PN7nfVFQ4tdRjOBV6ME
slpaiaW4a+U4X6T9+wkuqMwTFc+LaJMxDEpZ3qyP2jBd05OQC6ZBd79+OYycHSoi
MbVLI9WezlQ7I9nnT53CS6wgA6AhJtGz52mYX8XO1UI8c9IAkcvsg7YuM3tynT00
do1vfc0YPx1ft9gA1NZqnpVLm10wAm0rq1TCMhZIlB70pSlheCQE9N159K+s3YXK
wl4HHohkvD/btXgNvhb7QCkjXWXEnEWPIOxa0DH/TSjqGt4DNh+0lUWqpFNnO3yc
27iboSLySMEMT9Lv5IIVzfReOk91Uu7gfzcFNc/8MsIZX6xo5g1sS4N/msgS9m3C
LaniehPt5NEIhgxjfg/LUdznIRvfwwEpSxZCzghrTEPjsrTBUxkCRfIYw3PDLwxd
eEHTS50rSy24abggJgPUf+AIrvJFd4jol7tCb2bDHGfS2UV629ML/4m4JztrRGY3
wIgcDVELuWW3WH7hYuhnUuMfko966tvy/bFNKjod8r0ivRLYEB5UtfznyAGQ4dJl
72cUFtcwWo5vZYoa5smaX/CwDxNeQM4pwF0xFsohaqkaVnaHWAts6ojwxEE0M12q
3iaZFil+RD13AXV4hY4ayyakBZUDDTiBWKo4uE5ximretuBeC8sSWRe1s13dQABK
cqkz29ImhH45GkhgSScpfAKha5NeWIA5yLaHoiNH7aSMCH8b+PA6TTzf7XMbL2K+
jOSkKRC+xj5qPh80ic2eZKrhIi8xgwkJ/np65K9+bITMtoIMOMbKBH2p7rf7mKre
0GHXmLxk1kOCvcs6QASeHsYjxGisDPE6R/nQlX+69mxjs67QsyngpNYZlyoxPkY5
19xbx3afQ/ffu8074cKMtdDh0gvzqGRA+FtuQvxR4f9nY6Dg8gOlefqMu1I6pIIn
4xCSDJRSASVk2wKvFcFXxvQXRfWrH0afeUbAdTKel9YTYNWFDnhSx1HsUo6WQLJO
bZS7GSoHoOKupMGYhIgJ3lTJ+Lso5gsvnGEq69/c9TPSK6FcGy5gd+KJJ03TILl9
QnTAiz/A4v2X2XlFbiABnxKk02tKa7PrQVlLktvi9hsUqG0C50KYBWtqnnNBtYHE
jN+0SMrk12T5EJjTTTnhPPn7NuUl8tzMfS9ic70n7s2pgGjY4h+maoZV7+SJGmmw
H3e4WIamQgT5KQ/OV0BA12nriAj54U4Th/H/P4ReF5gUXb6QoIIomd5ndyYKc4S6
tz7hP7xYz8y9rnBCSur9k4Nv5TMO6IN1tgZK2XRTIk0CIyPTbsXvguEodpkcoICP
6OWO36dl8loW2ub/TE1uYcS5HOWJQ8F8YL6LWhebhsukye/84HmyTrdNKFHrgwvy
fPpPI1p8Nbh6dxQh9AelgHgl0yHkSJVzoKcZpX3HLlvKvk4PlE43/8yX5LQK2GTx
uk9nt877lQnjRRh0lz6ojfxdsrodhote0zBVN9L9BHVsV9hdr6gXFloQ1m0A4oE1
tT4rC8opOJ+Qc+eQmZRyH4iR1cQLdJ5JTfbfAFdBChGpQ7JkvG/l8XWE1V9PdihJ
l+/OblQ4G2+tsPbRcgbcvULuGyNN//SB2gPwvlMnUBZ3k4d3nYhbMdb95ySJRTI2
9p4vc0YbLl0c1o9B5S7R83mspNdcU7UdNJg+EflWTLRPHTxDLbWcPv/w5mfC0dde
rm9HcqOWWCC8DJJAiBtQlP3OejsaBJTLWj9rku/KsSQAGJqnm1d4U6QnGeJ7/fVI
Xzq3ogFQvOhic9MaDIYVPZLyAivKTn0n+fckOfW5Ax5fXobYLRHs19BpSgTyNGEC
X1J18GlBf3gGYOilqeEkjZ849LY65VuvJufWVBVPpTd8PpdbW/piAzJAG2zcH5pn
2UJ74FaFSe+oRMJW26gRbLXvi0NW4VaG3LnbXtmlxEnxGhY1eeRNPD7NGkQXjthr
vEuqvO8afA7feK0QiRE2KA98D83L8gkSx2zJf3d3v3l/qgAn/Xw+Oip3MYIXfubp
utzowURIg9hk1Uk+d8fAfhjv/alKoCvyJ6LwGSlg9y17kXfXfRLye0nXUzyRJo/V
QVA8iKYrVWdk9o/CeWaPuv9E+PVjIwdJbeAVYYimkeJhBNy+EFN0GRkxXNbZY/dr
tEvbfICAO2M++hNgaO6ei5oW/XBUduF4/anctyfBSJ929OBOhFe2GeZAO9+IhEfC
aArUQUM2zfU8pF/p3tHqho5FVfQIorHlrgWpvkca67v2KoPQCw4ykCivr8H3N2IS
17fzW0l7/YngpF8X1kinpCTuycZxBNPsO5TYU9oLLJabgyd5x8aaEAltA9Ij/FLF
xudWc8vmPVGARy45r5LCMBA3W89wgO1F6UF2mx8V+yB8KcVJL6Uio1dALZ8Ul0ls
kMWBGYd2BDgxznsyjR8HjrtBjA32gbsYINEtvumN59uBtAR7lfAz5pWdMGCEs3wo
DeesWjOu5Am76+HrVuuTGsjfqts824aJhsOzh2/NGA/qG2RZdU/CWBjO5oWerqbe
sYu+dcBpFT72hgbiaOdqkNwgCjNgb9dW6lW97bFrPxJ/wCv8vUzncMmgf/pTtHny
hqVG314wcuDrWdlhyS+8Fnq/uWilFeEa6UulC5EOMl5dkLQ1lfOYc8yg8JRMYNG6
BmJts59EuNWga1jKu6ngbQ1zguvMHV6YE3ZTd29BWiUAQV4FU5mH9CPvo/OxPqS5
sZl05ZJCzDMm5+OKWp5lgGSLpkgxxI3JbsgEpdu/hJdyUJ1nEc7UH3E0Awm7xWjx
jpj2aykQRjYWVjoPaLtPLaMlA/e17aP851xwgEKIA9CXkpUN9rCLx8HzjmDI8Sqq
QD2E/bp1YGIUeIeftRPloM6MdMZsaJ/q8njCcLOgMX6qh70XdBnbcPeXZNJ2vfKY
FwnxW6cAhXunwsjTWabsFwm7oOE1dw1CmiVRQAVjiwhtE69D66KKStl/1fltYm67
ny8tjRr2QPAhkdbA2Uo4Ts8nzYRtDXklsANt8sV8gQaZWB1dRHMeW2f/K6m5z7VG
oo+b4tNKQcLtsZigKqnFd9zAXBbuCezAD5l8lLxgZnJeMD4nceWwOt5rNMy7OoOO
G5KKsL3qkhtJ2agAbdT/ft9mDZQiiVJ+JC1ggYTl2qCYGV2ywH/3dP7FsYAkj3rS
u9isT/K1Ci2XU9hdp3VAGeuTSVVbciSMsCB/8J1+R3VRqTumLWQ2HtxPWT88dDZx
zLUlTkMspzrmt8qcfwR00DsS3YcZ/DDNQTMxbrpL+2DeOY/xao/Gc3b/iKMtNmEE
EgfG8jy1XSj6JEqxiM+CVojTBH6oTC2aO24TX6Va8Sz8Pkfkm1FvCQAQRgk0oV5a
P/hj3hOh5LbOsHErXVGPThL2JVl0rnaUl6K836y+nYf0+Lp5hoWEP1FGc3/jAo1A
4/Lmzl9a2uPQfYtJr7utDjTmGYp2pEknV/9f8GZGl1NftvHoVyrYLckJnwadR1cH
WisL90oIjw3vxscxPRp7ZMtr7ZmKlYPz+lSmqHipheOCoXfTdWo0Lsa2PBlF3EWC
YJbOahdNL3fqk3RWWa3KVwKY8wdtDtwJPUnUc/DY61ksk+pEGVZwwbuX5ECqGPt6
kLR2ynAMz6dZVIG4OKoRAyo4SwkgdpWCEPpmN84c5CjYZhQuZSAeCqNC07z772g9
KUvrPm9L6BCGRkQe8nbthgHjDCXAvub+PgfWwsvXcH1p4ABarRHGhxfd1ujh18zF
ZPKcHjpaPtZsy1sfYEfwed5JxASD9jR+9BZPNsgTw2Kd3AxizGcQ58n9PM6v4+uD
VyVHg0hdNVImldVCs6QnwnBfb63GOHJBFRXTKG1IxjVzPwXZubDkFq7X3Ly5fkxC
1Y8z/nmHub8C9d1xLx+oyIJn3msuJO4rnzsegpAsyd0HvCYCHQ6ltIPe6NlRnPUC
YqvP1BAKcDvlBv4dcJPbjih8pnmoaDI1MgY6QXWiUx6Z+RCIvEwVHh3cjIkZQ5Ds
jKWvZHw+RS1Z6TZfaC8QFnJgNi5iPR48XYbMgSxdhHDFhGy0HcZfIZBlgbxWlri+
bSlV2kwitVRIRVfManDpwFvLIj+UbeAhgVcJaorAkPEsBVD2A9Hz8tl60anOek2T
zfX7Ta89oo88xg04Q8GNcscZ70SKtmRqcl6YP4+g/OPzh6r4JAc36bMoS4eb6zkp
5OqbilglbmMbOtpfzAujlKPoF6Tlwnx1l/nxvmwEw2dDgcNKTBVbi21EyzN/p4qk
vR1BUjdWpj+y8iYE+Xv/DKcCpfziTCc0f7CSgowFMYsczV5WNs4g+X/oG91g1kRA
Xz3n9nXr67rjmnp+gM+mlWrxLFKxbosB75UWsVys6gZKZuEo0Sk2C9IGmdUlIp98
38CIRB2AqRLwSZCStFo34fNYeL8GLqsO99xAjqdgq0ke62Ei0TMEy0bm4Hol5eVz
irK+4bJfvofgufD0MAUGQus7c3/H4wy60HQdwMFfBL0gQkThAmhUjjnlB++bvfNu
pr1VRTQ1I/90JbAiuyKcHAOgSS+BnYJ27Vy1FXVDidnveWazVeAQ0Fs/fe2qKw5n
/frQ2lTVAvJCUC68cp6OGKJPiLN7Ldcu9d7hatfGCtoEFUK2ZJHpiaq1Nw62t5YD
RKjX5/JEYi+2228G4hlau+zIMkjQxpxn1b8DuC7mMEPDdSVuPU5wUxSbLbWp8CVl
AeXc+OuFb0GDIdlK30xs298DpmIA8e1NYFW0tn8KriGJmTdmB7rlInBnuxvHAlfn
qKQ8mReydgrJtJjeTiXQXRwbFHaT4nSiHLduldoaalWob5LO9nzWpRA7zqgON9hG
82mhZNfXCFPdOicoXtOuTXEf3tgSvBs1izlLdhV9oPgaRtMsX0Vz5xV9YFSEB7kx
ITWzeHKF1/ePG8lYq6/FronHrj+7F5+e9bO5e32apuPOQ1nTyZedv6snO1aiTiPK
xib3lOOsHtP4lujy7LcGfRxx48C2E172F9XSl2ABWeqqToBJOO00YQ7mZeo6rlzB
x6dsAyM8Nlcx2nPgHlFhjg3yatQPb8jgCHX/UspjBFGUhrnMulT51ubLJjsGxBdy
juSSjkYeByDWThoLMiOWMoeBiOq7IW1F80HKp+4JcyTOwU5LFB5JxHVAsjobi1Vn
m4h61kEeZYRYBx926ztQMAVrbM3wPJSRH8hIr9V+ikw9pBGFT0gENCbJPq1HaI0R
qe4/PlhZhnw/Rh6aLaU5UnZbfifjNFIGjRgji6qn6EYYbF7hAq4sJXDciwqF46gM
UlLDX3V/BXbpiWGNRq1gADCFMICx/UxrDghTUA2YptoXoz+ccABwzotkHBR2gUky
9OVuAr+1tx0Hn9ZuAdg7JoLs+w2rmLFaJLQiIeYjwf/PFlRYxNBgspHih9hOI6nX
zfTB6iDrvzLwRuN7t8cd8cuOZQu16yYsFvzYwBoz8AabT8pLa3X/vI2FRvbXdUff
dgFE4GCCCIiYROvsVReN9xyzdwBplMUDKrc1x1gdgx6PanGbL32zgX8ak545ZWaE
HbOP6yEgPaYC64JEdkPWz/E+cX6oH4VuQx8y6QAss/6bzCmI7bnHuROPxSEoTNBe
2myLhJyJHFVF+u5I7LFbFFuJAI8Y4cwxiKI4MEggQ+/5rowl0+IB7N1r860YHToO
VPBys6OT6AGkgH2C/1XFFR+9JwpadCKnA7IQJdqQlRZEIks5HNcAnfjEW+4s8RHP
LvxE3CFOQLnyMVVzYaNNW56OX7zzB0iFRU/2c5vzo94Wd233R9TYmHa1r2djfkgh
9Ew17uO2Uj7qgJZoTmy8fYHiT/XqEjinvkQgytgFVfW821THodcrOhWqmGG2XHg5
sJPET+pMd9LKnWCZKkv48JUFJ20l+FCCsym5JqwYoVa7B0Z+iLromA0RAdFpgymB
zIXrp1YnMAF/eas/eDTiQpBxTbKX9ww4uBP4KQ9tagAeOCnPPWcV04lcBDEicX3Q
Lx2r2Ba8ShqBzW5Piyc7qrjEGywPxcbolnP5BAjR96Dy2VOB88IVcsUSEiCc6xOb
xIeOcuJaEM1qSAnhV8ndYIThHnui61hGgBftfEZJIVIj565LVD+O6feF4mqrhch7
MBcTg3vjapFKtd/mSGUSf4XOal6vwi1n0rQwhTjqeir0IuoypIUAENLJn1UuomeH
uLiQOm4jhoDC5iKEjYyEPbVRH8cb/eEZxVQZMp6+oNmOM8pvCZ4QScujWxNfrfY3
sBt6wGM8Cf/85KOyfrL/B6yQZWZu/U5CgY88tZmVJ6l3JVIsQVP4PDe7RZvDpilX
M+dZBKxIoTcjy7zp6gtViSkDQmFCzgl/36Wlz2Q6aDQxkgH4cM1tzJu7E8gAhICN
rOKDJ8a72C2p5ToiLBg6TjUxpkFNMCpncMcAzhne3XYbp4+xXHh6DT/yyxcXNLjf
ZDnx09n7c/SxZMJigkQtVdkrtcDl19+kDFmwGJeIjWKfFWL2nTJbsF5p8l0bWwLh
G/EmUNIrQ3rjg9h99z5y3xbSwL+55oTG/HX78tcykFITwljI+c08HVlauo5fHrPN
5PWwuS1TmAcFgYvSXSNrcRyeTLnPS5n8WRCniYbEiWjeskQpnAP/MPUsFunTuXQq
QNNdjycsibDkfrLYYWM8lfTqyT87PGh4101Vjon8r81WEJjtReDj4NQnO6hRzuXS
9cvc/GB/Vvhct1BOLTHGLVsV3Y0BiHukLamQlEl8EGHz8VvSWcb/75nDnHyAg/AO
+Qtnxv5673aYaTCuLghhxRruiFNPh49h72+WMWmF1uKteru4innSgahCy1bhLCjv
OpOfkxAkNvNGjhrmtcsFG4Ki/7RO1Va/5hoGt5YGxHIIEFRPPT9BmOKGBJBma7kJ
12gausu+7vMeeS8YrCia6FZfDoGKG2GirXRCYDB66H3wWuNIQPZMoOk6ahcnIxCY
CIqvSpAY7XpZ1qnYbEiS7lUxZKrlGKJ8c5NqnZkEzABqOS/pnWLomMLv7IEve4hV
pkVPLbCPGGUCnHI//l3kXJtNxgi7mebvCqztqShUBLimpS7ztQapUrVoG9tjEgYP
Y8n1jl1NlZwBxwuXXIwY1t3CosVdsQbEZ0t/VZZBQEtg9iURHwW6nIj+XI8JXYKW
QW4etWaZwuPKOZDfGRttKHjUgY3leomXJuzDi/F9gcM5JW43cQmi3zNZ7bz10HUZ
TDpRdOgmIGqcAMTL1KRCOPHLrsxa1y++g+YmarDHsgfF3GSDoQ2/j/Nf//BzG6zo
rN05P+EtpK6u0heF4D6Q7UmJHH8IqrRZOu4nLxWbRRjkhLXL1DWUUdBNIO8fDFoi
PjEEWEwpUjk2FmlZxtzu/nywqDAKyuad70zLpDccs3vByJcqsuhxwP+nuyQcDwBI
jquBEmk3O0E1kZIdk1XvF/LXSeXL3tEcafZTvPrjNclrcjsM/h56iotWtJWNmG3r
WTWqA8LVnfTjkDZ9eCHVQOJ5EzB9CF/1dX6POuo7yVX7X0vZOztIKFv+hVbjsE1b
g5MdTtXs3Mz4zkW3wMG6CWG5wZo2UN69EL0tGxB9sXAmg2Yq2EJZEKlAeUV70eg5
emRxg/+2HB+bv5s7Lfdfs4yxyem0eY4+Ou6kM9FfeGHoD//8Baiox6oVEq0oAQsV
EGrR2sazRbJ4NgUfUeSEFe+jSVuvHZo3ybaSuTRh0gZXf2mpv87zQu+A5j/rY9mB
5+63CWbeA+RFKi6Rne08UIkLBgQlnkxkX7VTmlZsVOimoqT9iStxv5zDCvFnJJtd
/QyKUTuSED3mxgp7xLpB9HzXN6EPP6IH4uJeUsXkaBzYPFwCIiEKKmvWUrx+ldVE
wExJECL8AulCPNTEiBSn/9+ykAapRJM4PVJjcK5ilP0TWxDMPWFAlPc+BKRzpWJV
VJtgmZD1C9/ch1eIklo4swUw5yZkvvKljghTiV9aosiI+cwPu/Kl6DeAF2s7Cnfo
M08NhzQ6jK1CCe78fiD+6tlwrxwMIDMQZBIyHkzso01AyzKMxebPhMfv7dKq4+pY
VJe3ePLq44jY4stVnKtMj68fZTFL6ulhGG2ATVbfTa2XwvEUD1IyQ1IBQauvM2ry
zHmdapler5Ml1/g3sObrn8qph23MhBLgIclDKE98r/owFbLefWO83o6IF6W2FHI5
dWbIuZIRMss4lyDuxeBvewLfQkuKsop8dafnt28HJoVx6D1bpFH3TvhmUoaaKdov
zoKxXkGp5SWyoVtVEOVLWgPtVkyjvY2CuUHwcozJhOf0uWQMt+ECVdPXlgnR3rIj
HFR6aVKISr0NAzHW3cRidzyK7CoSGu+P/f9+K4o8mWpL1dC21lSUqUSEq37mI80z
epV0WRbeZ/joWdKWsKUDsWcoZ9GnMNM3Skl5pVEMX9sEHZi7v5vdP4j68Z55Vj6L
z7INtEwZhzMXDuwhp5u9n9lqrY2RqLh05F7gcrpY4UEO2t7ihvPnb3jq3uqtzNC2
VlSWN63eeqXYSlTrueYi65Z7OAbVqSgCcZbNLHPPunigNqo0CMtecXJdh2kt8RBN
SU8dw6p2BCikKb7Hcna9GGe/ZHhoLuZdY9I/USo7rtDpdrpuUdaPVNflidAzXGFR
uYJ8063nDTI3NDk/vJSH5jxmY0AD6CCjO17nOjN0bcNS3CmchUCm3xW3UD1UAsWI
XNHxwRhNjQtMg09i+eYTri0jztu1YRqT+9HED4rmgtn8DkRmrPW+1tP77zssaORt
C77Etd1eqCOdMv0yw3h8kG+qDtX1HDnGVytZoOwsHx9RzR06Ps2kcqaHJOMjMcZy
RFM5qg+xy9kpcLKgp20OVfc6ue5TxRqjBeh12EILTySvpp0tOzLYwQ1oDq6VNcyE
dWxNwr596YPPNvcGTYby9npTm+OJ4KtioNN/tTc3PDw/gkViwuWkxqqPlhWuZ/zx
AsUm93nADmKtiz0SrHRxkF16y53fHxu856CmnjL4im6lj04RlhEoCvq6cTlJ5ImA
5yzDlMoT8B9vxpnxJ/ABvoRTXzyMvhH4vBrkkNaqNppPAuhwlK6jnGO6mFsGzIgX
6Gh6xQf1qPu8ThWvZhUDP3ZLg+EJ1Id5mKPAa/kj55Tpo5/alf05DkRmf59hByQ0
ysdidBng3/Wr+cg9Iyea/gcZedKiiACFVPuzTFUDG3UGZGDYDcuU2fxDw7xtiTAG
rrDXutu6p6AjuCQ73gPJYE18vVHgYiMriP6jQtFZUxcPU97rPx2jPTOvoTN5+gHb
SJSMYKSbh8/nOflqg2UmpiD3Uuyy/iSPBeO+a2C5+M/RxcW9HdMJBtfik0aqJfSl
HTk4UXj9Yl3mS3R/WiFYG5vzyfE/IeXRSIKZ4Eyy3PbhDrv62qHSQLL/9BNV+YVf
DaBGOqHNgwtqJOfDZ+5cDOud40CJ5PgtBtiFUAbYSf1RUKQq9HmNEAPeWhXmDqV/
7Ge0FfkUiyhpxrXtjifPpQ8eCZsV0PxY0T9ZZApT2sdWpdqh6irZuYwPj3TVNlvz
NkgC1abHEm/Rryq/8m04XxidK6XMM0i5R47IKlF4g6Vh+3xW3TCMXbC5UguvAX4M
LS7tCHBVUAhhoIUVRoh41BvFK7LiyhrR1sRx9Gb0tTydtXGRKPoXWS39LkrHGlIk
va9WG+jry9l6hblDiTXg98c7/OdREWzI2V9PWU2BsV9QJCJVbtbB/cs5LxaczLwm
gSBAOu0JnbHFoGVko87fHIJwGieztOB+G+Zax6k/6VhCNYz+HSZvIWo93QIkmoLf
qP6yVCrjhoJTdUR58JWzwnu5datqqfYTEOG32rmwM5uwlh3DUTjjXYkKgn5osPVH
nGGRM9dxG2qm0THz36t7L1AWflOOctlt9ngbAk6wAIysC0DGxZf9p5bkL6jj9zH0
Lk7giHe7HsSN7PFKaqOAur1PBL49PK1VtHmmxYLSM8Go00RQRD4MNQtRwI6sNiVp
Yj4gu/IYlQiR0snxsZkdLnP1o0NQU+p5gD6vXmL5GD7MsP0+1x6niNE7eWWAKNTU
+7FZKnS6oCIn81fTbUuggssZ/Sbn0HeglYKwNkED750nRKcpwnFRaBNRGnQAN045
b5Ykx11k4e4z2TPa8l5YJQvW3nJtWv7bFVv18pFO+twJsM+l1ItystjboQPE1fCb
OmGG0DXafsFLIdiKDrhwHG/ktLvZAv5AThaWg3qi4LOYTYfhCSC9A2wXh4noVHzq
L6enADAaGrdKnrH42kKe6R7wMasZjoFjaAZxuhbvZVvgMGmYgxnRS2SC9jDuHDI+
VgOouGWxsuzhXLi5Z85DX83p84FhiZe4N8Ujufyaho5t50G/+NVVgrxa6c6r688V
LSHvtg/MQDVHq1OtrTcD113kUL2h3NyGrzAJzImi1vfQJG0sCy6x90on9NSRGVQj
jK2q1MO/uGHNNY+ERg8lXFHHzW5AdTyASGLQ6dr7rji05dGrug6M5z/qBgSUhFSX
EYibKh1x/OU+qi+z+NsB05ZPaAoquJA6Jkob+tq54XBf/jbXzuIzrs3NwwWWsMyw
zj1Y9eYKISMP0RJP2eDGaWSn6pHeSshExgJX4yaA9/2/owuwR0m2IeP44fjrBU7a
aah4n9MXqKm4MJa6ABCEOz5RfSE2GDOqvLRtA64tGO/UgaVyC9yEzxTJMvuRXNSJ
2INpg5CTt4CVBUUVM+oJmpr0RmvooU+trWCOp/5viqn8wbck4wADlcn53XjxZRbs
MhofzUzxFOFpo5BwqyDDCUrlEvXL8I9qG/UxW+dxduo33nYo09kY2n5eGEMe95ln
J1rxdKIsK6z6ZStvbHRQMOeAoGJDYDsTa69aFb5wQ+bzr3MNdEHS4zUFQVYdcb30
lvAtJLyGkIu9RjrPycRZ1zOBHD1OaOL5Cx9EPJLU2eRkKGAURs20090N/X6mu/qf
VZpbCO6/EB3eW0cCS5uH52uGnj6Vzs00lD9+taZAJhs2h4mh+Jo4CqJIEf9HkKZr
fInk1XDd26SUaPsVV+Jw85RZiL9LPveli6dK+KFVZdH4shioNpCVrzuwCpZPKEM6
MWBWDwN1paQi/INbWlFQtFDnpbPQjiGGasVo9jfT8tIjl3MKNgHELWVxl+RHfc9d
2DvulnIPx+QD2BBm+fJHWVobpJcejHcZaWlf956q7D0YpVT+3C1kxS/WLpuGxtoW
l35yCXP1NxG/1D8tgNzCC3zvP20Y11POuWJB7MgKxhvdPHvO37P2vLV2vZUGUKN+
0ue7hNW+6FTpHugtzRs9eI9OX2Y5uclEfPf5v/2LkOHJcob6TYScWe/h1vO2WtUv
3PQvRW+BaZ4EvC4WgD1Ba+Uj0Yprr68SsaCdj4UBfRFCeLIMYoN6nSWMf0//iesL
Nldn7bRlly/WVPrSpPsjS5ZUCLLwaqcUBGo68Dtv13s1lj2hg02n4SoWgZ7MYBr5
aLg7w4QBNBMIwTgb5z/hX2a4S0k3rwbpTeamuiaw4RwmxN+q66lhBblPhshguWOt
5DNgRt/d2bWXY7UyKBYi7hlFU1uzch6nfckd+wXDOUGOr4H4yfNzCPe++qUAB7GH
MqZqvKwiD+jnrl7dhfUXy1U4f1Niw80ieu0z+jvNaiyLHzfIY+16Vxcy5cJ9D+S2
iYLTLwKEvfVk+jUsbF66GdNDj8iEVgjNes4aAzT6dNpFZc1pv6t+7X2I7bV1fE0q
CsKI5P4Vqx9uEqJxLeTaoxweSHZP17UCnJfx1ZQAKQcpCiuLVJQXROnSpo3OdFxU
CFU/ItxNCCyXE5oylfYBcDu7EN/TOkHb/8QU9nYXXjW/mAbqSZxMHe4kxHfF6/ds
R2SRYgjTrWhpQmpdlBSdVGwGkbWAe9uB/b4ocNhCnKcu/iik8JUfA8zJvVbqmAY6
oAEJlgVkielU2tBW3yFWcoJ8fjlDRRPNkrh0/nvN0nNkIv5Qgxyy/uNHKja74G+B
xc6MQD8jF2Su1DyprlFVZmo9XAuARMf751j2xINTWZnjEBFMAU39Hjj1bmt0sTE2
oR8efWy/QOV3g6n1NVpsrrereMzzxAACcdw67uVjsB0KGtRJprnQPOEHM97DdPyK
q/+G6OAn+GXyydmmT2Wiu/g84N1w18I3RJwqOSO9n/JWk7iVPbQm+r+hS4Sdy9bW
/sqaW3W7yHa4fGCtaDV9VCtRVerBxv+4qNp3ai5nziCu0vcU854CakAGbZsRp6zN
mdFey8L/7yDBCsznKUpvnWu9UNRJGXgNLympBICzN+yR7Yr3G56B8jMm8Et7aFkz
2KCd3zcJjerGoZ8kFCSPg9oKFWRo28lI0dkEz+PZNeQQB1UE/BBJnck4n5yx0BXF
4z72g6ghtUE/FylhBncOyojP8SyvWejO593/krA31U7s0msXPNHcBWsKYDCEBgMK
DuOXrl9f54u+Waj2DRXgd7QYKWXJ+3d4kPWeHQddYn5rnJv+4E7a9b8E/q/rSLBp
WAIx7mxMVjEgBW4rsu5N+Oxbz3BRaaUMIFpFcp87oOiyHZWqRo8Id8RCXHRZfggV
R8v6JJyd9XRlE+sh8WdxHwcBotElr2AqOYIMQeP9rxgD6N9ASGTD17gt1gRqy05O
mGrA57Bst9Dd4JfcvzEEj0CsPbYzf5IGopZK5BHRxkNuVSVy7L7VazZnKLs2iO0v
e9CF0UHvtJbFfkCLy+3yyi1ZdddIAt1H/RuHDlI0A7mRXl4JTsEVmYrr/rWy/yKG
3gcgnHCwUlfhebgyAicqNzodw2HXDcUItMplLn25Qb+5gPk5Teim5vht6OuB75FM
QF+s7butXNI+XUfZhFFPAr1/ZqHacjpjtUejrHxyf+akUYgBLwGNBky03HxnUycE
bKCyhfJgqtgMmXN6j0mKQqvXM1YJv+xi8aEulLjvhUDXhtOZDSZYF7xVYg2VA9GV
ivwaSB8cra/QnL92esQAGcmoyGQOJcbv2gqux/UirFOAZBlpMS9WSftTDYD+Q//4
c7NtFg4XLk1qSHLOogzurDVkyU4QhSGb1qz3AM9gYURtrWcUAozffDqWlcz34Nbq
hiAMJFP7Bu+Z6TCmCDavnzDISfBh36eU5ARDhEp24Bf4tCh7QB8mp09ToCn0UkHw
Qp4xodGMHKzborilSPHP6KaCEoT9xQm8R0+jfzP/3FVe1m6woVuOqQuhiuHRGSNw
gWgt46R+iJaE9cR83lxEfXdoNVCODpIuafhSZ+S+ywsHHxXErUoexKQ3iwH/QnkI
DAjq143tx9ntlOrhwkI1ydlyMJPrkVFUkX+uu6BDsAQOm8fuO0KsoXSHDBkk3Umb
wlbWZ1Top8JD86r96Nxh5HpSLMluq4yfGf1YGxK6jtQJ0/3p9lXraV+D/A4UfFL4
6JG6IEbc4dU4TVouH4HTVxDZ6kyRtSr0vmkMeZ84xYfXytrLS3w8vaCxc3ZA9wqJ
LRo3Y24NbaC4IC88WiN3sKHqMmslxoB+LjKWdXHC/9zdeBacynU6pXQoqdkc2nxv
kFvBT2hgKGBbN3C0qIbjF1DuCksc5OLiayOLMY1KCCTSGtTAX8/35JimQBRJZ2nZ
XMYq7atxnl23psXNltU+GOexoW5effweOMSHmofeVIUcFFoRhD3tyCvUEe2fY6IY
MIpBMGJZP6fWtVpA0FFu1/F8STTx7Jr4r8BMiGeO+4CK942nXSbVbm9RcIsmdhwA
8zESh0OmrVkoLu/VN+ShGR6DVqtBY4y+tlDaXe8YZ+fbfpE01P8jXHsekdEfkqc5
pZD5SbrgdI9wm/bO7QYFuzkj2WgSRjyO2kAnF9c2ADaxqmZwaQtbQqUIBeaw9Yt4
BHBuMgaTXhwHtdOo07ofrgH6b4JpHGpPdq+yGJxfOkNT1g8ZzOLqPiH5ozEtf38v
XN2901RgeKeZzZM6sV+zTXAveeT2hYJg3hvkogiG9pekXd2sNnX7fBTpGCR3z/JQ
4gTxXS+M5aeams2c2lWc4oZv8xw2I7aqESaPPfutRu55/OnHVwq1IFf3IcyuFw3J
S+WKt0UiMAEYndvqdHNUE0egfX9VAmb37s6SvYowwaqR/fB+LScimlAyfMtaYREF
fe9UTlg+lxdwou8A9N/FG/zehvUFUP/0FPeABFNyFI7sEKUfFViUQdn+GyXl935Q
evTPLGeoyn0SAo4X6mZP9dz0GLRDP8CuJV0ScgDnLapqzZ+D/F38MPe7/9wgyGiL
8qVJYkofzqLeyBuzwcteILpEdZ4jGRBkMvinu3TJ66cCSjUy9OZs59rwJcWL3j5X
V+Kl0aJvRFEhTHzRTjh1At4lKw0GZW7U8UxBiQHXje+zQdOZFjkxJlABks006+4o
YuygGCzAeLFgnOezkytbOjV2f4fYe5JD2AnHRGQ8o+I4tgZjr7YWTMQCWQnwrCYW
+Xyu3lRdOo64Dky4smpvACz6Jp+gszOFzXXs4+T35L2yu6tEAjHNS3LI4kQuEjG2
oCjd0rxT/o/zYqOp9fIfyAPvBb+Br35AnrIEHMdVKpYkL7ypq6oBDe6TJydCn+nJ
E2AtjxXqX9lb/1LUk5R4EaWyAmUC+m9kF9JqorisoBFHop/hmHUKBhbcI/Z81cHt
wo9vcuxvFh8x8qITvc6a6oNUpf2E1qp7lNk9oXWkHmiDlXXXv4s35JUdEA3Ex8Rh
B+VVSXx4BGhCfadVo7SRIgcrUnrExD8Kr+9Dh9J9duUxSLV6GmvnwKgDTzjw1TDo
/sDJcTqQZgkDYwAiM61B+zkI+Q90xuPsVg6lWr0mtnVH8sHdSUtPknQ3Fu/6e5z8
3NI7CUZJhLKLpBNa6qbQ0FJveNhusfrSlCwwai0MPa6znrf8kGrAnEIVpYLW+MY4
KP1eULMQzMD3gLntplbg4KgSMpyyJ7em0nynccRwS7lkVpK4Dg7KxGvTszDarCWV
1AW/pYywOukV2es7epSLxFF28zQZ2iaaSHpRuNBqzLHNQgUcbQCutBV9Da3gEUcs
kIQ/3sbQx14AYS3PBYcmDCwkTKWjZH710z4h6MHODQr5M0PW7QUS2XN9B16Xjr8z
onAPGx7wzS3DPpa4pF/TQV0BXIoHbzXtXLZUJoaoMl9cWR4t9TKZHWX2L+BR2/1g
RKV7w0Fior/eE0mSMfbCXro4nuQXKNx7nRVf8PpOIQN3SS/b03O690IHmEBCsIuC
ZYNMhd30hY6iPicSuT0ukKm3RecfJ6fvRa00Whe9aCbEPGcE3Hws+hdi9mMxRRVW
vQ2ttoyjkQ50b3vOFC72GPX6OgEuGQfKb+7c+hpWiwP1Nf/EKZqKlaqs32Iqexn0
t5gAIfyY3gh1PYmbQBLl35NH/jNLNvYjuSUwzJR2GYMn/f5R0v+OFLWG9oGZZ0nx
8swZxBDG3bOtnpnlHGExe8v2gNRPdIUpLwQp8jly40x8QjaJjL9OJVAvmZdKeKB7
BgjvAIu/ZKykyRYPaLcIuh/pd6wrq9dtgjBiGyR2w7EOkXmjIvpjgiAi7dEl4DL5
dxzsO5xqbHKQlv9g4TVfGXMQH92bIFczCjU+UahphT1AMuqhEOfoH+CQbDSyBt/U
U2FJbbCSflgBUbJGehJHQkCTYpSDI5yWVyzhdj7N/t9lRZlpkRMmmLGrI+K7OQhi
1pu5ihYlSfJG82X7eHFRIp/jLRgUYDTqEZbSlX1IrLwLy1eP0YTIcVEhitegOlCx
mBefJ/FbL0s/6UuxeXszOCh3jIcJ0LrKcfy5CCspul6bxayn9p/iwIExz6OYOEzO
GqWcJpuMfeM7Yre9pGMf0X4VKMkPbIuzAE5UyDCs1jGZWLjfPC2JHkDKf49K1SLR
0xVksVbhVSN/+er2OifponLqL4jrigrdxQpW+Lv4/wAWRoc7ojMrzQa9+wRprIeQ
4A/KXgTspexDieJOsPnUlBpVFzM5/3Y6AOC09FI5jvwr2wSvarPtniY+6Xen/qKL
q6nwxqKRy4NdUm0Nfm5Hs/cvclWzVopGaPYvFgGY90r41RE1xVHFZ0SooiNy9S95
hw/swLx1WtaST8B1MBI++O0FxzR5zTkNfsRkjb0lNkX87WP99b3Du+poFrsZCUPi
UzAp+IDhnUa/c1LcUj3g9UX8UEXLkEJae5G8FezuKwR1vCBokH3gCJFdd/ryWby2
rGOIfG5h3EOLNVqBuwXt0nvxssUqFYh6VFOEVRlr4EwvkbTRXNelS2JdqaaBhwN6
xr+JyRdmGa4+1+BAsaym1a2xSmBm4ehPMNMugW+fCXEeuHowt07nlyo+VIsDRdve
7rJubKc76A/qwer3P3vqyLXoyh3M7+vRtVm57H2ROmDF5XD4aKc/4ERGCZEhl0Yq
ujPhodqVsQ9eZfb5+F8aeSIXA51txnpPVBPbQjxbc2+5/3+gWmYRhRjr/cxfNC6G
zDRD9CdZqjMQ314nu5wGGkqrraXLyOwuU4a7nfv6YYvCNkeneQM1RPvhlU8K9VMT
/u7O/4PpgQAjNcPTtn0Xb1i1JHlEtIP/rGp/nZxCVH1AYfuo8O+8C71erAaawQT7
W8HCffZM8VIZQK3rnlEtsfRkrz/lWChcgA/nkP88q9xN/q+r/mLBRfcwgBJLtb5q
nriR7pmBm074k9+6pBrCMA8DoVI6q8F2MqaTFyONI+NjAR5FGcy3bAJ8ODJpZc9B
q37V0vRwvj3FSv0MmITZBjGUQ+Ubf+VtjB19S2WQnNUy1SI5qcH+zjIBB+ko48aX
fEkNryQMwVaorUkTDb6A/rDZ9cUNpz4vJMIR65DbpBlg71rsyx/d/pdz8YxjJM+6
aaFsJWih3vnIOrDagBtNEWn1ebm3C+EcKj0f23ouesNYa+ZtSa9LSnWI13cdiSbp
xI/lk2Nfhy1ZhH5IBVAv7XR5R1MnTB21G9gwxuB0M5o8L9BEExAtJtPlmcer/Ips
TE6G5A0lQ1qY4uCtnlSAfRk9x5GXBwidRcWWh4YKttY/LYekWx9+TU/nUzUt1IJ4
SU2yAsMRzfard2AnSk28fVcINmeiKfxjgQz9ftGzKQmCw7ausoTM0BPfOQHh7G9v
KjOCdpHGd42oTJis9GN67i3/HIRpLtybhwDooJaYos/aLsQAS1xqmt9YGjMYcmAP
lt8YdDVulw/cyt2VXGJygQEhVJfmGKHpQs68+mc6zZmb6diJOp+iaZqra9tkKgbg
Kc29PgGI5WGN64d5+pQNJ4K8mgqavp2Ik5+xTfrwsCXyT+cBrYMFU5jKjwrUjyyt
PHrRwUWEhNIdmiByxPD9pTbujqA5zeRw2Nejmmbzkob7cvDrQD0eoUHZpYpH98oa
7j63KfeeH9FL/EJ6IUs+SgcP3jigQnzCm1QU9Sv8aTL6hjPfdY4hT73QlxcO70Pk
FAjXukBiozmp5QiQAc8tjUwcud5i+xBxdsJL9XBb26Np1JGlFN8FsBxhzvUqneol
PUyQcRcepVG32jQLaUB4IHK7tq0TnKlaeXxCkt5FkPiMHZA3pDg62IEZcAy4knvB
pg9diz7j5nDNxKyJ2wamRoXiC23q6nX1nH1dmojuNKxH/BOWOV8wWmXJJOeID7zx
1X3A3rlOrLp3HTQ2vDA4eFKXGHyg+Fdk+MUJrTOCfx7hGGy1fHHvQE0T0iU2+1+D
SJceZhof4rPqp/Z2UKDJVbK3/FcpLrsMfmjSsSsGmDgt1TeNhtddKn1olPiGdAti
xW0z7hg8UKMRy9zhE0+Y8kuAAHY09upSasqpZg2gQeaAv0Kt/9iEfRSB6xsBK5Tc
EleYG33lG6Kf27e+I1DwZoUrEwoVz5EeEl4+IT2UPKmDzWBhta8rnuDjN38K9DJ+
hqbG15XnwPfD6s0tFTH6T93SCj9q5QAGUx8kc9B2gFUV1yr1OsWYmEagfUsFTyPh
VmH1j02t9hxwKqPaAWQVYhejN1PaYJlCNImTelyPX15f6ahz2jX7DbID0G4dQcEs
NkUFkoehNngZD6CjU8W5bOeEn+YeBeTzLlo7I1nNNTRBmRmSAqzUGYuLNtjA0z9i
whD7ADnf4d17P2iRBtBBdZetQ1rXl0r4p9tFT/1EdYVg/Q/3A881/25zd82RhzjL
k/b7lstL98ncwKAlIOFr876GYQvL78RQYy6c3OM8KWQzfAr8hMpQIHE3nFSJ8GZv
lLW5Umx1NzSytVyoUpKpi1dIm/+HpgFxBxfgYULeeqR+PJ+0qX5pZaLBttozaTgE
evhzKwlDu/eiLYjYcjK8luRvHwD8sLQSD9wvRQvy3EfTmGLkTJSzENv0LVEz/wqQ
B6mnko30ZvNTKxujwB2hKa2ztiMRPTEHR6vLnoZWNBfKFHwkfgdMObdvtuC6cyqN
/PFGJKfjQ5KlnMnA9rvXUKXITvlirAH57eQzKoHsX2IhBPvRTQbp89Q3X3XQIEsu
mr0RpFktbkhqgVKhlTF1Jl4wNKe4dIbvmO5NYQjpSaaf5JYij5opNUt/kGi90hz1
pzwgLbKJ4vIrNubeM28wiCLUMmBTYCCHEcRUNNzp0I6jUfQ+ENyohLvagoY+MrPN
8qeYyDgJlcar5xITvbnTFEtjChFp6vDFZJ/SY/0Trd4OIMfm+ubcvabUBJNP2oyJ
qLKv3ujIEwT9dwJ0Kn9KkMGpnPfNWTx0JTSYfd/m0xwukS3MtIxy3yHwDDQYBRoC
mK52VMiCRXCpE4CgOiXvmZcM26keU8slv3TmwVukvIzJ9bdMfei6jDHxoZiXF14z
HjWqFsf/H1pfMdIWVo772Ve6yxEfyoARyBE4FMI29n3ilP7RVl3L8nfERNam2cfa
J1uEoNAuraMK5Bae0WuG2nQbeSwAtgDduY/yApSiFupqJjb3SncGHrQRk79o8QrR
Wj3v9H1i/TUDEmp/D2uYYJUQ96apS3xrccbNXKCuyNwZNxCYUF+8hhpu+GtPfgzW
rWVb61sNIp1bBKBbcLtdkxr2zXS/dQJ6Q+9wFVPTvQ5N3RSQS4KxfF/jdE2AOHMq
3eEtbseOewR1OxLUCEvf6oDrQ/MKnJtH1tG0oPzJaZ3ZHnXjo0TiswhNAeHItenL
riFb1ZZ0nyd6gcmIMUsVpQmymE1ntKroAF8VVNKOzE5lHEggdKmdUR2vGKN3zMm4
vHGIGF2QefwzbpHTKcFh8msX1bKRl0x6cvRIYs+SQAl2mf2ZJhTKEqWmHUO4AeoH
gkf8P+bhSjXzssUeVFIr66IV2ah3XSieqDDpYRDpR15PjR1wj6OZjvmsP/KEq0XY
hBJW7JldaofEc4YG9hN8Q1cjp6nuTUihsdLnWhHqXcTIi+Eabkev7RUrJ6JH73W4
qotQNaNGu58rhZx8Pt5eGG1tNvmiOW1hQrDFMfgNLzfOSLXlTRbMxFdA+u4iPSur
m0U6tpKItsRnNCn9/u4txY6+mU5o4baFXyDVkVGyEsOnnjKeRpNxNgeanKT5xjtk
m4PqGwrN6UpR9pOFVM0rzzTHKQWvG43Ow2dpWPKAzz/CnklrVi/SmMqAbyRk87MP
OZYkuCyogncpc7CTS/ZBuaO2f2gYBMR2qIbGO1q3dP9n5DhiMSNZElT9Wy+t2x5G
jJpS98jDyLlJ4c7E9Bg9kpX4WqqMuoY3a2cWktRdmuPLBZfT1dLdH1Agy4xuXymw
iBrmn3fsdhLP9hGDlAfTVKtkQzTUk1v7e4VbkCjXd1a+e599gLpYIrZ0e/C0zSur
Bk/g6FKrcIusamI/6zRh/GQ32lll2hFPeuXcWffRMG6j9Jp42R8COgqZoLEVJ1Qn
MaVMcQz41iNEGzIckA7fc6kzQI1yF9PtD2jV2kNEt0TneKMubVqTyQigqE2LAbJk
pRDs+022s4/OfwV6o1bHLPmGPOJEZHIo62b8jz491b3bkpHcbePCXgLn2Cpgy1XQ
mXSARtFON9xv3/ZRZTHvExjZt17nxYeNjORyuyspuElCicLhlDveIuZmyNyD1ZT6
47nncYbvrVxo7my+oUcFFihDKRTBXbF3hTE+xl12GJdFSfS4cFXob4Js3wtkvif8
QDz+5PHGSncz/e7ZqTrinnjYs8eJwkaR+23ZVPaEjK+HfzBAkpT8lTsGIK7sy8Mk
+woUU/e4ly50JiArSuyVLfSYgsCO4pwIoCK8E7ZOysYQsiqmLEv2iKbEmifbnLGu
EfsgRqpYvWXCs4JY7xD2us8ebLQpU3YOsf/GBLPih0Za7/uEWcrHbEskWKstTp5w
S/iFkdtzSDzeozWwgFPzh6OKqohugmD0w1pusHl852nGW1zcPKNgalvflSQeAVuL
8F94gt/1yB1yweAP5n2/7LIWZoMBf6ufBTeRdBa1086nKa6cp+LsEJA+uN02fPV2
s13r3JrlbV/za32dpPYgI0y81MepFlobhQKz8qKKqzT4/MWGgvRYP8HOZ9L5w3+b
73BEm4WsctpEDhbdepEv/ddnvrGBxp94NEIjqhUKMH4D9qXGb8W+A27m3fbq+KN0
ZcIsZRCysDlQh9mO3Fp6187btWcujabSwLMk+MAWwQRbcZtkjwHzqr0DKgq6/eRP
isMOnDAG0U4FmB0dvve1UA//IzuyJoyEFO+VFD6o2utaVrUF1eKTUnz9liRrKx9y
amnPTzs5FvFPQCGDY33sNIA6Yvi6u9EdvENz84w8drthEGnCzmB57CcdbthoEO4P
oPQvE4gK44FzBeJ2riKmuoVcdynKrotAHZwlSJ+H9msIHN7sJwwiwvmngwQJISsv
BtAVZStx/xlyyi1cvjo7+K/3WSk/H/Nstw9vou50fW7mKhZ+apgPerBdgc1+VuJg
3E7B3Yb8tYHZzKbtMazrLwzMCUrgqRcQxpmGAe34NDzQr8PsM41rNmvhC/4i0AdK
eLzZcv+N7kIyrwqs3QvO0UwsUa44FG++XQj89o9xPPR7gebWcNRogj3fuqx6dV9t
Mwl5bNzTPO42fmbwQBlSNTO96beHQUtE22z4q1GTXjjvPo+IKLir7OejgJ7QInAJ
+GAdJ/5rUxEeGwRTtwGGi27Ck3FqS6hpIpM+0v2FG0dZd5YV69DxazaKbfp9E9Dv
0hs5eiG0LsFwxmpLOsIrfEmqlBscMu3z7mxZuuaAcNGiBg6RkY5Sd2yhfGFIViIK
8QZiW5f43G7ViAUpGSzwKT4XOQMk3kDv4Te7j+ip9ZHYlcIbpLg/MLXDZ/uIKkAw
7KPxUgeV9iTwHisJiSOswtArA7gcH+eSjYByOR0jrsKuJ5U8rbRHsBlWEkG0Jjzb
WP32Y6BNVl3bEW2V4T1sZduR2rsrTzrtkbn1sIiACch66RAw7/G2mWa9qT3HO4Ly
jVMbjwFJjBD/6IWa+b1B9kvDfjIRxFzCli+P/Z17139yLWf6GbOf3OPZk5GFsn0I
IkyOhcq6DJoBATDuyVTa7B4SmLm++tdJxFl0k5ZFWzdlyeVh6jpU+qUxvyBRKgRO
VF7k0Q8AHeGGzQsYP4lhAe8D+BlRJsp3AK5Piv1MYrLsrB66PvnAXI0AcNsUkMPc
mwdsTSsspJe+FEidfUX4bBIeBCC541Rz3VJhDlfE0wMf6EF7UBhWx/OgSaG9X/pV
pnZoXiRdvSsAnX54y9RZe6D2ITb5DxyrZ85bB34WCbNl4TKNfX+7ZM4JGwVuZvfU
KT9by2fZjNfeFb98NQZuKFPNGq2IGtAYAC/lloKDMaJPuEcuOz2kHluumue++dx2
wzs3/UPQn6zWt7Y8eWp2CMblN245zOLBJzzMnnfkKTNsJeyfoeKLhlmu9a0WAbi8
B4eYo2ryHPPmqpEIPtrfRGE5Uuut0BE2r7Kw2X/TYa49MlNyraftuGj3JDLJpzWl
Ng4rlL4zdnt/AeZ1tLTdMHZU6VqUcWkOapg2Hz5EBzi/e5aCAljZCzScp9xggo9p
rsVKw8W+wc84vs9+jE6kq+GPUubJq9dnda0SPsqBGm7cnu8JZVDWrRxDVp1OLjEr
U4Y2Bdz4Ulh2wvweeYJOwxHd42RfidhYSeIm/CNukVS68boA8Nh1RiF+EXn7wQuz
kigYWl64Gi56+rsvxg3QMmptNx4SeA24AodQYtV26r0vTk9J+lKH3QMRCmtH3zV5
pW7o2oHgfOdJO3sKsy+94aSRjg0egbkY5mc+HrHWeAUkRKiXEuHO6Rk61i8Q+DWY
fRPdU6vE4G4/sHw15NAt9p5MMBY5feMcQ7ee7fPYHPZXLs9ibNoK3FO1jrLspfgX
udSu/nZQhJpteUUU69rrU9LNm9/nAaLlLG/ui0hFKeIOmSeiaU5hecRbb5gRm4tl
GRoR7njqnL8BP3mA9TQKXrPCcfvuV+ABiiNd6xQWvsTcXcNUs21dEBmYkhVqTD06
KTtrmm0k3DDO/BKgmwR6w8WrmGttXkBe9GnjoM7kXejFsRTCojSkHj3kbdJq3Odd
3NVRtobriJpyQ5uz0q2okAcwzroV5SLwsFxtC7GdOmeZ9UffOAuf2/SpggIAwRuY
LWtDbdzrWU+pOSrltxztv7dM650pBAAkvxJnBkNajmC+l0bRK88rRg01luOdlge3
jv2abV++0X+Z5hftVAPPvjSDSEVHK7M4oPaU/nzVpyKyoV4iEBqXpOa/P39BRlon
qwfw3PK78ppdo+h1BQp4A2/HO5ZIQsJTQ5NjYka2tdLZRR5WKQNP58zmX50FThmd
xorlymxiE6I1ZlnGvarcRx9fXuSKQe1QsnTUsnCa5lsiyXC9MkBFUGGeVVho5iqY
Le8OJO0knSOVI4bmbpzq/aORm6dyyFSYmFdtt0GoQIZ+LUHqTSUBrQeLJGeqob9i
7Jjp/ni9h2n/S/z7ZddMkiXuMn+KP3WxHuGjd6uJVsYpALOW/SRNPMw2LTRz6Wjn
DIQCsViHuSwFJyN4Qo+afplfF7ZkTfrAZVDNluZ8DEvk2C+h1gx2MY1SaPS4vTjk
i8vfdnlGNCfYInXt8PGlLGzB99wLDsr1oWDEcFaiIV8W6w9DHeAVOruoniSLhuqq
k/E5K8QGZbCFDdK1q+d6XUm/P2GCRv3Jw9OfBfU6qcQDtYfaurvlT1ZlMqX0LvHC
gHTVfnYQ2tx/OOS/KRLh0lbudbYY0DPCekZo1qUzhKgF/6ifP2ggZI3EzIi+Qyp2
lXRexX0M/9/1xryEIi3k34Ax6O2n0x+O8ZlKJfB4uX7CKU3aH3sZpNhWmu4j+4FQ
e+0D3T3XJ9Y3LJl6UgUHnSKjhxLILnJ+lrtS42ItxfN5lOE4/wSyc4ce/t0aySvZ
zKlBVW6iwHpoGjgKkfo+9X9pBZtGB1PCZoaoeoFjL8x30Lrr0X9h/+6HGnJVG++K
Hn8U55XeGtaF8qNPeHoz72D76w1f45sNZdGWpkgnjls5QDzJGpo32VLnrjdPDToI
3BM25X5Ca8bUb1I/RZWYLJEHqgbdekokF1O568FuUxALvUqglh4BfvSQ/uEnP0j8
Zo1oeeUICVncVk4yYgtINgjVuXEP+05CjKQ/lO20k7j7KTVxZL3lAcMdlhlV162x
4zt3ar1TJxg2Yjrang/nA6E9U9Kw3ENikTHRoFC+QRtXNBY4wXkN/SRJb1ZnQd65
i8/XEPTndVMsN9s2L1rop3p8F6671Pt7sO8BlbbfafcvPRJtP7vJH12UfoPnF6vH
3IHxR9s8tCwFO4F2fG0uR9535C15R1DnaPbIHdVsp8N89KjWlc31tXx7bncrxFu3
CatnDci6Ruwyg2E8TDLx1YbpCI11D+mVHQFNp47zFrwZ6XlB8pcfuFmRGhxALGuw
znxK33Z9G9mi2uNG+ztLMMhjbdPsnapLtKhpOjsgSsWAwAHPdv9aUA3Uq7liTMl4
0JkinnlOpRUTvXdfY00eVDG2bbXLZts/N3QJnyqsjYYa8AmOinSoLnETVz8cxN4t
CusaRVxH1n7yt5H2rj1demefImqY8KSBZcnaP4C+rqKTNVPz4hBL3yyc77Jg3ilM
4CuEXJD7KS4jQFrk0i5PsKSKJRHHuISp6TIxczYErk/cmk07ExBgcwbAYiDqpZvC
1Zm4esmRruk6ognUouqF7+DhsCi5cSg+TWzbzJX22nHvA1CIDjx2ATXIgg1ktRjD
sZ0hgYitCobN9ljyPbIDtBD0ruaZMFnuoDefVY153y0JJUX+1RPyXt+qhiJboTTA
MjX08s/L4Ye+ZFr1P4reTiuU6x+6gZBtjJEfkkzCmot7YafqOtYkypN7x8fr9UWa
Ditgq4fSm6bDVKeKiigNBYyGzHFhKHUJUOonoRPtM51y0g5+naWOagttm4p2cqsU
y1V27LWHyeMji6hON1FzWIdfGttvdMh8I9j5hqiQ4kzPIgEt0f6/rFp3+/ohGHkR
rx9dks97tdQQVXazN4tSivJcGGY53fT6HJIHm4WaWGAGPWyLJdMDztOXM54zDFoI
PlwjhF+hKnkPjk3d7ToVZWPTtfsTCnzuLBBmcfvzpfFGZTEf37DOaZKW4pCAmvsq
Byq+v3bOD+nGSapa5uVlRU24nNF/U+779LYfeBP+3TAmvEQWinGbN4Oun3Rqae2m
UxmlnsrUIrDgPEqylxUMh5Xhvn4DLVfWY4gRKZa8EqoNFC3VDo97/oQqoEFWYOVW
imtSGnPnX7IZjUCzwOGH0i1YbAMSrnZvna/i1KPbIrubcYRSANkmhibiDe3MNVY5
KX4G6oOEcOilr2l2qWmdk6FwLfyEvZ+AsA466LU26Iv/acdS3bNV2wz9NkmWB7wp
0ZjvZ+43Y3G1p5ZUnnW6tKvWZCTeLmrYSX1etKYEk7I60exA5dGy2XgzphEZqDwt
ja/OxtCuX1f+pGyoMVKpxG+jMY9e7zGZtdwX+SAX3bQtS/2PR6mkORBf2vZ7Qy68
rRiV/2rTd18n3OliqZpzgva3HfmGpTOmdYfBYF9Dof+18G0+qOgrNuryAOjilbwt
nFDDulawTte7+GFNkdZbZ5bqR4sbfuacfyAOP2iWhMENoUtowmMy7/qzPN481bpY
R47H6ITkucycrw3u8cyvORl6D4AVbBbk4kLzz6i7MMhbVG5V/oQfY0LbkYqrANQG
5cYj6AplMNiu7lPS7+pLJ8fnxrePfKWqry3TRDyZy9btXsaxAid5C1brJrL95Gtr
kt/ZICqSBYxoBRgKDBi5FlbSiesIEpYoqRWDkDbD3SsAhx8WRO829wC7kEhaZhKv
Q3i4wN0Lqvyb3EBpeXcDq/42pl4TPt3BY4EchGBfeaiF4XNek4pTESiJJi9nk0RJ
RTmeGSo6HWyJjq2xJECGIHFvqbZ9hs+Z7ELK9lmawwWCxpih797atcY9MJw1U/yW
mTFy+zK3LAc/5Usa8M0XCeVYGLYTO+5uYfWsCc7PhFNKhfENnYtboMSx/3HyoJwH
UEczDF7nFMYhPpWpfTDiqNQpHNULR2KjXiUN0XoAtP1LDwmRd6u7cZk0cOZGm43o
hl/khdSx4oD/gDp5BObSwzUsDAwL1aTHqYzmEsvt1YTfaISJLKuqfH8LogaspyX8
oa+Mcm9UCwXTaLEAJ6v3ShMyGhnq4qo1Oc3s2+06gfflCweghAW7abA62JRVqUkd
CoeTyIpwjLwoFJSXf5gSzG8FTldJP99dQZhotc3fWoaZF06i8VblYKfnYS5tgS8Q
gCjHCEfkOUmjIFoDrAQJKBgL9/ynW3GgsORYi7ULm5AuiG+kAFkwMQy5lFhgbso6
bNPt4SFqzGb15eKPa05U6MmZpNNycxlxbyR2ZS2FSZf5PNNTsmNaTUOqS+RGqWMj
L6jS0mMEXMFXrFqU+CX8duROCn3LW+ZqZcwAlXRyWBPWkcp95veg6MqxsoAIzLHh
o8htHPDQFCHPxTf3HiLAswDE0YG4IrsnW7iGHMNWxa1DSr2SvpY0SWRv3QQ3zC0X
am2EySdpMnEbo8wp2EIO31UMnHtihXBvdMFQ9tWyi2kfQK/dCa0IIKOIQ2oOWvDM
3Frjjty5sg7r5EKjHO6GQBCw9I08l1PoOseyAA18umeX7RejxclSMR2SSeDZ6qW7
oXN8ZiVzNNt0SG7ty75BNANQlt9HrqRH39/8AnKbTN8vD1mjiPANotOkiTP6Wjcw
fjXxqHZIdCx2ICYwDpoeLk89sJbrZ9exx6DkyFFptzX1T/Yd/bvx9oY7wHRQyYME
JLaBEEur4tPXpojNZXUh25li0VbpUAypTx8eOni8LQHdLcxpCbo98A79d886mAWD
AgP1YtWyOAJ36dGivsMluDz9Lcs74D2+BZS+NURl9p71mYBfMTc0VZqdNEy7ld6M
3k/90NN6CdoO7sYlFpfAV4oAMeonlg7yzj1wV5KrjOzJ8TF1P86+YUFpzgKCrlww
sIqQyU92QZ0yfOmdMrqrCAVF2FvthawiBnUKQAshdU1iXqkpYDrMdC1fhqN/StuR
JVMp7pmpBYcJi89eaQne5kQBBCHYRfphfKbxfg+Po4+nd6a4A5YOTgkiqGWCoXAK
8wzxLHDvTOCY+LA/KzoXRCa5Q/fxpmA4MbA67zCcAS8sQAF9R3YYdNInIkxhM+g0
yNJ9tQYkUKLYhSkqTLrrWew6mBuoS8yhlxk8CiM2qjIXdq65a4yB6ItJ6rsvzxdF
1GhOcaWyRG1W3j/i22RMdmo95+t1ccK7v6VvnDz3Y0893Hbv/ErnJ/WpsLpVMIOj
SgGmjLIu1KkYQ1IEVv6Wn2+s/0u5FlVfC1yluMIRfLTjZhrublucC8sd/kUHdkcL
klX8Vp5DKwGIeRcCi89smYdk7ct3z4/w96zKBaW5ziD+FGbmL2uNBZqKIz92VR0L
uyZjAhw6+SlXwjd3Fsr43yUX1wMbWG1fmq+eHD3HIKyu4minU2GaiOriGke4taA0
AfaZDMa1Ccdk2IOkL6Mzuq8SNmcpafgRuY4vwEIZndjjNcp67VHEX5rJlz9eWmTz
QsV2WgXTuF+DNQQnPG1TETFcCc96YG4jlmFVTHMowaaztYCZT0AXThq5KfQ5uyRa
vovubTEetXeoV2O8RZUHIs93VmRuqpj/zASC6ZLj1QAnWTIjqEnXQsT8X5DzbpFH
kfLJYAavPeuVUwWX0uDzu6WRQVEb613m0peDGOsuoscuDqpdBdX4quFuVc9yoCTk
K6Y7rG1TBX0t17fa89mgQU8GXwJQj4pPHSXEL+JsJBgIodp2+JFzZA0QEe6Aq/pa
md0PJuHyosRtmmFaGM8EFoxXshccwgZUL8FrQDRBJDNnRP+kcDyeYB3mLcA1zG6D
nI8YoJnQrGK7vORs9TIo4yWka3ScxcyN+FTETLeuwaIoPxURDasDZtfTvSthmnE5
5D3j4zrdhLHXy/pFVR+1Uzzyrpfz3kMhpICqzuhjWMFUMUfsKw+qxnsoU64PjQlC
b7axzCdHTHPQNPXcleHHxMVxX9ShsMKqI0mHNmVzfsjadRvcthP7SqRSda9ryIYK
Dlv7VmvPmR4XF4PkNgnrYG7EzEowwpu9T5Q7Uc4ETT20/DmmdcJp3qB/mFcvlTjj
stUmyMA7xFoqAWkOlSKloQi45lC6rHAdTgwWYaHCPelNzNT5pD3YTHNPpiW3xt8T
prq+H8GIWStLnOtEeuo0PuL/84nzHCIy3r/qpQRi9j5NOwOQnkcyppQU5tw9HidI
vFsdgfYfqYF8y2q+aT6Q7EyArv/c51TqjfxxCZ4a/HS5p9wcnqxzK0Ueg9fkRkuP
DukbconO1DuhpQxzREZ3HusbScEh8VMewAG2OAK1mo2RKm4/5zrMfrrDcHCtBy8G
/h2L1t9uAQE9PqF9E+lEzWtnsbBSltdlHfpY3m3ZoWXiZnAvtMHCxuKy8PwZwClV
U6Ld+HHtvjtYIoFwjL5yNwQVLlQds4wG9jJVghL2vz4Oe5YiWIgQmfzgu1ddwDKS
sMraKf3TCU9qsmeRD1OhCM7DmE6zKxXV1NgoOwc8U4X01XgrFqWHjZpjJjzrqnW4
u+8NLThTe/AaTyxOspidqNkktIuIlHYIcIXuQ3ecbiMrIgen5kKyor5FS+e3LVwy
mCxvxzBMFnNvBMRntqKXj66u4pj8ySwslYCEdG8k370oUJtQcNNRk05pKW3Lxhc/
vcekU4h4U+5C9Guru6r0SQ6YXd/j31Avgv0sO1hIg9rtwagyr9kR+LGN7RNDK423
F1VwSbCramvA4ZC9Mpb30BdE/EZH3iqa90sJAYK6a589quUuvrfH4P2vbjWiVPTw
6N5iTd6iPmXZVZvOe+fzd3uMFpSOqAhTSQv5yM9D2WXaeTKZhzVARr+X2nib+lVH
0go2fLWj2INzYQJnUb69K8cULy5I2i/fzFAAgCGtwq6cQpPFS+/Ar3I4v0nt1Axv
wjUMF4JcC7fHx5oNaYEuiG3DcOVsIoQus9qGUMBKTIJeThm6pljlFdjDOcCLl7N9
rUGasHPzs4dpdw3/t6vAGy5GAIcE5FvLBPs387oOSIimPw4IZqv2oijx9wWanXXF
8o6EgvTI0xCG+HE12wUzUPSOs6VC8oiLRXjNIZ5jYuR3/ePWRS8f++D9fZH0of0/
F65CDmd4BUIUATVuC0yho2MDKiI82/dJa+kYXai4mRcnB8b2zD5HIOMpRCAJ+muj
VI1xumvLkWAWfhs6gt+eyv9EgMFtqZiQlE6ZiETzp7PSAr/1luSru4IkGHYacIyD
Qs0+Z5QRgn+P5flsfMVFG89hDefM/nyKvXCzmtTBVkpTgUG8xwCgga13lEpgv+BY
iP3gY7trc4uJxNmfFtR4Rrg/dKPUr0g9uPWsm8I0i3RBwIVV6dQF/PJ2Rz6lTGmO
KSpXjOw9n8l4jIODJr82oKinxVdDDdx1vJE665sF/TJbJQ4bxF4hQ17MMmeG3YpM
CFMSR4zdXSa1T2vu5KkhKG8K3osjVHA4HSrwr+Qh5RHRXuThfOPpcEQmm6LfDf1j
xNc0EtHxcvIOFdQfiaOTSu+xCut5nqOFE2LWHsA1ulVkFh5zeQRREHAoJ1UYnUjG
Ur8+Jq/tncZRPJfVkz7HF2toDGAQngsdFDU9NL5RczoCMQ+hUL0pfw2fbwf364wm
hvVfigBupb2iuBB87IkpOmbV7ysmzvhadjxKTfdXrc8bYrZQ+s5wL8m6BMCtFOgT
NAA6C5jOfVs6epL3lBNP59cp9LVoHgTf6FBiSWgxzXmwXd5hNxEXo9O3S7ICkMTI
8gAWHm1jOjRf25kua8JBTGtx6yi2HYObPZhRSqJUTCsP7JFIO+a1BJYV6E5LNdQr
AsYaIUbV0s6Hiyjv+gqEe7esQDb/ZGs7hesaJ5pgmrpAYgVw91RVuiSUVeg4gMB3
NBwqlqZuQqA7qwmIxaU0sjV7wiQPGGdg4yp1ADInsnq5eGuFKQ19QYA1qgZ7wdsL
mSUXga4oQhFlDqFc3hTg1jDBDDhToOYzJujqh/U1xEUomIjBR2LpegxD7Rq30d5s
ac497kiBDlV1pCjdCLFlHkCsfh6LjHC/wV/B+w/8M2GFwjmkhqomAoh9fOxUlXmH
ZMhH98BeYIlUNwV3+5e5HbEoVhklk9VxDO5Y+YkuTXxWRBQZgl9bTGlz5T4R+GsS
2+S9WMqvh27dKRs555iNG9JNDWwRep+Vvsc/i/Y7lmAXwYeR9Phw2dMl7tAzWPa2
rPc02wlb0a4HKF5hrN4ZXSkU8rxItKOPoPqIBS9WoZfYWIDF+BjxiF+SX/r0afHC
teSUQR/safrdpbzYBgZQwTJRe7Z2GRC89sttaniTemPi08QzuwUVveem4WW2peHt
Um+JEl9IE2QDVyl/USry+JyqOt3xQSb/NmEQK0V3oZlOShHmQQ6I+A1uAXJNb6+W
uvs3+P3J5UgPhg00c9ejDl86/ShaFWnPhQiwzxxQT9UwGgD2PovaP/QTXCkT3D8W
kljdL55wN9Ljajg7L+btwQqJIdn1DPMXEai5q3WCsW8/6voHJM+Pm/LARLgjKDs+
jIQ8j5L8t+xUhwvM91yiJEaTkliieh1vMgwD8cdk2LCMoIROS4NOemmMeeT5o06c
oMclpCp0fAyxMwov3pju2Rs77dwQp6QyoeTcYwMzxLzU3ngVOROIrtyFTckjKAb8
crfHxSfQ9KFNwVUAJ/ZUjobyIicar93gBXuxog/cD3e74rFOHaE4QIsJPD7RqSpg
ZhXNmQQ3jCURvL226t27h9u+BygOJLFLxEk+0oCZqw8Q+jA3ZbcyQGMgjPZO2J9J
OwwZFh/177k/iRhXnrUk0ybVXVWlDX3g+v8XudoP0/1kg72ok5jI0NYru0DRambK
En+NlR7DU2C8bRMxf+AgEheSvVNh+qSxWARJGAfzY01jrNUyNfyjDrh/UxWfp+Sp
5P7/4tnieYwk/v6YoV92RH1i5birhv7ta04RLm52V9PqDqXXq8LuI2pm3Ilp1mo/
aDyvZrdqxTML4bJ/cRASK5EYBqs23MbxmYn7DRObxBm7+721TsjKNG4rtHvhYt05
dDJVmuI37/5vbaZ6CHbIiGJCPB6EUP5jdvcC4LNCwqbHZzRj42WPR+QZyJV+wV65
AMJwhCb+r0FqfOIrWx3cD1DGDemhgT1Ih8JLv6GD0Z2U4UD9cDUTaBCwswY5LJ8z
vhtYo0M1v/5731xx/ONjMirHpPqwiU9NBNSZmg0lj0ZFcc47pMfJNuDuD64sZR7p
UiKfz4JUncFXvDP15M+nsMqbE0v7NOAo2vhHnUspigqo6G7euGK5qSzgQH4Hv+1c
QxGNFsWSz10bFS9YFI2HndgR7vHyBH+Axw5lwBsAjk62B62/KD5dJWpWSVT2tggA
uYRNgje7o6nVK0+veJc8HGt/69F+IyBphZRS4UYsKkeZt9UmPRzZDQFTRSA58uwb
dFol7jHFOd2L8Jv+9D1g15M7vSM2uqYaOvIeWW3B6sWXuWaPfsVBtI6A+UdxM4X/
WUojVUihfBluLbD6Bp8JDk3Kfv/GDlaFW3O47NFuLrh08VZwasvzqai+lgI3l4VP
YhhPrsG3Nb+GN6J/hVijAnjftjQBVp+NjtlXVJ7OiuRo3va9T7UpiCDUoPsljZIU
qmZIMnCWk7yTb4zDkWp7lWjYKwFsmZ7UFUoPR58oaqd/hpQfJbNTVITOwZbHPrIB
kB1LmQJSzQBXsbF79Z+XVC+zdfoAJFXP2gT64KAV+BO422q40R8mQKgTM4C9JUXk
XC9ssIFHA6WQEuYXsFyXpdVm0F1UjPNyYrWvwURhp0RAvxhgmZss2NwU+9fh8Zf2
p89kJE45MNOGYRPxNQsyf8w6f6vQ3mMuVcgKYhI4LKJHhdhKbEDacvOyF0svy7Ke
Ry/kh82TK6DF11YxOfZQh9lRBf88HQCLQopBmjitfPRaROBLlmbuKAZZ6i7aSlkO
48l2CmNO6K8kx3JAzPORemC45wI06X/pn7ggOlmfSR/YCO5O1bvcxh6IbXbxMmR+
mxh5DxT/Z4aDVWaBsxItUPyVi0OSJc+sKfyuJtDUQMGHguBIp/ai3xMuUiIDU88T
xqpIV7DOQpSWAP88GAgaM0XrzBTlb8GSzo4F6zQIMXR0bbG6c3mTlnPDvhLKbUu2
kOet8UU1GvzsFQmEz03w+i94RYCO1x9HBi6Pt5eOxGQSU5w+sVRZx+vQHXLHAYBB
lnMFcpiaN72hZTKmGA6Kg8HLNhuGyRNQv2/HtB9m6HbgMNiYzKj1O2NklJaa5KNu
mLqLMfc8lyfagsqsFZusQR/rJ7mjeNcADDYHD+dfdX9j1OWNpJ2N3MVE+7MxvJbh
MLj6G5IRK5m/sRbIQxaAz5QsTmdr/5qfsOTdXnGg8x8Y00KhxLxCXX83hYkUuSBZ
NpFps9KmZ8zgDV6sR6hsvstrdfHeC5B/GqcZYBzOi/5JqHTRUOunk62T3klKk2Bv
fsuPq/UOZ5b8aX5bRurhiY5LOxs+EiCdiIyu0dZJxDm9+Fws11A15y04Gm9BrwGc
P/HJoSJszM1wZoxwcr69MVGI8yIy9PwnRGXqPs/rF8afjbmyHZDGOUZecsdLmAD6
HIJHL0qfUR6tlmV5jdq/wyATIT7J7MEzx92oKL33MH8AqU1gHW/EkF1e4BFcvgoS
UyQzs+5Z7trtw3TPF5YeLU0IIYqJrJ39NbwUdsQnH7JN3NJgHxymDbrTFpeXyjcZ
XBKlnvfW9fv0Gqz7GZsmphfquf51GWiq2Eb+L+Wr0o8WHjnKeJzDLGwjHjzkGRxB
3ZRDtyt97XHF1FJkn2D8BnFMVX86plkVaWKhs3vhJPq2yuUlQY6rmoJLEpvRZdBQ
AwJh/z9MfmLOB6wto1TXgOZqiAhJ5N4Y+rIzpRZ7Zk8P0odQycXOewikJ1RhAH8D
RCIRJ5LySlLWGlYEvOue2+vaPu47VZUP/kK9Xm7f+BNN+KPj4w/lye0iDjcWECEU
j9BkZE1ForNBHz4KIKoR3zMGRehZJB7eFgzP4uNn4mF15BxErBENGLshCJYeaOMb
1UBUcxc0/F35QmereZCKxmTawioUo5A/68FIv2JkxTX8Klyif93lyyZwYaKKEAkp
e0V6R6R+9wa1FOJQTW45A8MSZewYSqGeuDE3PqHCPoXDzj9Z2Rf9U7LRf4exGl6w
woU3N1AroUq/SiBlexW2JRctjRzORiq/GCiFfNYJXKGz6UlcmTvYGEJU26m7yMK0
W8M+2HDvs45XfRDxW7jXYp/tHjv7kZUblXvuyqylfy1q6ntCgMmhOdDxcOFrdvSB
P1F4Qx6iz/VvmOHvXeEEHtITgjgvYrbT9Anv2xI+WSXCdIrRxgQkksHeCa/lsbHq
6O2HvkTkn62vnfEtjUVHl9dWSHNU0Bgc4Aig21Rr29tBFvrE34y4K0r3ZvFzgeCL
YiLH8diH+NUlpYjJPjaVQ1LUu4mdatOXHqeaXkhJcYOHQOogk/hQJrcLIQt9cXnb
QY1sosQtLlT2ieezWIJntrtaVDU9bDVBSR19lkjGWpdPOuOPSeeUBnV93kgRyxp4
aHBMYFRLzC/9yYLXNTaslKejh79TRys3MbcjEewXBEDBs3IXjix4/AUpbzhE2Hht
mmhnqiQdwo5MFh2AvOGO6iT1yESLdRDZEObcg47E5uiPTm/3M+tIN6UCpn/o9jHR
z+QhFpvS+JX7ZIfhRhRfHJYPHwWy9muHn+q48a6ZbWOLAeZXvw3rj1G33thXf1iR
hv0q8BfXS7tKyGjA5jbmhr8Yyh4tSMC9h/nJXSYAEXQy14fIe4buWyokUpdgmo/O
fwejEyRWCiGBxaHhfsYZ8mIxeZ3oHKvszstEibyr4bbVGq3D9q8cUzl49vQIyH7Q
0hWu2m8kGP9EvypnDpE3NwK2XUDx+6RQmO/bCMM0Pq80v5iGDr09h31mtE97N1YQ
nnGa5bRuVNvjEeUlr37dx6nuFXxiXn9jEBHiiW2F2F6+we5tAhGiVlPnFD0GoKon
zEkEb36I04MLYWoh0KEDyuQcDZc6Q9uvc0NknEbPOj1+swnhEMqjeSSaIH+DyBp8
X+Cc09mjNaMzIWpQ6k2vhX8u1e1bP45UXz/obeTzExJOPsndJ6VeOUz5NWc7YKDw
SNyzktMHgKQ9CX9dlAgLUFkwExRNir2iAGdtyi5ENRijzyufgltTioa7JQIGIYfb
KB7Oljp6jNcwm0cMk2ztdZfZSGLtqb8HmkYcVk6HRnkNQl/y1fOAwEgaZefeF+hA
fwZitZ62cMAbvp4cnAEYOP7ClWCUUeFMPrB8G6lBIeAe/eJGmXof/miLZNcYZKtA
OW6nADR8PyV86LiCmxFBR9FtsHWG6eZDmUsX22Au1wsAhnkhG8umd9hR0yVK+gV6
cwO4eanK3C7fDTbAu2d+Jcay60WetASzN0Cp010NDqQg1IKPNHghZNkEzLKFt0Ky
DzOp4TuKp2BUGzz3qa/zUu6RuEmNUGN6RJIgChKp/dTthvMv6W3Mv03H8TAnrJB1
CB35QHu3S+MwlVxThfHYYb673JurkBIPzQ6imOdYEOSU8FZR8DyL2g6H39Nbhcv6
rTU5GyxGHiL+7YrKkRDvA+fJhPHOtiMuQuC7xLK2dEhcB6py7RE6bLTlZ0bzAKhC
6XvAlG/aEmJALkPo+dTOAkQcD64gVrtRSW9+EujpvCHp5/t5Hd3lTw9yrhuNbnBi
F34p5riiv6CdBbzu3BPheqplOgsEq47Lm3VXRuLwg5182OhconNkyodyrhMs/uBH
T+UsGEyvOSFz29kRTUWxla7AZzOmeqLXI9kTkLW7zwjwZpY+w7+5ffkMgo71+5D8
MZaUv70cFw5lQsIjX2Zbzikw0lSUTlamdvi2j0f6SjHghuYgOUuKSKV1HOO0txgA
0azR902iYwMobw8X3btUlyNmW+dYbXJPrA/PDV3Geys2AUZhwAlq6+jvOXygpnip
eGQo0zs5qRj7bybpLbD55+p88Pm38qM645UZtK3XofkNeDRqHsSXlk2sYYNyqJNB
SWBzfd+pzxpOMMCX3z/t/1YPjVlcer+sHPw2/HmLQT9qVL6ZgzerQNT1X+0joLlj
vEy2ffkeDewGUHHGiTfpoaRWkCv+OJuaofGlC3Lf1UWFU3JH9EQb5NV8mpaH3sIr
X0Gao58bS9JIvZfP2SMORceIdRl+NntlkSogmwfjZZDtPEbJuRyuSOI3lHO1ALx0
tyHR26OpEzjHVg9PgFUfOaxFDgRX/9pFkXEW47AE0zY6l6vL0yjRFj+p3+YSgz3/
T3BmMoYI+L0IuDV5HGZP7lvw2k86fRiq6ofcV4N8Q2Go/lsdhdkTUI1ob4xE7HFf
boWuRv1wYxIZjBMc8z8IlHys/atSZhklvyHH5pWQgr1dA8dB8pbpwI/sihYAYyy4
R8FWOrUuSgpDUe6IFs1r7eMIGCilG+omKqj+vhE4C3PpaLXmcJhrrQDq/e2k6QQc
WaxYaUTSGykiY5xO8vCybqsvefMW0z9SRQh18PZs8cQS6tc1kvN6AO5XqVm/HUAV
u64wGzWIWSdPsKM5OFoHqmwy1yxZ/A68lAXo8u8INLMVFCP79bU37SqWNEmr+Vx4
fblKfFBkgd01h4ELs4MAoHCyTfzgXD/+anj4ySHMxf+tLyabmcntGoRVCT1E/rOd
QmK67RizJmC6f2e8VYfPrCLK3qQKa5A3Qp9Vb/chA34bC/lBOJMooV09X4f1oueY
Axdo4z/AJq6MVF7CdaKg1/9zc8wCSVUUoJNOfObeTwvh5O38L+ZFss3gg0mjLWwc
s2ffnBxQcgQfHbeFSqgirFNkvjKixzzwtkqTY0+gQQbWAXgZtICIS3fz4iOP1lSd
MWzwv+yRn13YUv8Q2/rJDExGgybWwn301pAyBZBcbE4hr/OIiHjWG72c0y9L6/Os
iRzT2SQOa+PsSUymLAXT7kided9Ib80N/Pwd5phqiE7qO1oUYhLsgyBYRX7q2mVE
m5HI7GrT6ZEdoOObBAQYxQzHC5u/k6iT3edmpxy3rGeVWaiEexP47xkfXqZd/aV0
ui1eBKjMaXQ3tMUGp2CV7CYOSuJDy5c0kwC9RtcvZZAPofJRP97MQFcVA0LlRsuS
iBHVcRMDR9QVBQ7cvW8N1nrRgZ8iYYe/OT7CgcytPL0fhMzAkkAkbyPpfRn7BTv9
ACrIydDemonag5p65u2gu9kGmMsp8Qf5ZailSTnCWsXCn0rzbMajhR1HO3gUw42y
8FrPYabVTdcwS1I3JVMAb2cQUVcM+rpJ+3Nzmv03NC08rRVp6+mnAYt5z72uSWpI
jrQV3+2DBIlGn2+fmN2mezx+QhCAxXi0mTeh/pGncV8AnUDGbWk7grUY45RYboaE
nsc3OgOxqxvGWPnrsi1xOb72fKDdHqfATL0aF8X/5haKx35/IsZICnNuDFfkq4NQ
OU0xnY+3NUJWMJMcaTk5xvu4w4rZ/J8EdWJAdUwao/f9dUAzu53hQLqmUdMNJCy4
OOFOT1Qm3jYP16pEclrsYDQ8AWvS4xLhp8RteSLMZGHDlVKWNZ+OE2ytFil4HiiW
EBSRfr82zQJiKx1hs1InTT+9DPw+h3ksVv8opX3rl4rX+zv3iyqbUrKdqQNuzVYy
4Op8PTozIWB9+fg2efOJbdBBSqeGW4l8Eg0esi4SYXdYUbdz1CpPAlMdrm2RSJ4v
Q51+lrf+z/qs8makc/tVojTPgVG7sZPTmKSTkGyU18clF/qUFj6JTicra0YTatw9
Ew2/qufxeVC3VBZ9K41JAS7YEfVsmyW1rwwNIhdg10Wb440ePD/1XAYe3DpGQZdH
aFNyWMUfPKtyBdq3gK939nOjw2JkZCDBWAX4qj1GnKUjmjPj5SuY9pMT69/6Umnm
e2a4GRtrlC45A38sZzBBm65J/8vOwKhMyITU3MiXJG95EOVGFXC2n6WDYQNuH1EG
hYElfqlsqpG0MS6H1gD8bIq3IbnfW9Zy+B/Adlcc3aameP5qGTS4PgkCmqr2P53P
Up5gpUECYafo+gIR5Ok4hUE3a3BFm92dbqyzH0dT5rZO3ihy61Z0nuACzUgOSQP7
qisq24ujGD8uXfTu8UogL1StF54K7MAYnxEXha6NbsO8WqFKwTPjPFCiOdC7XTb0
i12HyqtbhwoIdUMnp7w7tx5zcdTucrQbxzzgZFkOHXXaMbbIKG+fhe+t4j9utV1H
ZUNU7hwp31rYJ3evrUGaVI84zoxGZTIoAgxlBONd860RgSnUWWASNRxifYn8zvIe
W0l5fQRXgmzS/dACLv5eMHMANd4M+UUS0hp78pXJu6TwaZozBKohRgbwTNgo8Yoa
sbxOMpAc6c+1YrBxL41Ga7y/TFdHepdpb6Q6Eysqd4K/g4vyI9XpM59VyyhbguuE
R6DvFixSF2t63jN73HpGZk9PysKBZwfbD7kewIKXZq2Apu+wPaQDWtYyEo29BFOM
b+5/+STa5IFuR8K5sFUmnqVmM3qwlfvPtS6wp/012pTDcR2kzCiZiU0/yiotL8u0
KPT4R3vSCWwGDm0rwipxB7TQByq1AKEe/dhC7pvynKVc1P5EMRbuK3R5TCEcc+f5
x8VFEcMYwxukUYCvls496ecgscDEn1kBnVkUkM7OPg5mh4yTYmfJWClhTmSJVaV4
DVcITQ79jyTA2MHSEpIAP65jUZON404aOj2+pVB6cRnP5INOjAxZolpBmCF1Lmwc
mU2bUh3hxV6ljdm07D4SlmrEiFYxjckuQ3wKctqo/L75doZ2aBnUiiTpANk1p4w1
rDelYffXvMEgYz2h2U382my0miCBf6wAlNrL1txqmbmx91dFDVq9bJ6VjyTaoa1f
EZtSESn5K6BKIkwkNGbeIHEDC4g1IXKYgwgkYlnUUJPFCCSErH4n5vHiFG+Hxzec
ghZX435uqQ7rRXlyFSafTp6bffiZNMTWTlAT0gl7PqCKLQP5BHMxC9k7WDsziryx
1yVbSE15aF0tWzDzvJtMbjhDqXfGd984ccpeQ9qTpSEps7D5G2rrfsZAaiAuPK5v
T1ER8qo7iTD6HONfzff72zdFxSI87a4pjQFlD6HXsgB0jSgH2iRwQaJn77mHQkeB
IlXNC2Ulue3kcL7202rUUmeiAfHs78Bo3tCB+VhBsl3CvJTpmcb6yryivqUAtNOZ
Wqe9EJuP8uwhCDMEM8lJpVcRULbnqitRFe6vGlFDJ4Edl6rSngd3in0bg9jIr9r9
I5ZhcF53Y1mt3WV2NitWcsdBe2OhillbcxCU6wy888+2kPpd6i7tAf0RZ+yVCc1f
SuBWdai06esgFz+H38/jZ3NfYlyJHhgR1txIw/SgxfvwKRvZDfZDqC+ccew86s8s
qOI4I2aHoJm1wXqlNFYTGV5iqoSsALgT6La/BhJqaHZKlRD48xKQyKcOmU57Ihar
qcB7Fbjhj4BgymbFdbhH9r4MsWYy3L0TTu2mj92O6jrOYwG9GKQs+peGS5+agy7F
UnkGMQdqlBjKVDfF6lY8mtR0bViTI4LMQGavlqhIyFcX5Atqb5OkjetFdASFmiYZ
ti7H6LmVJOZXDn5ykaXHHBvRDlsCJCELHurB9Pmvf3Kcm8SL556aH6htcraNRJI3
EOncA8nr+1X0myxdUTrjUbXn/ItDQtjrhuMECoLcd9KJFOI68TTAGdHBzewwSrIz
k6uVBS5/hr7uyo0lUq0790jPcB+r9l2c962CdUigWM7ql67vdNbPj9Ihk7WjHhpi
mwle32T/pfxsUSIwzZJj1LUPMvwB4qf1bOqdDmF0bSW1JQMfNNnXb9nG0OExEX4t
A/t/G69H5Wq+5MtT70htHUoyxCGRLkBPwANuRdlmcscLOF1/E+icB8kwbnm5IutP
HYuRQyYOSjNDrZZnB3RmXALIKH2Jhk97s30yWG76VXymc1gs7N3eJBY0MBolr9oX
0VbbJ70IuDiIJTUsFTI13fEQYtAVkwTyLMvBV2HXORVmISy48R4GHWObMiYNzpCy
5iTOn6J1UO00QjNRRoli1Ik23w169mRwBfIy0BVisAOsIhl6VATVumq7xqqHa1Ah
EXBV329xxHCtOo3oX6PlO+dD4+K8eCrGHJNrQl80LVFlNFvCSaQchwNc974ufV9U
ghtEA0DplPzaWJ1eQNYqbi0Gj+1fzMgDQ7VX0P/7G5sOy+EzPL+9ne8zySiw89NN
3GDsBLhQLRpwdhFYTSWYI91srwoRbBtHb/U5pNCjr6jsGd29IYCuS7wdq1AY61E6
UhMaC86XxPPlR8r8tgjhP1XJ8Kz/UZuXJjCFA4xugHl60uhuZI6NQD2/6qGo1ECs
zFQSppyI9IzarUKEbA0FEs28B/2zxKUCqv/a9Jd+lAc7eu3/PGHgrArkRs6mCzYp
ZN5c1v7AJH2oNlcM121WzxwC5jcnct9veOi6H5TXsY63cKeGsqs7V0NVF2S1FZgv
VdNsx6gv9Mub0VMJVQ18xDuvAoH7Z5OopWhcdqjO6Axf98GRgQHKO6EjMTa8NP2i
sSn2rrmbb4sBLBzZBMiNaYHn5wNy33YT6dPyfYUPViCmudhEO5aolAF/pJGdpI+v
mKrb3lPn87p7WoCaHwRK2FlhVIsvlKRXKjpEPLVju2OA2e0I7oZSPy3PllmmIHs4
F5eOa7lWFOyFRJKZyrNlDhfqN7zsGTuCIxg6RYKKAPUlMq3bff2zEOWW3yHJUlXV
Y7hwc5c7ACnsvI15h4p77BP7IN2Ps4jyc7VCJdTvYq9wPaS13EvExaLyI5LCryU/
fIhnnOi3lqE+iCqI1UfT1Flgx/g5lMXWQO/VGMJaKDp36qEM57JdckOL4uv51SQ6
Dvy4vubRg0P3VRU/z8yI5iPDxsYwj0SxZF+AoDRxZdbA9DtIw6Po/jfQN6ea4giM
DaM1h/2OricUhSXoNzbElKbAHAbDJIS3gFkzotv6qefW94Bbkk5XIjprYzrWe7fj
B1MvJ3wqbOsZF2S1c49NlmmEDSZYv2RhfFDYZNub08N1zkAUP3EdXjQod3L02cp2
Kdw9eXMRd9Iqi8rcxNhxFS6JMbLeGIp49xRfPtLQrWtHByyyIvT/CI63T9uxwJc3
pFBSQNPRNfdhK2MDhK/veA5Qw8MhMBqm+623+dcGzZthvJ499rCTFI664ZBKmLFh
ih7cpQ6y8LQqxcDEmraLhhu6gXkQSiS84HS5LZlNqCqBK08Q8loTqQd7A5ha9uWE
t+52wT2vfO5/5AKDkLm+nxMbY30QhniD3mMqSrcZJl8h8Ceq3P9TNVFYiFPA2uIb
RDuoA3qQC5VBND+1CK05HyFvSgg8NKnST1C0d2sNyuY4nszH+xNa9s6Fm5HbnwFp
vUuPZjRGuqCKhDFEQAI5tnw3tyTvG92meMLiaybG1qJigqa4x8zMGiElzJlTZCwL
8sl4f5A0G43x8JRVT7fCkjIW1j/fVvyaWq6sCsc9AwKpfONX4k98gVKtLtQf5Q0b
vsmtsfXC/5CiPfTfKjmj9MxMCcQCZA9bZsWEjQxYQreuaM5pm01JhYl0HA/A4Ud5
UFbzkvMPwS1ioOwBiGGIL9YEMZQoy2yt+XodtvFMhtSonBn7WPpIlq3oWUcvikov
OV5DBGEzhdYoFdNWGsG6loWtIh9TB1PZdXciNq8pTIyuL7nqU5RMKeR+ptuOF/AD
naJISe4jmssZaXpqIk7H+9LsH8M+47plyYw7e6zAQK8Oqqxo3v7IaYtSVZMZX5AG
Hl1gAk7MbJ0fpUdSObqKNCml/dg68YfmtdJyYjb7eVFTwGGTEvFD1kEbttalb990
GCvra10a7WYWcWJXI4SZs+l1K/bpiVmiFvb8sN9l1tT+9yZhgh6AkJ4D1dlSPULg
KLo8czhEBN+6g5VQJ+2ukJEndbmUkUuPZfisOWZu3yeDErT+kEO3e5rl9Ud95EG2
C08VUJc4gDx7WjFeZdC4YyVaXjRsCMsozBmQr/xsTs3FHJ9Z40vb22Kq57RNu5Ok
Cro0Uw4qEW0y6IpuZHUyxBl0uThzbiMg1RxckH7rjL9OAmcL1e9i8fqpk7+NuQS2
FmvK6boaoC7j7tMsdBOdA1G3CBoQgbhQRKWclx2aACkEBi5CBwLHh/AhU9+Ckw6y
nlePqPK14stbGdg3R15bPgoN5ysgjMoHMv0CJ1+rktGHvgjqL6TmM6TQJa5JTbuZ
k0vmMeo7GAK2bfhDLtYRmGst+Ex31QpybWNdAi2+Vx7AjUeUNbOSt7RAXLjped4w
BnWGsf1oUeWGmeGcqiluGy8Y6Oz5EHgbKvvn//VBdCJR8y29fu978+cX1NSURhDv
IC2zghPBisXKMk3vtdZNsVUyoxuaw+SW0lS/3KzFwy8E5dNW2bFI3vUR3pq78pzd
lmWbcZJsjcZbs7AKRV/nlzx3hCmymiCjZUkPnd5Ealv8TrKSw7X7PdSSArdjhIEx
+Dqt75cuIrXo180hlU+NSRRm0AOakSJj7hN4hg8dJpBEv5ZmXOciB0XiVTpdl18F
o6NN+DEKsNKlpT8tMgLgP47HpIEAqIJWZBPYQBUbmOn0TiiudFXcskvtk7l1fe/F
2HZSEIigLz8q72FgEPPic+1xCJevZ+GepRb75sYhgu8Bbd1oj4PSvdy0/UDb6Zvc
r2OndcWsAyN5Rj4hMsEAVyNpOMf++s/0MKnc5GkuT3E8nfa6UfsXNVTXTuDgj55f
dtRYmHoUmOtxfDwDDkyY5S6Tloct4tLY5SRiEYONL7cXfsN9ljVYmHXtChajjjAO
4v8xP4TPxwF050W5vRVhrj1bqqHbBvx26IAXZ7yaNm9nV7J9M3xVAOsX3EJa9z9z
UBg/BNJuL/MI3DhTT5iVJijP/ZslTn0dSFlvQS/ignTvh7gKZSusRU2te0D7zbF7
pojeKGgLNMkq+Gm81D0n6SSItXyS9TOdVmXrtRDbgVGOg36z7rccfCaYAonDTECC
ZBabhq9rtUO45nwdH5L10Wp2LrnP3HgWBpzNk8uZ8tRFuKIWZ0MzGqPK08a/aSJC
BHPokvg9/4erenKiefcjb1lP0uydeniCL63X5YVKygj9zLK5z3xbIkPmTEMq8HX8
g3YrLku9B8oB9yKZEBhAo/WjtOkiTwS78DkpwLybf6k+Hy3hQg13RFk6wbqC7Yzt
f/ohwLkPp7VQOgNbD+j45ITukRunfKQZu9rl77LNYZAZF3xOmYCzQkddLqYQ1Aye
kRe/V+K8NO7PLSE9LzrDSTIA5NkTlTxRjk4YNcPSKr4yhZ+lMmo2Z2WtgDIJ89mx
KBmDp9z7O3lvVXEJbk33iKuheMfwv5CW2EaMJIBGHqiijEl74lIVpWJsTttIc5Sx
8wKJcH1APLwzWz8tj2+Z9ZCoRQI8XSVUL3TCvGxSCB/2gjDXkb/yq7fFgG2vo/d1
IIL13Kn3A6ft4jc4F/YxUFrWOY0tvwLwgCMOe8hcisaePhxJkNXoobRGEBRsjBxE
q0FNEeAR34SaTpuzexQCerPvNmq8yYnOCFZvC9J/yyDC+o8ajket9cENJmdVve6X
85roLywhzOMZqdAaLE0MkJFrF169WZiWa1xHjLu4+AIdy+uaEZUde1yZ4PCceSV0
gXKuSQZv/ljil1gL6aVP3jkp9vFffh9qoi9Nf0FJMSibQtcqc4fKuRAvIPBA2hau
j9A/UOVO0Dukvtf2/S/4UQhC06FAyBBCJ0wetICAa0Ddo5Cl8QBLWIIOA3vU5hyJ
APP6zSGSgztNMdAvC7xM010m8WvpXp0keX68jhqBWL5euAWHORSuxRxqpB+ljXjR
AKz5jdfbMhfIN1h+wTWbO4Li50ZJjK9PMmOVYjyefc/0nFVJcBaMW0qr9iSM/tl4
GILiWdes37qKFhsg1B/npJ3XlBUMSTs5i6ocEnHhS1tD63s0kzZux/1YjDgnxq6L
mLIUmzDW3Wqwas1UPaiFd68BAKHBq504d9VQg2ztolZ7yyKqXAhxq2rsGU7M37Gu
GJIqGnR5tUVtqAV2yvTIVG7bDZbi0RrVmLiXo1SLU41YP5m2Ec4kapdrw5PS1o04
MZVn0iIkJuLmMN03/3ryqDIpE3F9/MkM2UU8sApKTHYieAvUDfa+J8evjYBdp4pR
+TC5TDsTxFD/7444jRdYKsotdHFkNyEmHtQYJZjyAUiHwiwglBPs+TVk7MRYlJq0
KHTKnLCgnv3FPtMtpMLHfdMeY7TbOJV/DxX4BGqCELXvDTIJQl3a5BjRFLSCq77h
AU0weVGUDDB/yMDRXebqQ83OSkx43lxMyhgKUS71TvrdzX+Ke2a7wUUtmU4BpK3A
+9/stxYo70TbTneBYWLlK6U6EJakrsDC1TNOhTAjA5bq6l6haGS1j0h5qo29PP2b
KrXSyYHJ8cT2YGuLYl4gl00S3AD4H/R7a/pi0duYSDCkA3NpomkyXmK/BqNB+J0x
rIrNO9SeQoOoiNfTb40O/Ry6HTBGP2MQKwxneqOwxVs2lzfVntWqNmy3rEFko4xv
eENoyADtpB73wPV4KDaQbzGXztllWvkcDByKUQWRkpet2beUvzAI+SdcNg3y5EUd
J6zxSZ6O1kT9GtQxpONvZzcNEYNFc/u53LEPOhTRSFjIZVkOituF9I3DM8xqp4xE
mi3uJJwlwuzF/EJqOhmLjqug9Vc63cdH5rK52SuYZPujZICNWSKIXYhjUjJxVQUa
oPXDVCF8+1U18wlPOU5NwCl5CRRW7BpsYoyfK3eK1j+yoIhX6ol55uA55d0jCKzU
KwNMQvUOvwjmFd/h9gSot1CLXfwzluCWzBHuPxiJjWNb1Ppn3rqgmzDNFY4zFtXm
Cj7aV571eKGnaVFYs7cp+IHI7cT6zMq8LG4CZeUB7LdeXpiS/e8Awf2rAV8Q/foP
Yr8IEew3Z5JT8zz0lloU/c/DeXK5tp0iHiBbU3Ls2Rl+NfN+S4VvvvmArSfHP3mh
LrYmUbcJ4UlrVWvamtz+phLrMde/4IqSp1/QpbKtzNk+TJOAD0PS2XEeshjTQhP1
7X2amaqT4lea2OEByCj9PlxqPCSTEsTUMsGCmhLrAR/fAptiWjtwPmIbjHf/N0Fk
nkiBVej2ybUBnEUCcnPGCsrP/fvt8xiXu6xfS43aKYmY+BlIgaEixsHgfnu5gDN+
duLLHkkJRk+WROKAlfLbcZU29vHA3sXot89JVWad9ZO1GpGH6UV2WA0jQ00Ub9fB
cCDaZkljPe9iOqC2l1gUQXCAtqxIwaT4TaEorYbHa9ZuMajv2wx5ZWqTL5bqmJdA
3kLeY52hlDhkOppQ41XamcLL+/FfTT+g6m9nfLirGupPRjSVVTIhh5bt0H09+b/Y
31DyOSO0zIUvfdLglG4tpFBR4lU4dXau34yDBe/p0ab6wZg0qg42bD8a19azSGiy
PmqHGp+6PwqReMcCY9YsLiQvwluANQ0XBudPrh6YWVEjz/7Is6vBo5VLDbsEVGZP
5kfm8bahLQdAa6i2mkngFW5pMpDOYoejUkCs1kj15SMHU4dsxBZ/dFSgoNC67+bP
1iiW3jpuQ5QKotrQQ6f3D0G4Vo/QPPAOg1Oorke0ANSkoovBBbwd/LgvOvzW3Mk7
J3ilR4KOf8IvGM6ZdHORsIHJVB/+Wx/lmk+lwGxw7wBI157gGxzbfWS1fXUOXN0F
0PU2dVWVGt8PWzi5U9P2XqVGM9g7KGnwaigeGDDR8xZsO1W37IdR0i+S4n3esTgy
yp8fAI67pTK7e82s4A/lAfjgB0Hw9tvepeV606as3Xm9yd0O1rGtxQ5g+vw+U8UH
fRUDDkUovn4N5bDn7BmfFjr7GwH/+oFoHpvjVXy/Ey2Y9hDkbyijTD2vcM8z/9rl
ZiXsNG5YebhsJC+ax5G/mPUmD+fJTdnS7OHXYUT7NQCD/ZPp8GSKl3NeUqx4EuLW
8gaVM9k20ldT9vQc3srD4vNhakqI3NlmIqSVzxGnpLpt+gTvYQraIhcDFGMGzI9u
c/v5q5OHd3rF9PnWxS5p8gJvb9ZnXhCWXWN/poDVJcGezGrfW9JM255nPfmBdOHf
U+sF3kJ50k1rXqytq5SSR74fEjeROFwWeUU7xorCjEiJsfUFVerm9hn46p/HRb6A
xvBiUhhqKC5ExpIJgE/urEo0y8J0yAHENBobmXIZehY49fuDdYqMNcz971RGBR8u
1auaraqTtBUUIbnumIBWsWcotc9TEYEp1XQmtUBZFnKtnbm41Ns6bvHfBWVKtsew
Gkb9ujSSoYk+xsE499LXpj0BS+Yj0Ykj1J7WtZn4drIUfoYd73f5QuGSxf93SP8w
M1Bq/cjUbA5XZa0z2w1bUQR9/+KzSy/nbyIK9SCO6jeKsJH/EE1GIzZuX0ZB8/BT
UNt0DEriiZeXv4ctERJ4uT4ALmQfMgVS3idwCuFCaI71jxDuel1Iv5zCm0Q+uMqn
U8h1XT6uyr9lCkijl9tF4IDkFmSLHDCZMj9iUmlg04sRvzWK6cvC5BMJmnsheQDA
wpiSZD6GMO+JniWBzkzcfLDs/Xpn/nSxT4KAO+PFJPkYzmfWGb+ggrhHIl/hRv/G
gP9VoAtjngb4nBYZyHMf3a7d8hLRGHh3GvB9jCs7nHGci5GwXcZz1jqZ4zl2NOSf
JbebSbeYbNT2AVc9uH9JsGUCCSRuFwIV2bBYljc3sQavAvpo/9LAqmQjVoeYU9pw
/yKHFiHiD/WEhbultIPA0UDIs+InZpaIVJiKp5mAYyUMVoxTPMyJU4T6sy8rkqZW
HWZplQwBLscZiYzH5mKd2s2Nywgp34JK3HZ7nsoVY9Ps0zL0W9kQ90oRjw9wJ9hN
natsyr6mIwmVU2qIysS6KljGy8FTOhhotaDt4MKCfngw96yl5CmlFvWlqSZkKaft
elYInA5HZeBzg9jf7naj70/pgMG7ciuPIp4oM5BUskB3i5MGBJwLvOzer1pDMIYm
okF3dq49G4a3PqYYya9fRPwvFFfTtyO0I4AIvNLsHOKgQptoImKTLrc+UF73s4mL
0ZvCrSiGxIUCfHWLYHdaQEgNhalZnIBNGH4AYC5guQ9P/aon5pcDdL3uxgWtNNiN
+WARiCJ0LdsjtUaJCj46ECeVwVVJrcXbeo061SPYTmi5NTEJ0J4uzlm1klEx1FZe
hRoasrj0ykGaRlscuXS2oSSv/OA1Zaxh0AF/UnkmsLlrlSLFoLmgJFZP/M+wGXse
1JLq+/hCfXV7csifS+SWZuQc/8qJY+K7n4SSbhtr/SsP6hA/94y28vKSUF97nFfJ
UQGxh5gh4ANSJVVF5stLqOdUyxBW0XSLs1v3o8MzHKpJ8645yaC2PGI0fAYSPbQ5
Ol8UEmnJdWs++35YZo8gbA+LET09OVXyw3aBTq5uRBwMw1PxApEe0GjOFfL83t2G
DsFlMKyatOtJomwxaUiOcsU8H3bonP/vQ/m+H/JuJKK4c014gWCeVHdh4LZEXfq6
4DKFfFAVgd1p+sku7+wNmgUlGG03isXMmLw7Hyi7PZuhIklDVW7Gt/qRnm+N2yBY
W3HHCB6j38PHA3T+UgVFiAFRFbcC+tYn9URasD8vG8Ou8yeMrGTQqanofZgewEzf
FWmPjJjUa0SS2JGcI+njNEdw36YP0CeZZZqT4xSnvXp5uVTprCuvQhvpVZCjLS69
NH8HSgfVUtxaZRdjmyXryVazCE0n16JZ3De8dXRZBwbElo86TdJ/7vXtXol7iKMV
JMWNiP9w1CItN9zPUI/p4834iSlCJfqbQGEuKw2Ge7p5+Eix+HqMF1vaK3wdJRtE
ESJehmNDuvrTyrzQL0r0SXnXn/bc5htn5dZEarU4FCrKWg4rgTdi8wd/eHSayeln
wvCO/frgbisikk0NivQ7fAKPhTesgelhkocOzcYLCKGZRFBHwQUChLgwTYszmXul
uv4Mz2zqsSS7Vu5qPtjwsH0NZyDYbyZGoJQL+dC/Mfgypo3bCXHOaUepat8JfaAF
aIAuq+BkhshUBz0C7Xdes7EIxmLO+56BROHmsnkEacKw9ZHsRoyJx8q4JQuwSmhl
uXVclz/5150V+ifItzgV5RY5pTYRYl5i15P/naA1I+I2R3kChXU5ujEDr7+NFFk+
OOq8Xy5ZBGB15PY1rI7A50f1fbkKUevOQB+I67TerxdkB7XdCSzd03XBbZkChs83
PcjDw8KCrYlaU/iYoQqlctwVtEEkgB2m4VYB7h5InimMiCyoC9d7bHA+7Qbr2c7A
Woe13Kfsfod+TyqjO1UXfG83TynVh4sZbI07Zv2P5gN1RfX9rC3NsN48XWJ3f+JI
ulXNEd1jLqy0N6Hf+yZB3WqVExner6EFJfp4lQLXcwc5D/dvr3Qp+1y6uuTEA60z
5SUeAhb+MpDj1+aDPZgnGSmn5oAQ0vQdC5p3/U5RpfgNS6UcldoQBCqbDftCx7nd
q9fceMdiU+b/hVafkf9iWdcSuywQg/Ibg66g+dX6ApqElkzCVQNbkud4teaFqg7a
5pRb76gJpuqhwsqlK2z6n9D7DJgC7yFc6GGvCDxp1tkCjmSTJMVPTrPyFRvpz0Fn
GtWE/R1QmxneoZN79nHKGe8OftJMG08JEr1Zb12//m97c5uLwLFyGqNjk3H0H5NA
J0pWoh2qIeXdhFZWJ0fuZplGck2Rf8Ep/xnGhaBRoDJ0VnTfkd57I6At16GlCYKz
cs/qukAO1+EiF1k3Drq3UfKhFLAuXsPgyjVCZgFNzyDaPqsO1fjcmu7WcZPmJkgL
0s+pJbw7qil2/kJMSQXqUE1aQRuHgpZyLwIq0rtDBKZzGeSJ7pFUQO2qTnIY9Kej
vb/sRWdjsl16hiZ7vf6rq5/EriAQjE0h8w0vfeFgfnkYNtBFGGx42nevpoUkRgXF
MdZQqGUrkuBta8enoysSMcVr9QP3QAivUBkOcVU4TpYA5rahGbXKk51BAtIT/JaM
PJLixGoZgjy3y4tIo9DavEBF3RCTdd3psmaeSjAhBczDYVXNOBjuUIZPRbEWvvva
5y6H1EVdJbzA+yfpzqVAj3OJknJvQjvnj/Qzb+afGC99uUQeTpwYVdPJbGAGsrF6
dhlfBYLU6i7PtF65AP262J0p5GBvLqU32eML7P1WTx3BfQjYOiJL4fLC2INdfrZ8
iMuLuXt1KmZgp5FvqDE6kMeXEN1pTKT8sywI3miKwXjFfyOXMKobqH68wi1GkRIl
0JF4URzp0ZHH58jj4P6lcy4qObw0IKTcCMs7kehQbSnGvhCIPMd2NWKKd6Z7TA/K
04/kKoU7AWqg7WW0VHwUGqxF/EGCn3tVvDPF8mVD5ghDaZu2lV8aGjshqoDnsCNU
XsTs3QqqVSDAhlXHUdwJ99jz13yPE6rJ0fAsO/ZydRhsC7rKj9xOvbJ/ZHkmiPFJ
wmGgmtVYlfkNWh5K/Czr1Ny6vIcc75/uGO/KziZcK/N7p3EIRERqfmtfosdq5VHF
4TLZMh+jRU/VhUq2fHzGYO9ZoO+sGaRep8dBDt11LqxnfO0XMBzrjAzLpDd4FXpJ
Q+chzg5HkMztyP83bLNeZb56u+v01bqzjFdlB41np5SoUirkTEnG8k3kwLnzr/+3
V+dtP30y+ee47BHAadb4v+L5DL2TBVt1Z/m4ZP3L/GP6kDBcyGtTDf+Iyb6YmOts
EtXER0ZrZBCqoLmIxCOruHsKrxKXyTMdZ2VDDuRvVN2ryKNruYFDMRGhzcPMDvJ2
z5Lu/vQ8YboY3MbvQq3a2G+BRP+7ME9xwhIxzdFoIu5dXqvW9kvlTbFTxni2P5wt
HyVEg8pB+cr4YCFrCa/FPOegUz47TunlwrCJLoyBRavJ0AIS5zs6Z6cRdMuEr2Ih
++bHQKzSorKVlcVO+eqXqIwQvK8gvB8JgEewaUMqh31mN5dsH6FfyfaNYQrznQro
2QCX+XdcP9iMT/m/aVpb8v10vLbkWqmrea07Gr9OFHwhda3BQeLfUJLKfVTwzZZH
deDT2ucI57bepFAvUe/iD0PpxSJgf5AsjLMLG3GsGEbHi6ZfUxRwv1OVo8pFqEYD
eu5mYzwEHdAb9JgMXo+WV8Kg1vEAsxeF+kdcvhfcnFhMfCy4VRu1vNXHTlei+lH6
SBixLTag7cVGYCky72uwI+/abYAMeEKNNllwH7/0QgMrzK0syvrF84CJYOGxcywC
RiuGiB4iCeEqmwsE82wdmo/+j5QWNOEnLv1HiUgM9lryzm4K5wO5xI/WIZj521JR
ecvA4y7hB96Iizz2oVDiIwdEk6wlxlxNSDjWyScvzMkIsl10+h2puOquXaH0LRoF
xnW3FBo/X/8DkTkj2KjezPkCUWBd/WYWQbZUp2LtTP6iCFpTGU6t9EZucJNQun0V
gudC3cYhQTixUhHHeKqMJIPMHnHRpZh8rZL6BthWlk1Gjm50AxIklsqTzc43U5Dr
tYgJrVfKNIiok0FIkuTLYj9/j6jghuijQkcc92QSRtV5NS3yHNRR+akfWBbzoW4F
aBN+060RvUyRhrbvxVMsL7c3/K4XIC+Rdt9V1lpXnU5bkKDxNQqw6f0u+oyGqkf2
+nRCvcH/HOUq1ZpboHeIQHX+Vrwt2gbUofpC7avLyNNKtlQqZpbVzVxwZAL/N+9v
qHIzItlcEOsdKDxlyjW8RY9tHzNc7ZLhA7cixvmy8TDxxLe/qnju0sijbgAWke52
HnU22tFYZ+e2ZCVvQWWRs2iaEMBu6scfL/BHEDuU69EIORZQ5rNdCCfIiD9bapqd
DBTiWkhGD4HWrpBNhJpxODh0tg8/ULjTa0VKstCQuMigXfHY8Mf+iamWWwM0LB9B
4CP+rEptOvmqKLwiuEnnLeN+1gFI+zepjGvupWxxuI4aG+bH1QrJQuP41XuDSAqX
89EMQtAgD8PK+E8s+2cyoxig5ue2UfaMQG49VvpZY7PuoBhyaHnq9EcF4Yfj/J/4
C7hwhXXWJohJZYpfW2xAOCnBhd/R3qAyPdnl5fRaK5do90/od9dtrUe//zECps1N
WwemtifpAWRg0boUJaszZnePCNrFJAbar6bfbGUxs29474+ORegv52LOzK2Xwx5b
PHiWrZVI67H9u6kRGZevFeCslanB56hPLAKecB//tjYb+yBrr/T7z18gEni/NXg8
iU78/AqYLFQ3cDrtqzZtMcMygM4AeqbwC8PRd9PmAKeOQ1zkn3Hh1c3NrpTkPLGi
iuLONskypQE8Ck6P5vpliRpeareFzFb5X+gaD6zov4J7aSUzV/LTb/WYLakWcrFc
Gx1ruBBxy0jDs8BZsFAhnAOxQi8MrL+qf0xQRBuM3WU67Xwg5Fy9y2wH/gaMaG40
50+9DZIkjJNc0CoLwlfqNZJAjjw1lvZdljDvupxfsGpBDu8711K6njl4C9ekejhd
+hr2OK/1VeE7N1ONXKJWvu3so1Ef7cHRQipqO1Il+F+qOV1ZFPkYpSI30QpFT/jt
yUrpKoOKdVAYCRe7snZMXZoZPQEKTorpG8b1XNOwQKTITq28tlUQQ3ecVKq1OIzF
k1CpiO++KLQAOJKGL2fGD4Scw9T3PRve6dghFFNO+9k88H+/kJDWVLPA/9NFAuw4
yRCMqciZiJV5/Tg39kFY8K/K0eTMw/h0diflS+UHUJFiMSeO26m2dsn5HeGDPf0H
wOsHZRMc31Am6ENmO+qZrByPw+kDkNGOIen7bvx9DrJFClq07cs9cjiq5nbWAATV
RmWB9E1VVEmuaHeW+XrQv3HOudVn1NiPLgblxy6C6LROKt+vBprDXYByReWLGRhn
PT5/P/Osiu8EuViG6bnhDxbvKj8Fbs7i4ApChcF/Qw1drjeFj8d9k0KMJW7My1v3
/TPOvEDeXLvqA/fiZT2EwECNJpVXcszjS8PNQTjjoheGnoDC0QN09m9o0CGWhfkE
h8T+/CTvnTfq0DwrDJReVWc1hl2LxRLBIeoa+QWe1/8LOpBU85cr60ZOIHOPyWhk
rYm3hUjLvBWozlUBG+TbV4DNENI21aLa75NqCUFCDDDfzJja4OqZAQRvPEUfHDPi
UDUWSViqWl8+jv1L1BaOqg1MF/m+xXygDk1mHTU88kcNNKQ4J2TsP/r3j+9gSg32
HSCVFVWJXzZrVWvBE3ETr92EoM+rpaacbnMZuocQ1ukPKsdz7Pu0Y4QLoml1mqaX
JpkMn0V0RQ+awf/y4hdUhjirev7iP+cwNIBWg2KelNOwTHEt/G5PkltenI884ulQ
r/iZRcG3kajOdcXZCzsx4GlN0miCg6sW+jIrMXKokzHP7+7nQQiikeJjGAOA82bP
oQop44UPHPadWMyCQnLnwe9StjGuxehOub37kMpurOh+vd6zY39efQ0t8Bi126SB
Std8LdYmsQNweYpPcFUy9u1Ld6S9ACCzrHFbEI/lwFoc/RhwnUM4ZuKauKBGcobt
rhxxWY1Esb9TCT7alln4ZA+e+VvPxfAJhTHeSnv5GQoBJ1x1nuPKjeIMbr1k/pca
ZXqP2XJd9VNbVAotZC5f6r1IXh1XtITQ5X+epvQLF71X7dVXHm+B4yJfGYTs34w6
QDYbqhCe5myJVM/8W0B5CJRu/JUsZsyKvp/6+azBPt64r+VsEqFB+ygTzrCdS0Oj
l7lyNXg4ktxEANSumQi8/020MMzMihF8ZXadfS5ujkYvM56SkhN96lPWuJopB9MN
B5/kK9XPMKckstOx9EclowRH2M8x70bL8pnzIy6byOv2pfptV973vBbUhBIhnvAn
MO++lccZnbpETI/bVuWrsYUraF2YZPTVOWxPFYMvKIS5Vdb4ABanaLKTlEIBEGsq
EwkNxILfrDP/elpKzD9pxJ12yDOf3BLnOYbVa/CJdChPL6xKkafekGOPE1WkOsnz
fO74kdb6NxffNU1ZRf4/JxAIKTAma4iwIowLKpKI128TrcWVmVzyZTfFtDik6qv6
/adso2nWHc51XiAVoOl1WkP9o5M0a88sMiRjXPFYTbLUFIfkSN8qCvRP+OF2eCwF
6hMP7oko+iSK/7xf75GKSN3OABj1Mx+JWB1RrJin4NoHitGmHa8yzeCn8ZTy/lkU
ASQxGT4kVstz9/U6azSFjCV97HbbM1JljpXV8BLHJqNr6e09QJNrppSJmflIJ13q
TgnlGvJascLkOzNDhhLO24RWnP/i5ad+pl0S5YSW78s5aiL1SvChnTfIMkdpWWCy
Ktcg2I5dgSW5ooW6skRRmitTuSnkEgwUOKNaGfIQwiaQ68AOoooFm3V0W+XJOVFM
bkfSKPmvCDn+Sfe0AExA5c+S0JF1FYruXkFjvnaJO9tL/b//8F/NJ1bpkf4WWYHC
vfXxI3VtDfWDpiTw3fV2IWkhvDFBYwVvq6P26cup7aySS3KsxS/AFauhWRhYN4gq
foap6v12aUXCFEVWlUK4XWdsluzexrLuuXrdLaF8EQ4pOyiAe8pj7r+8s1yy+J9Q
cV88XLtlCQuO+ZFrhSiciff/23HT78UMwN5h01u2DcBKe8xOG9P7dMxOPGYUtEfK
9OPFEUbzhSfN6VDh3MJ2bKnzN9V65+IzPGZf5Ls0L1Sqk+YORvs00zRdnIWEgzl7
AeLuqQ0EQFRi6URoGnfZP5EraDS53AiZCmdLlhfulAiqRujtdDMqr7zNou9UXFCF
lomOZAQL+uxhr6/6zPvXQ4zITufo826vHh6uBWES4RyO695+qcwS3YZdG6EuYSIg
xUsT6q3zBqeSVVg7Xh9c8hnxCTd0fEmtYXsZ0HR0UowJ2mouKPzfAIvmk3ZXmmg+
FTdJFrm9eQFerilKGLotY5R11/kmXf3pZzkWZdZ3fWzoTFjF8vnX0vIU1/JWAu+z
l9Nfjt6gkLdxACWLActlYZkcW3syH55IfZ8nwZNIC+J3z6ng4n6L1mUr8FhRByS/
cbjoLphZZ+8jj/xKzY7SPlvzB+L+Z5qcekOKNow44As2ZlkjaIxYPwzsEC/FRYAR
lCvK9v6GTMaTlsDjMnLlsEVkCfq6nhcbLdCRvK6RJunK9LfwFbFCONU72szpQ7fD
uPPJ1rOd7PU1Unorl7m6LfL1YGV1AR8yAAGeheMbiW/5QniiKh5QKpZ3r3wQvkkW
N0zc8G5mhdze23bRf23x1vz7g4vb0cIMrDbuEYeCD/Ssvcx8WDeCBYKVDiverrEH
35Cdy8LcARHsvah5+LaDkIhyyZuQ1+C59GsjVdl5fk0o90IKvy6Qa7ZSoroqRkXP
Fqi4dFyE16IVlyjcJ54PeyE1dB1JZB1Eih/BjAjTd+bwkALL+ulzUEz9ymhEK92v
OEdQNCY6py1AzKwvifZG+VT+7wtKuhcfRjO37j93NHLVCZTEEFj+3CSDksDNgMaA
iIFIfpNdTWZhlzhWKznZrUMvrFSJVelrBc9aFl9P34P1OnpqODJLdjjN9AcIz/op
nfNh/fXZZGEpeJOxH8wtTDoZPcWi1qk48D7sr5sMreAhwzP+ul1M0v8KurRcXiXk
k50+hln8WtXs48mEgjgy/b7RK6DKnQsu76FDcZthLnl0rV76S32VeeDPM3ntqtQj
smp57/MFjT34p4QRdag+zLBGBLd/m4YMJua0PnGqJHnlp+oFmwyg//VRLZkbRRHb
E1jbOdRCO54o1svuHVOeeVMUSumDiryYlnO1T/IG4G2pBbizfmj/G25qIQQ+tQ6b
jSXI2zdxet12YQ/wFoPRpEJREuo7kqOLvX+yTQ/x6MweW8tRfzi9whpoME2dBVP4
J8DppY+qaQrYMHamyZhp/nf3YZ9qn/xlSDZXU577sRmo/uPyhboLXNwsP9srnG1+
boMI+kF/kS5/Qxb4Wl1sOO3GWHgpX/6jZB58RoFiWstKXQXFL61wg3S96f9i5aEf
f4XrX9wRm/SaKKRSAyfeCp7TYkC45LfK1L2DFWvmMXfJoUeebxlHHJZKTGJtjSP3
dCnigy8hJ9NkrD3Z02jlP+tAWeSCuQ828cGXrMgw6zeyg3eY5v4jxQteaxm5EoyT
EOyZTHOHteWOmo08eTflqwTjRXybZ2wjzzIDfUMAm7cABCgQl7sh2WCm6U1eX8Ou
AKVg6/vrYC0inSmih9Ch9hGQBL0XofZ+edZ8iiyS3/pW1xKVCUOjsPP92XMXKRRw
Ot+8H5ErgGg0zdOumMeOUwq4bUvkKxGKPH9MeL1iNuZ3JnlrKwehdhboHv1cHmxf
9v3F5zhewbhMWIqIqAEFABMZiKtjc1TwezItSsNdOMj0m1DlD1C/zoCiNet7gDMj
h20hyw+GzO87LIJPj+2ZtKL2Nm0ubmCpRbiONF7IQdEMkW6mQswJiKx313rA2l0n
Khdy175olQc4cUfkgAXXnSk2nzTKP+naWU8aEX3CpfhfEXWBIGc46j7gObMQUrpx
MSDzv4boLfky6/4MfjVHSop/JYglvXlTSwOEQ4H0L5JGNemzSE/hvIGh6nZbxNu6
f0CIKQV1/qjeeEQ/NKUiYybVOB+pFR9rxsggvtZWl204L5TBfVzu9eIh12ALadLH
RCzgqnlCNT00J5p/XVKWtm/Av5hmWMpDZFFhpJiYqRRZvSP+KIzNWqrrfA4H/XIH
pLq13zCsgllyGek0TnxUpcwEQm9ahXm3g5hrJJmenU1Zu7K24CGerHXanqUXevky
sxTSQu0s3MelMWBa/OV3BXobnpsS8UzhKW/X/eK76LV9cEPwFkN8kJ7srxer4OX8
gyXgtgW3FD4eG5QuR7XnmDD11O/rnIsa8VtBqIFwz84xzOON4s/Hi7paReEmH57k
++TsEvcvg9afneaFF4Q/2FPhm9K+B+WwbCpAkcJs96jOqK1gtSXBX81P6m60j+0p
CdWoMDNb7unjIHF4TR7xZaZazmTpuuRWdyUdMUPqezh2xy7aLviZp2V1/VkMlY/V
IYuBdG8xhubAOQyBTO1JKSCosQZ+8N3j++vVy3baUy5d4C5pmNCAIXg5ppLhCd9l
h7vo2ZXzyNFd1ii/HYpEUWG7QkRWKtBb6UEM6YN6uFK5OQ5ZMMAu/B0wysMKg4qh
6fELMReKxRj2isHSGFy2w5PqYeOD1g51Ju+rDUA3ahNN5xrFIq5NWlCIWfFtt7ce
e8A/kRf/P++q6mNN8F9DbtFyR217K9tZsLziLwnRSn7QdcZJjJMNfechv7Dk3Pte
iMyee0R9+xEZVlUOy+OB9p9mjZwtWeHS0Sf6Jwq2rQzvpJx2t/27YM/2DKmV6y1z
WvC8klNecGtTlCo9vfNIy2sFpVYbeG+lxFa0102gvGlAude5M4WY4rWlTxYIfJRq
fhTSIR+4mK3VbK81uT8l9XM3YeepN3LDJTAl4iJLdNzhinB2P7aG2iCLU2+EanH0
A9Nn2qlFKpH0sXl/puQDwjrtioXdloL5wwNUtvk+f2F3WRS+HuqJuF/aknb3/dVb
u/6VSmxuJFvI8RB6tFi7athD4o72NkgFMsJs6mz5MRYNldRYKSGwhZav2/XJUlui
/F+zp0Wz4o3BNzhpx7D8QryBAcNMjHpqfUz+dadG8UV6PfnkNRRCTPwOTlVRtzbi
/Ettepub8Oz7nvfdM3OO8dVLCJWaPtwo8E1wXk9tpcItY8FJFf/LLjMfy3mzRqJG
khn9X1oHrE1w+7NH9BLvS0Pt4Z80lC/0+4ffDhaX8Q3Vr4CJefvBYFQFVFLCepS+
F8k5qnEvm0hlCXHxZrtp9FGYiOuB5i/zfSWHRttuRhFov86CrEhNCY2Xa9+DSmE7
T8wbaLLKy9tO0TTZGZOVDcTqmI5RetKJySx5NnWy8Qy6NOs9xerIj5e+QJcyfGu+
I0+3bfKVTBPL/iNjeEz0kDbGQhhlARWUDsU7TOBP/L92buHiCReSm4RF5LlkkbAj
ZLCMzue4aN+TIwxCO1BRmh3spcuIVaC6sCE85vw9fkpoQI/2D2B1kzbwhbgGWTJY
KEkbcSuB7ySDq4qE5NdHSqg7zsx6Ui6vRfsP8/ScUhLLRUwrqYhhS8yIo3PAq4gl
xijbW+usuNtwn+Pe/HDskIehmXDa1J301i1rPTWPG3iNm01mQ5eqqmk1zcYYGEbi
eIfnBzlHe157X6XVBg6g/nU1PQDf4dMuLnhc9q8N3KudsfmWPOxg6fGYpZ6bIKaV
YfWIVxkziwH3PIPZMqs7Arma96F2gsg759yo4v3qdZOmN+XJ8dHlpJirVGALI2az
GSFWMvS43Bts1UKmFb8zEj37ImUl1qNc0eK0G13G3WpjWDbo7NwWyk054KX8yy3H
adzyjNiqc+dcTXKDuBLY0Ie8IXzBo521dGKW9uSdp+s1HOfa/QZ0ApHjijyZmtjJ
JGejUERxZtiUxliJBgpFr8fkb+72Nk24gJRBC+U3Bzr0xMOwbVxVl5m8c48Bslkc
bvJoJx/gmFzj31UbHZYkE217cY4VVE2RiJhO7gSiUpGPp5QdqkaUiXlXR8mWaHgp
owS7jMrakAecVaPgSQOIUY9P8K40TSEUfzsggCpX0loS9yZMpjAi1Z9clq+nls0l
+KcB1/mogQ1XbVDiYcUAEBUMLDCldBl5IkAGFZeWfO42AuKhdCXYsyAu7eDRmumx
JAE/iLjiKz5pSJOxuDndOR1KyS5lFCRz366tW8zrqTwr3ZNsAnMk49tXaaAOqaUR
O+ZaG+6Smgi7gsvnWBSdD7k1fEq89kJOOquVtJg9lNCH12pL33mNutmFOZnH6Rk8
wsfrx/hDHVBcfw3zZkwxU7k8J0vcYSLfLZoC8uJQu8rEMAOeXxgO7NAnH5AHH84G
q1X8SRS090dNZ7fzRi+EMUNUWtxDWnLxYXg5vZ8eh13phfX11KJyKSPLkDblm3vI
K8BhtLJVwzjTcxOJoKTnQ7RJlXsKBdZepo2gqk91NJwDk4tC4mLDWSODTmrhSfz+
FuQGEpuazVwhwQZkNbwjfFhqCAxJRLq0Lfxn9uaH4BYyLWCK2FDdGAhFG//QxGMH
vIXW3AgR9lCVL9og6HWg3DN2miQ0id5BYZ0dsFhqc6UsKZDLKDmqCoWgmrlLW06D
vrNSEgs45A72JnBiFV85fp2dsznV41A7186II3GhaNV3/BrioBCUIus8x0mO3EVS
aZpME7u/4w7+QLcyRFzN1zdf3Wb3YZ1RBO5QXU30UDe0MhQlBZ5mPRxz3uSE9fFG
U7glrMvFVcPMl+rFu5NScW5SuDeITpOakBNMUnM2sfugvEC/Nw+uQlADISNuAbVd
VNpdm7StiKU9WUbLUY5pPH8oLOziZHOwM7Hl9KtCfMVzt3AAaUc15s9CxozK2u7b
OavyeX0mLySA2f+frNIhgkn7eHHWBOQsGBVMCNlAJyqtt7u5abdwfshknHB1BQj3
vc5jD+FUSKz8UAnNWKcKg84V4wgnThBwK3nA3QzD6Xnu+BfQDJXArtHtTEm7w1Om
fXcFGnPh8f3BFhq11nqCfyuvpPXx3IylBpgnox9Eiiw/ekKVEkInHzLP/Ed8z31Y
QbXNgqikJHlmWQaHs41IGxO23JdY+IfT15fKxdxSXTT3T4TlslUnh/yAtgPigEPD
BAil/ATLHof++0s0HVnkF6Mla7EX0W/BWRWayKmCFvBbz6j9YDcXd7vkNlxhbzjt
0u03G8OaMIY+SZumwHWsVHs9rHyWK9IlO5pv9sxwM/ibO4mHUn8TVkrHY6xpFY3m
w9NhtkQCxywNKooYTZI+hjrzoeeTOedQ2a2pjS7fTTYygYlH0gGjTOyEHMAkyj4E
ZSce0099/Lls1uCu3NrMb17UgJC/hTDadY3o6hfPh3Im5bpf8aBfIiE3QTYKM/ji
WaHmjaEUIe4Awy8yd5mLoRzVDp4P22R/a81vjogUmA1nXSUehwSniCHGvdbx6VGK
cF64r5uC+RGCoBGZeYiblj4i0o06Bd0GA9qAi34/FO66/W6dtThT1jx8CtLdx5S+
cOyFaHBsKGP4lFN1rDiFQm0lVIX056SOotpGe/U+G20aVF+MZWRnXPlMqX8+3BEf
x0qUiJIUREKNdAtAmHwwi9PY+NatcARXW3L85I9rOnELuwb6cI9By5qIyKoTwLDq
33RqgXJpVXCZD4dtxJmdaItm0B2OxwBoh9GGgowvPNac/8+I2mIdU4SuJbDtSVB1
D4+o4cgzLECAfoULgk/0WZeiZXQRcLcZjz5GS4vy/ivM3OpRMtniakVp5+4pSgu2
sPcubbUln/EryXLwA77Id44FlzMyI4mRwnNrxVqe/nF3/XPvvOj+awkCDac67Pjp
wFp+HGVIgNv2eN86zq2mJL9/9/BZG5lX9QHyG9sHur53yqfNRsu9Q9WAJTCxkAHX
I+2IwcGbnfzwYTu4rePY0IJLppI0ql4vXhQwF0GmuRIw52SFPkXoITc0U9jj+9++
GcDWCdr9uOxSl3kPR+KmBYNM3LsbfnA2SaM6jAw+OduR0StkVS8xcJ4OZL6fcU5n
51dhdJjmurn9q5qFN6L1f+AkwHAXYviWW4BJZ9YhLFQd/wodKg54fJ6YSuw8NEUf
S9aeUysT4FTHQe3KVsr196Vlziv7dwaRdXRsL8/p+8Ne2qNe433dvmiTlTuUOCG1
IBUYvWJqKz+yAi0jqtvfQ52H3i1eHATDVZ73MaR8sAYLGh/zdrBw78scZWoF8cAL
j7wi47SqSICGYjQRd12UY0XEowrrpdVLiaJlDiJ/42YYy8yIT44aRVzIF2sUHplv
+wYDbptHsmx8XenXzCyuiYr7yr0HsjlbVwhMjefQNuVY2YOp5njugzV5LxHE/KE7
CWtLoYTJwOpyojG34vR+nNFny+HVq+fjdegW3jSsrgxkLNAys3ELrDx5oXB3ajGf
s1pwlt8gI6M6Rzyrivs4uF0NZwDy4acPfl9MJ3dkz7e6SKkGZ2DW56fxCgLoa4FS
HmuTHDnCh2U433kCcmGumFd8EctaykZJEvep0h8QckaJUn1+7dke4Fs4BzW6IlTS
kSQAo3z9zSG+CPoveZPsDOy18VomRlwcIBuuQZpTV9x3Z60aWXqaCkAcJ0PK8kVv
VTXZ5SdgsP8vRlVjlOA/idhyiwfKdUsMsz+bOAmMFMiZ5Zo4LGBaFup6yM6kbS26
CLDnIymcvpw+3AyBfHlUIHR8eqWdJCF/BV2nHWhIx7V03Kr9yL3Sp+OGH4So5vwd
oQwq7ec5nGaFo8VdFhHrXGMNyW582TJMOYn2P/k7Wyn7lX/iLD9VgLTSQBoj0hel
PYZtPs8JH4TEyVafDJ6fvbdV+LzIQpddV2iUNP8IsvGX5OLSC74QwnQmBEncllWj
FKgGbn4MYEjpoqkJQ2Q2youeX9jV0Kv31Dj0a/rISVWinCXnjkMCfrxyGsmBItFT
6+MWckT7TWfHR6aPWn5IBW9BdnGxH4eEexJOMGdnrTHQYVM1+r1hdNSu7vlIKnqR
2QUWf7Hs7TDkCEkYfbZyTEv6HvSgYb6fWqqfJYQaa2+lvHHJ6sKBBw2NF+EhEwnX
XtL+wGx8UuXv9lYhea722qXB/HNvrTvMmtzwcUBCsB31o3wfWg3TJ/Ef4auxInUh
EyprCOPMHqOCaOP1Vr7cm5rB+MS6qy/eZNa8fKeyZ7/Nye1S0kpNr5IYIn+s6fBY
YfkfQdeXuegQKRx8ZmttFgh+iL3m0YDohe8NuBuup+nLN9t+67rwqbnifdca+EBJ
/kCMYVLqf+9ewsoB2NhbcPoySboEzOReVqthCwSJETm82v+PUWywBx9moQQT3PjB
/+Ntfj2PszpSmeuaujLNvhF5WbkhcwKT9t/gJV7a0Sa5A21LXswcHciDRAz1dcKG
RGD4GerimC4fZRvodkdq1r7ZujUbrieabM+nUciuAt5uSMLZY0beEF3kFWQuqr9v
lDUj95VYd6nh899Ns72KaymPbPns95V8eCDYkcvX84nYJTodcki4UtecG7CTJBdW
joI6IFIhjRCWgqy+7P6j+astkSWoAmF5TXymKvopNgUK0IUiovKZsltVCtfkyjd5
jQITLnV1w+1Kg0DHoHXR/89qEfjOb0iikTNMxaGE/rNf72xrma3szqNkiG6iuv4q
2GFOe/kAXc6Tn0B40vSFvLJa/KCPqAgeP6XVbHBwGcblJj5pY+yXKCoLr7HOChR4
DZ8exR8100jLEwLFG8335YejtXde8qteTwQmSZtRIYhasd/nqrLGNa71MCCyPtmu
HfSbJcZNCcGYuwXJWqWW+WfJd03DRfkISTKEYKLSvAD04Pu8T46M94jvMQ9tVHyP
69cokzu7JaHxcSVsKkb6LXH/Ws5JqV0C7GHmB5vmk0Xmd2uhsrN1Uh821XYFr5zf
TyKXO1azjOUz9E0OO1t3BBe35pCGeoWd+gHTkii25zTAw3LfBVg/1H8HZjmC2OOe
PS5AKvUK7qN86HzwYNiE90lam6qU7SGhayhPvRRr7QeOFxuBlOeE+iOFu4xKhMqJ
+DGsI0w8DNN4bviLX/fbua+uEpV5o2BnOpz7ZuLX+PYzeGMZy/hKkbCrKdQrQ0GI
NViTNZu3KZsmWn5OhCHzUUN1/PIzh4qxk6pDWKfHlrDKwzkZfmUszXup1NnJqsP5
8tZJb5Hr013YdMJbqZELRpkGpIEwTYoHN7G+JfEDFltcHbouhhwzHETEq4WztrCJ
BfaUDQ/ZM7cmyXGKZoHFnvsC3rqdH4Rq+OYoUrxmv2SYS3f/ZcClNBUD2PQYWEhc
MK0CXSeN2tE13g1Y5ReAYDBZFnOpbOPYy7zqTil0P9hJRt1msox+aPft/i+Fldop
CvqzBXEedCWqk0ahhjOh6cu14508NlLoVH71TcJQEG15AaCNWueLjH/KcWtVUmmK
LNNuP73IKqLl7awLOjZVGRsOI+HdoRbYa0XMVCSYaOZ8iBJXRZmTWJvV6u5MgdI2
XTw1j5noehOgBjXoWiMl3lRXJsUUIwgb9OBJ9GB8ysmnlErMn+zEwYa5bDTGzEJu
H3y0yOkr3EcChDpI17E/cIydz4D1FzT4G5i6eLweqY69b0wrImwFeS0b10VSzFiN
Qa51AVHJS66bBfGynvfVDpJhLa/Kcq8xD1diRjyfTTU7T0EPPTLOQlXVmBoDq2AG
lnVsqm64WyuKydSaUhNDoQqfUzqeRvXaWdnB+Hgywsf4fcgRTo834RYyWav3zJI9
H8lYoVFwaQyHWOlJ0DCSDCLabzyB4Rlna4cJeodVV2sr6gXlkICAZKXyZX/Z0oF8
2dUo+7VY2j8hOjyBycI07n0fIfiyerymSa4TBhbCgP1DPItboQnUVR7hi6hPol3T
7tYpqKcz/DxZlH3bZGB9Ogg3lgoex4gcjNg9qZS7jvbfJymoPG7DPGn5tq0roky9
37/Hv8IKOHXA/doUCjh6UwrY3T+VlYS6GkaU1841tMtBz22T0qn2m6RyVP9hKxeL
BWMNqgmHHfaH9mzYfHsiYwHrsK/seGhe5ziTIccjLnyukTJ7ikQwH2xt0cx9Mq/H
Z1iz7YYplb8ALvgAWiO4m7/1mttWBsMmYDjDWqdNuskVxuX3UBj/2PIC99ua6nME
FXcDxn+sbfd6n8WbXZdW/YPrxv4oFABn4sqPBQ1hwy+EppMCzoF/Fq4PM9+BtaaO
FAG0UZ8Bw6hIeq485vo/OTJhOxN+ZMEN2DZEeBc9bVtPhn1qrITRtClaTc30PVek
0vbw3bWkC2D0onLjMzPYDJXF9arWy0VEnM51OJtFGKolUWhkVPGgl0MqvJFMcbqf
LfOtcTCpYWTa90PZn45rvR9scIDMQlGyIVX0wrSPKHAThgkbgCAy2BLfPSkVfPlj
+0OzYn3tEU1XhZl3YTljSkeYF7fK4ZlX2dWMefgPF1N/RNvNm7sUzdXIzMNwXesz
488aTKADUL/1LCy2g/yh3vhf1E7ceViMKH9fejK+dJfxy61XuibD4WP1zFmC7228
Vi1vijnAyUJy8j6GQZPIFhpkFD6pFj/RjRwk8b1IGgP4cbwW4sy4EM+g5wdCPeyh
W1o10cUa2j4Xn+a3XNDl5B33DJLW1x+23ysMpiEPv8h6HYxPGMaBQELmyDnRNrzm
HgSO3U/XN1kYVprzjgPlZJTdOtPpzXEbyqjr7uuR7Vlb/o9gaux2rSqRqk5tz8uU
EAYGYUzB3kLjnxJ/Cs2Czb19VTdeLLVosc6UsCLSVCvhOsz/kpwWuW8D7sbXio8d
NbDnU5607bp60KaYOLrZWok5F+1ZTcq77256cauHcRnDsxTt6lB4pUn1TY4ExfuC
X1ru3BgfYr42YSt0bi0Yk3QjinugtQqifa9kdpzbA0dQAsXiEZjpSZb9/GEkVPqf
Vo/Axnow/poKuwIB4JVzE5i7DF7eYabviVuRE5rS4zBWvxw9ITnzQKyoXBjIkW8J
/XqNc9AjlhqwBQHV+pn8yCxpmScvcQSNp+LSWyico0XPXxuKdHa3/EwE5MUmxfDF
UEBrwmn0Y2Wo6D26lOLZPA1ijL8k7SeQmgJ2ZrTYUQCPu/MY/+V+4oCJzT7+kM1B
YQRP2V4G65cYsLDSB9/bd5+WfBPmz+NtQGNqSzWVEfq8MowVb68W3AFbb1RplHKz
s8q0FQVSfTLutXipkoWBxdChWdI45hf4Vu9Kl5LRUdhSDPoEerak78YgPlxAyyLW
S/cv7ex0+nL3pubfYgOJ7lxnlXkejXc7VjTFMNru03nLZ1Gz74eDXQWIBIsKE+df
7vPwpPjpKCfezQJB40QONa2I75wWOY4rk7jojsK5EVbdXWZSnPgW/VFGks3sVjWk
ZlO8wXHGKyBA6925dGR02O9/AIlzJQaxWAeokrHlnmZY9HxGv7zPhzlKjSSkhAPh
BDGnU4krw+bTUh20bK2R/ZkR1SxiAkazPDKrJ6auGfaskH2fwyo3oK/ipxkVm9Ii
yPm4wAYKSD9DStKhMbJ+TEPNgAzaWMEuqIJe2fmDHdLI799ANMDJX/JuG061+Xa/
tf3I336ssocyzcetpr3Fs/IwNoA113rwxLQcXeRoYuzF1FVgioGSJ4cBAE10AdJw
lBkZB719SCp1w9AKP3s163an2MnpNWJXML8JJ72v3z36VCsUb4xTVcTeWUTeAuSx
nOXxATcjcvbOQ+/bYbAOEsIYYK176Ncyd9QYUyi1Leh3taw5UlAyn5UNNPBa8nRn
Sf2fe7m0bTGjw2gQspPCz4+iDYUm3qaDdrxlzx/z96ZsOxbUo7eWt2YDF+YcRmId
o+aO2OLiIn4QNJUfnQv+D1ublz3wDm/QcnNE4Oc+KI7cLbahHtP2vT8u1SALn4u4
0XGfdtD2/vIqrFVhfAjxtJeiRJpmAnQOew+PH5nIRUuTyQyttrpiFxBLkH34N2hH
sPvbxrMiKFGJ0gPJjrIqP57OYymOcFB74q/EC5Fhu3igN/DfqM7XV3VijkRy+cq9
pGw5x3gFhUUm86MkBKbKYJq5r9RgiqjR1UJUB7KSnqGBbLUwqfLZzPhzI2rKI1As
tVkdPMXnusJMLkwoZeMRE4ZPi5L12g8YQ89iURDAJZRR1ZZCJop7VZoXphaStT1O
46ODwIfRW/ZX0lB5l30sQP6XE43AXaTh2AbhFFsuGEjKqN7H170JRGAD4uw+yNIi
HOG2sm+VRmVeyxpeONsYQ2XKmOU9dqknVGDfu8hL+HeBqah+IaMo1II+CEnk76wF
OpG+eW3thCEvLuTMd3JUqOJaUfw36YjUxihPCrZquiZl6JzeSzsTKA9nCLwdZTjr
Oq8bW8nRTJIKRR9nAQs4Oud2AofwLb500oXlh+t413XRgefDsAbsEcl3tm7xiKks
IT9AaxE7Oh1FiYue7E4kExOC0JaqsYHwIu8syx2vBWkvyVw6IYeXYhEQ6RX2iIA1
84nZme+s8zdtLG9FjKzt7iDk6+HrRd0QM4s7g5JyPTRDj8WtsupsX5oZ9T+xbdja
ZD24FZYQJgUtUj6bD3Zs7p5UP0UVAksOUnUKatYg0myeht8Za3Cm5wh6A5bDfmax
fRbfr0o5zPT4A2QLKyeB0g2WXEOlAZo1aygR8A6KZhZhyVpbHD4HMv1X2+druL9H
c0IjLFMcyb17vxiGl9Jshgjx8MBTcr2YEbPIhjrOq/6g+QF74TQDM1CoDzrj4JGx
FDqfi++IMugBS4RsZyqEr7DSwQudHh16iRBUzsSIzCdhYlLL16+5LbrxX5+3m05m
pxOGgCxuasd7TdPTGbns1p/qcIk2hmojLWhVa8/zQphnF+zAEUlrQl1cXeCd9SqW
pS6OKE/wadre2W16zJDhr+s/SS8t4AcysM+2AY1tq4ANetkuJneBZ0H/ogFzCXy0
z6JoAjhY9dJP/Tm5ezPTMygfjYf6e1Nx1BJQRINHYLh8j+ZDtNPp/pqag0TTzsLL
bj2dp1gHUmj4jFgLSEOGE5f67MTWaY/CkOQTRu0k4zvYbokXQlkTA8X6rRHrjdab
5azcvR1dTLztz4xtjjkbnKygv2mBMWi6ak3JXJYyrzWEJqtWSLZFJe9IU1Uxu5yM
ze+2jsGpQPUL6YOWOXWv53LzCAatcCqT25Z+4fQWw6ufGeyIMvR+IsYKWKbCcwm8
cev5zSKhioCCmSQ/piI1EXbzKZ2uEyek1tdLFue2HXblddjCLUd6PwFX5Wwx81c4
NpTjxy/5MW3EWlQigNOcvB+3Z4+G5Npx/rSQ7cvgigk5XPxQeiHjccr+ExWOOURR
I5oCJZjaO4ZMepKBE+s/Gy4LDk5wXDgw7CTjnjlZxopB5YJnyMk75LGKa7KiUSRF
/AyIoYbYQ2ucKBxWMLBxaBtHHTa5N+ISCpDf8bVFsxZDKs+tZNNbfySQZRNSuSvq
NneB8HD50DAO7ERpIjOvmexMYReBQR8Poqk1kzhICG24uosggHcpFfbjWxzuy1VS
0ljCLYnT0rOeQxTVz3mHoefd6/Qgqk0BWbx3FBjphFHv+ZpcuTUwggqV4KlNnMGm
c6b+V+JUCMLZ/1X+8GukPBbxx4JsLZGEf3agV7ObQvXnjSuSIzzvAXX1lKj0b5VR
LWe6sAsYpYlHSyaTHu7YKF7Z8fL9rDqxf3q9TYZh60G9xjJkq1DG0PyG5rWUPKP3
uI/yM0/OFqaGv3QhIp5XkNQlaDoLRxmieUYK3GvYcGPJAJZ9gxwiitCGQi5GHBbc
kocrO9X0c4AfmVN5uxD5zpEwfEswpqPCgC2o4jBtVwPZTXyz1FT3/8HqEd7JtTNT
dtpMME2CkLRmIqUYvZYsgqti5qMZvcvY2uIfqL6CAwo8DEJr1j0ZW3aN/6HUJRaB
6sBD2eSAXJxYi/NFnEzQ3oIB3XKbMvRZ8hw36XrTfEzKo+mkOSjTbwLlEuv5ITLA
g4wp+3dCAosP8+sIZP5UIvnhz7k/G69ri5teEjcycJRn/advmiUhEqbeSjSoIZJ7
cW/A0iPNHtBxniVDiYGlEKO0K2qB47hbxAsxze0FL1CKJaOK01BJM5A2caY0V5aR
bijqu32R3uSyk0t/6jNHoeap4egELF4Avc1jazk+BiBNR/fyvBKzxFHaN8enCjoH
v8+b8G9Pw+PS+sieG7EOtEAi2HH37peG3uEHxy/chBFuyTQX5U0TMdHDXyqGEU5Q
ho8l3nTk8TKm0j8d8IcGQrbiqTo0rlvXgrGqMm5En8shbR7mIGHfJoKV6EQy14SY
7LsbgJM8oQ0nVK54YtCg7gdVGH2V+/HnDOKgRnEkfyWemIuAgwqruXOY6zgjc9pO
ravuzPChR463EB8l6eaZ4W58MIETckSSetHhDzNkUmmqB93RjsId0I9rURp8ZOse
GgaPvQqnG8/Zqkpu+/BhExKdR0TSSZFmxL7seVKu8c0pQIZrHOiKutKpZAOJWK+O
llgTNZIHfzzxuud863EmhXORSA+p8dt9qBfx+oKzkKUEVaWTnGuiPocc7AVvWb6r
GhgRHhZUWFGQjLJwWBaoVZ1+REzwy9AGW328Bu8pdLzAMuGTHSqaH4KpUVoPNl++
Lt3WGU15csTHt8MyudVkzGOQPyeH2Vvf4hswqhL+fCbnFwSjCOBTK8eHJYGIcMY7
R7oj1adrs0VQtq53CSp8y3GSCOgdElw+pDezhQKDLW1shgeChFsYGtDuYgYD4oKs
YYdya6+yDbKO8W9DivIKPPDhClQ//5BhL4adaIJcdmfUwsjfXRgWCqVWoHxfhQ1Y
E1fP+BtcjcJ8WMKlnzx1AbC4Mg77fMLkX7SxQleQHSpihzyXgfB8wlJZtYy23qIE
MN50DC0yV/xQb39p8rk28Et5r67Y5X7LjUb68tOJnQHxThNrIKdyvbOyQibyYkoB
Xm0YY0uzk/5hKTaRNBjM0F/n+5CADZmNUNf+xaEqEGpCnJ5v3B6aFhbVTsTHJqff
Fehv4risevqMN6tyhyibSuHBAKE3igiCxqB2BhCS1r+NhClQsqwnBhe0Un9oTAvF
tlxodTNSWo9Gfqak02ySzZ5EO7E4oaLgtaVD4ZMKSeIQIqDfj0Dxm1vXA9g/K9M5
QuI7WW/vPUOZLftanFN5Pf2mkBsjpLY8XnSN2hs6FEK5TViGg0pqdZwPWPCKjFQM
+FqVoN6Vxwvb5psYPiD1e0Swr80E+A5ZsnD5Ydg3dy3gnypnqpFzLGAOSXUgHm9w
tuu4Ukv4w7O58Vo4xpPUeo8dgjFFwWaTwVG+RLkGUNbn/ODJjjiV+Bndfmo/01Kf
kvz+2LwdDXD+gq4pKt9HiW/0Mlg7JRCgGN2W2sgEvM2TLnJXvvksyXgNZJ0Le99l
oaC5tpuHiV6oDatxQA3Glek0XwXt18cBQbp3JfgGdDUPUgSvRqHuLFKAdYJrwd0F
cwAchlSnWeGhLBTzxQZ3RqkKG7w9WbJlnkx6cn7Fm4juU95fbzccQE95d9sOzxXu
2SpUjcboGa9f0N486err/F34lvJL9Ubb/bGXvzzzX2KuzM6Q215adYJtB+AsWJnY
+AQvmBELEkCs2hYrCevIs9fxG08CXw0sBoXeD0Nl5JXT1jINEPMO3B7B1zAVUeLi
fj3V88XMMJQw8FH/k5c0wegs6XSUGnApGoZfmXk9yPfqkP76d7BlHEFB1IqfUami
SSUPUJxYmgHCnlOVjqZRatOm6TafPM7ezQaDi4A1swBUf28j8DO1eFdjt8IQRxT2
3XVi2kfvjcV/JyO1HmyZybdr7N2zjzzvFi3+2Y+eKagmUxnxXglpg3CU16sGJUkR
LU0pb0iouM/mRmjepXc3QIuHIfO9h+vegR9HlQs9Bh18zHL2V6riXSEs52CVMXQM
05C211CEdDt3ov+Ruo0q9Eo3gUVCu3Y0cC8WESgJ/hbABIxqqBqwxYSEsfWWafYL
kfO7f1jmdr8I3XrblGdJzCNGRq7m+wlzE6sF3ZwnNLypD5TY4/bT577tdsilOVyo
hcnhwRsKhEsCHP+6U2Dtz22g3mWl9gttDzOXv454fDiGQ4Jg6EFzfL27jiEA5eXu
sh/vgVDRhPcxPdK0cV9OJvZqgBsfE62c3Ra73ch4n9fBY+PXd26O6vEpW/iQzVjD
PqOvU6a+irD9K3lwRlPMTXiWmRNEYKUZIUZReCIppNk3e/5h+slIoqf/FsF3KbzT
MlW3aRhXe0YuziultqQkGe1O21X8WFe+aOXPZRelDUzZhHq96Asg37fehQp0bYYP
ucXrCk/B+H/O8fGDNRVTrouXrufCbLnHnKVdC6d/NTSMUgs6vYEQw1ml9mOR2ubv
bOiFmi07sdUdugvrEddiaTmXkKBrGxjpDJTHHgvzlCZNpfy9Ha0zEHlWiDX8AY8D
QbFGZ5WB7zP88/NUrCY7HGd3EcXIfrU6XuSONyI1WJzZ52/kQuaevXWorjtnKkIW
/MSyzRH6FK45j++zPsrODRlh7RpIRaZLTZfB04rJjRkg1u7IEdyo+9P7v2ZgVWTF
MVraubZaFtpat7zCQfqMlPNwlt5VXtMg44EEYVe5sFouDhMUkeaHhs0fBTOVo3Op
Ti0s9rkbFcn3GjwhK+vaXQTAsuKCdObj1+lv+CvMEk2Vpr5nMQgdLZ+RzUTVi7Nf
6OgKBviZUcIqUFPXnoU43X0PSVHm7I21/3AjXbyRE0HiHIJuWqoSIfb9pMYQ549t
0LxFePCNaMr65dHh3gl3kEfVRu9sHhQmoLFPFTedNE5Nj+cL9hfOlqqofkuWd1jB
oO+bR66EiSQUqv6pK1DLKduDkelkK9ykepvzZU42HmrPGMnuvO4Z9DJg1HsEQmja
Jsp9mPPDNnds9AZnqppyyNLyfpw1Iw2pkNqXVwPfKQuXnMJjOykzMxDl40xbvYD4
uTrEN9FgMRfsBkMQKd4wu6UY2x2pq3tpYQomAcHZR+knisRK1oBUzlooueOZLW3n
HOVAhCguVVEY8+MMlG2bY4i6eSd4N8BngZibpmqsTkfbuLyTPuvPphrfXE9p1l82
PWeYPMkcUidVPtMYWfPFjz+cZfxvIbni+sgn7HaVaMyBqSDBheXix8gSOhTPfoOP
wXcHR5fwsizpqA05ggHIvzVFJb/YPbF7ztdIRjWmtURw+wXnqTcr4nCw4+5MXVpq
9taTrB4YcTlfd5s5UAWdxHKHpzYK1N4j0FuxekSng769IqVF/CN9G4dUpF9M3o45
rpIn/EcPJ5xafrsus+H7NuxNnaidgMaaGRC+19H1u9Fkv53r2phu3U83cca3QW58
DBnZdAC7c3b1SK2/5ljLzB6b9r9r6tQs4smR3Fs1pf9DkhOUBTRgoclzyZ6Fm4zB
UlfY3Z8/4wEjcgxjm0QvYR4yqkSOSIxg4fxmLmngNSi8Jj2NrRRMkmCUqo6C0EJU
QpY+qSG3CH9OvcFazybkln7ZZbdBpiRO3ZbYIHOPYhxOI+6D5RQRvWBVaQoY5UJm
ktnovh9yB5mkPLmnjLyb8GYz4DGE9TqwTbZTTIDqJZktirCzj4/WvcNzex+IWArM
FrriCOEb7JXL53UQCEOsdp+bYFGXDrHJ3R/yxBM6gHMw4yFeN7hLkq1tWi+D5gur
akxGBNvehHruxo5AXVEExRhXBx160GC7IuP20v6LxWZAKT2CGnwqV2Af45lRqwCu
pJ+Ryd1n1LuSR6/S5ZTgs1Cppy8sAxXjpbp9oJWep8KyeySX8SF2mFPaGXsTs8h6
J9AnP4U9Rv7aJ42Q9Tw+47CeYcXFx0D5w5TIdBaegkdLWGvA2HcKYLdgOXtHi2/P
6ztQvKT2Hpy06iyhHnhNF7GRy2X7Oxbs39sWBdIQN7t+9vcKDqqaO/FUOocalW0f
T5SNjA+yvDyz43vGspUc02UHlG9k0cju8Ggu3mxa1GOWdHiIJLjtLnGt8dJ8NGVw
vFv73PfYEm7uwyMPwi1dCTP1JR5KHHPgbz5mIU7gMLlStlGj+vPGGjWXsGzJ+8j0
xTSd83PWiR62nxbEzzoTZtsexsiy4TlVnY5R34jR31fj5FOCEOL2VW98AxElYkGh
8CrnUrQb4o1UzxaQMROjJFVvugk46SdlYMy7byxFarTcABCmaFAaa9sumBRykFDw
CON0QrbSy2LSMMEm65bJhcdRz/U231igYubXA6t+3AvFluN45SoMSMJBhyqEQeYT
9MLGOBiRLUIPe5rQLAGaTeWbEhHz6+eZsaavdE42TxGL7vcDu9k0Eniu6UhMs+xS
LuEzspfnxGhWJPpVpnvw/1QZ8RFL1xGe+LW4M0g5tvYQTqopVicQErEouw97YI8B
8Lq5m0+GyNDZQ1WSVM9WEGrVkblzc3UCzcLfOA3yuEXk6pct9gBTjXxkxluhHNo3
YVJ7Fymm29jeBct5V1IoKTrGJJ47AycZaw4WZrDCTFOtJ0MgHphdxbjGSKAg/eYf
ARih9SzvcfIS8zVHyX7OWQRP5Q542O8DNbuyTSvx/9MsxdObUuQaTkA8Aav5Tzyq
YmRk/ymE/gyFc1g4IhhQ3NrV2yXXEoO5/6T9bykMvOT85inXicZcPQ/DXSEdJg6f
2+D/6wuY+D7qAmjfvFHG1Rl9kXBSRPWqLRryUUKLcNnCMh+FAha/sE2xk1A0UJvH
UX78gHifOqAPDfkSmhei8D7C0i3ZnmXwVezPd4+B2Jp0KMG/vCpnm6OBU0NV5Fof
ZZJWoJx8Y3wf1ZJasjYq+X3PqySf9QE/Go4HeyaUgHLwKV2uhcc+KjlaLEyuk06R
DXy12JcqMe0E3XfCf0vJ087AZiTOk//lVb5LmWre6VymW/HBcUnn9uHIwjj1CIpQ
6K5a2vgeyfmtsJPZdDBmSJ3bSbg1487iedj4mBcgw1N8EHd5NXpX7eT1Ujz9W7Gq
XTg+NpQyTP3e8sSlOTVbKl/blZdry5AkslU74meQ7MrYyNk90PUuMvI0EBfcnh7I
sKbAivqWMcm2nxhbWHbcRldl6el17ZD5MDw8wtbP7mY502AVVoXByTX/8Nk5c+Xp
PNWL+/sceV6NyZQ7+3FnymisuTIMb4Pu/CvbdaWFBnYE0MNDyr94zT3GLnfQtVY/
pHW6TOo9l5DR8JRXcVZdOXdmktFdlqE935XGNFq31hla2aDIQKNQNk/Sti2x7aSB
BaBB4bH0g9m0qDZUlOAn3uUOPYHyHSPRJTYq2TRv3pP/tktVBOO7ZZ9AbS23EZdo
8yDa8VSp3INtOT/xEgif7wfwAK8tMk6C3AxIstpjg4+pVwKZb4YvVQfN77ie5Bxk
6NOETpeqr4YoWYKh6FhYtN4Hh+htkJGsXPbFmbNflXc5qA9odX7lf+wpKfR4QkvI
qghRqlhkIOJak1EhX2PQTmxT+mUxQXMC0gC+DLcLJ8T/dBOi8yBB7qI2exvBBmrW
M85nHdd9+mSo9i+FTfuiYN/esK3yf9rzGt2KFvYv9lRIAEKVpRmuG7hq5pciDis8
yqVU+K2+2fn4MifXKYj/2zV+aowowMOEN2+9vHXko7UR2urAZX4t5nKf+oHGqa3O
GIf2yrD0IcaDxbNTN/SzX8Iv1e2lln/8ozKuDQ9f3c7OsbplxB5LY1S9t24MvvBj
KcpR5pl4gfZqzUsk8AeMJC+ti8h/5C+3VufIBQrX1IuCQj5orLCvqjVICcBihPzh
vz1KFNDiIyKVfpNKzMBwjjDvOsjx6ISYWW21BjtZdzQdU8iafJ2JHQiBKJ65lCBu
V1gJRf5ugd6RVW3Um/aXiUwxlY3yue+O03YkUVRjUDMUNzmvttHGP+KXXvwA3+jh
WpS6Xos+jhyxHlHd1mF7DbhRM0F48yOGhhJup2WpGg2WhNdEfhWSktWdnYoZSjHN
Ciyy/eIrnd8tGl2N/o4Sg36nUlXRO1hHSMvC7ISmI6fddhud1lvaP8uJYOxd58lz
+y+ONoD9Cmw06R05/eMoF6cMLo/3JVLEgbJrOOHVTuB8BkSklODzcO1em9GAUbVK
9SnJrbxHxhmTM2m62p3p8JGlI9S9PbpBBuSic1ucbmTnSvfjTA34hrAfNo3P4EhB
pZXVwmg9/CTlUnnj+RDnSRwPcDIOfV/1VV2CI1aP8z9PtKCVNM+nQ0GLRPYd9yC5
SQ61C/bnvMZaOz/2uxD9EQvzs95FH8XPo8fuBn+3sCUnwdHOpe1d2J++rN0CQk5W
teOe9WUg+7n2x8SjXcbOPLlDdyiP5vdoG7iGM/HfgrO0pZtKTJfHN2rRlxbp6Njv
+zZgpdc8hPHmUNAMoE0S6RoM0Nxyx4fQG/jwcCmgmyyHJYwSEtYxGpNapfuh4aai
vIOX5MmvigDBx5bhX/VxPNqfkP2UZHCJWGY6MoxRKfqfK8iugZobL9fGAh2NYEq+
ngvKPcqKfgnj1B/3S9nFvrEvFQIJC5EkF1d3qoM248TN+PgqRlmVvBIZ2gBR4ApL
E8PIhg/kI3ald2ATlBhrVJ2WBR9CSP4GJBaUusE4++YreU8pjxszOC6VR5T/7yXv
hsTINNolbFK2FJBFOM8EzPDvjKzG0wyTFV4pQCla+Nl9rVb08X4gYFOu22tq3KdC
DL67lxV+SUVkK+ioRhsW3Gs0huiTbQo+1FhHOETCmYU3A/3whG0Mtsz6X4v1tpKM
3WxQIVsJWNQvTnBMM368RwqSxeZvdWZtjAqUH27KlraZJq/7sTOp1JTHIH77X45R
ZLGifL17iXTk7H7hbkJ1CqSiy0jQfHAn96RTI10OdeWJgBAft+JD2NoRXL2o9hZo
BQYvyk+LLTlO69uQ2zSPDhgkCIH4HGRv1T5FAS00MPu9lib0lH6Wxm0V+TVtcERI
23zQ52bSoCjiupdZoo8MkzjQCWlabZwaXX1EerdgIWMbIYkSKAlHRz/VBskrIyqD
pAo07yEySJ3C3oJum8Adt8d4tkLmYuC47bNfJrVDvUaJaOzalNBKltZZxiGrPifO
CtaE9Fl2T/U7v8g2CRuhCsBdYACHgP4lOa+5Hvb/m+oMcm9XI1oHiYg5FjoP3G20
PnhHRVLtJwh8krY8yQ9oiQReyfp3RhnA5ogsVCWuSHeEl41KZHCo2w/cDfBzK9h4
aK35LYA8Oc9UkVgeVHpMUAWAuEw7tX72XlEKhYdXOdLbOgE2RAWXPUOTzg6y7jMu
FgUWTXoN2YoZkOjFTBrphAIgmODVit3Z40sh7Z79mMW0oy9bTHQX30rkCX6xPi2L
I1GvmgPFfR1W5qyj84fbq+fS4Xo3cx5tIpEy8wbLrnohBDkM0ChRgDMokKe1+1ZP
q4ii5fEAVuVVj/d7FonPglLYSb7y9P7tCsAjlzyiw/kZ4pZx7jsQy+m9YTrgdBV7
UJ8oGY6cRaXxRPSzXYDIXHAzH0ZMXc60jkscD2I7WkuZO89usNgbQ4vkVztSXyEC
YJfRRrf+fjIPocd0jm6JHvF7bi16Thv0LtmUMnbOoRiCSGdGVSxD2v+6tG/9bSSz
KOzJt2VPfU4/5XNLkWe5RzqnzI3g7JoOe095x2QqFSF0lbCL0/cFi1cQXlaVLruX
TOSuv38FoM1POzMS1pe7YE1cw+kqi9AWzfC71OwDJ9144dJKt3ugtHIzWOfmmUTQ
h3fe2QPbMuMnagLofA5/RFuYVPr+ajXV5wPRLbXCdRZxUom5BCalUR6qIJu3aHiC
kEEvbp8O2Q+ZYDwzZhtpl7W690f7KQS3yFkKucdKwrQxPSoXvhAiljHubcj71IF1
g1QtcJrg9NaY2jPEbpyaZRzYp9Ccsz39BOPEFQ8RVSsQ0MAJXpkvFCfmCXKR3wOP
oqPzztjwbsz6OJXzrqBLyW8cyjUCSNJfwnI/PL+jM8ZHYhv0+ChJtHc/iGnmK35G
WqZc6lX3cJ5kDPHbIPYWFdC7HRcjch3TCa+DgNA03DZpUo3mYNO/v9ZiSaGosEQv
VQ+rJqYjiSB/Lp1bz7Oh4qhIcnt1t8rpI+gIrqPmdIePIf7hua3dn/7FyB+Ka4Kq
0MQeNPzEZ9DBXclZXwqF+sgMEy9x3zoSt5Q/4G3goHc+hwm9k35dGfz351Dr+7cz
9YxpG8x9tiqnEfvvJPHHxr4lPEFxS5YwJSSF3lsVrjxTIyDJzStyGgy/Ui+Ohz/9
mClwEcgd6TEKqjnVENMA1+YuCH8pt4TlVJ39PfYvtgO4D5jkzJD3dlkHsOuO3Pr5
gfbpEzTx9kZRoWrC+qhAY5rcsn8B71zbt1VEqrlWMv9Dp32sG4s+1kSbFhgnElBl
KiN4AtWkj+TKZW9446y2QB6Qj/arW0lccAkqS/Su6Mdt6lMEYRJ0ArnRlxZauTFO
UE+4XUKJz6nW9Y0rNNrKra3COq+RpgtiBM65ofg6nETAz+F/2FgfFj4pZUJNP/rG
qnMoF0CzlWR+gQYeHQsal+/ICEJG98PY3J5Budc4LzNgie1u3SDBMOCDXc1a/hgz
YkSF8VZoaOD13NRGfRfCqIMR5FFtMERtmZd2o6yUgZDBB1LIpvGQt/3cgHmXEilb
S7Co6dJQ6a+neVE7w6Ek50/Oje9DN5c5P3O4vEi9DsMFFnpZi2OmB28Pt5KK2x4w
JaIZcHLezk/h4PyLMEhDxmWaMK5uLwXnHjQ1Mrv5OKWlQFBiNfZklp90zcsHYVtj
7SFiq+lv82shAkxF70+6RNxncl0ALvSTfSQagWpOW2gBaa16WF3CgIPZ8nydcWBv
IYV21CsVNkougR0Yg89R2+ySc8lmXnebG1DK183oN5khSE6uFAN2Kgx4kzxK3ChK
5xnq28xZX4Xb+310Su45YBH+qxFFIMpWPtx4IiatjL5N95Qd7OqwQ62sUot7cbU6
KsVn+mxV4d7NnYykeutA/0mr2QxT5CT1a5R4cTWBwXjT9JHR6oLTbeuzeRCo8NVd
+LdABNLsIEkqyozKdmrMV4+5HDaIeKALK+3GPXTGkMEWvVwMc8F+r0bOuv4oYODb
OER13miyoid6mhvpoM18j254oaJACgCVpL9G0XETjUW/0gMcsrAEZT7ev8WCYEF+
edCe5uAHh3JmNjdpg/n4FzypNeSW4m5CkOJS6dUXQFt7i2SvN+oBP+ox04erzW91
oE7ufioGefWx8k7ZKF9iB6M0yOt3zFlopq8MKF2YWgffs1hB/nbv5JXn1HW2vz/j
lQF79s0Hf4iCTLaChK2xV7Mbv7QROfzpuRh7ZkUCdl/o3+me1R9wer1oZr3cjrOk
hRSX9Jc9yvdVDvGanpA/vftJke1EaY/vvJbyWLUPvyl4lHkebOMYipGlCJ5y8Zds
EXTg7let+Nd2b2uWuYIWeNsFKtGs9mXoanzVynewlKwZXAdPM6PQd+RxHPZbeG3D
udyptBfQorCmqbnFJx7BoVCM/vZG+OfWg95Ffbj33Eaiok5/WsL0i0QM5FSsKn5V
c/ftWhXA9vfvIJ50bJaUhNhQMQvdubW0qXpBdrL8RhumC1EqLLvYuTPtw/9qqHOB
LlGm6/9UhT6GCjmr+YaT/pEMj9LysQnAfMYdKWniMKXmzmXvlG60ZSBYmZ9uxXMk
b27tVEBbvVN/Rg1Gwxjj8MTr28S4ixWjUkwqvmLYSn2bWOKdLVuWCUscloUTRQEb
etyyBZu7aG+pkwkUJ2RWWGYKybmvj8T+jQlcl8Cbr170cpg8Frp/82QQfYvDY1KV
P0iid/b8TCOsXzmMfpOZioZH+7FN4MQ3VowqPVjZyG1Tj9Q9IaHWawhxFlMRQB0S
6yzl1IXvK9aPTrrslkw9jrodXhBXhkC+aJaXMzkIoFbht5vxWZmQtOPweEL4fB6t
JPLmSZIGL4YVITq0OLBWFzp9DW+Carkpu4x5wiRLooUhL+PG46Q8EStXxEBvaDkG
fAwZGWhTT3qRlvuxRNnSlU/AVId1+fUpktGLPVKvUt9Hr9GuUSxe5rEdNGPnnkjP
3upa5W9aOLFyTlm6Sglrbj9Xf4jvyBRUAk8MjQsaOi9PdzDvGew9ig/NGKjHyumS
8SCKpWp6B0E0c2KQCQcDqBg6dGwegxKT2EUh1o5bGBom3OBSGByTwlrdpZLjUtcT
eAvsxcxRTVaUB1uUjaUeV5KckbN501/R5CKZYs93ozuFChHJ3GWM/NmADHa01sNi
KbWQCQEsfsGWxu9QyISDnMR2Nf/upXlSHZCFFfi3PYT6/4a9JHVS0LhioseP3+T6
nUFtDPEq7DhG9VXpCKg8S3Lgde7HruhnNQYr22r5Qd1QeutRGOFYUsBD/k377oPz
d8nR3Fp9/YYAhbUT+yJGBokzjyMQ2pA9Pc4PgkDxQyWXpfMGxEDAnWe/Gfx9WvNF
fTYAan7TyZeQFJSS5OQ/kJbukVAqI/H2hD2NbX5r+qTs7/211FzY7Cncz/8+gGvD
Oid0K8FqviuJHju8CUIU8CeIFDOwT0L7U8MEuDbfcCGo8ETsmP5iYakW+MHt+ZVe
igpvn/UIJaFiLTaaXayt6IpuZj/b/Y/F9cNip5TFYXUIfIzsAiK//utsMPMHEIrr
2IEsNUgtsBSRruG2W2q7WdUTX7yWBkN7z1qbKOEbWIFrDSduPHGwUMlaEdTzD4jR
DmDpPQX6mj8H35D2aBdzafHqkJprk80tsplP+PswHu7BuK8oVXAeCCGDmos0XKh1
g1XhvdmXibX2ARqlIE/wTK0dVAwWAhe4XJkUq5ECezceE/YT4fq97kT6IHXqIfNK
0dae9dDJ8vc2tggtt+Utbvc2JfLyJd4mqHaKkV9LXHCnIbWQBTvf3PvBpQ55BX4+
aU53dMkcXGwjiVyOZ+pOK2SM3SHcaRGCeZR59MHxjb/NzlxV0CIncv4AGPUXaM7N
LjGx/99AfbivmmcLoqatg1r+bGaaBmeyX2cqXH1YoWxL/nuCij6zDYdbmre/k+a2
Bk5fy2ql72HMELZNlXqba/JreQMJx3u5OqqU9GYXg7rB31tlcTNjhDyoAsQIfPjJ
CVKdOiVakjToB4KWikIWiXfsBn4iRQJqzMySGCXLN6LSJJnJ2QLFMqF9atm5aQZC
K080Apk3CwrdrMorLtPhpai40J27pUxieZnxOYiZUzBDi4WFHyo7HGY1OcIAm6Ts
zTULRQzLEqA+90k7WeeUa1vP28Imnauz8AWqX6iQDvvU7juKmK8YztZyBrkI9IqA
XGkC6nBduzn2ioyMOwvOKun2uegyOs78iQUsyEv3Az2NnYsyElDI3G9Uv9GKVkkb
b9kWRKCyxupsmzrR3OEhhEIPNpWNs3l4SyzChBtMOo3qudL0T0nXrZG7Hjr6YV5s
OjE9HXcHhdlBDYylUKZKBLG2/XHx898ELFni8kCuuvhMVo99F0Vn4DJLw/ykbcYd
Q4NVYJjv2fBVynH0qSdSweNrz+Nr+Hjj1kbiAfO46VaBHjg/sM09/NcspQEefUzp
kfz+7TQKd0rwhAYZQnok8KaXR5BrXGLS6HUkDg1HJmdaehRZ2ZsBZ9FfylSVseSE
6+zXJ/eFq00sSMJkEVAgrZgPRwkRSEN06ILJ33dRRXMG4qVF4t07h9ha0Dls/0Vq
vJwFdXaQKLGTzbX8go/61c+4PZo+kO9hKIP24AlbTnxBuI2UId3YfcIgrIAPX163
2/2TRViLh3GqCKq06BQX6BLg2Y/e9yeybXfZiwjQX2aeG85S0uaY8zYG8r2goirM
Z/R8zaiDtJSsxIzaryYmxshyq+eIOPyUyuhbD/KtfFCmriOQRbs+alXzLC4iqGnd
mg34SL0w16PyBZXJixIqyyB5V0kE817cf55r5pvSfiKsosOB7S1FmHCQ8j79zrzi
99XtnEpN18qhYFavq+XP/GqE9e1UK7oHRGIIxNL9Rtz6N4BN6LgkyV15XAwj+S8u
pOpZYAdI0WS5+mmlc4hQPNqJumYQVw04VbdtkYs3WMtblZKuEQWnww8QbphmhCLg
F9SM26SbWdfmQ00cydUXQhJ5+qQkX3rfawOkkVpPcnMZhNqD9KdZ+V99GPJH8ZsU
aXtGSk/UeDbUvMKkz+qTcELGR/8fKHb9tjgQfRpL36nxYTO0uJ435lXuQHsBjJxB
C+iXQWr7/QsBtTgQvDecM1JNXriolUHXb/1d19emeVMlaCjEGj5Nr1QPZihfaML8
nVq9zyCKKHK+D6xXdG0HBTkElnQo/ZvW93tnCEyf/2lTJ4rAl4Yfang3qPPPAdgF
ZpYAoILthPUZerIxjds/DzQELm7ccJRxABELJmmZR4tfNbcWrlt0sz3Byp4dNAkY
HO1xk+oOcj7E8B70pdShAWvB/kJWqsYZcnaYCWnKxnwhEYxS2xiY9V0ua8iew94O
dsqFK6RbyUwcdvDBMb4JEPbOyjjKZizpqJ7V30UQsSCIOD2kBwSk46VpDPutu13K
oX3WQJwhaYHU7dsntBbpAb2Sv7H5feWydUt6/Q0dBy+SGOTWCk6qw45PhIDSb7kr
b2J/lQljT7cdqEQoLZBZ7V3qpc5UO3BF8GpEnlh2DfJ1dgU3LQLP+ZV46CKMDvZz
k5CnP9uTmRPC+RbopVQm4Yfhd8xU9yaAQ8291ve8zUeoiSUfNJAEH7xzgbkcaFlj
SRaFllPowORRmYVBuLWqOonzp9XBT8V6XLQWA/3h4ENo9YUag0kHiyIKb46ImaT4
ZxDwF7tzJ1a1XQfVk5z7LWEUb+TiYXEGG0xH0rQQhelQlOC+jHd7GPEtkTZoXvEL
uuwlmKPPFoxez+o7aU0i49ZFpCkklWZyD1b64Gb/CuYsDOXOw6G/YGrgNkk3ANVA
e/53CF2PrLyBc6qX60YKwnMx78UlamvidlG6woJ7KWsx+9KPSUCrZP+4tzbl1m0o
iJY53AWtFsps6a41WIQ56MsFY0B8fQS+6aC8aJbaIQZqa+QW8mC08IFfYk9qBvui
rJQAHgO/tc5rwOK1H8avRKCD25uvv/8RbQVKDbqG0Uw5HAnyYGj/ljin6tGJ9XfW
lasiDuCptRyn17ZsWiD0H2IDrazCIo4UNbjhHRWDtEx7xBmPN5EQf2FkEqyYKHzl
Vjr5UuLgkL4K7Ll+0fvJyEtRILudDoo+GOBe7yl7BuO4Ir7y1WcNxSzwIn1dbfzt
ZZWIdpcuSlfoNjH7qM7GSB6KoSPCsHuJ3VMrLYT2zV+sUbiCt1/oWiyT/48dpGrn
WPOuewmzjRStUSeLv9EcFqKqOWm0agzGs0lj/Ob9amsqdf2u12m1VYGSyIjK3z9D
QfHlrW7d91BfiFFUaDhjQKWhbRJRAjPAAmGksrWXSrM4PniBxdN8HCVDkFgWqeq/
Rn5hYgImNWS8QFbyNeVH2smJu7F1ocwdxfbKPi9lVqAC0ZovVCGRgMbA5v3sEZRE
EKNQYb82MSUSFoOUDwDo65aizVdTSwXUpP0IjK4sYWNsJri+xtdkBZhVz236W+IG
hNVtHIX3+Q6kA3zkhCmKk6Sx8b1jWNSVrLJF9QaNP+TK6KMm8SjntVpua+tKeBDY
r3ZU2sd3aNb563IhEggdua3qKToS25A+m/tKQxqf8cVXsy6vSToO8vPDHQOtSUVc
+iLSDy9WWw3EvkRp+CX4dyFBl7zTbOtKWcaWL3V9aDmKXmVnh7vOsIEtWXIx3/om
QnxltZy3GS0EXWF2BiLeDFHanes/a36lUZHWotOhhths36FUF2fMzwm4CgBnOzmr
+NIrazSsuf69T95hGpHc27TsSYOPRce3C8iK/FQxtryH/oDVgZrX3Dhw8pV0v/1B
3Cv6rNGnjpT9ga9GOveINKBFOaPAcPuQOUwwUKDnyxdV3FypWLMTY8QcbYrcaXHS
QzulMy+Bsg/lk72yS9Qw5e7m+BBxhhjCc5Oo2pUoePn+AFxXfEv0M4gydtCE1t5f
/TpRUAe+s5gWCYNiq5rlDNlZpplMv/P42bsVX/gz2GS3+TADR4ITHq/t5MxlK8Sv
YCfbMzFbsa52dQNJt7oZJxqmeIY4kpeGHL9/3ep/aglMmwYJ++QzHcAc3+/Qn6sU
blvHDAUlKZW5YdiYlKFyVkoiijvSgc+oAPMerPjxHq/UyPZizJHQVY2P8GIBWrPs
9W/4oRypS1Vg8gEY10NVQereYnql00Cq9YzuliisvT4kT8aqqbQq1B/8yiH2YKL+
5QosXprHjYGtjzQ7XsM32VMfR7JW42wzRav4Hrdb+aZx1IDX4Ht8NpeHsaxodY9V
jBebXixS5ylSgTjuDCoBVXXhpg/yZKBRzB6dDYaGaCx5kNe28hiaKhb6qsKy1ynJ
3ndJhGla1B9a6fhDTVLE6JnbF7cn/KkHpljogLLaanqnagQkLbJrK8M3ZwK8Mhdg
emz/U2VpskJDORK+no/+ZXfOW4Z5LS9sD7STNS8KnAMAMXWJNPp56Bwfp+1D5KG9
T4OrYaisMt1cnbud5TtqoM175KYvJpx6joPa2ZP1D6v+YWxZQhmJxcyoO1VUdGnF
xxr8yvtiMlRjXNaQWSf9xPVgc0ogdtFTJKdPqeRqiIVRscWqQs8gge7I7bPEBSSt
ohWpSe9HGZaZdAFXQnX0cytO3/S9/ZDa2B5txUnU818oW/3eghT3MIIxOahsEqg4
mARghCNp8vNvrRSlIDE90lZfpVSF6Z9be87mdcZvsC+TxF+eEPR4twRSvBlBRwWA
/7Xr516XHakSjG3Xe6sr1q8+SADq/nnsaJvVXf4VLcleGsjkTJ3WzLv1Swi1eyTS
UHBpJHiIhOLmF42vVvooDOr6aJUZqsI3znX6DBrzKA2Gn5CHFFA2AKCxDDwCSsGl
RlfAJYrDTSytS/7BxKPINiKT8n1WpNVmQdQ8Zl0DtmL3CsdcOCnF/j+l+Ykf+We+
icWQWi301WsnYex6bGXnVa/YnmOoOX3cLqZyRQX6akY+C7AMGo3FPtc7beOczV01
1Y9gzE0YL/UrTeoxOfL0567a0mdqx6b3+3oQgUoaB1dfha0P0xEJEumPZLQMX0RA
c+7xo6JUQUKPQ3bOe+Tsh3dMKJAPyk+8U4W71+WllCfWSYFcFBInf78bc2AFPzjU
ZC8f7gl280ooEsm14Ul4zuVIugzAAyMo6u+MMvul8oTL/yiFvhw0867t2Uqm663g
RwBB56bUaQmeECM1SjJ7y2/elP0zoJLcvie5KFJh9Qp9vWbJsR4vGpHLfolDpPR+
b+cxEY4FX7cOQW8QPoAaf2+tKWWX/mJb9kkTljk5KBEKdze8FCIug9tWmnd5am3j
KEiQQp1RtkXgEmcOuOhSk1u6rUHMrN7CNnwboMlxjfLO0A+EK+PFLnETMh1UF7u8
xeQKyf4VC7CFKp2jsgYKSz+dBtBzxXMkvPhxKasTpZBJOCD3EukSUXD5GTCtaz7J
CwkJIEsgVK9KiN07dYityW488Bqb/HAEQW0OSEc/0nn0yIV05MeG12Al1Cg9oM6f
IKxaL/18E0uuSeBGUu3BaHPrjp2Ywj0Qehu6dNMz5Twr+d61k2YSOeHCVAjs3KDo
SYQ1lMZGZ0RgtGa9j7B/3J56vC3sCking8AHt7yYu1MnrQp1PqlnzR08PcliV4R+
cvjYPI9xKykNk+Ygyb5uQ36U5TPnekQ96A+CD3JT9UJgGVXUe3D7AD9o5u16Y0wA
RGVmCOg03RdOnxJXSeRUa19bGCr6MhdHuqDTwH5iWG0fggU9KTET8vAQ91rp55gO
rd//ZmgTrX6IYMq/zSZg15nVNiAE8UYMGqtpz0mQJWlrG61Po2JvCxf9pWH0b4Rm
wcQP3AR9zo6Dkb8XVu9EX12CCr00bq7Qi0Tc3CIW41RQknhJZ1TQaJJ114L4JhJs
M1QCpfzXO2pw4EwW5cEJMqqFvBSGqEujyqmoDBdfxrGY5ylHv5/Y+Nee38eO9zsl
eS4hf+sabp/3TZJ4IHE/9hSZTPUalqYH+G72yN6hjftV+zZdnf3aLF6la8vrgOxA
JgXwfuMNZ2e17YFpCLn9XqTNLuPcgFoTtKpxiMTKHL7SbAZEFbVPrdA8SINcSN43
IiC6/ignj0GKkKTct3u268MLLHwFs64nXvb1KSmCh0Doz3yoquemsBS92Nx108MN
VneRMFdz/Ka6hlK8jML8aTPif+j6iqYcjeTDZ19Pf+vMyV288rZiY1rcIz1veByk
q37Txb0XASwTPUzrjKEfJz7rr8IrsqNbrcZGnTOdZnolP1szF/P9XToQXiZkk6xs
X8bNFsfs6SGiKbBwOYqO7U/HIo/Qx/8JyAjxc+d6728cLu9iWckM69ABsxy4PAsA
mnFolsx591gHi1FFpgov+8rLm+ENxYeLo1aYnd8nE241K4MyVne+19OfFBAp2HYH
JpXmMokeB7wtHiSTShYyQEWqjYteYVc09T4g+C6kWxA7vow6YRxXnEROTt/m7uIb
TJjEz9fyr9M4Pp9S2BqtYa4soAZKQvRRzyANuJ5DRUYH/++AbBqiSjh6SofoZt9d
7JlpUo34imsnA1XWq+v3JSr4xDAc3pL/PS6PKiEB3W2JZeomZH9CbeXNtK6i0aiI
dF4+PYWICbaYVoD9/B7VkJj5QmQIM8cfcgaBTZWuA6bl43TdvPlb4YHq7SvzaIDT
1SfFWVqKG5TyFi02xggi3bNQODO07X/xpqAC4w90iZFuDZlXGAyARp50/JRe4ELG
i7SGJGeqNARHOBmLG07GZPIUS/VH3LNQGvKgUcQokmRMLmQBTJ//wE9ZqC1ulNTH
KINjhebKNxSgRYu473wPh5Bc6iLjMn9iVYgV+B83tKH7WK5hsYPbkm/R5ROlLZyA
tegr2/PRJDSQhiQWyxS1HCrKWpZPdcBeB3t1FhpeNe5N+/RFM9+78P3aIqEn6HTz
In5YlQroiPWz3vlYiuUIy0yic80A45mug+ha7z2BSjMq70+C7Qxco6f3Zog+Vj8o
bB8cFTolD2C1LGmygl08OMuPjQMMVrhAAh7zDUqNuhto2YPFuHLyEg1WhCyI+6OY
OsCFHr4SIIgRs4QEZ2SsujXcbGnOy3zEr1y+XyTQ+sVMy/mOY6jjDgFnTtcHxLY1
/+4E10DrmA4xI+1MYS3TeLyBGGdgNXnLBhIN+iFmdgZBNZWQTwF/opMfsoRj19Zr
PSloT3WahOq9zDkf291sBQoVYRVJPgsBC9Xl0XsVKE2GaIII7lT4gGgMP+2WvhWx
5pFVOKARLP+3e1BVvdwLg2eQ/2/jcQCdP42sB7nj0mbhJ1jJv8VgVUrzU8X/apsK
Vh0bqHZ1BajDa/fG5+GF3Bm11gcqlOmX3G68B41RNVN00inEgHJkdVGX2e54la4c
ZcTNmep7ylUDsw2GpS8m/7UUSLu9Cl+R7LMJN46Uf7dIgEyNax4afP1OQmVmkVgj
vf9kr8si0PyLjSoK4FTrdMZ6yvJXz5hDCEWoG8AXiSPxIlWuSWE64TASUuc5pvME
kZr64EQl6PwgjYIcfpaiP85pH4+rBXJ7hbQpKM+KOkW62p2bZ/KdiHnOVH2xNDSS
+FmxzhMLCmp3Hlj7L7cNoUdMX4JIqP7AAGh0Ubk2d6QLJcQzmr50YdtmWPT5kzUp
5mNq87H0qxrSYODD/gTB/CdFTtzXHRTYVg3rnSdrN2gPAYRlcbwlmj/6iT7hi3MB
i4cg0TqgkD2onrddUSKMLZks39BusCgATvalxODGpJDZ2u3MjK/YgeyC+ffD0ceD
lQXFwGxgrdnqzn8/PtrqA7fUIXeBLgzY2SXvA+bdbXqMX2frrWpJMSYn6phu07Wq
IdOLNv0q4YwhrdQVKMSeb48LwhWQBurlBWhLZtXE2B4sXMlVhRgjqfaMzNvnVf5d
vu28GgG7K9lioDVDcsCCZqgn31g7dtxS/0UKdYaOm3aXuuo47juFFPvcW1M6RnA6
UasvHjcJFUkh5wGPiXxs3jPg7I95K3iSVIR8hwj1OntylE4YKZ+Kye0c9NWm4fiW
x22E+prRLk5RkP0xJleKbeei/W+3X1kjY7Ey0amXzRsTe+UVWfYH3Gl5Oj6N1MMD
k4FDM4mhC1/VmBfonASYFxeFoH6779YeMN04Yd/urZjk3q+gv70rCjO1YQ0ZsPoT
otA8gIjbVeeba52+lCG3aT1JgGNTtCKRJtGj6sQ2JequIRpEYtQsWCBknPulfC+U
KH0+zXdIPQzwYqm9EFW7PMIX2reCUYdgiWqguRkWn/oosVapFV+8/WJC4zWmsASd
vakCmvRZlUWYbf/lWKI54F5wCe11dgPSAOSpR2VvzyUkr2QjMDksnja0jFqQqje+
qdbYxx3cpI+RySnYTEiVE3Dxa2tlflYnIfxvuDHz46SwWGO39NmOLhgxw6Duw2ua
jSZHTZt1bJ4ENbEHXXCdvBMSRrD55SH67VgVsSwVHonChSKOWj3q+JM0E6BOgpUV
51dH7CKzBoZ1lHAh3/KQJihf64rbHoksGw4YAlbd4qmVpyDU3Pj6zaK77r1bMbYx
Zm/3qb8LrBKYpQazlXIJbss+5ot1kgAiPDKGBYNAatA4n1HmqIwh6e5DF2tBnwqd
NbYg0Yc/ZOYISZtVJj17NpPFP50akKXhoD9jFUq5eHRRfWTYT+hzbYbsy+dMY8tu
A6pZ/eT2IA87B8dEwbBDUMlfVKFJxLSDZ4Z/zO1gq7tX/z3QY5FZ4Hkyyb2E4hp6
r0auEMszqLRFZmQqYDWd2UFLMw3TIE7ZQW4xRoLQ3KWXpl1SNIFlWah51lpLYHQe
ANtw+s2jS1xfFFKmVqF9LsPZotjnuGQXe++6FcoQb6zZ1EHGkairiO7QqyFFhMGE
yVU7NRhfRLEF03855jzcE67DYdqodckuB95A/P4ToJTUR31+i/itomWbslU9kh80
hL9YJ8EUbwSGJyRSfdCBleLDlahzsGejkn8O908k18GvKTM9XTD6X4x1Uiz3n9Ia
HNxlPYsbrOHRgCA9V3rqIOSd/ZS136y6VpS7Cn79vEaBfjA91LHR6iibWonuioFb
1wydLanEmyCqinqQG940yPrMzNaazvAy0oOJa0OQvEhOQX9qoQmWiJbZF2RGQJCY
S2LhzlrcUa+epohcJ+6FxYErNjiBQmJBj2odFSj6N91/l+fZTrWIHhBcHKpvtHSS
QYS5eITSlVop3HE1LntuV9AtGKsK2KjuKyx6jFYgaA7+8+rwSdJwpKLucd+zzY4H
x1yYx57mfEGyVm88YjFYDYyYZIEK09YC3dc/xEPia5dfZsXagcHsMtFwC3JTrpGD
/jhhHu3Y3q57HFsC3UwjQ8keYwLqZdGq11iu6gzTYYb6iZLsBDuzotZX2xkp5Gmq
Guf7jB39QX25SvImyMXUjxEn0OkHMMgop5Dv7S5/R8FpGAmQTH1TMB7izAJW1Qfc
9wHMr5cfM9+2z0Y5f8Dlo5JUxrOud+86wXeOqv5yyQInwJBcIUe+QgxP3RY/jP6z
96iwF4mBrNzVsRw8ZeGZfDbfajmSeOcE3bcm4i4umW6kfA1BPr/n4WhO2FNGuR/7
sMxwhH/Y5v8Edmd75WH59ciNxYVlwYul0y/W62zogtSSVYzkBGOw1KnYydFS/5Zm
3LY7kykpRSOyIRn1fBso30Jw+hcg7z3yrMY5E1DOr32B5N2gTIcoYT9VNPehM6ru
6BvzADy9n0LBiJ0NwOQ2ZKrXhOJymYo+d0VIcWcA6CNhRpjBH/Hnnbx0HeGP6PDE
Z1vLHlKzsa22QLbtVgBnu5jIP0nRVE0LywKUkIZ+aRGFv3uj1HN59U3xXyGeuTwg
7MszLMm33+E9odPB1byGTs2mSV7qVR0duKAniAFxmCy/VEMMOAo4zZLwAkZ3V1nc
zfIWsYWOKWCnqQQme7lxYu6Y9wfHoEG6NYruGEOP8qb7XOY6pUMk47/dZwweJHtp
kp04IWExFPemrBpNDPAA3OncYG0Sw1vFwH6u7OwoOZeAb5dfCGM3ISNhmvIt4AjP
XC1Rhm6guKwFvo+MCSkuYxHM/GpgQ6CtULe6L7ytNqaCRvUByCW2bk3qokhq5Vpc
j+wv2QoVibq//8UdCww+yvN9DnI8ORdILEalg4qmEVD3AgB/gf5PLoiCmaoO+mwU
mUyCJc/B2HQ6WBs0CQMpQKCEp0Y/7NE1eaNLQYOzt+Fjcm/vlubgZtygmrOjPJ25
ryM939aGXbi6PkK49NmArBEnu+0fwZ+YnOw5Kiia5bVDNeCSdkpN35i5kFbyrXZP
e7KZiYrMMdvch2phG+7+ibBmhlePWZxyBDLR8mbT+TZfveCkmUfM40apleP0a0Y9
iE7DwqpCMQwzx3L5dpyzU2WQr2E1CJvCL5L1EpnwTvufuP8ptDUVskOCSwY/sn47
prgKm7bzMRiNDMFIGL160B/xJPxIjWjnbE+M2POQRH/aCvLVwsTDbDz11FEcak//
bcLTDORQpUl4vL4muyE8N+srepCBvNqZZbr44xrL4/hc2KY4ofGxaqK6LAGTq0HI
o2TjpA8fh0aB6TWjb0Lo9HZDXQkhlzcCht+54SuPOQOfHe4JkYvMMsemNuWXFV4z
OSr9vXrPNgKDJrctc1uc7qLX7/Br+vBb13y4V2PpP6cOCHlx/FcPop5GW3k2/AKe
P57p0G42TzO/ShTmGl5U1hRsZhLeFyRXp6weDaRYdTGORJXEP58K1lD900OFYqMr
ilEh5k3eoDXcJARwKmvHV7O/Dc/cJrGIn59EhR1KQbDjB1crx/5wxhd1YMEljV4x
Fxh9KwVSRZe/M5Hw0XaquvWu3nTsO+5imff3aaNZ+eYIkr+abA1jJMpqyukUxWY0
+bw9GTW+YBsgiNf2a4G2BluA50nwdRtGmRteOO8dMU3ZbEgc0+ds/SnXsi7t+yVw
bKsAcudNSvuqByYYGkc8p5CapNqtktLh5Sn5lopexanJKHvO+g4HFZoONh+DBcC2
1te402aOPRdQTNTPsq9HfAzb+CBKT+KaszfDVPHqFjLDD4MgdTC7Hu6C27oF61Y1
z1Y9zs+dJOdQjzWfjClj8vVt+7/IpWjKXGW9S50sgNrSVo7y/eqI5gVIQZa2Oexl
DvwA/skyClTV/7B3Quhkco4i0HvnWELzx1OWR1crmJgqoornti1DkrDq0Lyrijgi
vfgKeuDZZ4pWmHsmHfYrdBsl6bMPMnktqFsBYIEvodwVXrofBxSUoJVZDO9rtRWb
/Pr3LaYY1BfhMB8PXweWQmuZrnpwrDM1Aacep4A+bXY4ebHvSYWJ0NxoHkI9Kev1
sDiNkarZiuqmnD8O+fK7ayUQTDwEzMjkaKcuapjh5iK1HLjbqRX3oTciKNb1asjr
brpoXUFXe/axTUs4E3yCHEgbtXW/OuGkejlWsboIw0wnl03AHVDXWIYmi2RCICH3
5yozp1jL09Mgbyni77OyzjmbspkrAImZhP9y1K38loK0D828FRL8x+Qk7m02H+CZ
SGzmYMfU2YY8hGnMbhD2YWZlBUahCjOGpBNmWdStqpGl4P5zkJvpxnY2bXUt2Oql
w2lgpE5CxACMin1/DP+F9VaQJo05F0pBImA/MNXO/Mjb7xUaxrdOqoLM8HpjC60p
11EjAHRgreT0hofffK4h9whHU2O/wlAzljCTzEaOOlOio4k9q38kVQWFPFP3Ytqy
+wmiAY6jEt6QmxqyMsjY2CFfWyYL1GaTho9u1KiKGj4Jen+0R76L47NmvOYGNoyB
sOH6ni+Xs18Lt8v13KYqd3uV5+m/+d9bVSikPXPboQyxbdA4TrHtWne25bl8qFXJ
Pyv1XYhsde7eJg284FDNjGxxNVqyHMD9S6IWRxWzF0K/zdlhw354N0kVA27U4qfu
N5UloAETBXTfwjXWXUOhsALjcJkhRkVuwdygyReP8fvsRVO2AF+BaGcYmzlOlOzY
9Fq9EpG+E1d3QJPoiZdWzkyW9WEtVh7scCLTd3Zers0ggHX0nEgWw7po0L9XLEzL
pXUgjQEJ3+ay28EQEG5R3YjVaPwRVxuxkptIMIqfV+n6W7Ct0kT7hvrGAAsuK+jT
QqfOD77R0q5uF8lfWmDXROKYUrDsYKNDELe250uXvU+0lrfLlBt4nn+QKu4l8nR1
LEhiCwArpXx4f/aqqCjBEGOPiDb/9DNFjsiJzJ/BFLFBQHOsc7Xs/r3DL74t7efl
q3qLiP3ZK5R2rr9L7OSD26kBoj/BoGwkTXlztqmJ4rQYyPLTqrJ3rUm4sCNO7E7G
pCa8Uks8Va4yX++f61Sw8r2x2TitkUjR5/+5YrhzbcuZYsbDkbhGL0eFY5rjALUu
1k2amgZAmP/6mGEtu6inVudQhM1CFZJp895eJuOxQmvpIv35ShcscELDZ9IwdGHj
SyhLw+JPD1DG3lpSRy0U+qLLpp2cVMo9MoDzj9qGiUvl2CIURPGyiAsxYHtjEGnU
2YsyIaHeDaWVDX9txxgxsfndQhNmnpyA2GP7sKoVUYbqEWlN/zflAhtn8P2N/SGP
fObyOlmkx1xhIWxageQ7tcanvEj2VxkVECIVprh1zfO6Bw0ECZECdFO8IXohY5mT
xo8olQberh7V4QKzEzNpyKzmgUcF4OZasuQSdUX5rfAeDtAjkSchoghWVayGal31
DHVhcHmklFa3emg3RiZn7HRC2GT0cI1j0v0ncPjnL/XKk7//fGUwyJifT3+eI8ZK
nrdQDJlEst06efqUhyucJuYeg5ntNvPHGE1dqsZe3Fq6fOuA0CkVE26wXy91lt93
8NczznjjsWNoDkMtPvfbNWwL67kRR3iP6PS6LEa4lZCl6MQEj0HE669bQJrvxez6
aPL1y8MJqyjGkMuQ179jbXcj0edxu9ajhY1eB9mKOxXMSYmmywUH1i+FSl2/UvqY
CiEFAYbQ9BC8zibTN60UdR/SfzLvCTTD8QJCUNRgDs2ckaAt9mDO5xZZvAfXTzMs
jNADnxHjXnmGJIwWsKKylM48yzUN1lyI0NiHA6qDrIUs6jiMhQ7QlSsuGukgz7BS
/9DpYcQLXjRT6FygHqyc7WctEZ3LcdSB0egF8+38vpJ/EBSNBrvlgBp3Mb2lRwqT
/IdWmevEL+KgubHzNNsJp6uw/PPzkvbBsV31Zgv/dFH5YNl0YonLGExBQmq0tq54
+w5i4kG91AzQMFwSOgfYN+B3h7qY2aNtHI4CuCrgFU0AkFtZWaLO7dTO06twWevG
P+8ZDMvuY3hGl8JqMSQEnQFaQ3EAzdo1SjpjguSUieZQbafi0SuK7fsR/PiLOKN/
TB/WqQ5fkXrFhO21ghhrQg1/ut4axUJHkX+tagmyddQuY07/Y/sE+finB290zETZ
Uy9dlwG0KNxCo+PMHSlOIhEgxeHtXgVCxpiU0U6VdRg923XRHGO6DnX6+l2XiH3R
8Uk/U/OeWtX1LH15isnP2HC/lLYSKAtdl+8Lc/FGAc8YQZ521AtE13snfQv7/tAt
6iNWYSja3kVCK9YQOaeoo+PUi51ZJlHGDs+4JykzvAbMzNgdseGoU+Wgzt6obIh3
sFCCJk73f1y8OS9EAakw8y1Dt720jGZcKWMlKPyZwE4E2Tl1vFe0hiZ+EK20j0dn
LMg/DmimWM4eEHsgyIcIN2N5lDvL+CowA/h7Mpsy3X7G/MgkaY/p4Z+4Wk5ruLwR
uAo2OeK6jepEorUI5AbMRfqOauhgslaG6xQwdzN0Wj54Eyp4cQUeOIXIy6N+H28P
BZS987C9nrxFxQ3nJRGSRbC+qAXfGAX8WEZreDljPotBB3W1uH2v29O/KNXaA9id
ZnGAMQYQd4HEmyMJSkOX7uUOFbI8gCK4mI2bsXdDTskgI/TH24xzC8SMnfmcNrgr
idPIPiexj26ErompJg0giNVrQS1m5b3XKlpHPTQ2oRkZYtJLFuOSQ+tTAs84weVb
xIyVMxnzhQdc2YG9LVlhZeqX5/kLbLwjY7YqriYV1TFUNiJYJJJV4X6wFyE+vsyS
MDuRksDJ4lYY3oLWx5DUTZAjPJYzUWUqa6xfxat4iOWRTlB5fUfrfR/hH1U2uA9q
b4LI9NsrfZbTdu2b9QpKr+MFV6tmxukgTqQJ9CZottJxvKAiNSz83ljCWi/l4puu
zTRIHOx1Nmcli8vciDtiR5ylmHwxK9dC+5XQIC7lArluv4VM/vtOJ6V+GRRnOEmd
fm5xixwDHBCmVpXgkBix0ZFs9VngiNurivomOMoMysJq5OktA0xZ0prYuPS6/pFU
SfUFByGmw+meC+YzhvcfeEgem2Ik2HSkoJePlJTBldALuYZko4GOENbCNC08PlTf
mOE+086t8P0xQzN9z2L8F44gvinpZpPyxYctV+8HDh6SDErcOHbuM7LcaERb93CP
HozMtnHUfNMtw4Dp0k+ItKVkpL+zUM4+4xNnIJz8RaihEvSJe/dlU8qUXS5+Zjjy
pGnUwBxNg9aERW83+fMUVt+u3rnk1eevnVp/iqRj1+ZK2T6j4JFM+BNlwI5E33rS
hCNWz/oQMhQzmng7jkzBpCxmrBnl+s4SKeKq5nzuHEXNmoJx7Y4+L6K7Rx6jm2AV
rjhQnsQjNx9XJA8iaNSbhRz3Zx46GfUWWouNd6YEd8Tfoev/wONp2sUn3xYwqOsR
A7itffoQBXqo8HBw7jNPe7xy4NEjSJxXo+qmB9zaPfr+34yaTQqfrhIb5kBbXx4g
AZf0//viRYyrVjaMGg9lNiBaAqdmJ19n6JKGe0upeY0ZCOdxL1PG6kws7d3J+ylu
SsaZLHSRIiV6vTEAlwRwRnsPAJi7LGMHI9hL/cgRLKaSXFP0Zn6vC2Srbi2FcixE
AiQRMDa9mvARieik7U18r5FAAbCXwAtbiG61lnlWzwf0dbtnDMR26YtrEtfHiINf
xHFz7f2NcWz7USujL/OcwLjqeru4X27eXtO8YDvOuYPEVKcyhycVb8ODbEeQUGYF
KC+axvk0hAL5/MkFLHyDPZg+C0uL5xLOuxKB5RseYXy6IqAwetIDnsA/iWUPaCCJ
/Ycut2QhLtd6hrZDuFppYThUK3qfpZW9DdlTmvuLFp3hOiT/A0LBBSYmkYF74/iK
gnDFjUSS2qxq+QRaao4qT4JjhZJ2brJvfd4Vh5O3fSlVFLVcFE3f3UlS2VtUqy6+
dDCBH/jqNYulIYsVybdPjkeRBO5kSwsZYwomWtkGdmD0T2xfcA6mwaWpmSFV8q0+
Y/88vx2817oK7o5XSfT/OsWiitF4IF4dPLT231AsTcdwzuq8EWAotnC0XT3wDc3N
MnfTW0EdZU+QSfelOiqYuSH2oQ4mzCTGiUStQ6YTseq2LZUxtworsUG415XNwy/i
0PcgtacNb8M3H/mJ6kqCn8f8UyTL4BSN1IBYbXFejkUerSV4mXtaLqEtRDqVmqHO
HAfuF3ij084xRMu4vqwEn5XzgWrC35FXS+AnxP9xlhSUmAYUwVorBPV+xozRp98g
72vZWyph7jlRTOUAl+l9BV+0u8Kijhy5xd+07bVk+9mUPheZRGnXu0HAMHt1ZiIM
AufAze5nT9LFvGsrqGWFVKneBiDbaiPEUeXelhr81FHAScCyilQTbkoduxOLEP8c
x5CuAXWK+nkVs6ZB/Yv2WYOlMmM0xQcbu9+v2t9OAd86OKMpLCgWsrBlVbei6L+N
m4tKRnX2hiJuqh8rgEC93n8KLXQG3RHFESHOtKVxbjW/GlVhnUvh0Wp/amnmL1GD
nFBFAKiitHb8SUMk/IeL3bqM5CYZi/f94DWSF2RZuOqhCgGYCYncX98SpP9KAXuL
oxj4/M7WQ609npILXO05E/WwGZS344FCAWygGiP6ARp9dvnnlHaemcygxN0nx2Vz
C6UQNtDmfXdKf66UQWTSLXx0B379oFqKFqV0QW7qHgUZsC9GZms05Un+SNsVbePJ
TmUfjCsi4uZFvnv7o749nTGT3wDsvUUgIGtRzGhXL30SBzLYNk8ZLM/Bt6fPhHfl
Uw3jF54uGxsUvsmA1zS0SFXLKAVFG7+vOgXy1cbymC/Rfjkz7C418whoeMGYNGWC
eH5m2re0Bx486owXyV/DDKH7u/cvTWgDAtzflqBD9RwhEebRGWj+zYsvABVpYNUR
CRGUFLZjh/BEel35TMozUxEowmafD9gTgoj98If8r+Uwy3JrTDW9IdCrlv0vuipN
i1+XRkKnSVoyFFN9TxP3Ryl11AGozHcKGoZ6F2bcPnVkfjFPxGKUzJNH2nZPCK+Q
YKcepr5D5GH8tiw8T4jNB+jCLoRK5V3kW2bu2OMA9Rx1M14pcUJRAMDkXhV1JrRY
+EhimLlFZtbhX5+fr3y2SiYcW/4CdXfjCTrEDwOA9SZyKBpT4bo/0+H8Iy5HpPPZ
WDVErtnooFr4cDnn5jzzPhf7gfH9pxcYI9Ab5MGs10Y98qWF1eNmbmyQyMoGrWRf
Teu7CocMowswgi8q2LvNUT1oZMOmTwwm2ixeimpjRO/iSR7umWhJSAJmKsEeKXI8
qAHYpL0l22Ko2g5xHNr4qsO7bqx+AWCwqP1TLJpaX1fMji6Agb9jLzH2f6YjaBHX
g1tIReqviJWpgRBbAkK7Un/p2pYXodqGgz9hPsizJDc/4NkG81bIWZmWi5eg7hG0
4F5yhQt4KftSUztFVwp9/ymiR/Yc3exKxQOsSgPkHSVSOgTObS7SH6nNWQbYyHsX
BVtv8AhCWQdDRCBbmOM4EvvMxEXm1aA6yi/cg8/MxYNZxXY6CFJW0UbYE6Z3gFuA
wdYG/gAnlmKX+a9O1RconFZJB2UbPDWFFPkZnvxlMJK+LOYYFcocMj9l8oBW3gdj
6m0+bdHsrgY0brq3HfsZ6h0MEEwjQTfrUerxLkrR8f6CQUEC6XeZqfirfydq65OM
mJN+S4YbTTp15Cvr8Zbos7DDgB3D2KaQYeOApbaUWr8zvWQx/rvP5eeUyW6oH/gb
VkxvYCO44/929MC+0WFqFbE4YmsQhl7OQnHgiF4WQJ3a3Y4MWKFPfv9Xcup+radO
LrIB85s4/zxAcda00iU7eVU1LrL/biiFFUH066YrQxWrOzM79ZGxeXz9brKGstFC
q9KNExs/AgcXNdiaa0iS/THU6RkwnwGABg8qMKOzDYEt45cZup/AVVMRmuwyj/jX
q9UpCIi3m170M/FL4z5iFLIa0cSzDRBYQR7uioTgk0zG16YVd4/MkR+YLDfbMI7F
GxZstfO4JWdYanYLnYPreMOk0y5QfsovLxgKQ03gcZ/+DlbHnY9bCXylZZFQZk5b
hKnCXpySI9qGqJeZmu6+xln0qaKbjLe+hbo1SP6CqO3+5xphaCwTsM5ZGD7cdKPy
Ehs02ljKXrRCvlEgynogkc1FIOUG4yHyJzXbpvKXEjahdApSOAmfQo/Gp7N6SZYi
SX27R1nrrL/UkyFSkExuiKySzRZ5tqoBR6nyHL0aeaQWGqs6jL4aZjEAYtJ3AIVo
Iaq7Kzxebz4NxNDsAw0xhHcV/RDRwqYzXDiEEFDEDdHleoNe9z6XtlyfCOlAJlkg
ShnWhKmNDN0qeOBqLljceudu7jG3aNRBuLmLL/H2myYLct3id3E1zfSnGIlXD8Z/
PDpHBUIdnfgl2r13hs+C+YbXsTd4l5PKtSdmemS35hbYq+fACPMaPOcqbnwZY/er
Tbms3wCqya9gSls1sFdCkGTL+0HR5yXC5kACmIcUksuLwU1dCgLJWD4UZcfNodj1
J5O87fInfY6yr3WiyDDHJ/jWA03j54Ks9NRE6y46Fz7Vb5b05CakqqQLHS3uVhi6
lxlPq2IGse86njPLXuYh09DPt31GS3+jCw2AoZufiem9qQ5DDYzSbXdBU9G0x8ye
vF+Lg/T1EofJBcfvLXWpB5kRmdJL1X3lVZGadK1y36IprfqlKmpEM1JYeGew284E
KsBNmoTAk5wbcNss5fdI6GhfYWxOFj+lAAPHi4iDlS6VikM/Bgsz6fltJ7XLk0tt
oU3MAjRMTxojkeZcD7i5AJBk53TgphBj9XAvW8iDZ9Y2YQcgvuLVk9PjCkELzYcO
GIm7c3otr0DvznmD8aOvT/EHaOCM6KkupDBMirKcIQnd04frV7FcAlyRo2JOjGeA
26sbdSr7THZIvqwrXPLSaAphMsA9ymJqIAhNx0ALkmhS3UcFdOEKXu1WjzxrZuDJ
kyJJZMIo9ZO97dQJ+wiT6cBZE+G0dpaykMUmLHdshAf3IbNGa18dA5R3dB+rQOkR
Ti4x2sa1qQ5E0p2GREyjNP8wEOoWR9wnFStIPTqqEjWVGwbrh9dadpIPc6Yfg8bG
lSpD5bwVMw/YAFVgRsdse+1u8hgpHAJuN7UWIXkNG+DP9E30zW07t4qRo9+9znXP
G3EPUk4JzWeELkos5iwV6O4qukbTqwsbdLLLtpKKeXe4S/+9qiQpSGEE017vaY2B
m1wxtG8pdc6sSLDzyGFwDOjUbTZIP0MYnKJpGoxHZdqYYocVIzljMVT9NQd3ocEb
kDbUV3NCDidlJduKqDZH6Ypi2O7maGy2WED/JQL7CUYPZxCCStSUk9cbvULkDYqz
yialPYbj5p5UClaNU05n5YOjXWDuS+tBx2ItZHPR8a+/2DjymUuiri3zZkSM2ICI
FyyQbMs4XUpdL5PEVfia/ynbuzprz5bBvvEEhLDoItpfgNTf2L5dvfNzj9QSzdgW
kw4tE8B7aFrIjyiRft15Io1aWBuZDvTJf+qYH444iG5rSRxgWMQ0+T7lh1esIWYm
HLVFBf5Iylf95QSNua5ITmm7va0vzIDY8K7YYJq2KoqBAaYvt5RVH0QtKxAajpA0
rXSETB5SADJEkgEz2DOJ29WEKQvaz1Zi0sAi3DtjOiNlzFojIeeDDA4OlNFvuloS
dWrLOuXMVMVe+bXNipCGOMp0yX5TNoW4wEj0w4wMuEOdJQF7XN/y2GgaBAGCj6rk
s+z+rP4YKV1H0IY8xIG0OzE1LZ5qUrlhLvG5lPaycZ2czrhOP1uG16aDchPqB/j4
rRt4bgs20EYBGehwldG/j4mTKjc+wP0gmsuRXhKjQZC7gKTbiERtt1LlFCWm/VC3
ic2gckS8EvQhbvpceUBCPYvyaYTenaTBISLOyfBqMoeAlJ+b5SMPOKyuSfLYefHp
H4+oHg6++OAqup10wupELIyIo242gpl7bjbr7O7WG23gk9GBUk+0Iq1UM1Ucqb0+
TeJp0MFjBQHEyii60VI04SzlqdGeQdYR5Rrpnt0Kyui1Vdspdm1itZD9M8PI4OHC
vdcifRf0JEiwXwJrXZYudDMKbbfBnlXAYzxZsIZ3Yz/diU6hmVvA6mU2LTU6PRhs
JHMDzk/1mqPqB94kmvjVn1ntghNaMbirOZPK3pFmPkJfD2ADHuFHh/v1X2GYIyNl
VXXm0T2Ar6u4i9eIuDERKOXPPbJCDccGHWrWxDl50pQ2HTLBRbcWsi5KZwO57tSa
jtQQU/jgrBp9Sln9/8Q3di/zeoLLkCgn66vjtOk1SwJbVbwfNvFli61CdDkASgU4
R40DtlCiYme6UQ6bN70SgoSRghsnNCrhVk3sjrd0fSym7BKkBpaRXQ7etfRGqFkH
XFOInP1I81IhTCO/YcclVAuEXS+xsphKM0JyMV0GUHabYT+dFthirJKyKGQGTKMQ
cIJwBj0+y9Ib/KMev9GzQJj3hKgK55/ge15nLSm8rp5zLU0CMAKZLJgH02YFZsxn
pUGTsVyViNCrv2MD+TKTebPtlUMbRCiec+b39wQ8sFcxemGKNzhXBwHfIWDxt/sk
X2NbyRh9qNCMrxHfrRFgbF0vMOumsXglDLtn4gEUSOhVVHieh576vGGhuTEbO2im
00P4HWSgnG/V5y/A3TvgMe7yOZPuO0KewhCUkR569bJMQb1ODEDMkJP7EVrx13nL
/FA87ZDb1Jv1r0HjaN6w1OObTp38ufArGpwP/Tr2joB8X/he0v+Cmc/8h1aYisJo
uxqy3GC8OSrjWGhjiopOjma2xbA0fvW4wnMyKxFqnV8JrW55TU0dnsAyumKvsJwz
ZDaSl1cOnB9dPagofYTo/+2mMxLExzWJ2YuzLZCH8rKUrxdud0e018aS6JuG+sOc
iE4kfgWKLEv8V1CQrRWBciUxm3ogRqqKUw3TR9odeL8ESujVEE7wK4IW+hnuVaze
7Hdm7rO26Eim6kXywf1kZQ2JGY8HzkaAlrAaPBXvdfpwKdipVJVTPuyU7JjWiefa
eLiABMsSuF+YJVxQxAE812gN+P1wHw61fkpMLlJXj3Tn4oNBnGwbMa2LzZk93ZNG
grxXSYRWIIqsJ96gsTi0Zlzd6353lY/XspRmEDdpSOVkli91XcEW2av+N5xOR+E7
8hzk4zDx1wWTX9XIWD47D25dSgPXc1/NweORDFAEn3JUIpATpUyZjPIhGPu1cRse
5sxjePimD0wCOafmhJtBc0Icfnp8Cue0w2I78WhRjF48ss2nNyBfdkyQBxZZuXBd
ULdgAtdQx2W9FgvAg+0VOtsfRBu0d45SM6rzIGiRFPyYbnr17SYQx4VDJc1w+9Vw
BOwXYLRY4Dz8K4hXtvEoyDfon9zXCKQV5KoZ59/zRM3I6ujhvXvVj+sJDveps7tA
khOj/deTjhfN4DFeKfd5ZeYDmWPD+P0srrZJCKjEB9JWOY6uzxIYBbMWmkejw2JV
1d2PUM48Be7oTD78yAWN19IQIZUupMeDToW9JrQRUpwR5TYJDmfwnqVbXcgFGsRL
ETa6swUCelqFwiqCYyIY0uwlEKx1tqPgatk8jhMqgji4GdWkRQaqV01i3xHiKia8
hubKhCF23kj1daHTHRmbENKiNONh74vExFC0x/90Avytc1XkALnG7Hs98h5aNtlN
5y8H/3cssvEWaA5GqBxC+Xwpji2a7WQOwQcHqh11F4DSnsKdQKtxbkvnn9H72pv9
0Jo14MCnhC4rD+Ipi4eCfiPIQk4lgH+03dsZZWFyrwsjVTCQhvw+SGmal+PKKCbL
Gy7SmYHrujCDR2XEfZyKOz1gh/5Fh8JszX3RaiMsSd/3UR8erVUmjc9j1hh5ivb4
cJF/Owg1TK3JNl53hLS+Qgjl6w1jRVxWCKxLMBWtxylA9iAnpShTwMqk+u3c8x29
dwHgpz8uRVvQOj+bWiexpSP9Wj2FIHu4WVFgNNJlDhpiiAb2hxrZQhq7mSjcQ4aI
Is6quKReD4sAOWgpzDMOa11hBYRIe4IYbBIwege9VGeAhWNNbL69YqZJuXvM/lTf
1E2yhOsz9iQ3h4gNv7f9kl7kEie43GdNZXj2y2oKNqPu+jRrXyRxXcozY/wU8OfB
RCunh7T1A+Tw3JCdxorG8g9XezZSOVXDWnXrR6RVDbAXjRwDFVwZblj2lPXDH3LR
mWXWL/bj2h9ZPghR7dblR16qV/6LSvekgXjfhiqBFXvaFF9kjiCglSvKX4nILxc/
e5DfmHhmBApMjNUoNwdUV2+VzwyiqbdREizdgJjVtxtYS/Ios5WojSDtG3DpEV7T
fBObTK+UJnjA6UOFZQt6IBcKCksalsjv9SPDmAeDo+RA4w7xiqOyGAoje3RnlSbK
TdBCnZ+5hgZd2nL/XDARiJ5h6wN35+VP5iKlmwGxrU5P3SkigvY7VHMswarA+Uq5
bNNXGoJvVNdsN1CkD9FNepvth0hFo/lIpgO4i32ov7Dai+l3FyixkCvbKuVPE4oy
8RfLRSROorRowe2WiUtnbwh8KAzN4K531d86hArWeSxmBQP2abHKPiQZdTBvH+ic
9uRRMm1D6bLcQfNCBXsH5pXgKRQqfuxfHetg8u0+LaQwjDwVmOeS/jKSuQ8VDxnN
q8Kvx01P5I2XDuMVzundRNzPxgzB9V/ucmk9j3vlHRXm0dK72Hr2Ofi50a+nyGHd
dKwGdcIpfd94QZHWt76KQYubmljCT/3JAiRXP06dAV/yNLktVzyWn5h8MsMkW6GW
qoQmIwnYU3Kyrlp44BFb9/GJ0t2ol8zQC3Cj37sskc2CgWzMXh4Xt51/2tEEgzkc
65HDbUrLf4HWgfXLnyqxPbXPEHQce8SZTtC2KnFheilgs5nN/Z60mzhUk30y3JDF
uIhBjXwoNLnLbGDPn5mhwiyXFy++jPcRwMdPdC8iK3i2u29LvdIMunP/QDQlNZGn
Ut0VtELgVFL/FxMfGrIYRvQoGLjHDevgkrPRPRhexiCR65rAkmAkXAeTuxLrGbX7
NrrDhz+5G5C2E2Z9WnAIyQwksmp4M8dAeYRAvwyvr20RhD747YNQvnDubKX4up/e
QT4610f6eWk7czj83vrco/ujKw/xxjF3OBGIcJS7ezIt25nwunAxL1zXj66e6CcX
HC1cCMBfjxC9dHzdDr7oRx6H2p5EBxbrskyu4NzKM/rcR8voEJm95FV98w8K8uYF
YnwbqSsVD/R9CKLMfqJi4Q39FqG0TfKM6tL9txXajPi9M0skq4jQSnD6NDdk2n6H
fGMz90779+EWUfHR111Vqd1In3jonq1wwlqNNBhSGSeREmYWx8K81l96RdmWI+Ar
9G51Iy3a9IW35Ou8kJrdojFJ9kZs5EDzZhFu39hggVLVtnkjrge/hIZpbq9Smc+N
uXQ+Gl9wf5lt0UAYf4ZxhS7KgPk/Dnjnf5TQ7V/zwDt1PnJlLudlUfX0Frh7TQ4l
whicN+17fczY9ogIIFJO+l2hK8zsILOfGQ0yK6XocCkIXNLU4hjGYer2C9Sm4YUG
IZGRdGgIG4fLpcUn/4LhMMbKw2JpuEZia1dJJKW1yP41mVrUCMShzagFwgEPpL22
S7cOTP3RUIwoH8YOKf7gwRC29TAYscuYMyQPyUY8R+DauZuy7/DfJNkILZ/7dnUr
PsG7t6y1nObmXkH1sScoYy0w3Niwct3aAAue2LhWTFys1ZizTArIxrIV8uxa+OlM
w8V/OSA9pL/RWOrVL7+6oAe6L9xH0ysDdncXjht4F4exj43JsNQETHL8Vtiy6K/M
r0A2So7SwwIQbQaaG7ZR7WPPgYEfy0Sm475Bes/PAu7j6COUg5NkjXulnVP55Z0O
4DIxt00xaj/017p2Ic6yEDf7ZmxfqiyA5jgOBHATpf+6kTlvGO72F7ydkBCDNk8N
0r5Dkg1d45LmkSLfRTWvG9ZLXlwsg1vxRedLRGgv3Kj5w05I8iNNCKbDYrp9RWkh
1CKHIv2TE0J4jqt4SYvlmrR6GBwRuuQXQHVAfNiIdB0U9h1jWlHTmqsMWFnND8op
hYafHFzJnoanswARZ4F4OBpyP2a+BjEORiZu7v8aHPvjyQsOJc3Mg1pTwaizYuxa
cYRbgLYZcJXS8bhKB8HaLSgYyzHXejECWkJowFYM3YGPAo6xvDjMY5cIBcUOC7BN
PQeZxAkcufnSehuK0muJr7jqPYbYOoYB7AM7Ovt2cOKo9ZfbibvckaD+x6y2EmcT
ku0zCBi15QPI1Tce55JnULRYKln4Om14vlgNyjQK+vJawC25P6bDwW/1ayqDti58
fCDKiub4li5+/cCj2LD632aZRYrzpP3Ci9tln9O4Oxnflo+PtCILA2O9rLgo0PhA
pnkJV/AISxyrYg7rnqMOd/S9spR98CYiv5IAE1jSpVEJH+dMJMgOjD2EAk2FO7Ka
49GGlPytEV+gOkaedyoqPpqrJ2016wwojNplcRSepYYXpkQMHrw1arhOIvfyxCZg
Rm7uu4NIBg9ZzQtdtuKYRmAQgW1o6Nh1FsITntLtflGJDWQEX4cRtJ+VUOoTPgdA
/WYoAxITcmOVvAFBTaNlBKM44czOL4+3G6OrrH1T1RonT10zRpJAlcQ2v+fBauuY
1JfcQx3LJAMxKmIjNi225N9k5Lc1sqHf16NaubpKsfP2hBsEUzS395ABMPVTdYGB
mZchUdOyC1+Ax4Sc7NY0o2kIKxqGqjnn+9vd2aaakf/fzgTprRwJeGFJ6KJBn4+f
ru1PlklXeE4i03PWxyKhV3kt75rQrs1vRizPD8R+VIGfOTp8mlj9e4lNFTslSWEk
rzSF7nwGDS/nEpFfuZb9OuU9Vrfy0pVCOk1euXMMW6l2d4JPQ5A07hYas7aElGuL
Gg2E9MEgcWQOG5CJS1Bz3Ly72CN430ufdc3KTFaxRcHcyZ6saAtBLk2k0GlJJNCI
WT+LSQZliqylPCp9yu0axIKWmPshZQYLk3Ge/ar2lRJWhPeVdyM98qHueLqRzwHY
nglTXitGoBC1ab+gL4bNGzftsFP00m8U1Qs5BAvWL3bloKWAOb0IowP2QDCWZn2C
PBZRX+bg1Ilyeplr6Cs0aoiu3+uXyjeqOlGqMjoCZWsLCEbgJJsWgVHl+LfP4hvG
J/4HjEht6Z+sObkRJgC2U7mTpnawofEmL8Av7sPzzI+VhBP2BCGVmANQa/IoMoaQ
IZudwheRTuqEhBP8x4c7Bdv5wDyChU9EVKfQFRi1kX+qAHAluJUq0oglIqVIupkA
+0A7Vgt7ZlCgwHZgFYdx4vUo21hEcKoE3O6tglkW4ELemB5EHMqWgd0aFRmsqh7M
bCF3yO94BSFJ21Fexb95FhjvA1XAquNW3h3cEWSTbuTIiOsdY0GW0Tog4HB+l4eo
7Zhf7P+JwXIzCmmiiuZvSQNsuik8MK6K9gX6z/nltXTw7zEJSMGI7S5fN9cNS3Xh
3Zi1K1D9Mm/g1qWrIj41YBjaPbjjuA2NIcBxD7R+TIWsrAYurglwd/oQbdogGTYu
xIEWii1Seqh8vwhQdGNFNYyR5z0QOW5dCfxI6e0u0LONon9uQ1CgbnYYN9q42Fwn
EUOzfs7HCnGM3vwToPLbDxSDdgx7NaLQJPZK7ptykER/ZXjGn+xEGQ5SRP3/VLqu
a+tSajwCiTQouEJSnHa7UDQLQDtoJ+Si6tJQj9YDaHbVIfCYrmCewTgXb8vv74T4
UiFAEBIzCSyRSLI5kMbdprsVvkyY5aDa0bZvy4Y35Tj2dGwIBUu7CJmPkad9pwhH
naQTLiw897CDr1pP71iC55WI5hotttB592ONOxFvyOoQKtL91Ce+ayBhmDOWaSXq
/eXIwjIBjEiwfp/u23f3QUW8OQqJlPCr8kAdk0wAWqBH8E6guyphuA6fdydrRIpC
PFC9kzRP1XIc/RhPP4jM8VJYURHq/QYgQTHKmLWQWlQhfZ09tH3LeFD23pozjVaK
hQjGm6AJQ5A3C0lgIxWWW9UYn7ftDzMAZePxXGrY2+HzcMq0EFz1zzk3/TcFNpln
7twnyb1g7H2DMF51mF2eBrUQDLNHs7vesYE2QoqIXortGJd+MFj+zcenC7xsY18Z
AlalpVPRTo2oPJIEplqQX4akZX+W09iI9D+2cSG3iYDGqB/KuAV7BkKhlf4HxDQX
cKCnUrazXnwozgz5799OlG60UIqROKPa5gk/9UOyL+PIzmmhWssUPpfq/WLp3H1Q
wXW/JTS6h/cV3z+yaftPi+dxIpYQcStjiDf8APeXzf8w5HtDPbHaG8l4ukt1/rAc
iIk4+dGLQBFU3f80v4Tvh0jaZ3CfkuOj6jSc6hCbYc3PePXvCKayyoqDyb3NA7zj
q0wcR632KisHnC3bU37Ir1cxEgOQEZ9I2LReSs4CbD/a0ZG71uP9TM7vc6MQBcfa
3+uGq/kREGkppnMMfaLCncs7Xlfrw0SnVZPWelRdKlaD9OI6JwtRsbbeW5Z7gck9
hQjh4mUA647xeaZRSiPNtot9BR/Qug2Eaz8+Yb4YHZEkTMEwVGPtxkU8dK/85b+a
eazIguvYvUB1hMIKlawzXHe317IzRH42gJO40OxzTNsgHid4SlCOHY5+K0jl0oIk
hK4fJPOHfXSuKFpxzUYHyy8MagpGC49kNl6CQxTv4o8x+TJRgQg+FNAL0QJTJQZa
8/XtUD7NuTzhSfcjZndABac1iWpUDaEvm4iFK2nwXXS40Hk6DsdBl+KMBjVqPaG3
YZxmI+ZJUHDL7Juue0keGkCLfMXvBgtBjI3stWBAH2cvlhgv2U0L47KlK19mCB2C
jZIebtlP5+hJ27I1OMvGFj31QTbv4ip1+TLUDLiiirvMsZ5q8o2t+EemhPD05rwW
SblPZmfp/SFcryQT2aCTZjhomjSfOjMNYp0c/bgIEh+tG+qDi8j6VvVUAi0y/xqF
IgZJbZ0nMXkQRgLi7Y9DJAJLnZTkTwmf6YmMOjRDSC/Qv0dZEWLMIpx0RqG8zybK
WKmCPDi+jy3zIu21+olxQq/4zo62JhZEoqhCpZW5U9BlGjeB8ed5ZZ+3m5N2HwcM
F8xUw4qksZBN3ZyXqWmLj+q3nVpjFqHf0/fz1AshDDk0UQIZULqEeO2f8n4/Hnrp
OkZqfn7l2DYp2NwXOsAvg43SysASrGtZO+3HmDbO8daEJg9Gd5kuyN7YSgYQqDwk
3kYl7AROQ8i2WwRsD4NpWxjUQzt1sCvCE4MAKZ1rOWFzs+sKF4L0MhxQfckOAx3O
gE8drsKW2N9ok81g4b+16RTxkfy4rt0MHI7PFGVpCBJOGrbTa5fhy+g5Wj5DxP5D
P3Np8aSZ/RfxEMBW6eevmC+bLEtbpFX2Z++3olI7HNJWSlTtN7nQhQRL76fyt1Oq
pAr22JzN8CiY9i4ak95Hb0pb5lk7L+wA1D3l5jrd63/DPgkBwrQk+OcKqABiL7II
PD0KE8ROBVTFRFiV7EhKj7vtYWUyNMj+Rk86MRg/7enkuctvYc3uzjY1oNgz1F9l
fOHomTaT66+h17kXgveXD/fglnZcv12oqsAn3iTT3DPL8MaOIfL6bLqxBYdjuxua
zohr3BJmuZQWtsNgpRhtNDv+efKS1YWmn1zZXTH+ArH6YMZlLIe/VMQMNkQrGX7u
B9oR1lN0za65cLqs7an48RQmQJi0xpz/jkCmmiPTrb7KGsqq+2iSdHr0q7576rPm
1o+0kym1KOihdhvQ5c8ORqktVkCHNxvVkyvoO5Z6Fj696A+JbDZY8zuC41oC3omT
qWcgDoFrQmu8yMoAEc2UVRvjVjKjPOkr9TrG4+Ul5lq32N5e5pcq7r13vaX61Zfi
pWJuqkjR3jdet/9HwCN2ec23XjQZSH/PiavXirWb56trKPSBAN6Fra6PYndHCpQh
T8IGLP8RZ4MMDXpJpRK/L1X0DTWdyGYDdYIuX0osHGp/hr/ApuEeqpNMX4v/oYPh
CoK+ZJfsX025v4QdRQkNNIBatvr2kPhDNyludKojexE6QCGja5//M5fvu/0onVhH
qC5sjt16IMuYsunG6kosopENLZV8P3KfANAvNwgEYlbEftWtlMmkvw3luBOO7Bd9
sTVPhv8+erGWnXrAFqgg1V1+NQDPRcRhMj8O9iUZOu2nGRU0LUmO5hitZ2BNREq7
BnRs1hkIc7ZX8nnx0owCSJ5fx1XEuE057gNbFE+glJj4tM+0Vo2xTfO1AAjLQ9KI
ZTqWnVlY8wkKZZvTnbIWHHF2qpczXY4F83LgVgkkAfaZqILtc0BU7eMzJvn8FrUt
GUlBlmQBjxPEv+H1U3V8cafsEVls74Kp2+0qTkY+c87ayFuaewjVxFp6c2YSIoY0
hkkXeMSl1yvIWUcG2PoUvZeeOb+Pof/K9mC1cFmIV20kVvaHtJLXDi/lQjNd7HVV
STzPRbtgr1JeOvjUWrNInfqYs9YsO5IvPhtwAl8nUzMNqi58CUgnV1nPCxmORAlp
NwU/VuAwA6FWRIBqHcsvqGl3HkasjnlmvvW6CPYX6/XWEQPUQPw1ut3Yys69Td/u
MTsEIseqlmUQSrElSVpg6Y6nA71QNK7Jy/WiSI8Odv0XhXbtNT4NXQ4mtO8Cs3qx
lRDkq9QfsQdiYaAEfyPRW8H6rDQpjN89Mlub4GWxhHtVeo1ug92mYob7XEgaJ7cy
s+in6hotzt/GbTUE4A1fGV53gv4cueLGKAMY9+zoGjV1e7zgThJa2UBdJ4IbXAVT
AQpOuRy43AC9IVwF4hzHmUPBAYTUhRnyFOgH4eZV0RGIi2w+a8t8qX+x90ZmuTeK
wcRaNUNFUJZqwjkISQ5FEiPLeDrOs5IGwt7qEgEQq3uxvK4EZvhysWc5sdrkjVYf
gfS+qIdUjiWiiQzcAyaeX+xbLdMSjJAclNu+LmYY22kXKtWtZoqmAejbwygqV8aU
YnajWozGILECTPgkqZSQ2rCTWrTwesTPCGw1bHYhui1hoLFW7g3ENn6ivNvtcwx1
npbeQPd1z386U2XFLC4PLF4loigKp43otQHZHA2Fzr9d8/Ob81eNlzpsbBYLnWjB
5iDodt6SgA7uvrKgSpB6mCuosteWNq3Q9CHv+/aL7aRnW19YgGFDLxj/ZJIjhhVJ
j6CsXkmpMYY9kJvLSGpkxtEbRfZp0BqDEUIvX0++2ioiR2dUvLvmPRg6z10sWVW4
MCMQZlLdyQVMaCUKK7t1+5GxPtfyRFo/DyDjZZ1/1k+UV6FZNghKdJ9dij6vFDZP
2kFCMh2xzRuqH+Pt2B3mvb67ggvfV3C78Jd8ubUCwMN11bymyvca1ZuLn+/uceA6
ACRkyKO0PxuRFFm4VQDTUNbWlk9c5b5HWGSAdaC3GILsLe1j/bELnhH3tOmd2S8L
P6zfLYDa2QLahdKXcDcdlmvqZZQjfkGesDIkR/mfkk5z2gyYEOVXI3ELOhoCf9sx
O+8EY1HME5itKwt4yV+2ZZrjtVY+svSxX88jXj5D77Orb00qV1vz7qHUWrl4fHcD
V2tAwCIDU0Atr3OAKyQCq9eSdznSE4v3kbuKRKX6alrG51YxHwjUr0+6cAkKeMOC
uVUvOH4omFPzZKpM6/ezZesMt8BNkFBVyI1IkklYZ/RlWgAFBIQRg0X0VX0oP93b
xQTC9L8Z6jlKmJzkZLHyoKyodp58lb12ca5JgtSn19iiiVN08sGAGw0XoVEpDc63
K6+oyrD7b7dPWCTY+jK2bxODm+cccoSz8rjHHuqe9zT4+7dy3+D926bz3cXBIplS
GKjwoCy/J0Mefs+dFgJtyonhp6pwtWc/WHTF+YCSIuTAse5c9yl92XJytHvSXQyG
VPtR+XMg/MMgHGi+UzG5YDeomrYVavbOMS1mFnrmacfBoeQ459q2mhH+8yNzWdSK
7HNRFPOS/nd9odJd+g1FX4kQhdL5fYLoq98ZeuWd0v/7TOma0WBjf9sHKVha0tOG
kKtSf9q7IGZtHpkX24RMYMLxHuC9WpCDyQzfivJ3X4lH4HPen10gPu2BkH4obJOd
VrK5kPUwF3SYKysyTcPiMCW1Yfu5FmeL0IN003NND802cvcWt1fyFpuzClObB7zn
QU84ZBpFUW4rmNvXIJJST5MSJ76Si8npA7vHyo+ZtGD/4Qqbrm4d6WTHE6AVEKny
MYj+GdujXXDZb16136G8JHo1vR47MulTG/NURMOa0Kx2GcLn5MGQB60MWTxLCe9q
Ma+X6+Acb7RVhyMSCC+mQSPwUMiOI3ODQRMtHf9dhg/Nx6BtVcMwW/l2tweunWMl
QGmK44ynbaGeyuWsaShzW8jluMWOdJbVeX9fXAvNo7APqCFwKo68bmGsHYy06SOg
mnCroXNt50+eijEmCg6YUSC1APeNbz9fABqF1hIS1aZLVnVvpS4MX4S5haVPIWYY
duK4zoljOXz3HPijKg5Xt1NjmBsBHTivLJc41gH0tSwuZeW7/u7S17gdCC5WDu0S
qfk25dUG8IXIRC9RhiIhfAsCzomYCzto/cwYLy7CeaXsyx82YPsyB3tSh+HPh8l9
kv79p7Hp1Gs3/9W4XB/yvupMWbQT7nfv2I9yzzAHqRu1k96xBBhbbmlH6lcUDDgz
i8Smidd6L0cRXd3P+IVtv9E6jeVcISee9Zg6hMlgu9/iFkoufqcPwwj68jMxzKjx
fkrILCLxF7YJr/NPjqi4wMj7lu252u6TLXuxKKUSfNtlAe1rzaBDOXJ8vOBNK5NI
nNkks7TUIRwfschQn8CrG5GNq8Ue4eY5tYP+3ZyY+33Jf6jwHexJ3q1IO4JVm1D7
7ZBGFXKhDNHthDKUkL4rztMLXj2/ALQwkTuyNIgirUolcHEt86DHPdmkxQ16nvWE
IGE6b3PUoA24bfws6pQw8iW/mlGsGBiqsOKX0iYIlDfnJap12QPvk/QWwCpJVZc6
JTOaS5wnrSTDuZOZnS+OMdpkO0GzduBTTaeVAlXrbZJVIyIxWfMhAxva03Lkf5RD
DZL3Q/8CxGVFtX0pUWbfcWXRekJr29cr0j61Mga1g9K37janz06QFUeDGHOZD1SN
MwTRjpWJ5aX14lCXLJ5rgJzuOC9SxK9OiBJp2o7b7YenOdV9qLUvVayZF51E9QIU
JP/wI/vPmDPtd+9N85zLVy8YuGMvUShP/93AJOfN2SvbhkUOTGGjPE55kfSOW16+
32O0HGh9kCR5E4Uh9HnfO6snIFWS5SfxkFrNztFCDAJJD4Y0sVWqW/wd1r4FDH40
FKn8r9okMtoHPM891mY7PS77evL914g+2+XTzZctbgEnhZqH9xzNHJks9Luh3Y9w
NbUsyvVDofTJwraIvqLiY9n1gXShDEOxkKXWhSdykjlJXOVCO+bl2htL5xMJwzWQ
G5/QjldYFUsmr+NKBGJKmiEn62QHikxZZWtVRd9JlhjLKHpeZTBDUrOfI8axHe3K
8m9A1k/5fJQ1uOo5TfxgeHd2QJunnKq/zGdmXZZaTGytveBmjbgHNsJu++nBdZEA
YBKtkTDRT1M8ToSzt7x42j6DYXbpUZGnS3y3Pcf1UyglzgiYlMbx4c3vhTHnXRVI
pTSig4JUc+QuF5ysOtSENTsgZBDms7DBl6adEP3YS4HVcpsjQJUS7HkMm1xhQ5JB
aODblCRjSoRVxp9IdRLjuU5usjLPyhkHLnevEfFNeBBKkZHNuVwCQ8WWxWjstl9E
QiXSmvzettdwRjo981q4tNfg3t4ZD/oRyvi1pTefarG0xqhQzQ8Sj0M9jyxdFpfc
0fpic3BSkXPBj0jfB4TAU39+DzW26VS++WODFC2Eg/LHGO7gAHYufDUMo16jgOlm
r98bvjpRrbI3Pqd9yBLfnzqh52fqm2Rxqm1+z7tGpaWdRlesle2tHHmOouuP74s3
Ba93+klPBCT0cq9cwbkkqPbofOkXVEsxMeSkAdqA/DUD2LEoKW48CYwWr26QG3js
/INsP8LnuIJ3wFoSSmvUBNT93qFyTJxNJPuJiBAp0atvJy+WDy9RLr2siOKSXmcA
fYloKnr8bZyTaohTu26A2nFHEU73AtZsj7dOnXyk99fxaRbYbLNx+cN54/wY0x3U
S4k0wAnjAUc34MLR6s4x0bc1YDZeYU+zVSoUWdeUOSaSBsIfvfqJwL/RrVtl8yZh
S4+Lrh2+2kwOGG3XmhxLj31HGMcrKbThSE7l3PxDxX/U9aP5R/GtN21qBPxdV6fV
C/5mYH0UFAcegQrftAnSbVzme7FI/odx2EUgk0F+7HlYkhSEOHco7F39ZMUgz+ii
8R8NAwghypqwCUZuUyDWIJhytZQmuA+pdOeXstNR1myqeq6BJyn86dsHK5OP/ct3
BkpniQgCH+MR8J3dB7whXsPzH2p/apjUhBVLyvBT4sBTw4ziiE5gw8XNoQX+ZS8z
PhJ0mRzLbIC8zVgkWI1C+JWSVVYLmWRmJmVfTL21tvOAhUEIiI8gUa4+QgdMx/uf
E0utakI9EJNUzLWJkamTFm3tO4gQwYvikwh1Gwi8lW2FPNdxcbw4wsSFa429UGY7
KA1rDWaDPlljmd4fgNhAUi5+ITzTwmYuoURMV/6bUyj5fmngmPMGc01LwUparVCv
N3q51a+Voc1xMcA7+jJNLK5wcYEheaZLbS7Uj5GpsTGO+VxD0BRWn089Yt6QJytx
mpd2vp3MGYX8xn/EgKI6Y7VpWAF6+ZzjOJ3eu3NITmNcST+uYDBpaH1qJiuMot/p
YCYH5vR+2k06lAs+cIW+GImazqaoLQVCZlnbEcXMT5FSz5UIxq865guurjyYiZSK
cUAvkQnaU7mXWMDsobxrFN7+15hQRnUyCAvvfG0WUu2J8EGaxBEPsW+1eWS2okMa
SNGNjOye00F5RF/2P2TIWYwJ2Gk8vSPb8k0CQQyeqLNJYXNtbZRnlvyGP1fOUxcO
dUY6ry4rtZQasO70XsrDM1ZZGct2Wmeq0HI1Xxc2ZIoxTBUgraVAnu9GgA7/zrv2
QyLoKOSh2Rz+vaeeJOiDp97n1fTj1axlQMkPGBU+T5DT0Tx/T+PQ91ZjfXRbjcmE
+p8RTqPQlifE4BRvCk6X7ZihfrbMA3iBa49hP7EHNc/q4glSmFUOZ2Pv58Z3pZ/F
4O/bcr0UNn7DeNFIq8g2U4pkHOe8HsLXBioQE6BjaBeBiUdM1JQj8Ls9kNBiYs5e
Q1xKQ65kdTdnQ3pO9wiP80MmA0c1UbKWbXQJMJnhm/jrFkkCNddQ6uAcXDsVaGGP
X/Q2i+QaSkHHhEc9LOX1SAl9kJ2AJTZBAM0RyhZ1q7MNd3yb19hjK115OAZYreuU
DgjYvyxh3qe4sh+Qcravlx+9zjQow6X+wwYTbH5aoSR1rTDg1dvicT2BlClXARo4
jbXixpdRBksehjmWUxMlBvZgw89QXN7XoQWvxItntgIfAp1RvffBegl1aLbVuKzv
+gg5TJSvrV1iZugJ0hAKedhDCm1BX6RJnZX+HXvYczurb5Npowg2sqaj7bXHHOoq
bJ1Syqv0hcvfdLkwF9Wvcm68D0EqFM1kAkGr9I0EBFMFOyRnO9v/ZlMbL1Q0Gu4Z
OzDiTdvW+JvLj8NhkmA3Yng6QXuYbnWAYfLcrgDGdqrDwjBAGNec3cuRQP+di3mG
dAVXBenPv93GppUQoewsmUMuJzw5H3JYBmnlH/jr1CaAuFui0cxvPB1lvn6FWZ6w
66pRyPS1wgRtzA4h2y8ZECR2iVx50X6jzbsTg8e8dqeWkwwSmPGIw5EieZD6HusU
fE+CJpSkyUbIdgRhd8E2yw1w/UXnvYvbj55x+OraVozMva8G2EMvQDr7vu2dH1qy
Uf0fodIyQEKwJVW9ClOOUgN98l0L5ASBXtZog6AyJYdGU1mHZj127bb2+imS50F9
xqjqQVYyJJoRljdPrUmQy7KSA140cdUDPVPjxDLCL0FBid2jFvnV8reIMp4ZnWoV
16TqjXltXssrwGexivTOnPxFN0g1cI9sQyZMt9kfCEV6aZ4se34jI8ae7RqKwd4b
uB4QEEC9aVkf6ouwHhf4Aweo+oA/khXuE9Da+sI6/WHQyturXNFtnniaIFZqmBRW
gXxIPGJ/RYMDk/Vrupmgvyl8uGGHvX1a19YLN7YsXN1KbfA9eTcnDvNKEK4uitTO
0BXu2LmMmIcyyECI0N/YT8jhIldV3GiWRsgYkrjSMfdAxxhaH57GsawUVrvL0UJM
AIMBCHvaHgw/pWXnNccrEx6fDLpe7s06YtXQ1+ky9ncg+Lhowy1pB74GZigYNd11
dOoEKKRO/mGK50EQBj7vQG5uDTITeJnGEgXp5v1T2Xns9h6mmorPz8Y6qnMRs+QG
KmnDp9YfYQHY+fQcF/fvQjOD1GMf1HpdV/mjV16WvnfOJnGbKbqoWMhpV9oSZZl0
Gr4prDqZE/0r9fXwYBuJ6dDgV8Oh+vmxDuti4o4p1Ei9EsVXzLHQL4w6wEJJOBcf
m4aHE2UYaqLYrunABt7mWQYFJPm5C/XptYdD/6DYoDS6PqtsItSK7tsVby9VGFWY
WeUtLehMwuqS+b8ZTa5CGIuDU5D9I2QL0QAX7rJoXL3DoVbsG0rla6iTpjE/3fBO
EQDVk8mEnvQzzCNkpv94Hp0799+SYdmR7JofXm+E08rmxNPz8lKPhJSoHFtAbPPq
JvbzYJPIXUX+XxEjCCRqNA28EiatOQ4/dIjMTRwLbxXOUdDf1NYy3NjGbDLFdtG1
DPw7ywBCExlgQW6hW/t1VGT1uIQoLcmx+zlASxBa646I5Tht7I1ZnMz4ALEs37OQ
OxDQfNagIqVfdW1w7PuN773KXCNv/5T4q1MviEbja6Ew98Fn85jzzna9BT2iZ7jY
vDOvobj8mfFu+NJ9htyiS4TNIYmXx7zXHEnuDy0tDUYbrrzKKHlbqKhFyk6nMBVI
pFmVsBUN4CM6HrKJ4mzR5Yc89lkcmFTIVSncO+ALCnFO2Ym6m1FQQsxU+biYe1PW
bVB/p89jTDf79csSRdLlRFopLUrnPzJcOdOj50MnenqLAR8LuikboZkQGhtyFt4w
wV/cUv/7BEkRDF9qSN39PpDeFzCLH+J5guHDVW2bv7M6PeSBVUSUX1c++JLSg0P5
K28a1jybtW5Ig/lavoPUGaGha+YGRp6/9MViab6uuIjysBFl8se4d5oOrz9Qpp6X
/rf49xByM25UOZZD/oNb223IAnB3k5qFCqEevAR6lpnjUnH2dH0B8WW4yUyPdX16
kqKla2fqs8U5fBW7AI/PbAtyDdPMre6WGJJWFFLAm6yuAfhUEiQS+tO4IypPgeVE
y1ZpS94Ul1+i4xpXIjWoBo+dHQpuW4MA9H+O9K6C1ixwd5a0jyxRB71kiSI6VLZq
XeTn0V+0rV/lDLhI50pVom1Y71Z/cZS7jPY0jNt8Cz+U4HFs8AlqTzOrY73qO8za
oPuR60owNB+DpI7booAb/NB2If1RxT7NlbYPOZAxB1tvlaiWLxU4g4TdF8zLn2WT
duhbYD0AgsgljXKt/wva74NJZhIuPISHrpWaWxV0txobFjtDQqq7GC7y2V97wHVY
5FEiQ1AGGKjU7L8/v2o/XOF9cUYiimYjN/YrNxewAVeROlgcrzBUVq9m5maVv4Qp
1aMJ17npXWh+1BfOfQQN7O0aGQJSDf0i/11XlgPMQWoOgrujtMuhdeBz0tz8KL/F
asy5TxK+QCmqvzo2XNIn2u4SRiEX21U1PR8ktYCP6wt/o85x6XKFKwMB+Huz3Cat
K4XR7WyX5hRllLJSYVfnml+yPzVXY8E/6i2miylNn9j4cPQ16p6Pew7Ohk2uiUbC
YodGvhQ+BxV2WxpPwpyQa1mllGqjwoBYUYLVAewMO4Xb2uEufwcUXmco1U8ybj7x
NNaWGDKzh4inpA/4l8aTVRycCDFQcd/rQvd28h4KwENfpnJ8UsIOfGME71aNoHwO
uXE5LgOENjfw+lg8cRtEwzotoIpsubsEvRRjOkd+0X981LoGmIlce1Bt9XzVXJpq
0HH5f9O9IBxackzNOQRA3QJomTOe8B7eqMRpSGZucpShvDZN3CcoSrDAjIlygLWG
dqVxargu7U8Obv9WELoTb9vTjrWYFl9LGy5j+pyABettGXQ/5nizp5UQ3+08jlLR
EhtCpVTwgurotKQYsnL9KmE6IAPa1RaoCsIresRZYTK+4PrH5OWUtNG1Q2PMTCfZ
lfa24oYD5UFpwOxjHupaAXUOhfranY+BS7qavLKpFHTpsbRX4kOodK+1rfl6CDGC
ku7RATr9wj3CKmvF17ehqrls3dS4SDZc856htFr5SFHK9J4xcccZsFMO2fej1O8i
OYX34IVm6lMkcNA02VjGKuxuUGs6nmX1anM+naJF2GbKxOsMuGUfzFnezjS4S0fD
9VtvPlWu3AfCYnsYzuKOInGzLBy0K/63+2thngREjPP3pet4EjO2wfj1QrzWMVr/
bua4lxPxabjT6napw62OV2nfp7qUJF5Kqh5wrx5Ua7ze7tI2/0bRI2yxLGTqeUUy
c2jlfNhzT2AjuRoyKrqv8zEfNiwn8/Ep48IvEvV7Tjsi9KZp5xgMeRUfiFxQKEOR
ogYkDDLCwLEoG/UHn3KZxH7wwqfBfLbVBoYsJdb0zY2S6UXTKQ+HXXXjOa6UVl6Q
ayfIqmN1OLDYKyhJ5TOnkfltVMtEss88NvWa+C5EF8sNvyG2QMOagclxeW1UbE+l
64zBasWnGNFoFbJKeahzJ8yXFPSfwAs2r3ZTBCypnbNbWsMOjESvkMmldMovIjnX
PB+EJBLuTTO9+kv3htrE0FMvpQCurX7U0qb5YTzhiriXRKvRe1Dl2Gu+XSAlhMb8
q9JtXo7aFfLER0s7Qdv+fwQa+yf7dfJPJFhtucJsWr7ckNEYx+KykX5ZjmA0AmP2
U0F68nOBmCCridRaliVLfKzV+h5g9jPtRgInGAyzxVXu6uShqwB5gqURwf+QCGJc
ImUyvUsybWgILW4QU5epIQpmWOuGwf6XwcVRrSf/Wc4Qk/hxxTstM7hFB0fEx+rL
bDkTYhJsApOVAqxeICr1Vb5ZJbIdFdi3fh5VO7o/X2R6IVsXHyrxdRd3i7Nf4MAt
Adb46oh+L3lP60pwLGuEoUzAulCZ27BIZ/7BCWIZ4573vR5WAezO8TLigGzgxfag
558CezImXKsPl7GyMRHRYz43F7GKEjbX3S3UL6eEOn5SbKcgdS7+Ui+2AK1sCPdh
zxZoWnn3LBspgpC/NObn9CmYwvU4Q7SmH3lO0IArk8uoAvIkxl43YL91d0CVBrYB
xsmNJQsXGjGJBjV5YlUz1YPsBXEllEkteH5pUf4sJJND214LAdE9qcXIVJrwROJb
/Bj5M5cXasMhI3/DYIR1iBCRE0LQJ/vuqiQ9OakkL92hQPmhJLrYbXM78bQr3o0J
KL29SR4ULDPoHaRHhe3hadivY1Q0cUNjzLMeUFHwNpKCBtT9/mXAphyzxWZv/jDF
4rHt1V+VGOsu+tP59RdgAS83b1XBjVbfGytQCHar/WRZLLdnTRE1H0tMZwr5nR26
+/wp80LPiYEzjSAM8NWSFrz1BHn9wSY8k50Y71dgsFv5BHQNAvcU9J/+w19W0D0g
g1/8FOlYy7QgKLmjMOorOWdmSL9/4WOa/4uWus6qClHFEg/2VbnQ0iMfXAydpvOw
KI5/Xum4+wAguvO+/E5ytoOSke7me+kqwNHoCUU8JQH4Ff9TmAPPG5QUnHNgLq1a
45xh1cfFH6dSLX/GxvKY6pwgjjtRwf18HL2sdi60/2hxh6ion0QPBu2a7hRelY98
kW7w1zFo10nZTnYYupBs4i5k5CXoawFQQR4ccfp3uCacHoto0vUKK0z/hsGZwPIT
SJMHaIl9kOWqWwXwqVGS5yQp8hqnCGMPGjUwJlE7bZlmRWF+X0Dhi75n6j+pLjt8
Ir42tcs7rEfCUxOGj0jH+C1FFzwtNstYgTwzbx5efR5kGGB8E9E92yjwukhS+m6E
bAdDUeD5LxiKX0VnflHNLOEI2BIeSorAvUBIyPkPVE5Rt/QqkZNiqs3eWpa/RrTB
DYhZL86ByCcGjtck3LhhbOvzNrkWNkXLyPrp11/H/+LkTPavL/gt7B1JBDkEpTEe
TopClgpG/E2Bz7lwI0KnY1YLZpQK2t/4xcnVIrYRftbkESzABbf1+zQ8vONzTivY
KFqtlijcOdw6eGTwLgk97+idJXEFuV7ox/OV9AYEKC/f32ZsN10u/ZSPL2MSa2ha
huYyvNWvQMUEW+V7Kz1sJtCPVrH++79jci2COJThCxUapQ0Fij1QZhNUisgzQskU
41AjBgue/oC9nDledRG8WrQIjLjv9zdQ1q3m4IdV/Oo14P8rkGNPZxbi38KpKSML
cVLxjzZZWOnjt7nJABjcesYY4MU22/U6ZUsKAewfE90Wa56jBEtDnsylmKIA+Ah/
w+wX26sgmFJt0fnFg3JnmVkJWOdSOJdZj5WyLJWoOqZvGcVNJdj+S9yRvn2sva81
IflsSMW1phjWvnSGOdGr2A9Din+oGz66B8Bkdmh811AtBD2FuGWD925yL1i6/zwB
rCtrRI2oyAB7GIlEsZJdxqK3W/JbEejXJCzWrUWOTI070mBBtqiydX99uhU3DAnY
MQY2/MdrnU9sJFjZb5bwrgBk4FP8WGC9rjkaLg7QqPHPdx59XdcSSgN04fRkLB41
lhPOBwtGuGWddttx0pago9ECuggINdHSvLWXkOOWdAj6pe3EvV1r7924gLwZ9Qnp
QVQzBOEBYfGagOF0VGzlE4pyKhWl6BpRZMIrqzWYG6AbPFQpI2MUuvh+6jLMDH8J
0wbToBTtqsZ0OnpBQPUdBJeGmhLkmaDtENMY2z/lXHoBhkNYOUTsRzibyQPFubsl
oPLSkTU9e3MffL4zeqlqVIWbzoTkDTRujX8+q7m3bi2Ygp60108Q7WQrsLBMn8os
kpp826BsPDJPSOUYVP3zBqPAvhR/dMEsY5JnG5KU5p89ostDjQRe4CJYi7UfR06d
FUDA3Jn1GWwfmRCfAbkZ4fRNa7lYqQavdMLw5PK1ftzJdqvs6bnHtDOrGv716yd4
A4az8ElrDxfOMMFvRDsIQIwdD1omrVzAjms2bFIqW3ukFWZUHVcpbq1QB5FoIJy1
nfBJX0ZSK0sycMepaygXuXgTlfccKbwE1pWL4oTJSVslCUQt9noDcDE/1KqmlmOx
pkbXCq3ZfU/nk8x7MxTOu/zmxBLmiWNDDVa3B1zPh/uKK8VyHoOp2/PX2Q5OshM6
ByzvEuH44NiUiKRpj0nL0kfLLFfYEJu5Lnvo3iHMWlO78duPX98PuaGILwN2Ci5J
QE5I7bvaLH94s83bS3k5ci6I1Y5sz6Apg1ItBMapCot28tL2v8kvZeyse35GEver
FyUI16L64peI3Qo5O/OfBE18SLQsoWtllCSCjf8hxsQxD52whkQLNbdLVLe/xqqW
K2Xii/rrrLZi6pl7Wl1y3nMogbsX1ZJ6+XdFpn6bRiYs8EUgAiAGZHOHvvwsZxMU
j9UiyCia5TSqt8EdeR/3fvh2cRAq65g+J9VqcsLGR32vHt9FXCoX4U2klRyFRymB
GWksaKYzYTnfkJNATvmRpwylGRZv3BZ7uFVcSNm+4ck6LGay6b7qFhkSxQcG4VPL
IvNn61+JuKd87pmqJqind79P2bkCg7ihJzTcSbVj5p0uBLuGGzA6WfYVsBSdybOh
hIRtvAFWgdafsly7evNOt66eC3sNCww1AJNLcJEVDgzrb/sBOZ6yWc3zgEhOevjr
5qYsCrIAzNkcMU+3zw38efz5EZeqFnecaKb9DtgCeVmnRMixG9DiZscoB5K1J+jR
iQWF5y3naOguR5rCjGK4WEvKeyV2UAn5hDKJsULOY3vsi4OLH6ICQwSH7SKy4D7c
6lS82Oac2hVwqN9ICcQkaEeZZm9VCS6LZFhj2Tr5ymC9PJkF0cMO0eYA8Gb06KPz
qn7xLUWBUNIGyxC3WkKquBxlIG80+romor+6JA29TJvtavuBquEtZF3JuMfvtkwr
89PYk/0fmflBF/yfW2gDmbV+paHR7eXgQ6h+V9pLLlIUHaWlW5YTLGvmxESdeeEi
6dG50zI0EKZS4PrXX68hvWUOT2lNCkKdCaVQPgVYRnqFL9VgNZrAM7Ap/1XnvRSu
HQgWR5hNNLMZDcziNj8aliVtdbWa9eaSTAQ8czDnKjvGRxXHqj51bNZbv5gn2Kbo
yilBeb6EjXcUB8IzHJ9vsvNX/OLKaZ5YHyWVDSq/aqJRU0btDLrEORKJhKZ30b/k
9bfNUvG71+o2vZz+b9phCuOHS0JTJ+tHLQ94MgQyvq6FpIyeHndgWpvatwxqcST0
hmKCGxff2aeVQxRsTGGzlPq95lYK85DGeJUHLdTwX3pBV/3jP0wTEyYvUYf0GoKk
1gxa9fFa2Gah1L0G3LFbqwo51piHji8tK571PR40yf+yZH+7J+ru/uyX5pD74HBi
oDf8+er7g9Z1aEOFhSbph/YWrDZGfvZpd0jl2iTQTJn0YDteMGiKDWz2K/SzOGrz
DCsnuj6+vbBjU5YiYkZ0HA+CDzbNtPAugcnQ1OMQwEGrSJccWIviBDPIXFDxYFqD
D4wbViwK6QDSfPLgWTc9PNFlYA9WjePouo5J/kVuLEEbGavn97vaSAILZHBl665+
XEH08+0SLSXjZT7dN0vxQ7syRDZTT7pLuu/VH6m3sm1zA+tZSQxDKs2Lled4tBNF
rkl/EjWobR9g+WeYUVe3T8dxBLmEPE5lTjir9ysVfwg72ZEowKT4E5JrtoTDwDGL
BX4E4V90INWOSKU5XeJgbbIr1MmLTJie6UqPlvPW8FIwc0jAWocZFhufQtiNHpvD
+fDPsS0BVc4yOrnAg3a7Vfr9TShJL9gXGLAzacOvOXPH9cJwIz7pTt9HppYIQboj
WpejBCajHCS3VCGVQgKKaDt1DM6kccnCzZD2WEtSPRIrQlWBn0MeSWIpigrxRU9y
8/fEbSv2Trq+JbjH7oxlVC7RG9BAqjUbzpWKMyXxvpLL04R7z0qRwWbO+AGQa8y+
0EGpEfD19+kfdw9gwelrOZEGiyknAh2cyrUtDPGmyOhY8+pLFjafdVSAjeSRNUbU
q/+WjtDisdWa6hyEtwPbkgT7/ln0G4a3R01zNqkCTrxDv+1nJDNIYQYFrc0+LKD+
mlyDJxdgmBUEkzi2rE19dwd37gcFBWRn9kA4BatJJQyREr1YduFgFzv4dflqz/Dv
OiT6l8KSe9iCxPqLeeEop4ok/w0a2ahqC1CTNDH7nDzAcH3v4B4STLMyjgEjWejt
fEuuRShxJJq5KuTM5tBM6j+AFSOXT/r8LbqMuK2YtPEBIkR/8AfpH2qejc9ANaCM
tsOplkcgB+TQbVLhci7oyWxvM5GtNg83LLgUf6etRJNDgmcoFFC5WnJkgBgAxh1q
mG31ernD+CpK1E6CsS++IqCosqInh9X01+Rk0V6xX5FAhxpJfr9uoaBPJMDlJcA+
lPz1NHp3hv3NLKRXgoWgBS3IsMZyGf5k9Sps0bDY1uTycsCoOeDiBd7RpJL5pKkE
nvIL3t+lidjPhL/20GpRfDU/vtQZ2jh8dRIx+cPaHfOEhRFPcSgBvXXfgrdcED+A
a21I/vZ3K8doelkFjFeJj7udf/Etz2Y3u6tHNkvhFsVCRBFJpK0+5oTLmKaiG6Yr
7OIGuNVUXAgYrqMrW7mSeK8NqWUpvSsZFXNMRmkjoVGNdg7fPnkyIilAOyKJwYmO
o35c3zp00kCF0qRkYx7r6M2wANeFM4t3LH4b2yL5cuPgwuuWANG2A76sCZf1AgfP
12WIMWV2wJdyCLCjlzZUImHgxZ6Yzbq8anhunEjuhi49D2dYzB/2ilhVCnkLOOnK
YyHjOAtSDduzcygdwaTnsF+YZbpXbTKENKIvhexBKwmTbxHSAtPoXMTBLJOL0BvX
i0qmE1aFEFJMFbLPuifZN6jo/yLkVv05Qyjklg8gGcOG93QI1G4F9RZgJyjRQOzu
xRBDxjcrbX7hzyZB3uR5bxhH024YumYGXEXf88rkmAoUhG1M81KzA9fIcl1JaiNy
Neh8XQIzAomwAQcZE8p98gCu47VAavAJzwI1c6clk7bYuN7C13bkpoHuTm59tG51
2pg4xXIlFbzxJIDi0IiPj92yUUmHyVl6sjQZjTcPxjXiiSXzYnjB2ltqzwn6e/g8
0OlbYuyHAZ5qmceCYlFrzTDk8XLocVgtPDkCupUKZ4Ps56vpeFwKw7vi92Ffzce0
dfQbvcp8P6yK+OoYcqp1eqdB3oDi38TUumK3pLo7aWc9qnFNWD8T/Q9R+Z4LNCkZ
fza/Qsq6rNuNmWyvTkQl8LgfpJxiWk3dI0tz4Nozj/bzE7g0IsF12x1+0xenIByl
3bNMhxYtaVoDagHUPWLCbB917sC+fD7Q6p6IemBfTwVZ3ugtw3Nu5l97AMHvO+yQ
1JBhanYl9J4+pENz4EgxAESGRorh/yBrfZ/a1t3Ewi77gcJecBxVQ00Mmfnvsc5Y
MMwXh1PTDQxX2uKRvCYtd06dmjZ18SfaWvTnC0xapyUNbWJOkWKcav1HiyWoFMtC
x4Aph7OWlHu3/w1NSNlsWZrU5e5sP1q/um64mpUR3JdvgVM2GeyHZJeekm42ZR1Q
qxhXJWk4rNiASqd9h6+Uo0Z2QZVhH9x+tpeWJhrRLZMwuLU1A2weMwLEOUFL/XAX
PyjTe28pg4z/b2ErPy1gk4NEebd7Jusyg4UAv70RV9v8v2HsSURSRkT1hBHr1THO
PAU0nzTQ8gpGRrYZfh0DLC0kTpr6ucb9e3zx8JUetWMXq6VEvawpE68sgb0L0DnT
l0v11MDqH/XB7/NdGMktc9S0vv3XAwrpm6GdZ+o4GDbknNWF8/xBgIyBSmRaAC9r
LDa/me9D93WzWLXq4oXmdWQKJtgLij74Cx3tSNOJLUooR4NQ4Vq8g6vBYN0yEBz6
SeqD8r1Tg5TMdMAW1vzEkQZlx2ORn9I+0OMuIyIXb3KgBrcnhjpK2YlfQLBqxWOO
9TgcRE7d4J+4lgjplNRku0EBJCKgjOkueTsH5hfoNTKUQ5tjz0CKdRPW9FxRQLcy
o/42EIWA3ANKVle/nrCo56K393KIpMD+BzsKjTK9zg/LCEW5xsvonQQTj8Im4jlh
e45Sc2m9trb2+KCv6cPy/QvKD5xcSpIMf81yFrLl6FKd+VEMkbkJPiRlat2q5T28
9RTwS8eM9f5IhDuMJtzrbW2zr5h0JQIfpohTiCJM9fGGtnhd7kNe7+tXgEatClTH
NVdY1amfBBi8N9CI8u+cK7a90JDMe4rNyWhuQzQ+ESM8OkKTkqJm4u4ktR5tE1Nk
8CbygTO2F89/yR40fz32QKHboHRXGODitbutlsvn4FhnlwUwrTIhfO9nmcr+XlIy
QIC+FVmOlg3YBD/Vz+vQDhJanYjhFM3DPNY0dAV15wNuZv51tvj2gMYh3kvZQSQ9
eKrZlVh5tgxitURN5mLcyHTLSokzWdpFMq9adli/g2CKYzpGQwos7ZwbPBxH9hHg
drmubwbi+8i+Jf4qMSNPDl0JtglotcApHKGSMZDtF2qXSP2f7c7N1SQ1NkSjcAbV
kXj2rFsQFjwdSyH7AQWoQhuhUJZ5i9SNiFfr9fbnomyoT/03VNLL45E92A4svxwR
XTojdus6I1mFTM+HUldukI8XEPF6XdDZOKSYytiwlOCaTrqTudRcGkazuUx0zkju
AV2CAcbXx4yApCGfukSfAJlUNcLG00WO7PqdUiyv7+SNfnIB4suI3g1wClNwxQEy
Xl1l7DW/6SsKlQilQW1EPRqPzxwocEbajMs+PbkwISxrrTlj2YruSR/MIcs+95rs
oTAKcxxwqRu5CZx8xZ9gyYipnTiZIw+x3OXgEfhCMvUKBVrO/ywpJYzVbw3OzllD
P1LnA2Ox0ce1Jl3cQTKbWvKdpX52MPNskD2F4Tjxkyck3mBA74/lOYcVFl6Y/D6N
iFLP5DgOMXofUEezKejo/Nc1k4f3CrxYVV8bDHCzrHKAd8PjuYDOvpjnCeMb1yyV
rgIE2az7x+xPvb1QklkD2PDKrGc8wVG2WZ8Yps8IzxtBSddRZQEb7GGpP+J76/2I
bOLzUGvt9JmlZcCGse1dYUT4oK9GCDJRVrdQNfSWHQoSrIHBJRTXZqjia2Jh727X
z3JQRo565asRyLiF+fQCF3H8Ae9oJMwGhrOGtnNXYbzbQOVl+A3C8PxrdI1UE8dW
R+sO8UuKoIfAWlEx3ynYZZJIfSpddpLANDd7V5ByxpNbBGE9UlJLNS46irduLroe
wVxmmcPcMDxV6pv8/ZExREt0CdRASoYAt9JfF+2Rsj1OkNXfascwHWlEj/mMotPK
5mj1iWwtK9y2XQJhR3LQxQKmtl46jmpJC7s3HQOwTYE/42/XChNJz2rrg+KQjmTE
p8tonvotlzNBE4dw08VDsWtAk5JH2QG0De+CxHMaR70C/s9KoKxnM2v6xxAWIakb
4TnfJZYOKNKY8vqSgnU0Fixh7kMJ9fwThAI/pIOI25X5ZPiFghyy0p9w836zd5iE
6OGXQA6hANdZ9/RtNiDYHjgkt8rsi3W+LQktJbIMAZMBV12WxbipcwxNh7Cl584P
b3DtmL+qPC5KBXbTaQZJvX4ntflG7O9uhIaHQ0PRsDjyRBMG4j8/ZU1PNHj/O9Tm
y+/uPdbXgmEjlHswkToEpcq9ErRBajbRfzUa8LjLXR8K/+FEiCMfjsmqkT9lJ2Bh
NXm0IkbfDHUCLOX4jfTl1s8f2FJ7dmh/LOIiXrwu0nUKGikFVWkGPJhdTMPtVW8L
AGUHsklOJFpj6NLaq4vgN5dyQhd3lfFKb87PpvLAjWTcyCfqV1iRiiASvLH6fv/a
2hFsNyEhCjAw5IRPvy7J7uFQq+vxRawor2A4OuCyv4W1t/AEjxS/oUme4KRphB5x
ZR1TWJVI3NN5g0dZBTxN8v1y3V3hI0+WmZeKE1OhtIMruCuMpAEK5uNtOyqBbje3
bjQXqvs2g5gV6PGXXOYljC4R2LLHF1BXk5zQ6hCBzWbvI4SPCJJYOuHP+BCp9ox9
MUAnK8wW7CPpZVBORgQGjP1bb1To5c/ISqbI8BD8M51csUhxfs9NraGHbCEhtfy4
+7ta2ee0VyRD5tT9RJUZsgnpALB/yH+Pz+ZU2SDzOYQCAqVoIjYQRf6OaWFnOVDB
19GLXMD8VSk2Fyn09FT7HLudaIuYOEd6+QM80pSauOmk3PZSXqoBkjaud59IAMyh
9y/pM+53NCtUkk55xTf0vvBuiBJCQMk955WfHIxYxj/5og9ehGhYfSzZr+A4fKdL
cKaSwuZ0GDT/zmbvsbPmga7BUZe1Y/Ecs8djRuJ7cU33zcijpXSPBBFIuCFz4E66
0tsbSkv6i3hU4ABRt2zDQ2YjPAG8dQpTgy9KQXL+9aMfvxNSUO3zTLzdlWoy1HYn
wuqaao7yPADvrtwnUqR7Zjs0T6qtLJdcvs5/WA1aJ0ro78joMiDvNEf1vN93daPQ
0v2wS2FtEtf1J9ZNtC2y12XCmh5BxJevXmwncvEmLKKTn5gW6cZVCo8qF2kjePyz
oUp5Hgsj7NXLOssjCg5Yl+YB9OgUiv4mVisuweVw9ko93hTN+LXBkPT0NBt1jWPi
PgJfb4QTPLwq3le14ktczdFKVwYOqexmtc81QXlzh8eSokV+FH3HrDmfXCdgHsK6
U6bj81HQFS75+8SRbDCftssftyXLvR6Px680geS40GfQqiGI+UTQug4N/LxbfODO
/RJqdZ3+ggtbifyCLd4nrzlBFRv1VOS8M9JhsoVTNIyQgfl8WxcRh1jhqmf52oYb
L6+yXdID9dPiK6jdSF9cVz73VdBOLJlkVSvRpfCLEMjY0teJOtnxfpVlvg2mzP1y
gd40VFZtW6TgdxPMF84chB8Dx4w5bDQYw4TwRHmykAETdg6O/Z5EY/2o4Ju06Jvo
NaFx1o/hsxAAeg0wTTArakVJUqVgS9PeKUhxvbrOsA8quD4Mq6U+6eypbHYleM8t
uLB1dYKlpBlnF05KmRfSg5Xk+1QbhPmizvIH9SHjhAyN2rWKCkA0dYqrToUslYVN
jeQYF0GP/g5OI6JATrFHTkM9U2rttGdK2jPrCtbDiUjZG859/LDCLoW9y4cgY6TY
vIxfCeFuHLyF6xn/We64Q0tND0guRDQYLdmAERZRbZXOsh+M9EihL50QfysY02zI
er7hlb5mL96ngyxHCCVfbZm1mwVbwF5Moc6gf3PV/N4BVWFAYroaNaEkbwIF+wYX
D0YreTZRoSL+v5VIri2F1SOljiwtWGKpRLqHPddO3/eESTHB8+HSfxptQ615eCdW
WRuat4FTsPIjq3Kiz3upPAbn9UZj1i+8xq8oL7nQLeMsg0onvptU6/2u110WGxku
XmwyR8W2J62I8t/WE0l+3ijJgb58+NyiEP7bxOnSD3ScUHKmDZZEnL5d77kyRh09
yMow2IIigNZeXmPCzM6cDOJsgoRvY4IT3mTcsMaHUwyOoSAtLrIDv8Z4geCL2R/a
KxtcHfjp8vo95zSMV26R2RlvPLl8A+fp5rse/5hOYXlV4nM9CtP0HzQi1gSn28qs
YABAurYHZlPrrmgEY1bjSZcNm1w0rlXdm+tsH2tIvxyGOLLfxZzcUd8Fl4eeI0un
sROaCrLMOPSTZEOxeNcU5f4JgUZwqbq6JECMbbRw/r0g0nDqmJAnUuFKdzCzJJPO
uuMWFl4REW0aemef6spgGbUVRxxOyyhuNnKrslFEHKsbz12/yTDsGdh+mtm6BDAd
imYPEwVDR27Ufbzi3agtQGaNYfYE7EOUk0aAWE73ZJOR/FufCmQMMQCVSbCGQvo9
tvkSNCvV1y4oYlsYDn9UUDbGcV5+4YzTzMW943eoihYsB1gqHuJph2Nb5cyJrUnD
qMLDhNiC8FAzSLWMSLZB0b5E+EKioZ4QMlmaPuhoPAUeeMlNgcIWpYre1qihfSJ1
jIjQWfcOmVXAE2x4duij4dLm2/gG+lUrF3yby05yqZpVUNkPKpmf9utsddxpw5k7
vqNEu4Kfp8/j4bowTKlqQ5z7FprHAsNmO6VABPYQQwcFvv2EslbSOTTN4MPCMl6Q
xX9GlF3ryrtyQokTgQLcXAMgwSzingM0bc51wzTDy4T6cecaF5JNa+CeE5ZS0iCU
DaVhvUgjLYeeYAt8gCdaVZn7MwY6QJTJyr9NnREjqVn9PWvtNJVWKWr1yV4XszY8
lsq0uWq7CnwayCdOLx1sxY26bQexNoZ6X1RkRzdyaD3e3iFWOezBR811zJnUUGfd
tJQWwO1vgvnCwnoKdrpuWjcbbXQXkWaByjsarkI7FTaI393hoKjz1BQU8tlqZcJo
j81CeeStp9PXccoEO/W407YMWvxc7bW5ulw7aRlg+w9KZ5mchjLJKMiC0PtPapwZ
LUERd/JlvBdZI3nZqyj4w+9GyRnjQBF5zTjShWXqwgsJ8bkBw1Ts57Nv/6t65b/l
1yjZaYCRkX915A37RWul0xZIWaDY1sTTK2xksChsSOV3eIT+WG3p5zl7H71JPTo+
j4QS4YSBIczrp1DLy7/itZtdCwFG+ufYq4phyYs7Zubk1ol17mTMJ+UA2LYs2Gb/
lVHCMSzEI8mMq8ehYroS2fnpOQZhGHatdL+NZyLEwUtZ8jfjzTegvLzqxJn1xJHd
MBGHub+TCvI2kt96Bz0gqjEMzhZ2GkHl7hMpFDmSXDnlL3IXUS3GAoaBRTX73MOz
f8k8n8lkosKMxHYfdYgSbjKu4Ix2AK+ykiYqC4frD1V7qISKGyXkisKghB0sm4/O
upSM5kfNAtZDb7noppttE7zU7RBr/z4/C3E2raRhGkvzsnkJcXahM8SsWM9JDC8F
hj4Ki9tLO4oSwI6RHLuuF9fGzycC6zWDYBMMgDkchg7n4/RnQfdcwZQPFjJ+m1gx
MpmrEsCblboEzVdRn8lXcWOgD7BuOUEWK++07Y7AFGndFLf1RTahSQiPpbdL06XT
Q8ITOGn8XoX6TFnV42cK1AKThb0iUgdcJltd4vvuXdaPPZoWZCKNj/wkkF2cPBEn
DtmJt94Rih/i+lyJ0SqyXgqfJmXsS4iX92AuaMgyS6rsjrNopCKosQvvI8zKHQi8
X3lXg7BDabEYaxUT5GdAc3ctH9MXyNiw6WWXx5DxVo2qLCmnpDQYBUTnaiRQZugz
C+VhTPj4OnAur8ADb6Wb3OxQc/T8ZJ9jgPnDM2OC6ZLSq7iKGSbdguox9gQNNOHe
I7M7jKEDJVoxg4QnBYxZbJx7ITWT7d5miEcnQ9QA/oH244/c2zrays1g4rhxcYN/
NF9Bw5AtMepAvtv9TavlpUude/sqZd0KVEmWWRQAddmRNlJKo2IoZaBWcYqxdHeE
fX+yPqv9vxUI+0/XdWAFJwubIsQZm7M94oYCaXwYJJ9x6Lai5A9DldZmo+3Ni6Ds
VyjWPKX0hDXxIcvjMfaq0lt6OI7y1MBi8L2DXLAb5JNJxfm5BmWOUoz1fJmF1Fk5
7xscTieXWpIdzXIj3l5ydU0mP1Dtqrd0INOCYiA++XGkyIsNWOdb8fCWbx1NYkfE
kseAvIcJ7T3XDPkB2KtGJ04MPwD0OBf7RI0lS2MtiiU6lbfQoGpskzy4FTaly1Us
Xjz1fPt5puFNUOujHVHS+CzXtmbN+0jlEgrLyG3ECS58Nohi/YLbhFTaZkaQkofL
tFxMo8UInVz3hoIVnZVUGj1A6uu/SJiTBJHYVCPuo4RQJCbhamNUXjfv53Z49RbQ
K+LtqiElHtr8r1Qs/1JngwWAE3ERFcTKtQaJ33AQpzvU0I4xBjXLN2odLG3WEMl0
BHthQPp7oy1swdz8H0dySj+Gfe4mAPnxzggi0vOmIpbqs9OuJhBIsYQRwgKSaRrP
M7TGPdRhHOyywNvak+rPuCm7apdVhWmTkVzYt0d9AxlKaS4aIH7rR0pE8ZqecqiF
VMreLuSxYJ+kNdRLLLzltAXeUjf1AGZoDO2YiBvkbMEmZZKNmIPTUkaDcTRPwo3T
UXXTdKd2Jb3VVwtcstFt1/qIHKIAif8tFGA8nOAThfp4oxYgZyReu5xJST7HrRjd
3OTKcqliVXzwLx8SNge6Gt396IpehBYItINcjq+z7VS4uM0CRABeaHY588w0IUSP
aaRWc+XLfUKwUo8ZqxMIi/u9zGiti5/xzvuOshpDitrcuAptcSeDE3eunSDKSW2d
h0jmfvZ61/CmtaCszHCE9PWIAMgvpVbJhQWJCBP3vZxNUwOJCjZe6mzaOmnYD9GD
zSadyDSBoEmWeQVnqfApK4CNhtiT35EZmJTu4wOC+x5Z1fKanFjfPqtAFpPtwT6H
rvk86KALqYRnelBS+Wc/idUS1WICPMMDEalAjcHTdRnNQMMhPusKpDwDTBoqyaVT
67ajIWdBVps551rb410/Nokyp3LRhu1RKU/odMkgc2tzpcUWB4FDZW9AiuGRh98B
HwBod+ZJjq4WwMsLprd2Sg9Q1sOt2vYB8r34Ze/NF6Vs0y3d10l96hWyj03hvJ6F
4oSNuI5a8pRw+szUYZFZqI/PmKJuHKkrGtnJYZsdMd7JbEcb2lSMF+76IOtMTEHR
nUooTjrqhoy/NH1Ki5dYxKC1ffhMPQUKjyt3GuZcLQmnLslmVTztPQFFPZs0glko
UpHO6jZqTbuE1ojSxphLtLA7zhr6r3Hnsbd1AubyKagnQS7/Nyzo9dJynTf5oJnu
gLGGidXSsNlGEOPh9w6SNR4Iex0NMsGXYLvgMxkQPdPK4MHDrciCtLeT7CSkTACB
vVlpZzMqxC25HruT5Zu4uuAgu44ewCq5bvojmzhwWGlyOZb9GiE9mly4oKtSvX6n
Ly1vvWeSzdHcN8Y/yGSvpeMjodmZlHrRWB7InIOXzFMLb551wW46u2liLkgP9YtA
hDqTkpW99z8y/fm5xIaiA/fFDVmQQhI2uPn6iVbnxwmBO5bNvF28IhIfbsyi86F/
vwnTUCX7U75W7G9BvjEfbIEuK6yOwi01JszgW/EVchYIt6LaQCV3/n6lDo2gyUh9
Gnb6bEZcmCPbozP0EfKO58VKdUA+IgFTekpdp39GtZJHJYHkC2UixAAPuuxyOL2v
WUsgLx2SCR7dAy59T42DYpYv8cRj8fDvQwUr5B63Og3TKRV4ArLPwrJeFle8cQvU
4JnjcLi+HKgNQbbatdPuNm0z8Q3doAJ0ib9fpHRytb+7OpMZvauMz5LpPaCQ1vQu
Ft+JzebjMdtbMa1zvhj33OFPJ83iH4xNw4os6/2zM2Bm9oj9Wxbu6uZI3tJss5dz
5UPh+M4B3OpOBcgtbay1eNi3x6mdIxIyavsXcleJHBAS5ZTfUEjScoiVQVi8EjPT
RMyzF5ey6eAFwmdziYZHZVbQoCIpoLbkZ9B8NGmbxczAFNUADPIubzMFvIjwfQwx
h4mqNUNG+Fq72FIk4CMSHpa38N/lxs6zZi5TxL7R5Go8oM+Sk0dpXzfUWbMRu4qo
hlT9rU89skAUiBApaG94znCbogVG+5Y/q6C/hPJVLaIn/hgFy009oWXfAlBzlzjH
gYdU3F7bxHBmQjeGdSZ0D0mCRCqBu+HVDkdTCFWPXR87/ywGDwnHDZV8tVa1IzWL
d0ylDTg0ryLixDafFAMmN6zI2rNhhJlv5ZOgv1uz6gt6E2DlKIfajjrQq0qyYoTY
Hl6eYUCCX9mj8Qu2gfcyxJDi3wLsjhxIHL9nQlEA04drrCQqy3l5K4NK2+shXlMd
FUMKJlr16ldoiOG5ARBfzW++m+AkvNXVC8hUAmaF/7QGsuICaW2kxgE73hgKnGSx
whkhMY8X8qhylL6rh6F8Wx2BFdBKLJVbQyiEMAO1CoJGDfzUq8MJUN4GoRGf87ni
322nWMHFeGe3FxEB/Or1P5+9p1SWZgvswPLGQUY/MG22CretlBGT154zIE5OLq9q
iwVgUBo+hsMqPLH/S93ZuqF1Q4mwvcP93K4y7oJNRF6+ZBnnczUxZiy//zx/MXZn
ykSunp/DANnvFk4EzTRZzFvUpJ2d0uE4DUQh2TrqlW8UXlMqCn5r9od8oCzboMi0
DZBE7n1YE+ts/hKq5+fjdNqNEJOSS/u1STEtZNMef83LkfYVkheZLjxenbSwf0Q5
1xA0uGxaazcER7FPrsTGO87UuGrN+5mQx7dHNWtMKnAWaoekvmxX58oyX+JPTjZf
R6eKGerUjdV8GlOdN9ujTvgROlc4e2LkxPkfrjTseDTMzXiTG9cd+Xh8cS791jUV
4bnwbnP6IoZngyoDJ6+NN3Ae1ohFK0XZmq9Ju6keu/gXDFNYF7DEdqgXl2TmmH76
tYCLuEW/aNIOfqRT3gxIFStAs+MtTFNlZRG2qOhh8TB0PwhqZUQ96ijPB5eUE4me
93B+jThrXv7JqkCXGNBI9392d9MrPbfuRoQC8MuXFE0fTq41XeOF4jXwJdEBOdD8
/YxfdhqlRKwLYFGTXh6nsDFu3PZH6aJiPlGsCpm0bE/Fuy5WAgR2zcUzvEeKWbni
fEnzfaCk9o4733g0MmdvCBSjRbpoaHQL5zVHkcrfPmsjQXOm4g/W0erhKVF6RwD1
wrDm1rj1wjGE0D+Qn3y8s5kIm/CJdHtQ5orRcZoWI0TVYlTuyN6UIBOWi3w5vZ4e
9hXIuOqxD/F4OGvo/xLeZ0XOcKQnvt5JiWZJ/XOLno6qqR9coBxG6RevQ8oqy8Cg
XmUEpjTCoAV2kn5rGJ40OoYyHpwOtXo5XqtQUajlFReqAOImpScKHD5+6zTgS+PZ
WxVyDrOjfM2AD8JuhMrDXtaBwwzd1/8Fy0Ny06IUUOoR1YXw3KXqERwL0rGpjakg
g5HItBHeAtbGxZwoE397Yje4HroRT2sMe4thN4pXDWw/WfRLr1v5lupHYcU9Txqb
7uNFupXY/8iDmCWzg+hGnIEpUMaFTEZpUSauNpG5xCqTjMBCwcscQ/Y1Pqf2jjhb
wu3LdpXC+/dTa4TXExAt1AmES52qc/La/ZQuDgYqE478aI31CsqPwYKLpR0+DvQj
oHD78klm1RlF88aY3jdP1iNP0u77YFPDc3XWhTZXW2Qa+M6T4qugfWVdsYWysKQX
RJpJWHmLOd4dk4V/GW55Y3J6pMxCLrAJpy0KOqMTSW9ne7EWfbzcvmLd8tBZsIBR
vtIF9TJ8B1zNZeGp8gpCf8DYw7Fn4zPyx2ATEXS0vniCTdXj4tRCXl48Tlqdcm9M
bU7A/0U3lyWh2sOEIAIz9FVMZKEWXszs0zYBBo+Igm2rCKaBF1a+iS34ROjvugPu
vgTQLZYowJQlkhXk/xAzHIpQxLusTuXZ2ipezNcOD4HFfuwh9HTEVYPX+b4vPIo7
5vhrDqKtgeDyQJ5KnLj8lCTZe3TDZbz4LQHsTwkncXcQhQKwPboRgFu8zPkf6/Qg
E2DSQU7OkLKzrx+UJwHnKE28eNh2W4kobwoiCgAwRgo1xT78arU8v/iY4OrZTymN
WAgdHHyfbAfIdjGG0jNNJTcEtSCEltE+ASWUv4JJrtA73nNj9TR0cWj7+2biwmY4
3TGLq4W3rXklJhtn7XpgWDxEcMjKxoYua35/7PsPPgOu9AkbKT/omEDw+i7HEdx0
XyBU5mB3DDJtGMQq8b1p+NhIzBk8LVqBqL36Ir2dnwuYwKOgMljcRRsOiN8y5aVj
AkDvprvugVvukQI2rWWs4/YS+JoKv0rIr8C5IXmOyVPglIiGWFxX4nPAvEBbaQKp
BGTnXZPV3mPl9BHzTSiFCelhCXfVyvoQBDJbv50F3t/nJeU5Uxri02gbg2YXbsj0
mHcxmyDBuYOI1Y+P9i1MTPtALyfyJNaI2N2gH7Mvv+VZbeo8lJmb66mFzRXuzFvH
xVKvq6m4HgWqo2dpMuxGqG0ZaXzgdbhGG36yJaOrVC3rkmzS6rDYGs7l1vi527gZ
qvwnK2W6QT8u5YfSNVUdJRkSG+BPq80C5konwa1gw8Zt8yjMjS8iyKC7c3Ko3MMm
V936vigncyWCgYS/v11ENoQtpusbqgzjMU1due0NMTvwpIF6KFV9ou98k+MiuMBX
D+pCraxtqt1boGpO6yvGWkW4jtfSWb4hKSWTWVL9dDCifWMCqSrhWDXl83UhzqCB
sz3jbVYHl8ZhVLEwOaTVDqBxgF+H5LsDyWhhpOR2PPlVOhWD1rx+rIPa2MAiXq4w
8OAIgLxrzYt3uyDOrOr4X7AER9Dvl3lVfxJGQ1whYn74D0DjOqTGZPxS05GMGCX1
HJJ/TSCQSzK8ldlfyIXmCwj1rq1Q0r2nQczQVqX3xm5KRk5zl+G3D11qNrG5b3cO
I901rDJYNyf86b8V6zkEAGjF+Y9ad9GkP2tts47b4+sBoq6qyqyHxdfnnHK/BMyX
Jh+eUo1YXVy5+q7EX4ZXvu7n5PoayykIyffzEFWMYOSGOg3FSVKE/7WP9xYkUTHn
9XcAzn6v4BHcaywb24Wp2aYJXJOld65vvsrG2A2Y1OZUINZh/SuJII48kCdrcIaU
g8Gt18kr5OXl+EnyyFY40Lq2YytFQkmoFCZ2AeTzEcraoeuOLV5P19g12LIHl3aV
+hr3vfF1v2bj/qfznKRlofiRB7H/Rs1GcJamBua8alQiUjTyzthj5DuxgTACjSGr
1bT7PeukWWi4by56zsHr+11ajfndMRLJJUdDArUa2Q35tC4gGvTm0ab/M2W2i1Vc
NJ4RU7TXC+XUU7N7CLewrGNlK1n8L67pNsiSJx0l86mubE9Oac7444U+UFKvTXO9
nhHfBdzUpd4fXJIni9FXyX7iAUsnHc7oiHrZWaYjEwF8n1UZ3Ii9kpojFM78avln
Hm2wqWvZxyA6PDtoKYBoea5AYfxcvMIs2ANloVKr73WHK90St0QJCT3R1PjfD5ZN
t16aLIfViKgvTweqi2AgqOxQtLMI6zzK2aPJLzTA5PeT1U6+9rSSaJ4g/3a4NE1R
ZTvyHpGg6g3w2UEDP1Kr6IBjAkoPT07M5+SlcVasC991E4MqgE9VS+k2bvQHtqux
2+KHqC8M3T2qBnt7JrUEdF6gNy93WxaRgpnIWQWFfDXq7Be8HsiW7yhCdClKc/ak
6PrIiMR3/qgWGVrAxiVlADPWyK+Rg25bB38t2vpZUnhMFzk6VTihtvVXEp3SveLS
Cq8tGEHnKyWNuLgwHCEaC8/sCfuJ4M3X9CX5B21WshsZeOBVMcYcWKq+P4i7bhgm
NznVeHeGp0ZBg6bRa46yed09R3zDCtSdaEQGcEta8OnYFfMRc6zyECHtDdoivX+s
Bed8+1r+97+gXkqGplIRkf+AryOLNOKE45Ivy+lM/k02dP8InyNO80B2mYdBXlYi
R65UycgEI5Hz2SgtlQEx1FZQplpBqrtTE5xwStQq+SU0i/eOihjGGX3PFXps3LFe
KwDQ1KK/l1EXm53sWgIQZAT18FQrpXrjbJNYYsVJn4dnooNJfH1Se3UiHcufvfL4
QampfQnDUpkpzHgMaa9EsUC4RuesKJFdh3PCfEUFN6JImzDzLUd7toNMMgx9g5yR
ujjE9tvZFlxfYuCluoSPZTwUXOjv/NJy1QXUJJmEc9a4bNQLnmZoZPBtRcELyVGR
UbXCw0ZruD9mdTBr1CE4MBylrHGPv5eSq+EXuCGwJrmCqpOLELsKtYDVUXDIww+4
2zXfkdpfdqpdjrym3QP6aJzt/Vo/x0HOg8fIuGJkZf2d/Lo+2EHa2iZohIPU4kQa
KoqgrW7JnJTqAKG9nzyPTKDz2+h8SlvBJDMGk5YCqms43/7YipalvbGZZedrgOp0
H2MzlCE53lqUdVyFoeMHU16rPXg932Qfs+QjhWqusCwDHtcue3XsNjNRIXHAuJsV
NWylv2rNeHqXn4/ZjDg4ZeTaXdBnH5C6yHHuI3po/rhp2ET2U/oEM1HaMkwyAGbY
SeQTgPEJfZNfqvcP3ktOxBtJo5GOKH6bb9nSUCVJK7oHoIwnarOpEUFYlkSjiUEB
sgnK/pBHKX0lLmNkjFl4KVEXdB26QYKZsSkOB73eP//6yJanJG7fcexckqrE+pWk
V0YTszy3/p5DBoNda0Ui0/U1gpeThW/kt4ZcoJB0/tmBH6Q6giRoFisj+ZCQ/m1n
ZE31nr1sDL/+fzf/6N59WuuGYB82zlbsh4VhcOF69cQqakikKeOFwH0nQlO0BpyU
wZpHRQTp1F2Mz19zZn6YnVcN/tC53rkNJuHZG2LDfoUFxeZMRDZBD37Equ68slEz
eagErCc7gk+YhPt6YT62nGwLXIQToQWitCkrk+eyetPEcTYGuJhf7phjHlvxJGl3
qH8m4mVQEiIL0tfeHyHlt6sb+Ye+FMFU6b4z56CnZ0HZz3HBmWVQlbtZ//V48oGR
n1BXNzIWyeKcy7jr14y4f+vuh+1X7GbN0IeJeaIzuaqlskQSt5a7wxx8N4ySLcmO
OA/1Q+FJJj0mHPLvXHGa7D0cF4PeSiDk/2j++C9sf1EEJ1C6sStyGgYxyLKatNM9
kOvBJ4i+Jzs5Apnj13HA8gq+2QHeDHnDOKcANAMtzQfY42rO7xjn6BuxaPFySSid
P3FLlbWCqdyCZCNBm8hsMEPdtL8y0uObxbj49Ms88CJvcQuPtyb7O9IphhjsE9Yt
p4YZtpKThC2HP0/xOQ+Yy26K7IbxSo1nZuQ0tZKZzPwmLKCq3v7805eFjnz2Yxfj
4wy39Dr61WEAUC2iKDbucFoVFy4lAA/wD/zooz47+wY37g+qsI/iK4g2M6FT4hV4
KGtXTU8Fi6T1RzWW69ZkNESa5VCd+r3C9Nl6kh4qeNhgfEfu7mwNqq6aaWnKmqn9
Y8+oa6PbgyMVwXR1uSTEcsK7V8Su9EJAD7SgcWoGVD5/5Cw2Phkw1vTTPtKXhWgV
xAXDr3MMIeoIu5FZOpTZHirkYxFjjFG7KqYyntAkEJ/ihOtkRdfNhwBVlAEY6s1s
OsqL1t1ROW6m8AQYySg9WHVj4ppJnqhZN4enAyzsi9ac+at5CrpfYzT4UTduzF8T
tZIVfLi8zFS34PNnh1fttnaQ555W+v22A2oQuLA4lKfgVdHyeElqBu5h01dbdsOR
x+o77WpeWd0VBCyiLU+BOz7FDITvd1NvhzjTtjlC2CowcafU4TAnJPrMXdBs1zX1
hyuM3j3aU3ZmQTOyH1jYLXjqljAH6NSBOUlDIQ2yGfr3ufbqDkgbPNWQvCbM/q4L
ZoZYWOHaTsmvNACBMYpALJ74Mr4y+ngwSPAUgyZneQTa4J5Dg7JVcyvglF3W9J0K
s9nvNkva1DryhEgZ/t2C3XDZXI3927hmnGEXltt3Xdqw56e8WXS8b2JJQoIwfue8
DeESa/Y4QDjBQM1URwXPJZLvoIeQZmGAs/cLsKzQPqKVIOru4LT33Wey9slfGpoD
X9+I+Jvvl8K0b443hESbCRjrB+7u1YRJclOgRet3TXv0/w90c2OgOAwwKF1GPHMh
92X2HPBGwxBkIp6YXztXHeUzc2RAUQidaLy5Lea70wBAu27VyzZlKVg/ihvy0ZYa
+p76PuyADBUoaUd5Jk4PWNuYp+miR2nc8fmv74hUSXat9eiKA0BJpsKDFRhue94T
uy/t30dY9ozs0LfiBN7k4oTHLoTyGh2zBIa8tvMZ7OpVUg9juZmdo4UQ9PW4FTHe
qSwENu6b739k6QMptXCP/LBl4lQ4RRErDvycc9ZNs2DJla6CwmUwaScugg8Gdqdw
hLWBqx3o8xW1rnk5pFcjwpfkpuuv6gKkvTeCLeBdyj4wQ7D+D6yd6RAAkcwNGLUw
b/NGU2zGMtmEgrwCcNsyud7iZmj+EOJYrPzHoD7Xne6lmVo5X3M47TrDGlRwk0YA
sAMxmiHbjVpxF89mO0DPfCmdtuVHi3KIsLkscGzOgrZN2/E3RDwM8ttCNevAC4/F
Q7RjqHSQtboo4xakYUpQFJxrEdN9mDZfLchelSTk3XsgnDjLP1wTZRNclZv24YZW
4iTzBIecVkkCFEbUggcLms2h3SM9wAvAHSc4taKkv/xuLFyOl1SSmZcN/bILIIhH
nWdHvf67+yozbsTKa46huQzkLjwvikaFelsFNiUePB9rqx5IUOfR5a+A1CehGho6
WzbpmpaLJGvBvdEet7ZnAtaUm589LSsO106vWaAROXADUQzXC039BFloaQn/2f5Y
fU9wi4rT3jq2yhw2XTqlQ1UmdoNCt0BIf5aa1IF4TWNZXTkCUsqGljB6Mwb+ODqk
v0C1p+E2T4hy908c9XrXRIvu0NINczFwyW6r0OZ7AQmT0iysLJbtIY5B074fuSVA
zusN1jEYs4tqhX5lqSs7YFQlnVORZ/Lkpx10T8tyZRjVhXIDRC7rpPO1dHOkW2H7
LiKedsE6m+u0xjmty+XBn7v/UHhFdejwBgTiBDpRZtQgn/+6RlTq1TEUeDc2gqil
23UoWJCKimjsoe8cm5FDCJv/aja7l8oFpq2XwpMJzvWfLHPYIi5nWWYzrBVGvwnG
FgxHjaJiG8RIAZP6dXdq9hZvR/sCANgV0X32JdNln5H5nZ1faPK8W+lkLaul3WG7
BDS90lOrdPMiF/wQS/MDWT61jyZ2lrc+WmPB8dmSfXYBfGcytbdVgjsyDKSRqOSk
SkEHMnKHnEm6L5jsme9AvoHHWOzo7yZZCFDE3YXi4RZwQkU4HI4y/6HAE9hN6C1K
K0Hl6aI5EDvwE3Si1g/8H0id+YMLPjHhxJ9FqP/NrZcSdEIUn6r8vwkNjfivLsbr
tuJX4MuuoXxPeJvt/KlmKF+Uuytnta5R127wRhcP0MaR+DuQx1Zk64Ye9KchWi02
/IBtND2sT0oyNMRVm909ON3A7fKhQ/VfgKsJMpKg9oScESPPii0bH/sPo6/3ya1n
5nj4ug5wuf8iWQ+c9NP4Go05bZm10kaV2YTaX3zOaIczF2EBiTqA5JRfK/QypWQw
VRPAo3ey+Z/8DCbv7DL3NIR23jVrppj478XHsoSZdItwGI8V6gNq5Fbf5VgaXPLi
oNDOZ38TOPA/jVoUkEve9P7CglAuDkZ76o8hwQpWOd9pA4iUo570yraNTnnN/hkn
DzAL5XJbRVSWv/XhP/ry2yAg3TRQMiICmXrAL4xkef3oxAFPSV+9wLF8B7LUdTqm
oHCGCKbbKEDHaJTb+zFhQq9J8HrUs4GQOIhe3xfh12V5m6mQ76SX9jg/tKVIOhIX
06QqnhS7iymwbA3I6BjfOq6pkwxS2+lXfBXGQ8F4uk8AMjDAu4Q5KQV3sjsFjv8z
NbnceovMOyzN4lr9vMUYIa9NUUneUzVxVz/ztVGSKuyQH6rUgrvGuUBJ9l1D3jFl
6qo9qQJo+NxuT4/sZLWCKW50m6AMQUxj/934eGraYN7rYIEDJ7yjcIXdENAyw2Fg
Rygm0GDOQgA3EQ/fGQ+GrwJGHlQK5qvAOKF41WGu8mQ5BesUQxbX3r2GYnjX7ine
66IRZd1KVgTIPD4HqM5vQCL6pRoOjUKQb/+fh95qPPwTDqfH6uoiegxclooIitj5
Io3vFpUbd20KJPwqk4fdlK31BPnaQHLoxwi5D1zJv1O4qcM/XpbWJBkNuC/OS+yS
ZNzf6zz/VyCUqrXxc7ESuMAxjsTraSTA+XYagN3suSedpvGMsrbj26ReP7ydOl9n
jfCDOBGIDsCY+WDDkyqcujXFMZkmlZyhiZwkkkd4sNr98zxa9oMQYF9exjFexyUg
kQLuBDld1nYxu09tQBHbATTzi53D5G+fgkEPE5bDhfErSX94Tn5SHesDnMhjo1CL
kLV+ESocvitVHwDmqcH++gBJf/DB9S+M3Ydg5p8d5UZPkTwIdo3uSxxYtJGieRmj
iw3WYpY1+np/W8NTGjQU4k5HY6+nEimnqNnnVPyWHQ3kVUaKrig5PJsNVsXjq2Eh
QkmTcPJbSHzgeE2fLbwbTCugDhZH6gs8AjvH52WSkL5K/IjryEoiEA3BJCGJJl7S
K0oiGKisauJsDbz8VGdpZgEVzKAZRA6kQYi468skmaSQoIFCkGkqJFMABH1h7UBG
Hos/wQmn4MdAvPTFvXEEexsI6Ln0RBbad4Cfn3Pe7GZLhHSHEfbxR43wxFh6/MhZ
4CPSUHvA2sSvD4/EhWJo/MzQmTm/g+VG8Z7yqnqjuhrYZrLvPF2EsX9ZqOyWas9t
6n8jWyJieRHgTkms9OhY1es2Oa+5wJlCbXy7Hw+vxttopWDIzHf6qoUBVTRuEqJN
OZOWYhDBpOb72s3RFIAh8xl4fdSeVxvPOmc7lDg/O5R8ZOrMhGQ99nve2+5MHqaW
Fqul2m+c3EmMLYIGCTvQjetDOz0zaAkAU95E2ZyqqJCBZ2N+Xc98Vy/ZQBGxD5Ci
FAHz08zpaZrexS32WGQyeHPANzFAhKOtqOG2IleQr1txS0Qq6Zez02jjv5/7ffpC
YMBJSKyNnyquNUFMUIzbM6cGsO9iY+8i4pzug+BgP3fmNwDMZ7xwfRi+5ab5yhyW
YQ3DsZCkCnUL5CB+h23J480lvzU/wdlS5SelJgZ1OWSFoFKS6r5gdePQpxlrqvlS
SCONuPP0X/shou+UXVzjLDZ76QO4kY263/BoUtSe7QnQRTMDKRWgVB0Orfta7aY1
nO5+9Gd4fke1QKGT2jBbglUOLYWJTju/7Cxc4toMT8dtAYFs+U2EeiD6I2L1C5yV
w8PJqjpcadwOWFLiy0UBrbaZvdPqS9ScrRjllWLYrNqMyGHChm0lXb7xHMTi8AoV
12iIvfvVz7Xooj/FkdB4i+wFFxAmcdIZBC9ZYKnbX0rgU0hm4JYbMWDLeOiSr9Jv
Xz/skJ+B4axVUkRMCCKOzMpIijoGAc/AV6bbWMrnmWCVUAZfLgkG4KJ7T0J/phnG
+1OKEcrSmOubTBKCRw1E3J5V1zsFHkSJWIAitMmKgVj0fcn7Ln2nK7/2CvzdHMuE
g0VKELsC6AF1YDjrUDh0X9e3dilnrdX0+pd69jEe5I6QADI3duzDr8LS+TLpeCu1
g48c+jYl/nwuJQ6zmKjDeaShm2UB/wDglONxLDYtauiNEasLPlFY8YKdq4lavt9d
QJbw12FQ2JA3LO+MNR//5RpgGU3c1rIhK+hCmTwhk5UDLAqRHlZH6cL80hIIjxtV
TLsixr9ubZc0jhSgyGzNMmuxldvvzYiNwJH+22jVouxVOSfIvl+HBANXJ9y1wngw
ibeVkMDWXyDYgmsxV6cwa4XNC5NBz+6qPRbHTsAso6t0jwuuGr6q7+MU5y/o7lB4
n9sHMQvBsaF9Odzya5dNpLh+XK5XF2MMpaAa+8epNdHbm7AhwcI5en+GY9ttai5G
UIgkgMzmZx/8xjhfDuLLEgSNb/I5YloVbckWLGMzcgGPoGIOvhO9MIQ7jQGGYK7b
D+Nbl8TWR27iB3POazfs8bLog1rM1Y72N0for+GXRde0ctmc3kgLzcVqEIjoficQ
ZSf98E3I2LxedjtZ1K0myALFW8AV20Wd/Je9c7UjgO5Y6Hp6+bxvbec1NqwJzkVa
ZiNWSq7u6OUMvCb9ehoNBU9mLp5fvtx6zjdKTcgPe/p4TPa6enb2RTzXCqIVOOP1
VF5xejl8h7Pj0Ukxq9xsgdWx2FP6O6/cp3Mr0cwhWafE011VnS/tDbpBaQnRDyNa
c4iYll53QMkyIWPA3hQYv5FR455LAbkcjEFfIAh1e+G9a0ChjM1DON7/VvgqohmD
ztoW7WUL7qLMrAlM18w4ouybuYKbdstk+PowYgeFQCQZDQCpX4OlLYkls/8M1hO6
rlwZewBsQmDpOlCTVR8bXdkvUXxFZzggN2T4foT3UF/vGoPw8aN+9oh4duINMkKH
ob+IitlSAKNxFC9lquCsGrDARX4BsVMWXtt9j3Ps2mnBw57mjvy318JA6JLHo7AN
s7+i8ZOOYL7Jnd5EpmnxpVNTepYGyYRs/ocYd8IGrvO+5tziujIUxJ3GZ/R6eQQ7
0zzaB0KsIQRDnxoIYwgyRtFLVZCtgo6nH0fxyUSsBY1brkVt/wg+K5fy2qEnF5XG
OOwlyyklIAf9yGqvm9iDYFgiQ1Gc+qVyAp1cfOhiVSd1QcxrpZOJocxStGpiHiXN
jPbibklZXSrWEmK3ZXCnQTNA89iv+8dr2+tn8UqzCw8Rsiz89ffIulKdibmdmgWs
rzHbzCUjQcEs3udXomMNLvZjpv00dJT3IFKWNx5+B00zONenDYtFHribQsqTW8zR
JVPoPlUppcBSL3pnIqZUG7/1LhZvVYLS64EFX14U8Z8d3KJVjaQzW5K6OeOfQFu1
HO9szxc7aQTsKKJgGSSSJpttiPysz87b16gv5GnmL443esPUn9Jkuc2l0UY5CC2S
DNTAR7kycfts1E0VQPGAqQUZplyHW6gzxZNGZesQuLYL5UjMZg89tK3Ik0bhGd/N
nX0Mx9wcmm5/Kyqo0Xr6lb0HvD21NYp1YLuuL8JCU0MB72GoOGPSnmJqlAxDrm/U
zMJs71ffh06UjZ0UWRNzbHvO/8PX79SNJG092ZCLUuNYwBNhRfFtW5NzDPkp58JK
as7hwxe/kHSbyA253+tXLY7NpIDh7giOkiCi5Ez0zAHJZZe3O0jtsTUk2ng03qjI
hQ2V4XzkNvgFImyE2pqcGbvo8ujRYsndIG+IyyeuRLIVy6GN6lKpYrCGxpsWBAcC
K9URTnekcTK3ddHQAoOW9W/F2yJ0//vH/eAW267hh96Z6S+XbS0V9ReV7mrwaHu5
WMucxg6Ai4hbEDLa04HE1Gzdd7rhmwQKHClm4g+gLEeSTapb1u0iPBS5b9fwVbpu
OLklABc5hIA+giNStycz1XjhhitSU7Y6Q9cNuRq4WNuTWEk1Budo7RtNtChn2v3b
RaA1Zy0SnTbjoBrwi0mQskBZsxJBoDrTfSVlLxJ5/wjuU26rELpeQ4MPyn9AShfA
SunMt+PW6v3xCZitsk2RwdzWTXVaY8H+OoFlunlWkEcHp8+cAW9fZWCWhZ4t1HbK
sbg5P3PAgtuxdVbeA5FGKET4Ev3JXZxlUkp2zDES43kQMJGAdMgPDELwLID7KGf3
x/uAKRbbS8nc0G5fWC4//H79WqEGKp0QcnddvqR9810yWCZigHZTmf0XcpkzBIXI
Pn0ezWzgroTcISkL+lAc3gXVCn1QxTKY/dBidyMgxRrgN1QSjs4+k1Gzw4lLRmvG
N/TioI0O//h4A1EOuv+RB0oVZwHfqLrYdForki6bHDB4V13NN7ti74RaWvigr0F/
KAZqorO9A9mRtdy2UWHaQTtVmOLg6lQH5WqeIR9GD9kEJwGcCAh9PsnKGnAau5CJ
+L7PqyKAfwtahYlG6Zj6NnM8uU3YissNOWY6POvuWtpKBTFCzqzZ0x+HvobBGWIl
Qo+ExTErFdOD9gDrailzU0jaEBoF5wu5lzOCTkIg+hulqfryZ+AMTT2IL+kq01ya
HZYDl/fIlIUtEuR/+L95CSd+VulfEMXsTKnEMnub7kh4qUaC+qFt9ty84eHjZHcH
0tSYHvEB1tiPSaXGcLx5bECNs38ZK1sI2e5PVWnIjbJm8VCmQevGZDY+vvqWzY23
EITcZXl1zSVuXdK9gy1YbbktJm0wBB4jwXbmhblmwCRtlc1waZ7i5MNPkGvXjlFG
k84jLw1hgzfDjd5tnwvcOeLcZEAJFFJNiXhNZ0ObYIfPClbiUpW8khH2ep6lPVsu
JW6KyKMJZD0U90/MCTlJahSXKBG4l+Ew1JqH3FCxp8eyajkbNSLRiW7Rl2c3Jp82
uPOx8vcIdtIDJ+UHI+TGAhF/iXg3lN/YvTGiq9FmVpzJehE1jicObEucUWNPKhkm
jkmsj8gIw8GUAp/RPsn0h556Q3MjiSoct18bt4yw/wPVj7tKQovcv9MQ/d4wGaXn
VKxUF+YxJIFVAGdr602qYpZVvDhs0x1XFDEZiP3b0FaHOogYIK9RgLDySKucGfZs
zlX6Q6wVQ/x+MzTP1Z4MXgFbGpud9lvohxTfAxZCzuDu5H5jpZSuAvSy3+k6P6G1
C9wobH9wngLWBE/DRcKdZEuIK073OZU9jU9l8319FJ8ZcbDBaL7sGWWI8n+Fj9mk
/iHJL/F/I56DCLKTcq9yJ+xDHMhlLvibQviP1VZ6VldE8uOKtsAYTnGefktqDfvM
ZeCvC4NvM8OXSRLE+2BaEQ0/ee5lRgRpANCI4L5Mzog63Gg0gP+7NUA0q/7xFq7m
YOcFIRfCu3WRtCDI2BYScfaOy2xNh2ByAcprhNE38jLIdBQYTD/7S4EFCJL3csre
o9XR4XdhOjMJi+MBo6eZLgdESRYbb4VQjOLU08WcFiASTc1O1wnc05gfg9dh8yAG
ag9lWc/6hXaF/1iJQlqrsycSv8CH4Uyv/YHJ4DNfZeWwTK+1P9w+UZNJ4DeEJFyd
G7tmQ5GsPtecFbOAddN7W7e9nAw7At5cafIcObR1HkTLpZLckFKyY6KHiSXV5nXo
6NCVSwDAm8F8OPFtBsugmh3cQ215YHe+y8qySt5zmDAlRsEDmwuQRK3xk9oJJYeZ
21PzE9CZkv4F76S1Z5tOfBdiywnkslkBHRer9hj1KhBMCla1B7vugFotePjlp+V8
Z1FLWGULjl+4069bVzBGyTTnWXuKgFqibm1jsBpBG8U8Ilu7RutcwLH72YxpU9nJ
JFc6o1RLbtlzL7twrdAYlZdEPz6xI532DpJF1BpAyDKXZ6sCCvU9GzrQNeKSACbn
aA/njxv5LUEAOQOigmGkJ/GYsK+KqnJOi62eYtoBlZl/rtuxSwX1ZVMAZUPanx9/
HzTUscVkpjWF8nkLjZRkDEPaws3XdNLyT8vjkRsxuAA6N+sB/bWF1R/gfQnDrfxb
6woWtuU2Jc7UgXnIJK/EUt+UurTBfxDFLqguKNjArrT8GrQJM7FOamMLTiq5fVIm
R1jF66iJvu8/e9AAVlM3bYWC1tagoJwk1zZdDEtVHyIpJGzBlubmnR+Ga98e6RMu
foq6hoHAhB9LbhPoBaAt13/aLqZjlOfO7qQC+c+u4dn/ikwVvNZio2ttjtAPMK0e
rn4+r6q7ESUWG2qWqg5c8gRUYMAnxf8j68qvf/KBVaeqZQKhCVd9Rw8FCSsBijny
hR2ElKlWVabD3VKjR0rfbfZZnaeLSDjEowAqqKNQ+0S8Ko6UfFWxsVW4Gu1Wt81C
BnuyBaQeOFO94MKsziRnfopwIRwSfm/uyOuopFhr9q2ZDY0prozwNmLnuSbbS5FQ
uQbnrghgUxZwLW3V3S4tBvBkELzs99Fw43d1Xc45Lo2LwyM98Fsku0D5Jt1NijS/
MqyOn0OfuqQeRnO32jjaUWcYjV2l5W3ymNdRTdsWr3qui5A7Qlu/JVxPwWWsG6nM
8A05kmr97r8Xxk/cf8fJmlhvWkfv+nXdwS6n2Fi4M7YqYgJnEHqxo7rAd1kJ2EEx
lXHVz8E3xwmrhv0PP5aZVTkdNCOYqSvsf47B7FOobhUZ7OvkMzg7zQrMbloW5RRW
erBoYo3a65V87Ad/zNLsOOWlSMVac+JgQE3eNoRqgY5L50/Y4B/Iwe+PkxeoCVib
Bv+Gzr6HGaTxzxhn6+vx4UYgbST663hmu65r5dORQAOMSoWmKgd9Pkd5gs+xoLHN
I+udKecHLZ4FqB/EtPFVoQEPuMTChZqqJh52+xt7H/Q2U5OQvOqeaOtbw6Jr6GJi
969OqhXgfi4iAFiBNPQvv0w+OeeayfC59DzWqOx8qkdu94sDF599rXrKC+BTPjRX
nroU2IfFE1sabUpoee3RVG6In+CwHQnRW3fO6zGZrx5FC/74oxLEkC4V5UgDXkzW
8j+ryIaBgAWt3oYChR/OCAW2vMrBPFUF9iPL9VUt3Fl6kQjMqeqPxR+yq3xIU/0v
jJqpvjWqTYuLmUKBs87Jo7H2R3u3lU93X/x0d70yh9kDQ/QOuO3q2qZTJH1N6AUG
gzc/klUIip1iW764QwFLpGPbSaacVX1cqtbp5ds2u1bGaftqWGgkRllbxwmEZ8/l
wZ9pkDzCRGve/BTVt64TJ06zAhzNHoePPpMl1V37SXVbx2cRF/MQjxSv5WCPDl/N
Ocl7skxZssFLqP898KXp4eKlZ6/3gsdfi2KW5Chb6Pi8EHoaeKS7pnnh4BxRjIRe
wF5/bTgq+TCGNvQWvCnTvYiVUoah69R407mhiAO8y7rmAqE7Mpe6YNqmK8h/lMtK
QwORyZaWK6i3oQZrZ0uCim8kL0UlzJV6uS3TIR41Tbr0nhFHPNzdgvkBPq5/B0q6
BvNgF5nKioaXkUgxp9aazhrhSfPRj6PMTBUqNZZYuDGuhn77IytEDNDO0cDudK6R
Z1Csv6qafm0oMnwkH5HrZlP4bn8i6FmCkNIXaKGPHLuZM2067fmu9qG0oKWmmWoG
bCzQsK1YnV0hO6wF7o+efm1szWhGzVOLCR1ZaR7h/rAL+L/wI0Igb8dhYtcQ+9am
1cUc4utKDx9NHXNqZSdwQZRbUB3Uy582t+EHYEVdpfqw9B6zC4dT29soOBIsyqc2
qsiE+sqh/GXFhG9uBaUozinD4dUTrIR8NUPKpG4D8q06YRftOTqFjhRY7g2Ep98t
aZY1i5I9h6mkc/X4FJW7LgnutXb6DpLt9oxuv7frF493rLqJ7VPpD66VfVL2vOKU
jHyrzIvk5LbA4wcubWk7MnHNTXphhRwEeOGLF2/iSp4KVec48RDumrMCBa3+3Mzq
217gS2dA8PP/Js4Nq+PJzavD0sWPh8dOuWtHHweyW6LDTkdMwojdSMqt9A5AkY/F
8VSYT4WSF7HpySwG+mFJrJrwmDexRZtFXPSJmGyz9Ix7RwUCQn8aXMZPECj0/vmE
ZuD0UPvk3E8ehcEBnHOj2SfcNzVUA3v8eJmUpbTQJm2isQHRAa84c/EgN0fvSxGa
ZIhCYQj1ksJo80R8+nzfVrnQYn/ICC+Rgz2/t412xYbtqW9vayAYQlgMieV7Ie5O
0wF+XmfbVnJRydx2pG5y8IUqPwaXepRjMOC0cKycc/TzZyzif/wLCCYCtdsn6Lmm
1k6iaN6bUkSaLwdxCeAYAL/WlpRyOwlhLGFgQ3MKWfGCbVJX4oQAreWJcDbRwRFI
OyJj6xaCGZ27Qwit+ZX/peZ+Rhqpp6Zk78VJ8UVVxJU0GBdzeTR0tnHaKr4WRlR2
POfnwRVEvRIzlN62uxyd4j3elz0vD+fJZ0tKvzQMup/nBaB8etvfxYUt3msehnok
fOl4yyln9h6I8PoK5u7wDsIckFuyvKjjHwp3SEwiHIcy3AOlZN9w7wz+N4FBglfX
hq0lsto7gyFkCnV/fJvP1jMRm2Y6s6e5ums8PJgZsreixfuCOfOioxDuU0VWmKKk
7m1bFAHuczWTClMxIBjp3FqQKHWFxAnpdc0vNKGgMpTyOHSmJormRjQILcAWcHpL
FITOhQDUpT2w5BLvH1FQIGbjFru5ki7tos4JWI5Fj5qYSIuW3rs7wYHricb77k6n
joBXuENq7i0jlr5BD5FxO0cwdKABj8pUW22RQxFCctN+hFkzXQUjWxuvc5Rgnkwq
XBEq64FpW+InhBVWN9eoDujzDgZ8bfYqdlDT289ARn25w6dNTp7Nd5MT6NLTX3xd
BAUg8M0aXDUdyLUzJ27v+xpjEfCMkWi2AzbwMPzJzZj4CnUzW6mm8SZk5wZRVX2T
/hHqTP/Bvj5xS6E2jVgYiG7dOioCMR9RgcwSCHtergB8MEFT2BrMG6gyvQBO3Hh4
mQTTpjdPtAZLmFpJ30+wXYN2iX3TgVynbXnmOgJEkArkRmTxc+kLrtl2seR5skfd
UR3YnfpKIuKps8E2cyS7idc4C+nwTTRgJ4oIBRlHvu1QU6aHCjAtZT2Wi9wwFicX
g4cVEATQW2g2lhQQ22YK8T8q/4fdX54Rlay3P+iC+JAuzgzhLpZKpvhU2QzgRXXw
8eoPbfiTs4yk7Bo42CGf94CP62BGYtae6OtN57+vpgO8TPKLLK0kQLiZNOxMqLpZ
PjN16eSM+Wl8a5cX6uoNk7MhhtmgLWTm/WDcaAOMXSEi/4NdRHTGj0f6ZPUewhxn
h+EzaM4NSdLn+34AvGWSi5Z1aPYH2OTf2JtybBB6YP2H5M7AbY1+8F/t5Me4E/lu
u55seIEEQBbgW8r5tjKLkvVaEY0cvcfT4Mu3r0hqg0r31ap+ReMKUPY7CHg0cpMs
AoBkol1KR9OhkSxdbiRwl7KdriNLgd4C62CYxMBnhgn/jD1jA7QQp+JklrRN+ySU
FWeUp1Vzz0RiKmC+0IEgbOXIIKj5GhaaEIoEfYdLzm3eDWQQT9YKjLOJU8HVjvCX
ch0yhtuYLH7T7cWHF9EzcgBi9LebLatWBkrb/U/n7tumPkbDi4KWZ7Vz9nK/nAVn
GrXH+N5Tpno6yP2/cQ+pBHrGvp7nUsF2QIb2VNKtbqyrFGK83F7kpE6P34SL+6BT
+USXaY3sdKuzV/hHg06oy9vD7r5GO+5HXqvUjo6UbIHsQ8qRqChuevGNl+2biZNc
XcOqD6POVKuWE+/UyW+e9HIQms6KgilUaOxU8/Zz6T9mWS4i+Lu+WpFXNuaNFum9
PudjWq9dNCahegvrKSLS9381a4ikN/8DcPsrAHBH1WeX6YPhFSdbJTVLT1vVUkmi
GS/PkR/GzK1R/EucEWw+H8b3sCxxuDAOcNBf1YRoBvorw+yJNdFVYslgY64DsnaQ
8BYTVHc9C4X+MN3hFfaxiIkD5E6DTpLFlldpzNCpVs62GemI2kkr/5xUM2FNFNj1
S8aqOxYgpdtisKoNbl9+iGzbbSQBr40a7blV8d+aOw0t7n042xZKn/CG+4VxRPiv
IeQ9/9R1dO5hLxpA974IVSGwRoelGfQFx6IFls+hMb8ejtV7r5gPR4Y9Nj0jjXYi
kQ7/31dCulLwtByIEykZdzvklWFsLmXrWx56Gguxqcdjx3X1vBqmhWJ0N7nZn9Wp
pM8GD4ijMIirTWUNZJUBDtQUDsgRQVp9ZBG7xFsEdFs3k3zqGVNbMPAJGR750f/u
40JXZL8Q6fPIBB6WoWorSEtfYAXioo7MgE4/dtu6dAoyjfzAp2jwYmwNQ3055Yko
o3j9xh1vnhi8JrBtdOWT1OX16bbwRqWf2a9gdVnRoPZu1hJgKBdon/Jvfif4XEPO
Y4p0z9EOKXkcBtwGZhXLPO4KK5/qX85N8O/cKwU7y4VxsPynlR9AIls7GT9dEn4R
BRUkvEacOqa/LbDtUgj0ImDXI1egebFmAF1JvjrBDfCyZcPYd32k9A2uXVBBmRiL
m0h2u9CZebUor5FsMWB75XjAbO1qa8erHVSBCoA8fg9EoOIJAgm6o1/mXu6ryPL7
4z6o7ehR4teWpGjdjJMmXBRNKw5zPFj7SEvrzxIdottKN7OX+eQcJRPPOHkhKPwL
PZeiCAvDwZTE8ODJx+jNewRnxnQ76JwywoM3Zy3OfyT0anQbSAXiaBJkOu7ZGc3p
+n57RS0i2rDu1g5p8+bc58Cx9OCq3cFCIYgIidqCCzuqlzuKrQ33zVo4w2p0mPkx
AQaroMEES0dpOI7BjG1fO/VCvZY8n9dH7hBHdRNqmnu9UXlsqM2cR4YhUH8fWJKD
1GUakoawVQdFyX1lSCup+fAHCyUxAFq6o7E+/bVD3YEmtrr1HyoWfvl6oltwSn3x
N0zopaFO21hcVIaddcXgxBhJlJv8PAjVEheqmlc4oGYtbpcd7o0ODhA5IWH/QPeo
72+sSklgP7RrHn99lge7KGXMp+s41ZdueB6xc4kur7tsz5Hew7R3wSsXABz9QnGB
yBwl+zB0Gw3CE3qmGhymtU2T1dd+TiRDOkWHEMdFrXtGwdYfoDVCuAwCbQ87OHWw
Y886N/181OZhe6BFLS8RxaFvfcAprqxiyTTGIttTQXpMsm1h2hf3RBjR8aZaYc9w
NurAnRbLzaPVOy8HhSwQ6mLNFNXbZgUK081C5esedQxzWxegxKCw/P+6/UQc+kdU
L67CO/aiOkAyaLcZTYL+n99bK8pnKJ3sDfQSJzLKNwnLHeDZS83ztzxts8RxyepI
a08x0Q24pBPpvTCZEgVx23NaE9iX/EGBxlsNX/lttYZiGkWUbXriGi6zsmC0ntwk
2jwPpCR9CSc8ripE+LHb+icR8NB+aoIWKpBH/NKUJxDV3WlqvGHTxKgVdLcV9QbN
GoEmc9r+wWOQ9b31JHDTbs3sp+XcLfGU3YjPM6HfrJnimOSH+2paS1Csh3nnZ5Xg
ajqmM7HP/eZPdZxMPd/ewJB+rpLdhcIjh3P5ygmHsGh62ETkfGb/Uxg4bT95Dx+b
hFeNwWBjYpDAr0+sXromMigfWuM9zujd/J03x/BnbKHVa4a2bmfl6l2s0HrQKGcx
X2l4Jf8dkavk61O3lclq7zrw/7zPro5YOoAQLqpuqyCx9vfaC6kCBE3QjzTQ0bvR
0D4QBdVd7K7MhVKrk47K1vdXus3aR0MB7WZu9ELH6C9WyCAnX+IOVDxMwiJCdeBU
2gnYP1kaBRB1MWl7Z1w//MDnc9jeBizeLHp7R6eehPIw8iQ4jNaTgIUz6VPiKMyT
dqmkLgS2jseZAL3hUTnCzVdoWM8upkcVTxnOjx2bNthj3V5AL91dxDrAqlg5fXJC
XGLCUf5rI/FdG6qc0ZE+0bLCs++QmugJ8yBLSZXwxxLMRdqc29sz6l0NyiapxiRD
ktaITUoyOvxYjcMAZ6bchlbtqG0bP1FJe9u5g7mymKA7evXwkPn7+dTHXDYGDEPp
bYZ91PMUBavMdik0kkBjuDuJK8D7jaUEoDQljLV53R6tAenYjCBp14eQMtSQzUBA
UnGqu/X4J0aJpZbU7JmUMpQFFczpV9M46u38lxsGk6/vZ1XwreTryQqgROc6b+jn
cmzmNrFkXUFmDhrvWAUpcTBLGVVGYZIk0K0oZQv+cGPZXerjDZHyp6LblsSMsZqh
BSr2a2AuGYXVI/YsYD9F9XsnlEw1YN6y8sSMoZeris8+oGTTGKSHF+D94UMc9VDo
uoOpJh+eF1eLrcTKq3/+4DOWjXo85/RntCNGcuLFg3hyn9FqIL52e70mPM0gppp1
gHX79iz9eNRqon41GobfHHgRsK3lBpikayvstPpr4+wTGfsYWPjeN4sqJ1Mgj9aE
+udhzg7UmPR4I3k0G6ksLsuuOfzOv9diVSvsk6NgVj4FNNR1hNitLp1qQJiM5bLz
RFCs5Ude/Qqs0sSogh/vVVniqCTrKIpaythHan5fT7GozfZf86WidwGrkxHe5Yu9
YIXmlCZ4hnFrv/WxMFvm5PFnfiGyuKkRyKiTN1pWRATgnSP+rhpye0ekrM/J8gnw
2sis0H1e3B/UKFjyA/0Pu1t0QYSAHWDp9XpgrZEkSAKrySLycw8Qwe8UrNadY5Hc
ALdTOl9ZoYuP3dzLvdp2OmNrk0ZChOUdpANhQC979Rrs997uuOHnZFx8dH3uytlx
RllM6i4+XLzrJfpDsuQaFq2sicPb5PgJber2dp5P0YalZuroIZS1nzWqO5Mr1XaX
AXYZeuD8U1Jr7VS1/M4A8UFoz3useN+1gz/ueYvXy+nRkliQmdUeLwOOSHpIU8Hc
9dqJCdMernG2VYTy0UMD69ErGYLN+dz4Mbuxu0d1Qb2KBrmCgKAB0MBXP8FccpF7
yEk4X6D7niPgGVMpX1YGfRn/VIQTuEX/0vqfdWBM8eMQIRc6xhwnBymOVUtgiwMV
jiNBDT6E3gGrwDRsz6ROZYIoMdn3aVNV+JKwj8LBGkh+pmHHDRhlcf2EYm9vxN6f
D7uPLTcVem0DSqQ5Am9jWumukOStbpLa+NXtsH5t7OPWSwpyyDrk+8cU0pSPeFJD
GI+K0eq8iXgyXT4MNeDcRv/vXAzD2St5oxLzNud/1+vpT2yq1Ffa+l+ETjb0dvs1
YxSu7D/G82CxZNZIalmJqCHUR+FkYVgU/xyU67Pw/OfXA8wX+2viLHqoYBTXOBbV
puxwa5+KrsaJFY3jDlUIBpWuqzjIcKFVIxBhKe0wwnqYCBBlbgbMgInGZ32sbd8w
TIJSv5OWcZL51xja3sEhpU1wpRFYdLHSKbqMdpP/rXbtz7weXhq0TwU5dfsQwSNO
Xg/iCUuPoTOroZNTxjVqivhNJ08vFoaiTUDWndjBCOFCz/wg1BZFWRtudTp1STcp
7CH/zlxENfVcy//kqsIfqlb/KuoOUysk1U6OguH4fyhWfg4zMWAJKzj1/smEAu8H
SAu+EiuqUd+JwE7hbZkZkBlYz/lGmLpSUKeqWz3nnZd3oyH5SjllqRPQK3/7Ns+g
9DebTIakeh2JS20XrisJW/kYor8d89PSfVycAgWL1VAnTwEO9GyR4O2BUad1bwH5
00TzuAqgHLhDQxXvjzS+xSPl/fUFpUcyh7ngr4Eo6NXfsMYxz59XMiLuuf1uArAs
xn/g2PbuBeKLKP/d+dxn+uNf9TIhrFWAwTmof9ghicRUF876P5/PaLTKLEbJEtCa
aE0bzOiuEo5cLnekvHD7mc1K+Wuc0MykVpiUXPKfg/GDOThDIk2pYnLcuvKVd2bm
dekwHFTYlCn7sxjkNxBvAy6wyFdga4dgqoiuU38Kz8NQ6YKO1XdIQiM1WifZa0TZ
pjSWaj3X6vc2+VLyk1RoIbzh4Rh7moYEHNFDMU9xV6+ndW6z0dQs68vcJ8WAN9hS
69WcNU+DlPGarfiyADTawrVYqaq+fPiGRJwpozUJXtIRGGgaj451bN8VLCLqGNyv
OJxOcpRkZzgJFin92XNK+e7pcI2odfg6oZc0vt3vDk7vPjl+4HWufDtsynje2Go2
hneAS8QTze/7TRFnbNFuLg13XJ1BdVBroe2A5xATRTCQI2CSEc9d6YgGTmAqj1xV
D38/31vVlJ5YLvCNHoOkWh6R0KeRoEKsOpgzS75htRF2gEmSnz3f2ZLoNE0XDVjf
/Lu3jX3VuskTEn2wB08plmDaQCBDd2df3DA3U54q3AuUpKmaiU5szcOrihvEmkcc
bzBBUBxd7dGmhaDgUytbxcct5bQwQutlZQaSsT7PysFlD2kkAW/p8x5Kv4GVTagq
bRe8bw5f9Yhf3kgrNwMJ0dpyhm5G1ZrYS9P6vA9mQ76jd6cSBefh5GcxikY49Uaf
xWOKvx6AZGfFazFqp2OXmy9X6BvNRzksqTZdGK0wkF7lHoGROECL9m5RsxvrVmqX
3Nn4jiLmopMc0b4bSURdSA/9AafnMEkxSrL1RinGcjWwynMNSfV/PvCxgc1UdhHn
zRPaSlNR+RkJmluewD1uyqGrQ1Yg2+ct+mPJqHlwddxZEZWiR8da/dtfAB3hflua
X6xndO9zeOu0UJxVtRSxOBZSeS1kctGQvPq8QKluRIp0bHKMSOS+A+8d79Jtsy4x
mQusEHico4ofBJvkua2brd+cjXMPm1Ws3KyBErqH81ZcbSb7ZE2shgyED9yk8hMQ
orv4m1S8Z+0truygZ2Ve0aa/xIQwXoL3EFYb53f2sumGwPTHwYe0icnUe0PJKd/v
6737ldO0ztgkCn01SkG3EmbL8E0vQmJVDdtaAVgtJaMmDlR7HzNHH2aUwsr4Fjlq
ggYP2wWVtBEn0acYgDSxVrGsYmAvG+J9U9QOKwayTVogyEiNuDUn3MZhfZ7WBZSe
gVUfTXdQucABMKt0Aqg+E8xG6joLTfvDSKhWGzz6hV5g2Ai2nIrTH5V41aVWXj6G
v5tYIB1+9+wt9TppDwo+AihlLkKt9JRYf+5nctRiOi8l+2LrewPGpmRU2amWs2/U
MYlV6lNIqA6I4al0jJixiWzUL6jTnD3W3gAbbrYKQhUJJFKHwLXhknXMtm6BswzZ
93d6gwKpxRJigIxi7kqrJ31Q5aPQpzRDElUx6CHF0L6jpatT7a2hvSv2vtKHtt7g
Dlp1s4H7STyJarNpLQ5OHagsajjkaJSM3rF9PI8WgFdFlFwGqWkFJNE1BirLoTfS
4r3h6HmAA5EaXbysIZpkRMY6OWqBKpNR1X7BUaC/nlUPmJ07kKbDJn1EArJg5JG2
OsWZ7zglXX05Rn+6KMo0mBj9cpG+7LDu2olJEEDHWqKHiYRnuLct+W1stUzFMFhU
DFl7Ltf+hXxSa563t+1i1tAUQp6tl80y+3Erpdui1uwLZaxDs3BQ94HfT83P3Rx9
CgcTNUBPGsx3MA6RRf+iI5xJgjHqaUutl2t6NliU+9BzhwY83hxuBuFTfhZjd8C3
rkqB6fuiyELlHXzixgh0dYtc7rrVU+Xb+ZwkjMd9xZ5LtN1hICzd354M45tOCUWp
V6wemLLQh/zJUzepxQg7TqXyLlmCiedvFTc/+fqzy89X9LAmu8dwmLqCjl0RTNQr
2L+cd4Fwkk03bff9VDubC3Y8S6NU3iEvQ/AE8y/ZmDYYpLLAnTr4C5y52SS2wW+2
4uWW/iKgKdcEv8DXiEOX64xM8/ANJ3PaGRo30okswfMoM/mmkf1eRFJeF9jlZacj
RnRXAVFsE1ho4KqlXNnjhVZRvav7fLHoRSN+l+nGy+MKFLCmbwnfrch12IfhX0Bo
0CLEPdYaFq7e6klhB6v0sZWiNsuqL+sjCoOZnQaN7OK9zP/7yykLzNhPDkfWJ60J
f8KJYzs/vOoLYudPzaMDx+NJQquAAdtkh/8b5SdxFF7sOeMYIDMkCnuV5hm3N2RI
wbBxcMVcfJ/sUj/7PUGe65kH6u1Vugm/4nbFwL7W6OM9pBmUKX4Pzx4sbJU5X4a3
OsW8ryHVHtNfP7UyHT/kl9r2UziMRzJzI2J2OTFy266TYBzgmSttB2fvuJWkxj+a
yYPDDkdggqOc2hecvJvw3s57TaCQ3QzXTqpNfScUcvmBK1JBfpG1m0SW263SkXKN
CAopEfIV1c3vOMSF4PyxmzepLD0ZkOou3gfaPNhFvNA7u9x2dLrCnFfyxdogJ8he
G3hGdjt8h31DWCvxVyOxO+4FsY5u18W2D5xDlFL0Nt4gJe8zs3U2cuKFZmMSAuNe
FVVDgZf/dvKaE8d+LHsfuZ7cryq/uI4heV9xgCpdDZ4uDHSz4a7CMyOg7JJbeMLT
M9PPJJyxjVzEVSSLFgxCksK5O1jjnLtuO2XaE0GDBTvrHIqRfBVyBhvspEwlYJ3y
xXc1F+4ZlzsSzOheg0vV1KVjYpQMWNgsuuXrub7WGB4wM5sHfr2zHuKKyOau0ibh
HpXMM3YBaH66P2R8rK7kAD/kKeT0C6YYzg4aTbeMOLi54+yRM+CHilh3sn9Vqk2J
8TBzaEs5slPdc0YvXprHkA9s4CT5nJLK0Es6v15l7vfhpNFng4AAvIiNd6omvTQy
K8vVKvKGcF/KNb3zElfcjaL8STYbcQX/0pyhHd7WuYmKW+vyjl31ZiVVGwLrL4cb
NTx6PnqwP75pI5zy3ce+UnEYZKyvUNCdUaD1lI9wMsdoxZPc5lmRsY6fr5L+l22F
FnZS87cMNu4XW+ZdsSJ/hdK3yDQbhumXGAhiuGfsDCo7MyZWvC9WJiJ+buI09LV0
Me36gVB4snI70Cn+XbOsfFSM9HhIHnaUuAA+6KHiT/wPG7kbpMGrYWpOk7Xzmu3v
Jg+m5RPPVUOFIDMH2KaNVClcnjTah61nSxCj1epwU4xuIy9F/0Banz0U9qySl3e1
VZY2dHLkmU5Mh9CwBtV3AtTjqmaGY48TwpZ6xSIdnPCHCHbctIVXqVgxsJZpwz3d
2WiiZjTSqlomhD42W+bmaZssMTK10wT5Tbt6Trg2u+68J1M0Wp0FZvHAwjM/rKqK
aBnAZ8ouKy0W9iIlwq/pmpgmRaAoBiWtYS6OFMntMSv/s7r9pAZLM2AES4z8Iees
Fk1SH7zB0yNOSiCfdjrM3ak2NEw8WWgxQGz9ur/xI1N3IUpbo8g8gbLG36F5pht4
AF0z/Bae06pmJGLug72NAgCNUHs3JVBytUzMe4bF9D/QjpNLfCKIJEZ3ofCTEiew
OYfCp47XzLjwP2zyh42nuWJcyz7xZT680HfZ1ED7LbvMCPngZZKiPsbPFrlfusnt
o85yjz6B5ULypWrH8gOnCfEF4geCHpmXdf4SajDe3rjKMKbOVFkGtpjXanIkgvDq
PJetltpUUzuy5oUq3eh+IXb2cW4pM1rAfoi2d+2X/1oevbylD8x+/jq7nZwcqdQp
PSpt8fsPq3+r2vxgfquBk95sFfGdZVySPuPTcSsxyO6GHc4eNffutaRP25pQ2ksB
/eud4R3N2mqo+qGm2LUj+iK/e+Lkn6qfedJ7VgVLcDh0pYyloK/7wtTh80WM3bKw
UpvoOTmzYjn5qppB+GS35OGF0Mb+JvAKugOAAfjWCDaODPlKTP6lmNh4ODsu3rpE
WVJUYWcWulygEX31Tsk37+3HPLJn21Tf1KXOGwc7sfk6O7+4EH1QS6WTdXCiXppy
/o++JHrry2TaJcE76P4xP0NV2XpvLHGwyInTmpsQWJeR5pv/KwpOjaNxLuUv9krw
27qbGsq83ql9zKMBWmkzoqUb/Tbg/Dkb94x63CMSiNwBnFChx74TfmBY68qsJrbf
rcCdh95NkJQjRKP6wx6NJS+oCT8lJvIEboMY8tidfnKvlzlp2cmNqCVZQmImtdn0
dcfK/+3sprAKRyOc/lZ0XjZPnkvhR/ZSzLEzPxQC7vWcM2apLAeORJsV0wOi4RFq
UJwYXB+F5RfJeA58NfUstsVn3GIeG/jo0iBqPtu/6J9hC7o/KWuDiPCFlezwlUTO
mfUbn1PfghVA68pefOC5Jr4woFczVSB3nnp91Qk99+2adiKBQxoP1ez1LysB6Aej
aQrBv2uYjpvkK7qNlifmVVaOhGuvEAcDkqx2RYU8hdPPrqRxesvHog2f0t1mCV+N
GONKqmbjBLnSYnWodsoBi/1AprYVrSTEVkkKYDogmOKaGwvv8mIAMcopYRm9wkvs
Qg7iRkuO6qcKWJWlHZkuAvhpk2mZI9zE0xxifNPonb7zac/ajKlwxFea2oAQEY6d
IFyJ+mUo09lMUUcF0r5EyyIL1WhBG5j53n1hbonwrbSX9QJTQXjCIG/+FTvEvoNT
ULmzVfEbdZMpPlzNjR4W28z1VUu0Kc8VBd+P73BLWpvRtp16/FO78c4wF8pwpt10
5nlAWOCaxe4B5c+fq3KS+vCgn+OgiZl+YO5LYvw1JWji37rH+GSaPOl+gAUCDGdl
K2ZWiL1CWlCkzg9TmlJNMs79BLCdv453CCSAgQouXAXZkPbU2jOKZKIoTwIdPNDb
ZNyKgXWgysGsoehWTI6I69rEcXI/MnZ4IA5zeLVUGNCikr4YTQggNacy1cvaBEm2
XUJoUcYugLOvWEOYb1wWDSG/V2TZdkhGxOHG9sWRiT29QFkXYVSD3Ytn1tM1A9+m
m6YSH+c6qk+bXculiA4o+iq11PYOy+KidZ0OiktmlE45CjadF0O7SXKHKv/2BNdn
OKxewPidaXNr9xZE0S+tzjKdOWz4i84sF6rbSiB0DEB5ewDytKYJPIPJu84gEAYA
bZSzqgJ1GDA8/U4r2h1TBrpaTndsnZSDmKia4ymjwSQOOEerWDrs83gBxmGe8uSy
I6p7NOVpjwOH/syHfP9cHRoisl3Zrb8w4F+R50dC2wLIhg8G8ODLHl+eP76Ll28U
n6ugpFOSl4bWPe/MCwaf9PmQuaHfiQ++TYAYDp8VJXEEWhrkOJ+xmkUIrcjj9dU9
Wxg+LwH5jn1m+DBduknwcq8QUKNUBFDYY6oFb26IE5qgjQMu4UP7poEcw6INlB1F
Jt8NWMMCWp2wbN8GQa2i3VkN8IvXg4mBWWVDX+yuS5+XuDnh9gAsFd0sLb+tplUb
zM1fS3p8CRNkRyDqKvGmlcPs6eveBxWr66OHmqY4pWBEPgWMDKwZCmXVNHj1yyn4
jLUCN7voTSg1GGLoBknUnW7AS/J8iWRRJMlloQVkBdbz0xAJRXh9oUDWkt/Ak84Z
0TRB1HWuvPi+1BiWaGX2K6/Rq6qo8/N8EqdAiyslQ+CJQjWNm0/S1+J/jO9nEfZV
45lVAXdd/jzLnOyvxUf3S0hxzYKdqAHn9wesrSkRcM9hdGmT4SsrVod0JC4WUHHd
xbOlibKXwGfhfkqeZySbqq2uWNqn/kxBgjjQ5lYWv5kmwPRR8i0JyeQ5hni+2yHO
TXFftoTmc4Ot7Ch8WYztAhaX2TJZzUQnclZ4/5hw2lMxD1lbcyQrUinaFblrqJ0f
cXr5WCJ9wN8xH1vpQIJOnGI2+UhBQE9H8raxJIUVRln8O+e7RcLBkvwVKTjaYWXU
lQJrIRhVIwuy8meAfA/JcXg7lNze/6go4VRutIrXrhPSjpvz9WFJoCnyUGmpg9EC
sbPBY3R4p81GMRhMxnFgXNMqe/EIgscjgJAR3doHbTgwdmmmjvR+9bB5iDq+k1ql
QkwzJIdE5kGXNM4OQpehvcNpQ2IlByroYtAsnuasALP6sN6REo08W8Jeg59Xva2Y
RjVACxFMJVEEwpmXKhRGKJavHTa7bc4A7BlcE5pM/Pv8SdtHlcrVMEWsw2xYxjWf
q6riXkl/vg8KAl0sP0n+orQBB/VnpTfSwMBgwVvUVxIZPaz3/U/adNIq4rEOMe8/
Kc4f810d2dxjp3GwTzVUpMUyGlgqONsiTcqszAMfk4ImU6FoyjFVD1edA/njWScN
+bexWIQCFcLD2E6t4qezFTzJ+fa90z5cKOacg9JJrcS+z0v4L4vgsY7jwuM1uiWp
WFKdLEjmIIEeg+E+s/vo8+Lm/0doe0qLkz6klWSuJsnhzxQ9fo2WLAjw6407aiid
s/ykssCNjgwNQJf5rHEbEma+lrG8/WJmHZ7XroIYTJ/0lH1v9POZY7/I4xN2Ieor
bYn66bHD6C0Qhp/N0z+516DPG58Rdg4E2RTXE8Yr4iIgzM8nvgf6oQ74dR1eeSp5
v038pL73Z83k0AlHTij9mHafyoQSpW7hm6yGhXlIePaCwqxUu7V7NTizpB3U5rK4
f0LWKwtYaPhokMRKgvZ+hfuLCYksSjL+iJtirANJHG5tUBmyI5ah/DXFCtZQeSPH
+pMIQTHD9gkEO1ABvTFtGe8K0+hDE2zI0N5zhAc6ysQmQXxJbAJLD+L5a6Du1S7W
csQYmhaDm+9UKXuaKePBO5KZjrN62f+aYqYhVbBc9JbiM4VpihmN5Eli1tNt2+CV
Y8E6tZ1ByurYpvc5wiZzbymi9qtkq/Wu3AtRv+Zx5cT/stCFXAurfMsju53ubPoM
tGERllkiEZlYdgbg6t2GzEKyYDvWCntt8MMJc4Q1Zn6i3q8ES/7wkSZtfasl11Kq
FWEmem/ZFkcr88JVyspQPGJitmIs26xhxytyZQU50sbFUMy3hRMY6oRbROCfM9TQ
oIrzpaJoe8lGr3FyHmUUJdCCwtssK9rVIW+lEfjk2ZwB9xscWE98O/VXoDACuae9
EHV9M2UiyOTrdrxQZWaOrvxy5Yp0iW+o3hC7V1fNZ8FEuzFSYEbHuvApqSixYA2Q
ZRxq7k/x3qv6UsyZ4XUrAlunVZMBt6+ORp+4bT48eNzdoz/kyNIVvzQEm2G9e55K
6GSI3QWK+ULGY3QelS9eLbBiRQ4F0ah4iqEDXOj6Dx5dLeyodYiJxzn2aNlPcxEl
DDvrDb0c7sU283b/4KQMlbkHjYdT2vPR98AogIZ8RGN7QjEAW8ZaetTZ+fvVCzee
dC6OTDLNdvhi6B0Mv7kC1M6S/WrRXz22fnywOHDXZssTu3lSsKntTGhWJESn+y8l
piaaxtzUEyArfCnKA5/gLoQ7LLal4GTt8FR52Y9OniIM3uzJwx5RUs9im6peZH4B
MbP+ZBCbI9s12TsBF7PQldZeMFAR/3xk7IawZ81Rq0xclJ/RwWrUVkAn4l+GR3/1
xj4sCunuvp0a9bFd32fMhM7dansyrdkZbIOID8lriuhZBjbjFfFoQBteXUU46f2z
b93mbmEU1sF0WJO3ES90HPKekihH3fxzA+UedO261dNBclLDfGk/aqL5cpHQnm8N
mj/8UeUkr6TpoFFCr7ujKwX3oGJdcJi+PenQ8IPGoGPQsP6OmYrYofbGZ26GETh2
t3USdP2GUdLvP1RThz/HbWQvVjW5Tkomj5LypbyNiF5UVKJvALKWtHzlzwUiiBjF
OxVT20a+iQF18TWPwNJqBmQHAeiWkD32BR+dvgMv+r5UwnMfejaIw816TN9SK0+r
6A/1cEf6p6FBUQHNNAQDVmEBa9tndE04Ql3EcHBTtFH4EOloy7u3rz+7pRQXPO4u
Bw0291alBY3L+hhaV6rfG1KH4Kzc1lQyLlYAWBA6rFUBENthyBXLh/HRvT5vd/GC
LQisCNeNHOlP2+46Y6XSRt9glmd3z/fJkZX9rifeZVTlP6fbIq7ows9fnC2luB2L
8mtPqKRd9wWmcgQhnb8dvKGoSKNBlTEwLd6gVUfIdOCncYhJdhPiFY3NkxuE3mS4
CK/DaJmSzJtJZRkdEbpDTg+bMdJveuZrLgqYafj03AU+D9Pgv09SpwrJrs0yIiWk
mZkY3CngoFZsAOXx6ofDeDtbT4bP/8bs6JOGeOoo704DD92nBL6NhTc1mwRHfays
r9ipLROAIz02J/0epEiNhiT793+AF4AAGtZLNl2vvdrU6+kgJXvjUBODp+Cb1ihb
E97dbfnuPf9lohQnoODrpwFwyMIcTJBbyObPKwnltTR4q5zdcNk9mx+u819APQZ9
zcXCyr2GGT2TXnCn+ebRg3pCRajYowqEH0VjOViUftgsrqEuAfJptBNYTFMBSDZz
Nr+Y7MIxd9cOoBxghq+zLw9KpCImtwUZLbwS8RAZEM8y5/Wc4SA+/pRLQioK8FuJ
9tbk0aRXhHcN5QrnlkfVF1JORUHHjXAA3WBMkfgiCV3yF4Xb9VKSdT7PspPYRcOh
F7w6VQAfAi5lyh3tlMu9fvlXFPC0kqyiJDBqCBXDcsnVP4gM7MtmQtZQRWSn/BHy
52BdjRZ1EV3F8Pz9TaZRYwi1OU8XUS2DaBJHRLBOf0QqFiF037KkhYt9N4L4/dWR
bKUMr3pGiW72RLik0MKNecD+82xcvFkKi9WGY4epxrMUQ0SZY2LGSyIKdQz+nufL
XngUUqnlCmgfSIH03/H6RB2JF8tJANB0oMPk64dQA224tYGc/MtVYaWzdN806qkO
k+NJeB6SCLgWfx+OervGCx2WGrpW87pFy2teBQ+DJsphejcE++0T9yIZLPyzjmGQ
xCZx7oPDawvpIc0Cw312AR7PFVHAy3+3kd6Y13vhK5MfxXHFtSE2tVb4W88hUcYr
EA7rtOMrH7L9pkGRtdjo6x9Lb+oNolhKnJda2nnvpgWM91885H663wnFWkLoIY7d
CywfZrroAcEiKIcCXcqMM6rQylEdzb3HhGG33LBBzoDlAplE00mlk117HbDETL1j
FTdSWpBUSnUm28g/ZUHesciRI25EeuO9v1jvro8/PJkTUoucKHLmCcsx8BAIfp6x
7BitcCUDvM6fJQJOWgq8mMa2oXsGLpGjQKbUPqHWejAUh2P/9jevHiBk15CGZXtv
fzIeqeVwsBBI1/1Aful9UqP/gbeEhGujWU0HGGYtaCsdf6kms7ElbTJyAy8GJdCw
bjVkK/xbS0vuswrhLjWP+NSv+fv+C7sfAT3dMhhjpnYrks8YzAWpPV47EdbtEm77
OHgPihFKKAUhdTXLDEXViECkH3+5PWHQKs/K3U+CyDF0vgblxQFD5pyZ3bWsT+AX
hZwn4cCZbzIhC0QT+gVwxZd3K73cNnqsdU+XBIDMvNzoxvLDlulJO0w4YC/1gLt6
4UUJRfjG0zH+lvWP0oBTRSvzbni1N9o4mzMa3VZaR1QDTzySo2IkMQuRjo4zCzJM
AF6u+CD2H1xy98I8umMIPQro8Hk1+XwLF+EuK6H+CTDHFg7LhnaTakkrHrQaL8Eu
Ff4W942VKmNmhrPoit0PLhV3Pu4YK7A1wmR6DySc1CXwm329it9Pc1Xh/4W/ydPS
bzj+4gSDU9KytIiHQ9ZZBprzYfOdRvFLjdYUvJMaPz2h1akYnfboMERg48v/54Pk
kDIMTBC9lXxUOLUPZMarP6K4DMOG+0rpZQLMLDHMMp6N0C8+EwJ2KBrpFYlg5LPM
5fpc4A8DvOhFKIXpFPsdISrW+Gdqn5iE1rTWbuJZ5d6T7ArYUXRM3HC27ePPL1Ch
71atAGvB2WZUPP14i73HbQFjXtt5sPQQkMrbWkycFh0a+10AiOhODv1udOmatt3Y
XwPmScgRhVbZfoU1FMZ9Jm5ADFU8wis2aOnw0CatiRY5Vluxkb27e3jwVzsYRg2p
Wvsvpo8gedK/Weq60Bkt86lGRtVV3P1hn2PrV5OQ0mdhhoQ6rqIMd6q8mfiNGaYl
f04AcD5+ycGKyeg1B25DXloDpGuLkBj+ZJ2Sa6mYY6Pt70lpd/Mdtn3ilsAuk6wt
9V6a7rg2CrG/4BKG9YB1Ks1G47GPWhYoI3+ewbiptDtWo0SRP+1V/NVHRkEnkI8u
XrBr7qfXzaIE86t1UnOhy9bbrmYshFnGTqMWafv0HaJWGYUZKGvT6mjmL0XuLz7B
bjYU+duJfTZpwmNQPFZS3FKwhSDre5LgQpBjHiRQRLdd5YvYV0PYMyWwZJenI4Pt
mB8r4B99RW0pd9+PVzcMnfBAY6c390rKvgoOrEHKp9Hfa4tex1NlYV2w+Mn/xTN3
gNT6By638BA60BhDMBKap9gsPtl/OsA/9HN4/hhusYR/ZzbU2fSg2r/ycybT0mjv
M4sZngNyP1g/H13Dprz1hA3kXQ/pG21aNz9udFhWzA9rodS5XN3peXZh8wVSxP3x
WfKpTuJFcFBRaBtAMlPgSsP/uZik4b+MKULjgYK3nFCnRcLpj/aGyI1oXaV9STKG
xJV9ZkBbu19PDe0TK6NrEOlj/ruqtlU4cHGdtyy/ndrT9nmPNja/7TAuR1q/koZ5
garOp9gIUIt5ZDvAHOB1oBWNuRNOn0OiRz4VrcQ5SsRUq9limU/j1esDYDYNPtTy
5dGGVEiN4/y7KTMQbbYZhZnPUaVx8sJctggrifXYSWwx1PlILOIsQVKCft4k1VdJ
MkZvIdym662v2Ee+l3sOPR9JU2DjCuW2Yzq8dosz1pJIT7IpJ35+Evln/h6PBhTI
45ddBIwAKpeDX0IPsrF2Um7otsVCLKyaOZ427m92Mq7qSOrv0M92Sb2doPHeBk6L
SDxvPo+12CXow4r9DgQDXTjyXsT+Ox6KyQjYova+/1LxxPKWNLocxtGssXaJf5Jq
nEM5GIKhxfNDrJfJqAlWmJsZgJcEwHGZZQpf1xLs+gKxhfMAI7fif2hqxCJH5RD8
5ZYJp78i375OAYHKav9Dk3TOnTUW8IaGFTOJL/umw0DB+QNBxARMD0W3zI548WIS
OySR8nF0CEU7oeI5TPNeyOe4+KBsNKegQH5tl+bUCMlAofjFxV/0f4ZNP9l92CJD
vVxDnY1ijzkBCfW2Ad6A+SPEOafNHbj3SV/m+YYj3V/5OyeYZNo5TOYPIU/EwQgI
3JTUMH3k9vCboYxpq6YRDOWMkQHSkin1xkQ8bXlxQK2+CGA8i6Y3A7g2evSJiW5Z
7UFY78mAsDWcrd3XIZlpai2Nw0IoT6SpCCaOgh7hQyU8LsTyfa7nfDLL08o2EkRe
sL2DJ0A4FggpvouqhakLHuz0hubqMK91QgYroev93eLqB5YtUu73gNVdicHS4b1w
GJknsrESTEXyQsHOiW5BecA3Zu/iOL+BG5A571rC5hD09ySkVBnSXC84N0iv0m8W
1FEkv7YPW8caO2V/oUFpIiPyy/6nDGNQUmUdsn91ieDbymsVn5PeHIghuvdMyFfO
Su+/bIm7nS6iEy8NzuFTJuevgfj/Ir0C7f8b9MNmgjQwre+y9z0xD6scqTkGL9xH
YhHkYjR+PrbELAK3rTLrm1sP+o75QKrlVclg1D6Nza2Heat2E6usFRvTgTkw++Aw
lhhYj6Ae3QVBfoUneTU2+i/5OqkuzMyGnEXqC/THcJvTHGa97Qi3PBel4EMYw2AP
EmRhNeFA6HBhCxurHpgiyTjSkfu00FTVTun53hAZoV0mcN8EMqwBKm9Ecu5LcmRR
CI+Fdl8bjqevn4GxsXgYnxdXFnr7ZHmPkZBwjC9amQVFrjFBWxTMtFWU+vtJQx+B
BjbyyJDcRMC4XaUd9ricRhLFJJLW20xUlrd0EnrsvrvWRaGPBhefeOJgm0m70U0l
XI0lhERWoLH6Ao8u/sybV8wTzdXhJpNgdPv16qYgspvOrCdPlZ/yTIEGOTiBumNh
l4y8rhMlbirStU1ZkeD1f6EF8kKhMAiGWKiKgV8e73qlmtfwV/AExl7hSZZgJwcU
B4pQUvAcGVWquPZh/40uzeYkuSCXcFMQd54soXl6HJPsFHfcIzB7iZ4MQMOmugOC
7/LqKk02gZE494kxCgFrkSjNRaROgU+NRs7cFbu7RcSznIiDr/b1bY0ZoZ0tW1Nm
sEOOK9u6Sev78yiTOOq0JyvxEA3wet8Zc7cDfD/HsrPqb/cPOZS1sZH6hvcw1BTj
dzDDedH2K/6LAXbrAYDSozYMxascK8nCft5ctBmp1V978D3EAPRL+VoglyEUc/jR
t6V7yQZglSd8P51Lv8moYmbcxx9/HK19KGu/CWTqBJ10t48bSuvsRU+MRCnRkzLe
0TW5gfsMegkE+HEcx/pxXLzwOx9gbIcfJ0qHJ6nNSVkBuZZvDnifO2KmRWtxFrEy
62LfyJg7toYATOgB2mhFe+NVKWSpnbIb8LglM3CEu7B0eLZ0jjsbQ9NFKJYMXuAO
3O+QU+7mAC6Jx6M+lxcuqMt+qW+mQIaT6aOqde29qdLOmivs4OzKsJABgvnfiu5C
CW6Jlj/nasCYOIYyWpwoO+D9MqTLTflXfnmFLB/UrSK0+ZnQy3phHto90yR9a/iy
b73HnAao6n/XmTjOh+fqgAkawsLvPK95Gn/Z1vy+5Ka+HSSzvDzlXlk/lKR7QcdR
GYHga9xRw5pYniyhvQgW4M2Ud0ehxuwjZj5cq2SwnsOFX29lY+q7vmCVVy1TU4nu
EVZ3oNKuOq9BOc9LFfqYMvR1HVGQxfibUIFpQXV0vBH3JL5qTYUufOO9giqBzMNF
K6Wg2T48U1r7N5PNKBg+JtJgPqM30iAeLVxDOUJVVxzb15irjKQkpk4YOnNKksY8
vZdg8//jro1lNKgQWnE8xTu5MZ5fpo5WAj/alrYNgjm3Hh425IKVPQTojRmK2S++
lOZCLue5g41MHdB5e76+NWrMFwSTBYIyekXWzPV+UuilmRqoaUCNBHjMQho2O0st
LVmywopLa5NSh4FCYJOh2RmjIYz80tfLMSHTGs+t3CLs1qZXnZ1+6wWb4RSPgGr2
IkVqgKC88k8rFJnNSNAPGgwK4jAC5iyjid4ISdwZQgZCfDlO7HHb/TNqNu7dIMl+
yNxutZmOInY1iNSCpmqceWDqmfP8CC8NRzMbD7JbaMbFNR1Ky1eOkquVP72g4IaQ
leAvn1EXey3u8h83OHKgMP5fRa2nlExd92q4/+DZoqsS6ns9uO6w3PnL02hqAm11
q2I1lYbGyt/wmL9Ke2Viv3XFEMV/eH4EkcySHrOu1NsUQmvT08zPTq5zoOW6m0Ga
7cvAurCQCAA01doTvh/U8WO0jpghmpJRIukg60iHR7vjlSp1Sr470SZ3kYyL/63g
HWwtgR7fzIvczt073xdgHOzZR53tRVhKbmNXbWrtNwrNNYg0VIB2pmXKvCZVNqh3
Dmok4Yl6c2dq6+Fu4epb8ldSMZuy+No4dYX5n1QQr0sXHOeIYThRoLh1xTE4k9Kc
eO6B7gVtUEbs9VHr063VDKxPT4XzlEs3/7vEtydDUe7udrV5q6qVoiUodtL4Pj0N
swZ9ettihCio5uLVsBx4n5XInhJjPw/15s9sKhQpy2XJJzzTn2WBBFiONCq2JgGv
+asCjaD/1YgoKp5PXsxKoOBhZNa9CPP4Nd9Rtt8wLDu+U0NlAVW9LEPLcqukxJW5
D9BIpG0AZFXglecye/cqAbBBCZvXDt9APuX0DD/rQQgNCDmRnjSQpkaZKSNHF0S6
9YNmwzs74Ox5saqe//Yr3FFRM10bYNiIMEfnBq3MRKhCer3HXoFl3WFngjS08ij/
+29GrOOD8CBlVvEYoiyWzhG+yPPTp/4jLQzoQsXqHhsz0EvBpNXInzDo8WAwcaA/
brelo60jAAcOv9hkliZYTe8BQ1RlUSvmDriCt2nmNrRq+PT9KcgFhIRcHHTZb6fo
+UNK9YqQE9/DfI5g7VWzbQACxWyKoLRmf0UizzIHjPKTqIm69HX8Fgtf6/jpvNhB
iZj+tiw/vC+NUEn85u/aLJ79/GZQ2hWf+r8IBxREKWRIf+M2Z6tRt6jkBemfFDsL
IMikdjtLjz7N4KZKVOlKzBrC6LrxK5d9u30A27tFhQ8qcFYRgFMIVGU29UTMNiOW
5gUDsPyHOMzoPHvNZ846JJ3C9aMSOnPeMxQGEznAJ6Xdo9X7rZJeRmz+3LSd/f+z
35hx8zJ202DQncn5hDYtbbB/ODKMyxuYOAOVbWgBthW1PotrMJj9N3C95rV61i0f
tQeqWhZbsH/xaiM/ew7wfbueDKeITqpZEiuGyvwindB5f2jPCs+PYVltKkz9k5eg
kTyFSQxzHtBVwCwLHrnIIpm3YXzQ4j4Y6frNNxixsw+XNe7qhEnQP1J1QPWaFEpI
3npdr3ELJRtAaK1TRk8jlxiBmW3+WNUSN7MTA697f/7KxGcIU5e7L8QTf0kA4Y55
+6oirSKvgkCSAUVs9qoFpUp5/bODa7c+LCZWwYI0ODL51r2CN9TVHG/kI72Xze8J
zxnfHaGYCwBsgrKELiRuZ9a486SLIEzWmDYsAeffa9nc/9dM5LdCepjU4tBNZbxP
+JoT76wFhgvN8xiSPCbv1zTGa7Z9mBimaVDkziJeNvimzF9aFHh+1nEjbO678yX2
5oEOKnlpfBYhsue1irDJ6KsTMQQAItrjJsT3iREm5Vb2CnKWxR9qJtgOcjvd+lqC
yGlwc+hpcNLh7CKFaMQymL7ntXRSIJJafGcB2QrLk0hZDU+g5SulyheNgKV9nkLx
Jay3hJFATSF4RMGKnrvSKxVcu6ryziqrDbzytanbmGBHcRI34JXHgVqCibrAj5cT
E9ttGDlvNo+MlRpc0qEITyYnGcnydRKLhCPackCyDiis7QZHAtQyeQqhzHm821Du
6v0bSP58stfbePodpgcEsGlslP32DHE+PPkhWXQR+s9WMwkVNvQkp6R1PjKQA6w5
4GFhVEQugSnssd3CstQrvCD1VDLnjfv+4KdrUzX0vNreNK28gBW0JNRhBeDGPIGF
IFFBX/C2OWyEzdXCk9iGcFYtNR8/198pR59iJcq3HCYhUP7CzOd8XjRaGp+vDfcA
QISINvOVxQoGDdBAy1U0d8EmQ7WGKXxR3ujDCFH1m3kGc3Bz/IzU9P09ZSNp9w67
sbtiZszwULdZYxTgF9PIjbN4zhyAHeTVZsFi7LcvC782B2Z0xz5Z66irD78M0U3H
ezxuMOQD1SJrUFY9bRwvGjTVjH8KD4ULsOCgA0iIv5QIayei1+DmerirLDAvtOr9
8tOe8VMDPKLWcn8bCY/nuxXNIB5emB+E2P+184tsEiJoOQB7ClD059FeK5wYpRPe
3vG/P3OfAK2yuY0qL+XJFL/WbPRPHZ/N5j3piTLp9Peg/Uyj0cyoGGyg4MBHtX42
2ohf8qSuED5Ckotaa4+kRrCFWChvO7H65dd04w6lWpRjLnQtinmGNhtmM/1Ya3d2
hYto7E07rroAz5TuM0v1YETyH8E8fWSb3EiT6kiRDfjqIs55nB/0yEdx95aDfGwz
yqBcBS2GdXOSvumguyn9JPxszHJtN5IMjfw9sGUTFDFS6PN4zwFtIWjOgMZyIZIi
WAvd9EIxReYXTl40TycrNojvXbQg/zRCQsOVvX2btgb/0VZqnX8UYDFTUOlCNAHo
k1ba7irAkU8XE1R1h7Ba+0vfU2Nfwt0l4NDpu00wqacippViH3JGR9RkgA37BoeZ
umKP3e/LRoflgcrZjArwYn3rBqYyRJ2GfeJbxp/n0YFLV1EtvqCbiGaxZtYutjIb
hG9l/oOXwtQ1oVrTtz8ZUAdXKIlOLg73ovNHQZdjpy/46/bWiJmSX9UCjfzYEwEb
de1iB41wYh/qKEtcnowgyyQbW8bAw5LTbcklKqRplbdrxknzqHjoTo1go/1OoDnK
6pd9svqJ8ZLRldaTLvSNsLMXBZ4gXm5Wk2e1fwR+H/9PCHXU8REMQAdqu5k1UevY
RdTdtp5GFyGUNF4XFgtjawxJz5/mnksm5iDxJ5vp3KYlmuGKCYu8wKLSNGLzXIQb
ihaS822ksBwDRxjCjuSoZfOdMfleDWCE0lGrirmx2BAlRW6Llce5JftCtIueQLoL
FIJWL0+3eUxTAOpcA7qJzLUxTe94kziCSSNfDLmtJ12Gzh/BHotMVY9Q20EPdCy+
EqPb7NxEhjyagUelxA6Y70ZUGcCeA0ZUkQ96ng6BXzFnbFt8lXpUSdz6dPeH3fxn
yxUQgT2ZFFYmReCas1BtBSYoquGoCrXhGXz/aNTEhzQSNfaeUtlrqUlb/8MjrAl/
Hciw+GGzaDhbyQ0B9iUSYOx+KYAIXLYj7IKl+o/zGKMUXuLh5hgual2Q4kCxbq0Q
qCRmCjEK/uUiv2q6zXdpS/4VWvDHSuSLe1ZMB2+GwbNjBeAhF2FPYdgkoLbLsmua
Db+ovSxysbE6oJFHP06xiHFqQaMs+R35l4tZqlBp6dgFdTioqdbsLEf9UdNZ9j5Q
uV1BdGH44erKsYMXe+sutXxMxv3yJSX4PjJI+he4ygxg8PIwgnZw6LqdO3C+vTwc
O1VYr26KdXsTPccEipjXmMaarFrCyu8m+/WGlvYMlx0Q2HfAhKEo7iS9TZsygkwx
aEF9Wsif9BlMI4ay4AXzhrAHad7kRZjY2GoTdYpTOYx4fMJWAt9GyGNbmr5zL6kS
Z3jJy+8W2mEAo2JIdqgqv97FBsY1/pv60Glb8Q3FxBEagVJNZKalQbcWfyNjuypl
lCMyRPjee5JRV5UZkdJDO2qvc5EffZrFsTkGO0a0tsyJMqCbtuPREL2aCPVEfUjL
Qk9rRPO55jqWem7oF471H6+pu+o6K9QpFPNrKPCoxAEL0OM3eYmY5KIsZxxAo13A
HtMBMi7NuCnsaCRlKyNyc8GxvxkdpG3iQAmbuFl+8urFMnczcVKeZa0grKkwC/BH
RK3YlURJ/7BrSXZ7H3wNl0BYBI3TBPtklJmyQLLGrtIfBSOVojGmBnzmojWO1E3t
pYYH1BJ4In9S7dWl6Rfwa+u66lBFH6FX7xcKVPmLB8HyR46vvMgtqfys/s0UTY6d
Rf6yF8rRyTp5B1V6VZC6dpcltlO/2t8q5pBSmhE0bQx0hpH49o1ONEqsJvc+iHNw
j7MlEJN0nbcna/Pfv28rrT4pJcG452K+aVNSyr8gDsfO/IPmNtW9mceM91hlT8TT
jXChmpqX+QDbY9YiKzBYIjtYLxfyQGIWynWs62TPTB/ly0K2jsQTfJRzrUtwVXKj
V4u0sSwYHxWXABR8MHf4UX/k6reLM9Ucr8Z6+9NulPAovApHeP3HyBRByEkq/5Im
kuAIc6gy1/CCd/QUekc/n53k5nhZiyfZ3R/Aqh0H1hOB9Z4RRKwWalha4O1cUI8d
Saqcq/MXqPgvgZRyh2iBrO26ByDciWefG85blYzNyaeXGnLykKxuiVOlqWEw1a0x
xw9G1A+ZnhviIkzNrAJOxWPv7oTVAYt7hqCaMnzgoMrqDpRvvAkrB4pQtCz45bbm
IjP0zM0CRm+HDXJ/4uxh0KYo2NPXqiRVXCSCh707t1pisfKTSLyICEjtdX+cnbnb
dYI2qb1cjL/aZCvRDybF4+XPGawMhje3xSwrxGtQ6lx9gbNCcaU8Ev5jLEIVMR06
Fb+z5MWCQwSi1OnLd+gAJ62zmsZWE5cUT0chcZyDd39MeLknZ0FkO3GpbeQQNyOJ
sS2vR1NVxBgmDpV1psrw9md1cdYcyirEWOwC4hUSctTVe3IF+D/SlxQw95ahqndi
OXdMMgDLT6yfOPdLmVlomTkNBXZZ8YEcmI4tC3vqglPSkucxN8pY6MKHG3x3FvvN
+87hXTyhnhhE1CzmAFsoD3algPRULsS7OfiFG5GyYWEldeFy64M7kz+vmQ03iGaG
PQ0WqtR+a1vsZVhpjYJlOitrQ0wV7VfmB+sXLy6OyiqAZE/f3wyCr9EpcAeclPs/
4IAKpHlLdlwpfV/gI83iqrAgXljlH2kXnTFyL15iR5B1f6uI+1GnzF92Q67EC2Ze
MkRZTKrE2kyhbJcK0RO3+s5ts5HPOGSSxljwevOBeZhnWkYn8Wicxr0b6+WloRY3
JGjmXo9L3YikEq2z+nzjiusi1C/UT/mLYlDCdFNXYq0nFeai/dn10BkPgUvMum3Q
l/XJKVtwdq/cTZpDl8aWdsDf8yphr0nyZ5aStUm1AHD0jmNgEbVHcpFRG6OJTruu
JEeZQknTjeqsxscyxjVNB4WBDnOpEUxDJn11Y7AgN284RKGx3UYxrdPqeEA0Iqxp
pRAahBSBhVkn6L26aGCtNzzx1nt1fmQInct4lPDMWsbzuBO87ZoHqUCXLgMjiKBa
YxcKNjkz+2PyfAY6JoLTZAg2b6COeGA2RHwHQPQnIheqVFw67586dBPXntUe2n8s
tdWya4dXhVMoGOBcvtY3EycLi7Gp8j+z2TJtmzg59F+qiC0j0r95F7H/5CU7+TqU
n+ELxSMLBnvhnPj8yhXS63YPASQHruUHK9LD2k37626KcQbuq0cPmXivmpOG9Koc
7FXkCKXc8a33d1bcITVIQS5W1bAotrPUJVTvFNIX+RuGwVVtA1qCIzUDKbCya1ob
HNIIFQ6Wr++cN0UqJXhdk3zcMwGxLKGRQYwUlqdgP5jntLugI/JSQFka857p/VQg
5OBAZRajsAoN8BAo6mw7BP0STczSe9y7Rp4jErXA96qD0lXemQ4fbFy2FTVc/LVL
vqHj/eACr5RkneHZ/08AS4CssaLoR1hglX06mTb/kHU8ep9IvY/n8mFIt/Cdjg1y
JR2HjXAGViqDqJZ5Z2uYve8I1tpmjVJ0bH3tBdSv2kICOi65eOLRpsOJWzgLx4EE
H3LbL78kdDtFn5AxC7foppg18W1iwoJ104QxsHAd+rkZuTIrRmxze6LlWyvtW8Y4
lr8GLtDavKEPcWKaqE1L3N2t6OWEqkSHPthB8V6l591okqCEBu43bQdZ4RvuLOqK
HA/XUURYfq+tFO9guwdjJIZ6qv3TmjP5B6xqq/J1/HzVo8G/6914PCTu4O5iD3TC
RnSjvoBT1QItS6NFvpSVvNelW9Q1UAV7suhlmcXvPMBrcI+LdRbzyMC84mLWv/LW
S50UrwIGr23Wh9Xt995dMhl/vZJUM6IEJr73sHaengHnpVlBvxycvo9DyfVS/Ca8
UodMKx8MO0jPEdmnS93xRpDNFlQc4yr+JiVSdcwVDRmpAj3BnS/HKNrlCHMySC4i
/Ksw3imQ20KMpmCBlDYlRC+O2A/5H9Icq6HbVyLCdtGURqhPnH+tU4dRAWebzot/
puNGn3NnpCBHhh7JFk5GiGWSex4TwtJb7OGmQBMb7puLwIH2KxWvXVywRsuhlPlg
EwzEDcRmS5y7+5TCw1ppKdOnmaFCxWEY94GDsL7QYFfHrneTGnqoQyFMuq3Hmp6V
HccZUVc68hUfzKlmVJNz7LhV7W4A4GwA22aEK4cn03/VB6qbgkCe4Oyt+1rIOjfS
NtjXmlDmh69f7aYwMjcKFZGyRpy8CxTxgWm5WNF1EOhRSNSvpv1QLkymNa4qyWDI
9kCrwZ5VcHj/CIFosMaD1Rwz0TfyES9b1Lvmu/aplWHzswK++fxuNiMaiyePRE5l
mXoqMsKKo0bTpi05m5Scs/nzu7pQ04upEyhLuUaRMoFOxmH2QzFH1Kz/09rnsyqF
vPT41YLVbTwx1feD8B7lZpVDe+v/vlY0YeukVn7kXOsNKbm55rpoNxq5W7fJHOXg
f23DpwQTdWp9lizDN1if/635+q+hk8GBRLp5vZNzER60w14WGTRE/O5rkqFcpXxV
Ok3Jcl1NA2emk63K+E7PanGHBEKJP1P+WdBKhWW7Z5CA+2WcrqbWUBYcwk9z7gJB
I2pgtbHbfTu+i1eVxgO9Lxs+M2uEQaae20kQHzIm7SphBCWK3a5pRTq6pdFUO6cY
QGh9BymylXihtPO+SBekdwRio7bUsPfgBje+A+zph7AVsQwft6wFQ743nA++bcYP
fcQuUdz3CLXbJr+Xq/4GgWqiateza9bEI6qrGmlxqwCP3O1B1BIEd/ls9Aw8ILVH
ZM+SGggLnpUeNsMN0qhdxya68c5L3TWJKIRHZZPLATg3OyALdevArr94aiXX57o9
Xow2mxNge6xwyfoB2sVUF0ZRXUxVTs/tn6WtGSAA+qrFNcbGUOMK6NPsWBU9SF0z
beSzAp932oiwQUrt0NlPtFwRfAhyhqDSGMg8F6hXfqMUM2s2RpS4gk2MDcT3c/L8
55F0HXFA8NLqv1I++MtkCIsf191irV6pQGPSyljUfIXPIz4rHRaDKYfirXhn1FLH
9uCyjJ3+hfENVhtfVMOgqKgw4bb5wB3DFHse0IIBtYegCVmaLCNNSOBKFZnUvVSA
xFIpvUwNAXtF+8+ba4UO6Mn6l2DuwQjZR1UAStimhLFjXOLp/UgWaiCKbbmqDuSY
HWX5ZzQJU4h+R7vD/orKSWeMVWNREY9xpwqxdkbOXbVPPyb7TtSKITpgk89kWbi9
saNNZsGvchUDm9dkvUYI4JJWDBy0HNs4NpoymL+hCKDAfE3a84SvHYXPC1JvIHpc
wfTarQeiZTxFR9cDyXGzz2eIrnMCo1a/wH2Sj8opLF1SwgPeo9ye1By7BxA+L1L6
VR3N98c6g8S6c6Ls3PPtVTz3bEAVhq97uPkXxk6O/0CkLFH0zzEVmXUmUbcJ73M0
bg2tH8OW3wnkluFu3kIDIWBCxxg8FQIADp3zB17FI/bzMo9+pXywp78Tuh0U6dCz
MjIlQz3hhM+Bo63JY7J68qC+EuE/g+clrnY1olHvund/8IudB3c5i6ihpTVK1WZ3
V7NOBMOcaTT8mTWj5BiR6oq+DumePeF5u9f24W9C/ER27rb32l24grjus0QI5ah5
6pRZndFgXi6rg5heqSUiXwup0XRAdnknLr10k9HpuK3W6kpsz7XtzjIt2u1dIn3u
h3y/E5uupXQf1XoTClOEYFcXI7dxqt/iXt//wgYjJ/GJi+NhBcO1kaDdR3WxgpDH
LIblrVq9MxrgP0O4vbqIdemCYWw7ll+lAzX5dz8AANTfl6txPr/CuGrqyBDa92o8
eR9kecjD5WZvrpfyE3A/uL3JXc0ySeWNZPSBmCZBHPqup6i2QVt2BzpPzEcLW7gX
3odv5XmE3yBdt9Ko1v/tQp8zkKoUggkLXAW3G1l0+P5CDiVqFWCTBbX2ZHKEd3XT
FfIJdDT39lgq1VPOT7RG4rXCaO6T/k/dq/MI3qd2NqJLbPiphXPeV2RaL2H4gSk+
jYKpBhvauOBggq58aRGof917kNuGXyT3H41fBKwG4MiQ5buXrq09GPATQg+2kKkx
PdqjILM/c8nHgTRUAiVXrwTXwaEyBMA1UzEHYH4COfcGJu96uvLSEvoPcxHTp+1c
8oTkGvNecKfLCOOTjo8Mny9zAeDhmm8KFeVHZ8sjuKxiBwUbkgdQl4PxMy6Lbtrc
Mq631TEjDSlr8UbPlVJ7jfwUEfDsYrOekNPLP+TWRIblUJP/EFMDsqZBSHJ+3+JC
k/J8BlJw6bcYBxodI0/9KjH9tT3mobgsCuMPrlq8ebTWCDuGTFPHrD85lzpR2tcg
7ZEMUHBilQGQfjnVwgRnwW+hvQyHToxsSp7Su2TX/O3jyKOd8jZj6/S+ZK3SSuMz
bxe/UAChJsD+BugouqH8QfoMGgNWI7F3HfqnLxMCKbVgcZKr+3FQkzUzSzooEXK1
cnqtdKY4fm0PQl1MXthMftovnrT3hamx3FilK8ku8RmNFTTtLWlk6oyLufPF3nC1
l3NPcLTfGuxP7Yi9mtgMbBoaNXBXmmN1JKLHBwm1oGkRyfozq143Dhk3m0xbI/K6
6LSuPRUgZnGjF5GjGgVbmOvGBdFA27kYETKLq8xXNoI7nEFqIlqceHbsNRIXeSDd
1WyUjywVUTcWDcBI+QtRCGeq5EZFjHQ2zszWC2MbwcX45oCYKWGwLA2UP7dBiRVV
Ws8LFWMQq6YgI2MsGFJFfX3XLPBID1W4rLSJCNVfXEiLJCEGNwE3imxCJg5yBBHe
7ayatVi8Jpv5RIXpCLJ7G8/2R8I1GHTJ8i5sORpxbcacWi+4xlFLJcz2sy4q6J0J
QFfNMNLaxQ0L7mDOupgVo+gRl4smasLfOLZUAnuudYiwOognH44qml4xlP/IlxZz
FNbSD78n51Hd+PfMca+EIRuIQtIloAaEprGIP8vqjeLFXxyBm6t88ecKtJ6khwJf
DL8RmRotIi1THBKlKcUEjcbS+Qzfl0h23xnVm5DuRZQC9ced/P+4EvVWAGwOC03P
/nAIRD3tDfD6w6xYGRyVyrEw57qpF5e38ZIhVf7856wZYSQKE81P1Hf2POcgdLru
AgjD0to+GCnAwI4zyhaj/jr+KeVGQvoQ3mjwado2Q9bbZvbkNDAq9Ne+SvZk4VD7
Nz6Ci/CaMSCfD2o43mQSzu5t1eTcbEwP6OfskN7xO4vr/OC9X+xA2eXIvIIusoCb
J1zvfcS2M9eHH78CS+Wfl8ykuWzUFUY7IDYwf0/gs5WLRenB6UtI6rznG3bmFeLM
IWaNIx8n8FuafRnVK9FstVDuVstjZ/bIOTIaS5vsxx1CBrvNHM2lfDVvCVvU64Ey
EtA7ZlCpjsBdZ9v9GoLNUovrFChP7REL5nyckw9zCEFORYVFl9+Ka01XUBDMbORF
QAp44IHZW7w66ICFhSfqvwccqDYGp3RLgDazQu+HmcW/pl5RXR45wKacjXA7FcWb
3VCaQiGKrvDiraak389ChHFICFlZWfV3dRvlb/dAXqA6sQC5/7+hSG1pxBdcg4Yu
sdYyPY7asd5tpR8OqjO9C4hLLaRrZUwOuLc/R31TkjPN5dBayfwH7QTp9+MA7MzN
rYB9ubo2XhLEMPMJCVQOZ+fTj3lmYXsW+rDtRCo44VXm5yw2HI5RO2Lvashshx9e
OKxhsR2iynE9yk4JUtyiisyehCyLM0s5YRY2tRUGICg1vXfcZiCis6U7styRC96r
46ekpr6T4Rs33dFhul1+UFQt2lT32e8BFoyzynbxVTR1udYIHHrAaJyflMLLdmeI
PrQ7rB5NtA5JVqtLJRoc7YH8PLCNs9T0p2mtnohaDH1GZNuF7XD5vt5ihx0MGmht
uhVYvt8GRtBs+UCSsri8t+Zdqz7smPKHJHRoat4L9ZLsJCEnUIeyd93Hx4rkIQQs
gZnEXwJzXI9ZXoiCxOMF9GYsh1aIkQzb4FU4ftkFcp0qhaASQQ8oqRFAB7bbptG8
C1Mm8KtE2HGHmHKw3s/G3EeP0Fy8JLQr0UCTqKMweyip/IXMxqhR1aHTmOB7HP03
NtnadNykTb0gRs3J4tfIa0JTUJSK7KWn22GwjXY85jIzfSo9tXdhIO7xAJ4mz3Fx
HXcH8gUTJfucvosl1/rQWvEHhyudHjTO2OwO5MFIbOEagcSlceAIpWCtR9eaTlDL
t/tNep3UrRogDzd+URWgXPqL1kZejmukt9Jb9HdyTLdhQFdxj5S407VhNt5zyMlX
3bvlaEfvR8dUMtnTZhQ5DF3bDoJ5s1PjxYyUdZ14PApD6Jo2rqY0O6ftZlr25e/8
LHrguxJF4JU4VFt2j4byO7dhebE2Ii5BmuKKep4eNah2p7Tf9D0koHZRjx1ec8B0
lgdrK6Ch9Zp+0ZzXJM615uqz3/NIkC/fnau8BLBOk5a3SLS6cndwvNdnNUhsNQv7
rQFyrae8TQLKtzi+tN19+g+O1VoREAtJc++6Rbc4yTYnBYTpwRNfZtEu/ArIHq9M
sBYJ3urLJZpC6Olcc2cH0Pe3qYRkJZWnzgCGgf+YXC3zPyricMwJKFBMlKZWg0b5
kCT0WiQ7ueowauh8elL/1iKy100xAnUlUDR6MNKb+g71x0ZkFItFpV4aVocUey/4
E7g5286D8Xq//PpJcTtR+R6Exoeub7tLJAgNIKmrI9JOEn2p7nMyN0FEsP7rS0Cm
sPw/1QXPNvlB+mhTgxTNUWK1K4GA8uWSoyt2CGusFYhD1btPtI1CDtxIZT9yb87o
t7T1yD7/IfRcwqnfA5Xwi7TOcXpWKuMwI3rUXsF6nqZXR2IsTorIfNsfWplONnYK
dZ/kFQ0ckPOxtK7Dt8jCf3ZP6v5BeDhF3Nk2jeFzMhRvM6V/rTRhYb3TtCVw2Qxh
xhaiFEOfZ5Uz1reUB/vktbYuJi02juMPTlnNy9GE9kcwyYbtwhZl6OrjsmARKU9w
riNwBQq1te3XpCWIXZxgtB9T3hBXCVGydLcOSjRKTHfSmeHP5huF20zSoqAaMzS2
Lse3NMFOpSAcIuZZirHEtHL6Qn/Yg1DVF3X1LtXf7ca0pDaTC9KwjJFBdpCDxEo4
QO+649oHTSwKUyvwjXflW/teyQ5qZza5JroyuHyzqK0TqsnBqh0/xTjFISzbBUAn
jrYLIcDlDHUOiJIB0Ho7unFonpH9+ylgkRoPoXJaJFSWqvgkeRGxfb5IbQfHNDhb
0rn1k53E0FxFEw6iAslz5kpmSIRGqJ17sbOnuxj3djkBFCq44nDXnRNu7rWwds0H
eTqAVD1NzhmwZ2kmnzqn5eUPIBLVUV/DILXtUri4LK94xOrjMc0VMBvqwJBQ2xUt
6DnWHVJA4dpnANfTh5al2ogrbBBqTYSJyIsV88PeARagpk7xDd8PcAByfikJQi+n
p6EpL9uSd+43ObsGqOc4Wwosj5iJNFI4eyox7O5q4oVlrHyji4K/I+grNP4tuDd+
1rQuI+IiBNLs1IB1L1/XcKFX3YExEv9QbfSvG7QSezJnjsUhNKqBwaVhQefokiKv
czK9T+2qtkAdbNEWmncUciDBoP7Le+Tkyl03z/BghjxUgI0gDKvDaUv+JutcwwcH
ktcwmTOKdNLiclfhOlamhMi5EanT9BWU6g8TI1D7Ky3phM0TE117QkrhCMxfN8Bv
SNacMvvFr0y7YvU+20HoC+ser7qVZMTCoMTCJ8OPNVxLyIR4SMDaN55LBpnlPs91
SVCW77z6shvzC57zx6CU3iR13oQjlTEdl5olSgbFZR61Y4De1ge25KyBriwjreNF
zpM8PvV6uIA32zBICMBHWuqEqjMKM7Rj5El45PbGZC0NVvXTdiL5fyAU4Jap83zO
J+WKelC9dbtC/m35nfYt6KwsBcoXSkt6m4ua/C7SocMgQB870QJIoFegGDpz/29Z
Svc4hjEYnmUX5CecjoyUZVZdzfR0y2fwk9a5JOzjsPl6LxI+59KXVtz8yIFz9H/W
bohfpBIkIrDyNBvDE2AMiw2UCbe/XGP8ms8AIfNVBDESwodDxZkUNTL6YQn09C5X
w2hreBqd2xio953zvAdXOQUbj63Mqo+xdeXsTV3o0JtrkBOf8K/Fm0OizUQoHxhR
d3nSKI/PDf36psb3alfnekncqFlriAECTkrcKQ0g6oGtWmKkO8hqgsWqcv4GyaxI
Q2xa3Igk7DjLr5KbFDriJgxEFKrDAvmln+1lpdFU8ny1y4Il/I2i+2JPRFl8u24a
3oi+wg+FhZGFOPgo1tV7alvj6/f0Di5u0HEQ+215Zv6fxcxMpXIH9gN6gZYMFAi9
kq9qRIDTahE8LeUfyWjTOg+t2tQuuTrNej4ETDf2rRrEzGt4McT4X7XuhQN1ku8b
NvfR0WBULIbMN1pVJBd96AThLS7wiPhSChyw51s13R2eFtDPMtYeLJYc+zoonhCI
S7mkR5BUhXdIDpKj8IwO8FTxw/0CjI8lDn7i4S5qJzsPlriMu0Sl9GNjPHCC8yjo
XQ9JP0hGvo2p2DTpojWvc6xWe9UJnv8gys382ZfYYWNVPlu1t8K+M2xyym0VQOcU
zTwkMIZlH/bkD8NcPjXDNO47WNden5/Fbr+HoZBnkEZGdnLfSVj3VJenxjAGX69o
wfsoc/BUOgXoqzX+t3dbmvHI+4C+29Au+HivaInT/kUt6lKZbrsKmNoMU/hoD5RV
XbdCKZmMt3wJSpiGxXZvMQzSDzWsbFkG9CXtot0bSlaghN76s6nla3qBNcOnNuEF
rLaM8vULcbkhwGjWHcVPFpRV70EK3bufn0yGfh5flHWAmf0Wo0/LgIvut3Oe9iV4
K4evjEvhCpj8bs+sI3b6FFaHbC8PVVk/7Xtb59/fh688Q5/leSic9zQV5yEC0e/D
yNpsWhmIL3IxDvXZSRyI426JARpL1eNW//hMaeI4hWbo/MOEqNBXc+d/YBpCeJHT
EIJXiBdr+jd3UEwtegxBh29/GKmwc3pFK9q4Qm3UmOzxNYB62rE1sDswIEINubKX
GYWVs4MPSU6Te9aRar5TnXaSnNuoNNrdPxke7V4VyDZadzG7VP7Af7uK43fhEyak
FQLVqkFKpFGSBB72VOeCIO1Amiw5PcYm0jMz78Rn/NDlz2YBUJ1cNBSev65hwc6+
fOjo8TpseloIqZxLsFtYMGnmsyzUvZGFpQyM2iCc9UQLORQS761solIcaOF/+pyZ
UhVkZdySp4OOuYJ/lqJbaOKCDVV+gj2toDt1XnXTRXfmjR5OtkK3wOqn1TGd7OL7
qSp6t4e7gG1wN5YhWDsfEBvLJqeGfkw+DDTutdDE3MST1wt+20GdYYVLSqUgLfEx
qnxAn2XXpodplSKOgTKaldKXMjsBcLfpSoM0SQiPb7UButcmRpiHgcE/1bki+qv9
V3iYIYAiXtUdUC+3SrDDvFM0H3EfokAPz2JLW4NHkALTYdbXJ417iqrvr1sif7F6
SB2JIthqY9KNy6ujKlooAjpI65DX4Q0e/Fc79clPZd9XRTej0TVZCmqqz3yOymaB
7VFACrsMB8s2T7PQh5xGsDmcqQCVllNbwQDLNRrz3p591lU4Z5vC21YWyG9n1VxS
Xe1r6pOzNerQ/tJVVXkadU/w6M/HgCMRVn7sR5vVTA5imN628rT3p2nWbUrcvkMT
FMyTMbVeROQSG7qTaDX5qzaMwe21oh0i1FgF2LY9S0oOu0BZ2550UAm0Iqx2vTyM
RtL3tAIgf08M4ulEUbemDJXWuLO4KFcHDKtq2pCtfD298Po+ARfbCgiCk3ZxfgCV
h9LRwI2OXF+z6n+5YzpGi48DW/WrbsVZUKsFFx73Y9iRLQ+WHDl0wAOjhBOo2/Rj
u/YUJsPhfEVdGYpTqdjscUxkCkbTYHQi4nYQvr1qVUA4KPDtSOxS1VdirO3AWHWj
CuJp7hF5YOqEYjXcCqEslo5hwrDME7H64ZHHsh3OQ7xGYaz6bT3ZF4W+a71njsFa
Z+BwrMgY0sgB8H9mFqeCcNbkvrA02us3z8iuNg9P6NBQaD5INAzEAJcfZkENetlm
qU401BsOB+vFqREJObkqAxG+7hR4rxFIlgeC0KC3g2ZrBBLA84a9ExSzOmeEeL04
TsiNZsTOIRiH8UZdlv8TAmTPe6v/sE1x/F++lXlz8LyCQxgag8B50UlyZJT5D2+Y
0PHRUxN8GzXT9AOLlZG8iHhevY5D7IUo40jKjn7vqe22IJHyI7uphM2krXf2Uqjn
gr5JijAK6GhmdEnvrP8bzDI9zeJf2FuCnPGAsvks0urhcpwMQ84+ZKWeZThpQmby
OV+QWLcPBk2gfdVAr55YankbfyDb2tSOFuoNKLh5NTWizfJxnRYKB8k8eGl793IV
8ZSf7ivFTNGPwBGZVkiwvgePq87TrpALa4NgdHnw4fR3xqsZXI64q6hJ4vjs/xwJ
thjKj9P+C76ehKcM3T1kggTi2v0Wd+J39BODUvuf7b+zpfNBPutRf3mV98iWqqFb
XVeLs5pyoz+O4oYB49yt8YCqCDTRDIO3XXgMZbg6bhnA7NBtkqqEI+sQagoP/tCt
/A4k17sH4yawKAmdYqQwJR7ZsIMbyuX96c97ixwA21e5fdaicPkFouO/s7g2cL2X
ya9RwMewt2OgW6ROGAZr2FQY0TzbAxzrxi8Y1HllhCigV010CbIqR7eF3MpTfU8G
hOeD4cdxK2li9d9/o2GCiYry6u3VvOJmY9/c6ioF7zWrBJ+s/3Y3a2bC8DWsCfyw
bS+ST+xLiA5/dFUAyOVxhNnKHI8sYM8865yOTFcVXS9w3df1WDYXTZpxIL9XA93V
RCIW62K5S4swmtP86iVCJ3DIeY0cicehsS3xHkT003w0aVsHtZa+l0hiywvq1sYF
kp5RsEExXiSFavUptOfwNwvzxmtOuWEwmX7TtNbF8hNVVc99nMimsq3vzfJ/3cT1
zSf1Zt4XnF32csA/mQkYTpna5sOQsr+34uqvnp4sKPSXa2FbjU5Tpp2OKAmRM4ou
QcThjn3tJOmxKhsqb6rACsi9NV/tVGoIRfcqiKU/fTffWfhZRU0xvCQfV+g73wNb
w4LMVgVJno+c4M2yGsPUpn6OQS8ZaWdksDBjS+g1yhxdpNbwy8RfFzM6EkW4tKHy
lJ/8t1x1j2jP5SRkTdDWstgNQuvQgEoEHRERfwAPnN5dtQDnzZRQYdITcWRZEpVD
DTEG0MtCPRxQLdh5r8qlIHpu6VC0+h38Cfems5gGgd+s4nBLMvBY1GkzdFQ20bPM
ZB6Ba5IKdi2biCNB69Tpn01ngfAFZxnoHNFi2rgWFNj42O5bjU2CiE81VfXS59hR
JlhQ3jrc45E4WkH1E3jEhfizyiPTcFb7oniCttYKPsB5d4sdJHJjKN+WDGpfWxl9
2CF15AwRR5yiCcpp2myrapL0XMZN4qek4guWyhk99sMYfLo20c5CLG9HwvL59uyW
O4rGpyxWU2PHpqfUI2k8nMVIOF+8D6gbm2n+v/yI/SXsNC489Lo/PHddMeYjcb3I
LKO3d/9HNScRalcS4M3onzxIzZvwI2NE2DoYJ/YhuXt70oKugI7x55T9CuIjWlmx
FVafLzMAnO4CGjlmkZsU5CWdmd6eOzD/nLFpan7DhlHLJG9KyIGBhOoUIbNpNlYn
rxEb6yCr0tc5yVe/I34Cx58uF5r7R0/XG8XNGy3hp0Ny4rM/8Sc08H95YWi4McBa
GMBP1xjhU0tQc5nLgQJ3DuD/O8LWaj/J8MGNklbmse3Bom/Ejw4Vdt9RyTmXNkoR
zwm1oSZVdaH2ZUDJVS0yzWf0+KEqvgXKDZM8CLXSv5rpSc8OymcHC3lPtUyz3qTT
MQmIay4E7DFoJ+GSdrHU1BtSRXKH4IasZrYBPyTAKZXaiU+IbJ2kl45DH9j80UpK
R8s2iGZ/C5M5GK0QkO+RtU9Jdm0CGvqJkpdSYTBMC7tDZz00J5OO5J4GqL/MfAj9
32elNBqlFflFXoSDgG8XvV2KoYWWfBievuJ2DQnT6zI5d8GInHJ+yWGqtJataqGx
Ul2rMAGuI5uE5YykUArLmL2Dhr3hBgn5Rq5W0xtTawrgdVnalKGZSNhZYGaAfyax
UYIK6miLWxY5NYMwZ5dt7OhgM1f+Sl7lr90/hEZJ0BQbK/kA8KfLiCaEMU6piMjO
FjPB+n7/JFRgX2xYkF0J4X/0GZ5CBkENgTGSVskErD1FbeCOeXcGTgtXiqWhUkJu
vl7a53DOQA0pnnQwmo3RYBYvxtozR3YarXsTq7CAoqITuX10tpDz/6lXGvIgPEnz
WyqNOm696LKJKjvWN9tquCm3v+tda9RTo1ELn8x6NjIbRoal712clhW3RjIrGn8p
2tFqIBbcVFULM9yHUzB5a+nQGBCYeuQQGUyt49iXKdHOt/sw3GVw0qIfPasz64LS
wkiEhd62030jQIHDvzavXi1G031oDnLbsteZH6uu/Kh8i6n8Hlcx65vXe9HT7mJI
xsKglfDsQgO8GJk7uPLrlUMnx4eZQ4pRcafRg9F2sAGWxFmK/J2L73QSW+g8UjFo
zKs8bO4G7Dr2M2blLVH/I502FzXFdTUf1l0FurBs4Mfe0brHqV/fw7ZWfqVxLan4
iO2d8FSsBrZkxyKGc5Uk7AmxDNLFfaci6xsjRevuPVHloh6wGnf4aIrh5kLTFCgl
wp+rDVuERfoOd5HYGwLbE2NzuGY74WtqoKWV65OALEEuyFMvh5r8vgpzz3eMnWPo
NmbsXF789ZtP6KEYkf9dzSbLtRtve1lWdAjzFJeTuT3U8tRRzf9o9vS28v1Mdazp
zkJDvOqpjI2WwqcEj7QZ/vUQ7APUWW7wh+gk0tAizetri2al3zImut6Z8yZcN+R6
8yjVl+wvetNZctIn9jyT6dlfPw9dAZDwO3/NBdNlJbGKvTqD6TlGg37uOh2DZMfj
r5zLXb/RIPG/OFmnuka6NY+le+DydCfPoaoqR6mFitoxosADUy5uEyueopYAe5iP
fg4diEw/Q7UyDnzxcgHKJtaIbitFiiapv7BqLgj3ROY2ImxgGBZJ71Ykvspdturn
kxAatCcNJ/dvbMSk3hUcU1zqGsNk0Wbfqv0N1S1O1w73Dg9zdkes0OSrrekkAS7W
yEoSorTNmZSyORfYYcJhJLmousADzyrD7nRXQVy6jgAQJ9ODytKQakf7WZtwq22L
L7nDwtYZrSlHffp7fEwAnY2UtvAKE7yov6f8VN9RQnb3ShSwTHkC2AvsZs0dz5lp
THqM/tf+5NZKN5kuyeUMjlfc/RUZQeDzcPHldg1r0KwE9v4ydqw3gNPBf/b8iq7E
GnOhp3JZVDimwLsSU9gkyEhikQ9jn5Ue0GQRfiDHHgl0mlrIxopq5j3Gi9nc4YWk
Nr7kxsY9x6yh2EPY9oR3+lIGY+IZKqbXgBgfB4fQp83z9Hjt+h4fhkV8ePqjOEJy
muaDSKJIR/bGOF+9c87USKzBJ/+fKHpH60emfavEa6wesH4TV9Ha+WA6rxDRwo6z
8O4HIs4CKjmz5dQz9y4InhPG/3L9J00p6rvf96Ss5Iy5V9VD41TiOHpLyKVxzxow
+b6HlCH+0jIY3WgpRw53MfYaFD5KftMZErAwrt6LcuQAcVH2ovmFM8wm9QxAutFo
BJFjJKsp8+6uDrpccWlvT6LE9EsFB21lZeEyBijpkyOo/jZl/H/GLQlFp4IgSNNe
TAREEFTdVQB6jU5pUJMLhEtF5Z1KNClG6y44x1U3GxfYC0qq/atLu6y/9h/gSQpP
Z3RnkerDA3NOOj8dYBMp3XKkFNsSaZ3YqBByy2SavH8YqG5WlUD3VgRsN0XpIcXg
uaYLmH9/MUBTsEkDO6TITaa/8DLzeghOiPB4fXoZkSz9ojfgwbkSShc102YyRg1p
quXio8iasiB2a0eAbjvWW2NHsYu5f3ryo/zkamipgd2ZopzDNj96/uWVcqynIeBE
7s9i/2n2U9KJMAbPYNKKYB7sJwYYuW2+zyPZrwk5YnWGbDprmVXRyAlxEjl2qSq1
2y59FE6nO9HYTKgo3q+VFX4ByR6WjrV/Imu5rqJXoqzF0f1qzZL84Arqen59dc+C
0ziYDG2EaH2fD6/WoG6iNTBSVHcIdxPl4XujXYdp3yTlWUdpN7Evs/7z4gm6yJHI
O8AdkIbeok/biuw7nU3kzuPVNLpHnzI2aKF/fV6wigJ2KYLqslyWORhwwgMQ0qEZ
7DICajvNwpTs4eUpIYT+vMgKSI5qRnYC9IiG9beb4c4WfkgSlmRJa2TSTULUFEcP
5mEj1BmHFBU/4VfICgDjX4i9L4kgx9Gp4DHxMVKevnqDj5FE8JqJXYIYFmBGaZkk
piApQUAo/RQdkB5Ff5Hr03UMrh4zdQ/l/3pAt4zBBbuLYihOMxeu5Koi4tF8KEJs
op5rD0LvXeQveMRsyzsYK205hspd/7pOkcNnGxPbc4W+eASg3xjfy+FXAToaS7Pj
Xik4jeEjpNH+gGw4WljEA2EwNn2ny9FYfJlvE/UTq4I8aP3nMFNPTrnjqLh+UELZ
LWjPRQaF0FSi/o3k4rY4n/xNaXz/rsVAx6ZnjRXX4kptknNY1SL1Di4PEG+V3LBc
9lqNdzJz+VHmUkjTAwy5IUXn+iqR1B6WZw4mMOqTZEGaB4eHZHbWPS8b/t625SCb
E4JgFQaAk76IlymEz1dohJNQVL7W5N30gz+lTdBYNqi8F6Sww3iiKTP+8uVOXXYe
meZw0EaY5Qyr72Tm7xHcAo3HFIvq6LnMwCCAokEN0jfJjQ95Gs4piFhuJY3hHXMo
jwIOpi0pALt5nXAd6DlOeA+uxs7gSS1WP791BAmKZTS73w3qaqLyVSlFZTIrr9wd
4b4Rn9P61YwMxSuXsyO8rezRExifyV9mmFClRLBGc3RWL0m/Rpj6ush+27zE2jsC
J5jBq+YZRjx8tszaVsScWjO6khZ15DR8Nez5LhQVJTbkbBmlTz/r9vUz3LK9FPIy
5Xypnfdy5wRFk0OrTE/hD4On4qqj8hzz//0klllMItBcxwYoGSzjtwM9Zk8NLscU
xpBAncgKEhxGaEWT+qz9YM/3+DGwMiB3XkHvp8ycvSHu4h55+l27k6E377++xd0W
jHvvAfzINZjkVwEcsksbZtN1W0jt2BJEoaD5PsromaTvBmqFNM0pMXivEuCJ7dC9
GwovNVuK+kZMW8ZR+OKaZKiFRpKYQFqAdduXqsD7Kgl7lwj844QwByVhQonfRY1W
Ik0RV9b6NwoQL376+Lzrn3fI7NjPiQBq2E0VGFuW4gWvYYOdv50FIyiP1RslXTNY
mtgmXKeh8HvWyJmHdhueYWnl3Xxzt7HY/g2NewJ2D0GF58Ncw2+NCKmem4NB38Va
iiMtNcerPUlV831LfpCUEg9sK0cKENsMzqrCTl4XbI5uX3/ET0Mk3wBjKfp1sDUH
NW0S3JB7c11FR/VbxQttNiVZwRG5v3J//uSM8lChMGmUoALZ7+J1u5aZz2/G6Fkf
Tmq7GOf2Zkv1XtmocrlFGLU2MptDMb5OSOZUgIYOJBtOUFOwwqg1U99MMH2KXO99
dfGuLXDpUg2MeLi8hGe5Cr4oyT/8d1mqiq8ND7tQ1kanARBspbz+NlNbRVosROpm
15enqj+qkU8mJMz4JY+N6CxH/h6ctJ0kLgFjklQMcqWQZXfw26GZcOedadhyO9qB
hu5iC3g8Pu4Q6474/qL1BJ+8y1pdQFrcWFUFWcQFIL9XUhlsgvCNmUcf76B54McI
BaFCl1Jhl8Gg/AW7l4GeyzKJED1+OAfWYND5/P1OgHQzKwCpyIhw1+n2XPkEh6lC
exKSnwYA0uBsdV6zbYOQU8BvrJftaWwr3xv9a1chQjCObCWlJrD4mwiDInlf4XWH
g9u6Eqhs4SHRm+hMQotEH8Xz5r7AzA2pksSDzeGxp0PUh/lQKYhqt6DVq78NVHOk
JkRP1Inc0U/SzLdhllvNVtrKRqXnc/LpAzpNPe6u1syGv7Hjf44tMv4BewhxVdcl
g5r1J/opsHSyA+zRrUfN1mSqxB07RKDcQJSYVv6lFMIS0NbvCSHLQg/BzZMijb1o
tLRb8UD8N75JOC2NCBICe6VfHf/k2ZsTLjlQSY785iZAdndm0NWS9J8cGkWkkCUp
Kqsn/67AVafD1G2HdHH7eZYXmDrF3sPH0pZNjLa5+BiVFdY3dWShgy4qs3j2fibA
BxkZm98HXthumaLdZh51v8inmDbQ0A9p/m+WS99CiQQeGu9m6LVi1gFpPuIXZtmL
Xnjsz+oa4vShchTUL30euJEINIRu5nfeaKLcDiJGcdGztaaUlchK1jFQZVtTdfRI
Opf8xhISjdBQQHnGyODjMlizG4Xj3ZjqZONCnRWpqJ319LzlKDRDQUMA5ZxFQTnk
a729vfwvucHjt0Uyf5m0Jb6fzMzBGHqrZhk45PY+p06UjnuLi0KpMtaIRgF1BhcY
YN3YsDmJLcuDcSiWQtGiwZwSVUGw9AeLNrWlH9ltFyu6Rn0ZvEPG90te56FU33Y1
uSfxHVk/UwIzRXcJJVnkeeuxfyOBUvJ0y78vOOJMmoME7DJSrtMLmHSdWPdhlabw
KJ4og6DnrhCLaQykdmgSpEOGtlgIa69OBUHU7/Mr/0/oFly/0/StWLOS/9D9tv+0
9j8yUY96WVcZpq/h76AVbGMCwHn/YiDHwS4dvZOZLYOUcLCYnOVjR46MQ4oZPuFC
Noy/JRC1lgNVjqX2oDkJY2urLxBM0BTR3RBhM8duNmEXA0BZ4hHBYo87MJ9XlCI5
t5lhQOr0jFTM74R9iJGL82d1sWStUK+WknVzWQ1Jugv/kiUD5bYVZ1jkQ3zxqxaW
Dly8mZPERoMqsd99teZdx/QAyVh1WBGpiMda1v0HnQIr2/9bZbetdYDXiJUttLio
/3XURZV5NRaC+63iDahZfm9fdde/ScGgFMRwmwf09JM85tcOKLQ8PxPdKrRZk2NR
H3oBGX0AhWqmzfK7LCyMx8qT2E2XTWtI9YhGXl/V7Qvr7oI5r9uQAt9rLms3huEt
6d33YXldO5/sX59C0LXq1MZ1dyOnHKUxF5v2WaN6+S8BbcqtXL6Cp6MO2cEywH2p
vV3OOcFCUhekpn7p1ViQKwLsVi5Xfhjzcf4Wrwx4O91zHr3dKuzxLchwooucJAu0
JpJTK96oIcEiq/URlAtS5LhgZhZ8wWxjIctx4guIYmKYfDaNnE//VbySDHrGb49G
zD3HaD1pnP0dIvtwZTFiubcdSWS2OkR5G9GaTxTkjaPT9lkaByHQHognYmsPVnvT
kNaGGiqpclDkfMP3F4OgU8JLQhE1GFIiCkNBzq4wDB6D89Kr+gUEyMmvgAigS0LJ
x6VVpsRWOBif114dNIGm43WMD8jmblm0hJbl3TozY8hD50EDFiGypPs/HVE+M8dI
Q/XZfRnZcZSs4L8KMQyKyqRC+kwf5X82bsW0H4qboHG4ZyPeVGZTTvFquqJFaSXg
+CaAaINnIeBkSZH2RnSOTCrGPPLbXgeMO86xTQcvfd8SnJWjKkTHuepYjrO0ePQL
v4K3ebqdN3a47/e5DaYJcoA7bzPr8yt+nt3vGcDQhsMNxUpwqm3+0HZXf7d82t00
PXEd5LhbWbH12ukLdshvN3oJjwgM2+mbf7GMF2K9wedN324QHLdvIDoZJo0x/Fx/
HIsCs/bAmVmVuZf+Ed7MmpJGEv7SPsNHRn602QlcwoXTNnVNTrXRZfSTV9udssXl
T1u45UEE3tZm6jjRjPCQMv+yVFF53GzUMtCo8nkoFbz0F4meHzLBAaE9PvFrNQ7D
w3B0JU0xTNnvhyKNdltBR9JMX3tvZv0R5O70+RoAz9tNimQxqgptFmQN9OX58bZY
Q4UbOa2ZbQvzUVdzoFEYu32VjPCAA9eGINAJ4c1G9LuIEJNjIfc8tc6OVPEhE0M8
a6CkqP0jGVdC7XXo0AL/tSyTryEgp0CpBdXOSUSASxgCcIS0ZqlAxMjzZSEKEg8g
r8SUZOgCfWvgQugKV+yHCdTlTrNTQHViGtO7ArYrfsmh54xxrIO6JCjieLsosVyd
Q9vwrUN+T3BKhWsNFeXiIi6nfm0ZbJE7OwCplZL79rjFqLn3ftiPddZbc69ZY8h0
QqQpvCt3+fGqNcZcU13DyeywEgKkKffUBw6PLwWLNov097zf7bljRxFN8xnLoxhj
OivYhH0wrF6ShMb4XOxxXscJMylFUqLGQfV17RlRstNGdMQZCbEjYSquOr9ZSPlh
22BeTpsma7WZwkwYlfzwA25oUWa7PIWGT2ok/43Pxrtsfvdk8M58HZ7zZSxgzsFm
Rx58mFpzFx+Nzm1gpttQaJnZbT+b0EbF37A2GX8n5+xDiCWxy4dWS3QWg1zCilA7
dgXcNr2DnA9qrPhCybe4hVhwT+Np1XzMMKbVxiMZN352Zd7tDNS3QhnBwc8DrLQL
+7rFFWJHkpbiVm5R7UOYONLLRTN/H4HdCq2Fz83qYd+gNC4KJVirgqAiCBB5BpIE
0n8uXHYsgHopLdpcOo3tWKX+0wX1iQ08Wiq3DSxs++Ju+JayGPc/8tljii+w33MF
rMOU4uqUXFO/KwAA6eCzZahjEWIiDKZzpfaUmM/JF7bGC6QB0BNFpUEmgd7MiZwU
v8hikaBhk1FN3jazxUR9pyUjs7ULlad0yRXkcIkQknAd9eypQItJLLx6mGucL6QF
0ifngb++g8jN/WZAES8QlMrddz7VGccgyTmVqBHbSeclJs5nzDsekokZQY2t+OAT
EinRmUxaquotMMnPWcXfyWBaDlgnHkFEcjLkLsa41DPfIZHygLAjG3vCyGkQZqih
MJN+yMgJqtgbXpEE1W7dDbGIEFw3cYqAnG56V+TPfu7pYCSBaabFA9nJcZMMCvqg
71SR12NL+58EbHI24L+pyPBIh0eq2Bb5Hui7DrypTJ/hzYdZmE12ZuacvuTUDlrH
QLBNVRjfkREQbXj4F1VrV0+MUsmLOjShYe12xtiMnSvqQPxvDQuAwvEVFBAvdq+u
QvKh+7AtmhJS6N+mDfelElqlDygWIpKb5NP+DEArXOiWhUV7qj7cD406y2k6CIr9
WIVg97kRYe/jh9zfcDFEnq27dgfCed+C1GgeBfL4gXY0s/NK60EJZ+iptUgJc/0q
d9Dk8YuRwYV/3xsKlsLo0eol5Y4r7sybr4hMKRvhDZvYgbnM644zo1BhsiaYS75u
fLknd4FYEuFRDryBfbS+IxYE184AuuTriYebT7FlncPIDS2xYEQZuPoy/mzGWGe6
F+YxnBNrYh3pUfRTfYKtTnHwZS7jwKlArGDyvBcleTGKz21ibTdpvHC2dQiM/0Vt
uGCnjIiPAwNsHM1ClkwmUU65bbF+6Lxs4PWZCLQGSc8cXqbMZQu8PgZc+63FIOk+
c0vkr4b2tdGpiRqWgqAQIEKLBpRugWe69hm36/IJ7k1J7x4EQFWTFOjg4HFgZxMy
//qhQXqiXyGfxV/g9WnjCY1LVqZF+BirPLh8Vfkolcoz6g730skxIcdgFqRYOi3E
O0Eou/uwLW4YT7Q8JgG0ZVg0WW9o1naXjRL0OkAwFPw4o4ykawG9RB0iK7ISR6v3
0Y2hcYNtavLTKoF2Zm3Q70BJsYO0WwuVNZWUX3R4dP/RIGlSsMyXIqiPocsOZu+w
L54sE+/DNy/Muw8gkXbRPPTSj9vQwMqOTHfhnmdum1b9Uhnt2q3E0Ojf3WyUU4GX
9vUs0FgJu/9WATzXDuWCRawEpDZCgv6TNfrz/73MzaALGv97w73QmfcWUuaeA1W+
gUrcIga9GcTzAvHT2acXWxdRUBq97Cqd5G5D53toZzZhSjh9BAXp5Az1+F7erD6E
y+koxwG1F6QHsYprFAOfUMGs5qTFifBF4XS0+CEIpdZH7pLoUvOiG3jYYlofwBMZ
T5nom2wKKt8LYM3qUiXBk39xjbIOj/GrXP7t8T3YKy+CCdp29U3b8/SURPoNt6kY
cBpeCqRXSc3P9wczbP5FRExCW7qUF5udgBgMMHeydrlAfOeJn+2klE1TP3r5z/Uu
Le/3qZNLJ/JzU5NPuNNR66AcOs5MRTCu1gma6LRgImnWBGu/hmrKkTu5Qm/hRecZ
EZaPZn7KS3caEKAUNBNF4nUMYrp68DxmjCm6Bq158zndXEmJc0Zz0w8QfmJdjiJa
DYhPrV3sVEdxBlwa85mXLEBxu6S2USdmIraF1TJqrIHc1r2THDABb9N1M7gklhtI
HIBTrHxnV1EgyVXKBkgJ19onLyu7KN1yNE5sh6Fa0VQZb084Tf/XrDliDTeOMFU+
3tuyjhz8HuVtjhYrXz37lyjr0Z0QHzRyugyO3sBsQtoDW79N9j9WsooZToJZ2ZQA
V8ursSJ+QGEAgPzpTLoLQYfExiZau6UsePeTa7KbW+yQTtXCZ4SR/w1IcSdRuzQo
ccfKXyG9ErKwSI9BGHE35ILwkWk5W6MU0335sgtKrfrQy2sGV6V6salsD8Fcox2a
yGWNMvBSxECmoG1+x/qZZgGqll4Zncfl6AS89pMyuXWgPhxlbJn8Jqs/0w0m5PY4
m+2YOFN2BhloRWY5DgltFPENUIDwwhqnxONpKarO3CZ5X/Y4TVg9H9M/W+Zvcqm4
g8vcuWC3dd9pfIaRny69HNPcuvwufceSeHfYTsQCL4yqa5xNZC69/RGc5bPEV/wy
Cas70qjQQ3/Qfmm87RsKsEAIqXiIjHYpOiIMtF8Fm/yt8KT0NXRKsIC0gEVWnDE/
KdtSRGTqY/A3i/Cu+NKJaLw6NSqQ2JT1GoyDcB1whCloerfmsfZf0Ki3m+xGw6iR
5qii8iEbcGUPAcE8szntH3q/+w/870x6Xt2xcvTXhqXNysQqeyjzYE7DJnSrOZ7C
Oa8mczEv7DxGu34Vq5pRfIq4USrv501NABiHd58ebRyjXhGSuLhUacLA6m4eAhXP
ZxkGu07CH3uZAaUX09wDSPrBmYyiE001prO4FiC6pHRAv2jjj35pEfgYBlZuVXBk
W6rFzD9yUtUUIcBSdMyOEDK/bAhMKwbxoCBF2aRivxfP2HxcAuOo3QqnMxL9Khgh
DxPmRDlqvitCOLqK1J0jhyN25ert4wf17vcGvitL4QvKMKbQxCIyi32VNAUcC17R
8H8fJlIQ0i/3Da5aCDndgYoi2d231FmBMDNm6dwPwaoeVmPdZIfN8ASS5H90MLV8
gVq2A13KiNgdgMpcszgeDVodRkufjx0E8LYApGne8xRA7adcEt9+gKqQvKyCBHOs
tQDke2VIRc6KSQu4kOceMl9nxdvllPD97iqiuQw9xgQWOBWKX1BQ9SkMPmfgRHe/
g6HcG0xMzh/bW9YNoe2XAD3AaUYZCuEcq/jNX4qdO3ut4ZlxNCEJ6g4/fIVc1AEs
i9IXH69vvw5pQ7XBFflzraLgh4tMusBBx6+QGa1gEKlHLIq/ivUrGy+31ev3AKfN
aN8f3VMTXMJZ6wSB00+cJnsfUNLMQdo1p0lufMDodgT397ELZSQIQ8/YqTK580tA
5mXBm9ULrFgzJl+fA4Cu2liFdOr1W5N1KfKybIygm6UENQmXHikTbVCfdi2PKH5G
7/xIRY0cfZcr/wHmmiNWRroiT7DdVG2UtJj/qnd8NlrFg00vFdr4LRLZzzB2YFl2
w8DS4hmcVPCzO+YXl0Mi66aQtdxkHq1RAMqF6dUWk16lkf2WLxf1/hI5gF7oNMGz
THClnZkc4tB0Zxvjsv43VHARhRRIH0f2gm7cRVVs/mPfu0Gd+zpMZmaq/Le+VY9S
l/gQ8rOR8bJFfI34TM6ugMp+68m/79LB6qgJxtGZELRiP7QA3mOIYsQy0VfFbJnu
A415jTj1Y8g0LJwUSeKknmUzEXCjV/USle1GrzgKIkliRToKzg88ruJex8jcn90b
BnD1IlavlExPNYNiI0uVCpmRE3PxyLZPwD9ArBnJePvP49z/CvD9dmzhJkazlQrI
es3KH98VqkhY+B82c7CaeqZo/NMf0ooCd3Dyig4nCHZh+glx2zGLGjU6YhmxCRoN
9xCL+W39omQTC32y441+1l/YpVK0G2UVv9N+69OHJR81R3oaU9XJcN/f8ACxwSse
hk9G6AaWmc+4rr5b0nO1BUKv9FOv4nRPQBvj9sC0a+OTpkKlg+Na6BAitvbBmj+v
pmrur5dFqILM2BjX4xFOmdOY5XSLe7aWLZH2gi14+piGacvtiofOUHVTkSVEZMwN
U1bhhwznla+cSJ4V1RSjZB35XAphKDRlDrdyG0AVWqf/3eL/7A1cdk7bwE/AHGvy
oAVisw4OIGCs30oDShzlTu3eQaZld4r/oI1+X8o6pitqllw87FT5I9QAjIZ5YrD0
2SNLxVpMiSrwntKZpwH3JBCnhPHRz4ACIUElSOrAv9o/Z+n90mJOx1cOkmqmoxOM
rMHlxDOHgndmwRdjpEzKe3YdsOeqBGV+Fl5d0sgmfMOOfSaIDnHutMZDpSFeNrlI
RCQqWO1KWlmrUmCDJwWnesHkQOm+NLaseT7lZ3cRZrK0lE7H0WXNuxp4refJ0Hrd
XDnWBLvkzq2WAI0/dMGFXzSq+1AE9tiUwiOlr+8HPCOcIGihrKnP0aXXwa615v1i
fCaRadJRdqZFvCZ8AwFNwqQUfdq6eXYpvqp5HDyqjasZy5HChbu1mWRQrMzbgqxT
ELJm63828rEGYelg3kRSUOQqngtYXmdNh8as00oxLYsiFzYSWRZ5Uc7VcnHWWAzj
kntTb9ZGmg8eoCP4ylYIM5P45mXxzL2LJ96kIHqYINE5M+onCGujwCZ0JPZQk6f/
fhtuuLwoG3Wo0dSb7mQ+DYNjHaWWNHS9u7THMWZ+IoZR4TRT3IVB9jmFmyiRD39S
Fot80KW4zh85TTY/lq4XaPA4PwrnzL7dam8bg+iJh8hDbH1ZAvBuuY+goZgCYaN2
QF54+1jEZ8ids2jKOsq74fkjyD4hyiibwenALGxCd2CMjszLhS22+RFs5Ehoklps
1n0V+jQ31BwyI9iaTptINH8e6DATIZ0s6Nhb//8TINJOg4QcnFUJuuU+ypSjWINB
BjS6j/Xj+jgJlRlPfAEOPnKCq5SinN98AtaXXG7I88TG8v4M2PdNfI2lubyye7by
VlvTP1MebwHJggNwASh29Z0O7tcWkQCp0TNPVuvftorxT2KdgMOC9CVfUmc+RACP
HtolqJ9h/imfAPC6TOYhiTgbn4DIWcbN/un0qZPQMiq+713jk+eDCCrfwormaW5v
58+OI7gb5ADV7/f0AG3lBcx5Kf7AhqeuCbPe1c6ud9qnfXiBoMbGz1za99lD4+9x
aYGC7BbD/GpZ6OWZOHTBbcLU1Hp0D7nPY68rMiN8mBRCchvNIVLWuc1+UF+1g4T+
YBqMzkWXSiNiJfRDjg50T5cST4qN3NsW70+uOHWbx4Ib5WGFDpyaaJSAk2Cq6RMU
7I1TTf8s+bdD9Mcpj/tY1CjpYv70X49uzqxLYhXb2myL1NqWMh7Zk6d5w5zrvwNj
aAL7/dsFzyNzDDpAPvdvLZcqLMUzLOQpJndxOWqL7mHQP2HL8F2APqcb/yy5mqCY
+naoOJ3IJoK1MQCAQ6wzsp0co19ZWoNYG9WdmARqdOk5TE+9me5sPh5KIsjSUgz3
aaGSxzb6AjsL+J2cSZvL7Z0XyNUokYQab0ru5BOP1Cwps6s97GonMJgljEh6npe8
OIoLwCPGEknwBVm5xhxQrQaQIto2m92XhEX7tYaiy1BC1qYGzaVzuWRskdo+VkQl
IyhodUg5YPAEkG6jPMbKD9pWV04frlxnM3/TDTIGkrhSAmmugpnDt3/jhVMN8PW8
rIW6I7IUKbdNtVbCvGLvP54gANZtIunRX8zIbFFOk3yyGcPJEDhgKbuCkEeSHwMZ
v1jmlJGfUj1QaycQIzkbvKaEQpc5KKxzZrAxXG3Rtnc1QHOs81EjIeVaPd14WXcC
djVn3KuMK8qadtyd9b89/virF7GUjOy6RmXjvAFhqR1j41bidw35lsZeGNxEuYH8
j88C3oJoPW3CgpMhiQVMSyl8QCdiDW7e5TuI++RkbnHTxIspxNKOf0X68/U4Z8xf
zkdJdk9jAJAZNI9JAwJrmLB37tNE7kZJbZC2E9TH56wScAK1v7Pk+iGAwoYvMDkn
Gl1kTkEcGhoRg2Yw3QdWlQzWoQWZZdAcy3yEJ1aKi4ZjOeSIT48S+4oMwDLn2jwm
jwlSsLZE1sZeSxAvIhrLMWVPdckogCq7vyo/+meK324dXQXFxpvp3QDFlzly1PMQ
QSxk56UJTkVaWCC59t+g3zLiYfyuOJsn5WVxU6g+qDLjZLQjR/MjI7/0sC7BZayx
BLi0RCuOEpXa1SGFHiOfYUeyPTk8bz6ZN8rF5/eBzOdy7VHSxXEAUc4X8uCMCfW2
HU860X89mhWDu4tD1HTTBGVnUZbfZsYPpVZ0hXciW9/8YTpKMeEyWTt4wVAgSpAr
TGpwCQIdW/iN8Qp/2vpmuMMmvayaJbi2X9m5dRAvD92nxQ4maiozsj5nYZmr7KPT
NVJOabmXkcrhoZ3GzxkQ9is1TugIpztgjIdlGyLJySsjI2kPZ7JuLweAzHBrOhd1
qABhK7aDPZJ9LW/YrvpcRFiKROsrIjIjmImsP4DsckJG5VtV3dVTJeOKmWdK5u7U
4aWt27BI38+YyG0IyXIGfaEZtDMg9X3b3r7A0wJ30nI6kKtrCB0yGzfUVaQO09+m
KOo2XWbPx9KO6gtPMRciivlv7H84p79jPYWMGBqOXdnMQkaMyy1R25zh7hFV8uxm
ddp3RyDZ2faSc3yIQ3kST1zRYBunjKP7ymW0F0rmcSTHOxLhfpXbVisgZJ5ICAvj
39luzOOtBVDmJD69p8cAZ80w6wl6ZhbGpAgHOQZbokueR33kbFhdVaRfkYFiOJYy
jqnYiwb1VWXD/SU1NeYx9CxhjTjhsModqWwy5fSOqXitPQL19YW/+SyPTZGURAbl
OPiWlRYLTilciUULpopisBXNxKymJoeBIWMX2tKNIXlSE/oHPBWP/imDymaSpd+t
c7rwiRPRSP2MkhoOCMaHIJN4PAipycpJD27ENDQW0cS1Nx/hzj/CSbhxRJbrccg5
xNev7cJ6G1Xkn9qSxk2lM0CLDu0daKzf3CkrziWzajqP2jdYum+QPvCGrvKQo4vh
lqDYyi6m0gi8V6vkPNB6D1Q1ElHXjvTtuXyMOYXsKy0CM1NOMQd5t2D9ouQaX/Kd
EVeQdF+2eBe2qn2u6fn1OncPDZZLctVsBLACTyhFnmuO3dsujd76A8jhULPC4aLL
xMXqS/OmGclD8XY8CFXs8nLS4K79/yxFmHJH0H9DdZ9mrBaJThTZqNUGd2MaCoO9
cNRcMVumq+OHUIvJxJ4Ji39eFNfgXoF1CWGoT05M5jVKsJfTyvK77O4gTFjgGIpJ
qB1P74XKb95Ut6hXCBkIPkCO3rT5rdcsc591G7L30HLJUaCqGngkp46B5r3/rwe3
eTxft/K1YOQFjnUs3mga6AWtlcjjeXH5qP0tqdTWjlOkdY04nMQWc2lKGCp14QMt
3tVm2B+AvM5PP1kEn/kcjWMKNBp7Y/6xn/rnUJ9RH9AruyAvbeYwhAA1SyyQAcwM
FQSH6Oj/HABuw2TsFMCbvQh6+un8bljKqxfVQCvEQI9AdlYTS30ZyvCR/b1EBidZ
i+wOeite0bycqYrMt/O13AnXtEqsWxG2HUmUbaxmAs0ZBlBCgsr5BoMm84POVqfs
Fq8UmIuWrjZbu2FzCNXHgkZYoPHGBW0DSjeFkeZhMdlog4cpDcbletSvK+EXta+x
BCohhkJNAeEPl1r2rYHIFrBXEsDbmlTeXQOumj3Cy7gNttJTSnLGT8BN03Fbo1pr
vOX4LwfYzXGHcOnUpxcFMAb2Nt1NzgQ79vo6r/o7qHsM6BvyZtuCoAJfgJpsoso1
vhrhgwghrjIe4c2YJoPjcajXop3D5p0maTmb/4A9dRr9fSyOzCD2QZqQF8Mn9rB1
8pNRUVILuucIpst3l+SoUDKAkbbzXkD9u+1Pq37aQH0+I7yVBFIdbcguTO6D6OUT
Jw2jJRec8tiU9Px8sdfF7OMrOl/XZ+o6tN6Yvkx2A7pifs3TXj79zDfbz612sweV
HT3yKD4/5IBO8YAcsGvMy05in6cVhjJg3jEvEPNTmQfWRsQG/f4h1HeBCr2XIQV8
Btt6VjBv0m50LaNvF2YjbEVS4K7Lz9jUIt42EIleYRlZIHuiuXbg4L08Ll98S5p9
NScNIQaTjliZe6cFilFIkGt0Mh876wXuxFq0kwGpEofMGWJ/llsG/FINdbsZZege
XPozXpO/aGVqvRPM5VFIxwRJRjemxCIRH5TrO1RQfsvGoTBWQRkJa2PmWS3PSaEa
rweJEkP3TGtDWqIvpKnBxymlsYuRQy1VtrSFsyaa879ESl0xLwqnicelhasxGsi0
rlyIRfxtcAJ/oMuqhbEXBigVRYdwHxwmUumIHfQEv9IHZQcZ0/sQUKGy3xfCCrIE
GuG9mSlgy8l5sTSdLD75RP54reyFWU7imwKYhve1k0jvuuGkefYE1wFRE4fKlc8F
5DecIeLqyFaHQCj1TOsif19yjdzpkUl++cYRLcAuQLtPj2KSPcqDUQ65dKCLPpwo
0H6wFDbzbHhsWyhMe1yPj+BCVa0z/kWzofO8C0i/Y8VHDSmg7XynQaXY68o/byR9
epDD0vTNyR0zjEeXwgSfSy4jdUIMQr4ohIYXcfioax59HFK1FsyXJSkzXvk5pZWD
D3zTOKe6X865tCj+DiNdcvE3fpVMceOArYbwDUzZtn9vkZXBt2ca52lKAbAJqLIH
gXkMizwJQ67ZlJCcIitb1ujtypPcnrEwTDHiE0w5Yc5E4uBeIKmV2ru1T7dDSGWY
kp7/4pDovInzDsN+7lO1PzEUsxdeoDnei0H1jT6pxzxJ4vwZAUnGTfjAensjGRl1
U7RWOXsU2E3nxMIUNu7dX/YmvYpILQQ9rRPRodbMeVcmeV2R69AEo7Ot64Q3VLfC
JrE/4+y3ua6UP0AqKHHDfdiElS/Rubr4RDdf2gZrhYBCSdRRmHTkeanC3fC+2dAq
RlAd1EyoccoYHNQOTO3+McE4KlFn5gvLy5xos9StpV9IhpsER49rJ5Q1GYVnldJu
44/dCzpmirRBv3yRly+T7nhszWPA/pCo/0m4QGhKDdiss5DJckLAL3pEIG/WVR+8
n2GolYB7P9KBdFN+IGMDG4pbrEZ/VEbxLg//d/W0eYUhdyZzCz/y1fEHZ5IixTV7
qQmyRLSgB0HKlKn6qyNdJY8JCF6W66WxBuEU4GFXTGSFH087LODK3sBndCgusWBP
YS/v0/sfhEBF9yh8jjYmX1CR2v0JhYRuMp97Bc4qXoSYNaWtYrDrYdunjYtp9zPc
S3n7vuQNgX61IEluSVi7LbsTfFFyLN3t0hkRi/ZYZ3xdgAmpDtiiKmuY42FrBlMn
W5l8agEOQ7WrZX0ChxfGQjlxsnE4z5YhLq4Py9bwfUIaaVgb8Kk81o3DkQF0+P9I
YSIOEiJm0OcFk58f/sJd6TEqYuF7JLfVCSQajENYPrdfT9DZHOntetla0nALYoHS
MgG1wB8p4Tpm4O446o7iTcZW9JYomhX1omB5Z22AH8zyu6CJ6OatwOcIuLPEIj+B
LQiKtKmTmvuNIyWldCmLrrNq5F6IiribdUek1nkoQSVx8IlJaPXSet5FznmmSfto
d4Actilu5te40H16IbxXl7rofopqd4V5TUzhh2Q69tkJPACTCFoKMi61ywRsyiP3
i6uumryKR4FTmZv/b9ePsCTevdlhYibPyiIUeyA+/ieNyiNI4a10MlhAI60qmZ/N
UbBqWLE6wmWvH8Oppes9cUdRPOZ4Eg74yV0QAnLks7Hd4jhV1uG+jCeYVB/SXmdE
x+k6teS8x+SU3i9eijmdLg5Jd3dgFHfXzPxhpTRZlTDe2Akgd7gsSH5VlKbyokaM
nRSXLdQkqpVrGBucqP6eMwjiVtjnv/mX+4eMdOHc7qZ4lvtlBhrl22JtrXsLg2e3
+oeihAu+c+DseTprY7Xr7Tw4lYkZ5/JaL6VUp59QC0apLjCfpwjs7soyWGj++qtD
D4DnbfHICYAJNm6EuT+iWpIcnzuhXrvO/0ZyeeShDkk2RvWFNJK9iBE+cjgALsiu
2VhqQHd/pJjT8+jAFdDT7O3DKH9OhVKoUwEuXvUgOsvx0sFOq0kSBbqUsNpcXAas
ywZGA2kI02fyMRqOe9KIqiDwdyjSEdb4EG0jjXie4QXv8y54XooZMf84gFXStuxZ
dCeLTw1Xj53CXESWYZGWV9B+l3xLoUrG+GkY649dQTl1BUvhrr1r+wcUPa8Ta/xa
W4kdTZbaNU7+T42raG34ucn3TikGNA/zHOMiKy9g6KnG0fUg8iGgdzmkLO9kYyfr
MDX7m1W+bFveZ720PYj3iBlZaa4p8prwhfZf0Cedpkxysvibn43XuwzeEqg4RkMw
iw9mcdv4xp8JLd8MRkKtk0CMABTryXiwvToHj5YsPDrk0Y/mO6HjfDrXb8gLo1Bb
5KujrbhpEW17/RblSU9nBy/Roy1YGeDSlQqyhvuwBAtmYQEjbSMeo/v/AIpBqgrc
/mnaOdafcIkQD5YA3k4NZCFDrlhOe6bvmnQ6UZorMEIEUMbMG0We4umste5WmVf/
Mx10d1f1A4JK7VsbGGlcPAMMMpbxbugWBIlmlrA2Q7SorT0Uw7nmsN2cHWa9cGwN
w4ybk/cf8HdZl0swFn/kmQicrWVLFNhQyD8SOQaiicxSqypb9CrWWHvmSEJR5F8G
HlNs+NvVaaUK1KvlGjLDZwdPvRMImDozDmpay34Zo+AVq7b3IrJqTuCGeXlwn/dO
1J4qZFE4QNCK5unrIjChVAtlyO8cbJyaPLaOk2EnSdpyOZLYoj7X9MU3otTjK2vs
fiadYZNcIiSRSWdSzDTfgQVvHI03KT317zGWcsEnebVFcG+T6d1pIqMXOxwyMu/X
QMp48Hd9T8CTcohy0Ep0hFoamd8tiOuiD16VTnMbsHrzaXhrDLPGzHwondLu4Sv5
y+ChgM9KnZbJSrKeb/0sgytyqseHsJVdyvH99CaqzWkwCdaPrq4L9sxFDs2RPwJq
/FAXwhvLdjzNnZrBgabo4XMpcTa2zDTX2H8kfgiNFjc5a0wXI0TX04bfMLSE9pDY
YtPBLE1+bJCBhnEQ7d/6Uh3My1pwTf9F4ogCNImXfH0B+V2rI5YcElk2DRvF+PHy
7dJ6UovYoWQPN6Ce9xWmVi6unkw9nsx4E6YMsutooKUfYyT4hRT46z4iY5aHzvlh
RGJrYOkeAfksITiNdH8KxoEMYAhhfCnh2NpMM4AJTNkp1yD7j47rgJ4coz1rrqhw
ail3tMMeKncp3J8ZMBKkeu1fC+iiyINcX9YvA1GC14nsaG080+YUhAVy+ZwYefpS
wzUrXcpeZ8YCAI9PEZDudNMNDRD5cbuwgpGpW9H4u6pY8eoW9eErQszpZIJZ5N/z
LKBzL/RXNgqaLJ1fq21EvzMT2FyBSyGu+ui3z3Jqebnygs+Az9ywA3mtgyqEvGww
LM1OZz0ThcTFkeppVf4eTXipcXj73MG7uM5hvEcUaI/3Lj/cAGHqCDv6ZzZu2S14
Nny+mLKtvnGnpgJSC/WDMKiG2rHg+WcHNfoRvS1WpSeE019QBICXqD6LI1rfoWkN
xJiS5tEQchaaoxRDfYjJ+TXz1jZhcN1LPqse7EMlAkpR7xNbzu5TEU0/G95vBP4B
FaxE5uzRJfuRupTksi7xKg0u46OoiMt1mTTf1N7wrpxPsiJb65IpeuAR+yLOAd/9
XCwC7HNTQ7BE57kWj7415GepxwbXmFBGK9BUQrJKB/Dhy0O72cK59PKOb75vw6Fc
OrbESDLgtTBY3FyWHrH5bJVJPgVHRP3JN5JAtD7fzWl0/8ONEWlvhlHagfmIhegA
gu+MMSF2bsjEPEgwBNB0dHeCbQB9MXaBKFiyQW3uk/tvFoVQflAOrOsdDzENc3jS
3EfTcKSct2dVVJDUo+/yBRkPFujt4h8hEK2J+vDyYOhWrGkTEah7hwrm+tBUK7Se
H8RYdy6Ys/vik6vTWVtcqSkhh9J6sdVHcPkv1JHIOTI8iaHavLuCDlQOzsg3K/3p
Ub1tm03Sz6uWrjEDoeOjfHGvqndZ8ZBz7qkcKscfMu8RdJSpt5nDgDjRuBZbojra
hkbmLYoKxsjgZeaes/XQJFkJyv59kc1VC2wpRUToZX8+NjimXTbnogccHOxNn2mc
CyoPZgdfeWUKPZiQD2tEJX+qQwCYkp1ffz9Ao/CAH8g5oKklZlYIBaY700p8xwOY
hWAb02MjkJFL1Zo03ZmJXh7Fw8XkJWis3oOJh+Gv85o/FhOSp6HdLKOZFfG4NEU7
+ACBmSlW6omT9uYfzdLOZu1xjJKKYeit+7XA0HApPEQyZASkFRz1MfF1LHuqHGRX
Cl/Mj1JAyZbIUrl+JYe/g8Rtlmokun6FDEdfkx8FkOtLhCIhIdw13SRfAWNaonxg
pBVtnVC6RtdqFQCMqgIGfIrY/q43/CQdcipLcUjDmDlX0X212DrMy2qhF8/QHWTC
/jmGyBv6E/rx8ZTC/oYhTdfj4UI/ZDPajWmRlHa3PQzK+sgOecLwfTPjQtb2My3p
c1AY+ycZwFFjABQeCO3NO0Hh0lqaUE4M59Y24YHoABHvx0kcbDPgb3ok3dAsTLHd
+43dtkpWDf2lb9ro8n2pHHnPJr0FsMT1xSRuqdd19O2iym0LFntH89THYSDkLgOJ
Ah1Moh6LbwH3OC7gsWxjKVAzCCSHebjt7J818Nnrr7GYH3dkE+GvvWcPTfgmhQb6
fgJkfP6HjHUJ69qj9QqOMfc36DsSzyt4BAqtS+LCfoNHB41CVcRwn37jtIV3NWFL
t/q9b0VjJGw/AyDmsxhOhMneuYp+LY5mNvtMVWE6KomoWkvPXp/LGuZncect+6az
HbNpN//oyUGJEvxAsbLPNt8FMaxMFACC0kblNQoscBds24BNNpmRJ4A5t/ucCR/4
oYZJM7XAdwQxOP0t2Je47xyR75m86xDJNwb41R89ewMU2mA9hWwo6gx1yWd+ZYzC
wnb5bOKkd3DN8k7Zm86T2WaCyYrDk+Nkd2HakScHjTLuXTHO7jyBlZmC7yz4hjAx
0xfMaJ9bli3Bqi+qjt/afM02+C8krMCCGSF24+FKzus/Fl7ZWJT9zTmxfX4UVWaP
pJ0kKWrTe7I6MOIPUPOcSOlJMwldNb43tm0NLwyfE0IkZ/2s9rRtVGwPifxjp478
MD6q8PIEagUXhAgNldQEb2qp1i2TLp8a17DaPwyNAOuqPCVzRqKnsKpETqR4NMHB
pF6H+nkOnjwP/WGgAaAW6L3iREgs4vhbDwjiJO60XzLPDvCgmwVy8g0uZ79liGGo
6Trogq9dXxMFxj71hPWwO1N+vknoA4jglPU8sUG2Z3y3uXNw76Q/80QJroBbwvMg
iL/LXTTQYqdGIw9HM2V8GNpnUZR+WS40MMzizp0LUJ/gBTgvmWbN7HINVZ0x6ly/
ek6vy5184nNs0FPZelNhv7t4i2GplRxjLamRnzrI/hSGpIo13aEfiinSqggbYnI5
h511pwpJJRuW9glY3JKTLrXGWFaJtrh9AMxbvOi6CwVAfkiw7OHRVQBOP9eTrnkd
feVx+4G1YMUb+7xmT2T1O2U+A+p43LUUlEP5oOdLPt5SE/Jw6qmOvuPyUbtWAOgU
00oa0P3oVhXrpGpHFZHOXkAmVwNHx/53Xnj6vmW79KI0D4zgX+ir0CYpFXW9iq7y
V0leM6ZzIRisuEJXcapqSr6nFhpOBOip47HYLnyaPwkB9YLC9LRYeqWFWxSGrTK5
IzDSF/Uj19EMOpZJwAPFTblsV/cdlw7SsCR3Z+ULuMBOI+ItnPkjYTmssHfn+++8
PVzIIPOIw8VJdiYUgqYOdS9PAx68lBgiFbnsS1eF6Mu4PhV9JH6ClyB1tBgmGnKR
vXYXYX6K76T8pIF945b04B6UpTrb/3dxvhpFfXrhEL+w5XZ41O06aAP2xLIq+AsG
6943huCuIV7h7GtkDClz1p5FqFYfaAyN5noJCDeckVSPBgRGRjlPlKLCZ3q+PWdl
vBQcdoopwUvD7xJiJCYUun4SfAYq4z4VU4iYXkfgGdoDCBdk+4c0IAzk4xbfpHP/
tbOqEOghrbtAk8zC04U7x9rpbtNDIdXXOO59IIIh75f9kSkp7BIYtlnkptRWG6eu
vgoVgbgkjgF/4LTf5HmeZxCRIOzDW7lCnHWYWMr4mDT20w6Xyo8g9XoZkaGEI0Z6
HnNOKlHqpck3mSL/q0OBcRx6AZhZH3E1PS8r54CNnGgUlKV/mgq13gshG0GZCSyr
kDFuQpgs+hX1hnKAS0jO2bRUQpEe0dKSdIVwMhhFzyEdW2pJHq140Lp4c0E9zE7o
H22NLA4cR7rxTV5YyYL/Ao1XlFlxplt02DUiGgC9S+fjsO/7Cc4Z/Wxtkk6XMVz6
xdnLnWxqFyJJSwv1+N+o2SIsiHZrBGYsq0GxSINbYj7ACi/huxOG0dvIN0eEtrlz
4QRgA33EcaV63sp0HPg2JUkl5C4mNgsO7IS2bQ9MKKz91GzVpnziIKaqVcX8VmaE
CNSXZu9g/R9D2IUC/lyCEp27RPfhrvcppUjAsYxGjrxzWw7MpXnzCW4JCJECoJ12
sgQkVOebGW995o3nZ8/Z3d96RneEcSbX3bww2wuAehPCMnaRUJyMkuMn2fHscBBd
whesbBwXtHmDvWQNKGf+T2/4fB9+kZ9xrBRRmAECOB8COz6nrNpmujvL6dsvuSHt
K1Qj+b/SfZO0Puh8iwEbQulQpR/uCQSJY7IH84BPz2gHCsBqEpOgR5MAfT1MxsCb
o1oNI5LOjO+jWupqNn6GMFdz5QLCGDZDW2mXNwz/fzlSSJocgq5naWzq32cXtWq7
HLcOc4AcNbDbwmNL9gimg8xFseBDHJIYYzY1PflbdUdEWay003dlWLweQJMOIg0p
e5xvOqZhlWjUbt2N59GkeLgWN2y5I1BdDom7vH69z5s95VrfQWnC7g8HQpDxVe+2
R7n21WPqedV4G8sAixP8dLwznFwEMKn7TCO21CPhvz9sf7oRRFhhhNOwR337viRx
TEMR8jiWuQWIrqGsLRy2ANVqDCsJJ7qsK5GfIqkddl0mc0aMz31NiSlBRfR70tyo
wdoXpB2OS/qpxJLaBVvbt9e6lKCwAkzx709J8clstEiiblhp2WeqnTRzfZNdaWLT
q5sg5Et8KkVg/TYvMCI0lFNzRYRe/P6Fh9r80dWW4tdfrmcyxh75UU/9QnB+WCqI
i0OUvVv6BHzni24at9SmsCmn4jfwsIIwMhOF4E/Xkgd3t5774fVsRpcq4aeXuQ3D
LrXP/nfYi3kinis3/zfzuBGqkdNQpyvTYp/Z1mZV1G0DKnIrF02log8oHZz9lAuQ
rH2UdjhhGcA9f8Y/i/T5C20sxyJWH8Dl1oiLd32NPq05OBpusxvWc/hOtLZX6xWV
cYvw2F4AqfAR+bt7p/oQLAXAxnwXBx1qbq37i/zlPkP1HO2LuUxg2D+zsIO7Pts4
doNh5n16ASuOTKMHNrZ0gwDIzILfa/lSHVsXKCeF4NqWZyeM5Pj5G23P4tHNNoyi
TUGKE1mX7b8NMAB90wDJqulCizGoQWSxFbo5J4GIZiPPy7jOdd+uHfzsvnWbjbrM
cbEsDO8BJ4qTPlStUzKt9QTrLAbyXQaDshAGE+w3lP+o34xrNT6zqUgyLcbn2kax
lMW8iwKIeLnJApVbejb8XTx4Ko8cG7FlQKwHD+s8eGr8u5SWvb3vw4qrGo2Q9R8o
Z39o8EH5q0mhtubbpi5uR5FfTCopVe79PUdS3AC5OGHh4qQR70DGnuhzd5xjmyxF
PoX5pucSqwDdZUJOmxqwDSYWyBt7tLulo7ibEw07UnZl4CAu3BGmheZuphxm/2lb
MPExKvRvSbw8v2h8DmhrpjqepNQH1QNY/pAL4Y9AuaLw9ot0NO/Gmyr5QcaBP2qh
D7Vo5ee8GbRx9YuFnYk+tXHCnLnXrZto8KrqFl1fSCoX5zkNb95aIwi7xpSPSJYh
IgQ1xvvQxkJuxisW4L835txULKwYPArjF0O5NO6ctKhWWUCJgeLf6jrnTfsDWJ64
ESSEg0piFw6EjVfSiTxCs+lGjvsxKWzjMBmrMx2VVx1r0dRww8mjpqWq3kQhZuAi
XzggpJk/K1wOeKaWQNI+uWJaKSwpnMkioovXr2/pYTRf+UiSQ8G070q0SHcLw7ch
ceI6ByKbSOK1dYU1W50Tj9fB2fq/uxHTArOdmpD6dlNsq+8d/jZJdfSfi9R2MfVM
oD8r6uWZmdBwfPpHDyuOB9KvMepF/A3b7UWA6kF6PwCzHazD/gCkGjNIhsrYlbqT
BSasqU62GYo851OW5Zgc2rW29JAHSVfX5DMp7f5z8DKKSE686u6QYHsQPkLBYqGM
p27xvBSc4GhfO+xdhfMrvRprg3B+8BKza44jsPiNIFQOWKDU4TUfhPXtix4z5Oji
p3zylvwgdb1eN2pE2+Gbwv6Y10fA1VDeVct6ibUBgEo6z/rlIE7THAkI2hTaIWn4
a2Z59sqXJXIlrGstXOx3mDcIoxST49aY0ObdPt0f1JrkNXrPqs30jqYWxDld1o6k
LnsCu++xsvGpLWFmH8inaujjW5tPxp2p0AdmIfwiO7sbOH4xyJkRSegXvNW8luiv
LTCT/WYemB8tQqazSQVzuk6ownEK52n92wRszs3OAMcF0Zvb4cvlyJlXLjrApzoW
U9CdcGLyBu9luSrsc0p1J5ac0aluaEE3B+LpU7GmDjkVqeD32Dn5zMUNSEpw/i3W
/ziSLggUqB8yK4o48SM1dhrsUcyaaW1eOAaJC5G36Ansdcefb6HikGj+6O5MriaL
QlJ3soGPzvM7rTnymuIjgHOqkR5uFdVeImR+KdNjoNe66kL3fiZmkQN/hQLB93t+
8sXzQRYW4+ep6PdCib/VQsa9v7awtcO7vORUY0Ig8ZKjmPN9gJj0B84tIcRXNirU
amoxV54LTpNWUzLfoms4fkFXC98wQdF2vTZ2uacfixsrkRy7P7+5kx1E5S6Aabb/
gMRPpPPpn5qdZlx3Bt0F+vZ6WuQghk3IH1tsp1x1BPDl2e2rL7Vui1C7G91xXyj4
BekTz2rHrUFxlfJkMeX3+22SH7o79vmH/VpzH1U8lYp36rKN08pLELgIln82hUQH
pGZgTNLytHB85hZC3PfYTBST28gsYiQw4jnCDaI+enGBzWp+NC31RvIRvZcdozwB
fISloWb85MsBsEIOrVuQ2yhwHbx0oemwGvrYgkPhiImtlsZrnCLNz5pmkFDp5OCF
wmomFyMcHSlARoFxhnwv5/P/A/G8Sj2ZxEK279XWvOtF4AEt28TSqvmC2DeKntur
F+g6yY99nf03NP6kwEqIJsV44q5pS9C5S/oxlweR6g7f+uVN95BZotcGwHqqTSno
x5AC0ji9Wbuw+XOWNf08HIaLAmZMjb2vGT/ZfQpi/Ceno2LRt0G5ooVS7pfAIJ+V
dPnK2y9QwyPAeSFGe8n3s5S69JTY/eqj7ooVne2gFHPCX1BNoJlV0RFkw7o7U3x/
kdQod0+JpBrewHlUexCxViaA85xY3LPSL5NnaFqa4hOcBoJLzrxS+qltHlvKKQqH
xS9xi165fULXrWeUKO9kbzeHokQnFrDwE0iWa5pr63TeINWHMxg/LnagJTv9Kdow
KF7et5ZQpjZPM8pdCGLVyrCzj6ZZchu7e//BCuXuS3c2W+Sm3N1EZr5ObzLXXupa
MUo38VPaW84CQBHal7a8eSGn4tYFvRaA1gHVxuNXI7fK2QPKfPYq4Uwlbmfs6eWN
zQ5ihvsJOkexjuIQ6n+NGy78hCAxj1dnjUfvMAerInYr7eNWBihpqWcU6YEg9rKj
8a4bv5yfugQ6LTftghPa4BFhVTUAvI3nC9F5qoqqIyOP/LwxCiMMVrZXPvUtVbmP
RM+OPV7eekJJ/+auPaH+YrkUWb/Cmk3w/OyG0T9UzLhclVd6IIufY/llqEpAt/QQ
6ak9Nhzy7dpxcZpNVC13jth2+yXnPFRxO6hMMzt4IDtXkEze/1w5TCI3agQ1p7gC
x1Dn/iZahNsczd/CvaK9xNBaplKRkDj6kMsZkNsuQjUfsCXAxRJd6lmsQ47TBTNb
Hw8KdSD3Wjry3v/l3ZTa07mnS56EFPwd/3kkfX3vyRFySW6osb3JeonIp8dz8Fy1
FLH6FdLs7/E3cOv0e1NmaJpQv+4YvQ+k6bsa9wxwfueDE5/4AV2w0+CzbtiI+jVy
9MwetozZW9d8sSFxq85av/O1EyQapIBsr7SsFodNdWLsGdaYCryfkI7TNZuIhojl
oYZRK9+RwvaGs5aWRwqtJTolOR0X9OXQQkfcjjXHh+4NCRcQOP/38L5ruiDb1L3d
R/X9B9oFMmtW7dyc4TNFqqdr1w1DZAZCnXTONCyt7QmMFNTESreXuN6PlSIfFwqh
ILKMWfh2u5LiaqVn7hgibHNRl0yT+8otM2D72FCoy7HMsyNg+1K3GDas+4zYg3EU
Rs4jCjY2A+y6pgTWQbbVvY8kKLoCUQcIjBdQs6L+WLxD6bIAK14IxWUzdZfKGSXS
cbBNwf7eaJVY5TRNQOoPkoGS1WKG1IqLp7kXr4NwLRSJkBZ3N2m+6YTpSr0EO3F7
3o/cJQ8TvF9+psVCY7iJW7rZ0nPP7oXpzfJgdp2hrmJHeTDEnGrj6YUFnGoaNWcr
uaH8nJWF7p5pKnczSSrJSL8Rg2NkeLsBBVVlXV5BAqJdyUQCxtAOSDfXaEA1S+1N
dZPEowhbqVXFYrmJUuJdmnSu5231C/m0RA0gzjjCpCmbAaKu605kRi7gyB1BOA8v
bjrHai2BEHRyycQFM83NbDuZm0giHCQFv4nR6/PSZlavBjMyKivHyqTI2coxRSCc
KfvewQ6x0fCid9ug1d0Q4xfXdYjYcBe6LLlpeH3Cr84JFIQaxJELcz1FAlz5GVth
ZUcIK//TgrIWam1hhNb+hYBtTji0wUfc14bBhi8A8z19PbJQicmc4xhablP/927I
PTZAgPPKJpqlXfsNzjsRqPuvVusjcwcHEC2YHcov8GOwBfGN3lt+1K+5/Fi1RR0W
ZgEevo2BFk56Bu/ZMdfJLochh8P/UXKZchcGMe+eIZWxEhkOGl2AY8+JID7IJ90o
JMdW6NZvrnDaN+4vjowb0WQMH02B85Ehez6xSFa2w5INFgRq/k5tdDAY3sGlyifp
igc4DL98CWS+MAqafihZF2RUCdg7GnCMuf8ZQRfXRV0+fcOqlpVLsFsl/9mOAsMi
qotjfmEaLPiVcMx4Z9XvIHA0nl9dWXoQ2ZFKDmjbuvlJ9oCpZ0gLIiyLK1MeV/Mj
6Jcm2i31mUwnWXrkjZiKkShb/RCEWcmIXrgPEJnXHryLRAJCnrQQ+JFdjMBMue/Y
cW3BZXBY26vaCxnYH8haFNYZJfo3bZF4H3/8oTxvnaS/Fl2tDT6y3P8Ua6uWue+2
BxL/Mf/ggnBARhl5A6SjBI7FY8VCQjVCXN34qWfc6dAZ9hL9y+5tp0P4fqluoOKv
2/0oflWz/+fYKx5sWOZrLu2d9m6LEQzJ17uNs3FSOGVESXliW/kq0bpNZWVDciBa
RuW5qPI7MNj4HVrWMHcHogVZV9kQ7Dz3Z4HoPNvJ73hWrJ1HuOdks9pIb4Cb/poI
08kuk35DZ3W0S9htbJOHl/IUHa6HrBEMhYjecaznWCIQuc9uDdn/TIynC9ELE8GD
rpL3n5dxit6UIWS+IKKpzsUszVbpNb5IwMCerzP1aVKbGYL1k8Cqhm3zNREw99L6
c+d7Bhx3FFwVAJsaS0qXcPGlbAXEmHyl+IZ2/vrR0MBPy+ZcMbRoJ/J4wfd277j6
m2KPFpLh6gkPz5gUVqk1OnmXKbgYOte3tYHLXmHRyaNqe66lBCU3N+sl9xAJWOT6
tiAVAmSzU//7f5AXnOZr5U6gJKcpfyuQLWL6QNFwLWar9PNGJI7eCcExe8aGSWv5
LJ3orfp8uyIQlWkTFLCGUpnJN/IjjXbfRTkzX/ztMdt2vCphxhRJ2h8mj6mYdvex
ge81CO1roussUH2tsDz9QmSX5QjBvPShMwB/oFQKighcYGCV4kzRyGL7XPCtJZ8c
5qzi0iA+ValLcyhYljjOJ9VmG21SiY9w0YhMUnsCNCcBVrdZ0OLg8lGwn8DtNQ2u
nFMEa42vZwyErxpX11Ok3gyPeadGRw3eORhW551+0Uuca1cmW4Mpgt+HAM1z7GbQ
5b+W4VISwKnTGoC8xfDN/X8fzpCz9BHjqk0KA5ErY5bT8IdVCiAypk4CevaZN5jz
+apgj6hQPSOyziLjDhyWApk/U7kwqlKmT9+jEMrmSfWnD33LFYYNJB0CCehi57s0
ctUOxJVOH7i2g951L7nTizb757SkcO30qYtHI8DUk5xk8MiGtT+ZqFX02LfFb8Fu
Pv8I0bjHnXP17y2uWm0enM+V6We23LVR45w0pylPqcwMn9pcI/5BXBqOK96JrktM
Z3bgT2Ww+HeYta1fq+3MdWaQaO7ecwVDsQsppEwcG55OUomaRB3yyAYkMHPcxB3G
mfjaYGpBujN/Qy77uPKEm20xhbfzYA9Qg0XAR9OTTjPXw0pbllHZ9kTZsJOYjTIz
z7Wt9z4t/eQ97Bvm/jpmragW/j4qlD1oN0yTqaSX7F41sf1inIYetZ/Znp5WOCA1
jP0lMjmd+VattU1Vdh43jn38uCgfOfniQSR1TUwv82TT4+OglYu124mlqX2zveeU
JZz4nAwRKWbb0o28bHHhNiZrasxfube9iFmD7ZcoYM9cd30UArdcSTSqOVXCWSpv
eO+YuFy1JC7TGBRmuiPno7Jcs1jMVSjHzZmWMJPM1PRefPh0KmVHZbLayC5vlAgJ
dTWlIFV69wh9fwJ3+WI3HtKB2s5Zrr3kWTubXzY08YWB9we322oJB7tkZIjvY+DW
07/l9BUlVWeClWccPKCfQCCNoC7DJLV9PTu32ccsqkJZViFx552/dj9AmgOGMokx
sbZL/Hz8o89MuZfe4CJrPFOl4JTc7VzHwu8Aij6lo6NILpOPKPXYSvc/qvcqtyHU
xiqPvh+vqCmkw/KLh6/sclf4zOGOgf1VHISYrd2lrQiB2n3GzXfBXDQoPJGaLmQu
qt8I7wHO2kw/HfKcuYaUrIxFBNfhTeGep0FTZUB0VolY/vHlk0BE5qL8uS/OPFlr
MGUE5T0ZkcGXa1OgUi3qCBy6e5xCiXmWA6GWTWO6lqnkCQ9RVXA7ysV7IRrxQ7Kh
OjuGJX9fA1Geelb0JXRmREJwrd+mTz9f0BQrBIhly09XNV8DzDI69yMb2yjL6tjV
5i9fPm+mlihBEsMFkWBql0SZe/6sCLB7/LlT/Fn/dXy910dTJJ6IDoXQEXiDCtuT
Oq4jrGXo8anSZEyOkxIaGt7fFvpnfspmGzNjyd3HtgAEf67dd6SBetXPa9LUWAcF
7OIx6B5sWMaDh11RP+k5Mo96jl+yrgmkkc4kLQ+hzzDGl0hMZ11JsPdUnOQN72Am
mSAaUzFYVWyK0vOt0oefSI2UzgVNp1zBgN4E8cWcHP+EGUJpUKAyxyWNCCtd9UKP
YruMRnw5L7PKmY5tFxm2WUiHP8lVs0x0jhXWAWukccd2U7e3M8zXvVMPMgNaPME3
tCQyu5iZwauCDhHUQvF/E5dK2is8vk+Ey8xhYhWCE21yAL9JOdykCldmA9gPib6V
1h3uVqpmjiWjK5jQHAKqp7pR+NSr5J4nepbREpnYhoJ7sADPDOyHozMKXGqj1Snz
1mQOrRrdXVGXsrTRLSPmKYhxSYu8LMETzWWj+8zzcDVqTHcj1VimNOW2Fdi/hfwV
7SYxWbqqIv2CfRDgUMfsLPOokd3Kn6IESLZEMXDBdLiiiGDfM6cHmkUaLoMRSF+M
m9e6VJ+KUuTZmlxskjQ42KUOcIazs4tV5UXYSbJKoML8pJNTlNWuIVkD1YdsUObh
HrwN7SqejxsMPtAWFKgpnOkRDepnaYbc0dBlXFJgx/QJE0CNt/qPLmXIzHVKVtXk
cch3VNoLNZByNciQNhH6UWLl9lgO9fM2fONnHsAARH17Mf90XetOTgkrTWzN+HN6
23VHqJFX6kg+aiVQfy40KXfnowLHP3keeVBAW8f6/ksCG8sQuhIcobL78ORWR/6R
2izFuo54VEBgolyME0q6mi/6oRPs1PQDJs9XJ7+qiJ0G37uBlQd+dcvIJ7yCU02x
SRsYNiOWpG4CAk2G70DAIMFDBMKtr3HkuN8Lpt0aUSxUDi3v9o66AiURYTBZYjfc
ow+A9BQ0C6Avem8DIvejS1WQXolH4NtMeVEhB+vVrLhzvtpxTm9ipGFspyOC5fNf
o45wxJxcofzAlyu50vg11y47GfeWDdbmlKcDNp3mJ5nXr5owaIUKMm/FQ1l315a3
y8SWKj4VTrofvpyuOL9kl99itL3cIvvlPms931SinhWoPD7TKzoLJzZaoYOsEuk5
d9uHVh0N8VodxxFqavGL1bKBVqnAyAvd4MdWrKEt7tKKk7vvuBLXrEHsKWGZEPfj
YhGFjCvqXfwEUCUPw68SkfebcykOAa7JmcG5JupAmLIKD5NGMtsyKeCqvxJ9YAv7
4be/3KervbAbdfztW68r3Q5LupO6b/ayH0paA6lJGffXdNVaINOtoZyfg9gO+6L4
pkm/MnGwqBWtK7V+Xp/dQnAW/YJIPwbZUVnH/8GUfj+yH14e+ZdjGT7xbrwi7tvJ
TwLdtZfhEQ3MZumbrsUvRbcq1YNsHwuJkNynGe1rvrc3GEb/7AVwEeapOpNONJhA
UD0NfdDR9sBtLUyjl8pqA1PuOVa0vHPoAMJTtx66m8t/SADCQkofnqCj6ZTtQndF
baNKYVKG8+s/AAg/xM557+KL2gxGtfchaAH8K1ty7CQCmG2nvbQflaKQ6Wyrg+q+
VeUDbe85dduKaEUAZCfGB7+6a+BF7tUvJM850bxe6P6ElBNgQEWdmT3cGzuGIKqb
SlEDqNChS1Y2sUVVh6eSBVYFhY7U6tPQwU2JOMur0cS9OYFmHEwMKaZSf+vVj2Mo
5zlyhjiOD9/9hjQXNPi85n9oFHeJSnxXr+8oi+FnFZDw5qzDeFhfHqWnprDqbttv
8aHQlT5uDyhLgZjfm70OuXoPEq/qgyzoEAGIEqxHsyV62B1aTizn86maNmuL5phw
O+KWnp61o8CerI2FfBJ05bLxq6PoZJS+9XP0VFl1CdeQQxN71rPGDw8kTy/LEiuW
UWcwaA9ri+ZkOBbsQlYIDK1wxcDMGa3yD3T5ph6VqVC2Hv6Fts8FJNN7BSAhIFOv
ZNpUoI+jX1v3UJnSrfxT+voQ36TgoRXDAXiY4jlD8pTMHeg8f+szc1RsOUexiSxL
UU6EWW1ASbghegsWflvtSpmG5IyDEf97LBzK8F2XBYCyvS6Ooaab0Ru2369/WbuR
bl574uKNpyQJbL7oQ49AjxCDiVl515j8mhve2E9V4FojI6tkbiEm5KZZ6VoHVvCY
tJncjNFHs10nworyDQTq787AMfv+u1YTpP2ol4vKYKTMByI6XSzPki4dH1nm5mVr
Zd2hn4E0VJyI4IZTSlDlcvFqVA1ePkKr0xjgA7dlBU6jW9YY6nk24sriKdoeOpfX
x2/FFweQ3mAosl6kwh+dUzYvGSvhweWs/X91W4kjeL7JtDVAtSipAikRtVlS6JkF
NEhQguNkdOD8uBUX7Khdz07H9MODZKQ6HMZZjhtopILlc2vHrOakKhUbTpJ9sSBu
pDPkAXX8/A2E2JwyQ5GqFd9CBH4a2zU+52MziHWSu1DLJxsu2X80Aj/2G+cWNDKU
/4yDy2xyvdOC6H2u9Bzybv3Qvfu/X+11dTp6oO99SN/31QzByE/q1I3tg49S/UKF
FQrdIIN+QJWLoMMPrCYBcpNZOnLsrsCTkdI3TH15jb3fIwQKrFX1EHgOWrBiUcLH
vNzRlKxWrpfVr3q23fNh224afDVbJfe1gyWycfjS5H423X/RjiM4IGaRIvkIWQdw
poTrT2PKxLnWj9F/pK9EEMUn8Nvc2l7mbLm2FG3MWpwEBPmX02e4BI1I/lrLQSr0
bVnloIMKKXE9p90YsaYXF6AnAGSY0UhuBBme4h3l/bC4R9HLT6+SYoi1+R4FwuQm
HFDrlwzAyCf1K1w3nQWr/6pHmiBZPAHa0BkoADfrhwEV628R+6FTA7u62QtedM6a
Lc4NQ8xOCO5rpAfuJO7iRrAVHrI29gjzgz109doIPdT8mWGILA5zHA3ch6JKY+4M
njNGcHhevXZez35/maV/tIw2keSlWdp5H7A1ZR8Z1ZOKVP7UDT0TdL+7L7GJR95K
9N5IEqYYBXLeo8URUtXTjWdYW6n/e4e/a0AXcA5MZlpV/bPhXzLJroROKwTeesUF
G+iPXT0dYmnbjv6ZSKvP9OJJaVgZCOx8qqL63oJ4zj8NY9eT7ZlX9WO6yj4SFMgy
m5x6u0BZXBvfNNBQxz3HnzvTYXSmjIS5ihTBKmw18qb0fTDF5Y3H8Rwo52THUVaJ
XsUyoyk1olSQCSM7ZCt35I9daxv6Q3q3URnDo6tFeojSMtmaIA2/5/J0YZyOxRTg
l3kJuhIQwsFTmTSMdL5qsw3jGOdcOzsbSisu8eu9LdLiRa99FoUeZakBWrYmIJ7Y
cRQPxkHwfHWo2EXenWTg+YzFR5dXWAbFJSJ+xQb+LY/lQNEZrqS8vHiNf67YAgX5
mNJznAGehQKEI372D6wAl5IlJ75T/adnb0dQjDlZXjlDWay3PJxPu5H6KQwKGjQD
rVr8Ed+MRrW4XmRQHDJ43VeRfkPeoIrqC4ci0Q/73oAuA013XC7KXR0o+C1INfQj
tH3cXgltTG3iPtZyqatjPdAsk4G0Qvj0uWR7n3/lF2pX7AHEUbmpH4khM4UUBjlz
v3u69gfhCw8qiiE0tZ2aOQ00EJvYQoffovhszIqY6PijmgDfIuFzaGIa5uYA7OxN
e73nZ/xGxH7ags/hS3/eEqCOS3OzEG6+BCUQFsgS6XBJxy+b9gA1VlysLWujT9Sz
Pb/7zgRjAhJ+nMttPhMqjaDXgkd3GKH7/OJlmE2i9s3vo11fOEaahakwExFNBgRS
kf4zcorgYsIv9iCmqcg4EEO0AvTldigvtLaMiOazvHGa50n4u+4EHvdpHKAZP1u/
IBuCl/U4eg2/URuDPV7z5c2dShy00cS2XlMc+U6zIhI1AsK+P8Kmz1JG5EEfFGin
tLrv5m94281uLZUrugMnr9Ubi29agLnD/ZXdm7kJxH8Y+WUDQ074iGexRlQPoG0T
Mrlze7yz2yWW2rK+IPR7D8ATxAWrP2xCMlzFEn9sP4AaMj0tjwjRbzKuN7bFfM7N
k3RIAPrlZyrXwGsZ4EQKxBkpoV4aV5TFx8I618SKYn4IszH0ZAsigTQrV/IDGjfb
cFEglwbxMnZ4QjSSowK8YV9fn3dCgz/Pziujw2KHLwr1BYxJPZ49q0FoZmPbCt09
zvQaIROeXcyVF8akyTg5m0bHh1qgFFf8C7MdRoFukLIbU6CP9EN+1HApKS2Yr8wo
L0nhlaojhkANad2ZE7ql/DtNmzwcvJq5FsGYUH9vE00CS3u7/YDOaYTLOmtd9c2I
rd65RGRvnL0Iu2iTKBAnuLBdZkOxEGWhfV7NpSEKs0a46VXzL/zo/KJnalgh174o
feg2nmfNcCAQ5RIMsDRC88+Fijg3ZATJug4RhXwjZC2ueOIVy1ly6NB7LtVuhdOn
K+LVVJ3PMXQsoDO3hwtWNuAsoWCICVe7a9FBbZSp0uXAsV20twWsFm1R3/vPZK+t
c9rtkGo7S2UKNgYByUae47j2SFMH4TodH89lFam/jgY8CrTOSOK61MrSaop4B7pU
XTz8jZH7xkh+RaAAr2Jx0kLa4wGsU1CXqmUXGFViLLW2rWO5ViybqhIU1L4S5Slz
U+m1uUzhiZom3E7ixCEsOzVZwIOEsaSQq1U8ItYSlR53TrPnvKa1M4MBoxmdLXvn
h5jaJaVMtRNRip6yrSV0A2cj3MPyADfzMovu0D6e6JZODF1GcaqM0/EVtdzHtqOo
8ALUUv8Vgab7nb16DgCA6m7nwBBDnajxDkxXeh6rxTg62U0r/Ph8PuKef08DF69y
+y6VeLn5FxJLNwwUfi5OHKgPGOYeORuJo097T951flQvuELMBBnFvJlvVetqVuXs
PNiGQmdoJaefBXAm2HSjabWcz7xvvryuxeIFd7Jz48prXcGsfre8nVVzID5Z/PFs
JOFTyePtKUqycSXWUEdK6Y306EUlvcxhzsAZ6njm/MwhfHNldgyhSOtGhFskhA9P
kFHTkk1+EbLKX3JiVE3ZVOnknFAzv+T2qdUdGBVH9Ndxhm4DCABJOY1ZT7CvzKdT
2VYTHT+q9am5rv1pT8hgdstX+68upE3Cbfd+TN+gPalkU7x06XExPaafZB/eTLvt
ncvvmp9dhqcU9mDzD+CmpF3xhSdFBzeRpGFnpY/MatJVxC5ExRWYjBWXwKySRgwj
Ym9neyyhHVbsWzJku71QAJe7QhmFY2nKGrp5/Ezsn5EXKlZ6UsiCx9IajAx5gvyj
+WyX327dlWEXYf4WRX3DEyyM8POhipRiEC9t2P1uuLIHJLaY1VW1H73ExoAqPK6l
f9dPl14viGgJ32x5SObr5rCe/uB1M5P0KMF8xSfSkMCB6SkFQfSzEA6mBoAicn9u
HVPe4diPhx2fPIfzvLTU/cGuH6qoZXIKAW0FiA07k4mTbu6ez6OgszY8x0xgAN9G
zba/SBHNGweo7E0U+xW3UHCujky8jDTWUYNlEoTFObrvXdiHzRC593J/kJhApjSz
Gw6HMCmuqPKgX8jgtz/zQVq8cACosHu2n69ZjA5yTPyYw1yh+mljTRRf2pHz93pf
w3T2ZTCOJx+EN8Of7Ic9sipkzKOynWSnZa9TPtEHeqHYU+xKBrdt9HW4KuPCbLtZ
TG85vhBVNRKLtf7G/m7zBIlXnjaOfbxcMz/fRWP5aNHezP6QdR+nPnsTtBRbcT1D
1UfTp63eAXUByY4d+Q8ciXrnG3HSKToR9AeyF/0HPs8JZGOEi1bKfEvgVZUXZBM9
jS1COyz6y7yWW7Ls4ZSb7MwwUIdzdIvy6yEezAMZBXhGjJ4GwlIQR8ejuk5Lkw/W
cFnEYgmWXCra6mZujHdIYFGNny62hG4kLQTRED1NmKuM7TSXCFug3E4SH53q5rEO
l+5ck1sUTPKg2lX6dWkff5LrZzm53m4x+0EwZDwrA6lj3UR6VWcU74DQ8ixk0PEc
3oKs9t1QlHrOav0HT7pp/+CnQ8///mLoJdIpvUoCvyh4juWWUh8xULWlkza8KAJ6
zG9V7B6V2EQ6Chvcsf0deeltTrUWVK71nqQOAG98AHIhynO0LhvM4bpUNf/kYUF7
jP2aY1jrcTAteUBb/6u1xkE1PmTcX0pVsZcyAtuuzOAloa2fiZ/I48KdS5Qa93U+
+Vweo9bBTAAdYINBsvLAfmmttqEgOC+2ynZTfTGW9gZJzCZtHAXVprCCKOJNmyiv
ivHqevm3e6NqxPQlg+2GPQF2/CqkxYLRIOUcMnlf9cB9CZxDhQ2LoOnddhFqhFFV
LKzsD4I5mU7b/itoCEUW+PZYcx4K5MOLxPegq5gNAmf53J8MVaIRIDyITb/zrw1h
lFO3u0Wjn3xJqI7z3GgOwg2LbtflIB6lOv/NHoZ9wai8wZIpXA0NlMXifbHgdz0H
SPkV1H6G298dvNjBS3WxQ6ledOW3pjKmv4lbaeh5AmyIZmlXJVmsR+e8jJwS0neB
z+S5I5Xj8mp2zd4Y+8mVb1RqLq119bq634aMuvO7dKk01iqobJlNWNvFVmkPXe9+
XvoNN7gRZruQjI6+5z3uS21X7/FS4rVNrtg4chd0gRV6RuHJVERm7Q59VgerK9LV
OnKIEiOHAifLZoOoUJ0kdtlGnC2yIpdQxQbDbrEnprjVWIbS7mrZSNr4TLX0gWfl
+8S+th3t02MfAhqZL3y3EkKXRRf2nyErpU7KpaXXWEOOhnoR2OWqOCisvk7mAtFR
OBCncu08Pikmo2BTpflMQlyIDgB13COAFcmivG5iEt1JXVNx8bTxQmtQc3QWLvlX
VIPLuHS0vVd0MoW4WGwfNLwgJxflmzEMzw9+6eS2DwpcAKJvTo9wjt/bxkD7lA7T
Vohitkkf9asQ4CcFdx8dX1g2p4lObU1lC9hb5BvIPhoUkNBHpKHa+uRCMkZbE77T
ovkGK7kQtbxQNlYrMDpEYS/dCzJ4BJ37qv/tbiDByOeljuHlRlrv99wX8WHY7hqI
qMazyxRz8m1l6aaWgPB0zVXxBRwOgRLO6P+jfxlV0oQzyp4LRMWByhuiRlbzZE7t
4SkpG3LUlJvFzRWJg6mqUSJxcYcmEdODKlxKHQJm6a/zDFi5ck3qvKFuqkYIfsRx
/ESwe3GcyxLkpdxHyq3K03BBtyOiS/CFwc1Pk7/WnzgWauS1mShs4tYAnpzQOcm1
6mnMnyfraxnnJi53NT7R+Mng5linbU9Qgrq4bQUrSkmtX5I/Ef38DBEE3Nd6Vxb6
otgqIAw5o2bKza6pSh9tUnQnt55HmcqTvRJlKzMqtM/rmbldUNLv342dz1P5/ojg
dUBY2dXgBx+lFBkfGWm3EACNZ+5mcLZBAW38KRCsuQK3+tvOUGK0nr2nDiq0P6ek
LHMLyZqMU3p8kjwQuAeo2LQGtA3RF5SaRgdHdgx/fyJyTUiwk+eRZyzBa+6pGVbL
370fVlvHr7A6CGASOWbNY2Qk8RMlz7SzkCEdWW1aldUBNOZyaM8EcHEPXY2AtGbX
sPRWWzLSRgJYoQvk1DvMqGzKDKW79S10PPzMGfoEz11o69PQ2e11udH/8Bx8Ia9U
jZqOZtmJ1CCgNAIj1p1yZGKdTFQI0aob1f5oOxBj1UKbXZqOw0H8J4u86M06x23x
U05OsC3rvmimYrVtn6WCogjk74gL8YgXqBkwALRjn3Yp/moUOUvrWkH6nt3p/+qn
cBYkGrTF6eoYMaFC1aMnqPFnE2n+FuM5QxenBVs9kLJRZVGNjE3vqN/dkWkc8Wi8
Zw2HHmoKHoJJ7KQI/VOaqhMqzo23x5ZDqb6QRNbyT3Wzrjop2AMESJz1hFqGCQsA
NMgkznjoLmgY+q7fbARxnmj5IUMyRTPhI2A3zl7hhPxsah8947H3KR7ZwWFB2ar9
4YNOOQC3JPItTrj+HIY3Hke0q2sLQ6QhWdtybL3YRwgPEffJCEuJyS7P1V0AglVk
UNCujmFZ6AYs0AmjoEZ/KteFmat0OYmEmg4EtsuTjEMcyXc3hnPmB+pJUPtjGOib
x+C/WDXayEj2XngzQwkjSnT6USivuX9fYnXqjR4E6c92e57z2wt74KvG7v0Ofta/
mnQUsS3iDGNmGIGaP+9nUdoBZgXm4h4ZCMEhd4sn0q6ukBKnYfVPKvAY9C6z5n/G
XVv/7k+608oEpHsIU9lDY7DJJarD9W/vzy61LFfOr45fJNehgOU+zrOUVTn1NTyV
CH/eWVU79LTLQqwSEz7J/QSE8FhRlnVRWD7Nrk065chpZ1yKXUMv8fT6ljCaNDWz
CTnJgZXpvWz2BaBbUxVykueE84UHPPt/5lRQ46ekSxVcGGyVAThD1fi9S+nfWTj/
uok7GlXQjrLma1xViwTE2pdVJb6M7oT1DFY5R6zLRWYFpidJODY6fhDiPQu7Cr2p
m1mY0ybKysRksLh7OpHS8W5kVsazNLrcuEw9iCIdDwVU3MeO5eOhSkTrpIdUS7PX
K7NXOWkR+GXLwuufD7pv9cLELDxpl7AuBZSPZgm/ozp94NCODRzhELV695LW4GSM
HzrIsqbFefD6Cf0pZn2dzFwA3j3trz/hcq64ib19zBeP0QRJhG3D93F0r+9BZ1D9
c4hIp/WDNw2dQ3EmqHk+AagKuY7eVxZhU94BdeDBtYQCNi31Ov/HFjFVjkuPpfnG
l7bFszYT47h5AICz+7IeMmp/p80+YRhTWVZeB0uUWerHx6kQNXMLj+drS4Gf6ALE
0G1WL04s6bI4ee3/hVykwv/mv+UQ/r2Wa2B31rdkPVpQ9Fbi7fHLpAjHDx36Ibvx
upLiJPiu+jVTMqg2yFzR5INkaDY86bHNVq+Ybtdg6nwjXq2UdCKEpWc+kg//F1OH
zQgtE5PqYAukfis59QPvwz2c5hlep0o3TTK3kFdAt6hDaw4Ry8b+LHQiNT+3Zs20
0DeVM5bFYkf8T0BZl/mWnGKCdQK71veCdtyaLqUgu4Mye+0alZ2tB9dQdqYgPgzC
AL3CliHuZxxDNumBERTFusdl3vAEc4OCXZ18xflp84k2ESxyofJ1B2nB9m75JwzU
KtpJRPOu612hyKuq8E3HKGeDR7Lr0iE5ieHqYUf1X55x9UGZBw/mtUJvbC5mETF7
Xj1kp5dg/A3ri8/NdsLK+/zCg8IDkcu1qRk50qsypADhTOGQr0QOuA6zEcU1juys
5cGy2JQUs6oMzGh/JoWuU0yWmJMlHCCQ87Low9LeRirrd4sbDZ6ApjxqXZ9S7ZoD
twGmlHBa7Kd/YmrPgnEvKnRk1/rhPgyNyT4ZTHbBsFmyQwTvzD5i+AZ9Pd65WsrZ
2y9uXZFjgFWefWUNpXeEWsvmeCHyluewtKzMJaThsb2ZdJdEm8ysqYf4AmkaKgQb
PsJaRzG/p4PP/8lRqclV6MC3+gNRAzNCrOlgmuLqq7u1JiahAfcsooedg0b/e7Aj
trA+QehXtpPtHjSi4RyfTDQMv6n5bUvobHF2mXuvwKb05pWqrVHFS58L/dtutLAB
07epnEbLVMMLxBQG62ff21gJx44OQouOeoPzLCZzLB8Q/Cak4eIidjW9I/w63H2r
1k6oWlUuXCvSCwCgjeA0FpnxscsoeBlnt2TExx/GaAxu5RgYMSuXh22BdIBOBe//
BX/H2QFu1PTnzxDGs1SFWAWlyFenOLdxO+iwmhWK5MCSwuSNSIo7bLaplzAipR6h
OAZl4PV6SrOOraRO1eoGtsN/163Pbp6lgebCxSzIUM1d+wMpTtrujFVTLDRSeNkZ
+DjBxQF1ZOLVB7cTC+0p5Yfaqzias+RS4zgMcBepiDPbnMj6F8HgKxJja+HjxG+Y
vX67HrlNDR8ly63duzwlkXpUFV2NA6xxzoKsLnIDIBdHVEJVE3fzpOTETdkbtDrv
zEgtKGQxLlYlBefkjOTA2U2eV74LzGhLXOQxaWInm8+Ys7XmE1VjBvKbPI+6hYoQ
vFRLxnQnLuo3dUWpSYkzKKWUVRH5+iSFTc0jR1edplpDcsIdKeTYcK8Md8SkKG3l
ayXrwfpaTwpBaMJgONNLa/FQO6rCkGCbX0UaccRpskqrsA4GUePlCBARRSeE8s2l
ZrFMKyDaPvWm+W0ODf1t2BUCVwrpJsGmGdPQwSX7Dusgixm1CWbab6Ro8UUmN1KA
7bTe/wTAdG/2g+Gx0AdT3GcXOt3dp9ULdAImnr+mFbn/jiL07hgxn7dCdFLgYMoy
1J8cMf0EvmKDvsdaVEDVnU7aDKd14QMVvrmDyiktGphuxJwkYRbRcK86vqVGzUxm
/8aFhDqzpkkV0vNafg4gmFgD0GW/GWIvemYrnRUNSJxLcev4MhXw62kHULlEwU6W
oedSi3C2Fb5XNKz7qAWR3URa+pOaJoJFP98xs8GgEDK4BaH+nJJFbCv1cP2uo01n
qMj9ZvdYlT+qzcsUlhcJy8zjBMrXazY0xonrn1nDX01mdwTx1a+FpCh7Mrmnaoct
UqLU0hGMAqDGf2J1YuQw8zAfPzmscuTP4jb69kAtgtHV08URIOPuUs5bcq0ObS7/
zlRkMqAs3kwTga3cZMFRz53QMcPztfANjhgBWgc2ZXTEf3fMk61g2nFA/IpU6EMM
iCLhiZugYXUbYhN1JNOTQKqew5+RpcKCYCg4ZEV5lZhONvHhFl1Aq4OrRPS/tMnp
hv42izXKMjmzdEUeT4D77aOq46JGgneGXEQSGbepWuO9QeCnBBajFTg253eRGM0k
HfugGk67OvwM+8MIUxdi6bZS1Y7+jaOoKYgxSLfDPEQgn1cNklruoY64WwUGPe07
g8BvuiWFroplTQGE2wphoNVvWrhMqHx0pjtF3KgcUw0+YuEqEk0lHZE8DXRolDhC
GINAq8VxD4Y5aQQPd7sHTIceiUVgxJat52ICx42TC2tuUzE1CVTM+EYaAJU2845j
KuFUPkPkpa6EGdDfmz2UR/tBNxopGUDdKrA8/X55pVb/N987YntQ66QMbqTT8nrt
uYZiHnfUduw09vgCYm+mZEtfVmyHDf8hpiQC7bI0hpryj8SDEOj8DGllaVqIRDh6
NYX4glAY0ENTdOqzSYXZsYC8apqwKMBDNlszYTzrh2cXofGGMRlpSTob6N9dMvWz
wwDUjqyuUhh7rTa8U2y4QvP2D+0OKJ9aFkiK5OAh/A1nJU7fJM+GMumLDtMUoMm9
Z3VhOmclMjSA58TWrcXDy3p+2GXVJt1HX9v5mBO53tfx6UohyIWQzt7ut1jodROh
FWaAEszPOfihXPWyduVt3hWljge7WAj2feQH0HaxLh50kl+9yYv+nNOqsnES2aur
dN/aWo6QHRBAJHkF/RWOGSCLb9MbAKKmqn4N/F46m1xgeMKTE7u7dCsYP4OfEfF6
hRolFHFXC7IiHj9ueRNrbImHbLFOoKpwRE5n+YrD79Dje4tvZIc+wH7avLII0lac
xWhCBtvKGyCTefhYSzO65sGUeAW6MBfNCaCE7AbqhUwOfJ9rC5yeCgRR+K6uAbDW
FQVPILs6XdcSYc1OIRM4/limy5REWG3XSWYzAhxWOy1eHLW6bbQUtecOLooIY5lc
pvROyjMo6RBX2vIOhThAGwBUQtcI66XyKXcLGNLylMZkB3T5P0GGQzCXiTzdoVkE
CHqiRL778p8BDhBGRw4O8xF8mUbYTA5NZYMoeBgarfzHnWoIzh9YeO48UXhZxWIz
DdEzzReJfHYjgsQMwXQXfxKyJJCXmTd0vbLPrTYe/PVH9CSrbCzuN0Hl1F7A5krY
KJ8cWL+yMBiuMs67TOV1U6kiXbhz+Ahw5UpBYJ2Y2DhyylTZtEENPiChDvO8DjQn
1u+4IBS5Lx6+UVMIcU4ydz4LG+L9ILKks+y6+mKKN89oZFP/ymDbH9hv6GLTtmku
qQDz8t15ucqej+GYLuQmhiJk5fMILScdCRhDZz6RGBu4hIdlHBvJkS3IZSuKK5cX
M0YKoo3+R6KqAeNUMX3m7vYU4ycOBBNf4uObgGDVb7HGRoDnEl3DN/HgSS9Pg/4L
VsVYFvokFoMSruHZmKaQlvf/ksLQvFMtNZ0t3CG5CqBOkjVdwfq89jgIx5nZiY5y
FA8qX4gQSsCQW/MpFUSd+6rSAabglbzaXXvIsYv3CZAF0EO2Qyh5x36CQx7dg5fX
oIF1oDbzqTxHT4ytbqB44sQB3CWdITQVj45c81dD3kcrZap/mbA01qCcQIc5kbA5
HiTYBonaK5tudMtXzR2YJ3m+HWLfLcvVRMRZmLRvRUsaMLQbVyaERlci8rWTQD6F
7/1Xypc03/4atWxpy23DZIXI8XoylGsEbO76N5DX7m0rKKmfFDqx8iYd5CrAVRrp
fnA/8rYvtGUU5LEmw/timh4xW79wK1GUrW4KjJLAEwtFPQkf6/xveTbJAc9ibXwP
4T18fMZGxps1Ga3nidPzbIovtEDq+HXRySUnQspGrPUwu0ldq2dkbl9p9mKD8B0U
GPis68BQ7r8ol9Xs+GiK6h5yScTl9wWZuxoYShXMNwwTUWWR/3sKfeKzrD13ciy6
gT3b0xn8u0ChjpQpMKGIUUnErBwWREEbBONeV1QtfRH7AZtOjQ/LqCjaQcGbh6yQ
4yhekMp4yJlcHGOPbiiwlli0UPE1W+XaF6pBqDDn1LdW6iV96jhdMUZwEbCijcSG
99vP17CWexh9sNBuwnk31Y0DOJypK+UQMlAQ5CHp2MAap6hk68jgcUoj+vTWJjkJ
dlOHT7tCHQqc6SE7WD0JVNGeOihzLMbYQQity3N1RuWrWO3s1rZJqITj1+2eqX96
dfyLCD8pB1+TI3q4vn5B7gcEsu/DCF4mtR7QOC4RJE1b7pzgPwGhM/Dstd5OLOtM
aWmzAknA25uwqMZ2dRgUWRWlFzD9+4uHNzS7p5O/3woEHjnJ3nwTED1jiRPMTv+m
eU9uqVGRXbBqcEZotocUO/sA8e67h+PhfWkrQiAfDqGV7X9CM2HhoCTYOc/8mTQL
gDulAoG+lyu2fN4RS7g9Me7MPw7Qv8IwJ8DgIuuDY4Rl1mkFlNzxKq8htf1DI6AZ
1HmcVQxfu1KB2SDJXWTToVf8SN2Ez/4u6aPRWB230KxpS6oY3pPr/xZzKzuDFXxy
r6FAFygn/4LBWeY+iFNf6Ue5VwmChUOu6UvmgUnDLRUl7LRW/LyxIHUkRp5etG4z
U+KOaF4tVSWvK01uU7NM4RUicMwkBgrBUBFpzpyKhzuU3GKWFNqIb323JbnhU0PI
b1VHu8sVHDU37OOC4KsvTs8zQguzpHfls7sT2OWoLM9jJ1UFiE4d0Q7P+lwkPgpt
WEruE+8qODRNUpdgfDiWRzhOtZf9cdkr0q3AydBCA0OdJWedM0rlxP0VN7KuN/ZZ
+6FPr8f4R+a56jGMSSKGzCv0srpp2FIlx/C3ToAZzh/i8x1Mzlkei6Lo0fJNjXQS
TRfWg4lx+jQWVjHtjRZm3VQ/Oy0I2JRsqEJuP0+BVKPppLN6qF2Prg/SGlgWd0Mr
UgAEzVjgJM2lYmnIycRCJ+tcRRmaRLSA/zkduiVeWQn78qyIWYr5SpYc9Usc1nXL
dF5j8KV++7cwX9Wi1xPHuCqge3BQUhQURwKzer1YUUJxPxLKMI6FY5lWgQCmT6Rx
JLZfEcwgG0/702+8q9eU04BBAXcUffIJjNApNdJ2/r8zCbx3CjVbWeJ5uZdbwyn0
odrdOYHoOlY+3qhm2/VGHThpUbaNhbZki4mbp76XwH80k1jk1zayhNFuTsdSCEAo
LMsHKQFYewKnZmTqcDMJwCLwJRK3lIU3YznNFm+WqoJybiarxJOYlKDdYmoq7DVW
exBB1OAAdvsVg2X72ecDVK+ZWQs5YhjYo+7NozglF5ohtnC0UoiAzX1L2yNYfmss
dCLnBtrQ4Fg8g4rMzINLA4CwGJiu7mYFt/gmBpuI6eivY3XPFHuAdn3Jp9qHdUjA
QlRFzcc9JJZVwxB42/CdUJU5bOb28x8e+EV3Q2brZbl041w/Qf1jY0queL7IDgWa
MFO3cvpm1AVMJgN2WUz8pDM3QtfdIrtaDldgqq5EwI0v26gr0meAyXAqwj8XYCj0
BaHeF6ri17OvGZuzTN4eS8vL4Pt71noT/i0XtUuOEbeW3ZufK1BxB6sDSVvP6PHt
QkUwoQRsjG+/abZ65GL94alWQ8VvM7oV699fXg4uuwVLxFBcShWFR+zObHLpl2Za
bpl9viv3ySEVWOdhQKbE5q/QFGwaXcGteZmWzoO+hx2xwqRwRkkSPkdc0rRQfCdd
ARpjOusCClmvS/Edp7iz5w44yOuWzd5R/Qklj2LnzgX/PzjgS8dNjYucGr8+cQ/F
HiZ1frEfUjZHhrzwN3c59NPBDRW7L2n0sj9UCnuOf0BLkRvRFBJUYaNbCGFhKC+/
2hb+k/t/NNAgZovqB/6fPcEiQBMdtMhKCXwdWm8GoZWalA4qPRW7a5h4D6BwsBFQ
fOgnhH+ZrbcTxImBX3H7ruuWCuBg8KXB+En2o5/0MC49YaQeCjXC0Sa+IghmO3+R
vGx/joQo7bCrL+ZzPvXk+0iPpYR6zIt9sh5VRWNUbtngaOjkS9OUR1Nsfyc+nOQV
kV6VLOH6yalXwkOMOi3Qss0noYVjnWIx4A74esGD4XRvVDTHf6SB3llegGVSeLGa
gncVkhqFhbkqIr9qo7gCOxQf59VR7UUHcWdh3tqGykg5LMWReMncyyjZoNTOg6jB
hYIgBVQORMyuuewLEfWRq8tMvSBs6xZ/4khZVEH4P9cL2UGxCcyUpCob8/zIAnZQ
CH1tHSi7J787v4FCWFP4ayXHdSC+5klFcO4nQlFXl2bDQSwJ1ijGvz3jlXUXeSKP
UTP2s8C0x58EltibNOfJ8z0xmTYyfZhNovDXI+7fyKjbVHY8ptSlE4rrzZ27tL1l
nRsfk/Opge6QDpmAnVZv6ZZn1diq8NtVNugQ6oVsY/a3bUSBAKwOMOko8d73JP/Z
E34yHXrLzrzcvCvAgjOSF17ozNx9kSIzewZf3uU7MlkP0Cpajives/8ofDlHVK1L
dwRMk4riVSasTFl93fYxuGHYVS1EVarRG79voBdXVidb5fiyE0J5mUYq7Zz26yRE
BMt4a0q6w2kfxxNGRUz6LNI78i+ccx5ql8i42p+j3BHtDs7mobsJfSLb8TN5SxLN
iUPYUPyCVUuMWswWJbmccW1Z6e9EJ8gdeVbGj+1E0HETD3j7UNiG6sLgEpx3o9Kb
AXrkSB1yMKx6rBMXmH115sBY1ofpa6yaubvCiEIR06watte8Bq+sPTfRU/3NcYQn
PuD+e16F0TDcruvtLlvsCefLVnRlou8Ezzk+tQHPt17zYr9CSUNjRSPddwYRN+IG
O0h+WhISp07PmZCMreplTk02iVEuixgmv2cw+I8AxRenEgyNiWOTv6TV0UhAy+wz
y810ghNMcOcBSg1urRAup7zHwxhdagpFxu68JcweGNvjrBt7JhZ/VcUCIOcx+UE/
luIazi+xtPeIMlgCQj0MxqOaNEaEOgysrDIrIbO7l4uWhomUHATUn7om7cXzEeR7
Xr7AotmZYBoyKvlHMDiVHKkb9KPGSG1kCQFIV//D9hzm4qvqK6fZ9nvRmdHBNY3s
CLCtdePBYZg7uLYcE44zLggaQLt9kRbl8hQwYBbGKR2R05/22vICNBWBO/RutY2O
tLFZ3vAnylLGTE3lkDJmHOvSXDs0DJjx0RGziTOClzVrfH0PyUeijPl74RR+xzEF
akp5NMq1Tu6namuqBG0/uFllpYWtQMfsNCwud1UJnFyaMLSiu7L+qUqnYOl1HXsI
muqG9kFluhXQ9lFwEf7j/B0qJhF+DAeCtAQ97K92HeP839xluwkJ9nhM8vnYvJBe
Qeumm2O1AmtHCD8iL1eGuNiHw8FARRV3Zhr4czjiW6eqZlXyxjINcCTqlG5Ou2MB
dl1gJwp3job5luLZYaGbOaxWYtMHqNy9twZQXU3DiQPnt3q7NlJByK1k5pw9SsVc
9Qmf6RJFyK88Hp6nCpYePV07AaflIpMgU56UAfhlf8OjIj2ze+VcSqIxwqkE/t30
AGxtXkOysjDKr+FQ+4DOsHaI1bWiuIgjZmPDU1vhF7wWvgEpqAIzGLDcDKk1voPg
4n88bcAMXj2F2KLOuVXRjf6oomTW6C43yF0aXfLG+uU+ueF4vNeWXNHciLCbgMUp
KvolBUsE9RQlI1bh2t/rxz2Yr0nMO7YYCSIzDNckXF/lhaSzBsGXqE2SVl6hZq92
FAC4rrFN89LUpb2XN0u82vRwO0vy9RThfuJ1sjYkeD8Sek0BE07TYdPsVslh3ZHN
y4mn22cTeX7WfTm2+ldPW5YwSvaRfksRNyvdgYDy/eozZk/9UBFWF9lBaRxzNLFf
UtgtA06YPDCbAK6oKXmIEMEBPNE4AhA+xDAab6KQh10EcaItu1kXsD+cyVd3yvo2
4V81U6QzZ8HdiPA6DmSA+kRByaFWpupM69ugjr6q/b/kuwLHn1HPKwehCzuK+dgo
4MQKMmoRmDg4ilEUlONWyVjcUGIRSs9RXb6r/CJqiJahztmo4w25hVZkCVYb3Xod
Ox8ONTizYfFrm0ZEoDhTpm8k77rJkGox1qQVfLUgRinKVTauujqJvE3fQFfaLVhE
Q63Q6sCZo7h8B5YXmBVdRcOL6ekqp7LTzlz2Ptmo1UyqOI0e6gr1570fzRK1SPwu
4IUlx/A5/+ENfGnjKb3sog7Gnr/W8+M5FX/mcXnxJ2WRieHoFeG5haV/K0wDceww
Wg8KbHEHFeyrFCzA4eubNpy8FWg22AWCYcmIF/x+LdGfg/bU8Xiu0kFnsYT6FfEc
3Dg85hLrYbtxDqCq323vbt6OPisgtFn9V7R5gzD92sAZaBIhv4u4KRVQ/+3TIq/7
t9pAodQl1QR8MC+oPlouObTiVsuweRHLqGcyikyd5ZtiQyscqJNOiR+sbcIT981T
lcc82i3KpIg2CRconOJvOr+bZs8cfEcfWwZjIO3HgddaxiF7ZIxysy5X7+nkrXZj
2DdYXhH5mdepfxBGWRuv+HG4/fDFou0dcruRdENLKfUI0G/4T+3A+f8nFclOQ7z6
SxgZRjshlXwrcaxrrU7Ni1HA2D0RNCLI3roB00Mo9+PZQd9Kf8e8LofJeinbd5m+
fGWvxVkVB87MDAIA+HPO3VihRKYBWNPzD0GKMEW0zJEbt3zxULiyDD1/mbn3ESg7
iQJOES/SRZtdaSOEVKjDRSG7up4WrIur3HBT8K4Dp29nVPy5O0WLVjePPf2pukjH
EI56zMGqvM0RnfrEMsyntZv+Rg6hy75lRrFe97hx4ulnWjQYIt4DC449eZLU1cP2
wj7qyvpkTTZIJE8UkO59QWF8br8aFVqLpJHrYdHxuCNLqGFElZznz0c7drUerX7M
czy2lpmIle2kDRjqyS/M72C+t7As2+IKAdeLNBorKlvZV3cW9CHX7BO+hlmVBzCT
IutULp0lP5Ztrm1reGyT0ukoxdbz0v35/MQmo3ehzpMMK/ku5y0yhuZuCA/GwS/9
7i5DzN0DmdEZErSuGggpt5Gn1Abgdm0vD+u+7KOHY7Sa9S48lFi8UrYoJLM7KaEK
yRPwZwFBw7zOCc2DqqBm57F9hKiYkgE90876yXjLsvVxVijahqa5uT56Pu3iEDnS
S7vcqRHYPX0tTRBzJR4BoKjx1th1SN8qTkwrA/k3E4PKDjI9pmX0YlJ0eXtDFXB2
Og9CWSkmRyA+mhVclM7KJVMlXdq9HyTJj1G0YB4Qa5CUXvMKK+MuTholj1H1Ta+c
9zFCbdff0TdS8qU3AuHaiKXwYSeQajo3/omszhgqnjtJLA8KFHmaD7UuZmoZ7ukJ
7trGXao5MTxTFK5HHZx2BUKFywezAmjVVDOF9o1f+eyTmdVuNdc20DITn6qqILxp
m/4EbiHUUWyUR1cgKMn1Z8Rc7zlT9eMvZE8y8SRo+sCS6P99aPeELfLTrrecTkSr
RGSu0zTy0IawClSctUzz9iU3RSYGHlEig+sY6IWy/4jD7LIlYzpaWXmKigBJX7Y1
pfIY+VJm4t7qrh9xxAr4dL1Tlq5QDdhHYKTeWclzfs08sjI+v0CYXXQL4KtPWzIR
d95JX4w26UeM/LO/O+lwpsIz6mt5hv7q0i5gxlv63XAZvGkOrn27m/WrMGSlI+my
YErqBFDNiGTsSk13hi/vIQ3c8/I4z1qajGvCTUW23aieK5k2BzSnA+1q7vCgwM8r
IzG9NFFXZ68YdZivozXvaZr6remQIm3quR+mQMf+J9qylLpVnTkE1lsIElrhQzqI
Fbpk/p/YeHSUm800mW/D7mSk26Wh9zYKrl9Zglz8F9ncr9e+a0zbtjuQ/fzWVuHI
373K2yhdoq+GnjuWaZfMlo8GiIstsvMDFIi6a4WaXx3lUyL6vo7ZIw3AxVfSVTfm
wEc6l2qUnMMZ+6K2RJn4DrmzaP8zlja/Ur5dEWtD99prhSdmzkXruoiSbcQIpVcW
7BU95+iSY6SpejCiyP//8g8ECPpdiQbtDRwi6L/xChsppiSsCXfSNRmnrt+YKBle
ER0paeABv794ouK3HAnc2tSpqLliITPkzFwXpJbL6hdxMLOcr+gtfxl/6TgjpIdh
WOj4J25CcMoYVuS4bXH7+dmcYF+M0Vk/al24l2Jdbpuy2qhqFIuyp1CYLnD8HEjH
GSFYt+ntcnRSbNVNhwngdXNNGWJTDn8k1g1enbZDsKxRAt/5vno1vJwE4p9XmeKz
tWcDp2H1FoyLnry+pRRlQOgYfzZtfzLUSrfZQMHUqIlDV2CHvPOInpfor6bKk/CC
XxyAHvmUgOS5q1Ww+BYtwgFvifZlLG/6Qn9iY+HQWJ/saRN0Jnx85dLXR+NaV1JP
qpFQ3TgEujZLx4YLwLuUzdQ6jIvny8i9VgJLpeAPR5uiNUnfBEELxUbKe0NRTGkl
I+F7+vizwbX2pyRDEtDaHNoLeZbpuE6mDbzM2KP9sOeoiwxnVnlrjlA5C8mPeW9+
q/T9jxyTOKfDqN5A789Y0z1yk775wswFm2d4Jwwg+Jrd+mySMzXLe51HJ1i0l+Ad
6T3LCRtmfay/B6qB8OYN8oxt89hH0tMO6GE4eVGcDqyszZWoTdXccKisxj6hLN9d
BPM1jgWangxAYKGuHG0CuW5J4S1U4tu9d+y96O9YKDSSmZBEjdfmSpGdH6wp2nji
i9YMO3SqvwthSSxznpaUN72sawE9ICuaGmc+BnsHjnleYx2mIrvVouGq0I52oAVh
f5cAArdbnKmxiREuXrbYj4bMZ6Kz6pLt3OTB3yH6+AINJKDYkXdqrjAOOeXIF0NO
v+eYnQnZyR9r/1v/rs4+v2/H3wS/noGfWYXzs/L4oUaIW3pefPdEBKcq6gc2efgj
kIRFOvio0tSbjoYWs+CLyXiZyN6uajv3FKfxZndgHU4+z4HTIcPlpuRXJJ5Q3H9s
ltOkAjPrBRC4GIxapdOqVBONd1buLkISstfXwtcfF+dPdp+ivW1idqVSYYGFWZ7B
8ETcJ1XG1N1foRJzrZOIxDfAiS/n5+e3zV3MJg7DPdqRFXS0quDSln8YV09zyHeL
kcKh5loLX7kTjBlTjjjRYaK8qbb6vAGfMi7U0bAj9KbjrvYQmyya0PQKiFjoID5Z
LRCqIoYHS4qgsmsgfOJi/xJZpY+GxmYYWOINIy7sEb4jgogHcoF5Vto6ryuVkgYv
ckBOPK7m40JdztKQJPDOc/WpB43QnNrqT4k8GV1C4cCzHpdK1Xfrn3X2FgK98Ly6
GBRL8/qmmFXBMDAUGZ9QiRF5rmBqOSlM38XFnh7TPgspya2Vw3a0EVXyH4nUwiji
RKZxG40FULulZ+7/o3y37xjEKaoYRo2sXw3qdsNFUODZXfay0S0nHZktG3UO+Vbb
MbsEzSJCU7t8yieBjp52ByMgXGUScayHwAzsj3PqsQoGS384cRsLj8wb1b3C6/Mx
BS1uCeIhLm6i38AJCA/MkvhTwJ2h9SSYYMij2q7ELIN2ko/03bzW5abwq2dPBjNV
kBOa413ea8oEWGThG/ZSPvFq5eM9GiU5y1+dWEZ56ApLjkTCtc2QQZOGd7cYG5wu
viV4zf57cVj5nm7WXQa/dpUd48Ea7biFTQ+FPCocNoYh9mnAV7/bj0jLUU7bSjSv
bfWSGJFhno/uhDnYTDbkx6I+xWS2yJ9xVf9GGMul8cDp2Ta/w/yqdouvD6lTVMhr
KITg1dBukJzmoqUYCXkJ1KywnJaX6RsrCUblrTm6C9mjdGCXGkHfVTRAjPdxonYP
sXQ7P1jbBpi5lJ6O1SKBdHU2/D4611GTLQuyE+2X0NQfJvYKTpB9irQmHgLynH5X
kCOdUzxZIC+xc33Ly8x4YPqEBO1mKJC5XjvQXzgWun/cOQvEUAVPVyuoJNouZVxv
B7AoVej0U/EoTwQt0THE/yY/C2b+wIfvBu6nwwNKr5WHwqWrcB/N46slqp7MC9rJ
NzXEHEr9s076yuvEqx7dlKQny2V/5lSUSj1yq3Gkmg7IS+7Y/qxrorrHI3JtUXaJ
f4CxCufYkFmOkEFpViErCa35aIk22U6rzO37ol79KmJnoZLiODrOtkCNNvQn0Shg
+NT/6wOLccf1KzQC2+W8mJzYyyXsH82LLG62h41Qnwp7kh8eWxSIgO5fZqEA/v47
3+LU4HDmZH3z3mffy+d4YPDZEwTLCiJxDk7qNwV1aXrytm45efHWVqdV9qrmn7Fn
c29CAaAr+V7CaREEpttxsnAKipEq6FlXAadL24cbPTnTSZy9FekjLlK8EuIFtQPF
3IqCxjm53NKnY2Ec3sndKFrRH+Xp/CtDQnYWwXkAqHc4RbKTmvsQ3e4pfOjIzAHb
Xtcm+c5bdKQPDEz3Qvil1dgBQ+rGr5yo2TJogaiNTe3rl2hf89wIpCCDBF1K8uE+
OzJXkVekR6EJXGHJjwYJpxj1WWJZiqXd3Qaaek2G/cHcXAKp63o/J59BVGQz1PBv
n9vV2FrHKd1i/hHgIyq4qZ+QVyvar+iaIoZ3TfUbf5ucsfvynwuAT3RZaARLjgB6
o4Id64r2Zsn06v5JX6Lnj7Ly9ZkyNtJ1+xCZex8SJXJWUSCCpQF7RsguGeJiJkMk
wR8c+SO/7Q79VBGCGom34e0gzEKvmgEYpHz7d17tXk8xcth87gAjX3uuAPXWw9rQ
m2bkyoi01fxe1Q3K9xuJTyFRyWKKN6/Y4Y+vyt/lLQAQMDLTavx5nl7amoA0y0xb
kpSQZj6VyBuGCYNWjBL1l67VuwbsebjUmyDq6F5MjAVIsOaK3cKPfYj40UnTWyyF
r++82y31+YXxyLBG7hxRG0eMS54RvbGltvBWzQHSCq3S052tXoUVSQJyG94QkIvp
+glVJHYm6F9C6Sm7fs655ojjOxhm3aBcfraMY3QgN61OLTpRPuHbeXazUfSALvSM
0k3H4vUElR1Uc7MO52KSz3P51HHjyuFAobY9rr2/tSBpu2VeFzR1y+wb5JCGMgVZ
KPrV50CTM9Rsq1ujLmJElKN5YxD56LIBWWELCvEkxYMVNscRi96BJoWqxI73vRKX
LkOb3HHl8MZlDNiunbYBRYjUfDbxibSrHRGYOz14fYDh9iD08jSCVHqrWZaFFRd1
sRA0Kcno8z6zaOeCVPBZ7qE76YHUIF6MjymeyTq9BTphsMAYiKEdFseHuym1WQfM
9PdzuL3oy+fjq+tdwSnYrKarbKY23pZyOUdf26z5DHXMiH2EywwM3HZE4GB6jZtc
Skxc2BScHUKwuiSfWERJyMQJ8I6N5x/avYcPH/YJgXo8hdH/gfNKr8l8BMfK2W9r
g2ucKeuacKjrj3Kr/gix5jOD/ErGLgJP9iNn1srmO1kxMmf916ylVGr4lbhwC+5E
upHSsDjTazFngyYr8w9jeR8yC6W2avVSch5BM+iIaTFpCjQEnmmblTolHbQ7JOGw
2GXESkPoYaOUudgFa3fUoVDAOR5WpkcU77mV9d0KfBwna5B4m1RO4QczXKjixwmO
fXCJSk5PRg57R77bUM/IJZxhyO+uzqlfqkq+hQ95UqAf+C/CEFJoQvJsaFcsdkJ+
Cpldz7O92BcysLQBcjg6zPGIaHQj/l/l557oYK2VIZ812ABGW/gd/Xsr4m0bY/gA
GFSiGhn9qVukwSq4Ep6LcPGujcviNfQi76/YNq7qol0yS7AyAhZMlH0eReC067GE
kYJQebVNi1cGQuAPO2XsQx2hNw7ohfVRWCgk89h7Bdw1+kjYWXHTrkzwYARiBWhD
A4+BiaRI603kZGwI3cUWnunIoWnW4xFSRUwgcVv2v5fNogLZeXpGMPCayrZv0y7F
7Ie7o52hyJwe7GCaai8pQGAdBkExVzzg77ZHrJLPzCvSdLIpgAbuR3yrsV98m+Rk
LqxvXWiqeg0uKxhNtX/GTrc0Sxke8KfOIb7YdMw2cNk6QjBRfkzr0v2hPBYVVQK4
ERiS2gv6tjwYMnoEeyD7v6ZLvqn3ZRrfaTOujNIwNXq+vDpBdVj0IrzrjxN8tR/x
J2Ng3UwMIHo6oQHeqU5oqP0IKB5OxJZM0vnDiGybFUksL3OSdWBFu/TScnHU65RO
WkdXKEnA3swBYKuvlX64km/4TZUmcPtKeHL0uiGH9LD53J00FfJtzJJrkSuLxQwo
8l2xra0uAlJcqc8rrJm0GveZp8m697E6ElPPpqEU27eAnPx2I2uip/09g9gK9/14
c9SfOIG88Nz6YBJf6yGlDxBsYlEWyNfdYB1cwBt+NN0ujWe5O/XIctBu0ovAYpjE
7IW8wFtoDe7Vh/aUZZykVsUWj4rdlJBvrISXDVVA18dY5Sxit+aXEi3qLA4nwgVE
N1/o0tqkodAT7kV1S3rV/VeFUhbem4ZS5t68t2WAxyr9/wgqS8XHJzSVUaoNwAn1
5F6An6RsAvBqk15hieqBSX0JT8IaTOl1oF8Vqgy73upzsvDxnEG+fYM7g33o6Ujx
5MhSN3qKjTECdRdaeMepAd6m7Kc7WMNoc+n7/SEjZQNCyZ0fE+zEOrKrTcGaKU8K
TsQQClixghBe2q5GSiu74gCho79LuNR4Glg8QgKSXJVridOjq5XQbVgOMl+BqsWZ
CkEfOSi3keqbLFD/V9dWDjB+lW1KgchwK7SNmGUS07PrGjYG1RZEdmT3T9XDEL+U
gyf6lT3xF98mvVOGXi3kcBiiL6PF4Jk1LCzOQUfubDS66repozhbD6eM77wHzqpc
32zPb3AvPXF6FdF8VDQQQRNgA/ATyjxtaJ39TSdGqwhdIyOh1+QWSOoyOta3+OAN
/FeysklEsQK7Qntdbkq4ePq/Zn5R9QxTgHpOjaqFwcu22UpJFyzIF4nKpofXefdi
i5ce7q6NUlTzQkFok7CM+i5MltysByiqQVBemjBJsn2dE5nyDL8SWVE2OSoGwDjE
bIKYc9c/91xOrzzBvh9XMdLZhAj1Og3Z1Qa1O3AmQ9GNZMzZbtSAstMsz74YW6xD
8DeJUMk1XD4mY4fCMJpzLf3tq+1VG/iUy1i7akgwY20mSJOilIjeB6JOH+QcT8lk
0FeomajQRUPo2J3ahVqdW81Yd6ptBNlTQyQj3x4NTtFSFxmnJxO+l0vyh4eoclf0
CJNCEdZ0wvD9Uiz88Rw+P4wtEfFJRMrKgUMD2IjvXFCikY3L955/MspA7uTDqeIS
WiqD0A5P4W6LGb9/+GZEAc4FwH5zwx3e/8WrF4rYIbjQkfbp6fMZQNX5ZiqQOJMF
W848m2FkZoCw5+xx+CxTpgejM6zqc+jwk3vCZO6+Ar1fyH0kE2Zzc2MrRx3RKxN/
Jna1vyfUuWnJfh+Os31LiB7Q55JuJ/BAN39Lj16yedP8vA3zozTr/wbqXLo91NQm
RAtfXMssqDalGtA09LRPbRvO7Jb5pelctBt03ydwyWDhyHTm1nZOlZ3HnLIOGpJv
gCINUFBtPb1AWOSZkM9ICueowgIOLVET2iV+XBwJbHSxLnQArIqwWFUuWQEyiNhG
qpq+9oH9RZfpL77sFj4x8OpHAUMIIrzL43eyWQV3hE695FoYl3oftHJ0tIjiPUhL
VqWtgVtz181EeGhNn0TnlvfB7nUrDOYNmLH2VeuYfdelwdBJtVqfsQ+mYbAseNuN
I13cxPGF0h8uGTUXmKmHR3kKEUwTV7fEp/5DnLcUcmmHKbZ2XqO1sl4fh9VkBCk4
RHvGoEVmxc5MuEu8DUyzqCAK1bgkMrscUgdnza9XkzcnjjD6bzfW98Qiyu7g5Pkf
zuPiGvTos6rEIG1oNnqI4yyuF+OzThQIKTZIZeBB9a/D9who/M6izLn7FEuXawhG
0YHDeNQ1qkjQBpHkrnlN/dxb+hQpaFHFVjTfiOO0Yh0H7xWaUTI3p4ZGGFvv+Wam
Hd96JDmt03lRTZT3SsILbCZl/KMTdPiMoAMHB/dhtGlQ/XtCN66THDMlJ7utqqXq
fwORvYIjI/JrDPgf6t/7pzXRpQDZi+whksP7kiwIkIaO/jEZPaQrtBhcn/RZiOan
YV5vEkXTJslpM470yO32K179YFrOKqZn+A5eYOQZBh8Py2DnVcGKbUTQATGNWe2O
a8Izxy95FIwTazrvdBtByit+19SkCiYp/1FKeW7rP/LzK928H0rfB3VBjiNirjm3
1bdVyq9jb/DJ+vIr04R5oxt/FEWuxT8xXdMMKPHPvB7TW0nhIcmpcTyvXPy9cKzo
QftyXEhvrjLc1GAzLIXWY4fUT2vd0aYKImLDCPX772yojlJCgTIMGMDQ4L6MSyvF
XjGoxZgTmiKf2WIziWkSF6+w9gs/Qve3hcDD3rflEhzT2UofU99fj6FJr//rgjx9
LKYChXiE+mI9O9RYeMHUQhwukumRELNxU/wmBqs0Tp/qVEEsEpbIjGTsf2F9HPmn
DO9LpgHJNew/KkPZENcLrPnwtdwG+r77Xjo+Fs9FhcwBPhUfVB+pJ1zOeYGqdyJ9
g6IG+DQuhzROCyoYPBebQtOvrjrYekf5OYoIb2apB8pAx+qn0B1BoMJgbo0On3o5
zuYuTSWkDpz2LRZrgncz1oM1a5CE10/DNus9MRmOzj0Pc4QC/2jlcybgo0WBQtkj
Gc4V66lAk8ijoJweQ7BvXEfXfPuGeYI4jKtJMaGnG1l/13ag8R4SlF58nv6LBLQ/
fO4zrNFw27Hh6fFgkOFBZEUCtGoBNVTjJ0aya07JR+wwv1CK/eWdlKMCShqu0NyJ
fpb9i+/cyzgQ6uoodV25Ft1I6IwJyAtg+FY88RFB4TDS4ySHKWp5MyweByULtDNN
FiS9e/wjsplDPIVFglhQY3i9AvzvvzarhL/xVAXMNxKphevINBnjkbgAskd61W0l
pZDl1AKOhhvXtDKZRa9vb8Glyr3YpXez8PKvM5/9lqV/VT5KaiLVDf6v5IfD1P+O
zE5OjKqoeFE5UiaGulcbb2YOtSOkILsY8s1+eU4SSll1vmKFDzvPTk2r7Vx7kXSl
Bqr9sfDUUZxEJlk3cWvemyGbbyS5q7dBcEYERUpOW19zfOjiy+PKlomZ3Ww7oJYC
KuBy0fWYnpfx25Ny7v1y9/UHzbwt2AwkcPPlWeWs2xrEaGuQ1wRsB3W8ufhOzq8l
VcraacvTz+KHGktRBMzmD3OfOmkZHIFdkcu8bu28jU8rzIxeQKvrJnVqBdoB+wsi
ZdsCUgUlpXu18YP3LufKcRk2nYwlp2RU0iinTz1Hlo5HK5c7UK25HiW0vv6ar7uk
w/nksWSE/ejVHBSdd78NcTMhQqKl3c8gqSl2XhonCz6aL200qej3ZSR1fcKKEamr
kSXhjld64zc2OT7M29qTcLUyl05qSJmARUbfgJCzg6nUVMIWBsaNOmJAMe3wnoHp
pBHrU1sUctp42uqH9FxPL+chRdZc4NNtf+4eYt/p/i0GyWvlr2x6KInYO6a1ob97
MqjOcoG8H1mG2RnKXCCacP2hRJGP75ZSqaWvpk4+Cp1x8X4TlOS91lqV97llt5vq
9N1TRI3C8aTS675fx93RjOxNiNQVsOoatTOQn3sOLEMtHmUT1k+EUcaetU6bGpvx
eTaGW9yfdvbBBROQi0HyKo1pkyo4vEes16tzvsncEeGYuC9qqjnJfO/JzA7o8xzh
CIPd0Ge6FgIdSMyXn+f/wVAVvH5tuNOU+lL7AHIn5Q06bUwUsGgD730Fh+qxTNiE
IxpUuIxQIbQVextTbVESE1dHIkA0Ujx3rjbGsp089cADmINYjqr5VFOaF6mM39dQ
5yqnmvQtGLFR26rd+RN7N9HmjaXQPfS7quRtT/jPflIVWQlm0P1MuKmERrLGeo5/
qlob+v/JZP84I1T6dBCWYianmEd7VFovgUT6I0FudeHo3RqMae8D6TR6Gt2wSNoC
ABHmtU3pjW011gtjYvIwchhRfhiJO8xtKTEkl8KwfM3PYVqESrB2qAs1Zw4vaAnz
cL2Zy8xtF03Udkm08wSosCovZDicNrxvRZsPPJnkrs/1tnop6zoygIvtnFyxzZk7
q6oQgWYwEeBwT2f3Tm4JNi1Fih83g8OuKIKWaNMsBHN/fjKvjDh8qJKOyPbn0cVt
9lCCe+3kCuoXm8ZpxIkOfRP/EX8ujsVmqOeq/tWdUnNcA3ox/GodsfX7xzeF5+W4
zkfffw0bnK08ConurrfYDdivUrDjdKt9SuROwIHX9bC8Sgtw3GuAUlxI/flHX6cj
Lh37PXFoFdjWUSelcfSuqSA8GW3jgoZMk8VckP2yJxlL4PVBFfkOHaKgR1+ejwU4
GA+Ie0kRvIx6/A4JYv9mgQofNDEIpxiyRvgzc081CKb1uz2FeokF+B8N0EmsDHYU
x0nO7ulNXVA+4qrhOC0ws3SXrmDM2WuB7/YGbG/OUOiBx4GN2JQEiidWphRZ/n3G
hGrFwTzzgz6uEiMbUfBwFJ/FdJN+HrDWVo8Qq4ZAtbRwdtyiBaDRoABNnXCCEA+U
zw65bpcn+2rKhr6dBrSiR8HnplFwnfQI7YjikejWQF34zh05fCXxgubxpWJSDc9M
E7cYx70pKJFueDfkT9K3K++GFSZyKUPVaIHf6NQzT6XgCH4rw3sQdQfShS4Yu/2v
lYshPmPdQRPgksCULyTgKLqeQmjAjZ6T+qHlPtNjbG2FS/OEDZFitATWfu+3ew0G
vCYH3l1DqDC8QgQs2j3E4/p6iHVVMoTpwF/tOmhC4uUtGVuCLmaXb/NKTKsIqe/Z
j8lHkAaM3DH0ide/dVTglgg+UKjcS9torPGaqFnjnst/Ibvu4LLhrZ1JiU2V4BhF
UmYj4cO78W/XsWCXcCRWNg8mu+GtSgMHSAaOr6PzLXm5ipFWR1dd8olbzqER3YMX
C2RD28ZCI6wT7CIVxfHaj0wxw6DVqSaa1hRo4aIJO8A2fFcIqq7TwOMtlNmKzRX+
9D1Qe9IxaZRwbhP9Cs2959rFaGaDw3R9EUqW5o4/Q3fmKSJh1A1VNClRsFCkV6TS
pgR10iYr07N6nVJZUWiZtg3tKu9JlT6J0kipL8MdPkLGBXzgRnDJoj/wnt09KGsZ
Y8Bd+rfV3y8FqgeWmm9LvPL/TcEKKfn2Dgy5vpd7qdG1V4H5Ct+/hBMxVWcZDXq4
WNlU/GqwEVMx9AP1bbZuLVC4v0EzSaaDmf//lRrAH4lp4QFFcn1Z75pyy6/NYbO/
NXbKSqbluhqD9eiddh776reQEDhSLVsDMfiQ78h62A9UYvkRvyMIFKv/bkBzWvON
jPM/lbkrCta9qmQPqC2yzFpM3/D8IroCgwa75XZn/Rtu0fnLAL3yfsmZTCPylkO0
hjqBHzqffDGKl7ydyXUD4+xzOVdO3RXHGQ7r2hwTc/yEW4DxfzKS7QP8mBa1YDkx
jwBGypAC2KkVIRBJeYznw2tZHh0pHGcYnPPBzZGZh1N/Iff7k6glln18Ei3ToNrG
9KEIycXQ2XLkCDBTb6ELCCx6AffhD47X2MhjdeFwjQpAvSV7D8stho5Ffqpy09CA
EVrz0wOSSqUzDIymZuMHJ7Zdcyt0QqUk5MYtbqj646oLrKim3w4RiRms7d4cL2H7
LXqA3DOZKPLUBNYvqsNa82FQukJXtwJr+7ZFWxQJSZn3t2tKIdpY74U1zR2JalI+
2N5PLy+tdZV4GyCdf0TMkJycn3HVgr2m22Lxns/FEPpG+rUccw3ZhN/DJ/cla8hs
R/FMDriCraO9SKBsjmkOozjYGr+4p49q/bGbzKlAdkJNo1EK08KvrDy7Vg56fo5v
g9dkQu7HZkYdMtUyj1xgJM8IFwBMpe8fc/b7n0//94+8Ro1cAKBM5WGS16IokcCu
O93rL1r+nc9h089SKnJ38dyaF2bBs10KsalvPwXQl/DIXUysNjmzm9PKy6q3mRzL
a2oP1wUaxX7WuyC+wIHWwDj6lj6c4VpE3yiXb7e3ksap1AxFG0Npb57p4RglM1pn
vd8e3oWavXBy9AfCQ+3Q2I4+oCXVrUnBAfgoJQNOUkeD+tOgGID7rA7HDz/NV5FM
jcogdJNZjcTkTxBtjTgETdtOoGGJHuB7r565Ap001+RIRX70P2VWr0aFxiVZL3bR
ESV2s3HU6HuW+L320xqFyz8yUE8ogUBfiqmcI0JUaD951Pq68VehQJRKuxxVMKgQ
59lsrBr3CxZLFheX7PcOP+gmJ/im37VKU4iK2Eu/6KQJK4X2EOXpVjGVcW8gR4dh
zdsdjwTpfYdT2YziyX2RxBc0Bd1Tdwa5ERzCChm2W0n9cf+yGq7Xk5Xl166+FE0X
etlSQb9eXpyvollHYFAE7k+l06Xww+XuXcFF/OiTAZALp7ZkGIpxM0zYJIagOjen
yHkp7QcLIxFVu1lqqunJ8ziPwhiRZFCixpkS66qjTcQ4Jk0U5IUF0BYIEOjobRSU
GBIvQcwcBAw3JambAgrHdXn5bS9TxErFJN024/OzIb3LbMSnfN6E5mJgVVmO45wd
gdjev4ZPbJUvIFGiC1IeSeySgNvJRRGotjHSJnGiMzJcTLZ/RGoRro9pEfzaowsH
mGBin0sOm21+qrIgdCeOHIcj1ffKiQMLBbDXY2meBFSe8+f8ZbK7no1AX9tRtiXA
HGyettJWGNhQ/WsCJQezvpmt49S6UmcOsIGT1HiUg8cVGcdNHY8simI2JJdgwob9
QHqW2Lvq+gyLHysWcSBJyd4bsNv8uXBOERIS1EMdnZPz39RnUaSVFMOBJkmwUkfJ
oX1fSMnNU3abpFgZw1tQy5/q9EycjnrX0OJJzMaHrXgLpy5L0Ri6NV50XQbsOSLa
4P9CQeoRER/9lBWn7ule/Bl7ZMXF7BD52J9GFC8g6oUdqZ9da0/3eCSHMnhoNDCt
JwMX7DF3EIyXzFvCGSENDUF+Rqg6k3X3AAt3lWfj4WwwOyrBaowqGzWjpHR9KH9C
jGo4ijROLHooOOUHQsLyoxd2tZSC7dtPb7ln2YNuT6u08RXzNnaYKRKGXxvGW4jf
NQjNPggVfSzAdw8mCk3LVfCevIlBcztzdShGCvKFlEM7Vk4RYUSrlGrhnu0isb8e
OXJ6wCjeqUA1wWomXvPBH9FTVKraZs/+NtrUQkYqR0eCcD+qsITcvIzIucyrravA
f8Cuv/Xnim1rIYvNokmR3FNy7bWybBCo7D994EOhU5I9OgA0e9qjlHVn9XIvNEBj
vI5LjuaXCi2U5ClSQjKjPSzZRGGHUWtMk4fAC1ehcg9cu4ceh3Ny04qhxNbyvIrG
elJ9vJfxYBPIte7gTa6X8f59tLyDSOiVUNRVD4oaQlPAJlHAvR5Gk28Efo7aXb/g
oOdBo8gQhcyV1V0B9SesD7AR1TVkXtoK4L1QRw6bU5DppwTHwikUXv0uWnl5SmHh
LZCaMp+/W0Gr3DpiDPj4Gu/zzmL7aoY+fkgl1rcxZQeRrmZub+pWkT6H3DSpzTXf
+cp8ntxLciTc4CD2xfWAJQL/3u9ID96UCiXrC/djYvXJnIhz+H5cXa0wGcSsgh69
nTmhevEAQ3mFYqxag4gdIKdXRF3RaBsAPFyuNesf38/mrfu5VLwSXKKf6SasfJ/f
fKmdLT4JiJ9hgmNs7PKbZjg5DL6iX6yVuO5YFSILXKGbL3IY93+2pRiUltXPZ+N+
TlhqQpZcQ28hm8JCcd6e/gre4VpQQE7obsXqVRUBHObc2z2EyU3eMWflNJetGBYb
IXuyHca1ojqtLSpWTHDmeShUqfqVNml9UVKjriTviP2vLae2r+zmnXxHnppXPsOk
a3YW9N2DzkqsqDL1JV+F4lkJUSXKPSXyW+AWDTVBCsW7qlTseiQX1SqZEOKCmI6R
ME4U3xrYDp9+vKQiW+M8AQAc5QeLNpKsty0sRcUsxNC3zUmnj3WjZrZ0jWZLnpmQ
JMjIjuE9wl8gowEzhrbSE2BUItoBS0+0vZlcvlx8gCeGawTIENFDargmbLwMB6UK
LBSAFO9qM58hxpG9TfeZMuwWbxU3wSnjKtxNyv2ZjxwdBTRoLA8HHTflR4bg0SHV
vugOtnI5D23uDCleMvZT0fhot145HqUoEl6t18qTkaszn7izb4FIk05g5sGrYuB4
Oca4NkP5XmIyW4V5Bn0CZivOgkT1Mo8RRILg0Oly/qGMf67fuBrcC7fjiDEhxM2G
omzUNmeUpbO0+8aKYzmonsSthNPKzo1pKXZpw/dAtXcCR8eSor7eak2AVZ/jgkCP
pK4Wg0/EDsU9OEEgNC3IfNSWpHeKxGqBnTTdasS61kW8btntahiwgbrjD42z4s4b
ON0mI1ZBZMoDpwpJ/x1E/gMzMK8n/94J2G3L8BzHYacbK1fZz/z3299tjJHykT/y
OpOJmozL9jRPZ2DdwO5lTMzp5Pcb1yG+UZVxG0hRy6C+f0rIJKG3dKzBGXYvAOwO
Glg8nIq3S77+44P/MaVMmwLWFtSoABhoE/hJnuusdHV6bnhZUiM6YRYcyx2WvEiF
isgzvvI7CzkMAF8cNvZaTNmtCfUojFsTKjxyi0XItTpLNIFJG1bA5jEZyo3DBodz
kuNBKXpkhvyHrOZU2970D2kTxz2MS35O5usQNmiAMozjrqjNdJsxXZ9QkRccgb2S
oPWvjQIZMPLFn4BmwcuDLOV5b+QYnK7DvROiXfiAwQDsXMxoEK1mGlBY0vwuoc86
kO3FkYnqP60jDEFvgWHYfti8hdsxvYVg9YkYaBe/7G1PmiT/CUR28FaQ9hFFzp+s
44D5NgySSI7fxlQ1fwwx9RI6b3NoxKfjWJbGr1AgmQP7kqPu+bdU4NkXgx4/+Yp1
zH/+Ddcg8D+lGEsxyfGTFIBS/RUSIkdSOCoOVBQof+rNaIhnIdgydvAskL+UD4Jd
Bf061Se5zM58NFEjp902UEQ6xGPkD8oG1v/keHJKj8IvJWxzp+CmDVkiS86P8gLy
CbSiksbS1/VVYnuZXt9UuM+StTMYaYe8Zz/mP9qFA4//5oxoL0vPoz70/ObFMB2S
BMlwEGKnppkC4mYQMdigdtlmpgaQrprwNbIOG2yn104FRBzKdSR9XwARIaS2h9e3
Odye9cuJEaCYZCX2jBuptlAh4CbOHwH/YNAgB/N2fxu/I/0cywnKh35tZwMaqypP
xcAsDLTm/F+rMstq5MKI+75xWjnaOk+wWvSJlysHEcpvIUaG8KqmTlAeMYLA+Ost
B/akKI7rwnY5/S8gywg6wh+Tn+1N5J3jHMoHXsgPw7kv2StWUg38lSmXzMh0kC9U
nDMNEVQy7ofSetcLHNFxGvYOkhnExH3y+jPGVU5e9OACHOO+80xETLupRsJiOVD6
zr4L+kMhGVVIlE5PgUbSSNnA3fh1vDnOPFCqY9pR8zK7fZOn32HnxZk/HqVz1sMe
PgpN3QUlwCpoi/8E7SR3OKYQDq1HBMYJ/9nBhplVXQ/twuEwgU0x+SAN1L+1IhJJ
zmSYSPshSh4LOUbynKJboVyJnPnSoXQIH7meqdC3+uh5/jnA3WjXodMB1Zdwp02q
knKPEwG/oFJCOfPfHJMQIf1ezMFnCoQPDQyjxOpLrLXu7HzX81wCvuoF1GKnkbm9
cMT593Y/X1Dn8LveQQqSn/Gkh7fIJhROjPmTGJBM7qDJ++L6jmXKxFE+lqghAV1x
tMUgwsKw1QzKuzKrU/hibFcgRr17aA3vkP3hUALVHSESp/8xz6q1geslyH1zDc4N
86YRg/CJM01Z5KOM7M2m+POjozW50KST6Ep4Fj+GgT44lKaWsH1pAE3VJQ+rR/Ti
pxjvdKEsLxV4zkG3GbLGreRHtTqzDA51rZxeI6NCw7o+Ro/LR+AwQfXzV2Wkabc9
Bjf0UT/nswub9mC2wGeNkxRn5/a7f5vFhV3LlxgyS+CqFml+J0qArxnDoKyqVvZM
rac8BhDfWk6HDdG43jii7lIk7EpcMgWPKlihJN4WXdzDgdY5nxg5YHT8dYfozIcG
D2TtG/KhBLJ/lGMRlFTRd7kFosSMYwL5X4dO+vDuz2khWCH+IvwWL329FbVtZgln
eHkLpD6drtjWzYw9MQBXJXiN3CdWTFxzkB3DUcy5KzjZeyCAq98Ho7fJl2PKZzkf
G1mtnmw9TViM+pVYoZPVEDVnsejYzPtxY1wECz/LDNAgoZmE+J2VVenkljDcfwbv
fKrDh10/IH6Vyu5N8SzoZTy2xGP5WoG3AolxNCBhuZCa+gkPAHL/LsD690j6S063
CwpBfBG7RN4hpbI+YagRYQwX/05oucjQxhagjrMv5IgUMnbFUtQgm6tcG1a0ogax
1KnO6OchuVFUJCjawmN4fLVdczr04zWHwSXJaBVh+SDyrbBpdB4bQ7r9gxfOGRft
A0ekaTBN6ztckzWbxC8gjG3WApF/XIalZnpOGAzvpRBmHJLo99VGvBIfko2DP7n+
Jo650nzu89GHMbgErvIU2qT8vpApNpPGSYjFFdsZjeR6jXtByoma44AjjEzR1PsA
vfsx/p+mxsJBQRzvf+ozwq9X7aXRa6TrJDeubyKgXyIG5ZNii8xcwOX9H9ETzA77
qhMQhc+drJuLNwG95y7HJZVtoRyZk4ojsVrTwgM78zzlD1z1StbWfxBkU/QLlosd
AD05iYn1ELEov821U2cneRsVWY6FpGBmNqB1xDnc/lyRpycmacSnh6qAZSfsBOpx
8u2f3xvz4Q0MpigE6BacMzMnYuIC1wSeQcqZZ0lpdwWSfEsNKVlanqqWEXwq/UhU
8TWBOoIononvThB6i7Km0Be2RMrN8HgRLl6VSHas0yQ5MvwuwR/9vW6AwaqB7Sab
YvBA/FQUVABqcsNXwbR7S1tUaK2sGopEeBYDxq15Y0UuDV1APBXb/DStZLTwURhG
Iz7q/d5TzTO/4CZDXradWI7ZK1dWPbCBsUK4Uc4hxcUDGHbT6xa2On7iR+6cMBIp
wRq6P9h3WC0Ed0JZF/0M141ukJx80KCKXk6eTSNkqFK6H7Ct8OqI0BdW74s9egT5
awxXK46BQZFD3Lk6Y83/n8MkiUOGn0k7csdyO5e0Ohly6CO4zVlCsuRAMiEsLzU/
GDgUB5DfurTxt2AVfAmIuBwlmyZerFCiEiMcw5w5m4FqgaV70b7z+TPOAmK6tkYi
8dE0EVmEbj3RTv3AMdDglMijTyRZdako/cPRIX9a306ndGO6XGj87GeEUnqRiYN2
YLJxhkGgDW2YfSXeypaDXhVQ0k0e33wtiAx1RbEZhtZi/wtwr1Aqwknp60LYQGpg
JtWVSH7W5QwIhZ5UoYR+S46doq/gQaCnDQkB6WuPmVTJV6KqaIESBcxMxaKqZDDZ
YSUkgBtvCjw5fJCUfHp4x5lGzuErn5Eds6XGHNXrEfB4Mj1oQeCLAi0kEo1VxJC8
9CA0WEzpMeqv1+fty2Cz22/vvjcAAaqkrzK2q0Go9/NXxOU38Ie6am9T7BpLK9U6
FSUsiSwtCj0cwsVSXs9B0lQJUqSXKc7FG4R0fjOm5QLwtI/zR2hCarPAkacp5G7T
CjmXuLgghdMz0/5GZrYMSHhzOD8ZyunArsOjFPuyQI/I0g/27+0XC365bqT104fz
jd7D0bHIg5bG1dqSBKF7AifCdjcgkjia5Zm/5+qv7V3YE3uEieFnb7KFzDMF97Q0
GbpvrRYzw2yeGlRm95Xj/4x+W6hJTNEMVNFHO39qsYJ/HsuadIhoBZxzed77VvQW
y94Xy+i+51psJlhjyAgQwJQl9NUwEwDvkAmvAAVdUd1CD+1n7py5UrEjtD5M1gj3
7bV4zW70ZIVZKeXebGj5qYzMSABjs4aQJ0V7BLkmx42odVFUtSfUO49jz1CDgFlj
mvGKZBXW6Ra8dbtl2LH/qNjsr25LBP9kYtGokGjyCLEJ0es+S4SF9zWX6wRUgApW
1jLna9Nq5dHtQK4fp1mwwccCHxmG9J2aAq+UUWNKJNd3mmYSlJNJ8eATVm8RLveq
kEs9ioA3tzQR8CrbnPeJiqCHsyghAoFWBhI540CBgGntu0hBRhx6+iZFsGJsmamx
dmMtyxe1gQHhknssebpZH9dffdNxXW7Pd+uF4Co92yFEiE6aXrda9X9JWxhyCazm
p1HcMycbCLXuMntx1wxQSMtBngdH58kxU5RjO1naPtimT1yLWpJpCiUtTNB4XaQx
KvDSeMjFr0m2agNDrVrC28CsoZLRnZzBhU32BAALyAsk6FWa/V1KrOupmTr9rDyL
B6pqDbv3sx3kNG86JGzgWg5/wT7Bw7H8+MXMDLCpOzEthMtPvLt0rgdL41NhmMpL
aVAR3rWOtf18Q2WxUofY+89tTgwPlkwE+tzA2dVR6if8FnHOFyqS2+BPngHEe1Wb
iegCM4uNLQIvUIOERNa/lt4c8wlQTki6oiWiJyNIFQS1Lz8NzIB/j3fkmhh+5jPA
w44Y3DEgTYWRve7exD/++abtujgAMGTINN93c2dGGswSUMkyzw/8ZCybyTv6917G
hKMx6Puz45k9JIJE7bY6tq+VS0czcuCMAmeODBcdZLp0L2doVTh6IvaPPIftsGgh
NVBGGT/pIWo0526wtIqQYMvTrDfzHP7y3VvG6ZMse+s3mq/KwPqbn0VQk7DvsVfl
5+nO4bcC4CXG4yr/8hV39MtusZ9ooM6qIqi0+EaG30tGdT9gWCNMNpLCVIF4Eehd
i4upVHRwQWXYa/9N6/3ZVaF23lyaiaXeZ3iIbB4h5Dct/QVymPq4ktAwtnuPUEdP
qmtAbnIXq5V2NPU8oiyMI21SmiaxR0j/fim0YjDP5hi45cdw1Gkt986Vo+dV0j9Y
pyNwbuwfDlDQr2vQwZrnpecH9KVxSjHQbhY7g9+eBAJkSdqOpOYvvUge3TzY4kfk
Bvzne8mngbAit6A9Cs1WIpLc9faSaOCs3EHI/FV0XMEoYUWWC2vnmVJ8qqQP4wkg
ezUA3JROUR4TvkFQLfuC7gp+OCMAzaiMOvvk/V1amyuyQcZhF2hDzWFJqEtAsAJp
wGO1As2yOuoyteRNUqYoqFhab4ZFSr1CnfNNGlIjN2d4jo7+lSlQ37XL+7dTdZYi
5LiLt1RgbDGZ33NCgENsc4K27E8v++jsFwFjYSl3dCiZOO60Mcjg3hxB/bqJMfzg
3P3/k/HteISID3dpqqYXEyRiP0z5OS0d/2GSxf/8x/fURjjqfd0dyrvDjf21zjYg
TlvDDinOvC6HnmyXxaPmLK07D9TR8JJ1c2o8H7bdG2D5C7Mnb3IZmNMX/5d44Bol
NqQ49fOozu073PFWLgmK6Vy8yGc3gL/vVw1AvrnBrXxMF5CMgOTfmtOdzMCXBJ3P
49+vGx25yp7ZPns6pjQBZyFffj3ADs9gHwwxZJ8wnFTrRKDLIAQtGl7SGwJwbWo5
WULy2jcJZaZVet0uhXFZjhEXQNabmrNpDvb+QKoL5+AVysFTAyDztQKAzsKtrRGn
LD9UELSGZWrk4dk2keIRYuGMWJLHIBy5iWHtCapts83NUQLvDkeXUfV04a0MUhUH
EddJ9IUp8LaUtbBfZsdaZI9rWA9/1LtWV2HplObbJimhdIZCiEeCVIIJDfD6w2AW
oBLSmOvQk8/iZApztUpYXz+9PI11p4L5sQko+absYwso9dS1Glf3x/ArRHLOxFNY
C3f9ZDYQy1UKlmYzFSgJLqgS63mOIm0YIlGR4U3MRXz9XTsrJ6/yEkw9V+CCmLox
AyWbiovRrVh44BRNeupgrASwn7vPp1jCIO4AHuGWiRM5L4/4hmeki0RoqmWy9Ezb
xmjT+f361WzP409GP34UEa1lNLYrN9o0iA5Lzr8lMcWzfYwSuHyG//g6LKEAelFn
atAjvriGPo5SlVU5sc1A1RaAe+GuCNAFsHo8FyXFaOblRoux14NDThMEIXHjcFoQ
FBFmz0ZrxrN34Y+m+GZD4CXbC2QQJXJ47tlMSlU+PZlQTxuojIPqAmiPSsEL9HZ6
CkhC3pNvSuwBIJq5sw0//Fo+MpCI+zD7Egz3XX9oD3f1GPO4CXBW9xQIIwmIB8er
CdZ4lW9/BprqvlCK++cMVJcbx0A9/ZM+ignxkXi8qb94BrRhuOfB87dTsHIOw0zt
sAD7EabiFAp7xcfwr+qaTU2gWTos9slvOtESgS+pJ1HhtXfiAz/js+rBs0ocu8Qk
jhCdO8zzsptobzoqIYwvVKfLvvHu0kbJeBmJD1I+AVELXtYgj1P9jRw6OvNnpEdH
waheb+Jrdc5GOcB9Jqe85EaEacXg8p4qAkkw8eNKcj2NHgZqKtEAMUDItmj4hlFs
spgEE0x0VmyaUPEoSfZmYxt9Yq+6kNgRXjYoFdDfFUe2IwiI/lFyF0RxCL2ueO6N
bWbKea+hT8ycL/E7c1QiJzROnF7KojKSQA2WjebK2ZcenL/W9Zvz9VZ4p6gfZB2y
lljbq5wl+luljzI465xJQEL8tqcUFsk+e8a80TNsFHzcUx+O5QHXZ4iBExwhd3S3
E2vkxWBrWdQUEjxkL5Lm7YfgufxY30h30tE9hwjDIlu6v3Grf+Bs7zJHttRFefPc
B6rXm47eLpmOCyCQQxmgsXaG4svQlh13QKyYZZjDouA1vSSV7KnY/C7XV4NsNG+e
U1MEmxpwbqSJkC8rpn2Bi8ma7EUw33YNHJCF9wOoVup4tGhZ8RF1+ekC5KNeZUgI
39uWL1uU4CrUNOp0FMSNMxK5i7lGvvov2pa+GZjyPl4mjQxhbbAjKn1jAq1OoiqA
xVijxeg/KeIHG23p5vPzHk901Z9h39PCR6e+df2i+dqUF/LBaS0ngkNP2gDHNtH8
uklqwx4Gugw27qsr10ohnM2YWKLQdWBvWh4Wdb+kyOHhFIyGccK0ebkuOyoe/nJC
xJiRGI54N5mco3M3D+v/RhNCjPsNMkJZM98+7EueMJUzAxIfVdzC7tpbwbimtss+
ta0IlbUqPQR01i1znOuqsPLS13jAi2xeGcHAnaj8aFUBJsn/kz7xPo0AyehMGCZg
LHY2GtTX/KmbU3o90WEQio9mD4Py8lXhPUmNJslaiZnbyMOHv5KH2/9Eq87x7RZn
kSHKaMF5duuCue5weoLQWoCm9TJlpcBenMcODF4594DDgj/2HMjHv0MLkMd4Me9t
pdATmXsy45RIlX0TPJMGMXES/N15AtN8yAzracBQueJWgwP/wLzcB2Qc8PW6KxY8
weqWmUfMutepyQGObd2YtpKtu/DXI05ImFRXdPKicnQeVl99ex36TbuIMBRP3MyL
vhgVLOmaIzWRYRDn4T1luu+wdUTNRvQMKmo8fhNubYKaxDAuT3VjdSxf0JpM3L2T
7Ig8y5xv5NjH6vl8Kfo/x1MyRqu3KH6fAYb5HYq9F5h1WHBZI1Fo+oatwfs+k0MM
exapM/KHJFN1oU+CUfL5tGQ/38CL2TXfAVABZM4OoniLmPhvOH7TkHsAZiTBJpdn
AWQVOIl+JuwXMTc/f2MBN0Wpe7x6/dg6udp2FDI+heZBO0RTEoU7iVKKfDEAhHOE
Pj1GNyeLvfD+ClzLCOZ+NY1oBZIGT+dI65gIPVo7VhX1ydyaB11HMt45D4u5mFom
363/RH3ngsEHTzcTN0DUgcehRpomlWB4D+fGl61B0ey9m/bZ6lJbs0EAahYLql8N
8ihkHte6hvenNnbEXhQ7ve6kTuZXXr6CzU7WsCGu5KIe0DF/7fldDbEpmsvDhJOO
VPhX1vK2a6bJb366FqNn3QSbE/f21viz7cBEYyFkoAIq8b217+z5Kq/CFgpRw0DQ
ZwDbMqYftYhBqbDtBxScvdIyT+6AByBDG2qTqPmxwCll8YTeVgnXv6ARNzkDQVjH
ymU+2unjIbPU1f3czYU3b1+yj954n98762Ddrr+8KPeOsvxgH0F3Dpzfx+8cdGuR
bEQYZLNplszYHMbfMeBkEty0IYGhkDfYH8LC+0CEzAJD9svSt2VaXvRvwmx3amnJ
tkownaxEdw79xSnOdcx+44z27xVAfwCn4qI5Se8AMxqWVIsgNMotTyurRMnjxtt2
rN+S/NXsR6mxdP7KjS9PQr2es/MUlmwW1cBr1calBIgv8Kv/185AtmUqzl83JCca
R6Wq6x3UzKPYt9zz8hCGQ2Klk2f8cgDowjwdQlTFVJpj/WtlzbLwoOUxPPb8DYUd
u1jW13D7T/Yd9Vd/oI0vyq1K0kCf61IEd6sqsseHNcGCYBQPM9Z2xRMXsHDdqJGT
9x1MQkZsJoZwTW65JQSfALK9T7IitqI6fP+giHXED011/Des5iINePMiF8xQzmTi
FRdanPZ77KMXIb/fQmvX49IwiNdXl5njSrgbTRmmMU06cxI4BvK5o1UbZy/2kxOt
iTvTeXOWepLIZPPc3+N0Ghl/8xR39j5WCwPr6zHymZg/2J/MUtLvMS8GivD6LbaB
izLCmeQ1UfcG2uoBrC4bw1JECnU9ny6dgGuB8MmJlZcEFE49xqgM7yk051R1HrGs
S8BEHHyO40ma2D++24dGfalzJrdIqD6PKH1SvILmO5+Q5VXPnF/E4uw/4+U04r8S
kQmybUtRV/PwH/9gpQolxa6bE0X2/mYn7ndoItQ7GAk8tQF/tT0lz3zHNTaoLI+L
vFqWnSgODqXN5OkKQAASPJAH8hdtYDKju+/kxDahpq623RKNwISWrmHjKqC3TiLw
nXuxPpwgDAuIt1mP9gfIF77YHI3sNBKLzRAJfImRHhyWjuRE9QzXuitAtgIwRkrI
2FLw11doJ8Nc8D17Ya13sfM3Oz9oKFLLb3AKfKqD0FKEPTWR26JtMw9KMc3Is4eO
Kr0MSiCRVn2BXBFdlVpK5luWGYZolTkjfH2u5vcMsRbw7sOoDCWuOrxhOrAD1Z2j
ssZylJBSCRkE/imWilUJYTvhg3NNdhpwVliwgVpT0YID3kZKKZtA5l8Sfv96Ku5L
vslVZQSvyCiw7ElGoet1O8o1dQ2xVLXWqWOeUVYfLbzBcKZ7a1zMUYMG3nkVpO1+
Yyr0MkBfqOOau+q/6CsiHn+4naNAxd/ZPMDPKdgL8ypAFhA/xYATztdhTu2wDYd+
fhPxWf3u+EnisVk9gOAM4vkPxYsBffnoUbPBoTlHupOOhL6AwPndpQORngLn4PwR
jfz6cHL8ZUZL81dp0Iw26egQ+/efrrKp3EAXrmGwQXpzHt09WZBpbJmZ2ukIsWIm
KUZqK+5iX2Pf5FmXXbi9GlaBRyrZjM78vTfRJZfRm6JkcWGeH1GLxGxNSKjk/LQb
KHyJxHDbnfVGD6nCVrFG4KYX/S1WPGgbFhM/UySB7Jq/ieu+nkcOiui/U9y0Yb0l
f/wfeDhJ4X3TwgikTkzabYG67QdiI1kUDVmV2WkUX1bRI8LaxtUVMqP/zdvYKSeT
TvKvwCrb8yppZV2qOzWP6uCYc2RteAcyi2hGSflhVb/DmH7M1smGF2qY7/pYf3nK
2p1uRmETfD0q7D0XGixdg3/+twK+F0CbondPN4FAJKYl+QCdCoX9FsqYe06QXJ8/
KU3U7o0TsYOpqhBjss3eKKim1N2OurIjd3E+IMuUyL0koiCcXt2b3vco8BiALGYb
KIQ6Pf9Y50CfbnhccQ0BWhizVQo2Znw13VKga6oy81BhjBYBp8/AxVBeLhf2aLwI
bAZ3FnaZ/F5D056J/MUkDpln95DpiZNVWrtqvIlR3t3NKKoC0UeybBoAxG0uJAri
cujs28E5FFDN6wyYrAnjllBC+gbh+x9ENtNuL+fKWbEHJZl9fuLBFb9lNCGHv9tJ
QaVpr2jAILl4Z+t2OAKTk34WPMjg19Xf/NI+xXt4w8HyNavXgyUzndkK5w2vvtNJ
Zzx4LAPom33tGyAZpx0lqXeYtoJcwNek3zZFc2yZGnRZdJsMQF5Ss68BTzr9sjIx
DxQoCtjbbeMxs1w7Qn9EUjRZMsIVNKaoZgSxzuDhOh8vSIBbqM32XCCsGWS1KjVT
guLkqdMkWVo/QTXCXP4cRTHM7ilZGnUHsOk5nBWdiGiXH8MDBv2pryN0LUEp85aX
AteoOBVcJiPGiKTw5VmcE7TLketzcMjxzfHyDAn2foD2RJie9R+O/ayqAf/Uo69r
EMIv5nygx6yiYQaoRAlHPcV5jM/BftVIaACRDjgrrFMWNevBKgL3oCIrbTt/VFgA
o8RuTBTI1OYu3w6qZxLPwvfyBH6MFWJaznjZPHlbtB65aGbuL2lmwj6xQ81WV9jF
U5qlEL/lq9JF9UFrc1EtvV8Z10UR8FSjoibYkCdYAd8ckTUREhtQtnbIcW5RWz+S
8tgyym6/7qN7VYfncka/PEc3EhcuD6/kXo3RVmrrtnBirbh0X/9KSc1MO36qaoOU
6kyq0Tij+srqVZu0HuEvD5ET3Dm91F44D9iENjpUXT/EuZD/QBsxVJoAVp4V/p45
78ZodQnsIoEwiPnjnAXDO/t3lvXJ9/PN7Hm+c5eD2QjwTry+yAzPyioMvnFgb9kq
hWgE1Vf12vJ27449v9OJaFueL8lvIIMskX3sFjwj2Zneac8nW/lhxNKvlTtpNylO
sPCYqSvrNMVYRSA1Oz9VDr9HmPiaOo6CSHAe2BuWBjWyb1CSwKp2w5nvQdd1/z1M
G+Kf/47tEUCrIRJa8hFjOpafm78IP7z5f7sEPNP1Pk1c6TyaYto05Dlg6bMwwfE8
L9y6TGq5gt1JdbeYaSxsnyoyGeHRGgP3oYShQSiW65C++tTeA2ybwDgW/Qwbf47u
SKV/vr4Yl79dNb7ZMAsu5g21EPr4MIvQ7XXFRugnl33EYtsPd717HHMm898hAuyo
fYbq2y1Se+Lt07nEeBLKiJI14dd4o9TdFp1OIkgvaQ705HPlXTsHFaedL4psEpxd
alePzITeuxrAgj9dlv0DfNgZBQlhs0uDwJfKmAcBeTqdkstJRYZY6pd+4EZ5bVYr
FIk6q387EKUNH6dVT4GGVlPZ2OL2r0qsIPh10ct2nWUZebEvipVtWgnynALtd7Ln
p1RpoySvp8h9dHUZsPxK6Yn3E9lTQqe6NnMlIgS0Lau3qfQWBB/LSnO+aFhP9XHT
IwsR1B4wKw09jdvKPmnCVNRw9yjrkAfhpKioskWayGtTh9MEnjMQfMcQ1l4AJwxW
7rBrWdOOgw3cENbCcBMcIP1geViWE5ejUCl8wKln89tYzvTOsO/O2ZUhOFyafYYl
1Kdw39234rbJ8ItOiCvggzcT4CI51578gCQG9kWPd/6jX6T0Ra/0++k/BZx3pgaq
D5mM1fti7UywCD6cGEUvnhy/tvzoheAAZertSQfrV7VG8701EX5sYgDr6rUSYir+
sE4c70+gqFoUj+o5UuCLR86GceFkc4kgCs7nOPUlR6gnUxhlED2IGJwFBCCAY437
JulHIxAmW0VtY8e1LdANDRBl888nEYjb55xFschaONc/y7Vp0nmBG3J3X5hoC71a
CsuW9GpjxXRilA890KE7ztOeCcyHvU1OP6sGZKtH6DjeHvvBz9B8OIajvUvS8mBf
hdE0JWJ31y4oUb66hp9kc8X2UOHNoOcvHNWP7uXpgvubvoeZo13MIR9gl03kVi/H
o0CHso1poRZBUEzS0jzD6ZQltypH+o5o2szikYibxlkTynegZ5ApZDNmDaghMfoD
HH9gaOXQTOUPkPQ431VNSPaCtirHEbfQA4Bkboee2zm0sVwhGhdQpNErFTb2nr9V
tMIie3jntD58YA31XytW4y5d/AoWkngCO6F7tkTNRFAOjmUEOG1fiStO89cJEQbb
TOyGhac6Z+Bli4WCV4pL9Eyej0fgnA+V8HzrGMbvwS3BHAEibWCBOUg2k4qIjssk
AuMZND03IzA/zCkK1jkP8fl66RCSxK0QzKtcyXzwxC7iuGPHMdZYCeJwzbkaJm3t
1/gbl9c1q7k6jxuAVLqBO+bs6fgmsLZxjFDvQcBcrG6oM65t/D3OPMEr2WenGuZj
L2Jm00Xsrh2HO6xkM9Ft21rtmA+R1220LkhQ823ZUnjg81EkKTD11RAL6Icafcvm
ZwEPaQmlcJ1EEmQgl5nGdVAYnggMH0quJ4+uliSRxDQxswdeqke4uyhAFzxZGV1W
FEFPbY1YpGfznXJGACxYiWM2hFLv8hAU/CHfQMcOjUiXZX0W2WdsVuB6j6EZl+3+
UtvDz1ElN1Z6hqFcO0lodsl6S0nVTHbaxcZ+0f++Eab3cmuWDpaXHNXGHpaZMWMj
LTFSTrRit2HcFwPdAb4phf57lskOx7pT2li6ckOmi4YNTNHl/cPDpJGNMUCp/kVT
E9Gkz5Za0XuxLr3dXu5lcSv+wyXpxj7s3I1ewAXm7AAz9LzIO2Ux8BG3IS37gn/b
5u3ZZl7PV0dKMS0fKG9aLwTWsowdBtr9ZqsUf6SdfTgXv8npqNk+I10ZCJc4ns3n
orNlM9qt24wsfCA8F0lKLIP8kwKBBX+uswKL+xkG8Js+os4GwoPFBAj9haeSB61/
TtHxgd97UW7zJZM6pQWgnEu0NqIfQlwwlZi5lBAlu0EvTQ2aL3C8ldscHemaRp/O
FU251OKv1rWxxoTpyHEAKR6U9GiGir0xM2sVBw/PRLQByn9jMIDantrVlMOpKTsa
u3HBVQyWQFzJzDRk+iPCPJzQnyYn1ka6fcz9lvEj/lHZKECirVxNgV8iHI2+DfST
yhPjdXJffIdjRFzO2GFjEFD4JuSAS9cZxrRpBSiLccjpNZ2bItDKtBoQIYMGJmOO
HjsNlFmlSLMj2bzvD+SfcP2TDT/+SW789//0qGK9hCaW8Z8Q1mRxfLVTNb02furO
hoJCONaARvmJJuxzUx4zmbJu0kPNIPT/9Dqb4RmNokJ6yrzLEwFQznFU2QD1Elwi
V86hnwxViuuueKc+xpMmPYlOyqEFFwEIX/67DD3Kl2L3GUQgStl1ANkOEwiyt7Nt
MRhtf4ukEiTwxaObVqyj6ZTgNvr5Pk+QN5vpOYwgVcyanklrsktqlpfrU/og5L3N
+TYFiTSuBO7zQUKFHpQwYrSYom6kN3S/nViAd+ey603hs943Kn4fGxR4y+qe766I
plBt0unfo5HV4ijt6grkaeWgCoUqjOEPeH9DM5Hm0hyGKEKqlUx+4G3DvAds1nHM
Iu93gjX19Xgdr9rwUPeqJbU14FKJw3Cnqf+jNMs9ByMkCWTcmBPgDMbjFya2KaLi
DEZi3TarkWUIVNEjxOAuG3+i/nZWs8lBCExSSOYGy+P7Ubkpisfpm2/sKcGqxCsA
MS7NyTOd2Wr2YcVn6U5RpG0mZWH9EbKZ0+IzbHVOmlRv7W9zvEKLDN8hLL/VfY3w
4jpMF4E25/hyiAGQQhURQmry1ErIWAiZYvoKQeasnSaGUW0Bu4RBBSmOQNG8N6Nx
k1m9AKgYayYtd+ayN18LnYAVlsZOnFGyzuMJ99dEfcMeyDL6cFPfM7RQk4cq5gPs
yGYo6itxh6Wp/Jjver0dczfas04E3oumBnDu9Y6dszQpLW05Nqo7/OhlZtHXEgcK
rBb7rThrEMW/QSeIwfuBvBuoDG9+312NTotjCWP36HksBC4I2RYoAprYPp2bbMqt
hk9lRu2UJqeU8bNCEWfZ3rJbY1hFI5pF1pnW++fSShazM0GY3CU2BYzisxfPmuNa
Dl/Q29NmnQ6LAyYayybBEdZIlPIOJSUS+7zwgHei1lHBFmeQIDePfQ5dA2ILW7mM
f7mEPVrEk7Od8ycRlAGM/SC0qfhqzPrBWsLqsqBcYcRx1WV8Zxoq9YV8bLgaGZrD
jtwWO6mRhqUCNscW8I2rfZn7FWsi32ihA4isfcSM4BfrOml/ndTz72aBJuOalkJf
9HmicJIabEU2814T0hZar/h+82tb/NeTtMBOaAKiKe8n6zttmZ36ZdbEX2TRWWbz
Dp/49KjZCQeMGschtUQOOihwAm2OHzPFL1JPuiXYdwyuQyP456bp1ksDv5lbBN3y
f/4drI9d65jVWRZ83I8zii33fX0mH/74PdvHc2erWSF1TI6MFd1tDicxo8WDOaTl
v+g4l8++Z/grajq5Lv8Hz1j+len0siMFSfVUGtL6IsAWwGxavtR6KMBtvJhUeMQV
UQkp09vOs/C6B+RYyN4cbRuctvgX03wevwcWQhT1/7WvIMhjg4mTwkEv/unMep7+
L1FzLqBy4Wxn+P0PhOOM6Vs8gzqcaSq4qwmJkKqolAg3/yZ490jOwjt2EBuSzAOd
AFCb2RMURpfPBI6UhVxMh7z+CB2Td2tVLtlbVCHBlPx86tuEGO7W8Z4br5ZOCnX1
9gAFJcbPaem1CPbUMxxB+fuHMVXMCGOyDXcQF1Ea+z2QedZ1eARL3U9ovDO8Z9Ce
7lMXJWwfaKJJ7gynf3migWOYQ2rIrg6dg7axyAV1kQkByIcNMI3CihtbVsGyrM8O
nGVlgbLeniM3hLgP7E+DAcbTrlvok6rxC/M62IzL/UxEQs+eo0j2AOxzwsCsyur+
vED4iSwoyWLLSoMX3a0Pvg+Gp6FB4Bw3qoYn/60niuPkr2mbalCrWKIBpzyNqctQ
AD1ZE9w8x4lojBX/ju8x/OlVSADe9rLAHcAkrWcsfJrevZjSiihL3VptDbOrNAIf
5SGrgf0FQufD7IGrcmkI0jg34TA6j49niuSjGwo1yQfa+NHmyDOrjhQ36NKMan3t
uxQ04eSgQSTlG6Qh7c1+oaOOzGawNbLEDsIp5baR6z1E8jV4aHRBj/nFsJifdm4U
QG3KAaTwRMPgVMy+U3FI6Nk57QVAsOwpKVhQdj/REEOx+PIaHUjGrFXbWH7VDMaN
htU/Enzsn0qVNyAY6/NT8ewBrmiphmcjUhnXx22U00DKdCCp4VjHHTgueChnrWKo
2Fei+J4XSlO2+Cel6jAdeSwiTMeiF1xLpzain/NB7ceYFbaM39f3sPoTlbkA18E/
/FTblkjVXZg4FxQD3YrEhcORB8kbN6KhguhKMXgVjwNQ/FqiUpgNAXz1ivhsgHW8
/RGXzC5NjPFRa8PMSIjhPjX5EKg1/OIc8qxh3PZaNQBHfAWZ99cIQei7INxlQGLc
TyLBbbgCIPuipV5PsAdCNe6LkwKc65Zq9LX8UXasakB+1KU2m3OEOZSpoGIf+gqU
KT1qvTwD2Bac7AodwQbi+6U1+/RKkCgkb39Q6EuRHz9xDk6Rq8/8JdD1TyuC5ayo
NET22eX5SaBRdNMabjyq7gke3rAD5/StRh7QJeDKKR13lLywgemJLahAY6ji96bb
5eVQsXSQB2XUQzPMR7e4ClkIb7iDf1Cgfj3/+aXo6/KZ+C58nZ+yZ3Na3SjYHubu
amdFskiX1TBJo0jX4+zUld0U4Rs9W9DBf6uPuE3z3ngdeRP9wVlMxnRMl6lGng7K
QoPxpBRmWmmkQHxmkospBAMvP06eAxXa7pd7msPjllztjAid2QayrQlu1Q2N5aBJ
vhr4EkruS9Tm9wpm6+vz2Y+aQfaOxlVqyp0UUdfpCGNNJFfKMm2FZsll0kZOpVeK
EwMs7X/cFLCl6Owk01rhxpQ7OzX4mb55jG5J5S7Tx8La3YHQrWVKccBbExDCBm4v
+M1FHrTmq+GVHzake96Zt2DGZJtyBAPfUOCpIzTN3xDW7FFnsGBUbwmwk/JKSmV9
tbtNf1Wbzho9e698rBVlNN3doUognCcU8/BxVxaSmsEQvdbHH5W9cMfjj/Ob5vDo
uS1bRmkvkldj6ICIzZH5IsJUnV8xfVfHILoeGxInrbp+/KZhwhHAJbZSg2bJ7MvB
dwC/T7jpRkgek+LfeKd0zJzXlh9aQxphDObZwtwq0lyeJsRM/CfYz83fvYKWK9eR
gQqSimuODGeGQqMo32S3AuOEeGvOpxqThaLF0nbwqYwXidxfXw/8w3T3YRV7IOuk
NBf8UlvpltQB+sY1Bash/4bvmrw710FkDJ7PVxaPhNHOlGDzj54+Vqbff0SpL3U1
ojngFWEU3eteeGPfRSqECAe96J91eUt4UN5oHLP96QOamVdiXBzVwCym5r9HgonG
HXlHJ0gQG+w9z6Wm5YSwF51LaDb6rIgzt9TFATH9rB/YcuBxHX44oDH7X2uJiw/8
xuTGVOpkVaIV4iyYl68MIfbTbjk5xHOkAte9RxnE0QQsUSVIAHUJiQC4aiUYse1I
CFNaMky5lg3hwzCDBuZgTv7RY7TNZOBG0PwG5jzuA/kltei9wyJ/1XIM+NJHkyjm
60dENxlVwKpV6aSUnFRStrUrQcuR6b168Boc37XHqTkM4OF2pwgcLmvpVJxS73Eu
WUcgPVwnbDdhyvb0I69yExqrpQ8LHkE4FnfuOTeYVoEL5Bd54uhdo9b6VxMjlp8r
Ac09CS0i9HxYCh0Na77HGVrmPvAi04WWyKMaoDvHhlyORXe6HDQ7E/CWRSwDK3kD
vpsnUSKWZEGuMhvzxBEDyZPXJP9Pjzfn3eEEv+W8t6TRd4wVd5lEvsstv37gV/VK
gLL5Gruqkuu+ZYydKJNrvBg0AYfMeknoxq7lurHKPLD0n60UbJ5Tv6s0d4G/s/6O
962PE75Z8mgdsw4YUXcFsJPljoNBR09aThv6VzGNPCoiBl5fcy6xLR0q2PfoLw0O
yQtqYtVc/JKcIFcxmZTArlOxsSADEJ9FFjywq3dlytPSIhZLZF9v8iBGAB+OYImr
Fy+ge6ATL9aj4hRLclWthGk/Cy4RpCAG1SmbeKq5puicfbgr6OraBikDPdGi6HJm
xYRRrdoxCwjkpL2uPC6Iisp74spkCfyFVEgr5RJoN5FeFUzo1clXdsPCHmJUbV9O
qdcHKZ+sV7APZS4JjbO8oh53RQHTq2+w3cv90NJI2uL+H3YzDvEiPu8vGfdcKdIF
EtI1UGevZ6a7OpOsdA3QMRTzqqP5Er3vku/MYIZHrbMEGDAtyMcx/B/oSSGEiM6k
c3iENswEgRm9wayKbRUhizrcxDMTm1boJINkataLz+oqbuS3ectCCVDpYgtPXUyP
8G9MWXYfd7f9lnC2Z2zfi9Y5orqwmpHzh+ddsC7+tEI1y7HFPsEu+zmsAU/DQBCY
gE7jdn7o27q/K/ta73bnP5JHq62/nvonSaNHKf8mVMGOKtqYtpn+nbfVtTT9deLm
x4mw6RvScwyEaG8gOuKuual+He/KStbt47xmbxZVo273Ke0kHH4lERNGNLcyHi47
Q2JT0qVEzYCm4nqUZfie4d43FXMB2o5NRUC16R70NhoENDLmpAGJRR48NSieaNPh
40sTgspq9hlMiKUiV29IvZlJAWDn4nu6DJDI7Kg787FzfWq2E+vRU9w80Y04vW8B
WSgOWWyzrtaAd1fpO10WnW6wkvoHqoVLMHdK/ahRjUO+zF6+vk3/MPA0l8G508jN
su7JHmWiJnpuVQC//VtRwqPygkvSm/3oqSA/8nUHYxZoADk1TChxDQXcNFTBQ/c0
SAc9rHchHqXu1vHDYXUNUdDx0Xv4nNWqbkvcEFTAapXlFPxSwgNU99+S/Xsy1TEu
CE6iDKMcb0GUnnWkP1x/ar3r5ST0uexOCajVWNN6CvWGPT9E3aPs9LyySteH6BZx
vNyfYjaLx8OFxawz2EvXH7iXtVvT4RnpCK9Ly3S1R9W/fFzRa4wu1s4Je/j9S7dQ
L2VQ5k3f7MngBSkdpcQ3G9JjqwenKhAblAJjul6cztTT5rXoojLpKK05QUdxgGTp
yKtDHBjzzrPyDr2BsVIu9JrFkDRydTw4B9BZjokJm1ZPxuPMVJ5iLI/RxRfrqpSl
3WbQd241FHaEqO0B/sWFEMkTXOzl6smXf6rbUCBU8Z4EmEAWjqVNVqCq4mumPSps
w4IJgrIvLLiuq0PQfJ1Nf4M6WLsWVPu7yXBRnr6aukE5K/54KwJIlnpc/ukVpF/u
STaXKa5Z6UTwV1EbAnRb8iwzn/KBpZtP8TshLqnHDLlDz2WRZ84NqBZno3Yuh6xC
jrRsvcv8otfToDnCaEqoyy3x8K3c4T/vEKsZT6oVKZv6in8nPklB3O23J3oqNP/I
Q0wtcPaolb1xUUzTNt1ZHPh46AEcEluk23mz9jTiS+mktxfF7FAZFxTvZVcL7EJb
33z/cn+mzxp9iX621uTplpH33Ydqm1p/TOhtK/YSeA9CKlz02nWP/fTfHQvfca2B
4C/6LFrFx/Pfv1l3X8tLzJdDR3SpXAkzn2iDR/6jDdvKHJqn/eaXr6XRBsRABbW5
DQq/3FHVOAdr6XIad5sK8nqUFfrLjDliPEBOBszwfmsTiOW+nosF3+Hfwa97iuOO
7aG+7I90+hsbhIcrD+yw+Jxyb/17Lp0gZlGnHbRq1+oZvJE9PqlkR775kSPfCGbv
TJ1g0G4ksCbj16cJAY2cWbhgigrwYjKJYKX1qKbLWoANeQil8IhJzOZSluYNmOCS
DMDHayUl1dsNEzuZ6MB3AGc8iDOkRv6gAPqclW2JrrxOXnoVMyfUdcgtXHL7V5B5
atcV5TZQqJnXYEfUcj7SjoKG8mwihyylZojt6g7cAc4xQVWu7+6tMLm0qE8Uwq25
0+zSbSQ9yfFVoehFxmFAtcjXouAveO3rDgTUseY9uTrBpqORuf2dh22XBS7g8GEB
caoDpXud37Nr8q/RkfHEMvfsF7eZ8YvhZCZF4t2o5LQ5uBKDpcKUscyVzSrL805m
12yjNGkQyOMcPD+J7YfyzLStKFZ31vTord/CHD+xxQHdhFmx0J8QFsF9ulp3x8ox
7KM3Qc2X9sBguUDhpx4OHFzdLUC5ceVM1fkCOJQvdX6u4dokN5krzXZEmmKGRfOO
fpUdvi5Zs4dQ48dMziyWlEZL0IDM9kXTj0BXLbx28Ceuqm4jVm7SFIEykaSGdlEn
lYuKEId943ICjzzEuXVZFYa4tHEldgkZBPLRNSf7o9oBNom5mpmcQWpndKplS74o
XI/+iNROb8Ajd+7k/p5eQ9LjGGo8Z6y5DkgJSRlsdUyeAjH2hVaCrBbLXBli0Tgw
+CWwbSnWRKnGWnZLY9BF7CiRgDRpv17nT5LGZ9ZjwSTooonLee6MX7D7rYGzG11K
P5sWKMeZfuingZHWa1b3Vsai/HYg/cvZOL8hPu0VeMoLyB3rbmUj1D6Eicd4gwXu
KggDbuPvS9gN2yowPS5RkB0UEHU/m8Bu259jeffCFFFQhWG7RQYeky+S8BSgMAL/
gY/kmcu7IxqrVL0GV2vOd27senAIM25b9SpMBpZgTDXae9SSy+PZyjr0hZeWUumc
vBA4t4VnCk30kSZUJJtFAOxlyb6Yhmgt07oUD8IutS4oNNkgOlyK5VrkBIrpKM9k
L3BI/H0iXqyucuGiIb+EFBSyPzCE8Bbl+pP3BIGf7ytfhKS+/Z8c1BvBDcNz0VZY
PUAymH0z6EypvGFYPbBPmfHPpL3qRc8VNqTFNVSt1yZM6f2bFMdRR3nTUUR7s+/A
g5vkeLK2Ld9383hqIsKasNgwnAf5Wso/BDF6OiPuqTw4womM14xW/c7NOdqXPz3m
Qaaj+dVLSoCq2Ahvt5o2ZuUSQYW1kWcwNp4OwvfUR/xFuI2lsMg6idiqqAoCjw4P
VEKUgd+E/ASTV0fYxHilq/opaSipMvMvoyfc1i5q7i8lzNj9el5vEkipQmifaDZm
1a4MlKXV0QjsNElGJoWRdxuabNd/KRXuK4g2zL2nUp+Tx7iH3JmoMLG6ucV0yE0z
5OYxjjBP+gYo+GDrtCwmiXlFF1DnfWbAZt5UHUjlkPxuasgCUZWaaJTLGAOABATV
KIA5FVJDCdaodY6Vq7lSe7d139goXdwXPUEpHuTEMxnmxs8coqOSrrzq7jvbzK+s
GbgxXEN/ZXTqXUxUEUEPC4dsbvqSf24OoJ1LZu98sr0FiGfMjhj99Ahr0m4Z5ucz
Cy2SWbYLw92I4OCpixkovECds7GOuN+SDIre9oUtbL+bxWZibVbarvXHtMNCtQ9B
MzQahY5vYKUrcF99ezL4PqldtRX7HpAwdL6ePVF4KJOxQevv2Z5ZH/eZ1l9fh5az
UNA4i1BNtYbkWV5DB3qSfjPe4iR5qcyTwNZLGzsf+mxrev7ptWOth8ARJgRUnqqT
S5ztR0Ou8UFeyb7g3mYwio2UPBcZ0aVSy+nxKswXDJWCYC3tm9I0fykJEShfmUqi
gGnPJakfTeil2eCxHVw6DImCKxSoDZjm/+kgipSWvwKHCz2HHlDdwwjJgRmxW3R3
UQMa02fdI4gXf5w6pbjEdjbfEcsoCkqb94f6uoip083c7XLi2Z8+qeXFCfNGCc5w
7F1iXswxT3DTEJC55QKYBpmUI00F5gkvagXuKDr82fGfBtshqJUMIzOoXh6snst6
1B725VRaFumJzWMiC2pRnqJKNQHHl97pWV4sxmWW3pKOBaGPd0LIAT1ByaEdijHd
DNNn8BCc5eY5c+DPD2BMNNzcnmssph6pGC9V/PvC9sosQltE3gw9mg6mdX2zYPW4
W5muID5EZnYwEjV6bXwBehN+FnIDxNisbXp4hFqy1bXNF0a38onGSHzNcJKoiLfE
h2ggi35K3X0RThqV97s8sRkXGheM03GA8aU08fC4YT9NWE4GKbrf3B5K+QEZyDwZ
dSqvuvl6IQpGdHMw4y/0dulBRzSXs46F9r2IePPtDvMBWswJYAIt1prl+j7PyQeP
Y2rlojOQ31yfaz+fNen0mQO0KdDuI1yMiGQVvSQdVHjrRp/9j/cvRd1tDkjTv2CI
AWxFX3ssXYWJcobEhvTfS6xXS0aAjLs2zu3d8XgemcwHe0bl6dg8CdPIL9ZPrt8Q
jq4fa/DWHKMWDuFgxIau/bcrJCVhnsYmsouTeRDwgsyDI67owxPqkbvQLP7zCgZ1
y+t12E7ZaLjr5ZUw7zUloYPZmgQRyMypvccS07jkTSCqmzBoaq2tDPEoMhs48inL
nOo37eCpCJ4vhdkc4fX1J2WlAILGUWV8MhkwM3+MntLOEGFJs9arcYkoORyB0Xhm
vVnvHvz5NAHEBRak2MB5mBcnWP0A752qNJ9q4jZ8ErTqFgWyxIvq4KoczVKEfji3
txNUnYCAVe2DRJ86ZzUz4UmB30ygvIIhGn8aWQ5zvwyDwu5FpEsZxOzyYNBulax0
uRoeqnsAb4QFdnmTwvsAHD1VnTG0RL3d2GKMdiv8SgFRWisV3t4tt6clVj1KoHc2
P98SKVBzuQYAWZ+611DKbriwcwc9q37ngZ3zPc/WfGGfcRMsPCaQRHT7IqpLAb+Z
YK7+azsp/R/OL5Iqo5cVAf5ZP1PqR2TSO8sCk2JEvRkGrllB+iA0uoDYGKNSaM5P
PWtWM+oOFauQBtUQrZwrkLtNQet7ZwXabkKUQdc8E1oURWqPMHpJgz/72TVsS1kw
ToGr19U4/2MXvuLc3wHJWACryuooKOmFIRZeSPx75VcakQUktbGEPAoBOWXeFH8A
ZFTvGUYkG9pxnXO1IL4wGtaUZS0t1DHCznXwMXTFakpZZ0BnjjdMn/emcaxVAuJg
bPWquWdaywVcBeZNMYly9PhGiOfeFdXe0So6Q4NrjG7iQoQTMNzOZsIagbwktKAD
QDFsDY1zJjBx5yFGs/XzQ9AY/obSmhcMe3yxVTqt6sPdtxAZ6eqisqf2lYEd2V2a
gusLy0E5Gw4+6l6eF7AoxG2VeentUtsCce5uWLZl2ejftzjnzkQwiTGg84+vQbiA
RhuFwgwFTdnb9hvs6M9653oWjsE5YtLJ2yvsLTEIVPqVniFy6TNI0Y0rEwr0Yyox
YYTgo4ytVsrVlfwH3OxcXi1zBfdGzxEPamrjRHMrs5RD/E66vmxGOUT/V2niSYwr
KtTn3M3arZQCLcZTaCI6x5GyUTNg3u8+Iz2Jo4Kgc6I5i8BmugwKCXOkZDzzzUob
1GO9YDF1pKQbpw0DSh8cjYQ4XSS2jiJKbUOZiFIr74O474Xn/VEgZ33zkWeceLdO
uyWgKl8ybsNdhBrAwKa67DQtWgDFzp6ZhgWQPVv7xlJU+QuOEDknJ6fGfqg1fNve
91jKG6cmTQWrtQ2wfJ3rGvnANK7Z2ZWtlV4FEm4S55qhovhusAc9AowtzCWWfC/5
NcJucCNN+bfLRUT4tdXQlSplIImkzu7em9f7hUvf+f9XwZJN+72MoPKCmlRa32eU
G0VaiLKuS9GXp4wwt01ghWcNRj4fCjII5HVxbkQ25bPACQsWDWfisHOHusFu/Fj0
DyxmaxoPpI8N5fyUtMk5a4TMjqi3imJa4miRXLy/N6Y1bE9V7mdm7CYCSPfdFC35
tcYdWZ/oUvSDiPFBOtmsb3Pyx576yp5dVa9b4q+Q/nI8C1JaslI8P9j1ikOBy7WP
lqD73Y4D1NlH6o6OJ21jYA6IMlhkPV8QwZ6AtKk8cBhl5S3V+sKfbIVUD69QejvJ
c5cFieLo3wl7/YO/RHsoiENa/U9V1DeVWq/DwPvGMLglwOmI5QwAXhXzom7VRDWT
QbpxtpmVVm9bCrp0NYvUBwYHhJCPC5Fu1E4BUkFgNhfprR55kUDJAmj15Unmr5/e
TT2VFsaZAwChUtLigRw5k0kOXq609J4ap3bYINN9XDcFqudku00ZGKty//K3/SK1
4sdlOZ8HJ/x2ch6wmcl9sii2FRqMb0nQSNCm0xUuLHgOBQ4GcSgG3srdEO35a2RA
6R9y7LaDCRoXGKhiCmAvz0zKHS5PDLX28tISDb2O7fTf1uqgoF9JkGvi9bpg0CGH
QBgC/OkBQtXpetmq/5Q4fLJDdtvksYEI2aw+CCisoweo37EJoIb7Y6VAWlEhceqE
xSbJrN+JtjwTyb/1XZGLm4P4GTiMVGhU2A/Tix9N31bZaLD71/7djgk+lsHd54mj
zj47Y/takXe0QwlaEiDQCrWZxdc8i3sPJF3R5Y9+gNH+JLiebm3t2U7VgX9vqFgz
F91DcSo42LW8YVW+zAI8BYr0I+sjnqRqg5f9WGKqkesgFEsXU0vc5a2oRe21ztIf
l2Df/KhfvydVZg6j7kmUMfilNux9yandOiDs1RMMGUko2kUdWthwZ18TntEiJYDh
mNRa2SjyaxRrhZJu2GVLA1bLBVbFgKX7sc8sah2cb64YkdbzR2b5PT/Cww/xDWuM
dzbFaGRqIVr8hUOMJNHc7nWuiXxuYV85L7Cdkiu39ceAKulhyuDb1Pcpmbb4nH1o
lJabVVtdn+S1RxC536eTTAikV1zONkm2TglIUdbRTaEKh8e++l1jkT+n0wLo3eIw
6VEyrlD6Fzb0Kfzem66rpaQPQEW3ZJov4+IfiVrgMz5r5SiwYSAi3KjVtE5F1VAA
aEc0oVOylGlYsrI6B4V5QbaBcD9Rh4l6J3cgrV8F2hEJ7z8EsmhGmcIO5sZj/q4V
Z7uzWo0/aWfWnx40pPeEGt6zPVkJTNzTpgqom+zwaUEjPKdpzyE735tlnLnins3Z
3VHqW214HbjSZNZr2mpfxV6XkNiJ8mcn2NzlmByikNJs8fuWVqxLawuNLZ3DKYRc
Yvl/Hbd3Jzzvx94TzN0D3aS14nj08EkSyatHo0IC6Ol8V8Fx65eH/c37qUEqZeGO
kNV+FtxCHagxW8ngHESuNdJIDWm0rZIczlFMPGbMgp/nwgCt5CrDEdeledX8pt6t
cwBAhnRzhFN+nxa7Nvj5LGa7h28E7E1fLYHY1XDZ54qU+944I0jv0Fiqlx4y4an4
8j8T+x+tKCuC+5p07tieLVz+k/MKy6Mr7/haQ5mMar1eoNAQTFby9YGyfik7t7XP
qt3cwvlSHG8H4fWZScVLwi6RGxBd8FhCkme3KF76nzK5f4XU/XtGWknpc1FnXbNR
2jKXOeBudB4E+3rsrJf6d5RHOm9NVakTlmdml0okMMV+ao3SIuhinD4IjgGPU0YY
23iUmjkijhV5zwWHW69qB0090GLalNq44fk9WgdeFkt3q0fWqH9mvtZzeTpbjA0R
ZL7ngWHoq53rdY7nzYJP1CTMAOepsfXy7Deks2UnadJCg/CmXLkNWpLHafZgTiil
1Qgv3HeVKwQUj82wZndjTUYxKoLxJuiM3Q+pdssw69NRuWPe5wA+1ACE0T4uUE5c
A7STz8jgeOIe1Q1cquoNoIbdEyQWjVOMpBcfD75+xOyq8DhB0WNAZ5lDN530qe7n
255VsxoW8usWnZhovFjnVkmH7Xly3M/lrHM73zxfZEonRj+0nGDjCNlwdetw01kg
+RkAeKSEQmQKzEmeOUOuf1DlPLyyVmePWn2geuPNUTj48VMaD+y4puz7q8vioUm6
b8zdQk99jCBg506nu9STQKr2WpRj8hBHSucZXi4R/nP2THIlbUluXE/aFYEvHOcE
rTtJJCGZM05brZzQvItvbnPHqSBtC3zAeL+Htg793487Tgxc4WhDjzAlm/QoQ/Wq
fqHkcZlFChKtlbTqoTWZvesARPqTnVZWLpBizogAbpSR6wdQWuhUDQt1unUvmiW7
Otjc7t5lGn5vyXGIimj59aF1CTxhn0Hh3XUsvkEk0MZJKaalmmpC4cgO/Ge8hHTK
7R4k2xcqTU9cpYD6plABQcyHybELRrd65lYYEkWxI2AOLRkCXjvvslmPWvLpSfq8
P38t2sq3uDE8k6RQbRxXbqtKhST/dp5F0T4X/A4IWEAKhgh1Xb0LyhJWikuKQiSI
Fy+H3PUJd1OVnTwjSXD17hnbASH5r2IUq8TA0BG7YYTljeNe6xpo84dHfXwevEv4
BZ9Fi+6UAtoZEYglD90W1U3+sFhdQBRaBMgvkZrZnYFvnDpRDiUlYZ2y3VinMAxO
Zb6EbRVtqFJnOiEckJTeE0VrsgsD5Uvv7e8TTnopuDPaQhjCHjKkfV7hODgJFP9z
us2B81/b8dsB7QjtBxqN1i1YxwPZDcgIe/3o9IAMDXD091s7UZ5StlrxKQ2Qcsfd
MM0gBqtybiFDwPTIhieGZKB2XRMAAFdoPnUL2mnj8OP5mnDeo6qDfsxNdQuslVSp
cXuuvO9ILBLMXkoJGiiv7qGOI9ehUgbauVwHsos4ctuVl2aA4rH1EKZiHWyxrV92
/1OPbnwoyzF+wZThFVUQEl/COOOXZbc3QSsHyMWKn8i/UWCGARY6SCg9ke1E+VT2
gUhRRlZI4xUlpgAQooiVWDyKt52MJLQeGxj1QFtfyQ4sJ8Rt/a7L0DZ70EK3fJei
9g7QottvrSFXTwqThabCZ3xn7vyzi/LRuU7UhmuAj+TGmYz29C55aSaXDQMiqztC
SBjBuI3skrKE3Q37lJ6h275P+2bKE1HX2jwNakPfcXaCwTiENxpdikkf1evvO/Wv
1SA2+edS/QdIIHr+a2wok6ZbE4nai36SDtAlf7/Gp/2588/iJ/yYRln+0hG7wERT
ugEhyu5m2IgGurJGDyQ8ajU0gXr7WzgFn5G+dZUTsPqqQDLiB+Ir7v7ggr1D1TR4
42ObiRE2FdbLpNPPdUYd2BjGbG1zJrs+QJzuWDLhOfByNRxyeGkh9V9RyhL3Kgtt
XNZ765V5H6Wh+iResfjTLsdWrtDdFkpJ4pc4mSJqpcQiGNGRtD9bpX1oYYt1V0HW
ozrQs1aA1H6ta5gyUCFVCrYCWjNvH9PxSHjY1ecChRp1KA16dasizxjMrhtwSkJc
ZvBvLij07Lkf+QNt3wZ+MOKSGjkJIDeXVwi2CVInyDNxCT27Q5rfMiOZUok1tAyS
CTwehUUX3DwUD4a7sB3sfm3iVtnaJrpLXZhphdpg8RoOCTX2M9E4LbibnmHirUsg
Gq66oUJvy6ozZQPgTlaz21B/mHXQcZZvsnpIThg0CncjV/HA+OGRuJra7LE3KMyZ
Ht1TomV+Mntc5KP3S+JrK7zPXr5aBMnbDagbw1JdQ6oCFZP1fhmcuWw8di9WAfDo
GMgkQ42iiy/n9qlQsOaf9qOw09OwYipWiOEgX4SYB314tWKGWL61Z5miTJ/bc5db
V4oDON0SPAm/1ycGdobjNrP5R9M9T1FB68adbRK38WbHLBA/i1groCUlHOX6t+QT
oONrPh6QlqrgbWfwk4N+6lbiA4xTJXFcRSkFz983wKi937jkGClhNkr90mySjgBV
MNFDMJ4RyxqUWbEfTulF0dtMjojoiUqAxQkyTEW3NhCYSVKaZkJO0o1M1sFIW7cJ
s9J/zovKN3TjgbMQcll9cQyjd9bI7bs/CeUGprnTmDO5VJcDcn6947dH3U1flxvF
5gekYE1SURp8eY70rwOfzhL7JpzudSrh0XHXoZVW5Bb5VEYs61T/WvkTAXYU0Tu4
/VUnaoxmESItfCZjkW64wNl8aoLDRoiNfqsAy8gXg9qqJca2K8w2gtvGKAKmasX3
WV7dM0Ehrj5vJRFnwGFyBmlurv7GWufLhZr7sgNtU+4xjK6lFl4Ixu1447osQfvJ
jg9YCr7cuOrvZkoNmlD2tGSx7V4XN+HSmaoOFG/+2QelD0Cs3bsSsJ/5elwbFnGP
2snxM3HlEqNuqV2HNsyE6HMr6x28ncLniWf54R4zQfBE+xCk3Zly4LULu0LJQlzn
vNj5Vo+tkPQ9F63Nt+EigWaev2Ycl3kvm05aIpABJPuuhLyL+s2LilJfti+VzOvf
cEIQTUiH4ORouZWMMgmKTq0pTA9PqAIvkGk7XdDAm1ptwXa/1lP7yjCGpaWfDzLR
5yGT24G5niZowpa/2Dq7928x8URXL4IRSLgsCcNKm0f3mH8G+qA9tuKp9RavRaF/
aV2mdFVZ8tQ9UPgXTTmOmHB4/1rCTemjX6vpw5XzVKteUViy0EJKxGQBKKIQeB+k
jZ1B8Ps573zD25XDB+HVbFV9K8ae6YfGuAYC+bg+c2sUdZPPoHYeWNt7ZFW60+4i
JqpKL0ZFZOF5zf8GcsFE3IwXatKROVuyoJigJiJk+4LBVc9/lYgT23943QA/wj6d
cQIfb2kc/FGGxUeDuu5N9L+S8EEYpQELNA/rjJySC4HtaWTssXo0IvCuqcsBCo1H
UNrDzWCIfb55tK+klQHW7a/HPFeBxI8ZjdMCm5YrPcPB3AplZWvrFGly9ssjGFJe
mX71/59fQtaPWjCwYITqkq/ecBjh9Q9YFwjw9rpBN0980VlNgZnaN+vUx5L9CE8w
kMP4FVEjA7+RXN+xGqeEC9PDiGGqZh7KPpfjMgc8mfmS5vGpaOe67a0CLqyev/nG
C+hVfUcL52QuHYWAFSiSLkgHspVdCB+e3AeSyi4M4Syhovv0ns50om0UZxsX7Hxp
UGVt5bPUvAkA3boaMtTpikum0onmoE0cIR8u21Tros3H5C2t3xA/N/AgO6HZ2cFX
czg4sfTDKdFNOv1N8aI25UdEwNZPv2/x4vavK9spdy2+eQGuvrX7g5YoqNrlVJNG
2eswSuMheyaftCjyVo/8W5BnwZauZBzuO6gvWr6D+RlMwoq13jefXxdE8bImdHZ6
4x4JfdO1m8LZ4SgDmu5WfhDaAVvtlx3RIEJwdT08zLlrU4alK/MGu1PIpVg50rJm
yvBUUuJ5DIIZtKVJnStuKI8BvqNc21ERwDfVwDLGiRHB8IL5vyDtfyjyzbyHMjO0
OIUeJETo2OLTMJOn/qPZUWrVX/wpC30j+//JBeiMkKBdlIWyBKZxUe6+HdxPfiqt
bdSoAIxx+bVtYry85WSmxvbnHONsxNj9rMHaXVNYXxnhGDTtlrNWr8j3zLMsH9Ym
lXJzgzQA0SQGPRrhQ1qZFzLpAo8Rw06msfuBbhjKuSr9DVDD+ZDX5vWPnt8y5e18
gfR1bbMXCW9q5QPcPgF2s4jtBM/5ggwG7+BoytqBY5QAx9Jd0Ry5/pnQrai5M2UM
saFBRCCPWkfychzKB/1oM/KjE1HtcueLmPTvKAKACg0PvCEnUnhHphm4OUavpNPP
5g9hGHMG3hHJHtuE8JNoILJzTKe3XLotxZYXod7bMQYM65mwxagJCdyoYnXlHQKq
Jy/GvPgWbzVo+3jkDZu8iqv6wewQAuv1AtK8X1tX9Jyz1ZjfdEeKSZjhm0wB6N/H
Zmjfd/dmHYZf2BxeqhXaiGUUhdY5oEBNr27vtADp8iwou++JFpIBmtZyCMv3tV2j
aFf6xCZpHODTN+5II6sp6mbFRsIQyGhfHEBQg+vBQ8WjAb1Cap4zSpkPzSoSuwCW
6C0WBdmohR6pa8lpj7ORYj900hRMl0AzA83HgP+44wY8fKl/OzsAD/jJIBl3gr5p
EEKMlL0dzTUM4JwcBtIOcTVip30pDIq4lxi2ZBVQ3/sHK4YYY3m/h3f5EPuJScpD
sl9dVJnNGfnkgau2f6505pNHtlzXRO7367jDA9WppwaNBjRt4Vvaaf9/F3N6k15s
LBD2U+rYWq4s6mm4iFPJB5Y4IXFhAGGrjVXJfoXRTIg7DqoubYFX8u5/C1vpnVR2
T/JLFZ4VaGS3T8Fu6L0F3n0wo6SfBGEqLI9gtgLJow5eTX9z67X1fms18Ttof+iq
qDhQpXxDJFenim8ChWCc2dpJP6H4NojoOaAm/KR/Zk5ftNpjNFk9c8Qz0lMlQ42R
xAxXSYgfkNJNxxkXEK3lN5r5g04HSQm9D0f/CxiCeg8huFQ7NnQ59hzsopcjPzEw
hXQMs6pspDTQVQf7IzKWfygHpOmJZat+PnuKyj8uDNtiwsONFIGQEblR5oEtOdIt
AYPafnZsPmcySjDOriUciS4b4QR13w8arYKOYw+k0TbDMzUQYxCRdJzQHU1upHTm
K3+tdaRtPgwZKEuf0o473wWrJXqana8lwGSrlhBBPeV3dZdoR+Ify/u6IchwEQB7
qM+w50sXD7+K91oWKY7NGPYXUHcLU6QVCGFkTZdmzlZ0g66L70568uq1cgTHK8oP
/KlKXY/0IsrIT84zyZlL0ysPJ9LYN+zNCwAk8MoD640MRdkLXzdbys1MUYdyW5iP
VUOeGhsLMv+h9RUW1r8w1PwhKOolRM5zE0Z0+JWkQFc6X9dse/7D/F/sPOkDWsu3
utigXltUIf9rPLOABFNCYnftV3vaPQtewx2W4toyaunc1TIyxpXiiHzepEakIflM
x7tNMe2BlY2bA63vhp+NNHx0k1JZ7CystdDuM3hxtIgToNJohbF/xWz26wgleSx2
+bB6slNHggNk8hw8wlPN+to4CgtjXgFliQdLeghsPAZQm6QGr2UbL9XF3PmtUH6U
tm0ZehT5G74Aw5vqDypnGDf3mOoMo+qg2JtKNI9ogtXRfCMsvB71kP2U19V6QjNp
waUHc/SZxPvpwXFYYbkNmpMsuDbzOy1zqxr56uDHUIJwhpax++L2gHx64F2CfTtu
WBX7t/lNcZKKL+SB4FehvZnhYHjCnuwxRcPClcM1JK8X4jlWJ8f7r5zMgzHH9/pH
TXgwFAXl4j65lyju4q1GEC7azq8I194l1fATQt3d4oNWEtB15I78qZ5PdD8OKj2F
FjJudtDrwirLvPpwTTmQ2VrAtCIK5C/Wnq10myAo6BEx6rJII5PqEHulG5IVXlFT
YfK6CP8HEq1jNRI9gnJqp+jgnFRXFx2OHptKlFtaEB8H3TZ7Fc68mKbTWtDnYsm1
ji0bM15G9p/wbUg0tK6nusWJFrE+2ooJwQ0MZtIZQK+Zbyk+oMYpLAFa7C46d7/n
Zt/vP191dHw+bQYnO/gF3L0aggOXZ8t13Gwj135fJu7kmyH8A+fPF+AwzfxE+AcY
mDK/Kqf312sT3K8Z78pQDMMHHTovCbEOnA1WnSY6xQ5TDeyoRxvo9tHMZoRbNFsR
Ng5kwpTyCCbrdRJOskh4OKgTqNLLWPAAyNrnBm1Qv1f5KeLidVkodjRGHZLl/SSn
ib9AQ3CVUKZ3wKDKRbKpRlW9dO3E/zDgGTFMzTfM2O7MenQ6hERoQICqMugvQQAc
Yo2Gimdyqit9NHUuMt9Mnexy6GH+5EbtOjaZY+W7D2b9s4c0e5C2Ur36AYgcw1Wv
aubwLq6eanHkvzH4N69+gLK9wJs3vFQR2J9NeZ7iJ2p0HAhsoMu98HsO24XnSmtM
BT3pL8M9Wx5DaWigpQHUlFsjo+0RH87tcGw8c/EEdxwQVR/2We2XChRfdeOdWwZ2
YUHQt9oAK+P7Jkv2g+kl42JVwkEtkfAg4xS87dfwZmYDAORT7dNVP9OtuGqWtQ4Z
4Jzz8Cjz4250uPLU4P8TlyMqFR/KF5mM2w44NR2kupFBn58DnOiVvnV0h90yw361
N/7NImDmAGo4KdV+vhWK/u+de5Cf3RQ/AimndCfE7S4n+lYihDsDWj2/hn/gy1+j
Uhpa6AliFpfDkZtRX9eZCG8nNx8aH8rXHOkvb3L+7ix4AjDJNBPExelk7EVDv1wb
OPec/mJpr0XYMnYdgtIlSBvf3M8a2c0QC3JjQEgFfbLSW2ZGMUpXMFgx0ZdFmniG
T7A3DbOn8kLb/+nf8xznL4JBFywq1gwgA2kPphekTXISmCIYXznA3mJQ2avf3DRQ
sGpdNME/Al/wxa7JjesGgQDgzPmTTEPF9jyzK8E/NtKVrn6idnsGCMzE1tUFM6ps
pO8HXwCm8dZqq+/SIc0LvXg6GEENZVQzmkgmLEMFIc8UojAH1DMYdmY8Ncl2VTrs
/EKmxC5M8CEHTF86OTBggKniDUBTy9Ky3p6fOWe6cabOEd/SOHNEbJ0ojh7zHSRu
JWcNqeQi/G75U42Nl/YNUOdms9N6FeR3F8wCqkrY/SRalXfYO6VeKvVdoRHtUa1M
tXj0c+RfHCi1keHc6bBwWrToJt03gUm9tRpb5vHlVdLNk5PyQFnZppDEVYsnaibF
sCoUVaM03AYCsewnpbaipsNB1Tz/xVgjsCJrnIP1P0d55fHBr25iPU0QsomtHBEF
o3PFVVHlfp+7DO7y/72HvhxeLIWvWq00bqWoBQmIc78RZMD1XOEfdkdQjow/6mhZ
gYYNNwH/qCmF/6BYqMePc0zH0PDkDj0BnYAQOMTefA1VUoIc7vyx3uI4PxN3fgW9
Kyn7oiV2mxWlowtoAvyOvj32oXyQC5Ad6hGQ3jTwydLpIkkPF3zn4YRNLsnieJp1
2vs/8wBwS5n6/wY/581y2fWnn10plJZmESnE+gRbfNODyKItyvVj5OsAK55EsaTv
qJmZJre6xA+oXQiAaYFPyxmRG1HZO1Q5D1Zb7ORcOvUjw0pCAPyrR1f/O8mdYk7K
dJ1j5rabxQ+CO26Pp+FDUv8UPTgwlIEEybr9Y2w+wfmFpQRvmvu6s9o1Ux+9p5XO
hqam2dksZEfUPRH6gck1KaIFBulUPwsX8Q8V73Jt0hrCn3wx9f5ubsFDefInEVss
IuxK2doPCSzHC2ksT6Nu7BABi5kuI+QROn5deLBdTOdR3KM4T4ORn9bAs4DEjFAw
Qq7IYYxhycFJ/hQ3ecVBX8PdkasUtsMMwzPJKTKQtYL4KzH31jj0kqh0o0rmaExf
3Uq8E8J7UOLoWkfvWGjuKu880Gt1czz5EDLA893TsgstYQesMloF0ESkg9VjJEaO
Hn9fSb8gT2lHb5xYDPn8CUROXmJ6G/7ogfA5FhkA7S+f6/ou0zH5OSor4zVJZoTQ
2qDz1eJA+TviBIol1zHKrJ6sImsRw0VZ/bXvrVN/zOJz0hLSiH7VU/wrrIJKUJVQ
P8wVGtzRmys286gAGlc2+ozn0YSThP6Lt0cvLTtLS4xCEOdQxH+qxwoAp6J2wAIb
SsFUn3Ov+XUJ9KKTx9hHri5hEhjGAPmfS1ox6m2U6LMFEr4NRbHTu9cnlxAgJ1Zu
zPUSxnRh6oByHXxNFB+VjvruRrU+JkjHIroZofdKQC8zxjQ1N4J1Y0RHQPb3nDn8
3leIBzZAcnpRRp9dsOETt7KHOFyWuixBsNBhRVcR4nGd59IZg9H6p+uHATgbcIy+
G2DtMGaizoGgWuCjAD6rolqiAn06kjHBpu42tOFIPtBvhb3FGcdSznKkA1bo28Cu
EXz8/IIBA1y8qrXwWHKYmtOX72hMl9XWq9jA2YKFHhOu4QKyAVUa2xWkBirhPqHJ
+zS5L/xYgSfZVse6PFwmnQ7GJbuqk/CTHnEYU+4m45kQPEdXWIBTTC57TjZwKWpA
kzTXaMw7MFnUmU4JlgjoF7SHCy1eTSFVViQ2LODxoivV5n8DK7pev7XhoatwFM1F
2cfhg+XdYO0+uEZ2ZCLTn8CciU92vf9uFx2VxMCS0B6l91Ej5Nn64M8WxeUcTtpI
Z/ZhJINiJTSlzwdR9YV30nRgOgJS2kP9FVGvOTYXTbXoq6/E091XaoTh1r9Ryf27
i2KowXUHLP0SyavOYMH8fxdVSlsp//UF7ZtXtYKSz74dncR2RGFc7B0ivL4P1nk8
1Q+1LNuPDviYGGYu0DK40G3LlDI5rQm/6iILX1z6EbduxG0mRhcHLIYSXct73Xv9
kurgaZqFkH9QngWGMg9gRPGmSo4WeF9pGWxSeNgin9qhhwG+hPc0V+48ZcFHsJPb
NauvhvX0UuIE7c697jVBON3t8tvQhuZFAVvxbYiwhMrtf7GA9cV1SlopdAxRT/hm
KuLI72L+/KysKGuP5wb7iF2qf2MW1dKRIz8Rg7HyTTmqJUEPjmOzOX7elu3TIGOr
h2EpgP1hzHY1ru9mc/AseL3UMEMsboUsg/g0YhYwlLb1wNoKWbj+u350/27hPZDp
VnGu1x/wR4ZzSQ+ePUWxz5dQUFaO5EJdUT9xyQg33zhv9v/rmYzEGvPm1xLRVP2K
S35+xuwzZzuMLCZQWlbhwiJ8JDsp1xEdoMQDrtHF9QncmlRRavXzLP/AmxVz6/6B
0GzxQ8JMfqeje5KH7jTQmemnnHanYjlyJWC5o1bzlcdU5NqU0LDsNJ1wg4N6kYOQ
QnL5sDPLY0f+A73zSnN8dqO46/5QJbf7nXXVPSJq599beS8RFZIPeuOvfYd+/DKS
RAPG6m42KiZdA9QVikftFqQa6z6Hz91BLidmRUmZekfPPGKkccL+3vE6WTvae5O7
3L2QCrLJbZDbGkucRy/LvH4t1C/0rYnqSlBX6gNQQjApsu2/0t/H4WCqnyjunxWj
pMi8wLIlpelA17XKG5XGzRyZrRS40H+pUy3ruk+egTqoW1ODEz8kYZlid7IyUdo2
Jl5iZV0S1G+7F4Vo7E9Ff6oxnmQaHODbLsvMSaC+vcXMSuFGI+1PiH3jnW/mF2QH
mZ7jQjrZsqW8ljGE6nnmhbG8Z4unSarH+w+lw4bvd+z86pgExfyXwjHsLKBXUP5R
VHWePnlloNr6btcRbazUAPRnO4otuP2o2wnzfeKHaHGjEBWg/69ZlOMNoqme3jxW
hoEZ2qn0VoKT4/hB1zN0q00ITw2CsRnAvucSgHlR7hOa68h+LP+gtK26/S54Qfqy
SbP1cV5sYBO5UBhDlEYQ1UIoa3rjToaJJQSR7ebyh4i2x21gunYaq61k/8n6s1wz
+RA4lS7PfTs2pMe51bVsevEZS+hJ29I2fdA7haKjFudDiQ7QZ0yuHm8JzZX6+Xn3
mQU5I1oZ562BfQVGBIuN4pC/tXuws9yFWCMBqZDwE4mNe1YqoClvAzIVA4fDEnXB
I3eJtvTomls8OGuxwSRnDXJMndUeqZxMSyp4dWlzvy5B0F/Fo+fk163pZdwPPqPy
TgpgDvTukeAVpMtNJmURL96NZwcBJ1m8oK/meMzjxIgnUsJQHB1+VTTADDYT+U3A
GhPNgWc67WvQOOn5DBJKJ8ZCFFa9tPfA0TSnyOlam4zQtno2gr/Us6qF1oLR3Htb
uk1pRy0TBsT1va3MMYhQQxjhAJJkqB/6SqOnr64d8n3TwRQJmJuvMwjq8KRyjrkq
QmFimPX1GDAklzTbJ+wBlilU0cAAkb3PCOqZP5rvBVVoQVEBNkSNQgfBB+h9Xxag
2bEW4RaNCImAE1FJauHflZI/eR9fPUmrmcyqSGkZ3txC1YJKYrSA65OMKnx/0/dx
t7wk9fuxgpbIFEzkj8KEwiUJNNV3tUtPC5LMOr3wKD5PCUqD4k307TAxKW0JnTLv
7Ga18QACAYOf9vtXEkTjyRvOdFxekWOMHqCZ8jenKoGwqCfDQ4a8KAEnWqO31hzf
hX7sbl1lVI8pzm6vnhFSBLc9hqK5l4sPel+eJ5qYsWJJSlc067NRr0K3Pca0X9f7
aXY3sv37MoPKNaAROiyx+6ldZfENdoeeqvwWmfajtna7lC3qJJ2M+Os0zBW+lw7Q
KUHetIscO8dFaLk90okq6YmkrvlMx6uN4YVFP9lcUgdxjphlurzX7/dRGNs0ryIN
3iHBGgGmRDdhDAOw8K6beIGIQk1qz4fNVcpRzBNaTWKo5c2/deII26kfcVEAUp2v
hP7iNmYo88OlWe47TAKncxTrwLXcH/TuZHcgmE/DPRzvBq39k9JHOoX+GiGD1anz
ZYSQ5Vm8sbfKcUuekhljbWfbEyTU75pYLBNxtgQxp9iAKRRS2xsRUDrmgKMC35MG
uaRFvRHTRRO0XNruUIkUfU0dB0D2/U9s3xm1f1+JDMzJPI/DGvUhMqK9a5ZdzamI
tlKrFZ9lxrkwBdei5m/xMr/1OGIuB6j4GOptKLAIrhedDTOPBvrdGoB2CSj+gWyJ
/5r+G1IYBhJ8Vg9Dm2hlbNJ2JczdgpT+IFTv4Px8j3F9F4/ZmaIvW8XXfjaQZGx+
KfQT/jQq/lWeRWVQv+NgQQjk9lNgsaSn32yis2DbzSYfKNNLwo/N4GXu45WLaZQo
CYJscT9MM3jp/k8LDIBcFMENUwMahzjZPv2u/G74yKgEUY8a8qMunwFZdLs5GhZ/
Y9Bd7RmBItJVFuHE7sg3hSWVEyYyf1W40/0jU5s8NAW1NxmuAw4gqwQ8cWbVRjqy
kIgBEBDhQfduGvsv7a5ZrQiG93FzRcaKu+1O19fianBRYhAcmIk94tLW6GSp4PL/
lNYZkSrairAPN371WgzqC6xakUhsNPEazHbB/PcPWAatZhWn7K8j22g+5y3wAM9T
c0+i059UZZ8Q6EnqlRXjPJeTbxbPj3h5uU1Qd9mEddwEBgB50pgqPO+TpRqCx09N
/LhkonuY9yE1c10DU5u/oDw0yhXXeHp6BUXyWHqzmT0ZlHfoIzAuSwHDgNdZ9d/S
L/KkrktjpA+kzhHEn0Oi9leuAR/Hyu2f+O0H+4aRS/RZGTzptmL0Q1N6cbKMuiSO
eqCaSi+bPejaR7IDagjHJH870zzEJVxOWIb/OtADOsfDmwyLSAkGsgCqS5PrQU2O
DYF7yiLDK590F8gQS7sXHVl6zZvgVBCJdEVdTCji18PxvDIiTrNbY41F32F6lBUo
XdZAvpVDx/u7Qq7E2Ki8Eu4u0OmNjniTJEUqWFGlivt/mIoQ3si+NaQmFKjwTyEb
ShGoBjnuR88QazMP23lQwduS6KzUlTrD3wPJ8HJRWdlMmyI0ttLXPbj+PAgVR1Le
XYqdSVYKQAIgA5p8sQ5i0y9kmK95JAz6bxILugycegIL3tWZtK8mVo5KBnZbhZHs
SzJJCWeRi97eKYJdPizye8n3smSJP7HZFMJ3dncEoKUDGCtlRGVfaF26q6tELZNd
Ic2gcYzuG+SFvhYpsflqouRaoM64scr5uQW71/eF1d4a4X3Zjnqba45uJYUvacs/
YkThmaBrQL7OWPMqrDEsiw2HZ4nZARDbB86IOQcToOTEslAk1wWrFhHO7shogoSS
7Bxfvx9htW6sAgKvgBB5PpV7QlJumLGyQK8pV0nc6XFUOTylVDLOzqfJoTeQyvsI
dCGRCBHrGKQPS9UkpDvY5eotmP/p+rMgfffzovKeoisiRT3utqKgq7FCEa+Aj8f4
FP1xkDNFGrBqtLut9neih1/qLBHxa4DQ6kQdM1Hv7fTQ0k4zIknJOAMAQu+Ead+h
2BtsnEN8Sz9c8KgTW0pIqhPGLVA660rgD7Y1rTeLii/p9Ow1TZsKhGBX0WxMTa+j
GTVxHS9KZ0AovHiSMVZMxeVC9oJ1Gw0sR8c8oOZkYJgGHmRRWU8j7uU0ROZgZuQb
9ep5Pxbd/sT/eHwcvvEd7ZePTHKfyALgK+7PAkQqQOaw6z2YuAVEZqVblcpRZVmr
TwFc+4BO/ggtA/ORoZmhG3cEpObQCPtYgmnYN09NDIjOCvFzOpvewTLsg/pHEepf
ZtTGgdjgnUXKOmOfd/rL7GWL+bIz+8P/EEybCuLUV2v3HuyzOBo299/n+KB5j+F0
lvWTLUzJgaoQcp2ZpYojz8uMZYun62hBcl7yTFfQsFuhQDPRsqb4dlr/N1ay8fCt
wowIG6tnBhy+JxvAY5fvWFSVxVBk/nWkhKzAY2J5V/VrAE+6O3PRjhJMoZ3tsk00
NI5WvNeekow7KdUCIQcFkLZ8uXEWJzERVWhjvaOD7Ut60ssKXSX6a7M5gwZmY4Zn
MdND9MvrZyfNbOWKSug+7sQCslWrhM4y0FFt6SV+ohy1iwZ/4NjvHioDMkAnkGNp
vCYPBITg+qTIsOw5tMH1f/r4dvdmcKbHxmqJJkHLwLpCZlZGe23mJlJhfk0iMOQP
m+vapFsaB3BWpcVzhVIYullNOR97FMzys+QHwYbOtA5Ycr8NLKMSMCHyMWpSA7nX
U667M/BY4iJq24jubYUaLoAxw1he3H5dUK1ncu1DJ9uqnDxqf2VAD1a8+EDVXWEL
tS6es01XAwcQFHPgTHJ935bJ0yJAuCXLoLe1TsVpU2+Gn5HF/fY1ghuuBfyaXvc4
9LDd02Fekpa0Ex4wmumqBVZ/AEZgBH08sj38STJHkPIcyxJKTxlna9D8o3OhhNFb
I0QVEuGgTqJ2LErzdv9AxZbBpydj19CjMKcRo9pbCuTB3NiF4tgEk9lizTe/zhyZ
Mzqsi1AG5tsZoj0JIVYBl0tOa71mKgaFifMnn/H0CrO0U0Cqvzn6zxkRUSwIo5pU
kc2hL/vLseHSAri8QJONQo/qZzIfu1PxmctfEQGyp25iHAANue3sIlRjusSSXCch
CYUBm49/dgwTsNqpFKuOvQG+WKcRuklAhlOM+Q0TpWE2FYgYaQxvjsh6h1lOt3xv
BRYeXQXLb6eHvMo2mpLZrpBBjoPAnVJRetsvk6NSj+QpPkuI6ximKe8UVVj6y1lC
oVqf6UNYknDallo748J2uhfVJYlbboRuMQATkHmcPTVXNIVzD9axEicCAqedSA6c
veXkpm3SLebX2xrcZlVkZRrEzG8j0yr1pqa5MdPCU3wEQdCTWD6hmQXyWWY2N8Jf
rG9DGuqq0rxD32Zc2ufkMeMPNBF8Rf5peELOrOcaGdvdXQ1wVptJAYJxv8SUIZ92
+tYq0axcKIdaXBCDcoaUQtzmSVrqkXUiOsbCz3sev5UVLqshxLnvQLZk9lhqM2hY
c5je4K354bvKjlKOI68jiQanlhPZbRvVfYrrHYZ+Ctyc59wYMfsVgBn/P7aAuhof
lBuiiroypCeAXCqs9OA8uvUOOjuo5PbP/Pwomi3fFm2fPZJTFIE0DdpRsqD0ZSJh
9W/ANHtjBMOAzu1CK5pMECBjmddnRnjG9rY90RSKB5In88/Uw6MoVheAthAaaGBA
nWKN/BYktqJqcpR/FlOgu0UI1nlPNW9jywYUASC7snzFVDZ0pNfDLzmHXhxUfJks
gPRAHCunJrtgI4YF9UHkrVLUrtMJHHgN+lJQrGQ1+oyHpyakk0I8Eo72sq9eZnAk
NYRwtqtpuTxLLQOpPGSmRISiz/88tLJ8kAGlaJiu31yGuie2MvAAUx7RC1XLQOE0
nkk/0da64WusBix2WS7GhV0BIJQUqd612yezqGBBWEQsVj0qyjxtxtTpQX5yHzwv
H99VMdtacKW0a4+tVV62TOyveT7icKpAhEujZbAxyCEFECz4R3UchdFwc9I/QfYe
tXlc1tJz4fow5zts52XVRgRcqVCHiPfESyzvIEtLKRwPw681xRFSMLpuJwEGlktQ
oaNG2aj/ubdfUcDIFr81t4Ss75xn5rBs812Ebn2yDZjGnuK4r7i7NUwhRSsD9xo2
s6/KZMFrc05RSiEOJMYBpMF7JlYdIiZab8Bkrz7y0iVxYtC9r8ceZ3yKwB5nco+z
2QyAXXpNjEK4nlqs789kIvsYa176zQTdjR5hZXEuhhlp7OW31rVNcfN5YvWOFIh2
faHNCjfpc6qM7cphnG8kifwPAKkAGF3ygJbk39lxkJMnNPGv9lojIG0DdaWZ1+04
7vmo3kdT/tAtHXB9fC/EQYxx2puc5mXV3FUrNVz6Cz+epbyT/CMUdJd/CiJx6ApX
alEjWIXo+mkmGU8btpHD8+e2qad/R4/RQic0vJ8jWWoZVz4wFZjNyMkD237YGtOt
RRwIn3nxA70TwqS/l9Ev4rtAfhAhh9/XdP/EZrZBpEWc1qjJmDmrYisTxafnCybd
mHkOj1+iDVsdWm9AT7jcHc9j50V2OWxn79jNbyhXuoKmjQaKR47MOP0JS8GTATDV
UtFHOiDw33p+wqiVWamozlrn8CW0AQTqLWC5EU7nJS9jvOUHwvRRkF46OFphKKBD
qPD5NJ2j47i5wNobIPMX0vdP9aOGFtBRHhSHQm3OW8Sahdf+kiWQ+6Wgcur2Nkd4
5XqIrCDmx9DIRiRiB3UlDi9QUgIRMOKidZMi1TY5iiPM7mtqtidAKOFMFwQzhHGw
on95Oal6vxitk/KnQcHN68QO6xoxnBpCaOQaBjQqq/cmb/8TgoPEIRyWIoykGOP7
1kF5r5eGtjue1J8bA8j5nZP7Ro0Z9ujsmT1BDeWms9Raf2bEU3soSwPG+39d9xiv
N7K8mOsaTOqsvlQvgMEHI7g2XEF78tTe5bk1W79I8d2IAf73d9B6L5Suh//TMbeS
5FDEFwj9pIjEApdLvKvi+dDkuujagvKD8TWPqAIBXWen9LWjspwzMPaKRx33j/5m
8aarCkMz3YjlTEQ8c5MinQMX4CN+A04fc4LJdT7SDwA6gTgaivOQaxmVG3ECBpLz
yk+2ZhSaAzB95QMQN9lnuek00lFt0LpLcmTQQQ6XJyZ3szbbAq8Cyw2Q/ShMXNw7
9Oqr3/YFpvLf14Bv8EmNr03GOD8x49RINuu1O7v7jyqSZlsNrqfMJRO1FZOP2J65
+owqbbjJAJ52gNbkcINzVsBGgg9H147Xyc380AnI1X/q3pZp4LBRPAXNlrhU0WPK
zj6KJvzeN7uA/4N0YCe1pqYu6PRV1gtVRAPAqAYUL3xUV0EnCq9D4quFUmqYI7vG
KbTVf4O351FKSujtJGrO6+QPnNdRepATe0sL9wRy29wQmWT09p1ODxLU41Ez/SS5
tUQc5SBa911RLZPwPcv/OhS11avhLcmhGLBr8EtEOY05uvdqAxNuujQgjk/+B1WB
MOCY0vFDToMwxvhEIV/MBiHsYzVcWrnvDLJ4vxlm54tIFIm5aFt0vagoMOlUzgWr
YOLo+/gH0SY7bAwJheop8hBAvJdpidyIBt31jgUOA3rGPfnWPEUCR6uTj2b7Rz+R
I+vdoIGFNDNpAGHG93KcINVNNRntzMqcXuGUMP4e69ELz5iZl21XiqW5pVZN+225
WLrah+7jSsI6xwxrk3aXeYIQYHjqCR0wGUvKIJilpe9pJCT+eMehl5kdY3RUinfh
mSivG37TSljutb7G21v7HBGpWt3UG0Hvh5syPxIejXv6jzTK50vrP3GVhVCpRg56
U5NX5OeG4k/BldBoqb/B8ATwpc2/AnvYgPKL70sum9TuLYS4K2hTTh3ijWZTk/Wx
I689EBwFHivUoxJ1hy+PyhRzkW7hokBi7Pk2QtLsKw0x9KVBoxmlkXB+zmf5ly7z
5EKJ71SL+uzqFTGuwtg/XAK1qoP2RGQgr29n9XiHmlJPKaAUDo8bcms3I5SPExqA
ZBUpnUsoJEWKVEvBXuZ0UPp/AH/vKIWJ9iI2E6YRU6qc3tMTfy9ddCFvmOpXns6+
2rQzG1zp+uaFVu3aO0h98XtK8ngomqTkDxQSv9/Q/DclpsYneUOyxXIkOVloER4K
1k/vWsVf56cDHQ2re3rcv6H3YJ+7FWgKzF3pgqtzLLcsGhoNWSEDuGtoBot9Yk/z
vuEZG7dbpw0Las3OHd0AvXUwksQQdnF7zaw88ccvglQnnXExcAsDKaMIUhxltxQp
6ULxeLvoHSKzuumD9u/boQ6OGtmzWYDhQCRf5VkJSDNiZdRH+6gztN4kYrYNhZgB
U460HoZJMUwzcBvhOxzPnL+BmaaHZUxrHt7+inyiR/koe2qBKnwtitNcU0wtlDdc
F/Rfo5c9ynigNFyqg8d5WAe6MCcVrAKkdKsZ136+g3FbkPtoR16RWhoQYwiGEfSm
XEsRGK6sMXnyYw9YqfhG1OKxrHzMsJyAxreVvYYfncZ+dEk2Vad57Tb1PGJRG0Bt
wJxSKfyN+y3n6/5DI1Pf9eWaapQsMyk7/UUtm2jj9Rln9xnEojjZZiiEKtVf4ejn
fpd35T0s2ovAZhcAuM4vJJ6lxLHhQ4ofMqWRGMwz5BQOd8hTBTctio17JiqWy4VO
UWeyflADzUpkGhBXl8xVRAtMjRkJ3F/OOHolRJeXRFrxHVFBlRpLGrxW1sJGHDGA
uwLA9RUckJ+fll0TQOFqEKQZDkrbQgylNj+VMRIt+0/DI6JDSWDplLzFsdPgWHHc
IoGasgLal8KQCSK+zL1XrjLqYJ781y+qgw+DSyjWvuhyDgblGKEjbnXHTUHv8h8+
Q2/W6a8xuuWq75qIaN6w9gLhn4rYpLTCCaMmj7OXn/RFbJb3eMwt8yj0BkXHTd6b
hzvcVAQg3KynGL5Lhwsk+xREiRCSpdgAiA93P3v/cV2kZxju7l7f2NubYneQQDRz
Lm78pC3n3JOMDlwl3T0PiD7B6o6gnl2xqpW4xCZKN/FWfJit22MsfMXIgqPgEk6G
Q1MvCWAs7WN95v2ohB3+maHZ+s92VHZ75zTumKiUhf5KmS4Yx8ouaY0di+H/nVu4
cHxgBNgW0x9tCFqDoW5fziCJuTnpv2bLyC3/sER12U2qgbVwNo3NKMjmRsWbqI+d
Ph5smSeHlqtjATnurcTDckdJ2QgohbMFSnKFHUYmBmO/f+gcaZLSQRH+xFbdN5qk
4xoSzsuJCzqGvcSUIE0/fnMcTgyg/bWZ10nZX3i4Rv7+Y+bzi5nD9jwDYVbRI/hH
bOJ4HlFGvQ5aeA3H1o1Q2D9Sy0SgcpJ6MSqNMHHt8aL+bgYmNgLP/aANmvQj17tM
4UoYlMiQ3nO7/Nf93H8Wauk9JT1j+HThDa/iTlPqo/RDDxp3t7FyDs17Bu4u/QG5
X3/HfeybND4QXxmOwxxXhCaSbU5NLyJ+MkQLpcT90+h+99pb4gS/6WLIqN0Xmm/E
/8ToW2yK1Ew9o5/AxmyKomA95EY+kMqc6PZrgqfjKK9oKFHHZ088Ixt1qlNJR1Lt
N9ZI0Yyn8kHYsVxF83hifFu3geRA/3TMgirsRZaDfFID2SKg2lrWNPf9C9CYg02/
8a36vkcLpVTC5UPaXBS6XDUD7GfmbnKKosKgWev/61F2LcMwYBb4BJVY9Bh0aNQ1
e65EMNMH0UafP1oM8Y+InQtUkBdM6jyvUpMq2joT67jUjwxS0iYxGLAjdLlajbP0
oagky0Z223HogeJAFb3zCSyapxLPDAPOFGj6QLtLYji3hLcC5AVRaUCZIaEok/TX
/t2N5SUeLJLOF6A3Pj+vQSrqOPYiDqdrsa5wOf/t8S9F0Lp7hQLmWGNQoIaTfBRF
hTdJJs4+QmIWTZ0U8qtjg6UrE+EUU+RvXsTcTC0GVwAbTW3LHBvceLkUrI8eh8RS
YrENw0MuQndya/5B3lwOtGVmrt8i8NJkXxuiIK0+/GAAeSkaMsqoNsC/XCvQMrkk
2rUKVEDGCiwdISpbWYU4tdOtfGRk+yBQeTyB/yu6zEObo92buLenrFAN4haUK8ge
wi4lxkkjUOYlzaTddtuFY72MvEftYVhyFmK2Rj3LUuPTdNmBbdryjmJmoqSVoSLA
M99vsPlG4coyr9KMxcAa+j+SCaByuLdEfQ6h2WAGqUlmKcgvB3JX7VjcBRZYn8u4
lg+Cuq0NV8x+gDbxImlaIwdWCN3zhv5UdUOtDX/mzxUIP/kopBG1O84NCzbUdTSn
vci/q7/VcJoLZnWEjw1PECEVB9C59sVHGZ1MFuowMPHNGvHOVdK9J+paQbfQMAxl
C0FATyANt6BmATge2k/Xd9ps/A2/DwumliM6vP4kKfgmG1hQfmxTi8hW56t58ElJ
WBFW0Rf+mViy17vRIB4Yjf6WiAc1HWTaY/VyY2h+GQ00Vt8lM5zosLI+Z3Gbt82T
wkCg35mXq+9Krymf7Cv7A/Hu0ysDma10TPZSDuYQVNhApOTWc7ldIEIXJ1L9MDlv
K4R2OaWeHrS9AP/m+LDKQGnrvajMLGu/lw3z7NLtwEbuVkAw0xz9CTjKU78gnsuZ
Y0tLL1r/vJ7hPK2EnpHuundoYf2BiYi3sMW2eOP5XyzALHWIYzB+8Bn6h3c6LTFy
i/QYfM2Vj7G7zHNAZcsdYEraqP5MhmHfNjT54f4sL0N8cSneNsY+mG9hT4Gw6YW6
NzIMp65PoXQuQ2FjL11xdg2psHrs3taNXI8ZUWVxaBmpxFQY1nhVeE8lOTfTNdOA
l5efvXCg0NYx4secSqUeL0GFpiubtY7/dyrEhf/v0mg0/ZquBIyL613r49CuoW8b
/uqSpC8nNbJ8n8r2RRkbtiRJKj8LS1cbHFflRrJn0YvU++j2TmaZdHfQYAiybI0t
RUUDhJAQiUm8bv6CyXdQ1OdSYrwH3SeNuSOXNyzUihZCXwNQtzVjO8kgcO4Ec0LI
fmepziP16tVcKpRjtB17D9PPpFZaLE1itwxdsU5qiejeRPo6Z+TOFDh+V8CjkoJ3
ly3krLksARFjXtmGO85dUW2NYFGJKdLgAlm3KW8oGs6Lozi84ikH5xVI1W+c+xU/
uLgVP3eVX+nRIMzIT8GkuSdDUi5pS7Zpb2MPR9ENa10Eobh+UlpIqxC5kHYlcQjf
+M1q0BjKtuA+biBfZzUtieamEjsZ97HmlU3k1/Po0UTEJAtdIaaJ7ckojdnlLi4L
rrzeC57KsFbLTwkf9qQh1nf7hidoUo9Nt9eM4yizn7hlZ64/SGcXaWw69/WE+Z1X
Kv9BSuM7yuWMQzlLS7voaektlJnyo84iSiCYzhhftzFQJNkit989jKOfDZm6K5QL
nbNGAgvahdXjCcffOv5zSbJnMez5bPm/XiRCu+iCK9BEEatE6twHoBxc68by+RO5
1etpZvEMzBHNHy4YCvDyo3Ex/A7XHjc3BvsgiilREEsVCIwAaFOtXPl5cGr5MzX1
KZ3dNp0TPgEMlHZHALIEsQCWuIBHWmZ4jXYZcIQ2/cOlR/Sd4Jvt79bQETYsCdGh
cOk/AgTnXj3wkO3kpP3O36UBmXKauWSafq4l9NMHw/syeAckWLCYI/SNUaBmXR4L
xzSlPfh4mTbLsBX+5KDJm3PHacTu4l/fU3/t/aReLKBmPE5MJMMDDZIJ5vQxJF2K
Olb6MU5QDZl48r91ZAVUCAfXpZ2+attNNAuhjiovGRyzqPtmMAGVcmdcGO64iqSH
V9zsgc3/oKlXOln45g2yYR4AMhUaOq96s37pPkmX+x2qRPylOqZMtC0Jhed6n9jj
Sacl5km0TWSTeYCxK+Duj+GVyAaT6wGOxPEezAfTgoOIN9WryKw6gfYy+B8RWrP+
iC7SDQYL8STvN1Ri3KAJ9MgWcAP0498cjex32sMRfsckH+//cadz3v41wEZbod6d
ZBgRoE5UJYlt2M0qvxciRM773aUklam0wgiEadZLXwkQVwAr3RGG5+lfadN4D9d7
nnuLwYi6LIDdAWCJ9tqoHcc7X6kApI1Jcvbfgeg30wGjvuQnv5Uw7D4qwHj0rFHL
+czzJDHnF08zz3bxttxONddT8rwPYZTsCl+IO6uoZwa6OQtjbwocnVotnZrpohby
kJ15ZWPi3TxOGEuFdX9Uzy1VM3IA5S9wgdqE+eOZMbyPMrde9Rt5pJ1eRITctxBK
MgbNsCsPF6XgDeF8/shb/OELh4tu0Mrsd+kBB1eZyt+FID+h+pg8KpUSC1HZg6y2
OE2jPY2wpVse7p0dFUL8m12LPXuEMuQAEZ3NGNn7i57580/2GGO26BsvnvSfsHZ1
px6XNwZkEPvNVX4OOIXG6T6TRPQkee69ZJfNt5sblpRu0+qbsHYl44vouqhPv9bR
tfTXisZSIJVcj2kw6HBFl6p8r4rZvI94V8aBGzwEb+dMpjoz2jLxthOrSENX7MAk
fCsPa75tm9SwubDU/NS/GruQuffxF5BXH6S1nwAIJLlkCazW3SvUPn/x5aQMr3S9
v4mf4WykKCypvvqmtgUszQThb1Qi4pvOuakoGaEPxTkZpeM40w3lzemxMgCx+GSD
56vvB3QIrBIgQ0w6t5r0T6SuR/0kOI18YhqL1a11A2eDyL6crQsNarokFaTDF/vJ
D8cD5xn+XnXw5uYjT+oj7ymrJndnmOiy6Lewtpenv3ersGxE0OYWjQKA8bqhFrVQ
OwuwAA8ie/7GiHOInAe8kkC4qJ2pap17jfF/G+2X3IuYw7zdkDcGjbeOUnAUJVAX
SXWzp2Gebncst9+c/dTEu5gFGGtfTss8xzWr6Zq8v/7+iV2yAMRO3RowXU+fD8fU
YP9RvWgI/P5YPryG9OgCcgAZAQadsssKRT3BEWILLf35ut+3DjGjYHEOaWBecsDP
N43zx6DgAR9yqc7SuXXHx01bkDOLYWVZvagmQ0xCRf0MlGNIpM91OMjnUMpfwGCJ
afxNS2x1tJnITm5NJy5B33U5SOR/ZfnmaRfHrAJyfW68pLixaMeXEiXPipSRfJD/
K1TkDSyJMBqSy3R3ei6EfHEyc17nX78mOvnF8f2LsUy+es0j4NXsrlj5stal4jDV
jOMot4atxar55afP2IIQ/8Mxrbszw/90728IcJ5skVobDAKxtfKH+cUuQW0ea9er
yJSmVmADCtzUmfMeZH5Tyv99jgjq+RrtL1uFSNgofQFctKzudUHBOJOHA3n7l+z7
J1bqQPfIv48w3HMy6Sl+vaPYowAzgPjDTX8o/VUBBOdbGFypM7+DWSkdV8Rehv1q
OuvoJaBuPr1kGxaTVTofaGj2kfNaBaFaSBXO/ydyO3WNghuDi4hnsePwlSoAamBX
I6eiRnvj3FKi5XBc/C9wzHlIT54Uhig56VbCZvkN0CxJAlASOUPm7ZbX/znv/yHY
kXXLfFF9SWyeMAVdE7W6zDrS/JUZpaLaQPyfRuxnPSHIY3WfTRgux1uOHfzDi68J
t6+6x1c4G6Di+/Klnf2zDz9xLW3OugcQganCgL1KpMMMcjXa2ztfNZeevpUP1ayh
kbsa5yEjofyn3DFA6mdSmQYeD9yxQZrRfNRXwfTEjGp/tovA/z+s7jlMmH3+QhR/
2o/3SXeSf14seCzh1Or0kvslrjg7VZj4DWOBPyvHjkKFxkF4tbUUQP8zcevdsJdo
BO74jTtehyxUq/vDpnfO7fD3qeod2BTByfQhrk4f3y+Im5Di54uHnIYYHIH1ZTXW
cUjGAFfaCsBrkOdiZvPjrjZqW6Ca1Vs3wPCfqztFFERfIkiXFY210Le/iYJFZLHa
zU+k/I4iaYcZ6Aoj/iU9f5NRnXE4//0Z7Izef8erfYGaRoBsBN7EFAyPvjKFk5Tl
FRPoheJVJ/tLplYtYLHdzo0c3pd3g59lLmz6tdsOifoz3u8fkI4cE9QJeM2sbT8i
yM6vZDYTYgrAl3vU4oDzJOezD7Ubg8ZTtDrqlgtqg6SAczeDVh8nvwl/4GjJ8d5U
1Z4gX6lbONw7DCnFPkvzpV+An8nZnuqeL4YiAWNHSYRdi0r1Eut6MW0NVzKjrkJ8
5buGGY8YXTvp4LDkHbbV2D1hIziYgQTuhCEq6/ie0WhFv8O/5PD957XEskK0uwgk
oIbbfZ8W+yvLWN3ZI/D7jhJAklk5uRXQmrHs6GjHCP5I+R/sA1j58uElfcVmpBtR
i5544NxS7s0k0y6Lng6jASIuUrfWup0VCTZhkH6NM6uA1sp64R9UMk1weidimISs
t0qudAnnUWcSfy4E+e3ml5P9xPOZre6Nsl27l93gm5d5kUulAf5a5lKRFbvhNQox
vn4vR1qfASxjGbwAa/y8cRdLAXBKmbt8PN3Ew3Z5Wl04ACf/CcNU4oQy6KCYqXTP
gUdWZybSEXtQHJjnQiNK7r9nVWzDDKXzoQhrrYvWR62quQdXV5ZIvhDccSa6MR29
DAh+VuxLWVG5YdmCdgrQASqsT/DehsVjLNRJ5V0fWMsa9nwc7zvLk7m0uqDEy4oS
hGIs4dHGdKhcJ4qBf19uKNgN+xO1GFhdy2EvRoYyZg6OB+vHUz/zFhmQhWtZgAQo
TxTE/gR0nxGgshv2F/TwXg2kQhtuUXSZTe6+pFMxwliag1EZhOCm/KkvQl7QvSUd
sSMyc5Ur9oZQONrosz+E2xGipjdSfqnGIx916edbJUNdhX393hx2uWoJc2KUI080
WHDekYYU7s52saYRyF3IsDcT7Kvc8qftQxzv62KCM9j+mq7LT0K9fww4TKROs7ee
MwFuUPeyn1292bwDl1q+D+kitZr3Z2yXViQlFeKsSLyPwMlFr8sdP21nTCixCJLm
DRB2FXSsKb7Z/CgCJ/JFFRwGRXzoOqERWeuliVvyKA+EdIw1/1CwZxo9Xka6N6QJ
b6r/4LqHgoIKLkyvD9VliJYTUs2JLGUWW5htE/grl1sAqh3NZZxpEbVug3DoVTSU
iGiFEJbqlmedA4HW5TaTJXX9V+TZBWEmitWV68EmNjwqLb7Eep0usGANuizUb0BX
c/wGeLBIMqdCGzrXamuwvpTViPBpUdRhe7Ac9aB74C6upNEC7QOsOZgYP/wsA9s2
7tK0mepwGqT7YCJI2mLUq2tx8yHJG6MEmGHMvVIEM6XxbWp2vc7C11ZBzcuxexKp
r1tBknuSXWEcgfVKBiU9G56Xwt/45ra5P+B6X5/0fwhmoxXwfEq64k8i8t1rGMG8
29nePE7gng2gh9QMu1SmjTSf78dyiZxpW6vbULC/8WCyJktgv5HsZrgwu6rMQ/SO
LmJbTvlyU8TQbtcDRdewIrPz1OcrcqUOfC2cHkjjZ16tb4CEPk6G7DbKNuoQ5PMx
WcywriDEMLGL/ioC5ihkoX0CfBoGRmyeLnXJPhq8m0P4YtRD7wVOXoxCLV5DVTIi
YvueQLg1i+TbobG/wxITsGfL4iAlCeLCCzLfRM1BPnEeMVEEPqi8S3MKESAEynqc
/wPE5RIPodca/DxdqeJXguSkaWqK8f8AyUKx91iEFEWf03R2UxKA5mg4pbXfnh5F
U0OvFj72pZEKkn4aPMZIGRlfuKMWj8hVCecCvh0qSdu3DJ+VBWRUFNPnVOOPX8XS
uTZdZtP0xSar/LFBR7IWBYISOZlGBJrkfH93XokI52SGBWXcNX7ewuI7iHokE60T
wM2m8Qj50S7qyPV35197cE92mhmyShkFlBW7CRbp59wcfSbS89go2mdvspoTQCjc
D1ViYp0w2VsTxVd63iA/N60xhlV9XnaBhswbiUWvWYuQ8yUVMt9NuJBA0vC8FzhC
XrhNultYoRjicu2CsG0j/4p3brbc+c/t6M5uQ1kBBIA7r9PEKJwayHbt+dxS7BvA
o0EJ8yluBz0i17fCacCo3JTmG75H3bP735oodq9CbyEIn13O8z9IC4ppCqP6N0l7
GZvpih84JeXGqMJ29BOkuq2pDET+bWnKf9EkAiAmoHUNqiGATv4YLJnGZfv1go2D
T4j/Jv/qPE+LQoAw7uwbm8T6cUNNr/PPiXNIu+07BnzoQypH+BGpIMwttas8CA06
iJzzo8+/d4RdDWIK7m+nMMXKHck8aWm9GRdFV5Dk7FCla7NB+2jGOL1cg6/F4ZFt
GytjpPSpyuhgo8ZHbPYQYwvnwpBW1v8ynAP+7e4Lq4JtK/gkwLPdy7kToZBd5wlM
tD2krtGX0J7YQMUuCBLHlqxWxsV5p9RgZnapppo/ZVbmKC/gGUTe+MIpLYWMUCf6
Dis8FXht81+hxIloZzIhESEZNqNwCQvKMi13UUFPAGzvWcF1iIZtl+d1w25FSu5b
U0988H+BkW9S+eM8mcMN129iSUNwMWWJOZsnzteJZtf4uPkLQ9ztn9CenW2pIXTZ
dFOoWaoGs9JupZropbHYCR7a8x4DabH/yprY5TILm4iEgJXYS1Ojj0kBuKoyZeUA
670zmADQVoBqHuHTNSpNH3P++NexVI+2usUpfH6citoyubEm+i8at6NyvuLsWtgA
IXa15oft1HPkod4tvpgunPRjKT8wOKp9UwaK+e3caZbipMGV3DNiX4oVSjZKecdE
GWoX21hHPTyoZrbAkxuJPgTPxZmLLjni7dgt+s4megS5MP9VbdrfSin/XXdpcnKZ
GBrV4+TCKRxT3AGQr4x2YH/VlL4mY8mK6soyoWW7xVFPKmsk7icqlt0rzQSYsjmO
nbnyfNiA6iOEHKOnKgYhUlUwrszWJQZZ6frfVSnBZA6tvo85pLWlA9jtcn40oIMb
LzFmbg05vUk37rK4L5Cud1uVMrfj3Xij84m8nrinbPyBEDpSYt5vYchP6vKsLDIY
wOHKpwFB9BB1MPx3174pMRW2uuwyvwGJWvKhx8QQrBhBijvZ+tsApGhCD4A0clt0
pp+NdY3kN9Ycl4ehlg+3/vuzdA8a+3SPsV08iECaBmahdYsB9AG9eH3NhpZwYIcU
SjW1WKYHYunvgqNIfjv3jYHjOkwgfICaaNfDm6s1FAfrbu0/GPsDn32mwCHxO7qC
fv1dIAFNbWWZqQ4rsocBBOCU4FeC3nMc8o/US5uXG3y59krLvigJ8IlK1oWarVwt
H4A5lE2J8TS4/SOLBnir2MCDVub17KB9ED4B9AlTnRSgaJ5iVQITxWn9IcPyxvcy
DDCJhorROralm/slYcOnEZgIuK6932zLFTTXbDVfq8BH/fV3oWFs257iB9B01u3B
lHyywJH61zndrVjRhOrGGYkqusJ+eOhtgSdqNA+73aEYme2jnUJiUgmYvze/IGlr
TZYPXbeDGvHSRqK8bXWYxwSg8Uxy3GOkjJqm/qdCLmR54fSao0aEdtKw3nxi/cyi
jyaHUnvaOZP2q9zWUwce+Q422VqEcXwf00gvOPEl+LeDW8cA8S0rqp2D0B0BtmGE
bmYgMDJf4HB4iy5JCZSerqbtt7BbSxG8ASXgiW2AhQVJvIxVpbn6mqMlV5F1B7vO
H1Ud/0vzxZy7dS7kgO8PDVe+Omkg5lTslxcUACseRbx8lrT6bfebGtynyTXZsh8W
RX59+ty5PcJm49cwex/wP5D5NxUpD3+AFwwLSCMWXbbbqLqd985aLVXfSlINLgZH
kmbgGZkALsxjDdwf6Ewmya1atbxQRm2JNRp4diFXeU8XycmHSYMeKDax8G38VkMX
EWk1ACg/Qqy3dlQFJJzromtTMV+UCqeEqWjoAgD9eGoa4BYd3bd3qQ6pM7sZQxA+
WQQG5s8NGumFX6UXvqaVaQGMBGVWdBp72KKXl+qflZevroNimAVhXXepbqDmQB8l
rj1XKhIqQcX5xFrcA+uzf9+yAYVp7/VqzHkieXf8FBVGfkAgTDH41sthFh80n7UP
krUnlOjQVnLpPK73kaRl61stGyqgiqHMC1766Hl2RiV76AaAoo4x8y7eeripgi4Y
fL+nJyHrgUgQvz2luo1bf+W+YiqOTV6O/rnhPuJwznvIK8q30+jia7Ve32JbANJE
7vuauLrEvIAaYsj9IFbNqXeb85dxA/839BgOj7SgsRdc57kO3D+UXHMGljXITadb
X8dw7xwtrt1hGFItf1LVFIOCZVayjDNX+LmBetfp3iSmND0x+GA6WAbHGgeYcdJ4
ax614cEO0huyJQOWahrOKU9DEC68PwjOtidlv1Roca1TxmP+JRx+OGzDMWmGbmzL
xVqS6tpVe1J+cjhU4/g6wW6odQO2upvpkmeVf4gbVv+EifjhV4ADiRLibtHU2cFj
l1XQNqkgPloxVwi6uQOnLb0K7nBtkEWbkOYncj/X36z1G6/fnEkI9/4gAkpRLRoQ
G5IQKf1ey/qHXHDYgy+YijST9XU4db2u8rnhBLXiHBINWuGpvbOve+eRNCFv77Id
vphSucc4p31S/Txe6yrabPv3RCj68OPtt7gPgC7qiAMrS2/EKLP8ZODWzb3ND1Jt
U6MJpDEYBCOPWnf7Zxp6ASnwbxgVkbzXM0EGhBzoDzUFhQhxnlUEtc28vqP2ZnYF
fKifLg7hwn99kUaThLNArU4tE8pP35m9X8TwXP5qeY9o3MOyutO4kKEZlRK94aMF
iK6b0Iagdt10o/PoXCi2yRrQnYOrb/WKXW17EaYDYuFeS8ayW7sMXagbulo6Odgu
rfPWH8qJ6a+kFXang6WGIWHB5SMHtN1Qm2YwlvUVNE8MsWW0Oe4VGlCq2BvjFZUt
9fUAHLwT2NPFeYjeTxWJd3DNZRtpn1bdhXfQG8jXn+geYVl3Dt5mzwae51dbW5xc
RHMsy5AHEXEZjfC2QTbhViVgn1JpaX3mbUur7GJXNtuGg097zxpNHzKgHRb5b4pk
UHv6UUwPXc3eLhyyYmuPIEADmRpUPg3XHhH5WjWAdFETrO24CixquBxRWFI75cf/
LsnID0A1e9+IVuyFMtABM/8+9fM7MrNow48LIRwCBlUzluJILkX0uZO/5uIGyvc+
mCHiBbCGSx0vAzJd6OZiyJyyIQc1wWnnaB993mn88IN5evGxoPHjMmq126doM/JA
GIhJaC2KQ0owj40C3GpMtpdqNOgMZ/lR8rqljIb+U4tw07qATuMlp7snlU2Sa7Op
LmzMRCZ1nYauRblJ3qEMK8sF02TrBiEqH0XNDwBsCZoMFBafqsQsPaIF/ftZcWwP
hR+qzWd/gYpGXgJa+I0hq1dZmQtI78Sjh/PsxCkfUbesIpaYJzlA4JWDs9v3snd9
bvSbLjo7GPZDNaN8fQDt2joogQ7U8hbrTBKtSF3muNZ5gloS0mBDP8sO7WNh1j8S
wQ6CITfx4WGUGiOpS8i47hPvjxs1SkV+4b8p+SEw1A6Lq75D5OJTvAzwhwrdCvhY
5+rS89H0QIlWOFz/lQvB0n0dzHjEBdAtb1wnF6fnDP8gKCvZ2L9gU7aD1xsWGFKe
13eHK6wdrVm+woAqA0mYMlF4X0WuPGhla+C6eL+T2TiV2faw618hp3nYEy7Gg2L/
VWlBalPmhJNDbW8WYCQa73gY6NSb08RbHeYTfrF5CCTUjmqIMVOd+rGRzwXjE0NM
hUXIGdbrYgh9yfuH5r11V8Jy6w44nZJUtlM9LvmT8fZhtl2u+RBqorLAkqAnm8Tq
wVKGjIxTEaGbIqdO0xH59/8rQr9v3luY4hf5FP8T8E0NgqtRHj7qGIuHLED4BHHC
STc/F51ditU7+2bxLjS8VTf7nH/W4dSlpP1sBIE29i48i/URLCKrJALk5VoucJt2
ROwX7/pf1KqkB5YUCOk2U7InN5FSY+GNo7/C3F48AuxGn/XMjcbBcnkl4C69UXXd
frbAg7TBrssQJy0i1s7GxtjCyvlYUbXJw4hVWevfDullrBprhVSR3VvdrP68eGX+
XzyVUI5PkkehiaF/gM1oXk6y4L6kUOvsgQr+0O+u0o31jVVst68lRzcDi4sqDHtR
FHkNZZBBaG2mW8pZqCtqu63BZ3/HB4YLwN75KtPDv2Aa0XS/mwyKIMVxuo9LNt1y
ypDJRehgVEXRP5csmogCG0KM391dk9rmn6WAexAZllXTVDpgWuVSzmRstaaxTDJy
GVZLBi5AnihTfUqGPBudy5gz5iCNitIvntvOx5PD/VWxHIJcyBESOu24noXG+4CY
gqoN/lDFZAsbcQjgPcZRDNLzJfXJWcyGptcT17TGU3StJWtjcNNTek5oidsu5VKa
W2X9EUIee+oVOmfToAITGpxttJaQlvqPkdfr+j6EUpIJKirN7Qw+MeeOLE6WmeSD
1xhjxvdYaZJ68un0vXYOm5go4V5VA6BwHGrHczDgoOiGMczA1JLkSYOP/gKgR2rS
4EC4OeU09MdT+9KYp1f+x+F+3QrxWPkaWipJaWfDPrLEwANpHDtHI3r7/CL0lWib
5eZgOrvSIFcV0W0U6ovi7KZ0w+wB0MLxAHinM5pvcIJNpiZypSAgexvbghZEPvXs
ME8ZCM37O6MG8Rv9YF51Uvo33UHgyMz/jTgt8ip6Ip27ye9WRybxTKN7NV68/pVv
LGvf1gKeXVgAt4Wk0xzQtubkZwbjdQ4c99nvFOxFjyucTLA7AZjMOHbAL9w40uhx
qZh3rx1JlMIDEtXtPOstlH7naWn7egiPgUWzvF4mqiwRTZ7dXjJiQemqC3vuTwdI
BQ5lNWz5QB3VM2oa0lRX+A9lj5pIeazPF2/MFKuaTFRVBDzoNZoecwfPZsuBnTGq
QLqkKIWadnGKjbrwvx1OytU85jm3vzMRvYD1GSdfmr4aaDGBfLI/4xvg+s20FFe+
SmWJ21rSu+bY1DqkGlJg7sNWeAro/P3vacXgZWDsNoTTbD8hTRrsv2aAX6ZxJTVI
1KMflfmSSvMp0wJKf12cMoFzjVDaLW90hIUPLI44qujQwBscYuKNm+S186Hm+K7U
TDF8iRtgrhpjUUAwsdxQVTMvxrGg78gZ/DKZjd3X9435GS7y+2BH4UOmV3Es3p4O
Pn9YSZpKhb3A21ZBR6SbmZMgV/YfnrhsGlvYVelefL+jTR0LYZfUlRHj6OWPfnlb
vLdR2rRD+H/XV6qtSH+ybmGsgp2gj+BR9geGb8cwyKu11C3+tK2KhAYtkIoAqxuU
6nkx9KrBWkmqaKn0TEkIW3qAbj+htUPto1g7JHwLgx0Xm4BuqCJZ64oQqGtx5wYM
/S/Y+q9dy+tmpmZbPi3i9BDCQ4Pk3RGmMh1/xTfvnOunK3OzBREj0SBHmtcPrOJQ
RIstgyQ7Y4BpCgAihDl+l+sy70Uyrl8iYXTzqYuzPIn85qy9yJRPrK2f3O8BJWOo
IaONp3JAHakc0JKXnzms8Xr0qy+l+wMcb/GHiTs6W6RXpemOzIok4m1gklCacuzl
KMGhJQkQrslOoNcKijmQD0jU3mzLGBnbX4HNfRQTtshr6f6/4OMY55Vd21rP5Odh
+JfN+HC6cqxvHV6+Kvfs1yhA38lisFfPnuzlr/7FPFikRnzoUGCpDiLBcunGds8H
b4QHCzpJuUGp7g/tPpDxcDgWIvWuS8xtRHaa7liNxBUNH3c+MShtpepbgwJRxt8s
wgd+3SfrmMHFAJLRGzs0yhyN4zCN1+0PT4HMHGhRKW6wZRRtKA0vYHlRU9UAeOnx
x73xCopZrHGT6e3XtPUUpllOA2kKEDFA1Vt2rGA/YbVoYPdKQzU8XFyF/daP8xAF
XLIScqKyRCXBiKJ1efox3cVzwODzO/8OtIW0mvuHIlcMT3r/oosgqp/sFNd8dhyS
zNu6YAxVMgs5D6WXc0cQ6GcMVmKDgl+jiUO1leukVq0nr5hUvT494nBsedWOsaQW
HobTKWc/NYdTI0u8dCGI+XGqFIXq4Q2iwRR+hlvuT3G8lOFr6/ftRyoMAyEG3zxc
s2vIaU87s9vQTbc2JPT1NLT+Q9htPy4SnIFRgQTZWPB24LANmhX+y+EQJo2xUjOA
maBP/Q/V9k9JRaMFHsA2KHB+eQEirgbQj4QQLZn+E1Nm8EmmunksuXnvrrcRxn0N
qQW/rGk9bar7b1e8EIFS+5EY2t59JL5jF9G5wpV1NcG8MgXD+jqUdXyBGNmzAmGy
k/uzjlIyX8oK9g4KpY7eVbkcahz1XNSoKMcMkpAl2GKz3UAftTl5O27EInw6wcxx
FxOzg4owS/KH7WTZY4nOJgDHhoo50KunUzDTwbKQepJXnNd5Y0qpnL3lfSo0LVbU
eSP20kfqocZrxuzonK4ssnPeOCrCIccU5O5RzeHUAFFBqb+U5GQIDhCHh/KyXHYg
+4J5opiIy+gV/VFu+GcLOyUJ6Dd8MIIsoijbKLwni4BAhau7JR3Rhaups3UwLJln
TCD0B6taxk9bHwXd9bkZ9fUGtuQynKVkghrFNorHL0v7nZhS0n1778i/fZLBp2Ja
1K8zj/8mi779ugo6dk8jEwX+NafkjPYYiHc8I12Ig3MLnGb6mYpy934lH69JZtIM
oWHoyz42Szh+lEhcvVhhEQ/xe/OQuDiSisNVTQ/TT2dUTOxaiPBl4UXs9pdGbK6k
T2fvmGjxygM9i/ZAvfV110ty922deu35yAgThgSWrqbN4J/rI978HurQxre3Ys1o
a0QMODrtcr/tv3CEGij6smKkcECKgzvMphx1OLK/tEqxYdLkc5fm+XFn8H7+zZZ5
oewdmQ1a7vUuDXJYoF2aRUV2AMCUn4H8nlOIuVsRpzzq/cREkNxz1t1JLsgNG7k7
6fi7MSufUuHAkG0kKAfE/EkKLf/ajIfR/z2Aiz0qHvdTTyw3bJMcbzLeYuV5xnXK
B7HoMPeMN7z4ajTbGbE7xnSs1JYA1qBykzilKxkvRrvsQiBjRj+HgDaqIWIsRauc
KDjljzl7ZJsvS7Ijc6CboLmULHgIWUgkMscWpmW18oLAk/HbqmF8OiLIKV20TpJ2
QrUlzQpnBXccy5DwO1MOtxxBARt1Et8PEv1iNX+aZJFrEENbKKcmwhRNux6UbUzw
ojp3F8cXgo27saZE6M5Klbj4I/PukOtDSuR3XKCjCbSI5r2kVrpu0jBrHvhBKFWX
xz6JjwEBV8pZSUDtjKRnB6qPdgdFe0sWgoni3cAqwn5mcuAb556vJ9fvOwF8iiSO
9LAZYF8HOhG4yeqwijEZmhkEjzqoZX4RZGmh7kOtXQFn3gNmlCtkr4d4cEpHJ+3u
LD+rEVhhhYnJU8xABxAzDTG5xOrCUaj9yvKCgL+c6U1qgnemVoZ8Pn2sc1wAY6DK
6xGxdGrn5PPrtn2PSTUJ+x88dr8H25JEaWhNOjjjTyYWw2idsXuAPqR9JXHLjJMY
oxP36a37PPLzm2qC1I9vvILzMshN38jWNMS1p9/5DhvGoWORne/2TUduKtN/uffX
UZk9IwXw4RxlZZSIMaY1QIp5km/nIwUnWapl805U3n0voz09gngQ3u3nLmjkRXG5
/V5ivEasRRyskybQIWRAcTyLmj9gtVSJuaRbK7KGH4YPW3mdTH5vQewISgk/8xWL
iws48j5budCj3K3aW/q2R8LlCIsb8L/VVScMl/bM6SIEfHNwlWa7ViLEpDqVEKv8
1vuNTpHR1mbZh/JEilMVviJZMg5wJvAcz36IC6tfeA7xCgibOVhvyY0aZZvoMCcs
t2BQDrjJClA0dznvIuAAe0/1yTIfF+QhO+XOnqNDuR/WdMDcHO+Ydu3/9bwUu/jk
iU8T6FQ8PlSpURVf6UB5lNI9qg229UDqRsyQ+Q/4L6pXrOt88RheF/UvotDJVHQA
NPgGkwUOA5R85//m1CauzB6kDLnDsFQm0l82kKwNBsD6m7m9YH+canhDtAPYwwkO
COjXni1QtV/Nqa5N/AJL73600AEsDk2aNl8+P7o8il9GzR6+Wi0DlqkbPeqQH8IQ
aHYNgRGwbDyMifpRB2oMxfLSwc3npWJFZ9kOWbOUmxAuzs8k/qTqxgNvosvvGMIM
jQ+uDpv2DkhREchtUILZRbyg7SOrZZNvl4+zn7XSY4WDIkMcWrOWxzzaZYGOQHSZ
mXvOx/ObtXDGmDai70ifuHWfINngWavd4R7Caso4FwWZtCjuQvOKYHh23zH6QwAu
u8L+DmzGDmc6osU/uezOUUBnxYgwrtZ9TTO4/BSw5T3Ywb8/LvHeM4gegy8p/64b
ANNP0I9B0Wdcl6HzSxPd+ie+Nna2I4bRYcjQ0Zh6IwXkQHq7tY0o4CCLsEv7Er1C
5xpSWsWSixajQw4QjNM4WBe903SxkaxihadiEgK4eRm6vKu27MobRB0AeHar9CSS
GQYhB4cSMrc8F6HyPClcLahCCCyuKeF9nt2EoA2RELQFERJu7lFUaZJOkSB/JOkl
b4LLVEC36lwmeKy5Qk+rLBvvaaTV7/wKDZ0qWQ5ATopOfccwP0jZV8vy1yTa6pCM
tms2hMo/BbK+yTPousMH8ePEWoS8bQUUjXn+iCBbpdJHxp2UytoJ9c9rR9yg2wXl
EU9u5nPDZGVuhYhnZ0ydwD0U7biWHdh9OYznA01I9ccQuONGFK3HvfoDns8nYQ/k
nzkEtwNi5FPfUcU8NEg1/Ge7/HtotkAmmrzOu12XHqHCrYftkNtO2Z+hRmZ9uGjN
48N/QSPDy69ts0QZ93jT0DhKgkGjSs8DVDgL7tCogotEfY3n+eLxXylhBlppKXVM
So8UXQw4Nldde6djvJQrJMKmshmb0sDSY4IDJFBPDqPilWdDDOEDAAn0EF4ctGOJ
YsVX9tWb7wf/SgfOKlTbzE72w+JjHBg5nT/VEJGqT4QOGTZzPD9ub5Avt2UnrMon
CVMN+k9CrbRvzKhf2nKE7L0A8kJnnPMElEeVQOKRipxBrF26uvu4x73qXW67CRC3
nFjJl2//Fjmd8r9Y5WlExy+8eijPaCu/oqjDFv/3nbBCl7D2DUmsNRaaIuh0pvqL
CCqWpw/vQX3CUYQUSPEXdMgMoABxFN6SRzhkZKypQgnBjqfVhZJKok2TPAAKpxLr
R5Auc71yURvA9TL5Hz3JAIaXjlOwfviMxdGPUq+rl2jiK5VeOk1naX84Hm9ZQfvI
g/CaH/JjrTkPCA12SK9PiGr/WTJqwpJR9A+MtZ5qtl+v+2mPaxQOLGZ3lt+ArhTQ
Qf2FBVeYwwhPBfx13EgqXSSkryY6M+L+j/73zfIkTrFnn6+HW/PRjZagsXeI6Pvk
U370XWiwnRDB5m5aZp0YrwEEkUzWfBBsb1jIZJseHtkfOjaVec9OZQnGHxl5AAkj
YiwWrZ9U6lz2+1yL5pexNrtZ22PqxEUPAc+LNO5AjntrQuo82R1MCkvzrPHH2KjH
5uNDrSubF3xzRJ7fuOtd7N7QduK1xz1rNfVEzJQxjFRGXKEIdfHqyZ/tzndCXyW4
1ysJ6YZbQaiHU7mGDmVBeZFN9j815NkPAdQZNos3WiGZMk3mkLTWysiTFbUOnf5j
LzJ89MkiuyEuM6hbT4YDG3Sj7DSThteI7+0jxQXxfwSVPH+PL8M7nG82m+/uiEDi
KmOeE/tBMtOwe622z1L9Ns2VRKkwm/kzKcuuoIASKKai9ci8lIpWyyyqIFDhssnR
HyF5elVjwvNq03hImYjMKt2SKxh/0h+Jr4aBkEs0pvOxFvIgwOv9z8hPX8oAsosj
xa3ysvOavS5X1f/61yghh5AkOh06HD5H3wGZ+VqPhuRKnJG82crHeEQK0XR/Y6qz
CSmB70wn8HZoGXE/U5vK2Es16V89tZ5CqKVelJDKsfOltW/NrRQqqkMQzjoQzC2K
LFhPfK3BsNu5pa5xrIqz0eJYVjA2bIxrQpj5tBELyvLAkP9l25OgjkOQTgVlsR9y
yAXmkmiR2KtwX7gwT+hwlu4XzNreMsUB7+1atvj39iwWUz9VEIpP3i8B9/0lQ9mu
vtM4f5l0u6zB3kzYZO6wxIehu/RBRyE4MnAxEsMpDWzKhujCuV7phjTAHMTzHimt
Mx0LRXfV+BjT5traQNh9+g3Ujh8i4cNGLhdr4CFbScrP17rAwfYd2D7VUTsdbLsi
UJtkMul/duxrK+XRvGT3jCOi14LL+GhcR4xHnY6NdoVc23JOupSsqhmmwj5GTFI7
kylqhSHBDR2zcJT/g6+iqmr1ORQEe4je/egwG5eRtXaSJTRU17+hUpzVBjn+6ocw
lcG7G7aVmIbQsfbkYmbNTFImYRzunaDVzEFIr19CKVnSDli+4XMGIyH+341ZC5lP
Jfh+TpNLpV8DEMx8L1mo2V/jUNhZ/Fm83cJold+pmdW8lSAVLNG5FMU2oOPS9bDq
RaE2XGFP1IDFFUu9AKDVgM5xz4tI3AiA6XEeIR+wO5xMms1Kvd1Yx7146mzzY7AQ
DEXcb5KvDabGQlAOvZaVwe1C9KjPhMawbL0FVyJHp1LT6ngEWxl1DNd6L/ggw5o8
opSfS7TjpI8ARLZWzbFedjUyV7pE0o3TLBPFFRpyYiqWBajRQwlZLeWJlBBcHBFb
LfPxKG9Q6il6RcYqa9mrpC20lw00xSS3ip/w4LE5bkFSTCo1H561FePdkfvZiYUF
zfhU8NYWhwCTSeqazR/1xDwNghju12EI9+aidfEan+tReZXxBVBCttWnOqGQB+ux
75JprLkwnkgoXt7KCuCJk2jpuUHJjBncGYeD7bVrd/d5cro0t+3vv8rqnOTX0KLS
Rvx6nlaq+3kWgWMTX8bN7n7MLjjLJN5N3jd4UKAjZP8LKVGOjj32ZVS3JxK6BOw3
DaeVSkzbOPBoarJjcnY3U9rovHg/s8ezXvm8JHe/dRjLNK5gvir6sDlQ7/IcmfY5
KvSGH50NhLHGzu5SjaOlSG6uXN7ZFWWtexYyUcuutb5obSYWegDpHuZvBJpXuPS2
PxeNVW4RKu5XAPMwb7rrrM+bYwLAZhXst9qhHcoAQOPyXuSGUL91oBdh7eqjGTPj
i8c1USjsAmxeiRqjgWpGI9GpiDQv+0AP9T4Siys6TiylbKCUnYNQzbuetO8N6tN8
WEe+8Ma+aUKj/WFluXLXbtJIwxCAXk2sG4bMuh2QQ5H1Yl9rjDPBnTsOlrxEZeCp
BPxXrVIDUWGy8yZP+w6d5GIonk9xgUmUcoVUXauAwX97LsBshE0z70r6vnXBJIxK
E97Qes/hrUPY1Sndlom8B9dOCDTQ4jJK5uTbQN+0ueffHsSLNnWt8I1m/zWn0odU
9etQfAQ+fFP/LmyDl+Iik01/TLQLIc0rBXb2ycBSnbKqn8CC86xXhshOWd763he5
mfqqtkyVFXIDkE8oO5CCB2P+2WmcDReCGN/wxl9j9gWHClGLLzc7uA7xhcxsqlfv
4j9/+/IAoutx9o8wGtbMYvkx4hWgaX1IahIwqym76OW559Ol4zirTm06vsnQMox7
scFg7pGk1VGO6/Ik/GhO2gV2IFVBWjoyz6orICQ1+kHiEqI79I5guo8glNCifsuV
a6XqVExd8o9h70bbWV5lYi6D6LPbh5kIrBXLzz+q64A85MBQxoequoc7bGGyRH2i
C0RuG9JFCPXtUwWsOgPxfDZ+va8/3PfIDooYLBcJ1x+BAe9BZi1Q4GrisY1TMQFw
9mwLsSXdGdPyDDHWrvXrMebTezhEMntcoPsAXOwOC4lFGHBR4NqArZoGTyX6pdbc
cb3IR9hXocdLGc2EqLgJvNgIsnHRkDr+F1on/lwu8ZH9J0q7tcXzxOQKsORHzpLa
xyoq9Mpt+y4yDzRxcarDYCpmQvHI+Rxf9SsteyHf7eByMTYV3KC4jIAzSjtC8z9f
EEUtGncp9Wz9gVjkvE8bsv90CkzFnh+XEB+uhpLuOj4D9H1FBaBO3yQBVOiXdAy5
/K3deZqecJgD8MWB5lvySfrrk4K2M+tbV0aebLsWJPjj+AJTJ+MrqVU3NxzmcXfJ
JlCISO32JZFrIAlyuRF7XweRVFtdeyLNAOrALCt81MQuBI6oV0Qb9pRNPWLOO/T7
HyZKUbhjNt8+8V2nHVOOtgx6twCBEUTR+LMxPZDhTnRg23Nj2ev94zRMHnPncpNg
qCzyD1nMhOz3z7o3bv2zNfMn2WS3INlLt1TY/mKWewsXXpvKytSZpHHVPcgosoBZ
uAp9qqWSrg1JUtp+3cxr7UsDqNL/naRWtcHs8xL04lZ1b4NHK8nv7pG/voIoG4W5
hAmvBqPTL/h5vfnLmbimrxWJxfptB8t5m0AzLz1IgeEPLXngblQLhh9D9KhRwqfY
4OtRZXP9unbGm8hNP6pc8lgk5jxeJVNeQVixDH77/FZLiJn4h49psbWU3qOmjidP
dY4Wx3Edz2lnhvzP1TOG2enPXnpMjnakgmwN3zGGvyD0ihDGMCI+qdM/OvKB1lBP
6ZaAaOflCDNSPVjGBunbiVBQJ1OX7BPYz9jbHANQCEYtvo7FtA7gOxSbWNMnBIE3
tW63FBWyMI1XLV6osHureLIwC6mMN+quNww33Gk5or/4WVD13pFV1jp5MEmTQ0DV
+59FPMAD6XcgbYTb9Xb/H8tng7EpF3w8fzP6k0pqKAMJMpzz5NGU/EfwNqQlRnl7
fw0o13xwBBBDeRQIFkHButx9KZvN/CvksDpTFj9TsAvjEjFcM6CMPLVvU3r+tvhm
3woUxAUvmyn20cVLuhKAiiMDIywcsxE/CoUaLaYsGwtlrC4n7kCMd3oMhQGHTU/a
+FGGOcoYIv+C5GPZVdp+lTjkAXbbWYQubkcEHIc8SJCCKMtZyN4R7hy5YID+K/6c
hJoLB7dz88CNHWyNdxFFy5wUHYNNEsh+3ByCq27cwgCW7tnemW+iqpfbSfR+XheG
N13a1BDKTwwFk9WfyEwo/bogV7AuOH8IvD+uDdWs+bBbpEwcwkrFGE9zatxgVurX
L/pb8wgu0mLekP5hcvLNjCaaC7BF6+EQIY0m3r07Y5OXJd4LKl12SmWfVqdymZai
0EjlvjTjxgDnX5rpx34wtO+1jZ1Hzp7o3bIv37if1nbWmZ0u+2ICVPvOrLy/zQr5
Ei9hrl2mLZCYpi+PT8bKBwBFu+doXLmFjtsJHh/W/Ijxa6K0eMSCTkrO4ytPUdPc
OaHEKjRPwGNbpGCWIHIFnUVseHIV4QPOAD7n7xsZhJiqTO/AgcCMBYgkz0WGRGIC
AsbF6XILFkQcPsQ2poNJlZBvMJkV2LyNe8L98kCo+B8jpB2cP5xpsUzU89yDsvG/
3H1KgGCIxsVtuvqYK03PSFMMCJ95Aht5Oq6EoPlh1XrneHACfh+Z1jxrNQC+CyeY
l76Y5/h32i+J56OblcDNiZ/83WIFJh2efUeoJ5bqTMoHuA8rGYPmRjAFVd/Cpp+B
VTx34LlH6QZy0EKcpTV4TUS6GpwU6qQ4d2tSXoI05tLopATtGfIbIUM4jX7OFHr/
kLBh0WTOTBvowAGAFzZkIUAy8MsBaQgGSUGCoQBE0RA5zJpagHBXF5SUWqrgz/IU
tMc7QtFJsotnY5aEZUlShicFyOX0QQgY+HSDQJB1K+Q/Tv4oJOSU0YpBG9xnJIfk
pgiEGpnrD4xJdBNPGIlj8nwK1Fy6crBg9uTrAlCb9jBq/yiL4uMW7m4wp4E9LVlj
L6zDmNGlA+jZxNDHEyyzU7SFh79NRYPTo8StP3eygqIsbPPZeAWrKeLPHc8w/gt5
ruXJJ0wVaZGV0SLwHED+3pxifHDiiMIXzKv41URUm6dcUTM63jcBg6BcWhoT6sCN
IT6mZpVgK/Alps1H1QcUdcnhnhxi0nTkq8PGKnA3WKXJRa3/cnUR1HirMi1YqxJV
8pUiYnM2mFqU4dRV5m++Zjbz+M2cgrrWsl/5/bhmOcP8C2TmTwXUCrl7dRJj/CgQ
+3FV9co1TFsZo9jaj3dCN038GO4BP0YWM2pOZcJFU+SYvd+z5pSFmV6hSbWC4JP0
2ofnrtuDuNdXRRpzttNzaxFa7J6Kj5ltHWXkndsmyiECgK7wJMLPY7DivfSqoMoh
WufVHHbGw7AJNztZBDWwzDx3y5hHdT59hbX+hmHMB+H2+T5+QLqN6WLfK3gCetou
ZCVYcFzCkZbSy3/qkb/XCHHoFCKnGmK2rUi5Fwjk5aXZqdtjNl+mQMIAskpmM8LX
dEYdYe2gm2FbRZn3pv0YeYGUi9yZR66CNhAdX8OUUfvCpLI+MEzCtTBxiuexc77U
Cj+gkQZpm4o5Y3rCzmTgDz1MxZjHt9qinUIgnyHS6IVzyfPIfQni0DfkGNGQ17/+
O65vzBPkse+OiZ4DM7XghGEcdJ0xzdsrT3heKm3SV8rjxUF76ww6QKUVAZ6+0KfC
A5C80TuVdGf9StfE5qKAT3sp1U82ho1xZTlfKMm0kuUGP6o/OzC2eRfbVeSDD1VG
QPN02gt5QGAr4gVtd4KtIAhG7aDZHRrQ8pGJ3a2fPHJIYnO4z+OcsnBDGMXGcfKg
oDyDsdGaDU6FUGG1LV85agFrZE98mOhyVf3IBAIunqxOfX2diXQijClrgGD+fLbT
Nb/xTwNNYmf1V1btpspJMvuMY3gQMPbMDkvh0PzVeFR9ZWArCTIEpnCVzGxQjqwY
XTixT81en8wU7B2M2H52pHrASMaUfcc0nEd2l2IQctbY16aPOBRaUZsHtQp7Xwg1
s302HzGkABdc9awEnPI4238y/RT+HuJ89b0VM0CsKqvFA/lYUHWRatjoubHgQ4xE
9UU/4jnaUVEVxCiOFTX134DdD++thceWUT9cx6Y1J3XKFrYOzJeN1QrsHTp0hMK/
x45cajUTmCvibX4MH32k/PtUXbR3+JVbNobwk23NuxPEJuxBNL+/AumrvHLiFGlE
37kP41S0in6/E7AhZXfwfFHjquL2SK8lFStZSD+ks3ueV8qcKzSwU5z8EA/AipeX
w/ygIUP/IrHYc6gBTa93FOheswCXgNLCcqfDO2fVwRgt7RA6nNvQqpEPTmS4RrYF
Cds8fg18LyUXEd+WwGE28oBu8Qvyq+SYAj2OV+J1DbxhesAD3/bZ8ko30x4TiGUt
5ATtvFbMygi6RJMTV2JCYOkSTMH/djbuImiZh1QVaI0udUlcvw6NLeGVlzNpFoH8
+9Q26MtmyL+CRlq68+dfhwK9hk0xNnDQZ3q5acMZRjJWZY/bTGHgZ3eJvKOLEEiZ
PvDuciRjinqVXN8y3Sx3AKjICUIKjJGEn5E6nCSFcm7BkJ5llcYDUmnw2I7gnS+4
JkeBUjC5JImt8o23V0gKhRaZPLL9rlGKYaKpIjbVUYJfosO3fAdmy5Og7C9Irvui
DV+i6WY7zNc9lvngboU1OY0C/JnwO31AbN/7ZbkAulF4XosXgJIooKKg8Cqvrm2k
8uNs1fZZ79wONpRFxNYF58Zx1gFNIx5M/QevRYQtGav+nI439kdIl5ky/FwnmEJE
odhWjSe3nIVSyNI2qtuCegK19rpixQai1f34fTw2aXCe/yUvmmP7/fFLLqdwgu97
Ie5yNR6Tah4ge1Vl8rXxT9KL4JfDOOfXF676zfu41+bgsm99LhWDzZm28sIKr+1z
4kEadRDgjPHcSRXjxfplz12rKn4W0I+rlZfPm4ycAiCgfHY7MafcQPk8HUovkaPt
qB571LLqnVRY19tHC/GHuCR/3oLwdHumd3Wy1iL332EL8mXOknmBbzr7e43/2new
qsAgqpmysY6yDj7oPdCDGUSu+VhYG2+w9BtWnSZw4UjZhcB7kw/ZgDe05F1YnC6E
aJkWsYaZpRhIa2f3IsBQ+pABmgyqkbNNIH9LwNK2Jt1kjANjkdFHO6A+ABNwaOqE
wgL4BjoajpaZcIpTXHhC+i7p35lr8TzUMjWrqEIECOrwUmOGRbS/DVWl4284dRwH
1uwrzlBBIopTc/c/6tm2kSJfiFUQP77RiPcBlDtJOdS27/p5kUiVzCbC058ovXw8
pfUjm78ewKrc/QO6qWxhzasVYYgoPncEnpRqMulUDKMSQp7OfcIV1x7PDNpJbXht
NNkHi4y0smuZBcZMByLQP+fahEnZ0dSLizB8FySwI0Lqi3SevJSpEbHu871oquWj
JONojJj0DCDRlRBdetABEDc5zPZIE/W89tnNvq4OfcAkV70aNaDIQec6OTujkfs3
sKLx5q0aDICEbZnRRhY2yb/k5+PK8JauMwC3LS64TM4qWRJhZopYYgbNk0QNA4OW
IajQhwMHv4LnE7Y+2afSF3C5Kt1e+5IPp+GeJJZDMTIcPmV7yS2sEHQsseoHi5Os
tD8xjmfgIL9xxWxTdse02yqtHx6ABvVkOowjNyp3rdXAEttCDkMyTEjtd6q69P43
rFUQgRA2/YF92BQ5gPmEusaSm2jW+a6MP9lJlL9AiAjyR/ogw84hqVUbdhCTVwHe
UOWG5SEtV9OETFVUkt87rA8kQy44qoO3SrFmdu17Wk0x+t7QZKA9AOLAYsygdtHs
0hyhVn2stDlM7nNkol4Il0IyaJqqx40b5+mVq0n2U4kRPXz66u4aa2QbU8WZJl5u
Vfe+P1bZkBrf14Zy4HTLRXozcjeBtPf5NTDBZPAk4fyCYHtsDwptzqg0odF2t+0i
5DMNO9RHW8ffWRjA3fQJRk2PIWXewxWZ+yT+DitLNTyyL5A4PpkFHar1Y0qLGxTk
X7+p2FrUfjEbIMQNGbGBkereikZLl/nPLNX2Z+sj6xgxTw4oyrYrn4ya1Hn2ihAs
o7xlZx5MZtXkORe3urW380fzkzbG1/bSeTRsIKD2kJ9GlpQuWi9lUIOwIdS4bylI
nLVe/ZrDl8GH29SVGQmebDNwnqe1Qv93bXYhEyXbYeJVj9/1FKq2SJb0BvVAg8Ga
osQtlSh8e5L6pD1JSUpN5rgeoU/cJBPc3jOVOW/7Whh58lJl1ROAkP3I0JDOxRp/
FmswOWYxqiQRF7yceEE+mtaAfR1ZYj62cC84PegXqQzF97Fp8Mkox6ufR6J3Jla6
+pvTyeS3Kq3Fh57Bj+PHWb9d5r3jOjAbD7qgZXz0KgvJj1T5We8O8KQroY5C2Yql
QV+YQSdxvzxVYb/I3Rg7j7dJBIGt7DP/FP5B63uyEn9aI0Z1oAK2JUaSKOsWcky1
TpUul07pGjv3qPwAFyJ2CDwIWntj6C/vs+NOwpLNpGjejN2HkY9f4oAIrdqiseTt
haRv80EkofFo6NnlTmq0JCTXTbL6kFLJX7u8YdJ6Ja5KaVwiGczX0F9zAECanz3+
civQ0yJoQYHpGwr8Xx0BKOW4qFtaLVkTdMUQKbaP1c/v715axtlbfKdJp5sHf4/W
SRPtuoWfz7NkyUu+BpeKHvGNoI7RTW7+N3kZM2FOACpx1l7LZGSOJxFyO7eeAgsO
OSjJZmPXrDTAcUJLAsJU5XEwA/IL3G81mlZsKb3DQp342BnqOQWokn2LOa8uMo8B
yqF7fy/GC323gceI6xLvUZVlTeWCY6CxO6v5aiY/CaGLqe3mzILjdXhH8YaGqjQp
GAwfuOf9sxkU1K2+iJjb0kEL18myrLuEMmY2h52zHCZdKbaUQNadN8vyFRU9LcDc
OTS6nFDWuGvWlZs2vkQwmMo4NxvluZXCgyDM7Fclhak1SaxqbSXFzvc2XGh82fRP
6g4m10/XRrlGbTmvvb8RDBjnsH5GCkIJKycM9WewAwqw0BneHrx69u+FTxnEW/LM
itfdrunNywVeS6SKaVfWlbT8/GBDrICxPzgIT1nAKqcAsomJtZbFCZJkJ3QNtSfk
fSQnYA0F8Q2tQwJSgKar/gIjGFSsO7Omq8p5ofY5n5jpOQkjCm2+rdQvPFSj+B/S
Dwe9enhZBqBAUZiqGoDf5IyzfZootNng/LMSPUWzKl8lj5qaUs1wWybnugfsWVEE
YcXES1NrtAJ6ZG6/cIuO10OozK/ahXYlTU8eB+MlZJ+CTkdAn0+f+QRj10TDtKJo
kFhfjP+HMQZjzH4gR6F+kTG4kq2gH4/wk0XkbOQ0A5BD79B5su191iO8b0GzNwib
nNIDtgfPvSrijuyZ/UpJAefl02/jfzKFSE//vLIOJTuIdiyPJq5iozjUY112wFz9
4U+ENLbLLlV13QgDMCaaz+vSuWoGCu1szn+Uu8yOXEYPwlVlqSRaRSUg/njZpynt
Sk0xJLtGkwYrI+ZwVTlbzpFbLvptmDjMytRaa6jqzZNXnGb+fXedar/h3VH66J3K
xlO4wuc/YkQmkPUUKulxntd5gIVtuzr6iyLjbjBsgndQbK+EiG+lXXMFuXbELObP
kHWlJEgOPPH3fjp8UfisjDJZQnfw25q01WzwNHAJABgPtGZGIikh6OwprKfFLwsC
ef7qd8bWWkqv+LoOFUao1S0MWMf1ukwuV+dLPfcjSfSNduCJy2PPDH6VZF7OTRAo
S/WQr016mJtjqiEMX9l62PPpDTpfIY+B3K94NdIXHdvlVH007hVXw6LQPaBKcnjl
hlJ+vRJVsBup59pdBBjxyQ7zQO6BRRoMb5anCeM23+je8sPubVpVs8YnHz37ck3X
oMza6tSdP/+gdziz2ltpe3EVU5uGoftOMzJqNVOJPoAdebJ4iPabw+tgku78arTl
GHl2O8A9W9Zc/xXfo5VzSdD/1T1Blk3d13mZgWRvdIcVOBpwnpYvsSEIuUunj8pm
5w1c05FOmZgyrOIYM4kYSqIOfapTtfQE+EcdDW3A0Aics6qqGmgbljw789VWL7gB
fv0MVG7OSTKMH+kmw0V2/tjm8V8GLwGaNv0vImPglWv1dSmrMwoqEl+2xCjyTOAn
J1N4jVs6pKex/TFthBcKwYsUK6LvXhpUZ0oTu4K52pCRUmpc54V1Ja9L0K0t1ALQ
Iuqkrl6hf7C81vZAuiVKkH1aN7PRAVCtPdeycu1mz/07OX1ZgjT/HSR59yLV3NQi
xwq+caoN3+Bxfyy/ndCJF4bdw7zdxTEDaTUzFC38sJVmD7cGTf/45CLxxPy8PnvX
BFf6VtvQkqJiW79JMQgwW2wSRFIGrvioRx2sfU2JlmNeiycBQaiRQoN93Hf4CKzO
rw/Ge7h3VoKFLmjhVXXwpRtGlWLu0XjeyH36w5hmwFS4WDUhZ88oJXwqccgt3LLa
rb76r8HnKVaEZZlqyIyVrHGQc439vXC2z6krDWJWRuNbZCQdiP2QktgKsW3AIDAT
M7GDN2LnZ5W0M6ytrwXtteZ6pothskUx1S6Y3XW4xtZ1nYQsCPG7ci3bYMYVIxWf
iB9kzg6j2Nuzx4A1u4OidmfY7RqPWx+8vw8N8TaI42SVgr9NLQLoZvAdvZfYcIb4
SaPkdqnExR4WqflZvJoVqeYIgJbauhYyolptxWAmh2q0nmMOBlXNQjrnRTNcY3bV
Xn+memLNM1n4SBoXjmf33r7fKRdCJrza2TGh1pg9/Hh3jnPxf27cjhPLEgWQkKuq
iA+2Rv+CQWQYYIcFdVO9cfrXVUkrZw+V0lPpmhXziDQp58bR02pyRtWN9E662UdS
QjN/8oAJYAIsFbgHiiYQTnuOC1zZt+P5JSmXUDIc5ukXiryFX6AiaLI/CUucNoni
0n+lQpwNWempFD+TcW3/QVNwJnnM4iRtuCN7FmNCAG8z3msAIGYNbSAuAb6f+JSr
YV6gC1dm8Tuc5Nd+L6rb1lvChxQq0U6xcRtQz/U9//zdnn/FL+232ATeHN2nETPO
PuCH6LIUgQcm87lepbCj9uUV3W6ICtFkqsoEdNAq4Bmwza/qo7pe6/tT5Ucxps0b
xz0XhBX4KfqVsb/S1h3Nkvi9sxf0Bhvg8OUPPyI8BFlgMuoBNGPaA0FO/W3QISxR
hurBW36Kt7L8cxNrBaCLcYuoV99jw+WrPEoYyuCQ9Ya+P+wBohrsGO9q8dFXRi2c
flDsQFJ+78NBu2bt8CQUoYn7PNdS31KUI8LhH/8dV8pAHxcg4WrBW4leaUYdflrp
daEnbaet5di8ihIvYSPOTHtE8/unnQg2caFng0qW1kV8txnPzrf56X6eAcXnsDAt
9C5Fe3nmt8UD4mRBIm2MRMh27wYdKpL4EgDnye7dpI97KEGKDrZwqM6XFIjHq3yu
OPPej4H93/nJJ1uf8Vv5in7z/rTs2k1NOLAoEvLWe+XYKxaZigwX9VcsbTK/cZqt
yKBQNnofS6/5U+oq2+gHgUKPtxfGWK14Jtbw7Kfevqv2pL9RrpvlAOVGBO77sfah
yiMNz+xPVKbTmaCn1FqSdU7FZW7js/BCOGlIv/p0aKPJWBMuJlGS3b7MgR2YXOcE
2KsjynR7e4kG4OY4slt5gBx3zBcxqEkf2BdJ3YRjv6EzGQnlK8BpKGZdgOHnfZFn
/thJgH/qLSopg6SlbktOAWSQRDqgud+EJ5Nb3fFZPH9OSJTtHFSmJyLZ2zfs5EIm
9BN2W7OaJtc5b+LxEAxhpKjcSyz1Du7L86LpzhwYC14Qf+brRmpfwuDRTCh/Q5ll
5pND+kFepw+22zWCbjK7P8nG4yuLBaWS6AyTX0ZLK8YSTJMLbYzGrK376U7JBOqs
IIyzmQwzTQ1GnsPsT1oQJoMvn67ksNubLvDC24ZShLp5dQyZGZLHqMu3Y5MMKRxK
v+cbyG8CEDD+cW8qUKOQ83INMbxGeUuUWedDNooRoIB+3/9KY+/tSNkrErAyviL1
/cUyiuY7I9bXzNHFptgNA/WfX9V6MYfKVYTNdoijRuqIV6iuHEQATsuEGGx2FjRk
WhGc0dWZmOHY/cE/m/HnDTNk3ig8R954QjdGObhsn4VVZD5ZEUT32fKMIpzLjy9Z
gvy5mmmiwRHq4GpQV244M2vrzO2996ZnZk4RyVxzx4C86oqZ6JFaBZJP27B8c2Sz
RMdzJ4vNQPYiFwhQeHoDtC5unRvlQt4XYOzfq8Vjhx3RasBzvcOEQ3I8W64UlDgO
qzLlzURVKos5Et2c6OIIKGGd14kAEAXuIEI/o1SYuC0hPyTUcFGMTa2TF/qgPAj8
KkJ4ZyhGvYxaLbx1AbKekFZForL3MryzWs7HWLcR4A+mmT+O53+5x0W+/1Jiwa+1
uJdnfnc3TgYcReGJNAPHK2zYFrvKvabUlk7bnejAhdoGvelCoL0/oNDW7vxuBMc1
2wCA52v2N4UX1qaz1QFCLbEVMpZ3HvDIPeWhRfgrjNuujPxw8NkK1ZbsOiYRKv/h
QonCzefZVCoer7J54qA98b9RSnbj5OSp8EHvgW3EVoU8wdd8bXNkzKo1HTYkokOm
fvlJ5jsI/hDpRFaK+Hv+Jawint/FYcF6zfT27VolsVHuquDxA6Af5D8UhlNLy8KC
3ffN0QN2TM0u9oNHRifpGW+gne1G2NgTsYzQe9nRKxiuO41SvzJ2BWKLaZbjtug/
TchmTMs7ql18avKRfjJKD1OUJUFCFvAY3eraOG9ccMtwuFEdiClQNPXpijtjzgzF
TjMe4HRVJtEyGwUjcIdTHlcH8lM19yoGSdsIiNAJvrlPVTherkC396Axhemwjphn
L3k9alDB+iVph4Ry9DlbBVUX6SlCAK13fI3GazLogtNKrFIJcVcrn4rWpsVPsxGH
KsXhsmlPpYJ4vn35WyBD3bUpGbWcfIhicqKcJOvhCZt2NjvHfBP+zyoV5iUVPOIo
TtsBTxrrjWoh6REtWkmpX3nAIylbUf0aNdAB5+v6uBf7yKVQ6SCbjk3MvjMGw8X8
ezFkjuGtJ++n4uopu2pVETRQUUYocmKZeyowVAyVrCVoJNJKqd+ODegeGZ45aB5b
GWEwK4jTm7V7TDqNco9OHmJ018tnXyXhjC8UzNzSPPZZLMw5kH3wK6MMXVcDne4d
CBwl0StAbPl8F+4vq6UCOvv2h3uhXxRN5++kEcOGlIwXT0nn01f3MEcsfbAYwn4E
sswW+yveExWd6/vmYJiTFAky7k9eWDXKO1J4xlvNuRkPT+fI7Xy3uBxeQZi9VAYn
qJcRD+yQbYWhW4JsFiZO6THauTQ3SlKBggZtntFL4EsgH+yhgibg+2Ld4RGtoWmQ
ZfE7G6T/kIy/8kktosD+YnBP/FBBarOe43AaEJ/OIGlxeOkv9QmePCZqlwxqALmm
dr0AOxJ72uBaVVy35iN7i6xt6m5nuSnVZX0eb620Oy0XfnCeX/kVLZKggaCNTgFV
D2rnrzTUgMB52DZx7qQLMXMtbKaf2dlXZH0BDJVmRe6dNAYIB6QP7qDqRNoYbhoh
vWIMh6UP0YwPfco+xRnpYQxUdsOHqsiuKlkITkjcCsEJ2q27hGW6qN2qOYoTG82U
XEvLNMiaQ6atu9DXIrdtPq28ZB4/H4OdfAsnKFNdaliOOr0v3QczMqR5LoG4GQcR
X+Eb9nr4dQh/zAfbhpGFtBx0zBsaBfAWWcsTzctIeakYlB1QqBsqAHCNqL45yU1k
/lcVUW4iZARLGxSAPW8l+Y1fwlDGYXikGt2ghP3qmjyknyKLAxVT+8XobP8rGzND
VMnvGXrVkssbGNCnIXpY3+8uH9Udj6XbXOTCq0RLsSt8Hpg0UFWhwz6tLaQznqj2
oEUkv58e6leY3NkWLKRwk688FW3fwS7sAfmJyPP1kM1DlTX90uZ4VBiWgsO2owoT
iJ/3Vd00+Hx/oVlG/QCNopuVwFG96LZlAauHOq9Jf8uM3FYBiffnJZwc8IFd56vH
wLUgycAI/VZSnKF1O19MyYkDRwUZMBeg9YxKewj+xJRte6CYjSd1f0NiY+OJ163f
DsMk5wWlUd/s7GcX+l2W58ujbBEFzXttYvO3nmoXgbkm3lfFoKqnRHcVRf4PNBnE
TkyqRKHh8RR/xEh5zi1TM76MU+aXUG/wsWGMBkgDITp7S4okxnoEE3AjTGd88+z1
sKpmIFSS0ofTYzk8V/5p3zpy6fhd9NQK3/pq1hR+ZQrA8LHyektq4x+dLbSgqQE7
+7PO6hUT0XhOKNxBp67u3gWp0dXh2o6PogXjfLWtizDBl5IsaTb9AWIi1BBdIGRy
QLS8frhLV1jVLZo/zZq034KsMRcEV/NHQfR3N/uQBTgAiNYJtGfDZK7Tq4KQxQzg
XHjn+q2RnsYE4HUDaMMS0f8QULCCd+ksS3J6cvmhDZ/FkpL7p1tKPPNXlqhb90NQ
rJ3sNZHlFI9AjDxo2x+1T0KoLG9SQnvooWt0yVb0lQHyZaicHPJjhzody1ZnZfwf
gZzB658ABsEj9YQj1uZIvIds4hXvPjAM0v4GA6dTdwFF1EGQl72uCZCc9TyVVs3w
mFvD+FavOlczBtIkWxNlmHzid8P4C+ih3oicoLVPKCLKwqpDuFHlgIA93lmCAHkm
RNwJNwXRb+uzOy8GK2cp0ZflPnIKpEQUpSq2LQrn3v/KwFbKnRggyHMmW+9wKUgH
7wCKDlttX147ww5DW/kXL7zXvDXBEg+RctLroMPce+Vi6PR/AzTDuk+J0B9LmwJ+
09AqPDHgT99jCOg2lwzSMfrK5sztAPs52omR5wIJ9TNVjI9Dj5+gEpNb8jcRmQkn
vsqpW/hHf1SUzOBoPlk3veAtv3DSsoQYMvQr86ZUsoreIOHTmfG1cqcaK3rzvHAc
BU8Fg4i63r1HeLnGUJz0Vdl+0e3+7gmg+zldyPSR7soYX8dlG+1gT5XSkYkOHMPl
1OXrafgfFmhAzSaJF6HmuFk1KBecq+f2hShBAKC2GEKnqg76dcucqSH0y5yhwV7f
SCqd0PL7EJ+lZidpeETm6tJnwiLLjmaPQuA6RL7shoO1bXI2K+CoPjHEUiE50scy
utIJEcViPjFaRi0fqNwyYybQpY12pK4yn/YpIq23KlZHbmFVVWwZcy6LiDSQ/Azl
1eRMnB0xGNxMG9uQhreArCztme7P5YYkSIPnoxwDfKDd6x9vKpBH4UzCRVo5suyM
8VcGTSSKHYMIBOCcewx1vgcmfIAAmfqzhsHIVx5jwCzfIS18M5IUmQxNvpjvJQrZ
/eTGIEvuqq4ZIqvHQ3wgG34Yjcz7i8N8aEFsskrqul1lP0ggrJCjSkiJtdmA2O5n
UZIc/NAvC8a/cgTfHw3EGLL+cd6dWQ7wE4OV5U53j5mApLMkZenGEXNX/GskoTpt
7TWyKdYYqY6GBBwWXnDeVaGknfFCKfuLR7brwxb5jjhqyzJSjuU0SDQorLMlYRTT
FFhqzZ6geiRMus43cv1EH/lO5fz6lyLba2cj58BJQxJRg4aGIjKutiWYreu2PfLm
+p3l6pIIbfwrH0oENr9Jex1V/RBFhFQYnn58ZLOQxC6yZa/qVqXPGTqtPp2OToMI
yDY8jtXfDaFFawEEyhRdzXBxmMpHKDaEwVvgfoBE3ejtO1d+w51DEtqdm1lf82FH
/2iCdebtigsYWrGI35FtghPFDmCP3ZxeOv+nAMH7rK/O3QwoNPLMldWqYAWBJlLD
BHcpKQWQ/27e7RbRxtuyFIYZCVPyEsrQSdDINKy6WwxSw73XPq8Rakc+f/ZKwEZR
VwVyzRm4NTCNNo8UgB92o7kkU9efRPr3sDObzc9USdacCUPv4108QlI7C1vVVhER
C/Y7scBiA7ZR62+dyGq8jc4eoV5xICSQYngVftsra771LvRxhs4rtl9wOJOPcYk6
oiB7+0Qz+ANYzfVqCp1X4ByP1rWaTUPTHXJaKgf/LN4ytiYEI75A1uige75vlqXg
gz2/DZ+XwAjVrb6LmEloG+5qmdgUUpBb8pFWzvckBPWcUg+3FxbmAlGB5UAIcqLz
wW5sU7PkYUNz4DdbeMIPnTFHf0+VWyRKaCh0KKtSfTgf2Y7SZ+w/tmo7a6oy3ruv
rNFVwgbt+wuw2lMMKQ6ckJsGS9x+ZVAwIJSsMP/pLU7sQmW+Islht56rsEMlySyL
4hs2f9ZETaG3UIrGV/bT3cSacFqocyl0cIbMwhuEYxed3bUhOjPujuedJ1/WjtUO
K1XQfpHQEkRUr076czInDT8rNqRK0cm1Jy12OtTPspYC4vGLjv7wi5xGNbkJWKlb
pJeePQXDh0+PtJyM9K4NO6Lv9EMQ55qVPGBtil4uSdbC8XZBDWcpOlgjFAGwvwdE
1sbCxdDEBCxiT/3t41KbFzJpfG+16C7vbFQXv/RYEYRVcsi4xmo1LU4OXDXmkKk1
sTfbTtKc4xir9uE9zDG7fMIi+bnFjIhXtSc2Z2hGM22mWJFal5bOzOri0GOy1Kat
gZAnbnCdcU6O3Z2ZObLBuJ/iWDnBjCE4nF/4L9Ab3wXX73+FDkGVu1TSCsDAhusM
BAMxJoXwj300Ed+XtWc+rYU5krevKGrzbH2LHLKhYIFUvk8TWFAIduIImAdAhlI2
gRAgVeCXMnH07BsSOy8XWzgzyngo3v9Ob14ynACDJnTvqAy2H1ylNI8iV12QZe/f
F4KOO9UeepCJzFXbJA9tTxD/hyg6TzI62UCc2amyUqSACzxcotHgBRGTTOFZmPoB
jFeF6WZdRxiwpR2uaExNtOUIipyUio1fkk2fIXFM4zX+3hphAcGLV3Ll2Ixd7YSL
w1hia3sLJe/LV/2Tb9Fi1FdhjymnLZXPb9D5u1ck5rYPV3uX/oKnMXBug7nK2MI4
w2qn+I85/m8O+TljGTAMYd0Dp5fdLlkue2+fYfCxI30EWdQdJW2PGey04Iupc08o
cUmvY9lNTrxJVwnRRhUgBltXB9wyACotmk6dMBCyhNeTxn19rpGqwEPr0Z3aayd+
S2IgqGp4c3GprTWHwlK9HkQBvdPtcNOfS04mp2Ca5bSI2qNVBOp+MTACM/LzUs94
x5F4iHmKAx0uZGmdQRFa0Qc0Sew6924wzLRGByfE1ABaJJFIEmJ0fdjDvuhuj/XR
PIFdGXQ65VpX2jt/zMSYFqD4dWox1DoQYQllFCy0W4flqLuWbCwhqON8H9ORNp33
lDYoyeqZcQjlW3XQt1UHrGxKboAP1pmEo3LjcBn7uQyGoMkXmdOj9zNizeHn53m6
qY2WSU+xdwNwfkKLjz+ESJ2OKmwZ38pVY5ZN1tR2JJRccGWbdWf+dyEpiVbjQpYy
VFWIAwMpHHbKJc8hobKMfEx4a1zunntvxje+2Av+pNskI9vHy12Z21qub67Yosu0
uoiMjWUQtXXAV9SqSAPiuSRyxDFT0QeSY4WBTQd3oS692Z2VajQVgfMjCTZISYuf
+Ej3EkYbK+BNrIiDAlWJusjLdNVG9XcE8fzzxyrC+YIXQDVnsGxqjzgg5OgsDASB
qhcSM78dfuqaOSB0SHd67qFdfGl1v4YOWbrOsoW/hiFnhX2lIr2SXFDbt1eDgb1R
ygC8oZC1nkLOpcVFDQLX2TCp1AJ2velt0ifMUIeRGnYtQtdxh62PyiBwCYarViEX
pLO1PpymQOqThEA/rDzFuKr83qqNlLqvGittVBjeqmNthonfHKCJQb6O8zvFBpFz
N+0r6DMgB+emKyTNYl1Ohv/FggHNH0QBzf3ilvkFXFkgdrdfdmLKEDcU7h5kkl3q
zub9WHTMNFd1nrf4jwxUxa+n+vHq07iJKkfoIEelGicKiKiu5opmFqY1ILrNM23G
G9b/ReXkDQ0QSiIVWH6M31CT7Vr3msuaKCN43a3B8l9W6rfrL2JskLnmgdfJ/Cry
vqTsALXsdF73V3aExWJ1aNK8UMRk1ghMrIDYQ4PocfyCjrkLwhRvevpdl+Cfestv
n3kUSvosNKT1MU6ot3cwO5JcEEO2wSv06l+RBUSHf6Q73rurU9cSy3uk3dw8VFRA
jvswfZ5dVozHVABDCm21fwejCRit+TTen0Wbq3usevjy1REt7EcFTvTf0IsOlglc
uP0usrdqFF405X4R2hgM7J4YrUShFDLuih7An0ujiGsWXI4dKvXbv9st1a88x3iF
nxCn4M7RoV1qRYeu9lorSithsy133AN4Rps5cofXrghgZ33EgC6aIQaiA/5mxaiD
bXzH9+AziyQXjHg3t2jMwJkLCOMmPKfL3xERsKExS4kveYb/7zdMYQvf02xgPI3k
/4qR9cZ9cDmpo8Ss7vyxlm5Io71hQQbd7aPvxPCH7GFiUROEAu7KAavjuSTlyHrY
8fouIyo98SMxteTtAPEj7kbTvZsQ4QmF/9sRy7DrwpD3m36TqDqnQdYzEi7WVN6I
eehLOzyjrB4HkDjdUt8x+UCjqrQV1f3yoccJcyoo6udhZSmFoKjokTuJhA8Sl8OE
iMIONEW1NdGrqEigPb2KJ7pBi2tj5dUPMlO5/WGr7q6rxovdZmLsn1qLUBsiBTv8
4sDP0FutmcaeHoUmqeLuOEMoTA1Syu1WLh9ove53cFnloBoXqrmT7NCzTPfjFksA
ZBig93zGYMx6yqh00iXEjgPMIv2zHv+hY4WpBX3GkLDX0xmhzed8ke2Mat6QnXVk
/77h0zfWp/zOzRfefetNHV0w2LTdJyXL+AIZf6Lg3hXpcwEDq2PavKaVOFHfdKU3
OO4lZzBvcljYmRmQz5IqHiGz2k3T6VdOs/NAxaI0gywsSx3/UC9cn7DyakkidA8D
dynPGlmejNH6GL+rGmsBzQP/Dbf0+bnpJ0/1aojUSyWOXX+k2yd8bDJfwd1vuKSt
CU6y3QLRh3GsXYYMNRMeywChmMaId1PGb9c+bVQc9GMNH2HNCoaPSU0KXFyvyZ4U
ALXaYbq0hhKdu2Ca+nwF/OcNba5hTA71bPcXbJMnN6zFA3CQZdVGiCNjRi4DeQfw
Xm6ER/ZNNoy5WLTKBdq/IlAgtzrUTKxqpXWiDx/73zRSGui7cYAZBnbuspgzsE+W
gE2moQzNT9T0sFN5SmHgkA4/AHT6kmdpl7fSQ+0p7D1rXu98FYxxkJ1Y68S7nW/d
CIkNsCKgtrHQyeXIHTB+moLc/BfMwr3/W7LEEbUkdmEP40AwekMAml3SUUebR54X
9fcud9zixTQxKl7qZ1HQCKa+IAYPIxn4xxv4CSXedCreRCvhet9Zxx6s1wRzA25b
SQGCh2UCd5SjcTAqrkFpKWCxAz3v9DHatRlqpjZoLGwly+2QMjLSBEhypQaC0x7/
eg/GO9T9JLDpOLl/5WU5rOze+7YeJY7Ct+iEjXTChNmd/c5gR03JjouBMQbVCIm3
vjeCCamfqu/4WaJWJhb7fi+eX2LnX5lBEnCb+OIstH5dsNPoPmNlEUN6l6oLI3sQ
al9Sru5kH80SQrlz9RuxXj4n7EaCJf1m2pk/1hTlop+nNKd0lbB1c5koXOpO+XTb
EvsbeG2hanDvDtVISmX8lnelZGEUdhhlmnnkIYhxXeq0Pxs2rTbRcoylPk5YDB83
kyLfYT/6k7gy07sPYSxUxg5XIhbVppQ/eRJjZK9GycHD8XN8R1Jx0bC9kekb5abQ
UKYSldhCdB5rAmzKylLChIrelDgML/6J2cARnnnUHsRRRF6jAVhEdTyVtcfD++ha
gYIkM9sVfienxglu24YHk6TlvqlYSgmjZ2ZM8Ru8YR4REAdOcpnQxOKrtLty7im9
D9srfMWb5jMV1jjYid0oZzY2qpzr3A673GZXVEOzLCx5A+rFa8P51lO5PBT2A31B
oeZumyOfhK+XHIvL1muz+TJ7h8++0B+pxZVevnXeeX0discz7UwBXfNbfXBvC/zz
E1Km72fJp7wxbNQUDtaSlb56zq1FgZxJO/m+S9zH614qrPxPsjvexjmJsNaoO6WV
hW5LISTM8I5ZvgxBRvJUj/4a1gCyAR5ji0yd2jBP0Ki5JJOusn+CDyABNMtw1fpw
axGtVo8ueq9+Fqt23+0NI4GZWeGtr0SnMANW2XQvPzwTCtL24WrYYdF8LQZioK5J
c5x0OcwwmAxGBdQN3bKSeYFY7Ec8HU5FfIvy3cff2c+V+E3Je+DWevTAr7ZikpcG
qjKsxgg5mH8P/pVDJ9KkPrHDzBGutZtCYwRg4I3v0ZCSp3EPtdikjJxddE4wccIX
Oe5j8Ax0bE7ZHmPxqkUNKCAfezLU7nReLSsLan8DOtZQlg/0GpnABWKiZbbpBorT
15w6g7/uWV5ej2Wbp4sUJHSo+CUcu07FC+hLaoGyEhvhPVnV4zL19cXliIuGZkNO
Xq+xGYFliZI+e/1BHjAfS099Juz7tFOYCn/IvD/tihOpHAW9EXdSnrz1+By92J2P
OJd1tNXw8cv93IeVimAwvvjb1pORnY8t92e3WmtS/p+MVSafdtvVEgN6WI1o9oQm
PwETr7GW/0sFUbcLHUloatyubTw9ucyODPQY8+u3OJf8HJP0db9ZYCtXToWfNC4p
8hP4T07qPQDaJMq1I5V9ej9vZ+SXkKF0rZ2HzPEfdRmwh/j4YbIdPFtRqxaKKNrI
eXILsX0ZDqa2JxSNUVLhazybK71eaDaFV1EEzM+FLSkWB3Um1quOaOF6VpRLjOGt
I7GuUGnYRaXwIQ1LNiomCx03cNx63SH/QUp+G56wqWaS8mWq1IACvrT3/qXsyqRs
DxgKsXuPknsdpVRu44YxVtP//vRQRENa5mjTHMouApmBi2VNffSREk6mwk33QGPW
HVv+1UJg4rwGOoWYU1dctFd76Jf2HAdS0NdNOk6F8W8TNYk/IMhmr78x3Of37OjI
xT5uFAZLdvavGlnnPJF+cS8Yjnp+L8DQLuDZ29RBtYd054reHtvV6xbLRIwnxx7T
xM/QJ2Eehf99lB5KHu2vanduttHAx3cnkB5ihesI3es9NeW3GxCaAIQv29zjTfiq
GmC8UWXqeySDbl4aZ06DpP/y6hW455lMC3VO8koiEOyL2Jnx4QBOlRUM9EOiQM2c
NiluOSgoR7Hi/DhjFQMFgpi+3gf8Th6sOxQutaJheaIOC4+zWYGvjAtFieOSvQBl
rYwAsOTG2RY+o452+S2ptdfzcpcAjuOfYYpvbSbI2yGNh48z1B5nPGzKYY0F0u48
KF2GSkuoqcJwX+jITtHoglQfSoXu2vE5eJL+l3cg4QFChPKEaZNsznjYWfSQqEcv
6vwjjm3l9Zmjw9rUJ/k7Bvll4uxgQRkHLiocL+RHp2PrgV1+X6Ptj8EzeLjg8kkS
H0+pavhA79ZOjr9I+cyAGMpGV1EoXjxUxZ/bU4LykQicnH0GK/5633QivGdwBUxs
s3p46wQYXLErUSW+2WAzuGipbrufDiADFY9YNCDCPxzyAQc+ALQ+HzPBU8y/Og2j
OcP773yfXL0WOgyJb2e31Km8cArAsZWFHmZj+9i4w+5mQQyZ6PjSLCVqLM1VRqFy
eYmA4Dhp8JdnXFEnA+cgyhyTTN5KjyrT8i7f2NDUvoY2emDh9mXl4Uu2eT7WImPL
WGGVB7Kd01az/8rFzpJzVw2usmSQe/BElHgo2mM7lgSY5WqIB+gElZyuSLV1JLNm
PCLlglultn9/RybCht0nNvY4gq8Ahz4qRqXagggCDOXkENbo1acBxRMeLc4oYGIq
u0o7B/IPleVkYAcGJAmlIrhe4TNkFGXsT5bB/80viImUFH/wL0vmuUhEsGqLGQ4Q
e5XCMfc6HL3hnIw/Ki0ieFxXuvBgE8MqaZOohjbvKH3f42PcWKKawQGrra2PgZvi
pw/OAIZWKYT7WAsl0gZ+/onElx9v64FMyfWMKYEHmG+K3KlpyPIxL+kiiQaE40Uv
L9A7wvecKyYT+1jD00d2ioP7J+9OFrea9N3snDrHSpz+qEgNuiYkJnO8knb6tra8
obdw9lELKBKKnJRWgTf+CL9tw9Pk/zdhq715meQPlc6zBXd3ssC5eIiwWH4fx4H1
96c+mGotzAC/tMm2J1aaX2uk2H8BG2N0OtXUEw7/Fxcqpb68yIlluuh23e4Jng1n
dj6QU2xecsNR06cUixA2x/IDJHodQzfiw1PzWD75qqgat5oIiuAaMWItTZDx7Vpx
uFQXRoifyxk6bVtZTSrrQy8Br0ILJz+KrLHgwJsm+YQ+F5wDijUIuQKSZEgfIKvq
COWtWkgQ/YvE/SleytGdEua6CP7nBF2hK7ahlyy2WuubFcCp9F4qmEfepyGszrPd
vzz3JCC3c5bNPO1A12VCJNgcgWtAA4v7GtEdJnssg5pcBc9hxUWbfxverrAoVUd+
xTG5O7k9qdeqSWrfbv7HwoUug5wAVvQBYGSJ4n6SwQnMMXSD0ShM7mmFdJreKuMa
3AEEbfJvJ4mNAgKrTS0tOLfR4Ly7r1QUDLe5Jp3MnFiMl7MCv2svJ8m1xS+GqT0s
8RU4h8wEH1dT9WfB0T8liBo0MxDsnFvT6p09rlLjKVjP3FRvLsLDbzc235AUWgLD
JirnKuKU84oT0ABn56P6c8UxWNdSyAL+jlNy7ptbd0PKpgw/tKRkCEZpWbB8RV1O
V5AETNlg6VGZkLQpZZ4oW0pCI+4o/dJW+dsFHLFZVltZ/wCBFkxFCFKWFO/szblh
lpdpJXVyuGk4wAusW7YCaF5PtvyYqB92MSwcLt6yP2ZXpKzPnEQr27SHnl9dzDgJ
ewf4GPrXr6nbi5NMmsE+2Bhz5hJCXbGCJxYasx6Qwe97Kk/foAR2QD9j/MAMeF0r
Y2YnD3UYCHVluNur0p+siOxVSLHqVBDPgKPct8ec/o1YTcWKZyykTVy96F0scpBY
asA8HWXqL+GUxNJ0Be9sBJsCnDe4Exc3yVXYUVKgBhBwpWIosI4oDvP00uyX9mbu
5WGrratfbn3+9OmI3L3B6HLq94WJkVe2N8IqHMwotP6jhH+jxPXIpa0prpLS78mg
gvJGXyEgcuvi9mr2Udb3eLkRMzT0jWLBTVfrLJBhTr18hsqgD+z1SabXFSjX0uWX
EWEDM36i7i45Rquea/XfT3sEGJj/KwuuTRXQ8LO19krynqpDGQ+FP4y+yLMuNBTk
9cBVOytPBoQ5uar1+ErNlEIfRvqP3mXasrmugCg5pTkqZ8P2y/XvKwDaSoQRHADv
mgwtLkfRcWaolF1LO8heUBxKuhSprh20kT6jT/jXDQfl9z8sAIWr3sYnvD1wonvx
CZtWd+iLygt6DFG2k2KSE520VK0yD84YXjnDeDseLTikQUl1FHi+hycrYgFQ1W9Z
2drYMdBPNLKU9Dq73vqQKqtSmpP7ufVbvgAZwitldqLR+85e2g/MrhDFLDVBgZVF
0v4kVlNy3VGlaw8nPcgEKpN8TvyeCnhG3z1cihAv1mUUUitR2B5KZRrT4F4B5MBY
PNzbMpwKHZ6ezla3ejcr2Vr3+AExoTSHsA1Po9Wdk1SqVfc6PyjxKPxa2EuY55ys
e7Ye+JB0aF/L9cwpupynl2tBrug/vwDDaQKpWQc+TVzUV/SRJ2u4aJUXtH5jBLwA
RgxrztS9+b7jKb75XERVVIhZxohNmwgQ4QWU3o4Ye37iFhb6QKV1VaiUZxuG01nx
xovR0GsCmm0YI3mF5UkhzQ/tKmfEDFDgGTpf5T/ZNMv6st53G3wW14nUgQ7NkQ0S
dfqhnh7/A38sksSvZDVTCHJRoyHxuxV4yO69IDLu9zthMdEBX23nVy6ugCU4U5sD
JyTUOeG595dOIg8kFxa263bPrYW0IzH3YXyXaHBqLxNV9/MYJSnOBG4f9QKmM7zH
8COfUe6exLnMgyZpzB5igA5RmWo/nLCRp0DxZ+agmNMb53uZw6wAqMMDsloHN+o2
sgO5sgXh8U9bt7YcYUhbLwhhbe4E7UMvaopM47O60Wj4mI3xjDRO08iv8sFueZRs
dExtKvPkSqmY6/YYoRCTLKMS+oFTRRG/xKVf9qKqK96yb7KpfJDvgj1X8gSBl4QK
JbD21Ey9R390SohtZ3t61LrCPlxMriJPTIIzUNBElOthDgT3xcr6sqB8f2A9WL16
kqwy07FQQdirJhAwA15Y0BYt37P3tRMYE7gFwESnKOsFJRbL76riAtK/E2kHHU6r
7Ydlou+tB4ozBgkMmXGOuCCAAlIPvAqcysa21J33NAAWGmTFyigOawkM/bbNAaro
gvuPdiMY/jLFFu05du+o4rBtG99RypF/UJnOoOU3Z3h3YQeDBfVQOR8Vm1pTtKnY
fJoOjUCjHFe6wSmwzdDhZMbmcQSdd85wywS85wGQgdZnPW6Ng4LNNma/BTVQ0vZw
xOrSpOjVEgnZ8b+KqTTJ1Dx+zFxoJt5m/6NP5gIGRcnMHWOVfOrWlP6uqnidxRBX
K/OI2eUQt63n83meYwVYcT/eDx5wFahXYmSkN2ETCLyqAiyxHX8tnZpc+XkYxEvo
vytCCtoqCTERLHcvkhKIznmTjevWfQfIcN+vHUTeEhtUU5YEijz4f0muD3Tla3Mr
o308o/CtYG+JHwsu3mC4ILXJni29inZWgYSZy49EaokSSFC9QbSKSzQwRq3sEKdw
GjWLJlZqpr8OSYC0X7pimV/LAx6Auui1JhxGuGrTnw9knakBzvR4u7qCDa37UFKN
f/y8Mm66YFLPS2qPBlIgtAMSEkCzcvPa7bOTne/I5+N3m0EQ2jyljRRuDchuEyCq
WOhL5wJFyCDUfSY7GxmiWinu1hgO8jp4vCUzk3eD1jRY85o0hiI2MytsFVVOdZ2q
F8cabA1NLikwxhW6z4qqm9kkEdi8W/ypWS6lHfZVFhn6nVD5/FDdjbdJ8cJUFcHX
oPTWalfPfvK4rl2E+aO+ao9SO/xLCMiJGId0+5ff4b1RvO2R/mvsUpxh6H7qYpHU
4FwVKgyghybP9QSIVRW9v36PR6mfd+0HZ3pQOsFQzUhXM5QKGS/VaP9vHhPKOtr8
EnpkcKelJd7QYd2qJFnPxZ7HNlE9sUPb1OTVeWEAdRkZpGlVlOHWJphXrKFLxBZW
jwUeDNspCmko0YjztRVy9c1C23wyOE66gtESKFKXvkhJf0cToz82zyGd3Kt5W/oG
NRZnnqNx2U1IieDoiSrl+2gyHWED+Sujf3caVzMACIbUYbpzOpXHEuuwGotVpClS
Rbgv8Wi3+Po141j2QDfg1CKr5HGZPcQ/PhyoewEYZw3IypW7j/FiKKN7uxgJKJZt
VZI5Lf7foL7vAWtmsbrwrm+6NnTPruVZGlX4u8c1JoPi7qmpfL1xxbbSbCY7wRtv
ucJCtFIhp50HaZu73+JeeqPQ/BQzhlYPVfUdqz4UYz36uL43i4LeDQFlEDM8yMMs
qevee6PxZCCH8PwD2Bq/SZlbdyhd2CW7BeZADpPxYJZll38RjKdadEYPGvEHukbD
n3k01jiG/6fP2Os/5I31k7CkDW2d/WUmUWtx2G81gOyukPseeCyt1AQBja6Jx7Le
RpmVbWsQHK/MG3KxKptoI9TVJovI5L5xaSO8lsNxtUBl2Q9dkq+Mj/ayk3IXuh0b
vV7L9dLiR8Cr+RpFv8P0rlaFC/N55fxmy2nCGrek/40otrYMJtreyT/Pqo07M6Mv
VjN3wJXOKNAKGpkLr8MIWyiFm/JnJYba+n8xoOLJFefiWxuN8UyGdHHNdzUb6D2N
e0ALaO086IMBnFSZd0rp0GlWGGNGiTViUHfYIYx5NzKFk1ri/KDHiFraafMQtkzf
6GMMG6O//3BEJ1UJlihDJUMywx3UDBWx/8shpBHRYYoY0WVTFRRqVKJR5X9NCzyA
893in20i5j3muTkW3SMUEZiidjBHtGbehHI8z5KcN4t9wq8eGm6jY84jMzBlcky2
DByNdNuw4roGyKmiSfAi1YYRHDcmsThcQb8JGQvP/aHZ47uxXgYd7K7e8kPF8kfq
GmJ3W93ajObcdY0J8zeT6dExsi8bmJIZ5537oxP9exP8ZXGyzVkIpkzBp7Xtvgsv
FbQFHbIWwKG7nnQNy85ZA3DPW1WDksHPHlNxaGnHL/fcg8ivPfra4vBGY6bSoqGg
cMOCE0WZTV80yDgkAFG9m6zelD17oQfonYuSRgM2YZ2l7uOSxgm4Qgkj0hiFIWX4
bqpDgnVR6A8e078Bq9KMs8GqnNPre708CvTmoHQO7800w9HktAfUwjhikVKgS5S7
QHmwdjYQhTeo1n8mS2EHrx4beDXyD51YbaxdsLaY5jXgRnqOZhEHcAPn0LXfa5Yc
x3L1YdD/IjYGce0VFFV6if7QUcJo35DkSkqFBdhKocQpLfKvYAKlqSAG5pUUlzT5
78TDXWV1dQzqrAshU/uM53pmAHTpXq42TIRBW+F2r93Cr+UYEFy8r0bNuBdywZaf
t6wVj82HiUDyM5rwHuh+F0uCh2J/LFCwVGFD6PGUzKRNWpGCtXLnPG6Sx2knb1Jo
h1Xhx6Xwy4MVm43JZtNxV2GBVniJ3pj4BjlqqHmoDPk3nbyUzP1HM1TJ8q5oN1Ey
EKfgE/AKmJXDbTDCP1801FLCSNUGDWR79tWJHWHqUoGkRLNSkmHXzQb7pMcR8xOF
JvVHdt5VFyH/qhM1oa0xyQkOorqua2oC4pXd/DTByx8tBoUy4ola1mysal+zjyEI
U22Gz0a+pWIslXZhf9bKIWycDKwFbd5stwi8CFVplHaxgYM67IpzSzqAtVAm0LgX
zEM7ksuxZG2ymfQH1grZ0JvmLFS7fD05RTbfSzupRR4676snvHWgu1OxvdgZfG5i
/6qsw0LzkNxAtfsRzNFh30F4C8u9/WKOvjh7a6H4gxjoqgdOqm8ZpSeynIXG4YJ5
b9D+/7NIuy3lbNFz62CJHAp3CgORe2e4Za1V9zdzP14URC0PNRcUk7VhZx2crOUo
jUMquCbRg3pgn6Ah6SzVF1KfFYFJr+yhNDYqVN5+sLuODkFqMOiQXU7bx6Hccl21
IhYyJ0mUoBGOPU/xEdZb1NvMHf5dtQWS1zA9FvIG0E1cuRyZ9Io0Qo5e4ij/JppX
xvSGa9C9rAXQXfjQazzBD+bipTLaLY96EVgPWv3zHW/RKeCF9KeqAcZc0ilTK6vt
YX4UZe26ldWfn3r7+TcZbEUOMczk47mwf8och0ecSZ7ZHm9c5f2BYPaILPAB/4C4
0lExUHiEsUTxf3BTVPLnVfj1DCjqDTS31fMLKV+r6gu/jWfmRtWL6u6jo9jDCUW8
GpsmkqBQ+xnqqG9MYtqCXBCq2gVTgi/glCZBUNDnor1otc+ZuL3EwveEkMKuZL3A
C94unEbnt4ociRYQ/dwMwivXZSXW0hDXdfJ2riv2Dozfi7KrXooXz8Munjj9wGvs
j/KILdPE4Vm9WaD/zyN9FAv3vC35etin4tZ+EyFFqWcoS5uyEImJOOkp/xANJSrc
Rkh3ix8Zzk/Zkql/X1cJIBbxerapv3TGE8Hz8ssVjCX3AY4yhaMv0e6BuqOp/hX8
/EE75iaUNGz6NXuC5rK1rjzMlSMIUVJ6OpU3ksZdhUW+sW0X+FdhtoFy4CFtdnWh
p8A+OXiLZ4PrYr+Yz/ocXzDkW8xyn0VnkAAW9F0WqIubNLz7M2UzGKEpAmqn841F
VTBsAIgcMa8yuXMQzUBn/CY/BEeAsMmbZUqWLyOExUdL8lbt9nrwsB2Cb0E8+slL
2QXz7HWOCq/v8D1r6f9ToGXxTIP1ACoBNsuE2CVA5kN4QYlz9581a0wH/Vd6JsrT
k6Y4ZzP18gyV3aOOPMBw4ej8AoB4jNrvQOlAY9hE1W6+S5RcBpfAA936qyO5OHJ1
DCbvyWiJY5nYcY5a/SeUaSRuJlnM9xp6P8820rdj7j6oTUEmgvoOUanVcVdbcuOG
JylYn+IdUuLY5auFfIYLdl++vvBK46aeg7E4ZwxWAJcMmCk/Rv1YowFTtbMXAmB0
zIxJSc7D04a3XvaSwKPseiRP8sAB0IpNQxo2CJmTtUwLIyPYqd0+z2Wu33Pw6wDg
5tVqRoEvAG7XILGI7vBMYLgZOM0ukN05mtFj6P7nBGLoy7tvJdASac8dHCJY0ATB
jDOmCX7cGUXvGF0uhqZ2628WxnLpp4nr96CN+aNWqxyoSoo6bJs8vdA/mgZBpad0
knFUfdRA2CHMNheKh55NLHRT9v3mHjQM/b0o90owwytU7ze61Wt4ZBd9HTX5+vTA
IQtXBxsOqDF2hqsE2KPKfpi27c3zfH3ZUIOstvgAd0G24w4PMHmIhyicUxBSW1jn
OiG6wEGZOQtIGHhG1YtXsuwSLX+rU4bWQjn1rWbI5PXHqhplcq7YrGc6q0wDDgmw
lOH7Y6gFNnq4G1M8Qm5kgWlFEMIIj9UnPg6BycRBRydXlnBN4paK4cqM8sd47psj
nC5j/iCHhvXbxJ0pKTE2VB1QKfQ8OIG+WZvdnyEtalZ4pDXp9Tged15oZ/dxOVbU
qZ7pA+qBQ4fIZSNhTeOwrV0+o3yMUKLw0nUW9RskkW+fD6hWFStC+t53X3Zh0Uyn
cafegp03vmT0GD11kIsIP1Zr/LHPMubNm0n/q0ZrV1sNZdicl1Bs96AlKOP3Xv8A
D/MiljHbq3pDlMckp1pjR1hGF+2drdIWBG+EkoubY073TvsTzKvhFOMNtz5IgyAo
2PRTrpj4KrcB2/B0qp3bB7ErXC3UD8rJfuKjdnUVPr8nOFKKr7/B002MBZIzNQpW
kOAwJDKqHUklAsEwoj1uWxQvKqiDBeZxHfGQjZnwfs3YQzqB+V0v0FabIAqsMzYU
OoXdr5PQ+EwPyxsMi5GDCCz3vJiDTuFPKhMUrvz/t89LQOKyIMS1hY20w6YfS7JP
VgUwvDO/H4eNYSa8XGXBotsOTuQB7vBN/pj9jPT9sVdwE28hXuxwJFigTlE7owo/
3hAmK58MdXlb7k7xZJ3uDodtyIEgCUYGWl/1tCNmH2oyurtUWTOsRDXdN4radmP4
9qy2KcGajSSpSQEqUG5imz9IThmTkGsmq01daTVqIUEyuwVqMJv1NLOB8ga5I9G9
OcnyGkQY41CmecGk6OzU743hKOr/O6slnlOu8GYUYrlyDvYma+a3UD6WFtLbpAIA
ZaXGHSAyRQUvP4PEhai+e6dkwaOKtsfn/yfw62v6a11MUYnupqrqPKIN6DsQWVXH
lst4wlKNFh1rrvItx5CX3TaEzirbcdt/Glev132gKfDoYDfqQ3Znxfc8DyZRGuEd
fmEwEslRG3EmLQo+yYGOujAOkMQ4EFn+zJf6+tW8I+YMzm8+bu5RpppdLwqIo3mw
yDEEDsylk9TKsO2CiUql9qkmvjBubas5sUANVbBTTijrtqVSFpRR9CPR47FG9x7n
D+BSN4++4gpK+F+kL9LT4XE+fa46yz82zQ5eZAh5B9nIU3XneEtkf/fMczlYxYI/
ee5tG7jkdE8yRTCDVaj5dXmGruB7B8LYo6xM7QTqG//ZQN6mkhS5oztplUWKZaFO
9xQeFzf7vhx7eqUmxq+IX+4l2fIULXr6ELR6CSovBkdO7ZC8yAgE/LlTaH5xyElL
PsXHwc1mCi6B4AYo/+6BNgzX1u9CSGORK/etgwL3nHIhXKUkKRyijrGi4WCckfym
8eFU9DmTcYeqiEa/Z28uC1oT9vmS16jOGG9THUjgoqgXNvPBj8bXSBX5PprsXrpU
aUHESz1O4rPMaUnKuhCw6aqaSOEoWbHWsfhQE/VhKu1nmh+b8FUy2pyEFz0K08qs
7QOIY9p0JDbezEykzZmpHbVRr0Uscr92lxTTQ1T1yHrbNhKbuX3xLfnkkagIseEd
V9En7MqT8Mv+Wh37xFUfTDoOHP62z7PngOOhUxgRbWS9SjsVgwe7Odz/QU0Gapdx
G6oGG9dzN0PAWqnqrEnVX8YFylTzlDl9x8RdUqwwzfuNV6eCmApuw/Uk0CsjzhF4
3hR8pqn8Woz2jBhOYsSV4KL2h95/yVZHtxDmKJHJOZifliRpmT7hKPDnK78NouxM
6LCEXn4ghUCJOBenvr9JPkp4TOxSJ3VIF79NaGUXmuTJVNHTd8DY3naZ4ZCZG3P1
+S2c8dWU0okIx5jd8+f2Fn2o5h6eKGB8jfjlhuubZuKawqcFRDEZCTAHVjUW/KKX
mDe6W+zNPRN3a0KeUi8utCFjKIXUSdjzUMwiwVSc17lruxI3SRUcizoTgKtbUB0s
R2xZKR8r0i7SnwmEZUjVdwR5ed3EkMqsM6VOxLAC2zwfjDue9y5Vv2dAOe0DyfKM
bBBdMjj2M2qHMomN1Yvu+aeXVKkxrzxVKCsdpuYwhTfp8Ai3QLasOpY210NiqM4e
EefPvHaYHlywWctStLNtRqnMhSkh5mkZsIpxhIuA+JFEROIHaeNPo9tQb2LgE3Ad
5aP6WSp8gMLVMhu2+EOVzRmXVi7vinB1d9Dzr7LF02mcFs4jShKgf0flGTszXHYU
tCsExUXqnsSbDGGV7Jyah1wBp6OWkr5K5xEnWtN8l5B7ohNFvY85AWarQ8d9x4Fk
9YNSTVsnM7ylScmSFSxc/4zLgVmhGhpomiv+zFLi9rX2MA4dzEEaWO8dPj2Esx/y
X5hNv80ZpMUE3O4QKlUiE00vHDIJHZK0RK6DcRRGr1kHWS3y9UysnxUAWNy+oaY2
1tLMnsPQVy1nr7cwKM0LWzKt9LUTxAAkUuNAR6S45jtzqCLs/GSIcOspMSuxOsir
eR9C28xdVl2hrvDzak6u3cO3QaqcVUP4gofWZYW2qjpLWAXaoKqQYde6L20AupOg
UEHqANcAYKwnpKhQVgcKC+hikaBZNQ2nX9zCUG1FTRFsREeyHtLfFNP6ax0BZO3k
257u3ycwUl128aDukioznZz4JHb4nv1B38l008Hy0gFj/ZGpaeO6g8A+yZmrV1J4
RyJsNQ9XvsG1WnsFWvaie5WYfjHK3j47WciNaykS/ivN14UIZaBMPNxv8jAu2QoX
lKwiM/pYyng6WkalrWr1GT0nFVyIku66dSugxia1CTJ9bL22lrcZajnKuGaCYGWU
IUuxQBCXmFuJLzNqvhRTfMjVDH8OBkDZwtQmwyC1YQVnuJeAB5eTuifUPGVP4L8H
IYyzoJhwSgRY78yfR5ejV0H6+QzOv+vMFNkEjoaFLx0C9tLE5btqwgOtu8fTbL1H
2xWY7gTQNuAHCiVs71eu3RcJ00LlgGsWmZgEPsefLTjZYymEbiOr5MvTaGqXKYer
1VvsqvLesdEdDzOC9Z7zyZ5bsvIvViCJMGa2zSlb9dAp8n7WZ7JkpReijtdcxwef
PI6t63rub9IN0mnHPlvrnDyK8PboY5PlIzaUhm577Ludi9A8yAmpYe6PBsCFlnqG
T1U84O6CaFrYlY0nqOBAUnvRvRpoLNVuFUQI8RJtGFk7sc9H6zD0XjBcUNXQDLKR
SkDGnJLw4jzYpWpA5XMuiE7dIoBq5+eFvLnPQPkI0jhHKcSrBuKXPZymikbzKM4p
E6AkG9v1G5sna8iZp7hbz578n7NtdWs6PVBo1162d2Q8/9TZDo3P7cst6tdnT+bW
+L6NTIlvnrMfR2IBrQ5yvcfA4SdpAtnNZzWHjAgMWJ2AmRw1ZFkJ7DjrckgfpGJo
JG330xG+l9m+/ke5NJCT15Hy1Bt0OXjBOIwvs8qVTKy64ajcroIsNeJJN7Sh4Dzr
iSkNHbJ99ypRO3AQM7uxvbQz4ervforiOJliEylegEVhJ8gc5b4kiz7QcUaaN4j1
EFim/jpOQhKL/6X/a3z7S4kOvdXSll0wrg1FRbxmispdEJoOblfzgFweYY4AvbnS
3+hJaVDTXG+6qELW3TwH7G4NcUa1ffvcua8Y1GDT/m8mP5sMONoXPuwgJgIpdT9j
j5O75yrv9IgeGiU8H6H+dEnEAYz93azd2Gc754YgJDfTQFUU1pH3m0DN395cOmut
0WH7L07SIhkpukE3eme2JOeM5mfQUt2+1Nq3JzYwYDBhD/LnAPULy/mOjCrmQU9W
Y0VAqPsecq2GmRHgh3PGEDFGCNHLLPuabn97NcV5nBNf4fmh161xImGJwriifyTH
KRDIR6kgpWvmP+ztSmrmycfAo7I8sy4WywlzuYQHuWvLlkqVGLV28eaGotJfxNuW
ypj6dyPIvhaKBULv/r4c1TfsVqe8Pd9aBXpC789T0illSRXu8CGD8mBL4b62Pu6o
bpA8mb4a/8+UeUsFEYVTXr4BzmiRgbiO2XLqvmU/pn3X4/njaMCMrka7whNJnyvR
g4SNZ3muKpgxIN1WS2O6ngZnrjXBuBZsf+Nxhh2u40eNlKD6tdUpjluXs+xWIGNh
rZv3N8+dhQXoSY8KnKmv9UVFVldW9LV1HCHkL+GzN6JK03DS31nYWkrKWBE7aQ9U
S746uo+ZQPsJLJYXHJtlY7m77aA+T+GS0EKgRlHXAa7KW367GzXowk26ub6Doudv
P3vipPEYRsnUxuujqM7CHbWEswKcr8v/K2v57XU4RLtFvRYwMVBiyObVrGCXyyF9
gSouo7UwCw6CYa/306vQasYuLe/z/d0teWQaqXETmnJ2BBk+Tgbz66ENOhpBVUSE
2wOiRS8OAcF6BfdibczOr/trSQ2ZBYFyaXvDGDM5HnopfRlpYIgpyYY28wsgwbVm
9CbNfjFuqQOKh1bhmTtRAraDFJ5TFDpppREKDd9MbQBWovNU+9lAhmffZ/3iW8j3
1gp+ho4XwZ+MM/fw7tNBXqqGPDvfcn1Spu0ADwm87VYXyWjSwuTigcF9SltMSy/X
jLipJNIhVLHzrPzhEJDtaUJ1TW4aksQYEONlLoV8q0+JPWj5GBVcZ5pmZpaBEElH
A5AdmcFaCaMnIYw9c51QDh3I2jGw2zM+ZyxPCBoF1+WZ3jaxiExsyUj1fg/LZQky
3uQTdL9gnC8aOjurHZ0o+xBTqIqSWiOmsKv3W/b6sRMB3dxlIgnxMPaOHFHhEy2H
9/8DaipA5h68nl3DFMW1m4uxAdyXZ0IHCRkpdEA29esbyEceGoA8agkKds5RUDXX
3KZQ2GUlk1ONPU/D+FUOHw1t2BrqxtUISwU921vXG8UZpsvAsEMOs4hyOeXJC/fd
ukCW5eqxJ18EGvVkInL6Wvjw2c20xsi5ootBv8S73lSQrQYzlanZYYTN3CF8SGei
51lkgwk9AXdf6vto6xMDw3E4pLEyfkusLiV4MjxrUVPSRoeivX9txgV5Vad/9CqB
T9/57anBD2MsmMj9xHJhSb9x/dNO+viOtDcx7rJncHdd7ujwcBYGBuNWEvjIr8M5
b3oDoG+siTPOCIFYHgpPgw1tSH3AaZ/v4oL1+yQq0XFqqdyXb2MXBOQQL3mmSy1I
duK4pEJtjKSnMGoM38Fo3urbX+pHFe4+KDH/Uzi8AheLZTn3h5Dvedha9nI2cPNz
7m5KJovUICj4CR6s9Ps4xcp2Qp+3hAFWyO7N1WlqP16jNcT0l8IRIk9lNofRB3MA
TcwxzWli5Yund9ffsmF893tKxN9f59F4atTyTMqEVnfTvmP1xv+nCGJ5ObLZ8VHi
1XmAevsZScx7+IYXcb+RJ+F9MtiYoLPXyDq1hv/a7j5P97FB4fs/7/iwOXKhewYE
OeVpGzXnWq0SQIK8M27gqsrMsnOX1mJU7y5KoIu79nOEmL1nPVqeM2f2HALA7N8a
+CvNwmQCnSmXdlM2q8F1J4355Z4m62012RQa/Jziu8Wg+GUkb+AXaRq5MnqNMbak
iI4uohd11mQUMyCke7/lLjJ/UyHeb10OG9bhWopiK3ziIPE3kUSdR8ge/dqVDSJA
OjON1FF3I2fFszGLArSJbGyUHf4K0393E+MAA2rE4WZ/1i5AOz6LdvPaX6QM6zfF
8b9kGu6vf4/fj7bssOlDImlTnrw1ZM+e3d+FptNeBZOHP5DGvLY/ugr1QSpf7xx6
ByrMetfieS2uEuCVGADDqBoc+7st0NjJpwbx/KaIu3jzzwfIQ2ul8t3klGYRvoiu
XYUK3ocyYMeDlHN4KkX864SFVPOfEddd5iLx7tj/AqaxTpu1w+HAoGF/ZZjKFF8A
9gItRert4C4uf0FLui9K0iwj9Sqso+fj7CzQNsZA8dHEmgo3d6dfVZGpRZZxqOwa
V42RPWQtJkyZP3F42DqTculXBIkkAV+WZKWPSTxYc2YeW4EAZbFAiLdN/r97S2p/
IJR/TI4Ea4h0Al6VY72NNRV+6nIF9LrBrshIcSGoKiedgka5XbmkB4LBD4D+yGA+
HyiWMZXWFJ6UWSlfnRsRvZeyKXOdriM+RlOsGf1zUO28SgCVsIY0uTcYf3GNUWgL
LNK5GyBbLBf/rg4QvvftuE/nMiJiERSvDHldI+jckI671JKSpPq+bdH+Hrrod6LM
iiu/WK10Wuc/Zokgk3LpjFmrrpGMxOTHzlSd1H4pArDtl73NOiX0tWs83aUDLXQZ
//Dgc1Alf2kSGjYbGXjNT/35r8W96NR7jB+bnFEW4ZF85ierckKfPs+ildG/8Gnp
lnaHzKXun+SB+M2peciIUgu4ZdV4M1ZNZmsG0+3ULTeVnTb5c8v4nK6uaW60FWlm
PwLyxHbLe3LORFCMAnUOkrCZu9YKmQSt3XZ9vehtbH8eKvthOQWYQIOeCmLrDMQt
TH70IQxZFLpDh1frFlhJRZFjpBWFNADMdqng579cNk91QY5HVLVp9axfMeTVBZP0
Eykkarx+7mBVFUhFFSS6TCm5Mqr3guIkFU2Re2y6lEUO9my5sA61y4hGVuM2qArP
JLwou300KzjEqYXZurEXOuxGXuYqgR/nJ8VsErCTC/pfZMa8kPjQiTNbIWuai/on
cnz8zI66QZDkhm6kE9HFemi5H2Clgk5NQX6c250U5fAgbK1k5MJDwDXY9Ziww7sl
YNolA/cRHVwWvjBXpi+UxpygYBtv0Fl1TTMih8jU7EnxmqhP+dUAFu/3VuYydSkw
WK03lq4RyBWtUgHwx9pomkJ1heQ3kbzwG9e1Pqs4oETXc+P/DUR3dgZuLm3CxFNN
2OL0GYkGIeGg5brxDZNx9W/mj/PrifnoBISHpV7eXkelg3cluaAfpzmSf8MfCs+9
qWBjtESCKc4faTzfM/FJsa4ZREZc2FUZUjEfCKVJTWJ6xtMv0HrqkOJli2mWnCnJ
JSK/eDXTDqWDwLHHRFOKH5u6Tf/gP3mrLQxlqqsF3g+w+GwEH4IIt+cCRklQ+n1O
vZDgb5DykZZIlI7/uqWKOC5VqikamtzNgO8n88j1lRpr1lt3erNKFuMzrykJKIoS
/he1JWZgj74me98fEU9YxpL+8Irnm2li9gMc3LZa6W2B0vZFgQNyNZpQcOFbNCuf
sWwafxIPkCPWRw332RbAj77k6gbPzFWr3WEfbvm5BjuAtnST4MB1hDwk88eoCH+q
8u+vHMqo00DU52TzXx6TsVFI5KbT4DooKuVXpef6g+4Vnddugzq63OGHt8W15GpP
VDsH9/0iKRzpMiywFdh1enXm6O3amPDUmHXMqFH9iMkkVM0jalR8Yuw/HVisiqKQ
ZEHmT36iTBqTHGaRwKHuti53THPdzS4MLYkvHY/tAhBxVn9Q7bpkJx4dIB32VChS
tVJSbn/4yvl1hr2AjqA6UmWQKS9q9hzeMHgxP55H4+6CXRnYVN1bP/1+bPIqoRTK
bKYJL/KoEPGgZVfOTwGaLQy87KzUOIhyhadnAGl2ku8tLDUcOYcCt52A4elNqJrB
7AIH0b260c2KL1uFNbO1hwlFCpRzJUWWWkSz1HzABgjXMf35nJSbeIuoH8bEHvX2
39iVfHtL8gihOntLs14OgzBdtHmY6ExzQC9NYaqupWsyRgxhLkT2hGmyxFftBijQ
jucbU1bBeCISZMwa1xIF4ZZXx6VYEuHDYJofxduFAFs0Q54jvTiguV72A8G8zSGM
icY7b8U6ueukZo3ZcqpZhSQh2vcxoa2UheCwHwD/w4XxcGuk27gIzVZZ1lhdtbBc
+MzsqMlA3O5Lcy/o8wWG+p8YQLLssGxH8LIvAph+mgiRIhyw6420Y21mt7lVGV8w
D1et8LmPtVWOBrV2aldjyF4G9LeoJ3aXnPtcFEmomtlGB9uUXrAIO7I2Alt3f/7d
Z6SFQOotsv/dQnIDzvEkb/oQ2MoOIj44B39tKpmQby7ZNBrYZm/Mk3aEUMNCmOkj
HxR9aR4MRLkCt86Z3FOospuw8oPKfcjas+bStQD3hz1v0DHmJT3Z8j3n6vA5OuXs
CcXw9HaI+iV1RUVA5SVt573/dmmI6qV7iaVL+yUWBEjPrUMkZtZtzBs9lRzhe+OH
vUpN5jHMXaI8YgYgf6G9NskbudHtTBhYFZCZBXnY96jNRohP4zO4q3mLP2CBuII9
xTxm/nk3R5Seja+ekkmWaqAiZG5/7w4R5Y3A2O2I5EaZnbwYR/V/oRGxU7R8uMbj
dGZU0io1F8lf+TUBUYyCB2hg2pInSSATJEB2UbNGj5PTt0exZJ68fWBefdI9FcqS
+yNxZXz5CB0opmi5ZKlKxJEHLoKtkNxTdmXIpk6KRQULlMvBJrS1b4Ae6T7enrAY
p153wConm8m/ZOnaiPzy63BbebiFHn0SPwgq0Aa/yRQdSRHOu80hRwpxOn4L+ofN
39TJeawEgqzn7toY5d06lCXQSN5MJO4PyGz2565fwgOcgNFh/FTsndSd5N3SbMuX
5SpNqzzV12haWvt2ZXglF46PSGqObk7ZaE5XDJOZ6OcZGY9v8Xi/VQ0HfrMD16HC
CuUQDAAYUgz9DAB3WTVaTcIHiP1b4uF7f2kY0aDulGLGHIcz5fNn1pyR6jRmsgX2
UGdIhORHIMlfFyvyCfBsf0AbO0xBPRSZ+i+obR385pF7uSmKnmGQVpjgtLFnX9Oo
sbYaqBm4K3N72xGz6pqFMVhJqKwuSn9HMPiLvTu1RuTUBcUyTOU23tV88bgd1Spm
7oFyhMRi4GMMA5/sKu/XtaMglsVKMtZ+1CDCWktLB4VgM937/6nUglxyMRa+eDQL
BwTIa4hoOGfqOD4Ehd9wI8D93giqqWELps8tso7LzXmu8VnVnHvrCyAyjqtUIK5s
hLS9+mW2F1S+hyxKyuMY67t1DEmn3PRETohcPSBV3mPYlpObtmh3emgYVV6bCUKr
XWGSHUB5zu/Xbh2QO69kg88TfRkGWM3eJnKffr9p61psP4fSO9azM2rg85aV44+i
+QwA7MsWbvgx2o/runmY2NW7oyyyb6EhICspbErd7e0tNVuOIK9Sb211I4Bag8hS
6ieriW059RoNIRDNPgkx80AFoOku13NtBri0ZiTFuMzcXff91WqoCZRD/+n8H7XM
n7VllEqLaGIiu7oSsvF2s6zKFr5LkB0GDCZMRCPefMfiPOVvT2tVZSHe/AWTmvXy
2EWyV/9que0uNJzr0oa2zTNiBdlzE4ZkFokI+H/nsFd+lEA8xKlVH7/6QoPFhdPe
2kOnIpUuBesviiBNTcO0sh3A0KpRqymzlfgvco/LBY6QL0BlTQlkhADQT01YCJQH
6dXnEb0g+Oz7s46nzCstrmz5uu69DlUCL4kBEgAPzFopsb0sMvLxyAI6uWkw2rTK
BUsAEKG1AhCk0FEvwf+qupIqJ0bOqibvVCTSUKPE5aFvFTOJRnONunkyGG4/7Tj8
haXMO/rHoJBqM9BWtWVzM6bsAstCj78axnEHnIY3eUnljQx+x0Vd7iRSK1VBoppy
WPs+5pbY5smqSMa9H0qKw1ZBmRNRj3Ygqrb/Po8NmRXrZxcEC7GQxa0XKC/fHKL+
lGhgjAaG1I9FVc29uM0v9hEcnFTwVSlmKkeLLoI0D1/J47N+IEYP1CWJtq37WnK+
eMZzG+XF5GCZ++ZlbUo8Atk8mkTFl3mMj4RPAZK9QfFvEIcAQzb+iU8JfZ4ap/xT
rJp/KZlWQq/lebIo51slnOgocSSzF/qgSO/7vDuWbp8xqajxEcOtAO6qWXCwcAug
JCqMPnOPf4LOXr/VuXqA67rK+A61STgyIRO6l6UptX8aUTjwfXjwZk37hgC9h9Ds
mIXqwoRVVCPrOajSUbaULSwDpqDimfOKfoBAjfZaloA01Uugf9AfvVeln1yXj7Kv
xkKCr8jdbBRybcrb1tcdy435HlGWo/0PNP0PUClLy5IPT+iOObt3NEHB7N6R8Uio
AkT9MO2UgD5eGDsGY/3nLUkjmj2fidfOuvzLoC4l9lM11oUsN6znbBiEzEOUICVH
x63IzNLnCZLinVjuy8Ba4hkAzwDgjv+mfIox78WunO0wjEnderD8oxEnH3L2pLYN
eJdao32M7gehI8XwJCrUGwn74EXnKmwqgCZ4maFIQsuJEAQr/GGPtVnev43ZyFp9
jgaiQ5bAvB9xO05TmfJGfFfLgvek5yuaKnPqtzzMUiS/f7WiGDEgufE/kUNRP8i/
CHXvrEOLSfI65W7FjleidrplrTQ6Yf6KvhrXFmsHs8os7Jm/SCxn+/H1sJqQMKbs
Otx7U0Jz510DiCNbwHLKTc9JgqO2dmsY1prNn3Noe3obylZ271pDsivZR6GIIVfb
EDigE564vgeG4W2WyHH5j+YbqIjtQbPPhIhdPc5/9LidpPXZ9IxNsI1AJKToetoX
aK6C6X0wJOcLJSMovgNtshluZRI43KculG3p0TXzwsDUFqvLC+JCk7Sn+vMNHNC1
rJQhwMZ7r4pmZ7hg+bIuSI7dWZmknkA1hsvF8rlGbrwGGAHzGz+Qt0hSsbPc3UvR
UqJsd089wexkhQh6bPDH0zcOibQZjVfgzqSWlfdHnOI5UJzGl/zlpl8xOdUn7cYi
CWbT9G7EDKW3Oy+PzCgWnKuJ1/X1YsLvG0R88htbAYK1AecaR4E2td5df5hOD1b7
ncQP4KqKT6G0rIM1IJXxKMgP2Lx4pStZY1Pkcq9bWOcyS5JplDwPZgGEVVlwIWrC
Ztumx1lz9BAd9gEDcWaRYbuZBIbPo3qHlrVByDHYelvitcnpYhWHf1QTpXtZ3r06
jSwEhv7lmkNJOrFjNcsrizmbbajEmB5bz5+0JnIIlBYfLKEeHYvqb2I4CpJSuXhp
nMHqX/VuIEJGEv70y308VvgbtHk9PkWsXmcifbSZpoEg1XETlYNhiTDJRPoBrBvW
GZP1o+H4vGa9lQjPz2MTSP57iKz+KPuaQ70pgefeX9RXiLFtHM+AR3mF/Kvuia4g
DMhim4VDxL7BPki+um852wPiCnQGoiZ62pvs5VpNngmic2tAfedsw9lVXs+YC4He
4lJVtomn55oRppvoz0ii+YonOeWxEqyo43ek6oc7M8FeDmYJfJ3u6U5HNQdij5ZL
9DXbhK4FexP9TQZhPDpOFDm+D3TPrUw0qzXKRaZCR1XQhWmBdATpV/DbhGL98Zpy
BvlGYaqWL3nEsKzF8jqpmqxqQAeZIv0AjfPnwWSv2NX7JDzOYMBrab29WCCYxkfU
i5hVq2OE4Rwh8Syb19q6rEMusF6Ymrtt1KA9yTPK+vF4Z6+o9z4X549gakG+DUQv
rcoGa5WGlAWFOB5VFArbpYSZAx7WBN/ZG5ZYEVYlvkRsZOX0EpIYrNF25VcWcWnY
nP048tNvO/jhowmvTQaGnTq7RLvwD1rfW7uwxnk0txac4KPlh3yyvL/OyEdoNc3x
lNY17Io5aGCAW871SkB4ACEdoluGYYUL+3Z8MWAGSbSxS+ngCEmpcjVcM495HtwT
b2mE7lDSxpJTBTp1w9z2svzDmlKjM5gW7sKhswDdSef6aYtVD1H8TlbUGCxFSAlz
VgqY+7rjqMTr+VJUmtC+dAPRRcgAUTh+I+S5yHU5xAfBzFqdmNAPmtioGbCQestt
lSaPbo2kF/YljJ5J7HaFP/y0JfGKrS+f3BI+2N+8WdjZMkCOxMBcZZl1sFsWWrtK
oPJxXRVZQhK11KvgjLIUnkzoLSLwktQq0xdX82vppAJQtyiYZN7xrOwdzZe4XIU4
djBgZ892pNashX+LZMBGZMrVAiT25b8vnkIi22LH4NjHjNHogk4eZpx5DiFFZH3S
mP0ZAXici8rVWvp4pihD7Ycl7WWaT7vBIfR78ttNcF/EPtitgVHa8UbbJ/m836vp
Ig/YerewkHhDZsdeA6Jh1F2YBLsrtj1sAcajIuELbVrXlTnFzb0YuaAmESaBAKxQ
SGICHY8Nhz3Rlk30TgOWY3sYAVSRGg2E3lAya1u5gu9rOSLS+luy5colvl55v37q
FpfM33398nrbqb3FtzNXMMXCCAd0wsuWjEP8WQ16aROWzvJryWKah90/tWQXGa8b
b25RLmazlwTl8dYE44RryMgO6jID/8IjwWd6mHwoO3M3INq+BPjrHAMIQwSKg7qm
LFqdoW9UQhrNR0U8B+Mog3/9x6rojZhX/wLcTJXNRsv5mmn3EN2gqKnmbFrkOk/Q
Z+j5fk91akJUCnkWbX9fBYInZnoJ7iz8yRWcUnqfKR3ipN0TTBQTqxYDOgRwMs3L
TvePrndGKGw35UVI1VQOlvmO/Eb9C+kkcS3mtP7dl+7n0ywgjyICfjCBZAEXYHVx
mmVgR+uyZwkru4g0sC3e09KWYWGy83tX/EKohKNQGE5qjUoNbtVUaofilsScXEdG
EM+xjFpYrJWU4hsSV1U+TnluN6Bujl2Z5Xnjh1fu04pAoRNsm4cBwcdCjtJd/3XN
jp4ELLGBIZSMut+L2dGHqGSNggZiKmz4Afn0b8komeSGnAPiW9t5VWsmqqJbnxe4
zQSPP2QYZF7kcQ4JqYgIy6dieWPp+ZRodYo1IvsgAtg5MI1+6ift9+hWXRjhWIt3
6HB/d1YVROzos2P+Ocg6/jOzISQLR6AdMlPMTXKQSloTptLH4SqfRIKkPXz/C2Pc
kxNLRmvOKqrZq3fHFZXxk5uNWogagV+wTnUOnnoSYgNXw8tPCI6zeWk12+Lu+Zmd
ImYkZm8dP7bwR6XpIDd6JSTc99mdn/PtERbYF2b2TE0FulINzJcvOHDl6DBb9mq3
Po3W5AAI/6qXO+RO7UcWqeW2q7A9Q9IN+ZMclD2XFWG6Sk2G+buTIgTzEM3lv+DU
uPp66ZkU2Fn+T9ocHWvGoBceaqSQtMshU0hgMhEYCXINijeEPt4fB0YDg3s/jiEz
KQGI8mJikBWSKElFJUspRSGY43n5viOAJP7Mo4nQCHtoTdR1OHn6zvtTpPqhVyXw
04EHJ6cXdAtmJEFGwN/DgAqFR1XpCckn5QriPgZnPYSRkKbT5lwtyUnLpiasYp1Z
V9GoY21jYqilH7HmN0cXUS8FAIkNzPq8MV7TpneXQ6udjduf69NzEP7Q6u7gkXXc
gSzD/WLB1nOnfqQCHIPKN45pR77JvKo61E0VdJ7oxUlnjcM5OatwSAjzA6JPg8sd
yCnp5NRMTo9xc702La0cjpc3gVhX8jUd4Ac9FLWoyQWgQZ8gqE71/aHNHLcL4YLT
JZgq7UVNsssgA+QzVVGXIjl1p44hGCNAaiQphtFcJjFsptDfbMGOdgTbvWBXgMd3
Rttx+s4nacVZF18Q7RXe5ciEibfaTgdH2fQUhGmGe05rBDRRdsFw2XGLlU/t7ZTQ
rAh/L4uI+dQmY+rguS/PJfB9LwcFcXVMXcepl7R9EUHMHhHSuHYSTUwDjcBIHSVY
wrlYNr0LolwXSmDQzAuNcmlJp3qyilZ/kkMPOe6ndj1rM0WcAVruMDHSlfUnKU7x
Iq7iHfS8WcRM6kQ18EhNRnexvebenmtPvchXgqOgdwLXkCAIkyVyKTXOU08bzQrn
cIO+Z6oQAjjYeSaZvcap7WoY8E64jio+zpmZT8xtBYd+757upZSnkWKzawjN2mTJ
1TN+MuddI5frIBaasTFvOnqLLfoZ6NdQLbvpm/iSj4WrLdYS45s70bG48ApBZd/w
Unqnk0GiiOek1LfLftdReA7irywU6Kh9bs4Nx54yYDcGuN0X9zDP/N1BkroZtxsS
TmvPCInO1m7nAOIFP9LSUslUQ4GgsHaDrEt7q+fY8OmwG7jJzMDqnsZ52Z065Qn6
OnPyfhXNRzATdRuopgCTF/f4OVnB6jg2T0mursrAMuWU+3lLO9wwpK6R3WAy+WQW
pC215rVs66uVFum/JLh8PdGKvGC9lNwfsLPh5JzF2cAfyU/IfEzmCLlAEUF45ZkC
47JTgu5jq+e6xHyQVKYOCtoGd1nVh082t3rs0CcI7+beudPV7B2LBEcfcxLrdCVx
YU/EXsFH6N5XDd+RaBMCcNDq3MmI79O8kMVNAbfdyqP6DZAzYwFObw8TeQzTbaNB
FG16xJ+1uDtfVmL3hQ5IyMcPzGHPkYs/Q9GmNo1HD2kpiNx6UXDPS0QMjUM4bio2
azVZqYVJw1oLhNkZV4OlUowgGkwbE/zmTPhqSTF2f8+/SYSNUXtE8+rvq9tIdquv
HRxl417jdbHgaDzntgCJygt9t7Wn9rKT1qZbkxV8AitXqbxOQt+vyCsutERvS4eK
J6JtfN4QV1e7VxJYAiP74zwRQWPypmMkHm7yTUX/E6PiFVhXtHgy+ZZL3W5faI27
DP+eLBaA1aCIoyXAFY/YPj38X9terXurmaK5cuxlXwGhvfLhnMrhkPzdHtyM/rG7
Q93b+RxzuvRWxeTSdkwu1XAZTZFTPN09NcTArXzwc5ydEnz/YmrzAbsqBlwcZRT9
bzGbBmIL4oiuhQVJbL5pXrFxDZcIrVTPGgG01Z1RQWowFoowUpWwdKs9Tfl4G+Oc
K1w56nlk7rd6oVZWN/nob/SX8epICpEL5W/QhmkaOon3sLlf26Ess8LUPzE+uHUq
2rnJqetoyzziKAixGiewXIDdcIbaIOdOBf/QpLaTONXuv1cqJkTMmRQIloUupP+v
LxigZFUunYjxlIHMn6TZ6JphdDneG201KRaYPkV+MEUNGxqzGVw8/auADgThqMaz
GJR18eL2ItCIAw+S1Pz81YXM5dGBabY9IhtUfhfW6U2yACUDjskDl/MF1kyOa5V5
V1i1HwioHyL1XYfIiaNHCa6cYcbHVIo5zV40WtgrZGeKrvhSEMqvBlAw4+XhzmnQ
fw0UajAQ1B6LwiG8qFFqFwO1r0ZR18vxdcPuvOSkz401Ep/cYFuTkYoBwBeP3w6o
E868z/UQMgTibhIkOue20LGxQm/8b8GMGPN9p/DUvCZ410nL69nUm9GTjcTIJvJs
tLquXqsweifqikI1PZ5ATbh5SsM/GY1m/8FEjGSFVVlj5DKWPuDlY57sNWzr1GXn
vVjoBl8u096Xsowx/f3+pTnTUiSmvysmNb1umRQrGcP9DHbSdc0/oIPOK+FZWOul
5IXS6ymNuwJeD25cEquQg+sJ8LAj13O1zjdp6Z39X+KO3dCbSF0OBaCRRz8F1w0p
p5p+fCqiH/awJEgZbweWkcaaDuGGyyIJM2kjUVqCScaYlPdPbwlUssNIJsRKHUei
nm/5nClQ5cHdm0pxV120bA0/hEQSAwPuVNQgMYQOYr0HTWpkcr5YS979fMY6KwP7
uI7DVnxcxtqKOdsCOUV+IDjXdReycTrQNtDa39u7zG73ekp9jN4KDpgMI3tDRMon
FxLSb4DOISvGIbSOA+3thSuegPwgX6HwCfEcuUBYGqNAZt7el0sKMcTBRwe8ojjn
yQI/AqLbj4x/MFnSuz17tzbxTKL02R8EfCJVTFSOTasp8QnPVabx8w0/ecYdJjs4
z0TPbj2DAm/d9WxfPo/qmLBeOgq1a2i0Lfq+23kVqnPSlQJ/6MXqLmXgzHP7ss+C
uSXUitpLhuFy4NL2Gn/LwUvoRevBSBoESrXor2TTaEFbP8Xv0SEF/VNrtt0f7cEj
LDQ1/OdQIugJqih2QIKUXczMZNOEa7j3d+6qOIbkaWUV6dA5EpmfiLnvnxjpt2W2
kOmz9KsJlZgp5Ynvy97BWfKfx+e1TQ0jc1GoK4G8eMECxND9okwOPDpalOi4PNa/
34Kofl4NGKgfG+l8MumaGKZci0RTttqKvC5/6HXMGDJ62XXI2MKBCFxQZ4mMVR7p
Ft4VOFnFsTDB8yFy7MbbiRLkWcoTH7vJ3/omyv/6s8YmT6Co6rIhP8trkv4j0nxC
JiJj+mjQA7UbhXbXTl6Y9XPrpX6Qe79UUT9OTBztyeRCIGLFk3RobKws4p771R81
Sxe5FRlpK+QVAaQf4V1TEoFvERvFzBDc9Zkv86gxL12XdW88ANfn586wjBT7t4Nh
LtoSN7hMFcTJTsD/a6ifeuKRBLUfMmf4/H0hhHgFuHWsMyRI/YKjuPXkUucmL2cD
1wEDsAQ7KDATm1Nly+9+98ZBT1Y/3F83UySlyCKvTdEEPMsdDrv6/AEfaZIvHSVp
VZz6CbHfqG+lPD9+Lfc5wu4q7yhqhBcX3pACVqgZngKvbITpl65/n30KkDqTO1Rg
yoD/ig0W/GavtKV3cpy5gz+r0Oci2pGJ9preEU3FmSmkhqKNtWOaXQnhvTpJP3x3
gHuI/thgikerHDmNAm/G6ckmC2JW/iYoEwa0Ii+xdyCIzdAY9zZbhDPDXANRKB9I
uA3nU7I+RsqqCn+f86btTx7oar6mVxf8IFiK/hwBbwnkOIoNskZud6yuok6ruG3q
lQqFGuEN8iBfxhpOsQFZhEmJTerxsIVtTfwS1VDnLlxLlIItQkIbPyHZKYcLc7Y/
Hd4nsZU8FWYyALXWQ99XC5OaaFRBIV8x8KKC6IV7Xcv/uXw1XScJBxV42K44lGAt
yNYza1nTLA+A3WC30ZxaG2khDDD/yGtixBMMrsjhQSFfXQmgo06Cgm+sgpL44idz
kVtDpa9T3UKlJ+njNRagGCHLu/4PrG5Dd7CMMtXLFVmzuENuAiORYrd+5RvkUqKs
0UHpvDS+3VNlqcwb6agnDHQ9pNoQcrqbsFAEiQ8jdl36iEbYF0PnsfTkFhfn6vp4
PTA0dOFLKx/yTh/HYInk4FKe5DCm42rYDoNeQWGy58ZToCYorkMIwrAAIiRiGvCx
FNNnXHs8x4PzO+8b6a0dL9MbBpj8TMhoiUEuaEehhQJPPWFUWS9GTIxFs2wppJgX
g7vEYld5R63xIZVEHytERKHp0y4GuMQBOOvLmD5RBeb/vSNp0eLXQPBILm8y7bNe
Eno60+++/QiuRV2GG75oazFzqSNsOQhF/EXobwPn2ASg6jXDcdZ5DTk2s9xYNtRA
gKfyXYAfFRZgRE+XN9lKS7s4O66qLeBE+PmeIhcd2PK7CKUk669V3/aemmzKNQGL
+DY4bYDQyUMTRZeVgAszC3azWUb34xHhmsTAeAtL9wBfybHHLzQqYIquYYZOL3BE
LC203gzRst36YFwoTo/egHhyULR7IxI9kDgqQJDLh4NNb7uBMweQrlIX1aHgDZbi
1r55yIajOHsfQW+mk7ka5llILmoJys/AJPdhoI9SSyvzjET+S7Or0nTEc3SJva3W
FVrYvDZ3h6bYRmWDRWw3s86/AUhWZzSUfjqRMkWLCrIBOTYRu6uX1jlylglUrvey
3sJYclzJQjgyV36nwdz/j16WUKWif3927f9sMQx1kbN1mzXBc+9bJ2YyQxnA6LPV
FFxuH9JdQv6d7hHdSdzHxzGjNonzW1z2jUtt2cONOYZUcy3pwiIkPUSfJ7tIRICx
Y9kf7EAvNaKn0+9KL4HePWtkU5U8iWhP3LU9amXPwfS4/norkiOLxrpX4xmdGFn3
Ljst99xpiXcmZzKnHpB+vcj7KFJ3ah/qr+5siQ7sgrEzjeWSjPQfaL3NDuHcRmLt
slwrxsa61Xb761hghwje9CD44jksFIyhr9Y5orlKgMJ7NYZ/vMPN8C9EQ9nG/3yl
ssCIEOob65Xr5JuIl9i6yCymU0KBC6M3Yaud2oLAAqUAkgK9k2jsM5/YpQ/NPAuD
NataSBCdAssPDV8D0iIh4/RHmYODlESbte2X2r20/DAUftP/imyqghEP4NhNcT1f
jHPl8TcTZBfh4CfIu8qtUFGXegDa+k43Tk65W1rBGc5HcUCxAE38V9ITZKAxjhn7
TgkeO/sJ4/6walPWwVgxkxgGAAwzFh2YBz5NpW17w5tUGtn3p0Nn4Erk8rTe+KOZ
6k5KBdksfUIF9sHLZw0PrN7UM1Tqgbt2zVCkAbrnvIwJ+j7iI6NryAkS/neQ/miy
oDlYcIihaEGwJXOGzNENqNrH0OcJUuvsZAK3dY2v3cFLZOc2auoUCAtJX6iCWrJY
5so+OMkcfcQ+43womj5cMzofQ8b79RT41TcjvZq4J7QECuMUGWUKFPE8geos1PNc
Cxa9rBh/f08kA9kmIZgwlvKzXWOOgodFmFFSwAZ7m5ugYRqEujJWvFqYfG18j7qu
04gRUpIxkKX8zNoX66IkFKihl1ID0I/1xxtaG5KD2OeYkpZLTiz2yHOiXV1I1LY9
BkYFRHCogmd4LAcjmHUfW/CPuNbxYSknZNyr0XPF481tQoyo0vbVD73BrWwLAkmi
D2hhqwwyb+n31MUCZcqQdy3h4KDTAR48FGLCFsuBsoGsef+xXKcyYjsiVwm5CAIB
coZLvcpEGkwWkYGTk+LhIq9GaU+33dgGYeSAUckM3yquRzcxnsPS6003nvfXqx7E
qj8pW7lJXHvgZlinAoLAppsgAtcqKJ+YSxhQNtDxUN2OjZeDYC8ZPjKoqsITQ76H
3vISKoZaialh558PYdR0tYBX3kGRYxPegFExUYI/HgdTVh8Q5G0nYo2+Pq82dMeh
LNf5v2J2eq1mtPnks+urs//bd6/K1yJQFnV+fL7AxYt6N7s/jDV3SVrotnmyr5Pz
7cm6idQ8FYtvGZlKAOunV0iIUHZWB/UWuFoYWoZEsFvYWn22E7dHffYl+//JLUUC
zeOmJZ/cd148WRnahMQ9PK5arKJvRvWrzqlxPEMrrI19lHRe5vkmqb4iXbkmkJOx
RfZuDKLA/KA6TT0bs3s/pv81bYoNQMCNnPq05TT4nDSfm6Smqyj6M6MDEZ6ecP/0
/tv2UZ7N7vchbo9T8jgO7Icna678ngE6eucgBoluGmd0hs5oT64aPoPMCzBDzihg
/Mqqaps26mrm4gre9tWgO8OxUQhNsmrbSfgBUc2jbcquTfeHP0fSTPk5GcyCxZ5a
4ETVDi2m0i2aN5A18EpUr55RjMkdfvtCcXV+cyHG9F9cplrTPgEip8ox5dVgZ1SB
xgRtYFjXEngeNffu7PDPlhEVDqCg2MbZ5iCkEDr1h+IW35S2eWjkhDKsS/D1s/dd
k7NRx0pvmJWx+VsNsokqvZeUnFXHCBq150HQI1I29n0C0AfD+fbmmXmLQcMXT/58
AEquxSSFSghiBhJSUpRbmP0sHLnMK1la42P9S7cA41K+xb0yj4ZZ5x/5HJINnuvw
XKJzwATV6YDUfe4mzoIHuw6bV/M6CDvcqryTkUkxWooW8gES+3zAPt6TMoV2ocq7
APgthGrfCHjO/VqyDX7UXWZ2ezzqdybToORrWopgaNtinc5uI3Ku1Mt3q6RA1O94
JIDf71UbVJcs3yEbmt05g7InaRz8xSU4/tXmRERVUpGFSmyeP1p/R1hly2KjhbMy
8WYOwn/OaoiLbnFwkXlpFPRJmDfSLs/bO5ZILUTyPAMI4+Sm0ZgQ4m8u77CnWUQF
I1zBKtn7o+VfVqEQK+g9gN0kuWO0lUJSKd7JuSofDhoGgZ25K8ldff51Hq3Qye5r
2w94KQjaWuoZXV+3wzf+Bo4XSguLLs+SjVkmrwep2L2oY5TouV5gZvOgso8eoJLI
kQ1MGPkwcEt/SihIqJEW22nyH5CMCVoeA4zteP/kaWRYcIuHE7JoeJYZGGdsTeM6
E8upW99pdgDs+adsR1OtfRDK+I9BeWNeOMFD217n9vV4NxybYdN4WKX49p7ICTQ/
4lF1CxlUKrsLb9AZvWhVrsD074jtO41A4ZG6Jk29X8+mPPld45Ja63cMOOO7XI/f
xXeSNp6WLuXkvBOsud++x8qDhmYShx51tYXFKTdQZIHG53sSfiNmLBGvXMylP7j1
udEZr6hbjHyCZyQLiH17eBISHFOfUNFklddQ+3MEkYmHkrCCtQxcl5xQi5JyXC8f
J6NevlejJsoWwwjDt5iLp6W/2CA7ZIJURdlrvmXZvrT+/fe6h6Qop8OYHVGcZrzL
ZCROxDVnIvuM3Ij4ca76Za5tJPS77XOum65iLOVkypchWVEnwQUvhQNBM43LXK/x
/52Tljtebjm7ld59hiVBdlT1gpNu7EPbrBtsOAqVq2VixDwial14D7bAhQcziQmS
N5ZNwT59SoQMrimpbugsdeupMI+iM6Ad7Jzcwp3rCr1SYcqKL+P7/s1hMCwY0IdX
ir8i52KlF1U5fIkRCzU5H3xHXPFtnn8OZ3jSoDecQbBrWhEAV2PEUayd2Fcnl2pC
6WKZp0yDVI4dWSe1xvRl0TWYnrJQkHVWDTNC1zQJ6roktSHVidQAGOIFR8NB6SWy
xvufRXrU3vu9arX5OSJusP0pl4zc283izTigcMiqwYZcNQN7QLMRmhDL8AcO9smN
yXMIZiGaT4kWD3MoaLxEgyjiAkJA6dH6Iao9cbf1a2TcI565SUJXIp2Qsv2o1XR3
/yiLwejVmCcSkPVOT+ZBxPxwoUJoXeV3HHi8KxHnpf8ZiVX+aunKSPegrt3Pt5n7
svik4zr/Oag0WRL5aTQURHSKkNtD5iwKMKMAAycgNcnhV4L41b5+AZYK5K8JXpng
MiIFf2jM5fsXDzy68a7VlwyaQPLiMx8i9IUXLCKP6VosKGcRGkrupY8DrMIvAZjl
Qez7xsKGo2+5lg/3v3nwouyiSUca12SJXYC+IstUnYDl8Z3W7oNe/XQvUu4GAn2c
X8e2h5+ixUfSrjJjQHaC3pbvmAQu+EPqqCZKw1wGkcibLdi4torLzm2XY2Ejq50r
M+3lWoG23PJmsD40KLjRDg/Bt42jtO8y6vPplAoxP8or/AC0RV6syTQIqYSiCYPl
fiAZRkLC7BswVeEf8PswkDmI63WcYMozKkwQ1FruGsAZrk6RAokbaBubNjTl2Had
XpvWF71jyZ5ZoQ6pBf1WeISy/hzxtgwQLFrwghTUn6ny6HJRmxRkyXWXX55k8VSC
Qrz1NqNlW0BgAX9/P3yE8aGxZrDsfUuLK73PtRm2y6aubKsumk9YTx93v18ZCdxR
Jd1gvl2+kDWQQy4uGVKan5VAuQzVEb2VUuPAoekcVosjzSwkgLADjPtmOtdD42Wx
VEIvdpzyq/FBa8gdQ3vsPOYwBDElZRaTiVjl9rNHXUQeWkM/xoGcApo02TS0vZPz
rfnybSV5+vzoLR0vNTL+EVQwxcXZU9ZU+WJyijJydFymzDa7zF0Eajdp7mdZ1Meh
boI4015yRfDA7RG4e7zwoLkQQDkrxCRaXWbkCuFNMD71H2GuSbk/AsH4PEm2PmBw
i0iTucZTqraRkqwN2S7gSEStMv1CIIb9d2JxBw7wz7GGg0D0D3xbeJ/y+W0+bIs6
yDWygAl9eNwIxkDYMSqr41ucYgn65KZCWjNuVr3PbbDUkCQ/efeKEYIlMnl6UYqp
nsELEPkURVeZipZASW4134GWkK2GtGeZhjJECO44Sh9U+zoCXXINSoNexuuGgHRK
VKoO4NC8xXxBW/2EPYpW0O+KVjZjsBcEmhchER0JZZNPtLp2zYRXs6NKCGspDqVY
xkR+1/FtiZ1esA57DFzwgLxDtDrog0OHNzD5MW324zHj0S4tqdW3MCjQFaSJGM6q
8p9vy0E7KoqhlMBcp2x2BVXps3XfbaOLeGeg1vFBaG4F6+tj3GrNxufpRdJo2Jrf
5jv+szdOGfppcpWnqwTiaQ8nlB/gAN2paD0eYvW46JWG6Q0qYIm+J1ZMiWWNWbk5
LW0/KrQvX1tPbxpQwKZlDvKfd3FoFTNO1wumf/I0xHgxwjz5uLALWvQSiOGtNK4K
K/SpOA3YR5SBs4Rh/UkqoMveLU6IFn1SKRu8c7iT3/v+QQdKyz2Mfn9GnHSBxsXo
QKVAwIhutAH3GQ4ZNzhxr4rdB7KcnXOTGS87FSUGhoU0JAwxRZHXIcm8LQ0cvi9e
G8+UW9t+XD3Iz8oci8uS1oa0wTyr/bMTE7L+Hohrbm3eAviYyKIz6nebYBMr6TGU
jN8LiBX+wrHzSrCA1yJOUf/wE5WIpKs4RAs7vnLnwZaXRikakXurPz+g15TPRAEh
2b3NTSxUcOv90Il5UigUaE4Bh4xRxxbPBFbWAu9RFAYnagRWMc6pV7eNJ8E4tkoX
t8bEFnsN4ZQceM8uUlg1Ss1lpJIsSsqbaU/jvIADADrZJCpi2G7EPURgTCZNUzgO
VbWJzTJXj3n0xXu0ee48aNfMbigpoM0pVkOjmOKTXA6qjvasECOSWRv9psCK9HOw
K3aAlHpjsEWoHRJiKTUjE7Q2eX/m7ScW7+D0x4UgatQVmYjiLMXPmnmqG9pNSak/
WUnEyQTfTLKgRNG1O8/A41g/o6oYxl4/+2wgwGu6RoERdkNkzIKQOwglkFxdP0qR
sweCIa2fW6Dr/hvJVACr2mBZt/pamfGDyLQTFTiifrc5UvUALpqWXej56zVEO9tC
IGW8ZoOx1dF2vQG73kcErwvh3JB+3DuQ7DEO2/ORyJAzASpdUNT47vXjiHouthQA
65vOkxZyIF2l2W5+KuoYDgSfM+GDM1wjCMj5L1xcA2x71y8UFpcU40qrOEI429hl
c5ZjApgAYtkbFoZneQ0SwmuvWqOAgYOAXbtvQMi0EW49HWmXO7Ic/tLWiH6V36I4
xVrZaqkk9qcWra7TyqBdBy+m8PoY0GVdvxgeix0gc+zKIxzn08ruq4aC/Y16hScX
DL7ta5hKL3hHWVvJ2WK5Rit32Y+t8KKRWec3F8rdZrxyCxz+GOwFrCjCaWWImIw8
JnYRYz+mOJSn/N5Q0LPfDEPeb7LqWVHe7jKSm+F+EHIXgZyFexUq9jzq95T2xvmQ
oKAW5IHSEVdEaE6no9ERm6pzIBWZfkyBVXWYQ/s4dnAa50JjwGVYrUTLeYFVaEgu
0skMGJOnnc9nR88XBYadXmO43SjnxuhahM04j8yKFdBOXC2VoTY9IGIegjLcU9b0
BlqZvgKqYdJ4UIUvl+QdTHlb7GnjoZWScUzn7vRXjqKRsdgLKhtht7LvRJHDoltf
KOk9Qc8Q9UfZ4ShDifKj4QTSbVo5LjPtQFqQK64mLhEqPA6yYgWnq8T4rDWG4dDF
GQ7CWz0qbyfeT0IyevUc6Zq4ol5IeUvuKy+vnc5aPt7Ym1Ztq70gA4q+qFJAUg9O
m994Dx7ypwrEHkxbzmmvKn2yem0DKDj20/B2TyZ42FFiTZ8gLU0CwAOTRYTk8i3G
PYYVKIxP0Q0OnZmF1TnqSdT/AgkVwWrnMDrJX16+5xebuz8soqGJ1al0v1i65ElL
bvo8RPqdyewnzj8RyEO2VXUn3IlwvpGnVoFOVPotwu7B0mYVdDR3uzsawdivnkaK
N2OKHFFQS918ofJX+hg9IrJuj2IrRv1orxOw3tYVg6Qs3kQQJYoJ9PfTXbCKP1IN
jmpgQPfXqlhIwocr5Vhs9ooX1ZR6S8bQSaqgAzRURiup3olkpmWwZe2RLDs3uqxA
tJmk8f9A8/d+dd39BhOk24DOlAKWRyUWQAXHALLl9VmM/HE1HUzUkL4me44BCcvl
Lo179VMWBfM2rTgU35OmhgFgK1bTtZYF0FDt7JN6kcpw9NkCdKQoEOtnQb/HRtiA
SLobsK6WP3m/oD14JricWX+PiByZXSQxPswFChh8EQI/CohT2DrD3NtbnTUkOK6V
83+ydUolTH55/aMRTsu5x4X42eiQVrEcSHN8wbCWCAy1qoHcl4XHlJpVkkyu476Y
Uu4weBXIq5egWNFB+IQgvoTf6u2Eh5E2qQVUPcGDBUHNtUe93qeOpeM08L6YV2gK
bMaS7uz9ltJFMFkw2WQSSZah03Ssj+qa9S8LRmt6bsfB3HklGSb8bnz9OERTmVO9
Cs/exHgzWTWumz97+3vZ4nF8beuY9FT4bouHqSwU0mCYlm52CnAUmMJ9iUwcvcok
d7x5j0pWs6holOJGg8A4AZD9Nn1hwCfLJBeL+49FJNNkYMnBM0cv+KBbalveJfrN
YsnJY09xwQS7GLBcCvZMUTSAJcmQhpGLP2mhPb7LZeEARlB8/xYat13+KY4ueDoH
rQ1uAqow/eRDYowv/25KSBe/qIhYXiPDdnVeGHoGAngEtS1zGVHy8qOAP2dcq7Nu
+q8B2K76kjph1eEr2cmYy+uOI1lUipKvuJnDSG/Ict+juTwn7HPvw9v9KgIWXnO2
ue3fq5Yr0C7zVB7/KGme+A8CTiTsj7HBWXnV9BZ36SvIGMlowO5/USUYPhMhLwQs
CTCY6OKpDevKaA/51SpYErki2dik9k5JVo4QmPZTFDxgoYvK+j+Ro7h21Pff/jAd
d7Z4YQ8KIt41jIcRgTNAUMY9A/MRGcXOx1k1/0zSEgwwILDc8JfVoJgNA1CYoabH
pFBDgQhDr89Dx7qPYUycdVxp1FbJvWlsWNnngH99QAqotclMszAf52rh+QS/dRoM
kp373hQWivv/Iwx729kaFH/pDeUJCUyPkkoO6SGbxZGVKAl/MwsOsnfpbgw5t9X/
bC21+phJ9ow3fw4kOJYUEmHxrqW4t0lsdPPRl4jExNvxr/rFY4PvqEVI5wj53+fN
ALs7tDlKA+MiqOZM7T8BjPPODhVELHzUTcjWrb94eC635F6kEqX0IuG7d6LCUNgq
12VeTDxfkrnJ59/ksalUlMjepxTJ8b44nQi8+7MfGclfBfP6EScOd+ilM1/GvII/
flQbIulIQA1DWblN4dCf3nKvgao2jdv1TSsTnAnJluHdupts7uiVY5o50CwoeFjF
zC7BKzZBuN14nLXBnIbw3yf+55xCKiX/eZSts3JRBY+0bGCQApaHhj4UN/oLsr7/
Kzt3nqb7PCCWqsoMUYwhs0yfwwSj7jYdprgmkMBdnEgLaKrWyRBVTv+KlsuZKw3m
BjV0xCMGSra2FIO34hphv+u6IFYihHy9Z56DDBEUl6lgfOtpippr9b7mUfdjZH9O
ouqdYnZulwjNg7vs/rrZ4rShCkWQRhBgWnBS5kOy3k+LlHJsPYJZzwHfQ3AjoMwW
GeN8+uCSGFt+wxRh6FEsIxx9PkFoCwDiTv0UIRVlYitXX2sJ1f+YC0UUDgWsiiEi
WxfectJayqYW73yl5nXIgYP+R0sHg5V5F7phdzn9nhw65BNxAYwVHvkbRJdUeLUk
asRM2t/deWJI/fkBLWofg+vk/q/vWOcn1IW5A85JiDlfpHHQoAxjxKnvDEdGAVIT
N0jWL1veb166DoaK8pTOdmZcR+mTmILkCrWQXzgd+UM4yvxmbIc7EfqXN+4p2/qu
mH2aMQ/TqFYNB4rk189w/s5R2VyYsxCRd0I86iUucr7f/v8t1e6NqOhGxNHeRlU2
mQ0mjArPDawJaPhJkc0TTpuyWRo5XBJXRDGV+qQJik2s4aUB9gHmTdTxCkF1Ii5f
tRtvPr5tbdeglMj/D9lH5HDK9214Igh1kEiNW/Qmbe+vZ29FicqwIADEmUUm54C/
JJJ//DZlKqG/pJO2mCrqKY4R4oYuqeDVQ2cBivz84CHe0HAuNzJrEINCJJnMj0f9
SdxMB1J4swMYAnyzJ/kqGdatvC2EdbXgkERB6QlUj4fe4wJEZwFPk8iYBCqW5Den
t7N29ni55cNw5evVH20aD6aEEEhN3f2/cMTE7Hye63eazFBbNVy50iBYcTSfHEb0
e1Ayw4QPmTZb5bXyCM9l4WGjOibfj1/F4gRQsmI7u0ZAIuCT2CH7kz2HmRtMIoqV
awA5TWvrulF86lA34Dfa34A4qcdIF9N0+bQUqseedLiA7nikkP5QEuKYNLvCu1BL
Q78KXF7wHhdYhe0Mn56lYIOlI1fgDQMSmISt1YMxEWN4dSBgzrZf8iWql98LX5Hi
Y4doFocibPMbfy9nMYX2akyhL5iGaBhMOLWkULubNqDoCByvUBhz91TiPxL4aid/
HRabo284vHBAvi8NocG3Y1qFkdvSul75pb1Pl9iYsKkcY69NHVEUk0C9aVNX/Ebb
WS2/PbT1cis3Totld9jUKSbQcI7Y4M83H9HF3lG+hry7kcsAnt8wnvv/9fEsB1Dn
DYztcS0szmjeL9EfWrqf7eRZizntr0HmV+D5iGXISe+mfdUL9Bn9Nn+R00DEzuMg
7c/Bd1iMKfbWo+LRc2sVvDBgUn6xxw+HH/FcGc8na7txlKICin9MXmVFW/foq+e/
aJHlOjU3c7///q0INCbaZNBvPdemyKk1PT6oBVFHb6i9FR2O4HL2s20zU6peZM/M
YGuUJzbmpAtYGCraAiUAO9iluCX0p5YvVwwz2q40ANpALpWxJWL82GLych6FN8TG
wrg6dl+gDfF4y7x2FC1CLNK6g+ys8iJgZEYw3GTFYcI+D95BfVhNPki29f0Lp8EE
I2O6LZIgUs5ia66GDwXEqag2uSQg9139t4dXoDly3M2Qv4X5bHTT/pZrXyuHZ6OD
3HGK/7LgqKJooEgb3dyaaExCKvNjyYMWVHFdxnKjVR49/EnVUEjqezylMwviKo5/
YotiNiWVeL0rutDshl8rS9c1rBsiXzFOgYJZbvjeOBeZFb14spkPJDdQfrYwFMBd
seZm40tt8nNsNC7dAU91kHShVq6PAsVsx2ei9eceo1BrEkji2JSVSU+kxjqRyXNn
MT56h5rHVD9H6rkau/WSkQQqq7izKkrJ6o3/hAfEUAkbzSdhg6HNZHoBq548S+uJ
GObVnZuW9JCflpqwLSGUR+6MovQMga430ep1Qqc4gp/+4Yi60aW8G40q5CW70VMY
gWprqHwVHCJKzOgHXm8ifQQeaMki7jU+QIn/uzfOfLSbJHH6Pb9F/QDZYs4oRrhN
ivJ3fE86NVTHtk7i25VXP8LW65h4VX0fSP0rksAx/jc11PoPi1NavcezLKU1zcZC
bWc4wcpdGjSdDTyVrbCeNks0wDCPar0XH9F7RLHG0KuwllRKhcEsj7v0WeHI9IAx
TYKxypG92lqEoM494S3oBoXRvI3gz/RIo6PGseTAG1Cd/3UayBOzOtFUwY3GiXQX
wV33Z7ai3neevoS9aMN55aKuZb79tJKprlH22UypAFXHBe6PLXQ5bshLmG2dyQf9
bluW4ICuG/4gRHKMXsr4Cyigbk5W+X4iZaV5LkL7HneXB2gPB9oJqTvXcBXWiiCe
3HExVlFMgzwLOM9/v1KgL0gCGTEGTDuFE2Nf5SVNQcpAn8KTupbeCBYbjS6AYXK6
bScf+4uyYia29YPFi3Wu53YcK5/8JDqaxXQGBug0pP/c0ppJYrA7aI9YTjHt1B40
2z9P4wF0pu0Bs4uaND7VnOao4s01RWnFhLEqpQfSbFifUmxMy0XXYZDyJxaB2/dj
7MqXG9Of0zEdjRvXDJLfpAeuLpt0xRH7GTY7ESBvL0mYk/FYPjSbQHlQydmrR/r7
dzowt66J/HJ55sR2OItJ0VTNhBVL+AiSZpfafsrNscDoAAGMTK8/RWR8VuVVBwdH
nTJm3uxMYbvhrcP+BDimwNpIQkL/SZR9pP82wN4dNAPrPzkPB9w1MhoIJN7sCAWW
cHxjRiwkKkujGEs0IcLfhtmgvJP1HiBd9ZkQG+YbM+7dAz4D2ntqLB4Gd0wzJdDo
LC6dCe4ZjrLgmnkyU4/tP+ByedOFAEAsFSxSm3vAdHehirkx0HHbuyACsw56iygs
4ap504A9W3JqBCEO9/dxbc/plZWKiEymm0ytu4/yMvnUeRQX2stUbcKlNxXNTWgD
m+F9d1VxljC2TIDAB6QltLxVuSjY/6WUxil4GhkZQ2rF3D7WfUHgWjbQmxS4aDNU
r6/PvWjYSyI2eUUMBp1RiyFok2HbEQKCp02otpb5bBLplIpGrv12XtX5fCopuDo5
3aBYPi6GiQpSYI9KQUZ/NIJSGb7rcheldd9+Y+21Vnf4/Ayc+00RgsUAFsG/qH2n
u/nMI07KRUVmTBV9az8TieB7qaEdn1EwnXVPe77Ve7LpJRt8JuL0gfl5SxA6vx47
cBWWyvEkBlVAioTwUgOxX497iHLw3NCoBfN1wy+QVlMzAxnhOETLfUwgqVUZNmzA
b7VsP34+2yy+zSJpRZ/on3sGMnDTRDtJduFHp6ZIk+S0VoUxwCgxLUgBhNpoGZJK
8K5B7TfrK4gX/4OOF7tq37k87J2zzR/9l9VXgnIJPOGqzLXGpXW0j9ypsaIiH9it
0jd4y+54cHBD9Mn6pgwl5V7oYBMZl2lQGDLJwNCkvWU66kaz4uQjRGb+NkG+2yDx
xCo9TEMqnM4107UVsaPPXSXvbq8tTIdByDOSu+h5WjmEJBlCI0nkxt3mls5MgN/d
4pqTOCMqfTVipi0W0fTqTvWz5UZjXk//CNace7C8KD75M+JgwHUdYFtUAqwvx95k
jj/wAtwYwiYKw6XuS7B7HWA8WtRIIZlVTQ1UsCB0F+otz0IRWI6XiG/jISbSJmBV
/ympuTH/Kr/loDT2QRXMkfH0d64xnOQSugZNFTIZ2ROvHRtvAqsU31Zr2rpLYamB
Js16a29kZQn6Tqq1VKaZ+16aKLt8GrRy8qL0YpeUV6RCQu6G2VxzM/kNejIMIBK1
tFC2xsvFZUeEjfQeNuNX9LkiCa8iGa1oRpsVhg6IjO6iDkeXuvsXYQit5DkrHGz/
CgnhYlGRTY5ppsmFiu7ebGEdyXZT9MZ3PIcDmpGh9DvXuZKjmX9TOsBo1wyXRe0D
9+M3OZMcuztgQ/G0Ykrv3Zj0g3ceCb+8BoegngUqm1V/yD8OrATkJqwdYRGkHr9z
LdckD/bLcdiHM4h0+xmCBNOd0/QoC0mB1mXC8271ZDO+1Gyn2Sq3C9mdAcGv+NUZ
SckLZs/157NfyFZ8xmBEyUMEwAmtESecfFHFDgP3uFkuQNmPYuRRpfLG2q8xzgy/
xmEaiqVZGRvFaHYhpYbR4u7YcXxGFNy4cW74MF9HojQhYWzCPtqPpn6FYKEio3Ru
9DykiuOLjaRM9Bwa6qNEsOoLV7C4x1Qke96v8yH3L3vh43IPyHgoQWyV6V7clupj
ANDXNAv8NAqxoPpLytRL8hIcVZfbkiC+iJHnjJwpwYKV8ZLHoIedohrwbQsp9/cK
3N2My6aNd41sgZ8GEUVMnQitrE3yyGWwmEtfmz1RjkwxSJNgoBd28M3FCvQgWtdA
xENEsaxvFa4ugV+UacBgssboX0FqqtdvtM7/B8DFQyHZT27ssUPeX3ML4+VxAlHg
kh9eG4M930rsaO4pCoiEu86ZI6g0Hs9/y/3rF7aMCX3mr3OvHbcwOJSTcTO+TKAR
yHx+4U04dVVz8T+RYB6tc8yDf539493WHceDEXKMLPCXnKKuboI0IEh16OOyt0US
g2VSPdnMvYU9Vogjr53vdpozHSSofiPy+/LTjCwReT54y816oLTLfTlOt+sPNmHr
fwDchqHGw1bpaMc1zw+6RgxP6yTjBKtabvRjf8ZOhsFW7Ofj4vLJ3tTfW2U/1Cgq
40Vr+ft0VoTqC2V1y9CXISb4I+src+xkX9EQJDBvRAbkbAxI/ilXyGILIB/ci0ab
4q3E8tEZG7Jj3erWtIaLIAba7/Cxhm4MS/3YIj4+pfzCKOjDTQDcMnbyamRwSZpr
FMo9ivZYof02y7ZYYVGKjbpt6CvcHJFzsvrEplWIYVaf8VkMY2QunQC9r5qchtyg
wB2j52SzMBnyFG9jPgI3Bebf3kJGA0WCWZhX1yIXfkn/+Z3OE49qW0a1mar29cc6
vI3FFvR+wp5WCkhF1AYlMDxAfxi4QhtGP1R4NEQIYvwkok9I3eJ7Cl8LLavyKoBG
/JGtezP4qASpxml4axbTd6SrKVdLjL/k7QYsE2RRZiZTwsdxUH0BJh7JSzWiOWUI
R12CD1FDCWUg5ONTaeE7gPAWPkZnRmSxOE6THODtKMee6g4XiqF04v2Q4wSVWVvh
bN0028bs0gxuELBLyvsHs86oZRUDSvYT+tD4JhvDsoCLTzZebZqyJR5U10GPC3hG
8WSW7luTaH3Y2w3jLe2+5cRc0WKzuFC91J072JDquqSBM6E+0rcoTs++sUa8bL4n
NSv+H2q8I9l3mg/bpMQd/I9Oqm4ksNjjdSPi9tubnc1Xz2/wdQ9HYpozdHLfz+AA
hW+8nQo/ErsS+XD11R8YozbN3hedPi63TdYOY7QBjIiB27u3WlLSRnC3u1ifdsWQ
d6238b4h/Fru21uslsny3oCFCti5AlMUN/sqmOIlY4cFNPvCIL6x6pk4vID5vpKB
ku1NPie1xAcktuqIS3U+MNqcQlSSZ2E6GT4/R4ggGEOarcw1eRNFRr5y7tYOFEc2
UkO6NHjF/7vZqDr/JeMqNQU3s7zqmgqpGmG/07jj4RIptnSVguGOpwAW8qxX1V40
s4AZ/JvO+6t47qpufNJwf4Y12tTp79NlUJWapaOqcovAU32yry7hjO1vSW8XEj5o
MmOXL7xAE7ucapgfkPx06MMAGyqRwVAPAAg3Lj8EweDCnQuwAUT2v2D3K4xT53oF
fm73IrcRPL5fqHKWN/7lTInAdDuFKzmdbB+naH835jjH+jrr97XjD0oWUBXRzT9q
Ea1zBqLquezLnliAM547A5r/TcgZtucEjlF9Mcaw5IrUetR0yoKn50Hz2UHk7gkN
BArKF7fluXNjkRHtYNWzKGy/tidnUDIuIUUsYB7sZhMJt+XYEJkEedLMapxSxafl
l0q6hh8ss25nP0dkKqQqpQkDPuugMZZpil4PSQJtZ0kLdln34yOTuhSjZuJWSI+f
3yR5xmXCyzEyzPyYvf5hLFyGY0+/oOiNRxugyZNPW7HfEbuKBmfsK17yBnmqWJOR
tms/wEk3tHGJ84qObOhL7PojfCFIj9dO1YmbNsxr6ZZBJOcBKR/12B4dAhkVByfN
Zj76SHMA9q0+S/08iCDy99jcRjCxZViJUFkQ37LSf1krqkMm+hL7qqi8XA+u71lD
7NVPBttVDSLmRidRWGelGO3VL6nVxIuVy5kmctp73uxz9G30zGE3QmFQ3kv7RVuT
TwH6M7DRdWFwKyL7gSEAMNE00wVaraWheCZ6k7H2MxLIZJYuY6tYELRvv+eUqgty
fsOM62AT9oOHyhMrVjPoHNhk4ZOF7LLLfXDFmOjBXN1N2QXWKtSe8wVkuF/kU/39
roOESDBXeWMtwZH7ZRtw57VTAZm3Vh89TAIoLnuuxQ68h3Hs1jfQQirI6nCmr0Fp
cgyhDjhzhtQFQePEJ8hXm4Ej6K8IvVqw+aZs9DOmnjj0VYtDKdVBF/sxq6Lq+Le4
7FbKXmisjLiSh5MxRqqV9R9may5WqloKU1EvNj8JvohGs3JcGHUS+2OqfTMBK4NM
aV+/cbKeOEV9VO5dnP/8JTfRH2yOmJXDfixf4qdBm4R768H5yO67XmypccGe2T3l
KN5AlNVpo7xvgpu8Bt/Lch7Pa7Q5DQLFGExOIgwYXWlhXhAwiiHv601rBl4Buih4
a/du4kXRWbfGXsoOXxCQAm9HNW2VjSpYw5K6tgiF1XkaMp5zqZBfMUWkekoRpXdn
IpmddkjqFZEyqli87eJAfYSxOSweMT7WVZFsPUXalEB1BtiKh4du6nPiyCCcQsjm
gKAeJAGndx1mmFisPbxlOjjyfQ1H6JlLJV/Pa79AA6Pl1JJ0BhAlGBu62JqHVtgX
HzFT2/u7FIRqGQV69crNTO9KF6WOFd/aNs2kFVlUgvszZo/LFW+g2q7WG91T81CB
aeG++iDYR8XZj6I/MbSSMcuCcdSvT1Plg+6AaZC6+durBsHMwMzGesnGQ8a8pWxj
f4KjoT1fVvWlLIe9Nm5O1v9MQhBN9paVAdvUaiytivatmkbEpK0QeEetVXxqcsnf
0D1YP/LijIteiuLkTUmTOYIA8q+K+/M+3lxfKIBXM5eEwYcY/ZkqQxqp7mIfeWEp
nZ21KyJ1mjWvirZM6bsDtGGTDoCB89HWG9wTTyYvoETPOU4TEP2vAtJEBpvwEivR
/kdpNuubs58ceoD+kGmnn/K2ASrjPWzq+14A+XHVwdQp/l2brDT96t0XiwsMGOS3
VN56r15NZD/hxMMRNgOrLxKodmAbbNwfsqyWPVgDTOSdFZyWgFIgHgmmGZU19hNR
7w1OCM/sr2xeoXkHrTODwTYJ3gmHVOEvjPsg3nEuSqDfICRTcovaEVV8Ii++SWjZ
/gUBjHen01sIafRtLPrg6gNUHfYC5rRyeEM+dv1++Zoe5evGnISzLwQ37QwvDW4J
t+K//TVeM3btMAaqof7HQexUSbcNl2L48mSbqFl/4HDtLygG4eLaMKnfJBcTkCk3
MFtYul8sMNW2ekxqn9e0E4zSwPdIpVomj37NnmRc/tWdMgjLmZRRya/YcKa/bwNa
uxLp7LBeRZrUpUW8wzhs3SPAC3RWPnhQlgbhqdZwwwBTr0gmY+Xdv/eDiqA+lYov
0YYkZDgZ6hiFkgK7YXxGgvmfIC5xttooc5CqUbVZGXfw9xSINz65bUIMI0fB7A9i
4HEOXptTbsB3XrUnBjQU7K4HqXbWmLpUZWTstkJLlelfuGxhsMgNe+bSmXFEMY/M
V6gf1XsZV0yJliEMMoimwbSwwnjlqdoZ8jwH3bIA049VEGXF7Lbm48QElf8LlM5r
tMBdmNNY0wYnXLK6xBwPmLCSsG4/cNZs43emHmmu3l6RLXQ2zbicwOOd5rCIJ+Qv
LXZ39d2x9Pm9LxLVFbJGDJ5tN9dRd1hQHQQyw0OdiNCHOmVwow2i6Vc4tZuyo/NM
BZ286VxQKcntpuGXYCwVY+bM6zCYiE4EbyDhXh+1bfbNpyJ36sXZ/w1HJofFn78S
GzCcu3vetrQtQZhiVqHTwIvayLzkdZzwy5RuvHUHIrwVH4dm5h1bDWIyggOGSQwa
itdEHqfXNiwsHTsNAX14BjjB22Nyo3527vsIrbIEkHM16Wd4sUy5FqYVH0QT23dO
zVoM51zPvBqQwj3xZnQX/MkVUfsxPLO606EJUJtLNL1JrCmjazXlk0QNNeVy6wsl
5agPPLmVEzeXm15CByM+Q9/vVclXy/jYy6Oy1pWjHby2uB6hPyyF7IG1hqEeQsud
ZONQqdElQg4zsvLICCym+GvVIIuwdGdJtmiPFDWQUJkStqv+qRals9lkK5FmuViM
nEZVMKxdHrX8cuv/OylbQeU2T4AjMyxowxDwdirSXc4VyoSASUC3YhKXgwfWH3aq
zqRgx+Gko8/IwSfh/DQMJZFepIijeXvx+KDHwPlGQhffpALgLfjvQJdLJY2unm8I
Lkg5yK81GP85EVFB8K5lN012Wyp6C2GL29IJz44Do8GSF8xB1f4XkU7VDqZ6aQo9
/oeAJqzQMkDqcyrQctE+PsEnMDQso1i102+HAzb/lMvpsuBDQsLCs6cG+Dsnkkze
HrP0Kiq0gByTZ8fwSkVeBkWDPMUnkYa37PBsD5PA86kDp0RZcRfJ/300UbeJb4fv
OyceaUQydWGKkcikFdJ1yU5DnqleTUY3dJkvpP/I6thULrCm4Z3zKUNE7ny8Fnby
sXfoxk71UO4IMbq5ZGKk2Jm7Km92Y/g/d1i+1kf6Wwt/XVIBvI0VyW+ON2v60ysE
QzFmAUY6um5J4wn2Bq+0yMD7O8se3MaBaVmzZ/e4bN+pMJ9ENHi3VwHERbgsnFLD
UQEjJrO3hhUbDuNgk1wdftAmD/J+qnjLIKUjCZfX2kwa7/w6D0cP871sdSBOqVdM
N3OQBTz5SwKgoMyYz32EIzortRjKaf0zbOIXlo+fSDMK4TGb+aUjlZ8RFPPssKRa
UkfF/AnJnkS2/RCtAzXUAkVWZ+Msn4ty3G4pRx/sTGyVzZdfwSHFwmkUtBHZ3ESs
BdlsYQEvc42VxFDYHzO50wWlEQTrF1WKbeV/gehhgq1OYyDfxDaQ0AggvtB3W2tP
UYCDQwDa4OcZMVs8CvV4YnoHqFqVrZjf//4Vk2TeQXxeZEVQ+7vnkmDhNj7dPrTm
fGPH6/kSNoZ+cxxxYY8Kbve7WhhfTpa+GGldqrPFpLEfGQvMuC0Wz4MApEu6YtV9
JoLhu5HUdHwsFqRrLn/dguekFyW9wUvAIX4BjkWFkqZg00XtMAbYaLcUmSrD0/EC
A/2VXlHP3JL/m4pl/NpE4b+dPGpuVoL6LZrTZfrSIr5J0/5tiYsUn7I2h4kWttwa
Acclbg6ux5SfSfuJO7WfOTQ3Y6a0tIo7PtDOhWR6qQydK3NoEvI5ma03JKFl0vX1
ajAMcgmU7gatl9xyEj7c7rouc1IJ2SUW5t/f27GvUk4KQM2/DAEXoLotfawyexbA
JvchZb247U3QfXPIMYZ3unTdZUqRU3XloG/3k+YKY15r6au6m69L5u3xGXTwdJkg
BVJDuJAY9AsVvFDPuAxXRHHM8/fvu2kavb4ZYOhnRzuzDSvWdMrPuErVBd1CxiAr
S3DDPxMQ5W1A0bKSORjR1wYVtl0DvKJuI4emF5Uko0co/ZZ8xMZuGeEcso04cGhU
SSjfGzeb7k+OplFcsVZjHVQMcfKNQCHp6OVDT8CTy6cvtlM2iTG6wua7b72sUqH4
24Z3g9Dmun0fC3KIlAq4kl47kzYdinMeY1AfbkFGYDEsMR6VbdiW0B/mDgGsxPfh
zU2zbNe2Zt3nqqqL9m5Fgfd52kAaSjOYekCCyTJpSAeoV4eO/35WFVpuqoGHH7eg
lZFqJ3L/PMc+RjdT2aZMREp40M7bsS/XG/E/ZAY9cKgIWxuYYSqxGIqN4HwzOVpz
dHYUCyQwRZ+yyilhZje2XmqqU379QF06k/dgw9mtzVSB6lEeTcx54kdzbc/nI4/k
IS7dwEfkWxdzwpLzDkbk5Y1p9qG5QQIhBSV1j3WgLfVgzYRRRy6nVtyTL51cyVzL
vO0j0fJcThKC2dJuoyOsdrHtQismybN8YYOdecVxTpIYqx+mZEUA5t4hhNoAa6pH
qbT8mj8V0SEAZ4no9NdKdCLj0D6L9F9ek9SzMmQNFjrZeW8DIj5eIzUrE0VXJmy0
Dj9K8/2szEIg7yhNJuLPcaj+5pxP7VS06sliFUTFFy4T5avf/4NEAGNvogvbtCO1
lZPVJuYk5wjXTOf3JpPnyrsfIxtzASZ4/EMr1U5fWcjhKAHnK74IgmgP1OgVkUWR
IgraRiqKAPZ+sUCcYrbXLUz707Twc+cbMpMAn0oEhbvDsDbz0tBJGiRjfMNu+3Xx
jsAs/Db81WbhGI2B+Ovo4pIUJjMwLxDwenKklmgFptkuEsxkzynXyvyKNRGSwSOD
DhYkTqXMZzSf5GBlfahaEaWY01H8JvM0M3QqN2dROq4KjEEut0KdVDErPkUuFS9M
KajSiMGXz06RhKmJZz+VF8/+PVJfQ08wX3AONwQd/smxoAXu6bAwTChhdfQ3rJ2M
gnUIhV0o2EUtn7OxmQSm1wcqDaz9vNXhjhWF1dwMXX3UypVhDx3dtBKdD+NLRX/b
IsBl10YBhJ+6aBkgpvWIK+5vvC6Gx8zBwH6koicD1p17Y2SaA2By6goBoKJP75jP
lWzBDRrVzs4FPHHUqJCO3GAUtWgagTxKSgds3L07qy6OpU4z+dPo0NSZr0WsdSoT
RPjXrESYwKKMroQQXPSy+qXZy8rkDfK9YiGjTWmg2nxYY1TH7gEvImMjNoBtzyqV
lrGOCGFXcoAjqDVHObbiJy4b6VUvuplkqEhWFFJFdRxs1Iy2KGqkYdOzJmyPx8OU
8sVFAXNRRnSaPz5OlD4gCADEUnKApED7cD8+iest0y+M9/zIhBPKTG10trY9SoQz
E3Vpq8zHWZ2De5p5n9e58RZflCZJtvLtyAF/1nw3DStL9Fl617g5LmoxuajL5U5k
1PRNlxdJMcJ7Q2Ce8ZCUjqguO0yUAfG+2A7NIIXqoGcAt1kwP3c872rZWSbOZs1d
zLu50jZFxrDV/vZt6etjvX6MA+QVkEsgbn/jwslrlMUnCrRAZsWOTbZCEK5D6vbq
R4WxIskmgFUE3kZveFDrzbdl9wb67L/GszBbgNpN4VZXDlCEr9bY2J/rFXwNjOPg
JL43EhAvXbGyomwQrlyw+veIJb5eeP5qCoXNYG6lQpECKz8zr+1N9uaSRLZyvnu0
sJ0wbtYtqQBzyraGYS7ODeOxharH5L8vKWFhxIHxhWVWhdKJWzssI1TUfgeBpijs
BqSjMi6d081XhJX/6p1gb27KiwA6h6s6qKHpgn9xThF2vhGw9rbU65NUJ5w8ka2H
ILOOClOIErJHsp0fMAdVyC0FInE9uwd3itGlbXch6+B3+9zI2dKYAOhRxetP9jpK
TJkZ8wcyLUfOsJ8ZiadSE7U43m4OZxAlw5cpHW7L1zFHKaDKB5bhp64km501E/eY
TVmEU7z28hivd+xp2d5avNeVmg14YvR5PXUzakt2tthrX0MYQ/ZkTjxSCIbC/z/z
SHXcbneH3w8d4O1AULS1RNRhEtJm8E4XOByGOrDqFUKJ5rWpquHo8GfjUAIoTT0x
qFofzyP3Nxo8u5vB9vHFcMq2FJDuSSOJEpPggx7KW23PxN8wLxESGACchvQxasv1
xHRadnRoos0xa9LgSw0EQh+MfeAiYImIYYcHi5G6klt0ukUJeGKpLAl2vMavoO5F
wOwjYXwwy1Zhxn/SPfW7X5FfLOCgh1tHaeSimkYmR5aDAJVJRBzSQvaX0cNya3G8
CabqixL8sjPjHWCQTfHmiHp9GFldFRj3pwQCrZRKgJEdXk3T+HRJXPv+fyAI1urn
cYYXOkkcJ2kv6InMY9hta2odRE/BVl0k8JzY6cYTANK3c95TH4r9baGz1ICLWe8i
kndUb0p30OgdSg31dqvtOZaiDz2Lz+XnKiw0veX1LtcdzGCiojpFbUCSwHAPdqzR
oBW9Ovdm6NuyCtam2T5i/EQZCKdEZawxxS4NJnmkFO1aDiYpqYKxv3uUCZ2hHWpR
rzDigCJQ709yEYIvQSF9K2gYOaAYESTCs3R2b9Hekn7RnqVaOInjSXZuwBjnIx2C
NzrfBiC5rzjS1O/dbVx6ycg3HlDSsTrROxsqsps5HozlyL3q9Fx5jYp/0/Fc1Whi
9eoSFsePxX8w0k59wgEhV7G43gWe+enfP6ZHMiyFM3vOwKpofWAoQwo9gIgtrMXr
exKmjMVS0T0IEmCt5y1Sd57Awvf2tH4jA2DzKHvjAKOCJrYLW/7WQShEUjSKMppA
Qrf2Nxfcs19RBEOOY06SzTD3vzcvlo4Uu/E0HlPybgIJRU7gCvesCYKybpbvTqmu
y4JyO3WjmwG6qe0gDtpNBWLGoE5Rw6aqLLIwbi1tJagGPw77u0ApWpFoGC8msTWy
y4XpoJ2KNlCr4LRYz896DAdAhTfHGxzS5cGpcSEU92bmOQ5eR5Yc+u24JPF9X68c
kiFMNc9DNznEf9hqFG1vtueGjZVTSQLxxU7P9XWuvyiRxRM5EBWGzSfdK56ZSyY+
tVRgdM/jjbcVivxWxz84Ay3c747i8u97dGT5ZKugjLK7LwCZgB5GTY7o8cA6bCSv
3WGByGECz38CZv+JotF4LNG0qmz+XY1g2alntIRwK4Ra6BZkuXMGq1zcdN9KRui5
2QOcCplOgsjoqqg+LH8iuFvzpX+t/CpHrbaIYednfYu0MhFonp4TGERI6CvcKwFn
4JWsecgjTZw572VLzjV9dRlLI3Myy3iBfa+9Sv7imEBnAzstyOFuxbVWgenYv3zs
0g6+gxJ7MTB4316LWsZTxnQc2y3/s5Ks65oG/flMNP6ucE53we/8V3KEVhwmHIpW
PQaqrYQ2O0Uo7TbSB5c4VGRutafhydlpUEHz7aJocW8sojqrvPV9uZdqauam0UQ+
bg/2oaS7THikqT5k0m7wL66DMY55QkfTVrlcLuThzQk/nnS2nz/hT+TJwJmWgxwB
911YMnrN4RhaYMpW2nBiyLoEYIh0ny5bGDMjrovmt7LMopO4efihEAdSZS7QI0lA
Wgd9TbmmEAdN/UbiKsgNL00PdvcaXPubDh6Q6J30gy09pT2YeUsJHq+GNf5hfUnA
+iUDweWx3PGXFfzAyBM8/W6v1rHtBcYKYmRDrrpxyxm0nvyPmDJbrV9c3MOvjMVl
JEw3rXeVsFwm7Q7U7ojDDVtTSm8ziy4D2QSS9nmcTTfslFpDSABCGncmPi8KqMZz
SYXFOPbBaJL8kSZ0Nmctd8EwAfpPORfcaEEzRjIVrtFbiLfVmLayfR7Bsbvy/3/Y
H3jo5jYbGktelcKp5RoSO5oqEfSjKiKnsugKzCwaDzYUsMO7eQ3k5EBmBFykr59j
rdP6OkcEjE+Jlc9H5dFgoTvT1Lxzo1f1izq4eW2i0Fa4PJFZNSLVfZUU7N7FqFIY
5k4DLq/QXj7+nTtGiGMH7OepRd97+Ft4KWUf6TmlANsuOX1MbZ5NcpMTv6nQw3Rg
nkGRjzUTL5CxnOgJn9pa11nPHZJ/XIPIF2kBML+K4Qm9yVYVNNAd3lzr7DN2vwRB
yraUpcWqE3jWu19EUEpo/diL40we+dZIN/J9tgmbiiV2y63e7iTZSYCfcKu6U3Kb
y/IzXUY2hxdVxC7cVnNiN6KrkxwMmHCwJTRs/kVqEntovTVeWdGfoGFZE2GATlgF
bxnKErU87R6znJUHL3GhL4WOK1ueFyiXshLdfa5jocpAWhATys22HxBqHgzpu0QJ
hG7ZUY4iGb3GG4O83dZBW33XIjn4F/4G/W14D1OPSyFRcUQcALP1KqxbaHadlszU
Kn0UcgahN1xQlfiGClcCxrsNoMvtB3ifZXByHVWkRWHeFbISDVsdS/eTqpv17xB3
WV9fnF7OyJx6Brq7OVJT5AuEf3skNKgmunVOn3VYW2A9oYi8hmbG40WldvvPRNbH
Yj9qNZUU5hta6KsurZvWwOOm6wE/d0lv3Y7xRjG1ATUz8DfVULAvGukG7fFjzi/X
OfUgybhzkTHXxmy8yniil74W6KTjdZnbS2TSj6DGvfQC4W72rBnKhaoP9YHUXDki
yZdtJDrNvYUJqcjqeb8NeYnpXfnApc/grwHWzpJGRX0HOqaZGGXp4Woe3gYR7VYR
oNP6nEK3JyeGbQUK2yzCDPmlbAMBPU8QhvnlKslV217xL2rqevLTg6phu15rEKfm
PXBeZbgFzL2bc8m0mNQ7cAgGOait+b+jZhdK7ybZ64+shlMeNF10O2tJUXrBZH0Z
M4gnH8kXQ1JM2U9F0Ss5m8WF8lD/CZ9IkQnN/DADWjjvrHgbk9TYu3IvBU60wLHK
JOfk7zwNQS3L/sOrz6WO5sOvCKhJN8kCqm4SSI+WT/mbEcjSx8jwJcvqG8BUMB0C
9mMPytlQnOWVn4VFJyTQUb2Eykud5D7Tt47gXYUV2QkLegbkEr6CoEEybbG3nrJx
tzlnhN9OgtS5U+C4d0691zDlI656cfKwRLqTUuQDX6Nzs5VjI0DoIycHv26vdZfw
hLFE1SH1ld4yZDXCByaSs02Zwb6PoSaq6GHmj6wZK+3zJugwm+OEJ/KAI0FS/Xyx
Z7vtvZyrbRbR8n2cWaRpOrEvAUlguTTqnRZg5pSgZtK+TwCGW5eBXdUupmpOqEO1
CVly1U2o2d0KwWcp134XK94SWrOMzKHMvuOXHvhZGmrAVVnW97TIftuXp92YzHS9
31pstjOrId4vq4a2s6X8Gl2a+l7k03dAF/oKcAc0FUmOOPUbZH6zaGfbRMD5yvLc
IMElbNdt1nlkHI0sEyeId4YrjugqoBu2LhtGVxlRHBEMsTCzgmfyRs3K3dnZLBR/
j0LPhe/CXmk4Y6iPC89h9WDUOysBaEYUL8AKwy1EwFbYiOoeE1Z+y8mrw+iN7C6C
ZRfedPxnPVKGIWdNCFRjabW5ANf0mppsPj5l3w+c0nvXeVsUb/QYi+OaTsiy2Z6H
Ie4QB1spktbXgAPjROSXycU03C4GTKlcLZ5BYelOvfyM/CjqUcS45hynLLoMW6Cw
4VIZPySaWv3YrSidyST5hGpuv/UEbgpIJftni6D/u/6NM09fmGz6dFMcYAawm9MW
pR03/7njsP7AVOT0lVJW5tNb0r0nwy2ziqB5fugc1n/bQHmmBjPEgjoB0V0Hnp+U
e6op0roFTwLI86XJ3hGZdybgNiNBlpV2czaoQDqw1g15/mYUw1yPZD5EOMyTeety
VmGacAWImcXp0AzmfN1quRHkJVvkdsmnKcR7iXnJ1jUgQf24llmDV56RYzIV9+m1
pxQJbeGkPo+2NGgU99BkoDp1+vXKJDxZQspfeEDl12jqKqvwCsxW++MQ0xBssVg6
g3P1lXOdODqMiCP+r7op1eXpmbgUvL6cUTTE3XcXVeysHnPhZp8ELWjtm/vC/hMA
tw10ez6dwL5mmFVP6/HIgxRiekICBhRtLbwjjP0oxfZdiX2J3JSuYCgDBzMQoxb/
fDT81s5Yoc/KmjgZ7o3HhZvD9+T11zfPt0t4wCM+pdCckLeL6x6yUBrHKXkWGeUs
DQNT0bsxiSahSHH5yCHJhWOGcklEwq848HW4sojjti15jCmju2snZGg+TXPI5uRs
v9ubCRURuttbT/CtP91x9SeQEEF/8FvDeFB8nD/WKLAktvFJbJnYTaU5neg1oNmP
cnlW4lBxiYw2FyXdbuV8hl+39Ep+I5TlNp9ox5t5KR/dvqZ0UMy9tTBSZ9K/64sv
JNOLL24VQKHmMlqeP9tdaYZXkfFKz+DPk//lYnocFSbD++6FeU+qlCD9JQ2S1Ewj
YWwF9/0SsNe8cFO4iStr5LoNm6foxVnc1tDCu+KIMkU1diMrxdJ6kJNIwqx52NLB
rfTAgQrmkkVlQOGsK1JZfVy8WKIh/1Ox9FX/9YSaaqd1bHPaKncFtUKeuYAzzkMs
1Jgn7xrAxGhDT4B2/RfCDP+Vv3vyYfyc554NkuejMa54ofM3dhE7OKrVDPZO8Fw9
SaJAzOJ2bCmjlWoLaHIKc6gqvp/UCBOlRNYAfSfo/h3CR7BOtl2cTyjq6l/bsFFC
HJxjhRR3NL9iukew3a1pO26IrHgE4Huawj9u2E64zOVXsvg76mXlpJ/ILbKW6DTi
wJhHcd4zS7p7WH4wWoN5gK5fVLh0Ru05Jd3eM88QWu8X92excyxNydBE8XuDFbpl
NZmTL3uFZur/tzbpsd2PwioefGKLNlIewxk3KBFDN6ZMqY09JU5Xs0QTxtF/n6Jr
JYc76Q63g7ex9TxYnbuzum8vdujM5redXXJbOSyGHCDUn9f7eLH+o/zgTpwQ5CP2
LFSlFZLaB50y/elMVqa4fV4jS6mWlZZFWRDnALb3enVzjjzAJb5zcFeX/aUFNyns
E01/eJ6dj0/PR73lPJAk+qVxF52VNSeWbN1ooPwN6hRHAQf/RZtki4pLuLouyF1n
4lBVEZ4LKoE03wCtxou5NTxz/1qoREiL7ZVKktegrnuoK78MbakQ10qFN5eh1qw0
eCnvoQjMkZMNd3h41bblGCihTRGsFxRRkm2P6DPjnbZA5qS8c5g+azPfJvOJrhrO
CLxo2osGegWw9N5sUH1Lo2Zkdj1w6ged7fcCeHt6bBa+/SnEc6a2sgZnnAsELMU7
j/DM1OsKfcBeahBj2sEdictB8EFjuKDqteypTAYi7wav882uzO0oo4x4Lj9uRzWY
+o8fk3hspfvY5Norcu+BVuyHazzG1YA6B721NN+w7sSaoSZU/EyuzT0moRE3ss2V
H+EvVGzZiyohP6ODTqBFUGHdCfoMU3F8h/4maKTeE4pkrMLbM+uixDLUofuEp1jg
7Hg0yg1TaSdjwUvH5mBHC8TjFuacLA3ij+l+s89jOcKoviBh/h/ahbrV+p/MhhNH
sw8Pxy7+OFfJCuHKCYJr57v/agL4ODfQycm0brwIo4ZtOpOGGPYu9zGdQHtbdYuj
c3Vttb3LUhyzyTVBS3I4DWcVTacd5AzAu2S6wwOv25/xyMhCBi20lpXZhMF8MsvY
w6tVGWqsPVhCZNuJNkhF/TJmjb7n12QzA+Y27wxFrWXrPPQHXj36FtUkVpklCJYp
3braiI0H08636y0NefvXYiYLkHXYoKK3vXaIrldJE9bFRaRO4xEbvMgoK0502kOp
n7HJLBXgUnnPDj3rn87DT5YPywuN1dN0aYGOi0D245iCciaVx6JKTkL+lxPOAX6w
VKkyspyw8bS6bn+fm62YOBdhg6V4J9fcVhOe4QF/q2B+2n9imolk4DgNhAQaYGLB
0MyIzmlSVEia5rrRD0JRUZXulnSSjmrpBSZe2o0Kzltf2+disMzTtGCw5EoOq01d
JBrVy21+a2FlkYtsHAkJbFNlmf0+AuccHvSS6cl9fGq61b87zOKV4W7LvS1IHijA
n9Dk27wWYBSMZJuXQ5elux+gl+QfT3WZtaekYxEnlUR/TIOPEgcJHXZfEe0XN4av
Fb/Vgg04cv0NgXUbsYUCGs7N3JSkdCWQNb69z6/ecQ7DmKPpblmVFpKK36Gna1NQ
IM/Ot6d+vx7NdvuOYqyANVXbjr/v0IrSz6SbX+Ak/L3u7lI8wBepFNLGfI7SLiyW
PdVhjaNrmoOR2QbrrsUULO/CdOM99rG0D8u2STJy5COnr+ICJFxiqUyILi1l/u+n
ODEwvMWAM/KSBUEt5grd4oAP0I1i2HoPluLSeAZeEWh5EhCSpxIAyGovzuU4WXrm
sHv/Z1RXcbIs/rOlyWv6ackGF+X5rjp6nKJgYKqD4IvStlQabdRzJUHhXC4YyATv
70bV9eMVjXMFwa4Ni0acsquhGQS+k2qlQdqMtH/Yk9LShp/Me4VWKk/Y1nV9eNrM
qoZK85/xTUNYCg1LhwfqOYAMGThjOlYvSiHTRdfV52Le6bbKRtMOGwjhtVUEuWd3
vL5+JtbPcXDB7IeqR7ud02fse8Cuv5BnDPGDDVqsjQYc3+seE7YmRLzDb9W+lc/X
EmlKuemi/zmy521GzHUodwbpFBWv7L2RtcPO5Qn5NXB63bDACFrScdsAH6C36Vfl
gLCenqG1fLUW1FtnjGQMufSvG8bHkbZSGaIur3dqY+H+JVvoW3AVOlba9r7HC3qM
moDBQxFIrpBAbgt8CUWvPlKeNOSgbcwSCCd/0cqSu8QltQQyNiXvuuuSW5/5e6/F
qQCLUPFAGQxdb/ewwIvSbz3Zch2lTpfQhUoOPccIW2tNLWSvB0Aa7mOzf2iBLAiG
x4qKBu75EuycH+/AIU5fAGryYDRdrQG7Mr2OBxjYSC35BxPqpGv+heZt8mLOkM13
a3leZ1qd1oIWvRCZN07wW6XxR24NzlQ+nCFkw+uphLbtfCsXzz7whCtbC1H0OrCV
w02TzpapCVT/oncHsjXYh1I3mgy+b/RHuUfh+8hWp6JdhJ6eij0jPSXLsnRCcoq8
2aQ/Cy6xPrn4hJOMi06sWR1VF+YPe3lIbG/jK6yntboNY6Og5BzZ3u7yS9JBnv1C
B/T6dV+ZM96H00kWnFeNs71A0URRMonZ4LL4IVWj9NKhkuPRjrmru1IkytmpWlY5
XpK6RINd2TatCQyR8fPxfXEFbC3Zc3UkHTdSMBPM/eVLattmjWAjCI7hdm6O+haJ
xBBhlTYrDnCseIKhqN4YuqjRbkoLo/R0JPqRdFssc3+EhgMn6bLyFYi+1cdbb8Ax
9iOazvHR6QAptjWnqz/Ok2n5erxQ2T6noOhr76mnTLyMLzAICNP0F1Bldh15MUEF
azwV8x/d/UqPnp7sY+jntxA/yc8Um0ie50jQSkiZmWykVzUntdNGMTDk5fq6AqAy
PGYSJv5eORzqKUbPQzHk/SRtfwupZT8AgFg87dl5tvmG2EXe1CApzHJ2rmzAenrS
Irv6u5GtTzI1Zcl4Hr9UzwBpB6XpXxgbwVZRnCYzsPFVxKzrVNec30hIilkX3JGT
tZnfY7X0qMMrHdegm1qS2Imddeiy3oXj3lgKc0uActyUwvNIvfUcIJr7gD+7RwJF
SmmYhoxlSI6X2BFB07A46kIwOdUCAXCJ+CRv6qOK2BNoTxNnHJnq7qkPWthPLzJy
PjjeHtYohQXSXwybszBmC5Ku3aEAiiFCFLNRImqZikE/VS3d6EDXnGwFBMQOwwgw
Gy+pxxBFa7OWFZzbge+UlM/QjS1DLIHKFelDMZwf9sbY1bCJITtJkaqd+Ioggp/q
+zJ0i/iqra4XgpxlWzGZ1x8hd4YUmAS0VhL3NLnSMETqIaYznXrLelCYp0/KlZyS
G+Ga4phboW8wKCNK11wHBUCSlQMVN2TwCUW341+msjo95yelYec8SW2GRiVI5xqg
W9iDHcs7gYTNM247tYxB4rvstg1cDhu+RF/iEeNUoeKB0kaClvIP2CHMtrB1IH/W
zeGkeUxjMIjhWZJlZi4ErOBw3nY8vdDe0PFoxavvXGoD03hBAyq3gXFn/IXltOwE
0ANTeZlrQOczituP/C6CvdgJg3/gkEQpGvqZn15ZuACmpulOmkhCXGwYULh8rCWy
8/YoAR4zrxIoAKaZ3rd+MOrsnFq0ovNimQmeYOtJWLkdtJNaxzGiBgC3iFA7TN0L
SBk/FuwNHGj7zMPQT+ghDJioHHPHfgz7IHgUBlJe2691dv4UKY4hU8I7MQTlqIDS
sc1bHlXGytBy/3qiNLWRL1S1yEa9GWoGqxWqFC2gSgJYPl4C9Z4IbmoRJBf3otSk
C5gL0/+vKgJdwktISakQwDF7MdNfuQ9g8lHk7RtMnfslQs5gU/r+FRbFpmQ0MJXg
wCLV/7ucB37pu/7n0hgRIcq5UAjn2p/FA1Ncd4QFUCxqjrocQNGNfy61mf4umv9R
o0C+tA6QSe5ow0vUqZAlNr817tT4V3k/r6PpZJyJ1Zt+kdOhkakSeN/k0FHUWWnL
/nAymz8xgEXfFUyRS/WF9tiJKrXUbhKCP2h5ZQIoaRGvUAs5vCFyh43d30z0rCEF
nUPxlEd16CmHjJi5AeuJE2dHI0YN4MQoEj/LTS1ALQo+N3j7CRQWzWXNbZCWLyMh
+UMa0qUJlKHTec3YQqJXx9b1JT4iWV8ppkz/0UvF+JQsOdHnZIPwpWNAbV7nteSu
ddKATZghRlTxFo1JhwM0QzI+qBD/uTMmU60k3xRVVKgI1vhSLmvTWl0SF0rMmoZ6
HuKabQOwnM/GfeI9OLegMlw8hw/KSs38C0czq1B7deef/EyQl+QU7nbsybErE+vG
YmsxqBa0yfQ/2THb/gIXrvK+G+XulOMy9xn6LsEsojKBe5uW4qvvYgWBPLFTmlkL
PlhiKGdQavOKuU4gakQdzW/2a2m7z2gmbgF2nR1cUfyRAlwOR50abYc/xZA/QoLB
7vBWyKLuWA55+Sl4iwoDx7fdDr6LrxwCcg+wm2ibV1CP0obSGUtayu1Djjs+G1bl
XrQoPWXOPiXvpLF+o+Qu0/x3P9lRMG5+kpFtAkBPa0v+PrjZ0kZWNwBIsz5ME8VI
CKXfa/UReZtAAvSwddAEW26sRzaP4kvzURFiwBmQjD9zVj/mlA/fNm52I579zKEQ
2GrsLbFFAqLbYuEb8zCXS7DM+OGkb08JoKcvdrq29MSc/XmjxgJkGgvFknHKyehn
EE82DneicNEA78EZ2yUC6vlumozjkApW7xs/b9d94AdES3+5wYBxMrrc1g65YLbk
buFCBot1shaJJHNEcGWHNHl4sYH5K+I+h1HLVoAN4qaqTMgZgX2jVe3Iqu3DECVL
OkUBA7kvtKsQ7Ije746gaLuLg2fkWIMHnt2s26GMA9UHEltGsoPWq/H0L8pIIbKE
RfLhS7/kP8SgcxndErHx4zOShGt6H4cGo7L/CUoHu0X/zrsHc6K5ojrbtL4fF21z
p9YmrLu+WxEsTAE2ebhKMxoLGnqAew6CMV/uncJADxTjacfK+Ah7s/fhJhzbZNfE
buRVqE37m1jjAEVS5X0b44mYV06FkYKFju/jRsQxPJOEudGiMLYRUdZYrhrS3X48
yCwVwI6HYcnnEqe32/GIwmGR4kfhzcytdT9MV9Q/Cmht88Jce97a2ubdt8rsU/xu
4FQbGxRGcErHDjAvATaouMdhJTcMxpiTSZNxpEARQaRNzDom4I3MTnjXcRFM6QvO
tSy0V8GCuJM97nofb97ZPuYCOW+JOZhTCnIc5JqMQ6Fn3DlKtL0sV3KLVV8Mq2DK
KVPeEJ92ZRR1ovDkf0tQyT9E16xHEUtk1nJlZFtCbhFYDx3NxzZy5ONJPbFv//YA
/6dOYtlJmTElGzJ1vBdGZL/Z/rH1bWHCmtPh9Romz18E0XAuXZN380mERmZomOik
cMD6RRdv4d58VKo4JzGPcaVSQ0ohH8MfuUdyu3HWtuyO6/PK1PuuJ8FwUwC0ZEyS
aLkas/rG+1ZgWe3Jn2G5cEWwu5AvrmWIFa238jVniiCQuF0XqEsx14yLebG7DdIZ
YFoHQjOeD6+/Y4WAhgUGLKx+/pVIuI+isHgCuQcHbqmLSFUVg/eIaT6ot+8g9j/d
G7XXbzDX+kksq19guPMLzESB5j7HbbtlVsRleOo9Za+0AB1P2mAgM7WwZ8ENy440
rvIHF+2FE5M8qny+X8HECudk/hxrhSGo3uRHIv54HIBzbh6cvVv3lKth5qxl9+GW
hdxwxGCsQwWYFVvGaYs5YjTW4nxjV2PJOBW+HAy3lC6nKxqBP2Z4NTadtOMrfSTF
kkyvG8dawj2STkvZET9jVNEACPEIIUwHlDxlhEZg+3/RpnRsEKMX96dQHKOX0TS/
UkM2Ted2hf7x2PemWAfXDFnuyQNB9otKZFEXi6P7q77GQtEOCMkQ+0dXDwQ5YEhZ
dOi2VYAH9wiZc7Z3xTWAfXR3WUL20Er/WHUafqg9v72v2YQiVSEM68H6Zmh9EhYG
UgJeEKQ33eJ5kBahDZLo6kWXwLycRAo0L+7HW7vKnilxK19W4P3qDWTP+SJv3n1V
sr3D6MFKdv45EbW703WficvTDTYkH/RAcoSHNr23RPulsOihke1h5dg0sGol/+Yl
9Ki8VrfTebXetVfAh/A9NrFTFLz+d42UBG+vCghHx/azmtnS+i41KsqfgYBGSJa3
GVx+dxwcURnplHf8n2MH5D1AvDQYrFue71/1gEdCCWMSK4CJaZj+lYvoEnv55qMi
L/pr/u8GrnvYAXGj2jhxjJhN5jbsQ2sKe34QlWXeucpm0gBb3uiYNQ1lbYKbv9CA
3qrWGamCofBD9ifdePNsiCZhRyUekgHE6ggj3hpRPHmMfdBuWgGC3GiBw+EhHch6
5IymuVfJu6/CWUS7+mOQHjQbsvYDPz8Rm/a5FUOKemRvNWmUsIV6RrzcAq7xVmb7
ZexrIJ9WYkiQzBZUtVPptPY33W1Rf4xGgDzmvekvpo++SXDSvWEDLup7AUBq3N9m
5G41VrOhSuMcRC1aG2YaAc1xqpL57bvOHUQQoC5Mpj1yBshjJG1kGXa9bTdLWT6H
IRjW9quTkAkvvexKXdvaXVgsO+NhL+dAkb6zc5PxblgbVgyDnAOeoyXCX3aNWXdd
IslP3ETqBbPNuKbL6TbBDfJ/4E4vmcnSAvrxjME2bnzs0u6iy0cPvsQpLhEnKzaa
Oz1QZdbaYp71CK8RhbGh+G4zFkVwGvhv3Qr4pqgRbFXDrZb+1b9kP6cbURQlS/t9
vT8ZLsFhd1Z05n3iH6DEH0iXN9pbeR969XxAzr4W/ighPgI6xGgx3VIjBWksgnIm
VbwzyzbNcCjWVY4LUv1FfEc+ayEFlIDK5uuY5/gxludmpgbTEytDTKMjefreCyw9
iS3pvtD38GSHmGr+WdHvc1xn3LHhrxj6Z8F7+pBiZw4jYIwiGYxBoKQHS9KlG78f
D0xP3U1jNxlfcQ3yqXtc8HPsX+9BEzSeBPx8gjrVspZ7PoQ4mm+Xa9z+qECmUOiH
vHEfaeJw45cHIST3/BSAiYdsRnzW7e6feVlY7Bc8BrhUeOzCdhCNdhwu4f9gX8FV
/KP1PJ68TW/2laBaHaY14FQjxTtl3qS31Wzt6XP89XfX8+CTNrVPDKmOy5TTSls/
HXnP0Kxoj/vZYhL9X3U/u2fgLhM2qf+HERRLNMYu+tYJhwD2g5h8ip1oYtsxVJof
qfESme+QH4xkE4me7IeTbKq8ESqJ38XRx3oGiYim3S0rUCjpLECCEyI+u3bDhFC7
K1P9ur4CW2JHeefSciTAGOSgv99jmG6+oGF3jVVsELFf6nHURB9ETp54oLZ6FfTI
NocIiHkjk3ApKQgJOOI55aGY8LhG5wI9kxJCUcKtS+kd7MEVVAs+SF11R6oX272x
MlL+5PrfYIH20XoPcJAT169cmqe2lpbSkklXGQiJ4b3Ahgv7useqlDkM8V0AcWC6
lEIRZYFdfjD1axlGK7v8W6nYlnYDV+hbiYd54u/AKCeFRI6rQ7IakPVl+VLxC77C
WMPBLsnWY7A4RB17b5H/WTVI++zZ4lNU5VPL5K3ayTF5q6YeHNdnKMj4NUktNli8
hpzH7E+HKara/I+sX6EYzMlx3jF2zQWeCFm3PLONwuNFaQzR5gLN+KAh1B88mkDG
nCCgvZpIzScHV+wqdphov+F/jhbUHKUXDIlzqE4rWM9jLXHiU9lngIg3Csq5Dkka
9gOTF7l0aSbX+uGTAY97fhQ5tillk1Cbn30NSIRKKHLEtvABqWU7cOuOV54d5ss0
tlbo5i5KdMaeXCezDbNEQbJ1r3tG6klMJhdtzOzEdMFY0yTZVSFIEUFOslT6yXlI
zmtxyF8Ps/dVXH/W1MlDAlBr+nfpkdYnq395QafJBq8pcvY+fZXNLM0Ywn0Wl3Eq
XErOZi8OnYonmKyFErTiREg8Pjgv/HSTJkORIcavH2L+b+oeSPQF5ZEKW+DaO2cq
4Q7M3a1ShseTpqZVzCEOk9uBLpHY6gR7gL5+W6/nlIvJsL9t83u/UUKunKp7kGyL
x4aj9qMWf2FLWz9+Ff6mUOsPYAuqK0brMjrBgTSOPgFfML/Vo11XzQZMqR9M1Jkg
dIXT2l7ndGBxLFajBQvL6IC++yrueM+fm//vycBPh6YPDX7ZYhSo1kKSHMIBu7Zu
R7UU6OrFCupFyVYa4FOGdODEMZHxnvIQmByAoX9zDnnGAQzW9GSt0wCkWNCo9j9A
e0P5pEUh2ojilSXRSVqCufuXOafF8h0WigbseZEBUz+hSDuqlcTAdzHfwtizKIHj
+o/FlMsgziiptqIHlJiwXFglyHWcQKUL80aVw3ls9xaw5BFunHoawCBHYSXlOqHX
saoUiGmx84dBPC38q2BDxceQV4TZ68v6nurz6Xl+4bE5vPd2JKxitOg5yM8IJGMB
Io3W3iiilc2mHKUi1leSTym9ymgSB2Yj32bbMwyS5dGDwE0Qf1jqxTWscm9/nfka
yXFtY7Q/EWKMhitcTeZowx1uFdhRnixd7iVDbTO5Dix2mKVCbHGraNUhjlz3L83Y
hnG7s1YKMQxQdsSpwzr+6DoC1l5DM+2WBYdcqBiBW5i4ZvJ726lxK/royAs3xbIw
q0ldg7G5P8ktvYsQ4p3HjUaULEH5L5hwlvnDgAJbZELIvhW1kENr5lo0/XENyL6L
BMDpGopirQ6x6LWQ6e93xocvetM9jEqjR6xBdUq/JNw2mCCn6MD7lHbRC4fBkDbM
gzHZTse1qe0geCpp1/9+pHMKOlMbigVdmIvNLbvTigXG6lwFuhAbzpQUo2NDdzoC
0Yy8CkNa3e0/HTAlm7vuIl5ixxoUszgREnzGLvjNn0nbkcnDB8oFYgqDnA0Rr+uc
q66FU0NYZkRaotN2CmQwaSxJopY13/S7KgIoc5WCCCRlOTHFyrqJKfNP/GPAYAeI
mJuQjanG6l9qBNII8wNqQEAuDkHvMAEgwKYDyIjn82Z09QR8lkKKGS24oGgafIfL
15OOs9uyTiZ51y4QqalnOdILiweqyYvKR1wpnqd/0/LmWfZDjK+NJ/Dp7qjaXSf+
VAMBJwd+ncytGy1DmV4BoqbqLP3xByZB3TuGsalOpxPnld3SaK0nfq6bksUu5Tk0
mf75iSD5TNs6wmkW9tXWJHMwH+YdQVxWmKNryfcl3+iAm0fMUP9GiRSi+xgQfrJ7
/m1nJopAxSFVuybQZ16QWa1xCqpaB2VsYee1qKREQ6ymkYRZyzAL2jjkkcWoXbvE
vLkgvviSCFUQAyaGZNwWlZnqRfeIyTzgRDZbQspM4Vq43ONkBUCI2p0KgrKcvM2k
g5dBfL0ojoT8ivGpOkYqo7GfwQ+SC+EHx7ofi9U19dfzzgYrdOZv9cIuKgSnycb5
nS/wS+NjDtK0XCdOfB3jVrPYs5/y41PmHIktK6NeeVKju60gQsqSUyFz9Q4T69C+
YNtWzDtCisNpTmgiZDm67f9SIEi2wFH0jO/JHNiB45k/BMuodoKnTREVx0DlzCuB
Dfz3Y1ZWiPlJbsZfHQQHV2Irymx3FZS2nuZisuDHMw0eHMkZ/p5z9jDEOxwXb2ML
hFGfh5sfkc0nfO3CxoGG4QMX5gKfbXEIrdrXPo+y89ukRpNdoMEAlYa5/uh6qiSP
ZTeN5rvOISAbMfX++/N1fHMTk9I5CtlYSgaDfNcJFAVrGFkZVonrZR2YqXiioQ1F
6uqR+fg5GZ5wlKi3xixqvwve8ElIRK4GjtMZsB0cnxj71jmTH/Ttog3nAS0AOs2r
Kgd7TE17J+p1rmOtzDHb54zd0vCR4OWRizFwSZVNrXaaKgSZGuH0/XiojKMRd6cc
7r8NCtfXHzr+ArMWYWDMAaifJSx0rZqGRDXVMHwBj7K+rkiyA6KbJ8QDZdg4LDfi
p+TE2PmjLVq8x7GgwekZx24KtlamcoaQ5jjpYlqEv61F3qNLm2/yWVixENfhdsLw
FvQRDsI+CYcWoRr1nBFYhlQhAcnOHWMpXxYnk+0S8q0s9H2hZ76t2WY7GoR/C3TI
D5IAIt1+sUJ+HJc5wjwIQSXC3EUtX0TbF4Kz3Uiio6zp7CANJzBkR4TTwBydHQA+
zb2ZdS0CbThUy4yD0sbURoM37dYhhQm+2/yPHt/TTj1dDw4tGRakSJqzJONqkERK
xTLlYfZ4iWHZcn8XXjr6ZndrnGBz+SO6oEETrNSb1uMNvvg8nlyHiHJcL8zQhhIN
/6pIZ3X6hfDSytEY5dx/GtCICAj87ZmwwKK2/MwyjyxKrYoDjBp+V9ryPhJNvjH0
2Of+ZB/1B59Xs2GD/n9exd8t6qtb0vVJqYDuQTKi6dBG54Bj3UscGucoLcTJ9iSD
9PvzKuLiQW4hkf8DkTy6vDivMhgt8lex5Euj4GW6Bu2jL0dtPlJDJ1G/wfR28uuy
ww8uDUp1gcMGQDwfT8EU0KPZSdJar/+vCrjXqqJP1vDyMHReGDDZXd1Z1lt6Ovbh
sSyKga7LNgrbsSXudOudQZBbYEsy5plBOUajcL053Om07mLF3nYRiGNFTagijhL6
RCWLA57/rKsNS7wm8p1Mjd7eeT/MwUNE4+calg8P+TiHmadcqcX+tYyh0CMDc5zL
3OnpGbkTgJN6mCqeVdFmMV8V5kVix7ttMwrOKkum07fqVQcLMSWTHmpHlEq6LDwW
XbiyadSznbhfa97gvFhOF+ay1G/Ng7QlNDSL+WHQW05L4GZtmm97k2wozjN4oxKf
sH1ronBRtAPCDynsex78uxqsPEfXrhjrXpbcD9d2LWtmCrvHULhfAVdty7ZjAZX2
8pF8nz+p2hTbUQYNIIxYCiWAdoRtPkq/61cwsSY7szBRg84IeDGk5CsNCzaavRcy
kPK3QU+YlMpOsr1JNqjo/THuCmGPlhMidrUJeIEAd/3vgD3eUSmwF5U7EUXEiT+P
FoQ79qvZzyBmXllNiMBtn/zzqau9sJr6LJMx2RdX1rWUciuyvKr73MMeMpOAzJbb
wjylavwqRZcneuh8nTQc4k5LsjNIof3Y+eJU3Jr56PHAGXJdWkFup5Gxl7ph0Fg/
vXnA3DP0/nkU/LRL2HM/JklALsKNVlpGhPzC3DItkeNGGR2upYSllJocZKffU+Oq
wVJm8OSlIyVnnL+GixUjSf/kfwaQHx2IyMHEj40GMrVf0SdOH+eaXcsFtHesfBo9
4TRb/41Xg4rEaquBJ++qZyjJf4HVWEu4ZQNQaQQLz6ekBj3oXgVn37Kaxjmb9aur
3r9DqdQA5sK6B9ST4PgJP2+QF4gM61TgWTC1KrAp+/G5paP0IEhxBmWpzfQkgbtK
nmchDgRPE9f1aS2ypBsHlIgE7X4+Y5Xo4MI0uMtsQQL6hNFUHZXsji5/Fov9KV7T
kF3Mo5AUBa/PBBWUuLVW6wAc/ubSnmq1kuu7Zg6K3R6ApMp69hhHe7M8v18dPDWj
tkMebp/0uRmmOZw9nCK5fDD01a53aaTTGde89Pn01jDsP5jUbjGAElWtoZ8kvNv8
e/YdelautqPnNrhBMjeDqYfjjwBNgd0WME6PTon4LQr/eakb6mnC9y/iSMfNFs/2
Q75P9CU2mbFIERvRJ5HAgKWWYyqfyC32SKlud/iUKaZJgccX3nWSa+K1VwiHZv1V
5hdQKmkIZn7VHbsqz3D/HUYauH5+qQhJC4RbUPZrOYKxB/U2WXahMENV05eXbwvX
himpPmVjL7Itw9oxuE4zueDRPd8s7QgcDzF7Z9xYb4a1So+YhOJywvzRS2INFg7W
xfWX1efyZ2JT0oui62NqRvM22Nn7wsfmtPDev4GhXmYx/Zgpu7b8SNh+xqrDYFHf
vpSeXmCjiT28QkJPZoEMNELQ72ktplJG1rr9rl4RdU0Mgt6B+TwtT0rIlvADB+dS
j6/wbJUV9GHb5lR1rDpKMk3ghwOH7tdLPQ88kv8Jri5ZPlCu3z2p+YHvfaPtl7of
WgQA+xVcSCyeV0t7QBz+Lk6sXgkAyHKWpIr+uJw7wmt3QGtmj2BiqFji+IOAZ1Zo
rPrXnpZ162Nq3cZuIXtS9Jp41lemlKUW41FJwX7FEeYlZJ49ec6xAVwsVwez1xb8
zWXQgQWjotA6I80HkoP0I8JOr5LDEh22kzMZ2guOcgrg/wIbCh1qTvp/rBI/MLao
QOPqbqyp7EjsPY9C/jus/UI0jS9fdExmPWvzCrcHOnYznJzWQrwaxIBI1n41T6ud
a+/HMPvFqnUfPBktzLevRJoqGE5/NBpXpHrS9XS4ivln82qVqKYBKnS4chSEOg+2
IoI5XgS1Q+1W0zZz9ksxvZdsx9vvYox3G3pY1b/BGBRPmoFRs5JZF/fEZS1Pi5+Y
jrqr7hTNrBFJdfSiGgY5wTZ4i/GjZ42lwdTtJ261naCi6qFelwv7mB0rV5W+kQdb
GqpMpXn6M4jEsRrq7tKzJNf2B/Wq5B3JIRrNl9ST8FQKK1XVD6Jcckm4yqYRKr/5
cJzptiDeI6VlX6R3Q4W6Qu8lcF7OZKCf3jDFRjr6LE7bE/Z0NH43bKzM7L1UnigX
StxF2PvRzUthe32u0epJe50xgSZutZVDSBMMJBogmSpeGZRIw8iEwQAvYRAmYceA
OqYJqiThIiVP6sGlB5rkG9+aakXbqifuR99lTui5VW0Q24Ch/ZPQioShIDrOHWlP
Bctpfc36L1Lfv8AS8HMQLD7srLYDbYBhToLZSO5onrRtZyC6esZ15Sujxx+j/lfJ
Qi/JOB/FHuYO/vTd7tDtwtR03unf5kIIAZ7BVP004QhgZhbhDAlXPkvx7mZkEvtR
/KvaQpGvimQ7cnwGgjzxZkQOyV6IuKKwt2GbZbiLXKIQVlzI515ZiIBEp/6phNrU
MUiCgrKOoXUTf5qhmzvOABJYW31C00uq/78OAbWha6pVWb2ccAm+xk3k1JEM7MYb
w9fqgNDya8rsYE+0p6loiuXAEjBYH+XcoUi7gCx2aXg2kwkxfZMCh716WTsK7BTx
dHtupMNgVWlvDUgjBG+TKzA5F7iaIWVOpFYl2bvHg+c0XUH8arfG3dY3rwnWqHAj
i34NbN7jGvw3NVYo4wL/r08BTlz0EvHrOB3X4ol95zMILdYnCcQ/bSLGhVrQimRA
BCQBILVUPgPxZPth5udcdbYlw4fWpeMHr3XwA/JewDIpnjZWOeZJtSVab7hgEJHO
mx+oGTW1nVL3idEjf5JHuhwQ+6RVy7kItrxglURiOK2D6VaaDUOXsxcAsF31J1b5
gFWuGODEXgtGHbi/Z5tSLfg/dT0SHUHuwg27lQeha6nR7UkLB8xx2cGljskkI6rd
+6rKUnpyb76bSi9NH6jm4/S95+cDqpxYfKbJQvw6Y7bWRirzNObLV/2GxBBsqW6W
pwPEoUxdG5jXPtdoPsHXsAcckKDKdKq6a+64Nfzou7hZen5uSJJY0fTTKkSETr2P
L8+qcLpGflyjX+lljabs9b54HbyqOyuzWjoVALeTh5Sifg0uc73oY+Y5piES7pQU
klsuBLSstJ7YE1/Zv+uRVHQj7Ny0107qDfkuBCaIhAEzQMGhIDJdoHpvVVHnMaNP
shvfbgrkmQi68ot5yv++sSYhQ2llDjRCqwrHxZVZrZbGA2JiZo+nUr9C8YeZoiOG
BgDmindvmkoe7kIvpd5ZK2G7HglfGk2Oq+IhiWPJC8x2pSDhXv6ejh9533+m0thD
P5TkXlICJcqBRCybR5K6Rt9LhkYRUBRhzkIsHVBT12aKo5U8+PmAszJBDf9VaDzi
TQVTzOdgsu+VZoTUB3L4FCWViJEPj9L14PXxAxdMACakDjGmoxUedCmwYfq0Gjm0
APi6RKCOF3dV2PwdL3OIV54DPiOR/Q0nvLWVB/3EMMZz26XpkqFD3LXtpLJVbFfp
SpkE6IicrRY7PTYdrnFPCk5Pf7gBiTvUBsFSX79eTxG5tl2+AiuqfoFuuXmKMRs2
5i4mpUSFTm8MCByczroScAnLTNb4GGOBfyrTekCpwc+KfTGU4W3NAl7W/FPvorqZ
mK9x8By3gKa9bU4Tt/8Kz02rVkz0xgr89KF7Dr5aLvqFyrb1ywSjawYvkwLw46nF
VXdZMvXAJIiyqztb8fOk9l9ElWS6jyo3byjoezOjVu7p9tdJPof9FDC4IhOh/uPa
VWCSgX7K1mJfxETprZDqwZQOlzNHrVhq5IRasab/vkjuREJ2GziL3c9cyazaHV+n
oiFZ8xBPICjeK1sIhy5EN/mtjbGpBcG6NPFXnIszea6f4Y50tVG6OgYiaIwV3YuP
rNw8b3BJCzpBnztZIdKon10RZXq99Tv4vJlKYhXx/7gw/sD+6+mYOS8VlvgeTdGM
H4YDCYsDU9U6q6V0UnBPALLY2Mkd7PoQbIt/BdWiDwqQtLv1jbRLttFKWeksZFPj
jHDp+zkDqX8K2OhZTzBezGONIXJyDGiUQ8dG0x3e05jZY/yyFODlJJ4jfu/56bEe
hW6Q//y1guoF2FqI8Nm8MXS5QKyBicx+NGPYHLtxEvAJdYw0rgQR8Zodxdp0pe6C
qPvYwrmR3XUaQq2qqFaY5IU6DgIwo5oLdgV35HPJjdTdsozNerexRL/OyRBD595r
Ub3QJc7iBx8XXt6N87KNGDgCM3bG2qJLnduI59TgRsQribBvrWLEVnQ2XUHWPoF8
hwy2vBWxE+k5r5XvIYlZ3VbdYlRm+xS5h/AMGdXyQFhMWEmlocqgK7viKUjb1PQT
jL/FUas3v4sZmFmm2tB9rNDkTVp/eO+l+rDLC+73JhdzLJ/5l8NbL/Cq5/oWTKLm
dGi3Y2t/TqWQbfhwroX0ukS3HN3X52Ma+sPfZFgtmtOKF0v/1kRWPqkZAaFrwrRA
XpGxrlkI4BTa9YZUB3F+z9fE50ZtEixkx2hndzEVYynvP1u8K2+9FvBBlpCM3S9B
B8rXfgR8xoYihJASP7g6r+O5ZHtUmZWk4DHrWGXpGh2dRHRuotnpWH//3ntOcsTP
4YuSW5ghz3Qy04xvc4e5MMBk2P2YRf8s4V+OskWxeL/4IjoTLsLFeJoar6wk2qSh
4QzRswl6Uo7aTOWKOVpA8B2xQdPDrJnmO9dlhNLbiIkkiBuzBmaSeoE2EolsawYf
SUABpjtMNHbyYW8DEq+QDtBtUzh6UUD8QEJAuq/YrvH87jBgskigQmbLHczb/MHV
so62W4eGjwuGAdd7lJAilXLrZW55E7VkPo8GbXQRLlp6t5mssN0ykXyUql+UATKB
M0veft4EZArQFNpuLNa1ejq2tzyVHtWlXls/M3nTwDXjnZHx6xVgPDjzVr8vJr7s
NKXnluv+ogRRLvJ6qj8Ar92qxr9lfSTdRE6QkRFDaYIJM6iP8N1kIu6IMVFZ9ShF
NKFu/HiUe8a2/xHVAgx0hHmOqKjJPg4YuuKkFGSKqQEHq0Dqu2eQUIcM6J2NN/N0
PjtTiAhuwE67HAOp+TNmKcrOF7ZPh0mSzt9f3cS0ePjBkTLq5yiT99gpNgrvjki9
LkPXioqOGTjbgbliFwJ9wttnQd0smyYo3APaCS4mxyWwNxkePEu7DfGanAafA98D
n1zGbq/umQ0mazfx8HMnALS1TbXjH+rc9GWu4rIwEFHcEE57bSvSyZ40AYhHPQCU
FGcqcQ45Fn3l1FihEkunNJ2SkQE2Q8Xyl9PZVfIFtzIlFZ6mn0QQckw6RHrAdRM+
laLjGvZwpWA+yWIurUhDvizWVT/pIlKyMOMU3p7IoT2me+ck//1dmuKsAv10HbYn
B6NXJWGpIrhJr/BZFMJVZ1i2L9zCJJvSUeyxJpefDbhPHdT6Tx3+UhvSMXdLqfWo
eQZp0nL7pMmXhaKTUvA8tSf36Bs0InlaY7GBlCpHy1kiKoqBYS2LCoHCsb+Uy8i9
vGfAcpTYQweF5pFs4IEBNiw53hbhDGoI1qmz9eZQzc0Ez5LF/aNI/4AT9k8QCj/b
rU2Da8DrTX30dOhbyAOrHbg4GqDHBnqUGWicFgsMQT4AWwVR088GDME6e/7D5Ubz
TVFhBJwaRa9LqZAPrzEHlc8ImqJ1xmQ3EkMf9dnpyevlOV+no/cIvyZmAnU8A0oq
bGtXp21vIDrfFO+vgcNh45vfbCBn1Ux8oUjSBBUaSsZlPpkpzh7VjZr+naigi8AW
kDI+cVI4VL82B98VkUX9r7idCWONMVHh6rhogqo5Dia/SvOIsN65Uv6EnZ4lxENN
GPqygL9ARhFyLXIZNfBcA9JLBIs0xzXSnRTegWr1dnQc19+oLrCEhCkMZ9Gf8itC
/U1pnqTWrxxp3m5AXjehCdJjdQytAdM8xXLRou+7wCgT+W0WA/p+I4WO6U5xUYtD
WvUR2XZV2YSeSuXZaMhXbFag593bTHoTuBJCtvZkUA3AYPGa2VvVM8MmOTom2yBC
EN4jw6eYa7qHN8q72qMsbiVxa6d940vix3rui+cnhLKmebFG+fQYAu3xQp0u5hS2
EuoEx4h/97HrhBZ2Y6dIo+C/Rgc9qaPwyOHjj+qpInTqDZ1jhDnf1NSpCaQIAk/i
DmlSE590V/Dhk7yl8+THUirix5NyNcq3fXMcABKB0osuo1J+bSa8dwPwAmz7Qo9X
5kTjLLOA9UzcTMI+AkWsxxH0NIdQeDks054C5y072zQvArUnB8fpgDQWAlL7cGld
Cgge8yXGF77oQSYZsrwenNCfiU5xWzM6vMFmY4FIc1T/NyBLD104C233+dOxijVl
yt2LF6NRUewinK8XHMgkMcYmmIFRML97PgvZ1cxwimeJ8TQq9XvzcYcbkq6ijaJ8
rmCi5SJydhzpoRENQ7xNPkpz9dOtOKHLb3nF/LiFz8UJxxLjRy1KN4sgPOIJsS8G
NxQOb2Aq8uB19mXI5Uqrra/7/ZAuAmGxBh5qmcG5oNGCYkKh5kGnc+SKCU4QNyIV
mnbtNVl+Gafmqy+k3CwZwuhBNDVxzBxMl54+1t1eO9RwQznyMfyyVDGYak680h/K
L+chHEKlz6QtTJYt5pjfGukGd9rCi6/taBm2SwpSUFBYO4PatuEbawdrcPEjLpP5
x9TJglDSCbPNO95qXFtUi5ZnyC7iulW8c7N2nb5euBFGmo2RPfWvFhBNTXvDqWpX
N7cRFAJPb3MRkRHbz33p7Bv9ncet/MzTda2f8ip3bVE/7d3kkiXleEb5vEd9qY8o
U/D6Zh6/8hkWACsvvkSQb00+zfl5gxfi+LOYJjI5g6Vdfpa9nsDZS70+T8X8Rip+
jMtjgN566drOV7+TTte0saAHreB9hmt3bqC8+RQwYfIUHNhgadIjAq5FaG8xpsFP
ur3HnWjEj0Q4sYPfAxtrt+xPUKJbpq9ZmscoevwgNwInhegRB3PYtqd/n61Ygog1
DcabeyvEor3O8edpf4+B1P32c9CTcTDB5hzWiQ+VdpOqW6rXPRX+1KjcprA2tCi7
xrZNf6FMmZIQ9RH+WRWiJJnYEh4DCR7gLk4l9ZAusGqt4V3rx8sBLtLq/iLlmUcg
w06+ZsXureGCyy6iQCVLYAIixHhwaZolUs+bmJ9v/YMJ4QqwPY9ERZCO4ForFpvI
3/eUFr/9jNQmtKN3w4dMWJ8gSSkkxuu6xdk07E0hJMKdZuJIKzg4xuGRoyzZq+vu
PnVYnUUd6PCPVNZb6GwNN1dwHOZWbxOaqpFuwTgeAGA1o96jon2uLf7Weg+DpC0F
8IV4wxflBgVGXb1zuKxFAHOb/X+mM3YnONMGf0HDDiHymagjKlXyzjONTeuXG1uD
149sqAPJuc+WOxhaTkmaYOMVUfmWxT+5eIZmJqEtxq88FJBO39aBmOY0H/KTXe25
4gaQg3vyhw6yHnGpE3XL7d4Zd3s70/BXUn8a/jfD7L5EYAb1eZdZraLq0lGFW3pI
jD2n6ZTlcRegDntRG1TN9ePpLuFKUFBJdOvkGZnPaG3dFXJ4A3eHqjvw1wqVEMWf
2syay2h66e6gLDzmzAbUIDxWg9gc3ZOfapB9jheuWkHloU8yAUOkTh+V2KlAzjh9
uNS/IqyBdv6O6ncIL4oGCTZS/ZA17AUCasaHp8hegPaCWelaz2enG0DCVyTvFk1P
zJW4LrgLuFf8nN23doYGQwryRGiap/L6cnUqhk29FEX7tDfvucthfPlZiUtueyij
i+bFzrQeTrMLV+UYCRDq/F8lzBkjo+3aXnYIhMN4ivS9TyycXlKOishcQhlBufOt
OtJPsM1RqfZEL9U6xy7tHoRpUkYamWRrGtuIFbRNR4s9c3Qc46T8GCM/zDd6buMv
x5N80N9LnVXo3xzoaEhcvBzUiyCFXA+56ys/O72ISxQYghdEg0q+trNXj7g0YRNm
zXoBiUG/6gPETeiWOflCyowKIHt77K7Ky78Rjxify+VrIsW/weDVCDdHKpf37Aoa
0TvzTYaPa0i9BcPjGMLemoddms8PU+CzpFrHTJAGSJ1wo7aejA3deRMzF2s+R/JN
ilLKm8/ZIMk6C87t1+GgqVNhBg0dTjFhIzf6+Gsp9K6v0+CTzz4lQw2rotRiAprC
QYtNdpSc6M0CSpDOd6Xv8qF49Hl6Ae5kcVQnPen3xNHH6/RVoQQcN8IqHoS7AY4d
wo5eq0wJhoKEnZuxb0ZSi3luieSrgobaei2hOHKLiWsjbkpTyazYcUu6tbRViAxY
J/EpwsKXm3FvMn6oRrHbCuOqWdUXOe1FYb7j5dGn2K5YeFPdhUs0EcuHMJ3n816L
NifgvqKbM5Y3HUgxGyq0ZrewBXMfbGGPfM4u2nSOMsn9yr4iCWNPn34s0ePhQ8VM
+wocHBSzatO932oBss4hsAXFgaoJZcF5/fNZb1BJ8HzS0ROMA85Oe3gexM5Qq+Lp
uTtRfagq/zbAvjbGpqEr4hER2nC/0ffzoN7SUCQt/nCbAJ2r8JK2V+wYzeH6Tc0H
Jj1z4kB9+1nvVsqawIEY7fyYOKHoomaTJX/9qByiFWSPPLw1uRYtqsCKuGyTXQev
NiQVGLb5jw+rhBcdPbmUCPIzsev46Pa/Km9jGJUg5tPyZvRX2K1PzMSnoPkvNQQs
bz1h/sOSfiQUpo1l+fkcmfhZY//f1v5PJsF3H1cOcmKndnVQyoUF1I5SYj74n7tW
nKU0isz5Yim4guezjEFV7TrCMxemfmPUFeRMyE8qLSPqqasCUS9GzyQgOXMfXMon
YjHdSUsMgPEwc+ysqTcnZEdui/Df/ABtuMGkCyHKaXiwZcqjFXKO31MyLKRyJ9kE
7qqmALiUxHk3yIrMI5U0wsyTLjI77G0Wg60xryZ/lAcME5B6EyJHN6zjdk8kClGH
b7AhyyOTgQpEaMBvW7hYsqCqm8nAfkK5LwzTLi43Y5VViyMpfQibZBa6kBHgcR7g
EfoAY8D7juQxdHZj65o/aDUCNKBq3koy1zdR6nR9Xa9g9+U9kOCW2kr23dLfM5OC
xX20doGXdnUVExrCfuTZQjrTxwver/ApZfSyhxY4X9ZLSaWUAxlzmPYvfINDhyD3
BL1u9DJETNoYfu+WLqOLRPEmn2f2QawcV/jNLBp8GJe3RFWpSj/oMpar6CZYAdo4
JqxPjpGqM+pQftmUBuPqzNOUx3cospF3NLOWbyor1ewKRmpp9nCE6GTd/zO2Hph5
bsOFlILpposPC2CwCFfXtGw/Q/VlLeAvRr4BRL7M6kEsGS8Uunrwcg5C+ZsT0IWg
QravYuB+TmeD7dz/n1HXaIHSUFfchigkgk/z5SepxveYKeRuaRoIKOqNVo0UEnLS
c9CJ5rv2kIO8d3OX9aEXONsc+RkzJ87aSf55R1P/c95XuyXl22OcvyEhTK+0WkRW
HK01z4yIV0jI5rMPWdB6j5GnAyYft7LTwwigcwc2jC3FVhF9XJjhxL3c4oEFmWxX
pLa0ydBEFzOTZ2wI1CIVa2HTdiSb7KUjWgPXZ5v4W3PWKzrTDHyp9IsbB7/bvqz1
rydRcGLKWWm+HLlEDbB6aamSka2cWF4Z8G0vPd3O/KTA4lbxpHfm7be/HwvTpQHV
GAYx15ZLsxZSiisaRknTJnHtWXe1czeEwinG+olYH+6XXYanCBsFvHW4t4C7X7h/
UEDOtsMVGfOhs/tD4MvYVBlAIBBOXfKdKWtNLTNXbq8I928h4EklPWENaun152TU
Uus+jM+dUsad2RFz/hH2EE4Zcbdm6yOjoEYKFaC6/f5Tkuae6HJJH4YYzT2+DMJo
DDTbQm2CGpoAPG9fKlRbehPUzzHYSG2rjqf7BRGWULP/jXwC6e4C73sv8GfQuV/8
ylGza+GkKs046Wou9LDYOcfeiHLUUpukPO4idAXBzIJGQKUw8FwTCGtbOZrYfOWm
osPrfZKm8KIQksc4dLMdd/vdX54/ZyxgM3jvSaoH3jiWJ3PnZTAMIzxHzp+mtB0P
jovzOPmzhSLJJ3R+PQ6asCip71IzWIiXrtKCMOyUtEWkzDPf0ycAVYCJi6YTceji
+PDwg/c+EFz2wTyzPjKySoEGy0Rf4aZiy0O7C+rXDQ/6tRtkw7AO+3Fg7rBF3Dor
nhTwHWRAqjafhnaB1rCzRE0yTMvnKqeVhF3cxKEdnBMjE1B+mTkQT1c6z2vSLE4H
n6lAT/L4cDGX/kzGKg/0rIzuKXb5g4X6UiqCcHhOuheHMYHn1ya76JeBAepDUubO
pJtNbbF3ncxMZxM1Q4f8tckbCC/m7OPXhZ/jsKJzOZkbyoOMWPyAOlwKCmUbG/d+
LpwA+pdjOLfeNotOTPfzmvsu8xa/woEPb53esQXs4Ek+cPflph5ZVvPplF8vqF9l
hn6Ptw1KIHZAxL5WJmBSibc7jjdOlh0Oh+y+zdhAE0+l+Ysu6YCSj0f2QyvAz/s4
Wyl+ohLXBW7ZNtXBT0gPnD0gzJjy63X6NXhT3sWN59Vzqt+2iA1PW0v0d/fYLl5K
jr3dcD2jTWOT44uppOpO3q6DHvhZp5Ul21nvqov1JvopNbIWCr7hSlEJOhPJxIl5
YHb3P9GWhiizKb2p3croNDor6h6BPDRqcBZRZudfjFxBUg+h7uImc6++TuB2SV4D
GBF35Bf5OY7z+86/voR33ypiNnBEPU+JHGM7CfWpGXWVqUBJO6Bci8kN+yPt8SE8
IrjvQTfl2of/7RoOv+4AzEBAQLGu+t5VOnR3hn4B+RHymfsyaRk5zCVRE/umyygC
1ijrKcYUzA3xhw8bNaQEZiq9XjO4nl0AeafuqEX30K9BOUtmtSPpZUAgJOsG872w
RyFoIEdV1MzO5feT4qoUyHnBXy4ue1ySPDxg7xvE1/0pD1NUcCNPqTCQ5WFdA8vw
X+dIiLdipt/MikH8BmcCyk2zd7U3NvOocs7rMISOsbOhy+pN/zjPo++X3o6lJfhb
yuu+gwwm7zB4TVw9zJKR/xxcr8lCU6bt/wIJnbE1Dq7eft47wM16vON3znsHtlab
stjz58pH+qqnio8K3q917RGpF3+YynSMiUzm4egub2msL6+INjLi27o66CYY8+FX
MSAMXvotIv3hr+v8lpB4AR5qeXbkunPcEIAQ+SNxfMqiODtwsJQa+5/PY2aPNUHP
5vZ9FZBkFLliF/cd2U983L4AXbOoS7HyqM4xObJLQ3+j6DHwOARkBfSBSmceap0B
MXrC/Pyvywo1bqVe/UBWBEM86ZhAJE/+eeSDqlKwr9uAAsOGrpuzo5K/CDWvSV4x
0jfVCm/f+ExRkYijPIt+pG8DiQe02LeazknHY8abm/5BlMDitHZhhn6AcvESZF0u
2+Eb0Pb5hrFNzc6pNvL7GO/THHufhzal4VjoxecGS4W2Z4w+aPUAJ4J1j5zxPRas
RJosaiZaoA3PNwVW6AXYatVhEu2Xtrhauqw3iRgFb3RZB/nf+gKc5U+JQNhZr+FQ
ISw6qDEq1vhqjoKVlrQ33pgImRyA5r7iC1djHjCAPKE06qvg0EclqLCnBUCouMdl
V0sHtrCMiywJ5cCw+uA5Zl1NMayYHzkWZfaitWdSaNCjEUl0xil/3oBdoZR748iV
kZhEC38kQgKrAdYPINagKM/pFZOh9adN8kRfGN++p9P9Zh4AcdnF2w0CitRt/68B
l6/a+hgWipyM1/tiZfniZBu7lCTlzhUf9o+unl9jxUB13gtmIqUsSe3vu0dk7CXs
5EceOyQDAE4q2PXrpT3Cw7GXJtVUOW94ZOAb0f5rnXRdxdrYBP+OvHWSmagVS8Nz
tToBtSIF6ok4V8JoAdad73chhuFl+8owXkjvQa31sE4Ir7SMWhSOQtUy5ey2JFTk
39RNSh8KeIIVpmC6AmFFNGoMhmY719Vtl/kVvIG99yR7d/kQMVCvN9trMWHlQFDN
AuwJvxQ6L9v050TWbIzbCUeH4kLDb2c7+h6ShYp5A5XWetZcptahNflb6CVdp2fT
CaY4xSl2tveqjdD3KMT5F2ulRJB2MI7+AQkDbarT09lOZ44ZSgwtKJfCwRqBi6F/
Pczff5s+dBhA+t95k5daVN/HIFGe5OGz3r7PdViBHAO/mER8eZMZNFfaSEY/N1hW
UAanfFwcsauVhZLnqOUQCTU5OouR0ByfwPjNfBtnfm0adHc5uJwJIJhIcmmD42Bb
agicc4DtLrWNTKZii3YRXdDQzlGIAYJqeRfEishd06TQDbhm7o1+c8FwVSQi5zdW
+YUjbRFcxWDPNINMJORizUqDQwckmncePe7P2JeYzBJBcg6CsoKFbS7RwU4OEZU3
MadeUv80fIPx2bQg3j8lUNsNfBfPszJEXEv0jO+TxMEZAsX2QWjcQm5lVo0n2R5A
182jrZKNvHTx2kJujWm5/02dkqVYLstgpi61Qtlnh2mZe53wzNvEZl4TQaGppny4
a+HZ3e2SSNQ+n5JXrjkip5uY78QR9JvXduPnwhy/Z+2RtIYpSON9TxqT7+EzLGFF
aelcHs71S7XLOP0tujbQRH7MFUm4Xpa1sBE3yQDfxKPgCUbzyJ8jj4mi0oO3DHCs
sc05dRHcuuVA5TuY97qiGOm5kq+hrJsbcGaPmgBj9smBRkLFIK1Im0AV2guLVo06
2Mp+qpKnRJQpaBp4kUKi7/q1if3U/9bspcEUsJGf7q8AL+pM2pleVgi4K/qn5W/f
fcTJKynOCMhmTCFTh4A/cPc+dzf5sglmk2tAhCY92kaqPRSsuC+pmO6+xu3NXrur
k/CBkln72MaWg9cNZLBZyoxIzcEjN/9zKYYqijds3HZA2LTWMCFVFs+xOtcQZ6qj
mpv7jtfblfy1st+SZM1RWRCeub0bU1JsJJEXIEpwrhV5QjYRDTK6ZIxJ7gePIv3g
1T9dwj//3XzZ6rsfCCoW1PU/m1ukaTy7uLHSAY9leY4gSgvRVNKjjG3R+Dl3yNUU
ynwnKW8Oj4o8g+vFIX0qFV2Kq0NXujN80OtWPpX9Uix4hDThso4sg1Cafz+suBLc
06h87/tfHo1fQxAIcbyx5PwUE4/Tayu88QhDHbJhy5OezUbeRaImDmFxaEnwuyDz
7ZRnT5M6ej7wlF8FeUvvDXmnWc31bX8l07ccc/0/WcdyJXILEAsA16+uOtHLiIV5
Z+lA4BBLF+M4wAEVfB3/IewyseS3NvplKh6Whs7uDkvEvPj/9JzAAagGCEnucNoc
nG5fFg5Pk+m2RrinrzK3jvIiKdTwD4gufHdbp1Zx0ELlRPNET9yKnG5xA+6/ezZ4
bmw82Xq5CPkSQdGcOGSAzMtgCsrXYOnZtq7rCBAJwsKj8TOdOLpF7KffHFTc3O5r
LdBlTXpaFVy8eR7IBZ5F8tQ4Yna+iVSjoWAw9MMj9R6bUUvDMfmUPGV2DFsir5cJ
3eQsb7XkVHvAfTaihKLqclfK2SoOT7mucvzSNXP3Jm9pSxa930QDNMwTtZprCvaS
LNNJMJF8NoXD8T922GHbCp/qNXKy/2+BAkxTTfll8KvCN+iOewPHcYlLBfk4XVsz
LUDZBK5Xn4l5afQ9bhRZW61KbfyFBOkTyKwWxm9xQN5yZmf89/AdCINnNtUubiWG
kA5DbGBirBolG3qM92ZHCB5y9dvI7jMbezJAZ/Yv7xSusyY4VotHzMFIv4iGRhoj
M068c8jJZ9iNfHA9F0w8sdqhSajbsCmhwnGMwVjvHFOomwJOq2v52yKk/grejmin
KJQQ8C0f0Fx77lt1G7tX/QACPk7/ov/XhVqV4dxcgstREgx+oD56vjkM2zutz1GD
+7/CQGWUdYYhWxsYUvQarK9eNIpz/caQ2UufFvECYERtCbL0GthY3JXkCurZzZoT
GrAUaMvMmdMt03dQRpy5Tw088Vq+/Kzjw+D2+iQtQw4+TUkLwPjTeaHaOsCVigpX
fJNFbacQ8d/ek2Pp50XBiU24hiaUwAbo7ysyMaAM9+5zXhV46bPz1oEOG3C7GYda
t5FjQGNWvcRKaU8iREtPix5s5Etxnq7tkEjSEX8mPBUVPfTMxVShLn24W09wq85w
SSBw/opZnKixE7obj+ToO5WlfOvQ4YcWTuLon9nEKg4F+3fZZrsUlyYgMVnfexB7
r4Ha08JNl1t5RS/HZ8QwMWSoxV5USwfp6pShdidT2ASIFJ8I1BvmUndj+9VQZrPy
2Wzyi7PImY3aVd+YSWMF3+avonJSICJO5V+ijGw0UU/p6s8SWQXM7VFXhbhvFwni
WeSHfiSUJEZ+/twytT1IG2sWxYo8ImXSs8aBgJsGSexW8WPi9/D64aMgqmoZuJEo
tfSH1TJh1/XiULnrh9rd/ocIUoOH/EgHm/Ard7JXaUtH+fkV1mvQuvVv4Z7v8uhq
wZgnKxCg7yP7ixR3l0VON5jbeAImGu+gP5pdbr2ULJi1+TL5G1a4+Y42zqWSLC/B
xH/SVTF8IrCI7soVZMYfSjAZEV1OT3Tc+d20chcF9FgLem9X0RYqqtfuzJPcKm/4
20DC5qWiX1Gb3BsTf3MaAdUuwb9MoC6EIdczMxOEeabyy+8/ML+wL8HNYVA3cQA7
cUvPSgEvUDIHolYXPBlzvjjjUPoVvRM9De72fbnnha8GluHd7/UDV1TbA8gxHdkE
rZybtPiJkeD8KUaVUJjC2EsHBPfLK/11eY1gJXJ87VCztNfx9uu5rNAqFNtYzER4
gOkXWb8xegTisPVn7/u/9TTRfW+DovuSfDauepjYOw452nvllcEYCdHgc6OhRaNY
YxxhxNQs/33qip2edRsQUNiSsxil+MvDQ8olHHAKqgqbwlnBSoMS+IST9l8nR3wK
T1wcX5uG4OPkE41zX/EdtkL5dQWyw8Hp5V0Bi77FVVcSbLnVwkZYJMkXYm3CmfSd
Bsb440KmWR8L9fQkZMSLbf48JYRB4byD5C2LDOZHsxG8FAnOFiRxk3O3vyWK0Dpq
OTbqGXfxGjq18sD+q5fP3tIUYFWOCxNWqYqmePmZLEFkgONDh2JQKqP374nvjL6V
LCWhzCe+6kpG5QW7vyTRL4wIuabNyDg7dJU+lnZrqfS/FdfJQkIz5QiVpbVXShqt
qPOPChm5Ng5eofyuQHHs13KZgvLKsUMUMqYc01zibkfqlWn/tMKAlYbMbx1suRhY
GHLQ205P9hHyw1kxyAJjM+gI33A0CiSDdc4pAO/aGrKnlGobY/lUlOPTiNZNgFbo
BqDGtUlmflwCmHtzjVRxksVYGydtZRYPK3iGD3vw61TjHaFp+3/Ykwj2hVO6XzGF
uiNob4G02W4Ax6KdxXewK1iS7YTTPwHjSpM9Jff7r8dQccY7nVRGCAYLDYWWWNPw
ka3M1TfvAQXJdUYndiBdHXeHwNDE9g6NNxTOC0B0zAeDCtFbYoeyeUj2p8hgQE12
ToJXGNkE49BKeKgq3vdeyNLT9supPaDouPAOCuX5pFJ6Fe90KKGJEExvHkP2sjCt
uEfxwK6MBgHse6ts+45ywrlYvD5KxCVOI3rKH0qYSpkOCzXabpHGi+Dn8lMjOIAA
vmy4LR3hkaEmWplPL2uGPiePmdSz6nf2LA5AKq1g0UzCLXzdyDJX0yFr6rsEbzWB
dhRZ+f29/ywByvKpjHpA3+B6E1c3euEPNlh+saYFIoDqglLmqw4WkfWX9gnaNiuR
PuwyQk9zj/L4FqOBmEMBZ3ZAum+VccC66tfOyHE7jTaZIP98ilsy3g/mo8fmXYMI
844FOcNTFlZkYymlH0i1HQZ+sgEPGbGb8J5vGBNrDlH5Lv7j/G6fGQFBYI/T6cg3
kPIum56TgBXffloIiAWjy+FMmGr57tXZJTJx3fwbdQrj8sdDdMLQ/yVu66kgc6Mt
guTsn4jWJrpbwjcYHM7kjNKl7FwWtCwku5+KJWspeLzXbh1UMeiy8gWleDw+ZiTD
rl9bzTqsUe+3sL1QpPGoewNa8Vbmt3eb7z+rT7ZM7/mtWvUHLonYx9/olLpR9AKk
X30ZhiOf7PaJc3L55iQmUPaLz5+DgwV3cT8LNMltXrOJ+LdTYxg+kcJeVcHpwC/K
eEStlHYEx2+sVubsKc6C9kILqtUiZirAcz50naPKoSGhor65QfW8Xq7IHpv1oxt+
YfG0J86NhYUMEx1XsxyVIHi4ffxelhxBjw82NvmyaqlOIq/V0xcUxlIEs4gJNZYa
7Fq2GkjJ+XuwvKH923fvlnCPhEd/xjAnCbVxGuNF1+5j7JQxspULZItHXcJhBcgv
M1lEeFSqulhMixv9KE5cXhQouLc5kVo4w4C62I5SmDe4hh3dSEqzAxlC13dIvebv
Rv1NtEiyDTPvlQ9TSysvIGONO/go1iLbYyR5/OaS9i+uCfvzpAWC+xDhQH/eaWXk
Ks8GNKFV/DTTMAN7Q8FJ4tmMZFyOm2KtNOq9iiJ9ZymhYiPnjRsVTqvAwNEWtmtw
6hkuz4vtH8WmBYHzVx5cDJtkKlEJpPoBfOncw2RKcR4ytoRknyh4OMpQL4UpEa+0
ob0VfOddeajFoYKdN9fgj23Er7NFGhld2udbDJvdr354m3u10EgRAwUMfg8ajkDk
azjhbTfnYdlvGvwirylma6qScUvsxKvbI5HPNoOBZBlITmKK+bGTO1Evlxf534Ac
dj1acLbWvp7doqSq/G0j6KSBgU1mF9Pt46C8HIWqMmgRFutDyoak+RP5qpeYdxvt
ov2mmX+ednCR+uZ2d/f0+i8Nqf4y8+r/8q5SkBP6x0mg2SbOVpz2EMTwVe0RYFTj
bRz9IJKT1O4Bd+KNG9T7ylhTKZWGHltxMxe/ULtJY2Bz42YDA6GPdqVyVNbiPBCd
zJ+nuUJaUaeNAKVtJXunb49aGt7suA7lNSIyJoYc/ivgJXHUJkMbLU1IRSuHEAAW
tUwepcfmLakS4t7YYW7unVjn/cuU7SGNuWLBRrzx+o2u5NbcaZGrmcT9TULJlg/V
CD1lS1CP4r9fQ/tWuKOh79+KAzgCZNKQVqB4mFsjxk9RWy00l+bT+yKV67d7c47o
x67rZ6+comlyALvkULC+AwMH5ov6sP2bF6mMGdN8kIflPeXpLnSAdy1yyBptbI4n
QZ9S4tmyefbzMe7PCFbFaUDquRViInE3EEluHBrjWofaD4J875QDehXZTmpIkgxR
vx4iFQjCU1Ymqcalcyq+i1JGDzTJU7eILACXgkCLNLw/InVv5ViY3gvXsJY7CU1Y
eGglryUStMhCTN5ldTNG/L0hdVz8p+OCOYIsCV+VPSd5mD0SJ8HXKxOoyVumoRRD
jEE/lYDK0jGIHnbonz+Iv7wFoc38cndoAza+MaMfUK3WqxgYM4DMUgVrB+UknINa
s1tTxLoXBHyeMbteCdpMKUOnxxjAr5vUv8ZWIAIgVTkh9qU9B/yZ3iV7GVJu2tHt
7fOMC+YD86mn1MNjvh1DQ2w2scNjpfpwidGhdmSKn/ZeJ0BIrfZ2vzinL6u/kcSc
mjDFC2r5T9lsdqJxQLoPxojpWHwIHkVlbi1HvpIVVZuh+RhkBOf4qQhMDli3IrZD
EfLPbJGSdX022JAlCWNaSUZUkINFtcQiVGq4fWnYw2O+WygkYOUGQaVkNFElDZkd
hQPsAVeutU6HIe5Hv6INY7hFRq5d08+oGiEGc7prcGQQoKtYdwr13X08UsKccHfh
xsuNmUcAxXkFnJPkrAHgfBaqIKHghB+entPAULXKDLzF/fEwiyrNqPfBx/5Rtoxu
FOmHvyho4YYYQ1P1Jemuu7cGfbAGOuQFR2orCBM9ktspYuauroJrvLoJ6EczWYet
4Fl/MOreuqGQBMGFBJjdb+FyfjqLkmF24f/VcHKsNsmBhUMNs0kD6fTsKWcZx1t2
WzpUBo3avQqbXiF/I0n06oHUOEmn9reL1BXPBnF0xPRPuNNogvRr80OQetz2e16t
MBnujSGWgBz2H7j+LLnBMMaEO0Ouz0yq7csD0tIsTlQ2lSePJ6nH6sy4LcRwjihb
2Ld8n6kvn0ZkLGz3u47331NWqKO7RDxkpov9sFPhpWpQUDZJtfa5h7bE3ZZSt9gT
pD3Owcp5mxoxnZCcEB9LlGsx3q7wooWNwODZuLA8Q8UdiajxqPRFeCkSjIdX99TN
EZOb4nJfKkEEM/EqHX9WAMSOP8bkKTYxVpbUHxea0gxryfFjl0VBrJl981BjrkOQ
95Wb4nfZj2PjhW0a6eA4zKoDJfgtCihDMoqXPhQupVRSFR5IfPoNFzDrAsmTLebz
dDSwy9pfjxl0hfvUdOsYOVnjaePohCjmZx9BC2j/yABUVoPVt+2uAM8CEZ2R3gbR
8yVEJpKuLIKH8NfcZm2CI+L7Bskda+bR9OLCzLXt3kbiR6hi1wLLMCX3xMl/ZNz+
5pJBYzXIL3vxp6zSGEtCcZLUIv9VYDxht9bTsKZvGOYXR2jJkaHXpzg4XPHBDEcC
0PzCm3pHhPViPC79VvsNFtk55M+aOLnGsySvZj1DKo3Rrx7jsEo+JkZtDHasZnQx
7xKaFbBpqXxVhaGxya3foCc8nKZb5Rd/Ik5i6xehQHOVhzfyuobCmmXRf9mLKyp3
nLijfyY2OOhFi3L/j0KeO/xjks0MiscUktWT0V1dwUdXYmoDDOuXFVV+wLYZ4qNu
aqfFkpvaWLOnnZwUmfY73If4pbxF2Vpj88fZ0FKRKMY/CrhH+/dr20qJ6akOHUYf
uz9TqUaDO3BMZ8h0WItlIiEp1VUyfA/GSlnWJPbncXcp2+Ek0d2BdAQZ3eG/mIsf
LA3hKpHTtl4Np9KQ4u5K0UvvdyGM1TrMZpNx86CHYeQUU+et9ICl5CbS5Q/HJsOU
yy9LVGB8exwh9AfrIl6N8NXHR1PNQ8afwLJvtfSqn+taHbkdAX3d3EHL/skve+xd
3zJ6CyZvayaHmMtEwTyqCy3NMkb82tGVjhUE1S7XKBzymLpNRyxyOZ1yeNYUSTcq
XEGWAt6n3qSxyY27VKG3NFLGPw1LkDEryIvdCUDwBqzxF0R+SZU8FOFjSyKtyMzV
MKP4iCC69GneCxoOCYAtRI3CkicU4N5vwtm5VYH83prnK7Zo8+s8r0unMY3C77YZ
cfC5WaWwDIayPMg8sX0JfKEO1rptNlnsNwfClTfCKEkH/Girf6wThiUXagdRuy59
fZ6Ey6i345/ndIaVLuGtZr3pKuTDc5xs9c11UyD3b4FSREOG/eHFS/Y1Hat98jfv
12u9Gi+KBSeqKve4SaSCy8aF3oOknK0EowAvUqrgD4OHBThqe3U1oqnuh5CYPanT
tx2wZWn/CtpTOWvomTBZN4kdSXDSau4SD/SfgDkbiLOQ0sj/aiWDwVPnYL0xPXqQ
+jWqFNAkEKcJoIvHMoiqXovqrwN1r7O7Nmxmw/eGNkx0UKM4WRKQLKWCC+HBi9qA
WLI2DNGNcW69xMdfdkgy9fpRk+V/ys76uP+RXwAxktP1OMusFjJeiVS9b2YgxOUA
c7XcwRdWIYw8XdGkHdCaBVmZtxYNVS3N9q7s28aqy2QpAbWO0xqm51dDA5LKKaB7
e2an3juYTkm1RTXO9XxRVGz1hFB3RyDx2Rw7hMZlIeZr7nax4JcHOrhjqMlN5Pn7
m4RaOjnOREJ88NQP2+zr5/G+1s9wqRIvE06lHCls8hotb7bHtwBLAHCWkJmZDGhX
dvAFAfifyks66tEeiroYDZ8m8UUIE8vuJmipnd326cbzpEeLUhPRtsCWSpuuOmFK
n42LRBYE8TgttEkNJSzv7f576jF7MkVtzzpOHvDeoWl6EDaD+cRViLx88sroRZSe
CdU/97HLQd71a5CFK7xRAsR8Q9nzMuJxYnw2ufNX7QQ9QWEyCNctaxAEej14sYYH
ELJ3LrtI+HXGicv7FeVD1Zcpgi/BPiw7KNyDYSdsGAGhwQaPaGGKJZk5li3Ciaxg
sira+TAa8pMYi2rHvrvbFF06G7Isd/4bO8K/br8sw3cCgsEWbYtdtdwOaexWjIFc
OqVBWD7HmBXfJ0F074P4wp3l5X0QUV6s2LqEfhkYYG9RVFFmHg69Zi5sJn3J/zDB
ogDodxo8a3UPrwD+1+5tZ3q79ygB3vwjmNt5EtIepwOW+qaPW3WFpQJXQmNtibsn
OLsFCpnAJ/m1Hl/FSgnk8IP2KgobUqmv+vvKvll0au/o2740s7Y1FpEAuqIElmxS
lM7yDOoPeCPH6TBGocSLzCeJ3U0yL+7bg8f3rBxMoV0tiAjfG1GmjXEOIw7xZWJ3
OlcOCgcuLA79L9iFc1tltNcbfH0RAshN9VVAWbPivQczJuC4vJJjlUPH5uGvzhy9
4IAjQy69AGyf9nvgBntKRdHeGGWxiJPw0v+dFVD61uppNJ+TJQkI72hDI5kll2Am
XYtKxwL6ThNHZfAIuN3r9Z1+cRMtYIkkD8fWfiJc4nmy1EyLE5z167QIrklqRhSQ
ZfswkGoj6XiEY/1RdZ6rZA3nqOE50wDZHJ6fZiunDXv1tnqJiFlnXpJuRFWtENKw
+5ulN6iiD6r5xbCC9nEC+EtGICyKhta2jWybuKXFG0ZGmQ4zehD4gESkGTPsP/3r
/nLgcT5gsi4jDwuA4xwyUHaSl+siAuRq46G060JLL/RwAzc3o2HQ7wjWsqnkh5yr
TWiUfuK/tR2sZOg1zyiivDJZDq73wFBXCAAFs/3Vt9AsDKRvUhJsfjy4OMNAbNRU
zFOk+tU+PSi8cD3o8cM54nqv+qCrWqCqItUvYhLHWTNx3xrqjSJ6FZGaLT4++n//
93GKMZgL0HJT16euX2bCvvFFtZ6/M6w9OvMbQdYHfCK8vlWMH3khi8oipioH7wHZ
xqlOFCK+EfTR2im5vzsosbxCFOqA/JX85IczeVbkJLA19Ls04XfJ3V2sFJ/gIMBE
zXsqlUEGn2gMDIsiCR3bMHYHlLGGCaeUH6Y+QXOfGAFUPuSEBfgaOhqZyduQb9X/
Oxcx2jxpwHkkIDOs6Z7MuLxXiiJvmtENdGeXD7GW/BomBPd0nhlM12d5XHGqbTOG
H1BJw6BPBZ++/ii4vV0fLqWwqr2LVeUBn7H3H5/MvLxXYewbV45IBcemwfeXsgjt
cqlojiJNxGNtQRxF6nhKK72b+Cp6LINH3778eoXirGHJU01PyjCgad1Aw/daAClP
Z3Y10X0Dlifgoyak2C//GzVassDR6on+kAZYAZeaaJZa2ZTMuKV0mATt59ygRQ0I
0Rh268uA2cFBY+jeu8XXpq7jLjBDd7/a5RcL5Pq/SRHi5b6EwLEEZsnnmpl/3Kdb
y5F0IbdwiH5l09LifoC5wchLomnEoCPQNGaA6NWcJdLJDAj18vDxMoY3BWHeIuNh
e7TfHLkwiZlUKCnneSKzOty1hrrpAeoaVt10RtUoSh9tCk5CJc9iNPdYGoSJCo2P
Ufacbl2qYRRjPRGRU3POBZyNywkoo1O7N4wJ5hY3w5DhOy0/gPWY00kbYSZm67Vh
UunKrVxqzVseZ4QBd7nU5DeIDPivYQTuM7pZo6enm6OBylYwC9UfCzMY60UE03BY
LAHCLZV/X6MY02nGK1++ywQdo98V6QTJ4PVdz094/vDPsrDQSwixU/wOg+b49bU0
ynjioXKgpSHrAucMxpbJQHBphkK9okh4fCGqvb1i6Dj5S5L/+BjbZn+VDUtxripu
Jh5AEAKHkyT/86fAwvkGmfgQQOu3z7RA1bSixkUmcznCnrrDT8oYyys/hHA83kv1
o6HxgensO3Ikg5TbJIMmil9fmZMgbXNOj+vqKKAWitSxrmfMpt4KyehEHdZLC+QH
CwTDpnLrSV6BcCs4N0oyDXsbjuh3zJ8ByAcRegl9/WKN7t1EnPNOOHGDgaI+C01E
c2BxYYmkayzu019CR7F/5vqk9n0PpzhyUUJRgr01qC1z0bdDeJR+Honp1V7xLWzo
ML5KUaS28YFKgNgyyjcnz0K4hYLFcWoGPniIFD8Z8ZSuQgGhSWcQudEcNKV4Uu5m
MwsVCmaI16pq64YaB6iUl7b1XReVbK4oRfhaAy1S3FwN+9AYouG9FdeKdH/RMYPk
l+UQrnGQHjIM0YeLWJNlfrctibw0aUCbHf2YDVQkE2eETEJlDymykOv8monW6u3b
qVBOUwYPUcVWF6cpbffRtx67fevw7J+gZcrgdDf84eGf7BXUH27L4zX2G5y4vK0y
SORlhpjicJYW7mDRe9eBC8qLHUiEyEaxjtsyhPa+CzsGrfHQK/+Eq1N1nxOYdeWx
XHDSAGDdfRYYFarijEzR3ujGhSggwfLhnF72ivZ3vUyzcaFT5IRJrjDrHwaxpGQH
1tfndHL8IO35j8BT42ym2XcW/2HEguNHqMH4urmFwGNdtwaekefSy1miJsEJ5a5I
SJlwtIrzaq108+YTBBFWzbDVi+g5TjXigiGHq1k7HCyn9g97BZxqWuY8OYWG+AYC
/BPC3ffsR+Xt5hdvsUrejdwWrqajECWHlTWl0zKBnAKzU6vEIf3n8YUXbzYK2Squ
xk1ZE0SO9iJZ8tj268TZbSUxigvr3ojxjLtmkixmPtAWBqtl3axnkYa8ZRVmbVwb
EIBpg/LA80aDo3Rfv01Xpwg2u816Xg/Ys39iKZG1K2cY89CqjhMX888TncCpLcHH
hjkfG1RXu81HLDClxw+ABaW3WueZjUkg8CZhgMXfeIClkoM8tjG28V+/+Sitw0Fm
GktmeXLVAFZIJRWSIm/R6DOFjVpqlOwmIBGr4LxS87DIlCr8uXa+E33pXM25nsbT
3V4TdqmyNCN/UeJb+ABiAuSGYDOD5FQF6N5Dnkka3513OHUp32NnV6rzFdM5L+2H
4e9atfCTRIhRWPIZ8HDMSNW8UloM1RDoUwPqw4QHcppC2/0tzzdgYQXO6wre0yZF
isJoucLkSzozcwt/7EEGo+RCiL2PXlgz/oBSroal/3WgzkiTIxKjf1epqSOj/MLk
Nir0fnqyHLCCG5X0UNyA02Lm07KAW0WmaCmASDGAfzBL8NPlvMI74LKqVAWcOqL8
6ORZD2feQVXPEVUcZX6UDY0XKRZZfw3QzFHsIPol1XrTa1dXhr/CpiQoKkMd2aSS
EC7YkYJLPIcRG1nCi5/+uAr+dc19dF+EfHiUGg/Al6vKklXtO/slO5hfpqoGUGVT
io43ERU4nQ/SYAgDeKN2Yqgvg9HUbelP6K6tMJDJsYyAEiN2y2p2Gc10a/XE/sCK
vw6ctUPaHfEERIdGtiZrMEAeqDBExv/X9pAxZ8onkLCpLz+Vz5FdAcSTNSyc07Og
mt4Prr+HK9AHzpE2OkUS0+ROyEdMGVfGfYfaGxoPrRBMD279+WXwz0h66qx/J+Yf
8tqgB31A+2+pIgaRqwGRutH/X0ZY1RBTQJ3tbI6va1Ng5aOYZjKVmTWxXaIqV+5Y
dnpbSFZNuPcsGbGVCYzQzPAbWpsgDEgX5m80paw0yODJVQMsckV5N0vve77IpzA5
4K/h0mfewBYy/l0KwGGrOOUGBnVZS/dAhZyGYqznT5EfGr/ls9h8cj/bZZZxdPSe
xv9T336J1r3j+sVYCoGChOaTmmeQBy5iRSC29mTMoR9knvMOJU5O7MTztlylSsf1
UKE6ls1U52FfzOMjEMCdvtA4Nv4PQXIF9UiMXhqZJyCTnPJvWu44sH6MwI1EC1zz
CrJvGkp79v5SzHfTx3ulgwTw7UJsdz19BCljzDqvbZMMx3oRTymMKlk0eGGbCNZ2
MLhqA2lKIS8B2QP6pRZuIj14of5X4Ul5Uthfni6FTvO18oy3SmwK5IzYfdIn/0Vs
2t1pxHod8FL81gi0gX/G6+mU4WyL9DpirH28rHEmN9BbwuJ+Q3HqZOJIrmPsqXZN
cUzMuVgecpyg3SUCuEZE++AclmgafgwYAIJ+bRI0YY/RP5gCWG4nPjbXRw/djPnn
V2qzltMx3AVyakhOEBnjVChR9xo+nXe7MfwwZvDG9lzoHGn/0imwdVBD3rJ0pZ0R
qAZNw1CSbftsiE8SFJDt0rlSV0V60etHrbb2TmDuueyO5i6BLhqYamu6uxh8pniU
vz4YykJJpwovpYHYkh7gpdGnkpJjd+utGu40iJw4bG8bIfWr83Y7tY8OfmGe1CE2
oSv1fB+524n2jh2IFTIN1FA2Y3W7bvH+isv9TbSwcZEDIdbisduEGVYD7FhO+ydg
lvAYeZ/A1UEZp6gTDrdx7dEoerpBQ955KsOqgslbD6ykLQ8lxQmwCh1vaaTrKsMu
n1xOsYT8bR3zpXyawI94SwBzQ2CLlUVa6oPyiIW1thQhc/3fTQlvIK/CwPSRnMS/
ldHmphdCwv90ykyvGTUqrdnHRcdh7WjOjIONlb9Hnw3tdWBbh6ks7Wp/AOa6IIsu
KnCeEctjLUiNjgiv/7j7FRdyyZrwpHcZR+0p2uYLgDNfCMqFlZtkDqSSGXQk7Biv
NAHI/a1gPsWgWJus/Tcox6cLKBXduDw8L9G5q+aKFKFkXJcy7cxAhfoQB5mvhl8b
PcZtcB/fHvgfrWy6tmqwROumL3CWT1wwMWcXaNX/4QRBbhwjrwrcc6jrhU7lbKrQ
cAeQMtpVhUf71T2dFuo8JttiPLjG15y3rXaq3Sc5ZijQcfixxu3Bd1kBG3I0Qyqz
oMrokN9IkqqMgPtyh8bQX1xfrLPQYIMdtnY8boiVt9GAeCttHlDBAWwTdy04Rkpv
WJEKJPu+rlu4wPAu47HSBtJeDXB89ucClRhDWWd23ElEstA+sm7yCHsYllcu7IGD
U00hXmlSxQNLGvTfkf8UP53GDY2SmgBGjY9yJNycvw7zZrfFNVwv8iciO9VxCuIG
JUyiBJLxiUhkqRFwDNd7ehZ2dM5x9Rnm7lExcOEzA/japyG1FDO6eAAoXiLZ6APk
BuSYaYGzZzdtMt99in7h3t+HNxOwD1IvjsC50XAYsCJT0xWMVWviGrfUoBzvbwV3
7VEXeGQZejuyIeRI1CinR/E7S3b9KHnC4eIaUHzwUhfXKvFzlsXNQDOTmE2Ser5f
is4Jj6wOIDg1m/oAnKKbiaeoNSyws5OwGH7Fi8yPpiWyjmrxYYuPITVQCmjiGHOd
39NBzPr9hEwMkvU7AIGlAq5AdjJ47myJJdO/QoQFx812SBw3BaBbQc96XvDpjyst
IuhWTmhSZZBdWFbKFYzvKO9NSYun7QhVyakB8BqpF9/ae7nUH52Tqi8i2XC5Rgix
Furhjxp/4Cnvf3F3/aA+4pSVdaf6VY/ehM+xi1ogkpXNBgzcJWvTwC3I4Woxu6P/
dk5WJmHDm2yxXcouMCGeUxan2WQVLROZcV2syV0P/e4LAHQzNlxXWw6gasF4NgLN
Iav4r2JM4faEmG2ndHu2WKbP6WuFsQ6+FzvR+mtBwWSJq2tMG0WqYwGQHYy+OEpr
6j0QlLaxc9IlrkRc8iWLQx1kyAvsavl5ikrT6kLqyIpjsKeLw1/US9ojaC4cINFJ
VSLsxAxC+IPIrs3PMfSYvMd4LExIWJi3ls8gB1CPU8Jze2oYx9B4G/ruN1tF6xxP
N4BkXD7iwg2uAFUpJgyGA2v/bxrgx8ogf/Z/Gzhw34MEBXtYHHjKAbmoo+sRkvPr
/qsC6dF8fy7vcaq/UlMEQB4G0NTDIR/e8yBadPU+xq0q8BCsIkZXiTHhdXl9JEd+
pLKxSY1sUMtdDNbMqQhahBMUClzm4KGNyOEEcsZJcYi+UMngXa1qz8TIvqHiiXps
ApyP/jsujk0pZNyrD3M7zdOH7g+4ohflYHMQ+cZvvTRUg8mQQGzqOxmoUq9bvUJs
mSliH3170CrnvxGnyX657/dxb4lcoj+qZG0EZzIC4tDK5i6+g3FW1BCgTAyzYBk/
yf/sIwO/iIKltIan04559E3PSyou1vgKnJK+vGjAd7MLJ1P25s2mvAtq0fHCMM34
hpsqQSbtc5sRI6DD62mgbUvwau7zweJ91uPDeipCy4YzsxaCKIuuGKcYkyjd6rA8
ATlaJ9I2k2J2R10/B+3cL/sLIDQD8a+DCXKBK7PpMrXHWRUj1DDLzqIRitr232c4
45Y+gtV8VUeS1oBASBRX/m8KtAaCWAIYk0J80QvKfPgiK1Qpxy8cO3ofevBCgLyf
l56q0qszUZ34kh7uxFGoHBiIyR6Hs3DwehtaEhEHDBfp+K0gJrNTaFKX6xDBx1W+
PQyBBDVWCVNlRlGzF/jQuKFLjioJcpG36auf0eBQKegXxibE40SY8lOwXoBUbhA1
hSWP3mgdufSCywUjLyUsbcehpB74vURJ2Rx4JQtY1rjuZQaS7/A9Vh8eUs4YHL9h
v9wIsFAfFz/pCWpedzeAGNEsZjsQLSpPbmla/s3zyJy1zGU4rjTWob1qWHFFPrvs
ehDPyjwhFAxyU4OKKTTg7BkXmna+bsienQNXxBt0k/D1Lls9LCxoR9g1afhW7eaU
JT1y4gPDiLUUGEUAl/0szOsyt/cmsNe5H68wCzSKImEW0abXzVsfwSSgQyJwyYBx
sbTfRtGIU9lqaRDOtpHKfPXg3KEpFCJ57W2FjBb8HBoGu9vQ60d+bPcMHG+VNx+S
2fL/65+oLC/Pp0V7+nVc+21AnnYqylsYm7q5xwXSZ5iEsTCN2H1+htI698RP9X/Q
ymfsXb0oAzEnzTi7brdIEZ2mTcoUAJvvq6aB6R0mG633p+phsHFus5+K408u42I6
QfBXCa9nF4zgqC01haHpMcwFJEQgiYv9A44TWU856ACnq53RpmklEfHEQRkiUkDM
78nBHE72FHTzifFtp5uYWrK8NXW7cXzyLzv6Fz5maGmZWWTkyGmuneeGrKbpJekw
ahRrbPi0nSTMi4RSQ1l4VxSPJbHQLahTARL46/Tx40Ye5ErVLj6czuP07lgBQwka
xqiNiv9swLJ/RgpvHXJJvzn/+of1FXVX7Mo2LZKy9tWSlgACuNw4iWpBowAtib8N
qI5XGHuix41h/B4pDb6BREaQxzk3o0gvitNEVIE3747OkllbybTgrnUE2L9C3Er8
kDrJwkEyQs0E/3DSpAzrLzHVgMzirPcp8EUSX1CRPiz8qZXBtfpt+eyd7jSF6k/X
Hluurb34/cCOQCFOKjwaTwtdj0zSJ9zLxBQi0Xc3HoOYJ4AEMv0XlNCjUtUX0ali
ErSwcBiECKawhkbR6NE5F/CyefJx8YML7pdt9wBULbZGAQTPtmDO+1DXsXNwVC0d
jcTKWJh8KQn3sGnqTYZcm3hykol2Qdfj7A6S8XadeTBM8t08fNoJAp61H5GKdsvX
MhHR4Ayc1nCVZ/6q6C+ABzHLLG+jcjcU/jmsQsGSIAJORpKGvFJt9MExFd8uflfu
q2vFxCpL9AjoVppkQlgm9kW6oLHrlTxKZUMDFyPy62TqGj3nnCpwxJsO3R0BCvFW
M9nlOTuvWOkVVg6dVBPbX9lkYvG7RmT5XkEH+NOSCRAIFYEJv3Lhwu33Vd2rlee/
5Go2ALa2kQvTShfdYE5sldV4OmKwcqHnOzpnbDGIdHtLG84oBQL4ulTp0OZfFFqR
Zi0sVRmnF9fsvLdPGvTD2UVxcU4mJmakPxqheD8YhL6fPMb/CD+v7HxZHmcNNT8z
ez6GOBW3N6tzich6EnaQI3dkidDxGMV1836a4SaSiUZW5QhbUV7oKOpvUDa0oreX
oxE0wpT7JjAP5uHbMRnf6sGKZBQleSFF/Qky8ePMsoYCPSvR2z/QZWLJ2Tsc8/pe
AfE1pWzkDjwzGA81iubCD7ic45nFcPCuaMjANT197C8FoyRIM1OkH4okvJT8F8K0
fcrnwBprPQyB60fBX8InSIITFwE7L7p6L9kvONVjNbbsrjylAA+Q3KZ8GG8Tmfpk
GwRVUAhb3DwNTZw/agBKynpfMtyh2vULBRWKwxriyioQHBGpT7sBIqUPIiH/T/Hw
s1fXvhQangCOWU6WRyY33Si02w91QrfeF6y07yY3sANKmdXXJJmRBCYEaGVP+zFz
SMNCvQowKfVlZ3ePgeh1cuhW/g1Q/FJsaMsjXQnPCEAnGMVsLF5XrcLbyjurxnYG
4JeHvB4WLEnsqkBFnLdGUVbYJ+d+TLu3uPApcrzC/t0sZ/zxcxU4OXsY6h254NCI
2oYg4ZNf3Zaiat4HUZpLFUZ/9fhDLvRP728bXogamAWlmZJXfSfW7hVs/y4rXnPq
uy7v4PiglA1p+jVAvJjmTdj7izGHB6cDkJS4Zdpu8UUVktlTvZX2QShdu0tYoMBS
WX+UwxdX7I7yIpYhUOqHIGzf/h8SDuqnzi72gaZVXA0MZFY7ujE3XV966Y9TwxYT
G25UTIi2n1eEqpU3NQakN5Mn3yGvE4lLjh6jAJ5pw1Stal03+OftC6D96sx0UOU+
a8KoMWv9PojidUwhL1t4Iiezzn26u5x1Z0r3eD4EV138+njti3ZVh50C0QqtG6UA
9UnzHXGDCPytUP7OdNg1D4Vp1fDqcAMEnqLB7J5/oSoDFLLp5g1hykxyKzKJrJc8
xbyVFps9KbFIy5e9ZFOWzlBKkfR1WXMWMooHPLxJrgjc43CjfL7zELe2x64RGisr
1qMENyZsK2Ld/FtoetK29bsSEFz1DaPpCYDjdQ6uIXCIhFrBeg5uEqdxhW7vcSJZ
0180eN9slji9s4jK8Hf9686s8gHwrGT47UJ8pHvRvs++3U4MiED5ruW9NPn7ou21
00+aMRUd3Saf9zLFHiOrzSL2euBWrAe3xzyQmRz2KBT3XxO4mTM6m6NOysW2radS
IerW0yXYlenzR1CW6I9jiEKUqVevE2TLWLx+YpOLmffrg7oL3TB/JWX+cygp7JMj
NtOWacoTZVIapgsr3Hnl9pvKJBD9IfYfbg4plpkJFZdgG0TILC6XRiH2iaQ7Cqwh
RKXdKl0eGpisctajS/KoBPiqOgiqO0JHmLKiK2pt9IfeZsN8EnxKHx10CutOrPbQ
aMIcsezThuyAAYFWLS92fSi3SMvu6+uSeNx8ZcDe7h1ycWYSk+fJ6No+hOqIkhfJ
RrIdLqeKlHGfLGEuvVc3GbgWUIjkDm6lnjeuW7iHD1pfch0lf3HITlG1x0VYrFLp
gU80fZMgi1je0eYryE7sJkDdbrGexZgyW3zMiwkhm/rmlv+XduMT5nKvYGeFR7uu
4w2WibcDwWgMJLZYVrUuONv2LEYrZe5Va4xqdBu1wRucDzpLT1AhrGOWFj2q48HI
P9Lz8rWKwVI2AD2IENGihwuAqPj5dUd6L3q9VgbKm0knCB5mYhZdxaDc+r4n791I
M9pqaudczjamtwkagk9QKWZtJ6cLjc+xMmWaqD+ChYN5ud4r+5w+ybasWWthi5r1
3PUUMZGcL1ItglcBIY3O+OsPaRRhoikYgXC40Qm/d6m8f4ZSthcJKG/8NCXF+AVA
3dzeg53Cy8YG/bp2Ij8xMnWOvGU28kqKdcJUB0SPOrMWTBqbawfp+kSLR6PGzc3s
FX63XWO27ginAgJho639GmbxiBNbVAP3z2Gyr7fwY6OpklgOQcO549u4OuG6Pc82
S7OQoWkUoYz21SglxRewfY3DL7PNyNl/Au2rnY0hzabCqpyOHNZQFKIS1LZlthWv
kpTPlLQGY7GDa5HgSCrrb319kDnyLNnTR/ChJDeizzbpfGJ1D4N4aoP8nuCfLqbc
ncqAAbaujlc4qrzxLBxun5JPBPGIG/6HD1QsxjEDN7FRxHGzEuAWR8qQpvRg3yP9
5YU2/OWvSsBpo2rOB1iu5SzzrB366qse45QKnBmXMp9jvBc5fr6YshaU3IPJAAiy
iA0oKMTFMRu/pb55wZP1XYWi34/TeIfxHpPn0oh6JQzbrFWUnooE9Oc2d+jTm5Un
3VgRPHWHG7jJ/ZF8sR/6bDe3TltaPw8t/DYjv5I9cI8IEnD7RkL0mB05fKlizt/y
I8EFgDyn9e8ePsUptACdp/CKrQfcOSO/7PWps0/wdY38TlwJANXzYYDGZVVKoPCh
2sLn4zxbwpLhLmrxcyYsb6PbE/IVARY8uu5ggbZgwiuRAoQaEyC0Gv/4s99TPiCi
0TUCMR5EnuY9Z/OZVCaO6cNSNgsujtHj86rC43DDXBhWxfV5iENDfuRu3hQUU/xK
PiPt/0lIhuPtUd9nP1WYgtnI40efjgQ25BYbwQJPmuCaFmjLfL8J8JIpTENt/Ijh
ucSxHGaqw/NWoSlwomYEiN3GuxdzpwRQuKSGNpO2qznj5utJnGQ2EWQGZ/KGWf67
Lz3i+zPGK51wbAspkIVIjoopwhAFuXBZV7Snkjjyl87KBQTwe+mzA9O4wqhGU55m
t46kIjh1b7MmPOkylxnwfkNdQaheE4BJT4Ww4tlbm+nA0lwdN4OSWokvPLD+w7s1
VaoiP6ppKGGlzQf+JCJLad9Ms0nDFChJVzaCJcPKGBlR8NVQYeXYiqOAD7/+Xu0/
w1LihQW8Vh5OBvyP2gnhdnuG4ZEyhcp65LCEIl41kdjDWKv5l/tQOsZ38p+gmR7/
RrSsrDoJdL7hZVfVZNcZnpyDKfdgIPOpc1X0fcMjYsx+ZnY34Ud6eoFsyA2KrzOV
vOqUlJquYZlwDLI2cLiq7+6T07TQfDshsos2yFeUIKNcW4P36uXIn0kEc2CmnK2H
zOg7Al/vJi41O1act0MfNZPtDYYP1wB8Gd/rZPyU6BlXvJ2U35KVun7WFl3cwVlc
pbFoDX0XivRK6+5vAp0bXDAIZtOnwhGksZN5Y6aih8/iU+mrO6NPtbrnhAtbX8Bh
QxvMvxwPrH4iD+QhsKdza63PeBNbf/YN6F3avhz19jifn301yfBdpRpS5ssTblLS
bzrF8R4bBkFMXh9GEqxYUBgOSuOdT/rwarvovSzHOKDf5pU4aQnYOub7j88cMVzn
zHwB9Wjunugth6iIMjH7K2vsQcHKgI2YI+TF90oZFmhTsta1iS36HZ0ykcH8oaGF
m+tBqcASUPFiQXEN0rCzQ382p3B/hK+/3r+50TYJHYK4cBNfimp5up1Bv2gGEoQS
hpqyh4LrydUEk5UOjoBVUzsUWkN/qkfZDHkgV8+c8urjDH39UnjHUjviuxLzJowN
assHUYdKuJsynqRDR/XbAPbMvhg8HZXht9cvKSkOeKoZcq1GkiouXZN9ifn6GIkH
qIelFhEF+OQFyAnKGkkUBEXBMZXj647+BeuCv3L3x52nSthfJGsoJZFhnPyM+zgM
VRKHaNphBuyVxu4dZxVw/f1UsWD4CBHJkQ6yOqa25uHMY9PJ81ZhqaohoH0I0RoH
Qocw+2aqrdVDv6muMht54oef9K7uT+ymmvufFGWUeajuXZwiybWvETfkmLkLlKLn
1Z2vgo2oPixK7d+famX9efttMQ46J7OP2I5QWWw9xiuC/lSz6c5XvRJ8e0PMuX3a
fJJWlJXMVSAsvu5t0xnLOS9B3PY+vwbVsiT2wesTOVpJWxk88cK/3wYHc410U2a1
h8eXpT1JN+9yIKbl/hYrQyppgJ4PR1DYJL2YJ4X1yCsz4KeoGfQ4QLUOEwJ8oFix
altbYGf11h1utOuTte0ub4byfRt3zHFfLO7ZipfTWty8CFyePDo3JfwU287PV+d1
TJT0FdwAdjQ9qAOd8fWvDl5U8EUoaVVcnFYUWpy58sJYgjKA6VqdKMij7Xxc0leB
tzWDhinvEECZDmEmrxagJ6lw/u9tDAKZ3rs+9rw49a99l5Gh22OUBSW4sCuulV5Q
JCEtucVO1xBZA58g0OeOa4LUAatmS9ylcTq0ltqpBa0ZQ22GBWjN5mmvZhI1AOkz
3aCgCXyKF04RRTSGyykoWmN/P+7izmVtJx7vpBif4E1OD/6+58gVlC4P1yUOOdVy
JyOCA0A56KlIVN7nY2BlLkW3wSKkVa5efweWOThNFL88pAQLTlx3cHSImY5/4p+6
TAflJ0LQO1aK3i/yL256lX1iufuczoEp0IcSSCaS8ayE0XhT7gjD321+nklPDQjR
HGRX+N3o5Y3dWnOJuy8BHJU7HwTY8gJn9NTVJD73JSujXZFmm+xTf4FEGAEuI6y3
g2UtUR3aF2uqrhdITIGanvAdvkV6uFM+fnxUVaasx5b5iLwG7nCtqw7zKdFUVtj+
9yqQQh6pNPhq+wW9JRrCWRtWRCodJufCOSQ4CTvNwX2Jl7sc0HEOUqKnAF1PqdMm
+EM1iaeqOoxJxFYAGusrbobeV/1X2o9Arv+8P7QE202KSqlLWclf5tvrf/HKy54m
kwaxqLdej96nb4ieI6ApZFckSxw3aaNbfPTGsBQksghbibeGuJI09pnaASsYYAME
CEC+Eij/F3uXRJv1E9U+OY+19dcHkNhS42aGSAYdgAUpnpyjkzxboJtvbT4xQeRk
Vi/OP7bK5i56kZ/iaWog6PvFMDUjFzbcDoFa6gqstXbTP3yRhWpKC/rwWHCJJ88V
v9fa6oFBuxePUB5ZhgphhIuLhUoHEOpzXloOlYLdmsnYH+BuNGf4YAPVBFSkabtU
TiE6elbcZ9Ijzn/ZXvnS2BXGrvoDWzn5LdN0O2KNMLilZj0zEyFsIEkMgQG9zP3a
HKj1odJb/vWeSdx7Ls9NiNohuqjHr2644SmFyz0EKg+fT35VFl0Y+g+u46YidaWW
cJ/1SOoz6nUbDSgfqledYxzr8XzfMB/zyuWyQC7SaJ4vIQ5NoVwK3ZzrYqhS8k5K
yMDuROVYLVtCw0n8YHVqL8edqMy84rZUzvUBGOWyftGLOera3AHp/uQoaBCnZ/VW
swhSFqqgs/Xj404nuPL6LCZtiYnP0J3cdXDQge16S78EP2E+hg8hu3xlVdy26Yx2
HywmGFh9nTzFjNvy43u6V7kjTjwPuJIq6YbUElXk2LZxKF3kKAIvSLrL9GdZY8i/
mZJA/2vA7eAG2NwlHmzzf20WmKyaweSYDC9FGFCLuZEIASUvneQFGFfLeU2RIdKM
LUukDIFEXzpA+ssCeECUk+oGe/jyquIvaNKQadPBj8vDxr+wnYHl4jOWD5a8P9e9
LFpLbC5XL57ETj1JEVU/KR/4ZHioua/ooa5+0NCb+o7w5oukI9a7Vly2AwxUOQ1k
YDqLZjq4OK63P9/5+Lb6y1YdzdCtOfJsWjrM+eCcDllqbTutH4goIt2Gf4zdlLIw
88iboTQi7T+r22oLczQogZORCvhqoWCG5OcaVCPwPtlc+CvN6Ty6988R0qbczWo6
CXGpJ8hZSsNfcEFOKM+d7GUatsHj3AprGqLHbUsFekZlBVqV9UzzEP/D3K/kyvA9
VAULRUAGl2KWhK4C+BRfXGET76bdfJURwtasIFIJAX8CEMf+PzrXWruN9k4MECEr
+oOxKvDGyRr2CIJYyfDPWmFC1xftKwYk5C4WbuBzLA9y4yoBYAK3dMMqGH/HwxSr
bJX/n1euixPMkW05SVMDKqzGRUmHVxwEnH1mZV1FfXToNVlYjMvMJoYg4onqxcAT
bd9HBqEDwucqNXJg8+YFf2BfrHCBhYMtvMxQReAl/Qq1s15IbBbh8MZt+7pL8Ep6
+CZMLy/PwEXJFrBRgP+DJuq80FB2GJ1HOY9bq7ZmDwaUX36CV+7NoH6sa2hobLUH
GMZKGUHN0KrZLM26Ydx60wp/FGqQp3u34x0P4FztDt3YzEe/i4Fm0CScXWgegFH0
0Xe3EUsngtAkx7rSx0VwQwCx3rU7g/fHmbwbmZvBbQGoaQB+H0jgVq77dQTvVFN+
pm1xzbIZ1fOQOTPg53fBVhjsMJMiofXHmCS/0LIV/BvAJeOzeRfcp3htIwCRhei0
VzgLvChp67ViBOsyKag23YWlIK3+edKOO4M/tHa/BR/nWVaWpFTOl62oLxG4vB0B
zZgAePPSNoWWPCPql+3i1/gQnQVYQy3RQ8bmzuFHIREGjQAnOr9qhy4utzAv7u/m
OzTGum55jZpsZG7gAAgYvv+02mde4d9KSDjWLxWks1d+hn7xakHpZXz3kwlgXHdH
Il/GnkIqgGO5adkB0GL+FGhTaNlejF7xPLTxgGfZ3pDJ+wPRZqFiRR4JM0UFR++8
bMtbaz2Fm+3yVE2dbWQ4ir/mpr1YPYnf6xOH0t0PT6yIvZrpi4S5FaRgTDUuO58i
+8cVOs+/hqRWAW+jrmzh5ei90UDIZNIJps3ezAO6m4AC7MkKyDn/PT1/bqqiC+KH
5/44W1T5IoIQKqUFtNCBNYZ57WhGxLYHX2V5dUmzCaGI+7aGwcArvRLhtge0f2s0
o42VFB4Cm6p9lpCFCXEn6N+mgk+kVVYQjHarQ/vM382O693oW21OSywxk/kIP628
/H9sbt6z+CgXwT2v0WqcNwYP2/tOi88V2yEj5FXOdjwQhP65GXclX0RMxmV6XFqC
efFkYJjZc2LC4QSGP3/HnoY22yMSBGv8gaUSHW7kGDHPCY8KqyvFL2uDhGUDbAPG
D/chnW1v4O0/2Q6uEIfnSFQeOvQmp3Jsr0ChKUtJX7VLYh0bSGmPYjBQnVoXi27o
Qu2CusTrnaR1oEz0QbGvcd8fn2dJcuJAB+us4MC0phblh17u/nRNb5OsBkQoO5hf
9bTCAXjrHk13edxRxfVT7RBn318i3k+sEZ5k+oQAgIo6ruCuJ1bbZCF51krBiIan
zwtc6/EplFFsiyo05OzEF62trCppm1P8nFO7PORPLFALVFiVYwgjOTfWHtyIpNOf
A4piGCHEvdOyW+FgEZspEVOUVH2ngp5IhgtiflrwQ05lz0wPp2xmqmsDY3d6/MkZ
LGtaBA+8TeowTMPo2GJg4HSnJwiW8cbySJC1n8rzpdk/11LABGEy3vgMTLDXTMUx
5hGLfBBVeAzO0NzbNezXG0Ee4qmhc4QgGAtZMeY6pJ7SRR6KFkq7hdc0Vh0AJwpQ
b7wK5cfga61SD9QT5Wqi02izBjB/ApIGXpnSAQoXTRKZTQpUFRG5t61UrY2m9V8H
aUvqTA6k3bYkhDftul5M86etiWRHXgo/f6HZps1NWcjhx8BwQxuBpnDtHSmA4u03
UomZli/qhTiaCon4sU/zVeDDO9S+0oVBy8xSaE09ESgMMlNwnGxKAMTmToQA9sSe
NWGIGwGm3NGHFE+5Ldf5TLO3XMbZSXKaTG2MpDhJGeddnLqCndkqRTd3LCMHS1ob
I8vYMFtSpuCaC69fzMAh9OI/uCrn92/R/ZEu87ID3YkDmp1HFjdGg0LRczW+q4EX
ga16FEO9AhXyetzZUA7j6NqFCxJmCOhJmTrJyrSECxYky8/LMDEcLgy/+49pEp6b
MGVMmT0KfbgkF1LdSUYQl/GYxx1M+3rFm9RIs+Eytd1I792sRgaytzBZ45VLKaqR
aoIXTKVajOqZamRX7uAgSpA/hs+A/BNbWfNLFmvCESS0zSLfJuLWElIj/bJ992UZ
qRTQmSDoBwmeFb6Hjcf/4/reh3eeSI5tdSAnnY6cogJ045SnyzW2KWxHsYbUupyd
4jssl1cWsqb8GhrkINSfFUEswdFJPKSL4LK7UsiX3cjw6kLbKZ5Yuo9XEg8ZVQUq
w4V1pm/1SKX6dF+2Jx3yVHKR1lQhdR/K2e/t5fFaeepSe0Z+3Gbv2mtFmqR9xmDF
jwGmoJsVLFi3WfPCcZfeBiDBuBZInhL/2SCUHvyN/9RwZQm/5OBUO/dQkufFGdYw
9zVdwh7Df2a0F0KUKRW+2YNZSuGIU5YOjSrm5enclxvzOtn2w6jtscTUP7ejnS/2
JTOiwxmPa5bAholdLa3EhBDuc4pXg3BDtXfeu9wa1/Bw9HiXBcLIzIdc0hZ5xIjN
eMJ7ciJf8IeAQo3uNM8dGzt8AsXuUK21Tu5hjMHFB/gKRxFimjd/w2UVVexVPeAw
Cna8wL07FZlrX2FeKJ8CIWAF9AaemEY/YsDQ16BJ6GVKhf/BWFX1/Z5TmkEPbIk3
r7Q1M7HJew7lUoWJj0PQyD7F1SYSovNLpxnkh7gjnChlCLoq+uoz6HK63NB1aUar
qWxTVsgbBPPcDPeT2vfFCZYc/WVVFSd/76Dtxo7F9+T78ex0xUxndEBjKu3fcLnU
Rl2olioZNiY+2WDuxyE0vf4KIsnIPovuF5A59iNlJdnW9EJO06vorNxTtlKcBT8n
kf/QB9LjVOjyniBX3kdXQ0UGwJyePI9q/qsHVF7u461goW6rm5LxeZZGZqdZNXIx
LkToiGuvPyDrSFwsSptqFg+mtmBzifJB3NAc02AueFjpugKZ5bhlByiAZzJGlmSk
Jk9I2uv1I6JsQrFTSjvsO571fpMPJA+dzKmM7eBIToWlqGkIuXQzyfZY34vQIcbn
Wq4IXZVtmFfsHf6R0fpJa1l8wm4pwF4kF2EIrYdBNPtOHMB/q3cfmjGR+ZxcMvPA
F2viQIMWVAHw8bl5XiMJ2sPN8CyKr0ialYYVTTiwlgmtuVnmijv2jkpMF64GkwOH
jbLr3NFBu9uBVLgjEblCiHM7CILUv9VszIjFHB9ZPzWHjlZMplLWRjl3VADiqaKx
PeMueU7MDrJTPZ1M+SjrizkLr4nVu3/1kbxvoU67nJrtgV1JdxfrOR5Ow1eJa7MX
5jETOekE+efREc5yuiI5US4Pytvl+a1hQIVNFPTzWYtzc6ttlYRUbqXj3OPUzbi6
JzlkONOFND6Y8n/EgI9qEUPNr47Wvs3uup7Y7ofR1ZUWBKTVJbsO8brIAz+jIXix
pq9xQfjvL1srrI467sqgVs4IH07O8HGVBqbScpV3+FVkHmL3zGhmAw4s5iSQcEri
Pxh4aqcz5/7AkhdWk4W3GRg4K7c2Iz5vO41R8jc+WqwhO4VPj0XeWXHfZGYbwOUn
6Gv8f43Azwx1B9iQfF0yozeM188OLGOxY8/hms7+XNifJIw38HHr06OmxQIqsasX
mELiT5C1v5FdADkVTlX3+pRFWEe0WKXNZXSvrMKVSR/6ujI90ojSa3n9PKgoNiBk
erEjBqy6f/RdyBfBm5A92s/+PxAiPID+IM9jNgZCDB/1PE8OI70fh4hFOIYQFuW6
1HRviWivBFBzA1U8GMOm12ibfhW5Cpwd6CSICiTTxNk5JF8SYVweXxBxLbDAp1z1
7DdtVpLZMNO3arHQBrO0jwB4q+Z5ImCUXqll1stqbRqdo4WP5wE/Lfy8aDLw6KxR
rfmGr6NDK7HTN6398PoGl2W2MRKRFffOIknwuXXR5lKGHFqKX3sO9ZgyJBhiUT/B
aEegPrN967xeOSsvpHBdg3F07kM3TbJeSyu8FRodWktTf3qG2ZBiy7d6WdsreG6h
yI7vcGOyn6LMfhz/6LemtRFJGnWsgOsdrcnHNNpGUtYCHsPmkPB+S+ZEQRSgOlBe
oWIA1EWbtgJ2m85lolWRBkFBNltqzI59Q0pCMKa4jfZXcqkqIiNDuXa5bbKjVQbt
0RZlRSlN+HmYYycCGIWAP62Jwh4gOQ9kWTCpK2ISQKcia50x18WuFfqM3Ri4YwUw
gEoUPsk1/hspOaWQ1retSYpAlJ7aTQnzXWeoTywDrPvSGGcmf941bfijHtGqlaia
6NcPb0S90SX4Y1J77p/KrdD3bqYled2LbZLxkyx3xRKAAgj6D4CmoGn504MRtRX7
r1vy0yFuJlS21uQApRgrtV8y/VGY0r15yqT6FVilk20bJY9p+4jnhskOPrV/Ijmd
LTP9BYI0u9dnViFbhW9i3zSd0DjTIPD+NDbfHGR+K4OpabnsTjAh2Ts/BfJFaRrM
7sIMW0Ap6ynCxofNH5MTrPWgAfrFMJnOtRtTc5hmKHfNIno3WEOZqipKI+BVjfZ+
yUX9aR7GWGvyaa/IP2oRpOhjwnUVn8i2aytq8/k3yj+CyCU+PD8GkENYfTqlT4zA
GPXlazs2d1NJc+2HquEEvdCea7g+wPYG/lcSNUxqxyWPivlc9FZCKfEmVR9g2dKK
kRuT6L3uWlqbV0DqxwsvpGRFA8o9+3QR0Q8JG7vXLlo57lbRq9YbVaFLm+Oh3GTO
LZwl8eDobaYuQvWAtx4lcBHFuXEhIw2448V0JePhP6nNXJK4GlKyceF10LOQsNFt
2hGYqo+xgjfbapFHPgvDMQVh2f4lJ+0MS19azwa4mllNsn1lXbKZvC070dk/iNI/
pA+P6Djc10qxyJelPlQ+MRlWF4HRJ46idVwCtYrdAx6NtNj6hE+6LU2t9j8g8EuC
+W2HiISuvqOEs9WQDOrnobBRq/Eti2znDXDss2PYm4Ip9pLzKkSjhZLINQkCy8ZT
NEO0WfY1nnOfM9T+5iU2Vp/qs3aQnQjW3L3cFdDqmo5lWVFbYd3AsCqXqw1OIUh2
RcFV2I6RSc/OWW8XILjpMtBqcnB9AOnwPgT5Kqgi65yraOYUt2Oag9XnHIXsaUU8
FM5ikcjems0baj0rwhVql4V1snOO/9PGnPQUN/NiagryeWwZ2VfoPN8t1mU4nw5x
6PD4y4i+ime922I5RSMqsttHJrt5+2ZQaVeIB6G9ecilC54NJQVVoCXRYDsPEles
9Y8vsoJByVmS8zZs+WbIxwPMHN64/9iLXo1wUB1kAYg/jflyl/PbgtaZVEMClXCV
F4lXL1PnOt+Fq2vq2PBrQh5XrF+hdnmp9w/Qw1+43mtV/xZ9xyUCtYXBouI4aAFL
Ca5k3bjaNSAYPeWdk8gqOTzADB2bJ7I9USy/4Xc0NzZfJNk+nmOysDIY0gpd/7St
rYTq5vCKPUh7D9WC6ryD346tSNMKu6QtP3dph2EPsyVYFcXPJCV7HmM2It+sxrTS
KAW+8OQS7iqK45mE6HcbNeLuFvTvalvskEK6cZ2A5RpsOw6UiPfgRBZy2red7Y+q
mOdbESOi3sq4tg2JFPFNY5TUuzCvcSFQvOtDw8sVOJcrgWeDHfkiHv8tjkU31R/7
0Eu0OTKjVOBZffHBJ1PVCsMJPQZni4geyyNpPPuwaJaI51HCZEz8vzPyImeOgM9w
Urw0U3XIaXIwujSgV/w7OpFySSTMcm5aqODjaJcBPy3jZXiV9MtC7wxSffLt4jSQ
RaKeJqIsJXQiFvItlvloctWUnIsvTNJ6DrGCANqFJeD+Et6fkrZBxdBJzwL3c3q5
b3tQRaM9+Tqecn12sKH8n1coQrpsGycRxIZ8fjBq8N3l+HveYtNWQGmO9Mo8mEdZ
lPcSP0c6LC0v9Lo/IiF0Bz2hmJIt01i1qVv8TmqRXMm9HJyh168mTiqEs71YBu0M
7RcOuWH6R8KWVXplPEulIqqoWkYi4qoujsIe1uDv4FqMd2o+bylgS9CZyGhRaSlo
jmlOUFbtcdOKPfjVGabqC+LTGNmgpPv7vGk/f1q8pv8SfoW4micvNqMxxVaqLb/R
4GmKzAxKFQOIANMJmrFq6wfWpjGHa6BHs4S7JNBnN7J+Pft8kfob794R30x1R8Fe
6YJppAMxB3fkg+heCPXUkDV9qJon7j5F5AsCM328wageXjnveEZK/0U2b24BVDjZ
tpFZz2jvFuP9HGgONGxpcq/ZsdGP8LJ1Bxjd8nptHfJKhScdhiMP4GqVRWlFzwD2
LGw7vMn2HlAVksy96KuTzYVoUggr1vIDeqxi5MKm+Nc2U4CBi5i8YUNf8DZJ77he
Q2IxtboQT7zTpSSGURxYbzZ6Mn0vMY6aopBv07Pf+CF9i8/5HCenUfms54SvUHG6
hC1R5kahdgze+a28Bqu0XtxpUbVdktzzinJS+K3S1Swdwu4yQaqRXT1bYUgdeVZh
98nDv6+lTltwZQtX3cJ+FyJ4BZpg7HLWxflW+CK8ac1qhnkC+1Hy2xJ5BBKJdiV8
KW02oRjtlo1j/O0oZtXoq8a0n5YbjkAj9ESFUI1QzsE8oHCVXvdigMi9iEcDJ9E1
Ghiwz3OH7i6iDJAUvliejjaOdnxohNhyEfUCDYzFCFwFk/yvrf2mYgnD1wj5Mlla
SdivOYtuNadBMGDtRg4Rth3X3WhrK4xSEwybDujIpepXGeys7+0/MJFI2FkVHLDz
Aa2MtTCsPiCWYy9VL0/vt93vHvWHb00f36vNYAs3v058ozsdeGGre49CHBm/xeNw
uvowejHVtdok1WICiKaFkTymgP4K69ZZsSGsktxZ93oQ9NBqcVdJoGG0L2EDNvv+
AAVDoLPCHEv8OxLJ5WVPQYiRUGcNYHwNEkWp8hH7KWXPmYVjEN6puZoJ44cDmOkb
j2XQtIOqUKcY4mfrP/H513QOsWbIHQtZeyljzi93f1RHwuZRr+2YQ1RNYUh15ue4
HqAj8CiKd4UXblenlkkYFx9FEQ0Z/HLvsZwOezy3amx8VOGmlrfTnhmKiM12eW9/
vZEeFmogPc3E+vqLKkdGt+YPH5sTOyjSMZ0YaDrFs/3p7kbaCcFYW8pcF6Fb5odm
fcj+pW6WwC0FwCa3TCQZEleP82qi3Sr9CtopTtla0Yyt9fiRN9iAQy+NpFv5XDeI
zgjHeq3Aw0dq6xy7qbFEl7h6lz7dm2iL/3S9Wi4wBahksIP39hlZCpTCb8SOd7bQ
ln8ukz5YLoshm9Yqx7Jc9UixXNR7o1QE9C5owjD4570mMkU/yuuSML+JFO8OmPW8
hbeOhNGoOuIIrCt2/TauiyWhbwpIKmPZDocjX8K9H2hDSV757f/Bs42Lv/cfkmq7
55176Klygr5SGoWLRgbvDJv3wLo1vpQlz0qMUV8yB9qn29MyHve4ZBOyoCbyZWLc
gTs9VSfdfLMPgHNvWRoiHCHgwBKlxBlCcIuFVPu9Ecx7c3t/Zn97+qxFvQiOcFY6
a6klmB/pzeUeufl8GfhfYn9e1cxQ+sujU/bkf8R2+Gmccw9sfl7uHXtp/y24tpp8
W+JmD4wZ2cjq0zA5Lk6o4TYCNl5Cql9wBHvtePSOoGnLUGPrPUXaY+BSqtb78SmL
d5sagQxwPAzHyNrY1RleaG/KA4AO77gt6j6RHbacbBW66vG6j+g8e7Z74w3hxyUr
HVm1enkW8V2jiVPEuwtzxbiFMCM/fdqeg/Jac/HmzUoNEjHWFQF8MOAXdkUIGfeU
kyBZTGkDkDeazZI9Htrj8/eTmiPbxpQ3YdfoxpLJ3iTYriDjWJ71U30hqbz9QrmE
fkYo02nqJES9iKnYbIW5TVdqEQoRhWUKauiZSfhsWloheiCi7KgKMD0rYMvFXbWW
rdgtHy6y8qhGRJq6zk3QwLB8BQROHikdfqFdLaoMZc88lc0k/7fmXIwOCtN9ErdG
JP6GSjVSkiap6/rSke5SXdCjjKMgA7DetV9+I+1tr7jTkUwG2yWWD6QkRkW4FmMc
ngHq7Z90wE/JH6gf7LZl2+4Q+J9G0ZoOSQjdHAgmP8l0nsqz4NaHFxXSxWX4LxYA
yLAfrJsUrPmwyujqiyiBAClioVPpqxpzNV6Mn1sg4+LEEumQovPU3BKfcrNOMXo8
jfsrsY3lW1YO4AbzdAaqxuilSOL9PCgzDZgZifctRg2uy2deCGNrVw5+vsyGb3Kp
1A/6tWZXZlLFVqopmcMNtd8TpMUQZtinS2eiL12P5D+VHHNujLJBCL+GdDTx+Ggd
si8Mpw0CF9zJZbwb7oL+YhRaOP65HF+SqYJZ1ugoKeJs6BPwclW1syMC/4+bJjiD
BKAloD4dO/hEb8P7gIuJDyP7qRFbPoiHeNJKs3yTH1IZmtpOLaqkT0tlLzqTTl1n
ZeVcV0ufYgmEv3oVZfqdcQOQncfKhIAaFE2ACNa+S0bQgWEPzWl4mze3CFhbB/Ru
JQJ16Jxy/5SvH1SGDmzD8l4qvutH0OFGvmodKPvlRAV804VfoBcl8azcEv3THmMC
7B/oEQDDPnOzqLNescnb6/85WayuIc3hFyfTXX7BQl6B8gfEQEINv58NhatFPnWA
Vc53+w+UKFaPhJLPEPbFhY1Ma5yfAw1SQUaBKglJoxfEifcOkFMKjPAOMJ8SIXlK
SEWf98+1/R/boyAjp96dnweiluV2Shy1slchh8TJuC98nn/8hzyy4GpeJomD4xJD
cOMrftBZhG/8MDzF2U6ln9hKqvHrlMNhTnt5NBak8xG181Mq4AjiDhXtbuHWOH4m
Zq3ruoM2YpsEavVY/pbU162kRiapsmHJXQPnHRDHHMmR4C34M4ysSNrZirT/Wf6a
bEurwwzOr9EnVF4Yw9P4sdmd7Ip1to4bfgzXwqKQDC1d+7P99DNcJB5YJV7rBliy
lZAr6Jy4b5pyHu7NMO/fr+0aqxyUscndI+cVmUb3FgJjX6uRKmQD9x+trTmdnmXs
sTA4iamjQm4xmUG179EdukAbd7sTq/DBJFiY4b3ROc9qFAexEv/Og+6S9tNVesIx
iZK2pgMFnb9zVru9s+hZxng2ySWRosojT5isgPWQzC/jki+FDNcuuQU63d1Vcwhb
sEIduOHpxmNMHsJ1hEuf6FegNAbVMOoLt6URLMDyMMfUT/6qkMxNO/p2EeXaerRs
WQ7djM2jWoN8aYZDSYDwYPPZzqljt0+mPbPKnFvg7u/3aAl7t9FVI4oRHajOxFNJ
umb75RVm9jfPlKUGlLnwoF+0bNnwjlKu8x67PbkaQ0CH3boYfuLmjlEam2jHDH+F
pTqCyCBau3XKAuiAs+nC5T02Y+a+Re+0arWU5LYUGuwm1b8Z4IRmOCVLzNKVdJAy
EnyQK62Ogg7cqKG6oVQtVN9E+DRylpOSxuVQ7+9yzoTvGDJEykMKhJb/nF1wWPwT
5FGF8rWn3ljNh0wW1iHW94QPVuKT87akRoRHbywm8OKnBc98HrzNelhwHZAmrBf0
y05EV3164ff0sCBvFS2s+OsCMdu1exGAuEPD1dtsXewPO9RlQeWLlXkmkFaIhlq5
xw8PdlZ6NcZkAxmXYwlrozjeW8bQv9/G5RsePkurQo4l+4MtZuiUKwXsm9ylMz+v
WAVYv3XVKaG/cDd7Vh8xO++3KH8f4JCG9nvmMvvjbMtJ5zkVYtMvyEGHpo32wfmX
L2o42YvSLQm/MS+/MhdqdDJPy4yYo+a4xpDvBo81Afwnl5Cwvr39IvVKXrdad51d
mrPYEa4IlM8TUi2O3vyvfmfI22hvpqxvrDFdockl755ehACuhjcFAh6e6sXNOyWa
PifrwWeCGS2UKOsGS/222Ek8j+6GvrcaPfiHhcRGlBx03/UWNMinyyM64NxC4GBG
DXqCZggRBKyfuTwQ7XrdDyNFbK9GIOcqOjHItcjXYsaAIibMNSpQWM28brguHfnj
Dqkvb1cwsucQJOeUqcAmhsBAIrVooAbTyqD6dlX1WEH6muYgN6wSe6SOd7o2lpBV
yIq8jnPINChviZyilGt536wIWR3hv5GIn3WWykNBAXVGF5AHWbpAAjFjnqHRzMi3
16o0rw1EMExuQjpMsACvaMuSpmZM1UQi6aXE0KDOejT3+Da0C3C6m7df1unsSPWp
QWqx3XBKWHawv3gvioeeGo2ZcVq0LUSStnl9wh/dHhGmPeZNHtevACgkmhjXWoUO
mWCEyl+uBDYP96WKPZkvzPFxj/8wYJUJX1Qx/021YMEK65GFY8n50Urg7G19cvPS
u0DG9zZ/3RtkHoxb6pRQD17sh6wfhCUHl/wPWbpFuFnT6ECOINkZkfL+fYPUZdeB
UJYewWXXf7qKewinxuLv4I3YzF4stnVS6KjqSsOmv2I5D/Vc5nLBkoqpZ/zBSil5
ciJUh3rDi7cgkCqHjYtD6/zO0SfI7oU1+/L98wCuphuVmDPryRdMUewf58UBVjtP
gTOhF3cjBjT1jQoftvh1/GIB5F6KZrFhd9NKXoMYYP/NBZHU5+koCPecIwbYk+LF
/K7O3pBpuM/4PXrxOAjegkusqOjs0qQKwCFC5Kk55j/Na44LyXE/1JngC4hjwq5X
OYRhiPZxQhmkPse8q6MkYzkUuSGk3MEFlJ/ewyZafBOk5vgsm8kwZWHHJcL83ue4
rLbPc5BZJpNUGd4LQVLj7vYG0mPYSIEOSW37qTSCSsE5Ojtp4Z/I1l93n0ev6nuA
lQ6Z54ZiHoQG0U8+B6lJbnwVLoJRVnJyoP266z14qP2l2yAwDQD45hLk0o3tBKI5
uQIkSrscq4755N3tuQnBzyqFd3nnn9EDIhj0Uaugrj9KwO9Dd4/xC+Sxil/2kmd+
ePj0Aku1RnK9tA5/zc2g/nD+JPVzUekgUSexHIVegCVsC5mS/BqOns5DxbjUYBTa
OJ4I6KhgAsNyJvaCcj1an6c+uNKMIQEgiD4MN2oj83sAtBMV8GxfiF+BlP76ehyn
tMD0SzCsIGmBy2ZUDaPveodI/fHGQIAeXduyOE5YYRWJJaaPZOr4lWYWjJFzh76T
rLdv1fMUOOso4qykLjie2Y0dGnhu/inpGlmBeupQLNhjF3xXnG2AilM+EzP1lJWq
JWoCp8E+ldMFRmVjVW3pauqSrWyyjgRh3VIFpz+898l4/TGAU2S3N2TJXubInUGb
R+QpTk3Fb0/ikn9WNPgfrWnXmzycplaEEUYZzxWZPZ/Tl57liehmajbzQt7heMcb
SyFYEB2WMeM0OiTFcoZcahVBxSQjW9xt0jGTMbbhZ/EFVVsbjmOZVUAYCIfbXKpo
VSl0OO+iUX9vVhIsOqpMatfyQWDfd98lCQ+7RMlzosLn0wmNAk6v2nLBiXfG98SC
5OitI96w100FlJDI7fXhgiGXf+4E33frf2NdbRQMQ6Fv57BPsZaSmw4Jq+sEamYc
6tVMNQLGgdoXcEVJF+eRaCo9/dEBly0/4csXkfoI1O2TyIBYkpcg1a7G8ZKlJfL2
dDh1cMWRFVE/7aTYzKVhYUPcoRiQAlcwyIAAXNFK6NR8Hz0xrH5LUBwAhp/2HrtC
Hl+t1QShwQG4JS4yQktbe6y3yfENhgi2g1JSH/nJnnUP/vaHlCsifjPDt+DwsNZC
zh+8DF2p7MVCFZP7H4GAc3iREU3GE+z1vqY0e6SJZhDN+SHbvK3+H4ZM9BjwkMSv
hYwCCHyuBrh9ttORobzQkqHQK5tdEdAsmKjWvWGM5O529RyPHMQ9Agpn45aPN0B8
TcVek2WjxPRH6ROCs3DV4g+Zj4SONRGJcxPnDXpqvCPMMXjkgszsakmZoNegTgst
eqYixqrwkCNmupx7jYSjKN356V/eJNHa0aRgRCNHRvSYQ9izonefbD8o68iBMxvm
7rR+G7qU8UiRHjzCgnI4FKQm5d+e5+hO4AM/rR+2AMSUX1z9c0CbbMD+ez976+7L
bj29Ji3gbEqZPJmEhTyC4KNGUpyZxyCJI39l1FMHEwc9rT2k9mfhlo6XUGzL62Kz
Dj5rD50a2SWUhqXHtbK53yhfan5Vx//+B72/t1z6Dk99dwvqPBC4/Na3zwGfZ7RT
aEVrlobEQvgHK59Hs0eGIhp4ymgjdEoKVNu6XMayUqYWQ4HYmsWynR4vhTpxArTM
xaiN/xbBPc+kF3uZRpagH9vSWIJ9p/rK2ejNvH2Zr7h2huVTEzTDyF8wGMC70Abz
e8UrUXdy0KVjAgwkxTxozzcfXS3tKGLWbBAYUbmixte7HxHmTl3oIphUPRocpBqG
YME3S+f//PWSzUtrOM06yvm2kLLO7T3jDd4B6TkIMss+fHH0ORPguB1InMcxdiEe
y4qyhACs5etrvnNoveR2aaS1RQGP7Gy2ubPu0RBpNFUW4YyZRqkGusE0ZnhXzh5a
N09zzklUSjowDW2BksANPOZZTlEiIAwMXzP0kaVK2Q9Fz+DRF8+zYYjL5kiJsQWm
LySlk/kRv75IfwfZOEndYCghkwHQUeL7hPejN5rD76BSoZxBWlbRrCRqTAQTfkFv
pmv2hzarM2oS3XNd8pXn3mfeJj/3+BrSh3cH1mabwRgCtH8rJ0YCOJSt34pzJwod
5L8LkF2ESMKQHFH1NUMjFORYNZJm2XSsAB5yjjpHjzD9OFq3EznDYXLo0vWmDVwx
xA3HrRD9MiKC9BpKO426ksZk9MpXhedxx7DKL+ELDBTzqFrHW1asQfYD76DD0QTC
KTuZD8QVFuyNE924R40zJoga5RURKBM64uBk6FB3nxwQeSUOBzDU6ub7cD9DIqov
XVNpnUqsTIb/oCOjyXRLgb1AgCxejb7t+OBkdHhUVce0UqgVrjiaRMohw+/hXbxV
GpZe1NhI2sCJs7CksESTzwyRorTnBH9nQC2t6jZoi6Yx4G/QHD7deo8ALMkM8AoW
ROPKdrY2CfW685ZZz7whpdA+W5MkOjU8f5yreuD9PoahnD0Z+QVDzoLSYUua1sJd
pYrJLPvaG/Fw3P2pcvlLdxu3UftCbGtNBcziwehNj8OCg8gqaxoi0JMzn5Gzgz2w
GDY9ZGzOxE2GGwpTlieABtcTymOUcCdx0U2pIfQ1AEspB0mjdGVw0+ny7o7d50uP
ijId0kI2HWp8ZgdD3Zda2I0Uw7Cg5gCUvxtEZ4Whn4TJXGxoKEHKrZDYT2j4uIQg
Y7W28h6Yl0LMX4B8e3gwZms48t2giNUULm6vaRccGylpuYz3CoG5Ao42tsVlmVtg
a4QaN8gWHZOXFaXndIAVqgAXbZTE6/6MJuY6DpNm5H2lEOFEDbjGPrBmUDhY9YH4
9ca0B5Z7K9LwEWBxuIhcSJ51zFWKne7Fwm0ZGYxngifLjNF87KKozUq3Aa5q0pUd
SpwjET8u+kK5NaMqaHaLUoLJMjDIeFIm4HdpVwSd8uFb6i3cnEYqz7m+JZDUBj8m
CgC/J1C9lvSZ3MwmNpX3yNJCIfpPtIHdZIBh3AZ3Z6TdORe2B7gNuWdn0I90BC2x
iY+j5xANzoJEKOVsfjPYuENiNouNE7aDg+KvlZMvxQNmZu8/sPz+jZbIJ/dOb4pW
HpSuex3T3+244k6Qv7J6PxUoynuS51y6l4mnmDfo9S6BbqjVQVZEiq745axVuQvf
8Ku6yLAL9UgW6etZuxx43SV1pqTeDv3/b0yVwYXMF9hkNxFRm1tCxm7HR8UnqxMJ
o4UX5bx0jXT46xmTyI0vt3d//b28r/2su3fGqPBXacjFZgWTQNTqe0bjQmG0ufo9
7cl83r7D5IPCdWjI8f+gEw3/t0WmCRToRQ6fy8jgs8ktvelw6b96/WDlL73UlUq/
DNOaY8hFLwLGEvV6W7b38qbNYWxO/OUwhlNXgoeoDdbGFhXcs6JG5XU6crUahn9s
tdTWaEyiTuntX7FgOUgLFb2jXhcn4gyOUKlHTsSz9wSmwNxmz8RmL1FsNT0++fUt
ygRY2W2ZBhLOxKxo6IQyfqNEhmIwlN/C8rokqaRMd2tSqf2P47zCXK3CYORGQROy
u/uP1ZTC8+9+GZBTSeijnkhtxo7m/Vxc9nC+cxZicAfqjpHclZ7vwcruJvNdDRE1
bpDHk8yeTix2pStE9NV7gNf57Gx41zeV5Vuzk7Z5VmU3CAT+dm/wE+FAMHTWJArF
A9aJl3fzGM479ftqHalVlHvnnxDW2zYAvxirALhoi59kIqUJNL81PUY8j6o+UicJ
r+9+EruOF1ELEcxjvX4dlQW4AbVTbwUETw0xZKs8pIuN8dzyK9NxeiND1LJyAvFR
PS45sfL4on5gG+0YsEiG63AbuC2em3lgc1/zZ/l+b4qgJVc6ncSp5uP+q9vT7u5T
PL+buNunGadPsv5TPtUzJepPXLtU42EUQ2ssV7IFLQlKpmQQIMWTxfE/6pC9HwAn
umkCQ1gDgPAYs/4SWtmh334Ut2rH+/7rg7DAhcraM8mudDoodQJw4xiB7qGIBrOE
zyPDq5YcFriy06JNJSduIBIk1C8ROfDLJSIkSpMaw+n6HDO7XPwuLjka9pjTPuQ/
pPtnOddbVvNcVszbAf+b+ZnrrfWCnFhor2ZyRe07hIpfKyYO74pT47Lot2GB33R0
2/CpduP4FhQ8j1gf1EJoI0izBjtXmksjkleu/rLFtisoh37LT0XmyTlOVZWtn4am
8FUl5xmeHVHwToZubt9lrApJrUcdl7hVbPs7HTc34K+Q65VWlDqboc/Bo5UE08Ai
oc9q/FZUQV4tWsW9J5MXqMGlpq0vEWeVpT1Q3tZ6i+Lsfp64Ioqqlrdc+Vj2oc6g
XIys1kZRGbcaR8iRVqUXX7U6aZOf3uc3OHfFEkWLx5Py5e8jdIeC473rkukMerpe
4ZUKUB25QCZR0OAwS2j5myAA9/QKBBUECCWUCyHh6+K08SH808Vw8jekOEFQB6di
Ws2E7o7cXB/bs+EFGyUiE+FMZ8s1EjyPbCjQbDy4UlSRcGKJUdVkHBI0ZKC76ueC
+BLgLBa/0Jn+UnDrIUOwbVpL5RIkhlBkv3Cz9GMWbJYX6lXHZjsULrEekUT91dZT
tmMxm788MLSEjyV0LoEe9or0Xum35QPvdwXPEj915WZ2F+1XDn8hXkYKYMkwBjGr
Rsn+I4BpvVIO7A7Lp0FtndDxXOJWzavHQllLcO2mExRLqlNgCNegCXZhSz06ABr7
2On/DkUPHZpvKY8tVTRCycwxtj+ddrhLLrbY66VRjivnSKGXLX5+rz6QLRl1bPY3
zcdg6t+9ilc9UKpiX2mRBFssxfMv+G9B7z/1lHNnpYqGJh9OxmCN0+9VnA9ID8RE
btZiPnyw2LtRjkJ3CRqAT83kCaVzqdm1heLkwve9BElEBTM09RJfchTsv4vPN6Nm
TwQrJrr3WtevPOCouZDFAOCIZBQBNCV+/jw3TO773WDLK+0Zo+XSfHm+PeUiqf/I
wNv7BG9XvaB9jFVWVyuvkB1sfdMJIyBaVnOO1lhveI71kZKJj+NfOJOE4YR7j6hY
haDnXZ2kTpqAO+8QFyhT2UMSfDL6oi8hysrkD5yLDCSLoa/wLvFTOripd4jB6hpR
k8zk2lEXa6sXUiBk0xMgycLx1JcemGPAU21FkeXo7owxrxQW/NiWipTcTHFrm8ep
A77odXrbWZ/BczUQxT8t1YQdxctyA88WSKlKsrPhK4Wmpss6iXIXwmx6xMJQJFyQ
xsB/LM9ed0aEf5ASX+iDLUP4BPPlm3J03Z1pEu1kkv2OX4oU+ILPHng8jUEIntQE
MMD5uOmhvfR3sl+9ZqjxU9z3KGvXFrPv0F0xGjDw0KcdBpxaqyohIIlOLTSFJ9Pa
K5VuHKCtdY2zzjrjRDXKWZkByBWFEmKo5DpMW0cgF6s+b4LfxWDQySVnFHsgPia5
SW85RipnTBha9PeFbmjNr2E+MxiYUBFUWxW9p5496JO8tvz4gwd2tGVvHjBFvLKA
ftV3rlWIADcHtlalUVHdK5t234Hos1gUrVmX9yuRM/Szjh5JG7OCSMEgFhrb3kVw
A70zTuVtMuXn2gCfbkajWRzzr2O0UTiUBagjh6CSsAIGbmSQeuv4X+L/DfOk8+bZ
tuPIGv4flaEnOQt2lbpHS20Kuna4CSb+oLyv4iaBntspUN6LoJ2DSTOrW0+vKIqI
8sCWwov7Q4loT74Zykfp1Tsgv15lDckWsZrkUNwWNeAx+lFCDQUz8+jW6uNh6RQ0
/EWdNhGj+jm34lhzpmBSNF9FSFqZsXyck1NrKmVlIfaRm+EkNyE/wYc8CCxCqzDH
2GGfX+NnsoXBBklWMQ3EbH/mmrGyS77veH43hehQ1qQidQ47ToRN8Le2xMSG+YPd
5OYPjuMNRPbMdOLci8u0AOKiKSKzrHEZ2Mw5qun+H2JshNbBHR22Bwb9w9d6Svas
fZiJP0pwFMYrffYEAa0BsQ8QGmQ7nCDw/ceKQgMSV6qIlIqCMjaQpfqHWB7cvB1c
npzNrumcZdBBDxWjYLM+vbTZ6i4BcLZn/38t7rsVUPwufazMPAzEGuOs+lBXrxff
rdISFRJGxvmMF2tSAoCuMTs0lKBCG6jLmDDxlFQlodcjzy9ETVY8ZllkdhN0r4dO
t2eI3wRDkXM1rREiXIhykG0b+TQOF1V4+4vhmOHSnjI1HMtm1MWowFO11QxNbu/i
Z//LoAoDXERlqqG7Mpd9Ko89lJftJqFFp351c0kp/+cpnMzF8iN8H0SzL25ltRLX
ZQKa0FdZLd3Czaz+1ESJ/JiiBJ6TePQ9I8BnHFsL3mHdGmmI4WIBaENmjVOyCZn5
eubf+6vQfEpqUkkt6yzuE8BOgxwwxiwEEWGZ+LkiIWbWc0ptW80gVIosNYk2X21E
Tcy5h0KYHQUDXR4fhHQVN1TPlceAYfkkmNVf7F9R6ter7K48OwtC8o1VDPNUEMPE
wm0gF/+e6Rqlr/VGq/GVgUynOIylU8qz2F2usSO/BIu/7fvYNYYxMDPN1wlv2EBw
fJBSazg367B9BsTOW5hA8wNBjMlhCIsfCT8XadpyRmC38hfBD3g0G4vony+AveTC
Avg+rwoTEgnMUyYnq+JujgmU7qVWf3iTS6J0wnDLzSX+aQTV198a7F2jQb1rHYs0
U50lVdOCaWNl46g0oqxJsKpbLq6Bn6RBxTzVMl2B5ivVziXW/foDyNi6gXlS4CA8
pTFhLe5RCVxgNr+O4INiuAlv2JDdKPHAbSNlluQNnc72HH00NbFs3wTFWYQryVKH
nHijNxwjDv0eOYDkJAxDggJCT1NfjbXnmbF90B8FMfZCq2Gp84fcIXfoA2kUVv1b
oELw0B6M5DA7XVhUPQYRaI9h2ZQ8f/61QZJPxe2pDtEoubjLzPafhinSMYMDyCTs
S+hBeIMK77nuApYhDn/XA6UYN/Hm6NIZHfe3hk6oOQSuyPliHtoD+2wewb37OtTm
LP4ItGefy5DnLdp4cp70hFvlONeDCZJunOoirc43Hq48xPSpcXuYZrv+iVInclAP
DOI8frMESMSR0zXBfpGBcuyAPBxmYpwNNj/4pjODGOqYntE6oajpvZ3TawpYhlaa
/ueScE7te4aqLWI1NwwACjH5ZflsaHUcQHdpkQYU4i290P2ZMhvcu9OjhtOjoTm1
A7dakGajImX6PfytTjZ/QEPXFgGceBckHQOTIArbf9SnEsmQlE3UZuuy4Ae0Hceu
n9Sv2o663FYe0etpVh1l1vj+luqyeIn2WRbKlbABwxOnfoZye/M61H6AuAcTiXM7
zhS6EP5eVcSCXShmwvGisFzWw3DoGLVOJqLa5EcLW7rN5BY9dINKswE+AoLfvlf7
sJOLnVSLMz631nnaqBWoZAEgCAyzVjyibRpLibwM+1u3Yi1u5fQw7lzb0sU1gyp4
HoOov6dKug7dhIRM+lTj+XqeYaYQD1AOFAr7gwRXRSOH/Cyp16gIuAXEwlGvOg9R
o8wD9NmClSXaAWML2qdzF62KbqNZMoGfxEo2dkM3MdOx5CbaNESs0hcuzaJE+d4A
YuRcpzrssft9vwuSjWfbPs9P7W6nDSiD9R+ljQqT9erfcYgDwvAJQ82h9j42rw8h
j3YO7W4xkIvrGNeNtcxSvlkuw0Gba25+6YMECBcIRP7MeaBa3t1FPMLfYTc8Bul8
TxWRvsHkgb+AGpMKhBTLCzqawhh1ckfe7CPqd3dgDUbMoHSBgTU7q9L1Fx118Vqf
vaQxe1Z44eT2qEdKel6mJ21GlnnUBG/HPsKxQyLPlCN803CUiKu/sJ+1VdxxOv01
Dz9ZxaIdTVuEe5MXsE8OekedxkXNQ/H8i6CUh1xUeonBDTKbeB5ySh4BW6wiTDpT
8k4yuoWCjRjkT5w1cYFcaSuLWc5BHEo7a56mlpEh6fxIa5SXstjO8Onj7RnYWojv
mEeR770cjmJ/WmjkPtEdXYEVybpbnsenhAi2a99Q+hkuAl1lkKNqRXlp1RYgoP3x
zOw/LxT3Qu/6awSSligeYbm5keZuCIlO2fpjH0+kouETdnWOc2QhJ9zf6q4ZkNdk
GZZYc2lwDeM2nu+NtlNPWWG65ZMtKWB2vlL1oBEZnTitLRyD0FDak1vuvmZyQyF+
ifvS5Jt2T45Iryt2RJBS0X8AqDk8hIRo2KwLsVh1apw8iou7mnXykHRSyT1hUwad
6dQxtccjLUpUyyImDLRz4rWKngVsmNkhdy7TWYDH2um1yOS8n5VTtIp/iygwyUmJ
yhBfSyFhDXuGCHZBiPD1padcPJ4LX8+2G+lgX6U307bvh2sM5anPiyo3J5xqQk0o
vfTaNaEsRqkyenoAZWREDds3yXci3diOHraWVJxFOkqmKHF0gowNez7xIhYfQuuT
WU786BQ+0WEurr2bTni3s3NtjZFsXnr5wdFGDHZ5Jqx41U0hthcWlcrhzpOss2sA
tiFTDTqhsWhIUpX19vAzVYVis1vU2DhSadTF547mYpxh753I8Uh3WiT8Iu3UQiZz
xEMgy5ZmsDucIIO2GGSOMI0cc/K4WbDph7Uo/AjhZkr2lCXI+CJ/0whHewZxBbyo
Es1zyaQbUUIo1XM/gNjm6mdqRS8YusMqDwOiC86S1CfpGOG6eE9GEZ2H7EzcMFO+
5akd5HyNjwYTnXHDmFcJCzUZJ7qyhORw0iP1A2jmaXxW5hmR8rb1gyH+pWBEZCwq
m7U/d0PVvj6VWnOm6C9JZkN8nAOGSdqb/PfVADaqZaE8h3tJURO7O/7op4UtJ1re
3bEVHWS2SADwlsN38hlvsOTAL6yOklosJwL8+K+QQvOvMPOw/NKpz7j/007Zmw13
AlntKJbyRYAkRSXXOyMCQRxxpm7ZVN4+NCgZaJWWNQ/FuELOFPl9MEsWTYHrmL/a
GRZno1jp7qJtv+d+V8XmNPrJGqfYShO0lc7p9F52Fc/Q5l53Ay13riLomEfi/LTO
Sn2tBhxoupRdIVzfeKjp95TWzfenXiZsFIzl7HjscIZwOQsceIr/TTiU2h1bfwEi
P7VXPWaUD856j59fBXounBDw7vCs122/nZm/GhgiwM1roN4JXQ18cFmQpKkaDi1v
VB7BhRYkj89lWCbNq3kSGUeCpcfTqiJIfq1qNBUJUNsc/cPhal4HxbV6mGhr6HsA
unJObQSSYRQuN509TYdHRzE/H1BmTMSB0jC0UahzEOsiRbyrsfQOOxW49soZG9/t
ebTUSCQDZ5+MDDeec89GYEJ32pL3A3KymURUF1Grp3P8+95+aUE0Lq20ucP3AHuy
yh8gPjze4OTp3pTfHISI7I76kWADWbDD/i3AMejzF7n72NFN6Ek+XGvtBcy/mGqF
3P9MqmxCcC8c+opcFuD9v+dkEQZ8kzNeKrctnWTQPd5/kMoAg5BQzdm7qNYUZyqe
IGk7G99HjTsOsYhpG0HyAe8foJye08Lg1eqALoHWKYzVjp/wo/3yINEG562ibSma
fMhbC5ickBjtoICKrRVEJjgREiJa8xjyOB70//3xPt+P5+6fuOCZMqwEZqpM/llm
eordXYDC4TxdFTlFExvVH8yhMEXucLu4iTM0EqMKS7/Q6xoc+QdUbwIAx83wOhOT
eTgB2+5xLY2T74igu+4v3mguwuSwN7NsdqpAcRuWsZsMNBN50emBoyibl50Rsa5f
L1SMmnKGmjM7T6v+yU+p4gj8+qm3ebxGF3M37X42pNNiRGnlxNeeZhCpIK48AjJd
CJTV7cfyay5A1KwSPAH828SYwB61zsLXGN6MSYfMKfNSgxaSXMwquKpr8YHrrkgP
M3lfpBDLGgbD+7WCavHEgKFWo8vOQ5CCKOBjKzHybF+tBh5a7TjYuHDH/c/8rWmx
mBpfHXjheBhG1TdEQktVqcsZaHVhuIAum/06SD0aoCV0KVr70KFk4ye9hgfW+rLw
c+ZMQy5xxIDyhQBuFFeLq35i9gxj4bUK/TpYHtCz6qWu4c6lpwuQjc2t20WYWidr
24zGslrnHscxb5Ijlk0uR8BTKc2gradSChhEO414jYYoMJ5naf1XW8NsMh+sprr6
Q1CQNG5kpcbl+8RACwe1h95gbFu4g58NzIo4lcVEIkUdP3uR4U94DSGPZcFX7Y1X
RV5vkjPXV91s69+65OncCCeBgIFM/zCyvmzRUJ0ifB14OtiGxGwI9tp8rQ+P3Z2V
NCj0IfnPmghPrRTveOf1OHC9fboTYfpN+6UjaWPuE6agvzBFAu9jziO1Sd9g5ya0
Mgv6A3XK3ft4bME7xSMYlhIiTZueIA9LWpuvvEpn/aCaHfxIrVH/oF6AerR2CZ2F
wxjwhGzRUcJ31g0T679qKn52KCKkv9iGadQHxrFCLANd0KRbWsU6jCUINQKuVSse
ecVYky/WqSAMgLsV8i1K5Srdt8texSFqxKgKjsbKNUE6c4/694OL8ft0PBIwxZAl
QOmLRzFKBczxqpKLO+z6lhXoBqrZRhTkyyBWJIOEYzFIHb46nKBBY6eHxvStD2bY
KhpC707NqZ1B70oPJYkNRbkPdxUIKWXUbWhsTY3LWo7RERFMQeeRtMkSBSTtNxxF
XSUmPb+uE6JstT9tfvvb6SzCt8pLoe9iq+WDt6BJpOJr5QecP2y5cIVRfHFaSNjX
4Ez71/e90Ahh17Ssfvhf9Mt+i1eLATKBHrJFEGg3esFsGDQ6wUXu968DZ5NmzIgn
ieLO7xjcypLJQsDUsxN9qQ6dnj0Ej8fEHJlDLZKCVCKmGikiiRVeF354ZC0cVA02
buLGXY6yPJFYaBQC+1qUb2xhcoRHjiaBvvs3kMZyjkjCzj0mva1WdVdTQ3XgcJk9
eNRZ8P0nfg95HpimROfiLNo78sW73nT0fuNW0eybrYIEG/1KNQtd0weZTYuYPEaw
gwSVMnB/KY7JxA/7vqFIVGbEYkDPe3QPUa4yUQOBtpz3BqoQb/IIsLkagVSlYx9B
PthDhJ0/D/a8eINAHcBI/8+/rAMJhEY9s90ggVENZq3DfAZpOnOadBfiBsBJjUal
KuSfjuehSTgS+L0kSGoMMFgL2N/67Z6kMmZLE6JUkgPzgiYCdqv1DUnRCYOoEkFc
FnQE3iLXy4Da+v5SD9WflR9BrD48jYvUvfOyUJy1/yugqmAWa7YKh0AY5vgyDMjr
EThfncgDOQ82+PFqr+XyYs/ta12sCCCh1pRbi71k2JkhcY8patu1tQBfUmcOjyVr
ofh99qN/E90lGELjvaiPKKpsSCOCHV7IKcPFvkdbi08XsSkR7kpUEGidkIYJK+DH
5PYofkblnnov/TiDKjNfYuL4gk9itoLLDBIDtvPK7+Wm+iajoKAu3UZ1bMcQ3mmf
9Dt/q5f4UuBa1iFfziQVzoC15venx69P4KtBXMUcsrC0OXKuNNe3eGNfywbLAL6P
aNkhe+4Nz1k7CV2BI3BFGRm0AyPhc5JI8xDErGgx0RYB5lWyvkyoRwBWnacxjINw
a/7vbADEeWPhDyYzyY8VBVhSUOy4QbHNaDlksi4+FYGaouSOQkIDAfgsK+mkPGuX
eK3cSd/wVzSOnaMImdMyDNStB0OzcP/M2kRIxUBe9KNlC6JhbQSEwegLWisKYiCA
d9oAv3rKgSVQn3hFqrheAl0D8LxYRfrl0EWIHnqv8CSUdNVjEaCCG/WdM0VJuErq
8XeHTojr/lHmWlQTxS70pBn1aSNcTtMBGNsjAashMxxdfm3poruU2kMiZ24XS4Or
ms+BWJxXCOkPdICJpRRvjejTrqtWqZQQl7wRHv6jlJelyYS3S1CCAVqPEaOXSWQC
EW/urmHMpFnhiWKKZJTpe5YDSBOEURpYv1zqq3jkVkAEPNwnKqOBJuakDl5MCqgA
a0hM2FcN0d/Vh3Sqw3MQARzyfm5y8B/y3NQv/C1g9cY6bv/T7+rNmngzGROR0iLH
3VY85gX2kAkcc1HAzkOiPYd40Y3nM1U9PitUH9TZ+ct3HHNwjHS4N27HkRK45yju
1NxVynPHuueKESaMt92Pt0vEekdUWwFjswULk+6QS59YsJMJsSA1VUTvGtjkK4NT
wfOekqjdA2BIlUqLqneIHC2btFZ9kVuSIgi1hNPcdPW1oJxmOt7/V19TuyLXFRjl
39PAr/ckgersVQmRHaA2EjtmUTEG60aofVrC3/XaNKVSMISsSCLZZv66dqjwvwNK
FMtbk7zLFC7CVA/8zt7hd2UNVjgIO/latGv48oBxjh8ymyrrhQHxJEYoU3K95qzi
wsmFg4Fma6ieIyec1YL4ddPBaXcQzVWf1j7VyumriZMNEdc4uxHsvwxVCCcHBVW0
izFvW2OLHbTpSNLOaV1J2eUxWzmkZdRmW235K7dIbSwmAKJ5/Evm8z4hCZl+6etC
4PHMwdQbiFUoAr/1d/ptrmfMKfZP9rAc0+t2mGwexo4O1IamOjIKQ1g7ooe68uFm
7F1bYTC3De2lS8GtBJWCxN71yhc7g+NP/KR1ursYp6dTP/DXJ9DeTNzxDHfVM20q
/vLoB3BoPGaBjw9ENfXcQVmbu+na1cGNLu9QsMerh+hRjDAP/HwQ+HpW8RGT/4+B
cM7lja6cV1M5ek97haWNry1OAhcJsLjckK6ZPJg7vto0hdkDZCSHpeAFoxHkzJrs
gYmOg4aTSX/Gr+7e8EOQK3FU2u437oWkTmlS5C8eXIpy8NC1kNwP9AVOBIOuC21B
D1OqC0jzaYVo9ng+Rk9+buIBCZAHkYDMiNbGhjfKICpnpbygTgO2iCRRcLMPy0EV
/abrsc8cDxvHnz1TSQyb6rxURcvhGL+3m1TBDzkTDjGgdM5N94J3xvWvcAH9Vo3O
ncRDvAmJCvapVxZefgpL/CCe2sALBQdQB2eK8s48ABx3M+8VOrp+1oIP0r5GaJZM
lTSZPyBROLNd+ZP5njSZyRYL2zMf0lNfely8oh0B+W89iEIJnf2GC++mHZewXVMk
KQTjW9nWph+8eDacDlelvPMykAKF7wmqNRrZkU+p6WwjQlj1jGtZU5eI+tpx1t5w
urW61D3KZ0aTKrfCv44ciNk+n/nkxthZjKuV3G9lWTTxGy5Q0VWNmwZwATMakPV7
fhe4shYAIQ0FuzfURzrahm4PWroQ2E/b0MWIEtMF7XJwrex5nR904cEUycAbijij
A16oB4YYh/4tgCoSzEd0+neqXtDqOlZMUAt5MR7s5fpDivRdqqz860zduzu3Eutu
XB3HGZzuPe5Ok4d5iJLsIKG24kpwazCZjJpP5PBSGuE5E6W83TLi/194mf9WPfuO
gNDjTioyiil6v8Y65UNrcvzP5wAQeTyteLKVML5xliMDeVIKhKNVh26zReNqfOrm
38OtFQoWuZg5qqQFW5A9MYLPbndESVLtz9ustga6PSFF4UwlQWT/Ad+1JhBRHSr8
DvJxqy3m4acinx5oXQDERa3b8hhZLymEC+ZwYzyqCrv35tAhuc74sRkckvj2b0tz
a7AakTw5tNiZxiVR5a1+1+5ScBvK+hDJK/cVbvuz3LPpZjIYlakpfIRjr64aEmYS
H11q11zIuzO5n2aN4I2x2vMgYulCnGhH5DkiW2ov2UEJMV52utvgucP/EwtBJ4yR
wucR8yVg2HWeifge5mAP6h/v+1m0QWUFU/GAWSEttRtsZdCzppm4gRdPMfTvDqFb
QF3JzllFmgrcc9xGSD3xFV7/Y7ZB92bVLpIaRmhBQYpNXB2JgSIcctwhmW/cV54u
X1RAZKavnZG59CL4VG8OgKuOJK0bwTSOaQlDQ6OdQH7088+QexjLCOTAx6Z2lRmT
6kzjhUSZEVDOAiBOHpYncPLhha41CgskOJeIwe13cnIkSi6iy0BNE949Aoppp/eA
jUfu1RwqVrbo+AipuS+mM7dNrrPlYkXQYEx1by2KuyUsuQV1aI6uB+MR3b4yc0aI
V+ptCvACsYdvVpyCcv8RDOdyH5NSbKvdNow3rWMZwf7cxApgyXn8l+sfy4lIuMul
nSsuU1plaJW8PhZm1j0N3b3kYEK2ihMLxPqFgPjlYXCLn1FR59xWJ9Flr8DhmW96
VHA9zDgALXQDMM5bOkOTchGxlMKoNtUAuxnOtSLKrdPn0mElUTVWa3U5ZkLhcuBS
eHE3CGzK1oizYxZ9xINfoZ8TCg6pHLN2IMkay7ayQfreeBNXG+2PxTBURTEC+tdj
/2TWdBByahxcR5Z85sYMVsaqg+hZlsyziQPPOPSHZ9EKsXRlwDFut1IQuGJQggTP
RwaM+YB6URjrPOjRR3K4vdFP+tie47bW7G+XRsVwHWftOP4vBLblBbvWc3wlJjLM
7x7t40EKhBLaxMWLewYCnqJjbGGR1bKJAfgyTVAtqsLvaCtPJidH3/Q5LMoc7WVC
aKwMJI13/gHgc7Szp+EgktCTM0X3my7pXGm0ejSVCRgYGNmmUrHHYCxbtyiSYWv4
YDCH2OHprKzVFR6JhiMAk30uk02oxZ7KST711mEmdPpiqzwGazuRM8Yf6UvdTgNi
t27sTfLDDiWU6ESZPNqbeYVdpT1Tel5JDMzjYDK07EqdNgiDQfQglpMnkRcFCK2i
t8zSl8NNxgr2x6jvFHStVzvtBAALRufisxbexw8qwQhWxxW0sXhGEDNd26LRKMjK
A7uRG4b3HlP99rGqRpxy9Adt0xqPbUA7P5quEUGkWGkksrWPFn0krJYdEf5NWFQw
UGC3gtqaKDjBVfBZPH+r9iMad/bMWqT9NSPdVK4glDoHEqYHFn+f7SU76gV1EUHq
eFuWnhp9aTHdScnJUQBER8a2qcWcSVprvlG492QV1dLF13VJ3v4fqbjOQnXvQ3Su
SPSMENtWLRy964mdd0hztRlBRgOEanhXshYW7ZXNt/rnWBtMkeYb1p8vPiP5nlB9
ufbfOx8efwCFHSV4wrW5ytzUWUh2lU2zOKkFHA/aJrjrkAlPJKwD2G/m0/nrJ/cd
uN84oEce18d20Sm0Db9rBaZgZ5NtSMBt4J1NpPJFY0i6nPYiA9WhAIVaXCopwX9S
7FiTy7ikUsioVB5PSUJjIzsVyon2KZ+0v74xRWIwAt+QsqUxsyOlSb4bHWOpibOz
07O5S/K6HOssiZsZwWSxqxAt1JQ6p18bfk7LsvH6NFzr3drLuAqFJ8JihK7HQC+Y
v0LgZDIrWn9ZmeslRysvqOo0KtBCpd6enHUXO5DyafkX+usJF5qacBUJ0F2R04iX
5mrpM3xn0/lLssejKXthkDTXF5pvr7gV6cXE+JVwaN2qj/QGnpI5ZtkUNzS4QjM1
ehHLrXKAu0RdHuvWoz74DWjlbOpQsk2mtU9QtKkTWTGHcHRSIKEDZQxYrkr4OMqC
aXkkGDoI5gCAy34ECmJbqkY3wOOoJFeUI+4gAzBLQJjTFJ02eWU6wtD5LTUgeYEW
sWs3TQyiF1kt7YkGdODhtyG3EiIrGWcMft/iyQa9878gtui9s9aFMBh6dXQRCv1u
dGuvcZ1DNn2HlYrD73DxSvqhfpdr16OiigMo+HpenIZAvvQaRKmMp1drowfSXjdh
+xe6bEyxdrZ2izonzuWildwheTjfeMFmtYOAr+EYCKl2HxDih8Rj1VqHi1M5uEOe
rhS0qXhIQV/TM83yxIsPc+ro8cJh8FDb/9C73Mb0hkDQLfgmEpJKr6XO2timZ+9F
30tWdCWPmPGlfm3tnWegBe+YKhxb8PWl3mXh2y2qYm5eBfrZKeR8eDXZH02j+Gl5
zT/2ckyYCK3U9XDQm68xO6OZExT3zr/lyOLIBOHT01vcui/NV3RzEngFP7tDZqzg
w1f6I3NTFzJ1S61SsmURaoXr/W610fJwKe2PccE6iFyM2rijqUNapZbW8uA5HOIx
b0HBD7xvqPaLJrT/D14c9HWO8gNvpzjFBvSHzXLmzdbzjKWbQTq1LAXd51tLQgDl
EnqGn/noq+A7Q4ByYmqayvySwGtGRz8ZBHh2jEt/+8nMm/+Tqt+pYRBARJtX0ZX2
S5ZOrWvRf56iP57fL+SeqwkFy26iZIZI6Bq07CToaOxDzbT2xDCO2xYCNZRApxXD
EGm7LlfBeQRW1cysMJwtU+PhQ0eNUGpNyojdzDNiC0rCJ1jFr6D04GpThUHFmsX/
XPDgYR4Dot/9CBULXW8wBSuTTw/woB0akA+NapoSpSl+kU+ImmQ/W0Nzk0eupklx
4I00MJbMm1h7Y5H63+WgYxAaqnDhhNRlDbV8WoBQeKFz6Tf1GbfkRk8FHM/A2xku
PxRBoH58qPrZTiCacINWXxJ6dUQSC/t7AjkCqy93Lr5GtJXfb27OvOjBa7DcsT60
jGJkgbD0/ehaJUfEtgCglrzDtVzNSTD8ombBgYdOZ1MnVGWO+VJdMazvSungdShE
46BmRXKopxJCokGHK06IN2KSjBUqT/JxWCZ3YS9bqe//phgwbeNiqQbvkYTHaSgm
Ty0XnYWBoP3DVlEIBllk3cvARoyvx6YPYBEmJ2aIo+P6T/Zay4TBlqKtGEBBnxBt
6IAMxh62RfNA31RrGYxX+XKqgWcw1YA0iJW9AJcwwsRKWzdZn9NjFNon9YhrIiJt
nfIbzO47mtnLzJFT8eNVb3anTEDPjwxIRs7aUeI0SEjxC1UlO8CtR/SDtyFmE9eM
h+sXevdw/k0SOHmFOPAJmSQrt9zDTR35KjMu7eBxeAyW1BMT/ibLZREtXbAU6Z81
7ehuM3iZzWq+gjSlqBDx+YnPoGCqpOHCxXFQjGcG1IBDwGUcV2gI35crTZDfEYEi
qKXOqHgTCyJkOZBWW+FrlB5qZAMPW+MThjPTuw606QL8Y+1obq8nsDoeWaS6i7PZ
F/tX9rB6L4TtGxvni6XwJlz9Km9ucVw2w0wZEJU8vN1cZiv/d3JUR9LXHLUyWUML
o6hRX2V07yd0Ka0Sagl5xmqTcNKAtqFzFch3B8rfYfh2ysq6K6owmkXx/0CBW2kw
gEWsuwiNmQHZ0bZHk0OcUzZn7Fo4u2MSts1mxIfTJAuDafYbPqZXoTBNCAxGE1N+
ZZ0t2RmmzjDS0i5E/XI9v5OFtbNFI/rwHRZaRV/uC04gH0QUM54+HcmR2oVAYhVY
qdl8S7r1PfTAWnB4Y430xKQa2y9661pBKkjVRrinJ+tEJ72Gip/62H0cBBCcIh7/
B8MfILvnRyXGLEIfMkZOHmHXE+GlXUrNXV0bgrhrywB4txI5iDSUMEtaT/dwl9lq
mpKfeEq1NSYcxvG639N9+wV2HQLRKFM7rQ7DwK1jETFOYBRPpLdJlyUa5TcG+IV6
r32Ink6nQjxnIaSxoNJKcIiJKb2lowodggOGzoX+6jixw4iNFuNRZQ30+RJImdXo
eNpyaPoi3Ic31YVKQSGl75sAiSoFYKt3mZV7tsblDeyOFIUkypCckgqoqwgtm8WG
pOBLIING7ELd5eRIYuUBhQStVqaZed4f3KrXdoGYMxr2pkhb0qU6+bseTllWrGmV
wshzly7M6PHW/kBwPSfMERjCIoChfwlgmq3cHluTTIE03lr+dSi0GFDToJN/D+Ev
0CdRugF4BbfqIrex55T7ppCRFKVHcdjEU18N0G9N+WfU37P+jaMreQaYuIth8IPd
i3hFjjho8DkN1WdcIuuwHUVQg704tRTAJU0HW3JfFVZBIOUpV+uUSsFlZOys4xQ7
gmuesXb/NdI0OTQxDj/AYNdqZq0zBNUiq03PzovV508xCyYnmHOjUUE9YONwRBGy
Ce5dKcIIHQthiktB6OutWXzybumpNyOJlTnDzDRpZRdopuTo2sE74YpoFEKUMEft
PZm1DskDVc40tpIGkKiodSeFtTCpuw370FMTbWbEo3zRRoOkq+SpuFiHRjZqFh+z
EeqIXFN6fxHAV08ihorR8Y+Pkg3anGfMDMGAP3Nj3d5naskWyhX52AWSUmlNbJTZ
V6OBmPC6LOdpv+xzOyG1s7g1IOc/ElduP86RshR7wrn5M4wRx2XlgmsmCPyz1KJ2
kmD1YRh1cu1rgLpANyy4shiBFWrjPtJs1ZLgaziUJ4pvx2l9l8FRhJGlb4Nh45jI
aLSejFql9xxaVM5nt53fInpjtdZdFsd/a9j1k9NP/sXmKjnq2yzOnzph/LiGLkw6
9lTZpcIFkuf8dQMTxFqb19MwbVf2u516Yl4aTX41et8oESXfZ0IlfQv0ZMIcP8Rm
BdcKaB0j4HzTjmSmHeTycnHgCWaWDTSi1uLnS2jrcqSqiw/BQ4xQPUq4ZGM+y3v2
6UY25aK/7GYlgj1q/o7WVsV9Xpo8tkHY8A2+ON6MtFEX6bL0Tbc5ch+MdZxWuv/r
a7lD5+CyKZDAZ1U8xPCcUC5QOcovX0D/eEu1i/Ddl41WXEkee8ASArgWgd+nv7NF
2fRC9ftKDpS4wJkms6ZuWLwKzHIsQT/VHxPpeIZF0hNKYFkriEWAGn2rQc4f3NbT
RUBcmZ2SSat27rZZgMaNlics6Kcmj9cG2i4KOkLciIBcy1MGA+/7Kkk2uB0bNpcK
xO889+XsNlgl2m863oy+emy4eKH/9KSaLRQJQ6m+DLNMwcmxXgIzJbN/bAMVfjQW
9w2m9zwGUac9C6we9YfUDKX8jPlSDQknQbQIJTeDKq8ifxS+Vw8XnF7/wN+SPGeS
wnWFfArAMJpX7QpX3SyXmxcoCGGsqWQUgjgjNrcC52gtYDISywCmyw1+NSiLdr+O
GYhFQmERBU+XtcUkb1hHitkOsYLPYmIpUdACmpddEyW5B8y8ABZIXkE+jEOUuXTK
PVu34X95jxdcnw6eOSssY2S3dT1XrMdYBWKEf/eckcxUbbRXM23V3LM4CWjfnMaK
gEUqIJ2hFJ5Bhc0Q5TGnocEyUtT/eDs0tI/7NaMZCIhZASns700np5YLmQ07aoI1
xEqZwau5Ov7EwGjzaW9ZkPjdAxaicikTYDlDoYc2Y/kFKO6y9Y7j8i66khzkssdQ
GWP+RAKoqVyuP2+QEInRyd6B1v34Itha34fnucdSJI4ya9/znLbXz5c+W4Ln+8jG
UecFyl/qMq51/FAzKtyeKscQMZII5nvpqsGI5P8q8Abm1tqqHnPVhCfbB4oOgaqc
/PRG2mre4rIKmJbDEN5/qCscnzOf5rUyin2Us9Vt9fMpJ9P4PFiIppCcatyZ600M
ghbAX0PKC9SDmeS1LxTUT4Ii0Uc68rEWvsTOxZuZCE7MeukSZM+RHJjHZWmCkKAP
KZoDaHbAzpDxGmBb7SMtMlnRhTiiwBSRwZLpb/PRNVZ8f8uag/wxo3XArugxfEqH
bs40JF54/PTA/Y2J9RLQjQ+nWfuGixazDIrTiLJ8icYj3tLEabzGPCTUQHNXj/16
Q8tqKf41+KPxQMnC+LYDrWMGNiG/e0NbGK4sMOhh6AUc4l3dtIrIIcbBCa1+S3Qj
Kb9+kpUfhzuJHa9ZGkug+QFi2tCzxrJTX7wpZM1cRkorWdep8r33fDldUjaXgdrW
JqLuFUrj8EFilHiHc1mg48vgish6m7OQcRtj0y1ZPAvadp/GEQiiS3ClMRnrm0XD
iQBp4CNYnERxP9i1sOBDoxEVgfeGjeBodr2ZqIr+8MvRemfuxDx9YPjDvPcrUZCG
NaHYk3h/E3Ws0Ov/yulf0qqlyYin0Iv7+3weH/drl3EM8Wd7zOPjgOREITT9Qltq
6tYo7r2ApM9CSiidVx5FpdiGQmkpVmWv6NYtqqcsQ8KdZOegnFf9ZrXFE0X0lD6I
5fHUU8oFhJDfUcfB5JQ21JfntSbr8EHmvQD/ecGv1KqJF6twufdBoh9jJ2swjdOr
KOA6GnGiyEi6n8Er6xdTyhB3kZPa9Ma/bdMYgKg6DORTFVsHWUzXt+SmuN0TfKfb
foI5qsVteU69RdETZYBtu1WL5r1E348e/k2O0iRdhe48WHRhkeUhm8IvQPqxo+u1
5w+HBadwpyvfroTPsakjF3rXZDxatHPsUuP8S9ccNocYnXA4wsV219Iln4BuSZjd
DT8FWuy1GGi28XhgVNmcf5Hcj+Ymw/cakZ8zPZ2SJ+fiOlwwMMGZ2vfWsOsMePN1
PYqpXM0Fr/gzYxJ2cvlldvEDPYQnh7WqTub9FClCDrMhRtXy+D6JLAtaZdj+8+jf
qDcjkeaLW/eUurXVy45qmwW08Jl8UcXo4tiQDWiaZFmC39Y8hdrRjz7YMjyR68Kg
7GNpMlvtg2nMw23PkmcNiopk4T1qwcbVHkDBBsK0mslPvmF3j2KXJm/2X7XKrHyk
TQ4S+hOXEN5stCfSjpM7Kr+tpYkN4AF1eBpIMZEhzHIkMTyMxO9tFFmGt3w1tyQe
u5aUyfmncJ0CCCxz5nO7lfld4zD8mAdDilZ2WtD62p8OWaP9E6UOUQF+ByWduhYs
K4aNbkQbrZAphsA7gCxaysFPa+RUpBKTKT+hhEPa/sD1nTxI4hLqD9F/1cUTu1lt
FFOO4wFjIzWxwyQiA9iLnNKUpBUFDAaGKwXB2JHCuFy2PzEfyUXX2cl8GLeOyJ9p
qArFSRTkD34GbuucnTSLaudo1aL9iQhZSBJPuZXhuF5bhsNQwl4zHpEXnR2LcC7T
Xbo4oqte/BcyGnDR0dijU7e57I8xryOnUvFlQ9oRMEFggdh1BnLYtsl98pyjZj7F
k+dJyaLit7UypMsany1n+holcBrdY463/XlInTTZO6JPUOa/B95A5edJ+IA9o+rK
c4K3+SUUMJy9zMQ7lfFtfPKQ38qiOY++tW51EckGkhll/zqWqFLhFiA4ug0Pp+c/
9CeQkSd6n2JZoznxh0EerFMEe9L73t4VIrl6eVpOimf2dVOjr6qUYAnbho5wsYF1
Y+0xDiKuON/JESdww+l6G5y+cRC6wzkJYRDaxGdZlIA9fUA6dQOF30Ej6YXaET+8
xVEru5MwHVNWXC+7UBvywDLZcmUXknFU7sjDJCWID4TTut/dSUGUFBnevXD6nbK4
Uajx1ZQ0+h0eK4nyVMw/wXYDM8Mm4yTllP/h8eQLhwBkt4SOYR9jKhuqCIOKmRYp
v3ImgWUeFjs5GFGdL4SuU3Ix0DEnrhWkjArRzg8uNsNoGqz8+5mvjV8RClGhKE9n
bITVNjor+uqbrnpMa8nbXiZeWr11mGxYRq4Mw7EzCtOiALP9MgwtnaWIxk7ZGnuu
dN+on1avjv/PF/ZR0wDCMDh9Qm1VbfHY/BpPG0b4DY3J/YWJWnChHVzKKyDRYGTT
SrXsLXGyRtdPbUr3gXcs++CwqBuAHlRArIMNugykdb8CQ58rvHSxlP4ZmMPExscp
ZkhPkb8NmSeO4TyMf1EB/lCuoT5n82psgVVSc39vG24y8RAqtWsgpMCJlW5+iVl7
mh6HdaMkCAXW9uHwMr3QjWc02cs2MW3lmjxezyfIVR5mH7MxGJ3dwaa4VdzOnc3x
FJE4B/gv34P+XJpiOZtkQjzd4Z+/BZay9KFEGB7Rh/HbcI6xsCg4LErCdNpVG88L
fFkCkoXcVcxW6V3s49bItpmh0Dam4IPUBF32b9OEmbqpV9VH93eJ2rYDFrkx0IxZ
Hr6uqKhcGOEy5Cq1Yo4QtlQLW6ndmXTimS2uZeAl/OQ/3nfPyaUDp0YIFf/BoCXL
w2G58Ds6ZKE9kCIyvb8ZA7ZeNoFHQ/K2PuMjbEnyx3hitZ7yyA4bTSNr6zCAFEeT
drunjdCsGbj9MfZ6vHMG/FB/LXPD6COoxzBxRNMbmWKcsYjFO5TFQDtWJaTSMWIl
udPU7n/IRgRwrZCDMAU6cypOVLUOUoF4hFXyMNx9mxdgkBE2MSAHiUUDUcGueyLz
gTb7jeTRH6ehB6Le36sLawQc90/uRwrsJqv/WZobqKCIP3U5MNydxuRe/o4BrHfC
V/RFsT38ARPO+zhtIHxM9MTjDDDf2sLRZN/ySCJpT46/gY3MbQQzr2Xpl7gQ01SP
4MMdjBLmOP/NFwRvz1H9RvfN8lRMfLjefwkWra6EYRB9Ok1vKXVO4tqmLniq8Rqe
zBKxll8GhwmrIwSJxaUczLHYmPD0TOQ5+B93UhUw3Oc5KQxyQXMd7C0o/0ZnLJRn
dxm6Lv0j6rCp5rfqjAgHHtkr0JjD1WGSLhqB7dDJ6VbP4bOm46mEFvTsvg2PR9CG
hAXhOZrsenBkge10xsP2BqUNRYuExp8bYjc20DA07LNpM/0/AsS1v3yyGtUUzn8L
gEEwE8a7m1sA7/lenOuM+96EWw4UTmX8I9Pf3k01FWbukiaC5xtCUuEyec0oNR1G
3TtHfgW6hvdhO+jiGjFrfM3iL5oZGhyTklTGchM/Sh6Xx2PK0Af+ps1z2y7zYJfe
qJUOMCdla2N6MMCz6BfHLt4BZIamq1oU3rMUBUxk8TibwkuOuAwdRuyZE5Db98RF
7lzdy6hIZSTy0BqviwBwrci32JN3erkjNPY0PLKPKB39sHrY3pJoi7w/fHSND5EJ
GSXk9HrDYDoShgEbODo/0ma32KYh2j8D/4tFGhbmxAC2tG5l4oCd9j4r6kNmOqww
JCn83h+lqDNPvqIVaD4SwG94HBQa8dgbkpM2TfQnIS/0lDNi4tYeqJecNaXpIsWH
ukz3jZt8TIm/i0TYrGtJ4FYZ+64U85E5p+5DchQf3P1BJgyknE/WqvTtSCJBjU4E
kjzxDN+hKWt1xQzE0LSlSB03GUNpYSThPnvbnrOcCWatTvMA1l0aDQHhEiCQ0Aji
eKlKfcd3WuC8yri/bbs8AaVZB0MyFhoBCSEe7vryTgZhLGmb/h3gBEXMBoIyR7wx
7j3LZsNqsp+/8X82hci+6fvpQr2zzwOXF6o/eh2eS2o8dMOJkha17lYT4bjD4nca
g7iqi8bxwwOer8G8oUtfSaKFKFjGPLdV2HGY7eKaG++iEcwciVzKn9YE/uKx2rzZ
Su9SJ4mJ5cxc5fngIS4JfCNYodnfWgingcBTEXP1Vw381SIM2pX1xpg5vzaIytKD
f0i9TqkgET9kIbZR+foRSa/0umc78Xq3W3oS3FeqOQvSwHLyjbihsBPxSmFJkVeR
8xTmU259QidhyHVIS9LLYiBULIWR/Xa91BOO6JxDBoIRAQlqKzyhiTbjfacW764q
XRfao9jNhwWsmS+Bxqmcy7k7M2dWnnbvbyV9bNRKA+NKeRv183Jx5cbNytFm0Ezx
NDPoJk0QUQ4EtQ+SodNaqVjOiW+4Fqpkb98Buyck6mXU2sbaU6oSOBwcZEgJfKzg
EZYL/YL/wkN7/x48+OrCqqY7JI813DTi5FoWhbyfnTDwvxcBoMTZaoMQrFY85wkG
N9mcbHqPDq7CwDRqUguAhwsmVUuddmR19ZnwoGdmNPDQWaNLjOh+hBsGqXmw85HK
vyuDvZOK9MtvNbtpTcaHI0A9AWuGNAiN2cK9VV23YtaHsu2sj/FMkdhxD+J0rP2K
gWwmmV2+9wJC9s2bAm09oi4JXoBMdQegKKjUgfLLgdJ7p058dF+NLsUui7xm4t27
b5Clhnsvf4hUevoky3liPBC2JZ+saH9AX/Wr6hUVknMLSGWrZydbYI7OJ42bYo8M
Hdkd34O4XfKyRhCptzOO72S0rVzmjgr8dhu1HBpMtm4fL40PTxQOpGJMPVPyIqNM
GZXWP41XD/JguBcI4Z0DwefX5I0hb9kzJiO9ubVxXyAxU2CeWoCnSrWG4/gKvud6
Wn1TY1Lhy19cH7e/5GFxfB6icWoZyZly4IYuWk14IB3bELDVgJk02wwBtJOf4sUs
UpfxEDw1jhtCELWXOZsmEYD1m5X2RspvX1BMPuvDFJYJIGr5eEVuj0X/avnfDmLV
r96aJwE7Dqqze3IwSEygNwUWo/AYJ6hORZ3E3TMRWJtoN0MdOspFkUB3rVby2uhW
hrrETlVwZwDe8Exiulnss1ZGSmFglp0u2puA8fMsT8HDTSqzVv1VD8noKUBEck9v
rcaC4r6PVcMFYHatZNLoOB9vD8LDWqWc1w/jaMXlD5qUVq5lxzGh3g7xWGdbvuuO
AHERMt2HiH4p2prGAR6BZs7S+SAjo2qanG68TmfPuCIRRBWwmL7exi+lMCUyD1LG
wwie2pkXbkw5xwzdKgUGyPQyKxUnWwPfcByqA8+rfaale2FqvfcGJXLie8Sn+Etj
u8syfBF7Wfb/X+2P/oBYNngZ8ncjJt4bD+UYGK+aL0t10fsTEbApEsN7WMHRZo5d
mGM7SRqjtd/hSq5NINlKQIpjhmz2c04YV1b1UWsh49OT0fQoMJ7x+hT/h3wmFFEB
G90eGBNtabyz2ctwM8sOZF5++N8TML/knK9vl6BTskOVy4pmCy86Y8h6hQe9lKWU
tsLGX+46KGyr3pz/1Lpyq9mdclirUIzBtNZ+m4KIu3SpZEuA7icZZVCOpC9lGELv
OdzeSjTRBSw7d1190HcfJEb/G9o+Le4Ik5xZAcNS/scbMNRMXTNxTdf4B+IPu1R6
iOaJfJyJOMzpSrwe/Qbas0kdDvbWvYCH4RCKauWgwmOhEqGQD1iY3UdHeKCzmPxE
iD2pH2TMbo0ZHhzu/D/bWLQvBAvE7ShennTlvG1FNsjCqgNzI97sxmCP+wLkWN3E
mUIgWLczr93ByViC/jNgW0uGJhwSyYU9gAZ9/ktCsQhxnvpgPkBmgc27rKjhhsNs
WTVpig2EAdriz8cIBxLXH1ASikIq/6CskUwdiHANXppFLl2wt0A8jiwfX7dF3t1t
KKZoAnc4jZSdLVBlLMHDeY/prYhcWU6iAc2UL7VqxguUnOQ9MXO3tiYbp22qPQBV
ih7o+sY/wrXJFeVAa/kUj6VZu4i5rfKN9fZixBoj8G+ZcO8ExQYt4qwJ7mBmRZ+1
QfVef8KaSaO7AW14YJiuBcQ/O/R8qhSN9VmGiOXvSYgdmvj10QhW6Ub8TJMA7RC+
08wmjbEbcubVA5gxChmhsmAzlpSFH2ZdEXYPz2SvuUyfQmPKRpg1dWueOQ4SNsiu
R/zHltmCuqF3ub1aqRLVvcHinoEatzc7Gm6SrRwhM+KI0BMHQCEUmSCtD+bLlLS8
33VsFPSto2A2xM84hqq/JxPeajTKlfZ2fzoAKVrweZ3p/y/eamDL6dJM09nKXwc0
n7B2CDGPD7AY5uaomb2YF12As34xSfLboSZpkJZ53XcqOmxsyeJ5ibiDP9UA8f9+
m8ODreQn6VYEQWv/U/CDnfBnhfFWUvAbc68x4R3oxkW+5JSG2bRMe/BYRJp2iEP4
jxkPvY5TQY0WV0yTwGp+1lq5KXt7PWgHjJvSOC40WumUOj4uxuxszgybPmLQBCvn
U+K01g+CIr1YEz8jTj4XEBdq4U56lMmS8sP/u5+efs2xlMcCiZ2ReYC8+n+pC5Ea
w5e/pcRt5X/4cIYlB5QpLaWAYQsYbn7qrW15xUHmnd1eQBfXzExo1Qm4LYs83/JA
jB3ipFBcwlVCHQ2x0eilonoD6vvhe2xnsMFiXqcJSIQdJvKf3WPXqY0KnOeRSyrX
uZesvIBHH0STNKjPvOLciTF2j86PQgA4IR/9HwV2WsMU1Ze4/OttNONUPP5pdXES
uBjRX79NC8MqH5pjeHDa0rF5pcqZYYXZJcwKFW9aq+OWeaTNE8MVsTfnsiWWzYN1
e6rUf9n9QOW8gGiyI5AayytkB9bISKvGJKUnHsuSTvPyTGx4KjlJimudQBVl/4QI
1Adcetg80v5/f8uE3/JF5tu5eKsDnAcory/6ryVXgjOen4D5kGSbUK+p81tljupP
xzL4DKHf6iFlj8C0RvwjehtMxGsYPixizOy6NNUxkzHZYIPkdwes9LHmjeBlesxo
BU4GQ/vJNOK+XFXr8u0Iyo7QnXFR6+kRv8UQUEjjvEv0ZPpuYIqbljCpWL//zNUA
AQEbPs1PvXXZfmJ5BEMTNx6k5eY4S5AdlnjAtMsoff3npz+dheBR57IgbvfsMlMm
cGOJ3xR4nNQ9PzPo/b8UsfZHODocRx48Low/FKQdqfDnjKIY5myBoJaRau79jIk4
cTIk52ZA/SUFQoAQuTpgwGnE86+gwmPf1idA9EkEXP/9hGiOyxoZ608mr8hp/Tdu
9VOR+epoMfUgA13WU2D1sE1TdMeeQ77mNqxjkXPg6UNQx68rNt7Iifrea1jvgJPX
MkCeUqTdwS0rzrEf/tmlWWr7JzGcWvJxIDZ8e198rKHaVtx8ua6ko3E+eJmE6SN7
kRGauFvxR6l9UdcmiuPQKm8l8t0yWKZe+e6BvnD14j+0PO+vIGop/RqSW/TIa/JR
CBEn/omd4li7cMDwIL41XG8Fr4/268h25VeJui6qXu9AlpBbISonpBpa8litq/nJ
JDlDdhPftrpU5xz6jMJh4jQj35igVENRnODRVgbDHctGrajKz7rtI3e9aQqSOGy3
hywh+NmN9lgXinf5HqUNSt2dNe+b0PDOGtb7LyvpL69ZYKcUDR7SyPvSKCuS6Z68
zm09YEVb9NxCIuewWQPk0l019WWhYezIGfvEAJjC5ro0V/sn19pN3m45QX3cUNXQ
FQHBdDLBm097c8l541ZpFNs/CszzHIAo9W55afrOT60hkN8+i/ydiC8obSRQE696
szGairI6ErBfu2nd6vvUe68GJ3xi+BKub6a1S8dWNAqFo3bN9kunoq3mhaPO9ixj
DRf193Q31BtcPDKNEthxpkyrCQG83GWjT5OMHxnHxS4R3DENFuBWzxJ8UTWgJ6/L
8jI78fAgoNRF8DtyOci7p/SqZ7PqptCG5NcFvDWB9X/dCRQLqxP8z5W7V2Cv7+yE
jkf9YlgeZyi0zFq2uYzyJ4xdZ+8wNzIjylByxUl5BZpvjyuYk9x7w3rtkrFMXAQY
iaQ/LsMsEDo8fHdCecD2ETXW2nGhKC6bZvymQ4qiXX92NWHZ7N/mKAv8qhxgrShP
L4AHnT+cCrTSNjdoUig0fpCnDmh8V+GkkT0C2iNE2JAWEfYUeIPYU09G/+RTIppb
dOvotGtg0aJq+5fcNfI2NSWoX+4KRbUNKtX2ebKKIoVz+2iJg7yBz9uxe1XF7apF
vj0l6IaEfeqC7IS8YsPEFU9VnKiDKJs3kxEY6urlothh4tRVqLY/uq6jljfTboKt
+JL52ygDUioGWzJf6xSviZxf/yCF2nbpVkoUjuxxnozZaHjvItdiukBkmOjplVEx
FT71psptf6lOqBA7ekBSXg9Qif4WxRp/jOTEj6u9qnOiuQYbwj7tyDNDkllbE1Nz
WFA4LUAJWLKr2wXOCxRmLa3NsZ5XzJWSyF1LhdMyhxNp7uGVP3SRda9pjRTd8wZD
aIS8eSbsaAePukbhzubKREvm2wMqA1PU4aoLLVrWX+LjeEA8TKC2QsoN82aZ9AzR
hdKPXtNXLvS8+hByvh36wFqVoBr6daJR2jG8Z5GPzvVJAE4FPqWYmxqQQB8rOooS
v84LPvXYNlolN+WZoG4a//03XwRILizUPUz/QWhdJga9+1mjstBSo70uIuh3hZMb
cQSLZAaUXZQhA77s/gwIXBpScau2lU/JRdHxhWIKQKtly4KHUHs4SEoqJgtpzGrZ
5qqPdw5h4PXnWvj8Cj1vKdl6Du5mitCkGpW21WUZ318QN0a/W4Qp957hoeEQBmKv
6Ob8Ydt7L9HvAJ9sQpESTwBa/hvxKJgYad+MTf02C3KY5kCPw6K0m0uCN6ZGiU6d
1XFeUODJD3D7rtB0rNGvdGp1p3L5+Y3zips8da7iG9eKxbNobB3Vc1fhsXvMfWQq
OiPy+vSNzX1672DbZtIZuXPy+H44nGwC4Cj/8jq38cuy7gecIvxWDHcS8MSFVWrY
F3oPLIYdsN2WBtSeBVUWH4Rt93XTCEsGrMhJyxrvgBNknHmpK2E4KXLpAAQ2c5Xy
NMwALhi6dXQCcWX8HhykoT96iyF3ZmEEaKjBIM5IWgNR6a/YLhfZnckr0ZxX5GmP
2uDw9EOIaCkca5pp0Nu+hg/qoniQop0+9pU9yOpqDoNb45FYZeQAryXxp7BTYL1c
Z1b3Q/w/s9Mtt/d5MDmm7Qh7ZFPNFvdTFN11Dr5Hia+etD59+UQjOKuOSB/PbDvP
NJZr2jTQsVadMOGiYaN0GjmImrjXaQXJuewlpUR65leiQegzW8QU775uPx52nxLX
g9VaermCVYS1ujSn1WvI5HUe/zf/5l/JtCtRsC2nLuoX6zUSm2pEtpi7DT3RIAxQ
l8+o90jTtXX8d4ZOm7yOaECnXFi94gXQGoM3Rci03p9leA/tJKfIORmUdghoqGuI
o0vnFw8JKJaJk6wOrdthuHnRmZOngZHoJYRymd0RjRfYCbEaQazq8nlghlgxOvkx
OVnwj4Wmc0N3LDEqLcWhgHVyF5KY695NlKFKoa7BJ9fMBx8kvRepWtEWYKmlQkTh
qBEZtIzIhbfPpPPbmjqaRhKwgAr8nfgY5l0TPCGoM+AUA6ZWN/sQCRoVSWnn0n1Y
n2TW+0erugUMZLGtw6Is8Jngy5eIPuabigrl6+lYWN+tM8Y95ON9o8GCkYtqwrPU
izC5gNYqnmUlGyNZP5vhoSe4jYRay7OCSLTGpmpedst3XzQzrWxlBct+fsbWF6vD
o56MAn9Fc1lzcePmZnobTHMfIM91HiLTG6VZKIsn4izoVPAj30zMtFRto6x02Buo
PQXC73yW17gf3DihTMdFKFwEoD8zLgPif+mhBATGUbFaPTsQo33VoUQpwESln6ef
Z1t/HiIwcj5mTpjxYaLbrrX++u1qug8icDCetu3AflK70HfVBkeT1JEpGcA4H5rq
SEM7II3xgBSqwXpb/KJiU1euvQ3qkDp8JVZu2uHJDs8PE0ctrPS/VILdfwiWNywH
JIajIPba5/iyISNqcfa1dGLF0rjaJL3HPuh0QHonCbwTLZ5taCW6UHeWVnO+6Iqj
YDuvkY0gTOFCbJW86M8vtjkU78OvNTWH/NG0VboZRs23gRyCRr6EC/ikAViCZg/H
AmWtcXs9JyjgWQ819qc4DE8lCVgxhXhMN2Lup0y01EP+3RDuLu3YyhrmKu0/9GFe
h+nF+ed1wPPMve3aXyGRqY74HrjyNVQui7DkEulkBk74dpxaOkwlDDnJoZh+aDPv
zgOUrNDjDINJ08ks2JVEL2v7Wr6MBqiEc5P7nh102ORIsP4FUd5VJaYPSpz+vCwX
eehG9+pFRJcOPHdZrt/BdpUFgfL2VZWPL14osIZpDcGiLIBMUVUT0YAwZJT2elrC
1C8Xpcy6RVFR0V4Ok2sQe03QA7XuttEXWqqrGQLBgN2OqM3m5KTFPFKEastH1SWS
iykjGseguPs0XewWD3az8Y934nyReTklWG0XMEZRLrjSsJEdDDyx+KPI6+daaJ15
7Vbi/iI0QOsQQWh8uO2ChrmErpYG50UX8+aNMT9F0e1KLVm24OmcVB4psyp2UXRY
U2m3/eWgwQeufUKQ0w9kr+73pYW1O++eH0Hm4MIfy/88GbPiOiFw/o23ztfAbLEE
2KKgDMgUowcIcpJY9PeAxlFHZthdIsz8tzwlHVZAncYNIY2ppZE3aknZ7DKjKk7a
kAraDSnaSRsxbpl/hZCkZkK+XeUDrWsXGm/4vCVkTKsjuRPE3VhwinT/0iGVocVW
Fc0yNxNP6lcGgeK6uWiiWTuHE0kHcSBZ2+Tte2EiyJHTZY9tZgvYuwbRhrVef+nD
y0kSVMze4YKzC138AA0fuN1/W8ZbMcTqMmnd0XnFVyhfDhjVQ26dfEBE4X97HNYH
lwm4nX2l2u4o7dXhy+Y+HGdclRQNSiq77rl7JZa8jc/1MFC0ajFFXde5saSnsxVs
y8bSds80eNHz+V+bzDZeiG62ZYdp456pVgYkAmczDMKvMXXOqTIvRhdFciL54KDr
nbYiVhe5DvDNbAXWwJYp3bDIDyfniraQfX5/CrMnRM3P59bSnxPWycK1MDsZoH3o
6u4vLnhqOVUxwxW9szLQ0slDIBAQ0gtkpTB36xbjBBL3XCeUJwtPpvznfPdHzNn5
cnGT0ZG7Caa3PI+Qw+fxxIF8vSd+M1s2fkLRLFpHiyaVkIVODTOBGrdV4X1ZSf3E
GVDRknJ+4NwB8nBsg9sqGRdgAOx9DJfe8/Sb2YKBZPkMusK3ag1st8D+KQcb2z5Y
99r0dLaLTs6Vw11sd8BjNYh+6WOFk2Mn/0W+h3x4HOtkLWZGsFQbQ7XU7ULzpvO8
ToiY+2pn8TVFsRoPtlTO1cr4cSx7+VhjvIkQbKbkEBTKq4xB/5beGQDzDAVbXsHr
GkQLND8Q828dE7jqfkA+yldhO3y5nINjpVT1hAzXPFFR+i4i4NsDdkk+tbMH4o/6
jzAHInkzTy1zD2eHrNwrlnb2PgHEFoOwz1tAVRoSkvmxIfE2qQkv6zO6pyr3CF1Z
S8dU8Q/4AxkZXLbzx9Hu+JUVESwjjOy9YPxhoKmA0BwRvK4/6g79dODQElmv93jz
rpLUxivFAoarNtJ2j6KExxAWTJ0xp3Zl+ZrQ2a/D4cqGPlz5IBs4qZTPcRKPSqBY
vJXWRRZETahdfk7wxn56FNLRFGdDiVUEqkonC1/Kq75cNr+lCuilZ+OT+UIOA+an
5TcSV/sgqrgYqvsc99KmH9yVTocCPetg7OS5g3+PrEwm3QR9hp+np6YBAjJZf07S
CrFeZuRjr4SgonhUT6fpZBmmtLMPV2xwdeCnQQPMvQ+vkv65MdxOBsZ0lmpng2SO
DVZlj5C1AyPJItJR0PLTZvJ+LEXQXZimfbN9mVkFRNKShScElT+0dljEX2uYxpxq
xsCp2mHpfdsrNhQEY6dgmozJZbGblKi8lDGIe1Xi215ioYO3A4zaUmp7H5VVquzY
rue75pnizXiVYOvE3JiSh1qoJ+kUWicE6nJsMDrkMWxOGr/Bc7G7hdr0Ym9hNAD2
ZRmO2+UAMh5LaZrkIkVf4svEDtIiriUsSzEWBVZ5xn2iDBhVXLzCP6OqvivShIYD
77E29Ds/PddT0+qTLurRf4AOOrPdCpLo1YUe3l73MejMeuJaHZdNv53BsLC6zG6R
tIesIA7jGjMm43krcCuDsEVIeNTzhlfOGsV4SwqQjf3vFi6lVMVrDkHoPRi16CTg
Fo7hN7U0QLZjtSXi12y73rKdbb2a74wUcsDx9gSPYuhfl1X69o35FJv7Ry5kZV9O
F1Ktx5gi+1TFOJxDflv9jQzalXfAE44bf6XsVlftlnjtGSUFdQop5Mj6faHSZkp1
ciy5N7Y1NWfnJohrBSNy7aB11QpRIsQuwQPj1z2FOqKtlvuNL0kkCHiYSoYqYt2H
sytKaJ68zrzNSMpdEjosM3uDShNsdlOkypO+vqUXkN6IoOHIMgycmTBSMZ+1jONv
BpV/PCTmI77m7JXXrYbiFi2FtXoZf3nMH8/xPDVX4WFAgSvMPyHixFKd3f6A5+T2
IAYX6mHUCm/xGz5VCV/x0DbOv+44BysN/FgnOEAvMJF24+BdnQ6P/5m01WzhWKsz
EK7MZ2sJxecMlvOJC4JdoGxyxARkxffdFP1ylc+ujJWGHbeoPrwMTLEGAEkbc0z6
qy+L6srIhcV36q7I8Wt1L89UAtJh+1ZDQBm2CJrq3c7YmWKLHjteiasjbRM7m+4n
u5GOd8e52eI9Q0bfDD7ZXNrOls5hs1Y4D0rCmj+yg0g9lMEAuW4seTqZ1s5xCjRU
SZtN+Y0jEAtlnQ7Qz+8aOyqYs/nd8LRe1UMlz4pMuDZCUJTuKc89NwZb5hjLl7Pc
jtpabjLwRNAf22sbkjLIGUajsbaEuVYbl+4MEK4ycap0fb7mI+CaJ9pIfCa3+8z1
Ifo4C2y1aYranmWzpv9+mgAKNTyByJP3Qlk7wRZHXaAgLWl21WlmFWQkUbI3rMG1
+T+tc5r7JtL0Zv95VpH0B7XkHG/d416PhreMeoOlNLRD9SkWS8irlN/TQ1OlKha3
N7CmjtBEUwnppGGvtmqREOc3mFkpZmmNYCOVNe884pdhAktKX/p2AwMQLo30wgL5
I3Z6y1qmMkOM0sPya2yhjMuYSTRaHZ1m3ZdTSXqIW5e7P3hNEXX/nDkyTWXa9OXG
19hJLyOht6DzaTcC90sYPtdppP7YqGNCXj9GSL6EHm7yqtVByr+FtOg4VnIeORt1
Edtnz24wAdR+5vDg9wNcj6qX7rBAFCXb3WuchTVFSDBQD11gPhMvFBK9/Gzv+xFm
wbhheGwpTnKfm1d2DT5TaL4k9pYoZAOWOujhTLPSQWZeyJUu1uEan/sP5BJhBF9H
5vH3vQjRI8aidexmqYMCuPoX0OvLzlBa61//9Of9Kojt0hLJ13ZtXVFPeKzNtonu
Iidsj9FH1vkcuceh0ws/lpZXQo3Zhl5ofbEMBrQvrpg0J0o5Uh9ZaVoMQ6uLUu/7
4eEwaaOfdvdGkTi1hezzZ24kcUs5Gke0VfXg4YpxZBZR20saFl8f7UR8QrhCQ2Ds
Xk7e2hW+N9r+6MtCHtlVJvhwaC27Cbpf1sQ3NCmhl6CVZlGkPzfXMHE487MC3s7s
gEN4cJtu7khmQGvkae5+vcn50a9jNpXBpYS95lyDJYMHSs5PwdZUfEHgTBDEOARk
podqa4Cc50ZqrlyLUlRIkBSGc2uFXV3Ko9SK439iqL8FIi1btRUJx5p+rE8YMQXk
mnNYO7LHiqMBfSfDf0WOu2JCAHtyN3bie8Ie0yuaK7TH8Gkot7SmT5cCb7hOiP/c
olUgvlKqTM+RSrSmcvUBde9Y7Z2RnTgJCDaReEOjCjkjrH7TVRW23PmWpyYuSKxR
6ogJ2oaSZOg+qI91O6/IGKFfV3xA7EYPySpfcDd3brMaoK+SAUrphWKJpjf2JrQP
S1edMqrx4npO0+0G7KkauNVSvxCOAUKmz36lsTbd8cJLAemOtoQguyEUtVuqhY1p
gVl0wuTlCUWK1S9/eAyzGZQ2AzMCov9s/7X6Ql9amsNBpeRQjgdgtc6P5+NXuNw8
HI4USQ/eThjmx9zCXGaKjwt8fg+1fjDazoCcUB8JZHDoTV5z7hkMMePk6EdjT+OC
1dZBjl/P6xk5qLBF4i5ZVe25a+et1Ul0lYgMR3waK/L9vzdPu08twloYsbMYL0LE
/ESTE0zqmnu9qHyJLQ8/w2xvgtadcJjpgs9CSxDqQ2k2/47aFAv/wZh+TFJjCDZ3
q1jWC1G4kUezGlnZqjV1tXy1jE6gxKeKHeftoPQtqtvXJERdmkuK5G4L9PA8TvqL
9Pjv2NkY9gc+cU3XJOeYKCe1ijpt91I6wF2WoCNee9RNoyLFoHbM/99bffCAAZ86
DEWslACWZYKJxUucuI9EAN/atPjHXKuySRIt7phCOn9OTDl80nnWb2gqfI92F0MI
3JJydAHiJQutE6Crgibyz3sIgS3BR4WSu1lDaEWWffIUh/9Nw5FKAsfmnMhBF7FY
AzmZPxaUuIJwP3btUhDZFNdr3ESrKJNcb/WJT9W11DqJrtQcqV5gnO+eaFglBNWi
SsKtOmE4bPc6F2v0SVtPKsR7ZaU2xzNzCO4tXk/l912WENlwBi/qS1N4p7kPyAii
gMW/ILAjN87IMNRzEiVaSdm0e21IjJoYogZcCn2NmqpBU7/FHlGL2uMNwTem40lk
JccZYLSbVbiIQDF0/qFHBLomh8cO8RTldSLMu4Mrqiw6s06TuSvds24kWg1T4v4y
X7bWUmDiRbm5zOA8uQlcuh+W6F/p5/g0mNqnZO7T7DZ4YgNXeikSQylNajK7wAaT
40ulEK15Vtt6od8D7XCuKRcrVe6jBb4Ub0FZowWrJHuoPaXHkFd+DqwSZDnC7ea4
YYeYIudG0KbH3MwFA/hjJHNW2MmbAKB9t1iD8KAZi4ZbbcfFd2SycEOv3ePeMgOt
nDMVoXNtiVojtCdZi9lekzHIJOie9lxwsbmFRqWD+igPtyWPOaVtpIB3El0TRZpR
LDOsSa71Yxx5SXBzibY3eIhCcED+q+nN0SkzhJjWYvRGSjlxaUfVpvLcSl+W7jmU
AERtWyH7sc5uAqhNO3eWO6Sh1RzxtrZn/TbHzF4Lu/qYkuzpjEZ/q5qen2fgxDXo
7lO3M1T2p9gdzSz9SCxWnXlhHthUead6pHxxUbOaRmgiONS3h8kxQR+kzf5Q8eNO
VQ12ICccmholXs3x2N+RERDDRcNxu5YfgndON01O4MDUjyLTXyIccb6twBSDBkaT
1t+EhD5YHVtGMoHeBwogyMf43mNOkiJVZcSdNCbCEUugeyO/LKYhnjskfyIO1q/J
GCiq1a7bTkSGUkCdINcG7LurKViAw7N7+ueVQyxOkXqZnUN6hqgL7ErilFUvPuEP
ueY+njTz7A1hdpVbinBQtJ7gVzyt2Y0sH2Z8AqLSZkdCLXS/nNZ8m5JQ9o2hW7NN
p0Pu8dhXNW9bshsLGE+cxAwxjrjuTI3b3zctSbzMiv0ZNzSH6KGam2U8M+c2FhEn
c6pmbkmVxYLOkXKza3cFqe+lIRZcc+SuqRkfIZ8JHTwT4vIbVr/pMoOP9CKdfBeu
j8POVXp4yGLPt1Vp78jnB1+F5zZOqLs5CIRZECoIaCHZufLoLnz4P/kWihQBz588
3YdYMCALnCY2GuVZXgI+B0bheEZv0kXemydGbe7yeyavvnZ+sOEfUgejq498ss43
8QNeYerERi2PePNgVQbOGh1InK70inzEAFHFy5vkSKkOHYBBkE2OuTkecksMP8nG
UQmDhbQXbpk3YH1CyY39rXoGNm3x3dljQteDfSL3jnBY98GRKnJIH+/JMF0lLhIb
ab8HX0gPpXjcvt6P74DuEpLH4LXsc1J6oYNNn7IY2Mozuf0UHkcOCfzcODaqUpG3
WaYX5HpkVNoQcGZuCZVfj2K391O7OHj4n76fjMHxQ4eyYsHdz6qkVW7LMzhBY0T8
Q2DTnZGLERWWIAHmfMmUQs9oNLzae0SKKM4qNMkU3gdGF7BA3bKS7ABFXaUdcfEt
wCmyYS7fHHkVFbOysP7CXP8fXQtR+kgGgkGFAom4g4gzUhFa6i8hpUjzU9qECZVo
nf0F4yabMK/GPme9M6ryZQ7A2Un6jcBoqihVyjg9zpC2ceOZqLSZtkKKoXoadvsg
mUug7YDTOAg8NomwaXtzM2GSRyLzaHanM2Bg2R0Xe6BY/yKOa65CEB0nKSomOrbK
inhVnE4Rb3viZWfA+eWoFIv4wSMgY8YCYLYpPS29cUhBGxJiK3hgl8INub7k6yUH
9IiXN4k1134mdqP+mvDGEqaL8PiGdpIJhfrEoMvXOn5Z/SyOfftaGrSVtZ8ddUPP
+SiEf4ltbsZb+NeZMr5EiC/LaN06vXprymQ4x+7wUkbgBdbbJ2euQYhbqu7kw6ML
DiJtBTH03euMNekYVNw2cL2N0qt3Koeztra2EvXN62dmK/pNcl6Wfu17M/h+CJEO
vqVKfDkVAgLvUFWi3ZcX1zLrucnRY3nQbkfJYaQ9VFEsEtBIckfHd4RtY+qn6A0o
dQYlPOH65AZjqt7lRdl5kTwymU76/4UTfWhkAxfUUWrzkOTsqSHeKC5uJ4SQP10P
HzqfwtAM3Jxcfc0GD0B8agx21mkY/Khg6Dz0+w9+EVPxQpyaIHWJwcTS1/om0/tr
AXw8xxCfwETWVIdJJCkyZX0GLYCT6Yeug4rxUYJOGfKZFau9elbnaIFUPv5GpaNd
+W/HjVVBGfhLZfysUYkDPLO46DrLPHPP2HCds6nN+KCyMabzQDsGuJlTaG/3EjW3
2j1ZGzVL8uevtceXQaY9KBXIlVnC3g1dL9eYV+UMuKianNt/64zNiN0v7tp5UpIq
wD+kTasXTVk0dih6nc79HQS/OdkLwhCaDKlfWvAdjK5aUSyMuxVloywdlu9Df006
Jd8qbf3GVZBUIHM+lKGaaPW3TbcMoTWi1NWXIAe7scWtFPyfgxRJ41Rir+Xx5ynK
eMqvEuNjlXyP+a6XYrRZ+lNKanu0W6nRc1wXMGde3rcA8BN36Gaj9YlJhZ9/V/a6
kFS1Bv+Bwf5nArF+s4T325QYYuGAverwLqFcW+Woxb+3lrSrSplkQ3nqzpZL7Y0a
JUGn+AntCDlA+X63bsVEyq6dfBhaejS3/UN8MaBKBPOtQ4N+M0ycDm3gf8INWL48
0ZFmSaP180XlXarOQpEfFwAEIqzonQhinxyPnXa2l0te6VZJ4jcHfS5n60AkPyBt
vTLjc/5pvIULFGqTq8uyMlS8DM4QvTvNK3bkxIz99/F0ydcaHEaZ6JYo9ZS1HT4l
23G1sAwzAfx8Vz7+eamfJ3wfC6UsVAGA8Xv04Tapn2IKI1w4ZliHGGv3m4BKNScA
qzcz3XyQJa4jOyU0VFUKSvbh0Hf/1la/48HjFaf3WviKBvwJPJQSzxklDeErDTvG
acSqzIqtXXjwFSZHYMAJe8zmgrDhTfiv52hQXis+49D9jGaFl1CSKGYZmlkt1fTQ
T4UPFYQBMfG8lZHrnscdhFqY9L/GaGRy2FSz0bMWEQlKeQtvnAkaX6khvfoy4UA2
IM/kvWsfYA6LTg8NwqwenJhYXaBD4oX7cQy6RWCLFs9Ftv+RYceYZdAfKUhlpSFb
xz3MzAxQx9aGfq0y9NE0SHBWj6tbbU3oTxYcLFsxrsODcB0o9KxemhgJtuJ+mOzY
AJhSOgkQKHVETkHk2l0x9/yY5yLMsc1LGhf/e7j9VPY5iq/r2NjBR5YW45Fv7Kem
TiYHFggcpYaFjb5RMJI7D/zZXadz41rdaf4ssIzRyTnDhaQa2Xam0Ozn9YV+QWeA
85GUXH7wWnX6v8h7yqJfYePLjlFxe9fnOXJeado1IpbZe5HBN+xKEkimGfx4FX3j
Uv6Glhxz1MhjCnuE9RvlzwGU1prn0uDQKtcU36UUq/wKmcNegXdBLmNebcttXiUL
TbVOF6Br6dkCM8Btc6mYxybDj2GJN6uim51oVz0cz3QUtLS7ADyzApYyVBaScOmV
tmrTkAjdEhYTxYt4NmrlRxn18och5dL5DmkSQAPW6jN4hn+lvWiQYXwgGJMYFAQs
LUE0P3r6jsPSmZdJn0e9HLxT2oAQDF/UEQ8nqYuUc/PmFEOeoiL64RukZtOkjGsM
sEqMLOs/wHAQxm+rpHEoUnn2pLwKk0jYm8YDSqXJYjMPK1D3qcj7LRZHUxfBs0wW
ATUTbtuHaWRuwVcrRL1qo+jVBR1lhBTcO4WAxAw1NnCz9YrBDXfKF8Q3lHfo+Zoc
ygFFKJtpteU/bPmAcOUg6eiCE7fu4IzJySI8aCYq4wZ6vjVapqZWUhnHULryKELt
s3xqdV+vZg6OC7hrHpdsS7j8Jn6QixougOYeOuRvUqWczIpH5V9S4JWO6TQzBam3
LjztxkcOgerOp3l7NDjWcb+WjYkbX1dHfU201lNxphq2QPbt/7yOJGAMrKoOjzEv
V+8MhBM34+Bb2U1zGRO3RQrkr36NcGYMiVtYaFSg52Pn0uSfRnwn45QnbBf5iFcp
tdpTvIkvSCfQ6MG22FF+2AC5xm2Phj3QGHvCHiUEk4e/o0IsDCM45uFET8WgQVsk
ERT3rcpMSi0ZrOYetkwVuZA5X46bMcDHxwb9MB6yz3m1138monB9ec22QMjwgTku
8UlWvRddCMAEi39m9+lktAkidQb/CGdYIYq7mXurPDz1vZGNN9rJJAy3LTh/4ZXK
7QOfVMzv25Ob/Xkefy/7i9gzUtLc9I3xYpkORbiUWEYCe8yg6oXz5/dF0YxBS5Jj
0+awRF+TUXz0drmMpYDIR34SekaqZiZnvFX5Fi/clHqXbj0WLcz2BJSMjtlWKCxh
cM3PTegBer51gR7nEgJdfsmoZSmU6IGy+ARTMkFR6RDy1Dh3ef5Az8FlX+6gcpiV
CGXho7n81ftwJyl58QQeHRTxaEgSgmoZW3llgWvoA4p5HfLmd9UKxFLfN2Izo6Wc
uVKtpheom6Ua1obXFd9vA3BTQyJByJCubdQiOLqRvqcSzjUx/oFFZwdaPfmhkurp
ZFowYqlEbLYrBW1nk/aDPc/eGe9fu5fnXy037Zyaab2GBigr9sHy+VVR3WaliN2E
4JCDhenRXDzPWGq3sVF/wkjKqj0x++g+qR2Lu30ULLpwilMgpnwW9FXVpY/kszts
yjso2usRsr/8RAS3H2X8i4ogIBiZ81PCFA4art2IsAU1ONJU2siqvkXJ/qC1JgEV
Wq6FrP7p2dUCUFTi64uFPrzjI91ya8NaBH4qqV6fquKZM+czPjSe4sHPBoeEkOgm
9zw7jU6gm0OOSZjWR4bgJpkm5vqVtz85LMjWRmINHhBtVMn04GWLzpK2Onhn5a4J
bySTNQHFDpjX4HBH0k2n3r34f0KA4vxSinK+wd9x8mmdABdSby3feyxM70gz8k4Q
bHsdk2XpcU+RVxuaGnp+HhjJOrFVVspeYqWvlDAHoMmsqJNdB5m7ShQynK/e1e11
mLQhrIlmX4V95oCiyUhQFvY6HeDkLchx6ag3Ri5gtzFaX40s3Zq+joi93DWVB4sN
2TThr85fGRBq85RMQ0Shz0yygGV4nCFO4c9OwszRgEHOBZZYjtJ6vxPPRCvvTfAf
RvGZ+NSiwBwMdzEIj1/fu1ToTbuVj1dUPCVuSXbak6SWV3XPvXIQ3rrk463GRE9A
m0zlpfSuZJm4Gop6zEeppWbY3ENRtpG7QRWi60ktASDzgwXNlSpmIctkRfMlFr9i
RwZ7CF+DoZpIO3Rly7tSuOE5AOWsOUecUbudOGGe8rxxvOzA1b6ugCNzutBXCPuk
WD93WmII2EoW3hMicmPt9E6mifMdONNz1YIGpQZI6LX5kGpXGVDeeYHytt0M3f9a
mFAtpCYaNoDI9H66VhUaaNqX6PayNF3nHHxO1+r+jYVq5gMifzkfb2UwMKkjFCSa
g1o+P5fa4oQvkBPzzNnZe8vz/zLJ240n1XcVTdyon25YHZYJvs/AecRxPBLWNUOK
WHrdNltVyPwHRfivQK36agFOGfRArYXc90cPNpFpE5ic/yzeC1Uixtso2N2ikxxq
IapPgKcH8sah2q/BUBTe30zPOF7kATDF4zTg8gE+4BhC9yx/AqOsaTs1a2vDybR1
jV9Tl66g0BQd13g8oPbUKvjKtjcg+uZXH6378xVlhtuCrFcubraEQc0NwoneXcae
l2ZEWUcXw/syx7ZqVjZQ9kVi95OHowoAxzZG0lH8oX37Rg008xT5KOar5rqdTQU4
IMuHyinejeovrH8qzoweQeOMbI4zGOt78bO/lfWw51n+841TPdAdeASu5Uu/jRuW
HcK3ICFi3kvTuiQnXg5luQKLLSQdxIKuSRJHBcE7noKJzlMhOFMPkO+PTUPcg/l0
PNSV9ZXLBe6HFBRoY0fSPmpZVeMPtShtuni/CauzqfZ21SB6uQA5Ue62XTWfXwmu
WtEVX573QUrJtFuY2XCoj1U/QBB2NdrBcsX5v6D8hRvGVPHI01EDJKkzz1vKwDTC
7uvvigmIuNQhLKFtvzjlU0GzZBG88vFqmSl2zwiPmqy4yScuL5GnFfBPckffYW0z
4crDHpaamFlBzEPBJn01LhVlHY0QJaxo1Ztdpj2y6F5mmAzw3E7CM9GQnPFbL3AS
IZsIUOCJN3T0eAIQ/+vFrhU2sitzC5voeqS6Msi3Z+HCm7A04QhpUXJz5nHL8Qd8
O7dtj9BNRcYp5oSDBiaIo4bkfc7WxTuwYOjaeIVNsAmVVHeSxQLS8/iNrZhfANuF
4LaUDElas0plcAKKpMgKgauJOexBfvYGMlM+SzrGV4hfa4EQhqbu+63uelg0TVBJ
vf/BvKLME9lW8na2TkBY+u6W5TOVW6enqzv2hA7xKG/vLxWGc5dTh8W+XqTdiW1m
pn5ZMLOg/mTwLVUZT8D9ye002ClY6wc45UgNfK42/UbhR91SJVknySCxgLWxCALF
FA62k4dALWR8AopywSqo7nrJiOj/9tF8H8qVEOIPT1bIdQzOdEbqlcJeLXC3RHsL
laOR2Px0zZGaW29r+CsoASnOrxGsJ1pS/6QtX/m00fG2bFE68OSM55q9d/K+LoJq
GsJax19AAt1n2wh+0cqW5MSY6bjZfjUrjhDydVzden81XVkJp4CkuwoozTJVu8Ms
sm0cfQWiSPglG+DqeUJ6NQh8idA+qqaC1HhQXLPN5H/Hupe75OmqFO36wdqlE9F1
lHgIVVS/TUdoYYHr4MkaFLE4ZYUS56u3Fu6rfoDYZ2V3C63okOmHsiOnCfJjcaM0
4rreolJZGooaIh7jXRpjUKDkpLLxlWHjbz+Bgqf/krUhpWA98I3A0f0J2XShtfER
FhFFLzXkRghzz183n274TrjR0j4AqLEPgi6NTEcCy0mogAKiiE6RzCFG7ZU6kINl
1cKG6kVMXvckQAaAqocmbFwozuuVqFYL7axnWC5w1GqtFHTZvIknR8qg49a4MyAL
gPXDeW9BeSRoQKWqWITvIlWfDfcX4Q5SDckMId5ntguhompyjpeuS0nLuMm9dmeL
GNmtseHv4hMvGxhujwmyMHyQleKfZHKAeRrvi1aPKenoAC09zPkjddahnA/aQWBy
8RXoHm/o7f6BlKfzQj4QI2tMXxoZUrZnJPZeQs9hmfvipFp/JUrASgMWlUYeK+IW
pddV2fQNF2xAHTAsDixH/0Us+OO2g6gNXfAK2uG1nwp9nvNoItFyTLJg7uhQPBlt
dYLk/H5FXuGb8YtR69IoFBDgcrYi6tY0bM8W+1aqr9NOh+2oah+PkdbtxnavFiWJ
4Zz0e3lZjcGufDISdO4C4Cij7yozFOb/RDHkuO5aToQXDKDJxApmacdQMM6MKYLQ
w6zgyCOZ9aRgV7WC+ch3WBCAeliMRgL09zCLNaZmDsYwq0bJBiVqQRPh0pfSYBmW
Q2KjQ2+HT3RQfM5hORJ13ST0/grKgT08qzA/Dv3ilGCGn8hw81W0QE85ZJzn8DVd
UpuscKGNg5NSHcahWLz3X8cq/lKnrQB/Hwb0+Yea7lkwf3UqKkmGisK81ziD4dPN
DcaKMJRsZk6/8S+TUFhCmCG5+Ieq3R4fXeWgMsy+EIZUxwT3Vw8KnaFMm2t4OS/A
tnL42O+JFlQ/UHF/dOnpx2mnWagG5NcEiQuQWn8VRXMG1YfF/jq3KUhubMkW82t8
gjev7I6TRttXFSmqit3Wh3IZHAvg7i5M2NtyJbS6k4s8y9tgtxRO4ozAEKqNGEDz
ZJb/kVoSntxk43B9esHaTHff5OavjulBS+RX6cKvdvNTe4CjZsU/9A4hVSk/fysN
pcno2nBY+nIIHTyW20ptnDg9xH/pLyTRx4stYmUxPEE2lLdPhclg09PM+K8CiYD2
1nct94l0X5FhAF6r5S9Uc3+CJAf5lfwQ9tto2bEI/yKvgabU6KUWLppjKdN//AhX
2KEOprkX4ufGm2fIZz8qCxULr31bg7PgwCat7+zfGS01h7zPOES8TiVKGLpd8Fa7
6sajbPX0B8LB2U5WhH72HlsOmqxb2ulnsrn2hA6phMPLwgcIO6ThqlTfdcuhl/h8
vBfn13VXQZehAm3fC7cybRdJVfKnNXvzsfTF46Gkk0v79L+DJij/qm+ns8ZngNGB
j958ExW9r7EX+d6pP7NtAISNrPlpNog+d1RxVYkYhEwP25VqgLC/EM9gHeNfJ62W
9UIa5xNw5MVPC+U1WtlJ2fo5El5VRcYsNejCsPNaW4qIOKh9lGuiktq66w/ISbSZ
DX17h0Qv7TsDTcfnCQ0TBsQNEJ8sLCGxO7m03LOP7NegmX1xBeWCdbyROZYSh+rp
cXjwbBpldYkGOPOhY25UPo9k7W9XbHwb2iqb29tj28QTyUaddq1w95y4eR+5oEcM
o9NKJaQaAhHF4/BL1FkMJj6bDEQow4IrRtQA5ggpZFL5xUPG3KRK9mw+t8lhmj1r
KP+M/V34mPJgaXNdsik9hfjFw2WoA7sPnhSGbMnTIHO54eJ5l/OMXEJAraaeyomH
078Eo9iQiSTndvMh7/1Hg0MqX6qfKNqjIZbAy8RSZLLH3JsuSobcnvri3RFTYJHA
KqRe69OLKaOlfAJWhosbKH0rFGnzy4nVYYr91ShsFFp2yAhUNi3iUp3o9PLgzW67
ODeHgattJxy7Uqe9f900zYRoZymgNoXweS5+enO8I3IeVj5KlcOvJuSJ1bOOZbmE
jDWU39wLxPDiMDHNjnn9dBYSr+qwePJEEfaoCUZ20uQ3YY1t1l1e/8zAbDYQIQPk
+vadpRIzY8IvIfUoiDRKY6JuTZdhGHz7JGIb2wEfzeQwryxBCXP5/3iYA+rdPBy6
XoSdVdd60/P40w3f2hjuJ3gH06vR9Pzv4oMZRRNo24E83wagra+G8Ggv/oWac16/
cDUnCQ2XaqmfYAcFZ3iVqIYWG56kGUVLWy5XPRwgazceZrgdSyoHEqo+horQv4Oj
nAlWIHjbxc66jHN4SLoEDC81SA672B4HpR4zpEAAmhvCjpigrAa1HmdMuW9C8R6z
+2zYqVRNWpZhIH4rjimRDTGR/PWGAVatUncGNPbpLx7uRdSFJeYb6jbTOxo+bGEI
pTPLmnnbLt6rTcYtoBralcfhL2w3bjYv7o69ld8jH5bqGD1NkCTDClcAUa/Loc0Q
3dZKRHTCagE7jo+zMrijjwVsy7FSvxJ7bMu6jLrRL7cITHSZVJhXXUeW1x0V83q7
jroxnG72vM5k9/yVEVVmwdlQ1+e/+eX9tbnq0o7Kjb1O/8hfBggISCYtllPVUhfl
A92eC1Y/oFxSdlSScNmq4ehxy80jmadwofzS7dLyiwOr7iTcbVU/EIj0FGpBULYb
D14fSbVEAg4HXUwqyWiCrDHovMKiVoFIfBd3SowVH616yrw3kZ1oFF7Q/qyOJADw
6VsDTodWnmiWNm6kYcaAZDsYSueSNMKdF1iW2+TkqBrmsW/3xIZSK2nie5avumPv
7AuFRZz7SDTa2Ez20rewD9vhTcB6hmkoC7uce87ScAltpuXCqosQJzt8LMB5rXfq
VJVWIBJOjX8hqtBFKqP3XkQJoWXAc2fyOF5SPOdHjMnDMomifKZiLyZ/QJ2iua3A
urARoEoQXAeqKnRBOEDEKpbwmkbyJ7jaS6844fNZsPn8DWPKTwWNTeIup2WgoENv
W+NnL4rYp/hoIy6aCBoN9WcLE2jVcB+wrc6nPQrbrrOpnkm/JMvE0qWJ5Rx3E/uL
eD/Ybrb+h4EvWpQIdEiR3U5r3FUAM+ggU0lNo+QsNwaFGsFFJsrdczkpCKMGRmiC
RHOq6xK1GznD5F32f2ErE/kEv4OmV0Smsjq4Nr7krAiOKiSIfpySnV9mPL0ksEYc
rj68Y0jIkW/jj+SRp0XhKpKraYhu0w5a6ASSZWYZ4WEjev90UsHW7itBg8Jc+ok8
A6/y7zEqO+aZ1FsSlIGIOCMvtxb+2605H6boENTCKmJiJkQNEldNUNx2mLjeh57p
Y2OU6PkbxKpiZY8CktPJeEyJXklpnXgW+uBtrRgagb6NILeiNT753z48hMcZ7ju7
NGYOfwDFsTiBmBnAm89GbpzppT4WhL/jsCR9h0pudWI8GMQQd2LB+KewwiIssB5O
8b41KrOSF8B2zGdgbQr/XuhmlDA9jrTa3EBCuMIPB3k6yVr1caZoJ+4PbvttJ1EG
rM6d74or8Fh2TmNFgrhQ+VsxSbeKLIGHYWPmFXK5Kz0MN45eBEsPE2QiB4Z3B/YK
3Je5IyRqXAKyntcEXkEMSXo/f3ZujXj0fepeLwihPGVblaY8ZuyyG7RoOboBCeCE
KTTFVs/ugaA89T1EBKfnVkf2RZZKHHe1Y3ctoZLdLt8WI128/Q8vUcwHIDJVnx4x
ppsmTZm1Cnl4XbDnWYOHMYkyqEZIC/Ux6UAMTfHBXSnZ1QjacSxdAYh4LWTkCXg/
b1a1G2S6r08PE639fznl3PzQQn/mZuPgcy954nfLAP1IKOuWMcdp9U2uAv0GJe/5
GuKshqmIdezGo7ItZ03GUZ9hc+x3u7GMyYPGJUkq6SzBpbaTbAa8r4P+Yv6eG0GZ
5w1njgNnXXojoN8L3M+4+6L62ESlMMJTe8NlrhkB9Gzca10k7po5dPyT8yG8geww
Hi92vPVfqM3SIrcFWxVq+mkBsfeFMVs1ZGzia/wpVivELdn3ZX9wGyP+J0iuq+Xk
/dqC1vNUvG2ok9axPTax8n1c+HvVkVaGpT8oLhnHFd92e7YH1z+T0zgcSwFvHS7I
3cUl8PtYFNA98vM6+m3cIQWRWoQq6XauqrKxYkezC80zAxPHkFF+4s+zbdDCGCNu
dvX4pqsNqg7STTpOY6xWZEbH55JPNpojRYg2tKzQUpvIianz7xVkk+pV6NBWtrHr
TLcaNUPb7+5akf9d3OIqhjJvpuLbtdFXXgMZ3ma4qGzlYZ1c6cPWfS1XvuMSUml3
ixHpyiq/EZFDKt3irXBRiDborLcOLCXZY3bWHn/+UVi0ndlt3l/yeTGyM8RlW/yu
qVHsTDl44DoHDFTNrDKByQddQfvVCwasYRy+A0wei4+UjSoyiwN49NKQRhmBZlT8
IgoHaYto1SL5gDF5JdyTNQYLGWcffzI/zy95d7+4p4pjjJtWLpySa7/WXVxg9BqR
nniBOmjnCTNOUHvGWKwtJwAjdZ420WsJ4QpQ1pVl9wxBEfFIjW7beM4OB2yvpcvq
AkhCz7khgRWyAGX02vkcR8hHeqir4+bqYesw4sz29fAS6Pmw3jnjA0c3iqIVjp0i
z3kIPOXWKoif6V+IrY46FliF36bzClSMXd85EMhn37XtFt6AEb3knyhhqpS6SvTs
h17o/Jgd1zHizcZqsUcXMGhZo5U3CV2tZsMgTCINC0jQmiLTNJ9DKvr69HKydPkZ
ByETdObEXlTMxfSdolQKd9H8rhYC2wxENpyNogCoeg7RCKXAY7WILQCskf+1LuNU
bxW8nTA1fxd99kiaYks5C06ISStXgz4dQXuOP3V+myK6JzJDsnDK/7RPn6DMuPxZ
YWAv38l2OaWGoB0zl9dE2qAg9iHpv4OYPFSGL0F45I7KpS83V6i0IXm08syOHLr/
W4MnZnUvTw8rYxWxvn0kAzfG2NsNJ3J05DPf80cv1XrG8auz4A+J6aLLbvUvzUOO
90Gi7yZ0squ4twvEZvexT1nbC8/lDH4u6Qnu7Ad/c91CN4BSDF9QxQBZ3tVigZyv
tev+DJMDl06kJvpZierM2VoxcHmg5H7xax1Bo2RXUqTpxLMn0GFerbBAyseb3LCg
BaYhc+SsN1fgNKVUwkjNw7kM32+u7JozVp7FyjroJkiBHJtEQEsdw+lfH4d9HRd7
xo2ytq28INYSNuYQwlgPCCP3dryt2zDqprpW2gEhjefGeIkKQFkqo09cdwRAbUew
TH3dtYZJYly3WugLHVRMWa3aJZY93h2g6WiB+bRxIURiMy5aKd8pW2OEL0/CsB/7
b1WE9QS5Egz6I3mLaOVBV4QZDopi82uAeO0JcWHagPv1RrGqR8H/paXKFsd0ZHqq
URbdRODZLd7IDQYxTpXZNWvFQ0g0nyfaPdp2fzc9mbbXP4A31wWbsWoP19N2obYV
fyh4s401U6HN0ElJUvePUEQt+qNcY0mIyNO9B7PEw41ahI3paapumjUlfpZrgdEP
A4Njc0FXRB+SfW9Ghwp2w44zialoYQUJoaRBaOguGUNQDuK5Jc6Vm1wCxCc78uHc
b/G0nI26VGbSEzd+Diavw5Ms2/WJx3kpsz1SEFFQyYTJ96fZFw0KqH7L9dc3HkDP
GUHr2B7iqUisFkvph8svN+2mv1sf9oygZ1EePJ7F2YssHnGMxGpCeGbIt66HIaSP
zgJ6+X5gL2OvXbKz/OE/0OgYsRLaBkZXt2fmOQnJgN50PoOFaU9hhHBv7c/cZbMX
OM2KrjtrWqK4cZzGIIcCMdiZS8NtE6qSMl/J7WWmw+6PiXwLqzP+TmxHz6qEo1kU
v1+p2ZWbNFl5pHBhZjb81jfZjcDpmlyHkznPXD/DGF858k805gwD5dsq8z44Ye/i
uBEY1NH7alU4DcjIK1YOGaO/ZMk87PDPGd8NXaRaro+1JfjgtIJD4RgisxWZ/SI4
nps44tktDrYZt52+LavZe+7e7+A8WaEt4h0u3CS+BsquRMyZwxijWk/SrZVCqmSb
LwA8WLXnlLE2FGLQTHOhAwrlPAZDPEV0WSm/X6R9TCc43V/VQUC5qCVPiaHioaL4
4k17B9l64P4aFdGLbLyW2/ec/5e/TyX8ClwWJVu1a51YoYT4GloDmt0Z+JZcmf+x
wWK4EfAvQheONgKlnEHGxZkQpn53f4ZbOAynDXJFzaLJE9kmDgJviPDR3huMziLz
qosf0czPNgZ4sKLgY9gluJahkccEI5pyHq3SPWsvMgzym/NHNi1s9R0FZ5F3WaQP
uxCpN9wEr6jHnWE7+uWOpRcCH1dP+DuVxgZDoj11tJEScQLmnWWp+JFDbM+6jm5m
ZWTXu60fSBoWcscnO26VtLKuDSyOORLbkmT1Y+pNKNOhTVhtEarTUYaeA6jSJbCF
o6jxVH5Kp/+pm+9r11KK+Qmj+Di/5V3w4snnzYH+BZQ/hyvi8WWfJ9Wk5ccT+WA7
0zX9wOqxIEJ7wi4+ZlyJHwZV7deaAAKdss2MCzq8jWT52f7UJw0MrIEzcSGQgjyk
K81VNRrDZJVNrjkYE/xw6iIRMGe1SsS3BCeeE47XLG7+Ckek9/FQew65weuQ7MZ4
B8Ww9iDTvc5qKWbQWIsPmeMgrnvTCuz/yjquYW/pTkm+gcoc+q6Ds30nhSNU3aQN
Ir0yxRvkEE0n1zR2tAVEspdIq+wiYA6gQKt1emsenCrWpuV54mYRnkCuDHW9KHiq
JOyQjAcWC7tbLqOOKAFSDtpWUPeZ+rCnqyPWucLf1d2NJVW6HgZ/EC0wFsJqShpf
8ZNYKi7rBWbsP5a1tKxQlkHTEbxYyHIwO9f8SLFENmaPsjLpHuqBoq/4kweknA8C
1ZA8U4qEvlIw76s6D3ksXECk+egVp82Et5jq9HN9v9j2OGU/tr5ZJF4kTH7ci2nq
gPPz1JyE3EPIdv78YgJKTjn5criM7kMWxfp66nGwTq5IuhbP2UWb4iJLr4RF6i6K
CF6wUbNC9A9cl0vy2FpHkwqVWnkMZywaU4KgwYR4lgx3DzVVk/L7Tbgrm3rsWRCs
cJB4ZcyT8p/uaoj3WSnIO0DdiqjFEeixNJHcOV2onicqygi5GDtidPBpLjPD685l
15+brenUjc8yFk9csSbCu3sJnDKU99Xve/MPVQ7seJw2kmutlp0Y9CPMUYt+X4bM
g+Zo+W13sgxuE/JmwCSkEfxAWOuaMj5j3SVpxgbfFZXjucWu3MsipmrBhKFmbG09
AelzY3nfIG63CATRAET3h5jskkZcSn2DiTUPYPDr4agxq3bEQC2rp6LIuUhpplnl
1dlWvl8k4OWdurCp1RwcDcnIs9W3NNDrm46Dkldz+BtUsewHgiYimbYWdGUh9Mmb
diuUiwCRbUIV+JcsQMVbg2+YuMAoOnthqMDgvmYyHdAo/MYcT5A8NpqjY0zSQLle
EvVPwodza03jwAJcLeBMS+GEstvtIgexxbQIXbFFnqbozYlGzS1wQ8qcoavwfzH7
nDo87/mY/zTgT3iTkwie75zP6vaTIu9+1JhhER3QfN1cWpAJhMNRqf61WfOzved3
3kFPMhjPIdO8GwCR3puylc7fZgk0/ZAHhIyRznfNk96auPGawsbZJ5/5xrA9jJR2
9gQip9mQCyTf0mJTMKtcf+Sv9+U5FnXoPCKIDvuFzEHa7q1kpgPB34pbZwBwB8kY
63t6TlXdZVpNo0AtwLg2Ufy3JVi52Zk2u09+vEqkVbjtKy+o6xp2jSMlVY4gcQLM
31ZpkTpSX+rjId5PmvoUO/f53gYqG4TezayULMdTh5SJoaZjGcAikCzzrsTw2yjc
w1cdcIJIfQOawM+ME7I53YMy4ad9rc+DPfF37ToKstd9T/TeFxLHNYU6SY5D/Fx4
PVis7rPcKMH0rso00huLM0KLPFb3XuMUcikPPh7DfBBSsTmFmQyMWo++qmR3g6WR
Fi/21Lz2UvnxS3lqj7PNalC/8uvtCkEwIJ3sK0Azuc6htjczcvP9r/I9IZXSOm10
4F7Uw6EagoaeU+ncX0ChiV5v4C8r7LIidrgyb46m/76O3anRJHOOeq95GVwmMPWH
e9D6w7dzAVZgrvo9AAef9pI9zbpq9NrfnG5VjMU0QiM2cGaYICD2qJLkPDy85vBI
lVwhn408GrsCm721XIodbJppuz5oseA9+ko9CjdFUqsR9tmOuHF2glsYnlW49upm
ZKnTD9WKHESRyMrRF3tC289sFnmAUpQH76HLoRiIqIGV3FFKIBNRMLl+et2VT0vb
bqkrg/FsHqty2MI9xXEm5Xw2Sl8FCs/Gwk6q2SN5rOpDKXTcIOeZuT9PDbO0GqoZ
hUsZQIXUBvupvpxn/sPNW/VayMUVDxdrXtpE15bu1AW51KXm19PYZ+/I/j1i9X+L
sVYaytWaYAP0jXDa9AvP0c3IoqjNPlugrMZFZom/MWT9HySiBbhs69K+0WujqOQg
q5TNka6OMqhMCc3jw9knH2FXSgCUAFEJsdYAfzocCORUuer2nwNt36aSpYBNG91n
HrayHpjb6iVRax34TPH5u2TEx+D6WJfxtIzLWw2owfLsJ/00Bc4ydCea0NYQ+rH1
d2tauJF9PHKX2/m0EHhkkgb7G7JdojflzvcTBORlPchOsLCu9GF09GHsf7E+ssCh
52TgPPFEyCJYwTbeXuPaNQEZZjW/Ckc7g0FjCoa1Bf08h9duY0b5NEPFQiMvOJXp
blrfv89Vh2BQ096Zn7Kvas39nwwcEAQUzY8jiJY0UnUIbBWmnDLqdRMwfn9KFwzR
hr33nMReha49d1PWHEGikzoJNyfTSeu/peH9+VspoQ1z3ToyYB/Yj8AIylag9YSr
i8mH9ez22Pm1kaIiipATEfs2tCk/fDotblr+FxDLeXhRwKoRI7xQX6PZhIqGe+9F
ekjzCrL4eextLp8Kobutg7nqi3Ge79g39QnU+q4Dmj8kjI7IPsxA9uJHtg2XOfw2
JtDZurYjOpc1oJGqI9SBOPqoFNmMVOUNt4HfslbvZwT/N9ozHFIKGFeUZyenCF5M
HeZEW5DzvQ3XhJpGHTYKoT7VWNI9I4BMgju2VYugujFxgJjuz0aoyjYuzozVVbNt
Jm+4HUIhTEilx8Jmf7y+AIqXj2siciJuUzjEheFwXJ2bkeWqpcFwxWluYWfs7sF+
IcD009aMnxDLizU7gxJTWmt19WRAy4X5WtoVjwflkOMX04BJyIABJg1TXmD5nNVM
VATMqMDJ0WIRkS5DuHD+5FTY2goT7/oD8jTZPfPaf8dE8yeEEfY1eNM0n7vKQ7qq
1qvycEearkT6FTlORq4/ZJiyZ+7Cpfmer3F/spVXx3rw9kGj+Ns2xNqhrsgPTCTq
P5frVlIpv8BOkwdqwpAPK+s/OYIrGDQIDnuLR3EIb73imO8b7syekaSWBMIbvjo9
T9ijkfD64XbHU4wICHvw88l3oaisiapoMEPJDjG/P13pIGL85oQ0RPZ+bcgDgMv9
qzmwlqqDTwBDQXf7layXB9QiKX0WQUSzyL+JXTuSyGEf4lcDpxYxtwa7geePqePN
rFmQASAyInU9I4uh/m4oHDHIbUaq/SbfeWi+FRk68LmfGc6X2hwlJ+efB/E7jIih
pF4mLBB/k9vepdjBUtoG9QAEX6d5MGB67H06p0NXitx8x+puWH8dA6CcqD29kG8Q
kiCpH18JHz67T530tB/A1APHN/WpdaSFR0VQD/exFBvYb59eBWTjeUHXNGPO3JMS
5XmMxxVjNElbs8+rmeFbYU0Q1QffuZitv7/2LxFLr1DDJH8FSWbIDm1Q4OF+azy5
FVG3HLNQ8PG1xD+cca+o6mc/k6n2H0FfV86OEV/0/SBA83aeuqjqoxU6ppUNlpFu
6eHb2RewlRgCCwFCrd+RAgcgiPflQ75VSZiWjhDHHQbTImmzYWoSz87KPUc7jwgX
9O6CocbwdPlc2330xbpsZyWh3I5GjfZy/yX8o32ADz8a8qgasYmEVzOOlfLmgwDF
NeSYpZYK9d1HzmDMEd+yODNmAweR1BXQ9FC4Ze4MklBYXw6DZ858AifqNgaPOm72
5aGUVLFGEaBqbP6ayblc1a7HIkWE/rXA8YEN/5QdCxaoPv/HVqe7joAGx5y7Qw7p
Hl92d6vedt9wwzo8G0hcbFzeSkxnlpvMaGyGcdV0uXA5PJvQf2XPqP1fjzajw2/F
o+I9JlTmp4u0spVcAXaC4ZVbZxk8+eh68R18v7mgehNns7ppHiGQ0C/S1NS7tr6z
av8f1AkV0Mw93RNYge3BuRiKYUzMWkcCQnNo9rqiUT3Qga2zzYOWR7VwtYjqISKA
S01bDgD3I6GgRi0yG6gTURzSSAQpGgtVvgTiKMu7G8qzcHvHmJZQtjTOyJuzO7Kb
7wIVJGirRFM6lgpZ+Cv12ihtT/gEl32xaZJpyzirp0B/j6a8FjhFDAx34KAR75vo
b/nufeM4wE1QtLdLq42ZZ+becdXhXjHE85WSV47IhLa6LG9zpsiUykq5K+ZFqumv
AshKIlbBB2/7JNAzUkmGYBSSsakbZK8z0edRFzAblZ+8Y9G0G1G43GvTXdPBHgop
HsfjSL6W4u8ed7xiVt0zNe4zOInqH47ftixtJ9m4QidV5vE8L+PxyxVONZ8Xmzv/
Lu56evC1HTlhgBlCCILX7xagktjuLr2YAbdQJ6RHjzG2g6F5jwJVdz644LPev2+a
tnn/mlqDe/cPcz2RaYRpUgqQgJbfYsgb6zvlDukFADlBRfFoRsJhDotsupKt9z/M
3YuHuCoFtbuDXfo++H5DB1lZXyHgb2Ae0Yz5A8VwsNyRq5kAArvhXiiB6p6h/ppN
6gOGKHK/aEJYQwUDM6TjSUj7xi8VWqKcTviWzwT+1QRuCGp2a9MAGSQLtEYMayZG
vVTIQX4cFoq7Tc0hBgPtVO5G1+8ZoBixpuTK6POiPcYN61HPu02ZFqCxgAk4yb9N
ZgEqDpORz2eyE7Pg+pggkUa/0Pr7hMlu8em+P3DMJnZDm2Ly2DWO8iAAl6slMhhN
3mshSFu4BGdNeACZgimNQFMF8u50VRPW1UJuo5QLEDP019ku/yLmsyxu6OVJA8lP
hn2s+yDP+S6yY204241vXcSd7+wWUxnCp4Dfc/zSVNYml1Ojv8EfapaSSEFQho0o
roGk2gu9UiU/1Dzb85Ko1jRRiiaZWGwEvfolNCpbuIktjAbvNBZzKaL8rGq5+1S2
TiqqQMhg4mTSNSePZ0GsTiOiIA8JMDB1kPqRR1jFgVMVc5RxGQMyXMJiTogBHrPE
EcqpmPMVjIvNPyR69LefXCCUzhXPNvZQesqhL0uMVhLaeHXR6A5PVpdS3faldy41
l7g+1rZGFsdWYezcyWxLSUezrn/z5ALayZYkM6ORO6M/rtxR6mrz7ocKu7A+p31M
pQELki1AhSmUtNu8Xb7U6nagEScTdf6vUe0pU1A4pwaUgNNaINj4etFSrN4RiRAU
WGvoXm0t+zNNJ4t1PHuxVUoXow8pdzWZgu84u4ugdI39gHzAzlwcavIIJounBHlH
pVzVBv7yCmi5yOW6uhuVJGc/cSbZrQqRTQtQOVCLpH4pUkyQd6XXN0wOoCV0vLO2
soKjcxPkk7UIftmanR4Gf1kvXVJzHDpLmNGC0fG0hy3kCoP/YcO9/nd/vQ7XbV6+
6ENPfPde5WFJpeJ/rpZRa2lQjqMvyWMEwcis7XXQLJt2/yS09xVAdbMqtGpSw/wH
ZrxKVohtvpxqdYrBBGr6+PR2J0LMpJJQmbLsIA4gp/8UEtYt43NyP0hpofCmuY3m
giKuZi0Rmz5z8X1O4kBNGf0YyOxMS2VtDYZnvzwD8+W/pAevvVepC/6ucl5vwKWU
rkQ/cJQHTc6gT0aJRhyKAmxnE8zGKBSp6kigGwsmvDOKO4j/1TzvAfsHwNgfVJKd
i5pJ7GeVT4vsJ62+l5PqxPldIDB8kVaswUvEvdg4kcIrIS6Ml0iAdXAMkGwIsy6l
aw+mPsdZ4etPzDSbaRseJ3K74rPYVbeU5CpA9g7FMf/rG3BJgqJo86mNiFFb7qB6
exAPgb/BtmdbcoMdr+8ZGZ7ikTdUTNIhmjto4er/DjAZ0o2XoKSQg+VeRWu6ejSy
OO9jsGmg/lonASqLE9HiOw3wi1uVLO6531IULzqyi03TxJR8rWCOQB1Mc2JH9pH1
nY4fyfFPCt0IZ241pwEL+FvZscgfn3eU38uWvHVVsShGnGe0jlGiOf8JkjiVzn8j
pS3JHTq1ljtBJGx5Qj00apj27EOSqhZyO/X5QP0K+jImltG5DoHPgAYIFWf4rfvy
33gv4IfPilZX2SRqflBmUKCFbTpbyx3QkyrUnGrsWswwbSx9wwuLfpX+wH1zdavL
rYMAKO4jdaqOzkB9R05EeOmqZUNur8InI38sF2o16aBcDGlcZai8kSI6i19XcNbF
CcZLjkf0c6qMoSjhkdLpfj3o5K8qZYACRIWpsXg42bZ56md4pls/yVRMwLnfb+54
3GUGupZMwgTE4WgOFQps/lGDM6TtGl76Sa+btZUBRVSEvdz4gwE3zcv4alAdaCMR
ftWzSNn0pq/TC84lS/NUgq8S9ktQNS4KhL0WP7S2errqqwOqjU/MtEcFj6+6WjCL
iHkg+M9RuSJxUb/PtuO98PkMvmAaiNEIvzEeVqvdk3zsCW09QoKJHSimiDrU6EWe
LUi+5Q7oR4NPlA9kx6czbAfC4pv85/wLiJM47qAVt2I3IUcAif3WlLamTH12lX05
aft/5/7/WZpbpzrcNN1aQHyH2sAm2K9ys9kLFjB2ZzFEpLJfTI6r7q4cokqdD7v1
aeI9jb3bPjvYM25nouzjtMXqhYSytASYxx6hNhNYF3QffBkj2IWO5JM5ZEP4YrdH
4lUZBFk2vYqIVkSzoBmJZ4ON5CYPFa1+LKLEW7G/zxbQJSRZa4o42YbC2ttA8/7x
9cXL+9n8bVfrzor/Icw8dMOnvk4DZHA4REOSrpBZFn/+Ylqf7uQfZldgz6APaswb
eoxy/Qr1lc1ZyWwrJM8W5Fw3/1jYXSyrQV7i5Wh4ncds4ASS30FJzLucGK25EZJR
BDoA1FXZHodtm40DBJBihTgVtkHz9CEE3CNCRXSdX8vA37/uAutq+dHnc2fjvNbi
InETH5OJoWXuDjx5UxeIKGJsTMiYCJpJRiHOC96/6tvOVja5v6P75NY7AW56HuLU
J5+LJrC4eTevCKwU9GcE7RH/1flHwKc8FQAzW5vYcw6oIs7uIKkGEJ8cqydbhubl
c7UCIGIhBAayObI9k6aA5yZ+PTm49Yp+jPJtUZC2CHbmTCLE2ID8HfHtBznvuYME
jWgmuS0lHRLRrzek6LhGwZcwBMNGBWhG06Mn5jczAIHDu/SNPLWky+l1UqbvRd6l
lSGqeibqc306rCq18+976JZJ82DUBtPqtw3syThdDxIwoIhVDUTk5e0yInun8Q7b
J9Gl3lFLt8Ga80f92GVKPpaVb4BhE53xjdqZbM+UpXKTvgfnPpBpznCRtxsIxXYM
3onh6XWYFIjTdAYdkBhQSk7Uap+W/CmIFoZTNEiigXZr95wd1dQQNOcG5rlbZ+2f
HKwbxAZAlaw/QP2Aiza0EdAztpdQwED7SvsFhA5eBhVUoK7dvDF9mlakeJIJx6kG
qr4j64bp0ww31ZVMbDus2Qcvy3Q0L/rRfViuY7bKYtAE8ydQYRuNO6vo5eJt5cPO
9L3zbCk7/s3Zj7tpIvG15Cj8azxPCecK3YPGLsFRwUkcovqwIQgYNG6Gdepalpft
0zbOWPYwTR76PbIwTDkTm+xNF5QYu1SEkidCI7YoN7BZaGiHxWNb1Rq9oGLwa+SU
xAZSDFEPlRFV7/Qv4mfWakpZCdoaquh6H3pvXHbiqlsVib3tJBkQuIOfIHt3hqdi
nl6tBe3zKw+ESKaaFFf936vYvB1hzZSezMkT5nOaI0AeJkyi2FI9Ao3bG8PH/50H
z+lVARYIoWjfm+XKYSaZC4CVzvGvItYcCoDvrWxhYqWKSZAdh59rPmy+/AB92HtS
PdAbLTZ8uYanYfeiLM7oAuP213xMSwYC2xypnzmAASZZqHZaqS3g6wuSH7QnPBCG
rr5dMgxV8FhfNpkCWXp5bLZnBSWzdCeHI2FIzUioV54xqdqB6D/Nw02rAB9ayxQD
jB3ilbBBO1Z/M4fximn2fMvOVLPwpqN/e2saX/QCAy68kCWzTXwctdr/ydeC9kzS
mJM94n2aJk954XKGIwxAM4yRckXrJKVNjvYMAFnc2vzPt5nrqwEvV+XDd8GOPpv7
K29y3CyNndSUHfGGfZQAfZ0woqf09HwDREZ0Vf0AM5TCynbVbuPez7al+ow57MWq
wly8Y9razjccrL6HiCII7Y677T3eoT82+YKH7SptwZpjuXzrnN9E0dv6/anrCbxb
5/2vsRuVIExqR44EgLN9kMBsDaQdVUmAwxtFh5fBGAqPOFueJlvxz9COwgmq/9bZ
BparVcd5AMSNkoCPzQKlH0uov9ld1gJb4dXwVRikpLlm0I9Yb/83VHoXMOdJQkqH
diAC9aHgr35q+omxqhHpu90mt92uu4ul+npIvM1Up1e8tEXhL6TcU+TqI/XEXVO3
RQ25+bBbyt58Lnlb74ZTij7CT6sn+teJgmtYhoQQxXTCqCnuyb6RUrbIMo85Yuuy
yQicm1EqiVdTwkOoudCm/EQrmN+Ppr2gVWDi3cDj57G0Lumly5AIAAmU3sZWJMv2
QK62CKMHzuP41DiP8K76o7rIO2mpmvCzXLuXdbKvoqE6g64Ynsx+iJHHZFYvFQZp
BuAybHAhvkfigNwgYD7TK2B/HHGOPgvkZ3Y+sYMtxXHevfy8ztAPFU1/svPY+Wej
Fjw/SSpYVxvotWHzTj4mPt6D1vtbXfq0d/IvfNsI9wa5cOHf1FQ6AyBzwFCKzqUR
HPOE89pNLeoxkmiStKPCb0c/gLobkqBhjSjx939yWMHOw1zoJT8YhpqCl2UaLe1u
oZ+sPrXQcl940sNHnpbUZt17fcna5KQhUW55E5Cy0bar0tHw/MdvmgTB9hfcyQPC
zzStf9ZTj/4Z3FVJDv5Q8zzh0WPKsU0zvGpYr2CaeJfQs/D6KJgjpiLUq2KXpa7t
DyX0R4znQQu6i04JkdOfstVZAHhI2GyDUoZ3r+Ka1IRVRPb6pnpavvVMtQqaIOsi
eBZOEC5CnccfuLstd/dETIuMAZtpH/IpqHxQR2HozJcNiMNuVx1Ntvy6Bb7baUOA
naKnuAZhk+mzsl7GtbK6vjKeg9HXH5zAY/IqW7gF3qFiG0j/aQ8fmNapLav81K/p
SgWCofbFVv6CbG84FqFYcTgMNoIXbCbpv0lhpDhMc+8HJWcFG35uigzGKdimY9dC
8Sg5Cq9qdJxo5aoDIv7xayDQlZdDFTXRwGqe/gNSfE13pmQ3h2HvEvpGVZClPbZX
LRpUhFIc0lfZdC+ioZhDDWNDlEYaAajnDKMgcQ837ooIoK7QDZBstWWyVfxxd1Cs
jmvdRjka5WbX1GQIVMW/8m5njILRiTDQim1xblVHLMrLznF33CKLpOXJtUBEAvx5
vk84/n/xQYXxs/kDnWsd2ZMOvC9zjDIOYHPlidAvksqwhnbsXLyMMcaElB5zLJyf
GMqw1LXvtG/ROokCRqZcIMsM2dVMrxYCI4oIrVjPlGYwV0vsHRktGxM1TBx+gwV4
jEgXsECXRnIj/YVp3w5hbZN0SwbwXiCQFZgRcZ1o/JxNpgsPklIxzDYh356qcUhU
pLnSR8pyejxf6PfJIXvxRW6dO1y/3qimz+b4LTBgxektD+fss73bYbZQHakx+tjJ
P9jgpfeCP+8mtmCwtyd2RJPBXVrf/6/OdimK9o7+8lY/Ek/VPTrYTinPuO3Nk/3p
gWKxMMPEX9Q5LQ6YWzJMQAahPLgXe86KpfpjguF6PJaYi4toAAkEhaDES8bLqCrs
uF3aF+BNXyDxkV7lxNDmpdho+vly2MD1y0EfDwFAopBPPQsQBoM2mykG6HChbx3r
Smgy+PsuWeFy5VY9Penxk3yWarD+i6PoVIPVZEn1P6cJ+rOy9T0FZa4ARJwA30gj
A4KexCXjKfE/918iCUIN09BOCl+9k5yJRzTy/NBmS3pEmA84Fc5pj6M9lTayr59f
erMrAie7pa9274lNOtifJs27oAt1RQ6CvaCD5CsUdyqpzZO/fJujQsOWx8mh8nPn
b/szKfd1vbI7LygSXEOQNus0lNJ+stFnRquRdvvrtY+3F3YF8C8eIqXFmoLexFgZ
KIN0igovl/Df7xtnZoCK7rUFSjMnQMfgMc6hgZWvlAi0zIs8ZBwZ6FPR9mJ+kO4R
eeJ+0CtWQGS9T7D5ecqiW5dTtuyopMcjSTe8gwuuyK51QsG7H9bOzXgXLCJbPI9g
ZTP0WQv119ZJP+tY3zWbPvHC+lbj4ooaQ/5+KeFmA53AdZZqycFAdEy0Vyh5h07Y
O6+cM87zSeLlMfEBWqAx5jlmDpeOHuoQw3sp1EbQwcP5Zv0YA1M76owFb1aNPQXu
bNNpNM1vxELvpPv8BzRl+ne9Hd4rDCsFgQoCiAKsGqoHgTXOd8dsHYibXdFK+6F+
CkowPmE+ErJjZaHV4XAUhXvGBNCONFnnr4wtC61uaogbB7BwNyH2iogHoJz32djm
sJozUwkEmiYHaajKyrfHCFTruYuKxjgr/oE7S6uWrqXo9CEJZB7EqzjgbSYYnnC5
/je0JULz4HK2jsu4bXMEP8QJUGqMSpMB1OJQhuzUYcraFrGUApJcG6iGWoyzwUpo
lO2OGpT5XIFB9L+KQUVRPUOExl+ZsHwIrnyrX5QYXR6iQFY2FTJWNCCidtD8gKKq
qGqUUKXVgL6bqwqYb+CPdaZeW+ZeKYou10G89f71UILpOZoJjqd8Ze+NrDTSKi4q
q5juLYawwNdcp7p8WYDF90UR3DZWkPBdy4CW/RdQo6+ep1XP5L0pYJrlFnxWTgXx
H4Y+Ae6zLzjfG2+aufP4YzyrqSqD7yVvsoWH6souAt5F991C7ktFgLn9RRrOB0kS
dRGnQcO5IBnaCoCADDG/f2m+AKs9heaJzlyNzXVZQ2NuKRyV/MuK/i5wJB6dPNoY
R2Kea9le4L9tkino1UwQyK8q8JiZV6ylBInUjWDf3pJiJZg5LOSW8DofANvdMz3s
bc4Ol/t1mKIALoRXHBQ6Xcy3IFxuN2yaerryOpECQRX5P8/6+dTJBfeXejOhQj7Q
cDGjbjjX+k+UyB42q3w+blLShixjnkRQFQGkXOl4MohRKpUkr0gkSeWfWLeKezLy
oOEo1h7DvuJOqAu8e4gmfYKg9yZQTynGBjWXJCttoDcBztN1rVAU+jKI+nNwrp4o
mI8q+WoPZOa5mk5GUaC6wXdq5AHzrj7sZAJX84VCLWfA/5zdaXCObT4EPfjMs/l2
3kjT2fkLm0GUuFtU+CiD5MvcJO0v67Aidl9ODv0ISbxGIZfkai+ZEvNB6cu+y7k6
B48tHoWm1S11okmJFD+0GELgO73MFZ6z6t2KzBZEiqOVSdsR0x1clnphpTfzs1b8
hZM5pYv9YXW5YuP5CNpO4gxlXxFcWxTp+ZXJ3BC9A1qotY5REb1G5qPMKvUXUql1
hSDJDfa+gTMZz4nNWS5XVkfS4S7ca2x7VKoL99hkMDbcwcEain3TVmnTTbWnzetZ
EbVK5Dw+rniU2rvUAA6+lsgmpMKYxoRjpRNDftWIit/F/6OsEOEkIYk3sT/MbcT5
9wth8pf2tNs8uGpXiuLMB5h1fEENKr/puGR1hlLzyO+aL9mOnbAcYOkf/ixVRXqp
+2JDI/9VzPwvnCrRvSUcF/mSgNlDa8WWBn9M0cbfDixlj6XDcJQhA741WynkDKMp
BBhh32v7fkMkjj+5Omh3hA1dGFC8l5aFH0HKypg/6LWf90jVUDIHle6e1JakpAuA
SqxZBR3jIlg6l0mMAapJnirXSk4VFRY/XBohOp8zhPtWKu2YpVLG8JWCpkyVtW+N
vBhNtVbwXYJsgtAPg/uwFfpwBlEPPwemHU7yffJwYvzBGmXVSG0vghk/DO6bhU7s
B2B9AeP8+uHptyv3anAk5RiB0j1J54tec84NMABnLnEXZJOKrb4MYpgcFSKiioMC
3vr51Krgo454KJw1yjNZJo6FCbycRei2CYRnx3ZuYwGdTBtsbQBL9+YDt98eMGEb
aDmPYBKHrErA0d3lPbO/vFd58caoZ9Q84YZNyi4vm4vV0KrC7lUV+ycZp2h2k27X
VWAXkzTRpw5Mt0mVjrwRT6u6luyWdDE0/xkIu0MkklVmmd+WlZno4JGazrRmAlfT
wmtG5jRbmuA0DqVPSIOoJvfVX8+44QqZ0zRAcGPJsMR1P213euCAR8A4QB8chAFY
Q5D7P3gh5vCPGf76FBAl3UGUMyZ4N6TNdw6XYh3bqNKUzLQZh6G0/upI7XrWTagF
O08KP8HrubC1MNQOOWt12K/nJjfoSaAARPLYLUeAPgnzlJpiM4UOaYceozcbwjj3
rQTOzFDlF8INEVZiYPbLjeDXdCOV0SDFgSSwZFap+OWXBRVI4xfZw/dKJQ+/BM9t
jLijFiXCt801b4Xg1eYZDa1F8MEFZl6/cii0GVzMzOp5KEkdn/N6f386iPYvCnWh
qxdgKKOqdgWCRGrK9ctdwk1tImmcIEZWfN4hHUDACvzFSFtasko0ZikekFE4Omvw
M6aIwedBqe2UYDsYRpZYsYCS9Je829PtF6ewT5HHTskQcEgRxgzO1+0D3kl6/ia4
F+xqmMyzUJoHw+vZfLhQ2KVsaEB8z9M5ETsyZmJoJkn1Qd3Fpt3Wg4NxhAgf8bVj
T1Zwz9Oj9SqFYgO4GY+8Ed8KX84127r5MOH9X4WKImXin7W+m4t/+5go6TykxDj5
9n/Ybu3glKRG49SSY8H0YK2AqxB18VI+WAYvkErZXULz1GvGDTM6p5I/65FcqPfs
Bekj/lwZmgEAIm7Z8DVCz/D2W91IJ+1oXEPaNVJKXH0Upb0+4Afwp9Phx++Bd06p
0GmKS0YKCDnbI7Iy+N5j0KltwQzJEgWVeTzAfb3c60Cuc7uVTdTO+avTltlftMdk
FzpOT7o/hRuo7E5z8Iih9uycZ69T74xE3W/McGpmMQ72xOSkjQu7joLvM+odFG9L
ZhbVmH61QiqGy19mDHn55oMYRm+AkMRhEmnoGcNtn/VNKR6fEjLWxV9sy627YCZe
bM4wKEHPHsJyoSPEUAejRGG88RlDgQonhdV0zELuOKvvX7uYP4X65sDS6pVjxADL
tfMUUcInFWMZv85Kbhq7ggBi9Qtk8PBgLMTA/SAROol9+PFLHbitYDQVyaYwYuS7
P1jmzi4XUfs0PXflaJZ8nj/ahTjbjc0jjomARHtw9d/180CokWCImMN54mvo8Tlo
roUlm9m9I+5ny/894ZHB2rk1cENBKITnP2cgOgDDEfqbdUlFiR1PEnbzf2G6A0Qw
lJANo7Ac6P6/XsLwTComQPLuSd6wd8TsYVNnowM8hQ0hUA3IEYAgKfROWzv8fgXb
9iH6kyrX66RVCm8o0CmCRqqBG1iyLAeWY6/65RsFVHoIsySdRskRVhofJDRLMUuG
m0yuzZ8mLBrg/zPc9fQmrR95uuqfy9MGh7Ue01V2+fvdyQ7xRZsCWnZQhQg04c5a
45ECuZgkU30As2AIkpVPfdZBzLjruiIBcsgVVV554GavVgDp39Uzr06IvxnlKESp
VFGi4Cnc5nBrG55rICT2rIZIoOigsBptR9LDV4F2qVSCyTLDoSj5MXiBA3romKzL
vjWfkGhC5unfBjVLyA9BqPHV2cygfOqa8IxdC8FRWfnqi387yGFidQQHJXIiyg8j
U3WExdtp8J7FhdqBLILf0hLgbIX2qPQZnCVRvGWV5Jqu7JxecmyiP89S1sk9WVJR
gYZsOSkH3W71wvSpKWpZoWLg3YXM3VmlU5h0pom9t+rIzi1UVkmW7L9mrHyC4UDh
wIOiGYiOad0KU0pmLD+PmpksDuk1mPrMebK1i2nFd3iMf6l0vXckfkWLBhNFZkLt
QXk7wFo0lPgyeCU47HAGWYOJWmDqV4yGzCj9SBVx/8YatyTDa8Ju/Fl6Ldlxw4vY
MMOrunesifvoyzQqx2BJhLxv2aqvfbmT1Fr8UkXpNlC6X9M1d5eflj9uJBf7g7no
YsQ375z5q+li6PJLer6oil0yLYDeixJRFeIWm9/txaFC9lQ3uWmxZBcBpJIGmBTG
0gvNV8GLcZzCbKKBjzVGBfNylqBv7+j9vkvxWajwYTLD9XEsySx5DS7wXrD5eBJN
E2cK7i4HPV8SugALYPhpW9z0wFeE+8FBt6gME+TvgZz+y7sUOWMo/1I723atWA8H
NMPm3Y0litmOwUFcRZn5Hx5L2Zgew1FMtJXS0BCqR/tHQ/P5vzDarRxQNqvgBojp
6cCBM4BzSsFlhi4EBVuANLhd5WrSAcUueEv/riX74e1S12/5AopxTgVNreJAVSrK
v1L1PUMgjTXzG9eRo80UFTxQsQHoaimVoN3q0K3PSEbkK7n8uPsEyHN/A8Y/boUS
TH9rVRDCP7VJoC1erLcP+gOSOoM5X15wVz5fqQcFtgb+1Qoo986z75LJP9ecb2ZL
Zlxd5s53639VUDThcZGybKClOz4YuRQD1JMIX2t4Vq2cE1SQztpOqzR1QtzPSvZb
ocQGRY2ry/POqR9v0WqTX5wIt2Ymz//dVLr6egpjOxmF1nr14k//QYKc3NKgFKhJ
Kj0lEzzSCz0zyfXMLmgiaOsz61M3e214siZmNu7E6w99yhRjOm3L/AZ+Z225pVfE
arA2wHQWGcoJpRYpu8ZUcr1pDr0LD1HJ5q+7DmBPEIJoZY1Trlx3vt+Nj8g5Wsiz
bTKXkUAM9F/ajOnWTmASzlgaPDLnEm7Hz752h4xB4AO0hDMyHNynYxKZeLnOJ1DU
HMy+wkMUUh9qPZWVFAQEM/I1d95Ka+7y+jdE+jzxZfsQwZ4mJTsUT5nmRj3iZGz3
sNqVfayDcjkJY4Ha8ZuJ5/NXMI5NdKBCQ8qEOZW3ldFuMMHfY8uyMznmstvA9tha
cnba5xvN1aWPKa3foJ6Ue+o5SLD8oWFPjdhn8JjeOcXuAvvlUu+RVB8TG+PYByeZ
MyLM8GykbEhtmHgsENYXECEn+aCzblNPkRHqMxcjtkxT2pH7PuR51InxlVJMZcAc
VY9ZJ2YAtVpo8Cn7iJqsxlXrxQ0m2Mv6beJvxTw6CjV81cOi+Wb1ZNGQxzLWGVQf
WF/ZawfbTvZWLUhpfE2sfv41kiDjcPgeJNnxryilv+JpMcQbWc+VEGa2jyHx6pBB
JbE/j/WN7on8xKk/bW0PJWctCAYbQaNp5Y1bP3vcJm93aIBPbGfh5lbpJxv348+G
+cyJ+oCKpmerXdMBOpwqpOnDNCCajTlUddJs2zfowI0efHnmthzpafIEM2xp7fS3
N04/AgxU7oTUr5PfM7L/HRKmV7fu+0mWfHkyPS5RbrEnCNjWLRP2zoLYDtrd4ggP
yr2MD+skqmK1FPKmUuV8q2s5FXyT7a4Za1uKvR1n+AghF69Mo12GtxgLtvx7j5An
6OGT+tH1tfuxtW7wNyDKN64ILNF7UGvvfCJYO5W1jr7ui1D55MsiS5otEi7ZcWJR
OS490Exv/UOnMsRnYUCewS3RlGsNb2/ZhS8IS4Cn5cLBoMvQ2Lmk9SihalbpWeqP
8nGa7Y4opEja1Fct+XQatKNMK1xN2F9F28EXnkHOO+MSjDCMuwFKwV9tqX7P1VRn
gJ8393QJlI5ynuTQETTD1GWs2fEIEK0uVLTTofSJVAUiZjM0A/qvA0AcdmI5kiBY
xyeQWtGZ/AXumjoN3pNE3iC2p2oAqQhFsH9Fpl9XwC9L4f0SgPphytr+0UY6Sd21
hL6dhVOYeW31j7BLOmor3iWAi5Mv4s6ZlRp/fH8Ir8H3AUkz/cpWVbFJBX9ZCpBN
hRbKr3Z+HEiOmaCXA+ZwKq9t03zmATfPrnsN7vFnIVTuy5Ci2gnLvwK+i58PMbCJ
cJy9tue51sV6trSzaqNxDjcO3s39s63W1kOPL0XKlhI32w8UCbNWTVAo4/n+gLdV
zPVgmP4jmfM4wqZHct1AH2j5Gj59HCIHvx3qDOaaS+A0ZNSQfR8JSj8t9qXtITpP
14ba1R73Oob142XxhFxy+toRsxxbLO2qCqpLioFNd00W3hmRPRqO6bN05BBy0S6K
EtBbQ65+rIAYfuOdJ8hMoQPpum3SQQuVM5B8pKpOCjSUZlp72wGX+Fsr4yOH1Qgx
tEfiyu8/Ep6iYfhFCyp2Pj0x7BjRsEpE/8biI0K5pcrdX64GZj0riEqJXqnK8AAl
UxDuw9WrvCGKzdZ+H0nPh6IhLIxujE+E/TfP/+WTf2DS1uPjHG0geVqwz3pAYmpa
YJYJzJZV76YiIgtvjzVw3Tdl+m6Z3KS+ZE3VA1rOEgZjdfpUOMxRwmHKry4izSzp
zNgSMQPTov8cU3AdDq5KnaLnZfVGbSujeOOHDMuegWmTIM7zeP3Hrm1S+LslEfG7
O0Dy7Xo26b7+JETHVwSf6aPTkcBp4aM0FVxSfJuBwqvCiuU2eVy5C4kTooqtV0E6
/rJOP59YnDad1PVj1rsmLLxSHTYOuukR2KdajOfebo5c/pa1rLI2aF6DAdXgQFVr
mdg7kYjGieEp5hc8k4ArKWuhVP8xkd9J3LfMEo20cHNG7Vs2IIVsMvLT0EiMjPm8
jHrkfIgHdTGg7OouBOUHzevPGlXFwzqF0E370rqjs94gFanztyyavbNjSknG2hTV
eFPdLWewRDTfWz/ZMyGO6p17hwjtZVJMXZ9dAC0e56nohYSUoKWKXgt8x4YPC9ea
UUX2+eqcZCurmD+Qd5ylegfPvr+ZPTYaHhwqFPaRYcSqyPIeh2Gkn7JshVCOy8QQ
ablFb69V+O67fms2dcK7m1P9Ch4yGVbeIIWGYOG1dvsK271GGYTwy181vJGqd1wt
y/TEMD5ZPRpT07NBwP8WNyYce+v1C3rqTcyCVbAOwZ/G+9ofyvAUbs3Xx3nDkvCH
/iCtFBqpg6C8cqzoQyrlxhhDQDWyCLgReOpWOxhLcv9yVgtmud2si32gQL7c++FM
TOnP1TC8TPNyzbkWF5kAyDB0Aa0tTQu13cekAHDPMdb6N30zCfjp/pZi9PbGn2i3
+4htrcs+Enma2KyNt+P99ZS/NBp05gvJ1BBgNDBtUFPpQmE4m/z1DPCIHsoii2il
Fwakma2IKZ6egfWSnVTvaDr/J7qjGg+TrnP3DzLyuUcmJaDlrsnMh7Wl9Cvq/bBT
VfnvXmX1KH6Ms9YQdagr6E3OKDOaWaV1T85BnGpKwpR0m6LEM5V3wcY9s/dFFffV
U+b9LAQRKjW1GT9JKIJsUpiU6e7Y1CH6LJaXzBrMo3y2yfZ0RAPzT76Xt9uZvZuY
/MCErJOoVHnRxtw9GikPy9LeMKe2jI/3pP0U9afunViiF8osfePOSCT0D7QsmoFt
QuJM9hS+rjYPI1xdqZi2bgxgQF7Bb+JNi23gQ/1pc5d/kR0WbKPEteucPxai+5wX
Dh8tJT2oX/62PC4PUhRy52r9VWlqNXP1MZXhfB5cPi3KupsCJrEUZB14YotcUvUI
psEy87III4pYESg0XZ+i/cLGoZRKdAtVUzrc4AGJS9x6fiLhmIt3ZROK0zUqJuJJ
OWwwhVyPfZAs/ZlzR8tsB4jOACEHsrqULQjN9RX+WGVqveS+7ZdDiVTyZMMbEDP6
YEEcxt5nIFn176nsxTLVWH70+Rd5GRQmxblnizlRrnt7yWQQzySKsJZ9IHWVzE/A
ht7RQPV9768Y03AOGAPkD03YKDdbYtJQYYgUK7e4Ldks+6MrR8JQ8A5jQ02GBvn1
wG91JrpZ/9XZzdBZ2MVQ5zxX/0boeC0I7BbuYo+ECKLu9C2L5gSdcsaFaiHx1uGl
RzqYUbHwZNabUOgIwShh5Gq8LyoZEPKiX5gtTAjsym6+3zKwXuuPA9E/6HpVwvVL
8/rmnjtJSb4EAV1gvoSMDFI52jsUGBTAX3vza/FQriwR01V6QNwb4MdPwAQ5fWer
+fjxhANgOrBP018Diqp5dgRKF0MqkNdTpTt6iSYJOtCmvPLvpxhHG0nh707WeI6n
NnETEhmO7DsTUp63S1lYpCiBsX/g7fHowaAwvYk4LeBg7YwkuJWUScQB0/VfPVuh
P0Lb2uEBZ/gixgA5zq+I/I78T6o1bRweYJTx08WsS25MNkmyg76Zbir4a2JGL2sJ
AwsAlElUOtZgvvj767Iayphtd2iT7vmd1vJDLuynLLhEp8NNRJJej0MoE7PYX8Jd
zU6saJQkNRHvrA+xy8RNTOAgH/iBi2l2LeM4YuwNldguwgRZPsSZVAkXLSmu4Jmj
kaToYy5k4cSaTazpeIYvlSNlsZ17sR9WSmkeBwknBqOXv4MNA/iHFBomLjf7aVcR
rPkjnvcA9uOWZC9Or7orN83rVlv2z1QoY3QWSS0p1WDMYuvllyH6xkiUicwvLRRj
6kubG1+D7MhoVLbukdC0snr+LXtk6GnFAMyiER647ymOGNT9MlOezsJSl+cSy23o
wW4zu6z3Z8r8KkP64hiu5XctiCkunRiRsXOAqWJckOsGQQS2qU8PLfR0ik+2UdwZ
Bt4sfTRnWgP7DnzvV3j642Q5/+4Oawxjju12bt4gryxMJP/EwfshZEwL/bjvpmbL
44nXkR7q2g3IxRIDUQ0Sh/SSQrp0m+LJT3ng+3FkowjGjEDjpg9IgyUUUsq9LGNn
1Zl8Stpv3KeqsF4fFYner1JCG8ReZmo4HcpghQsCRUFGYQ4IW3SiULJjMDvEY5Cz
J7DSltXbiliqF9+T1idybfCMM0pcGzMEu2ED9EL1BZnIx3D125Oa+YBlNcAl80Zn
OdPVqIdP0eoSSYzxYFK8l2+C5jNLw+qIJS/36dG5Ci4a1RXm1b0G7/I4h65mNllz
m426DjOy/hQ20tW4XPy+sarzj4BYam2bY50p0UrRDVAoSFs7Yk/qtXJz+j7BT+mC
AMICotJs4AXEIAW0D2caYnwNDwmfrzZJef7+JhwMiYjafVnp1mvm2quduFEirLdQ
hKS0WZkqxDnpkMnORv2zbsrjeuat09WG6IiZvT5DuN5PzjLf/3DcyIE92YaOUHAf
x/HSgnoQXJ+96FEwv+dSkXWbtrWYNT7zK8L6QRXcUnQeQokvl9TtIElahhCSqHfy
cIHehg9WUxinFDL8BNs65sB3/JTTrwQhH75SR1ZYENPMnC7GVaJr+CIjfHI+3FHh
7KgTfbGhiM6VYeOSMLauN2KyN795RJ/3r9iuy2xctRu8y0l4I/+2R5lNyXIqXxU4
Af/rktTjuI/k9oxP8RhZGAH5qwk9m4+yXLSUKpuFSfY+LMjCA6HPGftPNklBRnnE
ThVGeLJ3Uvorvqm06sW7s9dtOMFGRqC4xADhHk6xjDlXEv3qAfOwj1FzSBv+4sW7
+5o8KtXkDFn+Tg+7zJgtv8PM16bkFdNbgPi7r4vv3vI//9HEuX9IwFexD4O+AIlv
jtoe5M7/XFgMHXWtXWdcDE7SFfRVsMjtYWrsSmj8J+TnsFmEcIK1fFbwRkqy36L+
Tfd00Hqzn/3hW9gvPBWy+f1x3tq7yoSQWQlD9VlrM7bp6Q0r+czyc4OvLyJLBsKh
DvXSS/hFvJKHVZniaNcYPN/CRAwkQgRyYD/d34l4Ph5uD7yD/1UivdWmneXjPgXW
dlAanZFctfSeY8XXpKgO/+WQ5sAJ+M0MlDDXcDNg1eRLb5LWapd7E/Jp0ksWnir4
UQsvHIXons/pAXJm88oNYz2ixhTgjyUdew5B+zYbVQD8nnqqjqXKIj8j87dpQQ3l
K8zsKnADVEOcuuuUmr+2g6mXeFFKjPmaRE63wfnAkvkLxLKICzBmOvV6E1ZPuw8G
7kjGtBtqP//Svoomm3TLe2/1pj1mouvsVOupEySqLDPO6o1rcgs/DZ7TcSjvwgmh
obVAgWCM2SYMUtKOb6lGvPWTQSpcUcU5hJI7HM2C7LNA+e5IucppFY5QxZz2wrcx
UJHsbKrNV2sGnirkv4ekxDbBK3iS0IylR/JBs3ZxNP1pnA+oEsEHI0TmaNlrK5pX
JyTZAVKuHfuPkAD4bLy2TwCYJfiub76oX8tWfYVfK1O0KScmpi4SvmU8bEJePpoA
J3E8zNuJ6LvEt7hThvFo+H/T9V+Armf/tVguyo/3P5fF6Og1Kj2xlbsMv7jxvE+u
Um+/snVJsj/h+aBhH1BldSALp1+YXeEIA4n0kAkBOUKqTAHnZ2iTbrM4hkWTmpmJ
nDfgK1nd6icYTtuCSQ4s/7v/qMyijjBudDEhfSBzKY3abTGniSV6IEy8KL6XBlE2
xGlEwizmcMt7WWk06vasy2Hdp0f2s3MBBz2apApOR6EDtAyHViJkQXoQrHdC4D9b
+2K7ASGgsEqoHnTFUvMVJLniBExoyXriT0KvaFUeXQVsFt+moDtG4AsMo9Y0EkBJ
kK1g8Nx0Hhk6pGprxVQE3XhngScExVEgNpXZqzxMYD57kNwQ0ydtYRsPjGHHYjZx
nyDVVLGR/1lIcNkZ937j9m+2duEt2IEYULMky57k/YUS9jgY2SztNpyQwwpnlq7F
vmr6yohkjRaFkDoq4Tw3C5TLVUXoYU4w3vFfS+6wFAq60KLxyoWgCB12YJOlmaey
/96+jLaaUsm1Tgw6aHo7iDq0pVIDc9fqMdn1z9NQr+5SmaB/zW/oqGoXVwInNCPv
uxCgdwphPZBovmGo6sZ+OqV+QMggNMedbUeiAQheKbNiSUgB3e8eGBowafIaavwk
UQ60rZoKYWxk1Dwp7tsFWP4Ckpv3tNALlDNHYhHDnlpibzi24RrfPyLyPNawO6a0
yOzPp4tkNVc3AMXaHe/PMhTWol/ZejV3+MyD+ppBEH3O4naGCebFMdiwB/+w2ziN
s/YN1hPIkFsZcpeVcOJNBwJ2B6Y84pJwh3nhUvkDulAWz5cxhyjVR/N7GEuTKP15
wqCTP71JiUGHTin4C1OcQ36Yvfw6waCR9YOFv9vyFYBiPOF0tYv7o/8pwIK5GC3Y
8V6w+sUtNors2WtUHbTIFKkn4s8snVI7biRT5JeNHbIfCk6kme8KmdU47pCZq51/
8HNjgl4rXo+ojXy1vMRHk+b7gKcyZkuBRI5B2oUGdFV3og6PJNhBX7OyIo593xtD
Ljc/NP983+ego+bBHTIgwPRw6yXN4Btxkwn0LzDeaMgzX0VjOuVrpUlvDZp4+wjP
JwtJMshpNOAyxJIchOxPcAF8bgGq6rnKyek+ksVgDiUrryVjva5KeFjb/2e+hK/z
g+w686mdOZ86Pc0gXzR3X7OJbA8K0YxoSDO2Oj5PaUOKbisbAAWnb6sTVgtvl/f2
vWtU96Rum1yhQgV9gLkwdudJ+fkGDrVBXwtbOwBH5V1NRU8JHGqeytSYOMQSUgWC
hsXqTd+S0y/I34h+MLfQVf2Yt3N6lLxH9cK0BxyUCmPcWKt5NGuV92X04N2yNh7l
WD17Pt71OyNtQf7VkjqqblF74Hv1cSloVSHzGvSuUxfPVZkCIkdUFuA4lCiWtoDS
n6gx42RDDLYJXhKaZmI/V1H7/gnImX54CixOqA1FUPM1WEkTAtE8HjPp8B/6vdZa
WJi5vIT3uizhqm9ru7FoJT0BzzRRBDJqKW3JK9z2RlW5nnoqIsg3PVwpDzaex/MK
ITsVqbc1kG7ex3l42h7/DZcgVVM1npFS8WUi0BParFNmyA2UX/zZ9z/+B95j3iAh
z7GZTlain4pdXMUlfr2lE7tsaMYFy8dBXCiKIwdqN44jo0g/I2KXWDfiEGCoab9y
l3CwW603+8D/Q+2PGaWEftGy9j2YZqwjQLhaxO6Ty1HVYuOFz6gUXVeZSQUjNhFK
n2hoYpYj9QLTZqAVKFhI7ia7Ip6ozIFEuzWBoCah6f4NxiE75jtmPvcbAntEBkme
2ouwARAnRyVnl9gTk7RfUrnMLmurzHjgwDooqG+XeXznkvB7MVZjbO2gJPKwdaVe
UCF4lwg0Ki7nOYTxB501DmaUtCLwqBxxcbWhe5NffRjLrG5UcMJ4F80Yl+Lkjinq
9fLpCe8FCZAWuRsAAQrqK9UNOo0IyzteAPoJgRfza2bq3mfyziv0NIEjdiNUhTeP
5KV6ygM3s/G8A7vunPI33Tk1Iosbf5eAPneWEm+E8hqPXN4dsf4hOU7BniOKOqQI
dF+4Fi+kyW8B+5fV398RSHQCWTbVTIR0oLGySuHZ9mh1K/JVKrb3RciHgeYO78zE
FhwWlS5mFun95dUlHm1MUFPZm/+BytnbEUAiEmGyfRPHCKRCjSgFbpQWASY9f2ua
djU8sOa3+Oh9jubRGrTAzdi6E6KdiKdrnig6jNDcS/jjV8oml763oaC+Ljxfcdb7
kcGJ6MPexB8Jh9GqNI64Su+uZ0l7gMgztwCCPAUYXx/l7OTeo12fhDEC0DOQAfia
q+NnB6fk+2vfae0qunvq47de8QZkln+hg81ptNUkDiyljKWzJrXZG2KhTcfbTQap
gncMNIK5FYe3rxK7493rU4Ssg3v143ZjnkIoSwN8pPnKc/p/0bOEddO83cXUuPq3
ol4avcUzON1ZyHSsda+LdLkGaam66LLu5oskdYqMRW7Ci6Sj4m518sO3c8t4+hRl
ipa29P3qkZ45y0I4vxh2RrKTc2PHR7RtwY+Mr80G3KWEk+6Jf7oVtmZz6S4Yuwdm
vm78e2hgdVdnvfGEO1Nc+kIVgiUjad2UN67z46FzDp2C+U4HARZF9H2gigx+NtP0
gy/80CHDCPfonssYBbP03kQrf+Gjcouta4TpHlT0UQ4la2gTQogMbyzGY2QOBkDb
5DZMf11vnLnXItaDMAg6wo3gnKI/rGha5usvQ5iDEaN0na+eq+TL2TlyAxHA4679
yKC41lE0cezlMLWXmglv5YyiYAI1Pz5JBfDCLg8HosTiVJvLGHc92gSaxLUorCgs
7AuFCTpbB9/RuIflG1B1KQBu3+abT/gvrJ/iHndccx49h+JaWYyeyBK9AgfqCuYx
7oEv3d/ZZnP2bteQo+f09gt/nCXN8SM5/BQkjHu1ca44mKvZr9m3itlY422Mdpg1
vulyZhNTdKR9hv1IKrnu4vxsFlGtcw2WmCkt9daRJebnfiYZkJZeqcHzQlDqHIZA
IoCJjmdWa89GLopba/FhiefaddPVVIVg444XROZc7fM4DK/Ge8GN0fJMmLeEWsfZ
UL8T2HBWzLzzoUWEc1kJJSSJnYtj+kNL9Zr8BEZdhKSZBi0u5U5Q+jFhUwy5MTaW
PWm5kDyFB9lnBN2qrXqG3CtkNj1Ortl5gnSu7XDsB8ONLl5jRXtCaDEI5389GhP7
o2AA894BAMHdPMKiE5R2324ill3WkHKV0jd9C8xWMGpD2nKZhxIhwNPs0lzD4K3T
cImlLld+WckUIgXsyNcYy1VpPM6JcKsWMoLeqE+qx/dW/BJRUp/980gDyq0XXcLP
sSLVEGoxbZDZ1yXkOvD38HHwXgfA0LWnXGq2N860C0bRNNk83MK0Rn1Q+qG2srGY
UxNYGohhNUXI/l+OxqXwPECk9Eh60FKLU/Yi1Vc0o2OfioU5O5pk1O96rbhrmLsC
QB03sqcT4WHJDaPw8bhFgJRt39jDLd7bu7m5ivrdIweM08YGCFP1sfBjeasSR1TZ
bWKj7/Ykro5pQ1JtI5WYFfC/n9Z+M7EFtaM6LiQ8E+sjUlluPu9bd7qIOgYWKdcJ
2g2NjCOZLC+n79XKUMvxL/x5TQ0LPe+aSL/NTZc4/J7VQxK8jNWlmcE5DbGAOxHh
pMPdG7vrQlUnLAtn0bBYZvSi5vl19mHitH2iB4Fj60SNtaf8g4P+n5F4tA9QiNn2
BH4HfjhiwDR7rOS9HvtAN1uQwD1E31eOGPVEHebRyTTzxPlLTVr/evvBExoAutej
WIrZUMJdv2jwui42+JjNgrfIrS2P0w6gqsgQlswSd7bS5Zi9vR/IlSdPhzs5gD7S
i0mIlsFm/ZzVaxrDXFkX82iaL6Vg59izFzA7hCWfzUY6At4KSuCy8OO8AKclEVG1
PPeFxcrvJbcYsl8vCpBP9y/Z4gEqRQEPGqdSd6pq3EewnooQWoFEQeBeFkgo9jKT
8ZEM1RMUqUr9qJC37K9yr/jKfCwEofrHFG1eZ5SJdEBXQguGeLEN6ltrmVC95Ilx
/iv1XYs07pr/rNRknY8ptmXtz3hMJWl9cBy+ubqWvBnfHEbw2kFFXtoQ7AUEGYiH
Z7x8fy6ZS0+zQJCvfStdPgvG2MOJKBOe0KIAEdhxoZjHGPa3pj7uFAH6RAjWDaYy
YD6ode1y0blCC59qL5ROGVCctnyT6zjHZrKtPK/ieXV0xjtg0Qyya62ulWEtcTHN
a0npwNQ5XEPvG/EFRQMO84Gk1TLuZzxfGC+bsydck0nipOS3WJCEILelaj2ntMJN
liLrrVqNJgLdfcDHe6YtZzaRxQdRI/OEPxkX1RV5jatyQDG9KKe44tbb1RrYBWSt
8Irx8ebnTF5Od/a9LPK38skp2vTlu2AzEOkns8h4BLRVnSUTaK7gJ9nTVuEyppR2
Ourbc1szLZFGTJttnRrUKxw9zC07RqAfR8IdGh3QkhtvYpvEyZsRA1tCg5qVV7nN
XLiAkxKRPBENZ4R2BifV5efOVvfyl/rAqfXoo9oKQXqgg4GMfG4nUVsmMOegOcG4
UMzOh5IXdow0UKf+ZbF3UFDlBWO0xcBeMLGGeXcikBj9kTbdC1wb55uMFhIPrDTe
n4m95isJcIYoEV2m+JGuJ8dkbr7XVeau9/oqc5BVAxjREuijPJaD3EHRelBI9oI1
5kIdFe7960Nj847uVoR8Fh+NecKi0o0FoP9/ibkOe561JtEt1IwOFzmRftlh7Gpp
LeHzZF+dv/ImaLipShyFc/ofrXbG9CHAOFLSlBgiCo60bl3A/MrJoxV6VPL5CFhK
VaJW21SLMoy4JQe4VxCdY/v/dkT+0u//1MmdBLOwRJqNavyY6xl+liRuRIz/d2j/
zAp0Exbksb5ZDxwjK0Hv3YLEed+jW9Kdp4z84m+cEVw13zuF+zvhExP6sG3GUA/P
MIL+ZhQkWUgEKZHK7x4jxttjSymTsnQNxYiYY9pOUIamu74i20PMEteUZEnT1uEd
ja9ZtFI2CAj8P83UxsPCOHsWr1Z4lTmQZKcnxwDBkEVmc6agu5Jqd+Pk2xo8LJ5o
vccf3ncJWKDxMsqUXbiWOYHXhNFuQo6blsxRv8J5j2obxQFWY5yNLOUzXAbX05+k
xVovGJPMr4ajYYlpEAJjhtXTuJF7hpP8c0pb0GgLSMsxkZpVqEB/Agpjy7O2NCeM
6mIRAtUsnq8kZnR+fGXRBr1icjNx1Ldz/lelGC69yC8KEGlnKUbm0E5M0nju+oIU
MaweZ9tS6zbCM33youqwh4iFDEvjky3cJHWrho3cd7PjHm0Oi53ZFfwpypqqxA8Z
hCIzEKsVrn/VtTBsRbw38u+bLQ9LiI+mBcvOw29quxTmWT35cqWa9VIX+aKJnMp4
JJo3gheMyzGwYsfDsSyrMz6EMcHQDEN4k9IkD78CigDb4dT1a+DKbSvmMl54kl2T
et4SEo2sH8Sf5iP7dsQr5vIfCOT4w/lHxmFbC8gmPxEvb/oEj2I+s8WK4C/SRG0x
RVE3QqG6uMj+3bFhwa0Psr1qXWctmiqFQ0+O2xi34n4ebK4PzVeUlz0N1fo54qk2
mEccMlf/b2OR6spzvh3K/adOkPsaTlA4+DkSeUFS22Vgp5/ydZ7vZBzu+MW4p5FT
HGotbnnNMlrLkGnBSiO8SW5QQAu2EdNmt5II9/x+B+aJT5rd8+pkbbIcNQDrXav+
+xwssvhGaQ+EZ1fzrLLQwN/rt8S+I2SHMrTaAJJS79oI9AZiExnVtEq/SE2fmNMb
7YzqRAgp6nfoIwjfQ9+eMil7Bpfr7Kn7Ctjltz3jFDNMJAYYi0AA+uZuv5Lhv/7q
JBg/V/YpwYIIkc6n3QyQks2QcPGUKiA9xsxD9iud9vGl3GJGHxDmce4ZYKTRv6SS
D4X7kpyCGRUsyhsH9IVamVgIIVVegtxGVq3hZbnknhpRO/4q6oqpzoCckZdIl2wl
gj3ZgRoeS8eUv4r2W42twCHpLqpiRh8elF6eKCfMMt3eoG4syawTBcr0hSk5okNb
VW4KCL1jOr3ns9mZ9++ZczKws72ctmXY5Y+kyyuPMGtz07LN4PUQ+R96bAjwiySQ
nLeA9Ru+q6WlzK0oQYEZlUZ6nheIRukfd0BQaikViDvgBDIsFRsNty3+dWJy+eJh
ByYbPDk9kCShRrDNkCF36DdEGViIwJrtpJy8FyeR4V7JYvcZxFrpdIuQ6a7lj0Zi
+or+WdBNH1hb7pmN0eS027JOvBFcxg+8/LsfUrMjaVPxBOCEdmYWoOyzRgKteui2
cfT1M8QCZl0N1SP+CJSvG8uzdZS9OTlmv7atssC2l+IfuokxvjBAe7ahbl26c13y
NM8rxgAH+8lnj8ayId8fdxrX67fNjuSMEokkbUdURdYhf/EgrKZ/YtO8D+Mij6Ns
GvWZ7OuT1pExxrdQMSMsO1dYYWKJuX8NwYF9RwtGtgs5YILk76itAqNHZh1w4eT6
uXYetynYI4x04G35+ifIF3eH/PqQ98seucc7RDlKnYqsYKpGjyyPMcfbFdnY3dEf
3vPTWjgeQ5WQktZLtmVUBM6FgLKdhr0aX1A8YrENO1lLGCZJmx9HUCIV5noeVp42
Rz7dR8KoGHkmi707/wy+HqrE54ZzgWgqR/OV+ETBNu9DYBgdoBiw3hv8NUxm2SdS
YL0bcd7SIvL8yVy7yYlglrJiGMeAODjVFEeetghLWywMqGtG3S5g+0mK2U9nkw3n
+7tL75fiDD2VBG7bhghc12YWTAp2rJ1Z51MP900ORcw11/QLbCm5my8lwtNtZlA5
73iSQIgtb2Pey050mt49IbhIQsInNp+Vw4H8q9FG/bMuOXs288uh2jChOOo0zFcW
Lc+cgxD3ogCWsd7QMzmeCU5jDwK8f1CtAiD0KMEMbZuzj6eixtIYH4gWClqbHxON
CHlsSxjClSnWfJb+BnBdsusQB0jLgHmWo2X0BLRZN4ggY95eGdBwD3yMyG7ft6bH
zGohMH+RLzuy0LQUXgzvRFDKzlDYDqbtbxbZe0nhJnAWg1fuI+jkYm2cDHEusvVm
fvOHaIiYdmbAhHLeMPBiuWBkssLIvR5uwDsz1KteU+sfxizoQOMNS2umiNSkE2eh
OsMKJ93yqjkpKLiUcgs8jK46ftZ5bn+wGsxZYMqQ4QgiD+WSC82HbV+abtFYxU39
i9Z+LwC3ZtgMQqNWWt3iqiwxQcSgYaihFo+7M2qjjkNOmuWl+zqkNUIDHyf7/yM+
Jh0CB4dyR/Si9gG8DQjfiA30WFQto1Q9K76HTghvAbamsu1LB4yZVWe7wXKlgRLY
9kurupF9KLBMKvJNZ7jjs00Ee995X9Cx0SFlF4JTLSM9u/1MQ4auvSRBlYz0JyvS
nCT2XWCCvd1zuax/2qm0YjGn7AieU3M150cDFfRfxn/0WAxHC/4KJjKG9tV3m3Ph
mDLF5KIp/H3FUXHxyGc3fFus66kYigbqGENX8hab9HT8MKYGX/jLZVcOfqM9UNmK
5K3U7KcfUL/WH/eXfnrjtY6JQonaHZeXhTzbLmxfL3St7CA06UYNy5MYcXBpBZIn
YTzPXy0F+aPTb4MZ2ws006SCMzayWhmo6O7u3smjxpFqVTKDlsS3h/6Bnj7uOBWl
tbDceUp3IVTs0hNnKZJurruXomyimEcjgZ1SIMRCleWIZTe0jwzHB7yRuN3pxw92
FKVS27M2YW9NB33ggUPzg9OitEB8dElCzLLRB6KwcM1Fk02IhCrF3zduIfMU4XQV
s87V1dTytz+tAYVbWwppIJ2m5SImS5Y4TC8Gxe0O7uYOQmwaJJC6ImiJjHmqX/RA
j3soQrAEUQSdGP1NpBF40/Sexj+HL2xVeUgnUq+EwHNAE1PpwxlRsRocSE821z9a
JOLJVVSinqLcodkr0Op74K/hdPmwKqZy/TqJikKrcq8UA4I1l4thEKMQcSMu96W1
bQfxSg2zx8slHrNfzfgCVyF4VjhuqPgOGSiovbFScsxac1vx1bKNQbT8Owhto8O2
2JH6YjVQYuMNF7go531tCxGxMtyIgog9xZvmaM/Kqr3N4Q4qdlhNO5M7HkOQSYar
XSWdNvx4oHXxNVJiBtTaDfSyPUTxVnxn6vMUU6pw5v91Bp9WWA56x0aoDg44fpVf
nos38kencZa0Af6a5BfLmSwYC1GLMZzziceSBpko71y62np/4wcWtLnEImcvLc5F
CRPCUMatDnzVMNgZECt8IOxtLhQ8up3tX1lachYS3vYW4zuzJQDsx/EKTF3Vr/SH
RNEIuELkHqnNg0geXsbLes7Swsp2nz6xa8j9n0iH9oGE2cQhXH2kswL68rQOf5zX
si51lXuLYf1LwwuRajm+ZQMKM0xcUlK9Nmqnu95VemPGIZdLA28MZiE0K3eC12g6
R6jMV/sMTDUsPxOjXC1vM+kr7Al8sXxRCd3iVqP1vou0qsi6e1ooI/gD0aYAcGUG
9TjhheU/NWDcHVmCGNksmDjfiIVLEMp9XhqKtEMudoFs0d51Eat/V5H1cYsryKLZ
7QZwtIlVP65hvTWMTccfWsK13WvCPf6TdweHp9Djwt65T8hTjx0veFBSq7SqXpaV
oNLw0xHuAxIqBMPz5Br8JQAkjYyavckgnzsBLNI2HfEi2NcMFJ9fbGnhSWvX2PDs
qcZMIt50HYe9wdJoTrYKdUWRAkal1Lvn12ycCnfoa3F+6NaS94kdJc6QBLxyt8O2
1/ql9EnAnhuJ21TrMwwsTNx6xu/SEvadbc5JM4dRpKa5BlftCdjw9CAkBQ1rEEfA
+RtpUnVZHtEIeQzT+MBBjNp6fn0KnbS8rP8Pvo3PaHRPSKhV/z5C16D4pcSbX6eH
CPqCHiehn6Tj2VrZMaCPz6AxKjqmz78cjQWEJC76ORrN6aUcRmFf93hWGCFL9M0z
FWl19XDPyV/V/4MKmxOqxxMVBKr3zZM/ehKYrURc7Fode9hFKXkoymJCWF+S4p+j
G8tzvoAYrkjhxeg3rieBngvFn+sVQVzPYvjxklSbL5+bXKsFHDzyesuQbVeZ/rih
qfXX9W1lug7MoMgIQGadcasa1vDRx7CebcnBAJQhCwlhwt2Js14kJq9HvGWKZNIP
nI1+lR+g6b1bwGSfZw4oYPTpTj02ULUdtuDbFH0oFNKXNub/tz0qClPnFzuRndMy
THiUXWadQtzzskHGQS5eEF000D3QdOfdbLSagH4pVfZ1kjzVPx2vDwe9H2je8N54
cYA9GgdCBUPlvTMXu8HDcxGPBUq/ncAVMkSSQaHR6gszpB048KXiNAHxfL3OC6KA
yIglejYPqFirP13brYrmCUTniVEmWK+lgzz1nZRaWYzzMc7ynP28ouWleBabSmn9
3Wd5Gq9c4VSO30rYB2jP9FREr/mJXZiylxln4qcHxfcGcVRMrbtlD8rkhKdqtWaq
yxj9F74UFlDSGpF2iGWE93f20NfkT56KxEwPGRhuLsb4YP+F5Ph1BZPnpbzZud4x
Eq3hrM+7RG63UtDD/lWKH8OMVUFa2DAgbvxFvkJqnPLLAscwMA133vdbg9ImINSv
fxtcUQAVHx/Oj0jhgZUvz6bOoLtl6lOABQ58yXM7s+Fu5tie0kUFSYKMHwZRTEMc
1YKiVJAGhvHpLgceLYbdSDt7a5BsEfCMay4pnGtiuCJaYV1kYJtAMBIYvs3++NvM
ZA8pY8a4mEcoEW1B1jacMPCENnwfu52O7zcxKC9E/wmQnTpljD4XrpdQyM90Ynx2
/W7q4CGJNW4sIY5VuaYaVygJE3NOG9Lb8R6q4ei2shG55lB9uCxv9ibni9g6ARkO
2h6OZE6pvi8Cyu3PGHxi6XF5KRRHJolUNYQnUqBrbGVKC3n3psaz9K1Cl7yPuUv3
0fx6qRKtJcXnXJWv+o2GaLkkHgjfwZ69b6Dr3C9wWXvoCpZd7dVftSNbfZCBI3av
zjDWERlTY7Rn+TfJdDjjMJhBosHAi5bWp9VcENPF1MN+rRn1mTTA0omuIoAT/AME
vsUafh+QdS/nUU5exJ0Ey8CLIKLKhd7WS98BwR6/K8iro8VEdWvNpMRx2w72sEE0
84wfBncJ4Oad14gz18jcjuq48fsZF7tGvtdi4BiZ1MJ4VX0m9cTthN0numGeMPZd
xtJ2q9npbHnhRzr4WxiZ1nXHm6AyUHKCd2yIpD8hhilSJdRwpneo5/Q+z9V5zk2c
r2l7PZRC7waYX5c0jMLM5fFuF2dxF+UJGejKKkkarLi9X1W10zGavNKY2xUzyM4i
C8Cej5GNtBOLCOpIbMKeKUzlRkaAl8sfQPPV5x1yo1TYp8jPZzZU2UsNk0TtsUW3
3XYGYxgbi0MgGP/82BttbCQyLi20AQD1On+fUq7f12GVoHkUFuXqwyY/E6TICTyU
6+2TWR+LzpqI8+Cl6cC/b03xMxMWrtTJ5vSSmm8HsR9HVkh3xoTIrmuY+sXxBHam
eNMdmHdxypYOY5B6LoHdSJm/3nASNdhhrEzDiBDfSmIZQKM+F0uBak3GicUTpKzW
V4gENjLLLgvdXZK1sT3KKzrhB4OGCfSLEgDlEQO51V+k4jtZYuruXFlGyLTOezip
oVOSKGa5GkTkNICxGYr4PVKelRClvrRFxgSLXa6ZPnvo7b4SvbIKoyFb7G+IEKhx
k7LwU4xyD6GEFTqr1sUutaJSYaTNqobVZBa6YTxVHIZFvBseSQuCqoWoz6zkOWvh
8brDgBHJnEfugLeBt5uJbKV4+KPuQNTRYxzccRiwpEQ+h7SfScZfqj72xeInEx/A
84HB6rIHh+xlz6b5+v9MNWTHZgyr1rOsykYyZ6mVjSrQ/QnhTa+ok8CT5Xwt+G27
RL89YkKuTVnrdr+MISlZr5QMP1UxZueuESPWtSdxXf6chvLeIamvcCm1B3lDaVhl
C9um1gbFOsqkrNeQSchYst7xe2ZdQbn5XKS0f0hpbXAXGa2+UgVHIFL4wF0tIZNn
VW1hU7VYALAHpggcRMJYck1eeg+H5+uGzIYwM/RawRG4B8WuQYqZKynAy05we++P
wuiGWf10BOl8QfqbRW+UOO4HxdhAU4OcFJh/rB/Cw3gPAjueGYZ/hNuiOnQ8TPeA
SB7+lpeOGLHtVlgruTO7xHTEKKINSaH6Mgfkq77KX/rVRsykBhoKFYjpAzLqcgmG
HPO0KVP2lvIZejwixItZqvnSJE+hEmVR/wXTeB3Sr0VJ7DZ+RyMsaaOBRPVWjP/J
t4cllJvFxjk+vmb0VIp1SPGBuVwy1BpOnT7CmyDBeLFOLngpd5JZpdPBdiCG7apq
fSFlyr2n0meFuCi38gMnd8OkROMnxQ8EDS9M3EH4Q6hlexzFdLDNbG/TojrKZiBn
TO3zaa769kYeAO3bBuACDf72IRr1+KpENlkVoyIMIX/eNKKkGFp+nLsKMNxbTdDf
XPIwfYyGizR7qnVOZDmVEy9jjwLr8ttrvemf1AEw9Ltf/EVQ4GMYIewsKo9M2ldd
EhBxF1YI0OwRssTLH9SF60DGwCURfI0xxQAEGDpGK+SysAj8Sv8KXCzBcPF2bWdy
JfPdNqJZq+tV4j6XsALeDhX7SerKTzhYfBeRPUwwmfWGFom+TtADkSbKS1JOyp4c
7fzQg8Ff1qQ9Q8WaFdP+BRRR2Oe9uzD34D92TcxHMw9fXARcxQZxQwvK52cs7ArK
4Tij13ulCkr3eqekZY2Lb3IVOreeI4iolFYljIsTRBPmemEH95mfp7DCSsSJvp+3
6C/aSfEuk4KK0jchg/5/ElotoFTITr/euz+U2D/MXNFASyDSOBewB6g7H7EOjX2o
qpqOxHtJ4ztq+M/qMc6sHWustJsJfEoNf5nONAlVoeTtIWGgITWE3fzYdgO3GqQg
SfkTbmJZD9YzxDaGNbpSYULGNdV6FWNSD3sywD4SHOVYwCY0Mq5GnNqEVUvk98UY
jwlpqiYQHJ/bZR2iCQ4ApGvUItfZAqc87FXs8x7FmHGoeOBWmBzbWOnJpBBUcxZz
ON5USpxzjX4ODCABB4SfCvwkGB1gLElpANOpkil7qirR4sNN3QmaLydpSUcPLeKg
lBLtm5/6F/kPub2FC46qxCX9pJVGyN/LR8XtlIbGz6SN1Mcz4EtJPNsBLmp6y5L4
yYcOW9t4F1PdsxteISs7yNWBoiJuccgEPsrg0CcKNzGv2CahDvwiVKfOoJH0V7C4
ZkZcXGwrQT4CsPCiYODmBrpaDiRxh2/KcpDyU0zUsCvJlnKztdlxRIQI2c2mpv/a
7R8oyJdEOuMqih75ZxmAGBf8oDnijQBpENlGDboHLQOQQ6dLmO74Duktg1vwCVXy
k3WylO9Zyis7uSU4D43wHmaeMLqSah90buT5ZVPbpm5fobqxr+OCoC6RF04RHcVu
HzCoCIy6UR5AHhz7npBCH6ShP7HTGo7BuQ1SlsTAtqcaVb2rtrJ39hEet8YrPNC7
VeaG874XMSuhg0AbElE+iPz8lDc3Zz/DHOqbfDdD6d+zh3G/mvv/ZXbVm0sUTLwg
D6QLJa7HLQ9iuN+H1alKbV0R6IX2lr0+O3l7Rbm2swxHh41HSbNFwXkJotgk1aDj
hXgT9cjtSJay91ukXe7r/5UmC2+g2B7gXOUxqG67r8azsokjBWl23wjEwValjPuD
+zLnRxK9AZo39R2ZdMJW6ydtMKSz+PZj6Lobu5s3bE2Dk/M4QW5hkK994gpPl7Ua
pk94C2ipQJvYwBjh6yXeDogVTaI9+9YkZ1GC2GhwE8zLCxp4wWZJCLjaysojZyE/
v3J75F6EfZcOdJ5e3ZCLArdsmsfVEspeG7Gezt6SP8vhkSt118eb9V6piEL4Ccsx
04szfNX0RK5nsaGf3dm7rvWvnUNmIdaNilyCOnN+2QokJy8IWjl2r6VQYuNm8bX6
+bmqL3tdI9YNRda4pmokYRkD3Tdf6B4bCE2x+GMRBVEDad5tErETyYvB2WTpgIv0
71Z6dT3nW/N3vFVyOZsFlsIsQZb16F48RCJ0u9JMz7eHN3aDAkS5klbk1bDH8Y7h
BXrLC7xjD5Vur74j1bZCIGYt/FTu9S8ICVmMlMUOt+147SWApAljiasBlJ02UH2W
MhE0OcTC/ydEXgu4IZD92yNNi2il64wn4JWYySfESix1elbwPvsDzIdHk4zZMIrm
bPM962CJ1VspfRLJc0HAyz7HEi5EInO+/kYIAJa+OXtc4vH7HlRwYFX+OFK9fiVn
KAYQpZI0Wz6jmEYYLkaK/KUmhynRHlpc5Mps+63tFWKhRh3Pk0w510kU0bOK01kY
mB90J9+BmcMF/X+w1UX5M0LMiIFK3MJlqG0eMqWJhCGbzWyqbVF+STw8z7fjIPEn
fA5B0lVcjUkKnTRnwvjYv45l4WdyR2IqaiGg4lAvXG10rz7JO8kikVWNI+tC1ran
K4UlKwoU6Ljdfq8Qv4RVuehtv/Ntq8zgyIYWoxynN3oQU+F/BI+4n4+0Udb8cj18
MNx606InbWal2hFvJreJSxgGmZivzvj2AS/mtEBthMhWhKhpZtLJbNh9bOdfScEI
WOZn5HnpgbSg/2/F3vXwJFTrrHvMFTl6WQJIuZGYGBc+hNuXQ2sRo8ObXf4si1tR
soPQcJedkTDaoN6u7Y/dE4QzPl9+QvKzb6BP3+80QbHHUwMtUjsICLfpkLFBALRz
uIh5InM+YedYlGuVSBB2zmYdcrEOI6wT47tFkFCPSHhDUd8YE+2uGQw4jVz0ixzs
eGbvvgdTJargM097i1g+QyNuYM1NKrPCtmcGz3D9Azup8zOGXBiLR4Rx1GQjJpvi
yKFpgrQJYln18LuKyOI3/m8eBudgiGaJKVkjDmh6RfV+g9fScSvcbxp5ZjPVX8V8
re4MgkC4SWggNlCZGgzicKR97xno55Obao4qEqUcIaw8Hh+pVa7bH0yofDo/oeWW
TKmwXNEFvcTVTwWcIDMnSc5BM5V2E8JkaTiOLCfSfI4UvR5w7hsCMvu+THtEAAdh
PCTV/YOipvs3ksE4UHosNcmoLr7PPKXqSzr5ScAWC2CzDqBtzK//oKoodNoniWYC
pyoKtEGieLbzeP6Cc+aN+vN9+iBxutt05mZ4vV1Ef63SACZ9DvahxINkTRRyPqqd
2AW8F47HLs9GBhghbXJrbXWlfoE/gDrBIM5Me9r8XmRSgnpDPfVF3Psk8rqEyJJ5
uJME+804QGvJwxPnERYgAjqwdRueL1efaMqVbvEBQNUeoKrakWXgOFlBjnXu1Kxh
q7neIC/+DARKaL2gjzVfWtwugAviykZNAja/gElRIGBMWlxJVJRW0wfRIRPj2zRp
/oVg/zdnseJPI5ePNNnfd1LEZpCQzsQ1xlfCLcnT17mG9YaRoalGclAtPDCtaGCK
PxR3oq2d2q91RNK2CLEuUU6vTIk9z4kzOe+gg5QuMSBsns24X7OGeJm2iHXs1Yh3
8yvJl+ndR9VqaYtrTQ503zXkVr3mMqpkUYPiwoVxxmwyJM2bDvhj0j8kTUAeRbYn
/ic7o3ngifTIKyV6OB0Usfha+TfDkzG1xZeSA4S4z4IJIDO49r+o+A8CiUcVRAto
53/FprQbTjmUveGiv6IEjXLvo2QfWFRq5Cj4e86pnwLHndUPERMSIbBzNHB2LWQK
uBOVAuEG/k3uo9Rp0yGCd/2GJ4H5TmcGoH/IucoFJ7D/akDzXJIjKTygEsBJvoXT
37VSCeGcFUDnI5zAuH+U3g3VeOLlL4RMdKArSKmbLic41SyZpcG9NFUf4iretv4h
/izAE8jBV2AhCjYg6kqP6y88cWqWKlKGlOqyg+6HYNR21hbxK1sWsSXLEJWpQzKR
r0+StQZQmGbyhQFUl8T5Wq+f3KD/lOa7+89OAwyklmh5tiQm0+Y+EpSEBhPE07v/
H3ruY5bW7UkIdGQyR6JNkFofxmh4cTD/MRkx0WgLzmxcDYu8tD4cLooa31aUeK86
G4Blal8JturnIaNdmwwOHkIPWAJryX4oVqyzKP5PVEqPwsHsf26l8K4/8Mk9KjFr
JQ2q1rZKiah8FV4jfMNTQKL4mbeUwKB7e9uVGGkz7TzZs71jSjbNKN6843uAVVmG
JQS/++zeWc049fggXtW3xcULY1VeAjCyq20J/T1kpG1UsJHrsUJA7O61HPv0VMak
XZHvm+f/UOczAol3Ddp3PGAgn1YfiQmGAweckr6FGPra79W2IKdMWhLe69rsX0T2
myYkkn2UCthx/JownB6zuNasbRaVk85LvW37XkTCgJ2i/4HG1dFje4p5lACf0HGw
nwcLrYpoE2wBPYCtcwlCEDdByjidh8VYpB28q5Sz9Bv/nG63QzeZyoOoosAoIGZY
5/MBge0A4pyvAyDEf4j6kfmqO45tL3/g18NcNUl0YO5cOF1W2cK+aVJJDUOzgnlC
e8pmPSwNpjwOzzLkxATJvZ4wEJOvO/CDVCsnq/Dh0nVfbpwvYG2janwiBjp6RfGG
t7k7y6pqBDMaJ5MiCKjUkZqNABm9CV3g4wqKVzznKmFUWcIdHYAHHjGXV3WPOxYT
ZL157NAC8wPpNADOBQQTS15M8DhGzf9BGiwK6PPw4xp+Ia8RRbzefb5kLtnxHe63
OZ6ynp9vtFSYATb+wBLqsjeUHd0E+2bRvWqqonTzRXcV9mpUNU0e3bJ5ZVe/kzmM
u/rJrC/9rPsKDqLyyihuQSCOLjE2/fu1bNGNdM1XotKjPTUbIHz3xo2NWbI6V9dh
ZrGXc6xuECdm1M5pt5XFX1PEroUzyt8c0Ls+EZ1F7X+5E4/dvNGykhqP3MD+BAaq
T0qUWh1NINhAm9XD31uhJCBgEKpz4/iCjqZOBpwDbU9GBN/nD5xkGWpttxFm2YRU
DsbxR1ChMj8WH9eXHJH/Qhs6w5ruyjuVoeuWN06jMkVvLOleyFgd+bHNrfRvpHVr
N89hj+363rP8MqT3v3yYKIWaidV4d8qn4h3n+1PYoQKcl+3BHv8D+t4AyWugdEMa
4rqGOWaNATeU7eeKfD8fTbb/vsjN2lRhRKvsX+UsRbhgixFuSxQTZdSjfESkCR2r
uWhp4guuzEwIQWl7ovOm/C6hDvHSCsD0wGqwHNHoAZfmy7OAeLTBYxOWuxXxNVfU
djpvfFyML6pI823zVWohZf0Q7czCqMSzswDou2zLaQ5lLyGfGLzAp07VWyBon3uj
WeoKH5cvg4ZFvXBydt8n9gg4Z+DuAnkqGqrn/UyfNbpb3927qTSmlyBe6C+2JgYb
pWjW754w9hF50mLJCXh4c4Heq8c3KE4bu9ZpRm4r5g8BAq9YiDGrK8qKsk8Ja8qT
VxtssZvYh49QJKTlbjQ3LPYKeqm3I8qsx3drxsy3xkBE80UMy/BaDAMkq8MRkwZF
cpdRADrYouz+MCd+zUCPk2OfdpFkCT9RifUTAh9e8aPINoJUnPlr1TsP6bYew5Y2
teAcI9NJS/nPtVu8pnizlQD6iNluP75akfPIbv+qQ2wLACDNz9n05WOHrpkd7Uz+
M/kdj+YqEJ1msa3fTlHpYrfQAJazVPBMU2+Tkxw1dj3EqI5qkfWhnfwWZMTJcX6F
wRA+h1HfGs4nujEN17n/KJf+QrJL6P6iMLjubym8OL8yX1CK/CqP2lWZjixGxw0t
OfrPsVifHo//piGrjBqwuHU8jpApalNz3Tg7psZdHLAA+k6YRrdH2oU9z2PC1hny
VfEqOn2kwXr2cR9pGEtF9laWyJYdN0O+H2LMPdVKbMXMt/Kmb0rapBd+kzySyElN
11JZIojEn8A+F+D3nruAGVzEjg9T3SNaem1nHCreONm3sJnsQCN+2iay4G5jIgEk
+b2JV3Z2Zl5jDXx43f5GCN6dfy0HLHbe98NsNbILLpnAkQfubvHwQuo/SpjeXRTw
xY+uhT0QKYkAbmp3J2D8av3AN8oH+ZADuLgsraFefouKTdeRaN3tVFdtN9r9bB3o
EIs17ZwJFMIzF0EdJ1ov6JYFjRnqnqsaeeOC2URAAr/2+s8AV/63bJE9TOnEEQyt
b22dw33BQbFeFZL8YXvSZXu/rvV4AdJ7/LQRJ3xQUQW2GTJDKdLi+S7ZZSbk8k9w
SOSAAJAgyUQMcdpirM9pwtc9642gUOB40QlZnMYipHPN76jZIXrouvReJ8W2tGif
ntS3TvAK2UTTgftAi4ITWnITDCWqzZDQeMQArmqKxBB0/ViQY+JCkdC6D1v1n54F
Pycg2NsHR6asUe9RDLgfMaKabpSI8l2IjDV/3g/sXyhQdG+0VEP8mA5EG0sIDKLO
bQucyNFlUyzNb3bOE1qj2dPlI0k2s3OIxIyhv+Qvv83Ac2MNEg18+AUEWPNIYAMM
wrGzrn+CUKShkS0KTP8XhWJFncTX90k6n9xDR/NADnxJPJetsl/QvzG01c5FuGE2
YVoqoEl3FZJqGHDs5KQJaNPs14QY7+okK28a3zAKbGysCaU6s495R4XMI+utAsLA
P/LjcmekTaEo0/2Rm+141VoQmmRJwHwcQH6hy+EEiFj0SVAfaPvAB7JM7b+Vebf4
rKpMktPYoaXJdfJJ19UdpyyHWHWmqzotdJzjq2GWy6r8ol4ulpjwCk9G5Hi5mZ4E
F9/6Kdlsg6/R+Dua5jE4fFENxobEHE+/OOxzx2ydQ1NM/UkiBTl1tkcTBFK7lMMm
1rHHk7fyFI74809F+XJwyPClVNIfXRukg+sJVlkgzZIYvAXXrFLgFn7WlDkB6YN7
trvoRr8y3W1XYkUN3rTz0YJrAZ9gJg96Y0TFQsu7DJPSUgqY2N4EDDAO7PuwKwTu
KCkMET15VVvR2SCmcglT9kmrV/FhM0iUiIDmhfSrIkhnXsoj/RD1B1Kq7AUVoOwd
e3zi2XEJ/yZpuMaxXxr3lGBP192r0BuD/ryu3O5hH7VoDPfa0bYIl1+INCS7lmRM
AIZ7mWuKQPb8pgxurOvi5t3/9cbLGr3B9Id9+5tVAIQrBKTr9wx6t3QhTF3MbJVR
BMzeb3Ti7O9QTl15+vF8gbm0X1q7nA3OPdkoxJSYJgdFzkZlAU1N0eSXQS9QCAjl
VMVir1tL/Ff+1KY1GvFxPCaAJyePREn5rn3mrWqxmK3+98qowCWdyMq+QwXYhBrX
5tei+8iFmvlPpr51dVfFWx23KP8MfI98EFylN7d+2k4ZGkbRUKuVFlH3kfLGtbFp
QNlo76a8qCDpsZHATfV7RbgQ8obMFkgbe4EvTRtwX0Bkpbiepiywhale/fr4qLnT
BJoZ+1YjYnomX+8/qpvIuNX/wJrB4nMRLjc7s8wauOW9+cCAORG1ix1mve/h4rRG
glnhpExdZkb/ZPetC/JOcmdNQUWsskiaV/cdmGi2FlkKlDWAA7hfHcGCILe5Ol5N
1yiZHNrev1bt6QkadJkBnjS0gFGewFypt3uLsE9Ur2fqsOU6fX+SeJVKd8+MWp4e
7Tjqypxub2A4ctd3+KHaUvqw1Ku+4pXb6kDEuQJ9iOqS1r0TiaRMu6wrtHpc8AuM
jfTMVkKF9bgAvjXuAJpEaUgezi8+Epc1i6Q3VOUlrwX1p/ND5nwYo1BtF6cuzYzf
Ydv9WUasZqICCRzLnYNydXdV8A9lrhtKD7QJn38FYAsjMEkx7NMHqWVb+SetYO5W
zzCSnos0IRcOf5KmpLI81u9WjgkWzzu3aybI7TB/mIBR/q7d/gs7VkcX3iPlryb8
2IlIMsyRPbSAq6BzlB7PgnVtZZTSAMNaNgC2rBVSCb0NrPfn8drFVKCpA4U0QFtI
hfKCjsu3+0EADxv52MzAktjUkQDOycoJwR64orTNqFx4GeypbjsRwpb38TXlgIlP
RBSrtffm7W7qcpkzxv6VSsH141ZW4svLuqGXwOW/1yC+tyOrNd1rAFHGar9mYdAb
UJdbl1om+3/l1Y71QZz0Cwes6hHQswqyFlnR38zjQaJXxW8Mon/ikdWpW8lqD9vI
BSLd0bAd/JyQu8ldrUGRKfABkFzzxBwe3TQuRMeiCBeCO+8YJ+13S3HKdPDsy26t
NY6RKIygo+eOfJ6EoEjzqXFBTpFShvi+pVmdsY6fFtSbPb7Lk+gxQKjtBIQ96bGK
BZisO59ICR0tmNPuc82kCON9HzxeF4D3zxnsCOIKLkGzfhh22om5lW2+l4gp13i4
mih7inEyWt7xEzBXsLDJMMfZy3Hsts4BPANw6Dh52zk3xxKIrh7FJZJ0a2iRvCj4
jAxR8wO/vBNxQXKKs6/AtcicakWLQp88KV12K/2GxlyVdHSZR8yl4M1BClVW7Ap8
rMfJTjhKxMSQVNeM551vTlvFGqQfeU71esMEwRE0yVoK1UA/G99AuFWujpk/iDaa
VOxwKgnYqb0io02R5YRe1tnGyyocaLHRPQyXe7CizZ0TxA3NTqduKSTZ2u/vTMoO
lZ//R5YaJ5c8W0qbDWtFQTtM4EAemHZlTuCmAKkAUW16cKJz+wZu6XxevCCrqkfS
+oCR9xLDxGTvN5xzjodMis7lD5kfqY/xF6rmQELpHJ6K7TPJEhPRbP3pz9pzSoFS
KjaAPWbRfQqkqQzE04VS9BBP+PHIRfsaL04woObYuE05KeDdODRCziZepFyZiRUV
H3S3jXc5jBW62OJtph6kdNqF0Et2CB8gBQNv+vj2wRLH/XpGmxqYMPJom9gW9/Ed
Nc1cbsgrwbr54qmaal3Pv1dEwx2y+esRWr2w+qodtWHU1rqXVx8Ufm4+znjYx8gT
2/4/WB/L9YUJQTuOlHRPGh/p6GsXLlEln7gwQc2KW8Rl8iXmuvy59aFfTPVF+MNS
fw2gIHC7y+qtyvTBFo4HhFo0eEj+bvGAzZsyGs+L/PkuG8Le5wM/m0EWV4TuZJps
GnkDOny4RHGE9Jw/8pOm3/Wv5hgNX2feh+xQyidOXKI3YpOlSXYFPiR3HwSby0LT
Tgin1hAbO16nxqOjVqTlTNYKyBz/vJvv3rPxFW7OQEg1S1Hn+PVCVweSdxGINb7f
qIf8iSWYVQjaFByF1DuyVBHHPxCH/VubYeFrc0TCfG+VX9nv9+tkwh9NwOWGpVXa
7WU5ldm/GTJNJCuZGWDt241byXX15prbYkEczyeN76fMuv1Rbqb0ChV6fr5pYRBt
hhDD+WH8WqHH0wdiAxY6/YP/xzQla29I2zWx29pEUI+kNYQcUZWZu2GasP428WTw
zU7a07IcyJeuUJhqdLClaYjlHdyfB/uDEta3cE0rxbE2FvmJfau5wKmLWLt3WYwz
TczEIrDIvQkFXDZ7RGMmaZW99An4MjmuWLXGkYWjmleWrRZ68BN2WICQOG026IHD
JgR8IUy0OjH2jCKSTMlMbrCTjisARevAWwoBLKQkzETLvxeO9hbe4zir9mHv7JBd
6+eaH4iR+cjholNsx5P6pVrhB3F6MtwhH5BxnOPG7yObatHYuG9w35woAoXhbf3n
xucNRtaNx3IkzskoewvU7ugTznTuejfkHnFKMVJAUYYZEFWa/NVazkTEZZs8Qzku
m83IwfGsXUhuI1N6y7goQ7zqbanOykpz2PEkINvUZ19ukisbGBCqYmXt5uIO+JbI
nB3X7zLP1EwA6FjZJ6jds/Pl7pEq9J5bQTfFfiSgtpxfEraurjrVjinbItJ6rdlg
lCqNrFGgodV88CycHAA7A7237qt4fo59u0DxK60wlU5a9QqsVrI9DYGWeGc3h7R6
WgK9lGTSxHh+DfanJzCPEGmeEERL3DfmwAJh2zgO5B0En89Y2WQxMo78g74Gwyb2
Su7+Y4pHPSNOQ6lawcNpJsZh99hlDMAUozcTyW/vQ/U4mEySvCD0r7JrFINnzYBE
zcy7IHs41IV93bTj8WRb9YgY3m/OMv6BZjyXF3QTFCsMhnZO3wXERKTIuL78wJM/
RyXJtUH01IryPb/qSnu5cLmKdUpKJ3CDFYF83ShzIS1ZzyDC1sADqvhDDBsmwNko
6CiTdTsUAVhdlWLuHKaEkUwvqPl2kSzR6Lfp2sbk2FlM1wGgZ+8TDkG+mRKn7CsK
VTYnG6GS2foRdQfajk5u2XTJw/KJ9mySMoCAGUR+MYaj2ehMH3VvyOMonTp91g9Y
SRNfT0NLyIWf5G/VjPgf4hqlWEYkQrkBQ/HWCG27rQL0e7PbH13uD2Yv4ukvKQUf
v+H+ARbJJ1a+pzS09OFy1oP0JWQH4cZxqi7rHGJpxV2VV+DhYtkWs/j/msSsIxuv
8xI5FVYnj00Q/wwdgyFp+KqIAvP0xC28K8RU09fr1RSYj1hbYtiIlXt6BML2XNot
iCfLpmp3wElhWad/9JwbvNVAsSjpY1Pw97vwb/sx3ho1Unsw2MPiQFeAY6JOdixe
OrvyFYwecDOsH8r7pcRjVNP+bnM3fWPgMnFcO18EbzoeRqhEiFRJ7rhskBksbtGi
LzugG2vugXHyds3ZuqkK5t4wImYFXlzHxbRzErWVZbcp8Hus+MJXewFDRNCBYEC1
EYw55yUOKTP7+ZvZVZIXEn3XsK6nMY9fUA9GP8rTWcPmDT7XSHQPzSwqynusMp7I
S7jF3mSeQ0ystyZqUCZsU2secIZXzwkGvApsiWr3OXw7+ynsXleYnqjwrEAowO8x
96wHsTUdUqaFyWJAJLGEgda/8IJBHx9mZczKBvd49xIWlomBNAfI689sht+xdM9c
MiLKYwWhDGygiRdolgqKlPhKezXIRfuN7qIAMdIPEFhuMzm8rA7L/1RKY9F7vCvO
xqp3w6RJTztOsvs1XL72cJiryoWcbQ3Fzo6wV/7/J866qFbVp8hlupwDGrQBA0M3
tQrjVAhWk7gooQ+4iJ18PqJKQWN+ZfOo8gfC0nhMM6JUJX3e7EWkgfFeutDVtf33
5EFHFVxCQLTXn5j6dQ9h0S7+ZqmM450WYXsB7VZR3m5IRGzNJMbMN1G/1H+YtVQZ
pK7AoDuN2N+rLP3AyaTLxOgRk62y9M4sg++WCmnv9nWJUoG3X6rBn/ewy/yBcdE6
e/pHrkCxZRA2nLOA1U/sO6vNG8H6zYea+5Yy0Rcb4Um97T/oW6TCpqTn7hcelbY+
nggMUR9LmjRlSvB4oAk1jz5fFUJo8kxj5RIi3K+Ii4ymO37wWQKwFbX1DlKfXvqL
yStR5JyeuQoXDssIrI7n7H3N4DbBQkJSncPX67wtwc6u+mQr8JrsW7U1CFyJcfWZ
LBVXsdl9TXnApRy7J+wagjCyYS44Jrp8A7/fb0x25yI5MH/zHkP7ohMkZlwho/Vx
6bq6rgap1Gp1grwwe+nAUNwgB/PPcTr09S45mEQcktZ34r5oswwqyaHFe42q4GwN
9K4pZUwXZ1J/f0hMLsqLrRZhbTeHw70Zo84IEk0Vyx+B/R4f2t2zL2fBKfHZQmhU
qvud0rg8jq4pmcSixQtGtUupresBqIoa/OW6rJhhRsLdHUiCjZk0PQUZ1Pkg11Tp
qO4ZIWSlOPHHFJRlbV9PmDSgdyKlCgDoYqNXpXk5KhdKntTwt4ap+b4ch0WnXYse
yRCW8kiSFW1RkBFsyqGuYWY7lSG9Ld1vqGxH5dkRuHV9PqN38R8o6r2iD76kue2i
i26j1cZ0gFf4L18Bin/WTk36AvAhaiVjvrsh563mteUXbThvW2P1vEWj2vXx4Mvt
iNby2ZSu5XLGJvpDIqSkzBcZmSs6i+9FaF2McVYgm5UPjI2GcxlrSyzk42hb6bUK
sdQygrsdTFrVvm4KnZFeA3jFqtwVCH+E44iIknRK/xtsKwtTCa0AM5SfuWclFWMI
xKFzLfKVmKZ2idCRFOM4C5cxM6+f6DRnt8MHma1J5Q3AgZL+OF+xz+bOaer2wIa1
0RYRTOvCCMyg7pyZlpDjmJtqgMmvW6ivD08rL2AFN88FrZguidKwwdVq07qd/CsQ
WwGMOx6IfApUVBbWJrf65PodOjZnYfE0QqWMdFcZyAcJVDpdDUoOm95Y/m+CqVxx
4wqx4YeVYqtrL7Hg2sdjE4HNy7X3EYh57e8rdL18fRDu8TxBOYmk9XhOkdpNPlqP
eP12y3aDDgVZ105Htg1UIUA5VO7DZBXpwHBN7BUSM5kRfgu4/AApIQxYBK1jIMs5
El9eLM3pH1LsmbVDq7eVyk03t3+IivxPX+fxaaLRc3v8S7ye+2TegGVmCNp6YDs/
uW0w2BK5M86LyRuTmAqDfBTKntLlLfpk+meMqHX769CtU1yLh9dK1orqiWykVpCc
zTmKGTBWCthoIo6cuemy8axyLSZQL5+h0KrNnMHrkEW7N59xUXJFyPq1SPVW0VW1
ni4c+53UnoQjNsgZvG17kJHvzZRAFMNQsuSsERPsWlaZkOVGl0sdWWDrarWD4R3d
ckRoArA0fKsMAfe/tmFJoplp2KIk7X9/b+2vv1/GYfIWTtPYiUDLArN0jULsmBWP
Yv6pRVoNUl2ej1a23rIWOx67dd7bryBNB+gCpiMDEtjB42iUXCrqP7soVB2OIhSC
L41bldiMCi9QUhAmLSEKa+DplA4Xlehbg21PutBcRENKDDWll1J3OgDew09T9iPc
VkSvjb37/QTsl6YmWJlxtAka7MKn/Qaz1UUfCV8X+15Ok6fEv2I3CaXo7CM64wM/
YM/1M0gpGD/r5YHBWBwGRsso11FdCpyuwjI0hTyz2i1aqXyguHsrN/VhK1VgCYV5
sQNIKyJE8n0UFT+xhInKs5OglNnGCFx/XrZbj8SyUS2K9NXjnW2m6U9TJ3xAbDes
dEdplKxUaD1EG9BWUZcgyP8p8iPU/D7grBlkRzfbZFetNoRd/qTmFXxSq0X8/p6R
/ZOf5XR3QpcC/4scmnLJdy+SHELOCk1B9vC/8E9FnV6SpjhaQlfn3tukhSbw6bhs
8GDxb4RZA9vvCY/taD0AmrWAvWPAp1rvh6DiaFKVJPAmpK4zMpeLwJJuHnZu1Twj
rlvu/Rwtzte3dhpKRSq1o6WexzHia7SCBqBwevyomXdGEO+stkvSZQz/5ucZ9DX4
+itHbdgFnXBj9UmqrcvzD7EnwoEnP3LrroijGuQdEIwdfIo9vAfuzravkYi9Iagd
liuTpdGxcObh96amst4kPqnAEyEcN8movERTl0TTfzP35uLRC+X1TwQyRE9tndV7
X1pdneMSYdXosR1OVL0wXmqBl2seKb+6bMvQthuDsqv6MkztwYCEzWwBm4YQzs1w
jt7LvCGfkZGLBB/TtpFGT3aCDb39WJRS1zSumsZ85+TCYfcJmKLEeAQ97HrLspTK
Oc5Q+dNylre2uE0jWGR0T9Vgs0TX+AZFzawMOad0jFjTMWr6AVqKDtDSuxcXlVSW
qQQsGyHE9vCeYwyYmHjBtr1B37QnmfRsiQyGY+cPjnvKGwUVP7NoNFNhwEG32yXK
9+12etpv26ve38Dt7c0yd72Tdg8yFj5AZz/DQkRIlt1pyvaQughPSrPo02sht/7d
61Xltis85SGUga7krIyBR3Bu97kEbjntKiHkTolJkTnwVfMZ/uJcUN8XDU6VTNfD
Dz0bP5Up/rz3C8nK4n6I7voqNbgL5M94CRrl5q38Oqy9X0NyWsNzKeoQZnIQgwLo
NKF09gTS/L1xuasuPD+1S+m5C6sc7lXZP4cde1I6DU8f7dNTlYyBucL3uQSyv0Cs
L8Y7rSLAnqvK6l938EF5swIi5m5fzS88UT7TJ0pfmYSMc/9qQiXsemQ+a555SuZa
iLGICJtwXVAqDR7bCevtkHuXic4bb0MBnT3p1iZ4bplpLCCNy6MlpMBTL5qmem6q
k6TKLaqUIHyiOokD4bjTkeLzdN86LikhQf4Zoqxg03AnaVZkiuPuLlRmpUJrlB7+
5qaut1DXy3KTEpbbzHpIe12YSdl3u6A9WAaxM8qDtqdgNQmFgBKAWkPZhXn39kKj
nGiHgjCnggdJoSae2vwiZd6cRYlZY1b3JJLWfAfUtxBWzG7k49lZRRSqvidgGimN
tSG+8rNBejELBTxD6/QJprcUjA0Cy6mAbuS6psg2GXKS6CJWZ9G9UEqzr1VFD3PV
EYU8YGmB+XKDZpKobA8Bo0ec+cnB4k3pqdHDwFK+wMuAoijKnvARZWBqrwum7UnX
uBYLMxp7i8nl3NZsySzVsiqkRycx1zilVElVTHyjNN7JfE1XCirg0wfo6CAnZ9FS
kcpAgLtICjgssJfHrmnVXmUsCgWSF1OFSMntNyWN3wIe6MJvr6lyzjnoNyDAt8sK
NLV0WODPvkY2YdPheAGAHpjBtBgwH+xBXRkhV4zJ2hIyOrmzOLiIiZ/Fcw+GzOlM
sgRgZX+3Ff5K2F7KQMl/eY1hD41q/BTz//R095iJQpZRT6WJ7r5MiapGtYEA9vjT
4Ij34xy86qRKeatmIHrZskycDjnb6jEGTrWKYfaH18cSXGhD84kRX/Jm5sFTX+eh
dk6YiRIQ0ptwMIKu2BvyRx0hV8nF0fzXg3lvypOTsXHgTQyCQ7HLFo0YwJ10pIcS
wBVEP8zcBhrIthgyckvpJfivQ0IvwO1jlFI0So/qBOI9ZkJyCSELoBlhTQlA+AAJ
Hf2QFVDv2+NsIrZEu6nHJqYZJIYXiFQemC0Rg/obOF7Sh+JpMJtmj3HIK6kklEPL
TNvu007W5aDgRT71/ZP8yb1phAFsbitMxltdXP8KvzZvzrKDj8XuNhc0S3gqCa90
BQFTqojmDJukcyTrDDBIGBhspZuYMfuenIiGyOGR/1IRjamvTuFca6RmOGqGI/MV
1w61OQfEMvRlcCEOmXOuze7F3jjNexsQqrkZw2s8DdUO3CawkeSOQ7NUUJHwyB/0
lr3rZ/D0O+qpxkLhOwV8hGkuXu/wcR0HNZozDBIhNBxiYBwY+ck7HyfJC/Pjjfmd
+0nwUFAk174u1mOE00R4WaYvvlHhXu219XzspkebVPJHUG4TcGaafQgdXegukLVx
4HLiE0rkd8l2PZyN2SE6ZRE2IQRc7e67syJD3OgfP05KNV6x4d873ByRlvXFml5R
vM9XXL2sz/n5ThoSymnyQu8sO6z2Y97RsivCuyPGR9Zg78F8yGnhoWngKskZsBqY
oqTnGS2czr8PbNrG9FFIuBkQqUCVdypX0ykEJ6nS0W9gyzgLFTvqx5zlvDaG4vN4
9DlkJnrybakcZrvtBXxJuli9yjx30x5/Y7eJBUKwqxxRTIzl0UUppJ0Onjy1I5X3
VWhfPRnVbNOZFIe8Q8OmXmGprs8GdRI2KJukk9+Fu1e/RrVufHHjwu55BtJLDhZr
4LlH950s7m/2nfH3coFl+oA6o+UpmjfgqGLS6wnqQXGEDgTyBFEYaXrzaxKSrZ06
3MymB5W8ukXSDJ8Qrp+Tc3cXcvmAaHXGT4ma4d5JswvOyjkkWiQFWLVQwO8VEWDZ
K2VQz0to4xLq/j2w12BAA9UDWv3rYwRT41jfmoSiSRVtUsAXbLmxORBPJw54IAr+
O/l1GKNjmMo0gexO7YIOBv7QC+iXx0Q6Rv2fB7ZLw6OrquCA5aptkzi4F/tUr+OM
/cHuBr8Fb68un2/K8T1dylKOIDKAyZNiQ8X6n89qkWjjeKn+1OHIxGKEHU/AoFBl
vgzlarwKvsd/A+Vlu5KzQJSDwVpOewkd+JUvvLviGc2yNSYHxOEHInPje5RH4OFj
d7oNkroUaXPTiwRErIm+v9m1/JmjwbGYw67EqjO4RbQqn3IY+8n2zfEyN/rxCA42
9NOdpBlEqXSLhIXwEGcwltv300QVvrJ94M2zaHBlA83s54i+zAIiooduCsw+CQlj
WLPott11dsadxX9lRKmyuyaqolnrbDLq2LlYuIQdq7WYC+WSW7gw5J0u9+5X5TM6
riv7xgPklOssJax03VJiR1joTx4bpoGYUhvpXkM4wdKshQhe74jlW1N+D5rab2Dx
m6e/aILa10hHKxMge1Ekpi4qRDlhprZ54JqoEmQ1eA7qiMzwwUK2gYxYNV2CF8eD
YK1QI/U8HpwH1AdTXpwPMrly40lbEYiKhjMnoqNXWI4JObIoub+24UVvysixVP7m
jV+EbeVO3nCDAybNMvBcVqVWIetzstBQGoLe0JfV4p77wALJ8SbF8hQV5azw3W35
xKy1xB9ZCDvW1reT/L2BDlcwCAJ9Y3ooqu3a6UEZP1m8L0xMj8VjBS/rJUJC/SY9
A6MCG3y39BMqJFMgsoqYjGa6QViP0AgX97l5hyJwcf4pytJkoVqgXjO7gCQ2MXFC
hGrY6dRwg/+2ioxSKEBdl3cYY/zvb3VkYyGqMIpcERxrtg1vykcJ5Jw9235KkVth
uo4oR9ChtMM7Es+UBl6JVWPulusctIvQe4J4hsxo5NHxaqKwXPVORNtHHUnYUUAR
WWUApp1Xpc/PhvDM/bpqt7hO3oSeZ4ywImyLEvDnh4pWfNeWGOohhMk86cTW1Y2h
5L9LwT74pRXZijjmXDaIlJ16rRxLT3+RfnGsWsR3FxwwJKMk2rYnobuTuUSvbsFA
sn1CcEZ2cnt0guVcBcPMRHCWAsga9YF5mz5CA7n1xR6+8tsvBurrv6QNBxA2uchs
x4r2k0jZ0L9hDwajM2Q2/gvpSCm0Nm0s/Rl6UccXPtREfMyRCbMaeU9+WbwDPhpH
Q12NQba4CrFhEBmaGVOqzsRKFr/3XyOtyKELNDe/5l68z1g232xyS6drMgbcM5eU
gBACEB0mhb2Lb2SyhcO8f4DRkJuVb41OjhlmVBQwnI7LFFDpMYs/DTgj2DZkFxy0
AXnF9qmpW6y0Tho7kPcwPlFnNeRHdVSxKoF7YD7dJ6+zzWuyKO744CUVNEzu4Cgo
k0nnwQ1QXuy8vqT7UbF56+wiHxrO78VM72RYi+QqNeVr1frbOAmcpaVTFop6QTfE
Lj7bhW1t4iPj9AopLyxwzeCwBJI2tPtjHFGJs4PDoYz3RaGcBNK6ZnlV1gvqlwHM
YQK23Y95OhfChJbr4SRI7va4ZzFJX0rCY55Ul5pp1fZQSnzIbXkk/tv4w715UQC9
a6wigiyTDjZykp+ftrTHKvZIb9anNeESSiZpXnVs6b8hJjx943DL6xoVMXeK5lW9
DffE6frkS8Y5konIiPLXxjcUcCCPxx+yZY3OlOeQX0Dj9jYoKI1bn1H+E87LZ1x5
gAZhje8y12BVjf9gxYiKKLKFORGDKC/OIJdCfBzysst1eCbZ9CaxFvoN5n2A88hp
cPi/xRqzZPI1DhdZX5nrwHUYeZkOBKaYUUid5vDIISU9UMMAcNpIOzj19nFZ94dZ
p7mQByMqTaAxNtMGrAhTzkvaF0i9ylnEjlY8drfkZjiMxIu9skQ7JhqYxHzO/24L
nfV/UQn/HZi4YGo6dbKgy/a40G63POjdQH0d4VACL1SKayZn2/W9nC7oD5w6y+rW
eZ1pXXXwqX6glzcn64e/balG0MCbG0h98OhABl4ju2Xs4NJxiccHCypnDB1SHinn
8Y1FWY8UYnc5FbUwY8EcRqklalKQGmE2kjfPLmT9jdldNS7S8ShQMcqTslZNCXov
+CrD9+u8wHC8TRRm/DENdFTeNZD5XT8976IHsSMZWp3V02Mn/3BjQFYyKQ4ff4u5
yaCQfNRhrWgpY3HiRt/sFGF+kh5OdRpIFHEHe67LMzddUmhO0Xbf/DfJuUBUAm0V
cms4ASAuAjdxcXhY3lj0rpWJNsVzHu7je67AvcuE3xFy8vy/eE2JX95UkuBkh7iv
N5KXynDXZYHcb3aAllAIRFvAku/ODk9OIw2POa+Sc5CJwH07CjEW5g4ai7MSnlV3
E1j+IB1wL/sdN+oV9Wa1ADjnLybt+EQy+jfh0t5cdAeSV4oukSPgN9+oy6l0ezpo
uhL9ZS0UvMoWz/rS9OIUYtbeJhvTH+9WSUlWZYRm4KIO6oHDTkd0pUZVOE1m9sBc
yHOkLZtUFbKgv8A0b77bsMa/jq9SjnSauMDIB070oWZqE96LL9hVeUR4GtQnpgQk
SBO1Gfc9nUkzfZVJg1yPFAI4AMALmo9/u0ZeY9aUWO9tcMyHENTSGo7zSevgXnGF
7FznD18kcNTQM8hmC6TW1/yu2blnx/Ml37LYyjqkwdCjvcA8qdL4oi1K/O7kTVyl
/l7EzNJit6uGp0CJitNkZWQ8ut0SCQnqjOojw+C1sraKuwQvteNp6bz9/SHWOr3p
4ekzFZBxxOpau3i+Kk/E30limQGSldTAOVzh7qlC0bAc4jts5AmExKMpZAam7myp
l+kNQkvlBFUg/kZkEFagZ1lQ2tnXQR6nrMe91Qo/BUsXvvrSMra3CwEEdzxGb6wI
X0v7aucaIQ3GOV7Er4ZjzN+eNqhLFwlfx9TvtUitVDJPcni9NmbKVLq4Poide8Cc
2u2XXPzl4Sk1Tjcfv3+3ZSUFabc3GLKV4AnKsycEF5YSH8fVRy2ZIQM6p0SPmmPs
3AjgwlGnXF5Ov6rpKL+a+qFqw/OOsyLnBWi1+lVncEV5kmwDP0BDPm66EOgMMwPD
AwoVrZQ3q4S9emRsW+I1jGrn7ckXsoOHIf3JevuKgOIyVvOVRNUAJjIEAUh4tqJ+
J0p9PjHFkSSFGPaxFtPWOhuogwlN0i+ABkK5nHfeDdHdsn0G4eMsJrwTAOzxAJf2
EWOZZvdHtQ6HICBTrKQa9DqiMcsK8gBDZGJhjeu+TsCJr5rm1+j42XiqN+eajAf0
Wr4wDSKl6Lzxfduc4YTw03rs8c/V0oEneFqfwtKU1B4lYyPdiQl/azQ8tbmlD89+
mk2ZMwsO/BCiJSJ92i1VYsuj8II6ien+x2uARqYbc5U9Hapr460GvAuqI8SkEuuI
DBU/et3OmmBVzgANKqX/2456x5Tk5iaOzL+8UH7el/aaWtla/6xR0PoyHV4OGSGG
UXTmeWmnFKJf7ufgWApcDuvhDFnb2J8ScGmFssyyhDKn0lFvuRGwe2+P8g+unehp
xuII9VD5RJC0eIIMWcDleZdS6QBsnJKdgQomWvRDYH0gvDzyGvwNYfOKKm8p6P4E
+miSkDZWM/zqK+JMtyrURlFAQG81LCc9KRv0RMiPtApkiTlqynhYnaiPHCqR+V4l
LiTg6/9C62HXOt4A0mEjV5yNiXqtaJyPi37YV3LEcWCMY2/Oya0ljrsY789Oh//P
S+wzRZ1wDwZfBYV4x8nuC+uN8uv+y0W8TRciOQSEF/TelGDxAzhST51aicfFguEN
ii8szqZ76Qh7MxqyskNPbL0CaZvLjROeJjeyYpupXu6ldGpXJsPUMoFyuWUJWeBJ
GXBcXt1VwE0k6tPcvHQF3skNouQDDf5+dYJ/IFcmJ9zjltGu6dSjG3+8q/8EXEj8
5HQ/2Xhdx1XGOyh/NXDI9RHystHv/mlE1Xyq/XLuvsOE3c6ugsADaHS8hCUOJOja
Ca8gLru8lqeataYSkHGLztq72FI7wqP7WXgcaP0mJTmM5BN4f7RA34UvHfc/QZpG
XZ0aWAgTAaiODJozoDjYAtQckjdzZKedlGh8ZfT1Zy4067hoQZ2cXyjcWa5It+1C
oMJ5TeJe4kyi2C9oVK5nyUJDGv7rhObZvkTg/r2Jrb5h8nIMd5mLm+WMdUw84xD4
lVXqWYnU/gBlAVeNNAcEfJrV4Zlz2LRuH67ru69120hCqZMp+0VL08LYvJDYMqMI
G5RBaz2SFdV9xYXfM9/GUN0YbCcumXFH/0mpCwwPQmd6Y1wvyC6xpOcHT7InrjO2
w2PiHafYqmf3c3nCNmD4XGVjUTVMOae4ika+ULwpWmLVn7vG+d+Z+lLY4OvmxYFf
0WEthEpZYOE3xSRJ1ftFjk2NM6qcKkNVPg8fIek0KYM9g4iu31SmudL0k1H6gs2S
MmsU6tz839233rkGaY26o/z2C+sA9NxdOv6aVacyYpBFj189kHYRrJ0w0fDpPxIA
v0Hs3sZf7mUGmwUYqpNfdNo2BnCCan80aH6s8RtTUORs9Kf7VlZu9/VZE86CszkS
BzzndtG36DIDAxYSWrRZOSGM7M7X+dLxwOvIhhISrys0+X3TlFiHIWSoR7A4Leev
HGhH6Genf1I0xky3BoBJlk3j5oGsjIDWiM5ZaFW8t40oi952yX2zjPdxYrqie2fU
vw4XXou9IUJGEmpxWuRdG3W960T81Q0gBRIXxhtrRgaRhkfUGMG3WIRQOWe2iK+h
MQvDep5vwsIxNSegiis3w6G3UWHrYXt90X0hpmv31VDNcyjQzkupL22midTp7Siq
KLDJMKxRAjTxDpDtyhEwOPVj3/FuG0NiBnaZMbAsao2YBl7eMpoJKKUljRpbZR1A
EoWZ5FEl8QIZyr2g3cqK3PaqunrQoYDw3W7ccDX1AG1M4v8Er0tkaicFUCZkRhY7
DWF+7dO5hsxTXTdTBHF0ethN+UbRQJNaNKV1WW5H/9ukWNGqHElb59PXZErPgFWi
oHuRDHwChMG6F7dOdI2N24HN1c2a2oBjnrCRqntWidWcOfyVmHHpHlwoZdulRtBS
LnG2B5mZTN/mUlYY2lqsFz/hl6Tzl7rZlCIyhBrKccBcuz0owIC9nnRuur9PoU0X
/NypT0nxXM7JOoGb9/vnraSI/C8TJhd9Id9oyBSU2Q6WClO/UJFk1AsBPsw/NbTY
+dFF9dDtA1a8HekZsfehjCTmsR6Lr7dfN7CUb6++q9MLnvSvn8xP5256P42jI/jK
ztz57hsz8UN+b4xIZeOp8e/+kjNI/QE8TuNI/EFKMPF55sXqnDq3oKi7WW1X1phv
KL6Yy4dzGaeCY1HkmIWMtUqXZv3X/F/us+jYZ5YZjW5AQqsm5iNk8a0o96myx7p1
Hjp3fY4CiwI/O9FWe43INDV59aorQ0WEqeBTNAz96oeQFJwF4Hu0vQh82ftLMpSg
nwTZ8wRn263KUil5EaWHJ2WxOG4dmzmWP+qTEPgjW85Q/EqRKjjIkFLWKm2+837X
cwrzs3XJGBCU6p4olxWr+vxaUgcAZb+Xo4/iu+VHcHWnmnSHnkVdck+DPvtqfMf/
xNTZIt1rJRIoNX7NEy52G9uZTOJVd22TzG7hS8Kp2cVZNUfdFrDd4uGjqxvZfoGV
zwWI1oeroRP8SKxOOUaWwk02pF3+8iC/Nbk7hSoo4bWFddTCLsuaEdW6VHua3CfU
vKGqiLDe/niZ+l9H1+UuBpQI6AtXM7CJo90HknN30Bq7EOva/denUqt5UxBV2c0v
/97rJN8NmofMU3jf58Pa4MuyrSvZb47TPsavnKOwUvQB0kbpFdje2zX5LM+r9+ZD
Q8mm+gbkLTTZXh7n/+wGuZJUnr0c+821+wy2zPOPhi13PAak67t6fsZEoUVPQyZV
jn2vReu3qJUZty6zTTAFzNYsdsasqCsqtDqjEKHx6lHftB3aUZG819MbuXIWAc4f
KWpHEd5KjP0Vf2nAGSs8EBAs5V/ICqoWCkgQ+lW55bJw2snaDJLFvKvZulnzYy3W
zq4sLvoQ9wfbWEOCRVqNPoqJAsL1EuaAqc9HgdIXSNVisGtojDdDtj0SRNbDlqMQ
bprxOSTi3DzADn1e6X7Q59D8VvsfocOX7wHouPbcXPDHFct8VBNlstzav6Q3FWod
e2XVKHBQfH3bJMeU5b6TavzIU23pdxlbONfTNmVv8HMH6ziWC6usSk8Mhpdc0Ff9
x7GC5bf9F8aSnrOxE5EKehY9Q4TNfoXf4IJFeNwrzA4dx0N/im40bY/7EtXs8fAN
GSmLzVeWZ/Q9wa1YaItk78ZmCZia2rYPTOXyoqBnU7kFBcVlICXMakScTPKryllj
Y/Pm/+YYtdFvTKOPUTW8iO/7F8Na9OI8rqNS3mV0laLoO5tM0FEiA+CrltpRtgN+
mG0Te4yqciPoT07PmlWF5DWBrxtk97xEG6a3iXNqJC9cee5UBN4QgFjUBOMSBfrs
m/XPdrxsbHN6m40NFTyVYOKG9dHjrjmGLUkcZq5G9qPjzXTpOSiOE2HgYgJbs2eP
rGLzrgAmtSMj24Q6nTpoSt5rOq+nOwtt1dt6NvJZdurxfF+9bvmiz/P+LAmRU9sB
SewBgHWt5h0XwglUsx/PkEguAMI9wZy+l7C8CARAsiAeSJMU3oZR6bvuwYVne1RC
VqvDlbxPlBDDL6StvpLBuDz2EJ0i6SarwgE3Vhgm5ajt+t9d4i2+6aCn+LfqX5+o
Q5rO7ftLbGxCeNvt44dcQ+LZzxSEZARn+6PL635zEZCWLBud6YXLpM0sOCw92TxQ
apQ0ymHdVchkrDWYVoGvJMAQigyLMqgHGoevJ4H22qF6PTEDTmGrqz0DdR/oyrDe
UZjc1OMCw3Z/hw4qOq1bKUzhr2PDtBSEsB6BQ/wNykOJ3eVsidvewJG6fmhkiqFj
t35uW0nbF+PDW80hW88yHMUju5xCAKiPKdU3wMJ8XR/N7ytA4PS8ORy+ya/nJ4uE
Yxe0PebTeYYab36yu7qqTHlr1zyKlh3paZaL9Myhjk1V3MnXnFI7BqAgtGFEz7tE
FYMjz8a5ZXYuNwJgTUkQFlM3ec83wkQFRUAST150TDV0TFqR13fAKe3VfJqKcn2f
ylJU0/u3BzOBu428+a+ay/k0vL75UULnYYnvttMw57V7YGxN5AXxjddLy7QNoE8Y
LKpXnTQi2iEYInLNp/BOX6BZHqxWnuIeTYJjwJ4rPahzRE1BVHAg68kJ4AISFqeg
5zFy/HXjKkDXOHtD/6yRdyJfDQo+FGxxiAUqDKJOG5xU63hlQSfBIEh+pWESrBNM
AyrINVh7FgKdTazIBxqFzdHYdUo9o/3mdfG7K+PyLyYCXFMWsQLycJG3CjhEO4rZ
5+rME9pCeiVVKtNDeq/Mp5Nv6fRR6P2bjI0xfUaleL2nxSywvM/GWoD9ZgWqAqSf
LGmABdznvlNFrzbYAheU4FNUeYymsqp8K5kliDHO9+r48Wac/vqGNzMvjFp6m7Av
mUBfJBC9ntkpe6/SF4rOyjyAdle7qwKUB/ulKSOzm4AFuBUFUNgDv/KvTB6Kz5WT
ROU6G4/9y7dmG2LKTi8RjP9VVxyT4H1f5G/wKqSvVykNRWhnLypzGmBpk5PMItF2
TNUUUmT+Kz5s0GuIL269hhGAjwBPMslSp2x9pEsZhZzTyGxfMUfiJz2Cjbvbquik
42/MojqyI/J1v1iXJJegXfzlgMlE/u8KzWX6+ZbHTORR4wGi/7synFuBCnZqmMjb
rVkof2/SO/fHoht8kVBYKx7YmNOtqLx2IkCGPl25XH1/+2QX3qQ1U2PtD77RKSgj
+WKpCGovH+rcqSu/LiFAPUV1KHmfJ3m/n38TAP69uTnNv+HeznDroU+DS8ZBR6bU
LfSy6O4EdT4tqwxRMoWRAlffTtUuAoOHzaAPJitxWoPWG9NcU9RToYy/cuOzjERT
6a1/tQxC/YmSwpCp2MiBYSiHOLh0JeQFC+hLweQ+4eXfCFIZ7PKjjwkXo9RWAKpr
tKOyuTOSCezdeQOcrHOqyRAHqfICbXk1mi7csFo4mpaANfAep2j0qQEMdCo4UK6K
/9RHd5snoxJG7gvCIye7LbPusFSNT7tVqTKA0F8tmwSijx9ryx+UKbZGyMJM5dTg
VgW51VAGqBaCLodMYAaFw8tgm07nlDPDEaBCWw58n2NC5lk+xxHog9ow+jtAAuxs
ZQBc741IoSgCGeB2rgjKXzyRrQeDWaAkX0tRUxmlnZa91IGfi6RQ6pqiyuFokDT9
bZCTrWGQRJLbZQsKVE2405s6uJcGdu9cJ8XO4YXxIGhoR2wyxHpbOIwDUNXHpZvx
vElPv9nuaYItxfXbF0x8u6vpuHYZIwAon1xktLIHMjmE5bKZ9crtg8BdvKrlCRbb
Jk684CAfmnGuz/E4XwzFPmK5gdmY3P8CcdkqaND9XLlC+deGprL3+5pGIEn3aRs+
YBgNp40HGU2MZ4vfxr9VIzJyfK6QZplGteUoy/OxHFdPREn5J6PiCCZTSUeWDbzY
MrLD1hDe7EtiqLfRr3QzxEbEE6ImBTt+itrPLP46ytzqEzP09K0g9/y5BvRqkI22
vQULOfMhxQGuL4Fggrk7+JJl+ZIKIwGa7w+gctD6kOfuJC6jJJI589gjBuIdzG+S
nMSiz6PGqlDz7LV8jBLakYbiyuK8SFV7TqVHKS88U36f4rutXRwUEQ7MECXgeex5
nHdRsaOdBaxxK4xB7zB3gih8+nIi9yFlJZz/6btwPYksyKIi/hXthDZlQmRYqzJN
OpEnjRS4vfje147dDiikYyFHiWb6uZa2MCexrE4yfuZlYdLwuI9zXzfRkFSQOFVD
xnsh+lv90ZtUdAX5wRw/QLUaM75eZ3Tp7ENTDSvRzS1GyzwiLucBPbWnVJK94//X
ytfSfTNshevn+mlpKXDBsjH/l+LEicaC0A8fFWZtLJ0UDK8xtf5wtcJKiwtbhBI/
POkSdjT9CpJhJdf0BuAD4qx69XVmAeJEerWpnF4r/Qvrbi82lTRMTCVTXAlOTlXN
HxdlbwNKgCos6AJgFynHRHLmb+Lc1lKpNgEn1qUllW97qePSRcHDxIZHSutAMDWx
xePYHpFqvmVFJOTOg1ibRreKuJH32qo9KSohUh48urooGm4NopH81EfRyoG7G6Dd
4sjal1YOuQV22lZau7JkMF1fQjTmq8di2IMnnTZ7JRgZ4G+7g66ZJt8OF9AN5RLy
faPEpdr5IFM/rAD3PqJMKhoNO0MAmlOL8SoXsGTYignbySGoab5BTfSnVw6Ssv9c
qOQhiCav8RtB+eoUVDVbJcFdtGjpy9sb1vsFaDc0bon9PBQzOq2SX/363rMwAcon
xuisRj2RPdjlX7/q9Q97YR2iwz+IWlN0o7vfPVPLgbdQ+bVDNLgKF1Kn9G9c6D+P
ePwv632krPpeW/wIfvt4J7BqGV0mJ8AKs7+UoDh1uZVmKoUoLC/Tw5EYqjGFSEvn
SRJpa7LfDPwCT3nnZyYz79ySUz9zUW/rW8/p6pYqeXcB9N5ygOBcxm+6x21PY8DO
wS1LwWjwcWBNbeTnaDmt7V2EqHjh/lzuyFMZadZZkAbpfyH3zqrfU8zZA7kBR4z/
cCDHH7ZOX4APE5VngTzLaUdn/l66I5f4rQiZNiMzT7VZQcBePOg9yHNHBM0QW2E5
/YsbHT9jHzA3rw+Ipa/1W/o85vUepYMlkoOWNrKTNp7T0nLUB2zTMc5HrEaasLdq
h+Jq32URQIbWPjS3wWop+yWtZKIeRqmmjP5F/bolduG2DplUmiDwRyYthxt6bLjW
xZKmbIg1iIiKzwt0XRY+oDJvPue4iq0O44PjVWz2YsLghJzuzrVW05pJp9CX6ZgK
GHhX8OgrkQmqgQSrQu6T/wYlOGNw9etrCxvocyT8wryPWqV9BjDx05mXTOtYD+bl
FTZ94/1JI0dwcu3kRfqZWRztCvO79YmMyfLV3ybK1TGzlbFcsedo3Xp0iQzkWYv3
50AN+jIBdAz22iCmbEBmz/4bVTTOWwk5IAVq65+fWsAZjRI9IC1F4ua81VaW8bUc
7Sb96toJmlkVhFpto1nZ/gLHez/qtEU1uIUjkLfK5qHhE4IRCdpcaEPeqwXA4s2D
4SxcyN1/pLp7mybF4J/k/7olK4eenFwCGe1e7KS9eLlc696TZtKFVG98zKx0fgSp
1ES1A2PqyE/wshwkPGXGz1qE/D0oXyq8QeoWfxfgCF98B+VNFPTgDtK0FFBRZsWA
2lT3XMc6R2vGzp90fQA8ndA/9PUDe13B3PDuipyMEDakueDFeQevKeRTpfxjvUnV
4D7PkJp6oMZmHErRXjwy+6veEvqHJo3EOaJhrKVpDFrtusLaFtU/kUhjO7BmkzTF
ANRbV73yuFlvFBGwp1Bo3pJh8nUSQvf/0zeVBLcxWATRleiYSHjcI9qYSgQbW6e3
KzNwvn/LEFnzrjn3r/ubU+hU7Bh5G8FEOmcL1GMVa3DgfIYbEHpTD2VgyAwDd3+m
l2Q346c7VAxR5V0S/fW1gT9rG0l4tRewFfa1hEhAVllcDDMwOBhaPL0pov7O3rAQ
2HhJbNjPwQQ30MJ4kuu6YcCdaHMFVe0A8PTj+8dG8P7WF6W9JsvOiSFyMh9+YoXS
sURWEZTdmOmvWCb0XncEfktAfQqhANJvh5QMA/2w715UPshVtI9IEJM/2Supa883
8sYLGPdnjmxo8nay1s3LB5fQR88CeL6fYjIC4H5V3OtRcrUUMUN+oEsdT5jEDpa0
u4wyBuNezFjLkvmTF6F0J1/vVovC7XpyqjUDGfQn1oSduHW46Cezv66/1w/ZhVPo
sWX3GxjwPrFXRMQ/WLWUiB4JxyCKgfyeCG4zzQQiNdVfuQdGVH2zQs+sHlXrt45N
0G4gpSUb0aALGTB3Q0Q/SYwnrP9SY8g0D8qxtLk3klIyiUdDC4alv7PxF4k6UgKK
GMYkeEqDic3gk57oB87Fet3jU7rwu3Z08S47eVXgh7bxiXhFQgRBby2oDbGLTjRz
s2xKW8yK9DrhR7ksze03puHOHM+2PzelNx3Yf2grQk7IKngoTJfTSxehqTcFC2XR
j2DnkI1DccudLcA/FkEToOZvJe4ueSxHEflCC0RIHv1iNTMgHEzn0NzFpQu7P69g
QGt5gZJTeQ4UO2pPFUr3IpyJs7Fa7DmBL7K1JTwcNeLtveuD7K9iZPmbKLF8q260
HG+wIQes+P4zuNl5eWCiZa6g2pVZZAp6EshBQvagt2CLnNMYcQlStiWemDJumlX8
YpWTQv+GGsLTay8ybN/ApeqIVaEql21xtXJtsGenldu1RfNQONKCT4XwTaTECUNt
dpkL7/VhgK0cQ2jpDZgdpcjAeIwd88oJF9u6L86bDuTeFgX4P5/KEaoJzAnFrLCx
pHkwjxaYvaLan32xw6xN9lYKYrwIXBuJSQCLGuIeJ3AZKbe/sY97k00qnVYOP5Gp
MO8QzY83SsZWrxQUakQ/9qXk30amGrPClsTM9SmI6pVwK1haV/0eIWiMxhQtZXrF
Qisoggrm74LszcAGPilpCzY28Cg9LkauMv64bJfDXWv5M8EI8KzpFnab5Q/+TW/n
6NC5Ga4zS9IvLTCvkQxy7wzUtm0i7CBbINBRlXVC9anwA89dsmCiinzG+JSPDM3i
jMyEv71OP8GVrDE0EIgeWjXtGH29bBRkk+c6JjzKijdaIe8Gh7A1FQ9adp01POwP
ophLuVrJg66EgB5y8ctr3/E9Pb07tM/keZEuFLhSPBD5Wo3ZQng34QMNwkDOGQoa
8SQ8rnXlIx6ZCwpgd7M6HZyoI7SCc9y3As+Mf9qUJaCunZMpS16p+irM9CcqdTCk
IL9TiW0/DWlBM9GeN34haOF5Q2gKO7ZRl/VPRxOprV2rz6MMZUrVrGdNKw1foZz9
GVz5DQaSD96hNuDIkqTdxxMwUnO3JN5OS6jXJbGvF/kTXzZoVr9hNuiUi74naIdI
DUHlD0cG/gsaOrqtHq8d0frE9dIjaoXTj8BRvhXvl1eYqqkBgXHYY8yGTEXJgG6I
LLhwhmq4TKg1UjALsSzUjm9/WTkYEalrntYqj4tpk35XXkUOr+W2FKklzEp/fk70
M6pCZ6DxpYIYHv1JR/gJl43rfB8tczlLwpDdOxQaS2DSCXqcdTfBCYlP7gFVC3gn
v6iAmDBkCV0ym98feUxnj4EnCStKwKX6t05on/t9lHwCb7LMR0hpg8CbZqQNiK2O
pKrBODPTOJMTcjTghLbxoweeJLhfb0OowZbMdF+JFL57F9IEHcmmg5KfGP/BX2Ak
I7+LRQpLAk77g0SuiAhtgCIRGBVNhx+UHFYwwM5fZkkOxkkuaO9VvuU7A0dj69sn
VaZNcA4XLrRk+wypZEioqP8vUh9phy1TGPP6DfIxKMgYTaxBLlZUP0XgjeKhyTKW
AwJzsLvlENGBtFzFCeoeDfr68owECv0Cggwu5ej0DdfgroiHjaPzd40D8zEdCJGa
6LVii3o71+6GSt1RZstDPsBnlZ/pR/QvEnXc0REAVnYSOsKOiJfIQRBr0vFSgoDM
/RriGSoIMlnE3qqW+OZ8oLd9uhDGht4JzrvvotGPeIRn9X74+FJVXa5FcPZW1Dnt
YPeyEgBadMFlMOeGbn1jG1EUsxLpCZKLOA3or4iKVncB3n9EQC3DOPMOJVYiPsgu
8BYtLdfDFjFLI2y+gqXZRmUfLnuqZHFpPfFSzzHA/xSz+6ZOHzXBGQ99JyYiKmkc
cp5MOZki/FNp3lHsbTkVDK/wDoxzsVmecZExONvcbZtFZMp6uLITgvJkjk40spc6
/Rvi0reyiKmyR8m/ZHXTbWt3oWJpRdH9inHJGwArK3DOquYtjxY5/2dkNxKB7Gvo
GjFOtUw/qM6K6AJ2pebiJy8hqU0XX4ChARIdJ4r8BcPNH+QKvGUxvnSE0MOSZoYE
5jP/w+IO8WIavgxkmgM554unIoV2XsltFS3/jFQKNPGDh2n96/eQQ8mUt21HWRAE
Ekxrup2VCrRckCQWgcLSzr0TbsyvAHx58LCj8n0nkwz02bs5gSMy9BcuxECABlgR
RStQnELfCQBiBpzJAu+sqdt7OGbFVZU3DIaYQk4eWRgapZ3iUwBa505i5EgSbVF8
xnFAw/u+tHqETaTULYIWJLMj2PN0XHy9BI4Aw84I5QcO6HB7HzunKAI7kjQxMKhK
X9LtvfvmumurATjmcrRsyzGtPCRUyNCOfIM7l4mAKGYjVjp9Tipw4Sx6xIkUABq1
l3Bx28Qze+ziwuAwa1I73qczXDwwdui9QY25y9jbQj3LWU+SMCv+x540dx2itZ0a
8HvHQruNPsDeEl8n76PdSpljJjsg+5RFB6Y/h1cxSCCWRl85AKqMciKHIdIlD3Kc
IhaYiydRBdZKQ7uHj+Tu15t6KlA1s9kyAPvBYAeAMLwnBEvshm3SwraiQdnS+axR
Psm1CWNpDOFayNaeZCuOkY4owAEgrXAR7LqNCkruPX/GM2vct7qUNCWDDUPpvJSt
hGnHFDVAWnl7+LwgB0WrhB6ykryumbuFKwJHYWmaC1E9Yp+bQZRmBK0Pw15QoAra
lrDtu2VZ4FFHKOyd2Cvv++a/FxgrNlQCXaLP+kYJJnYFly5TEEe1SVgYmLBaRPBi
A9G2Dv5OtnUfno4I1Kp1mSB8XMwmguUlnno2mQiQ7lnhKjRPf2RbKTfueewBMxii
BzZKSfrexuC3LWh76aOQZmtRHZj9ckwnHpfdCtfyqOLStMzbDqARKgIQfUGJL8Zk
vwP455snrmqf31GtHj9iMzFZOUdUiTFynsasYrQo2HV2WKWGpMWdXbyZtvh8ajII
3KEGMyFSPjLY0K2+BCwtzQKkoQeXdeVzaYMH2gUTCu0YMOurv6yWZm0/IlaKRuFt
+fiK23ngMIolBcWyGR/TBtoYG1ozqyLn9VPsuvdizgr4DBQoqoC9Buga3q0srv/k
WXyxKGhcp7ucbUA9WIkzJagWwGiI7T3Y4ahJKFzADcsQ0DZWKLd/V6uqfJtQBHYG
Sc2/r3JfGL/f66X3o36X26NiRlrnsUMV5rJqCkq2ZT6X1PSyrNGkU2HMTY2M7/XT
t9AyPcOtP434kqqb/v2Nz4uD1XXJ+BAlXh0bY1QAETihNrX3aH2Bs1H8dCAxX7zR
ZUrK/m+vnfiJkQQG7kt+FE187t+tIQcyKMxCk2WOipsWJglK8sGP42JgWanTlGVu
jyUECErjgoYRdYabnIWJJ7fwtbPLuyqWrx+CBlQ5zMxzuJEGf+ow5B4YFOdiLU4J
rLlFYlAWVIirt3lxC3rhw+pDNVJ2fbpASISdZI9T4j5bETwyhR+LfR2NKxdmeufr
Ttrs+BmbjBZrWiDP4AfCo25PT8j4jHoywIrcoBw7Oqol5cF22A+jI8s/qcIl3YL6
weZ2k7cyu7+oeTwoLgRRqTEIzHzFHzKuhDb0/NigZiTJLRz2HVcZDeovuLy9Cn+Q
kbOHmWLrIcxL/t9WAz3395TnmwupnPBDAA5teCD5+UEiF50fqX36uTLeMDcUw/pD
IQfA6ktBF7tkGQe6vMrrYHHRFqiEZTgJiWsVEBSN2n9xBM3QGlZPlPQ5K7+kcTXt
FnULlDgnaX3vOxSAKs25/Gp7UJDoWCWzaLJ0QZQpPVD7yVI87z6xEEmEw9MfBCPx
xAgUBgqIxo6SLujehSXHzoJ3bg9KB4KvMWcViscG0/nkzHZ7cfWSuQ033DdcVEG1
KX/FijVpOMHgVTWUEWZlDQtXIWhgdPShX1yOH8CFE1oW2RqDYblLhDyHiO5ycxh4
eiRlpIPSS00LpgY8uaDExDIBRnoOZlPbVrRUYPGCFH6S7+B1U0loU4yc4wJVOotP
e4KIyYEajN+qkeXoeUP5nQiEucpxOx6J3gSijFjWPGsqjGp4dgrbjlcYy0wLXxtE
Hts3IBLHOFwoe36By6zsbDTr28XGbz9lb0cYDEyjMjclZoNbLCy23gpeBy59PT3V
IYqSjHvwzZmZFULRHie8hld7CSvvnXzgWPhjZd0wtrZJTd2SzGAyb+lfXoMl4+om
Yt6V0xsiZZp2/brH6tcG8Ae1CkwPPuiiTSwbluja8zT5PAGPOxQR48aBHRH3aME5
FLQZ/SFve2bwai2OZV89xAoq9I2iS1C+QwStj0F9lNIz/A7FkY2+FsOaAF+dUT8Q
WU5OuNHYpg/mInDciRcskPLIlsvXGWTRUkM2Ga+wRzFXmTATPd3kkFBy0t1i3GQ+
kqHWVmGg/7lvCtnHA7JHJkG8Htg9S9hHT8C3GbvTuK7pNTcKykvfJoYVo6a8RKp5
lybVJbhotsKsG8Bzyt50ojOLMgNhWfxpMsakhAonxwousqiRTY66D9+hU5LqfeZu
3/FE20lUPdVVosAJBYqwJEBjC8tQ1C5/SLypZQ/S42a3oSj/aD7kvChBnZ0wqKlj
DmqMLdcihN4EpqyBEe1Ue3TXHY+ZVyqVHOPM1o3S/ThRz1SypzZT3WFHfzpUSUNE
SrzOroqSw/MRkv6KyDkN5ie8hsVPtdHsHSKmHpA56caRufmvASA9VFetzJfmLxK/
uTC0Evua6ndAHQQoItCLq+Nr0PEOex+N3l7p5OYUfK/OFbjyPCjVKux2LmGlOJSx
iXx3437dRJIII9rGsChENZ+gaLOosiIoIxxZWADCIYBq1/0EHOa93IwNORUpOjXT
nG6wGBaDZVjeir4rSJo0bYhNAops+tQb+2XYhFUMpwdsEvCNoeC1yxddv9nuZAqK
4hGhhyvXRzbioBDHgSPl8iAsFEV88ne1cmQoS1NcXPLD7PKmk1zbzrbwYhmLNQD/
MpL3NVbCfilTEBATfqEJO/oruGkiPGyWDVTLcHHsXZ97XXcek1595Mi7SiW4lgOj
mpey+B2yA8k2x+gj684fjPubz0XsDuY3DzMTdtCgGc+pKNTQ7JNi7j9k0zMOSAAS
USildMxNXlSsIyhyJHxHMHJs3SIy2yGj2fitkgO8UDSH9AW1Oygo0Ctu1XQnawfC
3exTiP0BBVuLdUCbinGsSkdNLbGZpn89wIyh47RGMIRd9vH39yM3aSxsD0sMPgWW
nMcASrbPvke/nkc2XSeJ+WqPBpn3TFYxXZNRbeFihn3PkJ+dnWjvo4cvJkt6Qkp4
pOBmDComZlzVNuEZEqsKRUWdGdi0m8wOKSbn1Rz1SXiIFymiBOjRWPFzyoNDHf3K
obaQvPLU2XG3wWLwdsiBU+sTVn5a6rmhb8cjEIObNHQSAqmBAyqZng6feoLuTLoW
Hrjl7erb4GClit3brf77Rp/X1UOOyP1xDdDUfj+nD5Fka6teWH9Vox+yzaz2ZS8t
xvtG+23U9j8DykcDLgIGGD/glSdt+kWB25LLy4F7fXbQnr9BATGhf0PdsF7b4hYK
pme6wGl4Xduxip9gphv4XNEHTi4RsGNsYdSbBm98d+mGN0zCP978jr6ORGllGfy3
0NVMYNH4QqYHuikhPy/7UGlw4hJJm+5TucfsMdiroQmjKEHkhTbgw1YotNQfufAg
SzJbA7dzSY9gZPEOwP2DR18LTpzf7c62oIVIDduB1nYj36/T1Oz5/JVRCrqoLWKF
kLlEUCoGEMAwV5UmHOgsmakjxnPfWYz10qZ1O+rrMo+e5QwCJinPJJN1uQQ9Tpn3
DdZr1eWhZ7eZz0qKxSJenbjFie4DkOj4mu/DyjzAunoJOkodmfhI5VjkJUtFH4s5
H6B8ik7Zko38OGfjfIcUhKO7X0K0Zb2VlkzijDfq2gxw5U5Sk1rAkwit15KTrPzg
Yowx7LhEvD+JbLektD15y3j9JCSM7+b5QxcmIlF2WVbAy9Qxkrxz9NY1wZKTTtzm
E3o2T9RWYMEHdvhVgzq2ogMglKFUsHMGCmHFrLfvmoGEfQmxCHfFDN90WI+jeVWK
LXFcCapuNCezsNTFxZcJ4SQU0PZjUx9FKIWW/d7AubuRQO/NIHG+45MVtPcN9A0Z
3iPdqGWD+PK8xPsY1OnFShUlh2jtUTi1+FwjEezWtCpmXg/mXrK9+4dQ8kv0CA6C
XV+npp8WHMoX8Q89uVG4nPI08xZmTzE1STN6V5wsh0+EiF55qKe4MSZgCRqz9MwR
xe8aZTaGY5fsvxGXhgOIUCOteH1GxVskThX4bD5kZKsRzegB56D92/achb4hGPml
AXBQ0bTfjgkkOtnlK+P+CWE32iJjy2eSc6p3GlAA6QWXWxsDXagzkDmjN3ybIUSJ
O1bDE687D+Yt9jKNNfoxMDusCVvZePdMYAb89aKWp2vb9oX9whwSRsTho69QM8By
XtO+fRj6H3mNflZoTkBQ++0BRmEC08a+RXFah+FjXppxCwtfDrCN7IsCS9ftDh+o
wScWZQl3WzFGB6oSx8UHmwekow24ieRhjCb79FfQqd3nknxXGPwWL4qyHZhnNEpJ
vrtkkaSznJBK4V4cpep/MOHkJ424K/RD/1o8iN4gpq3W/1z9zVffnmcA1IwxIcDI
MkGn0NTF/G37WwOILIDQO8yUgU9PArrLqPy95voXmzUGSH+72UcGrI6RTZTEOEhh
1bXbZ/HqP982jXIQX86QNmrvpjtc/j2gJAlY+RcfTsIXr0MUV2mFRW/Xg2bIbabj
uvvZl1MrtfPXbiYHzc6iyCExC40Px6s13jxnVbEegkC0xxDIn6ZYDyFMrD69X6SY
reDbEpe0hLkpWi2l7wpnd+DbmdNjEH0IQ4rimnmT2Yv6+jSvptClkH/mLXwLNexm
kXwQZGKMpV68hdJDO8xyJQEE2e8LRbnIDJO7JQpZjBxr8mMT+zK4qZEP967c4vnH
2QfTJNoK1bM+O0+i35+t31zLj7eQc4DDT2cTLZ7ombGomPe/gZHmFy897SbZJlHK
PLUbYik8ndnsUSe10kG70f9ibvCDA0O6UQPGQuu4YJP+5a8zMw9VbAnc2bGNQxmq
c84bt0NLoGuZEGDAKthRSL7EQCuiXTkPuF1eGRtqB8O6mXEgePnd5yqYVZH1aiUT
P39K+xAETXOpfkXGGM4Lo1YVOv4oyV/sotj9+DDA+SOGNRKoj6Jx77HKFbrUPRWa
1s3SVsbWUrNfgi9XwsNNyj6wGa0S9aXPH3Ml044enA/iKMCnvG8vngapH2fSdrGo
2Jp3WyMfICdNQOANyCJ9wGrZe1oW7pv1z4grZdtLzJ3QkmLgIJll+zwIyi2kKZ3J
+hKdf0B8pAFy2SD9GgWo9sxgGAHCPFDYeUmylXhBnGL8cugrbiiMiHZlRQE4b8uj
teVAjaw8/yWYKRMCkDW5HqKpW5IzHMYcZYb31Uw5isCfm4Vla/XTfxwFBSTBg7hi
2YPQ5nxz4QKaz6N2vPr6IX1xjeLCAUYYmLE3Ib78oF5N0YLA8A/nOjpiFYa6Ldln
hjFRVj18sV2bo4HS/lzdgCvaUVWLMfrvhuIGTN+JQ94CV0DMrZkklaRd1BqMSnCS
VgX0W2pMJvt0ctfOQn4mipsghlsafPR2wgva34h7LvOofTYaFqOF1OXuAHy9AJJ4
Dl9fbr2gVld9m9uPC5v8u8FfzFPTs51Qji+tnP30xeY/pqcc11LnuJ+g8ckaHYwx
hQHcY3oAgAagIUtZkQqrfn1tihs+AzSYdbUcmQTqXiR6Q3NuDmLcJglh5nZ4SG6E
4duUCNS4bMeed2+eK1FDKd++TOuVFq/VkEwjszFNSDHDUs6DCF7CgVG4O6MXqoTf
nAHuKuwGCtJFM96Ky0L8tPE17fAZs9bRd9WQf6v3icd9CFAdHK1z4GwfV03aayJR
a/HBQbhIiaocvrMTcB3kl2YcTzVdTyGud1wc3vnTvtGJLWZgXfbYT26PYLey8g3X
CdsJhuBUmfNkIv7becVFoVXt62BLTeqSWzh5ucncgyNmQTjzjAN2TWmGsmiNiylY
0imAA4u6yTEq5ej40fG8QIYBFOE7fdPeiMf7A/YCOBdSBKd+QElfw5gt6TBUdrhp
7GQqWU9+3YZpHFcrIvBoR6SG8+8vcQEDnrc9oIsyQqSPP1e2s3UIHaNtl570b0pQ
FNnKel77gVQhZgDcQzEgK18PhgvGaOeOKRt17HdJ0xd+jhq1yac3D6VPq3dplkpZ
RZC0RuL686Zvd7jvnYy7ch/MEUQMaAE7WbDWVSEG5yHfnIDPOn9ZHMXCyuyQYRMw
m7l2S9aEekxkNHhCifH1mqshWR6fVSJTdT0Hu0sDs73SOvYx0aOH0gnst0GgToO8
SFYPg9HOPpZFUfnqZTiCPnMQMrctGNvG3qL0OM2UKt+ulQiGRtcsmygKxTnOLllz
c6ga9CSFQZWlQxpgDBgOT9Lc+B4b22uc3X+GJ5YR9TrtuS3a0JTRKcqsYsGPqNJh
R7XMNaCl/jmu4KG3iOd98MgwJ/Rip1YbuTVQhR7URStG0iVMRRAKgjHF375zYC9R
6+leUxM5icMMuVLohCoALeI5RfNCbt9jnDfxzTtZv7qZa1Non2BZBU2Rb/lCQ7hS
dLQWab7HoXP+OQfQRms6nZ7dIiYHvcwYsYEBtW8PimjVwnJVQ7t7kX/W+lCseg2A
m3L6lNRxAfSz6qCwOqcACSmSQsBpe2ugrBz4GMGqslvJURINf0B8EgFtee67mCrb
AawIiKVayp8DyAIyJJs1JEILn1FEfGJB0gwv4r0F6TXUoO0N7fOfZGMiSyh3vZ73
+r+6hChYeFbTYrqTED8n1gIOAaZ99Vn+CcnLZTxgVxBiiWuEDlDDmEozlbYgxjUs
96gv+Xm2xVMIn+PQ+x/AEJzzgnjLo+lXWk1z+/5hpDQDtBR4p4iljvLu6mBI2CIY
k5GRRL+NrPFaG5rVdOAtbHqcbJV3T+2SW9SLUO75oBPSsirPFE41JtHZLJIBXp0M
8UxKIJstdNWAMS9AQaMMCnEwGwojeE/ii49l6w66yVJCLbw1GB9V6KVHcuuNjLpm
x1u6m2CtkO15V6aSAHGLBTQTlBGLCxcnwlsdY6Mbk/fvpRGBBlrkrqODrQbK06w2
ha4qOkJhgV0AjkW0tR2XeoqTo7AkhPWTH6TEAHfkkrxb6Wi+4yXrcmN1+DuTXvBt
I3S3vix0MKMgg832vPZ9ymZMYTS2zAcL3FQ5P8jSwCTNHmkfLweAhBcwa0m0GHbU
BB5PVoau9sakoY9fc8dT3nNEQNgHadbvIFic/0tGK8X8DaXGnjADutKwG+URxekL
UGsPkdG9+N61jvz3adj3IOYfeskAuVUGbfLUUZerZJI77BAQfCrNrvmT7wLneEEa
B2jRAoJuq2SCAfiLXcQRzY0NXiAYsDaP+1248ZsFs0Hq3i19RCM4Ic2qLbdT+6al
pMPN9ArPxihB0106KLYO1bwxbpBejpPfEIWHjc3eqMYZShxkBo9ni8n5NPmaVzcS
IE74C4rVgBJefTg1Nmd4LlvmOE5VylO53vnSMRytR1E1ReuUZ4UZQpmI7U2EPVbt
k5V+ktoNCa7YL5aWSPF3F9oiT5RuzyYAngSndh+JFh4BQkYhLsMBe/DGRMKyk4Im
bLqSUzR3ObmtKi+BUxiGoZ5WlqTqlvA9BqWYTd8MuOAtQcaqua5KLPUyqs9qXvTw
3LVIiGvFken7fRkGfuQPUsgGm8YwRvXPyh0uJ2ikQy+XSJVxF0NsWpoy55/vTR+o
xWbszya/+J5bQyGIJyCX2/6w+t05YO1A1qrapptEjK2IZIUlgbSP/v8VQiz78+CD
W7ZFOuobDLiOJTGi8VRvptPsIBoGEgUjtV2yT+q+YJ+PBYqrpxqYcESWBE1Sko+O
UYUsRVPLMk+3rA1HrpsugBA12APbP1E7SPD3zkPevo/5ML3P+4notAlhRlcpSnJ9
HrKzMGUc4v74mIC41ikLkfAvY8joYHkvHs35BZJBj6GCg+UodqHUosYZi2kWUEqZ
KrCBLwmXlM+dad2/h59Owbm1MVOgiolRLPxUEWJP6lr9gcO0N9aAzacnHQjf5K8t
eg1G3+N1e1l+1yKG8UmZRQUg5sN248ALBlhwvj7eYmSKxfjQti+1cHiZQsxJ3QO9
AfWF/K34Q99tkTG7ZcDTWy+Gt1soBaaniJf/DgSvCcBOkWa9+33KUup7Vhq634tH
35lDWb1+PArr/kA8BxfJS6ao1zCj3J6tb486rPpNaHTQdeiYcxpy2mdndwIBFbSQ
/jRzWTrrozdz/B4TV/itQdUU5+twhMSGPUN1LxsVPbdckDM1y+uQEewoGZq/zCOC
wEiFXXNei6R6NKXOXM/pDLrFa0tLx4FzcRdS4nTQdzBMRWSY3Y0GCMM8TwaGcS39
oIST+rXrDGkv2BZZyRc0zjsQL8AGdJZyCVS6Zowz08u0hoIv7y36wiJediJYekOf
Ax7yu6TcuilyNQ4x+om8TIF9SjmF6KcMow/GsVDLQ0fKh9zZlkEo0byjmVHKeKSX
+AmAw4BCREwVH6FRZLcba+3jzMMhsQ80arJKDR60fGSrw6Ju9lbDMzZGXQLm5k7E
mQqyR9Gum2zPdebtY5BBfurOnwc1O0sO+W00AESa5laayWulBarXivDom7mnw4R9
keRMTOG2juMlphS+/85xOAizWI0AYjvirEjtPikWXM/Yijv6WucyY5MVUyWSoQ/a
zqGyc8PCLOnWgmjHI4FJ+cw9CCk1STbAt3Hof6fpgSZhZXq+hDbShlECsoI/xuu3
fxGGkhV53ru5VjFzQ454Qcv77MyhF452gSBa8wco4FR2/vS+MHC3eAAug6DBVWtC
0YF/awNwQNS3pxA4e9tDfulGKY6zDfQjWgJl0+zJKQVVlaIdaj41I6VRGejrRRA0
tgRvM3m2QjmJ5Po/pxkmKAA6ho9mC/ddhAhA56Hyr3BegcmkQzNp6dYvDqmgBw4F
vZlXvktbNg9YVj/igG6TmKzYjkRIj8X3sVcIM1wLq2An+BHBKeOKMNUBObjbk/ov
/6fFhkh1pFwfmcf14OtJ3RG4v97TzkUE6iUIoAvEOJ7M08uFXYf0/0KFBXLK4bOU
dhHd3DkS2G4GjErpG+Y3L6hr5xrrGZLb6pzBq/kGymeoarlnBkAeb2eO68544JvZ
nx6oQMU68eLIaUV+Ad0qeD1Q6u+cEmCRq4t5DV45gpFtwL1pXM2KTcsg3kHURBYb
ZvvABGqT76YkH+XpJmke3n86WvyXVFYJ+oe2u1wpoUTofNQGIk6BUMv429WuNdqr
gzG9Hh6QFVGkrMr2YmXufnuwGiRyBy49PPiXXhFLvSRJuixF4N1u6gFzfD4J8Jgb
sI39Ik0MlIFWpRr8Wrr9m6r2yA/jgjWFjoxG4Lwt381TMAVcMHeIUflT5dG0D8J3
CPKujeJpYpJQoKdg7gaW1/4sQ0BJQ4pj5yEyP0a0CZETGXjrusjoCKlEr9jQjdK1
8bHJRQo76e8N0SAol6elxmE1pw8GG7BGzuTecG6dgua21V/skaeju3s1bKc+IDH6
e/AzUKYYi11yZ1NN3UqFl2zG3LjLQbaqbUcI+Y07hrAI2XP9wKVdL5vUkjoBZ9wP
Fd6/Vm+FU5uxIgZMwB7NO2TS9QO0n69+xQg3c56MRRxQm6wpuCC2JgjKYGczUhLu
nqlcQY9osanmRTbUTe9QVExRbnNPzvpLEpEsvS9Rcbk0+bXWpWf2hpsA+o2UEaIy
wZk4F6D62rw4ULav4nPrVmRpWfnFLXw3I0uaN/nRAfI4983h6dsXL+wTDJtPkjEf
MV84adNi+gKwKSDsxUe9K9WyVxf+S8M2xa2qrcGA1QepThEsjmyDDa+EqPnl07uw
3/qb00XYEBn7KhJTS/lLE3LrrjWjnsYJcctksc/k56gqYgnJG0NCgeESv8aV8sVI
XZuTllTNkyGH4I9pTU2eiWXkm7EpcylbE/9Y/24CPsbPVYelSO8PSzk3uz0wdbS2
9dJiRSyjAZbwWO5rgRaR49kOWcnSt6MMUiMdGMOUS/P7qbm7c9IKvUR8IpB9FSnF
NXB1I2HXfv9byqjQERR3q2P2a5XlhKUOfJ7qQx1ytA9uUKw2F6SCrpQHsG0UmTV6
dtvXHBzYPGuzcHTXfWUVQkbje3XMyyuPSd9mMB9EoK/fDR6CRCbUSY0Pw0nM5Uy4
Nirqw8syf0p/WVbqAuJaGMo3RiFbQ/ekocoiLK+000A2Suzpf2QD0vJnmEfuvjYF
jiGdzFKbrMCci0V1+BT5q+CT+/t1g9t6YsAeDR3a3c6hkcIBRnBWpgicDN+TXAbg
75y74UR8FH1HKGexYPF1OVCvnm4GzEGDAS+zsT0JNn9EhySD2Zft2H9c9VLllSD7
I342Loidskz/HWPKeboUPyiTn7IO9DE2SL39NoG9x9rred28SRBCp3bCFuGbwldD
SKXPb74y/GidQ2HevBhMtFhZ3rce4hUyMhUGK8pZZLNUwS7P/S6LlismTNgy7Xyu
Zjgps8ZePGPfkX18veS2xGnUNsw5WKlU/1uULdn1QewUQH98ECkMkfSRgn+zVu7G
cidoPgr97flxH4FJJlzrJKRIw1+/b/Arnc5zlFee465VEBOfUd3zIqj3L5E7jLSa
XyWzvUV/LmZY01ZGpUF82vsSqBlNGUGXvJyYiyW6PK+FK+kw+ZuaU7AUw9Cp5ZLy
x5TjgUzzdDEJ9MCCVxilltNh7dYc/qg3rIshWQUDoi1jqUY06+J3xNHMetZf+gPj
QfyEpx7kYttLriJZ00Xlelo0YgN0aSzBX0GkNEhqsVs2FL8duIwPo+gJx/Kab7Q1
fhPddPwIrgBNflDXElLFJghKQtSJYHvBYbRgwcQ2bKk4zYf9mxV74MjQ+fo3p0oz
lF/4/ub6dkKlgLTDS5ob5czhJgMmlGQspphbq/vbvqGxFOtEpYNDpOHrU1LFqzJG
f9QbYhr3zANZex/cO8PI4IuXAvyqpm3QcLGxkFuROH0emMJ8jSYCZjM11j+4cab0
enDEANVPyVbcorPHqc9bjZKB3G1S4c77CfX+6rxG1cySmlXAbEuAa4wheTYztCCu
cj9Y4Ggs6AtJ84b/dYMisu5Cp9xhp0t0ztLhEE2OFQIeUPs1/qgWH/wdRbapEptB
p6ruAdtn9iPitZKP5E3XPHuSCjxpFOoXLtHIo2UIaOkjOMZ59DCloMgWpmjhHiWV
bldolA3chBG2So7LiYUT9gNkmS4wDnuYzF6p3dKCSEX8Ccdj/rL2/Vv7SVUbOdk1
oemT6+iR0Uhk8mXU2jd+uBbv9dF8pzEs3goUZuaoqx6n1zCFKvLLPoAt2AihdyZd
Yuyf0XVR20PTC9Rb9rR26Nd6Y8SImDVtSgdvI/5Brn7diQPhM8cjBM/H44T6bhbL
qkf8d5B/8UWddBDoadmsw17WM8vJ5psohlius4wf5iIkoUfuA82/Iu4WztJrxWHO
Eheco0tLz4Ou+6TlW+ZRk4SOVgfbzE+WcUelYCN8HRKgrwAQpcxA3K5IH4+slCie
TZTeipayd9Bb1fPBRHMInBnQexoOEGNocdj/6ZD34BR9EW9Diu95YZfWFQYIS/Mv
Ud5noY+BnWS4xW0DywVMtXQJDQMx5128CmtFQNv+uAHPwEeNOQqhBE+68IU2SafZ
oKLUhCcUR+W2x3o6IgEgor44bq9jKRulYmYtlJsLd68YNoqabvIhSswzQUtSUOey
K3abHKeSVy8kus42yFMNOgaxZEE6huAsiadqoP2Obca8aNQVzi7DcGcj6Zc/dQqw
L/QvPx9nARL84LvMXjBQV6Fob1AggAMTipYUt8QJb8Alakug2kxJhh06oy1AoWHg
cFmVbxTc01+qlb5LB15MuetKnrdp+mEVgWOLFrk5RNAZso5k2ygXI9OAaZbj3kkk
eSmc+33s3TMq3C3MTd2+WfNLxOqtggJ01KsJWVJsV6Uc+LxmieDiWuyzCFDYozoe
tbR9ZcnzRNlvvTBKtRec6Jkc0/hULIpH89SXf68p5NBL2Eoj0Ttd3r30anS6NkQF
rGG+S8C5GFGuF6Lp41bGmM+CbBHkx32labbAIw4Y0NtCalHpL74uXmHOX39dch9e
yFyHg44gL6rknwGHu/MW693tJXMVonyI1Fb5V+Uv8sso+9STmjxDEhq9J8xybrnd
V/2GWwDe3y2bwQ9tbIYXxDnKS2ZowJkJumliDbaOkONfgnHbfWOhHNLpZ1dchzvD
EU+2+zdp8CogwyrkH5iHn/5hsT40QzwvgznTgcw8Kh+b19KJNywC1CiCxy4jgkN3
FBAcANH535myplEkgXJ9s0VPuVL1ZlhrqYTB+jgESxhiphEDrDKMN6qZgx8kELHk
VvVD1PEYMRNKrGb1BiQsQ8ywm3JXB8q5BFkT+39ExXepLuEt6K4FWGZKDU3QkCBk
A6gNA8fo/19cI+tRDtkbiJWPtIh3cTTKFPCkM2FLshac8MLwJ2bQJ1qOK54Dhd1Q
tEVHfsZXbx/cvrI8VjA5V/AkBdQ6/jLAihOt389EQoZozOP3Kn0LcQ0OQAuLeR1v
MBc9RLTPkPcpYEJ29J/3Vw5kCPIRgAYpdUoFhS1YCSpRSK1GTQUR4AkKyGas5W8X
VgnJnj3S7I5IT6pVHYiy27EonQjkOGlnXftm8vVz5cJ8rhmhcr1y1XDKx3GfChCP
vlCQi7MHAUK15ipCaWhTfZDautLFbAgBnad8tzJPZCPSS4Dn51iBP4D3oM2K+AhG
WklNkww5NZsx/8H04a7eJm6p2wGQQVNTTT3uCaewxggTISpm+IEjJ2VrrF8ateqx
ZUtsUYAT+Q12kxjJAhi9nwtClB9O8afz1UdU9pH4H8RDLCTqELVx7mMoQSSWY0Fj
fvIDTa3lQX1IvduFqziO+FrRwtZB9FkDLlESf3uS3mSC9ihnamnZN1NwbjVeNW5W
g4KtYxS9ujLhUJpEbvAW+SF/CsVo1X+vvxJfk2+udaYZUf2IldXfw4DmZqeg5BkN
nxMum9oYUnzE9hpw4gGHxLbvecXT2QaTglY1e0WOSD4RSYV49SAYO4BN0uQMfdua
5O0nMsvGExkL9HJOkIcaBgZFV6wlP84Pxeq6SetnbLU3zv7JVu95dwge7kqnqbfr
0TFI/JH5t1uERiphYFszBlcP5J+n6+SkGGC21H4cobQn/dfGPnzEzh/ygcwwEofb
2dAW0UbWUMnWMKI0eLphtGQ8IiwcRgaL3p49MexneBiBW6foivfFcavJgWsNis1y
8VcqvNVlEbx7+0HblAR794/eoDW+qLFuXH6SbxmM93WHXMMnQKLjJZAUrwjL4mue
PXQ4pFPqI2+0wHlqlkHvadzFQhBy133rRTUcnTY/CakJsQNoW6lprME2JUU6UbM6
KgEmc9pviSmI98YmsuerwVIlW4SqlIdhH0XH0OAAYVBJ9FGYgr8vwdsAN6tP3bNa
1sQvyvI+UJeTx2zj0wEkuxZusk0ECYCvfLwrJZVZ94CR1kb6TkMbr15G7ZgCraDf
GVPKFIiRAQOib89Qymn1yjZ9k8vL+quU58ZqzuiTZ4ouWpCKDo5ERIl/SVCtuLJ8
uSQI5pFKQY4K0WDWzlZuGBWXhtXYZB3nO3ubEhtm+sU1CkluT6TPWcb3p/IZplJ2
c7YPaE0obwIc5oGXOIzGWfJ6EWwkt20kdAUFL4m/dtPjIhHhc+J71JWLNpqfHXQp
G1nAe41bF+RJLJeSbyKZUx263kDW5yOmNH5qs4hXNl81rWtSlIA9ojZJRWChG1WP
Ere8hlP84LeXWeIeRbQJWEc1szkE7JM1KQhJnIPL6cpxZzjJNHLGW6Rl3++HBftK
uPoZWUIv/1qww8OzlMKgfI/eE0oJyzhG4x2jpagMjq8nGGhIevWQxX4yUMTp3g6g
QjOdt22OnimalyhusT4ugONibYPh+ydTM1b2IYi0A6nhtvB8pVvOqqRSy1Hh9vCt
oT6CnwcZKzmX2FLnZAMceYh3Wftg3OrVbphF/dHz9R0Wm7V94b/k9TsfcQVQb+me
03Zq90lbt592Vhe7Plh9FU8ZbVIrCl/Bybd593Ym0gYfC691udtxCfoJwhuFzQ+6
QBtd/S6AagRYyUgvyFqf6EBcCZhihGKrNJzAhvq1/6iE6W3tE9rihS+IWLyg9YCd
a6pbt9TlgIWcGQPxdHNXfWDWmrEJBmsPSLr8YR+CVxAL8YPfNj105Z6kKGM7VHxZ
Bc3x/t2lpdjzgLWaNh0/y9sKng1L8tyPiWXD/lgNsWErAA40dbw8bQyiemwahVxd
mD+xmVq795deSINHVpc9AdB1E0fhy7pvFotQE8KdtZygrAy5CjD5+XhQB4ByTq8M
7pr3tphmnoXeBvU7VLj7TEAIUI/4ybEA9epCKY4orkSk4T+kbj4L8nCwAxceY057
anFBq3tJHJJNxsrW+Bu5eL3Qk1SCfyykQYeW19u3T30KebMnxqYlvwKI3FHx6WwR
jMm5ukDIPGQdHDY5rIkFZiqLs40jln0SKFCbGEt03AKKsMBPtgpqBkPnPVs/rFFv
IlaFyZcBTLoBY21FZa9LOXaJvBdPSyPkxwhGGTzZQqjE9Lbaj5euph1NDNZExi0Y
1YsGmbN0QRS0h8c5tLc7QlRXN8EK7IdmtMP3Nuui18bSeuR+YzWKr5el66FwpZ/K
S9l3/xLW+p/0gT04c5AxdhQPWPR1+3r6lhSXeMd/KpM0A9t1u16pJIj1OnqHkXV0
jVHhSNtCys0LgaOmVUo7atkG+fJkn9/ifm/bxnw0zmA7igdDn/l6kIAU3ZKvQTQr
3WcytmfOytMle0KuDTDXUvGBNJI+LEIK5+hbkrUAXy3k6tQMYB/M2rOpR//K+pTH
H1C8FFubLDKG2H3r8cv8pW5QfaZJikyKbmY3PJYGG/PC6EBKn7X3tylIMGigd/5W
pRCUW1EGpws451nU3sw0xSEv9tlRpGj6tCxdfzyBHdylqAy0J9nXBsswjtgAbxvp
VatpdYv+YFsNfWnMo4r9JdwWiwyoxwS+HC/qvWOdfX08I7e2kPGlRi7eAVQZvqj0
6mT2bNYEoPMPCrF60Q6RaVPr4Ui/fbuEUTxWmyGFjUHI3uqnZA3OOyyh9cc/lt0i
wFJKSrxN3m9uXV+XCQf5NuoyWjUrpqx6UieQ3lKYGg8rFXav8uJvYtzcElxggJCr
AFN4OswmxupkGl5DQs3hLxZbg4je0f1suYmiwrwl41SPGq0eoi+Va4kzNJDXZ+mp
hXYxXQhmnwPjCsDqiZi6yycGCLQfmVP3Sf0tLh/edDpfuBRxkLayrMo8lL6fWFXg
O7Ll2zg0NS5YNJ0ctW51fx3i/4cn3zpT04hKz9wDf+0vaKqtdZWhls3u7wb+iLVE
GpL+cR7mxDXGnujGPNEOLAJwT5M1ODqtGxLMcKZXkudqv6lo7bZ+gbVpvP6T/GAF
h7fGRnnCxv8aAKSjo4DZnIKrzATRVK1rAvMjgpLb/8YUmKvkkLnmL6lj1PEL/brC
hOMN/RfOJsXFl4eseNGRKVTdt3V8Q2kfaucvb1zMBHMuxIK2K501KWyOQjBGtiD0
CFYlaBOgt/fbVDeJGs2PN6wJ0RfMCKbGfxGRlnhM7WC9r9ypCpFLDY1vebyJaJCe
+vjLo94kbY/ASXIYxgrsS2a657MpVfX5vPYQT1wT4E1i8+rdFlM2OFQ9jrKvuj+6
AwqvKwx54+f2FmtLaheorrQEvFnZnyE//e8ovxwJZauvCjgTirOpQQrdlrNEJs1z
DkTl/KXEQ/q4ouqR0n4I4W5JVqs9QKvIUz4//lfwETXQldwDCQ+V8yXlGtNUl7zt
2IZXzX13zlsyGZIijxlYZGv3xC3ljhcvDypeWIwmukYPLQLBEE9XcIBsSI3RtWhD
HqQJOsDxCpkd52rdb6NFMQleRq3ewy6hHbbbFP4iOoOaV/3l/9Ss5wsBk0rDJp14
zNuvckYl+sz5eXP54lW19FQjX9rimbOMiqY4xey/gYfKhD109HfDfWWDWE79Eh5U
EuoEzL089o5dNFGG+/Om84AmquK7O+XiUTXNE+loQNq1LUiNYJ2k/AXVmqw9EZvW
zmEDwId8JZ4JbZo9QLSdh13cfnrq/UhlxKVsdx3XxCc9vHugmqgZuvbUfLW82mlX
ScDzo1nL+3tWAFkbQfvU3LozUtCfgu0PAdlOU5QnqB1IMW5ljwBy3VJbU4J/puJO
r/GdTNhVnppd7py8oXt2xwqho+z+MxOVMQIOc4k3kXq3m95uL4OyvPNi3hpwpNol
3CO4zdDbIXAOpiv3atxptYNKMfXQfV8+2zR25H7HOSilJU+RoI+niDkXIO9SuM/X
E41iNaVWI9s5x1krb+dm19UzEGMCzGeIw8AmcRGdV1rH+GXYA2/xWM0jx3ab81SP
gUh0E1U+XZhyJRERcJd68JNcFiz2xpxUz7mSNdS6f4OO7zudxiQEN2DrpPELRAmd
r1osZOgvg/bNL7hERaczRk3PHmsiGiX9Wl3vRo1q1VaeDTM/0cCCuSP0O701T43v
8C+BnCB/ZAgH1+PGy8dDzuX17AStyr58jFh1OYC3j70eFZPL1wS94MxOjAJd0MtJ
sCenJPciSB8NzHIbOrX3jYhouOSNNXWNRKHIkZiYdQu89pk9td4aqZfEMvmso+LZ
rKPjLJjFJuee2zvD6kGRV8fQglGHPR8XXdA34tM8Ukn3b66b6rY02oqd41Iz4DN/
Ql5SmGDzZ2KtfoH2Q5uM/ZQGqkamUNiSQy0IvJm6d1OSpPjuz6f/l1hJZR+2mmfK
ZI9gaZz0WsBcuBLSDz0Y7Qk/lgMzYwjQFjEvwJUGAkF28anujrWuXjBWat/IvqLW
naBg3P7ShOGNYO6KhYtlqGtg5DwE/Fky8Z8zYfLprhz2o5l5O02Uf4wdKbyt2v1c
UXtqC47uxDMXbHZqQWbYI9EuXNZsq3D1P2yZt5g0kacsOtf4OFA4h6tDeJDmBxFN
18C5UqDoqKssQ4dttPpQWiI5ua7qXcnb5jWdD6xy9hALWn88hqXwoLCzfTK0hWSs
HRS5LhYNF99jHc78LlZqi248n28ul6KaTjgnO0KqVbp53pBARgOeSDvdT2idlA5T
fUp2kZJqcDSR9/H0uD2XCN6HU6iCJbC2St5ypCzupVWpBmGcOAT0QJPyGspVY6fg
mjdYbw9VY/vk/R7tvLSCOHBPQkgqjuvIYp4fDv0X/OUFXqSTrjulN18eyxKwV0sX
cdulvEEFkPyLhVNXuRrpWOTGVv+3r+rj56gSGR7+uVfbjGYf36iYyoRNPyZjVUes
puuQSIIvGudWn9zbXKO0xXUkiORTLZAshTxkltmWz1CnpaTIDSlBrizTs3uHQJh+
HTOI5snW88RVnjQjuYrZwWMAfjPj8Os5XaNEzTrfykTIPL93tQt2f6A/MFfjmYoV
YghWZnkmWLbpVSbgtZVEpHJnte/DkVF3FxXW1RG19xjgxLQj7v8Hnlh3MUxTDI4C
SeMwJ0IO6bZ5w5f+a3tJS2jGNkFHL6mtJLE3xDdEbzIBWErxzx5gWHpxTm4HsqW6
aF7MZPtbCflGJ3oiL6y3ti2qJA6W/VHDEazIvYEAlHBsUu3+C8NVSE3tzPDstrW1
W6FJyEWnq4ZXshMsdct9IYRuzmgrQiLf3fZgEvtPueYLgpuYtXUhCEnhK1nkctk+
Fjd+WPWSd2zvo/SyBIcpvPAFNeLOgRCxqCsO0QEYxorY1arJNsv7GEpuVYxIJrMa
XDBJ0lADL/dKM586s1scLO6185lr4FEd0641vH4o3wZeyOYZtlFlI/ldQ8jyHci1
byc+RhJuyoO/LbjfbvIqY0G2AxegWAS/bzOerC5ChL5o+K+xPJE4L5pCS5NK6+JK
7hyNQ9893CYqzX2WG4YSbDh2qwUJnInVx4jf+1nRV5dNOo3lxnTILpSmBU281ujl
xUi67MRB0Egtym+sClc1+AfrzAbOD+4KdYC2Cd0/K1QHMXPngwmygC2u4A+2OK+a
UHUjpWoMWXHb5a2YZgKjRAkud4yfVrzsY4X+aMkANnbfc5do6pOl+/XJWLGFo3ym
eAViR8GplVqxZH48k2xuL5sQtk+sg02bLFnX6hLqzMwW7gieDJEmLzmPZE9p1V4i
2RX3I8vVNXoFBumYoordjibfitzIvEzTjrXZ2g9DsmnaFlW7Y8739Xx6ci8vh1a6
jiGGai1NNcx+V1wpFOYXTiNSjvFYbot855pWbelrqXg6vo24wy23/CSmfu5T1Mjs
OI49LsWBIsfhmMQvffrzLw5ZI0ocjg/dGVMruQudfjZSsG8Cz1oh4biS9q86uca1
Cilo9gHBIR9MM4Z3cYHHbXuwKYlSwQNioIsTMUVQy8JEjj7LBMvyuYtYT+9vFx9O
YIXuuaC84mOq6DBdyLQlQQz1YZJnh/sPfYjkk0+dMkADyZw9qs/QekFKpxud8y+T
z6z0/SfRxE98oDn45k4WrDGxLQmkkZEJjfn4e1C2KDIM4GXUpUEPtnjiCx6PK3sn
scj6NNJxird0UNI77hXMJuHLq1LG8JuFR4txlTjnhvmQaD6i9LcCHFFXmwlZMIvk
X9HEuePpHuvOQME2/ouO2+tMwwk33wxDYklZ+n2gVq5nmBVBFca3V2bVriFEJwPb
4Dhpcjw0v9YfsrqPn7hv27ZCXgTvNOulxGrxgs4r21cg5pH5n/Zm5SlgYf1pfk4a
QOEzX3rRJ2/6jdmlpxfjgmlUdyONy2eqkPiPevRLp0uSzmFKHs+glhXZ5lxau6BZ
Zfv8WgMdn/0QUeGdaNjcPnS+2Fx6+/TJ+M5MAPeMZyGQYNjfVBz0S0okdDVEO3ja
W0O/Pw7riJPE6NQ+IZjtuWikNpCMXL4z6eTZ3x//YRljQue8X9P8mwUYBR9mU4j6
Eq/kG3HadLVt1FsYJcyTl0GZnsF6TbD0zfwyGuMHqzloi6dtbHVtMc43T9TA+EDL
u1wjJ0YoVYwr+s4JCeNgdINtqynZJafI+y2JD0oZFCa/1iv0M6sNlbXbxps7jX6Y
WYFnFqn85+01yVHVGbv8mU682QCeRar8zHuTSfwbvml2BVWeRUvVSlizPijGgLrA
dUQDmDx4h4exVf4aeDdM4+nQvm2hyPtIBsMoHbwmiqcOiau1MjG+rqdmDlg4vG8Z
WPXZqdR1zvxZforkGBayejYjJAmnO6tjf2zD0ZCMQHIgBuGIOnXIOfpTPtiOz0YJ
r5HMQfbGIfxNLoSi/PT1oZrnGRZIhaAtPIwg60HmziJhHIKzezQTvLu0bsRFR8pz
3vZEXYdZ2OdjnOsQyfPjpxTM0kI98IjA6Ff99htKJ8wPiFE+0Fu7uicmyBIGGjkj
B5zX+ztxKTX8kFhR2ufge3hDp/Xn2k9qoI+YPBjbpGQSL8snqJCtFf/DDJ9Mj2QQ
E7o4rm3kdnjUWKWpj2If+i3eEqXuQKT0J+lQDnhOaPrjKqgb44RkvpAZBRBdO06Z
yhYKNz+2Rgf+w38tAkgDClZoTeTL+VFHw2+kflE/JuA0qmtxrcxFXVVeSaBb36vJ
bLO9wLCuj1IhG/yn+i75iQE+NLWlNlH41JxwwW/TwkKv7MV/Um+QAYJRNxSA6S7k
PpjtVHHmJMajokXR5KqD5yF13XiIPvQDIpQxfqGMRk+cjaR6kpFv23xdpfKQXxgw
TlopbFhJw6m5csehe+z4GN65L9O1aigQnfe2D/T6nElKlTAkmvqVlZuCVHddlEC4
UiBMxZaEp77C0W1ITq2WoE9lcBv+7yhgUh7Fnfv1P8WfCe1luMIuEQQZiWsDR44j
iU+VPvCUxs964G8DNk4914lTC2kSGBS3KrBQ6msSCFir2RJMd0HYQxqb8cHdjw1G
upv9ZzUDRAziv5fNWqwfQ7Cyl02mHGyhdTppPBg9O08+qqVCxrrKFjdANZR5fp29
KRUE/sXG2UTaNh83EkheyNvepwccpnduFltT12ZETyAsqOVq2WLtLd04jR1llLZE
qzIIx13++32S3C7+kmdSstg3wxzpXOyZBPQIHA+hp4smHuFQjXMoDq0mFI/HOeJu
CCPmDF3/71nD1ZBM1StZq+dVmhjjjFT/PfzFPThq5o3pBfJEN72HwWqYHCQ4N2Kb
z2eh0RPt3Dn6IawozpqLCboSWDQocEKw8BXXZgYuz7bS0WbXf8BCqlWvvc3ng4N2
csnJs3bxSIEhRi+x5x5YYz0qjpAhQbSW3P5cWg5HzWdZ+BVWnPjJR9P6EO1dGi8u
8VpS8XwsZbUyO3J8++Z8diypxzQ2uGkR8gPdSg7ASH4ZXFkiVwPsWoicdPGIy/Zi
K2kyf7Q/Sq/xO8+Rs4IvECnEp3kmNjpNpzfOrS3umexhzhrdSx9O/K8zSYzAaGDI
UH2KQm5IDZKMFKBrbuiHbUMS8BfyNpYLSd6IzKzpCgQMNGUE0qaHHBR1gSeSdGao
AcwG9Ij58JiSvc8WIkGp7NrJOapzpnROkFF+/PvMWQfViOJJvEtARlUqjV4RAcjj
B/p9jZ1hf4+jxXY0GmG8x/3h2/YtaC/A9O9e4udtm+zn3hzZZSaVqBxMcJdkSJdO
/SmJrFjeaOWhILyNMeD+fadnI9mrF60aJdWeuMBRoHW6VshI5TfqZOzvCzCfdnaQ
7PiBeqR7BQCx938SznQ3ThTa0BFc+Ussh/XXKhzQ2H+4N6uUGO814WxpL3E3Mlw7
cyGubuvIxBgzxGYUFEcJ21JFg/zUOr3OOktJ9Nqe8k7f3VBHGSMKdu9zwqtq85+P
EAvn46Ghh3cXFHQd2gfhefxjV/OX//XrrbKapCNhFvjB+FUJK2/JMK0BeIMT3pEM
dPlq0+M+/nuBIblhLyULoqUk9fU/7z/qZa5TW2KJ9Es0alU08W3TbBXv5zbL4GZX
pGC7JRDqdjaSQyl9PzvM+rZk1AL6ayOI6TzLtMrYWsXtbCrIbFeYDiZ0qmWgLBFO
9yZ2vGsAi+dg9hb17wUZEagT6o+MyDJInTnvoEGa+i74qh/r0aZ1l4wudI5jyXog
l8lOqxYO8ferMV866fUKIH7MrljhPqHP2S3jVbjJW1eHOuljn+qa+otkHSpDbj3n
Gcq5+UaIsD7bMLhLq2rxQPtOpluN/nt8e/X4SqMX/Bj5Ad8Oarm/ZUOcDm4dRN5u
aCTLimJwJsnzv8SRJ6r9xME48VUyjHdwkrPtaNLOh2uTfgmiygYPpwsedB9zcLCU
3neheAToCM3BXWkeWZoxAxWKoLSGgCgspcx+ZyS5bKOJ8RO3IzZdl13hcggXhinU
Bj/y4Hh4nxkkvJPwpdFl+T/xpUSH5UalSPqksfeMHaIiCb2TtH0Yx8XdyLPGmTwi
3PSRbYwargy6lbKiO3qOSRUAr6NTBgYkNLhItkK6k/lh4QJRCQlaIJ2KQAK3Z5Dl
ARcBbTk4i3Yx1Ld2tRzplk+xgKDtn64vgb58tlycWbiDbmItdwndS0y+W4LZUqN5
E7rE2/7w5zJfIwOfX0b5BxdLSHPAtTRCZta8t9cTeJCUH/5cldTL+LXnmWV2UMHD
Oo+n6f6o68il2SPgWJ30kYFCK3487Hme3YzgVnUVaqa2nHkQf+LTNMjlqFVxloc5
j8HwfMpkLs1EAXShGeTfjFX3Vm1MXEMlDiMSia7JLOUKUr/Xkzt7FWQ2BnkGmORZ
4n4x3+bUi4Q8P4mrnXZxE3D0H3ocHM8xQiOrGihg8lR5h53MJlXdu4i0sTF2iVFw
WJuPnoIJKyf+FV7Sl55zJG/UrwPA3lmWDMYui1vG/0xuEVYjt/rNwcDqqOXM6ENK
TVjPcF17xRKXTf2OfeOy11vAAUsbG7JBaz+W04cyMInec6XSYhfUqxpG4JgqFUhx
/eoj1Qr7tQS4lFOMVtMm8lU2CFXQUCH9nley08qT0EQtgxGHYumqLnXly+0MSuFV
25RbzGdtjAkYapS55UPcCFUpTiRSGEA8pv0KehW4pHRbZ5UEGSBG6FZBQTlw05im
Po/bjWGAkOcuwZLBeR/eyrt/sGSs6cAjoG2bB7oPhv7FvBIcdSZK99n76asAGdu3
d6Jxal4maT/ohdaRZnNsdn/nnUiNNRKDcHsTW9bGp8Uqwxt6WWAS3ZPam7fEWEGr
ST/viE+7zWc3J9PlOHNgNbHLzJhdoaZ1fxMICK40Mkeb7ygGDlM3wSOWoo3e1EED
V74AazkKap4NvOKXq/awA0rmwp3f++y7CUxAslCYAuf51ZEsuJqSfH3BsxDZLK+9
B73iAO/3OBoNwtbKIdJXhJug5JjIiFJ+foM1Nn/blXf4kPmhOW7tgptBdoaFpbD3
XnIP/9xwHbmkYeeIJmd97/9XpvOR5voCOUD16Z3a61CzlbmHJyixzdOLgVgLERlL
zYqLwvoFncU9Ez4g5+effagtJtAiS/F0AQg465KMwapyWA3Z3o0q4rPXo9Nt/vOA
HvfytR47yAqr2XqFtuq5tvnMWLeJ9DyjEr4+crwj/zev2llRX7qpvERhKoOJshIp
WjYIfVJc0Z0Xe6VjwaQmxx47qRA291qtDVxyGsLQlicNHV1iuelTZ3qurvatSkdF
jACRjLS4Dlyc7NGDWIKWkljspXyBrn+zrsKvAe72t3KE4mtRZQ7MhDkJG2nFgOJ+
ORSZ3gjps9SJW4K+78mXyiFf8YZpJunc1kbnJkpnn7LyDJ/39fqnRnZBTqDo2hsp
XxaT1X53lIRvzK5myhorrUO5Zx9S51kT9rZzOucf6BWHLOODfNVtx2zMrdMS53+Y
VKg+NvMOkZQRahzXLLsJLRQZufMvPs387VPda+79YPCR/anELrZkFjOdlAPo8oxZ
R8hCK5wCzIhjzsK+IYgUQvHnAYr436fjmBovvneNYg6o8yS3dJRc/bpnKmVX56sN
PEINCapJlOeNLLhLvebRwGoVnE7b+ilPZD/zyCftK5wjZQyJw8wkvmPORCs/AOAV
+oZRuwfn867iBWjAVqTDFejMZbfAbFDL7l9KpTjZrSFISA+73QfKXFzc6M/sbYWa
0hAsFuR/Rgj/MOfi87os0JoKnC9OYuPUjkBRCfJWegyS/Ctik3r2HkhFrmnE76Q0
jqm4v4FSnPXIuDnePLAYf1Z7BeopOyzvEPHlq4k8hI0ObW7gFUw1rIPb5wV7CQhV
TjRbxKidRNAW1Vcg5N5ubuTtBRZL2iLEwLGgfr1NxTeFjxpYeZgBbPGzrj0/86zv
ONMz4TJ6F8zrBtergOKXtOenhLh0/k24t1tcENqH/za5gbRO9/jy5MkEPbhBSBUZ
HSqpkymRu0jVBhkF9y3N+APnW1TuAKQ+BTKd9/59fxkCyYFgfI8pA/GvhvvRMe/K
+Z2awN9XM2BKFgCZczT6MUhgIoMds7x+lL2BzbVcV/BOsIcsm+meFvG9kq9zlNxb
cOyYXdTuP+NdLt+GgVxzXf7iqh0fsOG3Jfel9QWnZwtlUEcnIj4agX+fv08sPnc2
pxyaEIyt9yFKxvGiFVdLFA+QIaEA+ia5smsXz27QUWPf0kR4MQ29LOlvQm/eLGG+
SSjqBRrRdgiw3ys2cKc/Zlzq/K4MW+jJBKNH/bU29T1WUaTE+mz9MtjO1AuYFeAg
PIzFQwEEevj9jLA3SJx6yOH506RFhs8os+kSiA2ERbMv7lw3xfTwg3cGz2LxObjz
xFjqdKnoBEkIuEhSKTUPT4Uy6Bp6sU1HcTwsGd6aVWiMRv6oRoD7M3BCuSUYBWxS
lVQVsByAgdqUNWa023XtsWH86Dzop3e3S0luDAlDMLjy+j+zbAEfM+CH+ywkfiW4
Byq8kshj90qm0emyNOSfu7n7giJ8idPT71UMf1RU+MXPNNv/RvNuhXxeEC7IrBrD
5KzLXE7v+1gG9JxKEmH+fvQt73HBdcq0+Qx763nkcC/s+wdnV0IWxGk61SKFTMjq
zGaSQDVEKS6uecmHtlqbVt+Vqw3702mPFmBXqz9vnlBXn+S/WYv8cyZQhbnr9wKY
rnkcRuy7AFTjMLFA0KJSRE/qmI0cvH8bx4WgPvJLBAJFfxqIMPgJjlK83gxEVL8o
NRqyX1jr0+FN4hUvzYgJ/U5xUotXX4ueihvG6Vl1xymqjZDYWASEymuApQDHV51B
zK9VATBYNJXqhTKgzG9F4pF8BKOBhP6Lvbrfkyh9cmFLoGCqB9YajCfzQVpwUU1v
wQxZKeg/9mQRNOcvRmzHqR3OvauP0Kw2S9UxWalqFfYX02olpVZeuTJF1GK4cvfI
UOVIBaDsJqpCUOnCCXYoNwcJsZlSTndxP+XqIcGyI8KE6SCWfK/BKeRQQkyfGB7V
xfhyQtR1z9GggvA/40WdlQrTx+sI9SeZ/VQu076DkyCHU+7ttB+M5mt+H08WxgaU
YIGtMuXrvOHbDI4JCEtMaaldEUUqTHdpyzPC9IOf4Eiyy1owAlB2KMSOsDEEGweq
x9e0Q4cOp2EY+v9iYVzpDdrCDgm3kL2B4o3KUI6sxWdz66ZFckfySuEmCL0l++dS
DyTVWzhdOBk48MZwm0dr6DagHwbl00gsdbOhGr8oCT43nKJ7SB5MW09gvC+VyDMM
Jxtm7ZZ0GbOiQinqpGByAQoVI/7kHdB4sB8E2BM7ApqpmpiIR98pgqQ4DQ+FYTAH
r9LnJ9G3ZeYDt+cT9fNA8gJ5wZ9upuAt1M69Op7TaaSNPFd+YHyCU38aTH2DY6qW
uP0LcnoA9eNMOGpR/dnsBYerm60yAWcZ7LoQG0k7XTsyyYSPqcL2+koteSJEnH5c
4TDeLbfQKTo3xG/S+w074QzFo1996K+I1o98j51hrEOVdDHqmSXeQMPUxwqitS4n
JluSr/z0VWdd1c6hCYb6azFcEnIwex05psxslKmHVx73MIXCem8THTiOGeN2BDaN
OVS2DGJK+soPo59L8UsDobRTPcJWw5XLY3TAgoM4af6KFMGW1QA6nEqLomhqvtBr
9yIMK9K7lM7t4ca1pQZxQsKyAworYv3xpqzCbY0OVMsLv79RdrFFeJenCmAg8Ydc
weNugyf0H0wX/EgeTtTt98dHKnPdoMaoXjSpANCo0SJ/VrrfFZGW22P5Ly2p9AFJ
k3JDjjpUMwCUWL1xV0ACvj+8HGi5CtHM8/4mA/MRu7DZ3YOdo7bDLChEUP4n3E6E
KkQOAMb3oL5PVtM2Mbw9c3PexfK1FACNBr0lDGZK83rwP2VOEDvyBf/7LYH+40eb
xiOKqpwg36ish9jaKgas/6idF9CFXaHFuhRsYxmO1kZ2pFrrA6MKmAy5iYHZdKjz
Ohal9pBX08DNnbGvqfKg8O2MsS1QDnGydPwZiBzY5POaj0W1A5TvZAZ1NgFlZgl1
sgZSHi4aKT1nCfxQRYZmWsBzAiHX1s/g0jqCMcxsVChueycgOcN9gqCdGp87IqMV
Oh2NyqF0MVmyOBf+cr9rzug7BKZwU9dx/VSzHNnPiZ5YqQkIt5TUxZLQ5BhV5wcY
zTaJ/Rg6IzzwrxkCWacylen75dXOd7wa1WC1dO2ImwXhdRzpE3O04Wy7ScF34sI5
czWZu2vO40IbOV+p2AYKkF8QxC+TDbBFE94UmRwMjb+aiNUBIhhRqHo7buHW5MAK
XUgcsGiifgGxAHVySdZAg3BD7bVyr+BdBnNYH2cI8IL2ZcoCGfA9OnpY1rqG5/ly
LxD06r8WJeNwDSuORgbN5EdQdzWKr+94DtB8QOIIR3TeJPjoSrVcWomSrC5cjhGr
2m28zyJX/24+d9SPGgJSmr8kUjh+A/uQ1Th4eDLk/V9ZA7tlAF+UAu/VGUI2zbYw
QMpbUFViTjtRacVH89BhDtg9nzHbKXpZoXGCzXud855QgfKBivFHm8Usu5ud5JzI
14vRbmfBuOXsqVeG7vr5SYiqI/5Pr6Dzit0zAGsrraiT4uMjRaLJkICYDqea81aT
Y6Unzav0NKhYDuEMZhS1i6b3h5T4t6slGUsP0y/KhpIiaSOR4Kb9WWCFfgZj/6tC
LwfPNVEgMiDt2FbNBiiZpH15NXq/qmFT3UtC5QcOl3gWACEhpfw/dDHSJpjyu7tk
+f6D4D8DuhQleDDC1CscQR8TVU7CJVNpNhdmGgXKhMa6NU2KBDc5T3upT3rQ3q0Y
fq4tQwwgGf1GnywVYUf5XmY8fRQk3+f+Jw/L81nGTPuHiiN3LSLFk7as70BM5sYv
Ab/nI/LdrSGiCxF47XzM080RBAyv7IvWr+WSVvI++UyPLXXULuNMyg12z49hl6uQ
JTlXz3z9ZWBMYrExmZsH48jtEEdHGI+cldQMVur2HSS8GOpmrT2KghGrTgRrFlml
TVsPNZGlMStrVE9Ku4gPpBBxzWr+YKco7tPw/+Q8kfqjtHK3fzU3zx03CNJt974U
TpSAFRfAFjjXIw1W6JXc8UFbMMDWmq6l/pWEIygP+Q3ffAX1+eI+JIGpg1rEuYEU
3juN5gcglu2V3uWnQcQb0RLNYkhjj251AIuxyMCICfnDn+GlfqzLw5qhu0uUNUpf
bvQN6qYyLZZ3n55/lW6Zz4AJmbA4lBNdJ5RrJGI/1YZtKUSI+Y13f7Q1UVodVUd6
AnlKkXvAGi4Kj304nSG4Mj8vz/Lb9jdN2wiQi9wSo1epkp1T+s2C2Ci0ArBT3Bsk
cCuY2dN9L+boV10DueJyOkQ0hF9x5utvj8bkph+h1BdCp1KuCxACGsv3FGhhR8MJ
EREzrhJnii6y1+mQExOARSHYBm3+63U5+ylHDJrgpRQ4uJwVAoZLQAAsE+rU4JJm
ZthnRVhWy28VbVd1WcLi1gJ0KioSc3oyhMQdU5G/N7jD79sl/ztE4U7f2OaZIeBa
uBzDHvlhqrzxkh6VZv1ytHiI0zktk8MhTdUFVIhmkCFlnEAdawj+JBGHiymo22kw
c3zcF5fQzsk7PMb2t4O2bfGEHGprVv8WUbA51qjnOcsTWlaRRVD//bK0FRxCsmBK
0xK07wk/3v1wSzvBkKTFO15EkQJh6slDNvWtCnRQ+olbkbXItW17ti4iR5kcfcqz
nw+B4D9HkSi8/ylUVawAKBoE7BUvLsSeQ8pgp1mSuSLVXdOWCSFmCeImRkMRjew/
sQY6TnChYyCp6V35Aoh/vB+voXSlDEcPFq+OwWhbhyu3TnSzrnqQJiodjS1MBjD5
QI+8UvrBz3VbsU1Nd4wbaA7T2gp6/5SmHKa7Wq6rk1W5EmVunw/+32J7uS+W935Q
95PeoiD+F8pEXcscx8qkFocb5V94DHyvIaV+gg7VYfMG6Z2sOrba2msOQOJC9GxP
+56gDC96OMFPbRAjmcqRpFKqaZqKS3eLXx56wHuwJzn4eGkSOLHnvzn89WEddbwR
AfcobA2Wb2fgXjttXIKFKS5M872YljO7nkPRRyv2Yh5lgSrSWg8MdnYy5IkplcCA
a57QzGb/XNUOd64f2NiQ9AVWT9clXr0zYP5FsMHF3+G+ZxLjjJhxfGyHdvS0SFjq
2apdJTqXw+Q/W9WGkyUAmevYXE1XPPBZ+ifFMxWkNFz65a7vEwngrXtEI4m1f5DX
hCmSnuaRBT/AmMilP+BzynnrW6rG7hoAd+ta8mfE2YB2J0FUgt4lVIsig5JV7z/q
N6Y5ZKj9Mu5GeGi9kHMQ3I05h7ErBFIQwo+FJFEKDOofcQENiNQaecIzMqf1aDJL
jypwC9h0X7pAHjL+xChrIQCuGtGTkmTlkh9gNu50HdH6W4BGl71APFEtV4SF2Jq7
gKlfXWjLpwdrjB9IrGj2Y8/TR3xtzSXBGQlf8TmXiJn3XSFeWzabmfrx1k3OWcgZ
1leT6cXrj2yuPm7qn6fhWoT7qK95qcO1wDkwTEKapB6stnESEgFotv4hTJaZVNA1
hu6xTkKfQ5qPzUrqGCyalAyNe6m8nAEJVfGU/GUvcr5m9Bmj5Q5+tIk2vpXmQZTV
87RTK1BSArZy6gTANa1jMCvIDiw3Us6/lGNYbrrJ0mNMu2IlKvKQa8WRJAhOlijk
u1K8WX1dUtdGVH5GzeyDfz1h1nFH+1jHMMIU4jnMIh5pDDoxifYZGj5WLJrxPr72
xx5u4LKfNdXJK4pPPxWv8eI9sT1lPzpDA6Wm3TlGA8JqYivOzrI+mDxJQuMKY9iz
NPc7/DwuNj1bNlKlVzfEjuvd7oWesZA9OcqOQX4dK4hYvWENxfV79JD+4j+I1zns
SL5RJlHA7A5KgYu2DWZf0BrTm502Ozrrs20/+9p/QDPOGDe/erj8zVyoUNH+UDw/
d2eu+F4aHbrOt24DF38gSNRoOs/iWfEo3D2/mdgjO3vz/YIHz1ob7SV2FdVZQtGz
cv2rc6a5P+1LBjhNYG5mUL1zuwUUolG3MGCwV8bwak8T9cCP0BnTTW92coXDISo6
NcsaTJxBquD6W72/bc5YdsvAF9fMb1O9LXYsexKT3MtIKkWaBBR1qfvlgNxtHcSD
qn51gwafTWFdh8WdjFfCeQHc4MxdwRyMq/KJnLWu5X1jCgU6kjB04sR0MGSKFBxX
MArS+5lzCR5KbA0SC1Zwze+W0z6momNTtHvPqyCJUcS8cL9S4EvtVPDuyJaPP2TL
s6M3XiVS1sCYIBOem/5+ZFhN7BwjmFlEKMPCRFBQqbgTvITRPCJ2s91f5gGFSxfY
cJSr2AnjNybsXDv0ENRb5Lh90Oe8cS3VK3wEsQsVckhy7DizyzoVrmkkbbm4z9mz
kzrr5lXHDMlh6nfJRGw/rbtxlxoH2Utpzmz83004HG9HQskLw521wGYLbynITmYj
4c2OKziizGSqoqDhc++sGpjkzh7/DX5ut1LExfpjeHOf/+r8DOMTWiNQH2QKU9Dl
K2aMycrkgVhmm7nUKBWqdQ+DTNI0GbOmp7uf/yAUKIbY/ve1FNzsw4lTCvZyHmSy
yekj5dfxc1uHiuKH+GMBBl5krtnUkMnNoaLqD9Fdvs6cHUeALzPRJh0wQznKc0tp
ex5D9vqVaECitRuA8S4PdewLnpRI+cPtm8NOFvV39pjMwLkCZ1oPokx7iioWoNLs
oz0rx003Xey9iKXQcM+ZlEJGCUw9keW2rgjx63gmsmR6cL5NOhf0wmIFSLkojOmF
ev1fXyUbRbT3gGJIdDY6DMiFw44DRtR2K0/CoI7a/QA0KPHyfs/ZlFhN8zc9wPN8
lsJoG2G3bePNr1PGnF51v/wBa8xciU9SPWEA1+LUzT8+dj69s6wryZOI3uKGDi/c
0ZSow+dp5dwzdvjvmGNuvYotdMEcxWMtKXK+VpCrAwMxGiJutWCUoG6RsTFsF+8N
2F2wrOS0L9zehMz4ALdiFMTfN78qDfG1s8DWG2eqfkvunG2QjpEhVh1OXWdLWGQH
poXvEw9WWO/te14ghNWas0EzZHiK3Z7l6CdstpUAxStximUYuUV7W/oPUmie2lfl
yCuv7Um5dAJl+Dgqp5xe0+423MbwqmdfcRG+uVRENK7dzrtSFayNZ7up5bQiS+Um
gj7KInRGzE69dmK1YXZutTzSlpU3QfGe6yV1Nlh66kBiysLvDVkB437ogGagx7vW
/QPTRY1lipcjqwnlW+uViiqEMe6JpRmxIsfSOGDlVCdAwnYFGAnLwswwyR+FdEZO
SA1EgW2zSHIw8nus04gNa2NVcXiDYMzMC9XPdY2tnyKB1iQ5h2y2grCEbKeC6lLv
a2Uja2lgGycg3nW3/iRn+/sZZDrXITbHmMK0EeBWfZNvjRcpVnfP3YDsLNcdZVBO
Ek4VHmv+PUcb4p/bArdn6plxkb5RQUYND2MlDX/8DjHTXq5dDJ/mgYWkYcgb3rRt
rGLHJOMS6+ab6VZ7a7p4E/eyoWnr2UjQVVpb9XHaBR+r7ZSzc7n7F0b6KBkHDwwq
F+b4O8P4LwjJb36hBDpbcTnRLIBcGz9p4gxPIYdFvYlaHSfo9ZQhp4S4KZ9ESR8g
noYYQ4gnVSm5cthaLbVddDR3am6NGObf3WYRoSAn3tiLtuI4S+eKPEbtV0EgWtkr
We6Qj2MwNdh35rlfvckcvTk5Bf1XldYCA3oGxK9XJpl2lIQGDRDDO5GDJWnYhBw6
5uXPVzwGpkOpN+Z23tpUpc4fiHLhmhJyqKYy16vrLjvkwcnUL7oGLy/0ng6kjYiw
EgFbEqOM3N/Aq9I1SQikGFrdbHoEN0ZtTTwML/iAIwLseFjCwqEH6AoPJ0LiSOHX
iYHojeOjbJgetjcWy/0BsIgCBCtiIf28ij4WFoLzm8+S+aTsbzF7LE7gbK0kqwth
jYAi846skQ08terMI6pqx9U8wrpN+8QCpCZBYDkRHhobcx9bSH/mmvsYFoXeWnSz
jkXBW7rsxXGVH94lp1tflTTLiGUi471TfDjhyhSQVui9ULCYIfb2TG5gAwsEqSEq
++Awvv+zGDwuavxq3YDkjt8S6aF4dWvNyRbsZICWfzP8DNrMdv1Lt5lW9O2TJIEt
uF6lWrZjjz6BTNSjn4NUYDq3QABXwXHg1xdjzLfdQJ1pipXwgqWi6/UL1MQxr7yE
9ekJTTht5ZMe15YT01jkj6rGSNpiI5C7KAVed8C+cs0OL2+AIH+6IYsYB67wJiFi
09o0AgNjvwtCb5UlFqB4L6VOmJiEvjcqVIQzhoImRXVY96TkNVH+bDpwBIfD+RIW
Q7qrfpCE5VCzVQ3lWbUjz9O3jp5pbpBPF0QkIky7SFm/x4fHdMlDcks4SnYcUtFD
Tf5HYrm6tDAKrjrs9eVviKJESDqUIRo06bfTiC+343CuHVOBYoazKkPaPQkrDlli
Fk/GSd6Lnx2KJmzJFQuWDBfwYSYwVH/C9KhOB6jGMiuyo6JMytntrUctDY8yuFhk
jGAbLobPSl1YVgF+9jzA4JOzzqSFjCI2+QloCslqDSpeKwHioaopmwMjE6gQLk+Q
EXU66OcjKkPXLvVglmn+5ZvP5GUirBf9ewPct02RO2BdmiwAKvrPI0WSDxwF6ns+
xRN6iWMIBy2DlzK2EGqqrbKkmvIc91euacIbN+ZiBWwXPP7nzK34RPHS0kckXXOG
vxfBohjlAthBE5JzZqkg3c2wu1uaE0oFM+z1RsFL1Luj380k9ScRnAXedUuZONco
Onbt32FjgvWhkl3khrEINu1pzZS+xNWOAUrgUVENGZssz68FZGh5Bch1DZlREr5Z
bzjn/j/yH4E24SrIVVdohFm2qFXMy91ZNCDW/s6xt47JXfieM7XZsoQ34TQwRikg
hBrA/xueWNUUoBEddJ5Gaa8fsUmLKTUThq9GycM2Wq5L6crsPdmFwizV322RMcTV
YZGv3QLfaqitUDjIUN7kwuS1rSeH+9O7VNAI+6zuFv0muLhGaUrOkA9mjt6Mdxkf
f4j0RhcD8iCEkAbJ+bCA94Xj0u8az2qSajJYv8Rf0PBDjAgCJum6Lrm6+oZTWtFf
DEj7kZkcb4dlcieNDA7oBJTHR4atBuI15Wty3/oAHsbC/Toda1RQFXckbMrNe/zL
muRKzG+u2UAQYvZrN8JMrUpsQ6fC7d2XwjJHR4J9JBKhMynPTuVnEq5EnVLrxFot
Qj9G9OgF8bx+76z1g+7Wiix/5WmLt5csDY9WLo6PBzXNhimWgkejFV9Biq2otw/W
qYUCrtNpUHMces0m6IfnxGmzgXHMLHAT7iIARftwdpu4cNg+JmSymIMtv2mCueZ7
eIMu6FvIBX375+dgQtvlka6XpRO8g73YBzqrGbO1bcRE6lZDiKnh0uX32hQNNvDV
SW+LOqbG8ixpR3kw6kHjpEceVQALCh9nDqhkLKhYky9xaPRC0YoegPO4YzN2pH4P
L1iWyWaRjZzqT+s+SDSYzn4qeHESEP8R8zSMCFg1gQeBPvleyjtHE1LRrjkwzXZ/
5rQ0yWsomTlyzJkOLGMLrAV6ZphgWEE5Wn2T1dNFBvwoULbDKaea9pAfefKABeXd
eBDhZblGSCyKHzjFeLzk/jkVUJzrYaGnHoREEvS1Z41uyTP/qkITq8m1RZShBlmT
U56QVgvE9dl/L6pl2b3luKv77VdSQegLqhBTvlSw3FtRYieigzIGTlhvi9w58SfX
tEHz7VWyn+DXfext34P68UjFAneGhTag3KbNiURduELOEV9iTLp4P8r4IAoVGOVN
c5FO5RPtFPrdETS8E4swr+p4/eLICkSbAu7iddpT/6z1khXxv8xkLy7gDEr6Grqa
t3AuEDjuniGBE0xrhn3Ntw+9PDOfA14bUT0R230xwfmE7ipnmuuFmTLDlUrBYOlZ
xbHdZ7O2Yy4Kz5FkVz3v6Z3ZhAuxklnq3Tu/OcJLRZpmikEaCRAr5v/eKRt/PaIv
xVdGu/3AHNsNJXnckx01tBPJBTEYQVoC3MsLncZeijFbop34ASDjTmC7lZSOH+vu
9XSTB4SygvSNwr4CMxYK+UmF6mncnIB8SnFNxtehpiJkamLDlhpmITMPBxKgkUOQ
EvXidksh1ClGqBDhWkjKIrSiMe4jgAS4Yce+gqfIywFg085SnCKMiJq8vHuCU+yP
DVffDa/7VO9bOVf/BmbIwctLLE7VGMmQ6WLHB2/H8YPudIXxXdbJWPgt7rFwHdKk
q0QxxvGHjbmpoLPhbsrB4xXPy9eo1xzyhyFVFVKsz1fs9gJw8jzmdAsw5Ri1g0NG
7wbc6MSa10AikdxBAiUGyh+R+hPQUr47/8rqU//2oSq2kk6+s+c3tLPOIewn59qx
F8gWN41LBOxsGg3XmggX/vYpOrFxH4OVVwc0leABuKgVtRYjh/5oZ6yut+nY5D5e
0aJwZ4j0PVICTTUr2NGCUnA4tKHAW2yiTfPfIZv/Xuba7XRSXGEjFUwALakUP/MS
dosviLxQWmdiH0I+Eja8EQE0RNmjTfQKaQL/3nmzxUeL4NyZfor9914v+znZ+cH/
TNYgqtOqd3r+IZPGQxmBUUCZKbSr1R+U8fvdicVoIQl/HTwwz9x7zGHUz0QeoeMG
K1lSap0VifwoMlJWSZfqGA8v5YmgH8bzYiAuLP9CAVkrEMWQVw/qwg+QuBzURhk5
X3AQ2Pt3+lCsAgcM7q0CGvn6FRZ5ZGu3ssgPhF58RGv2fDwT1UyLeOR6HZluQNGo
MvYZ4RA8taA+f2FPh9GmMcs4w/SadU9UXJ/DPuPaFncKuqTCaG1yVlj/EsrmyQyT
QbDLRXw2QQ0xFSg7LBYwdU9ZtoiMPQdwqLaabBASPPXfe6rZ8YzvYQHapt1YF6en
AO9DaaEt5bZ+aDxJ9Ruxu15W1LyL4X7YY3jVpFwbYHFCrkpgc5VoMnAF3YRI1fAc
SlEFw0ZPeaut6cdIvCm34hs6hZtW9KgKEy6M2k6JZvpRoFvc1QjHz/OM3cdI2ukr
9ZGKitSbVbSheY+tPl2nlA3EIILOqYl3SSX/A8dlf/3pP813PRqBaR1mc+TNWv8s
TdRHbezue2IwDf5/cdUSk5aBS9FTvEZFGm8Ha0+Y2lwFVrauxPKaVcAf2cXV7EDP
yQixBkUC3N7gNz6uipqW5/EVPTIi7JgensGDc5MVnR7+581yneXTrGME2NQR9Ncn
PeItG3mnEVYoskaEwreOrZ1SaZNYJpkB+QRlV1HhHazqVCzGQgiIZXFCreA/Uyst
7wMEu9DJ9Mswt9TSyvm3Eb3ZOX3K7v5spKB5tXrodgKl25qXss/dj1DFY0TbMvim
MULY9ZHQFgNGO1KSEVaaLTP5Uip2+8uN/lldBlRc5qZMl/GgWBsthlcwBQoXm4K6
EZty4L/WtIuQFhFy90rPsto8O1ZYF0xlgtcoGV+yizYUC0DNkvTQg6rausimshUo
q8LFCu4pHFPmgs4URbdlm4bntDVXf+2C+K88S5adY6XMd2MI08KMiIelDCxaZFYO
vJ7YxWXCd5O374uLP0sj8Wdl7/mXuXlig50McHLdxn1AKsmT+CZpVEm13w+Yoqv2
4m3+Ll3wO9EeIZT9hWtlX1rTD2LDEkNM3eSTva0AHOeEFFQQXghhTsynnJeH41n7
86rGYEdod7URBwxoKz4kH5JtF+QRhWT4+USVffyj4S9Kro9lrguiyImuN/9eYm50
+oBJhnHNcYXRneOZVVEFPkOC4mLmKie8ePEVUc1fbXL4KfM/Gs/U9wT/EoldxfkO
L8QXXr9ImgyR+0BpkCnhhdUjWHdQN5l9oenOT18kePc/mjNFNNgAx8CT0xB2xkig
QkmjfLxoxLmJRh+kC0L3evq4aiqEUyoE6wAjtIT1gVzXQ2r6JXDr401t7aLovNur
5RIslOIadfczYVR+l4XqiRSq2VxEbU297if0BT4P/BjGjyqVLLUfc5FkdkJLUFqz
Q+DMFVX4jufS47K8iN8iXI1odwoovCEy2Ych4LEG3uPCs6PrtYodogYZW6BwL89r
OMHb3UfYMlAU+0MrFO72GYY4rAniabzstMrhuRgsoQXApJvxCI5oFejNtw+THnee
XksIDdscfT2MoBk5aCV8Mp+2t7UIG2LIv+H0+U9HsCgpJiNs2+6J+hLZEWV5X38c
jAWvWPtr4koxq2N76jgfJWcdPBPqQ+c2xMT+DJ4aZs9hFBfCHoCcg8hW9tB66Bod
GLN9OQlN64H8wC4IGoiERmja/JJVwOdKJ2K2fzdiUO05JAC54Qh3BWUM9AwPAeEn
xKlIcCmcufiyq0f1ZT8jf95GRi/+RQoSBVQFeRD3CQMw+GXgaf1WaQcC+vExtLU+
2H22YvrUXxFbqlKbVzRF4SE9rrC1wZanIptM+R5w9l4Amt9fR1Uotqap8BpX/22z
snFVmyXB4wfhiO3Z6AqvW1QrrEDTCEOaTDWVtNj4hvaGbTtJJVTiZlX9IcfETAwB
Ai2HlngHC+1H0l6teoEf5ymckxofrqtVervhmXXGGRibvPteyajCXUWAwdQidD0m
KxVT+kjtFMchnDUuzQ4nwBwdZsNGL/u0k4v1bsesg8CZtakEl2LwXRuzTeDJA7Z9
N1z9DLNyg8WCqKY/kiCJxKJIrgEvEkNnkBmFG265ROdxPki0WRbp7Xu/nLCGzFwr
/unHY81JZu+B7vDPlkw20wgPNzmUUU1CwAWXrdBdJZTwZnvvIPzQ32n3SOKKZM8X
QKzkdbli/7K/m1xN8CVCLo9I9vy9Po98eSnOHGbX5wko54yaVwezRq/yyWtueLVj
hXDC2yibjWr7Gbw3/t/ek7AuPckWLQ2JsZT8kPDx6kBKG1/Up1TGz5pkqO0l+zQ0
2rKyyKzXWz76feGGYJcvQaovNXbHLQ9UT0lpJboKg21IOsGzgHD785kzS7i2ff5f
t4MpBhicXueqg0tZSFvuSlaBO9ElLGEZR321kA1sAXj8nyxL95c9BQQlb+ypS3up
Bp/yNhn5xHoOxFNJ3JXjOw8VVJcebgNo6FcPZsOBxqeWJVr1thr2p+guv805LPRs
Clg/GrHc7/K6Cay2T0Vy++q8D+8hnqSEDO6nOT+zpxmnplYA0/5yWYxA3qgcV5zW
8ooRXKPhM47RMigoBDdPb9VBDVrN6efCBf5nNe0G6jD6iRC9xnPoz0d/q6Fz7VTM
ynqSlftSRxyzUY6hdNqle2lIXwpAulgIm+WFxv67+mSMbzttS8KcLKenf5DBo5Am
uo6i8uv76XOi8CWezml2C9KlGt5HyBvB8dsAKV3rraUTKjw8nZnRhIrGUx4dMU+y
8778dIqg+3XmfaJdnJ6AVDkf2M3UyaZzPpPVknt8ffkLwRsEm0K4m7bNMnQCA2bs
4cjxz7AoYDK1k9mhXLp03JFroNcXDHe5qwnM1PHmB1X9bg+XK6+iS9XzwOVszvco
mxWd2zAXbrZnHiMAL+521jb5KAz8pwZPT/z7akD1/IQXxFt8uY0WDiCw5uAPD42C
iM1R3cYB9p9XgTNofz+85TZkAC+/XEWHhjDmskJTYfNBVyI6sug5iQ0C5Fkbp1oi
UaCPLt+xb0Kda2fiLo2hszjF79/PweQPGQLIRpNqSLhn4yVaba6ExGGmvtxRWHYy
AhlrPL212t9FayLzojmLXu5/38el5ZC2xTGQd6gAqbZGjfY4f+UYNTLmShEWoW3B
WsZQ9Pyf/bZv1KSG6xnK3X+Io8SXfFB7lqSz3vJyUdlEjNtlWavcDdoraGMR2ch1
sgHDF5KolEVtjqnnSsCfZdPEGxr8XxDPgm+KbeYipvMAInyK/Cn8o1BlSODYXVIY
ZTzxMh7loH3l1vC1PFLzpCiOHCL/AZVxNnEN2p6bfnmTx+DggyQj9UXE7jFrdyaG
BEiH5wd7M2DhXZzkxojaDFULPs7qNuR6BcsT3lPSxREu2NUHDDl0GLglDBpj7/xh
38bKPjOJSly7whvV7FcvPJnov3n6Tjx8hbkMn4vB42WvwjaAkrQgaeg5cfMNMZtz
ZPaKnwvB4zpR3zjUcWXrKuUZJnSeHY4czLzBf45cRKl7GsH2DuGnneFl0f9ngtWz
jIxRkzdHH/z6w0lvUTYusph6knIIwa4yWWbV6oMH0/kKwXyjzZOUtAGCaRkHyUSR
1/+gV1g7l+EoFNK6PvQ/rD+Z0xUFHhW9ro/yLpNkqKPUWbX7Xtnlq84l5DPR8EoO
FWZUTGBRYGoeYqiVJu/iA0cvp94B63jOSbqda1XJOXZZ3S6ilGbEPyWcwBP6iexU
zy33h63Z3p7GgEb4+wBdQs8hk7bDnkFVll3GJXSXDEmT0rRHKpZL8x6T658xXrRT
OVwbQDrIAIrAPtipgf8S6QI7FqGIkTTA+8hCm3FOEvG3lagaxOjbK55KLcz7nrQw
UWmXCn2S553gSTEvmn0g89mHK+QdPfVF/JWXoZj/U1eRWrn+8a5BRCEf41/laBpt
IMlD6hEls2rQvpH3Kmcxra2J3CEFP3LJg6myZfsEhBgqxuXTS84JFF9fzuml0weN
jg4SRDJR5BkW/aXdLF0jDv1vu+o1EvinoPawNYORpxNNV8VAmuYbUAgnG8LL4uti
pVS1zl+lOXe9ANDMFkKNAOiiV+dFbFpyeWI5PID+JCejNYXc9ZKBMlFh6IeeHrG0
2bwj07SN1tF+AUKgicSnPRXA6tlXGO/FG6ubUSw48fGGSVo6hZohjxqbbwQgTzq6
ZNQ7I5pxj/CUUNN8QD4U0qUvZkMmiwb3gS7riGAkY572p80yl33gi9G9IajbXbFq
tMi3Zyy7+aFkVQs30PZLGYxsuhgO+9K2GscTnEqqY+Ja3j713HUq+HZgWgzisNpo
sFjHHT5A9S0W4AYJphIdVoDsEFjMPXLSfq6y5TKcR/4PSKZguTaNzAmTY5v16QFc
zWF6pTCk2/CA8BxSLMAjpFfspbYkk7XbA5STUt//I4V5gN4atBI7qsewEKXnzCYh
kJjSlUXjR/CQI1rW3XSjbIYE7LNMfo3IuSW4fdxUWA8UuuAuGFaIMuX4oCacI54A
8E5Qt1IArTlmyDDNLdEnL8bSR8rYTfKXDa5kZtGurzkXOSTbbOZHx1LCV4P/A43u
63VxowNmsWtmAGhMZtjNHZJc4XOUeSUD7Pjq3kP9NcnIzgmDEWKSonrQ7fqcMEVd
6uc9uBkAFPreBxAE9f5zgh/US65kvtCgiMKoWt1PFhGUUIZ0qMKMwcQP/TDYmhYY
PrvXEGdLktzSIj4hVMVCigelnDYaH1dfdU4heHCDHX12MUJNwHVPeWDA5Vu5fVCf
OVo7DZnmAauU55R1wLCfJpfb08UB22cE5HV2gccLs3gQDBXC0N3dciTYhuZzWYV9
qv0D8mIOF9jVpbWGox2Z5sPDqIqWMN1zWooGKPwaPYjsoDpiZASQYZuoa7Z8sIiB
rjhjntiPyCsUzIHukM/DeOOMixu81xe56Pw1yGM2r2EO36dXpztJ8fwx7zUwa65t
szSi4WVpsu9qbQ7AYCQIbjTpnt6Oo4/WrBjM1SvznNuHOzscNgdhij+pvDpUALUA
diHkqQstW8g7165Nximncu8nRtT9ozHTV9X+GfgvnvOGpACgdfvrJ2ybR1whdA5X
YY6xxZss9jsGfMhrUqyCDquIUlbg+JusfiIKCrr4AafcnjbkoCpCw7/a3d03SbDZ
2sw7Fa2VEWqjOLGeXiSHe3fqZqrpCL3JJOew5mgLp+LepsgtKp6VIE6Rz8h0Nw4L
R6UUTKkHpLxnkaOejm5MYUtqRSEEvX6lpHqcnOrM5qG79xZ+sb8HZqoB/MKTWj8z
pHTEtAGrjApIGApXKkbTCEZ3ZaXJBUlvp0hc6HgdLaIdeh6EDzMXkjkPfsmFKBl6
jIzkYwkV9ZPwmARhnNh7qTYHQs8uvy5xAWvDLgOzwGpOnRHAAja400PSnpSxQqXj
4Ljurs/gGK3X55RtjmndZDm9bjmYFr1qF1SmQSvjrPYTOsyiv85s+Gsx/rRmSdXC
Ni5CISDIFfvCpLTrN7QPeH2KQABb0UxlJUa3aZsGzcwLGa493Bz+eCbf1XC2tn9l
WS9d8aA4wul6dOFPLOt62bQtjEi0oALuBpLBTv6GEOeIyRkfYbvobXcAlIuhmR4p
Yf55Pe32mNL51XyzwNTR5PbFBCBeDuRyEJ6M2gnZgJlr8ixno4Z2AhisFoCLg0dK
x2e1Ka4BKVFAKrguzmylkh5szJhthoTWE2089l2Iqsnroz/rxWJg685JbLQ+Q1SA
s//WUfxFMB07+1cr2IEefjtqY00nxcfhxG3iIvA0JCbvMrxurRCCXm/W7qdG3n/v
TJVyPVZ98IvIr0gM1Wwt+mlRjI/K6TUqVVP8QOJynNP5dE+dsGODxEsyhbAsocWN
wJitxrVg0g9Cmb21PeXFxAXvmnTMsj8okWWXYcNEDLwsz7W9VONYGJ84vmQctpF+
0lQMU++zQl05BTllVuJ11kggBnpc3WsygCcINKFRDrsDH1brOgiTrBmFFHoX2own
Opcevts6U05gxAil6sYPyL4sMS6mxMA2mG9YfpzEd+QQ3Po5ZuBX2wiIzXpIk6eB
vFHulZ+FdazFlAjpCxzwsaJn0nbdhfvRhVGGFkvPltNY/tG2DidfBoHAHOsZ1BOU
jXyH8Ms/W0mjBJ/FmLgxqf0qEGxOscA4QgMK0Rc4bKBCHBMRCsX7kJPTs08uHKCY
D82PH9l/mF0y9AV4ToIL1R0GSqF8nfqtGW6K8ZmUsmS1qlQF9JBJXiUHjPeOJY+M
0wJ4aqyEBtJ+wO7xn8zdJCcJVSQAsUvn6bd0iTSYIVeOGlheVm6ZztKl4wX9MTWF
JQkkk37ceAPFgR+xWgiQOyhf6QIzw2qir7i/3/R/lEQKTD4msNtN+oOddvTr9Ysn
o4+j6A/BV8j6w6rk9hPuD1UESUbDUrl35L8kZxc4ruVmDJiTOGXz+ZX2x/CBx/G2
OgH1MPfcn4BjGwfghf4h20FUuQMqO4xjJN8MSX4+hL77NZbYOzVwGeWwG48STs3/
2xjBrzurttrdgvwcRbbDuaIk2PhTnyEawEztiBJWpuwHV4Z3mEjN0EunZBZDxcJX
75zVjvsBi39RPLjH6j3cTlvDDQw+lEoskAQm/qUDRQWrCiExAf4DCBsTOJcnicVS
PJz52Kgvd7T8tZHYu6WOly2c7bTrRLG4K+e/Y1NBQct28TK0Cq06cmiNmf2JC6Nv
HMgAqy5earChZggNko0ypspMFoHY9cRi7D593gCATySX088XhZykbLOdoL1FI+Qf
qCSXDRMB9rRJ+6VAEKdMJKMfDOov/3PZ13kz2UM5S3zX3zxLNUOnql7v+aNiQH1E
A32mM5D2NhVFc/ovN0CRv7RBHfNQYAIiQSqzc3if1ypzffuwXI9NqA6yjwcSK25i
IQuTv6haU/quUx6sbvDzb+TO8ZejCpkI+SfHBhJz3b/CrWMVw+WTi3NSiif72eQk
aRSKXcTrXQQTBaY2CvM809hxiTBj5F/VPzBoXGAX9RZbtHo4Da2x95tu/HvnjUcJ
/XwBuac+Fm39Xsq1vi1+u0eRCvmYJBn1NbAjYlFD5QpoLFwBY+9skkhZLwFfIAxO
fch5qO6mecVjutL8de22eCHWoF6fQ3AWSl7Md9IEPZ0q6+UMG4wIOFh9UYmxn4Wc
RMWJqqsVDVgcgDF/Y6/cRFprfoQpluK3EKlIiElAiwg8pGhN3aagTecfElwAeJpG
0Qx1aY8B+8fG1cRe7YTZ9wYIGc/0F2Png5BWvDKYNKUM6ULQQXv1SFIoGmLbixAz
5OuhpF33VzPwEvKW3UZzygOUncyReMEJfl89kMod0M3Xabl8qYvI3Eqv+6gLpYOK
w3Yu6+D+7lQ4xAzuJRPcYtgX6gdMQ4KA2bpTgGgpH2u1/C0JrGnt2WGTivIXQ5s8
Lne25r1MXWOY12Daj7dfNuZQenvk5SCTi8RtFSFoEhOdeBYoPTYPJH3A0oHRQN/l
Skmw6i6TOhEDJo86n3G0uFBmI8tgAn160QEiRHaEm1er0En5bjS8aghBhvEhEu6a
IWMociw6RrfVobTGGJT7ukMmCiSXn/TbftKDpz5F04C7B4YmSc2ip/kWGwdeohG7
/gfVqrWliIcaaJoN2yCQuG53Bpfh7khQMP2et1cVURdIXE66mXd8iMC/qIVrhsxy
qTMmVzM4ekIVpkCsnGuP88ZlhhAWQWJ/XriZb5w8Hbj6XVhSz093XoLUhw888eBA
hI7IV9OEoP7TDvVWwDmwOBliu8m9I7fWjbbC17Wsl2jqbb4tb0+aYqvBEOvrUhu7
T6u9IjUSNNXPgcldEcyhFMQhFjPjOswkRWoSiPT9uWqlTzktHJubq2ivrvNQleDg
qfx/LR6Id+MvxolSsM/bsJiVDRg3Q5FFzRQvLu75kZbJA3TOWikGP60WFEcJmZCG
Rb8LzRwylZXLyGkL5FgZCqANstKGKqEGsuSBbrdLSgA20VnNU7rDJ6HqMuKY1pj8
MjhuH6349olnuBGpN1rq1GESxJ3TLVdH/bBfsg9YykARCJO2ZrANpenob+I9hGha
MfNoXN+07wejj4/olooG7k2JVeJheg3USKlGEuTtwDQSZWPY5f7rWBffXYPjPGAd
vYwiToUfTiXqfjwHa/YCo/5oiUVXNg+E2gULHTs2utQEFqH8G/1sjCBBUUM8WdeA
opNjJPAv5bEEIGyj3dQpaKddwEAYaeUJsa+pjMZANH2ojrCMpssEBLmd3kAjC7u4
vSVWb7GE3zYP+wLiuBacqAXv/xEH7tgCf1PpeyI1TqvTUX45yMUbCvzvA9ttRAKS
OwsUkWHx5AP6+t77ZA2HRrEHcvwzod4kU38lwOTJQ3FfDtiMQJzkgMthMpakfWWT
7+pLvvLPj7dJOfdgy5gf36p+Rbhu5z4KZtOQuhemKthWZ5qKVR6IJNuJd/Q7Mn6/
D56cYw6MHZGxA26fc1ZsI9v2leIZr7dAJ6pY4WbBEjkw/APxiAyGo0fjP8/smOCi
dNyvLsiroBhuoUitE9ttCTXDEGor/NeOeXB2oU4NT6d/L4ECqZ3Tody6WFoSHs97
PQ0yPANbhNOjlZL99aeKCwb8d6emqKdW9P/RBLXmdWKTJsmsaebBPfbUBT/U4mz9
bCmcYdf13HTMLdb4jteeGj37SZ44or6LibAwPnJoBmAZIOG7sJaA7G37urwIrjeC
w1KVpG3+ffKIX4iOg3AtkRoo/PBMIaPB3OfzGJVUhPdIr2AO3PFYM6u6xbOB8sFa
s/O0/qtQMP13hfuy7ZxMqjX+HAGRwt7RgyYPqTJv2GmUSY8cZzXKAffNJN9DcbZ9
IlSwxGUkgxRmlSc1ldZF+Z1wsOtPua9ytO5rz2H7hdzh9CbLvGBcUg7MP/GuprCh
H50HMzq5cncJnWpznQrgPj0OiVGaMATGebiT+tPng+0TkHgSmcLgPeTUVYnilptG
mTZteMfGXxDajQHUIRXsbATHQ+xozqv1hFQaH2dGEESavHPaHOoRZ028/6y6Vxwz
iLoSAI77i+kNIcB1Wg8SSq0nJ01/M9aTEVXkxbecfNOxnhVEv51bIiwcuk0GVXJX
Dgo7UPT9ugHLQU+NKTC4jGTy9rEITq4Wqz0hZc0QqGeFJ4sVJYLISuof+PqIym/F
qt9hjjU61g9bz7HjjSyT1Bg36oqIC8z5dPi/x3fl51HHjFrxxriE0QI6wdXcCIOF
kII5rMWLYWhklV4AHy9XiWMSaB02VthPpWpZ+P13YXFTz6cloSEXk+S5MClc5VLq
lvxBBtlIVbBJo4lvZ7dXKo65fu1yEmmwWSLNGXRVGyRLdBCCwU5z2PL4cUtU/6YM
UKs4g7gXjWFLhBIAgs3dw+7bCz25MHy2EpFmPaRY3cvdcVRayK81HAtO1AFMItIf
nYKSUXaiyIOh4VnR0EfuUgjQ27lCkfxhtYkGDgrACIPzy1CbqXybDTJ6jP8gaw4X
Sit4KZn2jvsa6qmbLgmJ5dQ7zMtsnht9ZVYQwasibS36Wlx0XTmgochb6KJCxwpb
I21NL2adtRbrgmFvDl733Z6WWWjhs4GGIKtFd9g/KPoZnV05CgYOsYuMV75YiBud
5FgZK+pmSZAqjd6suy162aMkSIjTvMy2du1VnynokbvPHLCeFluL6IiXzLRU1Os7
hOKca5Gcu3J5q85G4WySkOYuej+eHY1Z7YEWyxoDSY27VritZ+MdtALHFsl6Cxvh
PvZ9g4KoCd/drW1EbtinxR8grojfFqBK0D/qinGAGUGwcWLJo6CtcTURISdtpRkQ
Yta+eWWm1V9Wkad1Nygj1UjnFtIYXXfdE9LJMDCNBJ2VtlKSajceDdKdii6eJDYH
PDlG6sw6r3N5BbwclsTXQ65gwSPoT5CDgX3WhnJE8zELDk0hTqI6Ekor+FIO9s36
yBHKwDFs4aWc4rQ/EcZzuGRKw4IiZz2RMpNvia1i1sf4AhHibr01FMxO4NmiGn4V
N8MQ2U7gdlM2HzevuH1eYAP5hmgmGONU/sBZuc2yYmGsuegl1hPNXN8e9pW5Xk17
9Zyv/SIeXSPv6K7vYpIjaH14zS8zXniIlKo7uzflhHlVjaTGTjUb+/mx2VJVMdR9
hXH64wYYtN+27Uu5QK7c/kTUZFzMwJyxRF32WQYw/Xxm6cXwF3ncKTtJlUchlwGj
HGbxejr1Nkb4kwfJr5clrnR1Mjla2po7U4V/0dT3nMI2LU7q16kt5MNIuanT4YTv
HBKEnDxUCvPLXf+4OiLKr7YaLE3YMfavWGkvmz1s1+l0lrij+Vq8isUB7DCgPbEc
lzFJONZk6Xu7z/Ke8zlJ//SvDAS6CY6lwY0DuZDmpA3/EM+2H87q2efjpmz38kKQ
f7gD/37i9YUHWQ/vKjKqXQONe6RQ3SudnC+4cIhyciSMib6gmfmXxhJ7LuV/haeK
Ok6c1XcXVJk/3cflKhcyKr9tRF1VDnFwXJrUl9dKIGfbIlWMcHJ/Yxn24GalNzYf
cKiTo9h8+nOvFGdlP0JlgfFrGxJzP1Cg9QBWjMtaCTXr7slyTOpJSDpBjNvT2g3T
yiy5TRSqkIU7leXVPDLbN36+UKxZti9EMNcwis7o7hkAuSU+AHGtN+wm9suM9+re
rbVP1Ea9kAivoDsWEoFP8wXQ96jfObrFY6pIlx3fQHVGz7dvOIag9LoCkJlEKvkb
E7gRLrGS/ysPokoxh3/pPgkGA6y9bqRyXod/ldwe5cKYyIFuIMPyHnK7F6Og2ref
1AddzuwE57IQjbMm9m8uchXY3WBT+7LlC6UYk5ZvCpf1ehnuQzNc4JEl2gJZ9TNa
DR1+Rf6aIxN+Ny6eA3f7TUaewTU98L4iYRdR3TDKKExmnEWlTnCJr4HnlMEfrBN5
Z6M4qJzInZ9RUAdR9iAjDSRVOC2scEagh3DOnlHKwiEuM0MXyZ3Ll+9Oq20z5sfW
dgc2RvPg3g/y+lFLy4DKsrdIVyvwQJZISnTntMh1wIerJbGh/x+Wq0Tx3p+QHP26
HoSchR+HL2xssHIfCDGUulvQb6oSrQ8Qznk/DGZM2JZj2W44JoSrRaxrViymsGrG
h+IWVLFq9XnbogdgjXKuGn0pD2s4A1bf/S4/0R86VsOQIqtcH+ixMT7wrmXgYJUF
3iBjkfNTZ4oU6zEJZCe+lS6o2ripYSxqPD6nML1JEvMVYUvCnmCcoz1v3D73vjKT
tDTD+uoogpj+qg/r6cjkFslMuWcDuME3sQ5JibatI0bl2v+mLG0NloCUxR3vCFG6
9ReY6fuUd4Z5WMnLmYfXOBUmGHKM8cM0DiKpzOgl8ZRvMjt5aJHH2092UxqOAK3H
crwsSDjD82wsOXFIhYHNtvYvfNH94U3hjpIY/OAuBrDOaus+d2UUWWsFsnkd3aaV
Ai+bBYHvmzw++Jq1J0EveNIisTAMrHPoOLiAUCDfLesD+mvoaFFNICKYLQWJI61k
KrM3Gl29/o6X5+VARJocJq9P76W2qWBVGd7d4bbbbh8yPnXL2J9k4EzRfQNPFW/H
qw4068gVkfPdcsQIOpLQob8jjHJQpOr9YcHFkytGVsCgg7p8exRPXF4Yzq8lVrP+
kQ2i4nAUbHUxR6+JCjaXMAHBk9DuI4MkfLr7QYeFbG8kC5xJKvvauY/klAhRCjlG
BkDHgv3rhl01fuHTaNWhRcivIOCSH8wyEhSYSEz1ptoyRFGh+IBP99eF8zLnKjE2
gjVWlX4FvFaCO+Lmp7RonIBStqGbSLbH/7DZ3KFUP76HCMrklVbMJ0Weq++6Lb+S
hsIPDu5hTuf6jObZ8Q8SsWA1Nagdb/hXQtDd9tf1kh/f/PnOmvm2F66B39vyO2F+
9Py6eLhOzQ5JYVZkoJOTyTSO8qRUWjnAS7i8th3y7JtwoyUk2Ur+PZ9qy7SXiIB0
Fqb5OmB73axNX2VDczOnwB+YN1AMylWaKPbsHawhvbCV/6XdFWHtxBdh0406/+mC
y41ztj5uldGhIDTkxxaVY48z5WxXF6AGttaTQ5IRnpw2cWZv/hNnJ5LhPp1vwMp+
OYwR/Ux6Dihu/leGWqe7wlI4EU6oX2RkCgo1FOsY/jzpqzFVukeHuVm3uNTGBzoF
Jcz7nSHEgVBAGjo3VtJR3/xbUlOPp/ERrPcqdY67cJms15OAgneQr1cxFZiMDDEN
7jf2ujFBKcRcVDojfVEFYQWd1zXbwEJ+N9RoeNxf9lILeUEcJdjisB+LUzhzSUG0
WxlJVg4H7UzbnqSY6uXUEkP7SukSTO1zz+YGdTcPJJ0lUxrII/4r4OK4KJEClrhQ
AxTzQbwgXhLJ2M6MCkmTYPID3m3oAFeLfCPXJJYQqLP9QuAZSRRcnK2QF8pANoiG
ZboDLttBuZK84oCmNwUI4KyDZKtuApQ8cxtXFL6Ws7FpYhj2foAgOPqGPoLeVcS1
2esu5pefioM8en7DDq6TA1vwz7lYXBEeENP/jlwTR56rEjUWxkPjRVWxbWKpQVeC
UMB7QvQKkt4emLvtBmBXPsfUl9g6ser16RG+uokNxrn/hdGptblwAoDUNJF7j0+K
5aj9iDDXUbSQERH6Im+lgYGDlSzc4nEUBXfgTHLMzEatBXgbIiCMdpH5Wz9TL+wj
5hMdyH5dQ9acuvWDHCqTBT+3LU5xxqw7pOxBaPX2XUYyw8kgTYnWtC1nbVPkomP2
k3CWgM5E1PJ+xHxhUAA4su6Q8WNIwPOc3QUDJmO+mQb4aHn7h2cBQMD5p6GvV+yr
rKwrH7ITqQwc6HaNVO1DeQ7ovvEQDS1YkVq30DNlBwIv3BitzUqzbpmzd+sTB1Aa
ptopwabSgLGLb9RSdeaeEycDoxdnUKAwWvXKUlRPIR7qQI5/0bvnffwXJCy+Xczo
gOC6VBbDYpii7VZNLkXeH7DWl6BpC3ou0jx+SIhvS137nE5DlQSUj2Uhf7aeATp/
TOF4RSGs1/8gvmaTkxwfgIlAIAY6HOh9iQuuhMRmVBvLE5nnfBm5JenaYGgNPX+8
u4wViwj1yQld3FmGU3RyHkgXNBk4eZw1VyGO11h5KZODBRlofwyXbJPcbS1fHnbP
mMYIsN9E6wlX2inbqIZ65CA8meD+cU7YCy5yY3GuPLusXbd4xwGZc4UMdTiV2gTM
gwz6vf/OUTR/WlXT+qtlb5ZuS79ZtMy6NFBen1MoCas5l+gqi+WX8t6GcAGCWuWS
5+xbi34wpgjkFbtZW4xlT/4dEgyn3ysAsieEJop1Js35z0erB8UIx+sp5j/2bUG/
EI5cYisvzO8rM/5+Fd3e0mhxc4Tq/LDsHCyCeRZb/qmEc3JcL1s3IhbtUGV6RCR3
zShA8qejfuxQpStrycYsRhaS2T+wDln1SXfYhdWKUG1865+jDbrOKpbhyH0H8SFB
kZAKTWGgP9QnON8yDzSszRRJ/lEJSCbllzgeHNtV5JyX+p9sDxVHosITukyNO9p1
M67Gyn72RDPGDenvFqvuAuSgdtJZHAs+WcXrrT0H4FjZU3D3TGwKdFGBEbbybLd2
sRQPdKHsdmvTVEDr+Cauf/Ag16ZDSE1eRgDXRVhl2TviCsCMPaYGIw2Llj1XvkH0
6UnQN5pWCkbW5f60oV423h1c/0D+lV3XtyDabumfyZ4hen5Hjs1flbjgfsHZvRLx
ivDcyR5L6wJ+qrSWaroUdHCsA4HQQQTmqByZLKMHxiuBwwqi6IrzSTFhe5rqjS0O
aWcqYQuHs7LXjmDrtJ6YeCbWIyOcqbFvc/RUT3XV02dPkbrslnaPwdjyncsf9vAY
4ZQyvWBC7xuqAXxMCB6GRvWU2fMTdKXFWhAcBOfgOJUPlKprdjrMYI0mUYjHmpGr
DA8pbYTgFGzoha1zW/0CJ+xHoMYiOImLno/t0MTsSEiaC4nxuurBTaeYSKdCb5et
0rVvOrmYIoDuhVCFGgcCutexE0D0wj/w9s0NJgxHTRJSNdykWmFcQYo3qGP5tOu/
p6Pfr1PgwCFx2DWkH0yIitheejD3pPz3lbxsgYrcCEfpJKpLKIj8Mg5+ctps/OT0
Ig583SpnBwDWcGfLrM0yCITTgUK7pamtL3F2zYVKXqxe3ADcCqP3ckqfZoO9oMXx
rPT6dET1wMFn9ii1dg+Hed4IGeR1bBwbojuSP5WfGrJPTmuS9jba1ooQQ/5CMfvi
qmxtIVhNkLdt+kQN1HFkcIrPyD4Am47GM8NsRYZQEWYGv6P6uhpF5YVUJ11vRWFe
C/xix2md4IiZdMYS+ny4IBiudMHyX00FqJ+dPztAENJIR7Eoyt1WpPY7GKPx7kCl
+bu51OHayjUzr9FzhdERKsoSx0+8H710bxLM7Q3E5hDipBki4M1XRV3wNLccDuzI
0JPrVfS4lTgCIMsJMta4wYMwxsbYUzjdyN91h9Pp+bqymclV2hfU4/KUY+seNckZ
4pp/Rpain4GbX2l7pxNTPYzP2M3PzlweDPsxLji5YRmzuW94qVn8il1cfyARekv1
y1RZQL4M5iLkLi7c5mueYPv7q0HUSUC1kdQQ1Kpk4rQIs9D7HNrgsNrQ38CbBq1h
9k82KV2bpvz386vQ+8mQ5aC1yYPlO8IyvYIi/PBU/5C6ptY8ibl7beQ+W+QU/n1O
TMBQvU2Tn6b3/vRrLT1e/onxfNkd+x7tlWi1iy7VT0bMvHlyA6Mc6fx7ArNdX1Ae
XjNiuMPJOhUxFySWduKzIun2LjL36ykz4KhnoDDHEu/HCMKcSl7XeLjSpg4AJ7T6
uWH3jxCn3ptHFQ6xDOZ2uST8XVEgDvdzzJJXCHn1NMl3cprrltuookcoQ0bK4q9W
wmAFiOmRyyceKwSTD+HZQ7HqqPn6CNtX0mu8cSrq26ihb7VEGeNfbEtz2/7sMfoM
Gwsyz4GQFQsE2lDrumngYJqzuxvI/nNvgQNUKXi9Qehv7qbWzZnRoUVdxjxCurQE
pqqEav8ViTt1h7PGaFCypUv5GXceUledsECdDMG6f42jGLYlirK3a7Nh1e0dSRMJ
XWDSF+R6YSEY4D79aAOFz81eFlL78rS0b4Tugvu+wNobER3ZA3g3ZTZdrie37iiH
5eKZzJILLCXZ3ONQ9F5CToER2r8pMUx9/ehsu2lzN/ejbpzevdcOmz2d92mjpfVY
bq5TAJGwJsScWA2PP38U/vibZx9Qgn6mQkQX9SNXsK2cy2fXnsIm1ljym6k4PoXR
ud10PJ7KnQt9pyMUKlDqKi7pI06HftRMB/L59/xfVaDwtSh1I2wKqBrA+h5MtZLL
ld4+VZEKS+EoEqsUjxbCGa7kXR/dYsybvRptSGfSxJBRZdu5X1ACsuQBTGOtDpY8
SVhRnRupT31oC74u6+BYJOd01ezeZxwPvD71rcc4lIlML4P1HxLbfqKxzHoef4ky
DZElUh6mocmrbpXxHtqbONcUa5ukExFgVYX20JVXVuZLWLFEx1FG8Oe+BCeBwegV
Y9ssQAoEx6TAXdxfkHNLIQoo27Bv1Zpyy7dA7qKPMoLjlkEhff2MikgQOceT0Bos
CMGggH4mJYhGy917EmQU6GjeHz2zrvhAxmrCwP3Gww+sasNAtz2rxAr8/spu2SFD
AoaDwvq2ocO9SBuMM8jAgTYI9cJ1QGZcv1vFg7K4lzoXFWkH0bMyqbJmSyhBp8xL
ZphFltCXvSRXaasvn5UlE+UiKwS3L1zQvKz/xaznPYIttTppAHtfweN8L6ORMlhc
oPga6dwaW8KG/ZD9sUqajrvOdeK0VzB5ATpVRE+xO4yjUdvhUmSJOAujvOm3U8hJ
3cREX8qwhE/vsWB7NmZ0/Rf3fK1w9Wam4TCdWK/egbQE+g8xujKhdWd7X7PvXkT4
fdq/BQZKJPyCzvmmwbk6lS+8fQxHcIlEOghQH/kl6uUF1UynrkIEmiC+cwqy+6cK
O5PxF22NhioI42wHRvJfKSWm2AQ6cufVamyMVyOqmgmMkg7ejQE2NlK0/Btn2gIt
6Ahh/i1+EeXEMlSDewcbBh8IBvaf0J7ZgPIlaKnnZqF3munV8A+8YVAMj/P6/cLc
Wz4DF2Z6sqQeqjSC0zLz737wGwwMxqk4hYAC9WavhV0pJQaN8ihXfwFdBiqk2AWH
UmLfzVURf9TasKCaitlq4IxZskZdywmZQWVmJXuu0+RUVJ0QYpsKyK+txJNdo2rf
wGChwXBZSYZKzOzDMXNmXZX23+WHJseOPhrmO4vpvNJ5RKGOcej39HNJCZWWohwB
LCbIu/mW4WHgxgDIhobah017VcS4D+eER6w3M3Zt9ZeSKGsCrH6JXuMGlOU9v/qL
0bdSErkNy8mOaucTy/DFviOk3J54+IlkULBDuCHMC4AB42ddxT2+Oi9t0HFuzHpO
jV8Hl7moF+52IFdxZ5QMkm+zkhGYrVgReagos/uMg+jLrRfHjbtR3PGnUXnIAuSs
z8CMCk+T4c2+3UVvlG6REf34dwFP4v1LJnU15JY8JG5yduhXZNblgAuGKW20Jcou
A/wjnvUQKrMx+vyHnjHH+MD41P+daMtl99pf3TgV5guDyevKXnZmaPaC1hYDDJuU
hf+AmxMjAPBSjGeZzRYxt2hrKw19JIYVLEsXzxueShNM00ZGRJ9nChjXCbAYGwkz
AfeUUo5vjgDM+dVpXVaBpm/CcdYFuAQUdAXWxKw2Btqtr7k4yP3KTYhOJpO3g8OG
21JJh40Lv2d1ER4oV5zZGBpOtqyQg7FchyVejaCOSVMaxVvjszQtYEVAn4EmEYon
Vbv/PfxpBXP6gDTIaGtzjd1Zx1Ucnon0zjTg8u19L9l4FhiAc+9uVdZIZtVvjUMV
8cTrEfSfte5Rtc2j/JRwqdTiJgC2f33CNV7DrkA0uF8n6QJbUr3FwLhO38gS6or3
fliw9r26KKBcBYsRmUdEPXRn85HnaLhQ/BUlF3Td1UIMj/53KQ3vfji6zdrAsp/G
4PCLbOHZ9VDzfGyPSs04wUraqg59NCmEeygyUpJm6E5P17mLJaYCgrV2VmWDE0Cq
oe6fo50+lBrDIdJczAGpQwjrswl04yvP3Oa1MwbRQFdWbuXvYbjaEYlma9B+MbcT
J7uiUFX8TRE39v2ZG8NbEg/gQZS/CXlsqMLRF3pJsOd82J47ag/WWJo63gazkSLk
JjufgzPaWYQ+G+wW6Nq7FUWJbpxiz5j+8HOzNaQMuejv4NYnmUem3Qfvcc/1oEo9
IXehYizQgQV7gVCbzGE2qiHg4rQI0De0J28jldsfdjF5FsZ+b1GAD7dQDIukYq1r
64oTu+ubCEQqmfRjsFAlQ8eAbiwhY+I72ilgsfQizBH5yKWb957AzzQJLJLYKRtX
MuiW0CNtZICdBmi0Y2CCT/bu1uZOash0wZWtexwrmlxLFkQDApaHWH7jiZLJFCEE
ymDxJPF83hxs69r5F/LbnNER37BRlolgfh8jbwiwkwswLk1jHw2OCe9JfE4gewPW
0Gz+nRMdtVgoZg0SF+c1qnlEUlTX2LM4xeVFsieKfY1Sx4rI+YLwFGegJvigMuv6
NPuWUGWYPElGFwsX/9hQ8M/vFdJ3FckWs9V+W3G+dN1PlU41K7W2yqPzxAZ0p6Fx
+S06Xm00mN7omGgeHiP95+wi2G5RYZyMPdjfrHE6VIESpUL4tn4CU2Bsqp6io3Ra
3rtg2rzqvV6O4mpfJ4Uwx3Fl7S330u0iD8zsRnLynwIdjj+KC/XAdc8Gw7QaQ5GG
S3RHIkwBZCHW3rcN5gxLNLlTysnz/qPcozgFx8XgzIDTPjqWXT1V/37r2FNlBMSV
CKu5dk7UKq84R1qurIwSfWLf1Ixjvu9pLwKi/mDq+3H81OvYBfH2c/E7M+iMXTCv
mOwUXCGbEdoquC4NWyqCRvuZ05D/4D8S2hK7XIxQKX8hgM2e3MoXNU02o5RFTEDk
AfxUsGs65rxq41NptraUtypKtsLGmghv2eOEC+S0pDW6bWDiN8z9NzsOi3NOFJaW
5fdtDMlj/dIyA4coneHf9bI0cxQ0LarsIxqeTvchMgwT6aY98SXHA5KlOxalQb+O
ptTN1MkWfzM/YQaSW1UymR73nqwwfgGCII+nHJTbLvdP5psq2OcqcZ+Tz4Kz5G6M
fNAbO571W1lAZ4mGEe0USCVietYxFfRacHL72wJU0q3OVi3a6z1wj8zTci9HLHYW
k7kmJMU30tkUJtKOePuAD4OHO7TwerSILM8f1BPGWtKdrXMLg0oFhsMAIhR7YlJc
IhMJgwJp0HNbeNyJwa2xGaT/+MDFMiLb8dPdMd8fpVdbNg2UTVN5cjQEgJzQ6uJW
elEKdUkMJa/LaOfeSDAWCmB8YGe5+lIOqiXuPqpkJQ58TcmKrUDl9LT9EoMuL+AN
zPuezUt/rr7AN0fr4LyqxQo9xBfcvvO9KRHxYYNfG7Sma6FBZjoXAG2ijfSuG3X1
q62Xt1u91Q+q1J6e+oJOBtIeonjYKPq76OU3MNqz5NtpUCwLzVGirBRiuQdKsyS9
63n+j7E3HpblOiJxkmmfBJKNSJ6rUOA89E+205bDm9VgoK+7zdWgRt0hHGWAB6Zh
w/mMvOukNV+AwIQNCZHtB8wLMki/+OuItw6mBTwkqhD38rO1OJU4mrA552IXqk2U
R/cbvIhlLPUnShRtFSlZkA3gVXQXpLbLCfduho3L8tqXzgbMcJ6I8eCh010A9wvE
iqZGQvgAzzRkfOSYU5FQGZaotAuffd93sO7/gd8qbA+Q4TcIWUfWkmxbeVv+h5zE
lAm6yMT8My+QQ7BSx9meWWBkGsTCc0npuaICXES8H0vCPhVAZaOgym8tstZE28IP
cJYOO4Qgh+igRXLaQQ0yI3k4joaDsuXGdw5xNvudyis/+s+D5N6RpkbWrJgrN+vM
Z573O7h+Q7+30s3RH1OQ1v2kT1aWhqOGFUIfyFG06hNJtNTB6XYgX/8hCglEsypG
y6xCllaAfG6GlJkVkqgVYl5kJpZtU/7AebzkQw9uTUvweF4UPk+MaFgyDwrYbhzx
0aeTgxCIxVXx/cI4VbrastXGvJP/N1GxQwquOb7qZ2+8HyoNRi17DkFIy/ito3yn
Vgamh/zpEnXaD8NE3/jlgeofwwe0NhvueJwb8996MoNu7l7/S7C40LnwBAESdez+
amxi77/QntgzoDEy5baHjufjJU7b8yjKl3zDR5/XnG9L9QDQrnB1fYg7uVY6h2Jo
yxtm8EvY7VAFDZa0lTPE8AtDtp15dQZkykix27cPP3qBCxKOl/iMKQbUqJteDPuB
lfWevdSkXBnfJ6+OPoHCtlbHERz4taVeU85YBGmba42fdF/wGpdsPLCMjzybazan
fFeSwXKm1qshKg4GNK9Now0NG1KS0BViDBgFc1RTgDPf00X9s8tUWxgtr4ebNBmU
IXejo6/1yRSX1DeMEwiV6Tjnt68cuAJmhc4IxcI5iT+AnNrtBVdR+YQKptw6gbU8
gaCPZ6XbhFptrO5lmoe6vVmBI7epNk2ez7gi3V2mdEraQz+r+BST3IOcNLt4V5c8
2v1ZQh66QyhRvA23hhRXgv6GzLylNs/L+onL/q2lMnhARUV+Qv/FaLpubYRxd3/i
6A/TnZG46iwcwISx/AyEtJCHUggnhZgJvWhW/APn+CSMu9xEWNqyThdodJ6VJORb
bklJoJeclublTQ5QUfO/PGo0PDXVK0+NtvublXPXWIltO9X0nI3Z4kebARDo2Lk8
w4DjZD3dxiF2CXThOnEVdARnFkzBmju+g+WBMRz0Z1Q8cULVuBM7TVHaAa7JRXEe
6XWRPocT9LMNVKLPOUHKOo1VcT1ztcCNRpVVcTWMLZPYo7pNo5AlW++Liah8Qxhx
FXiANEfNM5Afq+6UD8YP6LX/q4E8svY6enGGqsFFk/5TZY6iwzQwMPfdLCVgCwu1
kkW8twcxQp8bGnxQFKAbjScQ0iu/9/SG8cwRETmzoqlSpKV/3aunPg+Zs89o5eu1
aQ4gh6RBqQe9X2rb7tAEbrEmM1F93ucTSeuqHdnnNzAMCWBtctr2PeQP/bteFGJu
oEHThMsM7S8eAmfKuLhzYFhs0fbfXl+Sj/1AJ66BWdY45IHcCScSKsBg3gOYEyJn
uIV2VYmIM3PdtImIeewWeWhX2Pm2+5FVyxLKLms8/xnDhTqi0h1SP+Zf1DPc0AxN
cHQUxZwzBR1renz3pz2SR/WF16jIphsWaRi20H9Jieym4z9mSZ36hbUkoSS2oei8
vOyZzHIhbHowZM3aQT4WLePPHaW+ImiRmMAOi9LOHPeqp/OPc3M6LdhuhBLdwe8u
8nNFrdtI2ViGwk5gUTBnh3uXe5dLPESP9IndVsqTPy+df5qWK2y/kOM83XjdXrzO
FKd3NCaOvL8X3A5TjJd7R/V61CNwVtjW1XF5iOvOdiveKbjA3Shx1+wHt0lvP7ku
IkO+mKDxheEYucVzwwmktLgQ+FCPMPi3LfLrpqlVh/momUBaoBNrjln06M6E0ZjS
vY7AvQdtw96s2UztmJck5c2ZC+cugw+s3jVN001qJaLtzMoZ1l1G/7uGD/qySB5i
q9neasuJvj01UHJAShLwfv75dFDSMBLq2ckKDnGsAxJ8pUl38hL9/MOhb2Y16ahr
Q2fBNafjt1QoFXsaeGYoYVPpB7sPVaI6K8c7mp5qVFphwZ7m7XfGdEZOFGhC6t5O
T+R+VF+UwNFnKIXp1Aj7DTdvHMAPO7hTy185eJ6dYb+qxbTaTMj4d24Tc6ySRpzk
aqyRs4siVQ98cDu0jN6nK0UKa7nnQRa8wehGaf54/9U6n9T+9/zSg7YqhtIl8yKI
CB430M0Dc6w7EDsMFueBEFsUVppDxTOyRhKiuqMgwWnuYeKUHJsQ5gFfvH/xBjdx
lFyK7vkzUb/cRWarZmij8eS0oCLb/eEsH3C9tx0agAy3WB8eHky0c21lhqCLuLWp
vLHBiyrpZwqKA+M64U2Nw70tXHCgpfYzhnmUEYzjRsdxRoZdhujHfCvWQ0YZRJOd
/CVPy+9ZFlwdfxBhEPG3CO+YTVaYu6YcRDpQY5yqT9M0Ar7hNflMONIPqyjw10Fp
mXnKojz3cRnc9HgUFLt7iR3jKwkW6BOo622iniMes2vGYlRWqsduSQKm62f4ctTL
npOrG9GTs9u02Sq9cSESBr8YB6rUpeuH/nN0b8b6qCENaEy5hSsLbPz3c5V3D4U7
4AzwHgqr2VV1MH655+M3/9TXtpnn1SqpXCPWjRjfE46ndpC+6fLSuPh4bFOcmqPU
kYn051LMLF0fwNK6cGgxSRqzkVaGwNc4CdMRNSf17D3nCmIXioTOGIo/kfOyozRN
fgjlpxZQF7ibQ6UpxBLNPDYk3Ty8rK5ozk7wPmnHhdlv52v7qOyAQKdBYgiSVfO2
Wl25IzKREHugfb5t8nqrhChaliUAAd9of07KR/1x4ZFDoK58tGg+o0O0csjNcBJE
nSdwPC9fxI4IaPhBz5G29CG6lVnkVshkCN6bd9OqeI0H/4mLyvgEw/x8cYW26HAL
PQmiy/nCjLHW6tarPQfokM1XMCEkUBbFmfa7nRTYvJDU2/UMR8N/ri6BHn437fOz
0MIFTprBfL9fCKJLd6ro8B/1DYgqOqmZ4F8ZThU8lnLNVXbN7lZtXJrBCtJfkOUg
TnSTD31kJDbDnZShs9lqYS2QjsPJbBgvPFRdv+LVT+E46ezrnKd92C1YrOrnmPBs
ntLL/Z6zNt8RRHQTyAT2QHI/q2QpPhMwdm5NAa/ya/t7j9dTf4J+Gsn8PdbcDvLH
ha/mAd4Bmply1Y0EIvM0lxveQbIluXn/9MS2NCTwNio8QiGIIcYpU9wzxFDN8ZH8
iZer1mJDDIiND6n8XVrZVXmaSoOWqBIIpYWsBvPC7e1DTkQYTNq53oIes6JRuvXs
tCKcXoSy1+TofWEw43cjlGEoPkw/LuTPAgj98TrNuu5F/vsTygYroG3BOCshc4at
anPQa3JUUtQrqOitMB6C1bz55BzPz3tDpLLV8VOWzZMzuwvUyhhBishzsoUfb0+P
pmPFrEZSloPFfrzcyWvYTI7fslQoPqp3x4WDKLe3kAO47HSbivsQkad3wvVa31rg
5IwGjnlCEIak/lx7yh7yGntk0EHMglyLBHzt/9o9gBr5i4wrZJxuFsT+nqW5SFPY
WoylAClFRvMUMzSw9EiN5KVNCxqVtJ1grFLptLzTr+dbUDIFnzmwYShiANpyQdAf
cPIxpKIkPi/YhTa2q9Kr9qvugFHWxmOwYvmAfEdVmCLDN8HS+0WyqTpOcDVh6UxZ
Tl+6YcYIqU5YrqHQpTR0S6J/Y70ACVrhRL2kVZU/eufiGshfgPpA/Jim3GGAOa6Y
ZMgN6lcKZDSE+xIrRULtDYW6ygKYs2pszI/mM4dVvaw934I8HlQJHP80kL79tFrS
2JNHkeHKnY7UCw+9TCTXeoiDuV/QUT7VJVhVkqnyOfd9dbrQ+wmjsB0f3yYdR+sF
CEDSK0wu//GIZrWsiBGN3YlLNFT+EptzvqbDzDjz4KpooScUOfTBxYeyyCJCPk9f
8v4SpROY0CknAsbgRrUejtb06XPsLWD51TH5nCVzQDaOA8bKO/xLtxYeW/joN73u
p2VNknsjhRQ+RE1u50+6+IH0f4q2M6ct8UxGlyHzGqKqx8e9vtVDsRS+TUlk8iob
zpo5GrKJscRO6j+6/fMjCxqbjSMWOw6Tr60vbDD9102qLR+vOs2gitrmofiMSm5T
X5vOCiYM6A+UHWvdwrGiw7lOBsOYc56oatrzqSAdinS1dPDzjnm/3PIQlYBFqZ6B
GOyatZLGzPDmLuT5dtDiJzuu3vOP11P4kfOmlCKp3/o1J4y77CMOers06pXMVPhL
nq9uCPl7qUc0+RxYqxMA202mcsfj7+HN3OUzzWpI4GJitsukP+/cGC+eSU5GWzfm
U7D0XwnEVy1VO0CsqlbA8CNX6LFvTAsvKGw2h6g1maxqBxE3B83+Kc+goVAnSw/i
A+PSa4fc9TEdIWEIGhOYJ+96+kDC4IG31+SZVktqYLK/2LLy3h9AGiRPCNi6jU9q
HKT1ANz8VNb3xJW+ExM81i/0MOgQw8lqegbD/d5n7Kf5FbAwztLIdjWC0KcSOnju
BesMGBNcU7WQS6OYwkWx9n5EuJND3LcErB29qNh8/0E2/oPrZHjH2eFPdkpzdDzt
YEJgJ4Fl68Lkk5piGe1q+Jq7iC93lUsR6LM2v7BRcT+EELPieeL5S0NRdfd4A5lP
w99ZCNC/2ZIGGZbkIyZa+wsLaVP9N9x24/X6wQBAsYgCKmrmtqTqrAgUap/f2TiI
EQgupRBrY8EfwfxYKd9tZEU8Znu1QU23IJFrQ4jxjDhDrlAFyg/d7Nr1L2sHrY2o
eT1pweoS4vOYBuPS9up9H2Qh87UU5YFhtEFG6CBvHJmS2Z9F9DT8PtDqT6CW30RL
fUOct+4Mg66E1K23b7XibqthbLrXj5kP7t5L92eVZ6/5n2eZa2gIzkSpxXlzcPf8
KgDi5eCMC3uDMnjPtzGYL1l4G+MPAl6rKCY+6Utcv5C/939OAZgDGO3Fm2er2PaB
6bqajoHZAboCSroQhUnfu1dJ0tl0g4a4A0Zb2W5Hg7D8qduL4Su5W2supbbfHj8z
/GFHuVKyMiV3PS5h2eHCtaZ+Lg5XcqiiJUqVeZPcoRmbGcSsfciRCHHvZuos+ZrE
re9lOu2m2JP1eiqlxBfn4bCUEEUme+uZvVPL+MEvSnk4AjW3vglVYuIqI1eAitGY
08G5RtZcUNxTlYkxPxk+WV1XJg7pmFEQ4RkgTV07WYIhuYnP61PzIA7OtVvlBdra
CbRe+d/6zoloy03+gmhdEGSQJ1BcN7eKE3XFCCm8fJF2h2fkB1Bt6Hv9RUzTVmup
G0he5IgxBYB2v37GABcd4THuXFc1DAnuSLyVJRol91h9v1jNv6frr61eXt+l0/CH
JIlfbGBmfknEFShvCJ6PMLsdTWSOwR72vpwqc/kr2eD/EtU8+9mAA7BIqDQiO6y0
DXver78cHGH1e+1EbiJLR8DwoHUeGuzsUJZj99q24AWVm+zumK/W0lMkOATsmuMl
LA7TUBbGRKTnbreco+yFceJMsJScAF0JeraZpT3toXHiXGR07ZONN4ZPL8kBJ0Oi
ul/YmuwmM7B24EPIJNzGduHHlohvIkSlehC0xZpprtRPkYN1RHieHmv9iiJUbljZ
QGrfheXPxocdmhyxw6iB8o3NdR0RJoLS46Ol2yX/L39SShQTBeqpJ42L6SZqo8Ol
jedmis0nuoXs3pnuy5wWIKvpdwt2j0mMYfDccT4w12MFQlvSLukmOSSx4X2ZsNSX
evqlN7haHafJKLWI7PF27soa6246iL/nG4aN9HadPfmNd2ldO5dF/QACfx3xp/R2
bWnQSS+8V+1ASdpW1DGYLywGO0BAsC2GmWViwTFPUTafQGQbAMCxVKtUFiVLZJCR
kSXW9YoOqPqfwSWXhHCJoc2qaJd67EHg7EoN5L99e7UTahMPaJOsG1wd99KE5AmU
sXcDou9zjeQp69Y4/O/VMlbjdHQJTX/GbXFOL0OvtZySOuV3mITMpJAVpcwyXi/X
3WUhXRP2oq+yFCZ/JsneIzlZHanqfPx45+iYMkDJ5oaNGJUWFFXnfyrGugTlD5NO
uyiOmVs2smUWbzYfSg8D9lrxOSktR8NVeUcvseI30vTxo/MEf0a2Sy5Nnts2kODI
zW6mraoIeGO2vmqh8qZab5j/lsFdXCafUKsZajtMPFoYSfUyLdWJ69Iog9lN2MPa
TXy6+56Eh4C9kGLeNjYfQkzHeNDjzX5BymSEDeJoEPHIyO81OzcgaUDkuRPN4qqv
PLHu5Q66jxoYlP2jZmUA4h7uquRbBWuvIT5UuaNJYE+wXzvjeKZ8AUVrjjU5dQw3
c61c0Srz1hnCTMWRnrlNi1nqQuZdiR2xrxBnExjn8h36npH091DMWbI9gr3wT0m+
CwjKheLYEHoGgTFq0kBgR+KUZe5WL+rdWi2mAsebXW/Et1M80yH+6gFW8MDGhFYx
NbkCp2xE5Mcabn0c4tn70hkK3OV8xUxLxzsG0nqzZkFY2+HhvPFTIPMK3TekUfsS
Ml0zFJrmRe1urkLIjZyZKN+QyZXeK1qUE5lR3LIqld5mVwomPzB7Q6yjyL9tbDNE
g3CkbLWOpKUgqUMW+3rVdNA8jNQ3dQMVYYe+qW7G34tN0uh/5QVN5zCAD8El4Joz
8aVznGJs7w3bONv+9lcOHzB/VeHnr4mx2biW4nlm9tTQuClx77vWDCbddjKezysc
ReUcX4VzKvazS/sfUdUA0ebuIjoH4Z2SrtivHa7yDvr/GlvuHGNCmcF7tEEFx1jf
1GLbo7AXWYvUcXvbvgA5r1Qvg+71/OYt6/NM18rW/+dAOU+ErcJhskaKXO4YD7xv
G0bTAXnjo1qno50oCgVpZrWEHKVT9gTkRl8VnrvEq8uSEw3sO6O0vFabgNYApSuv
KCU4G6PUbWD4IJkPl+6hpky0f+oa5XyEOtwhGj/+9VKdkftZPWJxDB08sq88fV5y
9toznh7qXIsQS5zrv4REHFsK2Zvq4McxJKO6ZVKegg89N3d1V+PxXKdsoAm3igvU
urYWkcSrP1j2UHo76DMD+8bddKbBLYNIj4rFGogrmAsAx41E2weVLuUzAWw30E/q
bfaqP6qllw/JO/Uh/iryhJZ9BAFYbF5zXH/QTp5BAQ3vazIdMpaC+64GELscsXDs
vpqQBugKQEsMHy2mJOqoksbjTs4OfsW9W19jLuTh1PzCpyx7hf/SzZWjBNnOjKDS
zrnPtkYaj4LmuHL3/SyOyvjjJklNMH7bd/hlCu96iKcSvcgCgg4H60EJb73Op0EI
o/VOilM9wnviZiHpQ0TyxJ5/B8EYsEHDGbs24mvFvnm5W2lYAnL4PvK8hhjVPZfo
fi0mL2al9EYrKoJSdOmVS5HO0GwWKpA2ZDe9ju7qfUfm7IPi/eLPuMDNULIJF7EV
b/RucaiETMZDJov4DrSN+DfRtTSvF3IWRiclpaJiOlcxmDPH1V4Z34H5PMGkvChM
dOYgfp4NBs/8dfXCZUrx/lkEvXZuN5X5Lo4/eOq57zeTG1syEE16DoPlPOq17pFU
puKaU177f5QhLUzSDSFoWRPjBPhkLqU80wVONS/YdkSbuyhu+QYtwSwOZJslPQWL
2qdFXHQrX8FFOkMiO0yq+wdw2e0h5A/pO1CAS8pN+qKoalC6276cocNA+/TSE9Ae
hZrDar57P9nKbAqxh1+n9das+gueuSuikMtLjXHKpmht8+BGKOPp0b0quCPYeKGt
YtPkqwsYNSHZ1uQmiX7I9nIOF8mlSBXT77GcpgUzvKsOxIZkYYoJIQWneAv0sw4x
c89s2Bn4gsTRdWtuZXbdbAxc1i5FCsJ9NuqM6KYZmXqZTg0a82Gg9XckRYW6wtUa
3D3A1hJlluud6tXih/SPf3K3t4oHWxdO7vJH/AXMciySBapaA8b5HaqceHp58yyj
gMH+NZLjMsNJlVXf9XhYyMdyxw5Ad/GIENSlR1nwTl+Peub6HgRUornZ/X63r4Xm
3sLg3Ilre3t95B8woEI9k/vB7jE92tZMREfXrM80UoBgTbY7moph/nAdC3b++9sg
F2wXhTiEOhg+wP5INkbI+183ExXZSj5atds4JkI5Ivsi9FwTGnKWZX10/dI4ecEo
oR1ozrZvz4MLi/Go25028q+BSvJP5NI57vflPZmtxeROhz/k/MI3k1m9Tgqze/FV
yLytzfwebROi+Zx2z8A4Z3WEio322awmYmg3CV5niq0G7gVHjYSVpXaff30m9tsx
asv6ldmNKcNhkJHEMljdOFva/A3DeTgEOtDsR+y/fANrTccwBvAqp/bylHs3Nu7M
vIgepoY0p9Mhi76xkBQBi902eoMYhppXHgzihlNKpjLlqwr4NEzzyOD3G4e7jKQZ
OvmZQDHDZArHf8MXEiDVQz5l+21yft8ydNEhLsHmkKvTFu3QkMtrIGSojvJMGQCs
Z6tzLz9YJ2D6x4t0DaGjUnlfXKlA+NDGolVyn1Ca5VbUIG8KZlpWcSxMSzjd6tpF
CeXkX3t3RRxvisWU9iecQkdPUMCkJ3sfKhiEpbn+/m5nPOFOCRXcINewjY/eN6dv
bQT2zrGA5C+c+uLXyckzPOEPzUPbAof3vKE/8lsxcitbD8Gu5z8NmOFBszultCmc
/Nn39WRT3gstv3/rKnHNGTsXYsrTlQS8c5alc8SSYfXJWkgj29nPebIAuTexdxmV
jN6JaF7IhR3FB2fwUy/3sOwpgwfuwWY3f+7fo9oovNvuxCOcTAJfDup+EFLNsF5f
1IvgvDPRCgJCUe5z4GAKc5Rafr3H8Pl6HSmtGFikqKgJPRgon+xMP7Krnwkhcemv
4d572AHipR4sN09xx0GqaDU5zBFSvO5PK19LRmWZ6luKibPQYj4bEt8H49DHSDs1
EtvHx7EKtBzSHEl4XcBn5QxKYbG7zn+L8S7phq0WCMfZm0iBzSh5UAr3wcOp7V6P
MPGmpwYkmrmY+8+SbMLJjdKfRxWREm7DvEAgAKfAB2yYsHxZCLZZKfx8/5NcgAhu
rmEVP3sLru9ert0TNRU9ixM8Fq6TTLkuSKAx0PsLtM0E8Bn+8IusmpnnwMAeJUE2
r2QWGLeOAKyoD160JM7SQmiYurr+nwph847X4VtQShAPjS8pUxhePUDA/b8sIYNG
rj5gqTjY7b9q/Fbx/oL0FetI4f6yQ3NzDzu9N8LvCOvyfiaVd2g5qDhscdL+xUaL
44Ok6kL0hvxEYRlWA85qrsKUWWpxniTDUHTUkM/MAllG33DDnKbUxi5/uF+oLjqr
Dc74oCAVRv92duzXexTCzxF0Zx0ev2FAs9pmuST/KhoxCqIlCAfrPFboFUy8XAvw
cfiEG9mnKUbCZnXv5xwEZbD0KaS8ekaoU5Z4YgZT5rGCQpugVq8Lh2TdcXx3xt/m
3kQIIdxVhecfw7qLrHIXFm6gT+Uv9ScnnYKfKsODnV8RWwdKiGd26ZBnmYlTcsJV
GC7Z91VtJs0MdrjRznl3xFZ0CFYKfeCM99LnZNtnALJaABJ49KXRMrDgCOyJOWAp
qvaByoWinXPH1iUSPoPtD3Jl7JCjKw+rZ08SDrOE4oEIV/JveoIFR6VInElqtWgM
buoToAzAEaMWwAHHwVrEO/6jrr8syyfrqOQMaL9rrU1k+WUAFVau+FkBqIRGfq7+
yYQCRKVnNACdHYT68AnQZA5h0CPqwcOU6AfV2x3CJF5FfGwekTSHCmSNFyhV2I9U
F1adewooSr2i3Hk5WoUIWGzB1tYB0RhaMK5buwClZxuixXBfrnTBIVQUpJJm6tX5
HnOZWTXcZQj+e0hxmteuwz9iEKILF/pE5gusj4Z4vjQ1DI6pFq0+CLNvNTlsOfK+
Que/sgvkVOUCmpGF91Nged/PgWXC7axoNVvmaF3BKK+TZubv0kdyezgi5QR4RZ4U
P984SJGYWDj52ye5udUdmCAmWeGcAyLlajceIzUOZyh9WN/7eqFl6Fp1sxUU3Uky
URYq7iEScDQdqlJqsnC8J7d+9P7ZzMQ+kOMTKkzqDOEQXOzJOt6r525vtGfFSFU5
nCMntC1oS0NkND+EyHazHac7Xcx2Sid8JT34EWd8tCwxu2V/JN+X/T2VvZqdN0L3
0UniF+YRJfhVsogzPQMgMz5liSiyvtXr17vuesQctgwT4Flr15oR6wvgfovkenEa
eq0bhFDheS5+lmbiQhE1UWsnxGPiWkmpI1mAjhFVkJR8VlxgBzLp6zskS76y2qwJ
ejiYJFmx3dELPcLbXm60tnAl7PdSM9Pa7HO1czI+aflV82x2RO5pBGbDYkOvMyeF
4gTwYaYjk2HlCIdjMveDx5x2orKDNzBzUygzJIzJh9mujz42JzyddbfgLgtkrY5d
n1ZHmzki05S02ur9JVKOZ0sNW+jqROaPZllXVFzIOKk15KCWkJtVubcvCZu/Or5e
sLu77U5F69WjXXKjWPSlxks1V1pSpQL2Xq7rbc6xN4YfPOFmKLnwo3Y3yLGlEEXf
TPeAUdRF5fx3y6GxdSPWnmpVzE0KTO+hu9jVD242LDUUBMuOfjZVc7wt1GAcITfW
qpdnzjTbQ9cA0wVuDGh66PHSC+8fSCQy2VwNPLv+fW+KNG+34/jP6Tr98yAImLs9
ruM4jVubR+aMv+mxjIv2LTxJC+abuKDWAUcTzqVvIXbsVNQFneWmdYfISykQtKub
on+zNri8g6Tl8TY22nAK28NH1+aNA69JPNY/YxDojl8eCE88dRdP+6fL3rA5jgxz
jxyibFgTb48RYBpZeu+QeWY/Cn2S4TpW8e/gEfqw5ePGyMJnYn48XqxwB1xNn0r4
TXYIwXdPUrkdWlajCRmHKhBaVddGiKZt7Gh/TTGhBkBtw68VPQjUgLFHx9gPtEDa
zN3bPnLDP4UjEPHTzBk6TXAoflt7UvYjm4Jtvi4SP7fJ2zVE9xMFPxu6MjwtfvMU
n3wbDQTqGUIMsRaD/VB3hJrZxW6Mj+bCoPBj+isNQkGmELtHKzUyZQrell5Nrjr8
cV9UtpPjWjwl8AQhXEHi7BxK1HAPfdqbSiLAFf9Euh97GCmQsvch65dN0NJaSeti
Ag0Nq8c40a2+elTBo4xH85KZXbiQ/HwoBoxPaXjuEcEZRCsrlyZ6fhDeIM4ksVZX
VDKTADHj1GLSw3lkaNnGZT0++ou/jRHz0/UR6YN8q1DDW/jRXd2k2nfLycKjP9l2
IO9fN8uaOxQo2RSv/FvWE6cKFqCKOLmzMXjjhPFzck3GH4GT8JoO4DBHVTcdys30
fg/Eh9o9yAuERtJY+Mt5wqgd/9ZhMAP8uN5m5M4z1O4jp7BS6CbfbYF7M08fEBfi
IWXWr6RScz92dHTiGxLSo4TGX95GyFMAcmxQKia6XX55SFNTaYmkz55Kc5ig1FEi
nNPA9kB1K0XDYiav7Iu4LLglRGzVKOd+x9iMGs51wvR8Xh9TrvaBJg2k+CPVhBoX
gI8As6dHlC2vtqRG+OiDz5myzZXjqnkPMjKzebRRiYZ7K+AEeXPTc1hghfxCft7X
N7weW+2OWf34VpET+mGuWll4pAnPRTsb/zgyo2fRP7HLNQRXlUlQXUfEyzVmtTIU
xCB/urGpliQ/HFexdzH2GLA9REyB61lbp0CF5ciwWiMD8WUY3QFMxiphdnZVAi4t
LgNUwyJF2dZ8kd44iIVZX/Df3EsAcqrAJAPZLkIcn0byzSp9kS/QCAV3l+QKYSoG
YVDubfwut2xQtluFrkxuO2PfhWEqrxUJkMCedhJDUcXFRnUCuWRLdMqvcytFz4aW
DzZGfyZoX+dwEgot2LX+Y0eLtOawRKY7/rh6Lo7Icz+Ozl5rCeYV0K50qb4Ia8fU
D4z+Wjm5OatJS5BKK3Sn+oyQtQO+A7RicsYg4UD0pXR3YjBkOYaAsD5vY1ZtxRP+
J9gB62DyxWYJkfnbhBmAvULLMYn0jJqnwNCsIkMe6G3ES+2iwveX0x1aJbqGxKiv
v7bFvqHLLgs4AcJQ0tDN6fJpgpTqtSnmpX50Psva91PGqQttx/nlgjlgMvIyPkuZ
vX0YiGJIAZjpddKKzcP4t6abNSpm9ZsPIa+Txd4fCLNteHhvGBsTGNxlHlUdqG3T
I4AGbrgWBBevEM6ilItkVnsB+WPDaLzzkF/Mwqua5wjTV5NwnMArCFiJCGwsnzJz
h1nP1koX0qqo15S1b1QBdha/MytW7TfziJPxZnF9BvF/yxF/Ogm3VkMBdhsVLv1Y
6zvRURRAKkJCfFNJbUrOEX4pnR5Gq60ZCMYdyEP6/Vyor/LUDyNl+C0mNK+tJbkH
Nn0nhp5EhgkvGOKMwFI3kBdIfoPKuvHU9o4e/Uh1Pu8hOYssAfpY46WAejiQMN66
uWHwcF4X5RLmgjNFmA24gUeCs8wXJuUAZRxMJ/UcHvUgDIR8CokrKCroifjXDrtF
gw4xL37vww0FWshOCGylNklF5PdJRGYI0BCkVHrgqf68ND5PPvVy5B30Ohrj4Bmv
15oaCda2X0idoj0ktIBuHpb1m2UgwL9oSBxocBfzMWFpGgDuDk4OZuVzgYEzpwnr
yDz7HJkOdqjgSeB2fd5+t0ZIVXh4XZL/hcmwKV633ptDtvj+llEvSQ+zvnE7c300
XSfRbtsYL/ky6mwsXX7SDnNhN+VyWex895PgmF+p+6hOyfwU5w4cRpoiQWI6Grq/
cWHWyjENLaJoQVLydwJwuQdf4YJviXXy8NnVKFA+Mbngz4ItsonLyWKdidH1Glic
cvdP0OxTpP/pnGG+Y3nN/AjLNgXNwHsDzMnBEX3qTrHGeUd4YKCIeVy7Cfj0+yh2
oMGa8Y/S4BoTDGxBTOc+TIung9S6wzFM8sBxwv81RpKp94VsE5xKa5QW0Y991f5N
+XrnIfymPHk7xGmXcKiK+PonnhY7qj+O5H/7pJrfxm2OcwsGgbvTWNDNspsFBXqR
oZZTpH/18Uv3UFyUsEEaY9Zkp+jVJMFZfW4lxLtrj0TWqgtHMCJq5VEo7hpNPUSm
KF32Z326CEzukp5wfTqC7MJauAmhLVxmJQ1/ZN68ULCGHiwKKvbsb/fshZUyk/FZ
CbqVITNYu3igc5HVqVqEoJWK4x06Un4qY7CDd7uBLBGeAKG5FdzSaoRUp0HCMf5N
R7biIas4lnh+GOuKeBUOigP03m1GuvP+0RWKyYH4pS3h6P+OTNxg9r8Qyq+a0t6P
UOnQ8YYohXB4euq4v7m+Q4BWQEvwLPrmoladXHyEHIhp+vEPqAr1i9G1eYIQPnVI
B8kbRowNGaQK00cCS/3Hf8HSZQOkebQsolwBpJzECdNg/CFD7GXzU0a8WcOTSBCk
8v7YUFK4+kM88GDCsI82I5dtgsrR9hbg5O3vpbaZUErrtemfiQKaRdSbSLBkw4/R
5pRIRzou71wIIUd6qZ4QWmEhSoZjiYuD09rGJNIsNjMre2T9jatGTcDfX9bOu2rD
iQPYydQVI6PV+AEwsimv2HkFPoGqWk3wcOjVgOQ0nG9JKjeVvGwE9vRUx3bDHWp5
Th8PpTOt3GnLJCJUmwTS1WuF9Gh2ed6P+S4WLwELLEbqCRZhlHohxKJqLuHfi51v
Jo5/TAxRbF4Oc0/yO2hA274NwNvyjo2ShY36kAymHO2HBkbjhUTX9epOi5zW5i92
9doQE6iPjvaZWGUD8eFW/KAmLA6eEVFZdPXvIg8Gox4oC4SWruEC+onkU+RLsFqc
SOekCUD5AAvkl8sukjQjAN1xOhO0WrbHgDSjpsZI+LhXaN0wh8hgjpSC1QNeyENs
bLlW0yfFKi/8CkFjvwTTFx9/IWJahFk5ojmIPqYQj1c3XbrYvsE+WffXgyQ1vAeW
ltPKuZDz5BoFIT/71diM4dY1BN9hgqOnKKxy/oB1b0w4fa+nLpOu9+UVaZJZNPaJ
FBVC+dqKv/83eAshIKp0TqMa801j+44Os9RTUvlI77xtdd1J3sfi4gN4BVGqGA9j
apYyAOi0u9aW+aY/sx/QDnrhl8LX3hTK9arMHH4SB5WdVVsDDxiN1UptN4ffMZ2H
jZrU8oZGoZQRShPFaMfURwTkTQNJwL2AN0eBzWbKr0ePqc/t+eqLT/03jEl/8hs7
RKdTnjjmA9hwtPP6oM+k4iIBfwQYCRPieyPEs2D0DkcuzJUVfuZsTlVHdvCcxR1R
3NsrngqnDHK7ZrxcR77k5y1AFnFpZm/umFiSqg3tnPdCFrMwcEJ2gxZblCqNfCIx
qsKKiW6U/dWpWIo7eIs6FuV81tsd+I+hYsbbGd58VkwWypTqp8yzg+DJoI9PIMRN
joPqwQ3Vf0HZ6Bm0mItmz29n/plnN/lxvfJRc8U9MtLqd/UmfSVlfJ9CgAmAeesD
ElMYE72eTGZ+JdcLVRyTgm9AmUNQgMc9V8n+WTl4grebLUu9z92q6oAlzBF0sw+D
7u4fHfAq2AaSlbEMr1f5tYH6MvIt00JsQA2yB18N/OZDtsXPf1eTM/c4rLLwh/JR
bhSUTtUOFVsBCKmHFXtsPI6JnQXCg12SBf3vskygJYOhUv6QmGcQtJbzGB8o8fRM
ExirQmkanAKcSUAFLeZ4lULCEqZpr2KT5sBg7hgkMxyIqtFHVWso796RzneM2D+U
2AstPku5ODditpL/C8hZVNLdII0QjpQUtEjDOAaarvUF7AL1vSxq0Intn/bmHzeZ
XUQy3J3HBhx/2k0m7F1MytRpSN2okkuJe11aBAY6s7JCWqKoqBI6v1tYGfVnMAn7
i/h8Kimc720CPyy4SK6v1N5VSGZDb+rVgJR5NvA7Niu3SocmU5yygphifkTDfp5S
2iPz/4b6cxGvRfs5zW7GEtohumdxKotmtE0noFAbH+X85XsXnRsj3CR3pGMIhHPR
aiyBh/ZgmpkdkkVmH88duFiyyOeZkJ7JRUuQ47FHmwrXiKr1ctatLRSOyqTbOFfI
Sg1nHXaEm5zgwYDVGaMoUN8dKQc1xPS3nF5rf1Wjq255YjISg1kQfWq2H2+w7rdw
TK2+AdsyYGD0D7mRVqQKM9J+BWzI0tKpKHKM6zbs7ERUlHX54mY2KIHQFZUki9bF
doEDZWUhUq28nxFy3+J9n18zRK79id343IXbCSziiL4rf6ZsWVcq2l5WvMLNZLQg
L4cEE9df6yujFzdo3iQAlJnjHtXp9MI5W0h6loZ6eVkv9D/im+FXB3nPQh0MQ8yF
ple93zL3djXRAByHcUjIFwaHf2M2rV7iDJhapXCNxHL1tqC61LJ+hVOq4NUKW2xk
Y1gUdjQwBDSk/5vRjNjktRaeKT+uHsszWq07gEXHMHC5xqQWJsvXXPQc7gK0f+6C
pDXy17w7NDJXWp7ChOdu/q0x+Puy50GgEuszHiJjLUP8AM4/TfoR7JZakPPDxcGu
OMXia97TZQML5mXWh84xtjcWIf6H6J5tbvxbyBqUJ2Es0sTx5dOLmr3Gx/3AIa16
kux3WmpqO90iFPEUaV+OyxOcCcWc52Yyd7Pr9AMeklVMvOOA1cSbxWUggG86fGua
eGs/7wlVaQRH0ZYg955b3um4wJk79V3w1NzEGc+bSQh35aJERBycOwju11WPXAlR
SpuQUpJYrwfq/KMZxpZENre1PkXz2UaXh9jglgdCd0GaWekGbbfO96Pa3sxl0mQa
wra9y4A8KGe/HvR8itH9f6yTD3llGbeTohU8XVfXV0QeDxHmshsV5mQmyh5zakKc
O7RtHIW355XYQJNPlfIe+d3SATN2ArEog4zg8DKtlUjbcus+/zvI1eoAYI0rm0Rf
z0ovSf9sJLvFGj34G7cLMLT2wa2O7vS4w3eYJ3lwAdgRsQU5hNC2MzCHumWgxzDj
L38GbEdlXTmBww3ECBEkCyDptUwKJHcySDTEKc1SiLt0AKfGfZwdVrsGge5TMZ1A
wPtiWP8QQc1JNNhoesn7znoPoc8JU/z+nj+Fgeblc782nqcM6VVDRYCuTOVHgwMB
58k38ipi+X8/8ujVIiZcTI85h7Je4T42I7fsJ/wpyrkz7JoO1KCzQcCa/5XptKbu
HwqD2gkVCnt0hL0GBG0iXCBaQ6ZCJYeUjJu6CNFmqteJeqyIAea5+LvWcLYMUKU2
YnQ+y9hiHnaXwlhw3btyYj7UF1K7XjW6tCFHAmBQW3gV4h2MsQxW/n/fT/Y7FtB2
GYnHPoSGWv+HaPPVrgTyMhX6GGIlrhliVVwGm36yMgvW2djYmTUmfUqTUa59tglE
gGuiLGr6ISly9u+3UgPd9iE36sBFaL484+mhMN/ir9ZzFbpqvs+OgzkQP2I9ZZ66
qLW9QW1eSRJ3G/DAXa6FlnQyPwFYXTubdnnt2378bm50uhr5fm6LEQSRbvKGqeNP
UlBST7aZHAmsRjDadRlMqw0cH3gXj7sV9yFb0TZlgF5qPUihHDudm78P6ksAek/R
ReuEdmWj5vC9zMbhpwaLKc8WoQOqB3JYy/Z9RsOXTjaap1/E7VHZrk6vbZjpgYh9
B/aVW46UADGXlz9Mc+fW8G7Jyw6jGVo6OmGNqrfAwfberWhz2Q3EONkIFZFZN+xP
2gfbQJdXjXvvSKPKgOFE5AYFIVrlJE0+5x4yLULZjNJRo9QW/Spo9cM7ZrWdBU/D
bjeOAqtxyu1NPEniUONq9oeUHdtzFmfJ7lbXRB7bGTFYKeltIsK33re0M0bufyYc
al4xKNT0CrLW9HNhxozKfe7uoKba04IMSrgE9CLlVsoYzHGx/6a7yLlmo2oDFBCa
wsEWZgLtD3RZBBF7WPnaIVph30INX4RzCFK3/3mE/iIlWcxA04mktcFj8HastK1F
KfBrOxfpmsgAtEgpna+331ramBx8tAfZ4IOeMRVZzJ0RomIjB9H+Yj9ERauFMRCR
zd1CzWYyCtgAR3v6f/RTmR4sq6pnzoEJtjHzvp7WXWCCsdhMt7aKMXUwF5cB95so
e5s+zwQgaTQNNkxIwJzhwAvetfGb7HRodRVwDeHAGL7IZ3fCOdEFEb18zyK4cnvV
doGP4zjzEzzZZ3abSXGpv9SrR5JiWUfAFiUTZTofasuQ0s15HJDCYrYULcn0BfHv
b1GknDL8AOawnDAdL5fm5doWmkTyTXTu+GtcXq7ZErNW1JJmW8hIoUW9owCesgEC
yIzUprkjXTZUiqZ4O+J+SamhhskAbal15qz0vjtBpU3uZnEc55E1Jaif2atKQpJ1
DtMO9sPzl1JGuOuBc+J+pNXmd5GOU0Yre2LUnuEjdU+jeTz7M/ifXti64tloFx+u
aHNFDUuEA6tpceU7AmCy7sE4FnDUNmYlneb/BcoxUqMdS3RpYIGPaJQ1gYdQ2/Q8
tXnP9JvzlNKuEErXitQy18tFj85NTSenBBuMUI3GDLTGzIorDikVqEbVIxpJls/g
NZM1EM+Gua8eiHSVRigL0ABjIa+EmImxa2AHerhYXKxi2Mobp1pBRq27ixvY9V5v
wAaulQZ+ibCmvVaR4oAYVY3IEa5kNsfCC+6If4BtfyNmsJVNfmphq//dx5FIJJIJ
w7zDzWfJteq2hW1UFdfm6Zv7QSHPKsoLA+/JcwOX2qveM8oojNdGAb0sICh6F+9Q
BFEu8enSoBI9XtM3cusSCVKkTSgg0st/JLgT2XQFDrS/KCzLWnx/0UwFClmo4VNP
e60a7KdEQMNx0RAn0IubDGDaY5yd9ZVesVZ41S0jiY1wijzbQIdoCiVnDTR2jL81
dN40KYtZb493o0lXUCduPbsDlalf0sQY459L2eU8/KgGd14TKgHAqWnJLV6P/15x
1Gb0w67mAYeP87Q11lZFYfFjbwDMR3EqFSxrqZp1us41O3VM3dcCrVUffv45b3un
NUPgW/db6pVzAx6z8TUj5M856EJ+4udIZYbsstSAYh6F6HMLTv6W6rClYVP8XHre
0PrwrUw6r+6P/XcnyZrf0JHX0+MupnO8bZCsYfC9O16x/sO7zDFQnwWYJi596j28
Yd/JaTxdmCeGlqMyb9ckyl6Z5nqgwx59CRfAN3I+QWrS0+AL4NnST5xBDX8tbk9u
kFNsFGRXsI2tt1NQE93QW5jdD0oufaJloq4/AnCZNoWohFuEM5qKecJNkgqsPJYk
mHueOYhTxRgZA5QVeypQbEb/Hmg7P59qCA30ngYTbHEY6pIt+icn3m9JwTQ2spus
AZtJbwJtkGt6atFQsyJ1V+i6zK8Hiu4DbB2e0eq57TEF6yXcw//2YX12c+R+wQmt
d+iQ06NmtRzgo+SYTZ4MbvhoDjScKP4Y4eRhepbYWZSsUxrr5CkxkY9XaZKmPYQZ
3CaUQ3ixPukOHrtcwf8frT5LYo6df0cY+rGJwbCmiw4FbNEVrUEbDC3zpYIRva7R
tHnDmT0wOMH0aEPRnOMBULdC21VuFRLXxDkz4uR/pSpENWcVBWc7aKUw212Qz1Yt
/q3Qnv0hL0IfmHVckt6DBx54r9ITQDKz2QT8T+ic7/7aW2GUHYw+HYMXLCelKGRP
Seek7KWa1jJpj8LM+hH22bUkkGL0SPc5bwimmnmyXQ77FxL6Edw8pySbr8dZISVF
dGbiNgmMTg9Ib07iohFRqHCCOfQpj8WEjzOR+Q1VSMVveJrMyikfcC34UvTdOWAH
etkoIku1oLBYzjeN0Sh6+0uQs+iixwe/KZAa1tpsJ7Y8qCOrdsHM3goswneR3OEg
QKatag19/NOlCzp6HdlzR0dtgV4BIXtPgb25ouHINIJSuc/3/VhsfqMOAinnNszL
b4q5o1ccVpG7jkAXCHXslLQfEAEIoYbUW5O8dGwtA4SLcWEs+MO4zoP0ydmCjGwL
mOSuCFop0TCcOQ1TzSeiqU6IaS9UAv/N8y1NDmiOK9TcgaC4FXV20KrzS4icfaEY
597MzvBDSHqpp/oY6+Uei+zEhQ8Y6IANPP4La31iKO4QuHjQpjNt6EXjKORS+F+t
BCG3qc1yO+wDpYmcVpK/v0j285U6GMjITD7RKOht6w626hfPHhm0BeGTfq1jdn8s
TSuqjbCnE7Md/+tvqzDE7WbwtCFkIR4os5+2ay6Qfyudj3SfG3Tu54w+v1MBmyPc
e06kJCl8ledjI0+o0TZGPgs3+o3fXZEEhW17gSYlLKXHkVKT132cN6KzwzQqMBXJ
KFmJUe4cDLut+k8IeGD/Z97wmQCSbvXhNbhvoW/8uOa8TQ58AvEaEy1xAYnjHSDr
rqJqkcTUzAsNraaFi6n5yo48Wfx/xxt9FUFaCD2ER/UrBfhnVksVVMDTT2mykoey
nc43epYRc9+/OZJsCMbePfXbJ8eramAyFdg6H4TVwsWWPay6yOt7vF2bC58WCLQ2
8/fIcFu4mBOEZI9IYfkOcbQSyD1GY1kTqiIEN7QwwztTHYCsbFyOzObSGHu+AmAI
tiPVNEUktpKipT3Hdluv3/ew7yjycJWPYluzazAB171vVz2J0DpAiMCWSjzgXHqb
5ujLup/4ZttngfzLs7H7BiRSW9h65RV6M596dWWpeZGXSOwU0Q5d0tYifMuPJ9jW
oY7+opxPf7dLQR3B224ayJP3NCwJdHtu7E28WNmWNErNWqdNiL9bpCLqbw80yNtf
QypT5IzRq/danTh0C361ZkVubynuXkhFMNlQsjxdIFdhMRgq9CnoBKR0q4igTzHp
AXnCX8frHhv9mOUzY3xPaziwEW6N7uzJD1HExZOyHoFQGGRwhtO/cOvNVrWyUQCx
zSEi+NP3AHrN1oMN7NR59tNFmpuiQ3ornmGdr23I5SxoNPeV9xCCyRMVnVJeOn7k
zgXvq6xBPzZiK3yRP4JDw9t7zFTAtzd09rVOIF7PljJ7DQAvP5sSiSVc30I5v9XV
bJ/nvPmmEPXV1SheB5vEK5k5H3ekum2erCjwJiSQyoaW6LBdm/HWibAsNDz+17dy
hygj8AL+M2Rk+9Nav+k2FKwx7P1ANFTAPAJ17L6MClM2M7cwf/aeZ2wwKBk8004B
+Ap498irgMFDILv3NptJg5l9CN4CewIhNYTc+YjTjA5tuepVE6vkPiB3/Ow4BhRn
VSTbOIDQzO6GpVIBgTqPi/Ho15Psw+M3NSTOAsepkAEJ1uDx5gXbjIWwQHPPRTOE
FgMmaVlHVU9j5n+Jqy/GV5u9It1HfVHP6viaTKy/qj9he9eJbpLyasW9QJXVL+Wy
al/9h/PhFNWlGGWs3QiVNmdIXJ6pAI1BaGOK30mth4nW6Oe9XA/llA4+JwgicpFy
49Mwoy1SXHS5guZGGEMSrRg0P3qkwaHoqWNcYsimV4in5mnaODc2iDZrejueuBOZ
qDRDQ1IHVTo9U7yfLvdpJQ801TbB/ZdR52zRi879YJEsb3osDJOfgHuDOAZmopwB
LBVf1xrcqvUzPYufgh8ccxBtlk+zU8qvJ+axFbXQrBFEBJEI0BhbhErlzFb4xnre
/uS0KVtGGQsBu6ef5XbkwzNuMD9SYBM2cTp1BAM+ljvNYUgQ1mMDuAHuzc3l8dML
XQ82R49i12w0B5oHQkcJAi4pTaxCyFZur8htHCuwNJH2tkTDpzfGbgnjt4UP9wKR
9qBNgiVOfOI03Fbv+vju8zWwE9UERyuE1bn1osb0nIOGLqeeXODW7t2jge1VVdeV
959SuyD13RlrqZWNM9Qva4Cj0JaRlqjcqenQIeJgonrxUykEN+i9Xn0QxxiXJ9k6
lcxINZ74KY/n4nzgXCkwBUPtTAWEomnbdve12eTQgz8hD1XJRpd43J6/+9+9XQ7h
KJKuvq0pVxxz7nRpMzXIvrwzL1yt3kjrnWrGhVnk5wpIXGTzgjsHOqu36+yLDXus
4bLox7PUiuicSaj6OFDUJxEjXB8ys4dfZ6nu4M8fXYv6zwlK33I5uqJkx9rBqXKO
vYYZdfy/Dvu4DF+NExlA9N2Wv14BQ/ehPjLSkLBmAL/aELowla9D9E8D1tJ4bm1m
kajkcWbs9UNT7j5/CHrDS37xEvs6ixzCO+VoAqXs1DYx2eBAItzTAqjCpx1IPgl3
8Y+MrymrF7yjWaIzNqwbhXE48dQop+TUcAibeFajSlEu59qdA8SOJvU9FIdkktR+
GcH1EK+d8MWP6SC4p4Gr+ZkHtbWPSZNSP/bnHZLGzwEODsTkiZ9NF6nbERXY4ld+
yRj9JKMp252/OUXfoXF3cLwooC6FS1BX4jU9iGjDolflcB1HQ3tt1fpa1eXQADIO
bA749tK20XHYISnObWRSAvpvZBGtVe0dLqIPGc5R8JY/sLn6S6dVBRXC55YdHTVP
KHSSFlzoVxLVIHF0d0LJfQM5obnZBMLRmkJ7sJM98Akdac08miYnawnSfOkWxa1z
Wz+IW7AjMYUu0qVoDPji7W2SEQN1c0kMC53ARN0mAZ0Xo//rWVweXZUQDNQHbTut
m7bG70CwG/oKsLaBQB3Ii8m/tTFwmMlWB6Ooi5wr2rih+80IvNtFuqdQ65stzol4
SJoyoptM6ycM3K+CutG2JjNwcyKBZqDw6Ab4GDaZ6fyYbUrtWk3R+CRWzKp4Gc6Z
uHHvG2YUxxkQ0+WsX90O+qiDA6Jf5qLDv//qhCFbtgbSPRQo6lMI5XCM/HNz0ryF
rj4m+xqP4NMOsXqA4bixx7QK1d63hGdcUBp+13mt7eBkSkMyQfn0Mbfv7tJ4C7TM
0USkrcJYdA0N6Oepp8Z6rA+3Ov3gKD2Bgdr+3xS7dv1bMhJQhRDJ3IkHqW97Cl1s
qlUO7i6NvdBWEcOrBTrlUhrRTXwFZW2bu/XCp3T2VQQqvw658wFfUgkHGCpWmLFG
N/L022EMtVIX3DULU5l6QZGQhADCePnw3mpgBqENpFoquFH2zLqQ/Ms7sGV6NvWS
B/w9U4JNSj3GZqL5gNLhWuKMfai1l2mYpMgkZirODHsnCBt4wuUK8PothR8NPE36
MLuBDyFmFmpuptA2AAWYFf2nvToXqlfTfoDdUWLzZ1dLz1vqHqqUhx6dM/T6X4k3
3b6RlpGS8NtILO5VoBArm13Hbs3GkyaCVgHayXhnQQpq/xgxNpVHeF5uH9+l4vyf
7mASH3s+CJW4LwRClXYsBn2sPOptJblAuVN+UOwYHoedsU8+Y6S86TrfCUrR4L0Z
oh3a2UKvc3ojCRabYEWa6CSdgc1w8GKFWfb2my6Ia2R4SiRn9MWfPTkllUcAHfk3
OZhOPysZ9ManS5jA0bBhR/N+1bsyXLyu7UXk5zNEKFseAGDd42oXUY1gTlQSnja8
KVksSV+Sbo1Y2YZR0z6nR6o0W+wt5yyfkf4k6hIH+FhtgTsaXp3UXP8XCmJQ2qAi
PF1b3Zh1KVFrWG/93RSuPV1zcOdG9UdeDOGgBU0tNw/HJHY5F/39BmbHYEMtPHSV
fhqxUhclQmfb/9g1RhYG0Bsu5YAdonEUZ3kg8XJaavMVBef/k4uauVel/pSv2fNv
JM3ZrAGdQaCajwBF0xRXKvQd9v6P5SMuOHgpkU2IEBeDTISVD55xy+E1HoLGY1i8
Ft+WhMUi6hRws59b3fpJnaimgifUsDRa2zGZZgOwo/knMu1DP/c8LC//hrrd0Q1S
hbeAGJpX/Vlo3xTkI5wpRE3ETvmU1QDmNI10WyhPg+12h3e0im40BuZPKE1FLOE1
TOyblG4ZSnmXyF1Fc7ShcM9c7RMl4eJptnBwyoTCB3x0/q9ubJs27Mout8sRKAzT
bNFsY4L+svIpfUuJIDT7XZeWtZKApGcYTds/Fl8t4nDKtjejqwWCbLbPR9SI2M/a
ibPOhXe5NOVK9lq621oSbGWqtrnFGr90kadszoYKy8ovWFV+/p9iI8AC7RoAJQko
hkhK2uR1At7+hlZz7AXO7mRwtJXc6WYbLMYZ7MVd2XiU3O2kxFC6WyU5sbOrCykA
7WDlVqXohjY9umLeW4uTxY0ivQfoFLq7aQ6khIAERYU2Cj/Alp+c2Nw67168XpU/
NJYO6k1GbkXSJztXbhcJKrKFOT1/DtwC7HcPumuhUs29nmxUDOhgMV3Y2XJvmmb2
ylf+wsMfLE+7YR389+xN5cj62KN17wO90h3/fWEAckm8YvNtLX7wJU8gWovZbIYv
RDSAPs9Q3fGuqhZVxn9DjYe1gUwmPcqilcmM+5vNsyjJJ+3guFb1C7sdeAID3L6O
VnamWkp77Ube3jqtH7lYiMXyL3aEUfZPzDBsI6y1TtN5iHOxXLPfPao5cZzRvFZg
8LqMLMkyWUtH4qGjAHDZT/bkZxLv35Q5Vb9JMJx8tAXeZffG8zaWrRzl4EkexIqT
xOp+P0HUVeNWtC9tPAPaV6LKiAmqIYOpgBqYiVqQ7oHCQlOMJCgSzjFM4MW6C0Jo
l70lC/9dDV4Vj5JESIPGNSXbGJEUp5ob2Ffe02MPirNBJhf0TifmlHmZxdzR9lUn
2CdYZBBV8l3a4O6nU6iCH0viIYBsBeJ6aKpM4f14q69r5//E2Ma8rKIpxR3z+hkF
g7cTc3MCV0bvjQh2mUwrxBKrxbiqpety6BqYhwMkF9quD8IgTVsWmyL6oHzelmHM
x2d0T2EXJAKkCKHM4muLv66EuyhMtzzOp09ncSNXFOd8cqwVtrXuRVIyJQyJKvGu
/xlp4LCwNpnKArkvhRH8matR3+U/EuYuqJWF4lzJqIY09rn7hXQP+U/4rJlR5BTw
UzCcPd1kB8vqfYwM5C4iJujUUxwE2l9ql9DHdxgtIw8KHd8S9i9dR8Y3MIr+lBrS
E9ON0WeYQExG1dVO+jkXQR90zuR/DEy7lhCNlosHlcp7WRjRoHtFT+5cKlIBzknr
C6yTu5Rou/ZW3CVBnbiE8FShRpqTOhfNAgyVmCf3GsLNai/wnYvYOn/4tpraobOs
wKQ0hqsK9Fe71watnIiZB4R4uGjO3IBFk/T1j5l5YDeQGVuFIqINAjdzZ3ydApTk
+U0m745MzuEQReEPjduX6dDx4Wk4ffcPJ4ywz5DnRpf5UC7pMlLprII0NXBPSueb
saUudEaM8UzaoMBVO6p7DkTa5FpFz7Gf0j8w+cVKHRrfvwPfIGR5oQLTJZ2sY/V7
0ShUnt9vALu/HzMaU8Qc6AvOLv4WPJAwskj9+qBQLHIQHNHyIwe2p81qoPRZ3Yxb
pR/KaOIqTve4sQr0IPNMfhtiRiKW3nKJCoLTmmhX3rBtmCbTtTmoBu1JcI0MlTew
71af+x7Ma+3QQ2uFBZ9cl+QOOyPLLOcUSURRtZbhtnlYhejxZSM+8Cjd165X5wkk
qMO4u0umQYonwwcbAn4fjXwem8+9ktDdyidTvbf3QIUdie0xXqNYzTd3anPUt4sH
4H9Ntp8mfzlbbvueihSBPIYp/WRXwQK5/nzgwLDx3vgg+lJD0FnPOGYH/ovw0Z4Q
Sy31tOa7jNORFl6jUAAdIxoB0dX6oiGJ7VSoEbY+9qDhQxu69cKUGoQ8/KbuxhB6
2TEEdCfxWVT7PnFZR2nIqRragRg+hSkQVw8Az3+DaC5MV6F5QyySTdyaYrBs6C40
fHJkjG1f2dCWuUt7izuNqqPCeFFBeidBFfmQ5kjLnKb70sUQG4T6u3mYi3FDZzE+
Le6s+g2Q/umrYAZSXBHAP74FQZREZvepNCm5URifVlLmVegxEwYC5HCEgLEPrL7i
dSq4Q2ilO7bu+ljEPkid7wGROyiFEo6eV7BIXmxAnE4jytzCylvH+LcDa5gTHcEV
g3lFRVnJjQK3shFDODrKNarksLc8TCJSVn4V/GgUFamOIS/1nwByLdnK723VIOhx
i5nBhWrChen+Q9xiHCnKDSuj0+Cnimbk/OviA6sBsiRDIFGCW8/B2C1epEavK9OP
xDaczCTPIh13DagENDcNz2Rh/wYqKqkh54jTbtSCcbtONbwgHXffsasq+sB+q2eP
xiDU5m+bzhYUVr1RHq55xML+1z5hUJ9Gs3gFcBX/S/lJuTM9M9X6nytD9QP7Hyd2
6aZKHndSWAFFcaeedbYsOlNtEOWCGi/3fAbsax7fRF63gg7g0g9f6atHJ8EiNR45
0ViKUxL+RQarrv3oiq0aVlbVBc3Bfpx8VckrN4eErZavdGQSyoN0Zu0SsM84/an9
gIA239X0pEENxwb/pcAJWRvRDIu2x7AjnCaxaWQ/U5WdlailabRxLpDK3McXGgMS
R43ON69816Kr81nIxrs9BUPz3eLJqcg0Xe++tCMa+nmUWM7VLiG124czd5NBARJv
AuvSkluPpEouwyey3KNJsfoCw3mp+287oXwucWMECFXrjZdiTO8lq07MLWS/Ltlg
Zww+5bAp3l3SKQIKzoa3/O4WJN82lRJ7KjYZBP4KF3iByqut5xcJb+sT4S4tQj2V
GfPJ96QOO3Y3++AHYToPcOelXGQPLVfGNIWzjB2LeIZ2YkXD91MU3kqqY2STt3ug
NT8bUDiXDDhio2uNslGb0ArjXiKb4/lhfGzm6NCk9i6m+YjhCLKcxoeLmfHPNh5O
FhlPspzHFLFbCRT+CK9N4Y6U2h1byywv5/LoAJlcrdTBBCXRFzpZr4cJdkgzvdtS
OwghZyZUZGNeKYWDwsPTwjEHwOnGw4ZrC/W5Jv00Y7RbHT5sMShGa+eVUf+j6bkv
7GmZyFvC1hvZjsPVp79cvDVuuQdNb3EWT6wQ5bIlqNTu27BLH7IBp/JgcuvZVGiu
l7pDijixl1Ax4Hqb7QKzdwYYR3vdDK3wAlbM1zCGAcJAtoF6V5o+sYhhqNE8QqLY
jKItVVmRxU4n1GLueW3k6qer22tCnIgx58+NcuKxL5eyPYWEYiy2ZHM58qFQxNht
va5DKLuBBTbP7yVlikOC/eE6itNxidCLPZS+cXwoXnWfDfb5vYFaayFaI/CY9FYg
3vuQ6h9ANZh4XhnLhpjuAf/Bp+aCOtlD6kR4iX660FnVfPYdWbO2F8MglBKNnnUm
CEMjVVuE6734nw0+63/y6a7zuYyiK154ldw4F1Mx7o0mYUJimsYXFRiTe94wFoGW
udFqO8JkIfHo0Ot1g7XRAXEEEzB0Zk2t6zzh/SCEHB+0ESdrROvbJm7lBgjLTpDO
WPL+Oai1w5BSS64iGNAtzSWNYT9TYQjr69cv8cgaF/vqUvUar0TM9MkZuFUWmIs6
VvNZBuaLSMVC8nCEvLMvIlbJ8tMLSWgkMHAvXg6Ih9dbXOaWjgxe/EhJnSPjAbdn
kbi4Ic3Fv+gdQFUSW2I/BRlGYkfW1DD94iyPbiYpsmDUfMrbd4F9BP9t6L+p/rtB
cPyQsFIncVIqFQ3hIKg48KB0eqOLx2psIM3fz3LpJC7UrezpQWTQ1c1xxjktyzxD
yfR1VPjm1NVJ45RYpjikSTUsF32ymVHQe7upo+k0UBnc6yvNwEClUsw+s4g1DdQ3
ofabKTJGGQCX5mk87CZnz9EcNsU9RietdI+60yL0w3D7LXq+AicPClVO7wuj7x+c
VUW/ngKQHudWpMS6OXIz4NzttY2uUuvIKrfwoiye4Vu7ISSnAVJZigf0vkKHtE7W
jhU7MLxFhceQFgy9XUldYvvvyM5U5OojvkyUXhL8xnXIQRa+hOoA0miU0ZjTwKBB
RWrGgsOugZAsPro8T59oVgBnA7UzAR3tjAEOjMo5NZto4+LQtVZXF4r8mhNkHdOU
sp22m62SAT2dcu6p7F8gMrn4ize2bwurJdmSR8J4x2PA4pxSJbfPJ5okdTvJzw5K
bc7h0PVy5Z9D32gpBW4Y9p+xQj6ttRrroutv4qmpcJTj7w/pJweNjR315LAPuzMX
TH1F3/709yY6F45waLvLXqTR75xccIQyx2JeQYMVxc+g4L3QKb8suSgscoqL63mk
eW7ttoCppGcizOi1VwdsDzzAg/jhkyALx8qrdNx5BxzaGmIfIlmgV2vyHM/1PBPs
WzHXSAuJ1LCGjgPpjhDEidmU4oNDubVyRpUjQsftO6q+cnEnpIJe6aXW9dSREzDZ
fTabjgBth9qGOXRzz/VBkwBWofY0KPrvfDGP9SZIO7HucvNFpid5uwWSKlk4Cji3
Nwmx9J6iv5iIZEWZu2OJvfAs+bLdRGj7IGTXLe13LQD3gy8TVtqppDKty3tqxacW
LcJ7uzQzMh1y9En8n7vwue6T/0jcrI0QYRWATj3RJxVk+4BEM8ZAbzMVr1XMEHBj
Ra+6RkId4ZL2PzY/DAzl5JFuODcjJVBNXw3VztPOkSPlHW6OJ3+WC0k72OZ1VGNy
8uQUUmYm0Q74r/1RQFCUa6iHcwLLvp9P7/6gjzBhLsCDeaBNqeYlSstH9imVctaf
aPqlx/K1F8UoEWQkyZtNnMN36ZrjZsEOIreeBybrS/BvCyCLPDlYAL07VJDcTQ96
OW0lU5mPrjjjVjWaU2zApI30a4MFG+4NqkswK7urFctSX+Sgld1TJEP+fPS4jDvC
mP8N6XNysmn5Y4tSvzDb6RXLzDy+DXR0cZ8i5kgDo3/mzaErHPWdRkl5s0oJf6a5
+s/oLIMaqo3eAqIdz6yfaAEu3wnTXuKRtpy3MpK7Ui0Jj534TH4vM8YOG8Z0g/zI
DndKDLSlP+PDo+Qv/mtDk+2k7V6Elpb/eyVrHg+K7E0uVm2eQ7Q89GHp378pINUL
kL9ggLiIwwanwLnB+ZgdhRb+FJCRWbvOrUowXcNq0wOKYG4rGgMxPYRIMQ/6Y47c
E+6Wj4EVYvTMh1G94JYhywunKfoVA8UPcANbfgzx0U65z6PQcw/Jk4CP4BTzP4yQ
nlAUJDxDtsTaq/XiuLkxF/nJ0ufsrjh6xDOFhL3ned/aO5ldVf+qllzSyfSIDATb
7b97rpkCJuYefMrj8f6MYIcBpmJeklGgTZ2J35+KjdlCgx5C87EmSjqwOEpKIfsz
+udJ5nRVQiugDHMNXq5X72IaP7PxMT2JSKjH5MRb0mM1UAEfqaOaV17fs7rIhtP5
U7iE+VlsRHZ3rB8h0h9lRikF7GWPqOm8FnCczZkVSA9filJDBDEedjDJXBHfnxFQ
Su0yf7C9qJfhgcVFXYJR+IeqmMcMYXyA0FZ0JfQ275KMK7v9NElCsiQGgjpHe6oh
2wZHaOPyYCYHVZltCrbr9zRgkZPgBK5O9CMTiiPCIMDtSwK21/Zj06TRqaHhAC12
zWp+vvAgOefjGkgRYFHRhSucXVXYNmv/C817KJXNelSUeelANRsN9epcMnKb8R4k
PXxO4aNP5T0KbgJ4bGe4FLHSo7V5Dk+O0+axKfw2IY/dEcRVD2SuU4r2q9Ao5ZgW
6U2IdT9V+R1NuDLQmWpix9CwFHtHvcwQb8nvRSDKL6K16yRO03gzAZ4zpztOB5gq
wSUCw7E1/5e5Ba2IE+WfBnju5V5M4ToCLgMc1X5Hucr9V/2kGyB7ks0yq39eVLxC
Sy0bRANrdJzFK1H38uDCOPN5vuyMwwiEU5QeA1ECRy/kZNAJcYzDBoohH7W1MxpC
m2fX3iFkpkrwgsfzrxTPJIvZTVoC4EgRjMhvQiBAofMGCSb9dUu6KZqbSxBh9S7o
EbTKmYOyE8X4sFdyWvVV5rhiusjt4/qUkSFhuXiAns+Xkg4akgNzKFvU1CyAdk+j
xjnExtXfQg7JuvQ4STaoiK7SMzp99NT2zGt1Y+eLAzEfyClRZSe+5XgeQeeJLrh6
HJeB54suxVCiOjYIbstUB/gWZabqpFfzmQvctsbS0cOtspNWZeJuTQAtXfq4DQZZ
WBO8NsF47MUlBRiVLyqs2WQ+UNIBng/11qsAw5YE6m6sC5ghHvvIHpR0dyOxVjz9
yKab+WDbn9/Qm73kVUpQhyzn0rGuGj4+phXO0FIJIPsrW1zztBn6pKhSH+u02yzg
lBB8otCUC9NKtqQzad8FUDnKG++mbuK/GLhNyN0AHQAiahNy9cWu8XON+X43aqJN
hCHeUH3iWnB85Vcgl5f/ZVLmcNKwM2sTTXUGfvN1GXikIGcHsr/OxjrbqCxpN7vz
Y3aHbJfb2HO8mHBicsHD4PxEoXwQjWld/ZMP2Dx8HOQbp9ONsQIjySgsWMv/tYE1
i4MjEu3HpUk76ul5sxuQnwK5sflgDVnk5U/cSRnaij1jwkvv3eh9MqoqZUWo5z8E
mD7cu65fP/sMKE+noqL5+dk975KoSfIfFU7VPsOHf4IW7+x0UVCPuz/nJxRJH160
SY0OUHjY6X71DwavUm2nvaz4B4CR5LkNLNziJbqPi4SVppq6yHr56P4CPS/dNyRW
YsKaKx6+E41X4g/UAMfGNUFUbw2xeRn/9hJnp9uWFPY6xJqYNOda+L6+rjv1aDEQ
PFnQIAOmem6Y7o9lvDYZL2ijfMC1zzV/nYY8/LDtjMPUj9ykYFHEDNEWyP+QzCVB
N1Uytl75T35x1D0CjF27PyX2pa4v9sochGlGnrX/JpJOvBtIbCq6GgWcm1rmSJbX
6eClMQwx3VtLyHCyXS7rEejcNnqNVErvrlIuGeXSq2/5UEZoe4j35GM+CJ+tCPpc
MabrW+9Os9DQeU1CKuN8P5szOrEKb6iRkBy1yRN9nSLyduwgsSl+rEzO8LKIDHlT
L1YYJSeZIqGqQ4jxhM/YPOMsRxjghMevIu43ms2MejpfnjlzC4UuljFYJUZWK2xZ
uTNFYWORQNjkvPSGqxbOxG426zOWcJiX4WE3nIvq09ao8r6pBy9mNbaF9+YA1i38
aR28F4/ZrNdAIe8oqWEmQjIcHx/kB5XqXEvRSgFifhFg0WrmhuuggS0KUAagvP3j
v9IUazEM00FwODN369RTELc4XtjGZxjbkBsqcQIicQSGtPF/kyhyoXK14zj3T2P7
fofaFW+HpdZelH15Kuv+nQ6X0DDvHQa1CxwJaJf+3SGexTM6vG2Csl20IiOaoZ4m
i4DGd0pyX/2ezERtjLGDYYu+XY+ssjAVfbfH4PJD4w72CVTOm87ypjKNdN5ZGyFv
fmOqMqzHz6DKDJYjtW7VCsVs198DLdPU2U2QjJC1rmRxvomtyJHnzguuJDqqaFdD
t3wAL98Ff9NTlUO+4Hn6zXazFrjZEji32PPegIb1UrwLxkTtxHPpiQBK385qR4xp
61y7h5AcnptGjnA4ywfPeqyP2RxcrTtOxUXJCu99rmN4AwSGMNcdKJ4yDZ99qMLl
mvTb983T5KryEMoH9zF10UGkE+rYsudoeSEtce7Z0G4Hf7udeth3f3duTXxbMLFL
/0JeoRy+mFBkV6rDH31ZqFvPQnkQRk1LkkykO6Cuiw8N8qvQvgRRl4KQTT1/njPL
Hc22J1G9gjH/2DEqOG/yckrZE9G3CBAeNHCcNpTB0VfwudYpdOSSxnJ2ZUi7HKkk
XV1MO3pnhhecidkW3CY+DVJ7SnKHHBw8qK/LukhCX+mgygi1jszdp8XVNNXfr8R9
o4npVdByv2SX2t+PwtNu6PymxA7SG7nOM+sm2BgRT7rT9bifAnjRE2W8UiNvy7UH
JqYo2KnyrBW7SpHbU2LSuNJ+aLMODq6DgY59WU4PFp7ADxMpSss0Yocq60Esci+2
ugSVOnw2T4QdClUKZIR+wdOYzexijGIow36yfNYSEy8RrQwv3wB6Jmo5Y3VWR+ok
rms/bNGTKghCJ89v2kycnYgDSrlgwmiDQPmFAEmLYEQrkha3SFR5t7joqcAzOw0f
bf04DXG9crtMU4vTLjE51Oyj1E8xBLMRtKpwFuwVi77y/U7I71OT0KW5BKev68X9
yw6bZBMM+Q9MM+kdqGaYr6CPL75CT0y6BCifBeK4RiAPN/oi3uCvxFs1SuEyd64U
Eius4LTuuZ6mwDZOb+rNvov8l0YUzctC+dpimHb67r2xTXoeBwEryQCp6L8fCoaT
X9t1ubygwvUKos5SH638Gn/5SD0/MD2PUicVaYHnl16GsF4GOtTlkzyrukE6oCA0
USdcF7YM40o8Owic2mgas52AMq7nCCRBXFCLyjaHR7uG6FWLjG3VwCjSnEcFTC9c
654colFhv5I67tpqVACC0/EBahnGDNwnV6yooLAx3c/5v576y4bLne2lTozAh4hr
NsoIwIb1xS0i56ZnubUksguh+gLdvM6l7hMwDdK0ltptDGWbXvndU0EYkXBKwfk/
65pE6iksEijjrRwrOPzAytJUuwSqcy09xy+LJrxzpV6gDWIex12R5MdTCACJcO4S
0mMTTI02k6k49kZEK/lTVuqYO7um5cGbut0SDKVJTZE/j7DRGOEB5+H3xrvOYHGD
NNbPbL3gAcLztxtYGnw+WTseyynV9/l4NopSemab0WDZphrUmljFYp9Ni4RIOxyc
B4asTg/Fu3xbccqdJv3UG/pgbWi5aBFTqZ2ZWxExYwIYJff/7ajpTaGdJneiCRal
nXJclZ5Gy3OckddaRifP5B6SLI3hnCebnmMb2Er/5cdhd3J6ouPxFwB4Yb8hav0b
YQ9gi/NiO9qNe8dPrs2Ygog31iaQNw1dWcZKt8iHYaIHkeQIeqXD8S3gYtdClN5g
llcx8CleItSsNNwK+7UDbTh0iUopyhffzL+p/XeIdq8WgpTAAPg4MpooSe7K6tut
mVNvKPr36EvvYxTOAyCFaoL4lWtDThdmy5AoExYAFRPTlMzCW49rHdfnng48xG/N
GDvJWa3oyF8ljv9zdq2NnXdWU27MMtik4zV8ze5Wdy6bCN9t0FHeysExp7PMT5oF
Ie6qTS3Is8bALLLjtejzWl5ikDXAWlR2mS+nlWy13OfXVCxcK+MYeb6Dd4MLn+uN
Z8rsDaF2aY+QeFb6Gkz8MazNOnMdnH2o1YDRr4ImJo381zA91RgZCXffJa0b2g3e
0zl8GuD509m5mjLUhUqLPy6qAbwvxgK8LLjyvREeh3VnrylBchKDI2LORU6dcA9N
Bn2/rG97cY32isfpjO7GXjY3umLJcdR6KTMd9gR6fVTLRvJ30sBAfs7rKCxUTOgQ
XCPlHqe9WWiOcrYYNGoQ9AoVFdxv9YQlKFCLnnuALVANEohuImc14bIQK6+35TeN
zJHSSbdHK068cc+aJ1zJy2e8OESr2p/wwtng16HIUjBFHBYGdsWLKSZtFEmTYojD
5/8QNkm3nx73gJueu9WcXdRKpS65A41M9JZmDV3dDZWglzE1MLOWHg/zBp1VXv74
cEveF6C7h6U+nEsT9lHIY+ACFguFZmBXNAXpBvgHdOfVIg4kKuG6tygfmT5/UZbi
COHvXaTu/EElFxDvsRi54A1RyddVEa5iXDdSEENcLEe8BOBrsQ64aNT2RJTGrQuG
xA5Z25cHoY8+kBEH2Ni3US+oRuL4DFx7WZ2XkWrIZBUAHSoR/1ji2SGQR9tbR5Qo
YtpAMxk+S/eVn8X3Ts4+D+HtELACMZOAK7lI85kC0szDnQ0gXsPFPBoDCrOB/why
40HIf2wGT1IFenKRoDWub3Jp3o6Frlo/De2k+J1LQYwyOEz4IxOzUf8COX1Aost6
9KEoA7KG6T36OwHGpYDyEWERdyQ/JvjFuzHpimKP/lmP3zHv3RqG+wnmxI8dMXMp
OhBydPkTCW+NXX4cG64Hwg1bQLsHEofS3nu41edi39As6OVGo+eg/nCGWDIfy+yz
Xws4RR7K1DfiNHgXaeveL9ak+O0dhuA2cBhfAPvU2u3MaKJpglKoBBKE5kInHm04
QgrVS6z12akhi+BaY01V1E6NRESMiLCJoCggiyCKj/+ke3Ik+B8Xd3u9IA4Z+90p
Nzr+U/AuBtCHaSUH85SmrO01FMfpMEUVrvs8S7TsgDV7oJdeVHE54pWI4mkkSLfk
AJkw1EPzpmWyrz9NFl2w+TcKeBUaPUsVJ++8z1QbbkbgOm1x3dt0U/uzE5p501zm
HuB69NULaX06vC36/+OJN2QA8EQ/mS2xzp+4MFrwH1ENHWuRfKOvHMeTo3BN9SBr
JqONfYT+sYVRjR+P2x917JBxyYPCYAjVssdunSGwREkfOjpluIf/RqYSD7IdJZtk
tOjSVnrjzamn54wZrDnOAVRFNKHNzJ5P3eoJAgqP6K57HrmYewOdpt6oFAPPCUHS
T0LvdqSuo5UZit080yHzacLeSR6+ReBKLFm/PrcS7Ttt8aH3ZQRQLKhv+jQfvCE1
PNlwKtfCaw3enXFt5LIv51C+4J2QQt1vwhLm6dwXeSPQlM2UJUV75zUFu7eW0ex8
joMlJkAAPc3rCQHIINr0xzGhZh4Pt0sDD7fFsBcxHkeMDeD5WjtFnHF095ju72Kz
uVblmeZrm0nwwXAE5adpRATIvFPKr+MI3v32kvYXS/iSlZH3J/7NOBUCslwPSAVl
0RdHOOuzTbpfXsQf+/vxrVSGdG0o0+u7O58jBPuZOXelvySUkd5HiicID3hEZmnG
F9gk4lctjtb4vCjvm8xzewGJFtx1Pc4JkZe/PDs+HcdsemuSt47ABua+MAp2xRBM
WFb8jqeWkhdUNye7Kg7uxMwIoaZ8e27U6R2LyJY+mOqIxpTlfvMeiNjdVXpTB3Re
8fvmja/tmT2yWfKFf3b4KNHU6X1uEk8JcWsjFEt2asa4YlesQfHFeqtcjDBZnPpj
cQHldLr4DHEvhv0d9onhAmPVk08ZOFQwxMw78TGPtG0NDyzdZ578jlbZjdE9Svi4
CxnhQ4oMfKOFWnAFaBj/sNqT4EnzmfR6UhBqHe2TGCTYGL57jNQYt/d9Wo2VTkiY
HZH+goes6gwZbBOLuZupKWcc5/UNE+RutR00ud85HbZ6NBTtaHU+LHqiEloH3jbj
qQwVGnlL6pnigyBYBqforf5eYOIGwJ1FNn3BIp84acs/COmxOoHtMBY0hHagxd4M
QXS7eRldnQEFiLr+HTPPcdEt9+eW8tVjXc54bAxDTOgHLDkAuPLyq35J63l6XUQm
FqOFavoO2andncgNqHlvEEuIeafPPrU+PHKXaJPKBhya7l/QXoFiVZzxrCJdHD/K
WaTXM8AxEhiMc6ABWR/6VAe+AXnnFAAOCDb5C5FlnWIZ1INl5hWleEcu8oI9Q1Kr
LyUnsACwm6b8Ubbki/4tBqBpXTFrOdF0yw4+I0mdAa5xicgImWieG2Y9+G3xwHf/
CzDsp7e216504phAFBpSB5MzKaRq/CDSfofHsbouvn6bVwyqjCB67iveBuwCZDD2
BGmDrpd1n+buQzkA0zoL+qBCbClZFDZhJktIUsEebaBd5siDmUE7C26C2jjMEjhR
0iPxQ3aFUSt2EBEEKd5hg8jdOR/O3+d7TFWCxv16EHBwzpEAem3wEAnPh40zrJLz
1ng4zZWnY+I4UX3udeTRqsVxFRtN7VfSeOY8i7WsVcwf+rrQxgCR8xDRvmFS8ENW
/88EsG7oB+0270se3beR1rtZrtolyFTvWfgPu9r9U6Wp5z/JEqgbxyu2e8euaOzX
wTWniLOBae5rKPfJHPEabaON18n5EUC2XehoC8LK0cD3/Dh3Q0IVNsq1evzX3E2W
lKypx1Cgckv9jNEBfDPqc0rlI13Iu1knnmA90LiW08l7RAfVeHXWCvIwyTwxD9Q0
te4A80JXU4tecBtSKyCK+XFZmvafXCJzIwVraeoeCkwPaYS+IsVW2lhSyNtQnT7d
RKLVJ0PkxduICc+tbTVutVaNU+7Lm9v5JiwXC/76JNPyhrNKNLNkwpwjh/1EW+OE
so/XwdRY35Kdk2nFem1rBvagsy8FMLpXJE3gs1uhCCbeps9K02Ox/Rb3Ne706fV3
TIZ3pc9+uAPqS41IFlF/RnIV6uAW02fuBVtkew9yKqwXBBjm5pOQE9T2PLvtQI4A
ZOrGMM7aBsjJtvmgn3rD6Ugo0uzz5qvDEIHGWwcazOWWfhN6yCaGpfOSeAkGydzY
zXUqkM/OUju11hg04RfYWTL80B3hi1WmUavWaONTn9qB3YQc0IpIpGvm5q++p5f0
1fWiQazpcVZXwM56EEspAETMuzru2uyFVRxOX79IrGSce5vuUxsDN7JfXs+XXzj4
+oh4IdATnkkSV0KLza+uy27uGgHRRgqt3shApcYZNRYHaNRxHfjPNanHkrK//XxP
yAiSq37Ox2+Evy/FOvKGwPcY5rMzIHxOALCO9Qm2s6936LhCuB2F+MRGw232lLPZ
ovHMuqL5uv5RZaLb9wkB2DMyYLz4r4xpfaXyDzxrc8oAmZbPRE7n0KHkfID7mFcZ
fqQXIJeEo/GP0UsJiFg2SR2NkVN2mbFna8GE8gyv5Pj3m393y41iYxq8H6ymNGA1
knUCaGxBEWNCMi5mHf392I+5uc0oiiB1UOw6wYApZt5EPVMRu7znQhEKzbdc6YJx
VCHcI294wsBgOutVbjbOlXEEZIARpv3OqSq7kSIosYJN7v+V6BKvUHdhDHrMJODB
N3tUYrlLYbZBc/v1+6vUKGjLek8i14OtXiFSUtegztBPfeIHlacqF7DuijzR139n
2lu19NDEW9oOsKzzVTz26TyVeS6ZL07wysu0DU8+Fh7eZlUxzVFUAdKpGwAUZ0Kx
HD4zcu9Eac7+xGX/0PF6lTw/mYj1+8bCp5nkN1GmI+b3OaQN1WrMjXRNiaHHlRyi
+RIjvcFehwS3ueh394LyX4vdsIZ5I8HTbn0gfbWbXJ4R8THJLK0XukFNRXpsEOz9
sArXHjXUxFqfOqfrKyyEBIuHXf10tADF+U7fLkvEuenPPHdqQd1jPWJfDMv9eEA4
XpQBReb9rIiyskVF+ujVWFprYII4WxSJ7rvLJa/zke9ZcfUbOL1Ysno0h+DZn+gH
VgowMbjg7Yy59KaCu97/6o1OUEn7NleV41LcnzM3/4qk6AXImoUTUaPacOnGRpRN
arR+U6xIHc0FjwVPiO/5BdhBlGbNbs5NbA5AkYyxBif3KVe51gtgPmm6EdhC+tlM
va496xmxdCerXvwQrgc7K+fafB1jSsh6ARt+wV6Ji5FHZwAy20ZL8QI2IbZs+SsM
hm8Yg//e9LneK8o1lBzKfGhrtuh9neCWgGwQeY+ZRPQlLoNq1CygqdqWcVtWlxcG
TloZ07rz3ZbAiNp80ZrB6isS7AxEI9l4Yizh9/tRgHYPqMMqGmhY+Hg0weJ0COVI
mUSvuxGzHUigDrsyHe4V6r0x8KBZmb+A/ng+f3YKDMSIZpdWzmU5A4RQ/WOFSpf+
dRWnK5SHkvqoAqIHrpPMDJdOyUsOjUy0izQky4zhpFU2nksAQFjIZL5d26qITS0y
dLA1c7QgrNeo5N2EoIcZJ1Krd1CzoM7AQwJ5+oJeYwv8VHdcLgrNY2d3ikcigCNQ
GDLUVUP0a3qZUlMGuLc3WEWmSRBFZRf/59EVYGuwyE2qved7xvLjhewnspLoel+g
j8DpJdEXj+sAeigu16mipMvRBXf2JqQCWq27PWBoNgYdVEYBdWBW0VSATILgoI5P
FNSMBg3CP5Z78JG0uYsSqaZ5XydSdF5Gyqfnlrvm1scDIHGseRSHdZZGa88nnjXC
1gy+vzY1eHzReDYpI528vzmgnnzbWyREFE7u+pdv3gp08aToWFJ6g0cshJk3cxbI
pVvodjOpLcqqdMDCb/NB505hnyF0EIvtt0ZBYFhN7lv8GfcAick9L1zeGjLY6NVy
v0PTl+rL9AkBeUXK7YRPWNSUIG1qzHZFowFmjHb8EYCIeuOTTFkA0z2H1sAiFa1m
WA5+n9AUoWCKioN/7dnwukCEmoMVo0GEFvMoaRVtkc8+a9/+YGpVefAJeLFSw/tU
a9VUlf8c7m3iZ6sPMxKSnJP2DwtXU4Zmi8zYVLvG40DuxePg7QR349+2okKzNAz0
H5gG8zbZA7Wbcg04nNO/+AjmJlfyncl1MPDu+30SLyvY/bmU4+6qWSVLtC6RGkps
REoK2kxMVNb7bVaJ+q4UyGlL/ki+dj0ssDbsaM+q9jBGcO8WpRH1lYCULkx9f93d
tZmqbs/swDZGKOpBBCpnfQZWmSFxay/mwyFrDTUK4hnHVxbyb3dxGq15oMN+huAm
93k571D63UNntRGzTODXK+Ymtn7RW10PgvtJ1ei7dStTTUO+qE5Y19pmKLTRxMEN
xVnNjg9BYo9g0KFwPG5bk+1CudoqTm/DB2udUP6da19mCdeIXHHdNiVvEB1LulFo
FJHV5i39s3bu4JIOBqwnDlTRO3sYUuIWMTWfZD8SizgOQPQD7AAeuXv4/Oab93Ae
qy8dH4OsowpERJnGBGc2bETGftJuUn4KC172mM0n5z1495BO3VtC28B33qPizy9I
WEp7JHfKVfEDM1Brx6r54JzzKUSkLizhPah8FKMVR8APG/HAlJwdSYPPa16TSzR0
HwzPHA9sS2PxyCYsoSdrJ9GSoEkKxZq6xe/rNPrnd67MhuZVdTPKTrKwX8ZgxHHp
Su/mmGSrILBsuE2ESewkghe7NQ+8fNiRJKF4UfRwjs1G768xj0z60WrM522M0IeY
61i8GGK4yo7nGoxZyQo7CBpbCrQlNB5Tl/5v/FDcZp04Q1LLPmeiepsrhW4bT1No
UXLB+5ELPjBoGMBbyC/MwdYGchc8XKmBFwnecizRquML3w3imtajCbd36zf7owaN
HuLnntzhGoRC5SkVkycQq7rPJrNk+fjQCxQeOiqhCEgJBw6XsU+meqgXCZRJyNEg
KUviNypSQ3tNgY0T3FwhSn/f86KBHjj7jvltWJQ6rxYzbMTR1Y+MRllvDY42LdHF
F5w0jDvP/YOXDULKSnkox6E4SU2SlL8iwxvUg2zs+P//+PAs+k9SMi3pPI1aBU2R
V0FEK9fBSozg8++A6eckobKPoy96jW4rdoIWKhHiqhwCpvTsx3m5oQC/3B2aIJCD
0kx4JJox3PPFDi8SZS6jZNxbXQLThRt0BNZ90GdN3qmoz+/eZ0HkFIjVVzylXR9H
fPYUKt3tA6YMJ/VNUvmNVvjCgaScdLtMMyRIBnT7+bAcoZKnHvHwx8YxxI494Pjb
Ooj7M8pgNQvNW2GTm2LAl2+9dku+gdgCOG5bLZbD83GOMDwRwZqJJIkXbLJvj2j0
FnCV4mN9DnxUKrl4LXm4n5+/pefz+hoO3JV19pu3E2WGvx2vk59Z+Tq79ggpLJVH
MFxmtGosncVXBmNtJqlyUAVLt9Qp/S+MA0WHst/ha3m3e8QoXNHqCgqOESnLPnCq
btqkcbBblSsARJs7G+IUDwj/QTvHnk7tVzhccELcdIcPyphL3Et9EE7xVvxGL+pV
sLhk3aRRFiK0nkgYsAAO4XUcnGpkf0JQtTKrY1LHdd44nlujaZZ82Cr8ydXGcbBq
6JlXjitfW6viejzNGrnx0UpDjbyqb29jXz9noceq1AhJ/vwOZ1LnahXr4n1dQi1s
dqW5SF5gi+djAetFLKtyLwS9xLNcjWKioPdka5wMjnWS788HwseifrDAIl79dHjD
709ho9+7LQQSobFoDRz5LnBnMmmoaOwu1YtJb41Dwvj3JAneaSo7eJ5L0wpCycmk
cCRGxrP107hnr7BhDiGxCeRIsJCz+YhNrArtubWhwJQW9TZi4H+I9KecNLrTHvQr
YSAQ80G4wIsgF7MhYV/iN1Yhl2lw9GgI9SMlDDb9N+j2fDYuJ/+HjS6aKRbTIQ3H
BLO0sDZbKSr5xNcBeq3XcYG0a+IVrHAKwfTzbjXKx+OfLqG8iqLfK0OgmI5V+Ol/
pNtJTt/WcOU8+BxhbrY9F1Fh6BRobOhC4lW0X5HoUWBzQCZOlCE68ArdhrRL+28K
8UKu0y4FDfe2hl8j/vakiMbwIdaTfFSgLJS5Tf1LmtVKNBykzWhvCK0ZmnTPfWvm
BS8Ua909tLl0FLK6O/q09diPZWJ5fYOUOqsKJGZssNj3rxWmx/oq2BPr+lFeORGR
UGS4yMTi7oY3VgOY8DYSglq5j5AJmsJA4pZId+qO/9I2DTnwCtSZMcxUP82lvekP
tdCA67qtMFdgINjShPuVarZNw7MX4SJt5z9BE5gON2RgY1Tc94bNYMZfgCchpuJb
HOQ6w3zy5fQaPE2TKv8gFg1kj8TxlNj/F2eszu2kN7eftex6FXlh6QN2ASM4zhMc
DE9GmKXQczmWHCpae++DIkeU+ia6e9DQGcETEotkpBROUxOx3rR7YKT39smDaSzs
yF2kcuCHne/72psftYko89AyNEaPn2aED5EYtdoRHUqwZ9PTKWT70l4SokkiZBJV
FR6B29qD6se2KdrowW0WIzpaSzh0TEO1lwhtj88SVI+eBJVJQKYkzk5g6Ha9vPC6
mKDLi4a74hKijllwvQXdW2Uu8nbvaXkwju62LVdM2Urqzx4sLSqn9IikJ5lKRY1A
RrlG0SEExsDkHY5ExNmltb05PDpJPGdruWxqh7CyxOeC/7g5XWgtHrsPjnS6Xvde
VPTu7EA9boKOBx71+fawe3vZsOy1l+SIM/+Bs93/8OcswhgLG2uqkO8Rkid8Qq6b
9rJ2gCGhB7WO187AgwggTmGjPV4RtmSYJO36OUmttvZP7rlVN1b9P15KSLwdbtnJ
Tg79iQBeNn70Ln3KbZ6P3pDyG0/oyZW02cCZWjapc3fvr6ljXaxPO51Q5RqeM9ho
P8zeVCLKmgqMduDaW8NWE4lLryjXB8CSJwhyPRExTh5Lo8iCeFp0yTxme916VU7B
VkxPdPTi9m0QZoAC3V0tEsOQ013u374DoeO1VZrCGtq+EUyKEmLfXX3nvqsgrFKZ
MlL+E55H5YhpHoi9wyU8lDFKAU8cpY/6xD927rIualECq63e5wYkES531rp/wnSN
kxsh5IJnL6vMGAmuYk74WkSkamAPCQHvYwDaI4n/sDstrbPJAceZwGXrDwQdLzsB
OxhCxXbgimSt5Myf+YMBwJR4ddek1G8s9cpy/om7DDr1rGl2c7dN3pQzVUQaz9Bk
M4Q2WngEQA8/r85tSNukrU6qhj5LLrS3YJkzLC2Au1ax2qwwGc2jhbU6RhiuqcUc
oHO7XTpYT7FzzFV3x6X7vN4Q+tc/duE8RzeOCJ13kYrboP/aYfQVJaDCF2gdJHTn
OM/zqSFITE8GU/kGloxEPDen0bQejMn/Uchc8tWYyeDI19up3dsyqVQEg3zDSDGa
I/4o+2IJMhc+CLWaTemHuCFZw42he3M+pG2S5eGQMxs6ybO58YqJNbr7SX2REnHE
LJVD/AHxk9HXFcysnXhJYJAnjjwizOCt0nGpAWyuXfm17WPRLPj7zw+IIxEzMhPp
pkRxsijQkQcwxyRbRKbtWqXXxwJQnhDp/UjpXS4libSUoqr0DvQg4jpbqYknBSLf
5e/q0d9TU4UOD6cGL4ndLuoJ6bZgCZE3w0e8lKTYE5ialGvB4uz49NTBea8RNvJz
o5X6Bl8ZWo/5kdrArMssN9k/MPoYRwEvhA4Yw35OrJ3IWW8EiXFCUBie98v6VUPb
kgV80wtO1GikTPPxdJXmUpXZqdXFkCpFquaQn7b5AjERqDzcq4bjugeYZWWxTbUd
4RxmXue1WRi6ph9uS4B1ZJNyGiy1ceZbXj+yYrfGTQaJOOTAxef1mvw+2R8vapW6
kMYoQSktvA29jUIkoQ5Vaj2zgLYUPhKvDvTtk07jvrp+ksfXuVSsnZk7mqvCwk+N
zF+/CdtRg4SKHYzjI9Ts7oUfltg2F8s2qbvYCkfF6raklSBS8sROTjwe1dIiGIUo
zVv1xFuxeaL4HjyrA9kGJp/5dEdriWOASe2KwI19iu8XJPhwG/neqwfvTy8xS+HJ
obS/xfuvGthAxuwWzO5HdgGVQ1h04xJzspPlslgGlxkR3OtBBm81qDCN0sx4J0Cl
xzUVnWZfplE788FWyWtdtgJy1kXTLN9CdAm0XZiS6wVv0+uyDzjWgREe2wVMZWWf
bI3ue0snDg7X83IWcPLH6fkmWSvxQ2EfPiTnHhd/roJvOELslw5YPTBDgPQUmTHL
2uU1rCiYWkWi5+LcS3iXr7oxnVG3n7Owyx9wzwv+JsYE7jnBwNSDY+InLnSqMAAX
EVCZ50PL/YEB/Ly+4dSP4bzvs65ODyRMUoP1gyNKB0lBnLJe+s82XAg2ZVNW5cWo
Pv0GsCP3Uu0p8AtEGMP6E4RLuuVjvyv9EtnHJonFaEsjixqfiCiyi+b20sdADcSg
QxOceiTAG7yr/z3bEN9FRQDhpU4JvyVHNR6H0X/WOugzy89Q7YKaldeUn1jx1FM8
87NgXrz2sKib0ou9/AHYGeINNQhJu8m31jtf5Jv23zK47CBu6FDXNItXYgcRicJH
ssVYgsXb83s3gkfdzhy7aSjc8xSkoPRzCrAHUON84bALWqTzL/0p7zT2s4WaqNTT
WkEeygfSMX3j9HVWGEcqio+g10XMtmqfz97WwrVWZUEjM6H92jxLjQjWBl2wY89D
kQFUBFD703FRHmXN6w3M/ufoYsmYpsxat200gSOzt7b+EzXXM5vwigywccyklslq
OJ2QhTp5z0/3zS1RGbUmGUHEQkR7sbY7JcrzN1xchSG1YXNYXMUer/G0dF3OiFOx
AZNsTTtA1OwXdDPx/wXISlgcWAkQvn/0AO6CZB4jvxS0PmywYeHIq1mKYP6i9/sL
Wo4Q1ySTYuwKvAlhR0H+ynOWbSGcCRnQ9oERnl3ek+ZR6eG1gHR0Q1sgcLpkil/8
UV9axjgnGHJJu08+5NYNe1Rh/vCz5VPqYLdRPKEJWDjF5yDEUgWBvRkt8K8p9Q7p
to/X67DwAeiQJaE6pXIkszSbOZk/OIQUzC86o7TFpetrqGJ3o/RgM/1dchWAzQVA
Ds4IF7pAP8uPGjJkboJyJ0W+GhzCQEm/whl+4lNIieZixHTxxHHKBrwkHpXJhsXR
/sQ9UR1RhbQnJHpSUZ/Gzu7R9kf5B8mOwZ5LU+w1RLCf1oq1TSRYanFXDLBIvrbL
36z0pTp5u6YqFJTkm+BRxp8ZrB8WdiDjD63nV+Ppk4WUmbuMPE+Bst0kq/jOfJnD
/Ci38LUHTqsMaYAA7Qs12ZlSBP94BJXknC/kU/R+QAG3xKfZ9sDDVa/ICK9b6y7r
n6vUkSueGP4iqLlR8RFpzYp4+JzBHvkaDbqb/ks60wLm0zRurU85ckMWLCtIPH7t
9M3OpVUrHko7Sr2yWpghK6E+FU2jgFDyYa6p8c6RB3QzQaK3DvjVZlLVubnkmDn9
OCqvikqYROlCapWtG2XeQEWaWDEKoIiAhJnG2oS2hBD4r9LdQhWMx763RDWb14tb
7lLPF6XCN5tj6JE8SH1gB9RofLzIVZEouvqts8rtp3fseWLBXF50oG/ZxDcB05W1
Ils0WZnF/ZGzUxMLgV/+upOizghDvc5Y/1/s8pE3q21WmN/J2ZQ2GsWkvItppZlB
gcOONkBQ8h2VKwwz7PPnvgd+p8DrH8oBBUXDUaBBPC7b2knUYtDqrQ7B6xOxPbTv
PE5bLe81yWhAoRTS9IWn9UN2lw/vEPUraQBiSRgEDFYxBBOh78+HMYl7OO2CrNan
J8a3iHbk3OXh8hgfhA2qdfEZ3HEGzPxRcAJW0eXhqBWm6eBp1vOJ+sz2x7JQ3eoR
GPWNvJGF3VMPkvkGlS8FYMdVKgMJwjEXN5yPLACtwYprgPaNWO75YNcRrGUxkCEB
TafbxkuyOHmHcDWTlaZvfkeMM2d6GRAAg0nVwZKudw792n3s7hFC2jybRHAHUwi5
pWaAumltQKvQfmooZ49kbLqYKUyFK0b16kkcqvO1bJLAhfNwlARRHdVLvUQOpW20
9VoEEk3ixPvM6pvdm/vmMxl0VSOhGyZd/e6NEo90QuO+SAy0EyVaSAP14SPvfP5o
QC05wXyN/kCKFuAgxn4jfbJi5lXpmMu1YKBvDEXAdhvIIDWFEEtEHzh6Df4jkr7t
G+oT/5/8PCaiCHn0dtXF+jAD9crj+JjoJga5El+QO+8vg0yp2FgiWNPWV3aJ/5pl
SDI2si7/22/5VfWBjFrvdEA2eVPLw7mq5w3YimyBOTgY8hUcbyMPekCF0bH6oRVg
2kJqRujWEJNk75fjtFYes/2YetgFbi8m4rrxI0p1tVTzXJqWdO0HFMUVHSCV2r3p
8/33BrPd5Cyly66UN2HSrirgA/Nko2LdiGk9BFdkJVrgCXfGshTlJp0LzOrkYH08
13YTBZEexg6JH0zxXB2lCULAvuXKs7tEvcyAv7XMqm59BWeuuYZtwqegj4DPhbMX
4K5MYF2GOfyUPPIV8/vz19p0MOf7uaOVctRhaMgIa9JfvstitjSyi3wbXOgaGhGb
FjqhUcwAN97OFjdV/v+pd32SCk6N2Tn7VtLie6T0hbSBXnd7/W3P8ocRKqPgAF3E
SM6KtatSVPBcUTQROCmXev29HVvUZjc5gB9LeTKE7WAW19lKsReIzUZifIqJMhe4
xetej0qJnCIiVH4n2pZbjUIv8pI9joZkHCUn8qBmsA+7tsNva8pb/SgpG2cYom9U
FilhUWrBnK4KlGs1ZdV21+KWiF1JroNUyHzDh3anpZnfAmw8sVRgOvFO6HwYFq9P
X67T8T+V8SgA2ENsMrmWwpN+Gu4lC7U4BNFCsbCn+nd98BA3VWZd1sJgdxoAvFgc
PZ4o9qniv7k52Kb+zjVry4JKyFrtgqbbEoZXyN9gyS7WryV9vr96EbTFVq0vfwiN
2JK8hNbN9GFDZUx0H2tqIb+pLvLKnwGVnmDmWTkSwp0bfMGoD/rW2eC/QuRSgmL4
1S8i09sbdK4spv1yGtpwI8nT0XlILEzOy912WrNvhXdNKnaTaxm5C3b9PUr9LY49
7bCBb6rNOSPAy9mJWin9XOsrdiy3ruseVibmhvNW6yBZOlgOz7OtEameJtSTXgwH
+ow3tOQCyVWwhwQPxYZOLOletqpIRUiQ1IUBCkQHtXSDjv1uaDh+LzDfp/mNRhHI
xQhrjqi+/MiMe7OuKKMdueZtSEdjs9h5fvz+fHqZr/kFC5sbKMh7u7qA+TfaLxh9
OKp2amKTFM9phL1EyYmel+dwnxkj9Mqj7+peYtOKUQaFkChR7f8nBTjXYDrSHgUg
3d1LOj0Jyp02QsFbNAy/DPjY3NhVZYWeb9kkaIeQ6nw5j5TisZXJS3aZiy7n0UHq
U3QRaajU02wVR0wxf0VkxChAGA03hO/Il+Hyl2wdMo/iWQmX15v/GPbCyAbrPZB6
RTyQswf3MgTWsg5Soj3CJ6+Y1X+qGhi3RTXHJHWe53HpnFtM7dUCrRp8LDm5ys/X
yekpD1QJ9Hld5mjNA5YMii2+6QZknD9Uq4H5kvOSzMAVGHR6qrRR7eSdKWuLv8eA
47Iy3OPYMT/qck+jSusjj4jSvZ/4VlZX9qj8KOdmBF7PuQ9oYzRAwpBaByt7gGT6
gZx8Kv+IUf3MDmQxAQkQ0bEldvnYY5rz8xO3kC0B2o38KWNOjNSf70WObVLMvQqz
WO6PQj0M9ZGMNs/jtFVF7Ge5yMv58SKkC6gCW72SD8r9GEVN6PFeLtIgBDsgv7FP
2nfGdAlG7XGboL6GyrjzHCB7Ku30hhokyBGro1in7puXwAb+nSbw97N7xyXGmtR6
p6Wy7ecZnuFSAbIkXEkGiGplqBOm8cFl2oxHi3aqxayRVwUxoFphgNTDvF/BgAZo
tQT7qqmpV+ITO2JTHOdSdnAWS29Dy5xEsiICH/VPHNsMo+hZdgbkz00NRK2JD4Py
AH0IkRm5Xn5vggVAwBLdMnfLrd3K+vm8pP2IxfV1PsI1J67icSG+FO7jmfEmm/Di
QXNRf3FivL4T4rYLbMdJyByXDWEmZdHJKiganPM4592NvIJQtYFKonXVlLqzcA6Q
VpMKDilpbMDWKT7xsyWYPB/hHzBvsNMnQqFkHtRhgIoNXcF5bqnY1xWNep9EVCvx
rohmyZX+kuafACwoRP9fwkoh5MuPiYp3tvwdGH4ePgKmqNO3BIfg6ilAskNebIuI
Ds6EwaosBmbwSzs4RYGCrCb4uSAgA3ghe3WLkrS2zCjduN+Wb1LCLc1yT3VKdEgb
etWcNImh76BgpsZTDo56rAlZ5R7rYmtTCImOewNICxrNUwdjDa+rpV9DCJQq432C
/YdVM4Pm2iA3jC9QbCdsOFePDAyRA0VCsxMDk2eU1bgfaDoh/OpB0AVu1Qy3lg42
sxaEu+Vl3lJxMK0J4HDjGbJi3bH6dsAZ+CSDzHxwFUA6mbcdBSGS+gyzoF0UFDGI
BV2TrIMmaGL4FlB0rLxAzxdpZo2qg8GZBOxvpcTZe1Wc26OF6QaMvg2v/67z3PQS
suLl97jxvOfa7TSFy+/SmA8vQ/4o9ECvg8fB7uUotLiTJ6ibG3JV+EwAunTnMv83
WidAqHOVnw1VlG1Vj4tcCapS9aeSLSO9EmuFejMMJKUe8bER8Lcu/sgplCirZnLr
5pEKzXBB4EdHBlwDsAdcOe8BBGol41IHkTlbXw32Dn1b385WwJqgwjSxdKD2z5k5
23ClXC5d2viGyJnBQQNu/caWZNpfNkD3eCnCvTIJh/6Ipf6NZgGzJho3R3qj4tlz
CXhyCTeU7GwadJtZUKxJcP8gElRxU7nve5JFLaA5d/PFDhc0y9kzHlRNqNgW9gm/
20PwNHlFQTWO+ktxBjXmMcOxPCggzj4s82uCL7hUS0+FvuWePVZ0Li05Nk1vhO2Q
jWb9sj77Y5KB95xx4gnOHvK3F4JGJe73Qm6Qk50lP1nXhBbyNRUQYAsy2RLDmCUD
v0ozDbtsEDOJysO9adFkWH+QRme2/vC2Zgjae9nbOzoe69/TZQ2vW4FJTP6kiY/h
Mkeztq6OOIDt7saM689MH3+HM0dihqMItZSVIdb2I+CHM/W8lqa/K+TXhMHwWjUv
f8U1cq58gykPUGn6kbKD5O3sJ4DjSiNd9hXjASVHnNLSCSJ5395myEI8MaKaCqPG
k62NP22KXcugcCg8L1qRdc532XzySOiWvsKCzk4fzZ8pLa+IeE2RpaM28TcMjhin
upF5j2DcTUkXdWW5016OvIGgiHsVjUe5K/2ia8dEiVUfrYJe4nYNAxoxZKtyC+Uy
wzGqtg6oHXx7SmRGiAIciPTOWgnyCCE+IdG2/XFTWvv5L82sdBRW9tMRn8nlCRzg
Cyuf3Cu/TnhdSPAazMZKHj16FlGhQsNbom1xGYw11UyaHZUxKhm5VlJvY8gGKRN+
txLRY4oRlyz6KDd/n9MsvO7yW2VA4chJEHLpAGYyT3lxW7Gp0o31F4Xiuf4Hatmy
abVWra6sPFnsCoBs4qnvWW4ZkYIMAsvb/4ix3dPhHQV7ZNab8iifVGqJzxBD0fZl
8tIRjWaV3Mvy+lmeuQlQcEQ6t+IwU0FnRY3E3yHZYo2rJ+79Y4/e4koxXNiPaD4v
ESLIe/VOhhblQ+5im0JHuRuLG1nHBz4ZuWRcCjaNKN7yNFHAaeUU86fiRv1FxM1S
72jBdj/ggPiwNE11iCXpUoetWZmfn2spEH79FNjwv5f5O+NtHPK62XZLXVxsJd5t
m/wwwXouyL0ZDJ32CcbTHqqgkLTytbAQJnUVUh7fhUB72vSkwkC438jECoLnWozp
Tri5RyGBu8iHhbH7+TFVLfrqMlf8NSXvgY3jKhq2pzkwt7e9yjdIbuM9Lb5uQrd8
9AU5L1y0IPOpF6o+CLJnt18xsJUsoPNlpRFVOpknWHDJTIyNJ19HPOyEV5YNKVCd
sTyqciQNoEZEdWFXx+HlLxanovXNWuRKodP4X4zRqXHtu3C2UFdCq+Gj2wjBVIbr
Bs0hcRpgwgGFOH4D6HwgwONEnnc28nPZjC47vYWCtVS72M7jj7sYZabH3pHIkqWN
M8MJ+3HCsrZzq7zKQkqydrKd+R7c6ddmHK5FXp0sAJCDQFZDXA6cUxqft7RvgMRu
OqBe/nVhT+VnlrzOO05gOxoc5Ev0b6VbGe/80auh9c9RmGw9y0QHpzcRPMJbEP2l
xI8HtlRu1bjMthbmKBD/QfLnumhU50FkOeP3Q3hufiJV0QKlGV11/d61USw+BnqF
oBWO6PAw4wik05TkNTrSbdeZR9iGsqUdhR51RHx88gFPOlEOKFy61mK4oAWL8HAs
IVACrkxCohTa6R7AyhcvTN1M6PV3VGAZWD3T+cAEj3eniy5SLrp0kAfMSISKAx9b
eO/T/sDBgp8wMjuSvz4BxzA2h8rRLd4+5DENje9qlZePWGF7OGYbEBUYWZh5uAPc
vyCnUW5xFH+guPr3EmASepTcS0HCw7N+H34pvUIJ5l+gMELvnX5ReZal5D841yS0
6PLTiBauY6an4rB++j+UtEMh4Ix9lRYTcHeua1pY7MyVO0qyrksu/c3u5kaFw9jQ
wOe2AhSj94jlMGWUuaja9EH5dLTwNLxh86tL9crMxOgWg7hLiSXr4gIVwquhiMng
slUNN5eCJjwnPgbGQ91rDRgfZFyOQYWys3zNG3U0MEtk39MfYK53Fqj0hF5TC7Q0
DaR2B+fyVnypQb5k1tXOnv0icm3/gJR/gY32tl5HtxjS1ViVUFoSx/l3g5qb7Oyr
0agMI5hDJjf5B+t8mG2J+kl9bbu13KSV/05dYp7RIlbxK5MKH0zLMbrrstI1/tur
+BP7cegudTczfpNMVSTqxljhn4rdZyY1N5x8fZBvCQ/tUH8YNCra3IM/RJY+PjHm
z70gYve9+Jz4nP+0sZ4Dc+4vRedaxWp7HO2FlwFQIMRY/kDia+Z95bG3PgF/9Ajp
G4w4gZj9Qx9xmgfKTme6vjW7lDfKp4kGQ9D0D5Xu/xulK+6h6mPi/1LQyLLESvh8
w0fGglxAYkbHsFt4BCwgNzPYw1lIBUiprsLlJ0IxjeWvM1qO8YdXqA/FFhVQFwc8
K8sHBU8G6nvTYbpyUJbZkaivqaSVMUpIdQSr1IPOp3yBhc7ZxIhjonja4ZoWUtzr
fwFwoxuZjHcubOhL9C4VerE200zPLb1C8JcfTCUkELxhmwzWewnzcj+FzFc8yM6E
kVHMdwfG8Ydf8+q8oJPMWZtQZj+2H7lkxTHizcs4LxbDfswQQM6Fd+ltwhjRDZQt
yY+P3jQ+RvCKSEGT4kepgp0uZGtyxfYeTK/vjrrIHi2MHCbSNMCh3xPWkgQpg2w8
vxq8M5jH38WemsYrWGOLGCG8k3oVMox7TZpGRn2dmGZ1xZCJ4C1WHwFqkf8/uGBh
xWvHpWhWTUmtTiBDG5OymPwoJQtQR874Ve0MZjwpQi4yJw3TfABFNAbKKRBI+VPP
lhO7CJPIci/YEJOXVJdPOjTGQuVc9IRTuQ2F2e2UaE8PInc5uljIqThTmOvqE/MI
aYUGnP2jJsmZCcD11TrDL1IdGoSAURbPHqks+iiaHrXHrIwn8B5KxIMqCtwfvkjW
54p+dt8G7w8nzdsOQn5SXMu+dgmXIfJBHLZRfHW/CVJVbKfqp+L/bxiu4EFYJE5W
hzC5VjmNjWPBMo4fe0Iz/t/VTCbATyaxjtdra9qjiWLgIpapKSuO2T1nO/rluiJT
JRRPNc9t2/8UGvQSFcBnMPQnY2euja/euvs8vamm2ijI9Z6+/EpQ5MXqeX34RPUz
grxctOtkAJ0zWzx+dSRA3ukFMckpu7QRfP/WMNj9vTeorpkGYcPHP5sY+lIZRZAQ
ekGqyoBV5QwyRATTqti2ta+5gmBWwHui4uo5Ylw/Ha/D+b7suEcaU215WcNBuwrr
ro1QbE9Ius4uPe+s1+JEw68Z2IwzA6BS0ezKpklilfUXiQ9IB2gewkEXNEjZGU/U
99D2fz1YbIdaEdxWqxgGGxK/+vlTJycbGYBv/89D4fjr3JYtIYwXhcLK6YlbnZoy
XIgUgcWIwxzop+jVmK/K/+pNqvpXiJ11VLqBb+IXJnuxsObKJ/qUI3u6+0Xa2xOn
MkuevBO2KR3SutVdLb2YOVITTr2oqD6nRqbUm24LFTCub7CoZMxJHiL8IWxp4wY1
kyc5FFgXq5PAgysMywq9ZtTiQ7ltxeMLcwRJ63LUAI6uaCLtcs9CBwdxvVC/LNJH
v/sqNxzA36Ut4ZiClFA2gG6uVLgjWxicGNtQuXhc0TqWU8nvJ0NfywP9157wznCW
fyV2i6c/PsOQ7FMJikNJS1zBXfz9lhGNbl3+LJzWGRJFG00hFZUgaQ5Oh/slvdnF
MG8XLw92cCpFNIrxBc59FRj4N1uFVnyzRQAnoYTdoOgTlJO/8BWyRYv74ejR+pUI
wu9r3tDE7MIMWnOmfrcBvG7KUo2cx1EZGGY9FLunzlziDkMc0Te5suB2uZWK805o
qwAewYJzvzqBUy4Jbasv+9QuMliYwoR1YeHfX3COaDXMV3FRRvV+Qce2OkdMV4sK
U3deATy2CpdLK6FEylRY3Fl6GQv2CogOPytikLdtss4cNtNqiuO+T7MOkPZzeC5i
4xUUQNaBOQocilvjPu4PKwo+1cJAdUxMJPpQy5Untq9kDPbFwJcWZLWKv1WhmsSl
BOJbg7FQd8yIGJWuEQe/Qh8RS7fSJezt8YilMkruQ/ydcJe+5i3Zh4l0E7U0ngdS
W/YRPbpKo6CyIymcwlksTd7a3PidQoTNcXqhMZVN3P6XnmF81MaftaZerO6zgUrW
R0Q/VWv13S6DMuSL7D8kTFdBfg1I+P3yhAY+S2WNP4QEKi86FnNHqQAsA5M8hu/G
QRTcETJRjtRq8O6X9YRMQ1gqsuBPtNHTWD/dpLOWlv8WAcEeDn3HjhrrBWZUzldJ
eZljZr5BastlEClqbgA7uIus67wW9WvkDlxsPJUtRJYAaTvyL7/2gXtD/kz9N4U/
5vuYiyvePZVzaKaw3aZxKIGPzKK1uw++s7xBHJR+VfMEmkyiwEdmb7c9fTxO1ASU
225YsTnzbdPscTVt8EVS6X9eitcEE5Cy//0Jiek501zMIOl2g6yEzlUT6DRgo34X
Ki89mthDkA+1kqMqntZDI2j99Tmyd5dJv6tlIzsNI9NijNF5nF2ZLpNACn7xGc0v
fxZKgMjSDaEhsyQhp5sg8YkkSGOVUA7pu7PnyfYtgJfoqHYQjoQ5k0Wy4ZMlhKBa
bVhSgz0gE1d5ZOsYWX1PYka0oAAR3ggsxo24lIRoQ5GQPebzP/sJDxnfZ4q8gzAX
hze8H/te0DXdBtyeOm5m7au3Ldmx2mKDwTjB2zt3urnwkFz1J0RfMJUIkBW7ZiWh
mLJYd2halBMX8GqhMndnlXjsBKTbxMbHrEo1NoiV4rIhZRijakUMCf6sOF604oFC
FEY/JUuzGzMe06GYRMyEVYsruAPaJ5XJ5mEuyIV1xsCCZ/TIzaCAYt0kuiHxb0TS
CtLi1/JxW73aYQ6kFT5SvL3ZxigvWMUwkrLq4sS37HoY4g4O6usgrNHj5KMMx+xn
yn73xaWJ4hfE+Jry8cL7HNYxL3JJB9iNcQV5fryMqXSYg5J9SJHF8/29Nvu88oT7
xmXTzhn0gli7bmPhh7M802B3NV0csff3GGEubwqUaCRKK4gyTaBNwgv70PFhzufP
7qIgQqFqojgROt++EbPv/UKHDhQn3ZwS8FFBzbXDMTFyvEG92yXMtrK4mEcvAMPJ
8iSOB8cFrHKrMzFf3t2cFkiDBx+qcg2TwnJ52dY7faNY5x3OFCSuTYhxsj/uxR0X
PR1d5HG0RUiFmlQEnow8xF4/Ykow7rC6OFfW7GZstRzzRaWl+zfcbsC1eSP5J94S
s95A9KEUrE2ox/9kTgtXSxbBw4Q3Ib3pTmZf78NMzL1VtvKg0+ibuE/WNPKbXjlP
WXWSZvtOOzrNX4U5nMzTWIp7vReIV5UTrXxvAdI4FafIuambY4OG9CS1pQi5fOK3
oTf8/kBTrxSvb7ocWz7QU3CHMqDQ5umf2e8ZIG9fPgmHxUgf0xLgxZNPj9cMBmzt
Fpi3jYo1WKN+QLh8eIrQCc7VyN7vHMz90RAGUQyIIWznmVHRBovMspF+B7prlurD
Oxk2jyZRaRJWm/kXgVrVPmj7pDNvhKxKFws8pfvMAE56LvVDy2/EfjUn3CY4Y9fl
tYmQXOVgkGHB9En1putuVuA3wgAyzc1HCSSe/P9OO7Bz7ME4x4k/WfD16GD4i8yt
+MkPuGvrOrofjAmtrl/UACmJdtqgvXBQ8UlkextgwCwKsYjK4xQsvvt+sq7GjZg/
JXgI48Hgh8Lui5CeBEHwU8uxOyvXkScDaOLH5EK21j1vFeIsbQDvFGATlkRrg4Y8
kz5XWnau/UFI/k24xdnN+zuvlCIGoEtzx13RPfXnFv1XnpsPs74qkcLiikX2s12u
9ChwwvCAoaYXxamUueIrTZiFdCZUojeIWRjOQLx9nidVSRvkCbPvI45+aR8WjJSC
7fOfTHT+jLRr6sYpjDQk4mjjKD0UNE3PbdTuAgN8ntDNKJ1qUCykyv1G7b1YsTvb
aDUowV4FYPnGPt9IAD2VjkgO1Bgn5KTvuxN01skzYTDPLCBWltb0cO4OnFYC5kav
PUia8km7Z7DIJZ0TzZ0pA71lkqJgKosb+uF2lsHe42GeV5mrYWCa7eFvV9CAjxzy
ADvpgcxv+F/d3yC9OpVuRG3eRk9U0ysMY54fnOKXQHLzY2ff5glqFVKcRvpfXFOp
aao7OG6DWp6s7W/cE1O5FOg3wuCJemJye3UbvUQm8FJGRxUy6XrkPHfFupQrtF4C
wBhG25OITpft29CZxtmQorsmW1I4vlYVE7WG2nyYElS7xFvJTvr57SAm0mPNlGY6
qtqL/c3mtQju/jY46K/p3AIAHUHG6MnlI4kaO84+ncJ2I0SrPAIz1l86YaK+q8ns
mxpWbh4HQ3H8W6yVm592eveoMpTJbg35+herW/hxSsdW3qwwYOfzXoB3f9k3HVJh
qsi62JD/90v6Qd7zD3AIvLM7Z2FD5SCaBu/dgeBgorm4vxGHm0QMWDo+iNVkRxfJ
4MEK6WjgrlNeB0g+wwL7G2gFV17PAHdCD8O5KkYI46cDRgi7he0j5nrFrBfJDw4M
3qmwXq9E5guVuxux0VfMU5i9If/qE+bke/aVjD8gARVVyZYKtCgkW6lREAbSrdSq
3HS7WSDEvnaoUq8NvHa3+SgmwyBCJnFrixT1grapqSww6XQlOgq2nLHJ+ZXf9C/g
0REO8F5PeDNE2WGDKeelx+LQe5bB9SLbslUdtcfR4niW/l868rOQSc0xU6jG/dvY
N7FITSCPeThivxFXvPPwPjP44MkR+CpHW1hsbUVa7LKG7ieF53wk4gfOr8LvEpgf
ca/lP7SLiAwbZini+mSyvBtv22aG6yd93l25hGaeDZ7MZIzcqQTFY3yJRr+uZ67A
GWvdFp5XDN3kfU9WzCbd7QpoWQOxZLKZrr8xfGGK+hlyG/04OX1Bu+X5ZsSRH/tP
xd5ejPywaId7PLTuVUYsnT2xfp6GiGW9dE8lYsOzCX9yvfhNyYmKyFeMoY5q2hyT
ziNKuRTfnQ6Ypb6ZBxJhPIaW7tOUI6csMsJ6V9GBxhYlYsmUVQCNdbWCzUb5KwXr
lnyg5ZeG50Ec+YbmQOQ3bZyvAIloLaEGVkf8OdC8TX+LsIAxZOGTTDQeC9BMyIKJ
NS4IGn3rP52dwx565JW8BPHmO0geh0/x7WdLLds7N+Q5B6SLNg+V7Qfz0EVNfpFr
XWzsT3KAXAcJFXiO1Ocm+A3if5di8r0/riNMR2EF5YCiZ1Tz9VSR7YqCF+umFQRV
Jj9cMBXsppBnr6y280FvvA+mOhIwlG4p7ChrKvCwTl7Golo6na0S/+ss8wnIRci0
ahP0wljtMDnF4eV3t+X/QNSEOR4EyqXFZdjHhu0Ki/+HBbcv8WvRx7igsOX4rRNr
ZczD76W8+jAaH/5IOoLosyjiqiBlyIrSCw/dK329DuPUCfkGK0MTiKl+MYNttO1w
7LBA9wsAY/sVtGDypjcCA6kIcAQYrnsF6jzHBm+1vAx3Wcw5m2O6QiKtOdN7Qdob
Vg4iC7CM/lCoctINt6+L5GmlttgTVE7zE8W4g5ONL4GpLfFWRANnEb1gT1BHke/D
VXrAKqmh75Ze1x0iMQyDYZTF6Y+IspUb5+ULzzC2I3qHnq1V0i2uV7IFzPlbB0vB
MA//FzX3I8bD/aMTqHh/ZCD9SXB3P4YxxSy9mkbL8Bgv0SBNcMEufGdhsyn57Uhz
kDOK9bZHaYMBBL4/H7dtGc72996OyWoa3nF2/kYKu4W8uLHFww8MkD5k8wc6yz1u
IO0ei0aXyIKoCKss0kMrUsusvzw1rT32fIuXAQWHdIIgvLrlEvcXZHzJHBvjUNx6
2RRmHB+YNg4tOqh6zFYxILrTCJocKYJ5rpcjRHbrjRaOed3LMWSyOqYa+WM86/in
Yll57lxjc8tQyjwAH50PFbVMWm+6pLVHFMV3CUEoYrTNbO491YkJluBwowHxrmMY
efD1kdC1NMLu+HjksnnUMNHckedcSBLABIGbViV7ulcbjzOcRlmMwqcf2cIVXzP0
9HCtEprCTM7lWoMgeUt4bGWVhrjNzi3A8yi1V1f8LTx5V5CWVFThic53WGjxw8Lc
nXhRicNzJ+FzzKte25gQ8fcXBkruMebJlm9KzvIXiU+OyH5qtSvAsEl0nq92rL+E
ZWkv65weX5O1QFd5HTqTCIYjcPdknpyHWEXo/Qv1iLK6qO9UgvpqxVAXOV7ivJcP
5YTKZEtJnz9I1g0j8cIqeeHckPBg3qid8XR62spZMP2zf3mB8eOnJyjYKuGCSd5+
3emRLJagMPzVzfWOmvjrR/DdzEJEyiBBkYOGtyOrKuHIZNUpVpxUQOkGlXSjUEZ4
6teSw+2MBjtLh/+iR3HaG6lWL34Nd2FNOqLOKzrKVNrefxCXwKkHbkmISj0XjzB/
c3CrYFtgQxij1s9dmEEII4bmoS3dXbJXid+SPXlcvK50nKNPWsZtaWqi0ufVo0on
O2X/n830qYqTWZFn6VMRFq5GImE8Cne54vG+sdU618AEnFbY4Iuo5eC4K2iJHU5k
dGQ+gYJblEHbffss+DX38zCioFqLdn3OHgqZ940eKUASlRVYNuQaK1pxdVSiEMfI
5bNfZ3LYoiv3wUMkj/YwWjt/ofztipfakxRZWppCYvB5jKAe/lm48AGrm01T3dH4
R3KYcCB4f0EvXJEZIG6/yxdzqCnHuarqgbbjL7JysZSRwN2ptVaoB6Rp3ob/+EIq
fENSWBitxQg+AZO4v1HGtWTMRN+LuyNhtwsCjvlyS4m1WrD0cnV5KJ8JGfdM2CBc
IwIU7SDyfEnNcv6rE1YEah2jyEuGNYzeW92TEo7hlPNEApKzJTO+gjsXIUOpGRc5
+/tuu6X8GiLgmWCgJ6xScoPDJGeooI3aaxvNJLj8okM7hkALnqXdR/ApQHuV3z1x
xNMHzrn+oBOToLCDJH7lIWUZF4FYG7we4/ZzjluvGEX6S+txTiKUkne7NhPGWIfU
PGedHP856AcI4Nkm8hA9BUHOETVlzfSqADpfQHXYAxs+zDidmO3kWWKBcnaLa/wT
EAO/O2tjrOVoqgGCxiYoWUPDCg80FrQznPqd2iRlo3k3YkVoB4m/xfYtEn4pIclZ
UZ5n/UfWyeAdz7c7HMv31UeQOHj7CCc2f7RT47svsWC/45gUTSjMZGUe/GmygQi0
vss7g5GL54W0fmaRU3IKuzvsxLGk843CBokiehs+gssAJnAObeA9/ihevEaI9tjP
g/Zo4geoXbFE65BlKuenb/t8erOSXw+YgQZcZjW5y2rbPtPEBHb3Z+3kDctpztIb
N1Hl3B9XCb2VEt+BEwDNzThD6h4zZEp1FmhpYPGxVICvyvpeZ01UvF8t6aPCm3n/
Hj15ThqMoHFehQzrzVb02OVkrb00M6RcvMOgXK+K5GxraFjt4SA0Tv8S2uPbb1mx
xFn1lpkI7Yz+cWbAfHEj6IegxyBCrO5btSC65EepWtwUscysEkILdJTL6W5a8Met
a7g8tnOwwwKDzvtORYAXRgu13rQweBLaeYuMxzt5krkvog56BCkPjTTr0cB3T9x1
H/oTWsXiy6qiXvlGMBxSCvxQe6eKbZUO+r5qNtPAEEcyH4t9LDsIaXqjYkZkDNS6
/akUxodVnaAL5tD9C8zZ4nTgAYNCt/dgLUNZhtm5SAncHNmRXzPo6sCxr8RGUAtL
CMCuAwGqeFL3rqbdCi2vWsNsH1iNeSjteeOVUor7c/Y1+cYWQM9Etm9zUN/MpnMr
R//0hJdWnRRsSqelUlvj21enhc6++1ysl55F1amtO9soZxfi0Tn3Sf+V3AO/8Irt
8LWCRvowcmkATa9GaTO+RlOeWyfDaqIWw2TmOjUk4XdzH+UONfyGinXO6IplY/bi
4+mYJ7x8eRT42LETEZSVpJlSU4ajkDjzaOE0UQtHkOzncuAnCxIe9IWphwkSdFLh
ve7aY/wH0YCbUSnQTzQLUyFoeirIqEi31oLKvcIm4Bwhw/SueSJ31PZAskdGUqQl
2bO8OvURVut7QRFx7nPpH1F+mhvNTGLEBSxWP2yh87zIPvpI/aO26OU9rZMHdc/1
8jNkjNe5O6c8AhHSrc/LyxKLVFJhWGj8smgSaHotZ3LO2iWlWQCgmmsDnL8+axig
0PqdyfmtAi3fiiCOUTT0Ew5e6kHN6HNta3cKv/dTt5/cOIgF1R1inAdEJTQkRwV7
MCINePJ085gE8mMBVpx/TSFQ10mIcGb3sNJ9l37LNBHateqUuQEPAhQe9yqcp2RB
lxudaSBNXU70sZJUEkACmXZ0Qp6B2dVE4EKOWzzvU6hrIWgHr6MarBoWctPHCxsd
vl/+REEedDVe79YuKtfrJWY+KzBPolE08MEW2Pe15K8vk1uAw7pEEIOPMASNxEAP
lLdTH3+WLnAyZCy0nyJ4uyDfpjo+8sxhPkh0z+GBkPj6nRd6HGqq3TnJQ4l7+Y9u
P3MPeMyq9rN5M+P9N8AAtj7q10p/2nsVrYDcmw9xJlm3jF6FY3cAwkJ6hs2Og4t2
ev5wBKhh9Z7ZT/ETfVVQcTlrY9cX2M+3dRyw2HsDrX23ub/Y8tFHkzYHZqnyfUHZ
/DROsZy5aERhf8O8geUTfS1UhXJAH5qNcSQ2vzywastWWAh6ninbLWRBe8Hklv3J
9uja++VFgASqqHvRCUHhGB7hjY1xsioo+h/T2HyVucoNQ1dd+PqKjAYRqKcdZYvo
mh8LzbLEx4SIF9CImS+2+0LQmBrWpuqr3x2Yeu02WVAzhjbwg3sdx7pvoR9R1Smb
p6egizsnsPgBZMDsfar4cClOa2k0BtQC8SyeIxYg0QGupZz2LMFqG7q3YewKjrOb
5x2TWx6UazZtHZs7w4hb+8bdE09plfucPqL9WSx8hefiil5zGldb5EUt7Fg0f32a
QEhFeb5uFezdXES4sgfg8bR7cyOOa6HwWT7SWpFRNG+iLqczgJa9AAvpS0/uDebl
kBWEsspX57hKY4Ws2lAehNLa2zLw2m1mtUIIFmvpOpnVEZftX0m9blTUE6Dx/2Hr
Zhs0DgRVc2cPq2if+C9babiARpCAixc8nzKmm5o9FQBg50oxmWK2Xuvg2TvENQrM
o41X9/wOfvKc313oRRjn5Wto/PAgDWRzLdtJuWe0KzVk/FATO7JCtqIRZ/OPGfOm
FfW+BZ51FgSmh9X9qEmzek7VAD3Rn+Ttubuf74vRQTJDpqI37XAB/EZ7nyhXHeTd
o+wYWvp+nhyEL3AjEbf4YzpUsZ+Ga6fG6/e0V6TjYgCQIwPsYrFDREOBHQgcIlf1
cCXKGsK3OHbZceI/AkNbBupGGL5971EZaGa5SGLf1sxyXh9FKohT2vBRVCkl3On3
33DN57wi40Upx4bgOMQh11Zp5vj0ypdkcpOYqdSU8vKg7hN0JzeRCVOocf0sTUx2
QIogb4QFHlFNNN1ynE+Bz2mVnkWhmhivSKMZx492aGK9GIMClF94wC9+DiuHS+Uw
QItVQA5lZapthfaRezLJk8e2A8Z0uMlQ5dI5tAX5jOzyTTxWi0w95D6zgvS4S18Y
Rnw9tG2TA8d1V96OkhZDveAuNnS3Qt2lZm6kp4a41o6HDG+hjSiP4lv1tZcZTgL/
d9o3h4djROuy+sa+zFW+oA6ySH82UM6SnrfX+nn3Z3DxXL1O8jEYEp4IT9rxxo/e
x4v0N98n1YE1Pa/VCI5x0l9UFmXThMpOCfzdUtqi84X99JJNI0pVA5ZOitk5pOvz
fqN1vfCLLYkYMo/ciOnhVUlwj0AbY1emIKrXCVpxmWHpeDXTyaSL9kEwFYaP+dAj
vKECmj3BKqNe7Y/LQcpYa+DtpKlYwlmScGxmXA9j8iiQOfy1DPtdf6r+F5HAz08+
xml9d/3K4cENomzfYyjYhC8gI0ERCkRBeQ3m+3SdqjI34/2fhlYjLHQZShVy6Xa0
lsXmlbP2n/kGz0ERCAguatcuSnNj5lWEJPTU5Pm6IeDb9LrZywl2QDSOrLBcZVVq
scaar0V/lp67Affs5tJYQnR5E/sTMxPJLZmAuvU53J8Wqa4GCKgWqtrwVSWFSLHI
Jc136AGLBS+qYV6Y0tG+MprKuC4okzWJMMOc30pPAGcG9Tu90ha+1PUb3f2yPmu/
Ht3GH3AjsxqUJHjg82vRZSO6ducJsms4eRonbzhOkdznQipho7WlbXSM8/xoqrL1
4EL0s6gRexZ7GqQTxC3pT50tCURQFYp8jmZ/Id+mb/XYl+xMlzRn9ybPxFt7dbs9
XPmVwF9bJAwPj5bmMn0AURRwqBKcIVXivOyUQ7dz0cJwlvzlCH6dd/refSuHkvp4
1k6ItX3Vj0kbVV+aPRf8Q81Y1Vbrn9gfGS1zl0pU3qdIvjVDkvjLfP2xdLtm141S
MkwFR+2NbY5KYWLVqxzPRwKrcjAO8gQI6c8UcNJ2/moVZlhMePHK+16WER+dDQiv
HaHL7Dt+usNk5XJ/CDnUt1U+eNDG3Hny0glEGqbU4Xr25kxZuSthVk5nNoMtnkqp
u3dSL88RId5wXG9G9l0mjDa0FVme9sKUu7facSxvNp/5nBhlmU9wrrXeilN1XJQ9
LvY81MKSBqymHLcsTRfLuvnuol8RpdhpWWRxX0cozd+oh2o7N5ln8SvtezDZ7ePc
DvFNHyxcNXN6tsXNKuZ97Al/dp1hEyiWU4COitb2VazP9XUnJjigKYOM+qJHTwT1
LRM5P0762KSRcMCdgqxt7/e5A8bq2EnOP/C7RQgP2BwTJPmGl1klIoscxO96BlbL
c28d/ihqhJXZt/Q3OhFzbv7lwbjbP2vWxGr49ua0Al2PWsuEzeS82rDI3tITSR4z
+9UsWERagMz6FLk9xonLHk3m60kNTNKuydyNpWTkFbIoegXl2c/bqBW4Xq2SoX7z
YiD/9Ml8Kutb7ZqlZAHedfAxvN3H4Mp0Cz6LlUKjGcpz/HLrtt0zRlgwHe4NrAtJ
kKoI7vf8HTJlJaqHVl1tB/xFWWcma+JnyPNoPZ5q0wh0VOAgrpTDh6lSxbenY3WD
KtWL5o+zT8ZIQsOx88ClpNCKtt8YO3Zm0HnqKxpCXIitbZJhtpd7hOkm4wFF+eEe
sXPKfd63h12xtef7bbmlQNjr87nXbmlZDI4HEN1cn/D9ff4Ai04BRDV8BP42ySbU
dCgLmD8KnAgsJUZJbTG5LQrh3f1jjh8RYEfJA/pEGt5IUPZedeyi3xVw6WP3xYRd
0NV4tr8U61sBaP8IAAete06hY9uFDDhdJVM2/Npl6eyeMlLtzl2DSnFnf71C6zn/
bH3MBoOlVhdpmvPxrpLpu9rGCLvjCF8/iuawE9eBy9iYmtBfAtFO1PJXjTVfeXxK
lQAywtj6GmvJmPB2UccwAkHEE9vwuYpf9OOUvRFoGJIu91VepeUq43VnIliUNkEf
B/ctBU4M2NpBKBdyWtnTMLMnhmvYTnvcvPuTYhZQsq0ZfWsNEbAYswqWuP5VM16N
RM84vHqMiZp+ttWBk/fTVmfaU9or2/lX9/rV5nULo2Eluf6i3XvaUAFXST+gfVNM
spelE5TgbbCCv75xBGOZhdbfaw9euqwe2g066UikbeVULtQkowfjWb+xgMWjP/Fs
4FzeOfWak/eVy0tCb5mSR+HPbIJh24acJf8kmVteylhTQnbqGF15xX6BIHYx7Nc5
uvGL77oXU4XFp/e5rpmntyAjtHPy1pupzMT8zaw1y3jpwgWVTfPb/gIth3NYpLGR
A5VXS6ClcWBAVRz8irJER8kAs6vpai8hO97MCbBBaJrbjfXrmThI94fmBaKX/gsM
JI8MxpTrD9ZtyBr/wcrknCrAideJY/uxOV0l01tRaEz4V28qOkpmkA6Ya2IqWVJU
0cn0AN45S/HiJZv00kL2SnlKkV/+4wl1oeyqjI3jjaHF5ew8J3px6P93Uk2jmy2d
Oru0SMqEaPwNrQ5UStEGEvkeglZXF8mvHbkh7Z1Hva+aZyR4bX+05Fu8DavysaBb
lKeBLS33v2JrEB6BoRPpBssupqaUaYjtgCfq2LlGA6X5er+vF56iXDYTmDjXMWNT
g7+N76+ngAxEiP4TE1E2i1sLXBgKauI3hl7p4ZyMTJYfRxs1O8RfKkGLdfzE34f/
wLcIikvpjXZw4JdemM/hwMreBfAHmK6vvR87G2bD+uXyrrV5EEZtT8H45YelEaWl
UgqMuv64qVJ8a3xhxbDaM1gBkwkgU6vq+d8vHrOty+NxdmRVexTde9us8URnxVLA
aQSEYTfhbneP+OM4evRVwKpaNlf4F/ay+xB6XQZs5QsK4scVuLzP+U9hqrVpM8JR
SBPvQaZtxPsm70uRyNJWAwwg2uNf4aPUc0ecgqTLDiXOu2xzmvPFRdmIjtY2FwfR
++L0amVpUVLTbplvT9ReCCPIV+GuLh/NP9MI6tF2cT2k6EQJAnVfy907xibQxY5b
Yt0MkH0F/08KKmhx35gpeYvv3K9priDIdZeBl8ASb5ycuFmdX+OimkWq9uK6O1cf
hDPYMhzMimKONYrpwxcZ/DbT8ooVvkc6uoRKd/G0srovMMkxSpWEParc9yBsouGQ
5lMYBJNayCjYev0bQ+QHOqVDwxYcPx5KeCnGUBFRhfzXkNnSwr+L7PqiPAugDlH6
Eh31KTEDu0DNBDcvCFhT22ESJmO6fy5AomuNTOkQe5Fh+IYwLbznbeOE2IWIGbcS
UuZo5Vfg5d5YLnyii/eW3+sJzk3jRgFEzvRVy8ICw4SOCCd914n0rOqwjjZjiiw4
sBZOYeWBTmPQx3VjtQKE3dNcz5Dd5jesip3R0fN6LCdNi22XGLUFmSYhGgzPoiBY
NQQf2Dt2N1fRTlbICY1idyn4gYUKNK2sUoatsFrq8Gx5K9JoDOtZc/+JG9LpBjxI
ARUz62SMgEm9BUbUwc6mW/n5NhEx2sDNOEZTV6TvnnlWBJzIsdz2RJd4ZcnnfdrQ
uyq5rHJjbwWw3ey2i8pQ/SmlNdSrQ9z+aoV6D0c67QOWld8Y+7eabEDoqnNsixip
zy18ZeU9pT+U5KTBEDBzBBO+pW4O49PtxN71Rl4TFMpOnJcTa8wTf3X+mBV3cHNX
aKtdWYxu4PGhwbSTprmEM6+LocQkFivUSrJqpMqEC5MTyl+WBuxqSxmh3XQAHv2+
3CFEz94E3oaNPPVOMnoCAky49tVIuvnkzdamipvjJu7QuLTjXz/vP08z5cUs8RTt
8LGhAsiriNfdAK9Z0WEjtdMJ3Q7SL2xt5nBWhC8AiC4pCeVTo3wijZ36tzHqLM2Z
9Go3/0R2iJw7u9Hiqsui+5s/98l7A9+sSz5r5DsyxdPIM/0q9Dq96FqD4kl7d6RU
Og7zIdQ+iQ+SMRFLTpN3Gy8U0AyB3nmk7JSdRgv2/1Es5N6fi+9j30akXK3IBoiY
53cy4urliZv75J1ziLEncxKsysQkt7zFC+yzo9W4+gyhfHzxCGYbnP7PzQwdCFab
ildpvqXTkG7TK+GGY3y2dKyncLZtVuIDkLfMu5onffKxQUPnfPjGBktpQBwYxVRG
/rxZzO7jhOKC0LZ8WJdyp4/DIcmHtAqnRfqzo9PeNjCly3A3bDdNMpDflr758WWh
zvGl4SQpHs6KmANNywwduoRW8mpNklW11NYRV1vW+uxTF70oktfIhZD/wodK1HtE
5sNGsSe0YbhWvgXOMj6RXi4iXPnlFwIwe/ZisXFBLgsXzdm3vBnuSTFUd6x2d6vP
1XGH7ZpFt9URXiS4xJ+1zDeUKZ3zhmBWmVGBnMp5l7AkYVmiBhGIFMbG6ioQ4KMf
6zUrGlNA9AXLt7bQfJKi4uKT0vc84U+7I7v66WzOaNRwnmmi1fEFWBdCcT9SBymc
d8cHE2G0V/uf/I7e64PkhjPfVIeYrV3tyZ5SShcsPUrUbxIQJCnGjAP+3iP2N0Og
MW3+RpuVwPd66PFbS+Och9X2edxsiwkjtkaMmSkAEvHzVg+55kjCiY67A+VgjOzz
DsTpWeTJBBZVa+zxaDKg8HA3EP0JWFz02bc76B5G5bY1d9N0JElx43O4h2wIzCb/
HDZHAMbQ2EvbHp67eeYt2pbW76EeUyVvG47OSabL6k4iXV29LSqEK8bLZf+KwMQQ
mO5WELy3zMGn/N1ccmRUw0XBvQdGeuHcltBdSXReMC2J6VlIJ/XZHBLWfjy0hWFE
qINPTN2qMLjTevE2RU1u1OMV/fQ5jjHeaU9ie3DpCT2qYV44VX5kNrmJkrP9tzW0
vocRAXN/jHkoA5jB0YzJ2VIqrIVWUWBnFOIC5W+yxs534V6S9Xp33yFaNl28BPMx
PSMBhJe4lhqJQ4gtSSsMAsZ4QCV2AJhJYFbtEqg/zgbrvxXUWCIzs+AxJeTrVVGn
idbqhzlCJ2d59H6tOz08ZQ67PkgE+q8/L+ynWi1Tpkj7L7+v7jF2zQfV5vgrKnQ8
iGWK8umKvurZvQC31ebmA4k7zIuyTx4SibbEm5gIjFpBsRgxQ5uaWfSmGnOVorYg
SY/3cxOmWAd+A1WtXe+7l0FIFS14sNYMVNcbBDHGV+Nf0TG0XYxW7uC+ccEVzg/F
+bZyypReBRHSGYHxCtA/sf8W0VKrpBaH6oxWQMDQhhdVi2G/HoSMKIMcy755U9GY
HrUUtzRLIRUwTc80AI2NO9FAIst4l1In82PANUzqG0y4CD4KcvuFXOXUSd+qljRf
Q/e6/1+wmJIsWPBIq7j215/XzwweZU97cadFRzWpOzi6k0S0EpN/qEyJEiEDLbm9
9/DrMvZ1ovcwfSRml/CGfsJAvTHdB8QOZD7H7d63pVPcttYAenOSmJ2BsRTuYkiv
IUUAIigwR5UcS99hppMxG+BLlQyDd9WN0jcS3csBikn62/JXmCEc25nHLYEH3QPz
C2MyCGh/wuSOzplRvA+Yef0F3+rfwgibNM7eegbUgUmSaMtAYQdsjAvWlPHLCJdf
dS/d3BfIIhq0eNO02Xj5RDHmtVb9H9yoE0J06Ia5GkvW/syo7QQk/CJF3M9ZILJ8
blx4GOAbBWCMyWo4+zr00Cc+SIZHIiCFmj65amYGs0dIkm3asO1qcKdLx28aEXw9
Mp4+sSOgSeYu/F40SoSJ/UoIwWt7xYlnOaJDtmXg9EZfpdg6q+zu9uDhwQ9Zr/31
aKoOneIXnrWGqmkQq72NINt4vi8rOfTfb5LvNYpp4E8n9Ec8DyE+78ANU5gbn53r
jYQT92Os0uaYOiH3XvmOsmnd7tBans5R/QNKVrgQ13LlIQ09w2/DbiXWRsisea6n
GcW0C0v25JoRRZiLtJ5erDMQR1hfTIRDNe7wDP1z+erk2H7rb4j7Dbfxtj6XUMth
hP3S782ag445xFBD2dN2jS+XLr9+aFhlU6YXftaq2aUWON56eeoVAQx4TxmtdJX0
zqnUx3uGzEoAxEa5D44j0dk9rRZ7AsbJarAZRokSwFXMJ88Eqe+MhKqT3B0wF/BM
NS7iQBBPvJ2kceMObLx1FoZ12JWAVh5tJH8TglK4+ehT8uYBRI5tRI3Avm9ojIFK
IdsvIu9zR2Tug+X3knxSOLI/9lexb4Yw6nAB1kECJu0hA0/aCPbXjNa9RZWsetfY
BxptgLjTG1uPx7jU7Vj8pmMs1Er/UGCD3Aoer4wD12NMhCjKi97ZH/He56K5KpVH
lO8JlvWquhSoroxHkCll4Bu/t5gROUj6yxqynujpja56JYwWsLB+n7ra64LEhf8n
bjgsTugUbm2R4D7/qxq1aO+HTMFov+eaRkomduGvErgB7nMmsFBtjy4ZdjK4kxk8
4JcMl/Y/ZYQd7fbQ9YIoODI3JoeAkW2zOAZYwfHGepgQV+uE5i9M0mP4vTYN2JfY
35SYJM1DEZgq8hD1Qd1bu+5kgre0AXVfUS31L8x9nPZqGFUxlgmtO0SrGXvC9F9D
X9qJRk59bpopzb+QZ0ZeLbZav82GAXGci/QkZluUVyToBO1crP8Xz1sdhgeHiz1y
GEr62ReB7JrqHh3/Wr5x0fA0IBL5X9T+tJOTkbgL8PRbHCzgeAZfEf6MX4trD6wc
yIaNWAB0fCN97SXUqdtoPBC3x2tVvJUZqlKGnQjVlHy9EDbJHWwKnMzxg5NSHJtc
mTGUBMdM5ia6QcqN7qtbe1D+k7XXjEAvejP1HUyDOaJrJHHWPy/yc57RRW63ldEO
GxNQXKfCaSlGokCoS1+bHF7tTuha5DucVGzUhYx6BFsBB/vESCZ5DbW8yJdppy1+
dz9FIW3g5jePPgJNUvFCRAZSJrzAnLTkPwgElsCsYTa4aYdMU6RguP9IrI/Eh7s5
gVeNrreUzGllmVdeIWzgHbsgyWcDQzPIZwDvmx07cuV1sHCckHodPhulurzsQ0St
fvorlzqyhDo9A8XSSgJNbccZKhrSrCdZXzPetURksORoUxD+ToZ7myy+riXfvC8p
lD/KMC+GQqGmt8jpzPn+HBIZSP+fCvmOl0505pCNbczvWcGItK1qTw6mmRGkDqsM
8x9nFsax/mXV3jpscklIN6U0ztQw2eIv+7h+95s3i+eCu+5vFWeosKrwHf+UbOJk
BqB6seW0Jo/kVa5f5pc5BBj5Ynz/kh36TpiodJZ/Q/ua+6rglSpVFCErRChL9/8l
YPB77zSPhgD7F8cj8yDuzb0L4DB6Inz1XIt5SEWVuDnAxv+M1mWTu50NluyP+V9x
eaQtvi3FPGo69NoX+ER5fypoxXVSYa5tLxcwHpyZsHe/UPWcZPPai6UeG8tOu1Hw
sG/g5FekRFWpp9H5Rg41AEH3wB1XF/KzWAZTu7qz1taxhJwDKyfLai03Jpp88qMh
mIPbm4S+gzrrio4NK4+cwhn0+rZzAE4pD37dYyKC1qB8h0UmUmbgfZgqPaKV0Dm2
cqQKYM1EqB6iFViYRoW8NTGIgfD02Dj6gxLxfZUzQGVsXkycidVzYlDu8jafuu4C
yvjbK6OyHz1EsEDUxUA1XbX66C00ZTHrALsXFZWzh2BysVQm3VYKCiw6sueTVjwc
NNxDqpzWC2NANBUUS1xwv+enIJczzipYqIF5Owbjg5URyTug3V+mSo69MdBMX/2C
G076XWrUqX6eY2PZ9ClSwq5oMatqF5UbNbetGuhalMRNltTx8N4ioCROITS2J9cP
BbAbb3abBfFffd/Uf/XYuB6R0gLVg0LQvFSYCuu+F5QMJPLg/+UuEfxJ3uCacZYO
a9EGuVAU/oS8yZhhFjLpfrvXhcEwxNG183OROSTV2XeT1ZP3c+ycxI6qZc/Q/hGZ
CUly8s3bwh6gagYiT/tbWiGEuwsBq7TJpsjQ7jH3KV8fM9T2q1WiY7lCVrfrVNS/
gPS3Apb0/anlO4M6WKrgttxvyKb7z/jmIlQ+qRMvA3fz32iKS9t1/JDYGIkwfWdI
b1cSa1Ddc0qqnuggKgB8U9BuOW/5Oegy2X96kHfY9z60HyTnmxihE9YFNSMugV2+
Hy3FbMbqfSHGY4nLJ9YZpXEs4tp/el47aCZ8n4wqzwwK5PRXJDUmb+dGErlYeI/8
Vlxv6yPglIEgTsXZPmc1eB0Lwq9P66GaHXDW9batb9qy+3Li/wCD2WH+SAUCD7MA
z69n6BhFmH3+ErKPm/OXgLLm05Nm8Zx5BfZgzLkQd/EgZ/JyHmfnubW/4/0btRJz
mb+M2TUf6ef56D2ApoxYguH1uOJ8baQNntkOsNYK/ur0Lhb6zmGy2QuoF7cWRj2r
i8SDZaYv8u8r4WpMAgMf/cJHrspfLZXE+sGUHXzzBFbCdnxbVL0HR2HwT1NK2eJF
I/l2X3Gt1bIv5Xqhp7kt8SEJZbf8OCL64JCx0T/CnTJz4uWYvj6MIEE23W/4ktTU
XfQz9b0IDRdbEHmMlbtfrqrJ4LID0ORiNOpiiwKNX/ZwtFRsUe9rWUi5QCbATcN4
U9rf+VByWfc3NqtF3qbpidPj2/vY6gzhhwRSHt5gC8Igk41Ha9KnU5glXb49VDft
VhrM3EC2VNT5WCTEdDINc2xrl7h07WwmCoLuNRhcA4fU9PhXJxpeY8KlMDxNef4R
LMp4puP6rCg/O+meOdJ45sPOu6y3iKSOUoQUuQUJ5cCBSSRFg3sZS/pL94A5NZci
tyOgU4ciGO3UqDmNPNCwnsJfiMjx2h7YFGt4R/S2bXQeKU4O2o7UjTTzfd7olke2
9TdE5rrmX6VgJc9oIFqvGnqQgKmm0B8yuJGBh3RG1JLxPcNZolofdOOK5SHoDboW
8xRUKuYAHsnFHFVO6zoc2ZkYfUVjBODmYXcpZvvyKh4j94uf/SbDAGJ7XA9PomrT
iVlERMrm01VDQIr+GI6s/2WO78voM6HONAsifC+zO3Ep/Q2ZU2QfnfhQc68rUtzW
bS75boQhU8xrCWbIBVqEx+Z/j82sM5tcEpQmWCm7CokdSz3dfn0yQ/j6IdlVDQff
/NlYoqSxw5qkxmVw+1g3xGbMtTzAbLVCzls4NN0Z8BN0O5YICGmObsTHoas9Uy/4
OkY2ZGlZMcngZMfHoNtW6u5fj5xTB4kc/9Ket55OoXReX7eqmiB1EN39EHFcfove
VnlivdhPq7mNHx/rwSSA5ha5XTJrqrmijbus+qcOqHDNh0fGfx7ws6gE4FY2S9Ho
QUR/gulTvntJJuZczgHqgy/BbzTPgFgrn/39d09Ggv2yqeQb6xO2N2Lv/PngvNnQ
DoBgvWf1qb6D4kuG/TPoVm/A2Nqdm/7gwigKhVklukZGmhZOThg2VcWU45O01h4y
Gp3o3h7jex7diBcpPGkPrCYN3O2eQtIkkBxPg6mBBuVqbdMsUWzoBYjteZFGfJ/c
fg3k/glT3GcIJyv3aS1Adj0/IzCNGi1pdLCntkzFDy0qmI7RQZTwB3R/hllUPDw2
TLEtjOx9/ykMbRH5jEA7lz+8CjFamfoiyXTaFa2mFaGT8tkidNtiusPihKMMReKq
g9R15teuSD5OSNeb8NhU7K2yeJpSM8ndL79QookPc/gJXbZ7GGtmPRZJSbs+a7tF
7jxkgbOiwMNVfSOWrv3W7oDzsYCy22u/yT8h/an6qk6JCHFIj+9TnPkUAAF+ESJA
aH1Sy5wqNwROFgjs1WnF3QByhVfRPcAkbj6EpUR9orJqr8+niGlDmpfXA6qv442v
vuE00cMzAsEX/Hx5yljjONtltZuaOn8MUsYeUQNIMFqM5EbbdihqhDrOlIqNmzFD
udH+RX5fmzXu3XgCavie4ntlDzXtJ6zJaNOnr4awACroJMOoQuzZ+lZ5D0+2vKPV
fsft1KEJs8U/8Xr0oinHUVO9q8/AqN2m+TH74pm50ps1nz2y4eCqskWuR6MsavEA
w158zPnF4WzpV3q4wtY4KDITdyxtexZuX29k9V/xbA812pRA/a+Q9AaE5/t7dEdV
3twb2QaVbO+36rro+yrXhZAGkF3ThvwTFegoQexLLgXrH2FmhOBwL1IYsUmzJpQu
WKbwFEmHedZBA6owrclANtTpFk1nX463MgiQRDtZUgOYhzLi8jnYQGnp500lut5l
pnB603lscTp77jql/g8xPvlPskNnY8KgQWL2JkBmkd3FKb2logJeUCywqvBy1Yuj
Bo+6J+nrm0q4Ge+ekDI30/H4f3eoWaxOBNQu9sH7h7nK+KeNyiaaCBFxTl/czD14
zEXC4gSYDSFYRRV30aquR5K7iJYbVqBTCFkwCjSKq47IfaDWvaBktzrp1S0KV/ts
81DkCvE/UA4a7hLhDs12VDrTiOef5yhvu9XMExiz3BndtGBaVaejH8HpQ/jnW8Tp
/krDx2vdAEbCdoA9M6/TCcghFAYTFUrbqXGGIIZomYRhiYFLjrTooJEQDvY3FfSN
J3Gzj+N23KOcxnAzlN2vEXXnV6CQuxHLxhLt3FD63e1f1M2o4V0NQ608dkJC7KME
Eoz0XMLfmynDJqP/iNucK7/Jd9CaY+dVNCyxDjZrqIV2vWAdzBIi3tyl/5Id3Niy
EWkCesh5nNFGlCSHRatTOccJ/KeJ7tr4MeZ0D8jVxY1EPftg1T4mjsODvK8xduOO
TUZj6Tf/kAblKtnzVbp2jM47clRCT4IzcvQqGNcyg9iEUpIbOtX4V3K2LF5I6Crh
flllZfIpMstd5FmGD436e2AxpilGdGGaKW1iN7F2BlMx9gYs/0AlfzB9cWsvFnvb
vEWZRbbyUrbXIHfcW0fBdOAGb2F143SHq4MBz3fZh81JQuO3BDQsaGa7jRxMDAkM
YMkjcW7KQEkKtPb4MrloBaVMVrVUkcTIjlDTNAgWtRgIbEQMGnnJ0sDL6nLhpKzy
TwhsS31OsGwzIYjUHICu7WxVRIBDmplqv+hw/48RQbOcFG1W7s5XgUq4NSbOyHrI
+h6/z3vkf8FRDQRDkbMFpF4NdU/SMFS4aZnv3mKi48y7TPexzGgXM4hXtaMCmBwM
hm6VkPoNHeZlst+GrCrxG90RXGV39476z/PcWYgLyyKg79ZGO7OETdJ6C6kDfZEf
uTE/Z3aZNzhr+BuYZGAcq7lYfZo7QG0PuZDQJfYBzIprliBujciiwKCHA+cgJ046
4xeafRy37SlHBp3n/+jg9JkdAh2twPg2aLiEUEEL+12dAJoCEuryu3ALEQ98anIp
7D30JzoEPopWv7UT5DXqvR2luBOKNfLtN1kmQop3WM1nTaNrl4gcKqNjsH6hUsL3
oI1Zo9dkKT9JQT1Ej0IIAhx6ATLhDwD1vuZMNBgIdmN29fky0nHAt/6fMkUn86PN
m60AfJClvhVOnmNjmXkwKpVERdnAMavGhgxb5Ds9zPYqrL86oZtOg5sHWhSeelh+
cLzjJ97QL83Ta3iS6bxrOa9TraVSaC0+DlyhyBezrWhUoOauFMa5+RltTQoeqX25
Srkjz8GbjeYH5AtLpq/img79enbTNKX5NxyvxPgVIq1DFO8pdRX7qJS31oFVAc2w
klAKlbgeccRI6nuSS4P4X2LIJYqrp3OMxThutYIxgenGz/Eg3rvPlwGEc4RllM5J
sHrXG7WrmAUIakFDtSRtgcwnw2LDLshvl759EninSxWFqXC2zlvtYVgtEQYgY+ad
wqErG/Vurkn3l6bT+puzKaje/BmrzNSKq+k3eetaXHPUAKtjGrniStsUM0qb4mYR
P2MkgT0du1wNj2yQ+kkVpzT7tL1z5LOZgmP/XnNiAhMuMUyzvMP9mN/naT1KszZ1
hD+EbxO9Bm03NgJJXDeO9LOMP2UwGWtphMK/I7SJPfLfZzVJBYUUB5jMv/cIBR39
REePfnaOXWCHDekgF7KRE/hgbEvxmsOEJf3LPb5aB8krGgYUK1tI5HG6bC2wY6Lm
GJTYfh881md8sIHhTWvCGCvBk39Jw8S0UGs78+TR1pbitoR/UoqAoxOGYPcdZE94
7MlSYs4fPyuOcnLwJsGoavB1wYHxmQrG9Puqiw6dlZaTATija5jTok9NpINAqOJu
HT34s+vo0tQ3nYuV6zmW28O+USOdZdvM/x/a7PR2+YQz87ge9ZCZ9N6eivUvjPce
ILEdnGamkhT8LB4SKUmG6TEfdJ1afuD4DHzuYpxxDwEIS/6atA04Cyjbdo5gd89K
6sF4FTJ5JM6nrGelOIXlJJH1UW9tm+ggUv8cpVLqAJ/5kT1y4rPKLTWFGZJlQaC1
/vxMHWZYgR9Lqw1gBb8ZX6+Edb8gdwIlM5D5aVGLTuaPXcJosD06WlbqTMSt/vxd
j3f03+IUK5hbjC8U7A+yCBriBxmC0K0mvuEXGJt1lDJWcxAssZw8859YeefB4kKE
5Sx/Gu90fnlSmN6xU31+WKmoMOiqL3aFyPEVDtS2TTWlvX4mzWTJYeEAacYRnsxn
qqG5ofmsWo7CwGOKeMtxXHfbSjIp5duoVCVwrRJY4pgyLVdofcav/9cpIANZDobf
Zyr+8WVLbTV2vBr+mFZV7+y1lTRV3Jn0Dt2LYeAqN4qm2ukbPv3MZQlCeUVJyeSU
QOSfDrXYt28xRPxU3m0HrAoQ6MKs+WS9JUw6gXsn9AsUcpeC3N2zLc46wFvHIqmS
VHGS1LF64drXmiPZD5TlmVsWiB2W4r7D84jmZtwxAnoiCpar5LzrlEySXHgu8giN
ZkssUhCiuW3KuWRyfloqwPt81w/RpIgmuzWgCPlmAOk0tol89+N/RgtsWAAgGK9V
fYmOsx6TfVDVjx9AsB6HsEwJatylAbG3O5WpPTypVDxq7V3KPYw+9Zg6JueBfHCd
XyPo/gYszC6orcnBb506qriIDx9ruYO6O8JxbMTflbnD4uQzhgeIfRQrrYN8mHPp
m+KMBKcq1r7DE7wSPa4szDMAQBcc01a0B3rTAkeQZ6g2rqMeQRs4smJAlnsR9i72
eUdWSH8V0+C71SRt9D5WgW8U3W7sTJdBMCyI0W2pnu01BFZXuOwvrM40XTBBEumg
TogGpfOJ2jUH1RJKBPSKcBCvWygbyJz4au2WpwpUH/LclyN8bb+p1K09oy+BgMOF
tXV1xugoTTAzFTkEv1t7LlB+GQeyorD+Xx0o792vEnvCaxpkzdt62oqKpOhFGWaK
8njBx9q8unisV3TvyU1wCJZnAgjda73KuwRB+hvFncWud53hYq04AdMOjOGDQTCq
shElmMvx/zhJY0AuvTKUv8xHYY4GWHeFwLDZt82yA2nMxPH8mQArujV/RILJyRqM
ilgTqmOjGtGricC1vEJ+kRNfpznqkYZU77XNAowdMPBaC1hMvTbaEDvn8lyufr9y
AzlB4ad5A1zYkexXrzzbAuxAexIKwK0FpC6tOQAfNJnjYUn96E4zZwr8vmVJJZhe
WOV/oRfNWtSlPBGt9aOg/xvO/nA2YqWYQHW6vpzZjLNVYGYSsE+FE2UlNtaJXrcB
1AmQeA7lRw4wagZFb6mw0B+Tja7e/ElsgYmUybd+coWr1RwxosjXpzzwic1nLXOw
wIOie48VkEZfnNbijJY1KKXc7kf5lab0sJIXZpAd1vRq4kpNXWVBQ8AKEUvhZhyl
uihpyQmjrkfL8HOhkvs82K9RGLEvdXAZPLYBqR2psOCRKGR2SKc5/R0wBrQXmu8/
Ko70TmPo3Hf2gfX7f7sYYZHfNw/23+tCiMkvMN6ALULCKZLZojUKq5AWBvxOTea/
M+hLfWd5RMDg6nVGok501z+1UQ5p9nYEDAy9W5J2rYkF/apOLEdS5wp3BhYeXRtW
F9ddFkl+7dRgcaFEyKN8qFAH3PGxCNWSP5JFcOI28GG0nDnzkWchucMvJauy98/S
S/XpqcDwCi+E6i94Em24j/2L5sICYvRskq/HSuDQ9r2JhgoxAr6iuc1usBcRopKC
MGFnRFKpK164yXp/MkE42I1rxScgidpaC/GbukpY5q9SQT0ZRFEbq4wHWeyyGTup
cYYr9KlvF1nc5usMHMKRxa3PJ2WLYsX6AEmcrSPjoK0O/m6c3y500/+ZgG3vVKGd
H/8eq2zjENBH12NB/E/lZOMp/mYseL60f3/6dwPrA3ipfkTxMLeCOGJbIpI+MLaP
LysyjuoElrqkCRkxfMnnn3LGdJ/aSGOOstVU9Q5wNsoDdxZWQhlfoAmMTL1FNCRx
6pokqVODi59DKUq5ov4x5f3XA3h6f31x7OqvwU71HoT/Nf14gGE2hyuDI0b/18JV
LhzwO2G6nGkBiDzohvSgO/Bfk3tag6iGu0MCnbt2nCXaxjs5a0nM3LjTHh1gkB1q
ht4rHmVVxhc70jruWXAQh8irIT2aKUunGhloiZ8xD6xPsLbAWvUFpo7ASSI3H1MB
fVBYVc0HIBqQorPbzt4/yMativAxPKnM7zZXsUMfMgll1zgj/kcRcMozmGInnXBc
CuZL1MNDUXpieqzI8QC0FBvXb3nVCuxFH0e1sOE/cM37oY0OVmYIfi9rfYaFJOQZ
hXyiEUwKfIUsgtjYn83fOypAfS3rXz31x65A5Y6Wj9nPHHCRrueSUZCOrM6xB14B
fwornPWoOCTDDMGG4B/MpVFSo4ybR47rVOPu4otM2Vr3venJimx0QIEiWmEYEctS
ORFzsJwPeZXmUP4UL4GtKxWEt3OZ7TGmLRHdyGQ57OXSDgdsJzhLq3vDaPiRLxNl
pHgsv415t+Cc5AxGpQXvmlwi8AJhK0vFPksMtMG8KRRGqNoFmTzSpcSe2eLNygbT
VQNCtERfpebYHZ/m8PcAAQqKKdS5PdmyQO3SdcBL/nPU4PG3odFEnh3DwEntRNdj
9/FMxBfa9TvMg1Xy/4NhQIf0HNx2+GRBaEPG1WtxTGwhlnQuIXlFX7Ui0ItZwn4Q
iyihrKXbHh5VWjLkBGHWE9S63HLSrVlxQAEuDWtZdm6DfTDBO1dIMqEXX1MWWgjs
rddSPnr+t4WXGDUvynuxBftqRth+A+I9spoTkkeNggrAnpTB4+kbXYwmCcUilgq3
lKfH1Rs9hE9CDBrr/6CFqnGQxLarqWadWaD7KTsOx7krMX9B4Kt9zOe1FYVebo9G
j8+/8YgY8znQm27iaE0Rg9pv5DfyvvukLdJj+iKjw40M5j8hV2OmebKNTuzmUQXQ
+Gw257hPBDHqKIqRQLFqQmJDvthG5CaIifY96Q+V1iMfzBwqHO6K6xQttCfpHxPP
uee/VHLq7PrYN6VNBfVEmJCnYqh+ECUDd8IOgasQp8S1/bT4uxi455wFUDDIvY9v
LzrGiPYJOoNh7JxjRLxYDLqD8+/b5s0kj07IaaLMq6rkt+BnJAba7e88lcx2S60o
rbNFFc58okBm0mx2sdcaYqCdxPOCNqiivb17i1OawxOYKGRavQuAvE71WmAuVqUB
Q8qaO16rPvpo7PpFaMSxuUo1FZXxqW3tWHm5XzsUOErF/DK+avQWeTfr+rauN46r
VyhPSD9M5lHT9X7xgL5tbgtXZJiXxOaDzVgvqCiEQ79dJDxXtdT2ljrMESO5xmvg
MHN3yjlsBDSvqKGsVRIqznfn+OD1GHpKFxBoTo9lQulCMPfufBr54+GtcX7zu+m4
S3BRTUu4tqwR2Ny9LB8ITR0MGru7vurje0v2AEPgjAGOoIE+ihvHT8aWnQtZXLkl
VXpYGl7VV9hZPw9wnJoYeLp1gMN2+RkpStSeHPjWSSInikKEiMNnQ/6mU0vfnzuo
eAumJnkjg2Mdg69ijh/FpNULKRggZWYv+mYxpJGsnSHmgTIhl0ptDN9m7EpS13J9
JVjCcQe4aoiCT+6Z5FlLq1yG0/vuHzM0HqLrbTUIesf6e50kmcOQ63pKrDweXOx6
Yn+CRPbWOZTyQxjMus+h03w+Gg4b3eU8OkBHXGS/asremkwQ+Pp900zXG5JVTddp
ynHOysOV+xZwWyQowFV1uqvvxMNrq118gI2IQ2SYx2yvY3iLYHwKVXLjLuxsxbZ6
1lj/pSptxrS3EMkMvTyYhYOwK1Iq8An2TLyFCUdivC24/Z0sjdpevA2ZDPa1KS1M
KKxaOsHVQUqUyUEAu8AE91szGqQs2NXGRUn1UGIIR//FATFGeh+922hkNf1BcQk7
QfBpP6vCGkjD9f7IphgiZ1wDFx+Tj2qMJyuCEtZ8F+VVCpBlZh/84ZeRdWVIRLeg
mAIzlbk6yGBxqiwJqY+a1mfgI2EkujVB2sLlFGealcz3YQTmdZZUl4PRs5Z3UuRp
EXxToVIPA3U0LV4cpnWKmNRugnHrDslGvI9xD6OTDYLGEmjsepjkUTQ+GTTGIpPu
Aed0Xvk3qTbqEaOmV8xJYg42OpWewIBWHFu8jMNkmSTYyS6IPt3C/pmv/NFwSS3f
W2Qvka96TjBxYqNLXz6lig9ITlKKMoHgM2Ser/ejN+igpt/QEoidtjTii2JJ/1mK
HGatfnPbwWoLCL9BHvasizobvYLeQCDyK95uS/ErgG+1mMgA/HeMyEBvCDkxktDV
d2fDaC4dLDfak0SW0FN2AdoaJSirwnhzt9a6BlCY0c1WgFJOz5jSOTbR9ffrK4JO
JBpbilPNItldgPI4itUi1q/ihgFJkPTyZUEqVttqxAPzh+tMRtpeF36oXQ9FZ66W
7L8ehom78zhy/MJ/mvJAlJrnIGRAawptdZXdDatlz3PIH8pmsiNqIioju0yldyJZ
tKQBftq5APRdlDPzwGZ0IKBGk+spLt/3eElpeIycBY3JywywqhOQVkEqqg5dwlEk
AoRM07RdA+mtUFSqSj55yXGjHVHPEIb3cZMskeuK10YjXV1JkO+sD8v+SOP/31Rr
tDu33xdPemjVW6WJUi3EJTCosO+gzu2M8j7E/uH7t8QMRm+7e41pJZh6REa6BVEc
/9HQu/e5M5QTP9VU5sh7PRLw4hFGhaBnaMspru+MpBEWIEx/7W7qtaBFvuCQbeEB
YUcdiQvUHr/DpbtsJG20uwsYY67cnXjcWCnHGDojAzSBMxLgKCg3fD/jUp0CgBGo
AkH9FNhinmjX8+aN6fnNRHDMrp9H6HhjPILK9SSn+bngeJbb0fzt4Yosmznb6tlx
j3kgh0DEOgWIf6DsVNb9mBwTETTO/Nar1qqYir6ggn0EPA+x+9/8WQA/WHj+aH/w
yYQl4cyEHG7xKtj0ms+oWiU8gwyQfrckTnuS/kuMa2Zj/qY85Yq1KGRFEBa/WF90
B+JaIPYI5tJBZ091TtEC5UQjZdd+ArI/dNMfQ/V3i7l4nbdgFr3683vgiyZsFe1k
9zTlR4SqY8qjSA2LZYtEipyeK7YsWyx4rCdOpRfMQEVFdLpOXN+IhKEERReMYlqB
6xmHG6IbYT0lfwDPp49ZgNcC3zw3TVmW2+f66Yt0HCFtqL5+scJ9lP6T2QhoiGNt
bOm2wNGh82OQe1qTEBhBnBvr6X+MXpEtJRtpjw17xT1CTNvqjWnb+dpvtVw6DUGx
gV9RAq8p6tQ765L4cGkuNBi5qzANmq+Ca6/o5oNZPICBSorWnRePPtwxoz6d/UeB
ILJU5avDt6yFGrLX5V1dEagjpvrrr0KhV7U2I42ZvtUehcsBVh/r2w0uj50l8ERr
xAs+cgpIeFBo6jSoLflROVksgjn4z1nCGR5coHpmulCljm8NlyTq4uAeDbUyqz+Y
N/aY1bb3jtR6Rp8/DRgoO9xsqRvgX/2q3HlPqMB3mZ+Qw/W8YevXvcHWBZX1nlTD
L6/y5toxZfzUEkozPYbP1Qm1N53LhWarRdHG2HiSmbhPUcXJ2ShUqEW3BcWO6TM/
McyE3f0HQZdJUQpN6P2yd/L7DqRlnZuj+O5VvoR3kQxCy6oCuIk/uODLW8rSCxJk
V7XhGqM+KVtv35mi5anZmBYSG1if38XT6XjYRmG6P6Od7E8Hf7itVU2crua/c5hg
UY8F9Ri8xbr51uE5/89djRKKwqbNeO+jPiEPQ/zy8dx1QM2W3cHBoghLfRRVq+v2
vfcOqfXynozUeRukCCvuxQifPOBhYVbDCiG4w3tpvBx6R00vqImhEZYErObbzYEp
FQpLV3iwaJRBTcfEbgBD1w8bhU869QsluZpAqu89nY4iBpNI6q6Yy5lXb88vbz+u
FnHnKuRHheDT0H5YQvqu2hXZyo7nTcaK8IwctiGg7aPdE4oBXe2Otgz7vHSmb/ny
TG+n/012x45m57/i4MG9r/vZ5wcu9ui5LKEJ8obsUdi/3qZJK5mlYQsxZQdQCu4F
aS0DkuYo2dMqqg09JiiWVDm+r3bohdUxrXR/4SlKbDgKTkJUABz1jy6uZL8mhbfZ
0irWORXIL92D3tjOv3xQ9lsMQt5BQ0vFiIZTVXrgVcFnh/iAUPES/9cNvLI76UyQ
txR5tM/U/yPMbThAL8asw38JU6Tfx8EOJtdQmhdgUkEjaTWRE0eaNSpznpk4BDtS
v+0m4sK3RWXf4/6LikmRWzA4x+8g4Lqm3Sc4ZG+DR+Q/RIwm8ZQiQ7mOxTOOP9kV
wa01S5U8Tn2gA8TCTm8xvCDFDyq6uCzm/tdpUA0py2k2Hlu1U+gYWbIBcEyNT1fL
iFoMniqlmtyo20jkqSzhng+JnwqnkS+dgDZZ/gVcJL4V//SP1f6xCmcCgu5UBxMd
6P8/SSOCv+o88WJD+g9O5YzqiN/mMk4bob4jQg4THc8L3F6RndVoW8jEKTD5BpYq
kULPOP/EHMLcomMUZxGcwKL6a9UcUNhk4lyL8SqMw+Gt8s6xJmf0eCTzEGTPZ1wi
A4lBaL2j8zyIH9KRuhidmuw4F11WD/xY5fNuiTV1mdcl65E5llaUaBuoZj+qa07H
OyYzFfXItRonEtv4tX3354mArKoCurqOnxyLrJ28YPcRH/snqLfRgHlXn5mYpTyp
7isxC18GuYNgk3oHAzd5GNL4GSCMtU0j+vlSq+EgfQ7M1ecTR3y/xjhAYL9yXWou
bC45K6bd4sofH9D/oAYaSqAD4jlzFL7AwlKYxhT3elQi1+kgk2FDiGAOjKlBrkUQ
oeM2t8ZymIAGKROnCu3vD07gnmAMglRuKXWSR6drABxt0RUvejrWInZZA9S7oOt4
dg0ovKb9OGcq9M+qfD9QXDJcR3WulAdDPFWog+2CiTWi912/HU0AOWpMR5R2/lwa
GC5fq31960TxwzbcKa+dy8/S6lrKoWP48VATq90+1iY7jv/NUnThgMMmdEVGunJh
h982o/B7BsyYThUChIAXsppdMY8SgrOuhTFFElCm5Enkxlvez9uSvZ9u8gIt0sPE
MY0j+fOm9gJSVjWlCu5Fu61TeSSQujtKCuEBwSfurEusBJY5nFyDww87jEfK1XBj
d2ZR7tFndFy6qa3NlqgDMZ1AeOTdUjA8YfHQxy09TMAed4IZKUF7szY2XtV2RBrP
eW16xrDELpHsCSgxLJ0K4XFD3Oq7tH4IgkQyueP9Ks7COjzwhyWUL1sijtnSGzqN
34GNeD94r43rGimWWSf2ZaCv47SFR+IGCL/7g8/rKs6PlY152eW3WvjFY4clckL1
o1RShjcWAiBas3Ja90lvHGlrsQ0yEXFlQVh0iz7GpIxUGc++qZI+yoEvd26iHLtQ
YWsV40iC0W6PkNABen3mFWYUW6ufm5rBQ+CMsqX+5EdFJCT0gFzAXCva3u2+IKa3
Ahoj5n3IVw9kCHGd2t0y2kjooQL6nK3o+bRc53QCGzQnmIBn+hBkerMSpBXTWpFY
EOEoo1GvtV7gCglR0WzLYIMzZq7bicY3UU4+46cwlvvFJBjaLxCsv6cPqimMQmmA
XfXHXoe+ur2bTGJQK4OH3SG15Xx31nzb2aNk/nLFlTxdnguuEoa8GPCY2OPSBAN5
++XvZBrNou51PP2M9Dfffpb3hD/iTzP5nylk2I2FVPXG1+H45bVx5El8OtNxlJSP
4nIicIeZ9rLqX7pZpL5SbYfKDApvwc/sobdjFrR7O1KB8mqztvPNBgnso91k1aXL
mPqqb2/j1gfXkv+LhXO4C2arUntwEaKxMcmYNAcs6SV2mE4geRypQQ0yJojJfwjZ
DtGugtJ3Bcf0QptxitamgfVOH3oCPw0pi5Ho2zmMvZGdZ+iXyclqgLBFjw726/Y9
ZpYr/PZ/W3hgqoOpYCWir+kS3sI60TaYQV3wCe7h7zz+C52pHN2o1yMpceVUU+rX
EJ7QmYq8XjBr61U8q+oOJqMT66/Qgdhb2AjoaOTwOpUxv5Mf9wR5b+rUq1wr3Ld9
yVD1elzrFO5O5knXvb0R9emCKcUlfQptrROfNStRsp6l4z4fu8u3uSQTIa6iRW/l
X2NxEvNC98bwC+vLI8fEkjw0bCPwaBbbeQFnyQPbk5hPUjimFp3LllzNbd6erhGf
Q9AYjnu+K/lbJ4C3Cq7rAL3Vdg4OcPWNBvBJLYRihvjIt+bjCnORhb47DqDkaEkG
fOHZpgbimsqeGzpKF39V88Lg4urO1DeZ3vucqYu+RuyVueMI1Y/8WufyPrxJwI4V
6GusyZYHjLtUwA2BwCOCdc3DRr0QsNaAE67Tyvl3EAbQoV7FtPsK8xobb2I/u/8s
ZVofLMIrKW+TZIUqstQB6APT10Lr8JGKjdFpgsVLgwkC7OEUMcPZHMVyENnoZboG
IH4CBifF7GM3GOL5bTsIK/09/fa+RJDvpFjTPQ/pAFOfYtclWJJbtugyfIaRGgJp
bvBxBDZ1yhRqM//IqyefLdj9NeKrLdcEOJp+JpezjCvITfaDq+6qKA0dSbiY2Yzl
WWbHQInGYj8R2fcyL4QYO4y38Fc1qKHJkE+7A6w3puN+bVRLTGz0z9eawyTuDfa5
bQXA+Chrenv0q5f6O8Vg88oWOGZWJMsaKYcVA0cwxRm5aAzagMhrH3weruCaF/+Z
WWJc1TJOEi39cjIcsh72xwdaA0kJcLUTXLL94koFC4skCb8u5AJdMRZA9NYQbbVZ
M0b7BJ/R8uTB0hoINW31wMW8uWbDvFTJfLdRrMmynB2/vFKAgedT5OW4fobXbzVJ
UUfT7102hZfTjekau943jHKRIwNRNkw7Q723nxY8+rT5ETZnByrot0ar6hkh47mD
2zijZuUDQJffUXlRbS6bEOzKUc+MIWI3rNn14lUJ2WNYo1c1ypAWp+vsPB6FIWip
Kf/oRzzPrlCy8bg0M/XunkosSMP2tAqTYPjezALyMuTuVkVTuKXkyzpg7OHe2fn6
7OY+68sU/phLLxLw9PKl8niiae/E8d/N0bfVwTtQGVVJaQ08BpVCDrh83qPXz3Ub
nvNNOYGwlXcB3/nc+9z02DYrSI6GncYAOP0row4ZLX4Klfclh0Fu/ELs1prXAqDm
KQO6AaFsJG0kxETGBtdOXLnYySG2IaUMRs8JR0XHFXlmrJvcdGmXdM7ZGZaEZWPZ
+FPo6R5d9KQdDZSp8r6i0MZcpgTHjmlR20nxIq2TKkvvB+ouZHuXwzY83bldT7CH
OVvjsyAJZHmEPbvZwKMeBWybEFSYwXQRgZbVIPT7YsKRgcHepoC1udfvs/dL+hRX
8wOUrXyysPw+RjrH2GTgCaexWsFXhJEOLIw/TN/0To5bMSq738pqwjCsP8Nm/Gr7
8id8vLTp9JPmtuKqhkvNP5RFS3UmS3JwelsCjwNzPlGcg2myn1HaWUwYjugeDpoG
zDHzQi1FYOnqyad5gbRHWim8jYL6A6U3uVqzO+Uc5rhG2ZeeTiQvxUciQiPWMEpO
/AKepeECnKyIK6BGwLccgZu4d56SwJ/MNF9hosp+mkLmUu2vt+rAXGGhEB1xQjoE
1Zqlxrufkmmau9WemeGgwDkS/DB2bxFV4fx0JkM5ODqwvRK32q8yg13jDfGll8+t
I8ujzolPe53c35wEp5+TFvex3CkKkPsRUbtuX2gzJFqF3LGmXa+rQE+Ar7CT2dxw
XmM9clgKxSNszHvhhFYZxvNcWkr+kRjeBXoN/fvYazzc5ufRtqIwjWkJ1W1Jifs3
w9aZ5codG6ql78by5zUMZ3xKE0I4YI4CZXgNhPRMLnT6yK7RlpRxly1TNIqZAFmK
KLJZ3Ktuc2cXERyUPMFJ+GZKgc5dTWvVec0CQcAlvug1oD6+FzNohknxVaREVBJ6
QL+KmZ/Ip15eODpcGgPaMKataAJuw25XI4egkm6bw9c0jRN7rms9O8IAxm+/t1m8
4wyH9CJaOkLc84ctag860zKquSXUg/sAFMMLakoeJauRbpdiDFEtDF+bw/nhGKNA
AttproSwsbfQZmtcN3klXbjpVjrBvXFeoHl9QxHTO5H2yIUvWsa4yUqB6O8hyTa+
o0bv6DNk4eVX9ve4e0Dbq/ZhyzEyhK9vOHL+FD8nxBEEonGYRM+QKcjvM7HfmJqT
2svW3GT5xqDMPcNKX1YG/D7olqRNJmcU1NR/zvt+7kDRnaJkJOJvO80NwlwWiEh/
UaHB4tNOLRJ1JsXMlRgJ4ILwIS8rgSuQbMTyKzpH+Jdw16Y8V+IQYcbxanlcxT52
EklO9jZuce0pa63ZF8lEW+UAF1MRysFhDPS3xcXos6pJwobNI9aNjWQ4ovnWyXPv
EBbqwUahAdhA0zHuzcrDdbm2TUyz4dnJY2DKoN3sh/xeSnn0VickPGVkO8LuR9My
8MA7YpuRk7BmtIzPPm/4wHkeWHdhm0QsBGnnSiGtXmB8ss5w+nAxCOkkX24xcp1y
k3+Rn+aFyi2o87wDuNga/Mn0Q2hlVQPtGaNg4LGoqSFhEPbIUlepyGetundVbqAp
qCSz08l8YugYRsSfjPwCuyc4A7igssy7ookt8tcowaGrYDDoJdMxJrjHSJrcrNrZ
htGZ89y1WA2IAIadV4CGzv7o+JT0LE4Mw2X2WUtJKMjVOU3XGI0/8YC/A04UeE5P
i396oCINJKaq85Y5Os50ZWeY69adX32yC70E32gJYt2abnYNjSYsW0XJ90n4GInc
rKHWhngr9+C+9/u1IomRX9w6ii79YY2Bcq0zWEyVZhlEbKW5VXmjb4J1QBfwtGO8
RJrYXVdhqaDaQ8kzklFbbdpAl338Q9idG0h19RzJoDIuBWY4Sdcmjz7yVbE7zpHr
TSDU+Bj7YQklOTXxsLzBF2eYktPgLhE/hBQmN8Qu5ZDC75b2A2CXdOWMndbrg4n3
06nZeIETcCXNq2HJdukpavzSXypF9suqIXZEPTcJFuwrBDui8bfLmIMA91sP/fDh
Cbp5SGfQ5z/j+vzPwpExW9Bf8UbvyaXxRdpU2U+FOeep0F840mUf6SzzBQt+GU2c
hv8Z6rPOHZbQilHI/cwUXSZbqkuyyiZ2si3OwpIvQsOvhO8moRP7oMyyKt3ueMg2
AvJ2xKNudIKO8F93JjuVjwfTwH1cxV2Iezl2RnbwvlCLOA2ll9h3UFs8W+2CrKC/
/OH8robUsKg8Tw8uM1gqS9y3b64JZOjmtzwDivVUaOsQR60jAJx0ebP02FB6k4ej
/yvxv+bOb92NTjoUe6OB2ivzCX4Bw/sWxIEizL5qaM2JA2uPJYmtf0Tg6We6nVBC
XwcUwzBYB0uzQwpcnCBdXWzzdO3FY7kYZYCE8+JIY3d7kiL6onSQG0RknFmZSPLY
7THACv5ubvYA02XoN0rKIN0+JSoAPClhPUPqozSlsCVXhd7MF8O9szQNSga75w8K
qaqsxORvrZvSU1TKXQrfxENDYMZjAO3NjY62FWNWpCMHeFhl2Pkp07XfSbS1AHZx
cBfoqHf5Wuih38bgmAoer8GqacnUuwDCxTSiR92gJQyrgWafTxUr8OpMDET9m8Qn
pl7qfno1x6+D+u0BHmRhIm/rOZHZGeXCXdyBgOcu+Yqru2d68ZnmBVu6ctxoFGsy
qi6atrly7z8gBvkXI9zGcsrP69VkDlBobJydV/5EQUHd7e9av8M7q/eTgF4yjyxA
rcYj/ey5M5IcTDn/vCnwHcP26Vxr/3yZ6Bo6QKcH/XVkzyJDr616C3oI4vFtmmVJ
4JkZcqhz4olj9tLiTQh0GxsMWjzQfpgbBuy7R4D/KLmLbZkAa6wyyR8RrEEGS0yU
mBotfGdS2kT27sloHSg9/eBbQOuPbWXCLuVkGPOnNZSiBpb5zZFA9bLajA/a4k70
01ferEXopSvjfP/p8AdXDeAB9XSZh8X5eavOGaSSxWdQ0AlN5pnAo7LtCxTI92BQ
ytbQZcERiKEkliCa1Eg+9vtntkeBzPhj90kwVei2onUnkRhPsFSVhHddNWk2lWsc
M3mZRYP1j/kdij5kihMaF9PeYpIz97KgAu2JP7ImUhODcm61Yr3aosHHy3kN4gN9
/5HY0O8RiPyvmX0MEzV6+GrrIHXhuia1diMotl7loX8oZayDdavPmq2fos1an2t5
SqEvNS47isGUwN6XYkbp5Sqcw/lVjQmhvqdJmJcOZVYQPcN46fgpsv6orVNfUBz0
8twwkfNxbz2gCWTsVYUSg4pSovvykSuZiufjlyqiUp9xsQ4qHMUYXHOtXTn0iwCI
RnN8ZUa1xskMci9b7Yauv/Z4DWeq1PUraPNyOse6lS5p3lcUr4nXnRv4APA+XpXU
BnyB8Zge8T3YY6aY1KgfDWGXKSm2lsLAwAtLV+pPKj+WNYQYafmKZoxM/yCJLHhg
nZro3K2FjtJH8vRdrhNo10F/NzwtdWhtn/7APLMNM+V3tg23LctoUxBngxGdsAhb
Sq4jHTchAwHmnjrSzkzwErstEi7/n6f7TwDlZrWCvQ7TgOdbHKO5s0+vVwjIvRhO
ykAKzOB3z3Owl5qH8crjhqzRQkyGvZ1WQ6E/c675ZHtT3/0c3RGCJF6whC0McEK/
u9VPgTW14hQHIFCHSzn/rM5l+POrPiig9fy9nts9Ok3bOFHg325+xTdv972oqaIC
xniM7SGaIXVaCOL80uiiPegmdKMywL9GJya85RT/ZIk+9ethGPz0zfDE1G0i2L9h
LZyxz1DaeoBTVoTqQs4jx4qZ23pnYBvvU3bXD2ycL4V9PLgHsgnf5Nu/CQdqHdc5
8yXkCCL2qoBvms1DjajOneWR+cpecuMi28fZyxB8q5l0UbMXmn0esmZzFw4ikjiv
8oL0ZLe2WVQvBddMGwuetyOL1dzCb7dyv/pkkpj2ePgGqPwOotpyiKTobQUlrftk
CVmzosYw+X2CVmImYmFC7DrhqP83Xw25ny6PhfwKnVulgE2pT8PPprKcvl23O6qA
OnwwSM2VKkrOHV0G3kcU/Hecdzp0ukr04doQhHfO/+RSPi1XczZCknLbhcSfeQJP
UsBetdOMEetuU9xj2XpCLokGD0i+/kHgCh1nSDLvSoRBQrWFid6iujbaIhJBmeUI
sYHdVObD5/L4wu9OW9Ohuk/CRhKeSptYPNSIpvyzZqgwQx2hOmeIszg6RuIl9ftm
jD5aL2M5KWwv1T6PVgRNZ4aVZ3hh6iBG+cN1bCodd/P+Flm3zJeUWnFj/LvqJmTP
4US9XBweXUEpx4mpi8vvvfLWapFJ9ebrIRi2PezlqNMCsDJ0LxveEkI7Jxrwf9Jk
peZnzmkG8/7JevBCrYbki0JumC+F3yhg6TGKR4hYVArKKx9JYQY5XVIq9mKEmnSR
ECnsbuRcV4xqTGV5kgTLimWlGXXs7u+WR1mdg3jGeZyhRnVnFnFK2G/rghMyYWif
6pfuJXKhSX9jYkjITCXngv7t/Lmum1wmje6wuGf9LDnQPlOMYHZlO59es54E+SmY
5xvJL4wdW9HjLaU9rZxk0sEXNtgEbovkFRZdgjX04fNeXzpVmnPaTZvNkeZMU5BG
DtriG4DcSU0gip2Kwq59DhtQO2Kz4ULPrndy87TbhjXqDjI68Cp/j2MtsQIuqDsJ
HZakNVBcrTzMFW/JvhWQyYiMfJ6CDq4EPpQNqBrS+sQ1ZUHHIMp82Wk+j/mvV0DG
PJgUnmtutIktHMbigS/TFkMtcwWN+vEC6m9o7ofOEw0z3lhoQUSSNBoHwU4Nw+V9
w0ndXhZfcvPcejkIMDjxiL/Xs+KPWjQSx42EUrIWY7sOl9O5AMeqnZ7dCzXCKM/x
Kv4HARobA9n2C68VMetmt1OVUoTaH+ZbZ2OepVpHkiaaBPa2DBXrxLQlDmk8aR4P
83pCeqUgAhW4iBCBagZWtqnwsfrGzTXhoQUwK5u4RrdgaO007FIxrCudS1fuw1mn
4JpE4ddODXDtLSvk1eEkUUCSquplJFexp2zIkLtfjVnqOKCpFqH0dnglCm8Sdb/d
z11+C/WLJ5wQPKiYdmBK5HABu9szXNTJ5tPyiI9WerKBeJuBA4tgXcL6ij/YnDsM
ry7OCjWXzLPSfQDeoCuiCKCfVLQdlWDhg6SseKpW/DU3LC69IFWsrfdzCfSS3FIV
OjNMihl4NIGQcMNrJ+HCEmox2KxrIP4j433L8wAYUDZlI5ZeTnyiriEVfCPPxApv
uhdauicZgFV7KJ2uomh4b9zt7/HqT8K76wksmR8vdbhkqUHRPbBHBaUKYBmJTRdi
JlYRZ0aQNWY4okLvqry82colF4atTgwGsAw6OHgW/7kgIFj1Wc0o/KG3gZ8XB91+
OlunEgRSY+mnTHGYPRGADrGF5iLwxaaLR7iwWkck5O7dVORe61yCP36KoYAY3YYK
dOa+9kOGoAuNRoWo4RdUUKGSvV7M0/XGZ7bhWYb6C3TVMsuMonv2eD6qX1MHhdEp
8E13yP7z8GKOf+Vm7aIdynpyixx6yZT4bvHHdFiJBeIZkbPNjXf/+GoqN/nVoyBN
CZKmPLO3JFe1A0Tl7gCsnDY6G/MrLz7SxCMtG7sIBocBwcAkvcW6HStQ1x15IzzW
LekPIO4u6Tz8smTGRwUPHkFrHiZ5VFYzELVOx28/5Depsmut+pRoccXQIw+VCldZ
tCtzUA8ga/Ti4kwYSG+PJIbisQCed1yLLHYEvuBSXt3UnvYzl1fsS26pbGdJIOze
sy56nB+Bs1WahM5WLZkaa8CrCxG8XXKkgZ17VU4ND8j6Ae1ve5unobKfAM7ogrc5
NDivWF/K1ZMudze+V2lo91jmmWYjUTbHvSB36YLAgK5RIKCgANGMgH1o6msSy60r
7Qe3xXkL36DFEOCXtHNnUKEHpt12IIHI9vtJrrg4b6sxGzvpz3OngCUN5tgJErMj
f7b/ZDkovidAYhuSXZIprag8x0lfxoCxYX/3T/TtAK4qGjWBQTAHjb2flKDVTihJ
fGPb+xLSd8WRkLsEIrNLMgeWd/Euy6NP5DRzFueUFIijaCqQRHgXfiC0t1xbzbGI
nbbnvjuxYWp/AUDzV84KT5mgIaX9cP77crWzlUREi88+B1a/vTsTjgy6N/nc7pkM
p4TSiv9eeBkE2DdwVi943FxKfmVZAC8nJpPkGbH1CYff4tuScTFhCJ01bKyWYeV1
n85VGUuDgLAQWIGYZTP+3EXzrylUpuRPl2AtBbwgpBpgicc0zUwX2bIMJhcHVURQ
ddlOt6+DB4Q9gfLtfAHmHCfRB/2lEHbn0/vOEmE73ZCaBJXv9865BMlDo8NW2WsP
lfQeQZYt036WakTTS+WWFGQTy1cDYtt5RrCb9etd1epL1sVPXTdmiUIj53qKXV+O
RVQaCkg0esu1PgMjLAHZPihSAvFyhR5184hi3cOTWFWe1EloENvxcGBJX85mkpKC
TK/XZJU99sXyLDe5HwZ6SxrmN+phUwYr3wDdut6QxMPKkQSz5AC+Qz+vmlWNqUAu
6CybCnNMD/k4WLZvnxDzUf0THKoXdbSJESzpbmSOwVJ874Dp+posyhiTthsgOdyN
4oblOT+jxiP0a5zjVu0as5D/rNgb0UxDLsMkqLmYlrC6WAt+v8EVg0gEQMo8kqEM
xpnciK7/b9aS+UQhp0S7B/v4FAIDwaBG0lwL3RgNUp4dZ2lTmlT7ttdQWbEVhJ5J
QqSmTDBizLyVgXxZ2d2hijzxO/NIkIyxBMHkQgZKUuuNoCZbQi5U8dMC86UKVn8J
QuXZlhReyGD66JdENObOG0DUe4n7/mfXTjllrjluGu6efteEpa0xHKyYM7pjQyUg
9x4NiLG6ad0L1aUJIjl5cgmmAxBLh0L62CNKCiY2wNUJ4h2drbgQLcvp51S3r4pl
72ivH9Hj0WhB4IHJVWSimzj+Vv1uW48Ng2R6zXWXdU7XEXITlaIdeq4e7gGCg0bk
gUr4hQrI3aY3s2rypTrvdTgGDjbk+QK3kXOj19DffilgHaWiKUEJ6gIpoImkTcly
KLyhFcaIdXgKCEaOIp2uWIYgv/uTWDid/vdRNqk1hc9OB0Sk6W33DPN/VVxGYSD1
vkfzvvdTozH1AZ3cRWyJdsvo1K8RP2u8SdatTQu3iEle2QM5mI4MHK437EvkobPL
OWAgT1sXS8w8pzgSOUtLUGnotxEBEdwh6HHAGDnxpr0/Btn0WFk21IiZq/TO24JW
5++AcSA66ETJu1YLW7611wlOC8szmx2zQzL2vDZtgnUphxxdgi7sDoxZJ0LhjbVh
ExaLDVA0H6QCEeX9RFzpyQ+XmMw7KhcceLpOE3koJ/7rgmKtvhkwuC+ZurovZ2Bs
f/q9YvMQZGsNIVdRi3lyvLaeWBATZbRRkCcaCG2nzzyCpO1HNZpxi8mr9sJVbgcG
ERwfqsnn0a1dRdDiHLvh5j5W2Z5/euYqWaS4KEycAWVZ12S0xXF1QbvDAGYnezKI
QJ28HfrFjWUTvzPPHRiMfy/uvJLBMaYnCKNnQ1CHwyAwLuQ9vYThD/JUFjb2NfEf
33IBwK45rSr0OWsVHBY1o3hMK8YxmYbn1kRcjQmdo75K17T4xaIi+A1rp4laCsdY
N6AF1VNoFEyMMCXgM9KUeXHT1+G37z7K/rYerCkpO0cDZ2t+nixLQEFnB6vpTnMq
94aD6PX2CC/8Ds6Qfkj2L9fMntVvU8CA8zg+ecvIXJ8wOooxgV8GYhaUioncse3F
qh9MaoGLkSnkD9XIr0QYV49g1Nf5zDxNkbIXIQPum2yFtndcFiGD3IQuXz7+4QwG
HBZJdQgtki31lStTvIu+yMKVC69ifhgPCHEX8zCrgATukgBivFV2JB0ULOdoyLwr
7U+bZPMa1W5VqTZFkB4pFUFwnR0L1wsyLpDs5bwTcXuiLk5CVnySl11uClq+cpb0
cwPZfLVADv/JzRX9BK4M0lPWKpB9XBnZ6FoZGsyu4gtzqwJZFg2a7eN7F9mJDROJ
neRom0gVg43T837YpeqVqjOH1ExoCdkyqacPEmgGGgPBYzI2PMRrTwq+XJwhxQC4
1EyIzLnhaJJ/4QJpCiYuUJqXE2J4ezAFQdXGf8BkLvfXEeLDZRKjc2/zYiwRSkFZ
ZZsdmW+HazTZRyHcwWo3evaEamXRkrXKadYI+ZCGXb+Fcc5bNjLnLXQGaro+4UEp
RFaB1lK9xywSqgGP+Xtukr3aNYmhxFnVqRfpfdlxXsP6AbOkIrrR6XCBa4Vk9yIT
4I7KWd71e/NjU37VUoW0ULZBQStJNohXIKzTtC+zOlh5qzaIIo/i1wLWd/m49E0W
K36BCEP7Fs2P4oo+RSivkG+6BI5zVJErBphjT3qGQPPabblBy7rKFXKkQSXinMXn
NxI9yvk9Vye4jI2gRpz6dRtsMIc3FmAJPfMC6FMXZpDULxvwooQNxlCnC/SeDzXb
Mpb00TPQ6qk7HjTiWtD3EUmOKn7BupTWIfDbosXtkMbbuw2tKSSI9plc+2po4aw7
1RyfvSM/j2aqv5A2UaRkUxOhWK33v+8ySND6ObTM4GbvBW1uvGm4QT2BBBgPXnD+
pkoMB8w3NluNyYqNBFxgmta6JMER1nDMvSzcw+SYT1Mh3tlDHsL5fii7PWbf8W2D
o2FD1NLoYtzmgaBFUfGm1u7qHyhJ97SUypsg2kP5MtCd/nu/uPxrglwlKMI/l/4i
BX3eU/NWi7adiOOj+UWct5gJGeCmCRkNnXSK5YB1D/apfOxHKm1fff2JLZGOSEtT
V5c7MvplPtQOlA2xQmm1PgLUWZGdfYX2UG9Nf8ZbYW186RDLAJ+IQzjhOBOf/4qy
TqFPO93s65X7fMuOrv9Z1yyuGReOTNQ+gtPgZZiESNSIW4wnVbJx6WH4M15VQDhk
/i5GrUWN3Frw17cYsPTcCJGP7ql4dION8SDytsrCcUV0MMc2wDQWmD0D/f5Dxi0I
PRsVIKdtqBLgXeIuJQtQx1kzJtviFMUCG19d4OymeJoX1a7P6+GTOdbf2SzFsCBh
xYXdNERi0yk0GErKfD0tkvL1g0b5ZAOWZGq7PSYSL6jzO4Jj4Brsl/FwV8HUINnV
FSVhte22SUxy9mVaW8CYsgMAbBV/+LlK/kHIe8F0IdeEjYWo/vL7LtoHF+MdA3w8
07i9aIp/IAdywTe8IcIfRU1GjTi6PC0ZbcX68OL+nM4UTVj9kAxMVQRAlb727E3+
Y8uHW7Cj5TxrF2Kybknh4HNu/zYGgCVGk2YfwcCJXqVGAY4f2osBrRB+wMFAuFKm
hUfVkstFH30CZ407yYjNQyMfIpGW8cP5iDJK5KAJqIFs0A5CVv1O0UVBczKgCI5h
Hf/5b9TqNq4Y+fNaACkeA35Yqs4SDjzgHCPyPk6mXkhcF4THLX4XVxllBRzjfh9T
mbXWX/F7YKrQ2qAu8MuuEH0Wa6Qmz7wNcBmZBqJ2/FUh3oOEN9cwZonRsxZD9HSC
Uj4hoyVDHUCWHF2R/PW8LMp1yVteGQAOlIU6yDhU0UQq7G5KL83r9fLS+Jd7EUx5
SQMaWR3MERWG6sk0/qca1Qe6QBtkpH2/SI7SEtZToPFpEmgX3FeQGinpmuolXfhH
vWPqc+YFPSFOh+eH0mgRfr1QZlauXE0CO6ImalV/Wm99CzjuWauUuLTI3EIuCMxL
e/oLM0ybV1nYJLdQsNNY1HJ5vieeB5J61URzd/aftZcfG/GhslAuxJf8AxIrM03R
wIJDPEWRpiv/HFnIplf/ZlUoXxrHlr40U+f8HYlEBi/sz9vSZUAquZduZVpo0g4x
cnchLK46dUx25tUVBxqYExzPJE6vYgI18jr4zvd99M3bE64ncXdoGjwP2PbnZG74
0sHAnqVgJ8g0FeWDuFTCJ9EbxmabTUXtSRL+81WfyIo9O3RNmsUPT1pN452tnd5u
vpURApf36K3sp//nnb6CHZGJVZfkplKSPycluoY/+FfeItlON4z+d9rwwcjg+MdW
bMGpN/l7bIQzlNNTsQH40FZP7BMai/hqRagVI5L4pNMzdyOr+PzH3HGsYk+kOf7h
HLspttxCijQNbFil2dIPXdMFP9kfWX0BMk/9tfD2qcRhsHnHA34Ndg5iKfS0snhm
AFnu2HEMRZ94Jb/i3wDlExt1eiovQKGKuryvuf5Duyy3vLMVLhFBRsyKfCYEm9ts
pb2krcN9X7lLdYLdKe4GIyMoNe7MjLV4aTpUvIzOQDhbzl4jS2StzfLOuAP9tj3z
Y9HmrVtc+0g4SPz9U6TshRaoEk9cPb8PICNIwqJNIISfj8QCH6SRC/ZUyKvrilD1
FgitdVp+d3uHLgfQ3SZYe3JJbUArBOwpgvY+IY38rLwd0qqBLYwLqv0+wrZEWz1q
go0Mh+OoXNLFp2jxP5M6w3gWKqKQz5ED8mtBp0XFJ2Vj/JRe3xXjDdy/yO1kl4x7
OFUEU7NbtxWQb2uaKRumy0ywnyP8LQmb3JCR2Ci5RSwFzG3NIHt7w5StFSP9QyWH
2BbAcbOlZB/MK/KBBpUxZ/uMAmTYCQ6T4DxdayMWE8GUbjUljS1OJgIJJf5gNH6E
X3FZch+csd93U6qhT93EZYInEGMrmrp5eQuTlRAqdTzojvjZ49gA84i7tH9jvEjS
H6MO0yg2B+2x0aE9e2MnmOGd5mud492zm25w4pvZC7BCQ1nhFX4jMn5kY3WLz33x
VE/Q2fIZZ69l4nSUB6RejV/oNroSqxpWSdmqnntc2sV9DwR6kR6W5Uf6aQOqCUEe
GTjcbnfM2Mm5xWJd5mjAmYby/P61/UMX+X0B0clxF9mGe4MP7ByjbrDAwxGSvnpw
MWIeVJEfuKlJuxGZtZEKKE1cknTA6/NqbEHozworGLCe3O2xhlpXRQbvaTSgGvMu
gb6RawgofBS1MqZg3P3dRNXoPFV3xmTj32FwWtUmwC3sroUAZB2+XBYu1TLBn+zO
tGz1QSisBrKnPhJhFD5tm2m+rQ+f/6cP0cXlxNfDdMSOGPyxB6Lf+XqeIVhxU6Ez
e/ECZ5er0hmgUSWqjqzpNCIzMB+1Ksp5jDtm1nC9lrNPS2GBh+jusp+pwJUBoy8c
1NDym+xc68efDvwLQk7FMSuRq3YayZXQDPE7o3wG2Pvp8vW1tnWEST2CZsTCz0np
XJFFXhC2H+Idjet3S1q7hPA1JPJrpmH2UMTypKF16GyCNl/f6q29CnPlV/evxukE
2N4+EUaycRI6t3U2Vi6G4NyQPHqU+imJg9wcpfNa8j4vyuFksoG/1BnWcou08MPv
kWzs611FkkQv1uRLW3xM976qKtIHl2jPW1AugAGu9e1fhIElrN7HYtv59bWJyBYE
T+3R0fzscJ+bf8kxb7iVPHXEvlR9UpXT+KBWGJyVmXVJbJGbEA38WcAOC33WVOQb
9+nmygDzB2QnOsVKd5thAFHekabGIgRtDf/FWCamXYOJvcgdo1tMUTIBlAHu4lYe
r1P7iDSgYzcUYhUbDxIW6oRNWF53ABT7xdSb8gcO/AUmu987QRCsabvdF8TqyJg2
hwa+SfC2hAKZbZK3P0Puw78oxlxXlxePEgUBlEB1Xmct5Ed2FX8tNj3BaQUUJxp3
3uXSf+F57y/izG5Oxodsfas0J4WWGF9iCxjIX7BeSo1i0Arn7DXf5rol6I+6tzQl
oCp6P/Zdj/xY+B/0FojwmU7OLpVgwQ//2RLsjagRVox2mCeyt9fShBhWOVpV5lPO
nAV9Cy7pum6AvnLamMzNReLjVV9MJYGLd5WzFAjZ12aBe2EWpJuyNdvmra+Y5z+8
LNGAiHNP6hlNb0I+TX8gEXIdDYkDKuJEM8jB2XQBvWOtJtDi+pNEP+5DGnpyM1kk
AX24SYxuJrDiCMXEJsbP5fd7lFIz7qHeNa9FrSG0YZIwd4hGWMoLbwNGQaC0Yvie
B3sdxBJIGgb45DJVr6ufurrm4tsvkmN0komqhS6ZCg9Qbeg8xzcK371cfaaxyx05
TiKiBbX3wiQ4gpy5uMSUBOpT8gMFOSFz5M7MtsTmxxECDawoLAH5s87F+xYQ/BnL
rz0xyIj8D92x6C4H/ZSMHcuT7zM4qJSaUhQgS/xLuFXkS5h4qGgqTHjxmYx1fWcQ
6m+HkcyBfPiVx8LLY2uwLmqOS+iEzjPV55YWuAK7naKyrV8QXqGyzx0KjgsuKfua
zLYhUBstZNSd64+meD1rQD0iaD7Nc/PXGYnLIEk4jcxtzR0vZobP3xrRhOsr79Jb
LsfOMZAvTRUV3DlTjhaKUi3KHR9rrLhx81Nxw4PJGT15rPo0hZydK9iWcVJJjb5q
7oM2PprmQA5bMy1i4635t6PBV/qgFQtBRcL2ug3zhcWrZaZXK69nkJOfOzatSb3h
jBRB3s9xB61wDVnE5TrnP2Y5qpTYesi2WN2FXTAEPFzxbDZNpeHX/FLCeM/DfZAH
h8P5ef8R10S9ld3z6XsXInAwSIYR3j2tyXa5WVhlna+3mO5fcKcvYFjlaECh9rcS
b0qQf8CIIgWOdPQsMvrRaiqbQ3znrfHzE+AY9EUKpg0UK+Mw13PAEHOSYjwamYiq
NhJ8wyKd/JsYdRvAv2c6K+TL0OSMQngC+2I4N30CA4Y6N3DuIRHN4qOKvSmTGbfV
AHeIbEr+wnSTNEbYhQy30fMXkBp5WCaVG2iDEZeNIuWn0MkcE+tOFZR34LfEfd9Z
P8OZ97FAlwtRMzaNwEAF6w5qmPIoKyooI7Tg4EirhzowHYI80WZU62hLV1OJgwVO
RGDUwGzOvwvfMXnmtXyV2K6RmKs7ZOH4s3B/jwrfQH5QNfFu7YRx8KgiMi7rnq6F
R5V6kCV9lrklBNRPJjj2RUbJsjJSCQLfDpN6oCbjoHPwsbbT9F2w6LW9e9r/WsFB
FpAHL6vHsw0yDHeMSpljGS+kYwcUCgN3m821LRuV7ktRMtkANTlkAg4RNdG0K/FP
j8yYYEuzlZad71PJ6gUy+VU9r7rTGYSJeKjThfRD90oIUFrKyCtezmEYgc3Cn0/H
s7vMyTeTqJa4dBHzDLat0NA9CF1urLKhxiIndtB9fOkzGrf3+DclbMRkkAtzMMD7
bHi+avLsFxuLtnPJQz27FvSbz8yMZWBMT0p81gNVGepM1U7XrWRgZK2U5A52QJKX
i86LBxzMKnE7smb2temZBWWPwKyQSL3yQbYik1atAUSyQ6aAyxuSdTUymil1ulmN
YESeOSd04VK5QcssEzSEP1XrhPW6sHnqpu4nAdXZoDq/S7vSwZbgrg8T7Bj9R+86
jqwFYEcLBw2M9tpQ7hW87LIBamKlHIDuOMvTHrlN/cTowCSlnuM4qVv6lB2niBAy
0joEM4tw3j5guz20DkIMipnk+b7tqtMOWZhXoVmzviCZuawjdZIxX/qagCUdeVIZ
yc8fxTK9KnKF4yzwTEYih0qqR9UEpnM5TO4boAG91WQLR4QZ+MN1uGvZc9pGqoeF
SJjH6dWmeUE3lTCY0g4x0av2U4qEJuwrmgkU4WwmnaX+weeJQCUsyo47r8NMK8Tz
mALEfQyfQYmxEzOKxw9HrD+NgNCgYCd57D9c+0CVihqO3iJ88StjDHB0CDjVToGM
hiF83GP7/XxeIdvoa02okH33Wwj+95agJgTGnV+wfhV2NjbFLxhQrr15Z6UHgq5J
FT3Y6EQkcv6/heUB8jLKPXVysS327JURpJcNcmSmfvZqULUuAy9W0vb8wCu/kvS3
yOellbYhfIqjrU1sXc/D/k0HnzyxIk3jf6hi+iCdoM2wwR88UNk6Q5dUYVcs4VBJ
D/Lv2Dvsi8MB4J8NeGEem9R/9i8sf8LxXW9TEScGD5t0BVQbMy0fsEfMOwPcLaOO
j4YiHEecf/FqzDZ/8xhdsboQI2FsSohTaXuZ0ESJfrKHfasScltwL4G+ScYsEQdH
1px/e9pRjwPPSe5EeqpxdfvJlfLEFmu3yOuN9WWfesbXQeI7Okcn+mZk0oqxBtoH
6l6kBif0M6Q42sAxvzLSjUAFp9fVAR8P6gzq1GZecONiefFQKFetTXrQArKqlZ+O
/QPFn2zFrRURg3lx9NAKbxPxMo1lAVQhSsNWi/gYZDqfWT7b/jyoOCEocOErT9eV
yNOWowHMhH114PO7U+U37NHv3OJkPiFWoM7HlPHzJ3enrvhSMoAFqsAupiQO6g5N
XGeLNeoKSZBNR3K+d1jIgI5HIRx0JHaKUlojGDP6786ZYPoyuBRuduoY+9lG1hKO
Mh3DqeaV4YcHIPE1+sa2amOC1q2ngLugyAWR9K9dRfno1TxDDwgUT0DzZWlmcDiD
vs8jUreLBuTO0nTj2DYI9P1qibrurgRBS8XNURDbn5W3feACaVqDo2aZOf5ow4M+
b28sXDWNzjC9GaBF3qN1+TbD8zQIeHeBJNF81q9x3Dfif4eSQCQiS6AveHCP38Me
mcqKVkVvahS/KAXPzOwza5tm4ANLe6UO/CuJzpRVKnzj8id71Y5Uizu1oe1OBKJp
ak83eowWNeL9ADkVVN7rP5I0xUgtHDM85IX+bnkP+H2BmpGGtXIOXiaSpCwQHOMS
KvzN4U06LhfRXPCbLFqo16oZDyHetM5rLwFMrLTDlHsJi9FJD4Tyl3WVEe85tfbh
71+Z2mzSLMW1b9U1GmCrYWX/c95mswkDOk/VMP2iRi2mR+HETwgpBgmqJi2+3okB
LLQJlVm1GAEagtgKPvXvQDjCH4IfMT5xW6cS/q7Y6ezv9e7J8BBynR289VieLYgt
05lOQz1idFFD6bOakJkwVNlX56Rw7NC8uTBRWFD27WfFeotA/58cA3FFwMc3V11R
eLcAnxq8h8QedwqYnTYjN6lsZxoX6//je1krnrAobK/Qxt6iXrLZcdo4H+U+Upt8
j7AfGRYeCu13DRNamX+Iev9rLApUvkmeAl0RY8zffNBdVXNMMiPjy2ccLWV9ihsy
0RNZGTlgIAjOrWyCWAog8aW6fcS1UX5ORl5IvS4nA/OtJYySChvfJjj4bJktOTpr
7wBi9I0nmkPdg/j1J1ww2kBANyrQXoDVRGoZ+bsgA9UJxmNjPSS+YF5RfXIZ8rK0
yBNmLet3LM/6rYapD6NzuHilQ8utcb02+YRXyXWbd7FrLWRSyR3BIYk2glaFb6T/
quP5+1krehv4BnmSUcW/hHeTWqIMA2eZMX95SclEw8ehsddQY87OXEUw6VsA00j5
2sxADeKOgXhpE3vxdEUP2AnsRQGdXL/qRRgEPuF8VCww2E765rAjac1vUWtbBU5J
yLgm2Acyjfeeaq6HKSoMLFtwetqskd0PZvNOPx0mYOfpH0BMg2v5bF6sbIm6abmG
eSzhtx+vc3WDywxufaUt5WqvQrdvFtw67SCIIp5IsQQ2wgFdn9UhHvju0+Mig2PQ
wYasTtCLG7q4DVt2t6/Dhzl7X442bHY61YRTbCI5Ru0+CLY3sLy9p7Dbl9wTC2E1
DTlNNS3jGN+xa9VWvv8nRHQZh9DH3zEjLzLEYyDUZxwI/lM72l3UFP9wHXCC2NR6
giW51VXOkDmp0LCXnnqaTTgl8/TKKHe3RroMZf56Y8pED0IJiepDpOvq/AN4h0g1
hzH1DBauofsmP7oxTI6NH8ZGi2ErJ81/MR/CJh1jiv3uQld6XPV6i2cD0YDWz9Uy
EXuoT0laOswIeL6XB2SBQya489Z0R/ogMlMCbw4BuO22qrq5bHtYwylE5H054hqO
frPVLpTZETidyhWza6MnrsSBUmOFoRxAq0Xb3zJXLNxLLS27I2aMlO/UzPgben0X
HWJYSVCr+nuZ2toRYo8Mp6OoulUTH5wn6HdH7rACQ9+Dw9dko2VrFWnrRryhzfcp
rH8dAxaJRFh77+/96CQQf07R/U5bRGDq1vV+mKX4DJi3afUqFqUrbMOcfddaSqws
2jRV22r1qKhuHwbjPaq4aAdpWUCcrrtE0jISWUpaadW9Ikz5hzmoz+YFUkNj07Ap
w96hvyUudhaRlHt5VV/WQgZrjoV2HdVKlmepniiRcKqh7W2UVV+TNhHTXi8K2Vm+
4dDaOO2u1fE5vHojkKVKp3sTkOgnN9zYTP3C9wNSjwT/6oZjfQhUSVa3zxZtg29H
RZ/hneonl5bMtYvBcPn/SIi0p8XWxupZeJjhAXpEIot54Jea9LecEbgXO63ukY2i
TAMY9RyHOO9LvTWjWiium2+7nIgAWtd4BV2yc4jGEfu+lAxzPxW77C5mFJvpZ0eY
lcBK6MSryvHuOaOAUqqbgpusXBFievWYR+gQF5XV/VA4yDmbfwxxppcNObtEqxL7
sPDAuy8M0CIJ6ThbGBbbRmcd1AI6TH0R/ZbSthwYry4CNdNMMNZfW26gIAyZzubF
jPU6AEqPc4Pd0oPMym6P4BM0bLq3MWmUCQ/bmPf0G5ymt/9NGRlXAgRaVhx07KVW
qL4AF1FjeWkQHJDYxzjnQMfTALYuaB8PoZ3bp8VAJN7iWRf4EgRAvCsjL+3irk0a
k2KFD/0dNOotKStTnaNxw3C4F6Po9s5UnoLqPGKJBNFPHw6xox58pJvtZFWjol8h
lqAyla1IeuIQohPP70wbO6+b4YLnYuJ5XDcMyH5NQLFTE1PBkF30JtIlFov1eFE/
yeimE3WyfqMeLp4uAr90Ik3/OavPAfoWMxrjRYEeztmNXyZe3Emr0Pz69nRYntPl
eknFvJLeRVgWpFwPm7wFQuR01g5CdKuRAIx9TkTRk78AMTLLjPJmnEfOCEGUI79F
dtEHhStZIUbLWxSby/M29ILZIBbVbdCbjrvkhopUbBeNHIEuzP1WnR16l8iRoH6v
tRkxJc1t1UjT8LPrFtIYtQWZNi/YEynvJBnXj30IyChs4eqre0wCratcz8SV1WIe
OQnPD64kOYkSRxbXECARQzO5/ZdGnkL/tGm50YfVs8PIyeGxGzWEyD0VNjlUE139
bBHRWHNmgzw8LhZHFJWizGJM5seAoRx6Geoa0VDVC3YcBQJNTVhqfFgYAj+4pwQR
eV8KIB/jS2pXWKsX5BcJVTdKnZbwc3/ehla/1kjyLMPIyJTLD0t+iK32+woIcDmL
12fN4ZkRx15dkUTeEJTxXa5EQcjQ25r3WH1d69TWHHZ8krQfbyBEFQlrrhQcoxWR
ya66srb8R7C2Mp8yXmMuQDGyUEAxrAb6AEF6qY+UNnRxYESQG3iZfEYB1nmEp51N
TrqjlB5mqghjhFrvNYp9o9+R+9PcVA162MlkM8eZApOjT312tDvfGd+q2hShTB5k
PIgPd7ZfC4So4/USDtE4XrK0JdGG2URWYbBkJQiptX6+BMh2hNt19nexLQVsBVaV
yw7wwuRoBpf66MGWdx1GgDxAFpjhrhqVPy5UXd1Hpxp4ONoJIoMsAosxZniW3Kb9
hLj/2ush9IU3gZedLmrFp1Zy1c/LQhBqChTkSbmSP6RK3vmjP6mOncj1AFpv1qKp
G6HIfOg52flV+ItRxixYWwv9DPIfA85TV6vBHqlq7/enrsX6944TYJ9izNUhiUp3
ldUA5VKeJL+l6y3e0Y0PvbeMNtNqIHjlzvrjaeLL992aOsBAI0+dLszoZuUb26uX
x07HKnQ7U3nuSP1Mgwe/d2ZfuRtbRO+Kak4rO+pG8O1Zl/hqj5WMfQ+ZY9cMRk+N
I06vjiVEKORCYkIDrzngr2irW3vJsUqDclDEME1TDQ+jGqTUitW0mSvWxfkuF262
CBs05vaINnMkfR41YWP33gm/M3dYafWZHP/5PI9MUHlNR9RPTkGyFaBdhP4uU9uY
bPqY5tITVSn6wm5wed1xBFj0qI9KZyyeCqKnu2WgJ8g2l31WNwYdjhS0Dh+hHynH
wateKdLRcXLGcVeNYzYS9PyE7VeZNJvXD1AMIS3SpBlJnyeKEQvUuSEweW58Bouv
yFZ0ocNYkOxAjy1XtKE5XjtFYH/9qcV5V0NiU6W3IgkNuBhOOo3D4XIh3ruo7e9U
KYWfgfYfz7wroOI247yaa080Bm3A8UnbwJM8zHRvFYgFY1P9gjgP0NIqNQ3spVVb
H9wd/fCvkbOx9n8pouZB2MM5k6Ptb/Wlxp4OhZ2kFOKXMUIQQu7Vy63y9V/xRQ3f
6OKI7E8xWrgLjXnmaBbvLflcVZQJxnCvmdynDqGNNGpUZy17U9AJN5PabZKbRxU5
vH7Z8UeIxLVWWtchVepinobRAEzHR4+DZdaPWNNHLOpdP7jkZM0kAZuFNGzEoswc
iT7vYdJVM6JppHKBU8GqRPb4LZolQAWXzTpCLekJlgcZBKrmwWdKCxFanfKWopDa
tnMPOX+b9hNGgwFQ7OJ9xHDxC9A6l/XJStnsNq3EVY5AmTpMZNI9LiOUZbPkbABb
ZQfjPmmFGvSYth6NTkxgTxlgQOxI3XDC4Smho1gtIdN+TuzG6BesUxTD0A5kDflG
JmCxq01jfQqavgiDkjvwq3+e2OBVtLwK7ZI4HFO9kP18NCtrKYmHu9hgItHYlkYM
cz1X9CM5eMUsyz4z4JYXhn+7pZFjZ9EXTKp1zMstD8u9bq40B4BxPC08Wzg4cbbX
YihJ8PxU6i7f2Ll6nEuzwYzrYXyNsLbJuGtJkZ6KdQ4ZDIMyFDBaR7sjAXSpOlLo
n0qdIM8DUUMhHAMkSF290LHIoucMNjy8VSLnCxHxm5ghw8GWzg8katHWbNHcYHiC
pwrnEwF2VdqZoJOza+kIG/3DCcnbs+PxCdnoUyKqpTIBAcYuJYd6VQc2DHv16ohl
TlYET1BEUIN2yqUY/xx9L9cSt2y/ZQFa8hwvGLZQ9SQhwKA0FZZvlVnzsgXomhQx
7JTS09TOpQDCDUChbeC5lSI9rZU69g29sQLfpph4AwO2rjdb6hFnhqFskpCKiNLp
Q8bor2nS0/dBQNNRaDwMpR22wiGPcHuQCMO45OTrwkZkPb0f7q3uIt7FUN2BXOud
JyiZ7zy1eSbo7Vg6Ti0gKaQKXKbrW+1VmSuwkN/+8ZAX4+jk8A9UQgCa0lgkA9LO
Qh0Szih12aXA7LQyp/JDAmVnAmhwMlh4Jk+hmmgXltPbvkFEBSGFzjd4qUbuHtcO
XF4yTfGH0UMc0FjDPfIb/XLIn5+f1KGCCSqEidoYGALLDj9NVYGjS+JFUU6ZhZE8
C2czdJooJUnYwpo/UB4j70uGaIs+qkZzN+x8+EHSfE+7Uiqqiq/xK3IAPUQxXyzU
pd5aPaNTAhLOfFYSfbFWkZZJb2jp5iB9UB4Om4XYNrSh0wePV23UFBkk9eAhy8ta
syVkWqhPT9smk4Sok7kfujGzijn+V2n5qXi8LPw7f8D4Q+HsPZVsFQNCDpwPgSpz
90n1D4U9H2x0QyWD76KvGRDNhoQVBYDnTFY0qsPBKqqYjM28doxPpV3eRpE1AXnt
X3tzHMhyH+RnsPt4/V9egL2Bf3a3YMDYNvCavLB4fM+Ma6wPS8XYZ1g1/t9xHU0j
S7AUiZv6ZibB02v3tye1L4tGUe9WifN61XBBw1wG2h0oWDZjpBQJLIG36qcaFI3W
f31ab/xK+LeHj5/iOffblC7uP02jHNYY1U5/mwEwTgg2teeAhJx+beaz2qOFdr41
GzWsNa20kHuBZ5f0R/b/QMQmV3p/UAQiJdXvoUtrOOOSkkLlY6F/1WlX52e/P+fB
8uA2YQpsgaKwxRfNJoR7HmEEAzljw+mRT/lfNbKOkaOqz8m7TxoVle1AQfFJ6o+T
3qV8o9GenZ4Wt1YQbZySJSQ1si0zWA64vQht31Ebtp7F6vM4y7hJ6z8jJggdvVcM
ZE/jTwgXR1cTPm0CaLxvRHsfqCEVmtV21Z5Dgi3T/Cuq6eM9dnE+0VzFYdNwW/Kz
Z1OvEHRYIvNmGBMciIMiMRuo4qtqVZFhyW1P+Ij4TM/QXqsm5bx5euKnaQV9H/xt
8QQzdDgYJduc7/vFha2NNG1Eyw4VP7Mf9X58VY4LZGTWGncR0U4IinW8mGm8QujM
MPsW46kuQuag6PxdCzjcLcdvTiYqlKnLIunwHOzsOWCexyc4ZcOV2tmKR3LB+Tpv
qm3exmTVo8aUBjQ5CpFDz9tPuYAxPy5M5LoJNytMF9ZpPHkbj3F63fQl+R6vCa9S
XuQUAkTkZFTLLh3zOoHQ00PCtjjuaNtk+3Bu5OkB4FSIVFcDKExCN9tVCNTgbidf
DFXEmo5sGHXndod3MNvkhFbQLqjQc1UUxzpHFtl4CNKw1W8dq5W3Ly90eCQw3srA
EjWGZfsdMnYty9XFunNtjayd/gQStaVr1qtD1sVITj0XBj2es3DnfDKY4LQAz0/I
ISgryw4KuVEf0b5/dquDxCnReEOtSc61eFX7PvC+AnMItlV6C5hiUywY4vTGU/Cu
kEI/UtIRYajaB2SxaZO5/ICTigw8tZNuENNywL8ytcsDwzEH0+vy7dkZP+bp0h53
pR18z+LwiWRqeFB8b7NyQZ7jH4icP6xslP1wukvQqrYMXyA8Hah9G2art35Z0LP8
s8nfnd9u63ca6WzS8j10dAPD91o2cvo++J8oR2xx3CRSflA/6gl/0nYhwpF+c8C7
SpGY1oJMkteQXOzGZeHaCVQ8C7vttxed1xXidIxNY1D5ks3flYd0vpVLlB1itg34
1ZaKZ5FSjsTh6ibgI6lASvTCu9yGQ2cgfoy3waQQ76NReaUy9oESUfewUxyY6SMW
zjkFrJnbYw1877PTIYQl63naa3cz0oIPDvauhajP+hp1rXo1x8iNJiBYEXoD7wqD
2hkW2S65FO+O62VQ9JR/0EnU3gaIc3NBw20yOnjaxanoOqgyxIxNQMO3DbCZeK4F
g8MrZOCD8S2R0oUyt6T9FU4jwQpzB39xxJ7Zm4li1hnGFRO8DReDFec6b+M0OSLX
G4QFPfXPEINx07qCzJNAVW1QM9QRfSP4f+bPGJQ6kSwCjHSRx7gNKSAduhqeDkSr
31KpXrq38/8yhXBmlqX9HtOSEQlUjMb2ljG39kwdHTcyHEc1eSqLB4vqlUCkd9g2
z+4taFORd15D4fz+B2x6q9azpKn7j7JyL8Gx4BtAQO2SnVyuFeafxz+6cgl/hVZE
vEHtaRC+sVz5Y8zBUWYhpgJGywAWAkCObur/pp1MuCiJc3+Fe50neYk39fUmaHO5
AuivZpb0ntQA9nz7NLkr2Uj20Yb0XzKbPMr/KqNHpJdow3/4GWoLwUHFoqQsm73N
O3KCgMDTBCII2P7CjKGlnCgDUXFm3ltpXePqfSv7Meez1EMnSSbg2Q6FZQoxY9tl
n+4sthwDTEPJr6Q1TwsfQRU00X0W/UrppJ7LUdwZCbclK0Qn9fa4clZg3011jZZg
KcCjG1GgHGAi/F8ixOwfuglPQWDc4ANd9CW19Sp0tH2/CNakNBAGgmgamfBjrHVP
s0rav2djvhoTfamF74zTBmGxwu+Q8hXzN2BLCspSvwFsKbLkkw7JugYG/W7Yoki/
w/2n0u4oq105+qb7ENMaXEXovMUddd7VMUu6Tq9Q3nNWt44oI3VfesSBSuyz8ODp
wLmwCN54SFNaY7JcYWVNuebc9zs20ybBbauipp5FSXHKVgAgWzMwdLi3RHd/MXG1
FzJVOmd+XL4wab7OCMTLihmN4JGzJPWqr9JWib0LtuxY8myTKHyvIVYzNv0DACx6
kHYJ0YeZezJqblXCo3zxo3pkmkEC/yM8PYh3s40tsG05rdDU9slE2lLBvjC6fdXj
cZWwjJhcXhYY1Hp+KnzGAM7aZ2I2Sg9t1SxTjtLTibX2+dzGXLNQXbeOjLpH1bmp
fxEiDbABxlQMKatZjg69WsXqtZY5qE4Oroi31g4TDEMEOOeOvxrS1WMd6lUUl/wF
Y79NuB6q4gahwUhyKjHgZmXXY0CaS7C3RVtEfdJNfI3g9gBecZY6f0m9U3r2xnV8
ev5hTqcFPB4i0NJzsGPPvPVpH+BZOkTgvXXfaJYdumep6/s1jmhbFBojjb9c29zX
s1rjzSTEiEiK6vT1iE6oOu6Ubjp9K6qrYrGRpYo326jL/j7iTJEH9iOgawGHrrIR
x8fY6tr9WqI+Y+EMwWvU7CrCE8Tb08MrPhSIge5d9qy2c+26ZIi/aNoHVcoVDRk9
uqIT0qOhtVpXBbxj3tghIlOL+1x2sCDQwGV9lfpjqwmcpuJ/iqiwDAzetG1kxcYF
NHc2ESYjqE4+QeeYXFKgaf9heJP6b8DfFtQBSqgK/wL1Jwmciso5W9L0jt1LPvcD
b7mNec4c+MiTJwtj2x7sTwvBbod4td/DVaQ/55ogKFDbM4dNkO7TPRIGeyR8y19e
25W94aURRiQvv7vbS9KvWjOxZ1giQoe3MxlnM5M/a4EGJCJs2sws20hgf9hLMeoX
5HPwZzg8LLAS+Q09yQaxZNVZcYVCxqVC4GNZ/ja4yMkTxtWRUZxLi00a1/bpe28I
+TCIXn/PDFPznZYmm5mU5TXJA0mRpIYcDTCbwBzBIRlcJJU+kDfCvNRVnp0vpE7n
7qCfb6Xeo9GmvtLC98C6duZ5JTOXgRx4Qte9C2SbIf/EEbN+EU2r2SqXZLNdje+r
c35NPR9d/wNq10kexVq8VYwQlee5MgrPumcXgcR2xEcb0eskhHd+pQ11skGt7aku
FqizSs7tUoSc6TOxi4vzcn64v5gXCKRDpuz4J20NmQny4TPiV4gj6Vv+hmCZ5A9L
FPCh1mtr73AId252WFb+LGoZcx4fgRvLIhDjJQkNDL0JhlVtLvexqxtLWumRy1Nj
tqzVzPTz4HylnJLVlfLMuCnuXUmOx2KCNVqGQ+VXuhkt1aFEdklbA+AoiuQAQC14
Xl+bnkgDPMGqhvmsC7zM6sXw90himcG6YGoBPHc5PN9nNTEgB5xbLUg87g6Xzl9D
qZsIseh+KJ3Tl+LLkYnTwodIHtEymff0hwjh9f6mF0htlVE6KP5rvGcSSBNFKzvn
Z6FeEVA0xBW8zhiQP+pm+g1NuymrVAKYnQTGWqU4OD7ru2xobyKJuu6arrg1gErC
EKoEMVirTu/c4P0hozHOW+Hp1IIwIzdhuCj9UveM0oD8L8jwscjdIC9kpmYPvARV
gSZL2OGc6y2/wyfG2GvWRWwa/saxjKVUQ15S7xDwG/MN+/cbGB6m+HOAIvEPXcW1
N8T5GrzKDs4k64Zym8IZkanOmir2l1JI7OAwAX4jypmZ5USSqGqlNzqT2rP2iG6m
/0rys/vbYLbA8mHDyCLoytUEWIH1TqXKr6jeRh/tEUYqHqAFvLnXksbXPPENojkU
fxkjxBQEPItAY6j68PZ0bIpZ+v4Ct6l5JHx2GULr2dnF0NYWr7aXataMPRRrXQsU
e0omsZUmIRcafETRhA4OJpGPy0bMJgvvqvznH/mS3N3aYrbb+3pBTzBNGM22MSsQ
DXc0o6H0TtCr/gsnl9Cbgf+bBlaV+ykn69hAW7M8mHZ3w7jqBiChzTL7bXdf6E3y
17ZrebqohYLhsTWKkI2kg6yqONPb2XyVsvCr17d8RXwnL5s5EiSAepdIXkDTw2aj
7EGqw1DBvAhMD3cbP8FiGfnQ1mI9pXmhsMmTuQqjSzEhUK9ZCi2aTFfhoGDjBW1b
eSUA8zHiuBJuqalDWwfxTM/aIkH285t4QmIXfUf/P2Q3zIx7g8+XbLVgfqwsSkKz
KfSxSAeZXjuSUvXzEGcceXpjlNDVkYtK1jWDKS74z/Yr2prH64BKE31xiBPoKlyz
s3NFexnp3AqTLacEpNo37H+mvpummXRtyZple0MGLvNGUDCzWrmksqdU8kPYj2KP
/9E4BIxZHVRRGbxjR5p5Z+GkOFpFrrqZN5YNWL32WSpVcibT7ByCByQDbXWw1LrE
g8s12dnfmtxixLqxc84n33fgoQkcR7Zc7jChr4Cxi3dxN7OJW82V3QRSx45ZTDq2
6OnDih7uMF3eCFo3rzjnIVkioF4w1XP64t20NCfwr9M3O9Fsg+5UYWMPEqVE0Da2
kEdxCMxifzD0hoOGzlqaKyob/AaHYSs0+Waj0eZhk9aK+e7FsgAahfk2tNfJtzUw
PhFXY1CfcBzZ1rsbVL8oswLdRxSYKGH1FQNuDGlgS7KCuGUb1gARiuFbhddK1tEa
A1QGdlmjlmVHUVghw3zIsodr2C2GpxsmSVL7cLyyxbdPTt+DZ4r/AzgvIx9/XkUF
3nYV77C7CB3MgaNSzAifFgxp9CFBXKTnZU/Pl+7xjprBLMBDDU+OatimPHt9+QbX
dvdWXbUohOQtjNZrbpu48UySMptNKIpH0EepiC8Ctp0u4mTwjwIOmVLm7Esc56MW
H2IO/KMbyf0UYY9JKKvKGsQOmJCs+wZIHQp5pnwrpXlr/ib4yfkC5tkRH+qN94KS
JrhFFCHNSiTQsXHnE8F78F44h8Rrp4POZZOojytbzfp7GFkOxQVs8X7MpKcWWq/t
lxWuVvTciUolFvXBFDoYdMQhswHZLgw1xJA7mgLUQuBwBSRM8Lvh8s6AkJcCMYkR
Bb4/EVjkhkU8nOzNjewt+KwnM1JTyu1IIsJKsgRsrULrH9Y4DiKQrxKDBu5yqVT5
TViAKA1aeUChpoFiCPo86I74UWosZh0dMT0ZNkF5mOSsppYnKJXRmg14a412WOZd
f7IRqnG0AjH9cB+mLx2T3Gqx9ezRA4lb765w1x+DWygRpqrPY/iFZZnf+yh8iKsU
Zl7rPCW08vqUeyIpfv7Cpvz6SxTs52n3p7uJ3pId+SSDffw1TT/AiCdSUMPo9vPy
RqDTybIckRkKFjBzhOU/efUeCvRUAW1Vm7REnFM43IIoipKOU9a8HdVG5aqq170f
N7xxSSg+1KanCXBmfX4WtzXwjAOo6sBUp+U0EVlNZ0ltmCeiQCl/GVCO+wf3E23b
bdObOSQu3yP77Q57KL3317yZtWrZYQ0cEO5a5VOTdizIJ9GyyVQznHiU0kBFrXlY
LaZmurYrphTyNMNnsU6yRnUOq3yaleXkOYzRuy6MsU2+aYWwKxmbEQAE1Y1LykZo
fEstrtSpygVoRZbRM93XCVqCwzPR2aDE7Dkpe8jleNWY0sqYNReIAC1FNTsbH7fd
f7QRyICgWUOdoCwihXM+ya0cKRv3T2Xp0FnmiPW7d/sCG0l4oQhiu9BOoL0cRVEc
D/4vKalp6qhrzhWGEqhKDAKpLPdsyExaQ8tD6bKqPiyhzJb/K+98+SMG3XtVRQO2
ry5RQuDFy2m4yfoghLO+uFM2b272qXJtx/qmKYcRzym5MxoStUunjwOU9Q3kP7nP
qkAy+xv8m3JC0L+Ew1mIjpU2hYUcgbUNCo6NOrdYO5nc8d3/cWfczE5pujO/YF3O
GXlQvuOgcw5a30UIpJzZ11dCAcnE5AUgQ9BD5EfLrwWLt27itmexM482zsN2qRkP
y5/0RCVpFfn7iVYi9unh1q/hLc3Otgw0tvehXm6srSa43gWVq2ll0GMbOAl2Sml4
qJCjheZuuy5wC4wkcZY5VK2sUlYy/TcdOQRqXAaE82rNndLQrbBMwSiMS98xLzto
Gu3S1468mLWFEMk6YiArYPnSMFkZQb3pB2015tt9h6LQCK/xmpsVonDAdDu/LP+P
70bYNIu0Ta3VIw4CP0zJwnaTe22URykgUCYlmHwfliBYC470fhYPmbdaQq/Fs+cb
cUMugglMCIiBWnd3qwI102csftbPR2866bKfsnZKdTQlwhIf7fwzZIG3NJRB+qJQ
e0kIAVpwG+OpHxHAR7hTX50HolKwrmPA97vKuMQ49NihLR3eKp+i+reADh0utVvL
rcFGDUSVWm+mttYuB1bLh+ZtjBGSCRn53ZjjpvjuwzBTPc/mG9+v7pdgJWrm3pYG
dV+4sUIMMIw7mCO5d1MtCMiil4lGA1da3pT+XXXaUa+f5wmLDKcMnCP7O+KFRaXb
wbCj6EUh5esFDXwZ7+fT1k09B2bm5bGwQn9uPyfSKp1Sh6EoDCWAXb+4g8Syc4tX
Y4YmGRZqjPp4KbT3Zw/hgbKJIqZ/KUpCVVPlwBmuRE81kH8WsyTDjtaj4lsK10qv
q7MMENW/IwZotujtlnun+qrmby6c316pCiu6udwSjSmSdM6pdZ4jTJAdGEQsSt/R
+G9oY1nMKMW+KhP8/+RSKth32uQLKD+qV3V8kT1ESRAsVhEetXIMTa0VOQkltEU4
NzH9kDfNHJMhDPbKAzqWmnVtHv20+KXNLMWa2nuRJ3yQP113zbCEqX9RSJrDM2MV
QmpTqFHXe6a0UmBZN3sZD9cdq8rF/UkLgmy/CUalqyaYOIjzXk/Kru+1SR4gxcTL
1XJWWzCAOQoKoNAZXFBRUkQPMV1+zHrI6nBuUucaijvGMVX0PY8VKfVBmFZrcnZ1
zNQW4dfXb1DcDaaOljZWL4XRj1/KdIVtNZ9w/BBQq8s/cRSnDyioTkU4qL3FqEw3
9StFAXzeNRggssRynQuD41AI3md73nED8wIrDp+oYDMKmIHq2vpw4aTDaF+i6MCt
AgFZPEC54mno3kakchwB7Kth53w6vf9AVhkmOwhC5c5RTcGuVE8oekum9TxloRNR
IVMjw1wPIzUTnHbWlrwb0LXagTW/CibR4jLXgVpk97PvQqCpl/qIKehOnLARuE/o
NFdg31vbDTJnlXoeUipw2VEb1H4BZUI0Olbx8KWsOxCxkL/x7kS3U9OJgDTNsPDn
eQzETg5BfUWRT/z/ZXzIMSXabkqnU3G5PiEDd9RuwhV0TNGpseN4gSvJ0oLFfljU
mZoUNskDjpNnpUjqQURukRdHEvWQpq7o2W9xyem15cCOUCZE0ZqQK6iK6Gt+ONAw
QOQ0JHU+QISDxhzR/j9zNmrnPSWDhg2VXZYhTejAMmk6MZnWpmvT0wZQ8ueM5e7O
RIJKKe+7YvuNSG1iTn6nbuAVkYRPYnrqzbR4smaDzhUxPINq0/3cswkiU5b2JQ2t
meMEYRtVmz+LrWf7geVZFnnAjLhvqNEqcLD/2zwv2NZAD9tcfGd4Nm1EyCgEeSSE
KdMqxkO50ZRYNgRgtTMX7S49SmDd+pzqYGhPWzUIFxXvRKNrKr2poOm0vwBRq5Ww
wXMY/XDQWGeC00SD5iqF2K5T7P2u5FDoee7DTr+ecRKYqB2jy5uQof1whz6grltQ
uN7Lqirhs2VCHErdPYbVn1Tu6H36jqb9+09A+e+briZYAO6qvSqES9eY10/tSZ1n
2Mel8OcQg+MYkjq0uC014xcS9CSnOfo+KrTeeZBt2mw6xMVDl8ja4CPnKB4ZmVv7
C9j/Tk7cign+QnUFZYEb4UBYcS0jTHx5GbEK1Yt3PAivUEOvg7t5wMT2vkjfDWJq
nyoY+WbgaqW7/eoqEagraVm139H1ox4WF3FmDX5UWn0Jndvrh2DLd8/I3LAbKRMi
X4HMc2MR7HoJqSyZmR6Lfnz+cECEN6DYjWkR6JS6caqCJMW6R8orUSfMpVfpPGbr
WmJr4d7FW8nIt3qI+3yGrNliY/TyYWYjHJnJfSKC1gg+sjWUO3048punBadWahKK
mj2qJDqQnu79Tp07IvG0RZ3bcpRgt9Qgr0Q7FASz4Cc7zB6qEyzJldV8ixPNAC2z
kAj7L6wnIrXLPn+NmM9edHuQnyopf9dra2pXChHv5N2GyW436+8cGSLcK2uOfLS1
gyEhLzlSEgprFDfpl8nD7c53cYwb+b/6IirSvSPxk0mVdLvfLvMErdcZAcDzCKQz
yXrJCHTej7u+seuOVji+4yjkJqzBjrFBEtWm0sYv8KH4oGLDPyUAq4xF4yjuLgDq
VfTMoZGDRo5aQwHS5bVEmTZk0LPQRcb/j86EQuim3oJcZxW9U3dOm5sGO6w9Dtc2
cpQjirVWvMSHvg57bGRARrnrB159Crx5ZCyC/g3qEtNh74mZNGCRiuaxJxcpsJBd
iFnnTz2NY3gMJhV5NiH00lAF+zY6qbDj4tUsdq9z2Szq8xCtruDE+5XDWVtMgj4G
s+p3j5eWiLXUk3u2QHco2KfUr/IyEjM0RZrsKwjCW/iRlwtOh4BX/S2ELKJrLWur
VNwbq9Dkp1TUwXAK29jTRuL6WPw6w9i+lUXy4xGrDbho8z8KOOCNwBznAojSz6vH
TwCX77BMq/gXyN8KaiDhUaf37OyzMDBzsYldhRZlMwe6HxeF2pEdv6kmN9PtRcE0
kNnvAF1vyobqXIgco1aiNS0YhtpckUgDuVQoTdv4u76CuQWNvPHSd7Xvwd2tUCPs
zostxWVJvn9H0+FIw2z1pRmFGTWU9SEOqiuZ+YzRdKedhPVdP76rJX/q9evXswM9
Lx0INfetjd2rkM+GdC98zmThu286ZBGfUoJkeMpwjymAsqBzquQwfZd6kj70mSyg
a6QUBzpIqnWnZh9XURbzHDLn6ZgeShExOOVq8psSPsWMsZ+WSZTH0Ksv6LbXKcPr
X5suUEicVGw8kcKT48KxyQTtvGpwbD8ctbWxRUMhJN5YhpNnT2Ilb9ZYWc2DZHST
BGeOiW1s3RkNMr38PZbVP10RaWGxDhdwy5JldZwYjTYJ41UnFozgGpl06eRrfB2h
Fto5fQuClCa2JhQmneAStzB3Ly+CmplWyjNfSIg8uQ2ZOMzEsHrC8w4HaQU/qjvs
0QLPOtQfGjsK3Y4665x9Zz882KnHwXm4/KBGGYlOnKqApfyB7CTJG+V0IoHL/hrY
xBmUOHwI0PdWB6K54KrE/ovTpiVQ2KHK95LeZ4qvYloZ6hTx0XxhoHyTw8T69D6H
Le4ztWAOYrIxf/70KoY3344zTjEQfh2ttOT6I083RPlApNedl7n4MtRE/MYScxOj
xrAGY5FGrVfCDGLRFKwPFp9KyHHF+HyY7AhNbOA9OIyLcayXTuJR5VGJVr8DxER4
bbwa8zzO6ZLYDnN2FB8B2U4QIpWRcFe5vz8VwdZ2IZvDgeIZme60jbp63L6jL7OB
82JXM9qQeVPaRWlPXEGYgGHY4ii2JuI68FdxSQJCh1TTcI6OUYPoPyjoRd+nEQe+
VwyPlgw9s5VQ21a3GbWGQN+xoqRvLpxv2lcwURdj7I7b1+nlnHAeYqu4KWaHOOcE
fBqpOQyNytSHBB8+MeV4MGfn2MAcPk56vDp2x36VFV62y1PlH2o6xdpmuiYuHf5a
8YpwsNueD9+8Fb2xcEIjddrQ2t6Px7PvyyyTNa/A8mDqHPr4uU+8PDn/nR0Yg35Y
CfOsln4H7NSPY+Prk824cTCUUIqNCqSGwf/eI1gjsWcMAAoedQRzmyI7LltFp+s8
wG33/FESjZjKzCWT6OfMc9Tav51WLaaWY064JPcYOHgYTRjwFAKLPR/KlnOfL7pt
wpOgACj1Qv4AvqL36d0wrNtQ6gri9pi564gB14YOlUQaI4DtWnQQ2U2G9E8+2sUZ
oAGpK4G5GrgtJiFViW+sZ4nog+SLd3AdljRdW/bbUIas9WMNOZ7p4R/6nOdSA/Bd
K9ueOysLFqLpYjsvC3gOKKWmwQ2EuuA2C6R+MI5JXIyfRx/eDJZpdi/oCmuepfJQ
TBDe3xyf3KHQrVUJdphpdGJR+Uxm01/Qgub23GyFNZ5HEEbE9MhJEsmzLX/shVB1
T7+aNQDDooDQMSxZaQ9MnGWg0NkiU6x7MZPY+uxiL3XMSfdIZxf3E7ityXXIA/uE
bHce8PsyrtDssG/O+LRjX+Xjl2cytPxm2amCjAaYAcjcOAN7+Phi3ReW61lEJAvA
KZ7byjwpG0sZTj4uuxQ92lR552LPIDL8eKOt2a47go8aq3swxGn5x/pYZBz8tkoL
RCY8U+8pZFCOFwirAVcv/RVpM8SAKsZ8pgv73dMCXGxePpuGSTyfbggV2r5OJQ3B
9mu/DpqO6zySncDO5kHryUIB4scSQSzGoT6+8EqqzrGAfs0ncBMIf2Bt/q30fSvE
FEmCf0SrHCrHIrZNgRaToxz2FjzKvjh6wSpNjiPpp17lbKFnGJ7NvPLS4RCigKZj
XRE/7BlkV01JIgKfTDupRMO4YAfiGxzMNM7ow3duDRmUx8gXi+esPOGVKO/9F65u
0CgynrS8+9l60AuSbQBwg/GyNvqlCwD7B7ezTQzK6bzftEKLWACvNkjZjTGxrWgj
G1xlo25B6pSwZ0UZd2btZfjhhHCqlT0/k/nVytJgWF0s+uarDE7CqBJ2vZbyLSQ4
wJB4UwAZCHq8JKoMFwhkAf35Ew+E04tSUcrf51BzU45LcHvWRDhVRoaVRH8WpBOi
Ls88yopkxRKPgpj52WY+yCbBEcLQuDJwVmn4p7UMNMXaxbdLRzd4lUlpd2AKOLHN
hgNTk9bvjVpydak9sb6McggJvN/9uzNuLP5iUOxAf0DMQDZGRG2dWkWSIRhOWBA+
WDBnW6A+YatSdrji7fNxEsD8DFmfHyqAIgcnv04HGVo04YeIoCKAeZw/GvNDLVo8
wRrUycbNMUOyVXy/VC216U27j0iO/aAQx34nbtc8gGzBLkFpdD52Sq5GhNu/dYTv
x0E6mVMiUeW+2Q0/TEPUy5jKMYDIlHeysInOdFh3VRPHDffgQKhbqgKuuWHVpDTX
wgHYJJhWSN/5utbLSWzCW1FK+NR7hnywdw3SQrQK4VyZ8J9gLsNgZYfR2e4I2BwQ
SBPgbUlcEZ/ju6F0nNCtiZo/dN5RMyk3S9RKrNmX+bB7sZaFgCAIKr4jy+pEq+s0
Tw1cXAvt8OjHqjl4PrrKGf46bio26IUWjVs5rfRK6w37tanjdNnT5CU7zjAKBYnF
/pSAO5DlmPNz53RDwdkud3cdj9IGB34jSDXaB0nXzQO5dSLBlf+j0eqNuwXuHKOU
y+9MYFYfJMKImcl9cKrk/h8dI+2NCxcO0SnDVKtNyvzcXUBd9lPeFmOQKZkiVSvZ
JR23VTv9+3GC9Fqo8Y9l/wLHYq6im0MHTN7nMn4kA0e4VoTBl76K6KFXcdaW7FR9
b3hxXCfD/cuHzrvwsUrA+sybd/Nh/gOcRywvKqGsjVeLm4RtSgd80cZGpnL9xvAZ
yWBxa9eJ0ICvSiik9nW/7IkDAVXfAETQd7jzOz9mQtn6XWERmqkSwOy4cxRclCPh
3z5wcP8voJT7jOQwLXNi3rweZ81mnuNL7Sz9Nnow8EoV456xD5G+NVZs08PaH1hd
S9Teq7/adfvilk6DCxszWKk8yjXF/GFRMnwnvQpUvqEunPrEp4dbY2Ks2ZddOsAI
zMVwVPrChXXpLTblcuCrds0tAUNEQZJWpsXA0FYswGWl/8S53w6IGwP91n3NTj8R
CGPTchAc3VcGwfQfn6ctdGGErY+9HBoq4K3sSuQwreY0wMSpHsShoCWw/FS1krT6
57uivZc3PPAgy6jMbxs8XSyN/RCYztifGvEWUR5zTa65EqpBjO5ykBIW/Tr4rvYZ
7od/H04pMxteFiqrer74j2sBNPPHS08Xbrr0C+gTvIYvB2LRSvx+kQFZEBpZrl+Q
qNebLzZxcw1uxagx0rJ3YVfsm3Hao7FYxPO7hGz2mclv0esLSktEk0PE1tlhZzxK
dE55rEzRjfFnO/oZk5XyJMkb/V9LIGwjaeWeoXlwXtsGOkVzDsSq+DNN/9x989bY
uEGTX50K53LV+AXr3o/Hq6f/UdrKgqZC6iucD6WN9Qp2YAB/cux6CryOjO7fcKcu
dy6qmbpx4/ZhplvQM4W3CCb0nQfaFBkJp6fDPNmrr7efSJWUSFrgdDXHpxVco5FB
YFA5ZQcdxUevsXsWKzzyUNOdJsTW1uTjyfwva8V+SYqlQUfTh0FJOzxWNb+xKR8t
bq905VHbV2F4xFb5biV13XLDRTfPuviLFBgvKtg/b/aPdTVzSZZowJE/74ipZNXF
LkxXusKB2gaI7VlqmsdHfEQeUh6UyO8FL6JddF79SnP/1BJlQjiXMqo1f1kshEPF
+9dWx1kAw9+1etssIPwgLxYqhmCFqK9AT8q8D7kn+Xa3dtmm6O/rjCcmULmqv5u8
qAtk7X3pSDYa9v0MiueZZbss8PamMib1eMqc4BolLwiXoW2/Ypz7DXl+GT5uL1mA
huhEQCJc/22KhNgFQ+i+W7brBehfdWOohFwo1ECGGPpdgO92d2CPSfsawMUVri3K
JBsvaCsFvfjKJxyPuUl5AdDew4cu07YYuyJxZdIFIV2oVkxWnSsHBBKw9B5bw0Rv
yzMT6VdpuGWEEuQ/ImyVLe6dO4uGUprjBF6clXM+ve07bQTsboudmiSuo7eVVSks
nOcaYXJcjTVFqFi42thbw9Kvj6S+2+F8qKLgUarG09Q96VXZTdQIutacxaMJHnEW
sXOFJI1ig6SZLKPyakTok9waU1qct6o//H/Tbsti3N/pnGfsdf1cJdzEpZJdzU8k
7nemXS+I8PJ4aO1KhOh/8wv31SfU2LI+TJyTqgrZhcDlB1JhL+deKfQuEmbO3Gae
7mAdfr2t8+j1wTpeQIpg3jxh/aswSrXqntPqcBy8zx/lulvnlI5F4+CSUBbLDjNu
MwZdk3v8LqJ8NFITUPagVjdzTMugVNIGlPp8OzQ+PA7CApNyCaxY50GFuakQdM+d
eOUi/P+3+o+h3Nnbha2UbrFZLoa7wBFqZOBzjuLZG78RVB0tTLBaxbc1XfJ17wRD
0Y6EFAr6MHNv8WXj6Lmv3stUQ3D9nDUrwO7RZk/NuIaJjRuY0Z0xEz5yGtKX/kS7
Q2Xs1nqXkpszZAU5ee5f3h6a3W2TLWcA1yx1VI1WURE94IVYb+BU37Q+xrIkL1v0
UZmGhJK1QwuAHLwUZ5MprBVZYghgmY9upxsGxNP6qqSAGX9shmBiYnrp8cyHNgzA
vYZ2ca+dKp/xJZZFLDDKMdBB1eUtiRaUpG/ziSnZ/hS8GOIPRwICwXjWItL0V/F3
1g1t73VUcVYcdh6L4aZOXCHB+giXfE2DGcgV3A7GsY6wLLHSOSZYeacyRm+97H5/
hfdQZGvt5EGYbpFYXBmsejhHO+OJYExgPVA446tl97e9SQMnMiVXIw63WAq+hb00
pheU7uQNK7T9bhSRJdltcRm8geQvN0KtVF+Wvf8d+1/fMGCod4UZV+vHrjOhULP4
gJvrBwxBJ6zWtOCRD70fo9COe1XncRyCRnen3e0NCTf+9HTXosSO+zEeKnvUfRfg
Hr5SB4stVT/ZGagBSgb1+3oZvClzA1O2iojTDLIkq8S2EFaZcNZqCo6H1qI8hH/m
T3/m3se61LqRUKlD1FUr7PCMKH9F9f4k5Fl9pjWuuWqraUIwCNSo8+CbJZwe6D3x
9G6oS12WRJc8+JQGECVdxhCM+HR+hKCjFrFkk/XKRMCFbUjJB6aOLjmJU8yeiH2j
Ergi5uDmFFGPhF1wvKZvlttS9KshYMiT6o0qgIq932MVqfIMn54/YQgY3jjD230l
RX2IY8iYypFtb6vchTape7c6n7sxOtiLfIV6zFrBhmr/ehu48gp9tsVF/QvNlKAf
1Ta2l+36A3kzcjZfqysidV0OXuHhMzYNdUSZRSvEpk6NT7LCd2b/zxokhrKXtZ+M
q6Tj02Nx52/lU5CLwAySEaKntaH6wWNcDZDaz+hZAknL891kpWlddVl+bM/6O3p3
LTFlH9ecgKTrLjrmtVHrvKNcF3C4jHTsF36PMgA+GyLAzKXHFQmuhZuhrZ29KcdN
t6AsfOM1dqVp0j28GGqjlzKZ/yha+1QJ32j0AuUTev/+OcnmBrUCeV/ldeJfyfRa
fms6FfaERsmF2Wzk6QKgoPw/ypvAZQ5wpa8TrkrHwgJximQIhxb2t3qPlRcOCytJ
m9EIYSZ9/8+yhJpHS1Axv1h2ABfMrqJuyma64uOZz974P8MG+/mSDgMT+BAow7Cd
x68Z01jtt2Ri2JMQt8LLwFYYQAvVZV5BNvJmVqkgPd3LACSwjNSkH/GGxD8eNiYO
ngTRKxr5ciOg+FMAZVkbONtpVPFOg0kwljMN4XJP1XUNSHXHfuEGZXI9nJlMy/RU
XFflzm8SayXk+1vt8VKQj66dOPswGxdhW//jOR6oNtF4ApxV8HXu28ykZIZPYwVR
VajKPmhLVjJeu/da8lu5mxQqYSgyw4vs8KtIkpspYTboNkmzyor4iIXmVsg1Fzw6
ktZeXfW6Iy9pW7vArfxDTJNUJPt+XHAru2TVPlVGT2dldUVG3jEpp1Cg11J6mNIr
hQf9gw554+3CE7wfZay52bhE7/gaCYnnsQhMJaNS6mUl7USfmHYOrP8sgCSv9YC4
Q7EscOi37958ttK1o7TQt29xqdUZ8gkh1gLzzM+r1As+mWLT68lb7era2lf1t8J7
ezCoNc3bJfYaNrvUbrOaVCTfIKps6OywM6faEmzvjnlPItTW4iLeDwJHwwCiBCuV
5dNytNKYxWJlIW891G07XS6U2Ab8O+7jSl1zcBQtyn/qdsIcbgFs44it/YAPjw9w
A3BYOTOLJJSS5KTLy4St/JqUc3AaqVMKMeuGEz1f+Gr2pumr+qZf1NdE+WMFjKhv
mhEP06aljq6Vlk3hmmHPMArQD+Xopafc9aV1k1Xq3foyMK3HexTs4LJUm+K3W4GQ
vk7qkpYpRpNaVZg6jm6svXewd4nr3qDgQdHtVRnf6WoBNg2U4K2m+km5SUt+nlCd
CM9/afPtU07ZMsfbHWr8NlULWJkUVVranSnuGTN9HiSq6jokM5jx2Ov4jsNyDuxN
g4AtJzV395gh5rEckFG5s88hBeTNt4ya47UqfDT/BTLd15ic38KponCVwyvhk2S2
yCjsUgCkbRkSwIldAfaDcHtbiuzbO7c4Qh4XBqMs9ETOtGBSukswSYNNnt8HwOId
47zEAFnC3DMHePW1c0up52cjCeDoGa+dgbi96oylXXkUi/C2kbCgl/A3yGTHJchx
9xRpNLUd/nXTcKLkd54xLokkTapMr88GmbWaJyb+5GzZ0jptC5vmOl6WEfe0c9wi
taPULClUXeAgDHa5kNCbT/+foXB927PFOOhrr1XEXeAu6A2UqXywDrQ7PIZqgxbO
StsCysr0bqHXXUTydUUHqZaJlRoioKBluVXiKYLPw7ut21/3gSxtF6Je2b+Ov3/6
t84tjO37kpJKX6X2bOimocRlGtEPRT5kNtt9eMyG1C9rn0UKspl9KxUz+sdutDCS
1a42JZomkQql6fgZbyQ8pxwhnDoQ9OYxP/NjrpJ58vbqLYaT1CruPuEtilOVUMh0
wnqc6LQ9As49ln7OCI2A+SjBGv5P2FH2YXMyVLJomdwLkkML6cA25XL7HFrKX/sK
AHdtiih3VRh7wzE4cO65RYA6GqVgaXFzLGkPOFHpFT2uPiiLJmVUVcParhy+Uv7V
KYVsuQlQxyJGnlhivVLze5ialG4Ia3VUzWI7tKsR3JeisNtwNum89yPU0lOMIlJW
guy1r7OKNQJ7xNnDHIzY3yDQPvGNdWfWuzFqDD9S1ftyNK4W2P/fym/8Dm/Sc592
CzUOhLZma9d7YILLqpbII2ad+CAiGFHHiGau+7VFZlogSmHZ8nTAlVeWV0Wq7BTT
27h47Xl4Uzux69Z+fOIuo7u26EYR4HfoOBRyvzZfaqAwZ9wmRuHVITIhfUfiRVQL
B1iE5yjVFONIyKLFvI2TrB0veRF99OLPzFn2b8/Edx0YLOn6zIZn/3UN3ULUvusx
1Qpmq1L4Hag8BxcFbVt3yESzOdp6SHV6yI0+/GGbEpDVaM9iIRVO5vGRQb3k5sIO
Kub428HzCX1M+fDYOKFerEsZ5VbRGMw198nFZYYezpHJZcchmstUNVJAiAQIKdmE
m13TI2tFULvm3s+7CY+g9kQscqrXKkigMEHMia8rctz8U77zcb3+OfuQ46LHv3iP
YEdmPGp4DV1cdcOyWDVhVCMNkVUAF5VgqTgkaRuwgkA0UqvBicLCMKF9Sqh3hXmP
1Rg+uR2MZcmQcS9cHgBfD/xdYiQPNVQm/nCLu9yQu7Qsn1H40Eo33vTS5Lr4hsvk
GbPSrAaYPBV3RokOnY/2P5I+i0ONYmuJKz1HfCr9xJc8mv7uUu6/ZptYYBN/pMgi
YPMFnykhCZkWo9bEVqiUlC9qcdk40mFnxXvYF301JJeviRZvbL/a6mwQ0lbYNtEp
VS+Zq6sW8EJEQQfBXuSK7VkmVbnqO8P8b7ghLYBzIRTrdCqePK4fQfNICfd1iKi5
p3YLXndmHi8+lCJW5wcd73IKnuneL+OZ4mvMIudiUcjuoekcpPFOIvhFGJlMzg6a
art/L7Rd+x3JB9bIfSQeyHz6h6ayITvdgk9r+mq+4mTWP5zHejVcziQ6A6T7E6er
EPqk+CXHG4l9igaw0DFoUZ7IhSffv8yMdg6iER5W+LoN1oZnvDhUsAxa1Ye0XyL3
S/WJ9Rq4RPnfNqgfWm4Xp30E3UonZNgyPneMBd9oshmQkJYxgEjQVjuEWqTu0ElI
guzzGMWnHTzbu1MszMvDcOwNi9KoBjY6Gvpk/8PXwgtBM51qCjJZGuxD5SP2AH/p
PDsmn9hIP1n6+ZMqydWP5F3dFDo0gwLWXE+dfoFJZPPgWktyQgxPHlOlXLXyXPDc
cbI3SHySecGTZToM0+ODmyre4VB2ZkcCaf/tHUxWQEVG88w6GTWSzwIHxeytkevX
cdm0XbNC4ZbL3R7E6QcRqnzFkOh0b30KtpdX9YebHba5GQN0Jx6IVUqmL4/3GyEr
LsmNcr3tfqHaYGzh4y2QGNz7+aAxnSmsP68AW4mqirlaWqFkBK5RiWYqLLSuoned
BudmAuQhbCuCCYA4khub6zvrJ3zkTcjRLB9m5ugPaiT8/OF74gjyL/RHb+xxG/SP
/YrGw0F8Ajdoi0/fDA+/pI2Ml184xcoFOFl9S98TFOq0q0DMmvCKgS80Za0vuzFj
l2vyDaJpf4HMqs2Gw/MDSqYEtDXVNJ8o65kO9WSWC4178jkMA2YuQWmOVutyKaZp
A99MAE/yicucCYKNeqx2NnJwb3hrC51+pSKjrhzMTtvta2IM7oHwT0zDcqaPaODu
pEFcopdbgupYAr3XoFGt07KLgFuAQ3S9bFs9VHJgfbfXj2cwniSUPQ9ePWQfdbtu
dx/8gngcNpfbmorurva9fNTTHTqaKFKNJC76i1QMR6h+CxnsnfTQnLVLfpJtWrNm
4ucF/VtLRM1Gz4S2rc/c68/XBxeT5o1scbCyyv0a5fBjT9R15xXVR1GXnn59QEhM
h1GTnCPBoGmeeWZ/fZFRDY1WHvGxoE3Pq917H4rg40P3tSkYco2JqCKgbuX9qQa7
ve1eDMbdkAHRcpmZJZlmryU/D0vghXL/ODLjjR55wgFsa1oVBjB2n5zNnBZs7atA
fzKer8Fwphwdwhady31hkoNlQO39fiO4tdKsn72d98Uu2eSM9+EfKERGbbvxyMJv
QeCsj+/1OB0+Be+3BRAuFKFQhjFnfmluEWi6JE9NI9+VNm4oGo6iA1WiGGqi97FA
1fXuTL90GbL99GJc8v+H7SrldLHPvO6Hcnx2FzpjmcoZNba5yncpPzHqjozZsBEd
puGdnObQSUMAWFivFvB/khtRIstezrR1qOhhj1L6WPESGTLeXIXKMvD2mu5gD3GG
BfRJaz1+L+ZzMcjuxqgpF4UzhwX7K0M/QEGuYfgitHFdTeBIbUeUQVTCou+w//N7
5ZbT54c5Uq2QY3G2QLthxy6VXoDz+Dx3oH+inYEiyn31uzZMYegpyS0PFldbFO9p
KV+OIaWHldreBVz0Yu5Ic9ONelQYc0AzGp0G4nPyrT52bFypHvKRBKcPkov+kWcs
D9XkQwBh/oXEL0orAI20QN3NRAc2J5Oa6bs7ZWaC3I9LkJ0Z1+UBUtdQlXbX7v8R
xmu44nFo5PgTLmeKCxwfvitCFrcX6H86uawQHknUrCSwKmRKTVx3FFfD3RwL/DQq
5TItEXddEwR9rBIHijW+pU/JUA9zjRWgPs9xVMuTEY22eKmm/D4Pm6PjpipcPgS/
+KGvfAi5RHYuzBX+lVtbdmwGm5NGVIhNx6WhXSjqdSBVCnzNt9oRv/nEUKjt90rb
WRXDZhaGL+Rrl//ZYyiArGDqKSdNdXHdlxj8aV6V9KhTJuIdBmlCIUwGWG7BD9uT
u92ydLWlCfnuDzxIk57hWNihGzjxobu21E+d/rOrQiOQEzyOCOP7pfDyoqeWOug/
BS4rUaC5guUkolLom2zw5aS7o5AcXhqS0CTAxKfsM0p5wAUmD6pw7u3v3d8KUZmh
N1LoywI8PxHjPk6NoxGLtNvt/JYW+eLQmav8CsDOndFbYRouM3KYeKV0zJ8024O4
bNsplWrIcLYLT3GEXCbFBf8kJT+5FUpcioHA464DmeXyzp5DH6VQ0meLoWF6iGkz
TZJ8KJfPOrF4a8z6iCa1bYXtLFMmIXMrDzJKzwpfJNKCrzfYPa/EgVk9XGjgikYD
ZFFUEaom4fsIdaRMN1QjwtELVsls/eKgVPuuufcv+94awOZOouSmRKRDO0UQ6cqt
xFqysQmdARPGIQ1mtlje+9tT2m038/sgL3LUFrdxL38HPVGXmlIdkFPQahaZiTN/
lgst7v4AhUn79eaRJigRYO+ma25CAzHtpUbHdtTqM1S5Bc6VsIH3oLC4xbDTbziq
XtpSxyd2OnKfGG3sCMn1UMucAJr7n4odb3mLA/wEx74JSqgQ1TbwGw08IUPH9uNF
pQ0uxDTbHr2QN6L6usaL/LzIOiJNYy/LyrrOq5TOQmC1uYAXEVSTnjWGRf65jXa5
PD/fZR6Sru9/aXSCAaIXc6c9Al5vNJehDsuLZUVszujCbWkcF5lnHkSj+mcg9YXR
h6wsu2uVSWr4j+huW7tBb+41SPQcRLBsoVM2yGY2aVCn+P+fcGDEI4LqWLaMKvYV
rwANJ5u2PxV9iJbvOcdv0Pb2MR+IPlTGejCGIhahM5aOBUGRfom+6DFiZqXH2mHl
f+VXVPUk9tIICi9STsbXx2DiucR8pMweHylLHiFJFIFhvuH4brBZXMW/yMYnugpG
RtyXeNnx6/ssRQjTY/eNWZd8KsL+7Mo3njzYSxk5llx2v3TFB+eaLxtFc4MJxWN5
i3CVjxV9d0bzNBCLAF8Npdb+0LO9rAUp//scp56AyN2ejEs79vj3mTb47Jifu/1b
F9uOMumrHdd9a12bxNMIv3Y7jbH88gTfh/xOsgu+C+6tJQ05MS84h2jueGpzYkmN
6P+4kZU2z/KcWlvJaDnMLIu8DvJbd+0cL5ai/AA/UoOI71HFQ7QR6T97rXrWC091
nUXlAKEuy0XC1FibeEzhy5wN91TWWp8GLxbT1TkgXn16BANhBytObiUSZrYIcYud
QDyTH7dalrMcsPVQyeNPfvLPYVTD1U/biX5oAtEb7A6rlUKMsFuSVLxHRpDrk4fx
WadIEEMOV4+P3H4tIFtFkFA4yOrbJddUovjDkHcFxxpMcHGjCYLhxOXFBONvzGVq
WvMbpjOl6aliNYkOB+3aeALhP4lGxSnFY+BagHYGOWGzsEAWpBirSMp6+GKG/pvA
XgeQybaAnpJ6UAyzJN5ql5MYYnR5YL6AccBrKiU5ho0TqDBngH8OXCRzGsgZa4hk
MPOH/BB9LNH4nKsvUaT/x45Zwp646hP5JSJkQQ9z2m8IpSLO5JHd3YNpgswsf4Y/
r3zR4qV/Fd4ceN4FJMJFb4niiGvVojumSiv3ZmcNB1RkYQHhaSpiMj/h4NyRW6ue
Gybg4+c7Xuo92fR95Tg5FmLyITi0mkBWIOUWZPhk0dRYhjUJUBIZ9wgg9nGsyk5I
UD04Pl4BMvvaIkBUgO9BgzIeJKEVbZ7vToBL1QDhonP8oaJsc7wn87vkXZbt+Vxg
rlb2u0H+FUKcPyahSNWWrZn03YkZmxkhIYii3TjReTnO9BDR4hkbzNm8TLg8rn4q
Gh/oiEZUnnnRmMJ1CGa1n3iyYFc8ZG3ev0Fyz3o3wMYF68wXFxlRabqEFCrins1q
cVlpi/EGqsDKutXj412jnA6advHNoQgcUP5C2PmLsvUuGfDLtGKAMPYjy7RR5A4A
47xf93qnNg8lxB+FszpRC3FORu+KKOnMQB6e5pRUT1MHuvn+8fTZVTVf6TE2EHea
0SLTYZDKrPie1XP7Eq+e5W3tFa8DZMcxzL3qt07pZM03pJIF9IUmflt5mooB+5se
YVYQHXLDYLcY/6f45EhW44gcMlftjhUzsaZgaPQOsC7MBB8HtA2SP7FTfWs/ju+A
POCjfrbRtLlbBon/g5xr0PexqK0mULSrV1jx28jIsB7sX1VL/yiEs6ejKCQllkgw
KfVs9srVMAQjK1N/VCUnjp5/8cmTs3od5S5KB2g/Hl2PZ4Ct7xY7IgDIGCYyWUda
+RPjrvO8cBexqpA40fsnYEkF7S9WDa2x6pZbOaf7JUIrb7ij52/tnQISkxqO4buW
Da7zOZom9jG6h7B2s6SqSEbRiIY/wrIqV1j4u8QXz6TzBSapC8oOAJ0Q4L/8DaEu
u6FlsHgXFi+c6zpaWtwvxEnp2El4FDKBoBPdxlFcQYcWP7/j77UUE9/XuiSIbURJ
3E+qr3IYkxZN2mAa/KFWD4UCOE+PCb7pDPvxWdbQfUGDK0+ud9JzhwF1QRWEpw3l
N6Bk+fwdkxPP+2OtzU2f5QjdtEoUt3k8tDsEvTqzEz65slHndyoItcIB2BD4sAuE
0g2gjbRKJZHQcOn+zUBCLuE657bzET+ENq32fIHcDQlGN+ubkL1Lw0yfE1nr/JpG
bU9x1Vn823+ls3VscUbPkr386ogjmKHkjaiolcDrTRw0+ev3Hz73MH4amxvYTqPb
mYTzIwEUh+VeIKoaTVFwvc2Fz2q/jG7peTMLq03qnduMe/IjUjMu8WyZC96BDyE4
ekSBOcFcvoswokI8T+QzRsnnmaJXnUSZeNZnQiTO+V1G79m9kSPgh8xjqy8IjbeO
ZUVtdun7+HP0UbUSkBEl8ol9SjCIkbEP0qWeQKWBlGWv6dKerRNyufYoPajg99Qx
tPT92/ocUkFIOwLzIMM6UvTt2gd7BTY+kq0d6rSKuOzujjLHmilVNGW36lXR/H/H
XZfJ/KgZd+1AB+jJ3R9YMFHuF+OaHN3GO/KLxARW/Z9Cw6cw1mhSmTxmZRkT7sDX
oejLAay7CFVmzrTLxB5oBp2/2bldrRUnLETGFfdHrUtc+jV4YVCOFMt7QtUvYd9q
d4iLcrDDm6LhhVVK64gf7Yevt2S/l4gT0z7hlNY9QXs4hzr3nstNVyyGmphxv/JN
hfQJvXK++3xbqkf4+KPALYB9zCfmWBZm2/u1do93cf7Z1EkTjg/1fUVNXXC5fS+C
AgExBHVqhOicIXIMHvNA+nRSRJ3M6Ii3SEivoQEyJ4OzNhwYljWO5cIvnlKCqTwR
BW5MSQq+wARc63obwyHO5vlcY40zBiuNl/CxMHBfBh4TVLMV72Zw4tfiAS3HCAra
eUt8EHor6i0x5RTs6Umcwb0UExfmzMdnbOgtbxoolFDSe7yrJ74bVv2XkyYKXNQU
IPeMnJHL2/lmsUcExqFtipdL1M3QFuSaPB1S8ZDDGQpTXKbwsFxg9d1F84tiUyNX
5P0mQVvbtbQxj5e+I5qRDpktLJhMzZQZxlJ7XHCeRsbWQypB2EKrr3iNn0GMN00L
bsT43PMismCZLHkMK3yDUucyB+1PuOgYg1l/EFveaFv8AkK5IlqlBG5kyqKaaxTT
OlYX6s+LvQss1VeteabS/UvvWXQfjTDtBMRxNspQmGpuspKVi1M5aoJPhswyF48K
Vq1z3t/B3gVnBGCz124RSP8gULM90scusjpSTe73tP/t/1IteZaCTEXIvBfzpQmf
NLFITA/Y2pUhTH/3y9APb7v2093Nhzt1Ywi6NT3soWA7Hooq8asjCeWUfYqx+88N
1zL+ftxCOO3Y98srCFsbrAbfC1jXu3ddxiVlEhSvqZHmG3tzx+F5aLiQPB9yZP3G
ET6tnInBXrBZ8Z1aw2rzXJyYr1ZF77RoACfElcHJa8wWMw43yCXLERteEh6LCQXe
7EYQbaUKOC0vrJExj+UBjDL//HaZS4ZnmuLrJn2wMjlGPLNVxgSTaphMhAzgFJkk
CUe5roXY7pmw8XE1E/C+68uxvUiT36OmGVhf+LuhoPusbK7tgTwQNPx+Lf5Z+tqI
qdBoM19UOLC4pngbJN8c1h4ButncJoTxE6RFEUaQwirsfI4m+Oi4hLZ02D86dgC7
H8CoCy14/kZle/eRes1kwVT58x1IF56IxKMpchYmTkUyk1HkvewxEG8MSKQEVenQ
5MTe8onvDhoV698CYCQ882Le/1fos6SjUm3ap6q/5SfvZu9FNK0zRi4vmbJlBFoU
vo2Fd3C+nzORtBxeGBIshq0uBqPeqgQRolLNshw+rlba3NcWyWrMcD0RP+WZGLLw
HtnkaeYlS5IF04dfdqaXhjzRviHpQrBiBwI1zYhbZU1RZxWIbuOpehuXTy3yQvFD
U2VgaiVikIMXjL66so5y2w0Cl6PfpZO/V0tKWtsk96BSLr4NedyLrKID+O8vVZu9
o9W0SCCMPeZf92ApLG2PHg6B84VjLR6zYlZjUzubREgVEoaNytaGHLQtpRFjNke6
Y+q9Obw0et+V0TQUv3Sw/d+W1f4nhLlIuhmT6EnGg6Ryji4gcem75aHJzzpmp212
ET89dheq0yV2bmO8O9cHoQzC/6f/3lkebPx76jYDGnbdwmN8ewMoGFU5O+v+kFNe
UZBBSfr+l2N//vJnTFzf9UzkD34Qm9wSVWkpqDUKyS3AXzP1LJbARSxT1kj3nYAv
BhwrYjBHf8HwnBHY50AI9I5t2jNSOmwdbu4GZ3UsIeG3WSv46tW+c0v6bco5W88a
BYbYWrBCFxOokRfCoWsoQpZ7XKASBjt9qNK6b1D2KqW07rgWL9Mpg+ahfkptwvIP
ZYHN2k3kDNK80EgEuJqA67aKCnmxrv5P1E8KY63LDR+OIJ+tb1CceygbsQY5nbTo
if+WnD1stEGyqMmvDQXDyQ72vODwkjs1Rm6m4aAgrISjzNcDxyrbfkIMeHIe3EB0
8c6hKGLKPT14+z7olT3hil7gUF50coxK0GnkNiz7CT5yMXGQMKkguYIhprbRujZh
zVZkqunN6ZmGPNzbdRF2nvVwreC8lF3aW28TQG0FmF5EM9+t9vKdg1IwTsoBdYFM
1Llf4u/AhLcqNbBX2zySW4RVltGI7mDu2OeOVdc3jAS6HOETKx1eVLYjutZ7NXPm
GPZWCPUCeegH3Q8B/SeiS4fVRQ8muWSflwYYgR1aBZ67Gv6cofgEojHjX+89qroi
depvmKOEVw5uU09+EGBcO78aMmixJbonHCZYc69AUAuNSn6ReYkdMMIs+XOKfamH
B9UlNuK1OCqIfym9fBE1y8n6ofich1Yvqh2USMeVcAFBH4pPmnGrXdcCg6SfOBzK
IFN6QjpGtwgehotRApJ4xmS/+66fRTPZGwN6YN/iwinYU49xyIwCNsGlTpVfK8yI
toSEUlJvl1L/uIHS+bcgMsrLfXUop0cd7wD2eCwChjEkiNStFBnpcTtjP647ZVSm
LDnU3oOQ6RpwjZRYvVQycERmS2y/cahfPTP84nlvJHl+W3r2YiKTwVGkxOXV/vrS
+BUk52xYoK25XQE1W2GlJfWIFfXOjojJhbgXZyXtPmzAUja0Z1n8vGMNGxPueT7E
GyVp2GernRsX6p8v6yi611eMwMLqRnXCbzCiLXKf8I7Nhy4YLMM5sncvNV21gU8f
xdNY2i/nMeQVu8cwmPef2yn3dnBayQoAEPBAoBhJL4UD9QQ2lkZkAdu/N3gjM4uP
icom2vA03Vysw3K896+bjIZrk28YUFfIKofSDMRPC+mOROBPWjZRox35K9KSp4c/
RvapyBA9SkGtfD81BrGFodx2KSsOTrknerF/6gopWjKexY4HnKeqJcS7CqmKCopd
6z092syeJQ2vY+/tlz7KV8HshZbwlU5lXsntgGGIxCSbGh+UiDZIUYTRXAr0rg1b
0uOCAjo/FM4LZa0X4B5XjPQyFj40+NZnr3Ve/V0yy0mP5apoZ2lh4OsOLBdOHRbK
v0p7qXp9r1NDmFR0dds4piazncGd8wr739TXO2s/CKbeOLIY+wFuNqeebQH6ddfX
sRX+ekQ0qYGbrvmiMTQYg4V1PXniF2jeevtUwKP2Rf3tg8LF7MgcmXvTIap1yz/7
Ue8ZMx4FCm6vszuXn3MyWpRTTTXgJx3yU7VpXLNNxoiE1O9Du9WMsdO6r0RZhGpI
V0w8Zd1INyw+buY6eVcjBHAEhqayF5GbIYMXL/HFqtAyKvIwwQ5vDW3sKLlrtkZ/
98bn/ub2V414XdRnM8OzsP3G4HOs8UsT+QKMb38yCLf/49RQTLe34YCgOSK2nQly
dEamTSvZhPanCrVDRcib2RimgjXV9OyZKhD+lrCRECYrmIc0IWmLxUQ8I4TEHiBV
2TJCD3QFLx+WfcZdV6CWf/+13ckhF1ejK7GxZEmKEbTq8FsLrM9nc70VixNJF91a
H6qpgRitH44eX4/Z1Z0R3COOLGKWbIBewVPMRqsDl373fPyjrmamSxKYw5MU8/8A
PsIaKUcE17atV6lyMEWiIX2k9QNza2zLEQpnf0zrb+1+lqZJLpPX3bjbpe6hYwsn
YF+jB3UailrGfCvz1WTIbhEHZ6Q5DuXghFq9lEiFGRkgWnoUQmHU9FHNsAGdPy6Z
s20at9fqMByP1tV2wJs524fdR9QQJ+gm5qwqAKx6PTaElJlhUR3h+0eEC1wxItLr
NA0y7cYZsFG6PkT6PGjbp8NcNuI9NtsF8qHkASXN1kUPg1Cfn6roum7IzUfMp9+M
qzcAcskjtpZBCdoOMEUlZ+MEpP+3UX8kwANfcLlPr48lyMPar9sy8sp4AEEttxI9
P37Ti9G/Haw6Bgs3T42IVkDE6PZlX7vtz/HG+mOZ2UIbJhLiWY1bKSlylcswRohy
E8Tb74+kKQEN9GwAzLl3iwcJMQKqzeRMLUyRx5vZCsYdXp07ZnD2cUBZQFEyOpd/
Fw15T6Ikay26g5VZO10hiEgY9Hh0OjMIpblcSaC6YDvO+KJ0f5tIS8mwzofvL8CV
dyy0OkDQsDwqiEmAONA6h/1SWkFGHppIbz5R4D9PUECyjTHs77swe9kZrO2XdDUO
d/Ge0iXhx5QoAtDeGWX+4gJv8QW+k/4yHhZZLKDPH9FrUjVBQh9RCYY+KwhFMXzH
/QrLGpcsehmmKALZUCwYMtrecwBp0SVZCXuZShh7xmSaLXzQyLIstGNz9P9tmEsY
bmwkcG6eH07BviglYmzMA69/N+kg2QuZILDFndnsKBvaYo6nrSsKqbCLqxldTPS7
HLE8K7TSzP4EAdEbjzZOdoWRKoQhy2hwiAf5Oz6SiJX/j1JbEw8PCAPjh15Km2Iw
Ayx590uTKXae0r1jOZYpStHWElbORPPEandkm6aF3BdnYHgCI4DwCFOv5berINJO
+uIXECu7+TjS2gzWBAoa0lchaxVL75Dwg0AQfu5ORKKzutzy8ja1sXCenaBSJKvN
za2cOIqrUgExsOu72F/vyXljKmmma50odkadeZ57Rt/OpWrzUAXWyxclY1S1NDJr
ZWhVt70V+QSspLG74aIvYuX51uuf607QdNle8BxvaElu0wyt4/wiR3d2/DMmbWYh
4q0VSIESVfOSpIXKT90aTsnPvSiOB5rx7lkJsXft11/IJd/EBPhz5Zg1IjyyRqls
H+M17C0klqG/x/YlU7pAfMrqsSfdLBouVMu10GGcnpMKGU+U4h+NddNlmFtkrzlt
RfLTRL0MtmVJBA/kzBWPa1g+yPpjZZLQ9KP1+AdEX2LQb+LjQ2vZe7df8+rU3hmj
fW2PKHAOzLdI5w8e2yOsjdPuljtddbUG8lkrwiJzTZ50cwXCOpFGgf7gt1QH33Yu
unKT4+0/83/K8Hiv5yZJ9h1uvQXqsdtb9XntBh0ttDNtAhv6PQ5065NZ7Tdph0kN
em3rXEuadd3Io74UBda6YlbYebm1XtwaRDx5+cV7G1c4d5TKwzAl8WC85nNQsboa
wiaZTzQIC2oIxA16jbrctRBNHHRmWeBy/8jT4YyyMpO4v4JsPTJqTW8sLXzf7GEG
lwEjxZQ91sKzrJR7COqerDHuogM3TVWfVrrhfJOI/+PeG9EbVe7ibml0ar8/cmjb
YswhGi65WSPV4D9cw9f/3GgzM1QjPp1zsHkQQunFXUDJAO9X+kdMaAfLuzmuj9/H
iefKcsclIHO1XVLggwbuMcRlIIFAGqFCHMCItxaagRo+V3QBXEnkVh39KVtB0gFq
TJxc7OWW/S4tIpcalfboMnQ2UnB4MXCdA5d27GneF/H/MQ15N3nDXikQ9NQ7Kub4
2JXsmjx+sbB/P37awGvUkpX/TRYwHEvuzFbUkCNFGsINmm26M4INleiaSZSat/B/
TCOIxFCyx3Tgrff0gZ77L8jM6NfLBmZJhZc62xKmuXteeKtMHyD6a3P8pjBQ3FK6
te0NZzvQ0p4RZeGF6CkgoCbDbdv3GTpom4cbixrxCqknFGe3Hgel69cUzzmgq5o/
2pUN8w00awrncbGwfltsYf7BAhM8w7L9lHIDqVMveI+FrBspAWIStMcBI6zYLOry
plbTRUDuG2Jk9NeubdnAO+TYyquv3BKPi40zT06/bq1duLqBEYf1phAcIExohvbg
VXkYZNhZYJFMBHsy7b5/V8pt5dkNvFCzQ9mj9+WuiqGQjeKC8vJb7FmlK4P0sonP
4/S8S4vmzPNoUCvNXI+GfeI77BoP7nhHd5Wo8/psH7QasFDRteorjxSWAZ0Peq/M
rfjDGIwWynjXoeHJo9MNpAJBeMPkgh4FK0HE0KYScZh60nX+hVXdBfjloR+FMcuZ
IAzPerVrhdkT+OCiN4KZ/frvfw4hZ73+UjkxuOHjY4of29icGPk6BD8KZe7Zq/dA
rYuU5rXfPl4HiX1ikZqiVlTR05SJp2B5XMP7QF6T3KSUNA/u3MOG6hWenkzgSJdy
TYbGvRTZbH7pCVHSZnDJAM6g+zMAs0Nhm0qQqQWC8512SiZHHF0RKxDpj2z5roxY
ZJ+1GbllBsAkGKgupj81S/BTrqBcImnxDc6MfeSL9f4F3g5hxCqrHJwsSEfSmHVA
/3bZPF8n4R5kmmzM8Cg+T/N3ZIGafg3mM03r+oq4bQO4T5idLgJfigbUD6cIRFlt
8BdmiLMRfYOE10+uHt6vPq4TYH8jnSkxWTan7snp2WiCPLYQwR1yOtMH3vwpTHQ+
hxB9jqCOD6MpI1XwsDgpYdGL7ROm6vymTVcmlo6+qSh/lIAtlMz15ngs1ec5DStg
Hn4NH2aFFdrtKjQXFetWpCaFbHnu34NK74TtYwHwt1gxndBW38ySz5uyb7jgtf8T
yvXzNTARVwlyiYJt0wI8lNeHTu56M0tZGZIiRoMm7AQ/MvrTbaPtoxrXQxgqpOHa
jJ1PEuE40fk47+eWC4p0A+F/O43Oyks0N0cY4mKjyDJx9+gYtgKPM6LZGTX9k6W6
CGEhzhBbcJ6oOAqv7g6h+6PteKuvRSAIxbWnI6YHfsKF+EbzlICNhmc4zWOwF9Lu
t/fCH+e1CDjEygAgHksw5GUrf8jD3FkSPDy6YEryshraAVgbeDD3Sifca/s1qfC3
fHtS4NgH1AcbDp6WNRkS1g0z2uZT3V/Y8SfAFm/3Z9gV6pGhI/T6IHPYmPwabIf+
5YQUfHq+xYlfWvl0uSpvlQhtFNvbJN+MN0mC8QppIoUt+Kz6gzHsLNYYcSgmAn1P
I0SKcqz8e+eNhVexyheTBkfHAZJWCsbypJd80pKtZ87IPb1MXluor/KGPRBDf5kh
fuBKVxe1Hjd+vnDdIU73qwRwGuuzPtu7OwX7xUeG3nB1JZwZhjKPXlbK+CgxnxNL
oI7vYpkmf4+B1+V2SmwbRwpBTzkWQvRLAjxzl5GOIvUhknK+gYiPlsSoGsb06eTq
oJ6zEXf9IJ7VA+Q7fXUjrbSjXd+UWTzIxemgIiWyJCEO4StyD/S9ykqM7w1V9RDk
vbRpH51CorfKLgr7I9S9yIsU8K+zuav0rX2lay6rH//J74JlzSOFsP3CTaF4+9aG
L4ggC9vy10mivGPqI+rj/q8UAwcwHsRy8Rl74UtHAL9F7G47oN+UZWuf30t2znEP
m0V9nHLFnyHOyhUOOPQGzNzLm1uz7hwLuDjQPhbo6bVFHXAOkTf1XHJpZ9C29oU9
oKngSkrT1NqAotQP6KmFAbgYc1zwNaPUQ4buYdjkdb/t5cfrFJS2rCgsTjLfCa+7
UJ0YxZOWqajMYOIBBgQorqMsCLicEMBPRORsotNaXRGeo/X96RON3YncMnKky4se
kSsY3L6lWN88Mzk+uItbyxlQ6XX1GMlto4CL3RBA9/Mo3QMDC6FcOQ3SpHu3XQGh
lVQNVg1YV6f8PSd8uxxgG7tlQZ6+VNS3eUUhTwhKZ6UX5CecXz1QOjJeXQws7ANB
ViK0/a/xXDJEC/wWglVm+ufhXzZUdpP4ODSzuZlIGIjLl7ULCljeFX0Ln6wRyfkP
nTPklvqOF5FDYE/c6JEYZCPgoLW0PhWKeCKBk10yNTCBnFHDhd9ziIWLmm+HMhWb
5jXKLE6VDbikj1mVYoBGPyf19TJ2T8Va7//yg8e20ONCzhcNJqA2hZ6BMRwJxype
VHetpKdpcooGHTeryNUpeiTS0YPwq9pESfr48TBls2ujj2YG1TpDYaBSje08W08h
W5tGiWvEcml9zC3IJ5Tu9XlD8sEsJiVDMKpiOxbQFzKimWS8TrU4KjaBd8pKe2rU
3apXIsLLIbo+ScrG59MTnKky2kxTSY91IKBKH+kDz39XxwVKgbSjFJrw16ZAWdTT
WnEKRRzGphGb1ASdeQt6GJdP+uPE6I4Lb01HpcnsIVG+j04JvqRWCYhZScAEeNcb
no6YAQIXVporX/xP8bOWw/3Tg+U78+l8X+44PMnASNungz81ez4gxalL/9dUvG2f
frwScWf4KYxwO4oJYcY3UPTvkFsdlzyn2QNKGIDIOXqPXeNjJhJLNTDvL8zhwvjr
MK1lyIXhJfXAyNoOmN3ZpE2YZjWgQpMTkfo0um67cFMneAMgQzQaGyrcJAccIJde
myM+qgr8x/WgAC9/W89CmBUk3LN1gcjyD6+1HoojZcmqiei/381kfRLWIK/+UEnL
HM0A3N8oXL6zEVBGn9mGPvBjybKKQET0JRJKy+7LidJA+H6+XLuInLkQVgOuO6ec
roDDQhuDlNLSPAqm5WrK1mp2PdNVfRLFtHCyfOFl1X4vtE1Qxd+ouyBBS/ePI6CS
5a/1UaOPMIf+0RXRU+UDRfaOAgcP/6MpAsa+AMQrVWprEfOZPS95n4uNbq6XOhH0
fc9L1ybJlUbvpNYVuHwaDU0pke8eVIG+1ib7SmSzSq0z3+ioWj+ISc+JP3EGiCql
scomV9IyqTZy2rjfckxe54dGSfAJJUcZrn5mNbrT7S+QnoSgQng5Y71aRABLtyLV
TAO+6qv3BYjZLEWHZBOLJPH+aPyiGgxbzVpW761AO5JhzYqioz3PwuTHLu2JiGDV
uc3fNXeCnVD2hDtEqzoS5a8Bz36XqCnZ7aaOX9/PNiyeuyx0aJgHUwEY9AyE8dsC
YcNP6V1ecBgVMfs9yee8HpIVOFZ7JdCPNcUNyvZUXNZT1APeTZA7YhSa58KUiej5
rM3Gc1lSl2ViJFsmPTic7WnZLJqDnz1bt8SBB7+EvFHyW7snFfVvpnK0jFOGRgqd
BdFCxSrfhRBRGqy+ikHqIDFhU/nW4ycXPKWYqbYxvb2jufjA4oYmPdkFc2L2/NIG
RhJ1jHVnHOmRGrHTanYX+9YfC2auWoFtDU5nzeisprvQbZGWWHa5EmQAMRIJmX6H
yIggrBxRDzD+WvBtWkGEhT3WB9RkC3apEB/nMg5nQ8LxCOIBBLkU5xrWhMFziz+q
a8RjXVA5R/47c55yTQ2Oa5QZoAQOXCc+tA9wt9u12a8SzQ/CnV7liuZQprho9sV+
bqBNVpyjr0rwo51NcRXzmkO0ri7vt7QIjqHqc3Bm22beTm/4QZNauYq3nXA9vy8a
RGtxs/M3h8MNS/Y3uRHzdOZ5jbuT9X64g1uDFkQgWR/JjJHDEsr1f9CJn0bSV908
JMh4RUZa9Qkhb0h1RlnR0YoFgnpcnd0KLu4z65ovoxq26ApQ9eYpyRPdRlc5/ZKe
udaKBy3UHQTsWq9lXFo8EKuoKTwP2GAJy7G5T/grE1cpsImruyTRSvyYRcP0shYy
lFqv5TOXEkIXbL4OnvNqMTE1jl94y6j50MmzMAGN4IxTndFwNpICd+Y+qraZZIyG
6O/h9a/fPLCrXCVVyDD6ByLvSBZmLABOOkRJ7c7hVcAEUNPFvwiJk+okwrE/Jnfh
8z51k5uLJtvtsAeHMvW+MNd38SQx1MQgj8dx47LRNR998O0Tu3ZftfzogUkBx9uZ
2IWv2ggOK35dkotWnIBCl9L5vASIhHgngx6R45xiYfq69M2BjdiSTRUUgji3dJup
53i4qCycx5fyizeR5BChuFvPUuMgtyEEjqDzAn6ytPA1hArxEy6hOtFuPstEW4X6
CGZj7FSW67s6lGjh4JqobftJXJbCHOhOnL4rBEZCLj1ACAGc3KQ4tOm0d9Lc4uZL
eIujHuXA2gtRS4pgQiuI9bgHCR9yI8Ug6sH56an+2Vxw9HAck9pF2TFk9ZKKyrEj
KFUlMnZRpcH/0uWm2kYuePJYz0OWriZMPoFkPESqzHqixRSXm/wpvYhlFh+bMriW
qEVrmWu8c97BhI9S12l018gCA3XKFjjYj4V4NzKp8g7P3JMptY+wnOWTffcsQxC5
3cs7ELD4Y4BkWCZBt63BsaXYMMA7NwejHTtuZry1YGJSoLlOCLI/g9HdannWe+tV
MZIsvJ22tpmZ6PbBBqUZJk5CGwjdP1YJtXyIEFZdRYCvZfftTk4gntNRoQ93S6Wp
08WzXNzzQzOL8mT892zyU2NiA8Nf/uPy5jrQAi4u7pd6j0G53q4e5ndZ4G41mmrp
u8iAzZ9DW4dk0/KMSMXHTVt1cz+OMdC9x+OhCcBiV1Ux/f96z4OqIn81SHL86vJ/
wIfbA9R56UHRLGoHlLgIAYImiyL2JHjjrCkVL0U7z5RkPHibIuQ4vldbvcwq57n1
PLbUynvP0S2vNjnfCvnQb9vH2oDXgpXocdM6dOxeT+NL9ejWswrEIHbd1274wJWw
YpNAImaDUMdmRgg2LNSk+FAEI5Etlm0nj6LCezuAt1vUpRz5chBGb9nJLXz0o3WV
vMYA83TQ1czqR6SLJAYVHKOFAZwtNAW7lu3UBuncdJajpg9vJ93KO2T2vFcs1ns2
0oT7E9WI0oJvm8CIKEDrS2JVG3o63ojPJSJSpt7IznsZfI1i+TaVffZ7suRFtCha
DyZsnlB/nz1/9NXl78l0HIb0HJNeFw7RmRM1NPQGAy73b2+GwCfRxO+ZZUHYCpMA
OALAV4Ln0wpdGd/MYjQc2ZNK195WMpRumgTPbXNv7xz4J0sFu62Wz4BSrUfHSMXI
Gw5DqfAtEODbs/W0TL4v7Kd2IFbehlxWTz2YgqGPr6L+Z9tlxDqnmvETWe4MLyy0
6K4uO6tebsG1IrcsHvmCgCsgOGjf7tFZ+oNa/3JOABDrKQHZsR2KCrGQQkBsh/jX
tiZQgm79pTlXBtAIr/5NUunFmULlI9zKKK3tSLjGf3Kfavk+2QZ+6gnSwA8+Idpw
mObD5YR2WzyRqrxOGKTk1V57zxcKpXV3HWZfomfo3sCMXeQVA9kGS5m4aLDvUNG5
6OXUNiICXTKE8aeX7HnzaPQOUYt+8PREbvqyv0e9BLkC30+YqBeSptFK2M8RoqZ5
oRw/omoXokpOxNxJ6ZY4TQ/1a3i0/6IrYkSxIx/NmBQMxPZaESg0gyLrkUI3l3u8
4PekvmkRvqUtTSRSH2uoSz+Hu5ibf4ngdaIfgFCPRW/gt5HyyGsR8XP/STSXQwBg
C1zkiMS/2WQKJpwwtC/zOmhF8SQD/wW+LR3gJ4oJ/U39HNGAtDF0lnHXbnngQL1j
wxsuVy8OtEkr7gqIhV5NHQSlogQhWyuNB2xQgXVl9vfT8L/6DPJT/ixThJt6g6i/
HSs+sme6OBGTfwUHCZa4gb5bQiiLkuGW4V5KYs49afV+OmdLgI4w0VCeMvHziZSP
XBUHPZYc8godZ8HFGCeJkhzdDLSM5NS+L+JLVQvSiwMRzWXp/y7+20UtFGufubMD
wUsfVauhtSyqdCEdN5dhTUcTGHEPZbIQKYT9vrB5TWch4uYcHrxH00YXjbjZP48I
sGY3VcgCU5mwbY/vsZKTYOzatAgnrv1TpgmajGg6T/UQ0ByI4RpGt/NYnvRzLI/M
CrZtJqbHU6cTOlAcUyLfGJGewrUxwKDXXHqY44EVFq8Og19vgOKDOGSa8h5tBTbd
ovPCZFg+4jZV4/kHATmO4sEoBjuWQt7QEk25fIUcG815NgK/Bd/rtN7irS8PntZM
49QEy58Or0OHvbwoSpRomrZWPQPI2nLRojuN+mAle+3vqYOqNZgTMK/o384YdAkE
ShOB7VfLhLNLlN4a8VR1Yx/94IPCb0BDHSTeGStH9OHJMKcKDGMlK9WKFBAdvToB
NYz5smvdLY8UnHh0UVT89u1LoG9kZtVte2FiazTDc68h6I0BJPzqoxXfTr9UcHfl
w9/OtGthMvp93ypNFUqDM9q9xGlcQpRNXFaehc4D85xRtoE+3Cv/4VVKDTyWUA0O
ofmt5qvaMiyB8BFcxyNjNBNHo1TmjuMubzC21FGI8tDgFp8jFpeWs1tIhF/yywnW
1i0dW1C+hY6g0gO9RazFw6LLZH2+vEZCO50P/9Zq3VatUU0hVah4wdFy2KJ/zfzr
ArSwssZu8ZSynJXHKY9AfJWEZaWmOnh8EhBBvVnT0cHfR8LSbwJw09ClrJLdNGaw
mERP5YlqZtF3XrxnUpm+HP9VDrEeB+wsbUndNcPaP4Rk6BfT/qGSx9NqD4K6hach
YE6vm0uTYYM/oJ8NxeKittH2FXKTfm0kek0GymhRlLdYJBDNPl0Zafbp5M2fjLpu
AVgQqCP7SKPTxDoJ2Fp+XxPwTIF6abck5g4PhA1ZehVSc5g5MIqEg1ynPxahfcBX
YZSSwDELPrsX5UrcRALpWTl7cwFDgo0t3jhY9az6GyXLDs7HqfayjExAeJ94i0rK
PIypqwkU1CFXyVCjBysw6Yn17F1Qkb7y5sqic9nYgBte4vi2k8K+La6e1PG5HB3m
KqxSpd71zx4Pa4xw9j6U6PqFf8mO8C7twJ3u4i+RxlP+JOAtwgImaiycFdn/RedX
zDZmbsr+s6ampA/4ExqI7RHjZVfcfQ2U1Qg7ISKV/rH4uZCZx6wubgS6XG0MBKL/
mQvF8JCKZen7CFH/roOvlZjDS8GgNvuGSMtbYePCgBnoGjGha49LVlWOfr2hEgL5
AbFDGsbt9l/Q/6V3b4hsK0PouIZQdwfEn6aXoTnb4w6GbESuhrIo7B9zG6vQX0DD
dAvODXsKhutsRqExvInZXv1AOO+3jylNFFhFBVUtC3Z4QlIbjYiifLbl/ItTSpGe
Mc/hXGK9P7rm/dX+6UAob4GLZ1TbpnZdPoyNvjSfL1mF2tpkK0ZGginzqxzvG8k2
PxgTIqIMRao1zjGOhQdwIiHIQQ90FYjt3c5MKtuQhyq1jEl08yC+DBDmWRs8guwQ
ILNO1aPeBdtg1BgKn/1tc7YDSGxnHaTP12I73BVTAb2qcBk9IIzMQb4MVhyTm9LY
jhpmGynX/4q5o/2kHc6kVs+ZfYih1krLcC4M8wXE5msy7vvgvbZvjOCLaB5nGevq
sH7+whjgVTBNrO2Qe7d98vCP7erH3mJxuwwoRIjlL3KYBeu//rAT7d/9hls2tfKx
QlUBdmTv6kuJVAV6bBoNuc1STXzvGt+YorSexjsNtDbIL83BIDHs7dTnX8E9l4t2
ofUfvtFPbwlZx78jALx4uxeHSaazRYXPQZwtNpoxtEop0CxNi2PKGkSLyD8J7Ygd
t4F1siG7rxxmpbPb92+pOq2edVVoCvwHq7QjltZ2t1WSsn/YkDatV820Tf83mk8D
i0kM6Zf/+45+yGgqYA4ghXPRNgOmUOopyXDq+UW7iouNSUH+iPdPVeE2eUfQbICB
dYVaFRtPAWGaMlBzFRKiJPwGIBhggB8OnzeH+5nYsA9Fiif7gER+lWv1mjBnQ+MZ
pjTL7qQDQ77MHVTq1aFH5bg/Bj9TctZNJhxyji8KDjXXSqT315dY8DkTHAfSknWf
3kWDJfrHNBamiSCP0OURJ5wvTTQHAcxUBpQEXho7xJnxUMlGT5FnozMqLVgY03u/
TrpI1mcSAI00xx+jQtLxx+Y1/T2X+v1mzPxuoUZe+COwZglDBOd2abESMq6oDBrt
kaqNoYYxUiY/TEHQroS1QiBtKz9YUUNMYGT7Un0ZK8a/7ABH8nub2Urxh3WCmMmc
axC38409BXogMTFBWZm54WomAgk2WH3mHqj+QCqzVsxpDbe0S5FZ8ha7EAgsDdyX
asEnP2FWQ+uZ+1HIt5rEp6LiW/k2TZP4hRZ1vPSTyEyatgRnOXwif5nUhZJOnHTd
8Eja8Bt8uhdCBC1u65IWq+rh+fFf4MORUdD/qZrg9EuOGFSadGWF5LQmGLZwYRVC
YHfzm1r0P0qbsAhNfv67aheFnEaIvdYUmDe087ul7JZNXHcXRUUdmc9qG0y6JLrT
dRVh9EgLRpgnhq1dQN35Bh/C3C67jb6V+4N1uZiWQEr0YJbkVKo/uevRGwmyYcxF
XTli55VJQdgS4syZ4a9TI9zh+d4fEciwt7xjWAc6GaZB+zvW0ur0abwSXj2plLpY
J/0lKMNhPsjUEKZktc24q2wBUREphXdpDN0MeE/59Sm3ZrIECYD4E308MQx6IHSk
VqAoOG8T6I7NZp2lKBMGGD7bpztRtoFktmaib5MPEXhbifgYCGqiyZuZyZSifYOJ
5QpwQMgmF61ZWDNEiWS4y5gxtuZF+Yr55Yv8GB+DlrvS3GDxfR2yS3T7q5xW3+NW
Qk/jJ825rr/Cg/W5AXfhqnHamexStDk2TgUzaBr9m5+5T6RpQAJXnNLqLcdqtq3W
NK9uJISFEXQu7DyCqgtNeAE1jUQjP94CHoezIuqlRHJ5CJfjP5qlLLcQe9pn3esf
8MK6N2/hR0BvYYK/4gi/RyVFVs24Pb/eNDMRY5lj2OqR7s5JH3i6sCT0BKbVWwee
weEE7yPG1ZmqeA9LCpE9/9hKW0i6PF4I9YzVzi55xAWSpAR8iPkWLgd/ftbaZJy3
d1YeKShOHJ6ySQkhchXAhtGMBkMmEKRvTl8yyJud9H/ahI0P1/EBsvzK9NIOTQ7c
gRxsbCPcjCcbSyyi00SnyuDPQZ7ypoEorno1+HeFJeDzG4fJtb1dX2/7w8F8fzMs
Pv7YR86zIHX9qA7O5u3cKaNnqpqmmGsAaB/L0HWIliWc7WPNfgFoWYYBNlwDZA9m
cpP1xetkzKCSGTfXazeMCIstJfkuyA852xd3SkqGufhDJJYJxq4nKACmmTvwq7sU
VMGkFCrbOf03kQ4b8EBNz702hUghvGlh/v6PXvcKfjZx0HW28VULpZH5aqdQvw9C
eL+i6W4DlIzZCTUp0N9fq6XL+gvscDY43HhSKr/f7jza5thU4XvR7aaUnxwG2b0o
Bo9H/3NzLekravsnItMES3C7/ouf5T6cXf2nHSFW6jEm2q3qus75CGEr8yNmzU3P
FJRSebmKXI4ncQldNtxsGsPIo8OmnNWfOY0yvPWxJhgErPpr+79NY0lI9W8nZuG1
lRQwIp/RakaRJu16hUqaPF7G0FSnJQMkT6496wBdx6ZpYyNgBJyUtxnio9KlATJj
h27vK65Eqetz7ock4hqe2/ql6XU583qvXcrzeZy5qZ5tSnxTh8ps2ImC/MN9DFED
Dui1vPkg79c6VJy0z1Q3INfjoy7wIo9LWvRPGV+r0PVrYZrFl0lrJMV6PEQINpmI
Wv8sJd35lh2HlCSbUo52fnNFFeopDGQc6VUAwZO8RYGz9mYV0OoOpm/GvnXC8i3n
G+kr2JIBGN7kgD9rJAuAM4+XkqLNW2ylAEsMHOvJrZBmG8Txu/rybtRe7ZmygIkc
cXZEJKFNMpNAqsZhxiaDb5fLd5CbZ6VHlAwMz4ARQs34T5glyqlSMiUgy6/JaQ5S
+njj0ZBD2nCO4k+yQ/rEoPPnoms3fWQWt4mYUgHcBzLPoCFBJq6hgDW3h+9O7Qx3
Lu09iHgjmPsdsxSm6gkzXjGSkUtdOGEixGjGk98LJJljayyRDfpILmjT4DKxsuov
wIAu7Lxb8YWlBn7BtnkAwKw8qBT3wwiyDj8DtqmrC3bW6wdtfa13PDlIOf1hzQ9X
EteCg/Q8vlmNU1xzP9zmBw7A9NzH3GVGpVpfGB4RZA/95HoK9gMctBvJoAh9PtSI
FUqebcmnlpjSiueVV5JTvN2KfToxfSZ0DD1IpH8tdsBv8d8ZtqxqSWJ2r+y85Y5m
Vb3wX0WYzkloGOW67FBAfxURpeLFK8QHXLICBbDfqMVUhg+oD6BSydreY4GghA+Q
sk5xVwcbwr6PF0ii/bAKXbXsFO3C5IzdVIpS+MYUxXqNGJl7bbXyaEjZIlIHN410
os2KGWB0BAknaVIPZ8BuhT1whOl1hXQtKF1TMLwOpe1L1jI9P7iDW2MMeNGzCMCD
i8eFLQJo4gfEmI2am4DGs53M72QdPdNwPREXE+aSA11eaZ3n3Z0ocyMxMUBEvv+U
WM0V0VSdWJMbBduka1aNgjJN6a1aiStVK8uOzk35mIINIM6iAbuPNrWhBDkl7D8C
lMLbpdwSRHDiosib+ItH02PGI4+Tv91ylVbvMwsxNiviPkkFwHPlxZrFwS29lC7D
I5MV68ZjF4APj0ayHINJkUzoaVH6k1UODuPJKiAxzVZ8BuSftcDlAaZAANinEaRG
ZHsiVazlvF99hCl8tpRo6YqtuG97IhYECZSaACIWiFScnrc1/9zYoWIVzAWxneRn
pAmGn7bjC53A0mI2l+lBEfnGkUZ+sUA/fkd0EtLq9W+kT1FMTNZt3PNagrErLcoo
0NAHqsgIHfchPn60anxfTPXla3+HNrRgQLxxXjFBFfReUq/ZYoPT3qXAur/ZSji3
tSH8jfKVhZ0jvPg4OFqSTklZ7YcZEaNZ8LVGNt0yjavPE4/y/DC82g10wjbthaoK
e2susMC0wxpKnfQDf1jz7HtU8DoYAWYJswgH0tVWMOdED18+npDfU5yUmXTrbr5q
IFO4/vZgU92COB/Idus1UQfHjd8LEosuTSjw6GNDmUpWDVR2hPt6nToCxQfVlF6Y
o0StaC1KAkT6OvohlGzcBGwH9FcYM1JJYJoltaacP9wdI/kt7HOuXW9eivCz6w81
l2dxR9ZkqJvVPtcEbyGTfXztT5bEcI9u1ErB45e3YdNS+EbM88tRExt/IQByDcuW
eXSABYutRjJkO0GLOpSQkpWv3lh9fv5o5+XEXz1c0MGEUy4wwK3fE879uEV9U5kp
6dynw3WuoZk4ZX76QvTS1XXciwvCTFj0maGbp5T+XIFerUepRFgMmtChqhH1D/6i
WBzN9IOwaE6IMbwhUlFm6g01CluDEiMBM1vi43wXURSSv93/eTw9lT/KFbsf+Z8m
E0EKgHvYuTnwLcaROPGzMG7fDsDb1QPAtEWdoWxGbBG+dj+cNiGKBIZGTlSiiRme
6KVt/Ar7t+t7sdoJ7vGpbu5ugjs9iwhZh1fYCpJzHjT9sQFXCooKoEfbO1vZDCTc
yn+G9dZAMvNA4Eb5pdnHPskowTIFmindJ1StbOJ0N2buplGYV0LJ61ohp+Wv2QZR
JimOBHffPduLTNQ02+kGGukEBrXLftS0WSLC+jW61IHJmuK6V1VA3TFszU1A8oEq
Q1dsfbWY6dTCLPQWnhX9YOn8sdo9mqj3sQ8VNKE/9IVTg7RWzXxTbxFXDYzqE43H
X9M22NnbIuV2/WnUPuxR0Hry1mLWJ0tKV8o4aNjxCtPxXgoLsOYU9bWZ3p7S3FHU
PD5mWVhodwn36ax72nu3v4yWiE6KwthNvSbAQ96oVbTPXauBEWAolELPolrn0fmj
/gmpZazI25zn41UmYXToHYXTC9JDqg0ytIJjH3GoA4gOkCVtHqerkdPZ5+Tf3lcE
Xc3cDZTc7WG/o2VvEFit0foKS2y9jxtV7n9wrgrrS+LXhl4cZ2It4CTvRYYYH9vH
DeDGSCnGtGrvldsA1X+YyAW04qJbFBG8itS6ahFvMoO/eFFM3rRFhHsziAPodeoE
M/XmX/huBuO6bDFbPlhJt4izWCGATK1za8OiC/+casQnhPwQRYm5mpSUOvkxvYox
55m4BNtTZXlYX8NQjPG7J+65Tgyuoly59SScmUgVlGU8Zp3eHPS87wwHfmo8LEpp
hiA0QKvWglEVhhY5GdAedEycyQMhz5gJQBN4thVB3YCd1ehSVF1xKLGh33zT9vWj
BJW2kJKTO069da59wvV0x12NTXrtAKr2rarVP68n9KUkIoMZhAjTcuk6pAt59QVo
6qof0JxnIpZZzeICDDc+X/VeF/vm63I1Lne5OIO+sGHO4HVN1X/f4SWFKmMpix8j
jhuYi0FuXgu4PIztyLT4npCtfqFQ8vK+3Kcr7U6Gl1tJy8RL0YocrRSnjYJFhqpK
gmbCtwnKtnAAIGs58ASJZFW1LYFtcgwXhiZxuP7WqMU5uqluusqeixdrDyyzQcrn
jP0ZjGRo3D9xMilBf7wpBq1juB3xOUPj6jveqZnDWehTysMnTbo8StZveAxIdlTh
r2dKP2nGLGxP+j/oEau7OzU6hH9Z33QvyDiB4LbouCWDLrhoh9w+7modiUQ9ke87
K8+YwQWM2pWFIMhzO8bzOvXPDqdxWwpdRXJvejCW2S268P//HdzPoKIskHE9xqot
xyGgxEfkFXc5hUaRIJ8An9OekBLQSKH9aA8i/ubeVxHXr/HK5Mwv4XsPbToErMkg
8SV1tUn+T1G5nnQSwohyQEinDdahj+S4o+LHOXIqj+IT1wwEyvn46G7SqeWXMd58
DjP/PDfxfQyjsJCq7/lzrwk/birwK1IcKAQStmwoDzVss1Vz1LzJctBOuTOHWWzh
rtygroHNWyVS9EVQ3TLn/srj16ma3hIhaO9pBxxcQZg1jUytBnJsmSzDsoRa148S
URlqfW7+VBzys7aJ7Bfe6Gbz/cxpKjwT2J/ahp5W7qMwd08suMc3TnrYe/WR3UwR
SUoeLZKvc0yRC2XB4znojklg/HuQ9Psnowco16NB+aGLR8DfGsVc46mHkbzoouBs
alt88QshA+I2zBL6BfiFWmufXApBvgqLr1ZETTNF1avH3SLKYVLgnG7bonqmLNf6
T0eWYJMLarwDHpo1PUoauu0AwZr+svvea0nlHOgSJYoulCkfWnaybHOHM+aEgdkv
4oMxxfSrApcGGdkokJCT5d7TnbaxAcaSU231n8IdNW9HkUM/B6zsLeau4oKPxG10
+e4uzBSLNdR1Cv9oMVHD50KqmuHvE5NBiNfHMjiMD9hCAchBnGUZN5uPODaXmD5Y
PhbESPWbD5AHEPDjWxINl6cwmF7NU1TJ4GaA20WRMOfO+5S13yqM3+EYM/TYnLar
CzXgh1V64S7YbMxwOVTLaoWfhwl+TzIL41AX5keoopczKDuXO74CfgprgzHnJxBU
oUdKLaohP3cjQQdJXqTrKc9L5AYXsRslg+znO/XrsZoACXJksSrsDf4Ot5WCyPnM
HM1kAHgvMGCLtVH0b+wLyrT+6dHwpHCRUC6DaTlI4/JMjjQQygYphgK1Kv/lnxlM
vO4RO+0DkB8f3jrDDUJoorDpEHPi2IWkrzL40MY/qJ7ptnhMR6SQk1tApxFGXbhQ
cVnz6IUv5tjU4d4f0lZzB4iP9m7jyJYb0fkUIHbTNZDUgWIrRDkz1X+I3+yYHV50
xrcnYp/psGe34iONjptAwPzgSj0z8jpA3MJB0z29r0LrlIR4cA/5OBiqoaSYyFyq
6wXlf+5LQEFneaeNUt6OgNogorbMyWuZkmflvEfjWLQ7JB2GNGm+NbqpdHVJjg8v
qOyaGzHP3XpKct8Wnq6IhsbJjCJMCgW8PVaf0JhedRc5qFVkgozneDOxDaagtYeP
oQEsi+fYpnCMv3l80JNAd0Uji59P4JMoDb9kDDiC7SVUHRefbqlQy2ChZzRmm1Em
iNs1faqHqrSEr9gUb3+BvlWtUHDv6pO6znmEn1VlO8Y/e6q+Oac0GXqO3Jt1sidF
ftIv+2CxP0dTlURCXrkxOU+Mt5aN/Jq5MfVPu2LJCaDVOOKIAhj9CslxPCGWdCXd
uMpe0nw08sy8VHpnZil5ak9ITlS2iOs78QuCK0rmkLVGN6KDYGJ9VOWiEppN9TnM
p3ZRr99AvrDWKYGYxr5Z5fjn2hy58kaQ7VmuxxOQq1sgke6TnYb8VXfnPk3zlgxt
nu1Or4GiVh5TSVf72IOkKi7lqf9+22nBW2hWZRxjgFRAfj3pFU7oIUawaGtDdFLH
rPWx1UeFJvKGaufoDPDtRnA6AMCfYr8IMgD6DT6+InHsAbhmOtnfekXyeJS5eT+8
x2xP4Uj3EIjNvUk2V9pUglxihN0cn7ssM28V9UQDtE8uVzLI/DtqyXfS+qYphIyX
Mw7JW99F14hkeywmnhXSBegK5HYN2qFIEew9dbpGmgasCthxGjsss3LH63FewuPp
eivBTpohOonZn5puObbsVzwJqqmNV6b66mTeZMYUWC3pm2x8fb7pXP8ChXJgLzMr
Jj48JUla40+Cf3jUXmUmrfBAouQdoQsBmYGYChV3se1WLP1svOYECm6NG3aMPMob
C/yzH9G23F9354IMdyfxD0k9AvBQ2BziUu/pA9lNxREpyuHKkI9b9OPsm4tM31q+
et3MvIyhauewJ3YK/GN7rDI0u2q52Ryu7gxbGVRuVbpVTR/4Vyi5X6VPWwGGdXAL
JeWnR5o+12cKWdsM/R9txc36A8faej16iX9Qq5VCZRyw333OrGT5CtbAjJ3EUKh3
ofPO0iPV89ETuPR+bluTeHrWr0fmQDc35u2iR1/k/ZPqCUWnfncIq9lIRz7L7nzW
J42+K/+OnJII+nMTMRsO1mCL9zpvHZmX18JSdlV34YVEg3ywULOy4r0HJR968PfP
c2J7PQyNHjIFImJEGxOOiMOkHFwzjk8u5xJTzLb+e9SQw3LX+5SEtPP9+BdWKFXD
rK7/sRmKKXUqgbw/cA01nodOG9BjH9jN9QvauUCtjSeP48AoIZY3TxYOONaUmv3q
IrsqVOSHF3iQ59OAdoRvE5eFP92nwM53criRNZCBRDzGqS0hgqVnqXlOfUeHt7p1
f0AP+bW5OAQTZi2W9IiKysb9JnTJQrp8nIHtz+f0qpBuCJKS/y6k5luoRr4S12Yk
0HkLnxvCiB0rrkf2We6u74sfHCqoq51oFHuxJH19dgEu7dERMYUMBFFZBglJiZjU
8Q2ggN+BD4SFnLkBZ4Tgpx0E6pd1i9tdTAeNiShnz2fORJffqeH2zsXfUyERg7l6
h7nC8SHbkRLuF5WTpXgVJk21WgTEb1BYm94kgPANE1b9V344dm7mnmtdQG7iDGqX
e35S3d5mQwF/b2v3suQrMV+LCkhnKlNjn+4HI+h98tVg3TcH3fnsCYytYXaUq43w
MQorZ05XCA9+C9EOdSgaBq39XvVJKy04qeWuSgQFuZMbM8jjNWjUFRBQbD6PGMr0
t5tM7+wjRMI4kmrFJRVdrRv7BcyncuNP19hNFcrjjN4nlgn5N1fuoL+c80/DDPD1
CheSSEINaf/B2zgTmDhkVHbMBOW5femJCMqc9MMpDJ1YpqAeHsgF7tP6O5BO2LWG
LRjhx/ACCCtVlekEIFz7Xi1KowJ5112fJiNBGaKiI6OJozBeWJThoRcKMGqFU9KY
gFotQ6tTEEnCBwOLZtgxvcjYRSEq7vwa4n/b6csMYDtwdM0VMTWXQIeBrCrT5X+J
/9l66M+tAjzd4AKPoz63RljvHLOa9bY/SdQNRbnG0KLc5SF58m3fsb2CAQGlGSah
vDf5RF8JKz6yCGX2BF7XFKjr9QBBMV68iNAkek0hsawBcX97amlTCnOYqZBbvcyr
Y3Z9qCvCDJIEDpJVU26IJqkxxYQSAPEsEItwa8J1ZnVDRMIHE0+Tq/xV6Qvik9EQ
CUKC8VAS1qVkJxgjIog7AFLCPaw/SlBvOBjdnuW+M9yAGhdZ2F+Gqe3g45x68ZwU
tDBgvSdYgnfDstSTGOXPMtX4gVNUGoY8RNmV+9zbjJ/KJtl28ZL1myGaACNKxiSf
2vojmgoBpMN8oGxIE0Id7hsU0HmrZz/atWnMhc/YIyvMWPLSjuUCIZqREB7NTc4B
/y7t+3BCWL264fCWVFBl5WGkVK3l4MH7Kh52JpXk7kA0VHnN91ea7/mxVlxfgitZ
VlR5W9xdVEsTGnT88YRej3H6F+l6LFy1WctkhxnZTsL/xULVWctYzLA1eBMdMtE+
z+Qbrc3dwk3TfrOHn9NLrmEkW1szbyKOLLsYKsb7k5KENv5+RFdVyQdB17ra31TX
SwN4qKOwbrTLtWJQW7/RDXV82Z8yXiubq4GOqNR4gGVx08C9kd6KPFRMCXc1RmsA
n0dKyalHUXPaWXnT06H73pA5B2dkK0citiKUcS6/c3gTCAEKWFP6pCdG3wBBFFZ+
9zzbHgLHB5OEWqu240hHSdyWYi1RLgNY6ZyrwSq6QEbXz62j/VRptldhKYNvfNdG
w9cIxRilqTVQbTEQbTYiO2xolBC/DqIfVi7QouMfTqn4eUNUejGWyTF/AiV/dCQP
li49iXKQYU6JGaleE7pGZ/8PzHUwcFxCmKRFDOT1MB7/SdyvcbqHCoGEAtP/nEP3
+NGGa3wufsWtfjdgkU0zCR/1hA4tWlYohcHzXHvlh+EW90oPjluqWWvTODZlsWR8
0w0teVgY/XUMGzewCR9zOArV4b889yVMOxQClx7X/hmfe1viikhKaW3Q9wU4V0BJ
FT9W5m0Ig0JjTEKWqGeFuNT9GEH77nQ5YZyGcIkq87vxD4oifOr2KjES5rVy8/9Q
I2CsgqIFJlD7qtgvMsS2nXZBUXpVIksQTx6BVVz629xAL01+xoGRvFpnPAgK4CWk
4hxXw2V1PvOu0+sOo6LZwl0/NG1YXfsUsRMzaM1lLWAtVg9YWgcB0v2w01v3xpRD
sDssA9MkbxU8ozDbuXfcHL+RQr6LDQbJoE7Vk93Zo2dct5C5EL4cqvyT61A97WMr
UxTbjBXQS/I61WP+T2vr42uigCPH/ngC7AtgxpU7CYhl9YgeDwLuHlayHyMnWGhz
E8TLXxmyTyCbuGB6LAC4gBG4rqDLIE6XMH+VM5Bn7DjIQv/nExGH9e/5wGyMeaYv
+SV8pxC9sMnHWBGYzPEmCrPVlWViLLZTKsPEU8q5UoTCxak1B/8OqMDLiibJO8nj
ME5SaXAvA95UgMCtm1GO2c84YkgUbszmKXURqiGh6pd+kOHoAIhuO3/slX+AXRkD
KSj1b4SGgrcm2VZWJjNcnqrbfrxrStRZriUKD1cppWtKLm0uo6C1OoxEHSom5Uf8
5UDFpy7oWX5pC6e2TeD9atqM1O0/YXGEwa2v7UWngDulAd3ir0WZ4zTq6SqPkxO8
5ckQPfOOiQGTY2FihW5yvIn78vdmCBUlQsRzKCMc1gqMP+FfdQWtdqy3oIdU76c8
E8cQwTCT+qbqyHEt4B5RRjmjHK59yyfDMkOLbN4851Xx1xwj1q6+3FHCypGKQoFv
6gpBrKUVuzz7TWFNNgz+MrONCPpZ19M73mvtO72YRSrfZlOs3oAXJhuYMBIurECh
qDrhozfe15mHQdtk/8tHgzpkDfJ0n1pKnSRKI96rnkRTOGGiT4/f0qa4UoHQEplh
TQ6gBpNG18ECDD+p/nXihqJx2+ei3QIcwBto11buq6orDpZmNOsJkIi7fKN84Lwn
4j/ucHFROlQIz+NzOXGwv29waMAlIWI2KKIYvGwSAlAgiQQNe/73pcVYJ30rWbdG
p7+eevkiAhWXpY1cKW3Fw1QwtW11yCqUSjRE6v9FbaCYWuNWhcA62BHO8TSiSI3E
JDEQyekm+gRExepj4tSzdV1aasB17SeW2EO7lDHI3juqZIUwlkuOsmJHPVvuOaCm
vuwmRmSDIxai2/hS0FzMyOCXus3zi0Oi5HhfdyFvWI4cpRdzlc+GEeGYXoPE4bD4
EGVfO8g8H3OpvWDfkVkqB0p7rSpQauC+xGdYPbfA1coglBmxDacXFUHJBnTIEJjo
zH2GueiseR13BK1V/alaGgGBGZBbw9ncwtTJLu76+6rX/rzsFlHaIn1mK5ELl2Ny
GonjnbUe0W4zAzrpY2lA8oYfgwX3dto4n3Bk45CGSPOIR2uSbhs449Fr7JrqrXv7
NjGbfGGoa73mkqBLi6JT4O3ERQwLHwhw0IkLNUDZjQqDi7s/91SgvA8jsGKrsAm8
79tamPlUrtKP/0qi+udxRlUh1IsxkxVN6fhcfqrlxTByjbQaKxJO1iTNt02ziKPE
cP5ig7YRbJtTbWNdkde7El16ozi5L7sFqslxNPj7MjmkcWGcQkV5hn1tV+2FLgyP
E93eWIoSOxCMf7Bl4G91laOFpFpKBeWbPvCFai61h4jPB1oiYljFOvgc/Vi0GTd8
vPI+whc2W/q5qD5/cxZVwB6iJjreXybLKmiovCUdeu05BYBU1cDaGxWF7zRpBTTw
ctYRcVgJnvnq80fhB/ttC9TUpwFLEmrPHWmi90BpXTxd2oXYy8ophmunWnB4d8OQ
w436KO23FYtwgsEZJo4FyulRXF/yZk6AMNGNF0cmdeHoBde0MfzEbRhjsGpR50Zw
4LOzOQ6tdOiE39gNxqStRvt2RMBLunwsqTa3zwgm/EHcdpB3xZjFmbWNz86OnGm3
79Mz88h7aV+Cgucqo5Qr2v9lhq3zUT/cHdgHeWUtjjD0MMrGy3hcHcb0jPqGj0S9
92oOyqaYhuYO8P4MIv9NKNoBqxVX8KoKjcOpvhtz2gbHlviK2AYIiIZrEkj5LI1w
o1K1+xPhIanm6sCb4mYJMl69nMJOaJcp8hetsTB9V+0hdbRK1qEZliT0k4Ogmn9R
dKB8UVAYCNePeXNmqeq3f3KKTuJsgQWOqECQKTvYp4mw7XdoeXUA7MU6ZKn/plro
s5fxlB1wDddgirluzyuqDzIGHB2Bz8dtBpAD/UcMS9dvS1M/G4KJvKwjtGY/nPJZ
gIA6OdF7RPBih5wxnDcQqHyfMbuoEAA55mSA0x8gxpX+zxcV0asyol206EPSEmUy
JhkaisLoW6n0dNHXDlZWLBU3MjJN7NmJ4BMmKc5+AJCXpuFNiqMS+WgE2EfFlu43
igYhy1RVz5TD9cTpfc3+vYQKH87UbvdjzbVp/0e21TPoKzw/36X/Q2HsKBLZmOt2
za9XfoOGCF4Yfyw1tS2BCieFe27aFNbJ8lrfEZP6XGOjsrbSNF8N91FAPAOGb27m
m4xQdc1tp7qvsyd/RXEVSqGX1z5dFQqmRBGTYL4nSZfRCMow1IUcGif1gEAc6qk2
PhK/Vh/AW+BWpt7p4F7MyxnGolxpsGEXAM5BkZ9HxlaMT/3FK/++1ZyGskEamp+k
arCrrtG6zxkZvdVxZxXJb2Wr8l5Rb4GXZgOnqBevWpuKHRaT5l1ACGfHMBTuPXo8
+VK/Dnxb8HCKx6jmhe6bvqHZPKnA3nC/uvdTs8vI7EsDaacNyehZ439JwJ3NdPo/
DUaWFsXnLad4RUGVdbJ1UcfiAkJpiqG4bx+v61XolMEED3kS9uwOhRCpaWUECpzk
W6p9njP4/ZMD4+CFZfX3QciEWWxzK0294jxgCP0Yrua4MZro4YtHTx9fjWfj+b1R
bQTpLq4x5v9UvbRHRPfA2apUj83wL7ls4IKUIF7KLLFbi4OjfaXeXrdBzRlFJ2dk
ZWpUx9vv4gdmiDKOhXJFSKOxuNnFioOHtHmIDCTt2HIQHhxfsH71BLViE0tSVIdX
OqEep+SNHNEzoO260l1m3s5uNfLhRG5Dcg8eQuwYUWmR9Q7RsMmunUTQmNdNrD+g
k1LJuv8KhJhTo5m1adyz3bJUfGYSfTMlyIP/2GYGpUDSK7X39iEqhtoElZPv1CBi
7mTsRH7KHaItRMTxIusZ9nQHsXOW8PuUb6tOJQR07XBLftszjI3pT/vx79JTganc
JwgupwF46K6W+erTtrqJLL/CD8vInU0i+zp9veHjjX1HiBB4bxcGryZW8q+pI066
LnCKajkIUOEA5q9tmKZVZSKHaFI9mjzk5DzJZYgT/AaxKeVjaAelm9tm3f2p5ol7
3BiAv30RMv7SxpWlSTl4YLCST7XnJxd2WjZj8lErAN/F8z6Hvxj5TpcIXpj9102B
WGsh4h2B7sO7WKwSJ/hAmNNNK8MFENcmVlpbE8lJTfQgbKKwlSurH5qD1rxGbouL
E/Tnq1nYI6YzTImRqwHzq1WebazT70K5BFtInxrkF9d89t/wupuGDH3KtLY/gazc
Bf9Ehi6NP44JJ8h4dZ9F39/iF8NOjDg5rLQO4ZHxv1Utj2YKjaMttgvIghXwuqOj
PR7hgkD2gjymaMftjNjjXqYHYjq0F7P4NuWxMIxRsMISQZvyYtp0fWWrjQrpXHPC
WCk6l1cjCwb/QBDooHKfaSlKOB6EwiXO6x8Ok43RaiV0+OLtsgxy9p63oJYzqKRG
hjE7/4k/oWR6psLKB/Lrpeej3xCTtlA1PtE3d4OXC/3vMkigy3UdfRSboVydBIZl
fFhrW5Q285MV0unNRCJi939iSVNgk9/HEGjvsRcR4TRZWnPA+7b42IbxAU59Hih2
OnRbvfQCQB0w0s/j/v5txE2o6LcqYLu/352y9+oJi+dMwquYY6u7+oSDK80ANwBS
6kvBSkz86EOH9cra/qY4Qge+AoZp4QaEroN6xwKiYNKzFpgHhtt8NHOf0Wqtk8uX
u6e9jQ2imb07SAqjXCGu7174XG2k6gCbY9FqZJ2qAOOKmJBHIl7It5F+vY+OOE4A
G/OySpDpBHYImVgBpudNyRKPFUYbP76SAxH3KXMVvcmwLXSOZOccJi5xghd+gVXU
vDZ3zS6JZWissludsA9LvV7lDz4h8BDZoyvoDy+34bLOQcgY6n25/48QP62u6VzC
EW7H5OPeVjpqWvhqZHYPzy4y/XITwmhj4R2SE4zIFm5b7urqaTKexBhW4TuHiK+o
z/mvFyWCNV01VPobp9b+f0TfGcV5dcdmQedUUiihocYqRbX2ycLIq7ggh8yy/Js8
GL50EtwaTT2YC/IWYD6yenwLa60pmvuN0bUhghW5OJpaU53VZ4hlXvBahKVZAtbg
mn8X0duoDX4C8kLoEpHdKiPcYKEEv2cxdEBakAK9chvhaO3tyAytIguWVvRX3/0k
hLXTo9Q9vo98EsjLc6ElovHBpYGBIJ4rQa+1mkLXCXdL4LpaUhtT0WSARBuBcvVv
6R2uBy7VmTu7gM+bcyeY151XHm/bpiQPRFzTzWMoARM9I8xKALZplFLhX9gzODKh
4DE1DEIMH5qEmKlLKIhDd3AprMmyA28MAtWZrBT9Utty5zUnDoaTo2L11bXK6HKG
pJhTD0k1cB2ADT2WsZfi0bfgxHb7C+v4qUYxDLabUjRQT9XJy+deQ02kzrMsgFvq
JsEh9fLnzbhjyvO75zLRHQxMAHV3ffSu+hKnrq4BFn1xgdTgHOoHBqe8Su5JsU0m
Cw/nOk57mwEUHzjs8vC9NOHJvJjPd+Vb64M/HFxF3f8UdK7PeUpc5KYygWCqrxn9
Y852Daj1Io9UOVoPk11Kfg3HHnCdS53i2qvj/7G8HuW1CpjFX9qwwagaFklDLdbj
mxilFWDNQ7rFRkmJ5yZ4kQWIlidkiCbBlh3SeMan6KGlWu1mTr6ZTQ94z+wL9y6n
cVBy2hQgpoDyEdtUZNK+O1h9QTiaPDSwFAyPEx7yt/zZEAggMp2/fP1rJbkfjbiX
+aKyX/VSFnSIGyfnqNMwGOwzZXcLaYNlhFQNjYf/0HnNCnDEAT2rNv2iDrY+iUzn
zqGy107UazonAEw3XFYB85mKYNr0MFEQaOu65NpGM9mz8n+mgHiHS6HxsNsD/FP8
o7wb1en/+n+NgHwlVEr2r58c2bCM2v2PbKubnSRs7SoLG6TOcK0wI5Z8BGyBTaH4
lJjhoLmbpbqJNlUTgntlN4LKdw1Hv6j7TVH6mAKbTgTuN8p8IK6SODtkY7s7mdfh
XBqfPIkwv1LG0mEs3Qzh/qlukOmtF1UuCwP1jpVNQYQdUtsaMpX/gYaZ31SjKDAZ
nf01JoE0IiYyojcJXTy77WI9wihHHcrRtt6AUWVYyHpoB8Qhx84RGHexPFLoQf67
h9rFeVU8Xss4PsGyJhontAlqC9E2l5cbSPpRLoFGYYSmP6rwH+jHRCxTRh2ueqtg
efFRudhFTFxAQruAZ00C6QIJMYYQa4tL+lPgsKSgFrRFxJ4ZLImbw87hO/WJQlQ+
cfAXn61xuviBHZ0j9e7GibKYFqABgMxM6sGmS/JMyDBspVNv51RW+YwZAiDnEOaz
66U05JGIOzZJxgVZtQQWy+6QSHZmUf1dFE45Ay1oe5iItj+YZOxnVMgSGDuxmkcE
kRMG77LIK1KQBmnfsUzjmUVj1te7ABWVas+v80VnKBw42Bh8Zv1IvW+QLqTyfmov
/1+oNRcqn8JqvMcJM48OumbsJqdq0NVYfvXF6Vv7qR66JrENO6HTe4QmzCRAOTfr
BE4fSuAsYRYYFL1OeQ9R0kdm2f/+LDwhwufcAAVj8aYvHj4t/uUd2zkKXFEKNNJn
INzo2f3SenCgVBjtuqo2XE6qYdwz+/ueebEo4vteXyRoKY1lImi239t8Krf/RuJS
f5cyXC543tewWrY5n+cXVSUigorNhaGOG8Y9tu70M/WVmnokItMjs/IbLITTf39r
/1Iw3VbrbJgvDZnil6RbUqr4Jyg2bkRefmGBjbv2ZXKCWGhCDxHA5A3ulMuyEObg
frl1+ZwCuNM/6+PXtWptrOUP6YOkqdXMCE0XaLzMW8OI6WeUEcdPV15CERS1yYfo
27IddSahYct3DcaG3LaRFa7WLBjHXVtpxtwbTj1K0gl52BUvVXFSe9W01LhadgwO
gvC+RTQw60c5F9zKv/9SBq7MkmiUEieY75Rls+fd/GE4D5CggCN9yVRpM4CHL9tL
zHx9cy6UHM2/b6PHh/wmw7sj3kanMcR9ydpOhpyeGHmMYJpAK8rhgUPyoagcyVws
ju6CNr+5T1nAOcOrzJgVcYnHyaFFThdLAM6At8JMQ28X1msiJcXZ2TH0UHFZGZBx
WLh6yLYs+TzfyF8XXo6LZJaycL1386FM2ZDbtOHto0jJ4/tvyiGCJUbM723YCXRx
fErfU/hYTk5dPOlOlae11yTPaP9DWIwU/OHAoupskGKMTY+B++Rqejmne7sktD7c
8yJfNx055coP73chcJejxq6WrDnHFuvgXyET5D/dkMasFoB9x9f70lZm1Upi2PQr
BFwg+VuEdr/wJntWVBApfmrHYZBWT9aLKTE/Gly1pSczYiNrhUqkLZJjyvmCT7Tp
YQL3RC03eBfWant3cKJHCUKC81Y26hRe+EL+19q3f0PrTHj76yzodwiWnXdCHmJR
nbQmp2VIxrMOUB+q2kZFyEYcKewGXifiKCGP2tFwRBMYO3sZItH/6bsUfS02kBvu
MlN/ewGASkXPy1+mzI3JUWYZy3t84bPQXxaamRw2cMQ7UF7VtZHKya6pFqdcGmQY
jLne1TSjH+9pmPM9TdBI8qPq9EALpfXD6cJaiIpFjOi1GGwkrlh1MEzB62uZXHxi
qjE0Ky3cXBw1Hxft1mV3n4+v0hagyaPARp22py98FSC1HZIjfFoL0AFkDMTX27xx
4Sp/OVoys/+fki13mkJxYFnr+bVfHnudhtfmmdo65uYmvrIgqL/7f9iYCfrWQiDd
n2RPT0MccBx3vPYdleQOPMq7GR6phEcSSziOK88+iKxPJnrQvHSz5PSKh37YwJuQ
FWcf1B1u75rPqN6wzVUL4uivSDtCpRSF4iJvZ4OtCWFCiF/R/RVn5M6HzjZuS4ih
Mr+o9Va6ZoWFFLnzIxMrnoHKZ32qR+m/5hqK9fsmJ/QXQ6MwP8JXbIGzmR3LqorX
Yk9LZJaBLk5jUinPHww7QsErP8ydr6m1lvzhM3vCeaGqChPcQtJW7qSYFeRikoyp
SOlDH8f8Jm342RKTq4d1xt8HFupYVsgjK+TEuV8tL3QxNFWrTgtMKVk7gGAjl5Z/
0rASscwVqUzpm57Q9OoGp6nLZ5cIfp7iS+6WKu4QQh28BcWSGrU9Sh4Ztniwmhvh
9WWufD5NsbcA1P1e1uCiXvgy/Sgo50jad8ptmMxsccv3a0RX5koLwHXMiOfIKn6L
Ludr6ElQs85E2if7nR1nfLqVuJjHrpzZbXWtSzd38nLyRRPJ/XkyLReSRlJVY4kJ
TnEGeF3JjWzKMNtvISwB2CSn8uJbxa3GnqzD6HKldCZxJdaa8+4e0gGhMF+OL3eF
6XUqbnlgLNdSa+VjcJ42bycO8rTzgXo0llCYPVTu1OBZirq4OmJcWSGlKWpt1ZoU
6XU2g3VikP4uca+YohpOC/ae30HQogRTdAQZI8iA4xm6aze+a4EkxZi8IuHYWpHh
lTVYd+jSptyoTq4gA2THUxMuGadGRX+tVppBBEfSclLv50PjAgZwSjv3v01PzjR3
uUGVu6mQYoTgBbuDln7wPBuzzpHSnDVOvHc5oah4B6fe12YSuCgUq/wf+tEzMrCT
8kBu5s2pQM0B9E4tgGF4Xf3+UVaVc183T69Yonx19J6GDxIEk/zKqw+rn1swKT4p
G5qp/kWrErsCOryR53LoO6Yu3EQSAVGcoLfFg/Ay+drn0yUUeT1oQE+Ect4P5asU
0HvR/fcktObO7+lDNYUQ7PETaof8DlYahRpU5Ict1x/mzbv4TgHtqqFNMD/Z+CIz
dMSGawByvmRzAo6lM8qCIRh5IoHDgl/UvJDWE6bP/5l+tyAtFWlj9f+B1FzpCMSK
KOGt8si95/FhYdJfmEvNwOCUB9cTVd3J2yj7Wku4Ff5C5ayW1z+4tTkHmymf1CbF
xIcV5lJE9ghBWBILoo6bTWSApTc8AndjRrddUhHL/H1LKf1uSQd6IdQRnD7U+0AT
+WOJS8ng51Bxap2hH8fxciC0fOQ/d062No97lPh6FAIkbjkpaMyGIybDJLwRTEOm
yPHw22zBre4HxC2SkK2OxNID/Bgr82RQ1Y2NNsrh/I0TRAFdP3iqnKBoL0SgjBrs
crG+yTuimh2q2xMv+WuruBIJ/baCAdchHdj03AOfpTQPsbjfQ9yZozmfXrSprAUi
BH/cUB0e4l//C4mc8X1YV8SiyNORBbzQ6yOpe4MvfUuwiHqo+w1VDZcKtsaU45Vm
JnWWW7hrxtoSZ2rJQL+fR0O2I32lnJZQXEsQyKwJhBcdZlS5xdNktsQhy6++mqA1
5nuQjFpFHpAuVq/jz8CpRdZx6UvXx9lrjtVOGF6Kc2ZAo1GyNePcIkl7DSXa4JZH
LzFNI7Uz1smilcnqYAEpCkb7+OID+jbS65psfk4FClFPq0/yPv2JwBlUG49Y8AVR
sthgj13TAr3Xy6p0GRh5q++A74r+ndowCgGkPQ72E8PjtlepYUGeoQlih9dI1ZPe
0/c7HIHJZxFAsHJygisLE1g7lWZCmSY7JEB+12gnjQRfiXTJ1fTMf3c+LJ4FyIlN
STeF2R8DAAThNmKOEnGEkoDnvte6qfmTMEPeb3MEEtKTNLLzshnQj6VZINvtRopc
o69PQSrWf5SGcZG47QlfjVIiXCYccy3aN9nQUGlCVq8gLfkb4Y5NulzjrFE8dmOC
6hYWLQdeTty5zxygS+5jCVXBJMP/swZKkgA8tQHHLdlj+wdViTPZ7f12OW3WSt4+
y5HSQm6w7cLia91ICeQvoA1DrvlTPr1lyGHd/2rhNPw2M71k9FIEgdJHOyZF4myn
6f9j6z+2NWh9SNxqqFo/HLERQ14Z6lF0MZ+thj38CIwFNCeDKo61hFV1+TOfYgQw
FUfXvgESfEKro1+4liqeQ6zoh8Z3+VpetcaPsZJ3h936IgLOS4isgic9/OV5hStX
+vZEnbAFf9uXCKquN67yvlJvMd44Middld1gO9aHHoetw7HjQc6B77L/zVIjcxHi
l/lTXIMn9Lc/bGLQ4s9TbLAiKRfEEa6Ld3VSrnFH7sULZlvndBwimCeM3bQccflI
hVSkJChmy52iwHRrYrv1tj6sATmJJ7sHHtsl3OQ1Z8YEt1fxH0K1XCtuhILckZ34
DGSfIFnv9T21ESMiB0HKf6XLzsh3z8DYEs2fSui755mU5koPTy6wb2UrSQ+WUqSl
XJPJ4EGIG8Qapxz9roUlt59k8qywvxrgFgHRxyxq0ADK/lD6tfE7dB9qZT3iiemM
RdZdBEgrVu/1Pz2ltcmbeL3kJ/4h1udXG1Du9oLlsAC82gDNNpCoTme6eJVXq4gx
c9yE2GLIus9yzDdhT9pn7y7yPimH8KBuZUKZpKHmeWbG7To2dnpKNtZw9EyXhbJu
RS2ejbsiHOkrIIy/PXnbAgg0bWtc9QFkJjDR2XbTmmTfvtZHSMhxXFYTN6z4Urie
M9wsYXCYKZ+sgASIORdqTjuIa4t4sYDaQRS+lp6eBglhUb0AImdZ3gTeDDqOL7Uf
ug0WnU41toqGnRGO8Yh9hSmrPBtON/AXfXVGpdcdRpe0i1OMSUzZB8Gzwtl7Rq1A
RyA+RCcyQpUoLmmwB5kzYciKLa6NQd8X5TSg6hlZDvoDHTHFceuKVg9OvpvPCa7c
UTqtaSJKoYr7pba6tVwcg+scXu4j5m0pDzXP3PghM0+vHZYTQPueB6vIF23basLy
My3C5ZJIAbNpWQOppkRKUGRUBeMYQLS3hdYHaNJoB9XBjmqsM5LwYhF1f1mnKnOE
P0ZQTaWtxeg08FUx6v/BUtfnzOcz5eX/UNVpy/M4IYcfU683uKM6KEMi5pl9K/Gu
ObjpDw0dzkiEcrIr1Bt/z+OHxoKsH13Z34Rhq59fc82UPPCjW5cwU4ewlg9Rmuwf
Bb/jLzS2E9ZsAJFFZkZ7ae/Qe4ZH0SmVSvxnA1OW3vjTkBcFXdfn4xl/xM/0b33B
UYuU/+IcWIvv2f0NJK79bGCS96h8o0dh50sY0Uok4xyjeN2svvJ6/1HGPXeasZrf
sJ1RqNyecZvlTJxdjzyEs2l19RU+/pUmj34BHLktWcPb9OAk3nlZzuBpO1w2tz+k
v92oxYwiz+QJszCfElNacz4wmlODllEpWPn7DXsLGs95XHubMwnQw7+0hiXO8sF2
ZuJa78pABKSTrnj9dyghvx+aJLQ7twiyGPzA53qgdCRvxlh4BHuBMvVCbx99bZc+
veihtijAgk2uXPIMa8IucB0ETQZPuhN1YT8hGVLwMZUeWgpgZCg1KPo/wt5D5GJz
Th48JXv5oatPx+zemhQES468+neVR+T2KZGqH+HbszAf/SEWewo5oLPeCvOIAZ/6
K0f4Omy5hVeELsWJ+xF+Sm1D2IqhmM7aXe+7sXCEdMqT9aQv9aPoTzjcCEqNpWh1
GgEmISJ3mlwJOTrnQsSvki0plF7x3/IeHboF3RmspIqJY/AvPXjd+ykxNXdaiJix
MGTefwpDnoYsF0S/4ZW7ZwYbuXIa6vZzvjKk4vtkIqqq0W6IE1y8wbcbc/YpqYus
rLLNAOeOqUwzk1V62Bo8b9qRJvo4HaVyocvP4oqQUl9Q7hvha4o87ttIqicwKoBg
FHqzVPSCGdZ2oq3R8Wf7NpQn40YUeIfSzOzJmaGA2/uXsMCp3tmfL2rXJL4qe6i1
gG83gRvvD7euuqjemsVyeoRpx9pQCZakUufhN/9sW9loy/KC86GAmn2PaHxkVTl0
286x6lOcUogi5DC0cWCOqTvvlBbvwYnaXfgVGMKqKhj7WfbKY12XsA3yXmMTEoCv
hjuiiURicRtCZ6kCMpddemgQsO5G+BIsm5R5h9TGjhm+UgbUucwSDeLFdd41F/hm
66Mopd49Zyi5hRRVRvZpkcv9Ca2AAju2W9XLY6pN0+hXay2e/t16sDcRymode3P/
drj4qoCZUhacl7XsaI3xmmDeNCIGU0OPtFeQFp4cG771AyFDe/bfNhVzcs52KnRY
zpVNZihv+Eni/sfHfgpAaOAs+axGSiANpV5JRVv70Brb1wjOHV4xI2VtxyZaTxhY
EfIczvT3dUfMSAE0vWScI79YmNpCFaBlL4NClFse7MmEE31N053SGFqhUbyjbF47
yykOTikNAVLwFYYtqa38uLBSX1gdRMMZhmXe+y5t2lLgtaNu3xeKIHYnSYY6+2RR
oE373amsZHE45Olf7aXoxGrW44Jtxyef8bBtmBndFsMZdohQMy4ohX8EBS5u/uee
yb0TMr7J/goygzIiCsJK5lT1wB8ep/Ke1RYEl4GPwm/nPk8tGXgPkJlDHFH1kOdX
b6KWS1EyYyVQXB7xooqONFlqZxGokUXr6hoOoyKf7Hdw/zf85hEddNRV6Rxqa6Kr
mm0yQSG71wE7JYGaSqI0GyG/2Po+q7TGZALP3W6qgcqXwKr3F7a2YuKq9s25Rf/H
TZHHkBQcOmkX7hNvLXWsM6ne3N9qsZXF2L/aK6WQ4DzwZxkVYpPBbULNNVgNLE6l
3TADyPt0YZRTSmdrFm5p1ac0dz0aMilW6QTOQrY1QU2QttsKMcdpNBhA/XPuvHun
c8/dhxD6uvic6x6ZQUNMGMyvCKWF1uS697qv62AeYIPgDON4VxDtnlD/GGqfwUCY
6WGXhiJojDmACOJf75pllqre3OQtDyKLyJO78Ld5lTH7LGXcoobZv6Zee4Cjihab
NJ2lSc6BcDZwqRq9UKMN7QvCltnHBpp9nfmaq9D8t0KlIDfTbJ053vqzRrqjM/LG
iJ9KrIy9xNKsHRIWqC3GA/1wIeWew2n+AZTcYG9efH+zICobyVPRDBBnGCKJ84gn
F/wTotC5DRqioYBPaSJcDRxnxhXKfIl4DqtOrZSK9VeuQZ67hPqaXLmOFDqUisEg
S5NKbdzPew5IiB632QnwJRJ1tUADXteF2XL1DwIvd7/nNoEPAEEL5jdlTW5yVu7d
pQGJMXIwmPOdY+ii8/WAI8Jy/2e0uu5QwLzSdF5pUALxJ16y6zpLNg3I+m2CbqhA
HTR6ZPUddpkBOSWdN6bUBsLGomrXNrsLaCDpCfZGfdOuDM3LStZDX6+npsrwg7Lu
sfNuBFJoVnCW95xMmdObppkXisIEB3Z9Q+cxCKQkYgutmdpUSs6v8R55ahFv6MHs
2sGMGud29ZoFxVFvLhDtbfkXkF24oAgzyYF0L2nLGfvuaWpW5VvPb7ZzEKa+0Yri
NQEJModkeSwFbcYEFbs7EzU1tp/pORg09iOBDeqD29aXAvx9YOzKcmSaJd0C9K4/
qaN1JmpX4Znhbde4aXjDaLSDiKmzqLydOXP4fF0moTrfQxaIIuQLXCLsah4uNhSO
u00VByUHbLPqB1fEpWksNUar7ukc41+4ChXMt7ABaW3lNjFUFH2ywCjH+EiDheye
qZJ62KoDUExLZDPOsWclf8utTAHATWIWg1RqZ28bosXz4+qjiBbASH2my6s3oqiv
kheG+vXQn3e6o/JWDIcz8rlYztK12ZGXKwAZKG6R6PvNwNj5M55tjJzWRNqc22Q6
4XIN29Pawv+Xp5CPmh1g/WuftVeD8p6YfYq627TxPShLEwo5aupY8GtXgFyUEFnp
W8iTiMRCQLSrYPG41vEjGzAsZLPA/GA6tRLZ6Z+euPopng23y1qkPwJZuPOReVCb
Ty/hEfed0krhJAlb12Eay0w7n3Tpx1Vz4mALaPSvXcFj3nHGdep2ooB04OfdcTlu
mkAaeR9r8zUpeR+yC4XkWu0SMDfyl1mrsGMxCOjbmc6VsMCW1y2qaKJrl02Z6WZT
k2wUxA50VIqmyi3En6AevYMgjWXRQhdOiZXgUYPhe27qJeoQ6brwQtQepGiUUHsF
9BPJradOTdhgG9nXDOpK331IF1zLAcsTLhvBoe7wRljaR1lzur7OMv+CinBq5Os7
o8SLxnqqPTzzC/qz+Vd30+bUJgyZVcqOvA5puvypENNYOAonNkGm7BmZGfHywi6s
lokKhGxrhVPcf/H8OYHVmQTMtRXNr+u3trGNnfUe/Ir0c1rk5V8yLOfeDfUVTrYR
ttCVvtnjBHPe0AwJ2kSUN2Hz+KeTH+Xn8LC+2HHJLl857hw+VvqnDlBwfMkHpXIC
JJjkMsNwFs4l7ztrRm4ySirxYqpPT7vM5X3SNRWu/syZNX5DX/mOgA0hj6iwfPRo
G3QT93yWpf3X3wicBKglykTyhmkFDB3bWZJlml8G+bsm1eR8W2JfGc119VrtF5de
JuqJPPj2tTdEveMiS29jjk6eh5SWtC8EvSYXP9Nud/gSUIqRMq31tCO2eE4uo+cB
Pa9DKsuQ9POlaUdsV6CaNIOpDKL4Pv+hc/GJG1XfUnZzvZsSYwag2HLknv+hRSvO
ap/iA7IyFF9QyOS3tP0pH6g6lis+qu/ak4kFVfSgCV2glLoEJvUoT9BQtZoPmcbM
Njh/pmtNCCEvrklZLAlU57r8ARjCS2JDjjv+EuJjGQwsHWr/gvwKz/YfC+rrswpO
OiTwV9ZERm5JqZ/Gr6/3isQGPHGx57HqPXdJ86X7OR604pRgIXg4b6D8X9wem1Xo
UMajd98CAiEZqRvOT2vQBmetK7Sz0sRc1XFjnSF5SCmmbU8PQvVUF53Newy0OizO
52suQwmFfAyrv6WZFanNy8msC8CCqeDJrRJLEG9qqfm+++lqfgaZbg+ZO8w/+x1P
2NSOQhXN6n99e5p92EfxIYt5iB8eu5Xk4dSSHgh0cjoX7vDBxNJ1jO0POnShoqTr
Dzf21ihqn9mhaCVoiWWBrd7eE0BB67un4wziWjtuX8MEyihd12iAcYgbhZegYsLM
VoFwxP+HVaSnOmP16WUicNvMFahV/EiIIEpo6YTg8mOTi9KVEaUGyP2zJ7GkOm5w
ZL02zrc9Oh+D9xDMO5ntTtRC97X6hX19r8pBQf2AJT8fkM3bykn/9dXGlzk9RPUw
1WPqm0WhuOo9ocdi1Z95Y2BnWZp4sUK4+hDaA8hJiL7ZX9EY9km20g5G0Ne+yWv3
n197js65piAqXgX1z2t9T0cNISQK16HYSlOoiyMmLXdoTf7iWDB7WjgLLZH2AysP
1iWztJfODGwjKka6s7Cb4y01MrXQylAZaIJy9dQBc1OantXrri1AG44il6vSdgfN
O438ylQbVcdDN36aU3Jvrm9Vaed8gpQ/uFxgpzRSNEzXr73ccCVwr2vV/5D9JMGl
8VxYJN47wVPistVH2dTJ30t14IkKRf7BKpg0nOiceU7PrtpzBvZ66kkUbjMGy6Kf
FNuK1tMLpLDApkaBDDuNvlN5G0C4lbMMQ4QbgMkkVnLh79YP9UdDF0HoiGKHYtmE
sWqYJCF02Tm+rmBC4mmiwVhC/X/SR4YhnEvfbB86C0hBR/hOhE1l9FGjgoX9hYiu
a5BxTx6Px/D1MO5IM7NxfbLEjcAtBuscs6K4qoAgHdPTbu/NgzCVPK3ZMtzx3RyR
t519svSOv6HpQEx1BHKMVtO1cWbDZn20qkSGbcWscOwBQRdBre/2AskJCz8dRA37
zlvWI0t3CE3x4kxjg5Rozg1MNLuFYnYARObs7CVpRLPhBaiFfbhryyS3UNJ7iUoS
n4m/ViSxiiGve+8IR1Mx2NXGl0fjrVu4Vg81wDjTQC6Q097j77fCC8OB6rPW/c1O
shJkjeT5sbI3asVJi6er+ro7isUv4JkI7SKPiHQZ7ketQZ93k/Q33IaSbviMw9Uf
Y+0F+YHN4kJi4QDZ2XCTHxqOVK37OCCON4c2Hxd/ZsFiy4fers9g3+PPRNeeKpRG
ehMkqE7UZPUsIKTwuoY3lIn900rpWQKOyCyq5tK/dFIpq3aUG/hCYpM2X9WKU++I
O+AomQz5IhXBb5ySwbNOYNQ9oYUgcmxXSbRfhDlLhF6SR5WQEDKoHw+ppn9XcPzi
kdMp27lMlEX6APdiR4fQMtssgR7HTtPCI6NfrgNm32kH8STO8WuV1VxBrvPAztWL
LwTHhzfF2qDOSzYNND8t9ukHB3pm5z+p81p39sdfxWik9reCgcQB88+FTrpOe4WH
iYWfRY6sJuGye9YKHN/XaFa2k7s2abv+wiOgIT4atXf2xHvL4g2ecOoa+pTMDsiA
LVj48Vt5V61jvTK2s21pdZTGa2ntP3BlBrEZLhwv4NpdLWGgZ/8nqSDqNyCObVR9
nFMR+U5N7k9zi6gYyI5baZEvzyz3jPPPl8HdnfA3PTKsWBDb7HO52S9f5VMDN0Ro
hzEI/uzRTTedsxG7htuGQsEavOr2IEiosQAb9lYcromfK3F6tu3AgYow3TZbb8Gy
30ZWQva4BjtMZtvAwKFoe8vVRHMDfmcwliNKGtmI7dB1hrYBu7O6VH2SY1rvneRx
O5QQ1hPn5fkZHhrzIMtnlGXbFvkGKRxV8y4H+JKPYw9QYVdWhN63HAXYtnZd97tJ
aEqOavT2Qb7+Vg1wwuaJ6ggI98ktdz/cw0hNVGPRx8n1WSJxJxtNY59TATEceOfT
zVcph+AQNOEpPS+oczXiZ/tC4APRO1NcQG+lDpivtoZ1dJJZcNYT/KU07tTdZcPb
LtERIkczpBLOo2iRHlKCkbrGgQgNOhDaGZN/VGlXyD2jPzuMFY/cTDrOLXdGGPAp
DgvZmQaQ+NDoNg77e29J4XMGnTXU04Okt7/TM0FHha0+BdEw1frT/iPEwM1ua8Ks
zrWexZqYMZF1qbCDlGqdUE/AD+v5fLLfLAjl8E55gllgv635siy6gJvbLKz+KUGC
wZhJkoPWiMqCz1K7U2Rj6rqy9Ea1wk+5w0GCBl6v7anonZNIQ4mQliQ1fPGaejB+
Ih8wcmrwU/MRfd4j9HAVM3K11jlJE88kcKUt2WCGm/rBx0WAuvLHoZpz4s6aB6Lw
St7VLGIOAYXGjKHTxc3ujFWGlQ7qSdcpWYw+pfK45wnHY8P28TkHJWejVr0+cVDD
ximrmK+t6Km+LumZ+AxgOFiVdrs4z4aVrCUIQeLAxkgSDTxgxQzRa6Bqr3+XH25Y
vUklT0lkTbTkfuj0a392xZqooBSVOgXKbtAkzFck8Da75iwGEWrNtRlkByJm6Z8p
1q2ySachwqpcSq0OvEFdtVZI/Iy4UR2sf1A8fmxkmEUJhXHbzW2xtqdFO97sLeMg
rucOOcEFdQvNuk2B6ZIKvk/Zs69ngJZ0D1pKPYZfWg4TJRzlBDlPqqpXybcbnt8l
CN6rnL3+N5bsVIyPT5KiDnsY9quC5GWBGPg2ei0/tSaXPMPdsyN2o5S/HiRWDBRa
Lv1gvMrqU6e+8miBU4rYR0t2qG6yRnGglLaTqnJU8T38VYcDk7GXij1GYmkHA+08
NAhfCtD2J/uc7QVpWeyDjCw0tl1iK+0DiJ6RSXyQk2+dWerIbopUl5gPKUCgSpDb
w+eg9x2ij0kxHh4X+4TpqnrObHwQ3aPbW1pzqIVGFnWgaRo0+QNxlmq6C+q0+xM7
nFTIEhrKieL+JOhv9zfM7yP2howNmf1TCNxkKnOVtZY3UYZGSsRmm5tnbLqb/tqG
7sVfbhhOpwux68kQV7nfR074aLFdjAWB571+U8uoWNYpSySEtxn32NaG7aW9l0Iw
WjxqYCRGFfIru+CjkesZ39uu2V9i5wYbuhj7kiLeL0m3cGWTU61eWRDIPzGz3kvA
/RjxamyGtWCqHNXCP/Ck0p7WtSRmTn/Q4w5hzfgE8o/Z5Ekz7v86DLee+xBOREbg
jlp6J5dHaUO2H1d77CJjQ6m868lbrgM+lryjaSAbmrVXmkgIQ0RrIvQHHblH37Tm
b3cthd0kycruuDx54wcsdd2cY88HR64fzw7ncazFP08o5kniTsWOGszSMFY6VrG8
7ipbNEtLecQguBeSy+Qb6x9O+uzUC7HREM2irTDbxKnDL4K28YbHUtC3fiYCTCcR
u/1na8QWB6/gJsHUDL3uwT84xrgK78+6oxInE+KOVCukyiWo3NfdT3xCwcMAtLRx
liCwnlnIVMwJgE/FHS3Nw/JyRujjqVHoDrzY3/nyA9pW0MpTVRomUtOBS5YptBO3
1YqJswzuEs2LE95L5ADkJ2UbSjhQErBMQx6BNtzePn7/7r47tuMIeKk+wsMbBb9h
g009iXukwAuhYrKrmEsh8D+/rBGDUG4ZvoPHFYgANWMCzBcY3dVXGkNhic+kkXR1
RtF15XEbLEiN9nM0SoO5cMzaGP5Y/j3GXFFgtj8q07ERgaDK5oYr6fs7B9tMN2Zf
f3vTst1tap0fLLAJMkbfdpK1Z5cNk8esqgITZ92OHKrwRSXLB8gy8qPmzAtA3nKj
in39LCbF8EWAVjMytHV+UY4RVPU0+DXKqW6Zsurz6rwPFIBHVMDx1pmR1mHLUvma
knff0RVm3MZmughAqJdv/mgOP16j2III+iyww4GcD63TaR1SZacKY8tNtBWy59aG
eDdAPExQ/6W+VvS5F8yk0jKaXqGX4VFs3zeohtJgEKeJ5UE4yDPDb5+zvC570/Nw
b0jKhCi+eYUEFFCzNIvBes6+8G1AaBaUTUqVHax4PCKsvSGNk2IOBcTrniS7Zl3i
ogPIEtTMKUulJZwB3AZ82+Wy8lACff53iWQr3G5N/cYvBW4fMvxaGI/bWZmLHBBS
nW1A6osnBYXxxlf8KjIpYAllIQ2jKXwm2Lr8ryxKAbIaf22xq1al7UNV1566bqa1
1a3SXYg1nzLcv8WWGV+l3xwUfkWTBWWgWhGtjZxz9iZqjtx3OumriXA0T8ESFAUC
XH7dRsCzYRKpSyk5CknlZwFCDNjR1kx5WsMGw+jn4igmosA+zjhJe3y1pT9IbLj+
gsj+GS0OokSTDsO6Ky9MTOeK70enghyFyx0hVQuNO24j5zO0M5ezzuM/bJ+0G1a/
qNuQbdYfkdmzzuBfh96va0Sjbk5+QuHCGdRDp3XJrTKC+Va7lP4p76jem05SCcgg
kCnFGC6oS+IgES7FIoxNJYbtWo8S4TK1e8n3LXq3btAU8kRkLXMQ9cy63gOnnitL
Bta+lPSlX1q+vFc5+ZuIVcfzQJQCISM7AqIAzq/lVlmvY7Zfaf6y2vog2pP2azrc
iUaYtK6au/reqaO51838cuFfuAp6hw9pza6win6AHjb6HYgBChK4gXGPXl6vKWcT
EpR3xCcPBkRPGyMTqrRCPj4L7p5HZBR5fBatzXS6JJORzvJsLVVnPIzcRExWBpcs
/hbKBb3/jxetYJw3yoDlBbxcLuN4oBjuKsZfeQ3/uHshKycpL6Gn/BUeXSlKty9S
wvKNQXoI4D3E6AaE8qo0El206PZDp7E11KN3XEGXd2rE0if0IriPSpGJyoGhc0rS
bnXb7dNNAHjHm/jWMQmhktMn8dl4BX/cLmiHG09upfsPnvtIr1KdM9DJ7SFyFG5t
W/9HppXlQTEugNjfryybVmHnFeQ/XUhHB7C6arpxui1BDzCNCLCFcplDqqPO7cEK
BZlJbUnS5QEKKnPHUzcS6Ifi/N28U76fRHLEFcEDUxNYTggpYWCQH4Ha82AMcFWg
d2F2uGfybe8bojndQU+yJA7hoirkWS5puwp5pMURHL71y4BY0goA58rXTHSPjo+L
JE28ie37GM+zZQAG2aCxQT2X32j0lq9MiQ4HCKdKlBmmeZyMWaOZFAoODTl2CTKl
fNqx8t19LR4UhiYIfyQ8RhXM2e1yCldjXpFrEYlkwb6MKH99GwrrLnPyBwyqnDb8
0d6aluhHj4Jgzef4pT057zDMGtTer7Zz2XBxPCukBLWTrG3jVnPsxwUZLoazLSSY
wDRnQpe+6dNUMdlF8CKKyGHvBC6kComT2CDi5qFyvhwl6ayHE6WOT1zDe1eFypbU
7MsF4acVlt/siFqUi++MWeEJV8/3NZGX4umjkocI/oWtXtv6uEXtM7grnbeYkf8m
XoIDvkkbKslmdSdUrNK04Ka2awBSG4s7H6yWEGalTAOhsjfbQO5nT4yuYPgA7n/q
yTB2C4r7RifhjtPD/gY4Gua5cmGkbVZSOX2clZa8UtWuDSfTCBnzuVP2V9AOFUpO
gkHCbRKdKenAT07zepn9+PV9DkKvP9DLybU+UNwIeRiQOmztMOvkS1VD7axEvLT5
BCEqzwzEyMdnH2ICP4YfFKZR9ETpwXvWw8c+CqHX9z3+rMLlNBSgl+trpPt6Hp2P
9+Vjwgq6VTlZTdmc/RcmCgHNo2SRX6S2pVKFELNp5uTDDuhEWpBHFSQVRbkoh2vZ
BDsOiIR89P4geXDXOWX/MVrYezYNg4Zjn5HjT+QEi3Q3yQoI0389IqZo498zc6Wd
OUPhTcwQ0niQ5M/QeMvxeOwlQiY6rp+oxefDOusavUk4b/6S/4Y9RqX0mklxkX+z
d2fo71Cz+ldGfDal7i8G7cqbZ+gOJTmnS1Zw8UCEyeR13YBeHAf1cSYv76O6zVfi
Xn1t9j3H2YqD3apSNmPhGEScWp26TP+UKoZr2nK45+414zHTK8zs0vntIcVJWG5i
Mcwn6HRm7379Vnu0bmFZtDbkblxr91q8SJMACK6EttzNLS0Bh3yznPsRHqGa8/+p
poScIl/HDxGzolStzslJdjLi5s3ROl/WuCuF/5yyNn+cJI8JtA8bQ4yehe0cG7SP
0dhqYR8+jtVJlgYM5NclPxHiFWJNBu40hKPT0GuHofPS00x04DxmYKfBRPBrZs10
J3S1trcfYRCD4hkdU4wVz6Irp8P22szJqHjwFw5xCDq9Tt7xrciapvXqo+f+j4wM
sykBgfmWvZBDaz7EJT0JagrOFGx/AQF6SAHNuTexudsyDzuPimkuWB9klqHTbTgP
sewRNPWi3+ACqOLotTQocnF+jG/LXskc2bsBArmJXUl4bnJjr2YHpJT6O00rSHPK
5ALhMywjsDAJere/gVlHDAmluXzpSaBXEVDFvmnqHfpmr+Ic8st3OYM29LmQ2Hbx
2A2BSyDoWVv62jdPILjnvHbN3gGTAVnI1XI5XDdNo1h7zuxOnJ0eycZvN3vZGK3T
dEwu0CCz8WZEb/t3PbiswOb5V8M2ynv/+qDVYkXY1JQW5gPGVukLrvSo0rC4+P7j
TYwkgWHODujtZ/iKPFGIXAW9fBeLNGoUzkX93SoadolYObwTjHprIOXvNoNanJyt
MiolOHFq63Y/vN472/BG1pB4JwBbph6MIX+mqh6wSRy4wkXj3aReLBLtsEgsr3j7
dPJtoeWt2N4C+qg9lg68Whkd0FJWshpKR7Rtn0g3HaPLqb1I/F93ukCFUUcaWksN
81QaS65m2xydErFAl3E++fs0hR/AY4p1fwfAOp/5SXpyqlcg/hckjo76qaTUG8Bh
kNoXxJwzP+LSCdy0N/A+yxXKhW1qQF1W77hd0uIecsT+xbHoHUTC1alq5lJvk0e0
3pCG1tkcr9oRhKSjQxsoRSmZMVp0Z+l1Orjhjrx4i3OIAwUglg/gIpRYc/Ef/rya
DeJqdNi28m/l7MoMpxzth/PFR0HPbKE4CJx3+sFGIV3I/dTq1w1c8qCc8abkVT84
ySilfNlO9FEBHNtstDWwV4qjyjo/0N33Eqj78ycxAGHQzy6puJ7GspHs/y7JYGTi
8Bd7pP3SYUX1WBhXLgsquWLzkscXBu/p1y5XXx2mCYkUiJbNdDR+oqSXQccmjvzr
WgS6SQNPcAlqvzgCQLdYpgXuzK+40yIwUfQIBVzJ2gbeP8Izi8ASNdUptoIT+2Pi
5SNqxxkF8VWdWySOdAbfR70PX0DUEJZIm91bQt7s8wpgszVfUBUyljq+eo5lrDvJ
jkQrnha+SXCpGHTaQsUqGhfXxd17uU7XFiYhY1K/+9uxu9x8pbr3hOXT0Se9xrB7
kq0tiTvEOwHgol8pLRtoYOKDfmOvGIJm5GLfgNf6xYyF3sowhSICsWR/uTahzznp
1Kl9wPSHAk55pEb8ZCluIMNH13gbTmoMWJx6NkBdaXq0kj9IQACk6zP952DKEjuj
R47jvd4LJbWwWhs9f6+LGCAKWgVv4UV/jmNzJspnQPs7n0eILpmvodBytfkd8mM/
XNMthgFwF3qVyKNGFheV899dfjSz4QLTFTXwmYFr48Z83HCijzpZ4Bt+69Z4gP2j
JJjCfEfHhtu8jTfSE11ey3mrVmTHALO5LGVyp5sQOeu/P2yAZLUnKQv0EyazVw91
99my5HDjSpk3VfEsLR2ge4/OxbvT3OD4LlOM9Mv8z3AIS/css4L2gg+wNNtMuKmh
NyJ6epVJLx/P1z9UmG+dadpcEHTzzRLogZhvF2Tyqzncpu7spe4yORDIK1HaupKc
3JTROwjRXOQqVuJGxtcrkQjxDBJAU3U/ZAtKLf9yvF+NhSqIK8DGRPttBKppYstZ
z+NJdZPJBw4YyA97qpO6czfJeYz+HCdpluGe+BvG1CDjHaE/w8QL+43CtE501x/P
9rHaQPcE48kH5lUUJx8LBpIrsVJ0Vd7y3auD4Z4qJZimBJQGN9ztdWERDcFnWmOE
HVFkpO/htP1s+NxpMyPU6SGn7k5zAfMLrf3grvtu53/iN9ar9WqG1q54b8h6HZGH
uunLOZJTWtFWSso44CXCmTMwulNJNBFezC49SpDhAOTD6NbAeC3hJ6oxFT8nBUqp
WPzfS1k7IARHP/3amAZE9NnR+wQUC6LnjbWSe9tccH3s8yOg7exy3p5E1+c8Xoo2
HcjdQ0TbjQdUzjpMNT7MDcCMYwUsjBReNnPN370ep0SnPX+zQcz4raId3jy3Ppth
FT44HxtOT71jlu8IavhHPQKdOK7y+xmoL5YDFcJ7zan8VVPhUnnv+HtIySmRTbEU
LQ15tEd7q/rHmeUlAQUMSyUfQtXBejE0DINeRsn6IwM5qMbcxkAgfrU06+Df9tVF
6pQFMw/qsskMPpJKtoHTi7Wm+VzFnX436ZUrxsiAMVAbq2vrdGePjRfkjXWIN1pM
AT4RnNf6Dv2xgkMagHtTOJYo5Q9SgcJFKo8IbEX9D8LZQPfXw5StzZKNO7zRFCvw
qny5a5C32BFAjZ8i9bsptX0grARQrESouY4JkUlM/8uZ9BQausH9s3jK+ZJhsBF7
niGhdrcAQ3ke1LNduNcb2X+vbKs2i1AKxE0+HClVSzf13X/Grur9AGZon2dJ7co+
ui237ns/omJYgYxT9x5cTuKXDlv34MIZ0ZMB3uGXGbpGyeJ8Ras788DjRxeerzvx
bxjN46llGTNWn6cSRPCgqfDKu2sTuBRssEQpnNWSOgvS7ggUak4jiRLC5uADUNws
o16ZvBoz+R+ngyN+VHXXkVizD4elS50DB5dFLLq0e5ZbGsbKrMjydG+o1iL8H+zu
Up/nfKLLpWrIy60D41lBtsb0aih3yrY7TAP9HFk28TtF+BcQV9VR1qfZ21cPFl3Y
SyiUUdA0dzoW0J42Cw0DxtsFnO0oxpp/dvKi1ZhZrzD+XMCx+/sk+h8NDqYjfKQe
fN7F9f9FslEDI7fE2WimQs5yZdNRbZPXlLApCVPbNi0B5/PnYeCUMqeKmwzdtFiF
blk7ZXGHtAJhrQjchHdK7mCE03VOLJWHKNW0aRD6MhH+EGEbH+EOQoUTM61dWkBd
K31ZzkZBVkJtxzTWyVZXynu+BPsx0cIOoaNtT90x6VlsUcHFDLP0ExGuqsGk/UUN
Licj1mr+j4R9Jy60niW2EMN7U3HN0kgm9HP4zWAxK9FAXiXPtoD0QUY+jdhZstgg
j2+2TxCGhzYWcXOV+2J1UVhTNo9uGLELRvRwRpjUTr0sJBuJjX9/RFgJ4oOYea7n
EWJ2/A1ypTXIneoALn5dAsIy2cnsLkNs45SdYCMD3fCybOIlA4n33G4LthS0YF99
clc3gSBoHmcMzk+NVOYDU01nnjX0ExiZU05f9smyeyp24CC/lfJ2Ru3sPwfVD3WQ
4Ld2ClcgTCg/ieNmp0mwhjIaV57Uy3hg4HQlNnFwAHqAA2l8RMtCLU5wGosVQ7W4
jUy1BVkclCBmkghS4hzaxs7wRLfriN+WWnII8HIgJFMPGgzfxC/WoeZzAynYsXjv
g/xU+L53gLYHx9kyHFFdYvUZ5Z7oEbhi/IRo9ndNGqZ1yridKWxYDjL7r6VID21+
rayCh41M34MDOIFh9Vl22ecGx+sG0PBlRucI0vt265NlFfH+VS+MNlQEN3HItJx6
zbFLVI+2OVfDCoWUm7DNmMum9Dh9L2rUW3ZWI/yGwlbDYb2mT6jM0z88DR5d8Hk+
UbMy6NVxTlIrLZYxqyFmBkRna9OKJBfrNEGgIkaOeCoRGXVlHVvbeiRWV7N/GlWt
zc9I09w1ftGafMTSHdEU0JXuj4Aa75TLAGXb+PFVWOGffP0xsMMMP4wK8/LeQAqG
RfTKYwmYAVFqr02rl0sYg2wj03HjOA8S+39WX7LLxZcPsTGKPkLGQ+TUDjeW7u4G
WQj7vVBJO3MgESQZJXCvTDQeHaBS1ifoNpEQ8gHHb7mSHM6RC/BXbMic46w+yUIO
i6KWbIqTVrMW3KdqU8GKU1S5syVltKikjwCpvwex7JmDigsunREsU7RfFjGCbxuk
Qpdr21OCtozk0ZipEkFBSLr255+Y0uxTwbwvxu/cQftwXmIqMI+Tc6qXaBXr/XUc
RzL9T0mV/2SznekfC0mj8DIqRl+WRfsN5IRQ957Byq97TAo4S8rwaevkefkeHFoA
yhzgaG4DvSSY2H1mDUEU2a3FuoOOgtlHyWiVmaYqdPDzf/em+vCo6Be4LO/SAMWW
GhoG6biEsN4vRhtv7XSrNLNkjBPFj2i6qGFDJ+WxfxMZe3hb/fCWT8q2r6zueybt
Mud1LwveG0DquaC5/dArICwxoBWLgNNUr9euao1G4kQwhOQkE2QVk20JHGnkvRbS
U9gIf6YZhCwh6qVEJGLe9hwV9zI5BrDlYQQGLoZxfdj+vF64iCCQAUry/o2JqWUi
Ny1rFoHNA32izHqozQMrNS43OOi1SeFpLL6StfdmzW9/IqufuaoolB3udNbVA8fh
4J5W0LMRKwHYeEiTeE6Px83rLcBAXj5QjfaaT73mze460DMQMzExsZJPIBzI3CFS
K2Ni7Ak7dvnqSuKgOLcEhRvrsQ7LqJWBZJjvOXIfog+VNeZKs+v6oFOW5awL+3Jd
x07hT0Oa9nK/S2s3WHaV0qH3hjiSQU3FLt0alfRBQJDWDB1lbfOrNs5QkphxU9tB
2g1YoHTztosv0dkTkkDtCAGH/gcPkXNnrvEz+Sud/lV3Zk+XkoyCB0Aeq4RnoDrJ
LQ/ctxZtf1H5x3VRIQebddTIdGlmELJM09/gUoTVnT1DjPUk8ugR+eoECf3K5b/t
CZm6XSFrPfawtdyJSaFnWveccQBiKwqsTp3r2i6UyLdPX6hrXpSN0OGxEGtO0uEC
llt5WxoSl8w9/VSn/58C1HPwpN4KXilHeZ45hA9hEXxDvNYSEYgq5LE6PGayx3v8
+0YTn2A3WMxrKGgdrslLBLPktJtxLIaT0BBl0aux2JTlWrHO5J+XGl94LFZaaJpl
jkYKJ+nJHaZLgqJ02LD31rC4SeOcdC0cpq3fJJpJmgnPoAJSwkPm1icwpUdCUk0q
zCypIKrmpUTpOKelC04As5CQiqYwp1X6kwHgABicn3qTm14WjNti7nEV0iMPAk4R
+bvMHIXu8zmSFdW34CqXP4fLqDkn3UOMJZ4ejEw2HycckoS+QF6dfC16LtLOkGrf
rcdCdaMkGR4z4veR3rnApUEVoyeztzAKiFecwu+5wtu00IGonGocThEaSuIVD+sy
QjPNSWWifzUCJ6Bq4dpV7Ob0f3M0cnF6SmGOFDdt9NpEg+odN9yk9lupeQqsjx4z
d0rgIj4/mfW/X1nEpc1rIzaxyuatraFVqFnx8bY1EH6QBDTiOGdXwPh3WbFcphuA
NYoGlFc+5z1AdHVOQaObQTuNCS/2Db4fdJvK+4NfuA1wEb2DeiQfQxYrjPUyn60u
1bWC6ZzJFN12vs8QmMuoRVMzWN8MbecweCFioJrGqdXRGo18yC2FtjJRl6DsS22U
AoNhblFI7QIIBt4CzB/VIzmdCeFE0riksB9S5AXtHoEb5I/2Ydt2MA3QJaqKddpo
z7/d0pwv6FoTplXaRRzxQjR6jm0muMG4I8UZVvY+BxYRpzQDFW0ggGo1ePcW2j8p
Kh2C/kBcjPFRbTrjJk0R16bduGhRQc2dg+ciIwI6GIDX2M1ClbZcq61wQiTAkkQp
chpbdUfbKjb7XDtJeukqnLO/BQP6trHUFpRW7uwTcydeZe31H9mhz85w0PjOP8Uv
qJLA6frC9BCdfHo32lrYoDQSgUYkjVoKiJr3jYJ/4/6XfVAGHZP4m2zZH4calm+f
uBryNVKUs66zMAwuRb44ex37xus1+CTzQGnm6joCT7vrWxagKGAnlQVk7Eu7ISNZ
fq/OTWI3WLpzbSEtgT1Wpb99agbIA4w2SlAa0ijjBHNhejR4YapWlLspFh1rplYK
ICvAJ7ruRJvU6V5Q4hX094d6ezmtRvIBZXXoAsuKua8A5heT+67AFPHiQfi1TaIr
zdNRCtR+5mv8Q02nnqC+4ZwsvljmWfPoh6wvwDp67npnfG9B3jpd01/L7LfQvwmP
h/vO6Ik1Ms/K4LCDtXkgWJSh7CiErlcF8j9PMpLwRLJkk4kNKq7WtWHF7OB55isM
R+2rTouWDVK5e6crdk/4CdNw9metC2GZG16b0QERxvG7bTSXlm9ThOaKaaNmoPc0
1q+CPy+W5v8LCwNZdo1a1JCUUQ7VXpMbTmLBw6EJusLTbyiFzVUMsHCUaokyDY/N
bcNXm9D6rnZh6bWup1nV5UgTpEa8xBpGAfNZoddyNpwecKyiCy0W65xzvVGDU2uy
t8HxhJuXte1NcOgOaD5j3wr8NPKpNLE1CQH9obLNF9koKlhk2tbtVb8de9IrcK5e
3ZHZq3AVVkp1GmIroM7cq6zt2wmtwoh1JL6/AQNsxda2+BsdysonSr4MJJherMDi
UndS2vSVq3A5Gr4UDEdv0zcX6p7ARQacL0QDwaURZeRj4kd/7MfZgEN3l1z52blM
nutl0L8LUGx9VoX6I98/r0Rt9VScmm5ayHfx1PG3fHAAgSLFl/5NsSH2HT0ID0/K
HyfVBRrmqsf9jvL0ltVFLlH7D7NYIqPb5v3QwoRsv9/sWPMlgYDIasfTyc2bGl8s
oLoehs1sg3j4HUzXLidqkSHeSQXZgje9fivR5L8LFHNWrQ4QNI6pkXyr5bFmxm1v
5kL3ZUxHzuMCQfS0RZJzbFOa2f9RfIonHzyFDmySgO/oTrzx020uJwdewf6x5ptW
Rlg2aOKE3L1nXJtM3wegYQBDimE5339WM63GdRYEbLoAnfPBZ2FMN2Ig5SZ02+oW
LoObAS+fiReSofaTMdp8I247mbRd5FPTgETmFHycMIlPeUaEelPW5Dbl+8y4cZF3
6XpYzIhugs8lXRc+O+Jz54ZC4Lby24qJ3nYtEhir+tjmvRd+b5DquLe455K0ypbM
Y2KgALD8ibJj2ivZx3nlL5TzWNHz5WPaFONEuiNlA9YnLLIit18AvLP2vHGwuOFx
YdavgUnmUzGPWe6pZZA4bfUzw1dXFIXFkRk3lNAIJy3sFDuKQq7tqetHM7ZdIqMB
E3GRwB56+57Ah516DDogH+G5Cmd2TVvMJzHea/8JzFvZtXWXCguPQG6aSVoPEFQX
HrYcGwDTl/CJSBNvx/6tV0SEm0PiMctBcLe+dqTkoQXnQNuaRpp8lsp+YIowTfO3
7qkOdXnXuh86WSlJf8DyWyIl5qozJWw/cscLeKd/mFp+vaPIcriEQ2qD/oFruUP6
303DZ8lCSzDyYMfmnLiF7XnS8QGDie9YoFkkximQhsA7db+WMWIK3t7hgnUIo75p
y5zR2MGVsgVp0cpLAj8PdDE286e+8G2lsSHW1lA5IF63MYwjnGFNUGa5R7V7Jf+u
PUoRn1gRzHzpRwShbs4UG1eU+dB1dAuo0ffuctiFBQpsIHUN0L65jCmJpjC0m/3z
2pFSY4k7BIME+lEgIom7/9tSuqi5tDgzdcIYNsNJ+7ac/w70bOVl77soM7K93cmw
67CcjXmW5UN6ZNZR65j2Z2lptxLGdRwT6XIufRhUkHfqHK9KvhsgAkeorbpuqvOF
ovfLadMHHKdbVcNeOAssjDpvgu59BIWOJW2cmQhBSrReQXmFIHdVBUyEOb9zvo64
Bc8fBTmWyBK+NcVZhXy5nJN8kFyzQKns2s/2kNG6Htd8bGKwM65lxTv5nqYX4nV/
vOpwME3EeOwe6jiBqNF6Siuver5NEaX+4fAQScJeKVtXENSAX+euhyOfC/d2k+Px
ELJXZnU4Oq3iYiwIEdapJ7lYlqz26Eqhbn3MyzjbukmTg36pDt/hUrIwfco09jyD
QUYGMoNF7sjAx4KsLbilUVqEC+drHW32FzXU3mrg6+ZAgdlYm4kWBx9wnrUw5rNl
5c69WK2LQlhjQ8AkmXS+jJO35Ld1C9HPpWsDjb06aWF9O8BNW2OfHauihDzCqJji
EP8F1L/vit3x3aL5Ks1fBRgNjbWkQYPv4JI6F1YreAvHwjw6vxS/tMUMxLgl/qgW
QA0pZMCfgfdjvrMxETmqLhPJnSRHtNfAKMoGWWup8QMKpCe4kEAEPn8z/iPZv6HL
LzYf/jgPzfIHeZ6q/73IU69LeNq+jJSUEsSo1eEM+/zISyAeE2DMe31UecH7jP5o
VqAL6xoBEc+/rk1yPuqIuIL5T1OJDrbrfDRm33O5qfZNf1RQel0tJldgPEDtg2nX
FLfUckYyA9YD5IGgZl2b9PkGKeMPp6hDCOUVM7DWM0+VntYu42wRIusQFfygnQ5D
MmqbV6n+g/PAp7ejV8MdxhHtREUKWKHwRElNS8fH9B0KdsU2uX44OWgXQUuxXp5i
zxegQSDVQpgbAGODtvbGtmKvhLnlBpVKFFrBCkcuCYEok0r8Dq2xlUJ/Sk5wSefQ
gjr0iIJJtJd4i+hdxi135SOY9mP+RRpSkozT/rvgybgkw50lDS0qEk0DX5iVazwZ
Nd4G17IJ3azCbZIVrFrn2sfHYi2LLnX2+lFbMz6Q/Kigx0bztsEAhktOOreVbtMC
Zs/BQWQsXlIx/anV1wK9kh2L9EChzM7Rs+gzdEhWhP+wNPlsKijhPymSPZ9C1Zyu
nXT5AYGy69OLO4nbpYkv/BiG1fezAZ+c49KMaEJz/uR0rmVfj9BtNCq92jHbpLZj
gnnw+CKu0YXdC4qNabhfSRXNCiACegKdTdCWLN2FhGseSeF3xlm5+FluDz/WGBuO
4Y3KqcpxD25TeSKQn3Wzky9gFGouNoXlOYkxMONnNop2ItOOnY97A5eIHBP73fwd
IGs2+wxJSDPt1UR13RpJDDuXkS9Z3XG+6b2pNRNRBu04xWyUzLOGInPlrYRzD1oH
dHkTtTkqa8EaPa5/2SVTt+bAMyJAJj7wwr0KZDabeayOoFvvss+31me/rPKeWNtH
mnZlavNW8ygSYfggr9xyg3vwtAr8t1iiyjMLTqUMqxOrj3Ku/BJN+yGPgexXGcm0
O+8SBvmofV0MKotsHbYGpg3TcojbH0omhXnLzg7tfF+dWUniKqJYxUgtJVzvDFBu
IHk7vg86uv5bW622K5svUnxD48ASfEKT27v/64NBer2AWqw7SKUS79J+gRjNroKb
Iiu07am4DP9n8CgFVmR4inx51au+9SFrPugOAtk9a4AnEB04VDEHoxtBerUdUfGm
zR4dpJaGZxrmqXQNtk3RXMwhEA8/HabDw+5qnqhfWqr5QFQ2qjtSb3ms667S/bCi
xXmGZei0fpgf68ZlyrY2AJ8Ik3xVkss9HImqNb45rl/BGFdvZ8a+TQhM8kUCO2ul
8q7Cv4uR/bM6cYI3j/sz5GpOXME+iEX2tVm/Lz0zXjiYym+aTY51zXv9zk5mfzmC
/qJ8x1vYk7DKb3E/8LOj8Is4gJsCJDEutibskaB0B0Nmj8Px/wuc1dMZbT56BSBn
tHP8hstqsrRMgRV5mUvzOwQFIxg2sRLnrhbdDGUeVtu65qZp97yrsyhugy9qhptI
vAXeXd9qe0RZJfUcJ6QhZhbpFcj9Wujb93Tx3nBStvkGgwMETC4Cf4QAWUMEjAsu
VZ1tcXRDPtsjoZWcw6VxHHB2iKvIMHK65irQNT2etpj1d6tOLyDaGzKhRqA9E4Rb
RlYx+jUPHpPkSCbZZDD2onsL1MZS8b1tnV+RuaueqiYHF3EOAftyucr9ZLxFmx2w
htL8uJjtHfvLETxkfzCTMjS5y5RWLQ1G3SLOKp6ysa/4mNwzJXQcQ+UfVlAziwC5
36xFgyYHnPGlQgeKSjkkgThtyqZy4qNJEvVYB30CJQlsDaJhy+lXuOh2zWidhdV+
iE+UK+H7no77uKq3AI5Ktb8O2wbJwQcW+c9iPAzRbBgvxBOV713516xKS82/ibaO
Uwzqd4/9DgSH0vJnpY1VQb4cutQrj6hfbjsb24Ta9c2ti1+jdTPDVxagP1esP7iB
lqeBlIaieXjDw0B0wlw3cAu/eZiSMOSI0eF+bKt6EVw/numTFhB+G6/Hhrj9Qypy
1ohPJtsSxkkjYKDWL0GbchZ+muWxF1Aknq8ReM4YUlXfcJ0HSWxRpx5aEbUNfjtf
6O2rZnOhYoCM1mbVZQ4J2wmxTo1M5TfrBjjUPeC7sj7P1vg59iuz5rBg/dhcGh5Q
who3+Fc3Vto5cyfvPTO273Ut3e124dthJSfK0/Dyuv+GAD8Ajcod8+EvSJ1z3kB1
vHHkqAAYRJmWpRWrgbMFmzBL9bxQi+LI+MQONJtqRbenaoVAtmiFcJ9cXW4zzVKe
9oKsQUQxvBue0IbL8W3R4R1hGzJ5o8XTQgQGWDWTfAgETyNdta9L8X54QWu4SGmU
RJJhOsQrkgNMNRHhOZBYm6wg69Onqs29upUjJMb1m35xZSy07CeSqEYJ1ZJWHMKK
TXndULzL9vM6Pl0KyMXoXT/j+u9Pgag/EI7YhjkxKTqV1GcpWCZayHoJcrVBu8oQ
4vCvoELhGJPAN2BIfPrnkT2yHhXDpVeJLY8/9vTMqvChc/olt8lIZUPvVya37Qse
g+/KiOOWKbzG6qJmbCWvyoyh2LbM1OWFrnxapkeKMmvBo9+I83iuzGpmTsDXvwG/
CvRhs1dN5t7n8m0jHs+rbfaZIwWng5oWt4BDjo8lEox+DYFiyDU5imHATHvnuPvb
+jA7sXo5nsKBidQOHnCTHO9GEwv6bz/l5r6/OaGyRYo9+2YNMQr1G+4YTD1lxUWs
MDHSbJK2//PeuikTRWgcxbrXtze9GWAArI4XMTYA/6PeHDXp29EtasVix03anLDW
E/XY+oQtR9yHbGuD/nB59bTrENc6wXN1n7tE8ZKymzZtwf7MMRRwLYEeaitfHhUY
+fUKa7tY5dp1sCMiCkAKIUauG74j3K7UevagKQnQMMdwgbobIjgKN8+FwSVFLamr
a1JiXcSE0quJFMtMvYknmQ/mQZAiUTqE4H9Q9SxJ5q8FsZygaDTuvchZJOaFKOXT
LFuaX4iyLrHrNjDlvKn44fPq2g7C7CwAOWVyRLVaMRVsLSYjk3TxKzOi5eLpVV/6
ll8IymkVFDhfHNtUYlhc/NH2jL6Oj8Po4RgNlsl4QJ3viXDZMp2tMKmc1NdjPBV9
1FR1EkaAUcbKaBbilzdeZiRgfOesBbwv6Os3edSXl+8xd5LrEUDILyBrOWMF5JLq
V3R6uMNxUIyfqFvkJma/RBY/J6rKxbMPHirPKjMcY4Nr5h1jNBc5a0WvXfLtKJOX
Sk0/Y4QRTuAoNqO14su6UHTDypjWmv2DiECwZVnM8ILlkBj6EHanaQbanrrdxGvV
cb1ygSuqgzuOlt1xGxau4c5VyFQ5d+P/3lXLxTIeJt3RgCahy0xX0CdweVY7G/2X
u9WvYMDK8vPgNGN1aGta/hfJ+MIWLM8SFYPgMdN3AmXijjg9bnkor8iIRcvev/NA
4uHXfkYEjz1425aQkMPZN3DoQ7NonJ3r6EpLcUbp/Z4lPMzP1tJdC+xF3pF5zlVF
6aHZWKtGaR+UwuQfvBAhlllSPaN7mzQH9zsWHOO+Qe7uN639+9/y5QBcO5WzAHpn
vmasGKHnQgJYwkIRd6y9a8Q2e1nVPGvueYP6Xet574QCobzC/vze5Sn14/5fdA1c
sSSsq32WqzZgaMVdnjzVgqJbvIrd46VhGit+HR5bjA5WCM8+GXN9t0KOKWr9Yizq
es5Gb0jlZMJfgyN9mnFqdtLP0KiZUq90inbRiroSAv3t94Th/aKLNR8U3XHODt4v
+1S6B/XXJ+ltyogiZkCkTgvMWgYeWM7mO9HgtmUe/Yg/hkCGDJ1U5+xx9hbAKRdj
kEiBpVst3E43flhvtLWk3FyWYZzXz3kjOJj/Nvf1fk+hd/719p41y2PtcZGJLw5m
wg6dKbtfZ8aOP0aOvgxLdumu2iwgDW7RmEDr8lsWHEOyXFjyCb4J1dnbY8XOiXVq
iMkUEgNXoYQ5blsqViq/bmcg3RMkH+PpcGy7SiWRRURSZwuY3J/bqIghdQvx0mUG
i1bZtQ36dEqzk5662/bKAxvXjcKTKI8mnXdgrjxXr4btpThnmAexOLZh/+dRZdg3
U2PP1yIZgvaT/UVSCdU6sS9YIrVPzilwEOFmKDld0qNWp5k3RTfFB1LCL7JEwc0L
EfBVnH8lrkrVSUF4VjENAYmd9/B8aklGPKtPVZAFrJ0jKeKMToq99JPkKtx9GDga
p2Jkgx3IrRPLtLONUODxxbbZr6pDux8WPOAmkdNYWVj4YoR3JZotohyzH6dXtdPI
nh6qRzEeX1uUXjdc4riXKL+3/OS5reiir3k68FPLQr92DFH5Tw92mhMj/G+/EM3Z
vu92QHztMxoCsJ6jKGQ6+lGThUXuJXChK2fySZYC4QBcAHyts30vVNbx/2l87gA7
s75OvKKcNJkKuSRzLMe+ft+E2w9qveYUcdLMP/+iL+38s7o0FhPUlioklwL8rfPo
clMj8oiJCCqw8JxytKlyQ3gKN7jRKj8MaHisZxc+UsYHKUdACYqpp+p16iKo8eFx
LNUMDwm6JlODVNqb1a02LiUQUdPRSsO5oBSWU8n0dEq6g0h0MJRFMXACyADGaq7r
TkFItDpLFisWiszvSrmOQmg5w2lC1Da98ryXQxtNkUnn3F7DrzxFqp7g/IjvgPEZ
9hql2UjFXwYRm66ghBWfq0rFbp0QvLndP13NX484QatsNPwDDf/yilMwakP0V5ns
qiyJcCxTPct09ZLgJBXnpr8ZgsekVfOKBXYbKkrMmHEYlHeSdWDb11zmKRBCwyMg
4ZSideX7Rmi8tX8aJhs+D6QGpZHJUvCtmIHh5EhgOgOx9b6rgrosV4PvKjEN+76Q
/5r1bbw05qZT09TboaXpsYYRWlzlZ0Xzcr4dT+7J8Ii7Wvvv3dIzxoBpd8VdgGnt
ryo2DEQPo1hFacSLZVvWqO4al+sAz8bU2XdvwUMDZI42ihNN0aT2phlYZooJGM/c
gb0Oj1YUfSnIplaa+jGNBicX10oKTANEF6oc9j/j0pRLfmIYlYJbHZJX9QLPUBIG
iLf/IUgthlw+Q9x0lyI0UtVgAdBsKXgfOJ1a5b6cYMc3FPcXvJ5pOZW58dd3wrED
ZkS1LlftEBWzU77iV1RgZXcgZG0it8ejl+sFkf7/ME7InbfZSZGh7+ZumA1FK9E9
gAthzp00XozJhRuQTOHbrjSSmDvNGJ1HoxEYJ2fhMXukq7S5Y6bvpKcVkBYyUhtG
w5sPFKzsQSIAzHPYwIyrXCemIpTbI2iwW4wtPhnY6jfbNFCJ9MaN89MynM6FRO1I
ldGc7qPK0KwWQUmtwE+2uBtL9ntUyHauZ9eKpEQmpqAFKwtA/z+LpyAx/d2ozEED
BUIqLuFbtUf6XZ7Y/N5vFcLjEA0mtRuC81IFHk9N/EKFmBACoNR2Ssp0sIozucZI
185u4t5Hn1KTssAImD/OyBtcHqKst0dpO8EPgx7EPik9a4QaNBk5SJAOKKHaKW5X
X49Le8DdXUpf3mf+GOVy8JN/Ca3VPBOWio0qPLawlzgx2P9OWFBvtFQVoLJJCKjE
peNsKl5wVnSMJwFPDy/a8VrMOW4DHdI3D6XFiVD5Kmnw1Z7fspZ5ySwbPvke/Kfj
hJWZ/Butf9BA+3BL72ExXfqaaRWK+b7CNE6Tbssact8KDPTwR/sBQvZtzRL9DhIM
0ymlz0EtKGtVE3BW+PPyxWzpUy7SucFttxBmY/ar9TgeFm0gzeCdp/Um778bW4qe
8RFaYrTRrJyhDzRSh6LunEIMTV5rdlyyBpyFRt75HSanrVpk9tr5+L4QFpGAQccx
ST+C61wP8cynUDni6LN+L+ttYPkhHMQnyO/CvNWyHOAxUrisngas8aN8Xjva6kdV
uAKRchrpWAes6y1h0Y8fryWWlLwbMr1kVskuSkp80RYi5KOUPL1jvBOy9rDjcBvU
hNZGHrdftQow0jgX92ipmEUrD9XaDDz1uHO7WwWhYYafWPWuMjXzHVE+9AiPNH4x
KlO8LKd4fuy83S7b5Pv78avVaFf2R2tvaIP4lTDyHbpLCSDGvIJiN5PDUNsixr/c
/H/H947D3QKdFVcHsc3OMMlO4i226pboIZ4lm85562kCLKMou6sdjEuRcuiETxez
zLkwRHP9vNy4mg41uuV5rZxiMxR1/g6m3jJL979fpAGOTJT/Ib+TKJ9wjIYecJnd
vPu++Ftreab2QleJVo+vbeVEhDotC517/jZOx/VDNSCTgAnllhirfO7litcLfM8V
SzeGhaE4EwlOgKFfkB2qOWl1OE3ea9Myo7a0hOqwKJJVizlvjhbn2Rk+T8aIa3/G
L7FIraKuF8izNoQvTCTCh1gLf4b+K3I6Otruu5jxWc+GLmz36ZuwKS/pF1E003rK
1jUu3Y95tYzDcGC0n109RgUdNOcKky5fzzRX7tyEIDsZgIueCzxBWp1EW97D9lGQ
sh6DdD3Sd1e1tJtO3YJvGwVIMvWN/dHLEXL8VOK3TJkT1pmXSr8RWRVq1W6tTqCM
PVEQqJjUmtxlJD+x6WrDS2EU7Vs16L+AYDlt07YMw463y/KLVJdM5Tj5JFP34VFf
fMBINX1JPvqZ3Do101VYLCc6AGax9v4st0ts43tPGq4oICIyJRpV8o9Ji8k22YOe
m9VLcLWMdfstcYXT+70os7Nw1N1Zfs91uymz7izs2nd6aAC4WYBIM5YTwLWLNmdm
qS87S0X254pOLQSekXT5IfoRLi6hYkk1JxUiKKL4Z9u5KRmgPqo46FdE2aB+rc7E
PWzqHOi0SO3HQNXV58AsR/aMtTEIkZx7HzRs5H+/f9qbK/y9zza/t17jBkxv9qwH
66dWahAEqih0rgzk59kvMCV2xllwg2qxZVOxvTifBbQNbrhops6aH9pQPMdFqph0
WtD/ttC5TFDWEQ112+/zBGYdyArG4n73Lijams9TtkMl8I84mI3/j1bikqPYsMq0
7yfI6SI8War/5PO/SSLw3XGuEhAacKZlvrjLch8c/D7lcgOF4AdyX+SCkrft/Msf
rj8QKiXfBBQQWDn11vrd6ggkf//G8hmY8FXMQqjNOrDh2EovNr0Npv1XzqPpkdgG
CcGw5fiWGK386sjrwoEyB1de8Qyjvx/6HIuvKNlhC2wMGOeIxQKKARas4/vXM+TL
TNr0520rVdhLDaJXwXgHD5pYouzCLmGWCGvyGo+mGFXpFvn+y/JWooj7AWz6u9ig
obBvcaDcFrGKBAf3KmgTOKe2jDRPCIvXulaQCx99eS9dO+8i4pgNyZs9w42ouWC6
4P18JFd0he2k+JkkOrX5GkALdWMexdL9Ee0oOb4PhoT+t1B6aircINHPY2D0ilZM
vmK9LsGFMqm86PiIRT/guZ2j3dk0tvjJ3Quhq2wAGqXMu3t43TqU0Jzgg6XZOqKO
DS/R4d4WlOS6Jxs8CmazZu9UGoCMXJKioX+dBFh9aJ4BS1V6hrNmo/p3SZssz8e/
fhV63pGRfQChDF2kU2ceJdfdNc8ONsvnIcSv7/bDvw2lKMqoAHbg4/3/5SuQE1xL
hquE3ooM909W86Ot7YDjqD7ebbFpybEwIaJF0sg7sRgXLOeYSQ22AIpA5e404Pt3
GvU5xDhMM4UAqXZAuPNmXGrvTWMfhqfC5gCJQt/TzgGalwAvWMeYWUl4i8OJRNXN
o8+cJi4dObhOv2C1M7IKywRMgXnHTL+Sji5Z4e4HQzd8n09I6tvY1F1yTuyIBp9b
R7klKLefyL6hgaTxfPPNz18G2SSQ9wIH9rhsiVhmm8tJ1/yeJbPpCWYFZLT5UTPw
IYGF4pEU/TXKaH3yMKU9Ua8VXZdlD+WArvIVzF8qs9Is3RTVxdpCFYerNkIDQg6/
2Slt7DXRcZ3QgO5jXbuh7R2xl2uw60EPBQ8mOeybMPOAG8f6GP+v+Z3dITeYgjdD
sqSjL0FWeL/CsnONOwWeiUL6UCgmJ/jr8+YaFfFP9gTjPopYc+sOH+t7+k0+bPrE
LX4YYKHWX4pWcA7YNcV7OgLzcxHx1Kng6gX2ov03O1/1YPD3mnnxl6inXyGica2V
k7YNrrzJ9Q64qLA0JU5HSKGxofww2PiVijMejDI7GMmColb4QZhvuE/fePofp09O
DvPHP67jDqIEHaLnnm+vBCO/1s6hj3eLl0zseOuKQsxKP/YPklGVblKE7DVHbRlF
wiHBZSZEMXk9vfQLeIEIhQf4o5iZiE2Z/zlsbQrpd7dyTXOzf4W26aD4TWuCCBik
b/hVMPrteNXcJs+dSiKRJw63duvILs3uC52wm34+ZrURZw2OztkPayJUehorrzof
zPwH9IWLmLV36UWA3u7TcEWbGkE5hf7UXjmSrWA8Jo6C7bYghjk/Ub3j88LWXH0a
rGZhgzB4L6296owiWAqiFcPdJYRNvr5mYL1TcvxXAC3XxMhLZ2oWodg/0uzwTJIG
IYoecWL+VvuDVg51LvVlexiJ0DsUZ1B40VQcki2pBc0gND/I63k7e/7hxwrnr/Aw
OIOxDK2gjcgkVKnjCsAIYrsipe7WCKTixzpn84SP0N2uRK57pzobsItsnp6VW+Q+
mfW6zV3mZvNCvJ/IbQxrCvd1l0TrWDFGmMSuGDjM0qG4NCjpLViiVGkNbRqE49MN
idjYAPNufw1kHH5MlHCYvysXxeELSnWDV3KFxleOuluHmoBOpqCwdf/LFT1a9y3J
6CYlv97zJp1LJdPK0IkwWeDPrE1UXMCNQEBlC+vV4AX6rlq45K5LMNksjr9LI7aP
zId9KxvtZTYPEHDizyIP5beLvYnhvg2SXvHxrquv88fBfsUWniGy8GXrUN8l4N2w
URVmMlRUxxBfdjKJMI/BTRScxwTiRa8LcLEGkBi41RzEvk4goWtNev57TVcBw7K2
LVQVdNptXi1/dSkJiGj9vPboSlxrbAhuKTfRBa4zuieZAP4peUph3OQI0Y1bQDFa
ceuLjqgq15e+Enb2S16IOAGtsiNOuNtq0K47S8Xe/HQFLjwN1OaRzxYem7CUPad+
kJsD1WECrghGSIJimXkWl9mKknuP1l2vNWmbXykjS0zcQ2E+/iGwM3gzf+H/fHAY
TnG9UeTAOZUeieOheuxcavoE+xMGirw7z+ZOoEhOXo/PHNM3x0pZFv/1bDcfRNkc
pJgvw+WDAR+dqfkRJfsPPdLmzknsLl6ZgFKIk7ph8B9DkmDX7V8QkUlWKPHZS5lF
wmY2kwBGaSB3mAHvLAnhkyMfaNY1FfyXa7HrtiuUUP2GwNamGRQbSLOlXj1qlsVF
FzuOnnzkaUKqcemnE0QrRlPi8KJi8JDazWvD8ETnPxYwr7v2EoSBDGmnXqRuU6FB
KHUvUxVkXpW3Pu7oANp8T9iaSiFhRqR1iGh6DjcH3lhWa3XBuYjPi74n96Bp6typ
PQLy6icYbwopUKavkoZ6Odj5R72NMGn/cIMYIcRl3Zj2BY0GtHqLaWM9is0jJoCL
BadE7z73vMTQtU9rPBnGTprVigaW5xMWh2YmY+WN9Dk09Cz47Sk1iCyiDb4LX7EX
fPq0U5Q5/wHK0ndPSrL5ixfI10qZWsyXVtJMruAhE26Yk62wGTAI847Npl7fM+JL
+rr4/7g1vsd5OUvmewOFCJUr5sHn1r4mZWDv5lwAiqsiYa4Su3igMpGpyEBqa7qH
LbfcLxYtR3wFSQm7Frjq4QbIYUN0jXDgJFDa2vFvoub+mU75ZchxaioGU0h1IsK2
9WNaQWS3R6tcC/1kr1RuYW/51kwEVByDKb9PAaAaW/vdAOc33Z3wjfUk4E2CAi8J
Hnmit6bWryErLj1cAzFIUjBUl2mNK8joLBbm1RRadPbTCdw6/nuziJaFjmcZxNLy
7CEkTTDp4rV9Vc+IjOljL5Yvr/BjAeW1qv0jrvsiGKs8kfhg4WJJaDaE0Genbiyr
8bqe4l6GmJWvQEyuFXY0no+ktMUBVquPyx8OvE9FzRrhf3gWo+bUCERxp/t1680u
QmvRbii0tlZh/EkBeXBdHLu6c7i1sRwpF/dEPHQ5cG/Ehv61YxFYkVXPKchd3baA
0Mm8mRCMcvIKQSIXe0xBvVQmpras1ErPZURrQC++qwhtLPJdjMRm51UUBBmjDBKz
iKT9vhxTFAc8RdJ5IvZm5WGYU/mZw2wB29MqwUmoifrk879AdbFXCbqxdU9oZgFP
iGMIbdKcEsIm4m5ylD6N8fvfo3MZ9zY2+Y1FZjO/YeOSn+4ERqQRsFxzKrDtvd+T
upH5JqCHUDL7jBrgwts4gmh8x/etm9bcAhsqHeMOl8E10i8JIIWpRESdXUX0ErOA
hO2D55kX62SAvYE5BkRvdoWHf6bV46tDasZXGu7Oo/9NNuaRBKjYS2aTKs2L7PjB
Pcnb+LdYV2mE2GDl8XvL/S7/iQcJJskl1gu9onknuwgy02cClcNGKbzPskZrvKef
fq61DCFpWeS6vbASCy6DSGEUD91d3ugpqPnnVBMDdETtSe4Nd5di2gjLUZrmQoba
rOxd2P22Ub/ee4Gyj4sc81FpZcy+cUH/dpfDAw+dBrVZtZDTicRinr4Ef7F3Tdh2
AM+H+/SE3R6q2nfV2Lb6chdH8VAfz9OdJ/G3wg1NbddY1As5NlctiZxDsA/MCTUZ
j+zuXyc0vGb+qR6SgLSkWba7VLui2lmWsDrP77vJCtAPY+sO8I8GSMO0Hh1kV5cZ
ZnAr6YYhXlXes60h7YFwQdl8VQEDnAdWJT/H6ZP7TiJ+/+XBpJRdouLkSfIysT9K
4kArg7qhKvIeu8bRM2Oe2Hy8MfzOwCrP2ihbWZJePyXI5RELTTBM21SwxpohkZh+
IM8391rEwJYq8xUrA9OYXbnKV0MuJ45ODp0p2eWrH79aY1hfV9M7OFcYKVLoTj09
AfLjOOLOCpMAEuJ6YAJpxLPsiKUY/NKWQAHRebNldwlUrXuo/iQqwrzkw5VyCkGO
21uqo/djYIdzSCpi98YfLWHJMoFMW9sopzkXjt9d5UF8DaOHh2UpK/X4R+vQp9ZB
0BHtPAkzNupQdseeZIKqIrJM9Uo4LERqYN9vUd/yI52T257ah7fk9A5Y4My1YKM+
CJ0cJQFaL5EajguJtJK8L3KQugQDXMf+sid8Mz+KIaF3+w7f9NZHH4JZ6tjSNJHn
MYriktrIBvkSaripzjys9pWHa1imcOEDsbxUow8CB1htqIovHXDBudKW9tlDkT0z
avroSSfqTB7YgV/ghqLHYbpiPFZN+ujOxlwLTXFO72nKDLPFuKSN29ThYtNAYk7I
X4UvvRpou5nQartdbnQPHFtHq3zMfGSDdxMc4UEBA3TgEFLuXLDQ/znjyLmVaC/N
cuMGnXBUmA9Kt8j7J3Qp7OFE2zotO+UWlmiPhlSjpJLN2kjGP9wicIYw9Txv6C9z
Tqyu0W/7EvDBmHFQzsprKHLZLiEOQUQqhP/fJZNDOvKt/8aE4WSsUjUG7vi3sbDU
26/nnDPAifUa3oemVHHHWQq3ipDqFWshQ55zrP6XWdl1cB55OAyCTvn76hb2IU7K
RzaXxLNi743QxfcXbL4gjwCSvphrU2ZQ1m3jMRk1Pf4dMACD7rAMb6zMjmYqDMt9
KimncnHmTI3dKolVmAj5k37ybpMJEpsl4U8zC2XOzSzfeu7Zv8uj4UMYdFPZDXA0
EcJokzc1QrrFpXkkkNS2upZxthI5ZYYTLLn8sWlyC1IKa4oRQZ+hXWo56SuNG6sV
uNUd25limKvkdBz77kLi34FY6dTPybyIH2xcSqPiBFNCfrESUVdtqmfnSnU909nB
xEcZwn96JBAKe7K69BPiS8FOGjCcKddRZ3G2yrJPWWiRrWq1896qJI4wSQrgE7Gd
ePF/5sDCumNoIUDcYAWai9aTZ8IDVlfps6C9OqMpfE7AQ1h0V/jOB0rTcqAWevx+
0tLjeYURqJcxEknAIlrBMiYlb/Kto5STyRDA8VPQUPp6FHrKRomcOj+7nbU+MX2g
77XUAMtibdNaPK68qxYpUXGQ4LFlB+jybvwF/lVxZrM5ZpsqWad0F96cocUuLVi1
NlygW/Bo/EidggK1iHtySTeDOAbFYkmuX6dkWD9cyQRhpCKlQ3DFn2PUakB0xIfr
W92CSW922V6QOrtbusYOCt3iY6phn6jrAR89eNx8qSDc+DevombCV5q26UpJ3Wq+
WqEv+I//w9nakC1ScuoBQTvB4aeX4L6WDENM+y7n77jV29lE/VcnEJ/ao1ojl7hX
UOsKg3EemIBlqHwACwn7NBF2NcISvtTjkYRZsUhhEuJQHCP7qcuTeYRmClS/evFX
T/HzwkFdIUlYmkPSmTThMUmakX5xcDmblgpaeqJHLTC7cBfehhQEwvUWeuZoC+5t
VzJSuPpTG+VrL2EHEHNpNCpq4FCLWnwWAtoIWQ5AueQPqj1bB32p3x5Xe5rs9Yds
MB3eYBD/qC7HX/5In/8J1zMOYLn6IzxjIx+MXw+Qw1GpzJte/2WV6D034C5VnKif
mwCLox7ZPotSCY/ZdteVNkH3V04awSaXoP0yKtehMW+TcVTRAJZFuUivPU2zwAIb
riOJNLGWixu7rfxpkl/TcVuWBTpJYKJJxeNeNdEzm9JYYww/D8fK8//imnDpHlYZ
SodzHO+hlkqcpKtnDC+nJAX6tkgwo8fYLCOaMBrfd8rJhcN23lEluOzgMBmwMCPD
k1krlsfsr76NymD0YHATR9Qfc1DkFjpwvB17I/3a8BUAG2L/neTSrc3K617T4uNR
dbv+ZVgmOnRj83KLZze5tyx4V3+fGhOCGe0sMx48byJ/1EyarWP+sKwTLbfO/nO/
WcGH89HeFmNVYnrRGAOPyOqB6aCb9ROpWNWv4U9Nhz5FZ0xtBcE9d0lkY8CWidDH
FTU7Sp5DROfqdJNksFCmy5WcCPJXELfT3du1jAd/AkeR257z7qCnCKOw2bTQ/Rgv
Uk7XzKuomsyc1q3s1OJZywRrsLeq58xPwbRMxIB7l0fpTWR0Wef6v0yVMarb5Hwo
lsOFNZIRLjpAfHYYC8IO7e0oqq3+Z7ooJmFAFDfETR5rZW+th1Jzp9UW3pLA5CtA
/9CnNmRvprbu4OBM7tg3q2uYuQrvsBZDKGnsjM0BKExAbSIyaDg6PTTfS/tduHRA
40bQbeCsPnmICnljA6DmtZr1kZ9kJFJPhwaDH4ouKN5TaBxyWAlkZMYE6RmkVarv
zoSVPcP5ibQe4SufA+jx66kM/MCDqbsVPH10b3vK/jz2Lbpy7fFR+waqOk8Fn9NB
gEXzR+Aw0bxqkAMM97amV+F9aSSzXGeUp1hStNl/lNzZ/QksAtx2giCpGYAMW9En
KtnnUXpTBiapneLmzHlBrsjoTxjwbHx9v9Ozk0vUwXDoYOVZ6WKOXfzVjBKSYYOW
LYszNLyp2SS9YAgzQHYNZKN+k3goxBUGOxDOtYZV5Klgk0Tm+CPfnmN4DLB0zsj5
WKNcoesoW05w1MUVvY+YCW9WOu8EZAdJNmNNDrHsZxROqQA/0il0p4e8NrG7NtAD
aWTj/0AvMUxKpFFzU6I8a508PmM1p9+otxg3OJj24UsIFmnRPv5dd7ZncNNngFd5
5HBRNnDTXynMEjgiGk4DUMKZPXwZ+SHbBwUGJsXKNXaXbAXX7b9vUHmbdbHjV99q
qvtzYuJbmrV5/j9uOEGktqiMg+dNFJZywpIM6UjQCqUj9exNM1ABDfexqD+4qM1i
H5nYWbddyBTEYGnTsHRof+6qZqc9I8BfwePE3cuLKVrUNpIfjy1pBJHgpXxLnqWe
u9KUn3jR71vGtUZPYTfWWLeL/U0kc6iC6myGEb1NTh8zgbGDsARO8J5wMp/2mtkt
bbsNJJfJvQo8LIuhyG4A+nAttARmTfqqdQOfniXsKNLIBBjBFY1q0YG7IlM8ULXZ
0MSa25w0TfcEsgOVvbmwKV9Gpb4m0ICpwiC3ukXTMfUsOMtHTHQ4cnl8+toEKWxN
RozmBzj3ZUeQAaxoGvummBzpSoEa3OyYjCRRmMsD9h9diKbur4pJy1rguJQrhFFd
DYGSoaPxOytMS3zGkmVvuh0VATrvkK/fFsVtzKF8iMkfHZw1cxWvQykW5oGAwBSs
kQ1U0fYj6RXVyQlTA6mf3uBY0qxX8ciyalnOIGPTandiikmJGG9VKa1kxSLIWPeN
EpV09fyK9IgD45wK+91JtjTPaWsLHZv+WWV8M+coKzSg7morjpSouMnBJ16iahsJ
mElJtaURgd0MyaiR1gXJFKfZgLziM5VBWrUx1tdJ1lriyVoJNTqhV7Vg0loTVE2Y
W2dkYZZhOhHrLiKcqKYJmkMSJmWx1fwglXf+W4kxBGxxdjHQvc15K7EeOJtHT48T
qmOBuNLqSYY8gpsSK4UGiIIIg2HdEkx5fJ3Fg9m94M7T1oy7qoqKDURgrMliKaTF
pgJn/4n08nHUcn1NHzGitvqWMKj535Zi5Yc/oZwHgbUDQVfKt6Ki3V6ZxPiKFXty
ie/s5W/TjIOgXQoLrDgkUxmTpivOPXupkn2BpfYOHP3ptQ4QY6CymH6jgLMyueP8
0sOkEeyu2osE209a032dhS7VhQtHwE93ymvL4XEajcjpK26TaKSOjxEiuKtCGbbz
AuuvyLCQ5bnUPBnwVQGEhkETulOOyniLnYIXtelhNiz+YPPkabxq7+B+s+rmOHb7
NkfYZ2B68oqntmc0qGKUTesxJqf5lqwgQKW/wxur+4PszsNlXUzdJAFVc9hszfV8
yZmm0L8Mh0s6nFtDSakviqvs6QJOn9yCUNFiFx+hdII9ySUGwecvbz5Vtru4eJMH
2k4OS41Mk2tTCw6OxiBsSHvG7vl08+GyxiQptqY5WlnsXhQm9S97SyRzpCQ7BrH3
yra7He4WEPLQp9E8NdXdZ1Tqo5z1DKQje9l0Lp+nrKPtNffsm1CczUxeV9TsiYXj
MubZPbWxrHkTMrhzfy0iWqQZxG21Dj5gfZlCJLBusHKSAoeVHKq0lma3h/KE/Mik
jKMI1NrHGzzBa76R/jNVwrob/gevCJz8E989SRQuX9Su+e3pv2x78behsh1y+OaX
bEJLTvLUb3egPaA8ytuYMGYCszsebYeE8c4tbp/w5Wql7pA10GfZ4biBHGqxZdLk
ePnqIIuD6NvQToocs4F+Ht8ce6VR+iGP62yiF4aGxXnrAWD9kFkIpD1EYtw5ISxH
o2+/ZriWEr37sIg6Bp9K7jjoU2DRt0efq20YSJxldyhOBO4jU2/tVbSbR3eFs7gX
/I/PWdcmjXtmz0dsv3KYDa8T5OYCY4W8994o3aZI/2zznUaaaP3HmpLOz7dGvc4b
/N8eRi+GmjOcj+TdmbYZYArDOpUJ5r7KW7bI8S6VlOTpyMwSOd6+K0lwIffFhMxj
+SpqD8vfImGtOF/CVHVXhUjTjZV+Jo2lgigQX/2VorwTScUufF+pg65w/vqmo61U
B4+k3REoLkYHUNC3OKfTU0t+wg9YEp3kgYM8NFXX2uA9Nj6zb3BvCa8gTf5Pb+bN
rQq9alr+QVnX+VaYwvT0Eu1ngC+3CEjlIFp6MR+XLl+/bf7gEaCHeHbYoxwGOKpE
ZYFVFZaWTRshu4sCs6zlsS2QwPltd53xUm2G2+VzFk6j60iOP5+Lo6Zp9V1HXPNL
e1cPHSq0yCrSIPCv7u9D8mJMnEymkCF3IAFoHAzWkyXGK6Dei2UgVZdlgbxlmuXH
+Z5dco8tRCXTCeSIcV2rfEFSmNQqAeUVdYzzgzrg0z2+9XQ4NvlNFtBSfD4OKL4m
XANTMQ1NfXsMOMydGteuoQ7XQRngZ88oUMzMkPZJsG/oYfGP+bwgvmy3UbWHrRD1
SUf3BHse4/QbEsJwFeWtbGpyQnTPr70zkP7ZWbDYsXQewqy9mIpGBM5Pj5JyeNvm
rxXTzg85wCkK5bK/20oqfzhvveIMIRxTOSre6BVANCFHDeYngskB/r94D4Jdir0P
svh773rgSBPCGGXm6MbY++yGWfrD7B0IxHXt17kdVywB7oBGP+YCh3IkA9h8wlI6
0UoE/Kw1wsTGcgoMg0aMyAwDDaw23TUKgu8QR6RV/4BCFbTG6TauH7YZIkM3bZRT
k2RA4Wz0to5uq8vwr+840r1PxnWRT5LH/OVDQq1tXRPtNWte7HVgXK96XOU7MBKL
lNin1r4qqYSBQ4ZJMUZJtFTg4ir+fk1nFsE+kfJhXeWtuAGhGHnRAJ3oFMtHPvdR
QB9JgAWb42amGuosxOsD52EXH/TVefOHA5bKQUqTOPQ+LBNEgdWgK6xIUvnkDrSm
Sl8/iWE1MTT8+1pF31fTd53rErHTsBry0NbrIeV01+96p4QQ1gEk4ma7KLJO3Boj
wndiQIuTJEajwA9wqby++lVmkitbTUZt7lQNGZ0PlpZoIw3nVf4Bymwr2HclyWdL
nKFqx5cHPBHeCQs965UH8ao0WnLSYI2Cm6MSJZCKsTXF8GapUHlYNohvH3zUlRih
9rnl4LqSxbbo1hgdiuQGKfX6LtWJn86N8r46kmet2YWuqeIWp2iUETZ7405NZ2gJ
Ns6ppmcsrDRYOZR6AMzwCISWaXHl5ix2U+NgNd3FVHIxMnfJW8Pv/o1MuZ4ElWSJ
9Klsf/mn71pkoif9O56lExIzC3uLZ6ar2VTlIHCcH05oO58OnCNL3kL2ceCeJkAU
jH/s/80dGRxij3q8I8/I6/AJYSP3JyIOKtWQlJ2jbV9N7uzDsGc22/e+rfb2pJfk
p4ASnr8YzFrrF6tS0/p1ztcwuyjmxos27PvsaDVD9wAWdIftQgouW1xlGlBuN5ZQ
pt+zEmocXA4QBEWlWlEVqBanGqEmtkHZRm9Yy8GnRRtzO14zcfYSjdxwegC6nnIh
6faP0G73lt5OhQ4O1RzlqZ81NyHB4XB8yGCytS18DkID9yz5HdOEXq0T6wpEyLd2
qXXxMvlWhSSI5ZiyJnjR/dps9176COdxsuh61wE7MQkhoXoPeeRApqHx+qe84EZY
2SscLIst97U9EN8mHPp6Z9aMkAgJ6XV53f9qhgmzEEzflnSuQmGYwcToQPrpVz6Q
Rck4LaPiH8b0IbycP5XkzGQXpvHtqF3zw9aRkXkLAMd7DeQMZ01w67zgdtr4nLZg
rwqFkRj4rTxLyqLEMQ7Monu8ZqlV7aJ2kddMwc5UKT8mGzloAkS4e2ytRmmP0TzJ
aA17VCXmiTRwZO+CFFElHRirNAKPowQgMgCf20dnvnhfKLIfBBg3VjFk7YRhd/Ed
Zvbx/w+Hlb3FWuWWLL9xD65IXoTJoUhSUhJcTW9qPY59hiJjqDwZM+Ujdeva2EC1
BdsspFp8dBv/fHWRs61coowWRvFaWhQ6R2qeqqrtBwZ3oh8+HmT0ipl8M8FQBLWI
n9EurCeNEDbA6wkmbqrXsUTIOASQaG6MsfG20QxNtNr8EjOb8t8HAeFewlOSwzRD
BfsYkN/3hoEWYKBBcneAzCvYAq/br5LBCYa3Y6Ok+U8oMOrBVO2vEJlAL5uH2rHs
Io2ZTjCRF4appAmTzqWq+vxlx8M/rP8gXJl+ae9wkzBud7GCuWYy+m3U/MoDJtzX
5VzuJwDvoVGOnHvtNgwQuQkpXlqlgg6EDAYTrCxljFwwaj/rXIymDxI+B+8uGKAa
ikmRFIfbwAC/5j/dhvmBZAu4kg/WLvNRVQZ6KBLil4ucj+c++kJG8q3+IfcioZoz
J3lHRKj1Z4lmP1bPHZ0Uo1x42XiicZlhe+fHWDnlQjySpohSKqJ4owz+oZc1mcwl
4CPuFZbaYnLVxOqXLoBJ3ouRkji3olpiUBW0PNfbvGen2RWoV8dAwLqlALAKT4pv
vg4ibuCHHuPxcpEv4YHttEq6wDnXCSkzLLNEaDdfVY8IVu0BVWtKrNgiRF8523SY
H2eqOoQnb3/fGGEuUUqZR1CGftkoL42C99RX8vsr2Vk8fvh1cNodevqMnWJggGQQ
Q2Q3D8TiVMujQhlWZyPj4HNHmPEvJI2LVq+MqQipsTpHXB8IY9rZGtDb1ZQzVVYb
SwOigF+t+7wHFfQ/ZVeSyWjUpLENTQAMxKQwDA4XdzgPYOQu+uRSQgyjGWAs/6lM
pjV5pfKcOZQ+USqj6vWjXAlMumHTtHv2vh/dTjct4Q7957fqyW94If+P/rt2PIYT
1A1jZG5/UGyeBhp9+2j0z1IfY3rcqC4bthoGxU4fQvi8QF3epgHNGZ6KLxqCP0hE
5AuPYY8aiYie1/rF2qskaRW085R6behMq2TvYIjUks/bXVlbZQzWu5sN9W2vRwbT
m6PACban+QQnNAoJ/02ijvNmt9rh+cobBS8kgd14WtrAz6b0Rx3FqkkwzZ1pTBQN
3qLPZrWpIbWniBwVwwAPEatgfU3e6fh/tfZ3R8dNLAV73FxdPE1XT0wQ/+TpP2Db
3i4oP1I6kX2P8hYWU449Pc7/KyXmAHpgLEE4+sAtxjy5fqgqaFnehJUc8CkWCaED
/kVmhxb3x+GbhteYqLM1Rhk8Fyz7+631mRUTWGj/RGys7mQFaFq3n/kUfQtcG7zV
WUfFvCqtSlDytkKSq62US1qPEMY0/AFlZ9A7d7s3YQwZxBiO7bClK6ktVPFDjOkk
AV1Gx9d5+4AdbomZKUJ009xArHnzW8zO+COO9eiGO2wEvVQrWVfU1VcVkbxzBxs8
ONT87NMoZx+CqNkQ32rMPGv2WVlg756Eu2IOYns7Ocg7//1m7NYpOXpD9AeVyNgp
K8KrXxf3Gy8NV4hBbgCYzFTJDWAycNLkqwXTG7ni0UxEh/u6Jdp9yxGdHuWs2eL1
q/V6YrI1jEeyDt6LBc0u7xL4WrSQ+y3FRRTgI6qc5tqRFK8Cy1ZwF+YMY7gYgGSN
ett5EKX2g3NVI+heN2Ifc2xmDE9IUxUYDKcqorRNV/mgQ/15ZegivBSI0Avp1ItA
iXpz3VK3Aw1nDQfHlgp7m6JSDxJs4yAHy95neu8yzSJf9T5fhtecb1dbjteQSMFN
WKAhxM2puBY8BEWGDWcsCi5B6mDk3B+BTzmhan7TON8IfA7ZFlR7Enh65zjyAxn2
aKDT+ERbXULP8yZt7OngHAk2VY0d6aDDlXonM3S25iUc2qQgmZ86EaAiI1c773hS
e71GsGf8WLx3CVywGjOSb0+VcxO+Jjq/6BjYQ5QfO4BYl999wuwJigesA76nfrVm
KUIEEPMrgqCDRoxZtCqB5Kx81PzDdqeMDbLux3V4jfXaoUtA2brozSuyBfJbJ98s
sCI6ooWyRsXpUZ7QWL3L/dTOc7tbgLQe2E+t0/m/n8Tdqqyef1XXJ4pJWVAA1a8s
6N/hEdijvnzhj+XvUWfHryUHaOiFx/EvNEJ2sue2T81rImFZsTDUpHujs00dVY8x
lzUsWkm5SZCgz+IRG1qyCBBJ33zyWvyL41vMJjEw4B2aSKGaSH5Ab1YS849wYg5V
yBFdF/WE4H3gRxs4XDsBC8CMVsJHI6GLA94sNLIlvu4FkJmawqmP/WHM7Z9bHnSc
rDTyozNwR9rMG+Cj19JRKPYt8kYDwp76ZDBhnfOGlEsSkj30V5CGEN2hS2RdMj3N
xSNQjC//Lq+JO+g9TOTHw21G0j/epWjNMt+TAHqci35Xd7kDSUs61p3JT7pPxQ7F
Q/TN4zn+DxyFhC0BZG2DBKVAMHY8u45e+6qo1WcEla5GZsll1Fhp635RvH5lJ603
UkVmwFbquOfCDW6x8q8PA9cxNnAmjas/mnXkSAAZ7mnO8s7bGaLlzrF7YGcV0HAP
a54mt23mz/wIRfI9Mk9ilDE63kibjWK58rjnraPVaCGjqHcIffcsqC6p3ytqMicR
0bTT3fEwK1/RxLzFlyYXqyGx3jTNq9q1KKlIh1zMCFmuYo9oteFEMxPYEVEOnFuI
hOQCjThl+yhtJ7hXnRP2HoG0+vxonLEq8opIfeVzX1y7/OoS4w8NCftHs4wwEPzb
oh/Xx1dDHP3FUScA5F2fWaUiI88P0yoGKuaP08WW9S+xXJwoXuoH4RsS0u6pv1Zk
MBAwHbLpI2gBHNJ/CuY4v5dmWdegPq0YexiNXa3BUeCSThPWvylrChynC2e7oTCT
fSkqJU+e+qTvZP/FSBxJOexvPrIThjpI8S07ncT8U1pU/H5VRphNwdiHDZRz2TsU
cpQ6gblfthR2c+QJhSPhxDdJbVakTx/7fBQ16/98Y42utCtqZVmCqZQysbl5yhjN
27LFS3hN1XjrcU6sAW1u7VZfFgN/A76fbUGiKbrxgvKoQvIxFRAF41NpPhN6c6UV
R4lWovuEq0wyITJ2OFEkg6ji1zENsYpqq6E4wvviSsxH7VyviA1YXycVu80VdCm9
ntggQ1fMW8WReWqQ43l8hIffqvwBFt7LPPohOva+xIvUjGG9R6yI+F4KCXQhImkn
1BA5LRhG+teWOUyBS0sJq3hr5ZwF2fI58XA3CO09jLzjl6g6AUpkz779USSS3fKA
/ZhgQefxsftnSn3FNKcPRIPEZ1hlmNmadcUEuuo1JaV7YKf5GsND5hS7Bf4EArvB
DBaqWqf3Zfo8eOr4MKPmL0MulTmfaIXTGzEkkvzdTTILkhoyjtJGrgXglAxurFIx
Q840a58jd1ZLtNYrYxJcdIYvCDOjWHCxza2QOWH/6HZGVr3u1Otj7CnZ5K/hT1Cw
0tOaEzpJvcIdC3U9CaqOVa2Cgg527CzrwHnU2ZE6H8zOT4LOBpN1TcfUE2HMtSni
/+QvTEJo5k4enEBj9TMC85z8a0xkHvA9bq9Y+Uy13NAFq4Pk+KCeLr/CE9bFdn7/
REGyoAFI6eV0RYT6Q5TEJK5kowqyjENDDYcI3YDovcIwG5oJlsZ1/0OeYwk6Rgpo
gbVQdxYvSO3Jiw1pyjRwFTb2NDCUMH0an6ACSB3HdCfBiiOddEmzjowBeYUo161u
7gFyMMua22otn0KOzxQDj6zngl6kbRf6kPXuzQ+dSaf/aX/AABDptKO66A1j2Fse
zXV7c5nU800LLrpbwMWVIeYXwD99SjcxkHrsZaTLmcn0PkscGIdZDebbB/LAROIN
Qzaq1lVnY+Tcw78yMXeTia739NIV0DKeeEDF2iaBXijRDyumljhCNkWebSbrPam4
AYnZkVHOlSxlurXdwziTTf1XliRzddbJ1voOvEUPPj+hbXo1nc1dWcgFXCtSYvca
vC0CI0oHK9l6VgUr3CwkwC6YZJcom2zm6tcPR06FOAJDEUp4peytIkPb7XWWI+vK
Smtt+8NTbZZlR6FMaOPmNYY75k+7/JccncymTkZiL/sG1HrEsVrUf5KfT7Y/dQDg
zohMdqQ6+5oRvgZfOI6jt2Dbt5Xp8YaftgBC1o3vUzkbGTYbTxQNrXkf4C/jQwz9
Y9PxsORFns55lc75Bf3vwCMO14rDRJM7cxiLXJFRyTeKC4IEqeSldGFArz7AunRg
VhaMctFmSRG6C7ZmHGiA6a5oscKYWS+9L3Zy3ZR261XBzuwTvxFJoPgRgyYUndsp
6cEJWlI1+9382MV6aqQS1n95pf7pNBHTyFsYBed9pk9pEsKI0nx6Joqrr7/7R0OG
zF7pyzlSJPqoPqRTQBFkyqswJut5O8xzmAoofvfLM8/Ge7x+fDeTz0Lahyshcz3c
1JqqT23HGZBbAWnXPHHLOc1MTbgm5P+YFn3acR+9Rkhvdpl4fDHaR+IaCd2o1tB2
kqO1cm34e6JVB3l8/a6KJrodwxxGVPzMgOPViqTV187ZNa0W9Eki6K6R/jrLeWMH
S5ho8RXqUYpgqfbt36fkr8F+duhLTf1dhypzhpnIdhDa9RmBpVu4UmaAHFq2OUYH
rqmnTab2uKGOt/tRE3vXQx44yg92nHefjHZX/6lh7FEcdLtrsYpCohJNCgkguByz
n59TZESrXJfKtlbwLDKFT8O5KGP6Ty4Voiamg37SRJl4gUKzhCdxr1FVzeRpTtwJ
aMgwUS1txw3h8Vav4V8ZRSQaF2WcsBSct6XYTEYOxm/fs1zf1ywHVpBS8XM+jK8k
wNekHWSDHLVjqpo/DHKlH9cnOrYcJm/AYklZrZTSrtnJ+TCipNTlFn93YgZHXaJ5
HipBMRpo3t2FNB8ax2QgydKLa6IcQSOgCyd2ISIIZtK9DBM9PKi9xTxdfWRTAYIc
1gEgRtnxmvJFCadJtc7sJ81PBor7ggWf2k29UXFyT2cSMBaCPEF0/KGv0fkwyh0U
UTdIek/GLAQ9m3gzMELVdrNg3WH5qz9Pep3EqBrxapvo6r+nhecKdxpnwW9fnIrd
SYu7se9hfYHP5zjxZL/iza62CORk500sctuwVR9SUvP1pIe20Mij2Ddrj0vK9aHB
unLf+JMqDt7N8IIcnvMKAro6qGLSBC7Xx8PrHk91MN6ycu3oZ0vhFNr4bJEil3qJ
Csklwqx0IYFSa8ZGrjo1UrR6T8E52UF7fgurwHniHp5upUl6Ivbj5O5/yeKAZ4nm
ul/MZLtMub0V0gkW4Np9e/mWK+Nv57zdgUg9P4puvb5XSD7i31lW/zvbCiRdi1Ut
kRKntvUfVDGd/xXmpUHwOZgr4Gl6oEt1+qjXxUVICtZH9DMxGWWo03SnXtMSNXFw
nhU7Z8ZzVIXdArgvwZ2Y8WxcoAiXyWEq+PYmIlES5YRd4oPmPsZn7q6+aQ+gHFP5
ufjIBRsoThTWs/56BW7MOpAyP/BZZst9xmRKy3c70Og7AnL3ZRxK6yuuDNVStPx+
xijGTTbuFMwTpCD8yIPLHYXlDycBA6KaO+qgOL2/q9nTnz4l2GurAiNyjlKAx15W
jsc8QE9ANls5+Hh4aiJkGxEH+XO/WbzT6k/QVYfZLUiVBhgCCLDOl8JIra8z0pqj
PZEel9ntQqaQfgekDucITLJ6BMzKNUFrRM6F0IwviX7lWEMqEAUdlIrNKl18354N
N62rCnDGv8NP7jbyAss3Fp+udrLcqXpMLYuPrE2A7axTWS1zXq+iUibOts4WBXuo
RK+rIyaAertL8cDct1Q1cvCemqv8lLrMRiAWd5OZwtajShG4u57uRp4WnS/2G3bI
TY/rNjeVdpZCInXvz9jZD7OMj0l2uunfr2hIS15A5fV/DSdOkU8nFDpnUlqYqaW3
R4z1wxgUqEsM+jUUk0wbw9ufmtq/f9inWxPlhkhUT12L4OQRticysoPOoxznz4IB
K4elPBAlGd0ZY54yyn4bdXqXNQ3929/bOxbsY77x21KTzcfznhHj+pDxM9xL494b
YUghsNUeJTLqM7mY1ZeiGLokymJusLkaY/SDufGc6EZ5KcNjnRIULObjK4JBSOss
iav1G4lxmg5THpzlKFlQi0IWVDK0k3W/atRt8BvNYzYsYglrgwIZ5yVs/NRgUjkw
kkqjYZgq3J7uxm1Fib3R6OpWFmryGGe2T0jeXLnyZJfT4lLGoulwt86njNbICX/i
DRS680NJ4uJvWVGySXYZMJVbCrsJbnN5CHYksX2+bCN3jdqWMP0jZd5xvtfeB6u9
7Vr4vbERMpxsCZz+al9irU863PwQkH1nVK846TLR0IIlfGwxVXNv7t9Kb3n5Dz9J
YOBMAXmB9eGSD/TaWkGw6mVETZWVW11k71abDo18D6rRDi4tJ9rYIscxFqAKcGRP
n7EVRNT4HP5TtfZ1XvK92SMe7hGSa5IAv3VNfhps7gzzzYmTWV7HZJ8tQEuQoC9J
rdvLCcpk9w/K/OJsr1894UHQmBKcH1TK/fUJ3t9qOLyurHYYMD1frkNMwLvFcm8B
GwnSrVGYmQ4S1rIfEl/SDj/9at8Z4gprlmurtHAmI0o552Men+MPdpyurE33W5yD
AGy0HklROFCBgEww9HsSDh8t2froC27kgDYRqQLDw4RJTU7hOe21+UYFt3E6Yajq
DY8NEl5Sqg22DroSTvVyJjdRdyvTIje1klT5C4u4ZujeM+OTv9B65X8fjqCRfvcr
kpiu6WwktmzADy3x85G+BKDZfvEoDRoM5dfek3fJXf6RKu95lrUd52HjxuCpECve
Ig4iHHoJ/lkGbGBxuiu2irGY5yarFYpFjE2uZFf+32a+3gHJTioyc3xy0DLArPkI
57Ae0R9FWsejpK1XfL78v0ORe+vJYDanPfjEkBuI+3dbYVX7UGmdSAlRGrH0a8U7
Xfs73G3Z3PDZBA2FTGu14mPUtO78gWC00AtQfKJItozP1XKEg87V5dX7VJXGCVbC
i3nrGHAaXLGnsDGB87s52L/2hZ70TOFnWdIG5PsrBp07lr3vu9URo21h2nC1AvoQ
wu7fOuiz+KMaqWu/xCWClgac5vLx0B4//WvOnbixrVrodKxkKZcNjsnN//HJaSXK
Sl0D4Hvc4Qgzvvu1eCQV6WJN6gqkxr6dawX8Qrvz8cMAlnw+CytAeDwDCrKYbaLI
ZezzNFXuYvXhTljSWs5Wo6TmXAIqGGP5nbTp5174/m4SRHWxA4E8zAuaKvjg4bcf
xpPFZ7dqCDp5aZIfWDdPOcfsuIhH+n7eBQ6xxDw+/ZCXZKcXom7FY8Kh8ePwp9F3
WZ9IMaUcGTNgSGQebcCZ8ET7UVru1Q3yexF6yEhHTXapD3tvZBAxtrk4s98RTd5U
MW4MQ7SqhVs2+3LLnd1bw/dJP1oD8YSl7Eh2oLQ5YG9YTh5CWMBpjN0VStxJ8cK1
7RMF5WLzbQPYoJOzepWWTUkuLO0Nat2md68DK0GBOAEFDLPao0W92WLZMdOONCXo
wz7/js3lFiA9wsk7k3/6HYG+6veDwRZPG387P2y6Ztqsxiqqn4zNInSS6BL8eABU
JBfIjGt9l/9G3Zb3XEf01kPZUxsGCRrvqgad8fMGyXjPTCJEGJL4TfU5ueFBopC9
BMw6p11jxCi8ZJ66RjCX6Oj22nkCil16qwo9UUDHPhic2vod6j5uAWIuCNlbbsRm
488H+FPGA+w2pBqceihcFpLm1fUfEQQPNgi5XdXvC5cYl9MtyZ/3YTDp4LCjUcWs
1Ce48uzfp81Uz9EQ3iyI0xzHoI0/Um8Z1SQX3cN5TIwIa4SVtOD2MPNmI4D9tvFp
5J4KXeaSNWbgb/lKDpw3WYaentPWI7a0OrSB5kguF0/FwvDsuhMTBlT8/EgXAZmv
LvRLjvgWhqjsBDr9o8T7+r/ggJCAxoUWRQ/beQWKOku6skM4/r+mE1wQCkiRvvcE
p/v+aulOw6TOgMqlnCf0B06r3HbMb+8utx34eBETloKOwlhQoumGrHeBr43iArDj
UOxQvhKB3GjvKDb8IC03hs4N1bruRPFzx7C15HXvuKvxT+VlNQ1n4728mrtq0F+O
NPhTUDQd1BPQcfJaoxaxqUuHkuFlqqwiSdlX4HmFMxRlcA5QoEYCtIEFiZGqriqh
pvKhSp0WmXYq9zdmeIRU/l0fyyousJTn7yLACOPC/ZZGXwOuwxctFmz78aXbTmLQ
l76ApEwmVWiapU2yx6FilosNKylo2zMn6G9TzmChoIwc3K4P12fHC9CLKUqWiafd
0AvHHYCk3yR14Xi7kSMCxY2EmLBIXM2jqZD5h4OAlPIG1jkwsnypLca9+pLqnayk
aUSDWUTly1wpOVJ4ANUMoBzUIrrX5cYs5Hd+GQwl8hLMTLd1RTJTn4c0lthrtNwR
hhsZxQcd+Jyj0pCKdOT74NXueT2yebTlXHo3EhdCCzwXJRdMfjTbBiMnGSYaub3a
8oE4iYhApSN2fYQM5X6GcalsCuhiX3Z5jNKWRCDlTR0ePS0n0/DE1DsleV/LigLD
T0OvL6+BTuNg1a37zvUSKzWjUSM3vNgVmWYeFke00xprTwD8y4XqYDaE5gNlgDPI
m8ZQcq1E1z6hTIseJD5aGgoOQCbIY0ymlDpCEq1IJ4tGD4zY9qKs30S+fUs5rJ+X
DlyYuImXRB1fs7fSdjlGexzr/J1iU4qdayVEWrgdkWfSWmrnwXdGHZPtS2ObsIuI
5CR4EzE4o2WyJ8QTqgy+Py9Zgtmhi8Eanp75qqiopvnqru2WnpE4GVY44xmzHeWo
tlqyWkpdyDNLMGjaUf2n/DyZAYKfufy3lAtwEnxuZF3XupztwVOdXwuld0M6L/ZG
FCWfQu6/e/IP0UVraOUI6FvewB9sLLs6/mwwKXH3desfyVZQ0TITDmjk4vEqyuAw
O9DSJLvJJgonBAG4ksc7FNTljVAk9YCna0nrUMuWhkn8tSVW1JevXV683ihns/df
vvXiiUwXUJGH6LoQ18x+LntWm5yO9pIl95bxQ/WU2fmKhlBrrE3UHfPdNzxYHy5V
swf1HJAJ8oI9tEyDfR4cOvnowREsY6QedYqf4EZ98d5QmfyPPdV6D3VddQLniNPn
vGzv1rPNHC/7tmsG/8gbB05qolVlmdv8lTYLoTjRJQe+ObD3/rHWCCQzQXw3S/Pc
eZ6VliS2YRbRIgzzmgzKuhgRJKNofPN3kizQ61V0fZ27rMObbfTre+HGD+JjYG+3
cf8VBLK+aO9kl315sjgheDIAfQDe0o4UHYQJ3O9AbFaHqQGGxi3VXMC1bacl/8yP
d7thvBMCb3FstbG7SOS9nnVjVa8meqDnwcCJsf3Oo0bsoJD290nsi6AgZ6NyrDZ0
qEpJ6fEEG8MdEyw5RIVm1Vw4RVm9hf8CrEAM1+5aaTidE0u3jxtp6vC5MUczXltR
0b3NLI7SuVY/AapJ4iaiKUhl/1s80W5rtZfaJ9QHWzHYpHVE2yJ6KKhaYjvQAiqx
kuv1uWvCXwyeHk75tQLIKYDyri7eohsMooV8yFziNTKcCCfzB2S7K65nPYVlQcGw
u32vKtvfvDSYJ2TYBJoJz0p7c3fLITUzFyvt25E8zTqOuZnZl7pFSEeDNIQom6Wc
0fXoaRorUjseba/Ag1Epc/UjX5bIKX0prklkwgNFt4RmioWIf3EOcXAEAjaKUjDH
zHyQ8vfmPbDK6Bl6EcNlbAGb54ozUZRZKNRN4SVQQmLjKu5WrhbqaWY3pmGiW2jK
Y0yVCz2XiyNw7yZLAPeDu5833MeRAlUugOCP0M85MhM05Qw7yKAywyA/Nm0SEMi8
a3ecWt3/RiTA3ZEZOpuK0oUqun7RX+FBNvbkY49KijdrvKr1jLh7R5Hcaal1ghyu
ICzOCUuxfBl+a8i8aiAN+uVhlSxdB6rHJ7dygV30onaFC7SqzX8akNeN4AAemfd8
zNVUqEjkyIlyDTzNKPdZbVHOqPXArgfdvUtzPycOA/+Sfwvq2ovsF4k450WjIZcE
PrZt+xkO5V96Lhzsc0ugqmFBUbWbFxXFTt4ZCo1vsBGith7VEmmhtgFpA0/WHjKx
PrTMqEm0LoxuVlt1yDfDUo+3YPCx9Cj6e0gwq7YyxJdxBE2Bv/4m9Ns0AujJe1ah
1Tre/tuQynt+IHS206PD6QgFMgWnXYBw972W8082W2mFtvG8BekXB+N6MOHKBGO8
957C8ts/sQ01sm8xG4osC0DMz+ij7KdpxOJwu9+z5eBRXFJ0Mm5RpQ+AlkYyCaej
oeTos61MpPOyS2zUpjxUVoCHL0pVcw/OK3nAhBVwx+s0H3X5saAmtOllF7CEc1/Z
kultQ1IYvZdNjTJxSv+Lm8YmUd6/2evu7Yc8rIlEpHX968yDW4DMiirdNFZ+mZDo
mjiCwUKdOHZt8oLbJ/Hih9fzQlmCTumYMde6cytO0ZB2flA1T45Hys8fyUWqEVDT
xPiHI0DaT7bEXaHYe7Le5J1Z5YakUNyw6WkrVRnwVC3g4V+BHZRLbyKwKe6YCqpF
MTOm74Khquogq4EfJdqoeeBjNm8boCTaQhYyN9Z1LWei2lgAZaBOF9UckjxYm8BX
D7rxyRLGCh+N9CgXEyijDWnIJkkk/sIVeDGy9WncJoZF0OUbqY8pUvsLdVlrB8wz
NLQNRDBMa1GboVEF5pRJiI04VLPDf02LEIuhti59lH8XV1qyQkMX8Bao4tLpH/Zp
IJ9mBySbuHXanuLQBJHBG5yFq8lRvHk45OIxSux1j38lL/qHKLphKmIJPH2rDKKx
XyRPvsuS5BaD1Wb/oJnJ+JW3WUUIqi0wHoWFSoJejb1yOKsIhCNI+iJm5yvtdsuo
3fKLVQppRWdJa2Yp5dMIAee0fpSKQkEAwjrEwCXSB/GyXhK4AytaTFSLyWkkKp6E
JV8wHbQJUpJTynpB7lFgn6T/3rfQWJF7bILsOYRUBN3dXm2pN3UxXN+KTnkixNLb
9nnY9JkAogRddt8JKVLslaK3Vt6zQj6RhNarjn6lZP4H1TKoDMveGldIosj8tID/
k1XrgxENdhBh9J7ZwHd9dld3N+0aRughSoaB59xW1DBcjrZ7/DQJdA8q9+TtfJp4
nc9PQDs/jBfGl7hkimBI0f1t0oHFPcdHvVlo7GdhjPrZlf1CKVkoC0x/74vix1M4
RGthClBbA14A/kuoXbD3TYZ2CnqDE1kZTKnCjH+WT3FepOwfns1c4H7FAMrHTD80
8896WdiZ6NPvLb9Ur9YAw8vwQp58h3SiLlIGsrId11WeN2e+sclWSEBKm8x4updt
qEQdcjVxiUfRlAqTEIwEld66DlfJOyyaTBYLoLwrXs6q3M/hmKZcY1o1UwoU50zB
+K1lqE6A18jtzuuTLRlBwVLJH4YmyY4WnkeHLJXzIDzDZTC5c99Itym5UOzZ0Gom
XvI54sfHQZ73VSjq/izEVqTPC2+5WQZLNxZzY7doCX+uQbMwRSlU0KZtjo99ukcV
ULasfJTPDleHdAcyLtqILd4X5SFaC1Wuy8ytlZz2uI+/SvX0/CJ5dqkZ5hmEcSiv
FHoykKSiqBM6NCN4V28k5nQ2fUWaz1NDKOJX+oh9H8Ieg1BZBjzczTBtrE19qDdB
vbcF2xkt7BiUGAkitibO/YjP2KXbQh0zBwCjDGvwZjZWfOa2qjfWN4gUSgXTLMog
X+5dIWfE51a9j1cYw2yT/IkOYet0ceK1bQbc+XhMlLEa0CNAOqvmrCYVdgcJMwYJ
W7seTIY/S9SOeO3CjS7V0CDVkb8Tg/hFKjvRdha8J0cDCCE0qCiraU2ntD741RUE
NdJFEiV/J5+J2Y1SlgO3JfyDI+8YM6guxaClKqwG8aFN87bh8MU8NO/JsEcc6V+l
htZkMkVqmkZIUaaB056DtkFDfcGCpQJ3M4Ydh8WogbF3ua2WyAGEaoMqjBuTaiqk
DGE1jInscgaiF1tVNlGD3KLcn7wvFwpMBfRGqIygusPA+mDDWAf6U8UVK+Oj6CqA
RPNT3FCEyxe81yY4LrLhgyMXKsG+lbQTXUpPUfiyhwOPgRePG7CiGfTHO5MOBONe
ZOMxQlzuc5enDRLJxbsdkv3hFGVCpgGrbd1W8b5rVe83IfdsVRHG8QC4fH6lXakO
zP90nM3EWlWCBPJAkjkF92xnNPaRwKtB96RHUHTquQ+kZQQZzJpKTWEHX9U4tUVL
f7ZOLaie2+4lT0o+jLt0rLSr489Ga1+dvFG+DN5a8BAxq9yngZO1XQCUvMiMvr4G
wvaw83me85DcHGCx1FRoB9LOMrP88/suC2sgW9u767UsVdMhCLKtAqT0XcvlCHFj
ilTgHvZkDjIdXoovXz6/Yor2lpWEVCTQl7NjnkArEe2n5hnzEskDKPJKSjISWaQT
iBKEnXf4FvEz4yyvcMbM272eacort0bgYF/ppg+p6QS94XaTL4+XUVvMsw4/9KPO
RQzxCAgG5jnDlFDltkIzmtrjAp9oteONRr/eYek/AEygkrWowwuTKFWOm3Dlxck6
7kEyCQ1Lva3PyXzyE4xaPu8Xe5KxFhc0Klr287wQsPu00D68ownaaFT+mTukAoX1
NYRsd7XyfqWBgTDK2vrH4qrzozfF4HKo8aNXD4lohedyZLGDZ1OrzffwduarmFbT
ZQ5LdGRqula+FpixKqAtva4/NYhd3FuTifbRkicRitMAjbxO1GLXRIzRS5acubRl
ts/vEoq/2k0KZFCO3aoCy6NJJsD/zPNVvb5sk/oOILwKpv4WC4jPHQlqoxOk+xUf
3n8nI1lemzzYuvnsXwpePJScPX0Iqw/feao+d2SjLWlFQjuv5YqNG0no/LsuflQx
o4V0kxl74Ub8jgQHbX2rtUT6/BH7GMPKSey33lVBD1WTUS41MCZQba5AhPye1VCh
OEJn7Z3LptB8L6rNlGBtpLwv18ZejZt2fUaGUttVlMViKgsaluf3WSgYzqCOhN/o
ZPrY8Ltuqu6tQT3QFdcC75R2CEewrKkh8cizMprL8zj6POquo9JwTikPIAwOimN1
zwyY6fKb9byKNYSrCt1Nsxj1l5RzztEdORTY/IaW3GUTtWujBxRefHSugqeCnxaQ
odq3sGi1UJzvEV5o6JIz0gel1hgF6g2N1tGNA9OJ1kS8BpV+1GIP52n+Tk8o570H
T9lSOfVg6IuMkexSvvsxdcfenZZjrTr/T2AbXXbyXJTsBTzUQtSfkrLQGveSsSXo
FK8rgy/Y1BZyu+1IQcviTUWXGBMsUnIWR4WkQovX1NenkeQCHaXoFzFqEVZt+m1L
bfqdz1NpHbS+syxtu5k7u0DyXTHisGGUEkGLbNMREVFHevj/36mcm2spRtKSjOxa
aZTU8yo1RhyaCx2Ex4OgibkfvLLHsNAQyHBaU4ndckBGW/tBvKzfqCg8SE+q2F+0
x1Wgy0cWxgJJDaZQf6rX7/8bv35UdA/+GE7QMqQbhcmwNdofamGI/u6Is0z+ckos
Qew6VNisuJhVLkmf/iJfOP8cen+K+eg63s6mViSU5MRESE8sfDP4p7KUP1vlwROL
ojLxoEToK4GXhsuCmlguQJp7NW3x3vhuv1Kc4F/FqJy/tesvYrmbZnIrL3gUTv7T
wZSIc+frIOiVhKXdSewNQ4tUrQWYk8fNmzJZWgSHhbrWeJo3f0mT2PZi+eNGdVv2
8hKTIe9QencInxwr+EuH25ULPIcvdFZMPC8k2dLKF60lReUnwPbAIkMUGyNcQANW
rV3Ktv7fuJmNcJlYDVYkVKuEcQOQh9gLG5fgC95nlR3QCWCzsuiw2X/nRbjwtSye
0j08tUEuAdZOEmINhzIL6jpV1S1rkxHkZYxz0ANd0jQtRn8YfD27RAwib8k4dURX
pZFEGDAyZGq13UGOlQ8zWPpA/UrZB8N5bZ9to1dIzwrXCFt2jDUZd59/f9kKCVsG
8gJTWrN8aRB+45kySixZQN/pYoGZr9flzXUa7U86G9D7CEgiMaWBDGy1kdXiR76x
dwpj69QXmTqZVqgX1QanoQYrkhfl0ezizuet/s/mZbmvwSRJ/6wYNlxBe9+4L+Rs
kNmiPREY6sjfSfMfnGDqaYEa8OpRbjGbGSbYaUfCGO8EVbrYL2Udqoyp7LBOR6tM
oPp/koi3MqZXKydzXd9gWEBFjexXRUmNCtegpWOA+rJqYb3t9hzP1RkmZPcNICm3
gDxxvPdpHhyE+t6rKFOd1UxVBqoWUqOO+f6zdqKssSNd4qUwFbrWFXThFnbHWvk0
h0pOX7UXGh/z6Fhf+fvr43kUMMhJ94Kp3A0Xa7VLZ3i/qARzdxKGK01OnMOcD+v3
Moqu+obEuNlImNKxWtrTt17odXXpJ/35JkhuLSOsn1AeQjsJNaNV38a4WDTKsqdJ
zPrzgCRCfIel2JEhiRdtkzZEntL5rPPdTz/dGilKvpOWdBdSKlU+hY5WX34HllIX
Ts0CD5c0BELt6cm6z2oL2yzpKW5RhhkNuhHHyYxp7674oRo9rbbyLILbXj1MsWhD
VMZRGz8G91xAF9HHC6luuHzBZh9RMp6ECJAQmmRI2GzoQoAZHvKWfDRhb5A3D18H
gWYCOzJwfTAvRSnr5X7EonYuWqvtEt4Z3wcvfNnOhx0+PvZxx7tYUFvlxlLv181d
kTUr9WxFUKDIP6nLFVyetm7TK46h0xQCejeOE9N0FWANvYWJVVmNb/YpTU+vuFaW
wIZL9aVHsUQm3zUJLl4zKyXPgPAjskUzAgvoiYa+Ksf7DP/a5B/+Loi1AavO4Os0
pMVjky8M8bdoYf66UKIOMYFAL9ua2CgUTRtGV88rI2v9qtmR9tZ0yqCcnir84B9E
Zln/W7pWGHmFKGHo5y5IrTQnplX/22QL9AEIGAiu/ntO52uzqx+Wm41D6PCasq2/
jAi+k/N2GKSczNreZO38IgwbVXh3GhkrxPDU5nEKAA1+7yxqnOlb8v9hG29fuKKG
KY2wdAGH17p2tI5Z3YDMfK4aES0u5010glIg6MZubprvhE2QQPBgppNtniM+0rf7
y2xeZ4lvQBn0pkJt7ruQyR0ZBC5AQYNuJQEGXzU9XG0AVamJfykNfruLHQg1XO/W
bY5B+r2DbaI5rSYYynwusyANdDrWZk0ONCWzC4cmPpVu5dm+f42IbOWGqg5giqi1
JnUaVbRwUUEjcToETJbYL57hcNfpdR3bPswTtVKXO50vrCCpw/r59j4GSig6SD7f
+nuGj8RCJyCKtVHH2cLvr38vwEPLdhXoi65RnLZOs4aclEw+Qeqhq4GUpTfvRqXb
4Uzex+lR3ztiudTDAGkeZy56uL8KavaD9YKeHGva4Bfd0SpiQNXlM4GvUzUClSCn
DDGN4jGWqABIclneAPj1/h+jUC90/4EVcZHDeQ6tvH7vg7ObcYhtUqhzziQ+leGl
0v1xvfOjGaxC0jMgBwVcsnwg7+fBBDWOPdWTWmuSb1R7jQC9Ddr4eQYUEIeYwPmR
6pGUD5lfPbeaIzP50MzXEl5I2du0W6508L54D2uruxh3iydkzWpdD6DQJid3Mj6F
PPnMf4+6O7NSMypWDZp/0vEzdwFkjmLMGLj4zf2pX0kE8LnselM1C1uFaY/NYF3c
DE88czL8t4+dxeDXls9facN4XHPl9pQI4YKDXfsBIYNtC3zE/VpbQLTS43TwaXaU
eTCQrynKW5B3hQaEWWWaLI1iYNhluPsoi8ZRGZA6DgS0ZQVtoyEmqm3bDl17AlZy
n/oBpwrYxuYbWeqB/3u5GLfLyWHoYDZwQksG2RRVmLkfrMtznhH4M21JYxEWK4eh
XNIdz1rlRAeskAvjhJp4wy+2ViSJTYqhHDLGvkxuz0wjqkv4Kn4nBAnjHcWw8lAi
dEPk2dBpfhlDOvn/5h0oT8XI/Db8pYWDVbSw88KGeuwrnHz6uC5xu/RyY+26f+Xh
soxKBRTl7kG/PiNzucgIaIp5M89ki7Ptlt2WmKHNd5fdBrZABRc7f8eYFGkyLGma
897PDDcTCDkwq4yYTxsYhgUsg9PL4ph98+wT3shDtr5bcu27xoyv+McMK8O10s/m
BBIMa+RapM6o8VxAJghAMG1KhcoEgFzLWnZaP/exvNnCL884ynow5HoIOgxBRs6W
F8WH16qnBGO3Qa59YqSLkfPtqwgk9nY0OqdJfraJsHwW1goO9Lw0ZC9NcbSL6g3o
sn2QwLsnQBSqFR+DoaUyACGBNzqAH7e7/oY3wJldOPRYIPN7i9TFRcIfvJLrXUyv
2sj8+guoBcMT5ULOiT8Dpe1PoxUK97rGVRSOIh+S62X2SLgBuX5le9NEDvm30Yjd
LLfh5TGV+qBb+JRNmiDzNj+v8aPF8lBk8SWm24HbHMG5qnhfNE9sijFXzVX9XcRG
rS7xg69fxah8PPPXR59gzw/Fc09ODEVcw8RMbIIOx+QAUo1/aoqDnhCMIzWARen8
UAp8ABV3B5/MmlRCGn9k8LegUUQt6Zl6HxEQ+6RIWNnRUOABVW7S01FXxFohyCmh
JQ1sXz4Rx2xH4gTRj6R/zny1NdhQ5NWaxhUCuMtNsIWl+5iPampQtT7eGMPhIRRC
EFVRn4KPj3/kbwO1UGFu+Suysx6buQXHnP0aj4EqkZuyJM8Ena8G8rSApJd8Qq9u
fS6HRsN7lNK1XJpOtYn3QiARr7Na9fOyUd9lVzK5k08SMfZti6MIMsq3qobx+xWa
42sNV/4RzMRJu4X6z7zL3YVBgASI/7zqie7mMXSvyRtyL8Rz6IXm26BuhtNc9i0c
vDw0agS+ZWcGivQcnTBBY8MBNmOZkMwthZc/6NNsLZQJUKFKRZVgyCWI+iQRMYH2
K/eDsoowY3y4+Q2O4Xhyb2C/kBz7qrcYaq8hN0x3tz1J0+HUBCLDgHsAu/uFg7yB
5cIEpH9N9wimGLWNmjjDCjOHAstsSgqgr1lsRmhXSGucU+Cnrp1JkCesre+V7A9A
eswEmPbhuq9krRoooNl8INi3HUW/hF/IsX+sRw0b4ULZ09bi4Z6e56Z8XtoRyV7z
rt7e57+3OCdSGkCHFBCFnvzgFWwFQSNbBbPzCpPUyYbzlSHUsLpOkRxD6Pa592+A
x3dKvESIP/XZau56qkdwka41CuXI+1LRH7Ty8P+QXfNaKgMGopS5ZgS4u8U8azbz
/j9s+fpmaeAowQbPiv6oucbALRqSNATlxvBkxZyWvOdJjAjfTi2edSKAXXG7FRrl
WYQ5vgW2WiozEr0KI2RnTAxiJLTdC5w/0nxsIRz8T/4VHmMnlod99L3AnGJgb8qp
Gadwy5yDBl5947MfRWX5rgIAc0J8yP0eqNxZ65gnMxRGOuAt0CIIiHddA4j1JLdZ
Q1kQ1i/zsFjij59naJYIhxtXtt2zhLfX7tl4a5o7nPjDQUwlOMbnvlWn2tRFZ4tk
Ci+NBDGPkmMV6XVw68A50oNTLQkI/W1dw3t5nz2I5i/4t1jnmRQgLSu+MdpaWxpu
tQoNmMsDJXx0ahItx4MrIrYWc+LAPhvw1Uoy05dLB6nkMimcmjoojaIZTZuRtQtk
LGxwZcK7/rFl5XRXKMm0zeq2DQcZOP3JQAJ+J0To27s/BLyUIp8CPe/8dGS4hbS2
/BuI9oADAE70r3weXgB1nFC9pefKVxpj28CHUVnRff17hbgLLu+2nNRNYM8FlxAl
FHVCR/6SzFKq+4Dh2g9baAmjZ7F3q2uxCMbAbbVGSALmNYrsHIrLBeAmM+LuNA3L
sqFR0ogMl1GrkwsgWCB4zju21x4pMLfBnRnFQfsSdUJ9l9wBnxAuVJD1+3AtRQ5i
VqOC85F99/07hau4i+XN+TLF4u4QL/UfRRzbvWeF3MFAIhhQAqLq20zv00ObRtyg
pqSfr31IStPn+vEhYqVBNNZSpmASB5kZxoifcmZfe5/dSs/LZFvv0QSKKx22Nc+l
6USJi3tYrp6tJ7zWUXxpJnw4P5uLyuPsVhetIlJlG9yGKYx5YVOmWU8dHtoIKxok
zduHkVcK/d4xlIhAsvu61vZvUvi2hn0VXZQXKgcrMcI3CrDUmGax0hE0JOh8ZHa9
d1A0IcaZX1UrcjKHgVYmqNiFieVm6s1hN7pGUP7SI876HDojYcNhm8wqWk9N6esO
ilIG5/1bUXl1XTnGnwIMIugSO4OOGNHnTS+oIRvBBkJhd/xDYP2FlSKidWaCFxDA
yT/oSclgFH+fz0hg8GV1SXhXEjXIXLSVMAVoM2bsl1dx9Po4H7eZL40zrywpGepk
inZ/Di6CaOT1zJkYTLcIeXtL6Pj8jD952pKPQtfqfZWmawPPAI7uzWIoen3D2/i2
ILHg2P9O3fXDafMsh0t0KAaOuzoOzCOELxxThQj/C0MTvqUD/7gez6MLeeV/8p5l
L3KBtE1ThXxeicaPgoSUpQ3BzT9uDFAlGAcsT8D0XjIukIJYQlTZVNZz4D/tuqsC
QyL40bXG4MvBjmaOTUhZG0FrjTlLfqyZNucLfEwBVrWR4rG3k6/g4BkIOzXapqbn
VYb6oIUCrc/GYOZ6PylLEbib4mplMiS+qEnSmQRODUyuuKjyFQuC9JyBxplTDJjQ
tIee8+2Dd55u0ekv/Ack5IpmIzg/ExRtWTb3fQT08TZ2KiV7YRv+vpCGYbD2vfHo
tqUf+M5eYkt3Du2ZV3Y495p+MuwjEjWdnza3FhAQNl+4Upgmo+4x6dcdz/LUOiy+
pT7MoQPyiJc85t9ryXOxTBgzx2/YxGnoeMxT6hbEv0nzxAQlbuM7v07Ai4+iXVPx
RYCpaITht7AuuVc9aJB+Mag+xdNhrPf4UPk3CNhm5x4rDjkNJxJMovCxyQGGWKKT
ZodI4WCvBAGjTnwaHHWq9Ek1s/crO2T722qbkGolP9wUVm5oJTgC5gw4QVlf+qQG
I4+jX6UwC5v52JeMnSaHJgf77MmdhYATPnwjcrG4WFKQW3DZn/UzAVpe2KAtnJRj
1o3eEwJ6idwISSv4NB1RfmdewtyruMVn0iv3VjmyyFFPpF7NwKYWt4vYgvSKbaG3
lV1nE0jrE2d5cMs6mBhlQoNproY+MDIw3bVLqy/tPjy03a92c4HaQAiFnoFA+971
RVNkLMhsqTY4EqEe3x2QRb7A6lvkXDlsGXT40r/BttALywhqDFr4B365f2K0Oszn
Pww3gVwCPTbDY3kP8ak903m3bGiT0wHlsLZYCQacLUVPXr/dEUha+VdB//IFJnAr
BGQQjJmkZJPqBbOvcj5asMR+1GhVzpK8n2mS8yfy+nRJ8i/N97XpYVpkrM0kRm2+
jMEqa9nH+AKDYW6SfaTdy/bvqsuzIu8aGsnec/bm+i7cFrcl12aB835J2w//W3Kv
W97nQsYxRBmAy1lO3PHKH6VWUuaUJz9LGn8bkZp8edYsn71Pqj7WM5M5si5Z5z/2
W6MwKe03YcxK1pe/lDWK8y0VjNdmZF9vRNfzGBXHFSbOMXQhRyeJfwzWXI+MucUm
9bH1R5XL8/BtI52fNM4Jw+g/s7gTcj9g1V3tcIesDci+9rfI2clZz7WnZOVScBMd
MVM6Y6eBS5zGSye98pTIGDCzWMsNXnFBFhb/tz7TshV8P1SRwYrDmtTlaHmA1XHj
gt4ULngvt+AqwJ+9ktrHrq+ZvUBuxWf+C5MP6wtLquIFK1mAxZAB9YuN82fJibcJ
agcIxjMVccbw+AnEcH/fBNtxnj1WZJb7CLFxw4phTi0i7IOVw8iuISxyYBdET9WW
oTPj3yfXsfAuFcTRyy97Awh55t4dgL259v2lzDJX+99MD5226xGxsik/UaNru3a0
59gnV8TbWPUXAH3kBKpbiNCjvHjcO5BGt1vOwesmodUECmM/E+jj/+joC6yy76h6
4oJTSynj6SNZ3REdNYYZQw1P4xVNQaXriEqVo3pVyM80Bqh6YCIFp6hECWHBPJ0u
gLklq7el2JbgJuXjfEcuFe+g1WSFNrI3sFeOWveKsVR6i/Y853ZNkqCw59wMvmJU
7HqgOn2w2Ffy4dZCE6RYikN0tO0NfWXKx4rFmXjoor3ycBoZsnyQbtvtKbOyT3aX
ia4TUD2dkwkHWgYzzsEND7d9hsclaef4VKB2u8pCvNj1EUpf4vblopugJH+fMzk5
o/+6OGMZ9VRo/DYFvZE15cCaPyUjKSzhzMLGOdcTdK3kk5wMd9LDJ5ZpgvGrQRTv
ACnswWU+iz+dfcndhEPMmU/YBLUn4qd27dFr/D8ea5hn9RtkdH3idRYTYC5K9ptU
lJaCsDxrnI+2MMlcT+M/uBEdSkTGQ5+7rlpkXvZKgtniqWeUDGSJrdEBi06rlnMj
XkoRqfx6YA9yz0O65HbNMjjszX5CKsNOHgMINrYKCXh6lGI9YTXNGH5TOMLxSJwx
LwEEnCE8wW6kIzie0WYnUPhb12Tfc0rSESASAiSEdIBp+qkKd0k8SNqw0NdsCOrO
Z4TgZnHTDxrHlWdK4iyZO15ME5VD0Pm/xdlR56Sg5jh8EKGQpzTuU35lr2/X4VhO
I4ogFuYk2nXKozMFHQ5GrKKX0rTgYnIZ+yiIYmGkh+Eo/8SOAMKUfEwEQhiIUeFh
zyWnO563WB1WM3GL/v0k14ZTbNxh+QuPEoB/KQ7gXZ9cGm8RBTNniDfBZRbh64fO
84fqWpBo3JGlYFY6B1aTF2LkhBSkIaGRuzpsEZ+4HwXiCl0s6QWYcEw/q17/6MXL
OE8+A/IcC0fjiMXMowhke0YoApx0dFFQO+RfZ5PADOPgRdNDZfI3hiqyAN95IoJj
xTePN2wdsqeSu6FkxNiy+VpyhzF2YDdJXkoPTr0LPVgs6xEYpEQ8uXiujJvb0xtW
Q/RNJgmCZuBQB2IHbTyITQjQb+bQDLdRUNLFvmB0h+yq7XJOLuvunbASzzwNyvdh
QTB7W8wZzRyBsJRbxJK4FVsrCEFxfNMeubBErfFM0HeCGj9AZsdb4zPBlja6BX9R
N2uKiqxLbHxA77ai56CqpnQvpgSYWSoiNVJf/i9mzftG/tIAYgn5T1HxSu9WT7cC
Oi4EKv47jAT/0hSDxQ0VguXsfjiM3Lo73F2AYUsyid7ZduQMQabL8vAcqhl2vEVy
/FlTqAHKk2KllXNgVVIbtHHqn0Jw9WtthNRKBzDpjJsZ5PZG0JzGIJR+baet/Y4m
6EnzAdAPsrJ+qYZ+KjMI6YmgH1Z9eEtJjx2CatS3jO3J2LmZUdKvXqYPovb61rIT
PWL8KPiQKnBZ28lCa0j5fAemxB4K7gJpew5uQooY5qI+rS05b/f/ssb5qJOLc0uM
Eel0o4p3+kQgPopGUgWmZKnle2k+l389jmtc/1LaJSnpr40rkyv62gmc5d+SE2/H
xn17Enqw58o4lHxrXb41GKK1O1ngyjq/JL6EWGXdEfV6YZvzM7edaZW31o5voiSa
09dsRscnY5FPQ3vzch0r5wu/Pn5QJOX/oRfwYmKOXUIVwx/GZFXxqv9Elr3RTriT
LHCaZVNdqmdVVkvtDoiGWVy8kV8DK1BJXjBInkW3LigoWpCSsScROrBaXc6iLuTL
H06yF3hOCbok15F2sIr9/I7FeoAqg1Gfl8caQIZce68LDTO9jInLaXIllFbm3qNa
kLyx/u/yvM9WlylxBIfczSWFcsi68dLoJxDnS8tUNuQO2TiCnW/HDSQ+9a1OYKyz
SciCXYda8X9bmDmI4SiFGHQ+0tPxA8kq9gNOth1VKDHTY0WqM0+C3YrJlts0TltC
2Jbvyp4z71HSEOSPbg2rADCdHUJ1vlicOPWK1Iq8cCXtDNSaDt9tU2H/AREA2RX6
ZqUSeu4azU5vaGGcsWP5RevISDD1PiIWhJRyi7xvzpkKV8JL7xA2vecCDhuoqMVR
LU6pLMwcBfh+AJHJoZ/Brbo7LqffKll3wYHK6DsleX+6XZUZNzgXY7ro+QB0bB5n
mSn8ahdQj9rcapvpVYJHvGXxA658LKBa9BUPpCIDJOpCVGGsmMwc41KnBILnArQt
owCljo4FCdaxEDMgCxmEI/n/WVFeKySt5qf4UAbhK8I2j30tjUQ0Z/irxs8JiTHA
EZv8dhvukw5BMbMAQ18M8EXXbpsEzww5ZPA/TgXsSGDbkIwk7OAdJn8qnhq6Jd18
3xPN0nnkEnDeD838J2tiidGELQGuQxQxbZbhVOMbBefP76eCP0diJbcgtSTfOKkI
i8MWelA/KfQ9rL9KihL3gcZ3gmFsMRr/FSozlzoyzU0utvW9kRRPBqihDhQIrvoO
NZWxsiWRq6j78T15hr7QPE6PExjqHzVj+APBW3LQ5p+VfL6wd19bF4BAhtMS/cNG
TZj7BP7KdkPkTSX5dkbGl59U7cvNeKyGQOtbqd0Fo6iassOz9IVeKHnaEuRLM4CQ
p3DHdlwzf8A26WMi6waERo26Abv7jeaMwd5qSfkbYB70QNTN+gX21Ci9oBlWqscw
9TAO9915TqgKMUyoe5fsY6FsexJXrFrnZp6XKbR63q9h2p3RCf1MbJ6moJOLKtJN
pY5smypVXOHkoaomrNXitqXrYBlRzJvoGIqnsD73+oc1Kp4S77gVM0v3Sc8X9Beb
U1UNn+Ovybtc8pdUb0tbujFS59Xx7aeBDKS2q2M05OwcMCJ02htRv8/Xewl1AZdA
AMB90hMAaVZ6/hFE025AtRGLPSkc0Or3ng8Tv2lOQG61RJ1+6x8SdoDxqajr70B9
yYsO0z8zKweYGbUkr5v46FYITZ0kFPNg+eaUf+lhuYpJEYDpFI++aGdvKgYVWbOP
5n25wWTy7YdkhF9qx1+tGmEMtx2eIU8Dr9pzJC6Sy+pvfcDyRr4P9MJTH0qxhIvz
KSRHDrDxWNtIfkNnLrf7yGg7p6X1t41xQ3vQ7e99wjitMGP0z0G3UU4E2G0URZoc
/X0DTST53Ew8z4OvNZ18JxE5hsWIYrC752miHKJv8tvnoW6hRrlu1wGAYGY1d19A
QbEjYAtKiEo1mr8zOVK3tNpXq6mUHXf1v/pyexCxOnGIlh8+HjUUBz4PvT6aAuPx
hsun/2U1UeytHFRF+z9VEUNPfDj5rgXnu0KmByAZM3qayVbsUiYVwPb4LUBQjckl
PZUiBORSiLds34l43G9B6q+aLTf0//j2apE6PYwS8UA0LIxjBFXSiJG4lctdZgL8
iQl1Tyg7++Sbra9kiXNwZLVzq+Uh/HxZ9Up1Peig9YcpGq8ZhcmBeVPFfa42ReAs
IvSH97TV1QVTMVzXzG8swGuc+7T8StAQYvqW4lTOkE33wJiKUw4cdC9YA9PDmFa0
7ynva1NEQiSeH1REAztvD4Tqtqy7VhSPJFnajwrGD4il/bRzY+4Yx+UXSIw1DrQS
MAfoaYLibyKH93mTfg1+KTOGBsM7TvSyUQkW+ANqN4GbDmfZVpQiJR8AERpw9/ek
I5L28X4Lvh2tpd9/38zy0P1yDvWRG8Bl5ACQOaXSp2sws64suzcfgoeM0XabrCkn
aliF4MxgEoNfQU8YpSkZff5C3Q7hiDgyjQqZlhvMp2XFSU4S/ClWrlZZofTx2aKi
HmhssOjcj37IXTy5w7iakCXm7YfEYbTn4oPDa653HOLVvEemU7UHjoKunODpsoy0
pSN0iiOseHzWzi3IFsqnD5Mui7SJg8ms+shuLDrG1XcIdvK9NPl8GcUcqlB6LCXG
6GKURQd71q3Y1HoSlMpQ8lYy+Y9Xocek1fgevB1SokjzondH7nXkHLAkMHc19w+I
rPl1NNx+OuLJ/LDKOM5ukMbLcl/NvqwYpGswUU9FVsIL+JeH660dI+Zlsr22PSZ4
Nqg3G9AjJNtrffhg4+2A2TVodz1KHEebcQt3AEaC3oNviOGdZIj9zZjaCgRuYuuY
hpy1EPW+8WW1gkmZ20TfdOOSdL7L6vCZceA8GFPr9wr+2jIP+yLSsEe8jAJ8QqoM
bXETT0hmrY/1+79Luwf/bPvNE4WoqD5a161u0x613EjtfRo0HvXDAW5RN+b+Fsvq
sNsxVVlXJz75NETr1J33Me/Ri8bmodokJrlO15tQVChNDexNbooV/AU+BJCS+Rq4
8DSqpPopVQxGS+5GIzeWnJAPi5UJuGMpzmCGK2a4ZQ7l89+I8G8IXIj5E6FmTu0o
hifcUr8rRRwhePI//hU89Moyh2m3ZGgLU2e3HHyYe1y6Uv/O0cjJwMY1NG3gAMSI
uSK8C+AEsfCi2n2WC7yH7sr+OGfmb4wERrWRKRxch3YCLeMTUB48K1ePWw/4bgJz
2u/i4Iy+/8PCjnRS2mPfa0kaRQtRrMestjenxn0iCLDOc5JJI2eqquXMtZ3syJYu
kwMCb8b1K1bqLlLRNmakKz0vmE2MDVgtOIeCDqF7eBK4KK7icSOBUzkNJoATgvOo
gdp8WDEUMD2pZUsIVv/QNDGKd2uGXFbuEKcBv0mvqf4F+dqzhsOvHpRQIgYqjVfS
JCX4ADNbb/lKOksLaOSZ5Mbh9PIY5lVi8v9v5djC3M0nYnEpeJFtFFrj0MFa9Swz
pmWTR90/q75mCxeo3MF2O9j0QRABYHQSxPnQx91/46zvg4CwniQMnBQL+kXN5hV8
CANsMD2AJKt5pr8/itM9sp8ZyCX3uDa+p/x5kxs9+6hbgGLyWdo2w9EjrC+9M6DR
/of34cHj7i+UY8Tvbk8HgIjAZOPHW6sJzgk8L/6l3bi1b1iDNrX0PSwliYVlkvVp
0mdiuwp1GGukGReQCtR214f+yoMcas3rhwNMYFJvZZ6vgm708HoUF29JqB0ExEK1
2z3WdnsIXngIoi63LKnADXQWST8AFlTeWOgHmh3lsbvy18Wi7ZAzP3gVpgITPV9/
lk6DSSB5d/VossWM++bKcGCPECFonllp2fDKI3ePBic1mEgKCtCs7DAju0Qx82Xy
JSXWUgFlncQCvNu9E5qr2t5wr1w7gIFOVG/DXDMgGM00GGHFauu31OHIQzvquMdk
JrQijTznF8J6J1um2/BqAsNv5sdqXARwbv8EF6maWm2tH8XvfG2zciTYA7z1oR1N
x0El7UUA1U8G5smoC3feg18oPO5tVa8EHZT1XyWROrHYkYmxApqjzMppKPyzc/Og
ZqHY9zOJ8aV4YIDc0XeLuk8V5WM3Es7TdSH93DGOIGdIuiIgKB8GP//b/RCqIVOw
K1NnJoy7USMtQZnO5SPirjtcmAPhH3NVhCXilkXFbAFRvJVJaonJPg5hcUYe3EDE
Bm11yJRMOp4GKGewJPuMPtCXRX/2Lp3S5+wm2tbIYqRJnR67P571jre/u1SSld1M
ooSJizMWPNxGIhJV2EWn0venQtcv49tIIcII9AseP3KE1b63+8L4XevTXs2c0lyt
2xhfWhfiYuqwPvnEuZPrtYzTLK1gq4c+c83sybxzSTcoagzCYARIi3pttsPMzq1Q
haZyQNO0TSmHCAo06I75/oyBpeB2x0QLHThLb98WBDflcFE6eaz0l7QjJcdg7FH4
ZC4diHVEc8WpAZvKAwLcQj55CR3i9VLlObSz3inZ6/dQ6gS4ssJehGpN9XrTM8JO
DsFMFzq2kO67EU00Fv5xMsWoceUQ/WA1bpzG0Rg9/Jj7dXxcLwPSOZhQ3WmnEYpB
V9RvRifmQSbXtN1WKw8SiQPhezyCiv4B9f3n4YPVsvY0drSFqFgdsCXl/VMvuAyf
E55LnExJpQkGCz5Mr27rrfUXRJypxqsTVB7gWJkI8Med/DIfp1ekWWX/4uS3cuXc
EMqqzVbJx2RuYR9ezSUZeAymY6LEgZKJvKITGdHY7Wu04S9C8UqJy+3f/hH66DzD
d8u0ijuIllJO5LEiIPhOiDOEi1iuLMjSZNDJKU2JxuZJQkyz129LDm7xdNMTXywA
NCrdu0jBBUqJzYdzdqzSLy/zv+SZHPtWgGnqGRtw/ynDvYknQlng5E9oQT3+F3PE
RhPfRxL1wi6dYFUUaKAYeJNGL4ajgaUx9Eljq8HES9WzbdnXJvCCsFodWnERIPJJ
IGo7SXrIZqILyIhXNVQNcjobRx1kD0QfvlMDZvw+8uEtvcurqs0nCahjRdSYEIu1
UD5SR+nlNB/vwdMPsw/e83shVsi4/Os6uFsHLW/1zqsIdCgWNqBcKQvpG6Eaollj
DymMRGw5MDwGCFK5vHD1U1SSJ0WlWahZf2oWqSBjQERlfTr8OYDBlFbdH3vUHSbb
8dM/wLkRyM4kZtqIdfzyHOdiY4aMEhj6Fe+IX+KfZDRs1EzRH9gXcNT1jHuCiOyB
DsLcR+VHTb8FnrHZmDP+C86aEkqIKQ0ObP8QOTlj2l4ochfRD4wWD5YEQDw6pwFW
LHnoBomoKO+qv8n46SHfmi+w9gUg2U2WlSqONL8wKIrPKgxeHErVR8IAZFiY1jb+
UtFJRIoaO9ubUIcMU6ubiWev+BoLxfos7ZeuwoYH0Tcl2cgDnkBU2nuah2SG8xcx
9F/5AlFbBFAiYcZA9BNLMwPZpX9ua3eMUz48A9yb+AQ4nxZTvP0NH/PnKCEjFxrP
qgvSiuAuX+a5TX+RtQdjg16AT8zUVYGd+J3uJHVmczUZxm9mZkNBKS73A0GUwU9g
OtsLjtLl4AQOTnL3L+38uQriv52K4wQBy/u9R2LytsvCnjSHmF0UBuJgRsgN25Dm
cffhuU0deDQ7Av8VpslKCFfKc5RimqU+olj5AtiBZ0aSL/6kBLivEjaLrF6tvEg+
YT8BWxAYBRl005jHBgGvF2upO7gsTWfN63hOSY2qTCyhlUjHTh+5CbdUUS6As9BQ
ivFTilJ0WYKzAp4QqhDYZloxXRbaLo6oiq+9djF4fuiMKY23555fiykbilasaYo5
FwIkoYiUxOPUfSthkpQDA4yfDKzrz6YG9MA8vxjjbvvWnnpB3HKEC9kWqHEG8xyS
6GVfRzaLgbbL12bN+mw7yLE+BjYyb3X2Gwky741VO7aHDOiuug4yWMGHrt+PubrS
mKxQ00w2VvZZV+105Aimx3yvjilmiiFmAN6HP/k8CmFWWyy2B6hrMvy33//EboT2
6KqDPcdfJeL8YQeGNoyEjMK8LY5XKT85VDBHz6O3Xjn4ZVFvjs/gg2iHraE8lU/N
UVWBE6nhLDsz/XloYY4mXsII7HM6D+B6HwaIsF+LaOmQFgDE2V80lybcmBmKbLG+
8qZCZ1QcZnq5hT+wXposeuIKrDZqGKNlL0848hSbERgpEhyvNXBdce4SkCh3Nwjr
OZ9AJcTTt4GOd/dP0m9k082x13fOXX3ZrBYK0bYLlLKYT+i8YzIsQ4ntcKxVNMY0
cIStdPrcJ4ZcWQxl/kHN0QqVY9pnsEwfBjdnGbR5dJZbXffxNZKOXjTQOnDLGsZR
0Ab+xdtuIryUhPCqO7uI8YZHf7SHBCN6aIlaM1/f+63GFjCygWUDApeBtDb0ad8y
4xPS8SA+Fyktb/c7+0G8js544QWAjWHqK60IwZQJwRGHstuigB37GmKLN+2n6CN2
KXp9L5hFvJH2fKO+uBAsxhYwdc3zrup++V0AMwgf3xDMXSDkiMS4VvhInSil6ByR
TLljW7ApjteXQ1VeMZ75qJy+oeEbhFSjLP9LJedvn7vc0cDrdf+PIuGTqTw6aCRb
kIJqjoAQ/NavvdF6Lk4TlgkrNaJrv3HVmlhNLxXFuKAkbMiVlTyVWOecxxiNvuJU
ysz/sooRcBBAUiwYhV8B5pnssy9X0eA46u5YHtAjDSibv/k+sdH6rHZBoFO2iVVu
BRAzVzRc84VR7du5WVQ8cRFJ6IRaks4L3rNOGiL9JdHJfb2fXm6UQ4Iml77JABSd
rUcIEtE3CGXI96ydtr8+bBbpwS8SZh2vA8E6I5LKoELi4F4B1FkLiRt6jda3sF91
eDLm5zzqBoPy8uXGslFo+Pjk54CenrX39Dw6CGFQ6qjHWfzlA/kd0RE8KLetWvtK
akPg+UhhSUqcubMC25zFzd2U9bDmOAP1/YcU3Fijrs05OHZziVGD+cGKfmMQWhTB
dEnp7zZCX6fPRWO51bJQGM17VFzP320UcPS82y15rIAo2lTM8RjRF5CYLk0olTPN
Ozxur2LFrTkeFWzrJKQyBFllrf69lpYizlFx+opm5DSLhyOR3RK0eQTV3cYIPJIw
HKFpZVgWX1Ayz4rsx16BufSYVjiUwTY2FVe96FWdE3lmyo3zEFFZ5FA70skVZfvd
eS8DW81yoYsexsy3u7e2vT/WbEpEgn+/gkZ3WLNcEtia7yvkq/7gvapiZGxRycsf
ri7YnBat/EpHqzeVfS4pWgy8J+D0M0ktywm9POMFqElESfUA0QSOzmAgLRuQOtEh
BNcuZUAzf+5YinSCVLqc7gZRU6Opdr0LHoGBVm26nlQnXZeWpysTsuSsGkSP/xYv
SvUh5gqXoaC1jH2MBSf5CuhQV9L3lVYDJ4MGmTzqVGU7SXu48ijUn/xdVEVNI8Af
ODo2yupYgzPK+l6PKraTR14fqL1OeDUan5L7wrlhmZH4s+LS4CxIiHXNo9GKvtm6
UuEZA32igw3XocYxVsGJM7hgzGiGPGii8Qth2KiiwJgUgt5x5UyugGoG3tvunDdV
U0jJN7/l/YZQhHhehs3KDBaFbausUjVgaGKSmHvknV0rcLOm+NVXxyvloYmK/b32
6K0k2t8jaon7RCTojtd/tCCgSBD2cwMN6dC7rAnu9vDqNDBB3QoFTh6H6+JUrWup
DOxdr5WEQGhPeJBpurfJz+VMFBWcZLq8xsD+/uIaE4W6zhwL+SyelZZBXXH02WIO
eCOWrtuit8BX1hwpQ0LC6e3jk49B9heS7YvXOUjow8ZKzxw8crPmsVwndbU2V6Qt
sjO7FSNbzl3wND9EjK6D659J9WLUXwExYGn/F9MdlfQbgfEmm77XyIsTGkbWrfYQ
/7Jh1mNNyI+nlYgE3SgFvvV1XXCoE7FYSGmjAfHPbdr1sKWaG4Rgu328eA/gESCW
949Fmujv76N049LPzaxErXcPLfliduGGp731lM5r8bE14GpeOBSB6KaLsq8JxxCW
wJhzQDv3QEFNyHUVgIGkPmE3F3RY3bUby8JGJSBZ4Jvr39FdGJ415BItsYlcVmxk
9gZ93/EynZ5rd1nihFzGnCTPNegLuTBnB5M7IA1X1c25ng4LZ/0U4zGph6la2UOM
SeZALpZqyjjxxm/ZqdKZ6UAgmEsfUjKpHfuQcQ1PCXyhYbWhAErbSKesU3Ye6nfl
ZyGPBwz0rwPpM+M/hgK5BbjMg1memousI905EeYEIoUwSUCIDNIUC+zoF3bYUhpR
f9AVXyBrGAsACoTowFVxlYy5DYIOcxFsjw4UB1KeVX4E4yAPrXM545pUI7q8vMI4
hK7qwIUW5+LVxHKOiR2bYHxco0omssd2Fijm5w71exZJBiDmOVai5ZskHXomDlxQ
SFZktDPUXUVRJUlsUKbLsWtF0kNmBYnBAjxMbNfTNatfH9w9ZHAz9rNIKRJhk0zw
1QfpRianHQ1LGO48eKmpMhyAhPrZULJNa/QTZ6byaBEZvx+eC2TkebbWqAacf8Tt
BNPlVGL/+KlHz8ehjTbf9TIt1fCPxgxd7S8521pXCK40NUjf3UG2eogUYnFyPZ/F
ZGFpj6N2r2ztKpCkblIuuzCQOkARMDauY4A9/LQmfpQ8NRtNv3O5KMRBt99U3+oB
XdgVl7yyAut0mZ65cV6MhURGcOjuZzyGhft6wNlfLT9rK3ztAT9fZFsv1nD+PFnV
jSEGOfgQz6AmjAbbEb4jBLP68POg0JloTv4PXKkUdmc9QrsBsS7+RximyjGwfawG
MOSrrA7mY6W7rf9PbP9SJOjC+HOlxfgS/XVHz2IKdb2t+z9gKK3UDlPYbWz4Fjbj
IVi2wERMy6B0NnvEG2bkqbVfU6Jh0ZFoQGvtXGodZpdjEGqZM7gLHZgC5NT+1sIq
er/zgrdXyO0QJc8PYu7bid5Qq4w3n+nsJe0gOZl6hHgo1V6gRS0M7+dUkOCtOqY3
jpayQ5t3ANzOS4Ghsr4FgoQ6GA8cQODkUoYEVxZD+di6uN7tfE+rGIqjmaB9juHs
fFhLusOyJXGOpbHgzylUGHXDDhzbkFZ2OJy7La8Qn0Mt1VP6c1i+s66KQoYMcKxf
gUxIxMkz/TzGVFuqPOIsLoBX0J8FAEcrLAWT8E5UvKPNV8E3/VA1hZXvAJqeoey6
Yv+jck4TWk0PRgJ0N4VHqlhILW929J2LfAWuasUwKkNsMfGlnL084+bf0LiIIczj
7A2zX2+5VStzSK9Vh03f7tHfogz2N8JHPIMMZuZruC5MLAx6DMWbJ9I729Np2zS3
TgulamGNL8nCfSJLl9DP/Dq/d7HkR1oXsnb+oR2+4iS+fMpvf+YnhpqXAIzvLMvP
44PmZlFvhCC/ne14AJSgzcbPEWl7SzWn9GH9tt4crPJfdgfI0A3Ycu4qxrgGCpj5
IpZo7svnHhGPDaPTyTAZsOy0yOgo/sNVn76O5YUmaRVeaJrDKjVdtsZczVx/rLxA
0sy+L22WSnMIn+2I6i+kveQXKv5xjtoZWaaTeOczS4Z4cOCzau9sAmJx6NgVWmW7
ySgsmq6V19Q+2z7own/nHnTIOJTKlJ3VV+rL9JOSG0ydCzO0VB3MVhvetj/uj+1o
Xs0p1DsStkwiYLKukpnEkLXcAtx9a6qKrSJXJ5q7AfHiY2MJA4B8XQkcRh0sRUBa
PL01H7UW0VqUs9NO+b+ypRqjtEhI11XriquFGQmajXFiIcEPgFn48O4b0+YIv8sN
R0kC5BpQMtPxrfqswHUMfM6AwllxssiAnaynz4to8LM3VC7pV/vrf9VvtCgBvey6
qYyD9RsFp9rM66GtaGUALSKVjBLGB9Jse6bEr22c1fo1L1qE8Oh+xhhqm1rwVubP
SdwG1tixV3qaMlM3eHnuS25GeK50oQ42udglCffqM1mIH2EoH8vfzkBXhsmmCtJc
oSfWt7KA9jR7XFiqu4pH9gil5MFtL+7Ya0OyNmb9q7COzFxoo217H3o0xm70DYZu
xfXbTeEtg6I+3HXY5dRCoXfnyR89wSXTZDFEWrkFE5EawioNft0JXQitf38oap5g
NhREiqp03yaU4POEdme9SOWQEVKUf0Gigd6vi3dPPrDZhpOOeZuqI79GUOMdx5jP
pPD78Mepn/YRBZs+iYMilN9VoNy3JW6qFNuDlsiDqQhFzyZR5yuLBQIlGPH3QVAs
lJ9naYXIOnLq+Hm1iUI6pWMktqsrvGtWCKBEbUoHWPJWsBt9jeFX1sfnMUsshwK7
9Kxp1NVfya6ZYdC80Mh38FWq4hCLpybsMHYIRn+b9ie4Z4nxiPXS+VCskE8NC1Hv
CIIUHan5mo9X8pDfzznRT2E4Ed825w61BZKg1oVfrt5XPsF00eLegkfFl+MN7pUU
Z1P++NeoWFbnQ+xmTmd7kQnQww8ohytbvwv8EI1jVX88sGYLXEkwHYpydFT0ZWlN
kd9HlSNGdEM8LDRvdQVLO7/Z6UL/gDqS1HJ/koKmRD9lbQHYjOPMdlME0G51nQ6N
N0cCsmdT9+VfaX7nCG2E9d2EvPfqhBJ0MsHPWpi09RXFwaVRBshpUXKUo5PwQkOA
f/7Fj1+SdHSfZVajJt/SFg30DbGMsYDAvAANEmDWzbTP9ERtyY49lwJxWkNhtfBW
pw7T1nvNM8e19jhtaQU66oaF0nJnwhovXRwfyJNKLbyL7bs2F60FCxdyfP2Lakqt
uIqAK4sJ3kIrFcq0hRRprjh/hsu6/hm9ToGJ0kf0B6l1Q60382AimKUt4eLgZq3L
QgrXY9SaoWwJIRrpU6B4xi75R6OMZA05wVutL3+fg4Y0ZaRxnB+SVSZwj54teLDj
biCHnMU+mGVsuthAHAwf/A/r7nkwx9/yW50iOMwA5dgPU4hZ8WwrnOwh7uMIAEJq
8fc7FzCS4uraBV715T87Ph+7PrjNsidaU2oC1NFFCm7GPpX1Vw7zG1TIVOL4m0rg
cmtaEiIgTR90wO6eTdfYtrMMXDp8O2j2XxdNsua//c5Iqp4spkLxii07B/gy5GV/
Tj/uBVTjTCeXpdurLBp5WW1IJe/Rz4GHiEH6QWuNejfI1eXNZXz51jY/D/zzuA83
0hhAx1tu1rXVKrVAtsND90o9t9oCotnXUMu8wBHVHn96Ga2TAyJHkhX0tm5sAs6X
Im1/tR0nXHr5ti+qNfuxtHAuPr7fzyQaPg/QPTk+z+/BXM4KjlexdbkzWz7ExOp6
+hWDgt+qEXr4k8/33by+4IW9Zdg9R+/zjAEUEyTeNHVy6Q2uHcT3wMYDwDK1HLi1
/Ks14/Aam4mScMafT+Oq5PgS5TLuzd/mVZIb/4UWsxCGLhJ50leOdjaKdFB4nIE3
l4mKy4CyI5AFqdOISJQ+FRYFp0xiCvYycfrSKSAlF22ytbrWdz/l56O/aPm+8bbI
Hfw0K8XV2vZJKsoX0eLIZ03p5YghgVAsuXLyI9/rQ4UVJGWgQN+FnJlq+HzIxIq6
DB5WBt7Qhc8lJDYR3NG6ixtl4yJeKojt8DsQhfJM0Iv8Ay/rzQ5rFt9Lt7Cira1Y
LrKUL0awGPE8cmCtVhx5xOPZRTSRrraLYoStv4JvmDB28+87ywkWaAsb+il8rw5z
PEsnOmTGMHZZmyX0R62FcPD/znbYG3uNrA3fHFW02L1vh5l+6OnFiIvvu8yvvVQl
4JCYGpbdaQtTBLMpNleZxH8QbCSdsGMaHowm0xIYEJkhqj5UFIGbNqMd+0HyJbUa
KJF8feOGORElaNdrI7sPbXRHTd9cOHAoOgY2UdN0mT7ElLU10jtvNyqqhXZb0J8T
U6QpJZ0Dse4iZzxUc2mQHKez/fjuGzpI6A9qg2OglEWLKi8wy7I6kI28Q7PWGr9S
HNZ1dfVWidbgM8hhGIaa0Irel1NXxpO8pHEwuguJYwEAOu8tDGyxY7GJFdqic6hY
4Um1jIV9O0KUFlLu8g5p/crElpyn543YIrI8DZ9gsjfpDGpTPqwe//NPfvuFkR1n
dFHTcTlY0y1P8/22V8DsMRNQ4yIyFp5cVVEk54/Zfoizg95G6MAreV5kd05wUZQR
kkobl8ZN9m0IW7YzHoUp/mniwo77fBW7Pt7tlLdXxDgOWZ6xB9Bf9cH2iCf2DrNf
nel/fScsLUTUg6WCWVxASeMEmlopL9CFtcTeXMpwe6LKcVbY4Rs2cL/34XBKqNHF
wHKCULOH23ahw368l97jwwQs8VTwpAWNA/BgcIbNtuQt8QAUw1c0PpS3m2EPf9ax
6RMTrj5yVIs768KA/TYefJ6A4eanRBpOBVXTkLh+SSrN5IxDEB4zzrrXEgMzYrFO
ws839vnu6SHGeG15hAjtxYfDoP/Vx5b+V5RdmO04/rCGZkiIsiVE+2zKqmYBfyBC
x2XpQ09SoT5vRzyVux+kyeUP2j6TIo9E5b+lcJJRDxo9B+sfgmk+Zq/KrCgyqKN3
YqLR06XICl8VhfZRjhgz5tPlKBGkG0/Gj5Z0Hd8qMWY2juNxpN9NKjDgIJnxwP9i
54lW+PYz4PV4K4ni5dxnj6b6O/bzqcuyMr2P+P29Ztbs71dd0Jt8q8cnqkmR8S58
qp5SQQl6R1ZoWh3ZD3En2GecJcj4sLYZc8cTE5JNISUo2J3viCZZBAQUXVr/lGTY
h5ngugKDf8cUWcHMYCx86pXQzgw1fHJ6F8P4399y1WGZ8g1vCDzOKPUu2pQeR1LU
KR770WzD8k/9kJb4jkANSdYCibLobcW1CBfeuXjwFR4Z1p6Zy1K95p7lwl68+Fe3
Ye8VUql4ZbUPLjEa6JrKDDFXxBvgoLsNjVe0bJvD2msNbwkbJKSoJe9cB4025zUk
lO3LESrGIYvlBv+lOkzzIUHF6GjQMQrNhDUTBPcqorkPqbDkSBNOcrHbWxMgvoml
UlaoZ1/qBS6YCRBT7/DkZLee2gTl2H/bO2ciVmsiH8vJLMtFZ6OUGjMpedVZaxTe
tTJLTBg9D6+VFtoitpv7qZtVItJA8oSFRJl/jhXrwmK5YPvcMAriVoXTMMvoTv48
5XXbX4fQ/KGA76Vwk+7yDQ87kTxIrt5Rzs2QlCJmixEBC5hcKY3BUEendcmuPtEt
+0Z42QNuvBWkmDJjy9rGUqiN2cABVd9FK1A0mZxamb6T7aXER1KUsgD0uIi4F5Tt
iskxNlV8S3JKzTFZVDcqIyyklJX452CiT6ke10Ajih3xILB3rA9DauHXitpBpzQ7
8pnUc4ujxub87Xc1U5hJ8N8M+2S87Rxc2XthCGSH3UZsF3R35YktOe3YnMijrFm7
N1yOLpYyn/tx5xsaCPBaOGzG5qHk+X2dkTuQrAYHh+RHdiEfzRC/fTDviGmob+dW
i8DmKoSwDFPEB5YGVSOUIGjLzITUnB6nDo8BahZvLHwlt/loJ8pHEM+nhZD51Q+F
5qAJVA8+hBgMsv/+ckRPkCpdv5v4CHyvBN1/1Gme9VEyZrJo9V/dCha55nK2FG4/
1zUc2e7tUyWXtuK86+Qe9k92cw7DkMWRleQKNYee5Wn3xQxm5KA5YMSYuJQC6oSH
jE7xwI9Gf6FRJ4mwBKxd75EkzhnM0S2J19vxwkysTN9lQlIKIwoELRTuYBhnRPMI
//56gu5lX+VsbDrcxIf8Tag4OapMmYu5O8kLJExRbfpaRfJ3SBJlhKLUtJvMf9WR
jQjh9qZ3KlItuRNWhrZzOeJxxaIXyFstMHyKp4sA1kv5sjNwqN07oE3IURKQI7Ub
BJ80vxBg7LTFbInPuBqHvETtpJc6dZgZ/cGlrnXUDGntMMPH6Xjtzilh6Ppy6060
BbDRLsgtwLbyMjwTLobriRDDzeEZmJdEQm201z1O8bzmgV5waBLhdCgMh9PpMHvC
AI739RiDjrsv3GCt+bBI2cK6MWf298FZehn6QO7UNTjZZawI13XxObXMKdy53krG
3slMgkP1zILibfvnvn8G12J4DT4Uf/Fbmy8jtYPhxzeETmWjmfYtBKdIbKbST5Nz
843QbNv6r/mu7vwh08KfADKcc21baPnXwhd/3ykZnXwy2xW9UpScZtn70lHIJyIx
o8zvE5THFqk65SGOs3JiLZBy1LOBpA5+YyEO/FsZOVcyKNvnH6ZpjterjvN8wizr
71wVjjf1lB+KWfmNLP3aWfEaf45PPhNmPCx3b2DOgOw6o+564ykTI6iVgWHO1Hau
0QW9yhyTQrYvsTWfiJnzAxinZ4h8pXrG/07xIQoikgEQFzhV2vEWo4ycvh14AcnM
1dLRogu5DGx++hTSDweCwMQG1w/7ufNh2hBuRiv1qQCFrwQQe3aF27xQB7NdniOQ
t2I39qg4fynl8vTVLf+6RoTfzBRc6cHqgSDpKR3NfmsTMwiHNu+POKpPx3zHBQnF
3BGbKJOKMBws7MyQbbj8ldsq7OwHViOKx6lko2qoqoJ5m1pl+0cIExAEd7kno0jB
uw09kGhQPA9bgv1XXRG38dXeHFM4p2kFS0+skGEFUb/Mwa++yzJAoeY9PgtaVtZH
V2ooYvY3op/4w1KxLpa3pImr3lajSYkMMWGR2AlLqgZyV/FNr9J9RzlKi116gJpB
8X0H5QvFlsnvKesohIIE3b7exGcbld67bXlltzxb2aVEGISOnbhiXpXu9Uhw2bAP
nSNPVmUni+IFnzoUL4votedNP0D23Ps3sbawn36p7rBhZc3mVHmo17LXOBIiwZF1
/XavgkoTTsvrqhBvXudvAA+6v+I+vlkWLZ8H84ezbNHdN69EKXDMzmcaTcTpor9e
atG6UXHuzJpAaB1mSKfw/0spOB+Z7E9tK09KJ5X/tudJp6oMuU6kwg9HhLjN10tf
E7Kmaz15CfMbGGSKXlm9oacj7zm8iQo/Ej9IxzIl8HROlBoiknOdJo+46L2R7MHW
Jf2ZTy3xf/V6BdfiRiuuhaSWCjoLeeCxFFzsoLx5sH0dl3OOuBYioxD1BWe1wqtH
iMYts/wmkhnzQ2NoANfg6rY/qlj53aSY++rlI1NrRn+rcZ9+UyAGk8+pwo8//xBA
U2N02KHySYXSbMT3FI4RDcCAmjM2HnkG4wDzNqwzgRAD2Xp7cIvGY3znHPJV8Ww2
eXbxLtQCOhAyM0WonaiIfO1cuwpjaeprRsKXZj2+LQtFXxsEUjxFaMgX9LcI2B/m
UrmHPKdZQoCszYGR/qwkaFQFLSLZ2BDVbTQkFZNi0R1YH5Qn+G3Gp1NKdDt/Ower
i0t/eSDxSlNaWGd6nlGsU2GPAd22TjkIonBywy6ZKHJ7jyc0RoKr+yYneteJOE17
l6BPDQ6DjzX5WzwzpSFY6tZsHMGG3q5HtmcY47RSYr/1r8TmnM93e0MW1ZHfE3JL
b7myGEt5/WZQCkwqEuwzhPdhJVjyfIysPI322+WXCVVZGmJatXQxHnzrFgC81qII
/8LLgqTlYptR1uXGlYRrpuqMr4Np3y0WMEfIMY51mRa16XBCa8aEiSDpLL8+R/5w
0i0ODqGVxog0wJgirmfvh3BtbOnuXwl0S3HhBZjQkAg+ttJsjuK65ewxWYGZ90vV
U4wltrH+vKHhc8Bzzj9CCveZUwf7XCca8cSRvTGidgLWQjjrde5bqIqo5+bmE1t4
Jt+Ep+QPAolXqAWll/uro4cUkSAuVZOudpyder0HOj3LjRqfOuFAvERFfzMXc0fL
1tce7oL0lLEZs3ixppJ0Z4AxKe53XabEPie/V5bKzDEZackybjNwaVxrIEqBeVS3
80TP6uhmWRBNEuPPbAvOlUWddiE+W9icHf5alUX5zhjIyaw/80FI0OjsEqMFnlQW
8jIuAgWpbvVOoeLkCXfaOmw0vPExDQbjNp1wER5iC194lwPR6v47LcabpEeewN4R
1Jd4s24IyHAf9mepKKIv+e8RdDs7/tjZYVdY3s/0hG1DM4scUIXDPqQl4QlgrAqv
WQQb83wDJVjD/qjhredU6Gu41YXwV1J4D5FJuXYVoSeV6dgXNV9PfSIXERhhjwMA
6omhf1jIk+4q15I7cuXiw73RfZgirYAClEqxx6B2WSF2blPYF5JoA613v8JiBMdZ
kZtFpcNMny7dtxmdWZPBbYF0vWKKCMEzNAQtJw46lxJSrDl2mBQ4unFsOri4Pvdd
G4rGe+M6EnL6eOEpdnNjdeQeaZ6m/2RF+rb3QKRaF/7DixoBuez5+XyyySSWCCj9
4LK2LHiPPgZ56lESCGa06xNHIwZKoV8RZqD3VIrl7WuN68PGZgAlM4B8LzfneUpr
p5uqzFddq7kA+9yA9Q4WMMfswwlY9VcZ2HvVDTr9ZG4iYpPdCgXQg+dXzQ7ExAkg
wruwcKA7xEKEw6QoLtf0in9/9YmzEtcEQvexhlvH7F0wA2MjabxLIEqGahwQtRiG
DhfPyA8BD6IoDOexLJCV86t8piRW1ZUFvF5OizUiRpp20jSj3eQevKso4HsDIDr4
/so6b/PxAys9JvJA9GoGDAkLHz3o5LasEgW9Si10XA5U+g+V0sMhw4xj117vNm82
b6KNgfwvg6Ec651b/tN5Ui3W4EOfMgMgOkoCTepH6O2CGPoD4+q672oo7JePgycx
n5f7rPzApszgDEDP818Rxn5DatRL7BA7FGxOZdMBKCUIJL80jKNutYpIVYY1M9+J
A4PjI5Ir0hqBlj1mQKngGRQ7qeAGhmUcdhwqBLgTKZqN2OvfJdUn2Si/pGIMoItf
GhtFa1dRTpz4J5Lego1IWacxtGkQczll46ifpUcm53WbxineeKDiKBRuXsR8S5qN
AyoHszUyppV1xZtIVhSG2fVzclze1lMC5bUxBsAVxLyxRqiEV2MaMoCgqw5TN7KV
nbcZyXGw4q9b1HPPEOGyuHSA7SAA1fWvLV77zB7rMUbA+0Qia0Sj34YRnoUEq8Zb
iLUac7KEc/DxfpbE3Slil3VAcGOP64pnkDK+0+ZyrYEqzKKgwuNNoP+/YOhY/84d
nYmHVhPdW3VSpiIsuLmyirVhwU71YodX0FfrhoqJeF/HlyD3l0MWR/+tYTyViEo/
v4CZWDmULqxxUtu7GpcTmXhGh3wsNE9xc0oT+xpuH+9OSVJMeN3SViVz9yQmX7EG
PJefUdQZDAfrKxBeGHNQz2cD7yDy0r+pZ/9Qa2/W8A8GjXDCH6+pdi3xVsuDRV/Y
9RdAyp59H1GVV9zg+vCencnRr7SNzxE0FUZKX5X0G8K6ld14bS92UKa6TH325uLu
SRLovqbp93zs4tjdpyOdjkLGkiDEeYiYdOZ9FrK+C02qIu5cbjX8W8sowNjtNuDj
Y9CGZRx8ilmXl5HVca4xnGctCbaRUj7nogXn97jwiQI53xvLmbQXXOksqFVjvysQ
EyJwIHiOerySo4bOGigoQO8IPoo86imq8rsF4PJh4n0/0Anc3QA4OHC2WODBUU38
xjkCm2fTQO0wopij5uZ/Gv8YiL0/K1j916w2ahLTC6+Fy0Dj3HTXN0B67tDOMXE4
lgI6DnjAQNxgnX2XfSWI+3LE6RJzjcXdY1WD4yUuvBrXcKSCdYCIc3W/6Sw8ZveG
CGmo6oW2B2A2oYi683+bD7JD+UnO6jNRvoa99pyBaFyHQc6uXVaejhn0T39u5ibh
l3FEY5PgW0ZrKnR2sCEwWRt7s6n1BHUrRsY4rmvYh0YynspZfvuqrW+vZy5XzzTD
NVGTdP922v9tKK0kjk9NCsxgWGv2MuVM82geaPw4N/Jbww/MEPck1EraHnyWwlT1
x2e3200bCR6VpOj8rLonjWsVHgFuUQBI74VI37Zkw0Fw4st2/9z8DwrevFVWqrA+
5YmrwQ0Dasl0h0SoYz4vFOAE3L5CE4bKwJ17t/7GaM15/irp2u5Pg2qYhijejcgt
fL+PpB1XeCltc14zkFGAYUF4xqUeYmHzBUPWxfqeskp7tNXLwSBvoZhnktNYFlyZ
y8rnEyanfun7CRZH3UkH1TdfXgQZQxZ7DMkuO7H+CLRjRuHp86L7YsteOqUguHEG
/yxmuYGVC8Cgt4/3Hon2pJObmbEzkvhVzjFogCoJ8+8VB0pgxe6vaTIGeKnUQnPF
/LhU91GekWN2eajsJyxzJ2TeBk8nOohHpltcgXKh0o5ML9+8w6je7H2hEux5hJRh
WelKZUifX1mmc/nKklytO28zt7/eZn9pB8sGiELUB3Ik9wTP2/3IAatvmtwBlymn
5O32oR4eB2iHOfP4kKho+//H7r9C1cCANbVHoKMDV3E9R9vBURR4M+SM5wQj1nwB
o3dRkf/k5bqycq2Et36qfxFs2jJudetp9qySkB+Q2vPpVoTisersjU1PDJ7yg6V/
LXGOei/w/R2Bl3ijv4V/q0UvGfHNqFxN0NAYzxvlhDlTtiGhIpbFsBjVGW0cOsCI
GcE5PFsKE1oBSYwrst6jZObsk2pkciOlmPgrWAVxphHlS6i0eGrvFucXpKOGgJET
JyLrl18h6pcA3vOsltK99pAI9nU+3XJ/4kVsu9HB+j1MHCnkIBlnAlQ+2HupU50u
nTpLGi5469JQD/BETSyEUQ1oOkFBXL8VZHwh2C2VTUOfCsbhsUE9ZfBHQE80Jav3
qiI49/1QFCjIc93jZSaN9XuZ1vBZHc7OJ8KRJWQUFBo1TiB7Ujn2YZWQNS9DEaIV
/mAAvK09vXi4oUjBXAcF5N2vfcO9TlfGz84vYVjzV3j4isRLCwNQTfKn8yXfU35V
mMtBv/UfmopQMAHGksim52jVGkz8AQnIrkhhY8q8o5lapMJ9clBJBS/LaYWKDUn3
OsVAWt8sfhPo0pUl+v8SP/JTlGUrx0EHtJfvas4s+3ocM5w+HLx7IKsFNWJMbTfc
jL0kLJbApVMjAQPe5vogdzORKql4wyHp1LfaWTfrAwmpa8XXQV0to8MYRwF+HgNE
8m87RZkvFc/oTp9G0CMERSpgBRnNGrzrZIcVDIZTxtvHBmd111wy45FOhV9WbxDo
2Hk1OBYEQTR6f1gROSKaNT18JYePLfo5hfrpMbeeGiyMjk761EYDWQBvklIilCuO
LzBGR6JOyYRpmTaNXH9ySOY1Un92Lo8RjvKvrP0QJDPg//tPLDGmxL3HPduba7lH
Jups5FJmoxRn+EtxndtmhQVqwghgwkdv9/jZLJeW25nP5Vms5y6ibOAe8mctIjf/
iqXBQfoqvmDFwJZJWFBhvExF91wo8EWTwnWqnBnf2ccCQEIWoyhAvqf/vQ9i0n/L
36+NoaF9iqftJYe9JChu5Dal7IFxRSjiqXtHyFqP9avscp8Vi8pqDXLVLp94D3ta
4fd+Yydx8fPclr9YizNVnQz3M8Fb4jsgnyXQuDe3ctN5nRXsuo/M6C1pJ1QUqOG1
NB8q3/sa0ZykVIF5VIfP+OryO6W9C0kYLOU2dSFTReQR0EZlHWbbAHrevPM8P1pm
oqRH5+jPRWAM4BVmKrt1oPFGLSqSxGZXNpvV8sP1Wmnb+r016GYSC3T7iYsOl2hF
OoRCTawnT7iDTsYYJ+4HM7UdArCS2b+l6YIyA7ORlelL/+t329elEBp7BaOidPkz
zrZQ/eVfWeeFcxRFRuba34M0sEEe3+phhnoyD+ZMO99L1ZNulax9/wVwePYPCaSE
u23GSjdxeOb5azVf2FK7bFTdeHdc2CTcUoYpkZKcfaW7TNeSfLWoAQ7V9sP+FNuc
w98W0AdxgFbxUPOOthqVpaIbvtbn4iENQHktxjKiOxwsV4kRYzqxRyEK9XZ2D9qP
BYoUt9XBWeuHXE5L56eXbPcmvHdIAviVjSiXd46ntt5BVdvA1mnJZC9+KNpyakSo
/ly8icsRuMJ0uI65m0pjH4M/03GQuI+C+o+npdKx7j6ZHx3Asv4wtcZvI2UsP+Ki
QuHdAMmKtp6lyVSRe2dvoetBGFvvXg9CsbkHg+0UsWMl9PDeiCsuLSWCIshq2+2z
0XivW5BSPeaT/bVK2SoJZv21wfhdAYjzkNp/hHwcdEqL5r1TO7oGsP+Jck0U+Her
mpbkk4jpawvFOLWmyTj/jabMvKpoEIOvEp1Jvf74NN582UIX6hwkcrXEc0vXVzPg
QbswglhbIgtyeenLW6bTgUvcCHzz1Fuf7ZfAr8XfMlGG0GJxHWi4nAgIRFbts2cf
G6RC0oDNloCmFk61RK9fC0h7ue3W6Hb7Ikp2u5G0TAk0yCO55zTRDOit817COzx8
qhyO8kNKBtmJY+u4RAwAMeraL8+bUnzZvYoApKIDco0bPxDWbNYFeEGrGdC8vax8
2zk0qMEzg1sVD2aIGqNhwLwUqhmaeNgoUAGFgDjM3supE2xMuP/amgN9cH1n8Spg
ESsEDtnG8HBzVgjd7dat2aIT+GTldkxpl1f4M9PBFAilMVL4/AqsRRfKqwVmnLXg
RA+w1/JgomZQVSPwWA0a4EjzsEWpU5b8dmBH40VYFgaI/4IcXudwQ1xAj5KrPpen
xIPca/kZO4UgEH720zFbs9m3E/n7G2D3AdLZ6waa6+ebzpP08ji6ND11QSCBFqAx
uO2JWeSY3bT4V66EEgKRb3lXoj3TL1KvEyGh6YeJsqb7D8EycS0mNyEfxw8lqMdz
Q752gEo4lbXAui+7kH8q7a9BAPQdPX2yhJRvCtRClktypHog+zsOJhr29I2bvsz9
eWtBggCQuqr/pRXwAbcCsqhhJfYnk5AEXKI/qTTwHWiFH5NijFb0U1ZXRyHgXlUg
g/+vIBJAPgeyIWsCoDUl7x7Usa26dmirSer+xXPWQHhH+8zVxH6GYJ3oOZ/DXDKS
U/NyzHpoxbyxu3IdEhuv5Fx4E6iWrAaY3fVajTDNDMtFvKfWFyG49lHb54D51tL1
+KGac/E24K/Ba77abhIo68d4y/y1BmDdr571fwxymPeYM0SDAk4X2OJ71O2Qwvx+
KErxQf+bwMmv5+FsCldFGirYKy/0Wk76AzvZshFBFRhytTddkZs47Li9774bGXi+
+KleVDky6dbLIJjpSUY+k9MWlGVCkm0dYQGIyCmNbIgb4tUEjWM20/TMqMVIU9qU
pT6vJhm4+HBb67KnLySSEAi/AFppOATVee1/+3V0D4dX1rd/7wxWfAodwxkYVXpG
NwmfwZn1mTmfmYJbKlMCQqw4zx13pymwYqSqtbYq/06SW0CtT8y0KxWIsWcWxdh5
ER+7XyVzvUfO8ltYpFxk6SqX5YXcaRuR8+3mJn+jvWPhiAdTxCXbgzd8pBUtPdK4
M1GDtgEg15BEZiRwNEEKFg8NZcOVuICqlelYCo+8p7lT638+YHbsRlwMc+0kDoDj
strZ+O58Xp0imoDue+DnBznXKTBqWLrFiSGQXIZMlPd6UzveRq2KXE6V+isQUCWK
etpqmGxXhRs9Q+enQf1xkXVKPLM5z7QIfDpQaYh3iT8Q0dJAXDaymY8zQk70zN9u
fNsygYG9pH9Y4wdalHMhxv4itast/oQuDEZYXo+fIOvaWOfY0/orV1Ux83nSiRPz
vkfcFMRHTVRAdQzpktwQxPCyVDSpoBDzibdwMI8NNkdy6iARThl5/id2WQy04yWe
OYbGN+iv2/c7bpyZKL0Kdo4jVetYwbEJg72v6xxim2OzjqaaQifttyrPMHTkWivC
+cWI2TSuFjLZpX8xBPNXQ0kICuTytRvNvJrMKwFXwgEme7NSeh3jNYQI27HaIqV9
A32alCO/65QCQLqUiYSYNiml8igGqRv92NwyBNNbn2oltWC82k+EfDBs7vekm8fz
hxTmHiSEZPVis+1bAvPWx88XGxFpR0cn2fmcJav4zrFmoOd8xYoae3UNBMNpLocZ
AjJ0ozRU6P5fCRteY9TA9WNqBtvt5kf5YFnMzUwxzNbcnU6p7yUobZFl4KT7ieoj
+6TmQ27CTrbEzwqeDYCGWpd7PcAuyhaKTAscRJXlCX+Rto7l+3NJTVDrS0NrytXt
PHoYgQI8W+WK3TejGgtY2o0zaKfoRZwOwBfoaWNFjIR493vmVh0EdYLMdnPFgwSF
JLdlI9QJTElscDrDckKxDqTRD6PfCexqcTr5xmgZw82EPgk5HujE5e0S0K381Coi
nfaEzB7FzCKFXdHTuP2UJ1PA9g7c9Nz9Qx2epqrAUmGf2/yUfcYR2TH/Sr5soXpj
6ewmIMI8TZWz1YMf0PcB+iH+hAef1DzGc1yanf/yIk3bXYrz8GmA/FrbvWrUI3wK
HqyfEMldXAp0D0PmlssbcQNOeEwSuKxMc4tTC62O3BJBbFGL03tpNW6au27qyHJk
6jpR1NjJZgfzrgw8en9ir+uNuPBVs8GoRPMnj93n6gGOlFajuOWbAZoX3Ovf9vkP
h4MJTM4YeP9TUv/YntxI2q6mQrIx6HNcsfMveLJ4bgQO2bFAIlbe8rVmqR0AvWu6
iZA4tuFecAvOCe9Jr17FT/YZaXFZdtvznRko1NgR5o6J7gnrR/2KbCe8LngQFJjL
bNyXhwcK3Gu2nyvTyJpeW0qPHAP8VUEEHy523FnAiqohIgKR9MMFng1E+LqlrRuw
L5HxspxfAKnLZD3aPmV9QPJuzAZD2J08oA1ZhNZ/wZslFlQZr3c7KtdKW3WMw8ZA
h30/b+3oQGzuyj5dV8hy2OAqe5tpXlemjBY7vMbTHr7eMr67IZ2uC0aSxSpwciYN
J2bqEHIQo7PZSi3S7Ko5AvjV8o65vel++PFPRI6aTKxNL8PdEW2k+HrAwE5dc7bk
PRYdkF/EA9TOJenWeMywA6OtUqNs+rlHeMMT3rT5OUmlsd9ojPyOym8FhiKyFTAz
Ih3uj77DH7uYdb7JPyLG4xg3GFgD88+9IlfNC3zX+eAzIi2MRMm95ug3dFbjhIoQ
vq6Xo1Agil7pAQRNZGhydFbY1tvYHEIh+8J7Y3ALNwpmOlAzgcGAv7d9u+ty92oV
vVXqi2m3FIlFYOYDNoHUST3uMOCjD9nQsFLCuvMcFL/+s7C4gvDuKDOOC/c4V8kt
BCmlyFnFq0eVqlxoKtFT6JydBkDxmZP0gbIMMvdyYGjlP9KFxczv6X8IxDM7hVoE
oT9Pa0PqtJGm9A1/5pj/CORpXBV44KcObw9vXI9UGBhJ1ZL+gS/NsotUZK5W7tok
mJyv5jx4/KYk5LJgEV5eGMoVKie3dxUoJyw0quAgvA45zlXA/+4j8tidvYARsvm+
NKfU/c+QFnxPwWe0ButRflIM9HTVE+3rUL1rw40I5JYtVe8EyIOxNG9Hsc7xza39
T4CvrNCEidEqWyotjJK1avPVarUBVMutV8JArllJ3br31NEqSX5oXqvQ6c4PhxC4
44WgVupIu2+qGJRijnac7uNJ7jQBfFJgBe8oTpNVC2NyxlCR6TWWen7rbhsZB0zM
BCEZ1KBZTWmuVUjnPBajRogjXCbddNlTPD5XXRlWF2vbPVS16vy2gUXfXH9u6qEm
ste8NYhYaft9FHchAgrYYiW/Qfnk4kEPNaDkf3U17EKcSZgJDsIj9fWolXex6NOC
hr9x7U0LiBG9GsDEJL3nTmYcG1S+s+3MUhL7G2fZd+duJhzjYWjE4lXxXS+rwS68
LV4rZXC7Wd+Wa4uELSC43ZUdbbk5S8Rv7a8a2l+brKEfIpWR0T6fqt0pW1ePfn6n
S5wd3b2QT7qahBkrzh4d151ZxSyF/q7mw0QDwWu2qcHsunM3pKf2wCxqXR9TXbQV
T17T4oP0WjCYnL/LqwC1gAKaIm7FaGEhCurX7WnooIWnPk136wRlLisQlxRk6moH
wYqsjXKsUInriDWzLO9ThP4MRtoR96MlZy8tRJ94jqG1NXYBT9abXUHNx6LtdZTD
J13MjYCJWrvlxFd2eI3zA2+1jPGckkxZFiiKprY0qpX7z2LQPUpfsQuQlW4nQEyx
lQxpXhx+q6KcM3tTNHwDsXlOgLETb1pebQZ6yMnLN/FIygZzLP1ut/Tz8FoAaz4j
ltX/KrilQq3s4CuiMF1kWBdvG5i78QKXywEPZDw7QfyHUW1DeKOb/KiqLdjTmGsd
r2p1tdjeF8GVb3MEeAiWVuQYN7IqJrhugPwMAsGVMm8PIKQl1bpo39irI04+hoxe
QGQJsN8Qp1a8vo3I2Fyuf87k5WwnbV/IsjjpI/snOTa41qBDKbvyrliyeCNs+qYa
3GHMSaRnjiuB+h6Oab3yoQkC4ntx3mIgYeQwq3vYRi3rN67ia5zmPxRmabwGXS3g
rt5dUHD7Y8Vj4d29XJGqmqb3TgBI4gn3JuuxSJtidJhUKvQr1O9+rm6mf9Oh8c2o
RNHke3bOEYgAOjdM79KhD7GJ+Ehyvt3V17poykx19d8kwWeYcGTAbKKLUPqOOlH6
+24BmHO50PQ/iHMuNyNg59uA2jOeMgyemS9VvBUGZGKQWj7u2chwr7wF8UolvM7M
96ZsUj5UFtE2ODWbbFcIevP9cK/NN9853AYnPA4A6oIl+IwqCkn1XHlgxd1fv+cB
GDzxrC1xvFiJonMViSnyhUNLWRRpgJ3RQ3x8kSg4jnjFt5tayRrHX7BRaP0DOnZk
mW98IN8Z7R5PT3l3u3Ojn7tJHyNJdLKsPymU7FImM1fg38DP8h9lpmIwQUB7EJp5
Id2pg91pXcKCPo0ZX4RqpYoC3AIPXwtndrBR5kKeS8Ptz9dXP8pzyuLit95BWPG/
LY+v0e5/dsb6T8QhehURv9uyajrykrQOlOVrypAxEJp8sPULIgBycDs4bkkqMAKx
RzSMuNauMy637WgjrV+aIFme5AOWpY3oShAdr+RFYvnTkt22WFiluuG/ugknCeFP
omTYJs6qZfPwMlJVi6Pb7vhDwcLtacijauOFWwY15+4EZAxy/BajnH8wLaTsByXF
tps8S3WF3dyNSuguCfDDd+f6eJQwkoTADUzFO+lai/GQR65Mm9R6CiiLC3MgVBBm
8LIaihTdspoJaRniP8sQ3VBcQmRxoeW6/uymfpKIlIBSgqOE4vIaoWiMZWU4gll7
o6tn19mruCL9YEP6NBcv2AdDI7mjIi2BBV1bOHjq3SWM8tLfMjLbpqt+Yo5T7jHd
rWnxLgh657JP0Zmg1HxqyCOpVeZvek0k5r6UZ+lYER+m4Ew8p9Tqq+mQDqWPlVua
MelmMhi038DQIFNQkwPlUtoP2Sq1c55sThHAoMDFWfFmXtbLVdVprjBWb7mNjgby
DlwldoHkted1PInYFhmGxu0SUP3NCxk6tclEToD+/JU6QJzDid8cnGLCKmqwuVM5
TBaysj3EBz6b4snrPXRg7mUy+jFsEBYU3UNYyM/8qsKUQy75S7J/eHg7htVn2oVy
XCthSnIEB20xhUqUDxh0XrHKIR4OmKgdVwtlpKNFaUgM8bIbVKiMtONzE54LamT3
Gl1W3WgY5EezEN9qrih/HQOyuhZff+nsc29OH8u4JXyg65pRoCQdYfL3naodmsaD
WDU77Q0cGoL+WGXfz8Srj+PJuiT4KTIo4xLZIIG+D0kghKfGVC2pz8c73VE3Ky2+
WdoDq6m3JYiQpqZGIB6RBTRCVeEMC6vz6odB/uSyTyIZvBS0Xm8FMHsFHvvfIhSj
LfQ7cWRIiT7SrQx0/8g+UKimxtxNycRkmb8l2t2oEaZlgBA0Lltkj+/DGWwl3dq/
fyays1yzZwCC4iG+SPhAyRorjZtuo/jYdIJkhQ4UzpMcboXuRDYY0BMI+jyWOnME
2EvpsL2Hnc4kyI/rCrPZ6ad3RSVaWEYeT4qktGvvgBZYniPBghFc8L8fgBcXRGlK
lPqM6yPr2/joLlaGzGOPPwYFOxfE+1Hr23/OcVQ+PyN0kxW1W07VpFB+mMGW/ur7
qZfy7dcaYEac7vOwa3E6L/6fyb3pJGuftK68Go/UcQKIx8TW1U/4hRNusdYuE81R
xIyqlBf0ne3UZ2UrUbBkTdoF6X5UXjgNreZxtz2eIxYwL8MiwdL8RFHJbAlCExY7
OmIAoyeS4/sa7wiFhMakru3OATt17H0zGszFCM7xSwCSgqVHc9pFTf6DuyAP7IzP
Ogz3W9SIUgecjVI5mNea3Y22JhK4Q3q5+5QNZrP0XQqjU0KWNphMAULiBFw+SI1M
SfLGZC2neNNNAXaSvPp8kzXu/fm82khgjAVKhOnAw/zXlAyw4O5eHyLnPAwPQ0ly
QAL8a8cb6z9WWDToSqXhOJttBq5paPgrO2rOxUV+HfPB1bas3H60ykA4lfOvqg8w
y0C/7+WxoluSkpVOYxJvfzgmM0TOa2Db89/EQz3IN71ovqULutQ+i7smu1M+Hru7
pxQfK+AbK8GjsMKPDPcOo15YrqCwSIvMAP8qpmIUjySj5aITJwoHnYBV95tMLcZ3
3RCm3iKpdc6qNBWBiuTahoTBk1oF/zjHwVK4BceG/VgJDTq2oa+Cyjnem5Um0p1g
KDTSsQ2ZfXU1Ss59Dt3a8qDUXT5/P8znYnbU1LPc+U8/SG2DNlt7K3eFv7YtCK55
c9/jfmhDAOCV63tQe8mHHk2sMH20gLm8wjzJ3LIovKMAHKH2HZx6HFC7Cb5q7RLW
eAWHPtWmQ2utsiuQwdMq/3GKuOB5f9imGTQCPOv/JpKZha2ehYjQreC5oEmgWHJG
UiBzLr0LSFDhJdc+Ph/U17i3CnYbJMQTte0+KkdH1UXrXiIYdm4X5acA8I0P+6Le
tzbRwspQfDTD1nWE7/nPh5oeMm5R04paBjB5Hv6VvQ7mv38bn5y2tUtC6W/e2yGF
b0Ke9Q5BKduSOckcp9G0dq4z7fvP0S576kmO/klGd1KRN5UxUPMK3yAQtoEeoKnX
4pCgHZxzjCq4RSrKtvYJ268DNkCzQw6PkDpPteLdc7xYEmcfmkYvGLvCu0DhfJjX
yeln+dFxHqlMbi+k06XB0D/wV828Q2XWTcBaU3/eG/8h4AsS1/JRbbUay8jKSunP
+KUXoSuYuNMAsk2ZLpmqkzfWOAz5C+u0agE1dTnFCjK0lvEIdWMOmO0qrjG4dwbk
yDGLHBFcQZ51//mqG1theAKaoaYjFZxKcJM7INUEvUV3LJutN13VvPUMsGyEEMrk
SKJ+Ra16ARdhBB1v7BOZPRiZYu240XiEGeb60Dcjytq5f8Tfxy9ijsnLRHYkENDD
/mLUnQwA2XVh59lTOT7xeEA9tBExLmLw0mpKouB7nkLB9ghpvMoYKUwcTJUKqC82
yqMnXC9DYZoBEQWa8IEOr+AGmUvQ44CYnr/E1ypaswvR+GNJaJQySfeugBI1HagE
1W1ikSsJdwUlVq01tom/0l2Xp0Q/1Bd2A6ctSeZq5PWQQVTN3ijMGzHlUdRTJ3C9
TO8n/ZDJgnoRH1hiiJXmccBgaaYkrrC88xiUXBm9IArxswYBg2UtSYMYKcP0BUIX
1Vdnx/k22Iu88TJ+nIU9BCjyk2qDoLKnB4a5ABMns9F9JbZgucvlkVmPvRd30Ij8
gth3zwWrRrYk2f48FmwPQ5dWS+3C/Xkj+tcsrAD1QqOkIBlElcbK9gaC1BBFQccZ
EtVx6hj0xENNYvokVjKsi05kRFWSVdzFXsgaytLq0IcgcPUv0h9BPoZpFOc/bByq
Chop7y1rDOb0sM5nuU8Vvo6XGCfAGkpGrLX7r1TLnnJD/4H4ydgEpLl0aVM+2S3B
XJ4f489iD4RWDPsjRV11euvI6QrRYvVtpdIAy1Mp7ngVQiEkYztJlrG845iBu9xS
MudNWl2SADqJJ5eMDDztBUY0LC9KPOkFPJq39CdnQp5r0JkLbqKxPuRowcD0+6OA
7khNBuMY9jFFNUnn7wEIBZoWLCpt07YZRLhV9QqDGq/0EPtQileJWrXiRWk0Fe+/
AgrWtCtIdotL9eeMwtU8w/SIhmETqvrSUO9V3l8yGIrKCFlrC6YAghUGi2oisWmv
f8bGwRcYc/FZF4r5QYbVtFJkEi9srKfv5NsADuig1GDw71movGmbj9NJuiah8uQU
o74kDX+WohIAMnwaAC/wFqGK43JwwKo1AB34t7owaGAKPMqO5xOeHL23Z64pUECj
ROe28hUCZOudQsbZA8QgehxbQXQWVNu86KmrTmFEPTxQRYQj5txo3GL8tC+2JU15
GkytTcZgmx9dJvJGC16poNcqU6A69kSwcQ1jEtrbMy8pJlq9w1eM66mrgFDQ2hIT
lTo6mbIeLYwF3zX3wqLSiGTGygsryzLfsr9jXrJUx0hDP/O+z1iVSg91hBS/WlCq
D/PDccbE4LNtyJeiS3HsI1c4UDQ/wxrN0fcB/zhRE2a+cStn+v3037aR3BFQVfKm
7kYPdGdPJUWqBI3CDkEmuHUuPlT1BaXfm1Hpur1KaTwKM1Svzws7RjRWo/FAR0m6
TMHQtrt/HuSlyjPqkhA3+tFWeTf50mZ2FaltbSF4OuIAs9SS3lIiDvonYjJQx8Yq
LsS6wOqtMIdHM+MQsKvx6dgoN9WFpCQt3+oGnE///5ZuPeygFYiNDA84hA+xXb48
1JFBV0j3HkHj+3sO+opjNFAX/qTLEaJd3MSfjyR8aFymD7R7M22R5vKIT+W+5D/V
1tni9MJV/5/0umCyQEagnnwhlX7fgeh5Y3BPcF1JKWDEESJu12uSnNxJCbLKFmJ4
DdwZkV/sqITsSzzQzGIYd+RvMdTx26F7P90sLC4jEffSouiWvQv5Wr7zOW9UWbxe
nd0sN7GA39Str17z4c3tcWho8fr0NUOxiG6Sh/8PkarUNyOi6jY2oPWvRrKsMpX0
gp3UMDxipEpRtKQfcQFx/7k4qv/zeFy+pse/HDVh2LQ/fqs8b5WsZIGPBuduqE+h
wlKjfmUkMeK7IhS9EyPk7gb6QVEAK55amSuYs5eJM5SWmC7O8xOw7g9DxWj+4B6P
/YnO4O/VG4fYco/k3n3G28/Tw53bEA8Eqt3m+gDNn0OgsuFdfCyfTc53gXVg9fs/
AAgRT+xOljuCVPdqfi2IK+6ipTOHbje5hdTickSoiW+RLtN9o3GqinW8Y0mjHqk6
UYW6jF30wHdr30lcrmfYdHVVpDQUHEaHL/bW9Fa6rZFFPG5v0w/GTwMDsR8Sv+X4
mvfq4MFjogVmYPDlzIucgrz5VADgXlaaRF0fG+wBIL1WYea7YN9fROYIcoXX5g/c
2WLrcJF//hWgrBjPneWDKtc79nYBGlHG7FP0LyvOr+kx2lL1b0z1GpBsw1A11lNN
umrNo97w34WKdVEyzDg76RM/ZfYVcdJhp5UvtAEI7eYnjwYJm2ZPaNWkVSDHwvWJ
qwIxh7TxXzixqKeDm+lAYqApvrbRJw/AJQ4MWRSrNGXbkEds2X6NuT+k1rlrU9eO
W+xlQx8jw/9Vva0k14KJk8hdBdXZGme4ynWyCde5pAqjBThKdUA9Vpqjkx9DEfc7
I4wD0P+97TPdZ91nQTmDSRqe2qa1iD8jNBazi8fbFC+snHatJRTvpwWR9vbLc0UE
zaw/pvsFzpNX/QcmvZsiNrRFQMxeRkS85znMIZTT0RN5a7Fw5uwWCYuCO9Q+kHYV
7C+UX8EhtAGysj/t99XYS7X6gguyjQekBMZK25uy4wuGkODgiH/COv7ZgKu7ZplE
oSfMcwkPIsMAd/++2orIIxr8VRnaRMvTd5UsXwZ9wFNC2X8vwSIHC7CE76Wd13R1
h/qxxVJGwvbKwj9FvAfxY5CXw45ahwkrQzEiPXFAbxw4y5R2+P/viFapVrVuueYG
TVaCxA0OKw8t31QqNo69h3U+McB5dd+2SzvsYL4DAqZOfXIuYhvVL5/isntU+1K6
SP8rkSql1Po3ZZXrjSRih0iimKPcuw0gyUwJZ57PqOfYoSwr/kMtpEQIb7k4z10f
O/HPczqtGtQLpthu27l0T6uigkpstRGitsqmhEs3CJetlUCeM/PCqHwba6R+SWD4
wAfrAL5Byxm2W3pnDbQtGRfbtlDiRsr8cwK61cjKzUxzChOhn9J2YAo10spkEf9L
7irDmUI2B0v0xHuARZPKQSWBSym0UqcOO1ofqzB3PyheiZJC2u2VifNslYUahsdR
86d80MtYWWjSYkjrNg27s6a30fU4LchdXqA9VMajj+P+HosD/+lYVDMQ0Y/Qz3EF
qR36EQP6C0hKuPcju+lrDb5cxtB5KemCJGjQt/Vlbp8Nt3d1fh5zgVU1SAUubt7o
uxf0EV6P2cBBND1RYJg2f6FUL7MbUMYBKfIgvKqauPCzpTvLQb/y5XJ4pGdgfwzu
Kzr8ebq4KmiKxmoTIGQkvpSwHkMRPO3yGwb9zdFr5mKWhH1xMFjP3gWp9+guLZxV
g7KCzOZUpRY6tYbqT+AC4XzLUoG1LkuNMjqxZlK5Hb9MihdYPNVGMD36v3FuibJt
Fz5woElZiRhlzKitCzPsZIEDQPBRrngep3tuxcjzkDqUkIF9elx3pJjqA1cwMw/c
4RCVGawkxL0sRZgO8oR+u1E+uSh0wgA6ITuBuDfGwMA7IPliHB34uNLqic78H8s3
Kitat8mCqqHD175lQULEkX2psplTRq9tbTvIlIeYBxyUgwcleuhMcFGnInW6lF5n
++49RXjcbXnPT63UFqfGmi8NGUAqowdEsaCeEXeTgDHcgd8hG0CaKtXnOuWY2s1U
i0vYSYJr3VcBr4ksstx8fAG9RE5Rc8TKLhwhj0ZPw0WJDQyBhQzP0nX8qBa93KwN
J4rwGqUcZ2SGHu6C/uQtdHRihqWpzK1GNqgPj4Qz6R3AV7+3u/ZmAoMniEcdjV1I
Y2HnjopdAGt4w/BRZjzDVwRBa0RYVKVxFUVfARNNxGzSV2FHCTwgbbywlb44YpZm
qeUC17hSiYCtGkQZ+Xjrje6Qptjmc6BsxKQ+09kBK/skDDMxZFDX+Yf7QTjc+6vs
uSoZvTrz17Zsh7BfX6kfAe/zelvhpg4N7FBkuwvZqImGwMiqgpsCFvcd+MPzEFm5
Qu17I7R+WtyRBZiQxkaPM8FeesC0AC28nP78xkVvhNzCSdTuf6C1g4nS2HJYtsgG
gM3Yy3lymTH57ZtMH3bcdInc27l7TWLdNOsV1I46j9e5xFou9QfuPxg9ixU8qpqn
K4zMzDHYKqb7IXskzLpfQsnzHliExWQvHKUjLa89uSEjJ4wKUW6GM/zIk5GwICpT
Cf3V7gg0jHdSh8GY4boPTk8ObbGQhEQPpDRgBPFr8b6GQV2hDSo+rB5BLZQ5sDQT
964W6WjTE7LTBhZDB2xUFVV/012x115D3CvQtr2BwVFXeKE3qcVwCUe/bbJ4vKn/
9buW2VKaR3uSaeuy4IB3ysnuBsqS7qEkF0IrGtppXg0J6uKIUYgX0pUeZdmep4DG
qbJFzq236y++Z7LfUAmtYBgT17daP/ccgwBHNGPUZWuoGmre7aVdNF0hvtFyMtc7
A6F0wpW5CRJ/xBLIX5vHhdDwY+7gWrcrOjxtDWAY3XQ6LVIsiR5mz9KeoiFOJP0X
bbABNhNAPpZq3F74GOc5z3+r6gY33PYu4G3QKpaFpPtUu0PAtO+6LbRFRLWl/fMC
Tm4B6h3jpBFrfFzufOrxl0x1GfIYyIGRqscfMvl6K8+mrKZ69ezYOjgZ8rKjawTN
sZr89GGq+a0mOEZPHrULktyCyF2NZR7jLhEja8/JX7eVqZxGlEmEwOkWjH8Lx7CJ
57Ck31WQmKJyqCtdAzK1/7uWVZ+dBoTz0HXTFNdQzz1XgCCgendImdAQ9NTWQGj5
DzyIEhMiML2W/CAvPXesR2xbk6ehIRb+svUHsRktCfx3DNuEypZHHDjImWYCfRUl
vovQA0MxCrn8rtKvVZ+ELTMCg3C/hVyzR5ecqypkNlRlsG1YI3JT2XNrZ9da56pK
6ZdtaFFo/rtNYBhxsT5ayYQ7qQU/WA2jr6aDQY3EjZrGUKnlSZpv4lz4BANqPsvU
4mWDvwCk+GdlDDJnxcp8YFGf9+HpmsnAp3jUU5Rs1WzvqTLhkDJxaFx/R9j6MAE4
EGZJ7gGirk0nVeB6qSLnych4A54kuouyGbz6GL7TnANQv0A04mcIM67MZpWuPFIr
k/QbNHR9fFMRvWxr+j8/FCenHhY/o2Hg7OLBl3ei+DGdeU9uYz1aP9F/M+sLC8dG
E27sIOWvTGnJmjV3YcBgBp75lamqyajjfcaDk8O5MZov45FacwjqKJovkaWYvxbk
avmi2HsCghFs+8a45OksMkwe6wn+FlI8XU+2S6XaUsrzhRQGmHayEk/PuqEoAfEO
nlSjK+nP2EP+EuoQZvP933VD0KRwhh8JV3NaDiZ3IEcinbAU6/EuCckLJRTMOyRU
RRPnH2YaP+4AYjtIg+drBNjCO3NGZ7ecG5KdRJzG3bsKxwXTylwP4Gv0fY4GE0/N
AOQ008Wd+NLWEe4QeUjAdR4y96cDorGI13jiHehBrmaFUkzry1Dpw0ZG2/k9aGW8
RXlJICzNcFO/4Onnemp+rs4tLaDsEqMRnadCfpMkxlkpZVOfyZwsoFZlo7Kp0Wqc
inow+L5P1R7o8GauG6c/SIpP/ls1wuLzIm3Ht+4mZ//nJAg74BRUb8Jfih+c57//
aCwPYhfnVjgg7asItjxmIxvqEPK+OWsVy1iU8km4KaJk+GixtTWfGjFua6zRyrah
Os3RQ765wowVCFYPoeY7oDYvSBT30apvF2YFHxeg7JVBIjQJ4xBkerV7FpTq8p7W
osvV9pBFMd6pLw7PqGoh9M1TxPDjxGSI+f+tA+qFFmyuzgw345VGdcwgZaC9CD8N
Mwe3+l2bd/9XloR9jPhzaqw+tSWOl/2EUfEH/WZd7vfSYz0fswUir/cl2dnumgeL
7xLqiJXbCEKYTmbj6a+Nw0l8o6X8v36UbpFHy0BTXEoFOTzD1fmI7NkCksBWVuTl
Z49cD9JoxaK5NJz+Vo5W/ADKn9WtTSLkaDZFDAmOV1ZithoGIPAA3os7gq3sV+2D
If8ndJfL6PE8vp7KQ4Mc2Pf9eVMSqnVBuoRVH2uAJ7ZmtU1DjDsPCNywmV038cM/
QPEV/6cNKFLaPUsK1JJPbaS35L2fK4W0McL/JgItsBm/NjClSVmdequcwZ5S8jAY
MLLuNkcqneOe8aQDiyo8UUDd3IHCN4YIH7MlsJ2ZGk3NZ1KAW0vjV4CTdqa9qkvV
nP/HN4iMSrNtTD6ONAc/AONs2BANcA2Mu5qGTARbalwoj9m2Fh0KRiuL+Mr063vM
YP11y5Loll/mdC9R8Q/1H6Hkj23/9TSFyuCgpshpJ6z9LvNHq0POLTTioxU2wSu0
Z27LcKK8ZpU4kzWgAbsN7hYLQ6LOdUjSpqBT9rXzfGT+H4f8w8ck1WsNVnX2J3a7
cHaE6FlEXrs+qalXb5lYp9mslaCqof4eN8+Ga6DjkfVzinF1Sig9Xa/u0A8mh2aF
DywUaYobbdHEe1YMCKToAsq/LmGzHIBZ3XMszqCoGrLtNc8k9rjG1SDzJfjnu5ng
iV1nVEZ//EUjLkOurQwTTMsi6NY1puC+bg/inAxQw3eDT1bSUrQjxHBE+H7mGC0Y
NXIehGoSvRCazCItTx771rkA+fUsyKJO6C+pxyAtB6dHuCM45Yr0r846nQ2ZUMmz
V2ZskQR5RdtOHlvtV+MUQBExz7j4lwf2VNCW6ffaw0GSVgvZyyZDWXn05F2UNXJt
2sVkh1uMGeMeKTYjTypAN5JAjC2erQOe5Rkj6V7mjrODVAwrYwdAHHDIHgg1+/87
JGMG+EMMPw9O9FPZMXbiZZUxds/BBwkVBf9WprO7zp0uhrNECAlxjn2zkyl4yrAj
L1b2xoY6nEsSD/nAjUzZHEmGHHm51xgQoMgOM7SB2Ik8JFbpwQ4MCZdygEFSPS0S
11vfcvTdK0Mx7F1UQ/LlsgAGMntS57G1mny4gyetCnqdtWp5Guhe2HphQEdH8u0i
tsPQ4OPOuWNdAW2Hg5YSC85/uS+GTYz4yPF2zsCZb59lmy0OrNyHDBcJbaZ/6QTP
SScykDBBv03iAuW24LXreNyXwnAIbgYoi6tsUpQLmu5YxVLcQwBRSEO937ajMEh5
8zpm2ohC5WmwTf4pTiID7Sd3AacDEk9a+gqZKfdqDUpYBKouSZUQAYBoX1Jdx9/o
cdeVj4vJxo8Hy35RygAif/h2GuQ8W6KdgyLOu/lvyRH7yHlFyPxIwgptzrikC+jP
1SP3ri8+TDmJ5YxuMo3m9UY2D+QE1hBW4M11sMPUtMzNuHWSmbM88uXtLqeyPqiV
aFHdG+LiFKj6osAzPO++Wxal3dQgJ1C6F7GlpEBETfPwI37RR26jsVGY3odfMpLS
0SZ0QGuIsaOUHJbC7XzglBU0ciQPePMeq00wWltwmgMgTug9mUxgsG8hDB9gc8c9
+ChTqJLy5H/tUqR9t6bmF0I9SH9TkYLGbD3Q8zWO7QHjicQWIJdpaN84HaxhNa4H
p08PETgqKxsdvKQ9+LfIBv8gafgj01luqxQuo60D1dleKsNXxO03emU8csfbx7dZ
tSMjrw4Uz7mFhThj0XQr+YnzZxFQvOqbOuH3RLUoPlN8m2uINvpCS3wvkRihX/kp
lecCMWkj/CvFylGxPWvc27jjnpbI/9F30ddNuwyWW4r/GQbiQ1QLl2HY53feghpe
H5kpY58A6S5B7KtfAoXAdRSRLtRUdlgE/pyzrQBnaOvArGTCNT8TUnG7toP9IqVG
my/sORHBA0AYWKkUAO6pkEriC8QWXezFYA/2twHsFdR3tQD6OEBGIkb8wByWUAls
Y7R+8I5ZeKB49Nm1bABA3Yp4bMz5s04Ej/mw9RqL3+pKiUc+CpwomvXzB/BS1jzf
ProwPyVzMRyruMKdRcW/mOJdrCSm2d8cQ9kLTlZMqq6+OxEmVhUC/7YouhV06/Dk
/ZZXGYtyJDcarZepgsqXxtSYwjffTU3r7V5IGlSu24UmkFiP4k+lIKqZH9h3R3BO
yNkPr4gc2oLM2gEoSV+w3zvYS3+LBzmegownQxoOm3hsLn2zOQqFGr50p1nOqjNs
eNzTJbEV2/zGc8tQcngSigBjIuD+hMxb9Euo5oe0ynCvAumvyfBoylywxD4JVY96
y4uLjl5kgl+XeNZyB5UNus9HicYk78x3jpKouEKpDWpgw7PpcVYOzSOn+lZIj7Rc
up90KWp2QWfHK74GBn0TP/JJLgEP7Uo4cLPhkq3+krq1VDALda56H15iHPoFbBvY
3PPOHXYiZddwMVMU6a6xPfS4PTfh0+r1/HezDwGsQypbll6pQFzElUbYkLDaL94X
yTcSZOft06VTznofcDvLSP/YPzokyZCTEaPzAJV3nJWYG3u+AW74fRYojVMW2VX7
ci5mfp1e/BXuxaMhz07REAcsW4DoSjeoitoXddbaiSFrl0Hmhm1a55BducsiT5JR
5aFOT4X+jnrdNtbQSjk7X0vpsn8TCkhT3TKO3ToaNDU25S68NZRqWY2UnvilBmbP
IF2pKP4BEzBRe+gP126xyU7v60S/R0IjXxVSAWoL1hnuUZL1VXTSehp1k3TNdurn
nMnS0v5ISa3/oUjHLnNa/FrRvKOeUQWjGASGTj3d9ZC9Kqd84BUYueftwQNA4F2S
wrWnB2gH3bAau1oebvMqY0msnjCkTQBfTRjn6/s3xDlX5f5TrSyBZgqWa0u8Raz6
klLnR5c98otLCY+FexzjgxVOsLVJd3puXlxsWDAQ/czX5E8i5leF5RPUPT4gGKkq
bIOHsS3vyEf1t7bJfQ+D/wIsXL9kOru56DO9Y83A7vvSfbPFlQtdwPwAytYidQiK
0QbteI/GXtTVupPj2eFPGx0QCjvoyxKFUwLCEWjH5XuY2cnJM9Ic/B2fj17cCbj4
M9gU4LCihXjJWaRUKVJXJB7C6M4AIWgxgTTSu1VD2zr2gr/wPxTWIW7zFRW6oGcl
tUfjLnTxWOO132y7YFTScs0eVfWyndpKosgm0iO31rvP1EiWY0+UY6GxYFPV7TRI
wV7sjrrROJK6oWuH1/JpzJYuH9vITLUvOz3A+M0z95F5gnxPnghFI2hDCXtn3R/r
BKycsEiSuN3B6rfXhLt1zpxKzmnFyOahmMTNDayClbyv9RTSmdbvFA66XmoZiuRd
+zdrchcRPy3E1l96GqdLySeLsubW3kaVsGOuG7YjaNRwUlr7D12FvZLnNnPdqL1T
5BxN3iVGWdoVjDlrccLcil3j62UqL6YdnPX4gJ3RDZt3Im/VZGMySGfD725Mj/5t
VABX6rUYeoASEt72tT2QzmAzZ8ChKXnCvz/+tlZWi/aVDD2/snTHSYsNUJPGpglJ
DU0atA9Pladv1fULmFQyL/ALf7s29GU7tY3ZdTI2HXlDpCygbA3KplxeE6zCzYVI
JdAIxWciZENL5520FsDlSR3OlwQ5HX5NslLHSSaBdctoJV8pLCLKEnvNXdFtHLod
1BO8C9DFXTO98yd2F4+N8/wPccZJFaoadrxPK9rgFo3ozB2bDQj/A1uiL8g2hxbg
KLxWzHsnQxV7We+QcduT9t11QNjB8PsCxDnWzZjs6yyxhdihEz1CZTXcy44sVVEB
3xsq7AxovHogU2+PTeNoE5n2tjLayb5yEFJp6rv7SW6RNCRVreXseHggl7h4K+WI
8WDnZm4mnuhpmPdMuN8w8oRlJ5/H+0bh2n3exxMjlMlVkNr5t3rEpkumNCydsO9R
9j6a5M40u4V8txJ1wlWMpLIA3eNgN8bqjMoN615kSMLzXNb4TUfMwbJco9xL7S+Z
OHuiH3jBAmMr3URhoCi0rQmbPAq4NnNeH+ZYYd/kUdRsX4r7eqHaw0oRoLwxTh0H
09bD0aJqrZctW2r5xynC6SimoYHE1afH2W2YM6QobDXfifAm32nWY2E1EN0iGcB8
NFiCOYgWrRc4FjBjod6aIJKtaaecx3pN7xWRB46ZqXXVneoI3FpA3vMJTwQPChHy
qy1ZOW197668/kBatJsAfCsLwM2liHZM9sCMLq/Rx4edCDal4HpuyWK6wWtVX/zO
86PKCs4azXzw8dEL0c1TU4rBWFlVwYHPUcYE+dGTKhEv7QpoWqeI7+yEVnrxykz5
AoEdznwPMLGqOqAnjoEVOa1eAxsJqG7zWM51+YuTvB/R3Zk8XtvepZupXoe24pB4
LTx469g7NCuHxa1u3o4LiXQLbi9avlTi5H9LuWau7IVSOQh3EcD2raux2eL/9MJm
QCLd+pY37PaTgsi9816AkJbS3/wJKSnUk9zMtoYOdqu3o++Vs7NwoVulqZFi9h5H
/9VwsvUT7YhVzq05wRvqbHtCrdiX925SkFCJDR5tBN300073ZL+nO9hWfmLdbmj5
feB7XGagfkmkDc2fZ/zC+fdZgyMiyPg8IFJ1v0sDaRfiUma5I51PADw9YA46LQFY
v0zNK9skkCUCCCw/xOp82QsDtn+scwN5Hje2JA2qTDyXt07Ft9ZMhUvX3hvM4tbD
/gaC8VOM33VP0rJt4/uTJkKUnZEoYetC/czZATErwqyfcUpzks9TvjiJaZnAaUVB
BklMZhnfuqSW1SXjJUMCptiwBa4dDcGl6PxT79dAqhbYSXLH5Tea5p2+l23NMp7Y
mdZvDP4Ppq7MfVHZAFZyN+kL3rebWw+Xwmp4JzED1gDNzDWPId+AozfO7Dp9/1r/
IyoYeY2ybY0sQXHfA4gfea3JP7rfrBOlKYLHGr4945hmsVgJKOjYO+h/EBqF4f5B
S3KlpoTe37HoS9jFFbeJDRVK1n9Yaf/skG5Gikt1B1BShofuC0kxSxnDIdalLYIJ
fCjrGs7glmdD4G/Nln7C7KgdG7eG7pdTr1HRtQHwgjhuzrVqE3f4+aMExolVJrv/
ZTetDCkqA6rNOb1kxHU96fbYtDG1vxOb72gqPde31kIh5VsHL44ZBZiDjh14PPlZ
h/TjLADOL+4r6kzhXMl7+alnUAEB14ofPH8k9K8Pbz7s3XBAMFsrRpcZB/TmQOi4
K5ye7KjulBW6m6B4MWM6bD5kq/hvhI0yE3KeoAXqOy2bjOZLakIxV2BTlj6/UXiS
ryVFnwWb1JA+Mze7EoYNF3imXKwlk5U5Eglzq3tuBZ9HCP5VchKro2fK570O+Zf/
Bnhv+xBliLWVxcjd+v2wB93031IlQIuVMnGmJ8XkXcNridQC4lLVTafwFw+GiAls
+jFjcIm1s98yCQyUdd+0hmqSjOM/hAm1/fmM+0pq3MGbGM4jTqAN4gWmH/Ul2kHr
ybi+UElwVdWAnE+Dj4qsYkFOgfWPIzcyRPM049PW3sG2QIj7P7xRnwRW2cuPNZX4
zX8jLnTtgVWUN08IgowzbjhEV+PBT6Ysbtf5SyyoBmFNv0xnYUZrIV23cEXaQ/es
8rFgzcZjLCfYjruo+D6FXzL4+myILAS2TV//b3kNKupf0b8pphs1DL3j/MTyEvEk
z++Sk3e7EtB08yizZHaYIItbsufpkXtTTR5bMoCuO/trBM1c8l4Qf0HTcMBplf7w
gLb7ctYdWzD8pGldTsgxWol91Jsi603TTICT5aHNRmM9mpG14QM0T10y1ayEsXhc
FPGm1v2SXmfxmvRWBU6nfEat7LdtHL9Y9Eaa8zOSe4hQ9HtB1g8gCGuMdrvUvC4T
ky4bnt1dHnR7ju1ZpKTh/SIjcJDWZWp/x/Eai25Hdjl5iKEGxpcemTKww4pOl/Tg
N3XJTeltb6f8XKPrTbEi2W8vVljOX6e5RRWzdmm6nA6ybLK1+Z4w6GqBx1/D6Tqk
Ea53YixWOJEdHh9vDS8nTCjA3jaHM6XNJR2AwKeJRL4c8iGqwNVdQrGfSnYh/Cs/
W9RghHElAxl54WC+TdCi09BfV8BxgyLG65CEs9hCKhHxNQWYGS3l2/UvNlL67OyQ
l2vA3pj1lnGohUXlGRAzgDmS/Q6J4u/B54FyVWargW2XFq85nAdrH1EVdfwLH6Ws
3ghqfzDlRgkS4Uu6eJLhmuK0i91AtP981RFfS1Hr8IIP66HohOPu9PLBfvZqLShU
rWpVKaEvplOlabAy+EI+9pnxnqA5lN9yCXOs2NmckV2kwvxGuYt5MWsPWuGHxm8S
qu7eUbkTmbl0NfMfQ37d9O5YvyXKkjnpuYi3qatKCxy8o4oPH1oE0+jFo/h+mmhO
T+krhwPWtYFQleBiqGfCxvMcE6gHAi+QeTihzfpcvdIASFl4ADUUWOtYa/IgkGeD
w3uTOkgo4pSIosL3O9sD+BAczgT4iMSK3zpc5pyz/AML0JFC1QuD2GtM6Vizs8jc
9UMtIHtJYnScdr5AFr4M5Q+i3lIVpMT8aRNJi9EPvDEO+uf6osUA09Do+iPlszIH
+GXNxRwxBvjQEBNFxU92Ls27xbo1Un+E3TsAGC1kCZ7m1032/DPHRUUW1l4XW0Uh
yxQuj3TqcIPGm7HZrYIMfEqdQXQzZrKYbnL7NrIvQIPkUIIrBp6S0FhlxNOhZ2WA
SswlVhqe1go97Q4HKvAXpZ1l3rCwnxnannDl7kn5Thyw5nanXqKlvZd3pmSSmSdE
hrvUYGitVFhv5iuuOcgZMG1/m49v81uNUZhofyF4yR1e85TNjMnRvEyDXOcSVb7J
YTLodqVPD5Tl4cCmteNUuRH4zZZFqhjY2PfDrq4wXTzXWjYMAZerERZd+gqc+zAL
P0nkgDeY59ugNKLnH0nkYaQRRrOph7ErYBKiD1FfGOYiggaLB2UR5tHlM71pEs4g
+u9EHj4wskL6vRIrT4iMUfeRo9WEYN7SRP8tUHZ6eYdIL6Gpn5sD09yZzZ5MpYYs
b4nEB8XXt0yEiD9WjL6crNE8s5RzJ1G7rwrTEyenB98JzjJAVb0Xf8HNH281g7ZA
L6TdlTeZIYkJA+JJqo4gy7LJzvsTnQ7DUsp5ceJqooAnlRh+OBATtQNeugfXyRwk
glmrqi4fSNpQAjr1NX+1xZDaNVlSfu1YX7MyQ9YMz90dZAdQFFtxS5W/CK32hh9R
boMXdYWadGym6KrYLg3kyFw/3Q2ZRZynOlgIFLmnhd0ysP2oLEvZhB8J43Rv8stx
1mJA5k8bzzLUrTa0S6Yc4RWBZGshiS+0eC7w+9q2aviSqsQJ3MokSMApCSupx/85
pmuQhuhR8MKcbVB3OaTpbTpJ5OFnkK8OE3zu7yWSYY99J+VzS1YX7afpMZY1rc3d
ThMGcGhJaKQtFP8hPrpYQU1ctg5rBLkJoalHef5P113UxUnzV22FpuOLYQpcOVpD
dhzP77tWJq4ghE0rwyqKoF7t32dUbdhjLJ69WKnD+jPVGMa7EZOgl5PsVm0gwOJ+
HgyBvdeP5krJUm3ZBe7TVdl4KYgfQzSmihaygkPC077upyeL0v+f+bDKz5j/lFkA
ruXbUFmh7OIFFG86RnZmQfuemijZaE2nQ2Uh6y2cBo/sTfFTDzz9MRw0+oIz9qxf
5EBUF+OQOCVqXBNkfTiGwBBJPabmg8RG00Wo4rXOa83elYlQdm9B0MY9TJXL6kFi
YeH7vJ8Qs41Gqd4lMgRVAa3gdIAWPEzgIFvURU8xk2VAfy0dYQJy4fhoIruzk4eA
prKf/qJVmQ+lf7Kvr4VrZfPJRVTzIkBzRvwgLNvTgL/bAJuWj7PdtWfcKCCMrB3A
y04axiRPxnTrp+FsIoYTuhPln4lsxWtYIjqU1NMcXNSMqUvNcbZy4CNHMpUkzE4e
7j6z2OlX2EWTZBRoj6+4saNGnEFaPGaNz/KX913QopEt/LeS39/Tbaaq8PCI763S
pO+tGV7PmTOYmU8vWqObWuOetK4dQujWusd040WAbAHmYgxZfC4X0eYGuxtMXXR8
Cd31FMX8UM8BFXarNosXaGYIgOWuYfADU4om9au6L3j3kZ8XexF/41LN9YeQHjE6
Dzb49l/zZJDNe9V3OMBcTHEYY0Ym8ibIm1cu6htLdIl2VMWm/V8GGcy+uYM0TYv0
vNAqBhExOkHKnNtY5znZq4BMsfyJ6OdHpuMe82falczOseVBMKyQTyq9df9ktxoe
tgq58/1p/FpxiMb/8E4L0jVUoMPYPWDYc5fbUKWVpfkl9Sn4v/8o8QhX5CZdzVgL
bkMUceEChnogrKLeDCmt7qelQU8PDJmWpI8jf9GWGG/g7sH7VtDQK3bSIfrLTzeT
h7EPmj6CS2yF6eT5zFAySJt9YIfm+1gAvfwyw1vrYQlLsLwSLoQSyTjHRpTi0Y1I
Jiaciw1o4Qtw0lgq+Wd1lX4nJLgw/B7Vyj1WsPrPtDNqBBTDEyUta81LOhxqqD9t
wB07xQK4CwDZw2x0ujWE/pjOmezCLNht81iIdG013qW2IBHIJJRQvBB888j/q37+
h/33+6jLzmAntK7O4AFSNw/qGTkUGiS3YP7fw+IqOzyrenNo1F6FMKTMRcoYJZqd
OezDEtgu9YnxF96osKFpXhmotskG0uvLqyjsS9vHNCgVz2WpzJBI01bQIyjfC1/k
pMHlAHJqkHjgImzqf+Cnzr62tmx8IhpglIqr7udqhsek7ySaBdywYDK0uZRiDz3K
bmNBsCzvv8S84nu9+89ENSvIpLqgLaSioNMNoOuZVjJr5DmYAE1PiKPVNaINYbxa
4fdRDBkoZrWkCl5A3S1l8VPXj/JcA89yULxdJJDhJtxOdD6w82nTtDd9wc6iO/GY
PfgV8S3qLaFu+pw5U07+T/E1jL/OmMrV+cw9ZL38FYXGXkP58Y2GAFBSrhlQT0XZ
7zBgiIjp9ZuweyuBFRGW+dxj/g5MSZoSj6/v0erB/omBtOn4uPWzYF4VewtwCaPb
ILUyjHtJzPcDE04Y0Y7jP6LtDCNRw5eNptdAYdOc/2m382TfpiA+sVzFBJD/nJTO
7igtWuzTAnuOBd435MeaWT1xVIjjg3PcwDkJF3g7/LOE1PL5DAyGpeoGzxLp3UI6
hnVP3Ygkoe8EHZTN7hJhUv1akarKqrOYe88h0w7dZZVd8Gl1wHgKwJ0ta4B87Hta
eAhp7Q5KVzCLJFvW1pLBWIorQ/e67ftmw0R2iwtTn4dwFJVjeQ5hicjFgx82/vyo
w+MS+1fusHeenPFgx+dinLqdKuzHc+n/KG79ao8TaY71tpeNYROcUzGlNZi3eXmF
eijLsOjxhBv5MSciH9/U/ddmVy3czrdIAmNfvoKXvzT0DsIXNExfuMbVmdDKYd0h
iNo62kxDYoywzlKUUGR88Hu6ojSLS86+o8EHMUNntI5VjR1TZjqEab+S+6mQhPCq
hm5Af3ZNoJ449VkHkuPFb101KSM98Q0o3AIujlayuTFYXQhD3awoSvysD2xSvOYK
Sh4yeVb2NX5XZOH7SRhSX6x+3B9asNFsHYGMKaiU+UpA5zEr0/IN3rhCG/z5muCk
ITs9asD3Plf3StE+Iiktmb6GCWME4eGBe/bEYFT58nNFevZAOtUTo5RkBy+2y5+g
abVo6q7lNKwE7ZBSHZDW+U9ESmUvPgbb96MtYI40JXdr8w0seWy6b/WiiqLWPfeT
8h5jNnalehbnFynUFRngCZC4UE/siL7uZvZVfdv/MOYO35LLnBh2im94DYfwkANC
AjorXZbDXvMGghBVXdnytbgDTEikQp9lQDsJf7UhtCtmo1gvyX/Jykf9RlJQ/P8S
lxDRRuh5cI18pkZ2T+Ygd9xWbCLYyMFZv6h3xdorRdp6Jl8JawRusQDClulOQAkH
eHCZesUQNO/UCGh9FpqFdHUEB7Kx70v4YaAKR6w4NgIP2bSpiUo+RPeQ1gN8wLWY
uW1/ZO9z0geqb1KikMd/Qp8RJow96eQ0o+974nLXsdp0jwHWGGd55xSPwSzJa7Zl
Zz98hqVCwRMX5tc1rukGMKolnT6OS4g6fl3slUBwf6oMtqse1MbyzLVFuIBVHmcI
xufGo/9Gz2ZEs1HQwPWs5thgtYi4KIeyZSZvTnBpowGrCd7I8zaZNBwPQBKFAes4
boOMLKmvj0nMdNiEISWjHI995d2sqiAFTY2wBxe14yp+dkxRAhDjh401m1PK+DQn
cR57eOZdtuj7SGoD2ee83OQUB03i0yN6Drgeylir5HJpJb1CHgZkk+z3PiS4lkjM
+e6Z99ThaZRGBEn7lpQzSDfuQfKdIuvuVX19uBYJBJ6Rvz20FRWcj5jSwaoOQ9KE
flQE/CkLa+x5rXj5ZIZj4hQs7yy+X024rjINoqkIRndXwyyiLP4mrzf7aWGlgNut
6nX+cjDV8AsYbxXqxHA5DvPAYqL/WY8IhCs48tOfYUmkA9G3ZHZtfS4pw8JBpOdR
aC+TruOPHBqxBozYGygzXxkuEW8VmUFhd79msfPvw3wectoSy1jGUYtjO2X5aSvt
NiNBxpFD7thFqPsw5jQUdLdDJ1k7Qf8pgCRDSW88dHe9oZmQ61LCvnD7ZRfzTBDO
+5ci9zNtv+8Cpig8Glfx9ZaW9xenNesvXWNEcHBQt79o31dNmNRs05bmTYBEB2xo
49AEF+YmSwBU/YRL7zxH/zT7EDUWEY1ZucRIBWzkhxeCpg13OlMaIEGIlM85Qzze
5j18FGU8MH1KEY14Pv2x4l/7ltbKT/g31q5PWxyLFGNVwBr/qNUxO9L3O4mk00lN
ys1egUKIlLNQeUxnrysnj4Fl53PflineN21dRjsucn38YKC9E3D9Y9sbFpwfdRUv
bVxKz8sceEaRfxDyQXY7JEYusohQk7UZisbrn7WX96pxtSgSYfK+Ey1xeyBrpLFx
rogb2x0Ki61cmtw3iVWq49Y4hfeIfapdc44LJRiCTfAD6FR15CzJcuUuX82e7gJL
w3Irawgf+PO5JNOi+fHeDajlIVWC3rJ5/urmcgjNznTrb9eAknSTqPFfnW2bREIc
VJWensYmd9yBWxYzHe1BRrafpsWYoi+FW8uUrWdZdz9lLCmOO67Ne4kMSstF79d0
HQJNhMVi1o8snF6/ufgaR/ucoeAKj3hbFboU9jGKUgcnLxzJKUGe/TvBJmAwULY5
kQDNcDBpsEFTU2ZsMCWx9ysfa9gzONywgpjjLW29gbs2rkMFFi3ddiWQOLK2B2wQ
5cpn+m7D8p0XwECKrTEJnlvdTJ1X+Hx0l7EJTYTf1/2fwnvAhL6+q0+uWrWbwl87
sArPkrcd5nM5xeOiz3vCEzFK2etUY+FVO0/oRsVlzFsDziAAoXbeR8UU0/lzIMbm
DbHz7Bl6m7wqboXu71XAtgug4aunYj8tKV9r0HAyRRp0NJ98ROZuVQksrHORgz0a
dXLTFlU+EW0XZLbZtl/iZXE+oT1YRhtvQgzMuLdoZ4YGiVyCYRHN3MeWrtlkP+1L
Agx+Pd/ud6bkVF1Y80XoBmkLQ4GAGxdSorojWYlPsMgl2bb3s5WgmUR1VcMPFsRa
cPj9CJWlIQ3Lqtg10RX1LeFpnuBcdPq4BwizpQMBHSlQEBC/fwp/qJUJseg97Qjg
ePECDZZvUGgTddfj4U7QuzbtoUSDzCzP0/X+vV954YQsk8OtY8zBXswVVNUFY2Ti
SpUa+Ici0UBHhAqcGRQJSiy/9an/rp3DaUI2IndZnENH3n7Pxc37QStZS8r5X9XB
gtZHDmPQ8pXdXs2fd6+TMoOYTPy0f4uB0tmmbIl2a9PBRf3tkmmMKoj0TkCcIKG3
BTUefmWT8KYY2G7XnwVWlOy7DFdYMDkCm1jpR3cwalw0U+jxp5OOKyfLahbsiHDf
NWI1Uv2ECsKEV9hRxL7GCXWl/2HyzIk7saEpcsvlRZjbXCeNqwhTUYpRvDvoBIGu
yWuvDf35FFKsGyh+dadhyGmfTxeaEpLsMudsrj9TunSmkJ5Uic4xb/yyfumj4iOV
G8qKpOR6+W1eowzhII8K29yBCBxE8Aucynff6MhwfhBHCOd50V6ayojP3S7iHIKR
sK+MBsWGKDd4+mJBkw8ZOioxNTaELvRxxn/9YtioXlTZtcKEW+RnKK1M0PRwWy9y
HqVMSnWUNl7JvdQpilTfCVT25BjrVDSS665YlDreFDy9i3Aww/X8KqMI9b5HJ9T8
2nH7PyTCegLbHkNnXWZSIfIVUqY408mvH9cRObrzqtgPDT+vhheYlgzLotUzszgX
ggadvm+UGnIaoDsWLgNt827MCddQW+KMolVdxt4sIe88yJ4/TJEkcBEi3zueSSoz
5kwRTbT/RAAkpzs0tIvhX86HY8ukakfF6laj7+mv7JxmZg4CdyvC0ZlP0l1SE+AV
nL3K7orQTVhpncO+ihIwhybRlIuV7/vLVWv4AWyvOQWuOVuL4wHSiv5ioorFfERv
wNkP1ekLJgtn9DKB8Dg1EiJstyoTTxsHYPb/JMMiQMbxreQ85vIsQ1z8+NpT46L+
rCGHwVbbQBrRsEBS20GJUEneAQQu7iRJqJ9SpDJqGsPR/N1DPd0jRDIZGPTj5ANw
kT6Ycc0R21WyUGki8POZIdRB75YJiX8ntf9CA1li8JWjUG19gTnloEUnqltnwmbI
jRUW+TjeDZtXGenA5aSP6Yyd5s//q5tOCYhLPFO78FbZDVtCHEsld7KL0GOXgkpH
T2OANjEIPVEnpdh5GLoQ3z2uKD439ns8JUatBrOx2BiLKTqENJCKeQ03wDv8GPAO
rFdSLS6Z9ti3eM0IT+2WWM6QmwOVHmP4kutpLItdW87YcLtvZTrp4C4GonMszp6t
KOZAQ+lFBawBqKJrsz9OgwLoolAtQhN51GP2G7kIqsWaxmGR7xqnbNAcG9xggnQ9
+DIGci74uKlGc6eJoPbrC93DbxGMYn9OkkwiBhF7T4O1hYl0gg1RZh6CYSe3qhbu
hJ9OksYt2H2/cpZMAazolJ40awYxcvk1HGr3ymnG67Sspgh1f3SrwE9wnC9dXubm
kBXHKK4KLZICxqRazRCF8bRq+G5pZozGSNVlCnJtjNofHKvXcpuaa1r7Mp5GYStl
8gqTaWpmDQYyeVZC79Ar9QYipSjeqWOUkMcYlnq9ExrOq3YJIEfX0E262+BNz1x1
Og6XWepnI7WBNwDHR0ZwXFVALG8MilA+c0kPlvbkO4UphAaE5DMdnBtuRR1G3ZWL
PpntDaaZHzkZCplegaW2cm7iT1rg9f9+RnuYsMJtbIEwcZooPUhn0vrPRi5VPjUj
G5lp3tlTTAzm5h4IQoDJcmO9AxheQ1zUhdKKCMeAKjH6aq8c98OjYzDuUhGR5PNJ
NijO6RIY7uF5JB+wls507NtnPjmkUb59aPN78jsRk9Br3/WIGY9fQpu5Sp8TpB82
NWOvWO058B3DKWIg4E7tMvaytYCcy9I6YRFg7ghpTcW/8S3JeaTdQcKsLePh7aFG
rpVH16ypAPjB5BpYGrVHxP/OH58kmwhtzDCU/MYjpHX2i6Bx/jl4cUEWFmvv+WrY
HiWI8Cl7tXuMEgnT/vklhrV97R9XLxxmVK1FLBYBf2gw5ZKqIpLByEBScTJkSvf2
0wlBlwH37UocuOEu0XFL+EME9jri4iqjumARgoU1/5iYRf+8geWdiWt7hxqDrmXE
8uZY5wN20eJdZ6G6vMv89NU+NZ6nn4LKWtwMSkzegYakrMUOSDATw3PBG4Y039rN
04vZ2BfR1kHsFMn6wcIBpmpONSCM7erg5JDJWwL7U8p/+6+0C31QzdrOuc4Lbt/U
Ey9plaF/TmMeup5r06OrGBpJvxeDBgNJUwvFOUfjzPjybmrx7MsWJaut9f4isEwI
WS6fpEmiJmAwGjQMsyL+Uyl5l20t93WkYTtgUuvh0TT6QtjgbsCJ28nWPvkpeRJM
ZJfbbylCub6WdL07IoRX32ijl6EEU4gSimxQXE038MopCuuiOzYJOG1XbAoTozb/
MSFW6R32ET8vXHZF05NQFfvl8NE4Kk0WEmVlmtYgao1Aq2US8QR6UfuQKlxAEvN+
zQlW5pxT4Bs49Fj+llWebSQUimnx0rPAhCg10UxmCnltSUeaT27V+e2oi+d1tFiX
JN14vrZmQfIgN9QelQZiTZVa0tCAA2jnhI/5OFvBa+pP/DdXVs7YF/AusGVBhocB
FE5iYjlUiiG8TMAbYJarigAzikWyVULJvOnvZ4IOUWEJJOl9g58Na/yRXoE71q8l
P3quBHNTQMTagsn+MhIwLy8DbcOdKlbDVQFr6PwGdfshhLAwloC3CCjW1CVf345H
XJRtTrICFJCL3VjKKMTEEbORuHLXyDrCwLxZ4/xgcsbVNtw4V60zA61C9WfIXkT1
eqlCqnivZly5y9Ck0NO/UlHMGjRXUgfAZy3w/dJsRu8ZAAp/IGBU/VneThshdE9T
U8CykxiCXNFaSUM1wvJ6NGCaJO3TanUsrJPRqd0jxJNQ1x4YJXwh6zqsK4ZZX+sk
/21D4f3pZydUL8KTQDpq5ldgm9feTYzi9Noj4SWsIuZrapE1nq9ZshbMPIBZY7xo
8oB+YtwaXUaIzwdN+0F4tm8B7wvb+nBZ22iwYlPAurhd82CZN6cMQv1jPHfnD2ix
YX34STu+Av8+HzPfJTAPteLOsd+Cj2jt7UT9buCd2Pa+uB2C+Wpih9ryLKAzGnBd
8HP2QKv5C6tXKKrriy6je9gq3fdtbaBKBgjx0w4jKMtJj9jyPFEbENuFxforeg7I
OIuLc9pSahA09Pglv8Cllb28MWQzSvYRFzzc61QBfFOa+qKGCgwbNVFXWTPyzG7Q
mMX19IL9mpSVvzsD2KjOTasNJtv2CEpvrRPKc6yu8hNqbyvGIKVR89gCbiZW/DJa
wd38ud478JOZbjULwcEMIFNLT+ktKZ4rUfDVoyTu1w2WgcXesBc9OJe9b95FiQ6+
c5bWfO+/6T7vqtoRjndlCs7sjk4wTU3ZAnwp/NTIHGCkmHYeewAIW3dyVVb557NS
AQX3FpmL517A2mr3o7dB5Aj4v8fPYkMIh8MPHWOMvEPYv8/GCXRCmFhXxDMJCtCA
zOhWodyE2Va4JUWQUDVi/hFVOU2lD1NkHo41oHGXPMkGTmaE/L6+28pJSa7Dz7Gw
K9ghNkVqmwoqqSwEWM9wouEWOLmHQ4Q2juErhqngFyUO+C4Mo9dK6vT5VTGIXjXF
bbEveN1E2KMqzoRZIlqwhNkcmRZV8f52vviTToW8j09v7SKfLVqjSfmx3RgXBehx
0/GCqnV1W82PXF9dL1w7ZG0m7UrSMnDfc2wDQDrvo5gnTF4UpuixpTPq5PqYSpkL
FelYKR2K2YK7tedqS6cX2Ngub51pYie2PlWHODcAXVGLzoy8/d6XnYD2jZZZVGVc
9YvKDgYJDOocL7/cNHaa1dsamZL0TnexfX34DWl9lVb4B/yn8Ek3ecZcwsuvklMy
tyFM7pJFXLmMoKQTfMAzHotaf6iUTDNFVr4p4sirEEB17BeBjohkUg/75Rsu9ITI
C2V5wl+xsZRBIDGqi1Igs/p9OyN0vJ9Nf9G8TCutnvx2d6iff1X3n4XJxLY8GLuu
OVqxGqgWJWc50BGCQHlkKwka9+rq5pth/5usTAjSoqxNpqPxV4f4or1/Jcg7vSA1
yKAaPLDm4yjPz/7NKNbhGB89UOEsFOWIz7hWkAdukcCeKyJHi14HdZKRbOo4EBYH
QLKj2Q1W8OU6EuoXNQp0BzlEPAARRdIqWU4ZSm6FSV6kHsZBGQun/cK76YpFx7xo
IbF9fNhkiVv8GYYKgOSIUKM+oxV21jP9BK/JwVxI5b2W9eMSlJoy0A3vel/6UhhS
HJ48neQtruiAZHr40iXdM1V17maQ1zQ6RZ/dosxPcsi4dS8y5k4iiqIrW08vCVOA
V/iNYDeneguQb4pHvmNwH1nBrOUx0m5uKpBW1uTeNQbqjar37c+tFkIliumTQU7D
t3TFwbHlG9zQ2eSI8flQ00lUN838pbFX86IsUVjBV0ev0GnKJhDTMwP4ILN6tE/Y
irJoiUPIcrDjXUPUXjKAtE7tY80YfXFhd11RfNUTAVNTeuPtzF4AeBOPK6oiUNxR
s8Tfa5zXWASX99hKcwgo9/4dyzgM2k7OOIEcFWRkm5bfRk/KZmoOBxM527DTh/lL
5USxPMbte2O82G3tHmwC0yUyWEDUVAmDUvKavpjAK7a8ckJW3XvBZ21qYLYucywX
Fr/raL1+pmX7ChgBk+AHTOpGKkMtVAaIN7GuAq73nspfsu+d/b8Vh+IGZA4pAY5K
ddS2F2ZW+uk/WfaCAfTMEJFml1XHQ8I0Ihxe4sMg07bSjijBmqjw2r2Tm6kO7fxD
QtO+MU7y6/RmqwyyPrsJIZ0p3aq6PPl0mswKrBQWt6LTuT4woZGy31VLbf+vNJrY
0AYZ+oWM8HBKyyDMKOkGau9FEG7zd+Vpu1ralraN0IMDLZhc8S4yH0PwlfVKSHNc
mJQCL0bhX8wvivCL1RqQg2g1vCuMj3zE9YPhDvoMTvdmAMBHSXZyCWo5wsoqXH/l
LJQ8C2G9ko5iOZ3lvot/886XYeNSMScyqN/GF/MiLM2v4DLVFe3O23I6t/GOcz5E
8uK4MQL5P5ycowWVdVGMqRGijTXY1QvYMROFywUEGiCPV+DwdANlqTHzpBD+q7+v
5vKehm8GBbqD2Kiyf+WjgJg/1p5cy13I2GCDW4EtDuJshLhJBnPhVLWeFDNd0iPh
oxuvTuJwiCTBrkp2yYnTA5bWQ+EEg+CLdPBjx7nGud9gZz8At2b1+Qvc6GQ3pYA6
0XRCxrIeFK1G33oFu68iuBrF63amVpSTWrxLW6TZuydN+5FBJohefMXIWlIMUngD
OnpBlh9/HTvblUo09/ixl/NXjY3r1VqZ+XlaM9KMwgjf6HnuNyxIAeFJRDVBsTIK
5vQ+/dHMVr40KMEfUMFEGF9SSo6GGAp9YpuSQH+ijZ7VNDGkGAkVgc9gs5Y9Ggq+
cHyCe/LOUEmsLng0Qmi1NPm4eYk6TxcHMCGrcPPKDJgbBGd4uYLvoQB67jlewel1
V3ykw1olgQmmEcL69bX/Z7vR0/7WpWIaCDUjtVlFjxfp6VWkYjie06L4XWlrYWXa
j5sVa0lLAnwxOjeDt3RI+S3auLdHMTA3pt0p6+nSEriWFa9ESjIP/QZjykbjjtGc
VL8Btn0uCHam3evAoAM0JwwMMU5+ry2e6dASVz5h6Zoozh/DmGuSx751ewyHwfcM
lNDWIKjak6pjpjTT9E6t2/03Jveg+OybN3TRkCocIIHyNbOthFSs6vYBjn4l5TXJ
3fVcVRzFYINXtHtikCyTjaj8OLMwIsrRQF1ycN4BKbbs9fmBi+v6MZr4ODdZbtAR
/V/t570kZDaNfLOjSUfpByDaqxML2oZsoxckP/23AQ3UWgRx/7bkvUWjdYhYFrPE
Vrxr1YQR2NKAjRMQpArCNfg7TqkSwHQByjtEmu8SWgd2fMhKYBhn9M7P+/h8/THq
tkRM7z9izaSGK1nqfHlFBfZwvXlgNIGr1xoHQ4gwQr5f+88zCEwvAP9thbxPBMJQ
boL+Eio+prmivi5x5obWoplQOaY8FRH5WU+vqsAzmXk7ImbpN12wzshalaKZOTWg
XbrfWC5d9RQJY4PLDipMKAC96mSzvJmLNN8mpgaUUQhOlbQQDozE/KcptfvQVPSs
fSexLZyOeEGHPo8mBuBXtBybBbssJUnti+roaSPjvt4JXB8QPEinmsLtPOCAATHQ
AO5R6W4YO0uGFD+xNDIcnOq+DQrs7pDRo4WP/wPYH2UaCm7PbaH5l+fn3XYlJYaK
pnOZffg2QtCVUgSyIh8y5rMNXgrbOYd9WrrDWw0TkK8QStcQUf3ficrzqHG6lxEx
ExDSwBK99/r5GRn56oNDxbdKxCjeUmggQIC8WBqpRsLgmNNXQ+KKk8te4XwwdZeV
h0xqLWGWpSdGfKd+c22of3KhEtJwbX7btril9iLmpmm8rhb2At1nfz10VUIuUrL5
9EilhmAuejIhNVKsSt1P3kwrxOuCvwnJC7IuWTVOXUY/z09yb2Q0Op95+nsWiaAC
KM+T3POGN0tHilW8J6u/fS8J7+dUFklFDZInAyjNwtxgjK1k/V8LdHkNZT9zLsiu
yLa9HMp6iVjVjiPpaEtLhH09RZqpKlrhuuHfHKOzLRg1Z0arNxVaQxD6gE2MYjBY
Dv1+aVySPZtpLV1ytUEgkXj9kd0c1W9tWIzSBKAC4AGfhCI1HlW7n0QkQMw3k2k7
HP8lEUApiyGIrX9MuWW1pWDN97y6sAt7NTyiBrz6ZCukRR1Dwk9zBhjUCgA7FXBT
L36HpccVVg797wMD8Q3RpftcLf7Gi/Tn/b6ytV9DScjBoqZyZAIbCNAJLL22sv7x
mlvnYRFCE+ryGPtn2p3ABUV0HkrYJebUBALnS+qBl2eaUMmuKtpXTsMbmbsdPX4e
KULVbCjO46kZkBEk9FIgChnt4jbLHZc8EUe6EphOIGqL/o3N4V+KtUG00UDHFmSC
/QvxGEEu1HGLf017zrwkq+QkFZk+4a5EA9+DOWq6+NH0km30dwWbTu6bPEN2pyIl
puSH1XCdgC0i31JTcqsmaUc05nJTBdznPmaiAJzKA1IZ9GD6z9wBrJ8NESuL3wJC
GVdoF3/Wtysqx55TjXY6a8IeDwbtimoa1DVQ3I7uzR8HzT/0hwAk1blAJS3GqR5s
TeMS1Z2FjJf7fPD1+4MGjnJFGrPMrHcVOG23jUHR7Yfy1XgPPmEVhNYdJWhum1k+
tL5lSHXzGRi/i3eN8jNZG+oT2nyxZRzajYsmfeAhaT8TurcVq0mB90smJ5yKhGyM
nTR6CW/YR1nLaxXkmmpvKgraPo3BGWt/LbJJHIdoqQSW7HKugEZlqwzTax+nxnRl
b4OWU7fN2tP2X2HSv707N4Q5k8hYTrm2KOuX9vzn6cMseIlJaE6J01xdwUrQcY0r
dInwXIvmQSnkZOaKO6V1Fmh+h/aKHGz+TLT1EQoR7W6gPh/PaHjHy0vX4878U7EH
mtpDqbbCKU7OJN8ibk1rabH8c9R4W/qlewiP5RxpApNVFi0i6oXk1vwQtkV7UcIk
ReC0AcyRTiVsoXe58TFTwtjEm9H5KCqE7no4RrqRV5oHCgfe06ANL2hzo5JDSgaF
H0SVw+zZm5Ql1nandqVYkbvrToHhHjM+Zs4mjfqb0O3ocfKRascVq05UP/gd93Py
Yrs4svaVuY5FbOjPxAhsaWYANmzsBfmGwzC+Md7Rzgj3u2FiWnaAeLqhM00NT5Wn
k/v/o944Wpjl6TTem1+pO4rgMU80PJx3eTYTA5kLKlOWTZ+CjMOd3flDMMHpMV6v
bE/gbNWo4lR1bgN+lHiyhoSaG9n5bQsHXBvMMeOuaYGGpMYiLvMCkjYRdo9xbhWi
esu//Cm9Ng7lIsvM3Dg7O9517Zg21h3GGXKffJ21YFdkSLZMdpJnn08lPrhAp5fg
FeYKRBAro3flORW1EZCNodIHLbYXdTw/Uwerb0J9uWvfr/VlvmqLrVyLmO8y8K9P
l1DR3GQh1tk0sqGyyDEkAxPMBOPPISkvDCCwvk2UhFFvQMwlWJux6rjLBmQZI2z/
bmEs/Qcvzs1un1UOy0Oq98jYIV7T2A+cvsy8Q49nXOfCdP3Cagiw55br1+YOPt2q
RzGnImZYUwA5b1Y0gYQYy5dke8Ma1vDpr/qJ7au5baLBb1a2H7hbkhw7cpUl0t5h
qVfZCbv/Jfib5CtAG/ubEeEuuK8Ho5xG+9JMgR18RiQStI4XODTBtNI99+GiVv86
7f/BBkuh7yOMXfk4mlCkNBs9x09y84HnDJnJvWO8RWyDkpZrH8K6cLq/OVMU/b5q
ReG0F5+gDV4w8bqAACUwmq4SmYiFzeKD1w+KB6caesoaLiNDE/5PGA3Azhxc/JlV
wDQ6x/aaXxM0P33MgNC9DStlKf8UQeqz2X29G2okIW0pTFqR/7D1uatdWJz7aZB3
ZOw2FVX+PgMEPQofGGYbE2JWrcY5ihB4GAE9zDHRVFa8oHS9+SFRHzcXkX6IABJM
misFhswag9Wn+68c0ng5RT3S4rpexUw6Nt6Y19VlziYluNABgVf+Kba4lse2zr1N
9rWkgq4gsM43GCYWx63ln7/wUv4wOzpzO3QcXWXpoT5lgREDyIA+9dTfbMQTYa86
gkLI4iV6TdFiq1lzb02Wz+gmYNF+HpXY/ZXbwuaytaPcjXY7VvbQN4/RiP3WRntf
XAWn5SVea7/4s4XWLuJOhnOibGdw+7KNtmZ4N3ronCTWK5zPHvq2y+8yimNHQNf/
54nJKcsuHDiJrURSITQvSVBOeOiy8rWMMZzOOo4b0v+u3Esiz6i7ci42fqiP0yH9
v/03gwRbV1osfk0khokPWP+Elr6DYw6F1yGqjSoS4nOF6jXTHXaEcbbDKCi5mTM5
qX2treFHv+LNHWAUXyFimtwzaGF5MDnBMcaRlyz9AocEUZM9kS3DnjfD3el1cRU9
0MkPY8YfpMf7QHCl8OJhZ0ZSZwlxcm2SDh2tV+57k2DL0e+Uiv6w8xEmnAp139dI
VFEJySNn2N5gn0QASxz+mlQ2JNjSsOuqQ+J+TC+C7nUIay/t4Yda5tUNeMmDWDnf
oL3AANfbK3YAnnxUbeaj8jzLUjwgT6eOgPvT5bwdKgx9+ONLP40FFofoJl2rDDYS
veKrjDARPe8NAvuEpeE52kIZwSo6/cx/Oz3oA0SiS/82GU0K4bTjxK49bZ8cFLQf
fC3a5/V8uh9qUKahOtGYcVWIUCS3yWiPo9M47YOxjOV4BMKNQh+8uW+9MAQAWuvp
nCrSwEnmvwR6HjWxYWcRhkTpjkNOVYTGfaB+UUjMUCx1Tj7iOixmiz09yWIsbS3q
9RXhgU9H3Zutumib100+DHxela41o/ySgkBbf21hFEJWYz64MUxOtJP+cc/GqPRv
2LLRbR1i8ibv9FUG5mST3PCJBZUZWnvTpzqEjuVg2M7c4iGQU7Dx+kURMW6OINC+
1lr33458N+ZfYf0Wj7txe4J87bGPzvW44R/c3Nd/qX3jWlzbnZTGQaCWRJuJCwx9
FahqXf7aL/5nlT9MKbiNBYSboOrq7Mp/3Z/whIr8Xgz7uLt6j7NMyfSA/I8OlLSK
H6c9kbmCStXhPUPMbrS9JCuG3Q/L8g1wadUaXpNK4XpF3nzk43GESRACetIpt7FT
7iUTf//NJJDZqg4K6FXdiEo17oxhwrmV2lfYUv5rqJFWPK8DUz+Pf6kzgdAZ/vlR
GNbjNmyYxjwedMBVtZ5WYP904KwZ4xq8M+Cthm5g+nLoDmHXr56v2Uu7Ns2Wmj4S
HD1UAB8qG2uoTMO/ZP46cU+ziGSUolq9fMrg+fwKIE0/EopHXYoNzDM7nSMYv1BG
KL74duCCrrShmd5k2WCLQang0oc4/5oQ/APj/AfPThgZgkGzdL+ASGyCDfq3CL+O
lQPOv08JSVJFerh0wNq4b9OEU4lnzC/hxFCFUWNGrTulFZGL/3kabPuJ0F7Wg2JX
4z+jnOp5dAn8YV5QQG0yP1EofJgZQ0UxQW4539eh/Tg8nDIuhZiVufGqvqtsE7Tt
qSUHEJ1T64TA47gSWQZBWtUTF8V7FDEd8GyF2HX9BRAHXP/GA1hdRJjR4zoBCee8
KEI2HELBb5Bztz/DF4VIrmZaVtxADuKI+s7GMU7VBYx16ZHdwZpc2k06zNQcAtKY
cg/wwQ2bvzXQ1zWVWxiAX6h7a2ZhWuqTY7AIPUsKhMp+Jdun4jig23FQJo7CKj8V
Kp0+3keOdGaNMqBEZx7gEJmO3KLJAxTx2s1eXE7YxrZoiOIqxvlJxdgrwORR9YUa
iz8g8rF1pxgLW+H6TNeTBIoz0s6/zB9/Xs+LvOn1VjSE7gXY9XdKQuZqTugrtDEM
dHWOghsk11YlVWnkb9jMixugLCoy+j2ZqyrcB4DcKNc7bjitBlOEeRdjP1uu6S6B
XZsAVOOMg+vbsqUKu9I+hJ7yJXcLMEejCzD/K9hJwn1S97Dk/sg4EyF102z4rgM/
ZtDmwfsh5bAQsQbQ7ZVjrFRD9+0lti39E7Wl7zmp0DZutPfrcynQ9fr/7V//WPhD
FBUSXkIM/MgeS72Dljj8SowNRyC951HO7XTUlGG/FG95BmdXTP0jQy1Q3yBNWyZQ
TggKOuiPBOiS0c4/WscVQcVzM+u4Ap3rWZJdK2404qJIrLxF3wiIZma8tt3GqRQs
m5+REFhd9FQDdimcHYyHBpSjKXgeM0Zy7OIR4+VdwbZusAQ7kFslrSG7n+ekUq+L
V+eGgX+9wnkMPfaSnVLjKMkAM3JnMR/ggJmm1lEwjzN8nD0zzLcpDAULWGCEjTg6
9sloig8/zR9dp08vvvixdk5J/WzYRfQZBOy/ukXrSmpRPhiUGzkSPE46+E574tIk
KaGaNF4RZFTgSXWiu4EzDNaHW3VjtCOtBFf+KHsKFoaWslRsqsbXl32UhC5UncFt
kG6a4PHiOf6ib+bS8FfafVcthM3zMBjKZBlXyqfw4QVLUTjj7JVwMFCXWa54eN4z
6nyqB5yub5Vi6wWuFDGWO0czsz3ZGQ2rdaL5mSEKgsDnWtbprrAqbetbA19y9wxW
9AWv70Oc+qGYX2/cBccq/JRoZeT8Wwz4Nwa5lpbJfjuW/UDL7LAw5sgvgVUNY9Q7
boJzlIRG8wu7G3PCs+8Mzlq/tGtiXGm13y87F3GoZ6rEVTXN0ks3BwDabbA+DuNh
NRkg6b2vwbuYcG8uv6Y7VgGnUSPiVk8+aw+rVWO4PxaQhI4s9UiDaNWuk6D3vTMN
wWKWyaiqEiYuds2xDFsuatEcDOhViSrpLSEevTWrfNxeKRkny3IHfAXbtvlLCfi+
bTw5q2AmRIziAmmCdVcg2TFuq9EHUBY56fScp89Md7A0PHy5LWdEGU4kXhImSET2
zptes1qJEWOCBuuKTFpju6HksCY5CLmvjeX8Y4zrQs19Ae4C6hmwNwMY0L1N1L8p
gnmnvkWbTod5DNlAsEQXI98ZlD0LPH0EWQ1cNda6yzsUgAzyBS3OAd8wls8yu+Iw
nwD5vivghWvHZdGN9W2ky0gMxKCeEUnQTkWYViZj0nxeW40Fls5V5/utT7aKFz+d
qvaZnBTIa2tPyKFXbifxEnnb4qvz0D83jPlYkfbd0OC8PSXoljAVOf6ArDG2CviN
Uz4VBASfDYEiCnjJfubkzm3xKHMr3S85PLAtfiVUh3PZ/A54Q9/c/EGG9JIFq/3S
PS/ygAzyuxLXXk2hf8mym30aChZFd6FT5m8ennJg4kS45FE2VSJgotllkUu6oNCA
jlKxh+HZbRzCE9JSHv/liGEbYCeREkB3gd0ahtSX8HU9VY/qpdt133iSus4n98NG
6oinmI5p8B8ZYdMJgAyB/pAlTfAM4zuL0VrInVKTRtnQtBtgjtn1iYto9M7T2EqM
BRiSph0TSyxsMIPraygUWlGLI0JDu1cHSLabWLVnROwkenWjM6/L7UofKJwC4EpL
KPo+A0yWBfgiIv3uuZzz5c6Tql2/DovLFXMJi/JiVdOlcQ8hC7TcZduLk/BUG+tJ
b4K3CuqisaU7pnRXpH5A58QImm9rpp2kMLENdFamgGYXza8yfkulBurO5zwY0XjF
gTLLTd16RsoSvAUVvr+JbEfdirzihS4yTurrHkcHcSI1MhmNgYkja3UrDN6E16QL
JMElihUfPs3+y/jJLer8LqhZlGjqiMrELnbuzv4n5zWFJubjZxRaKRjvf7DUVk7w
Kch5UOdbovbOcl9l7/RUcdsqV0fw4rCF1mbv6ZwtPgypdAJ0L5OrfhFEHjP5g6wE
vpv/adCAXLICi2astLNoyk+cP1Wfx63H3CC7SMoL8X4864oCEWOlXk9g4mzlBpcm
qbpRN1ISCwvIcsLl0UPOTUwNgnqwvVOPxBxQlw9Rz4cGWvegMKCtI0NKzvEtf5dX
nQe5He4xuvrNznMOm3xxJy8WAngZONobnPulyVj3DWtTPWAsBjxDTbQEvI2/awyN
XG0KRcJbjXzjkXa5ICjHh6ZlfS71rI1q6ApcmuAVq/6g4c+VZmHQX4u1eRLX5o1P
Z/qlcNIx6Oa/VnPkM14iY0gAYAGKf+/Nh4289vYJpALR+tYib0Cj1kypaGhacC9Q
Y3clMzyaTjXUUykx8U04gPxDU7NbiROioFW35Fjij1lP0pupSWIjvmX6KYW+4n/O
ZVk64L22dNZQjDgMfwD2/ZLg5vXnybgOpOIvkFvXJh/xlM63EpeHVU78KOc2P6WY
JLM9l/UNuIzmJaScPBdIWVQLIoUqKILebcX3QxXnq1117FO24ezBlU9KD98onAka
oPJ7iEAXn6pypQl1u7UQ7OnI7/Z2CJ+56jQWXnQ/CTyFLkHvSZMT1MsyVfr6cPAD
w42qWJWL0/I9GrYZfxHjiTWJrfXeURD8hmJFgqYbrhpKmAilzLS/UoAMHl2gJJMK
g4WaLwNLq/yAy9hecwUWbvUvQdZTxZLC+mdxolU98+4NkEhNtblnH33e718f1vfF
ctUEgsn9ty4AwSwDQ99cAXy3sd8dkd3xHV9k8Y4cGdORzvjNRy0ZFLpF1zfbMMZ1
YPXM/OCNTHVi+NcMSxUgG3MuoZVYhi6ogIwhakg+//I/BqXC2ujWKAby8h4wX4Kd
Gie7ZEoHKzFnMNda+z1ok7rWAepGXVzsZg+48ibFl9E30Ndo4PhZesW3a8JM+lvY
9UKSln+U5rEC23cY78O7UqHyGZZw4YYTKjESiSS4ZsNDPD8+TydGyfJUTD/0/Dzc
EYkJ9dNwR1YtYyvT3riWOMM4XpWYNHmRyvtOh//2gyKKrLhTxBXx47OPQuabZKh2
vnGfSVqgk5pfA+XTOMjXoe2NlcRvVP3taJozslWnDKWztrQyILMpu2ikKY9m0WtW
NPWB13yajuIR2A24SmMtSNxkJjyjfGHkOAoblCDpJrQZqltUDG3L19RjUUtt7dqq
oH1NtQNgylP9TyUf8itVsRKGTJqPS3FaKQEilrLkM//BHAM6caTjGX1GUS7rLb8Q
W+Sy7z0Q8aytIbEaMz6cTwWDLW7oewZV4zLStvCOfFK6Ypzfs1Ma5jduaFUe9Jvn
WRioa7NexKZAZbf2aidFnNYkHaijSfS+u5iiPk0MgPMCVxzg3ROnes2+2jjUe/d/
vv2TlOdLOTMWCoQUr8ksBnogNrlcGtWTkFE+oGKypcf11RsED+phRmSFEFdn5Bc7
yUjItEFBc2WK8vIUYtG1nyZvoFbecDK4aE0nYqBpEX3QjXJBboZzjUkPOhkPJUzV
8Diehgp2h5zQAjN/dysAXbYnzVhm5E0PazUegJz4tm39ZfScjElvKnqwYXl6sCkP
dW4N28/awq8CWtZ+KXSMhxRckSEfFBlfazDZgTdtfg/4f02T97ke0rb37ndLCPIY
e9EmxlnGPrgyXqpBMlBCWb327sC85cLY0b7rzquXqhNtAbGaybfeC20dbNAHXm26
seS2Q584UwAluBVGENRzDp20iydELqcZIibTCFVWMaR75adScRWjQJkW7HiUt1nS
zDMQ0HrxirGoqOf8mL77kFk1rZBOmjOPX3yGuvX9CO56IXMXyKM44xARoXUx5YEz
fFFRZw7s023y24+TwIYgWuIa71p+5D0xxeuSlsuoTKKh15UBplRjY0CalLVCd+jf
nsfIedTA4yYRiW6FJRMKU2DB7LPlUlrb/zo5aV6AEnmswHr31p5kvFlPhrnUVeX/
pMKhAHrtPK4LxwJqTkCLwwms3Ls+/3MisWJpE68a6uNnz8VqncY0o08TFEmXE7cc
b1NQzApDmaoYxa63shWxq9aOKEq5XDtuT1vY95EAHsWuy8duar7+Ot/Vcp76Cjk+
zNVc2VgOHHa0OezkQIMQuh150usNoTSsSeLegntgTfvazeHzUoIBRwhlZK6mEwDM
2W6yknHy/z2SrezmJJIa1uBY+iZhu1/IFsPXTvUCV1Mfdo9f10vJ78Ou/qHvt9M8
I3lj3OPaAfa3tu+Ab1+1NtGeY55+Tsww4iudOH0Wqe1e3qw9o3ay2ZUU2HeQPpLh
DNvYBKu271/eEZw7ubnEwfDZ0BY8q4Ogtw4z1PbVVm1Cn8geTPau55QzZ+N/oRfh
LvKdRdcLj90IDr4COCawONqWRpof3Y5+Jio0wiLhrfnoKOZ4YjC2mIKc7PSHuK/A
zgJT/Hg2hlGqGAXSOLhq27Gwl8qRTsGXkvOROIDB3c5tvfAhYbNZWUoYimOdE3Od
dA1Xk4nz/VpJG+4Bn62G1NHosvSrg/w8o4K+DCB6zS3z3Rx4EOaI/S/5zKTSqjCA
jy6u7DRJxEreoi81tgOHz7cbY9zRT15xj/3xp/opkc3wo469FEsZ1aMJBeVtGk+x
lmqNxP9zOX9QRkWwZMap08vEB1tFs4VqEouJJq3mU9FDwFwBV+hvCvcazM5P1Pja
1v1ISWFMsfggH4i/XRj0riccUyftyBDidzryBisqhm7cMc5/nW1m7ikbKfc75fQk
AhA/otvavpDNevXMpyflJ+Awb/Z/aNKH95BrzgemN1EcZNLpOPM1/bkgTqidPnVt
yC6vwijrT6EC3/CxqKUqTHrKZxbZmqHY2FVoC8k0jURzhM4py/Vl2Y7Y9NWuN1gu
GDqV4nOobiO3Q4H78XpkhwDPn9Ze7hg/py3QT+u9mPIaSI76MbSH3Yi5LYpZRRe4
JH2j/LuVuQ26eTEgFao+E+hQYJUc6kmhUIFhxXdiYW88clDJ/QyaA/zuMA/vL28v
Jp55Y3zfUXrZ6zcqOW+dmANoJl9qAiKJcrzyQZfGyxGhq7mpcGu4YKlkDMaT+vVG
UrtQ3srARCPl/Xbn0Os8nDjhSg5PeioQrXI3qIOA7mQ6Gn34MNFaa/uBxfkzzGj2
h7Sv12xMZ/uX0mfB5PBP98OW33MBuxR/dvg2TLYkZu7KVWPZl3tq5tXXVfup9v6J
LYPL+HK8A+g2cC6EWTLXNZnJhG2/PFkAkt1JwDbQjAd/rEzHCSbRkX6Xg4mpYsRd
UjF+FbqJvbvupFkQPPu+zhpVgrlNGr31PccNJ45iOWptmextRyFvDNlpI2N8Dep3
mQcXVBukx5daryKg2661MvZCRAoBCXskejGvPj+ZMjGJ7wnr6G6uzBFSX7CRJKv2
SuuL/3QmIIRaakM+Y672R6FEOYh2YV7mBhPUjc/2vZ19jQLo9HSlYhw8CA/b0E+L
9C8hCzkSBs3YRXLKc2jarT37Un8akPyBOToqp8ZSDWfOtLhJ/R4Wh66OhdPwN696
aZaojOs4oaIK3ZpzBLJMY9sEa60+HzmLHSlOZ/KVdA9FVLiYEQ055h9mz87KI09O
TuT7xIkch1CWRrLlFs0vUnJBEHyZLX0gw5uaVSGXDc9z+gQYCmV8c3G535WWr7ix
VSvxVa7SS9F6obWzFS0J3Er5uhEPVTGldytG6Ml/pe0CZ03R950pE7YWFj5L8pdt
XHcGYDz8j8WFjJZgP4tc7tOw5EnkMkm1tLPBGbNrB9VvsF1nlw+QjVbQHcLl96dW
L0fSyM8y5yxrMBObVTw+M/nvGUxQ1ZnHX5BGThhwLxwMVLUeo4u0+Zx9igBpyWuC
nhxtExPm+y/b8SDYgx+ou7YflWgNuQixce26PnXQH9SisBcPCDw/m1Lp3YJz1a15
pS8NEczO6r/Y0MTO9VM3FNfmbtyPzmE7+kUDSF7pMEgzLbG5ZZdopMV0uZmH14t0
xg1jZMiPT2c3mJEYC7/vlwpiSD0WAD4VB++Gq8HvBUi5lZdg4JiEdCS66VEaspzI
G4h1DjqCOOJLKRQxarLj7ZA4/6RxmnOkYnlcYAZahLZ4qhHD2PCtCmY/RKcT5GU2
uswnR911tEuO3OEHUzWQEbcF9yL0YADdLx6ESid/wq2Se6A9Ow/svbCkCmT5Zq3i
rJi2lShSDtPDfmqDwJoV99j0icQwxcjabhwLqDllVSY0YD7uiWVuq2e7EsrL7oMO
1PDGB0mJH4LdhaM/BCndgLBc6hhG1mHQzaHflIyqEiwGLO/FJd64apYhmuzjn0y0
e2QxMMCaf6fGjO/eeq0ZR/S/ufEkCJQhOLM0F7kyJUoF/gwtqMsNzh556r93CKR4
IITxGI2qVwqmbnF8EO2ecbuxT8EPlSY2Z5+mlKhfsWwP0xursBv6ZV7oP5g7V/Uo
GytuvltcdluHiW3dHPFgxpRmE5UFEryrCgWdg5AwvHCscgUfXMMRQKbwXgwjs/xc
M4J+8AiFiuQCyBbBe9yHK3QMRDk563LSqejXikuab4gnLpWnOL0DUH72QQPYFRew
s8FZYOvKIQikuJqzg4sp1tKLc4O0GUlcMkLilg+8Q4var547X3RVdZReZEU/WWWm
Lu4Wv4esA4yTNe+4WF6DfqCUSsFjlJpoVaLgNeuueYcIbKdczvb9mR8DEpVdOSGJ
9Gstb7FWVdRayUj4djpR4epQ2sGt1AkuQAu7I8gy939Od1CCg8z0WehWo58rLLIP
WMg/ZZcIDVnBwtOm9oRHzigQzJhg978tDUiOdM63PAkj7cdwYHbQAnUXnAdsG9+s
JHaAL0+Ag1vDsjBdZXApI63SAQ4quwFR3cg++nQ8+ARiNqOYN8uMEpY7ioCc2eVd
jgf2Qp1LfH+FNm7Hncq0uhCPFo9f+nV6NDO/0mfHzEmXlCY0kh8bhbwaODtO0NZq
Qzaq1rEwX5VJmWCrh6KmDSXRT2D0qAF5ZFyTBRep9BMa36zmPVXjgNNzTqRDLX8B
HdrMZlhtL3T2YgN4DCLVGE3hMVy9jBluKZBSqxb+o7V8+XKp+HGMDz0SCMX4HzAx
s2755VJo1QbRX0HpdfFztmLznPkSbRoqNVHb5HWy3pEcS+8di3Fk7z6KGTS1C0qt
qN+07ckBhkpCHOr4PFPjnz16YWLnrzSOj/gFmu+mCbodVUHTOlbkLHorFUV+wO9Z
Bcq4WEoHqXEcVuYNGF9oHDaReH6nmmRff2UjquL9zxlAHU4aM5MfOp5zJNsF/a/J
l9giXRHMYyXgTsyPeHCTRY69jFr9JyaiqlRTfMM3aOViU52fEl7NaIzHhK4PQOR5
c9ArN7NpgapW9wkR8kubAJSXkJ8wugLF/wq+S7zSRpN+ZCbFVdw9/WeGJJJvWBw9
QYYA1N+ovBYs3J4ebprhI+x5y9zs2qozuc51KJxVE7m7tIqwiZfFy8gWhyYqLipc
v0IDU29oOPlf4CG5k5GI3S5RUHYCjXsWDSm4OP0nGnX/7eeHoIZnR2YZFMuxa96c
7xxgvk9bW4OzBU/QSQHpCXUpj8Xt50Mfkwb2F41nMVUBHP3+IyCm7iKuTKfn5vgm
wnrxTU4q6Af6/06dTekJ/LolQrTVQ6obyn0DVhIbeiXvy2FMPJn1yqRnWlK/zC2c
qu+3TWmRSvTl5bK9yfj290WZ9301xtq8s5HyHijFU/fnXv1EXWXhAmeT6j/fqrTU
OsWMTlt/HJfRdqkQILF6TE7XFRYubvVta8iQAR2sFmj50U4yxD4xkI38oAJfRlRv
vXgRUn85qETn46FzMYLpV7qxd9pvMoZl5Q2bBXbdT8arDw6hXIiKaSowibfceslB
kcoJSvna9u5BmUfAC3+/phsWaW20EKRWkJdKNXUMZY4tADD0PLVY+ApdeFcxNLZx
oDNd1hugRGiaseTWKuLIfg8F8BNHYy6J34IgVi74T12zIkISGHzlVsTksVSpOpJj
M4WjzucIWm2qXcBfFXrndb1soMiwpZ+BXCcYz3Z1yplAVvpxntRZTtGotmDVBtbz
P5NmeCxhjhwpJZBbknJBOeLeG7t0W0XfEM0yZ/+PU078694liAX/i7/kH9f24hRa
sgauDDdnGou5uXfB6G2EBJkMu9dSMoh/npXNC3ZLSmDKn+wHMr/pRVYFbh02tLwI
qkONdpCweWGsYqZfPKInugzH8CHZfvwi1J6yUvmfg4bzn7uP65ksFOS7H2u7YRA6
nmFKvWmx7ugnJXXXajnaw0bAV8+U7EcOT2N4KmvrZEJWEKrI94g3Ebcej7o1Elu1
CJhwdlo7hqvC34uZjRX0KWTWpQ2JtUOUDhbIhxaZN1KcFb7ijaDuBtL+ArOV2X6n
Vu6E74PfX2/rEBG63VmqpBPbtldfqCCmc477bYpvW1mGEOIZHDYfkYc8j+6P3O7Y
m2GzHu2cjvVwi3Iwy5hb1Q+IgZd3DQZYKToNwETRaEnwmiG/YmK4Db7T9R8Du1/W
en8rTOTdvc28fQGjei0ortTAobmkotdNOnYONGhl/HXq48PQEbGvTOCO2Y8iDWdJ
FrS5HIIPqYFdzFgdrskm3kRoV8K+YcUiBSB1dZNYFPXGXPv8gg2muoaIDI3rvroC
H1s5YRRrMxFUz5Uol2ztfk4wgf7YsrIiXkWmjWgPtlZtqzRZfNZR2tZZoGVaV4YV
1dm/Q/hsUKZeiQ1KLPwaJaVqpIBeVTKohDpS9lk6I8LrCD3ZrnaQlHvqapS978d3
JGTa5L3RhvUCUcDGQs9RBLpUadb96vZzj8CFw0gR7vJUCWX1MaOksjEE8TpnTvIp
JnTWc0LuVLYU/D+JhpsSasjiQjbou1+ypSD6WUsWjS4JPKE3l92ZGTzV3YlVqJKn
qSByN3eZKrjsl4Ysh5Sqe5CmoBeKihSagG2T7EtlDj9tSc3k1rhH13UaEtD+w20D
Ey+DkVXovzNvzvkhBrL6Vleh5soRqCXOMW8yUt7clocWQBFlYHOgEHKTVlyNG+7Z
k8T9AKoqX+wC6DHfVAO/UdaIfzeOeP4YdhB8qH/MSTUlaL1AF5FHjvbuUX8TGaoi
a++AhKUqWWBUJs9eWo9e/gk+agcLxVotS5js21UaY0W/u+fya/mOHbkv4BE5udA7
jiiN7OOCm3jyqwthXNKxOuPQLKlLMnfjIbJ2jVhwzH3gjeVHRqFGva+zROQYOjCJ
YRz8I24yAQRVNf3DaUsvP3qQOrWgRYhpoWYEukRdRtJXyEYxG1EJ+cvqfy0d8ukV
ODZcFMFfug0iDl+9NZe7gWX5TnL7oEyt4N8vIFoN5DV7rYgfWNCmIQMaXXqI29wN
lGYU/wyw7TOWlRa3VQM2Y9SHztwcBfisLsIwR7nfndGg0MjZc9qdgpTFoQayzfCv
6JjEB5HixyqNXprh1qjJ1qA9ko6qiAZQK9v9P+No6/rTSNofmxjRuLvWRrB6sat7
ZRHSGtVSmR7UJcAnNY5OUfbJoxD0FUg7BUchfsyX7z+ong/6OHbla0Kpw5wY9VFH
oazwS325tJmUJw1T2Uht5kyuvB5owYF9L3hoBNaLiEkOMfnU4Hlr8aniLiyob8Ac
MSEgvYofu0xDhixZHEuE7ga5NA+J1IuQs/mKtuR9iHBlELflpw4QOeAmzFyQayLw
RfdJN0yC1K25NmFxPS+0Pk2PpclxSD9FxzLXR0m7gR8bkJq+x2OTAGA6el30MAjg
EMWBRMCt7Og3lZ4i5gG1nLmf3VVqLN7+e/psAQarZ6Ot+fDvXUL99grrqqhPrnQ/
pSDKcKWES7qEtQWxUbL+KZZHX4M7rJArECYQmDa7y3HVKtKqMyFiOXT3a6XwkuKM
XTg9cF6aC6n7+HbOrkG9pMv3HPSA8WvlDp8urGCqlO2WmIhZ1whe5ZmBT/EoOjrO
8aH/pSlj+PJtPuoRHBF1HGa160VDYXrYQlfsqSGKxr9h4uXaKQBie0Bpd/W6msaI
rwbprfjk/DKEqLFF3zj3yuDhAb04X8zW9YzW+T3aWhJF9cWpCsLgSOW2kRadJGOz
SdPexo+bUyvzEbyZb3JV9t2tOudjWTYXjonNKKpZ7uj7XaiCEulWdtTuXhjmzPF7
XW39D1On+FhvCMWm57MUR/PNRhl+m4LR7GGIBMY79InDWWfIHr9MSjq1PCQFTg2+
X3sHC/cCcz/gqzMpRBmBG+VdTwOmyVn4aEpD5Sgk20b8/U5bFMESogL2vZw8mYEd
GvtvGoroEVn9ASOnLCShnZKLiLKsH67U6S/s8g2P3T9+X+cfzGnhZTT3zU/AOEwz
BAEPLfy9szRWG2yT42FR+PV0RSmcl51sviMGElA8Rjlqxq3s7ndHTW+cbIlJLIOT
4CbE84fNYLJwxX9584fJ9OH7LYt+vN3AisTgnkdMLqwPvSNKLW/uHLeXeqdPrkY2
3G4WLlxXny3z8WdA7DU3rGTSIjvgHTQ0oJGI6FSqvXVBad0UsVn36o5vWFqoC7F8
vB1d6ReLOGhiZqWh/iWDOeCal9ST/99fQ6uEv/Qp+QKa93pYfxexcwjUJb6vbzZY
XI2mbYDUe/Fr7o+nuJp7EWo9/fAHdJQv8puZyaeLWgLXGQKpBmGom40xvYnlAH4l
ITUO8Wc6FFSyOUGlvqujS+UAO42kQaV5VLv1xEYqoqzLazCa3aZEl7WnDzyxFifT
KbuIFNwdrwgawuuZ0YJO1pxGgh0Y+mjow5atztTOen6flTowHfPLGA7Q4ZF0hAtB
74FV5P7t+HAfBjJfyE9Ymheo6Io0FbmaXvISBRNlOGr+IEuWhxhWJGQnfxVxVuDw
mI8jZzh3oDBqIFcblhLvssdPBqYWRsXGVaoxUQzvEAud7mkS+fjoDUVfieGm4oOI
57SgqirE/qJDFesgNSudrJjHe9iifF9i66226KNi/WIwiUZHeLjjjA3yt3YX6uj8
tBCdT1EmCWwX3Z336OGTyiZLCMXIEDnk6SKuk33U42eRYS+awgw+BoIEJbi7EN5c
GIaIyLGIklaKa1rVaRlfrvWAFLrxaCZL1dYNb6rdj6HqZczRGunGdf9BSy+nd8PW
8lRKeyWpiccjLLzOz4ATvkJbJh0TwudhDeM/Z4Jsa7b2fOLMY+Odq6Y/E8iDEZUa
JR+xcnWRQJWHyTP5stKIFMIg4gO0M7BYT4zmTxEP2/CSh18ljxXd4FfAeHvBQ/0y
BDS4owKfI0huAybBkYYzSrOg8Yuruyb7obiSRjEk3kP/20yJtv0mbwKJOPLyHfvX
T3dnFNjapQoTX/WCptQ/I4NRa3a4lJLL6hFtgB/5CCYqGoRb1yI16YAIvpLtpexY
9fWVj4be7ctXGibwAg0RHqngQV0BEFKhe+6S0x0hnWEc4oiV0UoRB2bVRSWQkX4f
T/Z6YEk0Fb2IgmfBOUNrVsOLN1o94d07WPbbSIWuPaG/qGuPKuYYpSx+m1vc2Eba
82e+EYI1pSBX5fQaDd0qqxvgtu8uGGgwUnte/mDSfwv2hCwt5opD9L4F8DKaWh+O
bR0OghqRsnXwzJMLYw2bzhT9hA/uPQZoOmaQMNVFuas2u57m+qSM5wt0gGCTwCxZ
fEJ2rJJNEIfrGSHhQ6seBHKbwP6EjEbXyqb5sZs1xAzbA/MVp03erbKVHahs+Zc3
R2q2heGwnje/30TwR6oUD8kN81S83qHvccNlQBx05/odQYCDBbyUOFxvgELxdN5/
SRajvAqt6wM3TbJQBu6vQIZFVY3CtSfcnlTdJaRND7u2QRxGE4X91TDL69REDxJE
OKFjroXLgD3G5sWwclr4CB+yQtTeB4A8cXVSWaezRc+Jgl3VxUnvo3gzLD568kth
8fwpfIXVlgexN5hDtUb+QZlmuKeBS92S7u8UfROApU48y4MhnGuFEkXEzlPJ5Z5p
6hEECFVrViYhzSLl+SWkJuCqsIUQhrtr3SxbzBOi0do5K6b/rRMRKxfulqvllWb2
JzX8TSDPqSfxSshjYUC4sMKucHnIbrZS5fUO6grb7hu1UVp6gGmjmuNfyihosCGn
f0O9kLvL05S2r6wd+8/78+PrYcdVy9QtSLSC7Z/CULgi9evt8aPNSjWNGzjo6ngU
nsPlvIEUvhWtlcj9Otz4eTB8zaWLIqEEfz6ATfoQnG6Vzt9yJJ5TINSVXFJFGL8F
2c3FBun7ChV92CR6UUNIlFVae7gc4RORw6vlzlMB8cgimaTO+Gj4raGG8hvES2BE
a8yBrgUK006V7UrdJf3jVFCMU3m4VBGDtszoq8q9DDdIz9EWib8rf7ufPfA+Si0e
QcldH1Yi8ZsOZPjDep4d99rwZbm8zq4Uhkn3OCYxGNFEfcIbeAnKPza50R29Tuln
P1NxLenv5wh0WGxgVetiBZ96cuGD1qHtmCZ9Y8AfSEvDqZ1M/r7HuXmRM0oSDQp+
W4rqBsHI/+4n/zHTPzSiSFMD3CwfPy4g7kcxQqzlCTTqHwqWCYIx8aYnaBAdoai7
lBSeC3pRO4SbotK32WMvQYg0tFdZGQpBa9aSg+u9fVRiE3EmsjjMhiy+f+jHzNs5
5zBW2IZWELroRmhMUkvB8gKPUWuM1IEcoGeQRaAooDuvNuIiDYHOlpX1C1MbXeIv
1ujCtdC+esTDREq3YgtFQVxvTu4bQjVOyKrXp2RiSpmvybTK8cwgEsF6+oojtJZ/
vuAYfGYjvPqbXBe1/MKatwiUCiwW4HCla67SrbqHRTPP0mOU1Qc3HIsvUsuxK7Ww
Doy39rAf8ubTHkTwdFlAerY8o6xLtBZHQs+fP6ylxqouSH9huy9RFyLSexOcgHiI
fUeu8p048TRovIuO3BFI5ZyRDSCRXfxjg346/32WG4b689oF1xaFmzA52CpA1fI7
Jb/lsDzmoFD2Yc6bVuLre33aBpmSkQYK18SjWs9l8DkhfSNxhRmIZE53a1I3BkPI
+iMeRSBjZNejM49JGNQhBIT3dkQbiJACPfUS1Wh/C5u9J5oGnUehDRUo1zBRVxg5
39rCXFtt5Uvc2vHGJXVjPr3bo7xf8Nf8nWQgtECnoFT9jUNftYSEUcaAi5DTtROM
3V9IrMOpFhaYHWp/OcyJIzjtINKbmrjECkRo8vQPvLnjn4gPTGZOzQ0bF+6MXcii
UM8HqotfE8ogkyfe3kXOfSjm9AwYifcJOGC2LFrS5ACyBRVo1OzoYzLYjpnuSx+v
1/J9ODVujiP68HFPHpTseEUghUAOwEN6X4/Ce7nnwyqax/hNu5X8SSDEjfppBwVF
prsipXqrnxNfkLVYsCIcUtCJr/i8Jq4o4neHWditty6ADnEDmeJy9XUv66VbIBeZ
6i2s8NS/KXte99mO7LX/AUXs2iNstU7J4PY6QDsszcj5WrFtF70l08EFU4wcMl+Q
7dwdrI0Vc+2ycxMmFHFO5UUNWmV4jBaLugo/Hl3Xx8JHLzk/mpXzYSYaY6xKaUFy
3wUZJpxNkJ4HYwWlODMrq4NKwUYs5TVUwpl/rIyTB1JSQXZO/JWwOBEFUICQLttR
z2Pxkd5ECgYxBfTkIFBwg75nv3dyJ5msOpH4LD1vDRAoJgLVJCJFh7ibOzOlNFXP
9OOn/+T9pyNmMy52SdxGQClE3ht4BPoIN9AQUwHubi8Vs5JC8P+4ZCrdiZM7SU/1
Xh8AmPpX+fv1iE6FAISz4edlk08KKxczDZv9Xc4olxoWV5+ZaDQNrNTpPdbq+TvE
CTeXqL9YPXwcSP+ux2jz7kgbjiqmwugZMeA7EA02FR9QsRnQ+/+NeOudUvXQgT4O
j/BcZNP5SkKrs1n36nVst6zV/F3hAbMFSorVZT8o7I+htnBV0tQLlbj3ZP7Gc6Hn
uMwwNwQ3SIrlv8l4VOGSBL20nkbiKSEhYVBtxg2seHrwasZTyLuVGUV/we5Po6DY
XLfQDmtmxJE9nN9NktVVwgOFt7wBN/hu+oOQ+yF3LuH+/vm0slncO61+VeScGUOQ
kL3OZSWOzui5c9/08BvaH2DeMNVDJb2NqBzTYknBW8NBfWEmtgdUbqz3y5mTdpUA
xxZvgjGPESOAjI1oVSFimYXIHHtFBJsnb/SwfBmfwkljIYln3dHrASL4dHooQiC5
qqRjjUpHQ4ii2Izgu4YeYTwRiE2EETRnTOUE3JW0dw5rEpn3cY/lc+Ltlqn4tnd2
heDPQzPczwS/OKRijQwosnrD2JDaM6W0Xniq0y0Bv9kPjfvHWt9f2Et/GBqABZ6/
w3hd9fBAEMW3bNM25y52vSeEgO54L4WpknFDH14p0fjeiP+MrsptvUN0pbF7IYhl
GFTuFf9ZSsXAwu3cHVgfA66CMMmpos4kmy9KUnd+6P/oMI7tKIGdZSXz7EfscAlH
VtVsKkTupDU88r2H7U4Kw9DwGx1ViDJtr80Hiz5ulb/pKsd+xLGDL9+kTr2d8v2G
BtUNWY184cRb8+rDqKqJz8/WRB10FMG3kL/BTX+cqUjnNGZAv9qtM/lQT6aOsuNg
uEnyLnTfTa0JkSmzs+aO5DOMfMjwKOk1v3S5Wb/dkUxYsIzC+nGHp7c2rrqoxtuk
WZgNM5x4sxR2EtHyCvTg234Uw0+yhp4EptOxG2qjQFUBrUU071kc2VWOWV1Sr4rV
lEcSF3Rlj8ZT4rbqMpfXwWK6gJ5LX9ExDG7UZq+UiP7woYyMloomBKbDaGyyNU86
0TY3bx8yTzT/EW+ZPv0ssF7+Egrv/vbTT0OlLmwLMT/2efx7fkt8WiIMlh99yRXN
9a91ByGght0FMGOvhoCNhLGuH4TXZvpXSqAVE+7cIZr9MysGedFbx10NdVRF+9un
FDgS7ybQP6+8ssOw4uBSFoogNW8DfCf3kdAsXQBVVhlb14WDkrsWGWrJSwZ0KBn2
XpfvHnEm7Jykv8rjUcVT6I1pP23+WnLY+HW9U1oiNiwfvVzf+ZCz0cVB1VbdssbI
Mi2XIMSBlZggN5X+Z+aeaWQTcMax0IWP9E+XDfU9sDDFyzAlVqgpLTcxHhBzpPLV
sSD2jPwiPxrVQXxCaxmWY/P3TfQ0ZEH7/0Cvs7V2bNOniwXOuEAeVHB9TIGwPfRf
ztG4JnVLhlXslCk+MA6AWTL/psSMP3XxXmtpZYB6eZyBh+fQJag2PKLHENL9Y/yD
n6r7N2eHURRu+82ikl+JRyUCrAxZaQeehgOlJ4SCUAZb2rwZd1CAvq0OS9JS1Cox
/1k6EOVLvdUcwsxm5k0l4QXcqd0bdknkmjHw+/tDfwOIq61MzJYp6tUh8nTbe5I9
4cnCfX6hgZMg8Nl4SowKtfHz1YFQy2qfdkO9S594UgGaSwAHta/apB6+PzsfI0eE
G0i615e3+T7c3+euAuA2Gi9bNdpnJ/k3qwB0tz3ehAnlfDx4j8dQNIboRuJ6+RpR
BcPrzd8S3iHMJMV7U0fpWalcmLMEX3TTzaww29ZJ7rh28JLGXkB/xbp34hvESanB
iNqAw19r5a5eb9MgTpv7qaB22yL7lGj0zI73tbhzlPcsooocliYXYvbKi4/2jE8i
bkaYWFQ4UJLWEBVxLYaWl+AUelunptzdPWHrbu05W6ybYUkKjJ29pJ6QlgJLWuce
iNtPlxFhbbcoJweqf9ruwFigUUXpbtReytvkkxo6us1OHIGKzhp9eEY1c0kHNUR8
0s5/VTJCspVh/jN6TQbvoWoh3lwKW0t7FqqC8wIyHaZ6WzrD4j6R6nVQarB1w0vl
xePZXPBJE/xj+Rze1Dz1D0xzA+DPRbdGt2HgerOZZ8UMMD6yLwfC5AxrvkJIqyZn
E9Xw3erg7M/86WM4YVL6YT3vBOs4jdn1UJ66fhOW4zurQpaU0DTSuts69pVxK4ah
mbgluYt/v/vz05XckbXlBHriMRIM/xoRfvSzcySlVnRuqHLDkXqRNq9I/qr2bcf9
iC8vqL7X6jYSj4V/vKRSR13X2333Zljw2hwmIVjigmFswKwxG/tXyTB9S57Ki+TJ
y7QFF04dOz1VvpXkxH0Lg9lJgicHvJpy58xVccckTtUW3ANzYWZCJqL1TsXPYJdl
iy0GoOVqoLaSu3IQ3cg5IsNthQEiXZyB8ITI3Plqt91JjO+Tf8GY2pQMI7Ft8R/B
L6Bk6MPKFmeN5CCQO9volNRix/2BYZfQhvlccHJYlzQRwgNxDiQsKbovOpjh+QFc
Egl92WeRySuTlrS+ciB6nSwpIbkpOdkMEoMhYw9RE27r7eS689+7ldPLWuS8/Blz
Yw+jBer30vxC86g6OBixy4NqxIl03fPeYB9kbf7xYeQl+P6GmNV/C22dh9kvf/Pd
Syn9tVoJvMsfUlu3fSNLEDjwjV5wjD0CBawbcgMTiaSKCSuoorvz3C6gs7UN49F2
SfcAdQCFMsfPtc8fpHkSwO+BOXG5LrypgrG/PCcWh8eaXO+YtGlvnPpEDXlaUoML
rB9XlXmOMvVl4OpuPQusobm+bt6oiay3Y0K7TpjTXSKxC8Fcrjz+2EX5OaIFvBO5
okJWVgqAODfVq6zAD2yiyV3InOIFMi1o4S0VycWYbPu52a0QtRw/FOp392WQbzMO
yMWhfm69kuJu1IxIu88StTq0AYQEMKvVLrkMyfC9BRLhZjdjcODobPNKlxSzafum
CnsvNGgvst86UGPxluJ5KT2dJnjNR4QW/IkmyXpxaVs4rGTA2qBBMuiHEEvOYd1v
o8m8c8CsWOj0RHBc7eDZ+l2jsEFFzwtTJXsPbjAeWtrh3UmAYm78jV7un5VbtGGo
oLM5bUbDD5CEfrrqz86WBKsuzFEwXA+myBFtJd1sj1AKLxzQ7wgCWewZenv2sPw6
hUT5FuhvirK7l65azgiUOGWm5UdJoGhS1AwccE4TfQIJcWpJC81xieDqgBJV2sq9
9gRP0l6katrh/pWdBuRbQ4h77FZK4jM/JAVXAmT7TatOIIJ1nu7LoxlS81joBIaO
d+6BRpTPqUfYN935yHa2cV1a9xn6VOK0Uww0GZDuxOUfAtYhZYZ8+Gl5qzh3trUU
olgGzSxMu+JB0tJqSpl4rT80q0sMwcjMk5MTOukQvLnPaB2BLeT1vWg7pRYP0k27
hr0Ip6JS6Ajcm5fmdShvXknELbsQI2/hqLuObtdzEWTjBldu1UO6HpvBrYpEgIe5
nSduR8uoaRzf+D22+km6qF3WFzj660S5InBSU/AxESG5PXJCtvyjBCuwL2NRGJKm
q5xfq+s+EW+4yRtRhZJ1zkPWZUxUQ1xQWlvfhIg2SLKl8VgwtNVCE2eZsd/YPkve
Bg6K/godEXUMz4MVJTQU/dEmai6wiKt/MDuvPsm1+rNaTok6VfqAyEs/p0X4dPj4
3cjoQAuPvZLEWK4Ml+zBpZWeFHCeHGsAudAmF81fmPtgvurMeZF/48cjGOS/wN8/
v1P6AIiXGkECmeFrwPWNuMjilVEbJJ/fRck6KFShN2n6nL2Puh38VPa+5BIRP+PK
bJ2JGNaS2JUFUjnpILg56WSzMMaOebEoFyHslJ2i9QV36dGrKhThUoSWymy1bPZ3
d3eX+toRQPfF02iNNOu4jbjO7nxM7CFZJ3FRQtjHBUGzrVRDJjImTCuHM5RAZTZe
krAECSUqs3WEn5esziCTUxu7jbFAxepA+Y4TeZHC+OFR2uI3BhSXCU6wN3oM57id
TLIBwUTuzeTbRsg6wA1iT+XakfwuPMz4aEeC7/EjNt14IMDMHIcUtMVbNoO2x+t+
jAJ5z+REQk+zhxFAfX+5SxWdgtPeZ4BJ0Xd6TfBCFayjpcCgzp5EQcVHMGWAkw0B
//ZniW5qBmMiqpJGexPgz9xP2eUkAym4arUWIq+gD6MdzttFf1djJNaRRrUw82aZ
udAUOWl7nsWkrulHhFt09crW8MxFS2YcJh5qh9FEpuIXKrOOIqtkiAdBiW/pjyqL
femC1Hus/ZXWLFrPFxtB4K+W/A+nXIcLNi0NMM4H+gshUdCkDUpuA63JJg3o8yip
hY8vvUq8iISuMCvkCHRUeIloZuo2Q5qbAkmIR87dpI6JWOWMGRNimrVlBcVPXqDq
t/odHvvcRHBj0vc8LW6jUR34dvcNrqsE0nICFdHMWRAiTBETDTcTvebenoZ2q+3i
IKLY1fuMkZ1PRMLTpfr/MZdEPwCpUT3JCUqUx8oQhUYB6xVGoHL9rj+s/rGiYtLC
HJ9oZEblle/I0InW2xw9nP12tNuDR0LLZ7lvlDiXh4iJKk/TF5+HsviN5/N1FKpX
2sOkn7L2fy5Z8WQFUEZHpS0oBjxoNAN3rHgGFvaZlNyneY9yCg+zI2VWmt7nOShW
wvL072zoejVPviQUUVlM/ieT8s3hGV74BTPA+vYuW7wrPS4/STPn7alYgIPKftMm
5BKmXgQjEhCKPYW8o+/M+QqA/Rk/ED+oQjQIuIJrMIhh1LQrNklZeVk/5s1SB7/M
6nKxb39CTVhG9ir0GUS+5nKXE+rNySLtilJQ7hauXQ28vzPEmlHqtVIgWciRm98l
GbIveattlQr3LF431eHTpFBLWcjTebPGyXlpyB3mr2t3zrF5a4TnWVN2b/Mo3XoC
KcE4gcldUh4eNDfW+okhisnvU4ZVvQmCZQHPj/UA9Cn5hewrnn8AuZsCySKkai+a
0FUT4S620ln2D+LJ0z1zKuX/Igxl0+q6mxQQYBVAMYZMgi0E3kDNF3UvyVw9LmL8
gG9a8iW5m7oodKxe9kVGMWKRRUaWOU1+bVmWB0l2aS5vyD9kQmpop/KxOSVc28p8
MvWccDUL8bzk6DnEf4XiQ5ZNqO51zl835sWH1M86IciwqkuRcWCTJ0/uWhq8CeIf
nq6goXBQTB57qwIGl0d5Ok3lpK17lDjQOXknRHMY3Qbsi2qrIjZz4gTf0GHj0ZQ1
000NaTp5xGuATKVEN891P8EsPV9MlKtkFpPpIYuuYS4BvyDH+BqKJNcQsvliPYRN
ZkNYsKJipkfk8dcvxJmX4NjG73NcK/RHvXIia+VSNpxV4ghbqVrH75z2Wh2U/6+R
a+UKhNpuDQlWwMOMVdRsRZezMn/odWKqZlQhhoAguqkXb16Ry6K7sH2M0ws/OvAK
uBwMZiMiNoI0OejfGP6cdtH2CFLI6Qktfngd5euwTeZz9cQAWrhoNCjMiKszOmu6
dnybT7K3cq0PhhyobQjxVaUlu4a/6XlyascGhJvXiznlVGMgksLiZqQ8rsbMerWP
gJsIZNZsAyltdHBrlpKdbTN7lG1u1jdeLlpve3ezMDnNdV3PKUu0bP1OKqMwCBH6
4RzfpnIFVuT0gpMLKXFBUBSNPPn4yTtrDyNwq85brcShoMdJ/6ZO6Q/cYrWShwWl
Bpx7PWwL+Px4ZHGB2/ZD81lAx1rkwiLPPoj3WCp4PeBSRRBFyxa8aWIf1/niD0/j
s4pWzqnAP3w4K2X/TdA36kru1WWwSAzYXXU10scJvDUgPcJIfexzzs1/Gl7d2aao
5zbFRArPFLj/NGvJ5uBIUaPVILvBjzue5nZdMz45fUwUy2ma1ChnusUyG7qYD7Mb
THZ3D6Ft8xzNQKbtJV0m11o+TF49KDMrX+b2XdgvhKUfwhAc4X+siQXyXLcQYjjY
Qg+XyO8GrTaVckIkyMGBicE/HY2lwM3N15NRnszrN5VzVI1nsar4QiP628hDTMow
SJu0O1OohrfVDUeXEGETUSd+pILhw9UOYa7+YZxYkM/Qcs8JpUDOflspmN1qMHp5
GEKYYTXj66FQxaCtccgWm3hIBfm6kV99NH4Or8ZxtDWR0EL20xhZ0y6XGP0VeYJP
72Wa67ErCEOd5HlZxAt+2EtMGGCq4DotwEfEmfcDI4P549a5Wzc8uJUeYXgMjwKk
MCzC7nX+/vcOcDBociOjy0PbobPFJZov8wLnhFAheMV6kWlKr926brr/W/ctPSV1
wgb5QbWc9wEHKvCT5wqTcpwzY42HnejLm8VWBsb7FHO4eo/yrSq5VXvxUUYRcBDY
tnlaPb96SGr1hSz6GaZGyle8Cec9ZuNOfDthjxSfXAAciIP3aeE8QiHnG27THuRf
+7q5WMviWtX2XKSEhq9DlYi9Os2fqGlrOnpyJKrV737Zbt1n2j1gMbkKPRWf+lzW
fH8DXCYUZQRVtYIQ3b8+nuPj2n+QMa22otVZrUJDyjgpLCmAS2xuKq7svqQC2gB4
8keD0oGvp54mL11WO4ta5qX97zkZZtY5RcBTziyA231LcZ5j7aUtIPB2G8WhdAIV
uNswwc/ABeOcuV8/oS/SYx7z94kfKFEz3Se2CLCw2VwVhET8B6RXgfEYs4ZJA7Ff
stSk0L+ocKf8aUdvscrzOsGGgytrzqDP0d289VYsB3KXnB5RV3i+I7+yOipyYJK6
WloeZeRqY8ImzPlfC/PTAGV1anB5/T6rL5ox/mLFubADITWRrjFswqPZ9Y6hQaOu
NMNj/Oyep+FSFLaDHsECb6FfyUoRl7FjQ2tBUcNn6y2eRBPb6OWNz5afS5ifApka
O1gvulrXIqSV8QX/+Go/mX19JpIqLFC2kFgp0ERQo/+KxNYINRV2T2DIfKZGXDPV
+arCKjHfJY1rXWj+HHpuW+99x949X5Am3duFlsy6v1wRCQ4bp3T8ycD786AIMRwB
K9bMHOCVRU6FFXvl5LXCjlVj4ydtrnHbypOffoG5hGmrw6TPdL1VJ5jpSYMMn9Lb
SrDY37/SpMWHLjwsuQ8EspaOGmkM2an/a21G5ArRsk+jKnumHVPEhh8szHTbRrG1
xt1MhIdxZ8mqaFD2l8gYS0sB7oVbmyVrj/2Fcz1E/mEzwA6dlNvfyj/2c0vKMEoH
0kYbtrsVFxqvQ/6PEBx58W+HkAwTk5DW8O/dAC7M7sOqCBm/k8DeJxrB+AxzZpH1
OhYAkqwHkmhAwPS0edYgfktayzxcl4iYOIPU6L/rfF7RgdNOJQTeRChMRQ23k4Yi
lqWTWxy8H71zMkGfftuM0IGCO+dqy+zxQDXEWoyi2WzMAkv+H+jDG3sUzoHB0R/l
H82IvO6+yxz4LaSkl0F4uQf2ZZc2aS99lFN0K2QYhj9iCkuoQ5gqTTIaerXyj9ga
g+vEfFbYaNoF7reXM3srIoPr0vfaTsC0JdI02s9vVWP8AH77OkqlDyu/kA97PDcA
Z+4ztN7bEAJCAgpp1u2L+dfKqPLLMUuGE1nBWdYFfSkiC7GbumUf5MaiOsvMyLbV
LaNMK5/L70wqbTBbGLAC+u1H5J1GpQE7W8zPm0IFJ6rtXb2zHQweFkW/OgQELiq1
7t4XXkkREs6yDZIwEOAngY6bkhWI/qhRhn3SkKMV+gNcYDvUbnMfGzUM18JRFyIC
vYNeW5Jrdd07UhJ037PE5AeVgGQrIhubhftViWL8uy2j5xXVBWe3yb6rq72aF40k
+i9CFVUc5Qqu/FxH00d6orA+60rJIrXK2uakwjMOvIpQVAKsFYVA8m/Lmh6HpTUl
hQZsxqYSJZyiGAhuZCQL6D5iKMC2ulo0tOv2gi4u8yR8sR25Fy5MSf8w8hH68tqK
R/1rg6hMnAHPn+aNYf/DL4c34SBAirIaD1mjGu4pDmyUh78UtGxzBMgil+6hDS4X
x5TwgAA5rxIkfcfoZ4qlyYYFfSAoKzkcHdK5Tp8S/1be7j05uf+V8+JMSqJcLm0J
rGuLd8dBu8/TasQlwkwA8UOez02HDLCvjc8vNwCBbp/tKU6sc7+MUp7OL+QajWXs
Zn80KtlY9eGz3ad5tEq0oO0/QoqsAtkUSSG2WgM5xaKs6p4uPcq2B1ULwppneV2Q
g/ZwbweK7WEhMLX5SA16SLemYHRvYqbjipcwEz57Ys4UYwpHA+WjZ31+Yx4Kik4/
j8JzaAesvYUfPEZY/An2TG4/wQxXg3NOPCGCFv3ZxtJrb8gCUaX/mkt5byG7DG/f
jK4uVr4XF/rJWP6BuxLWnjLgp6o1W9oLans/N3EMwhIeSgi+ECXAOk5vhIFxUtf0
DKdsKgtC2deMyV5Wy5OK3HtVqMb8xW24yuNsCyArMxFasxPPB4lhIeYGW/wT5iRC
BVXz36C9PSTnL28bsntxfXRcXUNBgoPDsOrPabedZl3NPnexodlO42CWN2dKRutC
lgl/MAdj8siRBQmd9kpbhFW6RC+nDw1JlMl2QbL8h4+2dmB3baUpbYTJ28x4V4EP
brddQ32p+bCx5bcEMvwv9XiydFu7+dn7AR4fiDN3DBfQGkBDNdtG5QGG7wormpLS
l9uEK6Ny1gk4plNipjfZqNUQrwu/b4xbamqe3qbPQeimnJy/c3rq+nRcf9k+/QwP
mTjNJF4TtdGukaVQLMSFBpeL+76zhYBUNNk3Xwt3ZxzszJ6qBB0Gb/kBKkxYVj5u
JMGRbrqlHA1RT46ZT88HF+Tjt/do8qYvbYGib6vznzljoh+79IiMBmRvi7OXepTe
PLxRphMaiTj+LDdQAhIB7BmSCMlz4txAcyOnUay0dLehCAtJXKSWe4XX4XqXuT06
Jdf3gqbZzEkDEseOSOQh+cxWFlN0vmKcOCO3oI5vUCm1PhSd4cAOv5vHFYju8Dsg
66he02MffrnKvNzzO1R+Q/Zv82KRNtU9g1YrcdR4cS9DL/B6Pm/FgwCAvP1SzNsU
GW5DCrAQKVKE+4TaZD8x75eLyHsky9NysqWo4acURFKWaswFABSGLyfO6ajn6sT/
S6MB++ymVzxbf2OgB3fAzLVZ1wEwotZYi+AASdlYh/uqRP4MJapectP6lowlZOzu
/QH9sCnZQ6TiyFwc6LecKT09d11o6GctaIua5r2eMJGczLWhmvAlYzYl7/ZFj0/i
ksJFlZ751Yye3nfTd38WN2jNU5OTOEBSdOyJWP5G6vmdQ2NTcy5YJCybzbR2Wf4D
uR8AKP1SPzSZ+WagEztJ+ZkSEX8YefvLpt54h3SuX+oahsPcb69Np97XJxAvDdBE
irmG7YMY5iZ2XWO9+jLSogBS2wSV9hA+RAyp/YNb3s7maMey7C1DtLBx2ivjb/fR
MekGJbgdUMhhHM7yFt+E5V0RyPqkCoIZbEKyqrzCGWp8dR7ZjmcIv4xYhULK5Y2p
b2TWsf66tMA4NrNgaaeFW08caJEBc588PsQEcH3Z/TzSAk4I844V+f43mZn3AtJi
SBnJOzIVjRYmp7Oe8T8GlsyN9hd99Lj8TtGre3UlVk36eGuQM+/cYO1yXAc3OjU7
/Jm2KO5eOSOlJL8Eg57DBxeBtN7cbUbHO1oW8zXVCEqXG+fbXD7Jz2o/9pYN0Don
wMFmC8nyYM83704EYkGfHGdG8PKc0bS4uxNRV0g6Ec5uWEV6IedjEk1tkiaBs85X
NvjYvdpclGtdHgInB3PHoTZFnOBLcUcKP+cdCTmW6jLQYoUWzQ6KN5Alu4twK61A
WPvQdLAwpSV2VxosgF+ewn1WBJbqBULDeT6LTtDYRgvFfASUleVakyquWC/i+vzW
R6pHLaWmslNp4JroQz1jBOJv4qRfjULC2LsBtQ4Kaf5D5xJWzDNcv6ohEEvFsvxF
QtoHdZzKVH/KzguAVuwM8ZecXhK9VYA8v+whgVPFdSK3nrt3YGZ+szfdVPoYPM45
l06JdH9+yYdsTNkbMKP7BsG7ynOCZJ5fgjRauPasvSJLGg3+fB4PYvtI9RLBBcCf
81J/EWWol+/L6komX5arKyRlaDCdmLw8GH1pd1OC00xaIiZUq2SoBHf+rggbEYJR
NqFK9ywmu8+tibglGiuE8VePyu2lNjTqjCKYteN9fsTJN8DsSOiMFzRnncqGMhPY
FDXnnPbxJLvJYpYkh9kgAt3VyOr2LLJ4nrSwHbKKPEWCWYaU5LopsFg+GQqiOPBc
8F28pzo+6ZUEXVYJrjZnLNDKpqpgZ54zXHmDnQtQ8ERrf3G2dD928M7gimSmktuU
3GwhVGBoqZCqj1eLB1LZqA6wSecLHTg1kbV2Z/iO8ysY6vhYT/r/ZD+8CfRQ2GUF
SyHs5Vb9LuGqCu/FDsVPsgmVOqbBGFBuGosjqu2ov23yVupVKWsz38fglrYiif/T
qSJR/lJe3d0pYDDdORzyo3oF4PLl6j1gwxyaLEKMUJWv71VBLIHMNo0NF014yM5s
1XYUM7RUw+WSGZzqz6Tm37DwVRLhJodD6AujF5EI2SzW+2KsplKcslhR45Ig4uFS
M+2cf5N8e7XknG9sEA0NYAgZxbPCLsz6MWGCCqX0FQCCReJMAw9ODoMrNvHd1kvp
vbiLr0JQkAKVhcoV5aSR8VWDwl9/39UHcb6N9javSOrdpW2l+fhpMlLFP+xZpH2j
vR/5CzIgh2TIgSq2wOKWvR3nS3NwzKr4VPDXv/PFK2iM2qN7fqDIBJctFflqRmGj
Fhp7J8JS/s+FvmQ4cbWE7VmTUTosZRZ0m9avTav5TUgA2mTPBHeDPii/T2GkPFXU
JA63n6gboY7iKhy1s4TbC6Iss7Xo6DY0p9XzdEVe5fotiuWiCtTdU5o2uVvJQ4Qv
8KMtehyM418tZCwCJ5rQw1e/STOz4NUJLk2U0ErxNvjSBaWb6vllf+hDzyVZryGH
DD45YsDU/6ZjGyweaVvTh27z4HEl7c8PzgLFyK/jOrpqgIh42MmEpFA3Fk44Vdhr
SRhWcyNzdY184DKpdDBOhn+rOwM6uXhDdIFoQ97XFz+QeU+UH4xh4DNCck13jt1H
oMbpf+++IPGz4AA3ckWhuVHtGPjN9EfUWN2/K/6lz/R4u2qbeLTbYGArPIVd9N75
6dDe55PqySCcHXzS39+mp2YxxVS5SHNdc7Rj+q+OIrHvkdLF9/EUhhTCzuePdJzZ
urQqHmj5t8cbyFzLLc12TJNEqtX+Quk/MH+UrTYkIUWDZfRvX21BlepdVGIRGSi8
YhnWEd7bzCwpyhu4wRgPU2qc8LI1oYoBbQ5VPhhf6GHjB5GJ+upVzbpVThM/kf1K
LGdSzZbM0GKtq+fmrUxpIxhYp1M9qIph/TVMzo6OQYmVb7tgbajM6PQ3yaCGmY+c
IwWHiFy3wWODcfL1rLHVPHl61+6riLHQReRC2LD20U3ZaXQqdrGpByUMJDmT+Qxk
wdg+rEbcHa6wldjfz/QlhY+5rX2WzlDCc9uG9+tY5841GVNEGuUgs1A5G1Y9xGvC
jlMSH7f36MRy9RUuZKnroGPTXy7RINLCgAX2/HX9ncsniw7UXdoy2+TUlIkRfGan
OgqyLwWHgjLpd566PLfhQhcRigeMIhk8/zVwWocl+ublrg1Iju4rmLRSS7v2958Z
KVzEyH9pPGMp2+QyZfYvnxP8Z+Zko8vOC9ASnHzlnHOPuLPJx9k0OKA2sH2m7fzo
d7tdzYViPIjkGvb5b0GHncsCSFQm3cQYyLmA48ICa+0SlsIJRFl9uM2L5hlTIkp7
C6yazYbPyDQ7mAYT7jbfz+cHJZZFanTLDErYz0UTr8Yi58wBjyUioHOD7JQHofUo
69QWSpNZVBdb+b0kq8VJf0aOkp4OdiZmKKJLlCH9Xo/+vrxcqAW4z1IeZM5EqeYs
w/n5JlBEhvcWA6q72DuNcRFv2us8sK/XfgmgSUn6mGL+Q8R8SBSOhxv5A7P7YAnL
U/LFqZsIu7AFmVsABZfvMOCHr8XaSgl4JB23Sr0h+Xv5SUoxP74PFMn3nrlxhqas
f+qXsj0DLM6bY7rW2zC6Lj//Dumorbvb6TCcsSTpZR2CyyJcOWw5N5o/gI0/MVsM
imnj9LF2ea0oRsmrot8evKudduispXzDDnUpWg9so13WD94KZXnWrkAVYklPRtMo
yMN2+a0mSw2IT0E7UneJrGjtanFpoexJLoXkdPPT6qHF7e05Cvra2t61NS0QR8vz
mh0JSe2hvUPVA0eOxvOllsmv4pYA/5Xovuw42bXrch5ZlXqwRU3pGeaqFVB1Swwq
svhXoFkg/aokhlWEExn22GtuGLjMNglpdMs233VxjtDOKaEZ+CrZHWIS2865vqMV
oPhLizMKml/I3ivqGXfCvxIvgEHQ/5GdrdSbnc42pn8jvbNFvEjCt201YYUo/54t
LtoaYYJi4ydTglPRy/oV9rqYH76+47uNF8rPS2hHvWjdY7GGm8Nf4WIQko2FzRtv
Y+/329g/kY0sskgPcVIn8q0dom6q8tHTX01mz0ucUyHUhSleDrKS9jRdVsI9GgRK
ZGBmUfbEoe4q1x1LNQHXKzkCadJ2/Ws+lyGg1fpMhD2YHTOdblZDwR3x2pW4gEiD
58++Huou3d/GRw8szW9iyJsRfq4oUkPooDLy6ZMSyGnlvUPJT3jIw1+JPXt8K/ho
oTFuoV0r8C+vdu9ccp9vT8Hd1XgqGMKAGKkDtGbHK4ooshP+tGPy1lEPdYx+OBE/
q3YPBYg7YGpfdWpTx8RFOWEEiswy7BCjZYpPjAekX71W+zw3oYfXZqM0N+XVvBlG
Ipm+XRt+/KWEDwYGSv9cyPLpnakTLOWnfFwxrIdh+cRKQI1n2jOBEiXxRA6AdKCX
N1epGE7EA2guN/2KgoHCogJ6e/w11b2HH3tSFCYD8HUtvUsDcy778KIrh6k0GVyn
T3v7oWx9J7PEBbdAwSC0LbBVwZn51bmqSg8IKXw32YUY06hAp7IUQ92y4CCo9Abl
uhga/kujGz69YmNkRRO+tSS9Ftrw8o5lmj6rXmRsD7nHKuunTn1HOUC8Li8e6TQ6
gLFE4Rq04x0HyrhtKN0znyKx4O0X6XZ3mvS902YE0uOJLVox2kpw7Hcftz4Mi6qi
YRiZNCTcB2Cj+nFcaC5VMogNsv97oN7rnd/zDVNJVpgSO4f3aFlIWHXig3z2dQRf
bHMBODpMhgimOJDWFJj5hRnw3cGIgvtdGte76RMl0nBs6ZV92gLni8P2aSsi9TP2
hbyKK0gXcQH5dd3UGE+PdABA1vELWJFhFM2f2CkfSl3FgIO8OqWaZabr76K2Y/so
/TnQ0CeNEWufjKA2vjnkH+eT6cRXcGNP8JkdH3pe4BgawOao5uvPIVieAvDvMi/S
sAeYrvrVecGHKdF9eoCllt9J4ppmBrmxGDaZGFr0+xKyp25Mg3n8z3QJMYV1ZZ2M
9YQbTdt7Vxhk5Y154Hs78vff+8d0m4HUr1B9UW2+th3Hnwajja9m0xdqwj1uZRkw
YKmtht/o87DGAdaozelNblVRjwuz4rqfWfrBbcbyFo2Ie8fnDXD8IXjy8h9rh1gQ
x8vNUko7pZkP0ec6yYjAj2naUA2vc5EGkyH/mE5FZzFz3/qctTHfQqLp4yNnRtGi
q3Sid1Y13PSoSpd5xNzpA5EgYkIyoXqxDn4+Jns9rJsbcbPcwfRB6wepISZsqqWh
en41id1Jqqu3Nkh2zxK/71nFB4mzsdAlG+EJJT963cR6sZYf89qeIU8jQYuXuI88
iDdw3GOcLcrksWGTbMew9NNnZw28jro7FKDnf04kB1E4wYyMWG8IOabbUlLw/KY9
j7ccNg8npHt4WrrYnw2rFWJROL3blELtOr9SKHWYSWZXPNNWzJLqogdW1srAuM+9
dBVrTY6YHzOLrLwkXCGjmu9MA6KCzDpgWDqvz2LuS6aX4bneefZjTGHUqT9KXRd8
mI1NFdlIE7FVOoig5eyF9Sj5EvN1KzitneHh95f94dI5957+Tr/w1xLtV+RgYrmX
Uqx9dYvJMM2Ltway9TdlFkz52LlZZs2y6X2un/xmptZPx350URaldYvk6O+6YZs4
2awMLpvNKTwSisi8+rheaySEasjrjq7t6/uCCLuTyhZJB46c497spI2fWZnr2Usq
IolQVRuSFCya3pfiqz/10oZiLL+PNzATDbIUGfRTzbliI9bdB5fzaLrdvPra6KOJ
GTmdbvwI9AHvn6l2WOtLCpsN6jYH9ooUE65kYliZXl3PI8aBjPY30A6lVHh7+baa
Fh2g6OonTUZj25Ajpdt1RymT233jH5XuSlZ0kMhMokucaALd94ezXo4FHhYo6wT+
jc9HoooUvAjNc+4GZqssDoWYUdCMJ2egPWPxwgTvYye93yFLWNz7gSGyx3lkMoLg
Q6T4rMzdPMXQhPQIEoKHAN2bR26AlkXesoHXi0iymXvxKb8BSOX+ZQ57l7vFBpPM
OjnpnVW+8aSTTGe5phXRd1gEfU2WTuJekhF20/NaoEYvhPeJMqI+eqqp5HFXJHnG
zddzFLwTjgTmCFnNcMSxVdXRfc9yp7UU65gytUOPFO3ivpA2eO+TghdR+GNN4nNr
pzVM3t2gJnNMuILb9jhIU/ze6JapC5T4dPYxdkjolkJ7lDo4/sWTfk1eVfotaFiQ
c00AjK+IPodWBktzmmNRJHCU5WDJf3qzxqwK8nwPMXFWB3qk3EIpHfqPm+WxU7Ko
38/iFOBXuhQSYbS0QgQXJj+XYP3+ol7ThL4cB9t/Cn24oUv7rG9gM764WjxFjN2J
4T7hL6HzW4k9WCv9zK6zrVtvRiMNJrK3Yg3BPAF1gXsmyWkXrOz6x/8UQEMXQ3fD
r0pRKa+Cs2H5FW0yS8c+bQS7CaE7M6ywp5Gj7FH+ba+dp7uHwEGQIp33Qp0yGKaR
BhF+QXImKmqWsWHGO+Emys90uKORLiivg4aM/CNLl5Y0cHl1fN/eOornWJQ7hP04
HRNDspP+B2UfJozLR85wPU9y3oiZfqEdpPELLUV0Jk/WbQv5egksCgzEgFdsuWQa
04tgZNww8LhJx9agrb++cD2P0RMlCA2FYrlPiOaKrMHEA6ynH+4bxWJu8lUGlaWU
l+mnamiyhoGIQ3xqBBzzw9uiqya2KRsVtMK20yu6TEMHaq1kN/+rGSv31+pWI0o5
BhmQGfCtfSTXQV/yh8/NL6IY27E0uaxPQIiHsk2cbV6aycKXl1eAyFFHhVRazSTM
2l5OtPcMPpAG3EUX+a5yga571vxTILQsHNglayNhYgFJ4T56WvapUHDmpZZN79zT
wZQFgy5P+sSvHi4O/pliSG6J9dupVz+JZVLZ5XbF2N09EpvxTNeiQr7DPeT6nRb8
CzHpVzhnPl0Zp2qlkToLclxzYVz/Xq4kBvgSui6RMgE5ZXDdFRSL2wHNgnfEK6B7
NthIh3F8Cz+5kxme+Ttdd3wJJKMiqo8Z9DUhzpfuu84ocUQhYYEiAgLX/EvqE+8m
it2fmO4kZAGAopRBuf/j806cpxPGmgnUCsqgrJMgZKrDuYCNMfBMe1IaKcWv/u8o
s0h3E1b72NICYaTwLOWPitGpGwoY6NXUzjbWT0IKxoXQZyQk6OH02sI3gBpZX6Hc
1Mwt50L6CdKz3XJcsBBUvBVt0qEWPoszXX1jYIF0RQsNs83S86maOl4wwGTnF4Il
isbvz8fq0JXFU1P4svzWJIfLOl/QC/2Nf/4X6HuV8azPF3tyt8xwuHz2D1CHzBFl
Aof+0Isv86lIiLIAwP7YVCacRmQvb1ewS2seLt15vwBRHAZ/YnFLzGRYMolqKMAS
QoRSJhpVrJaAYcjBvhxM+vp1JzsnDM0Hk1EzFczV1F3kUs3G1VEqQOry+u9tIdlC
eH+d9X8E6NclUhln7+BeP0eGq7JjuNUw0KNwY9SwCZJYH4DsJO8fHNt+EPVlpUHy
YxL7g3wcO9PqEI01dlc6gs5/O5bJDbZNplfzTkLehbFOGMNDEjbzAozbyYXJV/8S
ghUV9HX6wQWFQIWHoIPXrzV/JbiuV1tdCQ/qW2OFsPDB2Xov6JP2UfPPBrtrZROc
h5LfxD0y/QFb5SpMJ3uxJ5UEAq6ZUj4QYGpKXXlSJf3B7tWC81WKZ099736/fYhS
oECb+uYEM1prS2Vy7Q2xZe/TlT0CnYrTypwjKIiwS7IeFLjaisJOoqOPjEbc5LmQ
ImFvmvidheR7MLtjkANvTzkQhQf4od7uAfD3tso0dAo2gU/Dq78jzOnfIcACqpDV
LibWIjrb6MrmsImMpjSG8hdt/OzH3xs0iArizAjT+WTq4uBn6sWbSgssSxhNoaBN
x5yN1/vtQWbCAuZkIiS5/jUBZIFlj3hv3snfpxIWuTswBcTgLAByVGX45uZuVssj
9vYNnanbz2Jaa7go4Wgr0Pg7KjcLLvJZOsX/GxCJDOt+/SNJeY5npE7gGYeaK4uJ
Fl2OAsvltIvmLbM2tB387baCCaElBF+g4bPuLWE3z9z9ckZain5mfqoWynPc4nqN
YKw9jFN+TYIijez37kzbu5MtDMg4cm8swvPXVRWwe2WcRmPaQ7m/673EBtVFYLrE
AT/6GDnRz3tR1reHbrNU2yEhPfP2Ffd7v7N1Ay6k6HeH9XtGCIhFEC1hdIF3cQJ0
nUnQW5k8RiSVtMSh7qOPvqm+mFaaSafj4aPfmuLYrECExQ+pFdS5EGhV3xcVTekJ
DSt3OCsvlRgFTp2IkP5R5qQVDRaAzUFu1vSJO1RnU8XjK3AYOrXsMi8Wpx9IAG42
fukdIqRPOfoifyank1Kn4LLfNzeuaxfD4HE3D+tk2QT3xAtnzAuUQa7KyShCp6xF
/7YwD+mwWw7JiLSqKxRMej/CEorcNdIjVIDIyQIDhHMRSZICmhyXYAU4ygzL/ngp
yDRrFOjb3Bixp19RK3k9WALleew99WFUJjlHmQ1M9wAltJYGHx3PiQFTWuAR3BjF
wGx/nuYLfmFBQahA0z1CqFIlxKYteLx8qyxVl4heydSVnIdI6EmvqnvJvRRJfSjX
PHgxlnYeh4dk/IO2Hf9ygYAuoh3VaJn9Yn1+gdzYQGZ3w9HBIMuYRWF8DiuQtOYQ
6GN/N+dC+HKTyxMoFolJsomtxK3uNqkxJ+4SJQmV/DMPWqm50RA7uI38c13i+QqX
7iSMVi4Qr148KUEldTUtjGs/HVbYMfDWPdpbprZqiB4vOyLmKg3sr9r6V7w4mbvU
YAu7Me/lGOGXLi4HHCbR8WfODLLra3VkdMj+e3YxaRwxskiZy3UTv0Xa4C+SZJKJ
pv/szf1J72DR1eECIh9v79B1A6a3pTu1BxjwxOGmUYbP7ETJo0a/w0E/9StdSlgX
cq0Zmd1Ox0S/z0XSNFJwA4upT1QzCIyZXFVJTKfiACP94yVun8UeUUHjKG0v65V4
GTDD3Bd0uMwGWBjsBVaRBN1kY6TLZJ6c2i6jljJuPu3J2rh0XPnGfKBx2DBQNmOM
oTmDDlB3xFLi8vTNHYd9yqIYA+9TPmbnB2W7IhEIvBi0yuGZPupfmG8sQVrkJv2U
Eyxhqm5ZtzOeWEoLby3wa1pm3+LoYrvldknGQYMP1GJYWGaf9Qf3BbsYXaQ5xazy
1Jd5pLpQWAx2AKYhA2FKxc6uVyeGjJjv0BkIYCoYjOEKx+OwDcSlUhgNtuVS9HDj
MB5ixh44AKue+GWXHdTgUspBiYtWq1Bcx/LRbY/n+6jSJfYoQSCth+obODo/ggtT
nx7RAr2bdL5KIvoLBITxtyni/GZI3Ha0iA133mDiZDOkPPjHIH2YPcxcrSO2Z5aS
QmIPKP1vzmSxaR4xOqIFoIjRCyN5K75aMEp4df0NTP3BEp6N/ZjkTBc9rmQvQS5T
d1NsfSCfD5tUOr7wBTrePEqq7D+zbtaYDELts0SXWxMmz52PDTZoqekuHrt8WYh4
f7iIHad1ypX+4lpmZM5vEohjJrn91WFrtqMjwrkFin3o1YSdFBP+D7kJgabyob0S
k5c3b8eFVuUbqPaUhsK2TaK8FypSCzrXv7zjETrZxSh2beZI4z248BY+UKx43FK3
cuPSQ75HLKZz1SkV1jds1XDWkGqNZLkKc6+ga1+TjzPGE+J5DDfy5JFMnvmewZkP
bNinXbJ/UY2VOLXIcAHdgnaETSUAxIwGw1v2HnqtK0KGD+471GDBqc/1F0xA0WGt
UHDVJs2O5IoyUR0kDW6/Z16LAB2EMI6gUK7e7i0i14G/KfdT06zqRmIHBkI7QN1/
WheyOzY4/UvhKqphB09Rlxo1yOxNtpwdt2WzfyGsJieGNSK/5Lf6wXFaYW43zu5x
tejYEewDVQtsVNyPB5VbKLcboCYevjqIx9vdc+9xC54fX+Sod8MDfB3lmIiuQodw
IrpAo2hAPe/B0ju6lxI9olydbSl20q945u8B6K7r6RSZR9Rnov8zZL7Rdd0JeMPK
zGPNB7D/vtmeLGeAKRNg8zy/kye+NzpClZBQA9JM88h41jr159X3kw0B00eTRUBv
qWFO8HPM4UPGFC3eqY/hWa4ZITaLlo6Ft+ugHdYmgXF9IWbATua+U9JAJ9PNe8+j
HBPFIStfxCB/lPEPSIItL45oohGTss65n4rpbh+NQxIR+BzGpximNFYU3VJJpPpQ
RVH0vnKNIdetg8M1Zf4kgJAaIJoWVnQkwCSJYpVuq/K9qYH+Upvhk+ah4sGjLoK7
mXFdoP7yudUfBXbUlcRHeIe52n7GrEpaF55lQtYRy9ckxGtwPnPaPq9exIqFehqG
Y2ck03AHi+VhBz53F/6aPO3Vm4+o0zrnJBXvt7i/rKkhe3CcTRLZUiOPHhcKIj/f
DqMI/dETfJ5SYW1kbjrfnRJZd/PrcfaZGBtV1vYkfKv6QpAlvqe4EdJ+aClTNIOV
GpKpLvnOVjtiwJFM7dA327qDlICdplt0tx5L1T7X92FESiTCOZ0WVwzZCio+lcae
xiqNBQYyrEsOp5LtcXowcH3314A79psXFOeeBxdvIXOsBL2YTGYY4V51/y/4typk
+IaKyguIenSa+OydulBZUFCBi+WsDaBfq4FEulaGo+0Ba4Y/RCKcZBhAfUFF4lOW
ut7jAAQHYEUlcHBap+DcR2WSm1QfHjYr1fkx1RPSwLcekY4FoeG/UDKYWQzX+Kth
z3Cbcmk/q7GfKTlL9f/PE5aXuLRP0/vIWTZpr33OxkBuyXdMPSu2q2aFpqj7JF8Q
HqwD4xn5HvRY9bDT/Tn5yPkxmg3MXPTFQl4Z4/dWnKffqa4FqMsVBpH8gpfa6d0y
yLuonb9k9UViZXdJdzzd7N6F9raIkKPsR3DfLDMzYz1Q8Z6LrPTtVnKkYTn/IG0x
2Xa4sbI68qumpECYB/TTfrfcsMo0kXczDi0dYs8QoM3l2WdfQHPxkTCm/+oXZJ6Q
coxm1xNCsiuNQcvZMfN88nC0gYAbc0JR6RRM+3hHJMD+fkPcFdrcAf/ltdD4qBYl
3nWocAkKUPCYHmbVnXS1iw1WEeOx93ch03Wtr4N6lsMYc1fo9cOC4D1fTgvx1GfN
BTo8CLuvNn8Fm2dxp0M9oEkYuvxh/AVaVqSNsO7gIoYL5T5nR32fnqdA0sLXt+Sx
FGBSbVnV7z47M5WH6taE7Y8pHK4Ekes7Dx2ZAH6vll4akmZ6SURLjTvpxmETSk9s
iiX6kOGyZLA6849pV71636sS1RA+lrHpshgnuOYKR3enredJxMNhBqy7YiJq8up7
3SXNic6Tu/RAvsCgW8dXfAb+dZXCcDErU2LMNgWen33GDtE7JFqzALI7MC0hVUxE
jjexFrrHxHzZwecZJ3gjGA3pYN0pRhKzO/U4aLK7HvkMsQwMTqw6goCxFWHaBs1t
BNYSfxvvNoTQpyiP50wqHkOFffssnaKIDuM/2tZ0AWEZmZfgFbpUon/W0VvbFxMv
5pFOWt9BfAmWxWQg0DvSCUjfdOddWvpD16wNn7sNlwaFwJHi0AIqitetQy8Fy4wE
lJhifiPCQ1jG16P8/O4y64cYNTY+pDi97LsqH+tx+ybsy15aAx2J/e1ls68xaBSV
9GUvIgyNaDIXctxIdEl4PUYBscUSABupTc50T+oUuYZafTFTj47PbLsaPaBMB4V+
u4qtRrnn4EaObrOwkPzs4emn22z20PtElWlOgGkMKvSrY4MmLBnuKznaqqCbFX64
Ojis0YwKoN87ZaHIisP6br+Sx1gWxInQjNNNyjZxSFHAJds2DGakDBWKpfKgvRa9
hWt5IOhnanzcijQ9odb72XspiMZ+xeJ/k5MET+epNOhfH6O/ScbphscD5WGNUIlg
JpBGdJgoDqXaNr/Wr8tFhXvv2xlpoWoV8FLEPXIxs4X0NBYp3CXs6d7QjB7XbAAn
GI0b7pt4xjf6z+euN8CjOONxQ4zg3vWEv9+7BOvfqxzlE3k71gdb/MBd4FH4EBEG
qlruVVk3uPiI901M12i2lrC+4AJV4fBu6NRxnlCsejGRNflo7Vbjcm5dNs2O7pW9
4F2Fl8/SMXCxvPdKIJHGxlIMM8eUNAAxg9eKbkH3LtAFYxYhfZ0gzq2mHqBWwiIk
8regYGcWeaIV1tR8DhtRpwZBvbzq1Js/keayyEPDJ2T621pSALjoHUVtx3oMqggu
t7KzAfUcPbiKRixt8HHR1r+Ha7pVR548sr2vBETWEnEa4g+ndqfONgP+sRjRiJAu
kFTJFwFFgbkuSAAJo6961h14xpWfNmKMX2AJDrSOF6RQwZOqjYDti3qBXpR2ck8w
UqzMh51I0Zqzy+Pgf+jqkhxWtJQiG5QCRkSq0MQioNKpQalCQH8QFpu5fLJ7ZtGx
r2WojW6lfflKJNZLxyhZpQs8TWu3pUS+MUBxbo6pyxFZ4JWExGrlXr7fBLJCBm0O
3XVRk1SzKFEv8WRofAfk79+DYue3y3nd6q4woBVQlzZYzv1e4ZP+/ZXJUsXDw7d2
kuI3Km1BtQhTDZbC/3wc82FviwT+Jh1fq9pi1BB9aN2RnwvXfpIcMLafzfr+T6Tg
oMCLztMcwmWYpizU2NjUXg63fzqCesbzkOGPaDnQ1QwO5Hym2Z/EVUIa8Ke2xZBH
OyIAxeTx5DbQHIRV8vxeY9D2l0ZvCUkxrdENpWmmoquEjhqqNU1Vz7zUO+8EhAUy
FDAqBqP6CGIlBN6wnfu3i3Lqd49z6eAlg77kwtLRtqx/+YOtrctB/oKN7Z0EmIm4
PV26RL6gvivHV78HhWyw6KxHUdm7IxlZiuIlcqu6SaiiiMM2XWJW+tIguKMAygwP
eLGYb2F69r6XZ0xIEx+wcfh/JqAbfV6rVfRLzConpRZHT/o0gHlAp0/7xq0Ysn4D
bzBKx9z4rrZDwcXII9DgeTl/gPjGRXiZmYMgu9Z4MdPNQBCc+i/wiznWYEFFt6/W
xss9lkZ9YdsJBzMw94pmCji9WDvtZvpxDiswkklrZ3DDoCMLcC87iTv8y5u82arR
Z1cuae3yPqRQIY9rd/TZrY5hlfv075QoL6gyvy/x+APOwaOd4p6zCH0SnWlWflqB
8AkUq0tMwbny35qEQmV4oDZEH4rfiw2+5iS+p5XOqXH8enKlk8I0a7MYIbpEIMaM
JE8XvyzuK0lHyZ0qXI0r2fEJJXhZscWvoTRG6jfzKpQxQXv+Hd+/OYGTQHVRgldz
UnoOGTAMYxtJ1kuv9nAjyYnZU4/3/7zcSpHQUINe8wYmKLjtpknNdwph5DTywLCQ
VLC9ABHxAschCsqUcI0bXW3AP4bOnbPRfLrDTGKT2Uy1v+4ogwZW6dwHK5RFXjzO
CbT+kYyxHPVD5o7J2MzP/9ctyr5pfFSYaMn4OkjAM/NKIbFnltWkY9xrpNb6hNPB
b5XYlPtm0g9aLLUNEm1OoLiteSicnxv8JFgibBSsFg+oNZV8irA7be42FVL3lXcW
MoSsRmZw7RXBafKknooXHoTb8culvqSr3qNA8HbSHRsYl681AhxOBE7XhGEZjF/6
3ZP57DC7/VGcD3hgIaClDM7VpSMkR3kW0AavJ/KbGjvAP2qCePXmLuNNHSx45B/c
/e6ayrOV09nTU36bHBhH7L4CDz8SJpRrvAWJmwbiznEF3J4vdR6QO55hi+FKt9vc
dOFygoIO25tO7+KKtwmYoE6UEG+foD+Pex/2NN4za6erFQnbrcQGCorqnBKTAEVT
FV9o65DgLLwBe2Wq61xaeH6Ooa+qd4sIFWSOj4R2nJXtt2oqF/vJQAmTt3ooIY1+
//9/AmqEbQm48jvIh5G3oiIzcrU90l8GDHVh+JUL6RHdajZI8W6cZUjf0A/dQLcN
GEtV6UqGvS/xH2q2jUAzIJ/vKBPEhIw4Oy5RgNviSOSPdRzkt4KDRLBu9Gr18zHu
MPXix6ulQ0SSZiD2CTjkH4IqhWCw14+roggis7dScz3sn7DOXB3VvkZ2LMxoSEtV
EE/xxWjWBe9NtVX5J68/M1GSq7uus+sVEsC75nIY9z448RtTNh1P7c1o4p73Kjn2
9ou9TrGFYAm/nwHFd0UCu1Q57myvvxHacq/WqzAyNXOxDXEchjiwIdbZZobeYBtE
bh5O1fNwyWZ8MoOmyGVEq8XJg8fZbBCbjknhX0uT7w7RmR4LAg8rBhT2Y/LNsN2W
FlhCRhkDynMxe/mRvfDds1TnCItEbKd2fbiNUaLqtRSMcMxRBaPf26KKk1K/Th0F
W7TvKxbXLhPuN2cPz3kGhtXk6MPiI9nu9DAbfG4SwDz+mS7j/kd0i6IqDqLTqFjp
t6oRur/QYYCZvlYQwB2tKgi/BgaxBadhyisrj4M9ORzXav8ywvIQtTi600k5YnIp
mKOYiRO+t1e9/UL+ERkYE3DlW1zWV8zeifoRRgROvp3qQV9J0kkAxiMZGpxlmGl+
TYML0vlhmXWrzX2vmxaHGk/9HhQrnW9zxnBMQB53f05dcGvqHiDkuosIKZsNCGVR
PT9UIodNpXMngRwcvTFd1vdEfxQquua0MAT0Sw1AJrUqLtkiW1nLOXDUix+euTPB
F4nrAp35p0dmMJfaOwEtnVG7UQxmmRnBwGeUAS8swmnfsVCjE/q6lxmH5S1p6IOr
mw+kdpRidf+1zBG4GY0lXvNSog3HoPJPhcqAYOLRM7mvKjCdsqAhC/oYN1fKNO50
6a8UjuoDkCL+apdvGWdDsNdnlD568kQ4L8K+f6Kr7jCNRMI2HsCKFDFcGVQPNWHy
vNju6IRHUhzzh251VEmeIOvz5xY1IzM1EusffSDqPG/GnZBzhxsBwHi15kXI+qsY
RIakt/AgBdh6ZhnsKeC6sEPYI+2YGuAdizZaDyEWVvh51C8Qrhbk+CPgqzEFkJmB
a3KDHI6lD0jQiuV5/m/iRiZz1s9ro3hGSlhjywVmWKkvqGRxud+Ma+W0OHIOvlHZ
PZT71KSX4/cuUnMD485sq5ANETjC8PEgV/PP6lvn1i9ol9Jsiq5dm9XAR4Lo8LX2
wgpJE0lZLq9CHSz04IJO1CGSZrc3pzEsjfXZfr8hSUA4CANB308V1CkQEoQGPWXJ
KCegJNDlDcNBMUHDK1ZA4j4QrVQaaTvXxPz+hGByfbEHpXR3MnfGFO0kA4aPyK1O
UdvUtU3Bjsk4N6ZsjlvSDVAzl7Uhbd+zrtwVTkl3YtPtlMG5whcaduY0WI5wzwqq
nuEh9Q2HUzsODgY1cdH8eS2SZbKnkzVtiPKdPvRLNp3Woajdft8PAwHU9CdMSvpo
fWfagjsbuvj4HNDR+4VbjYwdmxqN1s6FlCfJudDuLRkYl12Wk3KyKpnabrf90uDb
jyqFAf7BcDLCuvSrmVTrxwT22ooCFz5HSbaKI+0W0izzH+aDxFMFKhZ5iBMmX/1p
8Dalg30iAMpZ603TOnUbmu+EoKQ2ikYZuSj5ChD2/KpvPil3S/9RVc5IV1T7g/kW
rBzghkE2WlIbuj7ScfbRU4goDmlev/zMkvbSDPXnn8HmDIJNSJxCq1A0F2Xra3v0
vu58rgNbrz1xZS6F/w7p+42Pp3tUxfcIZEyPmqDkeEPe/wOB0Bd3W5hBACb2hyFb
F1Bp0L1DZHu9dXtpIv940yxO/qPymxFiuBJiHIvHxf//sW9kDnZXNnRunEmADkID
MCHIaPL1bUKDatqnKHjvRWSUEAIHJY97rap3/bOAbwXqIiKN70yOfmWBS067M6b/
LNB8f/gip02e4dS9VnKOUdIS1Jn9OESQ9MPKeOCYu6vGBLtUomc5Mt1+BkPfkQlu
V7QlpC9Li6Wxrvwylrs299oI+QR2UlKW6JaPtn9bSDCNefqbebBRSxBwd8p51twb
M/gfULzBWCpeTd9daqqzYZZsCJwK9eSaj3mH4Ma2NN2JKLa9hU4iuOWGOYH1OvhH
rZdHZgVufARNhHYkSGWfZW7sFRy6wfaDcIF5kUW+o7e810rQmpN2kswlMWhGet74
SwNSl5Qrs2yhqZTNkby95xpVazu0zSUn0oQOoiVrLZFoLqT1aYdNwxr/hncmSQRl
6mAlxhnC9LHCvapJOTpYMudtKt51EY/l5T7r6Xs7vzPe42Y/IMb1ZB9oTXAQFeT+
n45GSkeaSLuchToQxMYJs7L7F2TfYawFV0qmRH5iZWE9NfOIpxrQfuxv01lFy+wT
/vkqG/5C6n8V4Gc4paZNp7nAfJ/5fEEssQblkAQMr+S7d1/G6D7yFrNrzktPAHvB
Eey0XCaNaJ3D9+HxPkrU7ZzFexdbwMLKVLB/hetawocUhZ58iIDObcyKm7n9ig9J
qFCXFIuE+CMXGSiO+rD3P7f8XSpd0UlBQQF4OajlfgfrYGiAgjZePvVnbUw7ZFCY
69VfUfQJp+kDoXWvNVrtIf3PnmTo27U6SxjxkF/nSsqhfwQGiYsJc8VV0BhCjkI6
jFIjzo+1tjIxlUvDHBved8k3P4g+NgUDws0XhUE0fR0B0BZlSqGhxZwqj0LLhXTG
nyB+dKSPJE+2A5jhE48TasF+LQN15GVgp1nji7jLaVdtbifN3B7kcm/G7qQ81PaA
zsQR2Nd37vfFhdZ6Kzs6OAuQWyl1QFWKKiPaoJlqIQfaLxt2aj0sj+Pn8i97Nw+s
mW5VcEakjJEiAErsok5NcqMdNLJOK5OHrvyCdNiu/r1tS0MPpRqBVXGvvveo1JCE
H7qQzpituwjGAlHBjX5GJKqO+9eW6bt1nrKZpeDjvTUiRK0d/NhGrbMvt2Pk8ZQv
ALQ6lPUlDoevd351s/QT7hJR+LIfsCbaRZBsbsnnI/8aVkRBznCTnbFljKDtsPDg
fhjhh2EXOcOmY8JWl5TeFkJg8CT/6sC5LXVk1bKT/VYT7GAvq1Fkr07vwj5iSkDb
U/HpY1AcGWfDCVhhSijUFbdVBOyyVqW6Gd6k7oGLhQKahlJFzjiqcOuZ1sS2RFGn
/orItjugkBvnwGXOyxLu/YBo7vNmE4NwVfeL6CVG1e2zIjAKLq3OTamcbAmhdfoS
mpRtOfBtAwlWPUjQf7TU/cwhllvQNANGDJ/ayZml1LCH9BBX0FQyY0iemPWMB9eR
sXCg2ueuDPpeuYwP3MfBzCUN/8WRomR68uNMbSPQKuL6qiTYyAhwSVNnQBM7f5PY
qQjFMqRXKfsvJZHH01H3b9z36CSNf9PdDpzk3OCqFPqRWuW9jwKW+Z/S/UBMXW90
ox0dIHU9lGinN0J1SbVsz/t5OYcsqhOMa1rxKtdeuUkFry67WRNo69cXzIfFnLE1
8TDKaB6ZX3elbhiqruCzgO758/ki9SVg1GaD7pBiwk5PSe/gbAJrcukfmBblPHLy
+WzQ0RzGDh4cW75C+w0aOtXFrxZBHzrIQ9rOY1+h6sZrmY+O2iRzuZRWi2hxpmZc
sBJ2ENnkT5Pi/OIjGIR3f/SNzLu1Wh6H3glC++oSq6LbAlf16TCXyQL2qWGGvQcu
TfsxfrGZjx1KPZ+/O9htkPZ5ev4l21Wy5K0tvPOx3D/4RY+xygLoWMmPfRHYOhsx
JVmJUz9cv+lS3I2IfKA5aHywIXAPxn5vtMX6ExHk0/zTXzb8CIoi97s0EbgEyvJe
/CNy3rBLg20fdG0mXAvv9Ox3m3I5hOpBZHscsJmaXMt5QwBLYMOPAePSlxjxlEuu
Fw9guiE9XJQUTXugVoVw5cI/raIHZYiu0BIr6qPYEtjy2wxONE29EYXUjGfSPN3D
LlSF1Ka9jPYAYor9iQCUWQkTaPbBjFp+TOqzQjf0aTeJV9XChybm9KjocoarLqnA
TGZaeQAITx+ZX1sBNsn0oSJcjXy3jP5YivzZ7tljASr7uOGJiq8Pa0+5Wr34CnfJ
MpoaBpiovej3JU+rgO7Am2JAeNduEEMQkgXWyWuoAxyeUkCWuvTOZaLNZlxNJbGz
haplbM6WhwelGVV8pX2L8xQKz3+ljvinNWYgq/F7e137my9dVaaN7CKTFAJPjn85
XHHwny3pknwujtK4t7uHyKmrz4Sb41G0XFJWYHJQbeG/Cuu/X6RTZknt9c4K4enT
Rko5pwFd1ivAbBzju7yWBzTdFYy0g0YQqRnxYMWsFOpR9IlA0JvDeXwIYIqV/QHv
+Ds2lOuqdClc2dWkZoqQ/xo2CQUKK1Mc/8MJbkJxkZUt/47wlgsgRfwWALEhOgHx
wPHjricYOoRBWFDpFA6xC4kSOfs/5AyaOhYXJF4qJBdzL0zxKywMQG5cpgCcpx16
pZqepnhVxc+MOzzFwX3WeR+oasf33CjxLCwD++l/sRn1z4TRPYTXKHyP6GOGpkzo
O0Y23TLqC1gCYmSlSCbo0ja/ZIELRvCzQJpd0qX+RezFerwaYD4xd+k66IrHv8cm
U+5dckKia4G5cef2G9loU37jl5kWPxZRzl2QE4q1Gqx0wDq//kFztmZGaUpBNWZ5
O0CcG+ujFUBuSUOMhUW+pqh5u+CGOlBJiEDpa7TzIkfhskdRQXL4jbb6sVYuH724
GX/kUZV0PgD5VzBk3PnK4ZKamPMC8GJeoi8mN74Tz5/a50AkkmnDpZTxcC731CUj
K4g02N93c9AP01yDUN7Hb9QbpfmGNDJBl3Ix6MDfy5f/7AruB756Zizrv+gsD3kP
SLe7B3yPbwuQkp1cvtXZIMD9PtccWGnU8s8CcFc+CVsceDI8l//SqXVN9b8uc1TP
Hs2F4la3nzS1taw86+b7A9ER49+ZAngfQeGheoxV6zCasqIV7rIgjV7NmJjAhYPN
iZn/ZQc4/WbktZneWFWaJhvAJZ4YvS3mAwdbCE213SGILIr7t3DadzHxibO6sBhw
ZqlssPYKoqglCpliWGGDpqAsH9LUZi14j2K3iR+bMYB8J+br2gFpoq1tBL8tnAx/
eThcAsv1QQd3tI2vJsjHyxc9sdheromiT5OLVXD0BLWklonYyxqbITP4koYy8FCQ
H46mrDlusJOKOmwAXRWBOCGYy7rVevQXacLVdquWBnNS6gZQ3lnJLq1GL6QIpSvg
UteTFdJkB6svqqUbkrw64OFOG2Iz+6nqNq3x/9yJ7CtdWen24TTN6g6tJGOvrrRS
3sDtWHppne3jZUoxEPUZP7nrW3q5ksSW8ae7PhBYiCOBeLFReYXLuZ3bS/NW3sJC
rcVwfDuTP+P8sTfbQvQalHytU+l2ULrEgJNHHAFnwS1Mj3QizZJmVIrdIPRkDCAO
dMF7tT5chktozTVsKpY2dWaczG0j4yG2npQUUNtIJ3W0m2WalCYwU+wooVk6+5/9
nSX6OT4TEAbNLmNWs3sm6c4hgpFLMSxuLfXtuT57wbK85faJ8Y7MeTriKkvhEBTb
/d5/GsO+//woXOVxs9IKY7NkE+38xR+CcFDdicGBwiQ+e4xiPhZFydkIDq7ng0Tu
6m4ikwJsVsvfsoR7gwEwNqAbaQSdKOMPpsCo7sxkSLihrGxF/gfdn3vzz6t6kD8C
n6qf5hxtu9ossy0i64X382EnnshA5hypWnyNm2Mx4QaGNkeiGU7pMn7uSTKD3BTm
+lUk/4WwWuYk/Olr5ufksNNi8ucfDOAMw7Rfel8YWL6EJnDCtjSYl7EUO/c1TkX6
/+mgB32L6u5h9dXo7noFl5CjDZji2lrlHVIXDtA30RZpYGl64kENQ76z0NBuMDfz
fgVyQM1gZw18cJEEI27GoEDtNbOCUN2MYdXxfFeUYvEHN0mcZBCT5+0s1ApAtBjU
CzH7XagkX+4t/zIWvtS16HkWbepE3MPEKKNDwFAtzrMhXbkQRRfw9vb0Jc4WgKYy
IC8QdC+JljsxApJaUbPQYzguSDAxcV4V36ezmYV+tHy++sKXPfjPXz3cIDcyYv6q
lcoR7z4L54PDZEiKBXr+wQkRzPTgoy6PKT1nW0t/cdJmER8R2nXkUTgu4TPgxqG/
5smCegVOX2D1CrZRW7JXzXjLE39rW6+qdFNvFXpz+Q3J4ddBm+U/UgJQNBTVnwXD
M7KwCV2jPlgVXz6HMRyWgKz72SED0xuB+EFyL8oNzsfSIQ1ZsVcfvclJKpdqZDAw
N7F3ChSXQzlo+kIYx+uVOXj1lqzNAb+/1IyiGigyg6I3LoUxQTbsy5msFy4J+v7q
rWY5H7oHu8qr14m3Mm698EB1yaErPp/+gTZENhOaAt9Z0FFPAEW4mBW27sQn5QZh
gPARB8+FYTVdnh4WY93POP608dG0yY4kTl0Zb2Jz2vq5lgO/UjsYdH55Q27V/qfI
OatTcQ7XFHaeHV/mWV8rDSCYITv9iVr4PI0wvhO9Nw99PUXTY7K8p28CjhDiEuAY
0FaSz0mu2HtUX315xbgesgjAjH6/sszVUvg42V3HLvs9hOOH3GMAhERmg3PHv8AP
p46wu/IT/8M6HTkeO0QTXH0vS2DJX6prl9cQ1VPZJVwvW0Z4ba018NKf1yaNHsmL
aDAcSvFR18eFExyg/LurBgUt4GSSrNmcsCJ9jwk6pAU0JptIORwa2sfQ22vvNRsz
YHu7fE/yr+iMu+ElOYylwjMnj5hzskJbfgPMTWIBFpkykQZCOO3cYVNx0kVo031T
SrJqI85GqAUs/7sv3ef04Kmq/JkqXTuxlQePeavcouRK39xtbaw+LEwnGUn+PG6G
8SsfKoOSHtSIbVZ+Ns9RAB1WkHmsulBFxCOlRq/ele6xAh82TqjDbFbtA7tjddT7
u1LKMUkARNh66v96P6AEih73YvnsuIudzro5K8YUm2/aX3FWvv1D/pAn19p8taly
hMBUjGTz4+bYnPftrtjKhnOIhgKONMhdFJb1UnPXp4dLsP1Pj/qWX5CsDc6voojJ
rbkT1ZnLTM3opMrE1/PNVk5aHEWrR0y2EKRo+migrFbMPv7Gc9K/C0RjfyZqVJkt
nuJybATvHFWTS8rAyp884YEIQKDBnzLEjNbt1RR+7YWsC69fytplsKFFxgvarSaM
z7VFJzQgx/mkr7Xp6fnFMtZUQ2tF+KAtW8DXMEyQ7RUB9WnGBiFqS/gSKPY+buEf
QwKGcjDp1Ji3RCEDew98xxrbpy4SzkqbqLc0EI9i8k6NJP45E8ldakxv57gb+xy2
cFrsOdkVAOLHbvNcVEroURo9x3f8W9X7/pTXVG03xcocMjscvvYtfK1YmLjefJpJ
TPrE79S9TGkg4ztTabhwHUG9e/DYzBrKfXdelJH9v6ngUguh3aTyOCdQzq6iUDSS
Oz+wZC2q5qQV1JdRp3YkxyL1EeHh/JDeCbx/OBIEXXxuVlvgzzQBJGFsGV1B2RrH
lXAVhPLsbz7oQLhOw6FFt+P4Uz5CNyPNl7LCHG1SabXmSqF2jPgI9MsszefmRflH
iXqWq2XDpebe2yDrcOUjH81C06l4XVZIs9QtAwFFO5Er/N36kKsr0kdgvKA3U0/B
kmbm+DsslYFSyCG3lCgqHQRAPurI28BNg6jSURakse5wzAHTq4hso31OS9kmIYsv
6gGHyL4BB/v3y/EjywSl/QZ7OwVFO6ouWARMMiJrcqtpa+S/fAV02xpfGbeAxQyQ
83EdF6KYIKiNyMLcH93H+z7JUAYjKuPBNmM4laVjwevDPhRChuvaLQ+lNMwqEAc5
VxuQwheC2fEaHvhHZzYj/tWl2hVQzttp6hVQ8MFA3qB3OJ/vZkiQZg7jpi7kgcOg
G5MqaAC1jOIbabqtvbc/SGjO3nmr1tPcIf4P+9ADT8Gz+wPvwiqnrvhWsyWLKZ2q
zNICFMNXL+6Mpv8iPNpgbuLA0pQXBI8Tl+gXeYGzWZUy4Lf5IOXHY8i7JQU+Vh2D
eH5v4GB2rFUydd/buruNgA/rwkEXly9m9MQHGKjRMYduqcUvIMeSxbkVroP2+ZBY
UGiJS8eqxX5xLSV3uPMWso+R92OdW95ouKa0VUmS7M5mbJ5Q5dLh+xHnRcH2b/VB
IBh9NHXgdx6dRXpS72Mc8clnBw8Y0ZcPmVK7IXc1VNdAPOeP4QkFRrhzaduTK4aD
TvoaIDN8bFZ3nN/rStbZxbpfi2kWqHniGA9Jl8QstEri+5Jc9Xo4ymj/iUNy5Hxm
3tPVjJghNvYCMY293yW4tJMCDuonLjLpg4qaum0Ucwe92kUjsCWRJbuPCVFSTZTL
gjZQRrJtL8j7pQArCU3XCcEuNUqUMERin7SPTIi8le16J+GH5QPtJqEbNm7Lfzzg
pcP1soofe46MML7cjM6XcJTGZkSi7VMrPfC+9Vu6iznpUDLgywD7dpvClh0IztvL
roIb7D6btJepoEB5htvN07QlFuwrS/HawkvogP+mEdm/248cYF7i4nHJlpbY/5ah
XWzkTF7/02bx3cDdeyU5pvOwL6V19PnWyGcD1FR5kfXrvn2ybSNMQLH+c9h1cSmC
sXr2bVx5ezA1hBmpHoND1UeMfxsNsL8YmFmAZYfwQgYMGQxz+bn9wXMJpX3+ornt
fvt5ACb2YpnNAmy9oCauEpMjeoCOIuIM9ah+zFAa4KS4UW3wJY5k964H1U7i/7/j
Kf/40Mx2dJctWXwc69isIiUUq+nFdxvNAZAeR5EuC653JiBOjbM+etgM8gdUw9Up
ojqMAqeqJtXgzMcJT9Ael8dRf93oE71KLJ6TTYdGYfCPWNXHR2cQ2Ctw9BmRZpQ6
BNtKd8l/mLdhcyot/8oqFW9I9NlcY6eesIFEpbFC3zQcsGpxRIcjMy0r8dG49Lh7
tO99rmC1DRpWSVMC492YvGhkghK1Z4MnIDNLFqaJBZJAqZSsyQsxjFNU9JjHLxwa
wVOBHzS8I1kHv4KVBiLLwpwhj6VR1sZ68wkMMo8v/Y+h0UBkblUexEg+k1G0awlJ
t9f3v2V88Y+OmPKFt3RUzjtI5Uw+Xa//6kyNxaeRJLHmgqKl0H+tKRyb9CJn+bv5
aB7u56y3uhv4oEn/5o5bDp71qwQZAKHLAm5hjVBMw3k8aKUUHtomG0Y877AVSaMM
rB2u4F136h9EMFprovr800lM9oRRebR9bjaFpEHbpc4VWMJS0o6od6KjEp0LyjXN
LxNgPV8fw7FfgiDih6UC4+aD+c5dUqGkmpbF3/Pkz5bamLpHiwl9CqgmPP1BrQKu
NI/2juibvD5U1UMJfATWykmwHSkzrfqoClyN3M2nFOzqUEqsV02+Dbqvr/9yenGC
bPY+dQRxoXp2paiS1QENOUu1sJb4gwqNiZCS9L7Rz1aOHaiaZAl6tDZRrgyHNZBu
lCkb9UU0/C6TI44yQFdBoAMb4XhQw4IEmh7nicY20yLqNunR7vrmICPGuZg/Xl/+
4bON9Cd5nzfV+T0TlG1gy1c0S6n3mDSDk0qObYRw0X2wgriUKAAKyvc3uDNACwq3
F37opgAzAI36qUn9b10H9QZqCtt9BUDcuTU/DmEf/6bcHeJ1hRLLB6b0QAW0fz6T
yCqLtmvWpHBK01G3bymk1yL4scoSpQWF6y4jY71EPq+kkfdZxm+/EU48CoMlgWyf
PQx0RX76mGE60w0z0WCwcNRyirRIHYGtbQ8UDqXZqaQ3LI8Yrv4aKmZUs21L2pni
44TyA4Gh8Dm4QcFxIkA69In08RQCqt0GF2twKKoOI0qJhyJJEMN+jBjsdIkbqXuq
p6e34TKrXn+Lkpe0E0JRKaah6hpqF3sQYwxuMRpqlsYA6hWFHRUrU2pZ1MeSB0AR
a1st8n8iXcqnfYkQ+MLPYxwXVZ5evyPufNuVsjjFyrCSnn54LwQR3GYEp3EmcY/o
vysEneDU5f6jRqAdyE/kwMY475atzFyG/3fS0OF9X+3Bk26Ov9iEbPQ4aB6e2XgI
RHpEhOqZF33JhDZ9kUY5qaIFzNQMGT5TasYwvYEJSwlPitzoJLxdF9oSXtXYbIpu
npJLbyF54h/eQSloid5rbvuhy+zsTPrUQ59fpgz2CFcMNbBD9t4mBbxWQ1mgMgCx
Git9C6wN28EeJWdkFBA2UuvI8y/i5mroTmYlKhwzA+diAI/nJWxHRbcDMkXbfYAs
9/KYi0jy8dBCXukipCxwGPICQE0lz8/oxugePBoJMymd5XhtF62z9IkmE4WBjLlD
ZMqbrEJQp3gCQFu1wkSjlTaD2hzzUtiHWimMGK25Ura5hEl1Xd3pXXdWx+kazkuY
fQFu7Fj6DHwxEhfeVd07VxCoR1Fcro4rBJKvcDpVXpb64ZLIKCZC82h7j46qeoG0
+NInlItTUNqlASpn7Xsygv7N5yl1O/IqQ0J1m1nBvzh8hS0k8rV+blS8XCoB4WR4
zV82kI8XzgWO0HQeHapwpMZ859Oi4lOmFUx8ig85PdauK9bVghs0M/iEMcYU/zNA
2DWqG6uMyBm/U17Vb9KXX9sr1uxfXlrzMjYefNH0KhHv7WUaz9hIOS0oIfFphwg8
796r/DlmaWzfHpp1ogpAetl14ibprnk7iqpS8cgxX7nR1n6vNSQQA8ztQqinUI99
N6bepMT81RvC0Sub+GKiTLel32r52/movpapVRGSmE0eAtk2fx6O3ZAODzCKtb/j
yngT7EPfLdIIHBajPKt/56QxWcRmibbUkdT/yVWSvMXg2QAGxHpkimVHEHP4s8lf
yP7uU71QrfF3y3jJZoUW/iQKzwu6p9Wi3nZ/mEFrEAvRlYLtjYBxRZr0/HNSt8/8
3wFfWX8u/f+WwexnGAta8XfhjxK5otJN08LvjmSgftoLlH8E0Te7N6RP5USDtvmM
cb78PFOKOQFyLdZLnvmSi5THuGAjCEsaqaiuPzYvIrkjsHCFzowzytKUm2QOxIl8
YupIGQFBIKrFqCJiqbHZ+IewZQ9Fq4Ihi9/2QLnGa4mg3YwDtOXOKy3t1Q1xhbtm
ciefnPD+FK+CiOZYnDKyELUpFD4vVWb9hGeOsPRXmYXGkrWPqaL11oINRcjOfKBg
oB10FfFQFA3X4dsDqbjZwahIwogSO2bjwmsZPkfX5iZQWWAiJ9yw3CFYLYlvJ5Wz
Pu90Y0THOBZf0TzmeA/YEu3HWWeA/YHWBvQyOdAOR67K9zr0rzK/7vkiQXoXVzUo
0cE8PV41RIivCpbM86fwKbGC6hIppwH7EVesmoTc5f8AaQh4u7Tfs7tZdPFdI+sv
VicD2/Zpn268QJCJBjmrId2NtH+vHgzDwxK7+29RbQkKSub0bbFXDhIL9LSl1rfP
SjIh+s7+3yuWfQJybjqHAWcCWuUIO5Wb/2B9qn4s10WcRzSPFOGhD19M3CFoapU5
0z1aSrIVTCPO56KzSP6ywRakdWT5tZKxTVdBwP7bWo+3Tmaco7REkpsaQRyJYBc7
Ceebmc3tMx7NgvGqj+4ocxopmSFstmxix1k8pjGdyU5q+JSDS/D+FKaPF8l/IS7h
bOsb9x9bJYy8slBkAug66VJY0V0w4/ndo/aWDp5JW+Xlpd1OpUJ0MFXqD230dNfR
MIq5FNi6z57BfVbnVqQsuFoa6TDsz/8qXqUkotgYDHgmpW5PacekRSDkGBPtCMxY
Mz60pWX8DbCXARLBHBPCdqUOiZKHJi74ff0Hj+P/YO0N1uTK5hffzPLwWzj/++CL
z3jdJQN2yjLtMcmooHWUyQAXcmmZw9fHVn4kNRLpXI9AFbsdDriQM3BR/dVuGXcD
NPRC9+qX33sdQ7uanRGomq8fOTfnjja10nJqjLFzTjL8GDvusmL330d1ou8huoZO
I+NHyNDthIiyqwto9xAMNDLaFJ95SiPnwy6qtSt88jDLwEwrujNBkXJHXJoTtg3B
2FcCifKQnoQVSGgEjYplCbqz0lAvNAb/GPs0T5JQS6K5W4i7p4SQzTmfd70Q65DN
jA6QdJfzsGMR95YkePS453W85KPJUQSXfJpA6pPgwA3TVudcKg076bV9z1X14XiI
vzWJHac9k7N1rNJOldfJnVQ8zMmGpdDhR0pus25b4snFjgw7eWiQyzHqLXEyzkv4
WTp9kMhSG2PVgMUDre6lbKIGNTqBEjql4NtkOo++okm6+Co8p/G2D4s1vIYBmawX
zKS6AlC421w1hVWvrCheRUeiU+FGLNvhmfABxR5/PyNZlKS50Wsyb5XRO63ElcNg
vRfZquWYg0LVK6C556fbI+oEakBA+YjWB6DmxM8hMCalUQW0ewKhGi12/KzmpmK6
8LkyXl+VZkyCYB+T+P0EIls8X/faMFwLI3AVd7h9Xc24tVoma9Zyu7aJiWwgxC6q
vGkNFg0IKTMnkuV645b9EwgN3TKhTrKzOsNq5YOp3HfPqi7Dz+PJvGZdW6G5H2rU
ye7Iogv0cpHfoquyT9HUG8Mm2CjOGUCV+Fs8s/rGZfZ2BsozDJi8ylz9sdpTTDSj
1Xxoz/3O1+xIKwm4PiezdH6dEtU8P3l+RlMEmmmBxxhXtVdwaLxsN9QfV3TtB2us
aDzql+DKDD7ObYD+TiAX2jSMqE241MzR2HALK91gXzIATpaG9DpeH9q7A2KukHZs
Uulmac+VYM0sXoUZ27F8pPs9+VVeA8ByCyAbPqmeEpXrE9CQJ1Pgr2e9KnViFRxm
IX7sD5fe8vo44+aKNhg9v7qzGXcIzZl1b6MIUBAKsxrnRiNSingczKFAlPr0f3be
nc38Wzlf/k4O6G5wC71lrS9cRdDH1UOO8PpXJ89AHAcHKnmcHG/iEATBlXSb+TXm
1IiPGqj5/OE8MrBg3pEz+OiMwhI3hNj1Csnwc6e+RLyxmz2q8x9W7DoNM6byhLyg
eN/qMX6KgbGBKAlmifsJ5akpxcu6PNym5UBigXqsNCi/pJSK/cUaoPt7gcK+tXPo
n2kq6s0/LNzsLg3pINsWqkc1DZH8TF6nm2lAT9fD0ueNUBAS2ms0UTBzi0KUocKG
v7wOLMFGgOMJnZnPSwhkptxSyqGoN2tj+suy2RKJPQTyUBIa4Ed4L44tVnmk41V3
NbBzukoMrgeLQDIQj3chaWEvjd93f86W6dY8JrhGTxlNiD1eGIX8XsR1Np2l0l8T
P+KyL00fZDHIxIuB5bI1POX15SNPWsPDtxqhQSFAeuv2E7roUCUc57loTyZCUO8S
aVmWTESongRJctwGXsPYEImWn6S27wahQTATs8DkG6L/OgRC6d/28gjmVb1AQP9Q
kLKv/ROQAvl4MQ7YVQoM03uxJq4nJ+cjQ8BTyaB1s0FcevATmIvq9tntNMQ2dqP3
vNARtAsQjj7R10iq9RtjlJEYPYAseeFeEB+jWdL29zDPn6F53QG2uTiMgCrFlotS
4tk8zVRa7lMfxIIM6iWOh8rFhQw0nbtXFdJaHmCIft+4OzF7ObywfQMKp/73V28Y
TYswNjwDsSJZFSxSPzXJflBbAUb/DqdcJdWmVAkUYUhVDOVZkGkyXeGeUkr9vjhj
UT2e0JuaOfT2Q2bclckSd7PWgaYS/tJZWlOrqgoNca1t+pQBUqP6F7W0uCG3bpLS
FlVTp9UcuUN1VtxQFUlmoP3eZtHtfmomB1xp5GB+AWnUWomCcPHO3uZx86XOXj3z
H5q2ekK1abomURaZ8BQ+wURA0tN0WBDiReZuZT/U/wgmPJvGcEpIIw+Sr6xblkPT
KOoc9H0gTKrht1aeEM7D+mR0dnbGGciZWCcPg5UBRu7ZsOm+vO4PNIHAY8VxVFQe
bpkRM9d3Bqq8rV70w6o788229c6ngBOeOe6pMDC3T7QgdMiNG6QfBh0CSlKoKD+M
WTbumiZIC1R75E0DAVfrLr68jmjgvQoJgdNXazdzJ6IUUpQFnbqzx9FApkysBJJe
bkIul6f3NLNpOJ6hbJ4u2+OZgaQwqLZ15vEGDp3Sk4ZQxOFq0GilIPpdIeqq7LG4
ip3tnHSGcoCUi0HIXf6SM/bUmE1SNpgRoDNrAckzlFFmD+5hmyg2n6AjU+ZwxEr0
q1q8LhN+sLwe3Xp8CZs5TWJkZ/R6H9anToAmK98dGwlzD4vc+uxkCmAQAc/PQe4v
LEribGXhebGHyTqrVTOJ5oWKQoeA6EvBLwfFDnNPvB9/Yu6d5u278JcyYNn9cm1U
xNyIPhRnEq9MzkWkXQ7fHvFFQvMNtKB3Ttv8NP7ZndSMjENDd+PNRd8397p3BDXh
vVVDn5hQIe6Ow1/IC3ugZWZ7uoFvBM1WH9OUD0SNn7qbsYNnufIpRt0AeCdJtvrr
An0a8XBl4gddV9XGmJGi5rBu43C7ATFvRsMrAYCtUCJL/Q09DTv4surmouCUm3Vd
/L+jROegZnwJXWy2xdg8BjFffzTCxNUBu84fUAtxETQVMe6KgIekGhyInOktpT1H
hVBtQ66zlKqWTVkMGvMTCca1Zeh97dTCdk6NOQX0YlmCS61WUWyKJjRVBdj6yXSZ
9VoVsJSibtbHEVFKhTr3fW7u8xctbXqZpOnNi+ZtrATy0kcvPNV1hw8SpQTdW0ul
tWqju6HCum2yo9/pjoekiSWGFAB/dEU6BOYFIwX/Loen7Apxk+hUa58dv9AwXbdq
y47/H//lXSkfvx6H0Fuh7M4yAvQT2Oe/C2KLwOrV+134VZ1zGcJh9neXHleK8Wr3
aIxZaQ2hooRQoQuLhyuba8tg6SJtvHwXFMw4/rHSa6rji3O0x4r/NIhz8vlXhvW+
L3CTjTapHnHyqxg4ZsXrlP0Mkhjwf+26meuTYMkV2zyIOgYeNqu6kSh/WZ7CmMZF
2zgEbhlKMoU33Ji66Oai9E58VjnqMexbUJwS2VZZutK3idzUsLocovkYhDYYPLAG
qSWsBDbRSuCPDASCiEUAwZZMjo0QE78Yq/brBNH/kjQ+9xteO7W0CUhgCZewbifu
dn3aePj0Xhd5eopZDvyabvAVfnR/eS3C6eKrmcuCS1iPzlwKCV+gkVISNsy1Ncof
5eI78gRSoZRstCJ6dVNjmkjaeoD9OrUIf/N8Qdwog2pYQK6aHeWtJkf7OlcNk6Zc
EAf/e/H0bcD9KB/TSsJDIlN6s84j+YC2bfUsogT2X1WVNMivBU+BQS7hbafgZyQJ
dLloCoPs3Wn456Q6rOOgduz7O26K4R6i/Q9kh/6hrcc1hALi6TWdDczVvSlIjorD
lupVhP7HHoEMrTkUDru16Z4crJJukqRUWYgpR+iU0BJOOipvO76VF14ueRyjG2Hy
gkXQeRP8Bxxz9TNntcrpShGr8kRyR4E+y+PWfQsXPDOGXob1makZ3jlzGPI5gNEQ
xgzPPV1UXvR6Uzasc8sv9fH8FQKZ7B11oOYbgALERDW4w6fSXxUyvYeILWs2rjkt
+nrtyW8iiKheW/XhVugS32TpCXDIXHIXQIldnqbcTG+ibl+qBtUFLfBhUfPXlczF
Jo9AaXRft3FK+f2P0SHQzmvfgcDAI0JY8FO3ugAZz39z4MlRkwIYwgiRT4wPAWID
pGzm791bPy/SlRoIC/zbTlZ8kNBGi3m0P5K4hhRfK2xmaeObUYhIzfRiQ/NJ52Rf
6PnhcPG6yMppxrEYjIF2Kx58jPUU2DoyYtvNJ6bTQWvHCmYGg7+RaDHYT3oKvgTz
NC+uPlTkOlob1tzpE5Bg2LYjk2V0lLzQXLJwYevyywdN6eFPb3wxJ7lwHAXeEQCr
v51CLOB5ETpb93YL/fIf1cZiT4zXLKgZ4l2RDsE6C3WyuL0ERA9I4Zhgfw5d8onr
hIKkeo9PkqUyxRybuuipuB+i5986SmZFv0jtkG7XhUr+M4qEqiDGwE89EIyhxh4W
bsCkmLgXWoHdl1Cycd4IOH40y71/wrgcKdWaxGYaajQhcf9udo1mjZgCpiVdgBM+
9NQG09cpCNvCrsoAXlXiP/JVhdr7N/z7GzCwrueFfSY5Zhg32b9dqzZ8pRKaCUUr
aaIUypIt+BHXY9sOS00rHwCrOB/qFVYcI73IhuuDrryZII0isOwkVPet0SuPq+S8
PjmWPzKtcFqFmh3qQ7mZ6yYStLnzOvvLRF3pG7xuKskBwlYlDJxlTW4eL887f2PE
kvSW/F1H3fdR6AUeRzB75uvhTjJU/wBmb6OadPHHNGyrMQxWwJtRA9wr6DNn/edi
wXN0ACmpiZMPk1KaTtHSUpt4AlGvhAOrv1g4KopcNcGmCWFQ2YAoj/ZFqLBWJ6zZ
tb2mrqwVXxZLXKEY2jrjVjFQhypa1tftxuxaZu08z1KTUob1M4Zq9skcBaau6Ia7
w7TvXnPEb/Eoew+W5tPqfFT8Qi5WeDaTS36OnOxksaEL8wjurQcwEjEGHLxagMrz
kVrDk3woWqSv7dq+ooWQ3gWYC24GURxf/laImeHwXzTNp13XR06V24Jcy11XvlFQ
WZ5XKtX6atDYCsVsdIxaoeRuQVsoYrGE86IAmdfn1eSqdWC4uUwMPTbQqlv7Vxj1
bZ4JuFWoVFiCeGqSGEL03UzwPwQjth1gN656Zrep0iF8ZELoAhp5Vpo39/GGh/hy
PJnUoz6pjpdN/AHUhSDqMM5h2aASjj5gWWg7O0qLv1BbQAZb0ZllzEv/kfRUBJr3
bRfNNQPHwbqWboLXQ0kQcIEVVo/OL6N7w5eRLmOZFzCiV9yL++39dAe88RVyXurP
A6A9KAi0zRdGPhaU50WQdzFwzmE3Y6SsYQVAqIVkdcQ3FJ59kILAjITo5NrX24XY
ouWcaE0VvwK3BcN0WwhQQ77OkFABLeTHZmegjnFKObSGX+77zkKvqRUDyuJjfEWO
6hgMk4tYAbM9vAC7EQWQa4ZwVuBOwh+jj45hek1X84Uls+C2wxdQRsw2LQ9e9++Y
8YW+4o3BPfdFwJrgKFK18JuASH3tPGRuBhhFYgM+c7mgPK7Y4TLjI5N/r8+c87HL
iJsHYZ5iZIXuqMzK/0MXDKxfONxKxUnUMF4eUAopfkgqZntr/cRs80byrlHC95gd
HaZpmEsdfYMwz19TBr72gyQ3yvpF6bGuEsenWoH1uC0G1NOQn8+fTaSkiv6u4b7x
yD9HPtHd/mZ6zHEMaA3BgRGvAiGvsAyp26FZSpHv8xd/zQi0ECZmr0DkgbJki5s9
jW85hQZYCPu5G2THrk5rQpaTf5cTA59vPdrvPwahg/v90rhZU7PTRCFmdD35nqrO
9SkZ3SahMl10nM+5CQpMNp5GoEUeS7lfRymmnxdfh4atpKoyxMUBSazsN1bXMsx+
NVJQXqMMmCODIP4ZdRz9HZJBdBRVTsUrAJDXInMQXUsy2So4d6Xlmsr/ecJyyQoA
607/sjel36lK09SxwYg9PmbxeksLSA7yCStSP7vayzDxfUGW7bmsWVfxNizsWpWc
bk0j5SnfUjibARWwmjq6egFXip1wuNF+D4oftLBOtRPe1BjDRvTcjFyU4s1OS2hL
MnxNBIP/ejS5zLA+9xCzbCWth+5jrFrD02NsYjU4STYzGw4Ni1rZv/mBbcgm9P5w
cbnNwfGJakgrv7h/+TFr1GLxCvrxhESBfE40szDjIdBxypJfl/JLKIgaGfjsKbeb
+xsGD2rL8smFSDfOlU+gC/4z8hbdlsPFW8GERxbfJGY7sMXVgfKwEkzywxXH1FmP
Vu26wijc5ocq3rwrGgF9l7R35sqX2MxqiW59lu0UMPNrzDwjteHIFBl1bzNQclxh
jMDhFWNgn8jh/KzabMMj/Y/pJ0NzDke2hVI0Gw2bbe/suHmO/hnKtG/toudNm/BB
E4GHyMc88vtUmB1CNX9CgxtHU+ecUyeL+gViB0GvQc6PfyLd+Essgf3yIaL4NM3t
VEmj1K+EHTIP4cMC7hY+nmP3kgYziY7jmqcdxujj6OCqOdflNaDYJp1ZSFFkZYGs
O3gpWSpm5p+drX8l4JLro4BcilFoKXbpccnlIpzaOwWVfq6XuEYY4tx6MU6RAqAz
veKxh/Pz43wjXsGIjli5ygLcxgSH9nwUddB/j08bOe8kN6j50VKx4SZ1yxfmwK2P
iS0Hc60xs8wmQX2FWyzdcq5CLowFfKcsQsKFJhPzNf4tNgNxd00Jnly4cgARJt8o
I9DC7fq4YiVpzqvouqs5h4e9QPkGDwp65T0ISIuEoskG5HvQnoyCoeoumQ8kWZ5s
m29GflHh7qJf4sMMGpZQkBRChSfymwhYkV74kMDQMmQ/gCtNagSbyTUSOX+1MuZX
WhOg4V6hF03pZuutMzLDkpN2RdJH3aqfxOrpN8EYRwcs7snek52MK77hDlD91rNf
BLJapwbCjW/L+vmEQyd2ibgvZxp4lx4MkXqCHmtyus1mIQrCLfzr/DreNOPnakWX
SlgwYrcFQ1aiPW7uIDbhPE5sKCvRDlyzxKWt5Ezri77ygDbZvwDRZxlN9W9d2XAh
VVKfVmK8xlWvs+J+NPc7QDtctFcdKENZ/FIV5XErMwkIlrIsTC+pB8jipqO8huKb
cPgaJ9qDpFoNvPJNkKEb+wT/R0jP1Mh6JPz0H50OrKPMWx8wagNLz72Mk8/6RP54
VLxeNy0OsIZjGntf8e+M8jsFaXxySGb8GVUOSmI47EvQEWzMsZlQ4PO4cz5IvKSX
V1FsW1odQ3wee8N6lWxicEHRfBDA6hZOgS0d5e65eMPyUcdkIszRgRkPouMxsg2+
jehp7J9ZxERlCNVwb7qUmY9ReLAMtPVmZOJxxPpWfJfI6zlwKmeRsYUMGWiIsVqW
bq0cjZ/YZMr68L2lwocd+93kUJS+pQBehUZ/YHRtLXFO+KaM6UjIgHLZtoXkOByA
WEyEPUWHYSp3UjoEEjrWWHT1rw2cRde+xMZNcd0bdBMYtP8B0l0vy+jJ+ndEUPve
VwkvhxtEwDyzbT5rq0glEn9NNZcw+iSeU8aSgTHlbfUNnY3YE28rtY/h6o/SqG+u
qsDnn1MSm+qKuCDlNmxA5Q1Il8nxtLaNc53Q8xaVZJna5bJ3c3cVXPqmUGd+vbWr
fkcwpJu3BdQyyaGxE8UoFaiTFlDmvQY9ZYLXTC+RZtC5ADqU247D8ZxpoblR0asv
ZRV9qyZguD0FpN5LS+7pEXprL687adjPtjynO8jLJ8hdvqNd2enb/M62yBdS4wCs
Rkty+i6EHLFCgqpgkXxf3mb3YDp8B8fFqsjtfwRVAgmknHPzUSrgZR8zRumN70mf
AZiNz84Vq97sv+2GLKdLD/uPe32J01EYQt3HyCQ9F10lRsTMzQRLNOsme2WY34Co
JweHaygXQuuz0+9cYWZ+MxyGjyanASL1BFyz0FT8TfXEkKoLExTL9hN9H1/ovre2
1FbJy7C/dGdVXUD6kuNVStiy8hMguV3g8ZvM9S+eJT2oB+tcqRJb4Vu8EvXZMbkP
jdbfwFGIET9IpWCKCSI/N7E4JO25mg7VtnmYosq5wSgRBvmzlE2AVV/XBLPkHuz0
P/wc/KRfGN8N9Lujmz48JRZ5kHv6bcjAjceTdvL/jTCJBVDfrrkeo1r4+a1gPZeD
lutfNd9KdsohXxHuH9c35lXl6QFkRxraCF4j5vPS2VuC7dUqVuXHJXrmDssWT6WA
dlxjqSoUigFOai7ZPLVNLFTetRMGCLKtd+IxdwPTXJH672hDL3f6DJgdkdasJOnY
bWnhy4uz/fMWAPHu+vg90+QiqyhmIlEwxLdzmfoudnquwARXYjy2iV69GLuCgVrC
w3Q/x2PmLrY9Sb6DHEm6ZwdHNC19SRva2DvJdb+v11vKL0Q0lyQg6QzAgJbRCBeF
sBjWzajrOoUdpr6R2gMoxrrtaC0NGYddHs6gieirYOvkCc5t0v7mD5tMFF8dHM8p
maZqojHwctTwWZi1d0LasibDG6Pbc9TpWsKM2/WnF5WZVDZ1PaPy0dNzbqk7oP+C
SrZ+nw0ftSzJWFbd3BNQyMpvMpuaMKg8X0oZUCRct4h7JCFG7BP7dDPLH/gy/xI0
DTUaQXar+V6xXPCiUuMCTUFvgbs05NZ7lYTiDdU/5hbH9l2+j+H8x4Gv0tZ81NIC
CjbMWTwtSGx7AIsqW3F6X1lnOIZY12BhrjV5HRsL8WiK93HLRWG8z5GNhl/JiMnM
TKaeq6AN4SaFZrfPxCqE2B7lsgETTt+dfnb/cUjA1mwBCg5FtWxl86Wq9hKtQvcK
4CuhnslDYMeiyw3k+538oHuQVp2oGonFAwBYankya7R1rJvPx6u01vaMQjFOi1gy
VPoWYkNBIpu8VrU/hQgV/XQiNZ5g9R93W9lcIxKaUogv6FpDTb5hzE1RT788mATL
8Xu3cOD8wNiJpn6jB5NOVYU3AkrZLJDq1+58lu4mZCDxdyLxBHYFos+TrH0fvuoe
+amqlWJFA8IshThXAaXZ6BcrHGHSQErszdfzXHrLcdcpfBhP2KBJK3IU3YoCzbAU
Sh+8CXa6U6XfPZSyEFCjVDJJxPlH7suSG6NLXqOg24/f2mbx7f+VTAiEzu4VmxP0
A/8jFFrXdM5VAmK0Mpv+vW/ue7oBQA1ry+LqHxSnZnNvVNmss2/M1Q7vc3kb4Uhs
2hZ13zWX8iM7gdk7vW0HQ0YuVWyZzjrKIVQUn0UIyFN3WmCb+CmBS6On30rqHeGd
39ohj+tRQgekjLQmOPlPzQS1Ce0d7wQ4V/LYmY3azAR9H/Q6L6ud9/feZEfDsxTa
iOq8LqYlnDXwEULlofhDFIKsm9W+mI+2UtWiW6VAZ/Zt6A1X4jTjRnsHuAGoSxuf
UpJFLozK24um1VS1qpkzKZdpg1Eff+W3DmsPPd3YIb4Ceis683hs0VV/35BeTStq
BohITODgLpqgdacdCWVZhFITviHI6d045ZcIzNSRi372RG88vV1+AWBhF6aAFFGs
CPFRXDf6kBVQJKCsPf43vyG7lR80qJ+zkH5OXppEqrYh70TQPX1xBQrISXSXM6Jv
2VTp8jAgBHbc3hmhlswa2YDSq6N0GBZWqmsKZh1jDGEt+B93V7a1LD1c6/mMFokr
HwmziLTX5IyFZ4WZv8/lYsRKaG/9yD0WsT4X1VfFYoDwTlRICddcdU3qUPOJNV0z
mjdsLrK8ME6ebkV+m/M9Jux6eaPEMwUXjv+nhsmxjlj+47/JA2ag91KFirzW+gSm
uGlLDq1p4voORxRLeeUXDHZN3bOByNMmxMQicDaREsLvddbTnFOj4OZ0AkNQJUvR
DNUbRzdkjjjagI+7PmCheMjTwRfcBz54g6Rr/9HjOPVerDVQzvpqJpVcxW/ZRhAq
TTIYtkkqWvo6yvn7JI82k/iHP09or92mIyBuNWBQM4xqEZBvxsTCwaJv32aF/B76
Wyg8A/xocFlhLY3txqtKSv3AQY972t4yw0wmRKGLUuEGYue6RpDN3xbErjPbyGi8
IYPWkhZEifzeSl4GybfX4505pTZzZoY6B8Ou+Tczz1hUnjA8cHaoA5Hz9IjGe/Dp
4HSzre7oz5jZWRw+AH0gbWBv2nfIq0wL/R+PP9ZOff1TYSn/dFa/AN6exoeIpohv
YLaYAhmcB8MsBfX6UPIGsp3iEyBtB+rGcxD8HBQtq1oiz2ZCy7AjbwTXiUI7QsY/
AQ/o2SIR7s7tzEjphQaTsY6z95g2bV8S0yfB06iwrLdrrb4MnHtVG0Jr89bDeCgG
rZpI/z3MbhatdY2XOCGcrgmdke/zov8EVUfCzmZp7gMQw1aKy5HKyoMT2qKKFSy0
UPRX+7Qdnr+ULnVT10wPf9uSSaH8E9ohCPudsFOR8vGRvdKrugdhVqgbQViskXea
5+RLV9bAJ86IYfD7uGpZmyTXXXmEPFqRenUl0maJOSHGKsfxmOMfjn7fK04k293D
909OWp2tfHfTSqB3KFgnhIUGZ9gKPuy7nA++3BQJntacj19bfJtM6sw4ck9ZCNvt
XUZgJHmwkr7cFiD02joty2+CimcPEmmTphzmO17QbrHiN9BRE9OETVhQlfZSo3BP
8goBjSV69TmE1OxXvSNhJvz79iq9OVUr8aBGQdvXPYHYE4uIZWQwb2Xm2j5H2f33
pg4XbZ3PpV04pnm2lY/gz5zATfisRbMDPoOkMlAXksrRAg6IDg/GdG5C/BhSncV7
sTp7utfturnke5O/aEBSgp/B5sdZ3gK6ySPvHdAYvu+aEjmBBeJJdR5weeM2zbDD
gn+ulUo8vS9GrViMsOGA2ZCGiVOKsftUip6hSM9oLIh0XJsEGp7ygm9V4E9xLVLX
ANNHh6cfDwXQvYEblZskcWBX/TpTAbKuCH56+ew/EL3ydrGDnYDGTZrFgtw71FbQ
mrifQudyFZPJC8zRZvZfM6FT7xpectFLI9aVUxaPJGBZCQKtpeQ3M22/xS+BYn4r
oY94vQ53XtTcU+ahfdmSeU+HsEUSiCymoT0V+0e71BiE44QkezYreX8DnDaQJVse
MQXKTHfeB2DFDBY2nszONvGoBtazxZRsa8dbx85EtQgodUjt2rPva1Lk0KEqSL+n
aY9eQUag8rWxyzjYyWP5CCH4XcU3q+8psY/6+aQFqQCyQWo0r702PD8opzWVGtPj
h622Nj8RahAs3xCgw8F3Om2KwrG/mnLmboIKYxwHyj2TUYj4xRM+En8njc1tWVoz
IqziCagh4Y+LKI17WSqGwi0Ydf7iJfhY4c/jKbX/OnsJm6QJHm2h/U4iOI/gKqrc
7+WsFcMFoNpleV8tl875gqlc6UUUjUM0K9cH6X+uJ3BayT6WbY1M+IE8X2+KXzKM
JdiKP3pVVBOnvwNADWq5ruZTsjeJv56hl+o+GFxwH4EXvDReSTWtgjt2bRnhJ5au
AxTZkecLC2mcaT1rDqQV4WGbmyOEjYiKZPuHypOTjIrsScEl+571/l2D5xYIGhu4
ExQi24NQfp+He6dm14sXDAG1czDRKVb0Az9s/PCzDdDhmAtBV0w6pNgvjM2TIs9Z
Ip5pkwVo6rvN4EyAIRYDTjCeO1SlCMzzD2VeZ718C7Dz/cbfAgAaH/Vw/DbBqe+8
O45S6fRTotDpzzUMSDx+3T4FuG0NeDsn7MnHgivL2eWFaxZ65uEDZYnwyWKuuYQ/
DUDNxC/vvR6SUL9g2/tALrh4XH2LM3WuFwGGhriFJp261NNrKglCKa4qViNHsqYw
6u4+CkDaFhnoH0IPrSMuME1qZBTJXAb8YMNyC6zdk9hhgOzqQgAIN+G/FqFRsRUq
/Izf1cIT99eCboXw8tVttkK3R5vTsDzBGcHunYTzIHxnqJhvHXu+hJweqtVtolr8
5wkvemO9hrtSXAAPxbaS/6xJo+t7+k9aNZZTAJ59itKe6Gwa3WZZD4TaIfR86VwS
MHDM2RgqSyOw8jDxg3JPB4l/16pjsF0CtOtBzweilgfdqqD5MXogR1lggY/Nl7sP
YtE0HukxZ04C/pAAzmOmX7YJnZ812rjgekaob+Iu5KFc1V6yOe8A6l7qqC+trSEI
16cpUFh7jP+SY9PXqLOUs4M48tzYlgivlUPiB+97fufWffNTXFqHrGiKyzraFAM8
KMU4r7iuIcGmpr/lKypsGs+WFu0jCt0fgGq4LgqDMEGThGx75D7AfBw16XL1zRpI
ZWU+8BI7oDsQt6YR0b8Hs/Sz2iRgJHaPp0BfD5nIq8oy0OPi+Xga1RAeqGWSV0NT
pkhxYRJbSuxUS5wx21AQQ1WAYI4KUMjXcq0b9QyqC2vqdyZxKNqd7oyTAtWmsKly
0v8YGf2ivUXzEv3vLnXmxRYqboNR8PYVKc0Et2NSBkMLU3miMCRSpjsm4KePe4vl
6SJ3ilu3TVYqXkZZN0P/V05Z45+7LWkw0yB3BPSZ302iU3gqoVN7AvETMLSKKGWp
rhNpF36uDwlJdSymTXWg79eYLu5tZG7vRiZV6SkFq1itU/4fbyQ1WNXu6Q5dIIBP
RzKYTG7Ed0aOZHjXcGycRyTTzPQklikYNJadBdC1gEfMMH6PZoh5VwpPYrHLwkoS
9uDMb2bPLgqJ8oCJNu8x4rjsPJo+hnRaUs8i5K5XJK4U8qgG+shaAjVPmE3OZtjX
oXkOdNagQxrLvqYjS7HuoL+JqN01CSzs+7z1FQSTlyBzjU63k7l/9lB5PceWTn9p
CIrWCKExNj+JNnLsOvwutqbEv65NefOf9MqDiHLSxabl05Uep92gIT0B5LSImInW
DGTB/pnjNyKWOzyfwWbqW2vgiPihyG+Ni/OdKm+eFG1WOz5+Xq9yeWXavfzZ3yMb
MXc6fI9ovB4uBHb66CgCby6uZE9g5CiCechBMkuR1Tiu/NlhIMVJbYNSaCt0fH9T
trdEpDS7X8yOOQGzkCm5ePrJxICbbdoGkLWukldEnUdaCEAKQIuglTpk0DMPmZkW
W1mHzjPk47x3dG5yP0jwYVaY3eA/FzTx1VFA0TUgrPHXltEJXjQDWMr2aiXicEys
sFrgQW+73lAwlLuNw2rscRhn+yhz9IXbgZC2wjUTecPKN2SitG3x/dtO6Z/1RSDJ
jp2H6EHR1U+2nQtlM7gWHTqB/fLJ8/CrCZlTiElOcVHpdgQzsYS3xSHogsfUNP/a
GvmCmzY/HAp0cGUXPeevxZVc4zwOiWWN5uDpt7cBqtFnchWe4u9hOw6pmmLR+fgz
CpXcm6lqVVGK8QhQNUoEWgZcMjocRdswPz2EtV5+VCplDCRLyrKBWRVCJBwzq7ut
4geh7M0MV/Uxq2cZXlgLMKBRJvj9RIHBWhX6h/QaB+9HPx3+hotWNP2ZtRB1/ZOE
Q2PKUckXDaahpD1lkAcrTO1x8MRN6RoNTLSh7VAx6+iyVKEwuI5rzppQg/K6bsAT
34vQ+QGjUCxLb7D/lYtjPyKk1x1vO/dKQ022vzV6arDSdUyxusbC3W6KC2cDGDIA
0ebnnYbqNvvqAs0+8jF8KebzqUAB6s0x3nNwxMRKWvH8Amc76l6QHqDIWCrVXVaj
VqmKFEFPLwlhS5wBw2TyPAawX1Z5anUmiSrEuwu3T3p3y07HFMmNe/1m4tx8LFhJ
243I/S7aFXylsEJtTuG5jssDBLPqdJ7PiNMJ+IYfytJVdVEr3L8LT6wy3GI5VpTE
PmgIk/hNc3wI/CFKJ8NDefnGrhNEw7VAufu0fpmHOZTmmG9jaXm2HyKbzdmQi9bb
neZOqjbShe8u5j6qLSLCCrEqcOQgAjiTx0P4SlRl1SHYZl+ciPGSgsBALEO/JIC1
pXKsiHG/P7scIyPf4qW2p6vPbGKu9+mnn4tHTT9GSbQAKNNAZbI7E+upGzw+nign
k+LXsWQLdk3ySCz/F4xAStvd6Ib+qWsI6ii+u/b1vkFHLW5o7246ppd9bmkuQqNu
FQ56yMcoYKlay9Z7IZoPHy26cnPIev/YLrwteAdAeyyS60y+T1O5Hg46FJZwzR9Y
M+p5WGLgT7eaoQe4fmlA7SZ+9YT1N9r795cg9B37YsnQkGwA+wlhVH5GVH8ttd+h
TNcoz0hlBawngd8T2dhXZtNUGH8FTFkWMFjbDAXySRV5nD1Lw9jMR5ylbJrA6nrp
W3xMUub2mkGgZlLgvCqNqzI+h7UO/VYb7mArUPch/B+2Ji3QpEIf28CDmR856V4T
CrAhWezl1lyFT0+xMIRYO+BwHeYnParNB+5abb36l8J4y2JiUWIlCcrWqil0jOVn
T4vuvHq7pdtORHvHyHZydh/vQ0/puFUwwrqn1ay10pXWn/XjziUq1CXSDeu9POlY
lE7FyCfdn/Fo/3HhK9xcxQZft/rICmjpv2r7SnaBerCzv1gjNMkPodCrZ+L0z4bt
TN0MhA45r4j8fbgR7S66yCxoy8dVNBFB19a+6dCnwupXKaeHLuHz4Dx91O1BZwEC
v+JAAqvOC5I6eLN1ssC/Jq+0V4Qfuy2aRJ2VHWShnPea7zGO2dRE249I5cpmQeGe
p2F33FT8UxIl/SpG5w5o1Bc3MFCZ6OEDxvrSvYQUQPAwbrK1+76cacPGsvVhJ0iE
95S+mm8xYmUn8zbVYM7adpO9g6VE0Uf7zSuc7hc6JAI0QbD6xz5waKF2QT1PRnyr
9cHCYDKop4iPGIytuWp6bK33K0a/RFCPVPba/lzYARjrOxS6FMq/SmfLjrTKjp78
e8jBt1ynFUEgCF3+2X6MI2ZcH03jYEQ4y3gJFUPPXjvJoI7GSctMRJPf0VTosILw
bhcVbQfCDPpg8w9LNOG6WE7C1zbp5Vh0Iek8bWD3p2vAlBWjy4Uv44C8kPJFMKEL
CQeGDy2U++Q7vBLl+hDncBIjl1pwcTdw+SB4A++U1c49t55cC7HqGnQE2hARu6AO
+VpHzo+T95zmjRBcBE8gfFmK6f9qZq68nYPnHoO1XhvHiy81zLBoCu5rfk/MC3vP
XU9umfceSbv3VPay5QAvzq1YD4Upb9T1ov2NfKPgzuuO3V1i17gs0g9udnAMAjow
/XiRKF8k/yqZV7ueviFlLs1MhtITlMPwoRkMWDkkq1lXlk0rZxquwfX6hTKNb9L8
CcLH7Rq8LaR9Nd3ZhwRzk5E/d5TI0q0lBnmSAwNcvyIFfo2L+KwQwpYhSYcSnUyE
CNQLbrbl1MWPfMIssh4hgmCzElmR+smxpuKcfndFHlSrkvP50Oi3gkVLZ01kiF9C
r99ZOs4I2qbpydPRkvL+lb1lKaLv0twnLcPZI8fS+fc6ip5w38pc3iYusn17BDKv
lzaStsk/B2IRw3aKDfFXZcYkmwjhdWuKyB1cfHayTR9jn+JI/ItNsdRHJcfQeu7V
OCk3hGbfF0SGYl0e4Gz/1TXWOhBB028e+BnTZBNZ0L+XexZSSvuKOIx8UC6F2g2/
e3GB3ojKpb+VaaRF4bxQtkaYb52hbVHs3ts3zKnRBjF4HIL+PpWwy3HuWydqPCHd
rxssFHTSXNJ3FpVE5uLM2umked8FzUTMxoF2wd8e3eSq9c5wMKGumcwLLfkN/HQM
B7NsENr6IlUq/vtO8k12mi7dwjs/Z25AsXCAs0r2eOJgVEYxW/bIYRM4GnZ4xNNK
dvUUvfQuLU7ibYc2kDVY5vczRbDpCLwDXY8fgN8lad1Ob+rUi98gx17Sqt1dk+Xy
h0io2RO00fPQqaOBZO21qPav6nsX54Aa2Pbyvx5x7EFXCNkmO+PIC0fMk9m/4wQ2
fssjmQxOm8san2eDeFqqoPMPKk2msDjW+rvRcnWnfYajTzd4FdhcwCYBgyRi1PhR
+4p5GZOhbYfL9qpVbvWb9mMiGk9k9tgCIsVZ9e/IOeR09sNRF+voirlR5nGQoXDL
MBKKN+LXMWAeA7SNK0LfQDLASVvgVRXspfdoDugoHCIt5yS5g+I5TqPs+F7wPdpj
QKAY56jgsZXE7lpmQQ1O4flL6ptvMmcRc3ckum0aRjwOghNxX59a5LRsjPfQ98j/
PcNpVRtVQ5EOky+ndoo5H/s2VkG1xnrgApLLY85hPGpAHJWRjJzm3MnE1k8tiCvL
VHLBxv9ZOi56fDt17Lxr0A46+F/jAet7388wUYIEZncuKXYW5vqdKVVe5aB0LS7f
+4qukkFQ/DacwxJLWxTHRR2PXJ7htcNE8jm0SU3a37mc5dmLljvnqzy4o2+WHtHv
T42sWqFM0IrSm9DR/dmyqDqUhLTcoGVPsotzynUIn7q9nzKve5H/3sMPxhgo9uwQ
sCiBQI917QXsNQalaNNpGF8AsX2zbnVzPq73Ys5JbZkLWo3cnsB8/vi/b2KSYWwq
qmbmvwCRUZdPdYlWigb4ZgoYlM1gwwO4vuYhDDcA3t7GkQl0zedjeMSOI+PvMXAR
i78P7dqpVQqqbtnJMWKJMOy22vmqNxsntwNiAZHpTkYGQfVyMCc1uqcbjaFL6Kh9
oGH874JorkCE4RxYuW/jKedm8UgyFT4RLRVshthM71ak5USS2hQFDLown3EJTAan
XrMMxGyp34WDsfQRTYCgWjmQUdxbXdRd4Y6CWiU2W69mUj4pwC9vmYBICuRP0+xO
HYEnSeL0MSYQSl1h5SgIeEd/wg6+xBNjDBnZjKuLhLHoBP/gyaXogepivwi5GRDv
0Grq9GdFOR0MRhhA2phvsKtRg2G73sBZDkaWHvSACm499ndQwGhyv/QVEIqwYAck
t+NuLka7+mU33kTGUuxEMbOhAigyEeaXVEkFgxXcCW7EJWCuoQsIZLDZPBDqizKg
i1CevaBZqPMZvOZrUexyGg3D33Pdw9ygtrgpk+VTZ+44muUXNgPGp+vz8+hZqyPC
F64fC8orPLeZ+aY2vsJPvddQdLOUjhh2zxOUndzluImZn96+qhrXmotFcZwtqi5F
Y11s4yh6dVZzlRxiN3HCiYRSjQBeWcf5nbb7WprFfvY9nyeCnT9sw6zC+oU7Gi84
dQjxT+L0xv/Ll0Z0G+lHekb6TKFV7ome9t+rHvNpOavsB8ZTlNBlZe/FkL99MZNJ
3w+xIPaevJQ0RtA0ksAA85z3QifQ1MmuZqljSuWTVPTMsmSTmIlZ1K6wsqdTSp1Y
wUpjVxtfJmM+/D9ciXch4DQkz8tHsBUdgxg92Ehnj3pxKCBNMrm9Vg5bTiBuF3LD
eq+yEhesO9mgoNZL3AZbQ0H8T8jD+zwt/LHCMHecZPXDOk95ulpI4hw3NasuGCsI
H1lIp/IW5x4EkmmbWW5VMPe+G7ZwEBC3ekDtaFYGQwql416lBpqfhPPLUEwUtOro
ZlHtxgbfdVss1OrlDHdi633a6PMLsZ+OPWxWqF9iM0najbk4MOK6hBe8xWVx4uID
NK3jMRngMsVQbKBsWaee8M7cuUwyMT5oTvHL92RsmpImElxNP24jolKYAhhptr4u
V3n9CoRmXS0W54aWjHJUB821WLFXso1yYuhjalAaHSXBIb23Ac1w4TNpym6SYtr0
540MuyZA0U8Kbdwh7xgFflKRlJdAKQFPqULrgdwuzYMf5W0PVtv97dWTtNpYavkR
X/65SIty57mQDo+v9E/qsRWlMeHY6/zFQdGhMsOHE5rkKc5rvp+7hg2uU3QhVqeJ
Kn9ABQPI9N59L65/UNTvidIY3n5BXUgJCKtCqqcjyRUT8iJB1emZkNrES8pvo/CP
vrnZmiwMLNJfx4R9StqPqcqHNckuXraYpnSB9X+Q4b181HURisMz0W4oB7N7aRqh
pCRq5I1F0qhr+sM/Ez0bPpR2kAE7c1Y+bz8bPxMv4RevDPSOtCh0gFFuYrr4jFW2
pGQByidv+Y1yNw/g7iTeC/Vp9+t0qTUmw1vsH4T5Fi79y07b83RHpUWXCjngMZn8
EOZx6dBTrkn55r/MB0AcdPuRGiRsGDXlHbNG1eLE02BvjAwpEvrjEaG7EfASizQS
yDhyfyykcL8XPcu38yBxyeTdI5Ss9JnJM0xJxJrBIU4WnQnhbracHaWqumzL5n/E
Gpqro/ewpRHV8n7XhKltYL1+2MRR5KFgQ60R2jUMhugGYRy0gaQuaNn7muvEj4Fk
qHf1Yp+VJuYPva0cAmslb522lmWcLCXWSynYAJojFF3V3OG9gy7uvLF3ID/D328i
hXjKappEitvLfsCvzYlIeUjpeuLEgYkzutD7zQgGQjLpqzymTAia0Y1heK+OYj3O
Qapnx1LSYkXJbA01kxJc6D5U7Plp8ELpPS5XiQnWmRmXtI3/rnTlnBdXoKJFME2M
o8Lh88lLJLul5iTVnKK8fMx6AKmsHztiWG4lCNoL1ozWUtaiTfzI0Y1bN1pt9/7A
LWyabaVFiSXsMkqL5Kra4mNXTwFvL0v1DQ3cFBAOGigM9i3BSZg2w22NHQwTkcsA
vlco2ZfO6kgffHj5Eim/SuywMtpFNZ3epwOXkgXT72t9q7mF+SktO5NDWUSwnZta
SYEEeX4TSJZEnhrXkOK2QziQ2e2nWiHVjKqZAuDNA4y/75rqZ0Tr7ZDb3COvPG9f
j17qKvrYbX0Zp28Jj8Il4shZSIHYuxNqhIyQq3FLFwx5lmQ74M5/SWmQtnp6ZUmi
Zz2uk4F/RlJjEMch5rGGI/syZcBrOVAk3vr3uOd3MMGnnQjpgg1WLSEOoJwtFcUF
wqekfYwSqig4DEF255ZeCok/Ide3Dmh6z3tadS9xlp9zGm+WsJsPcFqbejLuOWzo
05IJXwE4hXiCbQmAA0YTszoK84Vt0ocjOYJvpzI24JCx/KBw8MAeMMYM6whNZnni
VIhOQCLYGiS5NaT9BKNN1b3eHa71UgvbUsU4hCXCSi9BCLmTmxCgWCHDX/P9g89n
OMCTGcZvMXrv/+5SoBXDFFAszsnN165t1+TUYKa6z8fueVgwy9n2r0krBDifLaWg
14OJDB/ruDsmG5TUNz51hcHVz7ZPAr0lesrhBL301k2UzcaGVHNcXE+ztTRwvYQ8
ED3XQVcKh08PhOPQgPGY1Bai3Ggxsbo6MVYuuuEWr5MmPwr9vJlIKv5QMvDCfRHO
LwBiHWC/+qYwu5SfsYfzSw8NddRGdCfngRoSZctXUUVYHbtTyq2P1JlcFnU8QY1U
b4h1og74sDWQ+slRNeLQ21p9uu1D4OWTecz+cWts2z+RCP1PFUlYmUQ+VP+aVdt/
0D1pAsY7RA1/XhTXFSnuB07VDyly5N/kUC/fYC/f0FUpOxIzOPgS7O1Mmi1vjUAt
U6v2znvuASDxXBS6ppbDl2rgF5r1N0vh43TUC2JaasnZ/Mk9BrcEP2ZfxoPFMZjk
MIKF0a3BSYTf9qZxwj9dKrJXp4+FpDDPhvqaFOXzgJTVQLX9xWQitYWYwD5AiZ9S
0U5MN6SJXIOLWXmwsRi0zfrjtMeidR8+EnQnCJExKchddx8hyd9fSdnKJxZ6YJWz
eOvmVzMZhQ7Z7TqzsdhF2WCwuqv/FbPUVXjuzJaNCUn65PQolIQXVynnMx+IXB4h
lT3ReuIHn2eStyous0DdPX9Ia/GD1qEaRjm4Mg3Sl2hFBEvIvTKH2jRZV3j+Ic5f
q+DGs4muuPoYaOFtUDzFNzQxzoFgEujiOcnuhF5MdthED9yHrJeZZBqkacdrklnX
7TLh3H+NGw4T1cemgdryQWh8v8uJkam4vAKBUjf2sQk2w/V7IW0YzeE7BFerarvo
bQClNSRWSalsEkcE22ErqUcyLfKMLwCEB89dQ53T2GNr1Hbup2ZswMK2Dk3ALMmS
95mzEfUSgTif8Z3BVxTJ9unmb2y2M0HfdHlCJmAaNcBq8wmd4bdUDIBBPrOc/hjW
1QVkEe8M/i3Fu+c3U+jlQHrgMkiy061BPhH0xKBxhIm7FXcquNeR8ghCDNbmA1Zv
b5bWNg/lrSPDWBaGr8W3NMI8yWcPiWCwEzJMw11s0RNiltRlw2hOatPl34gqFz22
ARHtSzlGi5/Qgj94H0CgtrAS7KFDsh+3pgHWmPxVvuWDxuG1D7mLzq1EWtiz3M/8
m6/STx06t6lJro7tu+RYlZ0y/XQAuRLD81ZNtpFYIjoqkRJ037i8KCdAs+V/Jo4q
IewUM4syTNol7oo50OLc8yyRpR2Z6OXzoOWajv6qixRS50FbB2zbV5TkC04wxT5/
5NrZ4U27wUikpZmlBgAvgBz3y8JH1B1bf/WyQ4ibDUS3j3tU6BU6KqVH17gpfvY5
QHKQAdX7h13jqDIEW6U8jw539YVbcz7X+76ogFIHi626PCNVaVTla2KUl7cV12BW
s6EDxrVaJyvTMRhtZqRClaDyCuCHpIGITQQ4hxHPYgCUa6bk3sKDAkczoifSR55M
WwUQ4pizv12zlPzWrgcWzC2ebNGT/raK2nJyrRJLCmGBCtB7yAfeqAa3tpCb7Awq
YvopDU+jZTWH5jIik/DDxe1rVfwUZZjGPLfKc5mB/1o5aK8BmbrqipREztZK3SR/
p6lMkfPfruV8vzYXTk4O6OrknzqRfj3OXDV8jS0JMjwPw4cRTZRIo7E4hl/IUHgp
BkGUB+zAXgBiF4LWkjI5XlGEe22qtJ1wa2xCMFl+MLmtdKY1LmV5wIci8GAn9zNE
C85s3CtJ6RVlyc+PM4Eu4n7pmK06xM90QFQtIoGjmqN8ELK0nQQZRNdv2WhAaU+5
c83/jn8trC3hZ9Wip1BimnLpF+pdhEHam3ZLXqDLP9Bu8Uy5745JZb7DmaWcIG21
x38M975MufWGTBprvHgacGGRMJnAbcFt9MLlAqd+WxZML0bOGIk2V6KUU/Hi4BQ/
4hqrBysfwsXCZdxZU349bXjy5VjsWuoj3kLj4imoSShgDORHPPSWvKFwonIE1m/r
XH1Lk4ti60ynK6/A6OREy64/YqLhy86XDHvSEIBhPY1+jqTPq69l6uHL8N9VAicp
kZ72qIGIYX4UsSrwe61tpF1CVhckG4RBfcugCA0L4Y6fxRqr6c/eZ3Qy1zGx91n9
GstrtP468JPTW34JLr/H2+0i5IGqQPsbSo/540lOBoptKco0h2DpZILKmO9M2Rlp
PwSI8iYyyZ02trdeoEkSdTe8S/d1AZqcilXA5J32IvQBa8rh1dkg0J8SKHW7EgDR
hAK3JRPMri/KxNnxO/gccZoIR0u6SfCRKryXMDegmdZLGuUfeyFmesA2mR50Ed2N
YBgZtEXW7TtK9yaxy8U7+GvX8FXGpkAqq63Jx1meEfv8Kr77rLW6CFMf1+iDY/PC
ULPrYsFHeYZ6gGSR8bHb0RZv3IjzTwfoSfpPHDJXlctoq4N+ss7cYtWzuKh3bkqP
wnwrDyARXoUd4wXdMTKsLPeqvmN7R0e0uNJlKiMMx1QELqsyA6Zow4b8qdWhZfU6
JZPq7PCB8dtfoU0s3NUIRAaCoz3GPzlUhOACNgL3wzB4LtLnswjHg3C1iTobXxab
iLDhWCvuOQkDxHHBwEID9EM0musKMbrWSwsmYvEOtiLugjNUwFBYlJTkKmy2DQk8
XIhU/PBYuNbRqlOXHaQcasrwevAoCLUqQf4nisD+2UoXSG4TtLYj4e1NLTvCic41
UvU9wn7u9hr3HpHCvpI+uyAQRcLPglHGSLn7YuZbDQZ5QMVz/wbnrZF4KwvJLKdQ
Ugdb195rzBpYcnEMHJXm1t4v/xIvNxxxgfrRh8tkcWJG0ckl6WJI9qzl37ehvswD
wEqdyuLZyKX+korfU4Isd89kfB5+bKo35bYb9H2uB5o+PiAhb2JK0WD5/mv9K93I
QU0bqmODX1RYpoe47Z6MS2DAvG701bc5x3jvW/H/THzOSK/1pp2rN7WyVgsg7Ith
FmttG3abYvlT8/v4rioN02SUqaDCkUseGbKqZdJhBHoz6DxQmRHVOgIPP4RwRuOM
L/ffFaDTVcxAD/GRr3rLNFg5/1p64hYTv/xtMx+wk5UIxj5IxrcPsu4e/29ILm2H
BBlNEP55tZb1Y7dkBm7+hm52VPuGacAS6/Gj6dY1qdCZwBVIGzxk37byHqzrBMPe
ZINvRzY4maVIY8QdThrT7XDVVcgxqCw8puzt5j43wBORimav6pccf8msCeizWKV5
UQPuIfaWCSk3BoUt3EqGdttlIefmaGcp3F1nhcbmLIM1PS0qwuv29ZBXkOryiut0
s/Cm69ru0xjnitd0ZQyIK5gtcyI37EENMUOvffqzZ6LtOmckSSCVoOgTtSvfFfB0
urCw5J2ghUMfY5y+8k/MvHD1KzpQoQ+cfjemfeiSGiyHjZelek+k2KsYNiJRGjs4
DSa/MXNWLXfUuKC5/UoRc/AReHiDQbNx18hB4VMaiMubDarOo4/IuTEwHB7MeSHU
AGq7x0rbDtfTKOuhwEv9aN9gwcKI8biJQK9PXvxM/e+yNVeliq9nZsDYSLmLLsiX
ynLi/WNI+/Hv9R9IHRwPXS8TLVgK1ak/nuJlHw6R+0VweMbdVQPkPF632ZxwSsYc
KYsm2CxiSChWQUx54q5SnUl8Z0LLxvalhTW5mtShgQnKDostPcTlMOJlwUiO0MYo
NEM89xhaIoGBAEVdnBrHBhQOmTLEp3H/vY2qPDDKx133uuLJPSiIYLcY+zuVyLAq
6CGcVomGD66vXhTweMQTSzVq9rbUrJFpxMtaJKbfn4Ksv0bm6F7Z9vlbFsjdhWka
V4Q8z/j51gk9LtKlUSEPzrHntOuifFon5d+/JuK/E/K1JwK4ZycNfNVV1pHOilaB
r3tVuOYCYGmPHjhhK4TzCQSwbvS8F/SeEiWmydrdpvmKFy7V4isCIUw84sbxLdsg
BTBx0Up2Bg78KE+tWP/VOgfAp8sATo2aTt8MmDjqr84f/K4Eq55bCzVx9xQecEcK
UmkcwsiB+Ij+53blWzPDX1mA3eq9YEMECmQ4CguSHYFvt9sVWZdMC6mlHNquzumf
5k9nWe+qxU1zc+UDfR4Pl0fxOUyGyA7SEyfoLNKZJOQTNeS8ZfXeGxubu02qnuu6
Qrt0LldA9L20K7+lBsQSL1qKCzIDm9HlTXAabqBpbk1Nn13j7ykd7hLNnX7c+uoI
xpg/lcyHGZVWBVoVbQXocF23GNTMrrcfqBozNiF8aemhVYCaaUWb0nmuTygy9CJ5
ON/3OqI2I9FmzPyo3syWYLco7AxZG6Qz3HlO+BPcAztm0xTVb72AE3+fLcza25ws
eVW3p/f5ZNY7KQ7th77jvr4fQHtR223Yl0yiNMq067dV4OtMGSl7PJ/96VdSCSDk
3O/cGF4xAfA1UpGhGzHQ01PAC7IYcfy41kRprFZql1pEp/5dGJj+I/XtN6I3UMNB
I/rdMJhBkmHZnC74ZdZaEVHftz+4rCVk59bVGw8HdLRd2EVI9AUgEuwe8U7LfV0v
4qs0aOd5tl4MThn5SowjXVVxU4b/o6g/46OSF7s50g/wsdaEoHBuEBZu/7j7k5vG
CerXSF2j8mLEfWhJnGcuuSbcl8VTMRHIM9Nn5b2NF87rRghNbHqOVBb3HEz8ZIpw
dCph09/HJWebRlZI3pFwZ4pv3/2IbOpGoDqvIqYarl4vUy9f5NMk9W1YZFw4M5v6
czINZYZinrwA94NLsw0xzjr/EVDDqkuXwmvAEjFb+p8afNqFji82xToOMjBRrPWl
nIKkZj1+lhRaGOcNyvj+VYd19wZFLVFNl9r3eNmqvafscuQZHn5BnRdTgOsUMiyy
ZfNIDa6EqgXrK6r4/qwnkNqnSvOZlEcd6lBtMLTfFNiNDAKY8sEYIT04hswLW0Z1
XlGjNER9N28j3Jng4kNE70QAE+utSMUAFSLUVUTZHis6fiJDDj2E19F5EszT7New
a1Vh/n60pVmZrH3e7F/y5DsbBjOyOLgD5L/Uy6JS05A/EJG2bMx+eaVn2QoUTJ7k
BxWIp7pY2L7ZufQk8hzFhBZH0bPfNLbsu+Xj1/5wbAb07pQKlf9q5GRbWitTq4/N
7coKNMnHDrqm/FAjF0oyNHtJk5ZxpV6VC9F1y7n/XmWQ0yHUYVsH7dfYacQjVnPR
sGdUO5i6qLMqfTlFEsFKI9N4z8PHqonydgSSR8usaj2explDxcS2U7WMHYJmj0YM
8Q4+lVBqyIsg55mBLeH3NWtzsbdFckRcb/8PYanwxZfh4nNfrRRFi/lXrQ8RIKUt
RoAenFsAq46XmpnkHTZMfafjh1v/Rf3SAeyMBd5+freFHJf3nJVQ5/db2y7Ot1Sz
yxo6SB8J3bqHPTeFyL2IRvVxx6UzYUQXFyj29s3Xr5J73DnB1LslF4mjzBbkI7Oi
Ue2vOg2HMeDn286GWb/K6l8UdqDp8BtkcOdpeh9gL3l0GDdZWpBi+ZNwOgLDdo+r
36FQSVjfjknRCG1URidS/IzHMfGXxBd6F8XHVtc/lZEqDtMncHLJo/t4JzWDjkri
ZEy3yhV6ZhyjMWqn4ZqPkLsEUFRKRFpo4A4PG5zn+8uBGY8cmpoJm9osjqw++w7i
v2LuUW+krL0XvebYCTMlosG6Wzfj21TsB6UjKWGy8Lr6pqzDAJQkxPR0vh35DgGW
O5SLZxga2te6Qmv/6CnGu2Gy+lv4ufXfOLEjZrveru9+U7sqUii2s5WKn1XllqqL
hePQsA5EkfVwGy9g4DZCzGgmvr/SpAfeKY8GlmvXKMFbxnflF88DFm3XE/Fh78kD
SqkpUP+Nsct8AfWkPCRF7JedAATkvCn54KAH8PPH02tybAtKFZyMTt91jqX1c3M8
1GWzioM5/CWyEjURroh14N5hMnlw7a/8/YmESTQFiF5JFLx3CZ4tU56ISf0GMcc5
tMJk2828blD3O8zkjkwdOtVQ3Yu5FJPH7NzxeUaJGuv+AgsOWZ1+x+gY7dOEtZsY
YR1H5zj6PI8Ft/q+BxqhwnHsopk5FU/aA0mblSNEAt8R9ys/6ostR8s2KBMVjYAb
gy/Fy/P7WO2FlZEDtVf5QgZCR03H12bOlFPimca5ng6effIezUcIR60CIl9KWsyz
Pkoba/WIrEOttvVpUC6nq2+sMfk21cYvkYKF4TNi9pJb/JvckaogDnRKo+q8t25k
hwES13CdM5S0oLf+itFdYLYJJok/0btsZPLc+DXTTrUY4CPSbmswBS0LdmdygJfl
77zvD0a0qKDwNsktIlKu0lbXaa79i3z2nHcerPynj50bZChq4gCDulTXoUl3QOgr
lLa2TqSEYPzilztTiRWemjaeH2hKD4YausvtN7ioi8wU/PF/LZT8PSJomgwgU3EQ
1pFsbk0nF7Ra3k8uFMmxhKbLfglP4hP6hmgLDlCaorjwA8XCP9kvbRusXt1STyra
gqQVt0jTNHGqZVAAHyZ4R9ZaoZHxloDfSh736CRcDlDWE5gjVaRpPIEdnIEGrZJA
LDT7wt+/EBOv6fTNh7tr2yHtJitvQEAZdKXGCakiiByV7PR4tkmmmN+rHp7lH6t1
ZdLmO98a9tEDOQSWSqS1KRAoEm+ArpAiFF3xR24smYdHNsVIb/XDUSFCFwyFsH53
FI9GoA9/wJdZlEife+fNyxAVx3X5J4N3aZHJTCS/jkYApB5rLm9GbZbir1clVOwy
WML28EAHSvtvwjQYemkzNs4i0aK4+DNu4NnNWJmZz9ar+v1p7HZk+Lk897sAwDV8
3y8mM8dan4PnOl7yl5PLhXSbVlLhWMazGvfelnVGqqkiXccP7RbdJiF/SCMAsBd3
RhY7FlPbfjjulxUUfDvpZ9zCWwVLnuM1HdzK+5iLr1JSbygQqnmvlR6DZZ/4GfOz
//SAg1flUGfizMiNzv9h1xfZuUiDUPzwulw4CiChDimu2TM1oMUeExYII/eaWM6N
ZNn8Dg0S1gbUm4leERDiCNq1YOm6Nw6V34AoXn3KZarpMTreBPAWXcTNV1UExImW
sOc3sa7ZtDRSErShmcnWuliYhuRizsVfEmguJUxEx6fZUdZkC6l1/AnDG5XNCkxf
oZkCUvX+j8Gn8bCNz7i5D9HdUtcOIuS+hCMnMS1P4HQYwQNi9HkAgacijd1Z2uES
ce/ZqYOMzGnu7ILGNUbkIeIK5xIdLrv+TEGECjuraI2cySnhSUJL6GQ4ekRSujys
yI1uh3uggLeKxW9IdwGimnlbF+YLM56wrYnPfSj/RzZYGoOjgDGNKY2kpjOFp9A8
L2XAX8LzMFU5bG0SHjWSOKcjz5G2vbKoZ8sYptJ4gb8vtApunRmXRRlf+3g2VzzM
QeA6FAb9qfHFDh0UcvnStzZ7WDyxbiIT9LnNETG2uVePr9ByQK0diQLyOklflQ0J
fzvh4Ui3sQi69tSFkxa5N6oRAGoknI6jq5X8SOFjFyHYSC9FNY5L/DK6/okqbiv4
Bwo2CJgrkZFdeU6n0YNDnVLlU+RnMXIsoMrQslUTbtLW/MxEjyq7eDANELEvK3wO
xuzA4G18EeWJSBuu69fT5f3k1s/PPvwpdw6ZMFgNkw4kkibOroYcIjBdQweCK892
E17lLJwipZwNuugyunfWpqFjO4OzMLqJqZZiHLMv/VDrajz79oOHAmiwy6XqtKk2
fyMU7/RQlncdw/Y5bCI1CVKnAS/UybGJ5EJTIBsKu+D6Z3cu8wBbZTNsUlRRT38d
asTovvJDupoXYleioiVxfs943zohK3hKXvDcHBNTqY1lYIshDAc9C2hB/ToT3VVW
jnj6nBbeRIUuQ61c9bu/K51kJRMUTa/ZcN/5WQfdOti6jxcKMt93vMn86PDLNFCO
KMYVAQnf6L4CGMxnrp7kn4JsC17LRHDOFHtUXINqSGp7GTWVKmq3mySExR857MLD
7gl6ungNt3T7xpfnAsAIQKO10Y+r4WfchITFMl6IDbi1vje3oKrSmD60zTF0+9+1
meL0uLvwdIL6sm4/IxvRuPVR1UBVaQ0Ccll5Mx1vcgWsvExKbpXVdU+ua5MtbMXd
DESed/0y5ZBb9lBaUdcO9Xy36MjxEEuX29xxRBlX8f3EN0Ps5FYy2KxiL9unKcOR
XLKsCEUVZd/69EJ8zFCBpIrPAOlES83meWkUp6WjHV8jTz44nR5NnRugWHwuBL5J
FmSQG5087U3/YB/snd00hLc+D8GCzgmq6CQbNFGRu6JBP8VMpaVswjXBjMzT6lQz
6fKaeRnxrHpUklZ+zYoiCDNzl0A8/a+Ho8aUtMgk8faqhDiYFgjdn/hZf66U+PXd
J5+sWj6BnykSuDETXF/An3wpxDX8eNw8XJWh5pWtZ/aDc4hBPORhQ/em80vR+bHi
FtVjUgrfgknPwb4QgCgzS8SRErX7NGRhcJBgAgthhgmmqu1R7micJoMAC3e3aokr
2pHPROg3jYvG4NTCpTLjfNNjcVeZfMBKCyvBeaPpRfB10mbLF8+S51A/wniepLWb
vsDDt5YXlnf300QDbbyxM28ZlCdWjd7sI8fO///T7j/8rESp8HOSJr+2dodqtAAr
1jhosoZOQdgtc0m4s75cF4c85Rw6STNhQylPY9xQt/4lu9yBZiAQSK0jX71NuqiL
gpS1lS4O7OF17603lJuJ2uPcPhVjfpws6QHwbQE3Z/jzTvu1PplrKQYlXNw7g9BW
Iegk+rJnJ8boURQ3tHS9OLXrkzjAfVAKIh4DHrOvJt0mmhwYwB8fDndklFPOWHZ0
DdhQm0L831gQZzhbANlnsKTqurQHZMMRiTpcWj/l+nViZGRhnLLRX4yoQnWAL3Gv
kncyQzlQPRJ04qh9YZAX2cXeam4VRNRzhO8hSIjF/WkuS+VZABnX5GSTvmiC7d+t
RRgd7MI4Ve0Zoa9uDxnTqUMrYXj2MRCXMjhERjzPQ2dwfxrdeJybGSDI34gxXNgc
LgcjKJphbSwZHD374vGrHEzj9nAMR90sR7G7KEvN1DVtvVIFO28LoBDZKRC4m9Gz
XXEDrnVRzWWONQ4EYONe8kGeQmfzWM0XP82+7Os8f5FzhrGmAx+vRQV+/08F0knm
k8SW7qydZm169fhrRJJkuzz8TVBLWKb9iAh3WG2gULiV+s4LHci3ngqi7nLQYYOg
jXlDOFhHk6XK+m8bD8VLvGH716/NllYCun2qd+UijyY24GPZNI/hDqOLfIS/0WEf
u7upEFArjXNqRfFgsmlV2jGqbt6Z2JQdOIjv79x4cyfJAp3sz0Xh4VAHYuDyVfGP
m1rLaoA0dFMbY7xXj8FMDTmm9U+6BI3euxhX25xPngfCu/pFxaiL00yVq6E1bv/u
5OM5/OJLfC8wzVZKwIWNdfCrFZzLXWLgNm5gzW6a/q1nwl7ezKIoRPbfp4irgl/t
DBnFkAFtwcZE6x/p4YikqnhvCSrqSV2+UyUMcknNOqyX8akhq9Sx02RRd3LMqLWx
wdl2FClRCvjvCsGGQfOAkK8vGLNd3NrQ8iB9s+sn3SbUd4mIwxJITAnuHIVFqKo+
4WyTpfcaMp2UVmfsNja88D2otsey2KwOOaFnAgbWcrXwO5xs7YokpU4DaG0TZegZ
6NqZzFvcbD4Uah6YSsuZj+YpXj2wGVXmPpITqInL/5nAPXEayoX7RKyiy+9WvgtG
U9OFaFM32Q3aZu4wqkudmou4jhmoWL9rka8P5tq+BLB6nl1jqzTE8cKbK2tmkxNH
k2zJgyeMJb9/TrRW+cj6yHQoTAoccX4/WdaxrlERSKRPcz30if4l70s2gxYVDNlz
FwXiP9O+lUbOmnyhmWWQvWqPytm5A0ofwsO69uWx4n1bZ3iBVIvDLSggBt+JA81h
3m1OzDnGP3I+oHAPWb138UhCZ0LcbbfHg4N4VMgEl0NxUN4rbccNwzhg02vQrU+H
Njt0eWxo41XBn8EquBh3D9HZ9XrCDl/sn3KMpWVlikpEAv8E8M+7VeCloxsUFwqs
vcpU3eJN6nAqUI3urE99uCO7ZNon1TjSAYUopHNEPvziTf43yFKo/2lw7c3MVJCF
pMn0Y72JygHB2Ufcf5MK9pTTTQg8z8znboxWriNbJ+GVFKxelYS6J5Evzb4rbUyl
UQpw+bMms3vCNIGCPC+Y0y4WfKa87cxywmXbs4KI5Hh//6SUI2FaZCq4zMNcZgnO
zBXpThvMG6VIS1PIZdmPTg56McB/rBH+V3weo4C621CVWf7h5oSVOfiMiERtBRJu
S1x3Nzetf18HVT6pHUl7LCGFRfnwtdGMYhmImlZOa2NJD3i2p2iFhMM8dKI4D9XT
nVCfX2MoRUXSRQb8KUGwX0sNzO7tMTdp8J9ltDios0CZH7N9YeRv8kK5UxmrzC+f
VnD95NDB6OOYpzBohpQ89ESyp5xV8S5jSx3kHCMtqaZBM17rmJAe3/lYMaOB0Vpp
L0Q59gdSP6pcD59xw47K56d+qmleFOWkVlAN2V7rLjwtIFJg9gjWSIVZPH7W3Api
OJko3lTzC/5gsDyQsMYzSuqfalkQVEiDrPI/zJNeCoxo2i1gqRLTqBuO0IdgsdnO
ewEBjVdJw0zjDDUK2JlAz9B+Puxn8CDtvqaGPO02MPov2XXWTRrliL/oPBKbsmVK
q+whwfLKt/i2ubZnRgftoqSsCabjTvDvd9eLeGokVF6z6xetxqXXUGp+bVAd//wA
HkRQFkGz4H9IX+FKgECoZAPOwb2fAHfDzEN8YeIxquZcWEjXe8ce8p4/8Kke+Lvx
Nfm19C0fsqej6YchesdJKQMuWU67hWEzPJCYNc+5coVVnTdnlcAXI1sNwqeclyu2
Yurf71lvv96UPnWY6t4dyDQwv8/dcvezDRl0DuvK8PJB3i37jPgZyjtBjy6JUD/z
uYxeSOJWjRRz8lKEq5N0vrOi/Xwa2C+SD9EKjxkr/BiYvHHjhpKxX2yVWU8vFqKx
AvBiVZVcQEjzpezTUzrO1aQYypTaSv72KQ1bFuzWCzlb4XsBhTasTbhT2KaiFEDa
i2U9JTp/hy7Gc2/YolaNPtsVohXhMjn69+P+9nznqp+9emuMB1u7E4s5hvhy16KJ
ojANnZrOL5pjAksJuL3eOPvf6r0Fgwn2fqQ5mlR0GhR/5q1aY1aFy9jjKosc8uDH
B20i/0N188bGh/3edESMH7wr1wZMahPqnQQapg1tgVL6VrKUq8XqPuCrEAaLimkT
ECe5s0LbkYu/lxYcmcMYAstBL5DnmyP0LPJ0tAl+uElTKMwt8vFQu2wnsgcw9Yfw
mFEEYUjRvMfjnSRKYz8KRj/QtL3B7570jYTg6gvTYwV7OmWMO8RSsOKmplcLswcW
lCC92YZjM1t90+yWVj5zXrp/q0p50qkcQ7JMPDwNYUgNC9IECVRlSt3jCjwKUKjr
soCnKRHURzIQW0sfC44ZiryYGuQblCY/GMDbay73jhUKtUAj+to1tV7n6zr88bzf
9OPF2t434VOD2yVZuHScGK2+rH9FDvBk8mK4Fjxp7pQRoia2vEuscDinK/xe7PcX
6135Dxcu1TLXHtsk902k3kOKFuS7JuxaMBE/E3S7NxHhH8hjNeITfp9n1nQyAcQH
n6gt8ledd3sjMWXvSCjW87yH7yJYUvAawSbynN9nEcDMGnhvZgI6VeTT6QQHAdmR
usxv8vi2H04GSG0CSb6V8V3R9xPstCFnPbRhFuWBoepDVoUHCHeIpW+6e8Kt9+ou
muDQ1xMZY/NQi29x99UmYPb/YZgFoGyp6NFk08hrBrGsYSq3T7vPsi6mEZU2Xkvc
3Z+wg6TkbR3U2434ggrBuFv0vW/3RePK09u63vLz/6Zp1n4pErYNmbu9Z5iry0v/
M1P6TleNIs+mmt+CDDugRItJrjg+1E0oywQdoRfDERX/hapZfCNsC7H4H5/8ywmX
QMDK4EQFoWj8r/VEoMUfyT8J2z1Q5eM8CzPC6ynZhJRcxGWG0HWBdMWmxlkwt9jp
a4oZ/3/JjY4ZRtAsA3v3VaXZx16ySKLOqKwjrSRW3O2fgsCeoc6jyH0hUHr2SESs
wRBVL2eUQHLSnbbZbsqHsfYG2jMgMPddTukeWMHWWV8qrLgLLwgiBjgXYptEo605
ooBZ8FSMhykUVQKVVxNhhjfM/hTEdQiq6RfY+TnZp8dXJt0rxRnZX5VRLkumUWNK
8kmDzhd7SC2VyTF6qFni0L5SwXy+OVFnz+aOuU2i75jCE/IhrDZ/uTe8WnMYb28/
l75oAlULZ9uO13fo+d4aNrxCXegxfJgaRG+lo8hzfUlqB0wDMbzvwnf3Y5ITMDf+
c+Cbu6ObZrpHz7h5or+PUi5kcIznqtcxxmA7dQMUZgpZWXWBdJ8RwyOc77cIbGSG
tZN4trJMcJ0yLL0IOueyLyNiK8jqJS+HV/AQKTk49dKUBiADX8VY0Q3Mt5b7Noze
30D0wL1pgX9S9yO5dRSA1Rp2ttpxQgRxYygusHn3kVx/ue5xiJ1+P6IdMF4mH3HQ
yc0KZH9iKaoRLxKeNyEAxqYPKlMfa96QKk4pmUHdHlpWMZapXcspYAnmAwP9Oadn
eCFJnh5jy4FDvdHrm9NrsKy3l/xmRseYUoNpCaq/dEw+JM+23JdEJa6TeD16VT5j
YApgBRAUSfwiWt0T7MYNDc++Jr5f/fjTYpB8KM70UA3BzN91SLdgyUB1dTlvm9t5
hP4c1liju+jJTrVU7/L107LULw0rAXliAKll48MKcaHEPSw0BhyXd/C/CnE0wEn2
FrTbE1oX6DpuFrG3ctO0rTBpVRT8XpA4rLiNZqXCRMMXMLse0Jc7OjQXRoxqZXop
LwR0JBdMPOX7le4uZ/rY1/zQ1b6AgS4Tp0y+5VoQxis2AAeoh2q7zORl3xH+v+7O
guf0ollvNHVSHGs3KgX5aXS1nVdh14XewzsJVaPt1n1P16n+kQTnefzrg8qt/f3e
ln8QDvka+MDlkjwQDHZBZlM3h6ftuBh0nNB8HlMnJqo/FJMkZkNCc3HruFRpB9qY
RH+PkC4Fg+Ms2Fr9Y276gip5jrjXJzHZSLJr3veK2couzHThHp7kFE+TBGyb5MK+
a6vegGeltKevtH4w7fjteheg621DanN9Eyw3LYnNKu3ozUkqC69vjKkdq1JKv1it
/X+7S/4/g2uBIVfVuUJXuEsD4bAfgnX8U+/O7G3aIR65EaaEIuzfaV2vqm7p+1lW
e/Mi4GZeLFLkip2L5e2gd3jfuaSaXwu/nR8fqRfUdgbQTkoDyBJQBVi8MKFTfvWM
ZxfGqGMJxjolhKnSOvxfeFf1iHK28UZjKt4UI4Yr8GyFB2K8ncyQGxdzkbVzqH6n
8qIPYVj7yzOBapfrfd4LHwg6VLGAWZsy9EGB5U08GzQGaz9a6pzyuWe3HzuxSH+N
Pss/MwPHFOypbNq8m1GCBGJVef/ZgMk+F/zwjNZiRXJeaYJDDtNvsELR1LOKwY1P
WQbHyfP/GGwrMDzxPNtMSqFqYkCx/6GJZBhFclRbMPAfdfbAYKyjSeSA19vfbLbv
RhIFQjZon/aRauHAO5P0opWMen1wSLowShm4cl8WGvhPLtETQ/97TbBrcmPGJsIf
nLiMoBjOQbSMJV5Onuh7VfmYBTCvkKs6TK20AVB4K0y6yB9j09HrG+k78rEBgi9f
Tala8HDQSgV2IP2x3rR4ie0uU6ewB+Cq5CRy1AgIK7DLaj7LkyI5CiG9Lfds5DaC
bNkN2gBvkVcJCExvqJY1hHpKy4XO1rIyaBvQ85lyMFSeerWgmDXh6DlK8LBml3S2
P7I43Vs7JsqVLdlr9UTPmv8+ec0WO47KYFit3Xeb2Svy5qKWX4MkLO8+60laEEZs
XTNjT0FpdHtQXxCZy2KZXJ+HbgB80MXcZngDy+xehFFufYDX0Az07lTIVXMX3ilu
YG0if/j5DJ8wpbs7HSO33Z04J6F6cDxl2Im4qqruLKad6AR1qbeHreMwVfgi4bCK
dZKT7mPi1LMJyL54ELXAVQTohEbgS4PDnPfNdgvaJJOyoQgNEjeyKcbE02kO/4w8
+U23+ksVCCw8NWpcJhzjvdoqWOuQjjZ/UPkDisd/SMyc/MmyB/hNK9ZIWx8TCrGk
J67BybrX69qwCNIXuf54bX+rSTeeTKm7dBDonHcKwnFen4ux69WGTN1nDB/hrpkJ
tVZc8WoAqe0JGM5NBfmcz5kSHKJ3JveqGKpcVnLhkTthD2SGLherLrW3nydzrahM
cF10WoAnoJ48fORcNZIsowy6JSnazl6wFhZI6q3CjIiTBTLbYXUo4bqfBYZsT5HE
ClMgtp8M6Zlnj1yfcIuS3v3jca8HTIoXO7xD6QJq7czCAA77h58YyY/Vx319vWsK
lSEtQPxYBWWzhfupnJjSFfIcsmwGDrDXWfQEGmsiBKTFr/KccmT22p1ZLu4BAFjn
U/md5/YJCn0UX3UvJlez7nCvSJiGjduptY6u/DZR7uF+OxOH4EQUlFLLpD4IoZGo
VJqOFNe5nsLvdz9xaehQGArJ7e93wULBr/kTu49gF2tDLAftlCly4Iv86p9Fcs2a
6Crwxq9lHjtDaIN3utuf7DtuRqP/ty6h86JOTlR/H4fn4vG3BXDchiqdRldpSMcl
djYEoqBnBMT56dAHuc+HhkGME5ZKV0kXk10grVbgyTeFirpwdCQytygiXjvlSjlw
ykqAzfF+qepQnDYMwmcN6iuzMWlG8hrdSZNBjfsRmbccg3NhvGaaAQKNaUKodDB7
SLSB1ilI/9nH5ZAu95FA8uyBhvBvh+ljLxTZSlG7b1eeSGaETYATwRC5QZdW/Q7R
Uut5YJknm+bChmdCMgExTIeDxY9Uf3uDPBXsDPyZysZb4RpCWempCnA7qPeB3kGE
rb710GS/vTT0GAI/+fUUFVK+SC4v7J/bhMp6GK7q/audOlYtpfty9kFXLclyP/5D
ArQVyAOaU70L+ODOAnQT77Lgj0hBpb3UBFbghUYe3USainG9ya0L5n+ARhRyE9+J
Wpz2kAcEB5qpFJcUGys3uhvGZoXsiVp4f8mqUFJ5YdNA/8HUryA2cSazSByQR9xg
Tzo32Ob7ETgWpzuT4XRlmArABmVD749YauIXtZgtyAgPaS8+gqdiAeeDcUtVwRmx
WeGl4IaJmAXcsqZ/ZzpmaEw06it0rqT4yASVTE8/eDYqMP+wzpMdZL9oQ8Pksu+d
M2VYCsLgggeIWIb2R9NTv4IOi6+vFZpuHOvTUbf+AVG4mxtOqm9JFRVf7zJXu8aA
YA1Ay8ET2YhTKJ+IllZKGD+38IZwlieOqQmVKeknX9RzsHjMihyZAN4fm8Z6VCfu
EXHkMJYayPB2rZrpXLvsi36oty/yryzFvzXuWpnbTcyBcV4B0060JOWHwPsmqqo2
wYyueE3aZ4RNE66KTXqXsc9ENxwUvPWnjMyfIEJlIDQ+9qVzG8Tto98gAuBgTljb
KRYPRRjtd3t1oLKPs2upYBrKPs8wl2Wpxv/HhGX7pab57/8CDovp7bC9M1nx15nF
OOwdjacI4AqYIIa6Cod/lZi52AVrm3uNRGqJAR6HpoAUQbb/J3xzp2LwuqEhLIKs
kK85pV9orIdJMJxxDCMgji8ycW0PzLQcfV8l0KQvFiDqVyTt2CwPT+vwlLdVROfF
Xp4olNu9yoreqr7NyPb0F/paR1bh8LYomSwfVOCqpuQpcjNIBr6OOxM+175bwq6n
5XzAsO07okfiTeapBQTWHxsyTZat1lzSYHAZnOGzuwwW0t8xHR+GiVO+w3TGrE3W
0eQy2dIILL1+LhjAzcGIlJZ12E3uq5lLiJvj4mcx36fCPM1pu1zcsb50X9Ru8VlM
RJufJPPLIkHk3gl5yRmneqHspsdfmuqwZxEis6biFW2gon1IpWl9dCDeKURyibLY
8BSgM/5yYiwGdISa9/dElfLnGFhs+pMVQYSv1yCJMACd+7rxjpDHudnGGLiQX9J+
om6f5aZuv9lwJQ2TT1u6d94Iz5SlGHwIakdmZFZJ7OBlcypYC++bht/+YwzreY1S
Yf+iDdUd5bAjsShXHH4wf3Zh+UPCfv7671qGBgdCfF58z61AaoTKDAv+YllacJyu
018Gl93qOf94BtejCjBOUT5sTKnAB5RkLZ+HGmLfE0RJBvI+IleE0cxX58MUDLiX
0IP5MXAnWksLPMwb+y94fva8IdW5riNlIvdK3ulBrPibQWbb1KnfCTMblvBdd5Gp
oyA/ZjB7jjzwFBPtQr0kjyuLtZRQwd0Jn0FdAg0BCrAA55UEewCLpVnxcPDP8n49
mJu0M9YCoMGADqcCrE7paA3XuV+rwYX/Opm57BjzoMnkpLQzZHO0JFxtxp9EZm3G
CLODwXBVawMoRtyzRizfsYokD2MxvDZkYEcU8Sogi2Fc87CuSY/JEv0Vw5vveg7h
TArtyT5yGqdeR1S5XJnwVcw6X9zywTaXuagkcMdrs47BuZkF2KUJbI3zKNPzodeH
HUS4hHGTey/1Uh5VNNRhfo4OjuGXqigLHx4OJuJMfn391GwRAUzZ2wlzscF2qr4O
FTmYlaQD8sZsIyue4Akqyd1GX9mkbcIbd+5t2bqMEXEC4ho9YAzwVRLG89U0xOEi
/FSnnw7QV2uSiXpTJ1G0ioGFtEaJbignYksWySxgXYnpyFn6K6M+2YJ95xNPa5vc
gC/JpOjuQFiFXIunYPOe7h5gQcDmjzeL+3yQaWEoxbmD5qJZXYlqNGNfySZ8jz53
ChNhP1j5sIw9f1avH9UDUrfngQz68/7ApIAfKJAImMbIC93uHQ3ogYL05IDg5ip1
GIifk2k/j9qujsfdGI1d/s1vc4wSEPkUtQbGOkrBKzojcHANAHKX7+Vbs1B6j6uT
qKThM4SKiDJCbLDb47OSu2oz7enmealqGsQdgLMmFvkuxSiss8aDpVrsWj+DjJJo
GuowDTU2zQFqe4Ln+Rw6gskhbyt/jZzf+Gm66PFp+FVM13NhVvKJMorTnH8nifpY
OhBhNbW25+0lCJaJvcQyuJRIaJqquk65aaiWLfn56M219RyHeqcJOLCuOr3Yy2zF
Bi6cGvBk2MoTm/PYdJ2O3SM2uNZ7J1MbtnxBF83JwGCmx3De1xINFkISQzq3jJxc
TfQ7q9GLkUFNaZBkZrwjjSh2yqdgoVbjipte4UIjwWEp1ztGrcyi3qk3ROmKfch9
4kNljFaU/8FP8gwWyUqukC1mp1UwRDFHeaSYA+MGqInQZF4XEbJDM+3FmzjxTCHH
AzgtIHbXrCCR+t4K+clM1l1WKcCuTNWlpsg384+xxGJulLOCSNyky7Y3hepoTRMG
t1SH/Qhc5Er9xSvAo4qwOsdSMk6CyqAf2bMni9jojtMD6k0E8u7exlPeqDInx/SO
g6cC7t4sFChrlhOzkClkMXsC1IdM5X8vpmUZVB5nvtx7qjAsy9MXmpjpIBh1CQzo
QcPhS9bP0x/Ne7oSoRNFfpNCjIbE+qSMr2hWtRmOWx7+DmzFnSl83X1aZsU/mrQy
7AoDILBLp2nmUDENX28Htl8LMDjlw8JaYkw0P/nwkfsNux0ikhJ93EON/MvIVfqa
/RcgSEHv6hwqYayVemXM4xEagRYUfApAsGT+3/zuEzqVR6OcUzLVnGqRGo20PoZv
mMj9Pg6Tlo5nI0kKP9ETZNl6rNLmr6MPHB1Etkm9K4nTrhlHvk5xQagE8PdC8uTA
xbhPyvFQK6rXGmp4PCfCwvGGnzxGMcvnkWoKJmgTcOCmRT6wY+hKADhrniJtCN2q
ch8B2My/bgJGCYFoXfKGBkKMeA9Bk1WMd1TTICWKiv9p6ItaGD+2UmHFhHfjaNgy
2VdDYVGzOVZGjAsO9d2RIH+tgBEDLU4Xe+1UzUFhwtL22SVs31e+lVT7B9epl+PM
wlnwCWTuZGMfIGtzOrwSdR5FdQPhj5XHiQ8+r2M8T/GkGCOvEBKDAw2jEg4kT3YQ
cQ3MZuspjrLv5BJLHHBArHdJfhmHDyJdbtpUg95id7Xi3dcYKAGfBhwb+KiEdjtG
8jecZxSdpQsIhMDQqHnjmgYtDKGpg3yQWrgh7WVCC0ooIKZdohRe73XwxWqwbby5
AtfD/dS+rqdCZG4bGBoIVI+lj7ACFF1ab/vAW7yFcj02NG+Y1cxtu212clNUtsL0
e80FXzjYyazf2veNsSriq8AMxnUiBUePQqw8JeKOduoGOQQhBbPWCjZYSdmxjhFu
dzULIba/V99wYs/MHkY4XKZIK9fkWm9YWZcT3+1TJsB6/OHUnpCVCBlNZLBa4Xsk
lkKY66PvsR5Cy34Z9cd2+gQGR0Xwz3vDi2V/X0Qlc2TWTIUEQfIrwmePMCcl80NQ
nsMW2k+n4ojIECgjsZa33fYTy5R+1OVUVahIlR6FQT69BkhWRY3Q1MVvS1iCi9KU
DmO0V15Iwui8SvC2p4Av0eKmKi7+0Ctv9UeQmGrmOGdTsqHg9eJJlzpQgAPHEJ2L
ui6qMUW3N3wvpXTJdjuX1iLSWVUXjbmjhwqhmxXLA0dbXadvlQuISH0ZJ6gRoYQW
qRG6B0fAvuIi0/m13y1DmdzTQbzrVQgFivqDET+qF1eICj7df+HjaFN9GTRAXA9u
CXl68QUWggTX4EuhhYACubMsjWWJ/RGp8MFiASD/UF+IcFdZYj1xoxTs3+oZBo8S
2JWhOqApd9h1LMd2kzBGb6EYx7RLRiIIFM2Za6ySm5Oys88sIPiz/hkFrFVo9sPS
EAKLA/sjxCgZVF2wgM9MU+xBcQrhMDGcvQcRZP5p9hjdelJl7/o4oLJjoP4UdD/H
oWCf5FjXC0ge+DcqvFv1XvQIzzTiEspbyEWpdLQB9/C1pKIDzMYo2wZagnA76r6K
hcBHme2QDTgxA/mRh24c+T0pYqSe3nPEhFwCN/09Uq0zHvKnlqGU9uIa+8tpwRNc
6c1uoKQSKK4wqxuMYG1QWGA43Dufw2sz0gwLjh2RNN0AJLR6PUMNP1tEM7JalYhT
197HhuLeDrcpU80bGuN3DoKHksEByc1lvOViHuEpwb+QzgiGynd7gQt27RbBT/lI
KWWWDLKyFLKawKLvGI5odDG33WoKBgV4lzS/HG2L6r/fDRWycS34BqyorXZ7cu+c
Lmmks3i5LLUvawR7aFpwVIoaFYtWDL8mX0Njo1hyWS1ScMHSACyubWunHO9tXRs2
2GdPN+yK0RgbKn70XkYufz3bfJwPy1LeH3/IhxxlECRj3dqBJ4v+7k64OpMSawHM
MjEQsaP0Ory9Ksz/edIEmyGSIMOknTEBDoTVqk6dzN8Gt8xjvrR98GLsiPKkMxmM
Ia9ALgZdfwCgcZT+z0heMIRZ0+cUfxkeKDDyKqGydD8xgMq1fgFd5vCQAwaOYTTr
WWeyZQYZKfyjFuo4iw2Rpm9H2jysYmeW/rs74wUlFtNWQhgLbXVIHtFrOttGRn7j
NxAm4J+zr/tqXmi0ZyYhZfkwkwN276svEwhWbj8C1ZU4/oOiRPVHAuCxCFnREKhE
s7x9oDSrzj0xn70B3QshyJALasB+DItgicGE5DPUOzouDOZZTSNGFl1nZZC68vzr
Lhr9a9xXRCLou/HH0PTwFQwYj+rsCF+EMmanzfPlhEk8YB1UxamrJfm3U+W93KUr
lJ332zztEJQPXPHYGBA++Xl1FOHiAU/FjE7FDNf5xzTybD8xUXOHhAu9xvci+B7c
BEwt0n6SVLPvfUnLsDy1l4hGD5Us9CFo4ac7j09qIX7EoVajD7vQibdH3Zl3IhK6
tthkAgnGhuWSsse1b6ekF8knVId4F9yZDv0T6TVUl5nHC7U3R77aniycGLkflzBT
W3mBIz9eCbStFqN38XNrkvC708QokmwbLIwHTfX8yIjhLSBi9u/xNFSmglKxmIiC
36JHtoHc5Re+8VCEZxGSDcDUV3nheIyjAssCsRB2CghO5028LdOkr+dOZmRetsdd
R/bNJ4rXBPH3pONktq7hVHx5QuZClpGy6TnTwOFGkTy/krmLyzW/sWvV50S9wZvw
jE0qB4Zjacmfk9myjwSs9cDZVkXumPRXayBrT44J+YCEFcMyxnmGfBpmtQ1jeGwB
TtA0rtIrEOq61kpSxtsYBdGfVKX64bl9Y5fJzhv2zCSteBiWJdwA4jFb9dCCO+zi
ovY34dzZV+ahD2BUjCnAEl0SvB+IcltYPeGNWo/8JMt0fPYJpsqHCT20BnM6c7ll
kZjZVl/NZpvA5ML2fGZegNJOIBi7d5q9/4s4jjsYmAvq3paB7sqVF/rmPINX3FBK
Rh/G+bWH8sXbt23XBnRFT8DQ2+s3aG4+Qh/q3uvQKhZofVeIijfDvSxSwQF2vhwy
EfKMiqmRZNDMzgnVKRV3kx5YQskZZkfKy+lXi82kX06ZXYYhJit6B1RWwzdHC9fU
lVaridgm/6332E/By/TMge6qv1f2ajzRus2ib/FVL1Or8v0YWP7u6wprCF0lY7t0
iEixlk+C1zc2Pr2qw9XTxjyolg3fSarFStBSJb2nA4xPsPVRHsv1zPj0Sp2ix0LH
mqwFh9B2/khsGhHObdCL7/R3LXJ3ISpp5RGxPs79OUQnBBWfmuJE/gKQHAOjg64i
n5hPUJ9lFCsh+pGMI5LaAwMd9QVXU/oKPQJOV6jZNvhgtZcK5TvVKavFgCDQ9Fnq
VDlPKyDNTwFdrf9cR4EBokkMGZ156HPlLwB66js4Iqupr70R/dsiv167vBWFgbxT
iH+yKaHXP+C3nJtXL9Pf5AM4Ip3jH1qDEhsCVuGgGILHuZ39+i+CvdrSoiTnFqsw
wQv3gkjaCfesUYglb52IlEAglLu3i0b2QtEMsjHwCFh904UHCa+GYP+IwHlzf8Ld
RViUyH2saz87/BGfameWTzxP8PpO7iX1otqz/xn/jODTiS+pdOJE7ToiBsksnnTi
+umsfcz0TpaqM63n8H9bHN3hLovupxVmVWp9q/xhq6SeEzCRkBGkfTfOMFJsem7p
r3OAaZzz8uqa5d3IyRLyYhghumy2kp/KT5gOGuhsDyE+GE0Yrrlx3KhaLJzme2SL
3gMxcxMSBrHZ29RyTeYLE2nQnElb/VuZ6lC+WLX5AanWHZ4fE65BKJ1k+vdq8RYT
ML1zNpfTv+xiuFDGSl30XQgrJrP/M0qFGgGBMWXCiZlnOpgAZjwwt1rmTyZKELf0
uaP9kdPVAxmYh+oqLL3HsASsC/0K9RKM1jCf5Sq+MzRlGFyDTXHpOAygcxEMILUh
TxPSRVDH/LW6YPriFJZfqYv1oY5MlGI3HoLmEzxssGlW7GWZAqI+8wUlRXA0J29R
dfUQ2zhANfXbiEcb+PzerDRaL4Jz1h6MJDlcbHKa4G7kQgHSSijKK0iOJiam7AyS
QRtqluIMA1phPno5KbyuTMQ19bO5/VPTmwoUT1AHBa+MWb8hzBbHTFOFw9Uw1okN
aRw8e4VJ+P7aJE0lksBI+EaMkD4e4bNmXi8BCA4r13vfOLNEUf6aZFEz8Jvmjq+o
dUQA8oqxyJE2am2I/qbFQ5mnSZ78Sk115NLCLOMwYYHkbmeveY4ong69aR9jesqu
tekF0IwbCdWu+JC01TfTAZnLnLlBCmtH4A5+0OQatl3jvEr9kuingfiYwKlkzsRh
EHruD+7t0A+KNj19LYCjwKMUtLejH8G57KTtlGR5SJHOhEzkHZmtLNBK55V0QhYz
zmnmzb1Skp6UMZFMB63vUgWoDaz86AVYd3EaBcBH4QO6BIkdoYpy1D8xRDBMMVk5
+nrGYpOJfRP45FSzDOTBtD3/ZkLH3UbmIDYfeoKAFoT5BTj3NkaPeIEpxfqAbS80
IEKdXn+SdFUeTgXl+scPZ2RFFgRblCozblx963KvJOAqnwC+kUZqaae0NyA4b6oN
F5V5JEXEXfWXCAoS1CMr7wG5rlvSU2SPvtslJ7Vtd5Q+81CkQmjCE7MXi9TELThQ
Ayy0M/FKZTzGIpSWB3hPRbPihFSvVFVRtP1GurGWD2TWNsF5igHH1i/oNaCIqC0M
ewH22rYuzl6D7kvuelJlGvvHC/7wqdKNDye2nPoU8mvRvxHZNdEkMzKw8OfqYijA
xiK1MQKLZFMvb1Fqf9UD7+fz7XMQ9VntL5cJZKy8hADIxA4F4jVU/SmkgAfnkmB4
dYkm190fNTNHRE8zRZrRFyCZXDU+GxnVTslyaCQK40eesaurt+AxRA1YUcq11uYZ
MUUQEvLjYu3xg2Bo0GJOA8Sx1DIl2+hAXXr1WCUcyjO+dXjz6mdMZLEqUsyInokO
sB8WTjblDH4euIoDXXUAVah8wrPog/tV8Pl0tpgCnH8E4l/5ZdBpXcAUf/s+GBNX
iSZYL4fUCwZ7Q40KCKiAp/U+UhjS4ye53eEN8ZCnWrycpTJmjQlV5tnDHjOq2NOi
VT6VZOrcOB0bcF6zA9Va4lOtTqxgKMAmh8cmiyiunrrVMZ/NOODXrQZwnqYZ4oXx
r81fSJUU4N51TQmV6Y0hYom3wCHePyOAvA0RTDHEx5vYUqXpXKY3yiUAXk8efASY
5kvVT9/aKtdCgnxbaJazwpQEmnIaHe19Jcb0MKnJEijNBAx8mZPN0YA44QVrmU2Y
J3TBkOoseJUHSm+JlmHOl493FCgGjiBd/wQdP62pdrEbRdE+Si2zHGwZR/YHIcWy
QoBAP8J+C4ZoCBK1e8ssmU30/0ocBmcCsx/pJSpoB9KDfJlZXB0Ffth5qqCzk6Bc
/3akhcCq11JwzsX0c4LjnWk9IBFimbgRwzrksubuvfKLy0BFyewsrSFdNWkUCP4z
4cgaBjy0IGaFW/hdXNxoWEIM6mpIniNIkQvcybarklQUsqgdURmPmGYPlvWmVWRD
sz/Qqkb9jkTMgFD3hEfrGyEqoNo6++aPyBNRuEE9Rf5HHK7cfLNFrPL77fCKXOA5
I7KtKa1105IBIwYxaXGJ7jBxz3WGvmzi9ksylclfhUzYvZ0mzzpUt1EhrEleZeHa
cnnNJTDLxOIKVMuTuMB+astB/3NnJPbMFJnb2yQIEEQjJLrXjYsxH+n/3/ESXNd7
WBUjhMuGwU31KBLp7DLclLmQZBfjDUzHjfw8D0XKT4vuMnJd6lENavW1evm63uoP
f8b8aMeZraBHHOLJropUEd+fSoC7UGH3YBmOcXRb/oWq2Z6jfFvLE4zZqlgfRrZh
5nSmKJIWCUnyoyFZDtvhGRDSVB9E5QcSPz1FM1l5rE84/DwNcReQJ/e7mCuRGlka
sXRYMwGtweA6y1MIZS0LyNrKV6X2nFewyVs0jqn5Yfs9EDC0ROoHC7R3i+PmEe2r
Mnj075Q+qD2FTlKWI/cylH7xLggMH4D20OzL8qcZ34mToMdZZCC0FUfUqFzR6TRA
tisISUmkd3WJ/sls/LYY0zC/89G7OGG5y0fO7iTDKBkRdMNtd4mfWVycElLLkrXe
OJxrpRIPb7fJCNi8FWHSsixNg8EwhMMHJ1e8dbajD34f4nRLHyJ7DnDw0rYMxcJq
q2iJVhKYpYwoVMhgaX2m9Cf+Oj/b8WfMcXhTHhPAr63D6AEM88m5oO8GDLJDApLb
wKsc1c0/7pQKIEX4S8uPhrlobliM0ZqVqRDX/BMxbd0ORUhGiTYmFyKpLx5lca9t
L26EEL1WIoX/4FsCUIRgH187jP/EtBLPsIsJJxlTniG3i1pfOQ6mBjr8sot4PXJF
YRshCYXV7YTmSfCGm2LE4WAdoPVRFLmwaQ4Yj+ZI3NOmuxDKdyO5w9XUPcJ7V5yH
m3y25pm3CWuiTt6WLhwW+/GH1eZL2Balp1BAIUauxXd4l9TJqVj3XO3mJJFo+Vmj
vM0Gt0GRPicvJY3CH0vFP7glrW81+SareCsVBq5+XNXo7+LCA94N6tlZ2qUaitaA
i6tPeHR5bYzPNbvRt54ZiuD5hqidrHaE5woww//zpiOvYt9zqrRuwGykaLiwyYNW
J70ixGc+TnTS8rYkS49btwWl03GneWWSZ3XWoTq8qbXVNNFDBlv/UuTRZ7v4TMyl
pEt+ciH0eYMg0AAaxj4E5kEtIMyTwjRAcsvqhgyo8/1ncMzTjrx9mEh3jj1E5Nb/
S8ES0oKJG7xqHPayhvE3LdjhEhmE2u9pAkl06NWJC97rHlV/VXSAqacSP7No7CmM
H6u61+OQFn0m9A8KmYuM2TBQZXsflpImr3QievI5h3XkIql53TiJLa/JXJGGBeql
W1myAOA0izsC+4N4NsQ8JzT/hZbbZgjpB8DxRTnfTTeK3AmPJ0Qei6vcdQ+wspp5
k2OGZ+8QttkZwG/y7WazdoFjSHHzKP+tcW+B2AYS37O59zbGdq/GvBJ3ptvxQs58
C7fORZfwhkEfdTn8fnQh+0oo8U2y2cW61zPY/pLm759VSVs4wYY1fP676/1rs1+/
R59YVb6Hz9apEaPLLoLvfJ+hakxBg8RzcSI7Ul5/RDY0cxxyYmW+GpUNjnGcE6T3
ivm7GgkJ+yAw4yAnUoiPqY6RIoUuE6mFnacEPVrk8aNMUXspO5Zv0AfMN4WDpqun
+RWNHHsAuwExmgUBGYndlQ012GN8KoUE2PcOz52hHW/Gw3LQUAkSdYiWehU0GRws
cJWWjdV8l4rVG4GgaEIZNWZ/FazhhnIImdrNkmLhkBr2fuCTFSfkEOjTuJKGek68
A9XLVF8dPgI75Brf4FWTBRGVLJjOwS9eGlB6oM7WxL0EsWoQN+Euv8gt7mzTXVub
3W0I2Tbchd432mKo/CFO7DL4z0ub/3OuWK1PzF00ZpOXyyFvgDESTrEbt2uGG6bv
zJdFjLT7pqT+UwcbaOUbF4fHaDEeniv5Z4Dpf6hZHpe1DfrNg4xeKjEtFt2wwXDY
cLkSQXBGiAGriNxqvfX1Mjcn0LJPIfiBm3ktCn6bYljTA8zSvRkEBiHjf9+l2gZL
eg630F/gjeZcAt2/tawgs1j/JoN1BDQIvB3HFpXZRA8Sr8PoWMOHYxpQlfjb7tUT
HyTA7g5Jde6OgHewo+oTk+RYEKZ479TgS6EyetUS8frlr9pMOyc3T6Ea675OQn7L
gWWcrS5f0QiKdhvRodUZscyj3IWpG6vAXxYu6pMP745qECNHIhuxjBbWJ8kb/7A/
H3aQBxaomXfrWuMXotKLftjmV7YTkNecGA1DGuMwQTRP8pFkikYO900WpSHViFAu
IV9um65jQzjpYT3erYgMtQprcdJwoZMtUylKZ9CfMX62wdnjbpFAs5YpAfsKGace
FjqAO0cZtIYexBPm9wl4x+vbyUzXbF2qMmzAi5IfBTURxjgvR/gUup2L3LUX6GCD
4mH4YYxMYh0Gurs6oZsFLq7bZZre6dC+hYIY9AkM8Ojq9/CWmsmfFL79HdwUlMmO
M5FRR9HxEWFw0/pINhxr7HuPshiXhwXTFfoqI+8AvPlIUypWZGMBHZuTQnMUJx72
xz6godC+JDXusFGBN/sDHncX/+UdSz+aJawmtv9L7nx1imiB03vOhc6L74panEdF
JEWCTDmH94yAy4eAzvQ7mFSLulgMNNs4//SXvu4YxTwFkI51fW4Asi8zDo3cwPWj
KJliKaDVqKMBtdf6xuLzGlEotikK7dkuV9iBaZwhFtgDmrQe4vabpxA3LTSCuW+0
1CwdWJiBJubu1GKQBCxInwNI8eBVrEdPDVbTZDRrEVQ3/8uckNAafdWFs47Oa4lZ
4yPm25hABkhzhOLXDntRnoG9AFt1z0BStq/r1Usw+YY+xd9uFwQj5wFCbqHg4liT
SrcYI/pc+wHdNzxkzuzQAanwQGrtlGMJD125ne3XdSaoRTWlTLBJCZ89qvSq+v6o
dsxEEo7Y0yxJMljhMpV9aOJP7xMXp4bpdZaVUFcSwRQk5z1Fy+Xr/60EfkVcgcEX
ocXqKt1FdhzTA7AkYWLME/t2YpCUJitrqunv/8g7DXH9ni14eA7MGRUdo2b2o5zc
qBtghYKC+UZTXuh3c2nQzugq3Qo97XYJD7NGlPSi6yzxLIe+q+rbx+/5FBmTsz5m
VIm1Fo8QEdTMsR5oqAz/xSQUc7rbc+ac7/d6SMzVTpzdB13Zjve2QqyS+jY5cwcx
ZvlVr4LkaQlMzz34aOrUG2kBy+M0csQJ82i383YDXXfeOfHLpZYR+I0P1b1l47kx
2Ux9894iZO5T0mTUnMyV61WvMPNlYYaoaNviGbhQrScBbvvvK9gnfhbqbjFzXLkk
y4rLXj3cE0P5F8DL0qbHTgKJ6zCtB4ImfClJN/k8vZ42paMA3H3Y2L7GlYLwLomi
KkByVxMth6gwUIisoIlszm3bDgmPzpsaVspTk4mzzO5Lg6d8vlodMXCWb5SSIyDc
wlv6FbC/eKPco94L7AnXGOg7DkAbDaJkUBVmvAG87V2MGE23hc0/L+m8fHoHX/DD
xkp+0FSUlulWrcPUlvzNyjUvUGvYZd7UdkpfYkhbzdYZTFd8wo4uE308cSB4Fogm
KL7lcRir2LaAFNpe1mMb6a14DZ5m6MJd4a3uQycBuieAz9/l1EhSj8fhhf9cUIk7
ukYP7SyKh+CVUshzirr8bgyKzghJG0IVBGmWcYWzDwq9MVK1V4c+k9Jlg+7OhC1l
NMLOAzYeZoadICLilr30phi/p9XLyk19g7B9+QNr7QNcEMR1BGr26uFI1og9puIq
zjQhmILL2B6406Cgt8Zd8uP7Y691AxYF/thbc+K19jyNk1sE1+T+PUcLL06f8tWI
rCBZhZYUUC3JW7wpp0FaB5rl2JWtNdGRLv2sqm9fNHHGzqD163OSFlLDAcaeorl8
1EfUGx27bEmUlCdhrxmjNyXHnTaURfbnUgsCy+zr782y0B2j2CFpmSmoOCgI2mQO
5saYmdvKab2XFWOJZPz/NpWfZ4FMdfJ030WZX9vnxDaxrjInIsV70fPxgrbylosb
0peIMZXNLkTXet3JzF5c0IhZDZIFEiujsDViqdbYQ96Oe/Ycl+QeaAiVM8KHc8yD
YfR93T2e87Vqe1ZulpAP0bZOOngn7xKy284iSFAIo0w9s+4ycauU3rRf0qV/gJlk
tGvWVJQeBUDI4phr3YG0UacwlNUKq4VbZ3PPR+e8g54Wk1VoJ6aCZ9CvoWahZj3D
hGnvEWDH34sGYYAACYg8oWIH0wPXmc+kxnbw2NCB51HCR9i7AG5e6IB8XfpMouI7
ASBReYHClqrQ/3qtnQw0oydF5a5RexY+q4ZwQfkcOkL39hK1bTV383NQRMiaMpKH
FF1DJKJlf7UcYuBTsvbl3YMKRNX5h2S6YgPSgBsEd/m1BTj3a0uWGeY/Ux+NNCZZ
cSY8jKDLLGLaMtVU1jRHBxx0D8vuOufZcC9Yc4aDW6YwKjZQWYIs3RbyGbvPwuai
N07F+v7aFVYdV2RjtLzN4FqDXhFfXle09Cse33XcHWuBicD2beU1mZhZ9LvcGqge
8l/NopnduSWK1N38Te6qGjw1Cm0wD1dpdLBYI7mqkqMh1gTvrYpSMub+P/oWZyGh
+RnT03RKf0P9Sxzb0i5gszwb7CL+fN/ie0eWitWTLB6GdLmAe4POM5KhTuv+/wF0
B0Ia318FcHNdbwOEuUlukfGrR4bkTRoFu8AQzX0IvUGsHk8NYTgtGb6LV/UW2YBu
+9mrJjVH/qZ4yQLl14gTMwbQoMO5OvV4nzvhJqenfFSQMt749pYsqiAzBKH38L9R
ptYGy+vbZ9OoAS8iMKj29sMkf1FZmgJdpz0YTGPzQI1gKjP3fAxizmH48ZFneykN
enAQ3Q8kSjsYr7u4dY5QL/CmFJbtYjple4fFXs6rNI9ayQn3s0sw9RRrVJRXKJiq
goIcExLxOirBnPV3vi9BU+h0a8qH8smPueXGXZ8RFhvEa7LuALui4pJeAKqDFQYO
SXnPdVUq92al4SSGZGkrRkctJzxmTtkX8UwvM2bqUVrwSy27YUfXIh/WkUPZOY6e
o9XcVWRf/c31X/EhgfhPvW0+BZfDbZ4+4LDI0qMWnh4dDpt5gjfZbk1tBZM2eGaq
nojC+sfpz+mvTbok6UDlQh89JiEQCzGqu6qWNPoxBiZxhs3TNzGi2GIO8si4A5L2
7lYhsB0IdGc5LajUWcQEFEAj61fBvNt+zv0L2RW+i3gxBo/w/DuhdqtACVNigSKf
nYuW0pXYsJBj5PwKSI1u8z9cabqwhvE5lDHNdwIpqW0fYNxCRUvHV6OjEz2x11U2
fAMTS0rZ0XmB/eC1Nb5BxWvV/MFq9S4A+LggEmyySj0DDrGItpeFSRZTYdSWlKeC
nFrO01muiIdtcASGEKwVkE8jhMryG+vQUXuDb2GY9Awg9rYe3K0rzBw3eeqdHeCC
5Mc1X6IGF+rZOCXY55P/QMbcE149B1OPkqwY8DV4HdVPXNqmThpkOkyjpXY5rCnA
befgRTDLQFGdbHwOcsDvERx/yNkttPrLpv4fb612HkO7rRh3MVaY5FtsBrmZIpIS
nwFYwV3vf2DfbMsEg0S7lp5rIeUZQa84ngTHU3ItaF1hi3tjwUJMGa/jSL5Z/Bw/
FdQDcpWf++YxoNF6qPIL4E61ILnymJhYRTAeEkK96HWerImEHoAFx/JbK6kSw710
6BCpj7Tfqmv36RYjxzTZsRaTUXnlX/f8JdbfynPgxkAu95idJhWOmKlat3arXwsu
/7IkwoFULRUhrGH62gFnmty3w3Kj9lA6NO9pa1YrF++0tEKyMVMf2/whnQ/qPs7Z
H7nN2pWo3YYNqIWIjVgfy6h4JKDrccGz8B0nvd0WWGf11prq0ynKBMV3xPoPTANX
39Ee2orp7x7EL7GJSHRBkvbqT2+tNiHIkW7VLHtMTy38saLM4Xa62IBf17sEKz19
3FLjVCShCHtl6nNO0S5g43o9KwWKMZqnrDmjcnP4ZEPKdUbiqD070vtEHZohQlyV
ulcDfa3ekm7Z0FRoD6xOgsApepPV412uJPFtWr+mmpEKI4Yy3T3uYLb4e1ZDg/4M
iH67tuRcz0g1WBKeZ7ezcsuLTJV7uW9mrC65P9+HGUb20VghXJjs+zmT7GZCQbez
0+wPFyrRJCDpQk43kNVjX6QQ3QsLgfsHie0+tjcAEjaJn+qOyCLn+5Z1EKYcyr1z
k1LKxy+CIslr2mgRKEhnns4gBQ9l4MDZ9EtosxM345RU7d7rNp8U1lOnagyNuqIF
lEPAdU/8YTDg3jlzUUw77ic8z1XODetSozu7siiF+qFYJ8MjbF12M8+5gQUvCQ2W
g1bAVXr7P8A4Pmb0f1D7jGsuUELdruB5A9WsNQUpArt6Akyf+x7jkj2a6KkijuQN
6EiZeEfjuaHuTwINo8BBo+pVczslN08S5vnEP4toQyhzRwDHGz95FkvFfiY9AxTW
9g08d453RRedkHX/OZyG0Hy1lnF4MZaQ2ZbTxs8+JQaucDWdYal4ZQQWoyeqNmax
669uzoo/+gHRX3+58h5TuLeFOg1SM2JCtvH8/7IQS5eWL3lR/awReTwqspNYm28X
bbC/IWaiBdS/Y9mFbToJs2gU6p4U+aX2ZWpp96SpjDNJL4pBt0ypug2TElrJV4kr
950SvjIT0zbVFRB2dy7ejMdc39bJBr9YxdC7GVe73fC4TG8JC1/3WyOhsDhf/11u
iYaDsuxao1LyCCeB4R93wMb4EdlNj3M2japx366i0QHF93nKUXNlWJVHcTEWglk+
zfUYs38dtCzwPz+ZozDODA2QPFdydtFRdgWIE7QAroS9i4KxFnhj16x7i9B2Vk22
mY3WiPdwQtASF1Hb/JrRNUV24oUQB49Kt0h15gNoY3uIIuur8l78AyXUGP/qZzZY
ZjKluru97B55G4+f1kx6qFKEe2Ze4WZlYAPtDesU4E4mAJ2P3MhncpIlb/K3V1rk
bmWFqWjwKYxIrPcnxok1XAt2cDstzsv/IL/9Uqg00lFNQyhbKe7Etns28U+LzuEz
btj1CCAsXo+2fy6RKclDj7nSxHQYyX66KZ/L32s8L+rdp9fCf6mFbc2CFYXWNrQK
ssIrtWCGXUsagmOuh8nQOf5R7eqALQ39Z+MFI8m9WPEpGVd4dg8JQtP+ypxiomsK
HzXyBPYoxGa5haeiogLruj6e7vfjdtCEWf5equC4VvIG99A2rdYS9HNM4ioEaQXo
+kha+cOAevsCtyVOK6CYmfCrSxY8INEYdc20COo9/KGAxuwaqxQSj6qYbNGOlbvF
EXEibguZQi6zQPlrUnv9/DVbr1CNdWD749ONsjO9QflZhtF/VDo0Kk55PbniYw/r
x473fFY+zl8KDQvtESIUm7W4NLBdBZ84UnYkLyjspnzsUFg7esgsziw8ejq0HW/k
KP3Z1hUtlkLVc7RMxDl1RmpdV9uDMzmZrMGX7Y6XeuBxHK1ZxGKwN8cEteXS8dPK
SwbBEi03yPCKuS6v9x8CPLKMU31d7nIMK8u/dtMXMyS8em5LYnxIO6EFFiCqPN/Q
VXHL5W5/cBSmKe2w8suAEFpIXvDZv/bcR1ZlDQI9zVCBFs+Wv0FuSIiarXXQxcoI
LPL3rzoVUfoStVVSMb3ekrQDWPWIYMwnFVA8FdQsfA4wqNDkPjTR0wCgae4RQoEt
BmvYuYxcmsEhAj3XO0CKoIgXGjGvAFzmhS+3c3FMo0b16udJz86WyXA1EU1F1KVC
X+MQNJ4O7KQDTbOJq+OFfdHlidgSi7gw9yT6LNHGTxlOTegySEDlqN7y6/jYS8Uh
LJrIkn23CTdgAd0658Xdx8Ib68XV2jsMdfcxRd6+RPTkYFuzu1wbdU3MX0lomKAK
Z85tHlvuBxMv+pe9LFMEW0w5Xw0hKEQEOE9r/zF4SJvhYt8dq4hXASqjcB/GuZ++
kUXW/oeD8ALvFN8wlIHgd5IhlwNgXDx/7S69mwvNfr8L3ULZ+wxiRuUBk6uI8dFA
5rNGW8+IUYr4u1XMmwPe+Ep6Qh9lPa5JdxMETQa5nn0aMYHi8Ga31Xb4DP/OFqAJ
iLjGYM+909xRCkinHdY98TkJXGSnwtXDVBF6S8BRc9mMYlHQ7Opuy6hgFo3upPQc
pwsfURud7r2paND3UzW74UNIOffdgdUuTIZQ16i+23B2Xv30YmlcQ9Dawax64p7O
ksxlPJoScryMV34lqXitOESb6vZFB1F78+qn+OfsSMiGwtsRMxEdhg6CwlaVtuhw
5Cd9/vxLQ8tuNKoAmV0nFBXor+BRk0ayPKcoJQLDESq/Q0ztjuQlTJmwuyjZg1IB
nc6mJnENMmQ5Hj5izrmZOEE6+SQij1mzCvUHz7Ikz2zmo1bI1LPpeHJSXRT40c+X
NWenqLD2e7eBefNkH5nuOwrgQ06fICtW+ka3Kl8tgptRoP+XKmlIi/SoQcJeQI1w
xSpg0LyVmcQLnAHFpYrrKxDta9tlkoCurBNOIh57py4nTsUoT+FPCPAPCnr73FgF
tW+xWaTDcGSXJCiDEZVT5UJI29rU52HKgEBbzk96MfHZd87vmE9HKetc/5Pe8Bjj
aknXFkJi8z+Td6w4TsmuxK5ltNWH6gOCG9Y3N0WDFXnr63yUElJufdy7YJDZbFtP
+N2MWkke3cH6KGghNuCkqhiBzpk0S3tavkOaJhmCVipIvzLN082RTfQ8tIcVlzMu
pcsyP7yKuOjlTlQyOyH3HN6ZzV1lQecj+B2FxsMzp0r4+MJvd+WVXfToHPAJyaeg
bP49QYxguhTFH8xZKysH+UQc3nmTmY8bVEdt8Kzq0qiH3jKmXNpzDzuT+WQ7vRMU
nisF2K2ASXKhJrTgLQGeVNpseyfM+Bp9lxS7gG5O1tAl/cpvAOxhOaWmv+B/Ro1r
O1h3AnvAtsFccECcynerBV4C+pMtYWzCnmHLPWS28oNbi5p73f/MRiISye8RXbnd
4QLzyMXHflzLoHELxnc3MAg+NZ5HnvtQjVNiwDlAOaVgVHg2kNjp9Y6YreHUx9Mr
SdCBzA00uUtZtosKt38vu2Aw+SxhvuGpmbAvpPKKdjgWDBwjbgMDod2HeAgORZWr
DrcKGk6pDbDoKf4tNPvlSZWKhv4SR9z4+XOUtslhZi1E/+MXzMEX+iN4FdXuU/EQ
Ij0GpqUdStt4xYqGM8VT0mWsxVgg3BEzXyVssnAu4+mu0h/mAXpm2ZW8HpeUobT6
HtzMHcQb8YBYq9N/s2e2CsthOOycEb/O2S89TGWqPzrhHo6PKgI0dM3lh152OplS
FJor4X+NMpUjvGSnWzySbgG+X/ePZyZvBZgSgrr62itvlO5/vHDOpXmkAr87W5fR
BFrXH55ae+hG8C2C0iriSwpiICDBtn1ejW4FOwsBwUtx6TVkTn8XQGduxzptjgHz
yuSimCKORP+7/Elihh0y/lMw1oM18DII6aefhorYbLMywPakX+KHa2oB5dH7W7Zp
wkVncV9Nqre2ze/KKWJPLEcVJHtBfXsp4sRoPDTCPg1sQNgEfyaHplONeHezHxq4
FnS4JwFXOAeBICER6skXL5P1K4mAuIsqQ1n+vDy62espHqFOauSRh0sMVy0AU2kb
S8acnCMDClC2r+WNavg+ylz178IPK1k/5Bcrzq29gsOWn4AZjFzcUjR349+i/dsR
lmmdbxHEi5lvAihrvq+bSlUxOyCkiVWf/J9FyqbisoXXQaZgLXW/1XPRSS75zHFm
ieEQ5IqzPpXQW8mepd2ItUDaP1mLD4Rl/imJ489Cewxx7c9t4RhQylwUhCPAy9Zv
M/Ly4feMLi1lQe0r7LxHTT1OOjNzRZdt4jlDvUS3+HmJ1nmo+bssWKWFTDfEKvSH
nPDgEa23pPDKKwpYiMS9o9/IMkHHu+/kX4obVsL5njsniH/9GiOGjd7B93PbFW10
RbRSLtLAeKb0FJd2x5IurypUPf90bnnPu7vcUu/p1bspXb0wBFM1qzOFprV6TiNe
8nGCrDM8uDfEnWIz9icnBrIdVHYMaeX5GyHXaPFr6vwZ95h94wCXlSCjYcGUc/tr
/MliMJty0U02CRlws2Lx2zQWu1V4d5Ue3oAN4YvjU1bekivU5FYP+fYeuv8ql9js
n5tRynNG6wEgmRbHCN50Y63d33oc7g+DTrRYfyQOogF6PvuXdxuKYlYOWc/gDSSj
QFuUUxYbUs0/S8+PvdEy6FOy/+twFGOudTX08xbRmaLFswdsQVHINf4rGf6qp7XB
xhWgBB0+Jq8ShOe7uB5OGToP46UwrgcMdGriJIxunoVywJC6iioU+1QIuKylOHRi
FsrMqlwhG8FDQqepkqooSGaRcc1v5QJbC9btEnlCpadTGdbeeYOL4I4Zbq1I9zwt
SEQXWDhF7LTfUgNwryNbOoWaHdXaYhob8a5KVRGxT+ZX1WkzICz2A39qzZf93hqf
m4URvxFlQufxTjyFlZpGqsqq69BzeDcfiJcY0PSUbZoDHx6W+zAOknrJMoKgg/hC
yuBlpS8SJ67SA7N+WCpbNmFYjjob5dPNXHWoVG9zjavO2He39OWsxoYRR2jJCrvD
tHvB1h52iK/g7lgqa1O0yuWNIv3rWhuYj4QCQaIjYVr/YBhSGKBPTSLacwiymK3A
YQJ57Sb8lMSGjvJeZcJVDRmWiV0CFZpnDZRE/jM8mgqRyG7zPZe4ppESPEUzTFFi
E+lC6VWUmcqFMVG2DejPOG7BeQ2Fcb4+D7/kM/bVxshlgn4T93jbAPcB5oe2Nr1/
/azAJ9tII3NTUQAxnnhTKFTJbDDFFEBee/HsTggKVpfYMzsoAzaVvioB/2RqvvLm
mp8qPLr5NSvQ+ZiUP0UE3X1l2Bsf8gU+iuH/GSCJ1arko8qsk8iS06U9iZlqpXnJ
+7FHCb+kg2WpJI5mxZyXHcDve03HJ2tu/x9tPiy/iypq/uaKGLrbPR4sBmPveSFJ
hswwgEy9jzHkynjSWudXpLUutc8GncyY5NOnPUdOfz99DL+UtQ9bHXBzckhKltjb
CCRwhPQeK7jcAzYt63pklZAW/JkOWlz+mwsPP8CvTctcjhOFlHv8IEh6nGjhRDEd
janAnzxXk+KFtfzsd7dDd9oO6jfkRVZH580XvkIFHCtVZAAoNVwIdigkbD0JmBaf
3TO+JD/CGqMQOm+S3ylYggiBSJeEOpFN5KRWWdd7XdRzhUIr1Wc2L9h/p/moiVw0
h/h8eAjRzjpJq1IE95XnJex25iMNCUI95nWFdokXWaM7ys2SpBXkww4o8V+D3ctP
S56TFjUARR1Usuf5eqcLq8Z3/IK0A0ti0pOUTsWlmqOBew0jQeupR39l0rmGAO5h
eq1515NRKSI1Oj2ipIRo1Thbl/T/u9qouZp/nn0WY3HLjS69oPI5XwVhbUqsaapd
Pa3RO7CN51m/+ZSVFEMQXhUx0I9g+b63ODOgiHZKorXg1oI3ueaMCw/kttNyV2/j
zgoz77TowX+MHXVVjGAgTqmJTCQcewMosWeQIzGQMNxsLknWGTXmQOrYPKiFFgS8
lNuLohHLVHWQauS0WDTcG2jJkuI3D5Gj7XMIZhzxEHD47vOwWA3rud8ay80A/JyZ
EvU4Q59tHRxH0AO08f9uBrdu15DQrYpMgcF2wX8lEFqtDuDQ6/du1ujHhoLHOA4h
hDsXP3zZjC0sGA0dhskUyAP/hh8CI4ULH1D0tLyymglan5iaM1eVJ+yVo9O5CX4t
OgoRXg0EcHSyELmNPQOXcvQTyuMnfGVlkcP+SwgJywhafekI0D1OIbkJAOxnMiCJ
2j4RyMxxfLtLqM6q0sItlgOwNsBh7T+baGvbQUJcqFMCYfh8FKwVWSpBrpwNiOSK
T9wFaF/i4kraWH3EhRsT7KrAF8PIn88HqaeycTSLk2NmSKBy+QnsbXV/9X2nxLXT
zC0Jd8wSxRaIy2qGASOrxdbFb0hclQNB4aHLl+SxAS/iwPDhdcZWfQUldW7f4k0H
9ctbRQwcNAh1jFqdHpSpK7dZtpNlu5WJWHdF7da8IIeZDMfi1KkLCi5o6/yln8G4
juU3ZH9BRs7DL09xR0OnSjQSmj3FZCIzcIqeuCYaSdaICRpozpjw7fIIjnuH0u2u
T3qOKyM39W73fpKNQGYGgeDvEQwNlaRllttqgXY8kQPXVldwLMCG1V9XZIf8c4xC
aZi6Q54UaFXNILbq2uyiw95YHgMtinXG9xXZ4khGwKlWnTenlRt+nXVdApHP4WZd
HmHK5VPpA5XxiWSw/ncVu+ruZUiW4D/L6kJnCW4unCx7F/ypsh56jJ1nkGCpFq4Z
jl1i2Is8DCes4EJqnlIzaR5oiy/T804rwQHbHY9FUI2SBPRnSJzMkkIlPsQOSsv6
dLoPv7yqjtgABfbt0aHOefc1UGtRksyh327+MymURGRj1aiAB3gTuNdy8L8JoCY+
Arr1WXiEQMi+hnPBXT0tlTxYgPQpSpR3O0T8UWxJIrN0ixmln51XyLA7XhydAKJ6
9UzdysLNMw6QdpVMGtUI+OFM021UIXExHtKx5bVlBmFayyYg1PaearzhIs8IPzM3
DCJJyfZsEvzLCSRzFNZh75qkVYnHYUHSvCEFl1XQ1/zCA9weov/2xiF+jGosku12
rcuaQWYcNB1IBPJqrJ7M/v3RLndnM5lDIp/hR3s3tnbpDqlZi1jIdRGtmmIMAWXE
JSAF+jhsm1PzjGGHkE6eCbVbPkq/DI0Zjb3Hy48GhK9WqG4GxCAASc4NcVg+Vxrc
lJONyWJNPRTJuVN209zKW5m7b/or9UL8lFoBlNJH41E7oMs25xx7sdkIEQzAxgOl
BB8OQoTvjY1zjS+E73t8Fi46FLbnBqiEXvhfV1ZmDPGmSRF0d+12cGOif3cFR/LE
OfGkVZCug8aYr3whFudXxXCD591QSYVayVdbN4mEcGwU+eCIKiIEIEBwE7AP/nr8
1Mz1g6bZD+8oTwZAi7X5kuRko8gScfhRrJ4c9iY+26zDbjjiKQCnd9qtTkfdt66F
5jvyrxVU7UxomGqqqtROUmCm7PPFu7vKkUFKUz8b5jpiCCRlHy//b0GqqARCKYh0
Eecn2I4kdBxth7NA/q7KftgQD1ah3q3WN94vpusZBsCC9XtNOzb6wxgsgDDnUKuU
ZQ4FIpG6T0/6dya5bPQ+dpO6L8B28qney7Tu45CBXR1I4impPGMbInzVJYYXLWiU
anureETD12xv1YUDBcembkUVzxTTa1Txew2NWu2iW6Dw2YrTojj/Cw4CFQY7n0R4
1TBTKNph8PnNtkXt6ZmqrSJNU+XDBa0VjNUXOsxSR3JWd3LWQwHRxBLDOknsNZTY
VU1TLdZUOu+aJ6Uv6y4tC4Grn6cPYUljbioK3tBOXBy3zJhSMue+lHVPLIF1dOQj
pNExQMk110FcfKTPKZdrbvxt+PaCECLlKk4QCoi310a4Uf0uD9bxK4GuBZCdO2Fl
fYl/ANlP1m8nc+KXXNKO7ajenEZYLlLhwx4kAD+eIdhlbvrSm7vBp7Zg3I6tDX0J
bBFXjmoBAmOQkIo9R3fpWNK5MQi8QY/aUWERB2rSeTGSGnCC9JYihvwnKfMOCjef
TCn6Axt6t4onY178RiyG2k/PD3J4Np0WSQAL6kB/VtzAWbGpMRgFkoZ19QWUn5jl
RKGB5hgQHAJHTmkNye5G6s9K5U7J0py/Zq1LfnugrFyp8rNehM4X2gmZovkorRo/
HqDxsCRgRB5ybFgsF8AQtlpFhG5c+YEOkdyqqLzupjG4eBSON9Ks+D7UVnc4iZlN
SAmRY9k4KbMqYU3XDVt/R/qI0t/wDc8qzsaIEW2iH+6u5PdN/Y3I6yTbeFRUqTHc
ODvDfMZwEQAmDh5dOCXyQjhMFaZhCvc/5eXn/ZG81SUIMZGu5YZ2120Q4zt+c5cP
ywHMYJeo6r40Hq4xcU3g7kzwns+qGZ9v2/XllTHdNHZI8ovhGG7lgQSTsJR3KAY4
1iMnB6RcUk7ezmner8VC/2GlJsHJKjxDSHAqjNOEdG63oqhS/pDgn7m1NLeOc1lG
fIP607QOh3e546V7FoaqnVCTX/LaLI1rbarjK7spxCEC+gyRBn5xE8sgS41L5/as
K8DODg8HqEvG1T0qy65NMQi/nEhLa9IuvF8cpuBzNcwnVfvvbCDWRtxaAqJaYjLk
HJsfzWZzeEPGBxybU4mFKbuMplO0HdjIg5KI6BEJQWl/s308XbmstwUJaa7fK1Uc
mjqfkR7lgsFE5+jtOk5kbFGhD0HMma0NJ63jOuRILU9DFfoaOPND/pV+YP2162e6
7jsLYS1aH1+aK4JJ4MXzzOXc8tPrz9Fz2G+WPSMUn7y7uIEkITzp4bPXIBDLu36g
UBu0Qa5pBjed7caTwkRXfH7ay8ckV+zViQ0ngKPaPDn7WhMgPElrQrOozKPGvldy
J/xMg+ZSUO66ANeLBwytFC+G5GYCkXjOeW7PXIFlHKAAMDzdE0c2tN0TdwEka8/F
9OwLePvwXcRokycZWseTXJGGhL/PS0zOv2jeyR62VBwwSwiOz2dp/3eA/1hHdzy1
oF7bbp4rdOeUhtr6IH7qq+xBIziLvGYLq/Jj0xuCMFrlMZKMuXqPusmX62J9ZsJ1
+pvqo906l+FqrxHfbzqRQXTpKdlcyotpbENILkUaxxiXByECwTgnyNAxE+5+KSV9
l/ikbzEuJ6DlAWlHiPmyzuZuql57ZY3BXqTx9CDGsmXIn4M0LgNJ4p+Bkwik91pm
nFGZLW+myZximG/ODmgwA33yrs2pqJPqd7ghYlwdedPMmnM2RvYjwyTewO6vwMm6
S/sfNOKpSDz0uVjLS/1+3GESFi4RrXqI+5GLMNLz6tDHdQaVbGHqbVwVVx5+O+lh
1+E4con7LPPjDZOwTai1Hug9nloYIJE0bQBf5DCkU9MpJlqF+8MXEKi7OhfpiyYp
3mGhaK8VHzeoaMGcb1BMPWPjQbRIp9I5WLWRrie8Ek7ETtFRVY/r+GPf87UOQ/Us
iOVrfgqAnbqUvVR4w9i2K8NQ1690TdlpZ6hp9B/yb193Kb8koJAby/SGq02dBypm
UBxVARFRNmgTzgxHauGMOxNVI1A53z2xZefhQ+N8ni4N5nbqqEdeZdysA84+Xwoc
4qmbILznr4n8pS6g+ezAKM795jjlJttkhbx/yi5DPtY/rF1ZRYJrRLC+PCDNajKm
IwCnUjfXE4wBkWlzftUkBVTNgHx6PXGk0RFFcSKcfU+yz7uBRye2xD6aNao+zRvP
GDDcb/En8PRZSNayUqXw6NgOG8ABWnV4U/Q0KKpntYxSlcyUggrxUXmfSOpL7h4A
tXwrhAcSEOXCxCsz5XZ8wiKfOl3sr+EW+nPiwVQL2hmEeTC0gZsnXIKIaug/TWYq
BVA5Q6MHz+QTAe1i/Ih9yAz6M5Riar1sYBFK/0vOpRVBPd/ehLGlkjdzr+Dk2FDB
YlM/l93AF579hjUmqTMgZYLdb7WoviHFVHgLtGLJJtZn2AwQIci7R9yY2GljvrvH
CTM2lT9nu+Qj2imCXCw7kcGEPrhdaRIUoMiNFExslJyaVnV2Ug3M3Dfr2QVOJKM+
+yYemTSMCODpYe9iZu8VPS697rfjokOlvF+aIBRud5Amc4CY6N1as3rHi48EOObo
KBX7pahDTN0WpdNzutPSvUFcU/kF64E3xA71GjtWpKSMZyua5KFg5TBgL16f6loZ
wiwbmknpI1+40PJlhxxCzmRw8fueyoqA9TejrN8PcQmEFlykMXJxg4gwN6VyiKR4
QjRtwriBDo09HRDQBC4KQw6FN3w2M7dh355mMglLReDZq69oBlek4XTMX743DldH
hfjFFJOVn2T4Q1S7CarporKdZ1DNubpqO6dJAg7yg+zHOuNBNfeUF/jAKTcZC3e/
7Fz6oMNVHc3lMkjJv0KFVAmUz8gCvwaJMRmzBK+Z4YmwuFXxiaE2p8U+LVOkexFH
J/VWCUiUf4u+PXxpbZ9UbyIy2isAFI6mhD9rd8mddo+Jm2PG+U0sv+ZeIf3eZjqy
KyMjdgpI4VOJBocNfvgnSiPj74CnrlzplYlENTiZcVuiwCaGUr60x4dnWipDrDHi
OIoKgQCL5IaEcX2E2Z6vtX2/v0I1HbPyPiWVTS2QkoID3yfPW/SJRoH1fEvKCQiq
TylS5NpJ+92H32M53YCoC7GSDfoQEL+bli2/A/qbgzzEFsmpfCSh2sx0PehlTV1J
Lo3iYuJE7++Zam5OGlIpIMEwRlK4tGEx78H52ZJdniM4no0p9olPIb3YalEEvrMJ
X7Qj+reGKvZRKLfKcLUYnDtfPnDVG1lZ1JdHsG3zdUWK5kcdGc+84yxWUzoik4Sp
OdWiqsLoFgeGAe/w3haZ4AVBgNUSL86Cifah5ymDQA+/MFT8lKE/Zdl2RaTH+9kS
5NJ8ge9c3OFyvaFJ8bbRwXgc/TvvqRwsl27hYMtMubs36IloFlY3UDGhFFs20d7i
6lGBSg1hFWAeOC6CKGWDOIgP3+VPEYutPMvK9U1x7Zng6r/mV/5rfLLcrNBzEMMp
+tvtZiDYs+2saDghxFvKma7u5350mecaOTVzgecSCOpGe84PbH2Yn5DMnHKJF4LY
d6nzzdorg7TmE/kJ1rcBGRIeRnv1v9Oqfexm2CVwG4aFp/o3TkOcGpftB6ln5rIT
jMIQHrK26HSHvitVyz60ioPXjnLNcjsSwUXb8kKC2zMEMGAzvK4d1rY5JzX9W/e0
UDdI3+BFungmUk+0Ow5I3Gxu6GAuOGbmHOsBn73KV2Lu/OtlGOMrodcjnU6hjdQ5
7FPgbeaWyYkYTl5VeeRbYSydIIeAIdqrFopvZEhzGU4Y1AoKuC+W+76xvNhdRI2e
kBtdgdfBqiJSuZjzYLO2XB51uejkX51MPtAIpojKcCLs7SYhmoDYGQhWTVqIpdvU
HbLJbGlEuB8MHJEdOfd8T1e0/xcvsklUVYKSjI0AVlpJybjGiQS3qCS0tBv2exFr
+AIwkdCETNs7YYlOZOc1mTTwoBIDIgKPgjm18zFDBj2dBU8b6MgDwU7yn5LbXHu9
6ZKYhZdLrS7tAaw4UV//V5VAV94tM9f3Z9nU2mQQwrvJxeahD1GqnNDyP4PxNTgO
hfK7a3UDfeahxOe4l9EQ9zULOBsSga5ylT15xTh5VHstrLrhLOxZHjdd2j8lWAX+
Ddwln/EtC45T/GSEkkED2KM0ubamnt6BKrbG/ToelM/TBYH1vr85L17XRh21AR03
+n8PNBROZ0nq124f+z6VE9mAJemZ08NaJ+BeRTshCL6b/N57C6ngv9evpyFMX51Q
LVnxAkcb55J2ltO8Xe4dg9jbYe8cxIMjhf/7zBySo4TZxgpW534GGdg/FxqObCOT
YM5wiq3nvYHeWaD77eBm/WneCIhjG7qIYrFsH4NPwtGR7tlLWg4Y5DREOXKZfVKz
uCNq6wcRzqXg2ECLZWRQtrHAcizXrVtHOYLh4dFvtnBwGZ+GXHOpYO8oUMBcvpKW
cx3+3uib0jdpeXadvEGyLIwEpvYImv8+G0M7MMSmuj7rCZ55ZkTot9GjBqSznyxn
u5BT7I6htPeQm1PbSDC3E+z/8pwAlUZRf6rkV/Sz6JDoutB0apeerB/9Vrr0bv01
Y6bu37xXKixYE6KxrCEgsi9WJxwquPkZzn07x7Mh4VKSQVAyiZiQNqQ4qDeDMhIX
c/3kQ+6MRW1I5n75nCIRKcubKECPBW4NINGpFn9sTSRhYPe9FI2naqaRaTbvbind
fs82DKAgbDvQmR2dAuZCKmGVRPGypsRf8WvOuhf6P6nv/djfkJYVerDwKzYIsB1b
soUJzE1VyAG7vGRc/lMA+87/hNO8kXVkesl/vIcY+6++x98O1HiaxpzgyMxYDkvn
eHa+wdMB04vPU26qg4kq3I/xEiTVT6Ii6zsOrpY838MYMjtdH5qDNh0p+Vd7cVGG
6cdEDXwSZSd41kI+AkQX9AJe1/RXfaaMlRuRV3+Gp2AOdk6ku2u/FZGsJmungHC6
SMFnTcq2OSd+Lxfw/hYJz2/6Op5j1sDkjWxnaFFtDiQf6/b17rK153LCx/sf3DKJ
WxJhBwluecAOb6trgeTaOc5jbNfreLjCyVSPFGlkadIjFouju4okPe5HFZ8uW6p6
NtrKOMlBNvboRumVjM97uXNNF+Vn9j5j86iqRVW91g1Zu6uFMz3ZAl/3hbcIrD+t
01Q8yojVUVfMDVKTve6rWoM+7pYYSHDoWmiq7QTsBBjtLaCjRUTuqj217E1Y9Pn6
qe4ireezfvFZepuQPHyNkR2ngJzLm93zWnSBpWWIEWRD1wGJWRb/lpoHKKGGjziw
a58s0QiYkZEX/dXMB84+VqdVBjRC9EU/1Bx4t4VIdGcdMG0IjaxSEb75wf6nNtq1
J7kTlzwY2C8HXmEDJFv3PSryPKAbYcJ4t0DVskwJxZcOPfIROUHVSHlueBv2Y81j
fLSQ4Rq3hLz+MWX08KHdi40Ref64JMiuBGxyglQ0f4DGB3Xqx4g55ihjgS0GSNDC
2IsgNKI+qKd8yZmXmCP4TMhUDfc27Gxkx5Q4xHIGUa3BG/vErThTU6agZniHeOex
asSeyZc71yNSSXbNpr2HbtQQ3jpkYzaVkhJkx+Ss10Y4hAMNVM1ga8/5rjoVi4ub
oNaqNEC17wWE4Atw7v+CJ2elMZx8k8YA7JIMrA2LfR1dfWqhiLnRr+VSDpNgmykB
ZiPeB8BUtjSpDTxmwPDBBXtFHYl9KdwltMG+VCmyo6p3p3Yqb9MSUcsZ6fPqgIsW
BEGUuF9HbI8m7Jk+Lfv80mtKt59Vl4twVJE0w9r/xOxmulGtEAYKOAKSvswrhXsW
SLI9uevXIISnqXt6Qt4gqd1ciHkpcEcEBzbUKDXd1hdORzHz/sK0f+TJx2vmDZzA
XwQKckjOml5euAL0xLZBJCs60PtiJ7jBZ9m5Gej1k6xzQ+2tgLtSJuXJgSqXzYnR
tELY+AnfhqYYi/SgAt900b9w0CP7aexwkY8LDyvGlcVHVkHKp8yxSccadPsmPaI8
rO9J4NkipbAWG1YohxX5evyBdOEk2u6E8zOCGg/RSKBh23ThNmfEI7ME4tVArQkB
AwqTlJmeKXC8fkQywGnYOTNuHCQd+v2sjrJIQ7+XVgOYAh/6KCNbhhHW8TBUJl1N
3coSUYqIxJeZ3n7R94OO4Bh5C78DA/ckMkh39G3P9hnLGuc2gRUQUmQml31qp+1y
dugG7CGRXuAx12y3WF1MX29iBzCdv00/klWrtnZvbvI0Juq23IgOmmpHBe4/RYLi
e8wq0kKIiPC9BFfQtEtHOcuaoNw8b4KSUTWW6y5fueWOF1fBOezLkG3DGSecAt8H
6aE/3cxHUxV/eHPwrFFuNCMM1ia3JMjMK1/WARXvIrNU5hiuKL80E4tjdkhRaJ3e
ctWl423jXletpS8T3+ALrRv0vaPIqnhyFLEQFFkgbCSrnubDNfloxo1leqGn7x92
SRjk1wTbQ85teRsjLdgH4UIM71T5j1iqDCW3918ZHZ+MW5w4ZgQ2s8EUp6LkBgut
6ut8o1sLWtAa+qHhdStd9lv4e2jMbkD7hQPIgQdXZelTtK6Q/5XULoN7U5ZCfo+t
g7qwM9PiZ1OgtMgFCQTnlYDi3KgCTCorHURHYCvJuGTLJXA1ApmOWv7khtlF2ft8
AotNHDgvNP/Yjgj4HAMgOF0xEKGklQkcZir4RwUf8PR0bOOlSQwwZqto+zdkljbH
NtmmEhkukj4ykwS1Cok6ODYD8y9+EKWVZzSvPLBIJdFis+CRwGmk5z1pvsz8KVE0
u9B+i0URf+XrbRyACo+gFps9UqxGdacYS1djFFuO8G59hA2TbGjXBaD+ThKpVag2
vPKr+xLpn4t3glIyfTKnSeigbhLunt40/Rw0xkrHwrKWABtyaGE+Le8uiZpGk6OU
BKGMjlyyrl9jNOtDqNtr2zTmIrKbehcIGAFqFpHlUgrQBcqXXdxARRfOxBTrH6Bj
Dcvep/zscWd+ZYY8t3q7p7m7j0P8MY9lFkbeafZIZ/Xu0MfmqjnK6X1eGC2YRh5g
AhROEJQReEBjNP9kOz1/cvAsKjgthj9va9UOiBTjcDdwta6DsyzSzXihgH3t7WLd
ocBZmK70S6KH/1yaQUEF8cSj7riRwlD2RT4Gfo8fpF40krDv6N5MjI3ucMPt1L95
vutdj3N32bs1hjBMrqkCCobEXf7/k9e/jkKsWOgJx534vf6ap3zdYT2ngAeisc+2
vpmDGVJWJxV1TgpoUHmBOv93JMUxIwn4okO+xmU54QNN77XittDvg8Dj93E6XaaB
WQOUh6zHaao6uVG5ogO7xfYztHVR451Q1SX1O2x94stZfdUe1bXhYVjnNmuZ7/OC
Yo1Afq7Yfdc0CesCb/ktzrL7F5UcN8WWjiOFauuJFqoqx1sqCI1uSy5aS++Mhg4w
txveqmSmt6U0NsiRTM0zLeWXmlVhkhjOabZNOg+uf4dALytrM6aBYDAmsYAtt2RS
HTl3W2WJZrfoJx/yESNmCGx+7mPOayrsKYNbES1BzOp9EcCYq1Q+Rxz2h8T2xklm
ns3UWg+GY/hF5DgnPyWnudKbM9XjzUy4VmgzIHFTxR2cuIdQa6sH4VGxZBS+a8un
JBgHA+2RZ6KnGtrUY2tQuTylzaBJszH1ByxpL0E98itbtBahSUNfBPotkymi3Bcg
gTt1yUi9GpoCJFz/tRZ7Bni3RF/cthID9sUbj9KekC4N0E82e/R10JiQ1OlZNpzg
8o/mFYRi/nLsIqarcpyMOTX2KxMAUqO8CtOQafGNKnvG9lLHJOgwma0r6zjEVOMC
rzT7wpVi+t5kRWGLjzJwgm4JKb1C1Jy+o4FkiU5lX3WcV4l8HbZWRvUAUIAWj5IW
doNYJVht9uh3HFM5QRVAPAFe5MXFjWRXU40yfbvFHoDDfqynLnleATWOo+rmbA3J
bllm1fT1nlsHJjYrq5Z510Mt/9NeqrhZ/CfXKyDv0UokTQcr2kgteExdaVbuSCK7
ogP13nPcibelkyZDnfBjlbXqwCiMLTCqM0r7R8RWYC76Ev3BfhnjUYWaGiMMwieA
85BCnKGDVA4ZU3XJxXgCxrXPxUcnwF6u1cA5clcOmYg83GFelD8OD2bKA1cJRvVj
UALdTWHnFDJ0ypKyMNH6toAQcbaF0A2qbCH+L3mLRv922P7AUd8v40OBf8UuqFBk
N/Po9og7oscmMZHZjZsgHZS47b4vWCAQhA9OoS4OmizW79PclhiPdGY+EzMp1NAy
fQiYMx7yV8JLuwW71jVIyd8V4MHSBAp3JrFH0OfoD8PzCUDPHCtYaZ2o+zcUp1A5
ly6mztIbbIivil/joY6OLkprWXuhXkER22VHasiITXVyP+6bfZdx1nnXzuxfM2bu
PREfBleS64xVKecZ2IHdkJZamholiq6tgbFAOV1duE0W6HZ4BpeOgzqKZossdS5i
/J9e4qkgujpu9DVvItd9aWVsU7uOHg7mitY4d0Z5Rtg84reC6VzX4LUrP2+valXU
Q8yHtx8v5+Ipfwej8JbzdBKQ7RD3hdbAyKAUqH3lvotIZ/raElJF6HS/uA2CvOOJ
WeUg8sLJnR32MbyBxOtXMbSYT23w/OhaEDvbMy8gGuJWxf9lm/9Nw315Um3/0lU9
5Nh3bExvNKG5tmcPw8f2E1LxMn6hPv/GNDDxiP9N0gYH5egtnjqH7n4Dawc7CRkj
4R8S2d5osc40m4G21TNKqpea0E1+uI0bT+tTosO6WDkfaBT+FUV88SDYOVX7WuLU
XUFnyDnoVIRv9Im2OYVoska9MekV4+EKWe/z2wSdKdxJpvg3ubO18L2LWEkwmoq1
7eOd8VTVgl2e9sgnxH6FD7QqeLcs5hmDnjCR2ktbL2uLeuQ5n0Oz+QVeBL8I2R5C
IZfu8paAitYSZORTzH3suy5HhFuelWc4DXFvCir++CTq/KHh/luwxc+5bSGQDVk0
/l3CzdKRqvCo0TUc71TYzzl2Hab6VuN8KQicAzceWO5MxCmIg3g8O/ZbBZFee1zt
u7FYicB4YLGxWZdiyN67xEQNwiQRcHL9yR82koCZXu9/Cz4Erlmg9g+ig9f0cP7v
COZ/Cg9exr0+JJUL+nmPjCrR6KqAplc3uq095t0Mkqf/OUG8sKRdwqO2GMY5+KKi
0ZxNTVo8WlPxYHGVWeOtWuY4HdNQCgAeFhJTDDzwQggBgTPKowK9xXSswAfj+2Gy
n3huLdZZrNke+LLwAQVAcQ/8pQme538l6sPEL0RlqO8D6fZdJfk/WprsvyQbB4Zo
Q+cKpXGxqmZUMZxNZoeSQ916lGes3vEEElnnYdeDm6/biK2XIGiy10MSfB4hE4zM
GSv98aQ+xFSU39Zah2CKutVnvWNV+pFgrVKoAcCKStAxRIHe4ZgI5w0o3f7MlYK0
sgB1w22PTQKRhkkRDhu8+cwgV7u0CiN0bLKcs3po1j//znXvfVDB4CnDo7h3ri89
tJrIccrnpnU1qrHM4RyuSMX1WO5lvj+my4fmnQWJyuHIZjOHq1WjkrISrtvlz2jN
GmOY3tYH92rRsvfwxz2d1e3KV3NQMccGnOpP3QgOf1DZAVz5Kt9U1WIe0OzQpVtV
yP64tWjnXo3iOVP6gH951gDLwHuXSedTCtIPzjgdMkcoaVmjw3T6Zg8Bg3ACSzWi
zoFeUL8Oo4GzTVKI7nRomn+XTH/CxxzsakCWOSLW/biZ8unonJF+05obFlohtk8P
cIBIsHwIJ6MZatU95galSCpwuzq+APLDjgr0X2qRxulzasSbEu523OwHp+eRQ0U8
+h1Y2ylNNHS2OXxykg46j986+Yvkg7PxlD1JTYnA7AwVpz3gZ29xLv7kk5AG1Pwz
iP6iEbYrOIqNBf978efFejM4QgYqUPXWwGiIWNqFC5n3wA09nldlxjQUd/FS0Fl9
nq3FwgGX4UATsmvLDHCqKpiRa9JgkTK1OEzGEK3H5sxNtIzl+etJgy/mFa9ShsCr
jsxo+4OfblD1pTnvK1tZ0+0ljd3gEUw/Td+sFY551a78AIwJQys9+hJIQyyoiik/
0m1MKk14e94ca6Ni8EqjQj8r3oLQs6q4aJSGpxier2GQ8qx7JQCAfBrRAUhlANP1
Vu8Ap4Rs3VkmxeZYjrbV8GXDaLlTMvmXYzCqySk3fNeDdswOXDq1iEeUZ2+YNV6R
a8qcF60rzVyItPTnTzFGDGlxYQax+4jtYKSXm4pGw7qF0UnLSrdodVrF9xtrR9Om
f54FPdLv5oOeBXicGuYv9/vFTR1Vp9CURbhuDl+DUoX82Ic9VMtuk85vOCJqqG3Q
XfUstu3RW2rIG4xHRkOZcgtffDPmrD5aP8X1gz/PhF01Qs43sVy3N0wWQV/gCBm7
lmW384QDOgKyPMEK1KPYK6j2UnIWzg8arkZTdhiCA29VSCiyi0e2UAAF/pzzcvax
OtJNtrxHnrlzvclxLRP9UPYwt6BBPDonDS+7wFInt6crsjsgPtkvK9cN7F9r7gyD
t5DZ8PMXAfBLk0wDCCFlrAn928M3eB6iKQEmv8gM+ZiMz4gWakuLi9OqUvgoorlh
RoXfMTi9Aq8UJy8JKYW/U/cr7YXSEEM3ilHVXnqe/Q3Lj3UDkRoW0aBSqoIr5Jsg
dzI/QVCmKbAzt3O7eyQWMYoEqqcmz7pQ4YfXMMIXFNE728HCg+yuXer+HKErSE1q
Nsvpkss75NqpbiZzqmemL41a4dim8D+4pfibO5dkO4121NaR/9eD/6FY0FDJzA94
2+7wF6pC2OVzM6QgM3hSSiYsyAAX5GtSxepiX+w96V/uoZ4i6WvYrk6f0oT5tLbq
TYMrKQDFwnJybCgIPkaNVDHq26WiWA8W3BpGo5StCmINS87HPSQwir4S2qXiRhQS
HWFdyHawjgIqgTivADvl06PrwBGjV3yLNasYNElQUaxUB1VfgWaWi+13W5Ls1hU/
AOj0Do3S0ybhfSs1Jwada4zYKMDudnoOmjgZX42YA5FH4L/jS+QCIZT8WDQgsF5i
7/1mrRkwom1OxAIH4XiniRdKlfjzn+GR3/icP4L7p8SaBY6V1cn/ILO63nYyDyrP
H315eE7Dgf11FojkKm5+raLKIih/5QVk7G+AeopWWDRU3zjJsezC0Cdv8NrABG+e
kHCCHEAQ3E5Rq4nEe1Vncx3rDfmdN0zymTCqh9h1lyZcIadGfmCdKkzz67rJDCbE
TKVO5N9aBLiB/L705mCha7eNvZ+IbEFCqyE/PX1AEreZ+MDgfVxZV3hSDZ+mLTFa
1shAnOi/mVKUaGgPzllAO/CgVEoN5ym/0RTTJrqbd8ilVaK8JxxdNIBohBG6bnmR
0fgw9nkaEQOdLixx94dk11BdHU9BeS9hfMxdI42ViEqihmgaKKWrKqGd4qk7Fuu6
YSJKipbpLlyn2hLLyM/qhe0/Y9rVluquBvhxLZgB14w2GF1NKC9GRTdIzfhE+WZB
yU1dbx6LmhsUmoCtG35HLXyGmdEBDYu7zUCcwKckwxWGWHgjlANQGGDnfo2T0U6B
zXZkAC8DGNNjyqu7yJUlmETsSnBwVntEivWeG9+8cju3pD78ggjYLlxNBX4cl8TH
/68EtKQXbZtPDoRVWwXJ0ptw676LpMSLbAz2oA61jWGDCnglOGXFUMmGma0Vmhen
aaOv2r2pHXPeUy/PzPjR588v1W2H6w3pEToHTW5XIB1fdTgHCfEHpmBq/DKtgJ5N
9CKckgaRxAEdqsA8gg4zTaHKt/aAr+ZaX3lxl9aGpZUjWLqPE+o/78xL9U7L6hWe
z8sl3f7D1m/QKMjxBQz2nj9PC7yAwBAEr19Q26Qgljqf8pnULrrR4+o/LsoFJT4R
tjue2xs4wyT5rE7U2l48vUnMtsGbOyHQt0OnhjvSzSrBWHM1Qn8y5DT3TWjdsIDe
dnhyhcWq+m7MHm4HGoQS9TsEq+liZL52z9nqgcu6StOsOplF/qjJGGPqqj4ks3mI
HOX8GDBfu34RAeASbXC6cwUkTOI4vv0DOKBUoS3p2XgNrPvrOMSo/i839HpVRt9u
kbrRgNu650cb1+cn5GeMG7M+irGIWTndsTmYIPYGjVyMMVbvDGdhK+HG2bHTpLw5
nzZD2YA3/htYRDmVaNrzu7gQJBxMPg1MviYhvmOz1nj/QYxVGGMir6EgtlRwN9cb
CFDTws4etUYauWearevt0af5xENxRQAv8hMGYhiY7Z4Je/xQq4WMYbT6aJxKdxwk
93YaI3OO8ADeiDGpRhAO5jBZWDwN8kviocuPRQ6s++BDl4Cw95hlqeYcSaGg6QWc
ukmDLMDFJkym+AKymvrUPwmuIcRfFaS6Y4Bys5xEER/dxKM2QKn4JXgQm1d1zBps
ZaAuHMCjR3eI1j6lk84un+Ryojfidpyrin+iBqbNqBgQRvgSx0Acnea0t04i3rrV
k2ifeEu1Seq4CtGDiB/vniB18TusOvOBZ9OieXztx5gd25Gp6DWmjbwM3mj+m1VB
zZuJYf4QNZwIuwS/qz1uqUY3M/7x5J+mtpNJE42lVrMy2Ziq0B9xC2hxbXzULE4r
/iQDv4C6EeSZNr15O3+/CCU2M4tx/nM6UXCgJS5jlkqWGftRzwnb1Bkdyj5Q7ciA
Qq32JszLvOp92gnsV5lZB9ZU+AVBV2Ab5Q+fJvdwXV1GJq+OrsyYOFyLlWrj3Jx0
zkuiWSJ5oA/Wxz+f2dUian9uYVFfy0CzsXlQ7Y9c/xWqjapufMZN7299CBkpv15k
BSfn5+IVTssMVN1LzioGdJaDZOlRHWjScdrd1JkEjuutaoKxx2XB2k68dhmgdodG
Tl3tVsU9ZtBvl2JmtR83wOYU2hhy3qUOGa2zWO6GBpS0YLH1uoenOXFY854NwAJK
WnRWOCb2NCCymb7ZAHIegWeK93eq+pwY11Qg6O6Y1P2QmW2Ltq2SW+pw4PICF/2V
3t5AXaS797wVBj8+MAOXDOH46HJMLjcvdsrmv6icRA/7shqekpNZlYvvWITpu1Bm
K6LNIGUJeO1HrDS0F0NFoxrVQjBr+9IpXV1u41tUOVz4H/f0zIXhr0TgEARlhj/M
YJkR+S3amtI1D2vid4MODEobhWNwE6Xni3n0PI1+HOVKZ5ykFKikLom1evlosyHM
8awDFk9MCTDA4kqz+D4wRYNEGIXjLPLN7uvkCZu06yysFbPkPHUFcBFSdWCujQII
Qy3DSkbkPTUkkxQiOBuC3S3NQFEMKI9etaJtST/L/vaItRh1fUTssppxFjlNt+j+
N8iGiLkDOcEU8+JfEfOInBjN99j4vILeLQiSy3zJ6Zz6EVbh5OIi6ToijMx0Ia8c
CQFGiZffj9yfXHmP6OqtXQEAT3Iqc48IUNb5mHkoHIx4K/uILSjOf4on7G1/189j
EaCspo5NBNGVIXu/3pIyHwXx0DPunKJarboBEBWbbYXh8Bh2sI9hsGUbCzHsSu1e
9GDsxb+BN07qwMpXx0geLS718vZIsZc109cFeuVtqK6JcpPnFPdfyopiZNzWS1n3
8zlC8nnJE3HxQLD4PqUUdUc+8uuFXa3xEVDxloXoAWsDcHRGqveFkCfQsnQ7qIsz
IFw6ldqRCNaqx+FZvLv001UMNpqb+ttouJtl8DbDuUvY8y6QFUDTT+CNT5hOUWpk
Mqsa3d4ZWW/k8sXxT5VbbLdQ65XMbjOfPkxpUYh635vgtMGSqepRF4Z2WqvVA6rm
saGg7KsiIKAYhiSHo6u4qDKMF9N//9hTAd7jWkPfBWOmC4chPWBZQpuSLxXtGrHG
miRj31WNRnzykSuza24sA869cIvnTwWqpUIRARGToIgi8wz6Rj2YFkL2Djup4w60
o+HqRcaHJira6xs81BscRH9iuK3Nau89kf3lETeGNTeXCVH1HnAW335ZaJUeRuTI
PB/F1khlMX51sWjxkK+fdhoezrNAZ4tEUbNNUPIpY1Isi4DFwPNIZHOp2fl9QSqk
csRFtcD24WJOeewHSr5//pBkc8Jwo0AhIF3N/YWOkuImDXiPlGAmHrIPcZ34eO4g
omSFeMKfNgPcIbgqE9v+B6/KvNnrhhKjTIEwuMh/hYsho9gfAaLgy+M4kpgEB4Jm
q/l5pwcZ9XQPDT2A5laRf4J8ACdxpD5Tua499rI5+yfeRnkUNODjNzRYK83PDFTt
DJc4bcRCmBu+1ehzms0TJkQOhuquVYqpPpe7h2YUDAGh8prnMGjpyed5oTllRaT9
qBZVEaRe+1PLFTp3urbbhj2IXwPZHFRD71XtH6PcJehrPSdJKGh+wYRmMGBhGEj1
aXSsYQ7pambHICus2ilFFEtFhmUnQya9K8v+hwThuncqbY6dle2ofwg2eo3xjkbw
Ur8Vz8URufEl5Cf1R4O/oR9GxMR+RPj6Ri7G5KyD63j9iXhgTUxCiaFmvFRBKvcH
tT/rfEqpPiBo9czU/EoWPvpDLPE13YFe25DBJP2hySawKFCYM+9GiWvYn4bfiJQa
imwwri8lZPderUwcB+IE3b1FM96bakweAHRwgAi+Lg26t4MSEP9r3xm6bu3NVve0
RktJTwo4ZMKtMHp5Dk1DIaiMwmDV53iq718IBZUWhm4dt7Ids++N/DyaFeBolOoc
0sSeYCRHAT6JCdO8R7DD5lBZLzZmf1bUc6eyLgH50Fek2Z7Ge7BLy6Um0pbO1P5I
F3++4mrIFd9BTbuCckidq97XtPIVjW9AKKjMJY+wnymYl2JHWK4T7nHMGCv/ODK6
+m5/7XL0S/Wx3tPc6Kq6bDAUuRn+H2k4D7G+bs1kP3rujcR/hA/F8sCJaPNfc2Jc
HHlc4TVu0h4SOsyMcs5VTNP8Vpvt1D8GEG+UU7ASQRKIJ6vsarNsW5pLPuWNB061
9KR8BwSFoUHerFlOUpvY1/iBwrqywHR1ZB+sJVC27vOkZL2ZqLXehhU9Nrk8aUAe
7LREzbRgotdo6F8+CEIPAh/QIcWYyiMIZ69gczR+a9too+DUw25eVrVRiorOQfHW
0dklaQWGOlmCcWS1eM4R9nE8ElH7orlKJ1+5zI3S3cABvGksWztqFzVkp81jSmgF
5u7BGTBF/+Jah5/7+lOjLlSR1b6ObUyOcVOSzG/nd0Yg9idYe9/6caov11PrinR8
JL9+Um+rk02V2YBB60modEs6HJ2A4GdtWazd5Am39NhUFQ7V8mRWiBHEZZRAgQM6
hCZKkogSoR5U5mqiw1kLzc9aTMH/Ut4qQLwJvv83Xvn1FKZL6at/G2vtCem0CQsJ
fsItYDVI+Lf0Gl4vdRzBRK28SgG/1U25q5CTzNEcTAOIL7eaNWp+u64rljKreqwk
pVQ6xotNwKwSgi+x2/1aVZPXYY4oXtFIoVGL41y8hUE/ld29YAsmjeJbZtHH6+25
l18eBdM6RZrm91myDCSGGG1XReab4sceLUrmfmKfP9hR7zj3v9G0Xswx+/PpmpM3
CRAUWt5V5KSJMWetXMFlDx//WxxQhnD3kTYMjvBM5k+UaUj72iB1o0ns0oMlxl+Y
NN+IPAvrT/gkagIXqpvmRWtXiIUdmkq1k8l+G+vZoRku+aGAB++ynFmj3aQjwuxA
GNsUWk5REePqEE1eQS7ivAaL1Ftc4/ltP3wMWJWKkBCzl9Phj2hUDV/U0ep9uC8X
fqr2ZO53An28WykO5B1ftUv/OMCAPg8qPIuJIBLnlahHHOg/Rmsrg1vxwgzf+xM0
ilVPnwwVomPZrsDIgsk8qOC4kP+JfNdfptG/MW1WjdkBZKhal4wQc+TKyTcK5S0i
DTCL8XTJCWQ0ncJxguqKyBYveofkWHx0ffH2VgNkhtKq4MnVCCr3TlzoLVY4VWLw
wAgVlcjZsOElZDU2Hx+h7PegCLl0tTy7QxZW59Yvktn3x/Oie+Gfk1iLdYvT7ICX
A9il0IWySFFtaNLL46rsviDnBPcU3CUZOJZGO25nlR4UN/WZHVm7CVTrjb1tXND2
A0gaXVxcbToagCSlQ9udJse32r08p+PPL/fsQ4xR5cs2cmP7sZao3JDEHn5EohQX
3+fyh4MvEixFFmURsDBFQBEgbec+eUJR45k2ksXKDtKsxCxQX4eMOWEFi8X0t+g4
dekr+XdLE6QfHoT3E5UO08LuwiakZMb6PgUv/n/P+J7jT9Mw1ZwU0DVh0mwYkGHE
dUrofRAVBeW1I+6HbjYxQ6ul/622UGMLm2AJGxUvEU6wqJtKOQfHH1tZtQFnVEQc
yFzW7HOL8x0Zi9gdU4Op6xBmOhrRvAJ6Pr/rZ/4h1tXIXmyYVKFrhO43zEXfqLg2
pnh7fwnwpCato2uLbQyZXIVUEn0gev+0AGF1yV8glE0Hoc+SkRkJ9fNhBV+1GPQh
VHCELtJiiFRCrl+5dq54NZ1+PQkyYEFyVox8wVVNBmS4DQPC/gkhlhhogs++QGAn
5R29e2vMKhk9qjrVHK5WQo3HGW8/+YMfdN5i9j6et7rCm+kmEhG3YFp6Z2SxIFoC
tf6nF+udW+RCiYcDU+AQh+ShzLaQxIJbwkFce+qK+9vOKYri3/Zfy5CX2XYtHPyp
0PqxUVWEwJ9QsFCYCxguLfV6UUfOJP5VGqbn+10W+kl3sj9k+iqRHNGE7ASRSJzW
kKPHXSldj2q2RjeX6YcCwZCZ8Dwipg8x/nN6ObFVB3a6DktVmBQIsUeDJZNJLkKG
CrDxkG5fu6e1OEFwz5jkZQQoGCB4tAQ1uEv5JSWn4eVRXmRn3epbgQBONZvqh4M6
+4w5duY1ehl66qkQMYhXtyiqWXIqlOXU3KekvAehN2HnIRn6fzWZRJcaCv2F3+YH
iSZL3YmVqhEA9ct1MnuFcW55U94BKJL44WzXF+Eh1U9B0WkbtCKT4j9gTVNycsfv
1HMK2GmfoA47NOG72yMktUe2fq8cIuKaJepTDJTMmIuFM18j2iAZu5ogGykibB3U
t2p+DFO0QJA15yNTUxNCIYFyK1iRxh8Wn+U5lX3tsBzh/M76buk/bYhbj5gZW/ui
xm8NmdeFG+uiY/GuS69DGXkOTOi0uA+PKGnbuX/MMWXdvOBZF2awDYdU5BoO9VRy
iTdN5NFi2ZO+lhkmmHuN6Vc5ITugTBp68WRVv14GsFTuQFxf/+U/9rxBSyLC/9wi
b7BCHutB+xw1yfnpl1uiMom5lXEbWEIQer7y0JeheHs6VNks4Aw/uomVR7xoU7is
wnzKBmdaiRmjwWyjRk5nYR6jBpFbSuTWaMtcoy3J7HV+11ERRUhaUpzMEIB7LKf2
vN9bG0SSQTGRCFNiDYupri+cILBrt3QMdR0eoxg2zLa5KpOLj2oU3OFIOv8aa2ka
vRxIq29g6I6QquRxAcGBHAyrX5rB5zdXkx20nRiGbnHQRohkRqoygn7i/8SaY0M1
q8/6VnK3EzFJbGePm4oheJhIyM5CJk/5H8OSk3tWCde1DqaDTPfdGbKSikQ+uQ8P
vWZXUytuH69aSMsHsH1cFimtJEj02+X1TRF0y9/tIirJey1SZx4cn/h1m+eI7SS7
QhN11/KW9VcA0brAZPWWir4gyBnymdQzmlKBWYRfiIV5mL2jnuwehOb2/TH+Y6s4
go/x3epdq0sDYzWx/mVjSXjsN1ZZwtRLVBxA5/YNJRvZrlckfNHcAP4wXhg5IaRc
+s/IrAKKIWDl9DVa9Hw3bas9/FS+WzbQ4kKNcJix4ZEQaXUiqj9AdTJcnclbcu5o
5bXFKnDMteynJjupvYNQdG8dS11kHmAtOdLqOfbAHTG/vXPycM+zauMY8+Ntqo/K
AH8AStJrQR9+Yb60zY0jY/fhcF+NUn8U4HPTDclYvWy8SCpmgKZf8ZCUlvnc+8qy
9uANay+v5VQeJlfEo79Z4AhVRR5rNgodkooVH05xP3X5BNAhox4UfxtOJD7Q+97M
P94RK+ykMcQWuCugu026sP2y31swokS7xlWvOXPjwcGwK0Arkr6YcY2eHNJvwxaw
2Zubnan89qFtJRzDNvfni1wueRiOXybIAbDOLbPZPgiM32t779fWeSkhx+IVdMFT
JRSODd+sIeEnfyv8fLNF51zZGTneCcml2Qyxkzln8SehRb7I+I3Y6kHt5Jx4W86B
2YZaa50UtWNU8wGO4+B9V+QbdYh25Cubg83qG5npsf+SSRWKRlrl7mmOBM1ETWaj
ISJBMIEHv19vDgGcB+XXm0H1i6nZ267dCPuybkRjI40Ijl49UjOeDl/IWJVh6NZR
Zf9iJG0zAXStZcbYYVfPbdPELjSdAG3UqwWtDeaaVoEEBCavvZK61LAYhi8z3O8a
S+FPnh3oz7474t80oN5yrwP8IyFH+olOAU+aEaRNFj44zNl7Zgy+eEmste/4ay1d
It23zamkK39bQWAgqM0NdZ0+I+lKQIzDgyuIVwcGkKeiNuoDwA5jDmUeapJyNHRo
XhYg1nWSRyeQaaE5wx2hf3FFDL7cGuHR4DKo4SqFZcfUR38u3GVWyxAtF0mfVNgk
OMWM4lqYtXbA73NtBzufqKyOsWhJ1mWcOVbKj7o/CILF784PBK2Qne49o+R6a3st
sFcRwigr8OG1B95Asnm/Dj31oBqi8dw2qeCaMnSdtATgiKUJXABcxKN0rymEtd53
PvQdgh7yCQvGsvsU6emiK6zB6XAjzLN5soTpCL2IHdqrF55h5cRiqHFSpU9QzmNl
IVwYyJ5hUaFLE1SPB5JqGb+79pvJm9CfSCqOUnsqc7i+k260wT8bOCxiXjP1Ungs
v2Wd4qxGZ6GX5IIJFFGEzyuqjgci6xyonofbc/Ybo7e2W0wszEMRtQktjLJlI4v7
YhUm+tbUnCfktUDrLzqCe9Kj1EiYNCTviBWCu6793fiRCraAQ7qaWxAxCEBuMBA/
wHnNcmQDws0V9qhrFnxFHu2wcL7S8fCy3+G5CVE3/yhXybJBypt6kknuBbMIFuSh
189ZjlJyhJ0ZiTs+RKJVQTaehOm6nbzZQTYDz56IJb+58tWBLHRumVkH43zQMZ9+
n2CaGay4FJSH0o67/jJBP0fDm2CBSDxWtCrPachDCtMJTS0qSzkafbXVLS2kxyfj
VLEjymHRZPx26tkSavfNOCUcvMJAwi6cGZOvc1zrLWNtnP38ZUAid9pZWJvlG2eI
6KQyxSWGO/HMYf+dvTbjD+INMBXYhHGHWUAY7zviq9jcHn7Zsd+MKm36pxV1+Yqj
dknwdsvjjWZJSA6Bb1xvDX8p4crcRX6uXUXVNsBCFLopUFpBYLupVuLqpQ9fbUIR
LG7tcrt56HXTk2uKFK/J0jICCNRWNpF6eR6AfZ93DhB4JoWWf4tUnuIwL6BL34/W
R/TOD5fKY2Gl5iLUSy+f5hpjvK51fCBYuyeW/RAvWLrxxfx95Zw6PQH23AEPTfon
luDprl+M0IlKWwNwgwoUaK9UMYVscRoRsI42sGoFRlZscbcVIbtPXprHfZpO/tFP
hzHUjuAf9WJJvAHgc7TvOWmRg3TA5VLKrHRGWhZ3VbSUssGzeCmxnewniL3kQGwA
NMf9RXYR6PTtOlSr3Yt9+uHNzA9bWSrmf6+zYtGRhb4Z0Bdn6BBbZOKmaPZ2YT8r
4wvtdhfPH4B8BqwIHQiLfyfu1gtFUDrz5D4RHuJiqpMqk55LFyejnnc5V1vpcfEU
bqrjFKPC0H980uwXWw29EdsMLKJ8JvDAAzSKXFfpPYluJ2H+Uuyv+AUqGMYNcfA9
7uEn6yyPqx9RBH6QC0Nw/8+PTkZ7zsa9IVEcO6gjQcvKFIKN1caX6mEGruNheff3
OL1w1RKy8EvVQkHNME21IzfxiyYapvdfubJQd1SQR7HLSHeGajfk/Z/jCNAw55F4
wYQLVhzyDe9REj29Mja69Jub4K+zxyrqZumOFvpu0/mdjnFb0XWeZxaYUZScqqvQ
jeSGGgv4XH1tpID40t/1XMmUe7pQJdI12nl5sH2pW/N1aU1/hBkluQWuNbqsvvU3
r56VsiLIjneRorTCAym0IQ2mTuknjbXwZz/z2gxsR69qGY6uNo+GEotpoa25+sL+
zWyqbGTuA0Pc8qEIBp/gZnXRWvhPyGwFybPnn7iT2oI4lD3z+MLIy2EdQLek+Yff
RiPmmN2cbGOZoYtwvoyw26M411RIqwBxRS/QG6i24ka0vqIexwUXxFCBy89r4CY6
omiTK2LljfEQwXcYfjaPJIMrRXzk68VPGEs+TsVkyRddIa/tkeyREq/HuyCCAzdP
FubY2/prRIbuRw+JBMIrKlJwnyqJOAgedlJQ/wzqScaxpY9dCU7ja5hEHwMgFdTf
bXSch3I77Ux/i0ZE7c+0xhs7WSFyF3WlY0dZagI/hxVAT+LIUFdjsFlF0ASKkpUd
haATJn+iWdcK/iKQlXDIaiwkF+WfQcT6IOJjEp2V68gjCmJoGzpuiHJYCQt0K+C8
36JvTAXZyP2fYO4bMv9zPyAc5rPFAtC8L2Cs7sC7VBFdU6BbOjOxYzyCsgvbnEYh
rEY/YNuU9cSwy/PvK7qz5ldankQHeQMNteMa4r60S/HplaR3zD+f9Jf7/Ia4wr78
AP59gDgZDv8PYGsyEbgr/s+tGtb4k5iY07UF36o3AA+O50d0NFZTu1c3qAcQ1vDJ
Z7TSh31EgyG3NjlDFC78Nfyzq+8u5z+SEDi4USaqWzjqOs6YMCsDfVKFG3yGgKNc
H8j/RAc0awYCp5q0gEhi207IloDAJmAg7b30Vnm+vzKcaEAj4kHOOGgC7aFYCHZW
p0iCYWdrzBAiUPcW4OFiJicJfyx1qaPkeCdc8PNUgNwq5uv/L+YAzFINKMAQxFuo
bgB9WFPWcl7c0W5+aitsQbrAMn4zHNSCyM8IKQJCo/MIto1zsSte/ZH/FgzYtsZM
qNJ6BbRjFLCoiwO5Lhoi0FJhORZ3h4W2O8UFYNUOcOawS8rW2EnTMU/41CHnfHll
PtKAZ665l/Nyi+ypKkWu5PAhXqxw9PktM5W6pOgqe4+hAnnLJPadRlpTeciuwX6N
FgaAR5O731jveqtGVN9FTK3VopGcdNrTnaEWx+oHFcCmclIwzDkkz31p0JBTQi9Y
FgK/r3ndgrQjCg49j3xQXddJDu6UHN/Ofi5vHM0GJUs6vXgJTwD28I3qYZg4aBOW
JtG87ugsPyu7abhAJ0+LA7lIDniWtG6qAxzl1szOqi+dwc2e9dcAMf3eg2Kn5SNf
T7HX1FsFDQEnKf2RpQCE+Xq8/G5G0s9fEjbgJtuH9bLxtLdnoVumk+RIbmy+2n54
PN3Lb6SiFhJxLaltOR6Y9h1003o4N6uPOjbtLJFZLhF9Qes8ABUL2fkqAhNq1obm
3oAD+lFrxUXe1Qt2vdopVwFyNKw5XXkQ/G1B/tIPcfbxv3jcrNEJeURa08mGUIos
kTsJJ2A4DDsNzMa2NWsutKjSRg7cQRm03psZlFSjzZUsNdgzHcforJWzn122vWZL
72AEEtdGwY6XfazCDVmKpBrkxpIW+J7dF9ZmzSKXz4BEMrDoPtOngADYSW973wP/
tAdDD6b8NsQZYyy/dUOkFUSLfIIAffzm1R5KEor5L265HwMIjOb7BcXSb3HMk4zX
iilUVPDpC1+2UtgCacTejtoHbt0O3Ke0yq4sxkcc8r2dG2Qeypy0a1g9XdzqRAu4
Tpkwv7pRJy54mbNZkUpboF6yfxj9WDOS1UbTDhQmqkoxWUVVllhO0GPQXZwYEGNo
Lt6JVQ+F/cJepAhBzjrW0oDjHBqwvY96KBvZcoG2xQB+7FlIwm7oTkzMkIMrxtBE
iHTrY0VbkkaQBDfI2rHn2EvjqZN8Iri77dgcjI5gPPCzplLY4VvSLbe0U2wzRnsq
gLT/bt5J3HPrqxREqhyprAgrpmvT11naDVCS1wWybX2pdPVSKbFBN8RwqvvIJbuo
EP7FW3tZRBP1Mh+H+LSDUqWsTT+zOyR0trPLmVtjw4Yypd7Hmz6xKcBMt5Zu3q4Z
ewa+RuhJqkRyvx+pYKSCeHYY0SPz6XPud8rZFor5rriA2rsqZUhLMy8+Iz5nBHTy
MH1UlQsKsRh66BK0PFlhJD9xiUauTS0QoPDjHCTKqW1ZDCDRz0Ik/V+bezMsybhO
4yyK803L0QAtl1DdkFUVcqch3kApXTcJgfO1SB/8tKwEkZtcsoJEBamZkAKAlp3Q
2dKE633O//RtaZoxPW2yubNmMRgC+YBKYr3RA23gSpl6SdHyLz5XVtKfMrf1EP4Y
y6ZmMb4Y/kGnZq6DNPgX5GRL3h5P7k3Bqw4UWSSReSH9hZ/xMNSZyJsI9MBvvDIw
EPg+Us+T4QXYONTB8eJO1CSOufPNq5seegJT8v+xaWvEZ7CyHqlfZC5OIyLm1jZn
G/vmM9ALC3/DZ6aOFpEFW+MEYqft7oyfku0nkaE8ykAIjuAqOlHU+8gsrdqgg+qq
vAwsRXYwSO/ncq5NgScwNgby+4UOqLpSWgknprwUOArGlokgj542vNnXLcemOtP8
VLKn9EMGl172fw5N6HbeNpkrqcC0e0T8Twe6nHJCETn9f+buyOwGMNvADXR1Mfid
mD/GDXkE90ENLhzWGs+pGpIAfQFH2h0MotyFZ6vQ08hjWfwnJ1kKQR4qJ+3CnJbR
/FMF4pXgEzv4raZAqSULEmUmUcYqVxb3hqwk0DpRVy1oNPY9FGZqRBbeGMi15nHJ
zKAMcMdDjfJKxfx0gDy9oHmq+rxOF+MrbwSdvGeU6dkAxVCkqGz8lzypjgeF5adm
mzlMmB4y6Kiq2OXgy/ur8gc90tn+SE6o7n0B1Iteg8JMyPaO+DyLYPscSv48QWRg
mpQpbbdYnCh0gHpfShgIgAwbIh1fJNSfWZjujYfnNcVC1ZY1c33crKa7+cYJmbRD
vSJSnIxOs9NbnhM8wQf34nHWe2LK0wOKC1Z1vg82VO3Ek563K5mxApMmh/AmRCrE
YXjjz75q2rJw8F4eNXVi2KO/bjjfcvzOj3psg9xDuyrpJoC7UOG9svoQmRRKOU2P
o11JYG1CuNSsjb2bsJMCoGuRFBwEcbdSy0vSJIr4vSWG4htgZVaDccDR/GEClDhD
59DouwwGHw/DkGegVjYuiEDsif/DV5DUIqooUhqZOBAxHTTLbKSmHyCqwJBkiTum
zZaYa1vcevVweQH1TJCkZiodZ2KgVy61GVSblb3YSi0K1FNaSIXqsA//AASTtTP7
exC2MsO4vwm7uotRSQn9ubP/ANPgEYFYwZVj46hiOWBoD97UboJ77+9/Le3GIAzY
xSaLBt4jbXd4xDyoFhJwF02bDcve+R8D6br3JHjK//yXfsJ94h90GqOjzgW+F3sg
3m917ySvRuyKEw1GC6aLIUI1qsQ2DDW+azpsCR2vxfeq1+1lmwM602KJSzyDc/5P
PNOOisLR0PWBXodkmMqnDLUqH41kKUhVOhHdtmxhz5sENcseTCbGTXj2mGYQ20A/
FMhLtjjx8tUKXPywRTkI56/Hx4Hogrpe39tLg3vWR3E8GsAObp5mgimO0EI1FaVj
FRfvaDqIg/LTfg8a//JCqJww1XJBxAKfsJa+pfq7/iQzqbuT8mVYSEb+IkjyKv42
ZrcvPnq/srnwvd3r89xJ1ALnScsVoMw2i3qaRH9OlEBfhxscXU+ALC/EDopht/1a
5GcdNx2c5inNIYCgNeasevsh82lBmyOPTFjytIPgkQLKUHLry+vfI4Jz8ybioYt/
0MqlqfVBEX6u3dRp6Dn5fpGSYlc1h0hr9Q/zjyBhFYET31PU/lgQZ+ChtITnGISq
wZqBMRbNjV+0qiDiwKICHmMPVp2ba7IIOv1ZNd8rtBGlc9XmWJmORK1l8knWqQn2
NVzGs8LY3Yu6fOvV3KtPAkzqMzVfIR+jctzbCqfn5jaSpoNeXp90lj01eaWL17tu
QSy4Z6b7Q8fKqfbw2A7sUTXdfr54byft1s2Unh9v0DdMUxE3EczRUP8tKSq6L5Fy
poTxHB7tKE6qgboPWKxQZwPYc3nc9BQllSpdGi1bpMEGsfCbKPvO+8PqmyVY7trL
hqphQUhjsqja2QQ1c+Bta01hw/0JbOzBgsPykakaWpJKdU2riKqiHdOv4VMQ8SXo
xlEOa2jy1F/K5la15P2tflZ1p6aKHq1q3Q3/FMF3wjwj+tvPgl4LfyKwDwjerw1x
Lo0xLsO5M10ivRgWjlS+0jRjUsgrtF+orPW54r6ZatK099/uUYFxPk825dlguzvs
5A9EWcBpdJ5qmUXLCW+kugbGe3SPaVmSN2pbpxteZtux67y+6swa1Th6Ftj9/qWy
ewgoRtPRsEZAmrtNken+zL9EI27w+czxt29rdbOBj32RQhplAocnZL5YN8J5SWU1
ppb/XwhOrJufRXPXHteGbRSXEZdbiXjm9CdhxnteriXNVo1JRgskM0DX/rgWAMMx
eKGfEpsSpUSwdQXAtlxKTacSAwT6Z/RpKv+UlWdqAz2zGQgX1kG1vR6lHNykFHNS
exHp9Lfoe4xpkm7j08yLkQIt5wqe6He96iZ34YgHKWwbEAg3zndRX2Ol5bAvqrPZ
O+ekAXtzGbUsbeboHtZBvdrIS1MMRqAMSyS6bJATOw0Nnv2iq+nhkZ1F6215IR0c
X7CzGz2wYY31iArZKZWiOxPMIo1UQ9FfshiO64DqppR0y8JuQSqwfji9z6bP+gaR
WmnJ2ddigpsgEo1AYY3tEBshG1Jl990BTf7JN6nmOQZczCNovLBZpfXu78P0yjIr
OWCne/Mqln8rAX7Wv8ThH0HnuWox1lQJb0bt0DaRBSaeyAN8N1cFQNddldQH4gwq
7LQeqWia3O4NNShU3Bnwtrq8jV7qSjNqrDYl5HziXePCT8r13tDeqbuQv0GsMB6W
0ba90xNOH7Z8mH9SFgn9DXoWoHuav1sx2cuVS/03rJqDBzbIBx7YApxFGlGEKh3U
Fvmay1Ee4an6zu03k24tdoxlrTu5jzuEXOBq7xFl0z7qv5W7HCCUuQ9TQfnIzRZe
Cxs0zRAJmJhRFLqI4Omhr5fE4GfEj9Hq4NC0GAuI0D1RbAIXCR/cR8FX/fgb85eC
dHaGnIABwB2n18a+UClKgyotwoZ+cl2B9tg2PsZ0ofQlqWFHz+7cZ/TFt3XowANq
Yd+xwfML6VPr+1m2FguJGN2CjYOC9OQ188bZrNWrnIPL13V+LIggpmpRBVdy6NNn
drRK7FtALvnR+unwnSdi8RT0iweBeGKNC3oI8enrBJKRkN8KNiGLHSKt+Jj1j4Fd
4MkTOw7zc+k9kr9zzdij2hbwMpetKaLCpD2y/VxafBUyuxNPAADKwafx88PbV3IG
nSbBPLcCw2xdb2U5rRIRkCgY1Ef65m/D0TT0uIHEic+i7bHrKFXuikncAZ3qi+XU
Jt5ozHoG1qggE8Uw8RJF2rADWFPL4hp802tOibMOlzRmHzrJuAEZeUePn1d/EXGc
O4ezQ14Zs1NLq+gJtUjOei84zEFahIzRRdX/ZZxqgagw2ls1v6VJlkW2RwRbWoo1
0E9h2XJmFYjREBY8CiZJuwElCOZQ5a7y04r78LjYdFEoNzT+fz9xnzs/XLb5p+/C
8/7pLZrBdh6JKqm6ilH8OgpHEJvfHJD1h20XtOUoQQT18WlF0mScS11C88MBBVAz
m4tDGSyfzcMKoqyZX5HybMKMW8RRNUco9CHQaR/cDRSha0bzQlGqY+oaeyNYqcDn
aSsG/XWcjDpx1oeXGS2uz9GqGOUzmPPTX8VRlq8nYDVHlBHhKFlBfwIZN89wtFKS
QUJMa9Hx/KTtpSUjdz1PS3MRZ2I/ELJAuXSHgUpP2vvZxNK44UvP2tckYw7VLsoO
/w8/GcY9z0glKWTcIT97Q5SpUq+HKWu34sjBqyHLYF8Nnla9vOe5p2MowLYGtcGk
21qJ6GzDbbdC/dUW5sWWr8Avhm+u9xNhY0Oz/b1qbO9zjDS1XsdsEhQY/7w21tVU
EUsOFMpGd3u9N4DFrZMy1TQIXuE7d4GVfcxJq7PkZi9g0lwgaDvmmnQXvuwrqyTf
IueIhRsD79uf0QP2Cz9dPj10f0AZfG4qZCXtzIILBFtnhK/rkI1HffWxOG3qQ6v9
hYf1X2ykuOFlFGzIsPmCdlvGNUG7UpBQt22f5D91SksLjnpPiBWP6ZskLczmwfMg
oMGEWlvQMrt86Rz31WUBiKx6u6Is9nKvMKQO1UFhR1/EBJZI+Mcr5T9z7WJnefRo
jy6s4rq9L52p9Hd6im5StXXclW9MYJUNEmnCmAk9Or7GWYnon3PYEVns+DQbnDbd
Fh99sbRHX0HSRVisUwxHaHDby6S3bVfgnZm+urV8Mj3Hfoz+FznStZzXlvNwtiYB
CZvNEYAnNkqK5dJSRfx13czzk0coSIIjK8lMXMMpnXma/WWxNMiADcwkeMYpa1M2
nQC6xpVo93hjdEc1vy7WKDl2dARbKpp2O1/noQLSytLZKUlmCy43KA8Aks/tD/eU
mv9d7roe7oSLaQlclJeJd6vKyvIGa5Gis7Fru9By1x+h5uU1Du/EZyey8h++Jo6J
kR2X/cq8AAwsojo9E3tco4zFg6gi35+3725Ene01qO38O7ggPFSDKtd38bWOnYoK
15gMc8EDqEH1+kIWkqp38RbvyUyI+1u4g8fFQxub+JLeTtH0yKvm2+zwCH+4OUbL
XOtw+zEasW9okFp1Msil+uM7AcMHWbpAmm10csn3JayCHmWcxnSy7Yw8n1wAR8VT
dDdFvSanIFTMDzt0Q0tmqfiTtynUti4UFMaVejIqBY2kurLAkUwXYfoZigUHrzN1
0ZIa5CPFXEZdYRVB2rPiZJFjr7dEVowNWgf4/BBuS1EDo3gQaWE4b84rgPVBEf46
f/+9I11oxKQVBvQEyAmpyR9KHRWlpgicLPRo756eTAGH+8XD0tcSvt1Qg5BO81ze
EJI7A/brh1hI8KxDwvv9WuVyFErVPkeDFBfe7fH+ri3U6kXQhg95fBDHqFVc9C8I
ssMvdH/Wu1PMaFvL3zi29iyCA0rsQK3CRpqbZzRd2YLVzxcNEKw06RjEQKSWDpt+
oeytF0mr+Pz5950Hc5raA0NU4pGls9ZVl3+UgXMAMaaBAWe2PpaOMHComVTdaWYK
pAjDelkiDHNjFOg40wtHXVfWTE8w1HcCSheJrM/tLXMWi5f4BzvMkpSjbScG2GcZ
LX3PmRGW5dt9ucJyaL6yQcb7aY2YrcmfgoG0J8gaNq5CJenGtOIaf+30w25eLGkd
opvHIq17K5dNKNAkXIzqSkfrluEyqP9/K3CV0WNkBLUhf64WMvSYEC86wb4swBMs
r5PQ3kjSgT5RqLYhFn4qkrhdscBhX6nqmNkvkQHbPSdhUvI+loL+bPG2NLXW0D1q
tLKIl/Bo+cpV1+G5YPatizZv/uKbbzgeQLGl8pTze2kHngU7Yte8fiQtM8Utyz+b
p+AmfN2yqSaeR4TLJxSH4vRSedFpBsovMCqUMS84LjJI+G/T55aUubC4iohY3D9H
KAwIG/TdzCy3pjSc93cDLXAUWHPHei7QcWmgfzrr5dDN8MDZSqCnaO5ETiU5dYRP
MLRjwnUaT42Qei5BVyWImQHJsTgR9Jj27x228SztV3fyr8Cmr6ZZ9s9V1k3pCTWE
EMYPqZSeGiEYFHw7gOQaZwPiR+vop7xdo9AvNG/njcr+cW3fpAdfw9E9q+dF3N5a
opIu3fPtqyCH9Ly9XdVm2tDwhio6wtdXcLc4llX0JToHPXAQRfS55SIlRS+Q4Jl7
w4SZcOPVwKenerEhu5vuje4l1v+xGD6d2zjY3G0o6s3Upal/4+C+fCnIh30ZmgYu
vKEdMAsu5Oixdjd7xchJacQjoGC4vhx3Bg6YSkh2Uqwi4k3V/L20+v2I4EZCRCRG
FxXIb6iDsB/77i2RE5CQQnEPSW7M5zcazvyrQ2lsmiAyr5hw2bELyiLiX/APCa9i
PINAKkIOF1X5OmUyXeHf7xrcAl9u3uvTBBp+ZYAThk7czsWK8a2JgeQIIfJZp+in
vst1L9+QgWdBqC4QTThuwL7dOR0Uzi9oy6XG5sX9gcM6vDXTvjdEK0hWRXX+0E5K
aGljMrarYSIbHPO7hKf652KmWTXXUmuz1jsDGxh65zVrM2fZ9tk5Xut7x9+Atp/F
0ylj/FxV2Mo3hsYQZH9kAR/p+WHgjc7BgyX1QDKweFhnZrFODCndGG6A03sRNFUC
VPQAi/By4fQR6KhBV+HR05klfrE0nDs6hePpyju6Ln+GUzWDSsWgJ3EOiA4/dh3R
ERwfNQSRrdXlbF1Dab+aslj2tFl8oOeai8qeqPo9A/mzc6qqraM7byBU0wMESIrt
np1AgMneZVZvlum6G7QIB84Hqzb60ipnHfuID6zSLiwHqcqHKOLz0H7qXBZ0mdU1
0ZugwKfBQeKv7SxMFM+I2uHdUsX7ol0Pbf/T/VLCm8eH0sOi2AkZ3pQMqiRRIgUZ
PJavT+0ngObmWjpRQECz+nMaUAafIK71h2lrR5bjGPfI+9zw+qTmrFWk7wrESycr
ABjLxmEAwtIYB7yChQcI09zGF4fN2skEy5R2ZWy3OnhOvtkHaE83LbtjC1w6fUS4
cxncBwx/spwqyqGyRs8kjL46TkXJ++YlMSVdFgQTokq2L8WAUz8seOSWze9rcUh7
fU65HwKMhqHaBVzLbk6Sl9AZIOIs0Ud6OWwD2/DemHzBediruqcImODEKKbvw2Pt
a53f/bl1yu+V7YxI1YcbNMbHzrGc7X+8ZROg3EZGEKSv0xfYfUVnKeLfupoWyqaj
7DfdIOILN5NcR7Jok4PZsb83L1nZ4uBHmGGIK+jdZ50p3o6oxQMKxCoCBRuafjRK
CEHqjQDngjGgeRv57H5Ur/cjgn8WHeI5nN9r0KTHvuF6fnNqr+GlmyGECywauL+m
n8PftJCc8JtxjJ7AymdwCuw2MUfjb4LI/pFnMHb9cIzg50O0xV6pOyu6maP8TKni
sWtXKMbaHYgnG2UWxut+fk+9/eGca1ESHU3XYIkLjXn70RhxqMQQdODjsSZdlURx
/deGZzAoxIbewZ5Bd+SQDeHtx/bwMifCWvD5P8jcDBrU7iTAM50IPzMYikTnbur7
8dzj2ihgqxVqA4owJNpqgTWLaekYYZqdK+nOCkMPt3n+FvAaKyvbxbadE4V28TGM
xvll/FSHcy0VwAXfA1iV8Y1AWUTKuhYbe1lpVvNhAD8M7b8juFcPSZXUIzVTD4Nh
CDkJUspR3oWzaFs2sl1oUorFQ2XletUWCtLjjJizwqhqfMue1RUl2isE7E5Y2Jna
LEYuWP3xc0k9uoNzqwWSNsNq7utbXMUqH00lq658Efs7v5140KW5H0E3b+KtmF/w
mI1OuNN+aLaxW5R+SII1nCvJw8URyqRAflms9H8O/aSnb3qeMbUHGmx4wulc4rxo
Xt+LGjFjbCT4cRfExx2Q2ZW4eSxjqLKkERHWlqWQoQ3CtgIkPtMM2BY0Qq24UPVC
B+Kn75p+kFiMp5Bw+NuIsYaVGcn1HMlF/5uyTiuDMnsIjz5PQauffJ4WVOqoWwYw
W3qnvvhTGCz3HRCbxxn80axRA4TAbceo65jTRSe9v/Yv9RjMfnq/UCRxgwyeEA6I
e1PlstuIhLIFYkP/ZHChyGrSDzKvYTncSDke9iM3xomXenDhM/b75u6jcxGNiG6v
P3yJaetLP+VSmYjLMH/oh5E3md+WV4OasIVYqR131VAkn32NSc8Z5wzUtuuQhnjW
/Dr6ZTGALcFH/tJ+QOnDotMiWD10bGkSXNO/KvgmWWxSF1+MuJsg1vYsJvjXV+ST
CtqLeKLjeU3s70BxvDhQjiK9+bJ0xe0mqS14Z0dgJnH6Rt1CusyYU9Jwsj2gbaEX
geR52INqmj5ytaK9i1z5zyI3airr5muGsu3fq02mMldINkzIsxVOTNyqz9jgbc9e
Dmi+WRwJGtThWgGa562DpsK1rXQZ7fjkSEnL974R3Dmm/Vf45U0wpHYOg6hZi90J
Bx2I7Dx6zwRViUdqET5wuOdgUrO3j+qMCTQ+iGdOYYPm4Opu+Iod28htBcf487hz
21hCCubvUmbIEjW2StNilRvqnvf10mD+7WShzmxNgBXCzvf8QmMILxYnqYThg03/
tRRASa4GMbq/r9bQ9Np7dDWknvyrW53A3f/tmDIi3AQ7biTNVdIRJwuzz3gHicHr
sooBQmq6quEz7r8r/tsa+LVAmee96QIMwHy/a/u2nzZ8OYViSMOFa5Eb+8tUpbLb
t50zboC8tKCwfWYxqN45TMCyJXuyIuVneDqpEV/M/KmUpRduZVEq0cawysakfsTQ
pRj6cwul3TZ52XI8AXdpuyW6CzBlAQJ65SsJfLtSh6NowMEL9Tv22S6UpASxee31
ny7iRPqxSuBZYidOXmLWq3tV2BieK2KVwdZsGgjLogNcXSzs+hZjM7xTYdJ1ucuK
UhccHQHXPnSzbjpq7FJvNF0jVwrbAAe1NQOvc842jqPzhfdLmHZvBb61sRe0EvI3
cSd4Om4+ubyHxcTK/dy3XF9qmOcSMdKsipFnoaL4DYOn7F91kyGGndsmncHg3wiL
JPJqrrWRJtV0kW+QQjzar/jOOmc+UDMP3YqtLl8MDlkLjBvegjmqv0DL3V2MF6xA
jYdRQXO9eOEk3lDBGxTLib5GS66o9gaKjwhVctU0c6E/zc4aQ6BrWbSdCdotdK+m
u6rCosaxlaU+AV92HpKKe+h3V8Tk+boGNGyMdV+a6zbJZ0M33YrcBm9/p5BKPval
pGPtjmm5MDhsyuRe67qHMPrYrADEHJ9HHMCAbMZYH+ue7y+OcQiJty//+b5/L1/j
dkOTfK99R4ZTm7K300rAc0UyGHGVn3OcqZix9g0PzssbZBBjfxSDxemCkZE9fZLR
zUlXZw8GyOb6pHG9lRh26UE9kOBy5LvjtP6t5yweEQncrW0awTK9dUropItzHNCB
/f/IcbZYZW+9n2WxM53l0/M5N11l2H8vHYzO20KREeluxqvQGLdhV38nSv6FsYC5
Y5vu46dJVxmMRE0LKlyQJev8Y2YrsPrjU0ywUMOMYEsgbVJqdf3PPRsQh07KWRPf
kDGgPkbmgxOyGtIAGVCXud3wQkPyL1Mx1oNH8hgWw+l6vZ8RQyxE7OYWcPaUHhCi
1ijj4HLvMrloETn9oqNiLoZBXhKIZWEUgPFUSBh2IlEUKR2RDtleLhDAMkiVYxiN
z5KwfolM95whG+XAnhzBZ9UDATR91WqHc1YaIPuhZwMSUF6q+iOt4G6gGlngnJUZ
EJyLy++lXF5OfDcu2cq+j9kQM/mnOUfVO+Cmkeodh+ybSKFWvt5T5WodPNJ3Livi
Vg9JicCkOk/oBZ7DM2EeB3Sg4lFSY/un0BHN7k15dKpy3LCtdZTCXFi1FbHfDi4M
fWqr/nMkrmw4qVbLMJ8aEkjjx+/q08v5rOMyDzek5iiyHELyhrM0btejmz3aYdRg
s1Y/77ffFKPY8cxFWv1q6WShR5O/VYPHfqFvSdODxm2bww5AZRx2gal6cMAD3ULt
ZgNIJ3R36jpguxyDINozY2RcpLnl4w+rm2jqdTsBK5EzCs16C6etSBIv8oAsiWJG
LF7ZWFFdFafel9vDZXZq/o/nWvR8j8gB95tpqgPpX8U7Xdj+IE18YU3lIqLn2YvT
KeE4HLnX7e1NNO+5cv5J6xjrLn3U2tQdUYoXCEMb5HIaS43vFOsQFPG0hvZTVuKp
L6sLwSZIvsMx/y3qYElZaR493Fc6nT58XLqjFB5EGqi+O4yerTy4k4gSw+T/3FPU
bw4cSJhmOFA20Myw1WpIaAX0ZEclB/zDM6EXOU3lpilIaicDYVlKFwVESpxJnHVN
lYMvxmg45qOGx9pguchIC1aCWs60tYx8ALcVqSCHRAEcB2TpnrO/LJ0HOhQyhNC7
GWBsZtLiXsrzZC2KQZ0KxpXoNFQnlUjyO3Pvn6WD2cO4u6AecWqA00bTGGOWj/7t
rFJSUa2LMzl35450WjVpqK9ekHDvHOz69ob4XoMszOEdvFykotnW9hjM9nAV8de3
eVYrK7hav2e3/QQXf38TqSWgJPHHcWh6hsbpcdjoS3Mv63/3AvITK6oP9khnCFHm
lZGoQllKRoldpflkhymrWf8C/VdLUxR2nhCCtjiznlh/j+FGr4hNrhZ65go/HNA0
vrP1lTCoJpeVfjfXXfAbfeQxsPJU6Yz29tmtCeTPEIf8QT9p2FeTtkTIGybsKsUt
zumNZtff9Q08VWsyzGdncH+H57VZqOejH0Dq8/uVkOgeguP3R16nTM4IaWeufsHp
28rXc07YLj/zGRbJs67rOSNh3bk2/iHA+QxBzxW1y6dNNdwv0M+mE2kHn6DZZwg5
PTvfG15NJFyOCUSI78Bmpt/68j+njYxLCeW9II52iNrW/9At9QWQYXJs9bpYd7dO
Z8fbvXYSKCheVozFWm+7fYDDP/PGUEuRcffCM4MD4k2AKowHt2a6+zEWS2nfI3/M
/GPvDh8qLRiTIpuLFqOwWMASSLJeSlGPQXsMVdnOMzKsanz8DyZ/RX9veeO+R+/L
8erstuVWWaT9WHQtpnZjxaNA4zCdjSYuqSZXlDW4o8D63A6zp20X69egLDSrFTUr
ZULC0SC/Yen++RQP0IW+Xmp4Rzt4wvkRisZOViY23ylLBEyPLwl4s+LcjbW/4ZA6
pNFHaPGzDro7k9kA3fU+MShmFTQKeyQDEd1h4OJD+tM7MYmOz7JBj/lLLbAPVyd5
JnUTbpys09rr6AebIpu3JSfGkK54XUG2r2NnIF3FO4d2BrV6eIpWLNswCMzbjJGd
DtOrPiKtBBtiVCBtkZwfqiY19JVL5skyEEdZEAqeuSnZnRKwEklE7cnpP+GXst8B
3Kc44rqh21BdjDLTrJcooK7+tYeaVxUJ7+9/dBIkQsesl0BfMWgdwubztkOntbEL
O+UNjcEi1fkNq45QsRn+uCLFWe0jYLGUgagB26qvRxZcckz09Xda+eXYsjBxlmvC
2ek4+c/pg0A6E9GUtmDYgyjYEyY+VMozZz/Dzj06aEL3fPDDd8ezPB1nyHGu1X7o
pvUomfRAH7xIQo1B9KvygUEo6YaOZ0Tl79OHfZBXr6vsuk5DhpVIG2ZxmJl0SjVG
XVnppCdvgVFilzhdDIrpKHJN+Y+Vo92VzuA0eoDUaMF/S4pqjhne+9HtSnbXj/e+
nWaVYl9Ds39i1ZCMvTgxJhcdMhKpuxDIY/M1fIFGo172wSSqfOYcnYaZKUnQDYsx
ZieJ60m53CpYKBB3f4Kv2bdKp9lWlD6Cay6wmGuOj0SlpmDBPlWEN23G6VQFBh+S
RbmK3jbSkwOjTOmTIdEmM/VIWaomukNz8Aftxlp+CoSOy045U8cUDnnaNizI1SP3
a01VsV2M8VeP0dLDh242K+VeBR1Vo+fArXZ6TcvdEcIgZ9tXdXPRMYYPaI6bbxE5
XAAABGHM1JlESvijMKDxhxcVoM08LPIeQrHQvhOaEs0UhwFAQtDhq+tWl0SanxNO
Sv6KK5RtXOsFnVqjlSYrzQKIrRKB2zU0sfSl/e0eHjjnxP7W80sMG9jr+em2QZCq
YEpAU44WYxQuzWn9qkLTUst2Cz3vqNMtH8YjiOjqbm/qIoPt0Sal8wDRyadJq7Re
LyTTYgL0EA0vF70w3BU1Dz80Cpo5sSpgZ+kJ95VxzG55NNwpOK4sVyr+0t6VMBlT
l736zL7iAFcakVCibFFaxksPfDAESk3Oeq/TlCTtONR0z8faZRpPHQv5KL2bV8TA
u6cJOvs5y3riGebwHoIkSbfwDCIdrZKBIczRqhaLOHNvLRjOgIVXPMGa5pDhaHrh
IlQmT5mVVLa+y+y5iuTYYKGjSsEf5hnC8z46Yw8W6s4JQggoJNoWyIBbQBXXtJR+
ogf5UNDPGW8/4bdPkkdD0XfqP4xD92I9iGB8vWRJSXwg8WWv42gJ4fzTo7gng9cz
eGI9qxMv19yIIlj8VF+4vAl3hfUM2PyZbqGydaIsLXuPWwDQADEpdQJ2YEZO/jTO
Hymsj6BgEbtOTDH4Qv9qJxHVgjWIyY7GRyCNxulqH2fJJ94DeYL9lg4/EeFFAgTE
DRDiseYaMjj2eSLNV7v56hAWpdFQ36KXz9oZBPxZrZNeBKxXqkM1y4gbAcSqjwzR
XqMwkV7FMB4mn5XJB63abpgllh+bKXs0XewNKQbPG3aCccbGKtH8n5cactfWJEb1
3GSWYHGQE6idoFAhrOaPgYUInYprP5/X+0VmzaSH5EYWM6SdyaVl8MMYrTgX6Syd
AZd50RKsVUvsvQ9rk33RRHhFiUFd/tKyNj91VGzhgEbifK9SQrfcCYSEu0BluQbU
gR99a4rnaJb9jtjFJdqKlgWhihN5+fqbQsoNlg1IQaNrv/LOmeW8//FOQewgIvI4
2BZLznM21BdrVJqfT4PYVtyJtpe6B6BtjUhdr7f8qWiDEH/Uk51yCUKqGFwGOUgS
h+7ksFy61oKUwJ+bmdgLRLzfZSW/S8kMMGpuHnfeq0hUF5w4gyrC5Dd8mN7CXuQ4
kMB1fAtZ0OmP29xKaVPiEYqpwVG+nnTqyO2LyvCOZoraDTudggytZmgGeQbSLHZP
exxqqQsjeQDtudpEr78UuoMbQRXp6ehi33d1SZe/WcR8X1DeJp8EK7KvyxuN7prW
mEBRsoW6L+94SmAlSmZxTsIryPt+E2XqpFiFdkdyluZeTn6N+BtNvtNDLtdDV450
ai28uIcsm1BPcyy7/TPYoyJLNx6uO9LT1ToDestKF8HYrJ67EUreCgObj4a2PmkR
3jS4cP9F/YMtWb0FIzlW849y4+UmDDRTYPPLsB5kJVEWndBZL+XTVodIsKYCJxtl
GYgmeSZ5WS5TtORDWo+eaGCcyjrJ+Ycb6FzxmkqVQteKwug8AGVKbszvj46ZJItA
t4J+G29RqLkYoEl+oVAtA4C2+FLFFQQYEZoT9RWhnE++g7MARk0ZzGJvgxauoAeP
dKfy5ueROlJSidpx+ceRD2b7FlqucxueeC8+ZCB5KKdbtzsNbtmZVVgxG4jJ6jf9
lTM1wEp47ERMGISMJzts9VGAIWMifeoTt49CjoQGETxiRSVBc8v86giwdCEpLI23
8s+oI8wBNHdbxOiyF9LuAR5h0V6H2zrGWa51+0p/8wPSKAci0GPHHcvoXvjnaA84
1Q0K9pbX67JrN7QVVCn6z+6NNn6kDZflGEojbl7KTkuTj7+J8gkMLXSWN6RxuZ8w
wJKavJtzbHjdq/I+/qF7KLZcgYD+XVu3nid7FigTmvXMLFSErPcI1QOeLKLcg+rN
ojw3buPuqZAMnANqOpUmzdiJ72IC6pUMcuLk1Bp2SK8IFdEqFOeyKrTtkJmjcq+o
PrXgrsUVphisFfnzbzoVnUMDDQHySTbcA4NjUIgOaGJWNA5208Cp7wvENupm52lJ
t8r5k28gH/MNSTaTcZg7rQvXw7Hjp07Kt7VTIXtfRYJCF0cIsMPIceZYeQLsuFZM
EkTBnfSRz+ARqPYclWOTgwgwUk9QUqGB6oSTyU0g6wOZqLH9/ahxHl/gJrGjr9y9
tsQQN9R80GLULRqaiE+AXu1Z+7xOrrFifzPHKwj2nfwseq9IAsQpSwIfQ1ui/YAI
UBzpld2xwyB6XOaSpw5Hmcpq7lbe/wLp0X5si4t2r2N0PNO7zLRhvlg8C+UOf38H
K4Wua0cqpv5J6Uuvw+eeHaGAnCUNoxcssKV9IntXhWkRYuv0dFvVbABCxE+7e2lp
a2gME9pMcoyhrje4NzTb2E4Kx9k5x/k1WKBCi5uX405O6q0GIhR2NNxdjU6XtD42
xy6futGvc0pCKGgF+pIq426h4jqbTBfT2Seo+kTfdZQiAsVcm90HtnLC/0Xlii79
RTpJeN7Jk85B/Vr96U3p5aE3vlgnpB0vZlLAK88EjMwumWZnbR2NbckENJHWkN5V
e6jTHjnoTlLSNrJ8kYKIcb5F0AOAO48VWDEifiWwBBFbaiJkLhuTVu+xw1Hx6Bwa
1L3xq858E+uCJXXhlQCTsN0LJPdsJuAUzh1n4rxj0wR/SvoZIgsyyjRykpXVUzCx
VlZKKTCmPHyDmUMsuGpsxYU7aVkEtsHrCkTaWcTk/mgQm5Y+JxnFbYQ78VBqB1Va
Vpn0UbLqw5d3EHPgdOGOeYe95pYutEYYyUeR60gKqMYZb7W/hFGxnDF55Ax+4yO0
uJnMKzH8E6fkcmQqnkE7AC7gzrkni1VEbiQpFDh13QNX51gsrOoEjU0BNZOR5ku7
e+GVQ+BbxVuLtAUFrCUFP81T5G8mZLU7yEUfzohuNpwneZJouh1a7cDJ7bAG8FvO
fUXnwiydRqCKRCty+bGfIMpzUt8+QZnqvSMMtVunq/gMBF1wGGjS4PDLmocqjVn/
UpzNupTT4USN83Km8aOxsH9+4i3gBc5/vO9fPxQffKWBK28jmDSyhRRYWZ3OFMmC
tr+C0WPomvjAxk4xJfeZyL7inwPxJicfIx7KOh80jVsaRmJ2FjiN/bM3atX8L3x/
X+Y7hSMOCGVfuRazESyYq2LVGmTKUe7v9khJf08uBgCsbF/bk44H9PzKFuCSf32z
ILNLdlRuyYN0uW1FW09dIxef6sNgY7EylH/pB28YIgk7EiQherRq8otjjHj4fopP
FVqgB6MYeWst3A40TlL1peds5XFFjQpTU7TvO52zVOXg8eswJEmRtzng01OxXjG4
xmv7I/jvkLkAE0VFNSGIlu9uTmy41ShZYPEnLgXigCLzP70MfWQW0Malv5DtQdu9
8Crc1iuIFSz0Gl/KRBj+aQFWMtdY53urPFWP0X1jbMuBB6zFAGO1vreXL04XEJel
4rkhnyw9QtIU8io97w/VYfyab4of6n/I6dK6J340FXIa7u95Fj8VYEF6NkIFE3p4
FtO8lLBFogGWKp0jbWMMk1dvWOqC2ZICqUxAv15XZJteRZUqEsvfRgX8D67Ii/17
dJRoJ3bZQVQV5HCy5xioPqY9Toq5eSYIKQljO9M+MwvrYguaxnNeehaYnu6ifI4C
axBK05fq6lrMZKFJG8vdXxsmLqraPrJhunR4MoOVkoikgKmZDByZRMNi79b3mwQ6
vtm6eJI/gLseUT2122fmrPpDMHkarXBnQYHS+g9hhPle9pgfW6Mscw8GTS4QvSgl
c3zuFhDjhLZkmTSem8UFG1MiIwaig4VzZvR4xkTN3d+4qMO0umu6hByx0W35TR41
NczDwPIoGIhW5n/X70PldRtl4evcUi9T12KpeTAfv/PYVyZiwW+XA7bmzUOHriJu
n8T6RmjVKK8tDcMVZRIakBMsVs2GJSDjc69Ot0SrmvIGbblKBsnRNRVYDQmgTSAs
gZ3yDkptVTEb80P+ZR3xNw7o/GIE8pEG02XX6OAFSBC5yAliBbwqg78tIK/c0lkm
UBi6krJieHf5n/zEND8WiI6YRvmQnYqfdnm0lk+NBizCrf2YqROjZdfLHV8v8lDC
7TvdzybnoYWSxCvDDCLM2vxxG8lOa0RYkA6CH2SCpl3yaL5ScdznSTCSUZpA00ct
d5p1RGxI0AeRqzZPu6pwHODYfqzVaxOSUaDG1aa6ESZPcfY60nnBRNSCR6RgLN4Z
xcCRwsglxa/kNLmqLB4pRaeKccyMJEgyR5Jz3ImmJ0vgIdi1fF+5b/uRO1g1jObq
ujDfIX9Tp/W9+OXV4arlVr4SkXP7daSFg5CKtY4HJU6AHK9f4ENBpE25842/PXkr
n7yX2aFN3WhYoXL/4AOMqDNsy9Dj68UWsrsq759sRmjfZ0CXWutOz8WP8rVfy56Y
kqOVG4GQBGpr/RhO//y2xJgF+Mkf1ANAoPPplQLxM9PgAL60XLp8XVte4s5WRsuE
QZE233gWokYFEODeIBUpqiWNe/J5psVM4BT74wi3QTLGroyKL06BmNS2A4xlNvVM
iuxBRYQXjrUVmloNpBgCiLyQ/5o7GJwy1KF+geIpur4oEkwtJLl1HomwBnrYFA49
mevxekQLRRuzfBTkqbjL4Gz1XfFmCNFtU7cEZqWQg8HaQS5jeibGUvM6r46mdpcC
aB/YJTC9icsXhOE8XwtT2bXxvmifa8uLVuj+n+149oRV+UyNQwcKSOfQGe81yqpp
i8EWWxnUDluh3L5Udhqt4JRCQ9XAEbbzXpLRSy4VZzzebtYpfpLFB1P8BH/sutnU
tdOWTIhqq2kIMtMgwqHMgN21sWh70xiTvb25CFn1TgKkJuWYneoQOzJ6xFgEvZJw
IL7LGxyq+8InJ4fpR31ZxHC7nW2WOhI39Q2IvFT5SB9NoBlcHWVDs8v4r5JtjVkQ
dXdnAar5TECyZnAoj0hkcjjk2JasvxE1pfnDmGuqGhmG254xhb9RVfx9w/3UU4g+
qbVZ+G10alzIWorFnX5hGgIcpSeGPSvUDyLSEqNh9HM2zvLDKQHs3Z7ucNTcyxF2
tXIPfxFDPuDxzX68Ni/2K9/DNMW79zTqJ3CPLfxvQ//+dw1NoZghf/jWHxe7SnCe
tkW6kZw/5WArprV37VozF7jxl3Fyx40yD51dgmkdVy2pfuNiGyJOoKQ0mtY5saa3
89MQJlLjbUJfkauegADeRJGQD00ZCMUQTZVXQtpJFTMxImcUNuJQkP6MBGUfR+fM
fvL7grR/ToCdDAcpVKDFQkFLNhS8oUHzD3zva8C+BZMaElgLGhZR7OsjIpxMqob2
Vi20X2Erv5IP0ksXXbbTJqwb1hONGDXyyRrSJo0JEchUFLVgc750DcMMMypBdO64
s9SDUlXCJENopdhKs72dCsuA7UunRjQD1aSJ8xhzWdVfS+WXenZ+KcyJz5FESMtk
nnvIVqS71RxK5+eG/qVSWtktv2es8rzZzDFkjyKT0SwNgQ5Oxi3Gsesn8fy54iOI
5HJ0HtRHnGR/+Y8Cp1Hj+WL2htT3rPDfq0pyhH+5fj3t7c4/XH/EKebzaeuwPkFv
AYdWvQBn41QddCwfZJqcmv+ra7UYRAxNK2X8gDF1vPoSa+uAWvHvTUbiFvEUU+3P
f0X6WIyvmhWrlY8tLyN7GWMwDm+POpy3T4o87xGDOYjpejcYNtuiC0Yxwofm/fqQ
H2XLvuJpiIhbMcZdKlQdNu0b5eAhWdnlxNq5tsOYbfLd9blZZpOLBSL6kbdyTgdY
CpAwxw9AskPHB8jvun8UbkYzftlwxvJ8aFmlxQicLxHQqHth1JJKcuCuMrQSQfIQ
nwRfqxg88monGT3js5C0RLivXJ1LsoSo68tv+jO/xH+xGf/PhbcgH0iNSvuSo9oj
CIanp5NplscTD3OyLS0IFbnef2SC3RwY5d3U5F4R6IScPUOMfY8RW1i93OcvOKXB
Av4fIfoz4krP5AbVLS8ql2D4fNHhur4VTTiWlDzOzGF5GBMsZCpGbqPc+cVgNlxJ
/1scOUidwhHDuBp+yfkcq0UQzsCx/2a0AFEBSfmKMmXLMg6Rrfp6Gd+nww21vQya
eGH86AAmfQYDgTzVu1QaaErXT7X7aay0oMa3GUr50tw0p+/EWhcLBFudFe9vali2
Rk4XThfyWsRqSPX3G3vqcsTDma9q0ZPYNabLZXTco3vHJHKavExdO4ZI2S7iQfZx
CXqOz/H31X7BXSWVB4ZlOhGNzfpae1SXCX7Xat08R7S7TEdrI3IC7VLopk8pjae3
X2JLcgzBW/j7Qe+8WvSVSxYcLa+3fRFAFKPIdcpRe3IYuXsueJ3wov5dKEQtptKE
U+YUlUoruf41PH3qQY3qwSJ7YSW1J2JuMIvT9zHtDSKF5hdiESfxzqTeA6vXXiAm
PjQ1zO0oRt1uU9ekuJXEPMb/iauROY/8NRsTM0t8ZPRztOIYtYl4ZnemBKx2gZ5l
cFawB8Nnu9g7X1IIV/ktW8wA+qOnoq7QkDNmBpcFElaKaDNDnOpP5PeervX30avh
LI1RTFlaukiC8bz1d3WjWw4Z48f+/D1gts1GlvBLFVjKW3BQxfhkxjtuGvm36gg6
EWN71VtThpAAQfNA0zAwwCrKSmF7ZWodKsKUjsGONAbb5ovZo+M/Jzd0ClWIYovh
e2N2Usreee2COdkWkZWCLXvtgVucAAryoeRfQ4E0vvRuytpMxTzqhrVSOKieAZzs
g8jKWz2V3eyDMR20xnbvubyWgYf0BUbEhtXwvI2WkEloPICJil9XBxNQaOEg2xlv
1L+BiNyObK677EOD0uCllWO95VPU0X3uzdVVZql1BkZpheDKTzoZjMSEDD6l+suB
EjN0pmuEgoXva6y29aZ4Ulcn2V9qbOyloU3irxS0ytoExcq9FrPOzZO09NpW72fC
tlhSuHQGUYuAoVyanCeqWFwb2QFqYQA96qr6pd4KCbMKsj3cP9U9Ovb+a3HJHbnY
FtqUyKAptZbC5VVOzeMNYDke7XHwcBUysCytUSqJ84Oc+yo/BWKGU32e7mWkT7kq
iFKyz6goit6e2z7M5Es+jdKYZf3hRR/1mpLwFMxnUWh09/n40VYudXKlt/q4zxDa
O9ffO8YdNd5bbKpTaKiXjdAeNpKLV5DrPLR8YG2KLOnImPzWzrSge3Ro3DYQhaog
UGeBA5Psn6yEuRy4R0kGSwf2EP00HUL+zS+xkKrItrh7jpdk6L1VyZ2Hf3/54kHv
bxN6LclOT0a1JZ1ph79Neq7M6xR4LBA6298x73IPnb9yOdcUCSJSmPUlf3X2EkFt
aErF3o+tKq2CaC/AT9cXpfVnfTTLj1ZWAuw2ErI1YK1HiZ13g1+FQ8lrwVLlesHx
bV9foGjpLn+JmnRqxiT7ftlt+WLXdXflNMUDHc9loOtzURPu8y1HvHL6eE+1wN7/
03lSwfsTISkz0INwUVTjxHUZ3PXaD9f+sni+weFDHK5rmPNqMonPu+VkX+brmZdy
j8h3lDSK3aoVWvc2yxRPfBr867zx+TlPcsuKKXgWX+tYuSduDfq7sD/cC+6MFcEk
qN+GAtHws8xQprJcKLC6cHWzTbQODdu9rTKsBSkSRfFsHtrOZSeL7YU5IDrU6Tdo
0Rr000SPssBPsjI9PlrUFL6vHsBFqUk8SBoJnrD50vDalA3RmLihYUZFbtkMn2Er
kzMUQXNifsXJFwEzz6vB6/kIm+7lC9v/yIXgSBJzHstlGIGsLC0nt/QptVanjcme
7rqNN/IMWFGjs6W2i26WUYcVnULL+O6LP5GrB7PZwuj3piJ6hzOqWIg0tqE2nUcF
zpSDkFINzD5OuibKuXSNnHAVwMivc0MNyt8xVXikNPUFlZzxbJr7YbNmX0eYYz8/
KxMo5PRMIs2PCR6h2XXtcR1vjSzEbUZsc3cOQxw9HnWnXp+0w0kR3leMBKqYhBBI
e1dWrL2z3hqsPnzwcn+E7EvHcxNpZa5SJ4C10Tb39owwTK/f3ESbxrydlZXhRqmQ
QsY9AD0HmvxgghMTFMexd0ZDcMh6sSQ9g7ex/ONfrkqza90DD8UTuujCb02phTtV
c+ez0Y+EQw9IIUUGyxPrANOx97v1Tbpv1A47c5/9dwshShW+SrrY8AVWnDMFPsNo
VAfxrblw6y29chv1iFlBt+HuCcw6acRunbMJ4JuDJPnSiQ/SYeT9NiXbbsimtlxq
mRJ2CN9Sjfu2day/IGaJbFRl0uediP9axLBe61rpoILPVUCZZgkClUb2es0S2c89
neIRNqwWGGckAuvMoTsDPKqzLiD6acQnctjRSNj3fBRSqFVMg301K5RzncKL9Guf
FvGdhA09gRHguQUrLEED1Z7ngSfbtG3hX2/zfIe+ZkEXFJ8p2bT1V/d0UiKSF4y5
w50aDRmjuRA+0KPs/NtthkY6lz9rdV+EhU43Hvuzs3DRv5Qz6KyyYJjx34NDaZ+h
LuzDqskF2wuR1KLCbyNHyfOmsIhera8LUcU3ysyFDoeeZr61Y6SeHWX4EPq38Z1g
4ItKDTYgzSPxtDACu4W1Ff3N2grEYtNeV0m5UojJTYd8zppEIQsZFRbifly06fIy
IKA7Zq9/o5Xf8So/qrErGCnKWhCPMSxG2Og+4Mk4YYnB3rc0zAVlVzXGuI/JxrNS
Y7ZNVENwOZm83XSx023Zm0lupsNjWmEaW2wPs9fgRoJP9UrGmSQaSmgE/CaM/txT
Wjc4zPuvURh0mKwqrK3jyUezennrFZxSlIH+DZrl1xh7mYlkj3XiXLf6uV8N8Jtd
UK2Z6aNzhc/+MZlZUc8AZ5TpiOkhaz/wyEmxQlmoNJnsln+r8Fmy9r7KiFKUfra4
uSRep9xRwMaTRbXu/oi1g6kWZxkALgGo8x6zhWO/O57lTDSrJjh+5bxSbaEbhB3h
09wtqDLQQevicMwjEp8o1ukCQy68IWNPDv2TFatBMPgKnBjQUFsMT9Idqi5IK4AF
p54vG25t588U3NQVATtLsnAYJIWCm7LTePX5bJNZf0HRUxoLyZtV0RnAd33nKyAG
bjnUL6oQ0c8y2rdcWjw/ISjF2vQZ81jmeEKdxtTWSUN6Is/rR3WNN6pfhW6yq8gt
PIzB2yoQHIueH9MFekKudwVl2kXNoBmTFGnI2l52G180sG1tTeDWRBlA84sQORVL
5IiKnRPZBWxV534qMdVfknIHtxHZJbz6xxrgNnAF0U5pHVcwUa4ccZdQ1fvvLeDa
SPTlnPafB4fXkHUyQKdIYscyVtkkxEQOJ9y1dWma8Wa54RvbJ0PCQcjXwQc4D+mg
+WIXNk4vZ+j/QrpEqgBLCOB/BNtadClROcXIWlakQMfCJviQrbHGPDDt3/Ua/rS4
Oqk5Fn13+kg/B98IPoIYcQXAHriACipjqo34R9Tcu54m0OkSeC++/lskTqo7Ju9Y
k2jk6R0rFQ8zqYbEVKLyEXrgia8DC+6fQWK6EkTBiyjpvd7AIgaOfSQPTqT1+3YR
5WFGRp9mKrO0PWIlG4+3sFQLy+Bfko1g7NtNZyEjFMjI5SUcJVkGq0xsCvnPPGSU
5iuhZgJfo8A7OPA3Cc58EjiZItt6FAMK0ZP0KJ8/ZdKyTXEXMQuHIEhInwWJFoUz
ZzYabkihhhfQLhoUxRaZ/3fnaLQirFvPTalgB9JrFdzU+2I51yDSr5LNniba6xh+
hq7AWlFtN9v6x/fJ22X/bhEEGaSZU59sZo4BDbgflckR7vyNvjEDk2TrWx/FOgmp
/0DXkxx8sCB+g2iJmgdDQy/Itw998SsoFW8i87dHX/Q7t7W59E0y5qNQ2E5mN6U8
AFt2CTo4pL+FuRimtwDGitaHetCuwjkkFKnPd4TJk9oLfyvTnvzIyPerTBnRbfel
u+x0b423XEEu4tPUPQwA7svzBHwT7+Icbj/XI34+bObx6kWpqvjuwM8EU0JiWVma
RnyTBPaipHns0nTBSJMkfLjGw2Pkvos1X+bE/QINvtuK4siHYIzBjGKriN9MQ3T1
AkE7DG8+Oj2Xu8BOYBuiz96ZagovNFbM1ugnbeoLAiEFSsFcmJTpgTB2mI/P1OwV
J05wAg0g/CMa96hx3EIs1hndxrn68ApLTLv7Kp4Qa1utfa6hgRq3TE/r/jb8MqQT
NjbzqcVrS8HFKF3pEaadRbSkDOHjY0USMGNNlObV6GbP2bhFs1lOLrjaIVqmo+Z6
E9vhwYSxkJZ0MNUGN+4yOenXSRV5tzMEBjNFwJ+oTpzGcm3Zo+AEDABkjpJYMkxe
7Or+QP0sr2AUnGfv7Gki7IM/XvnDJVWBzsxOh6FHiWzbu9Wjooo7NcLCLIbw/NlP
gzWYojgq5Hp82muJZr4yTPu+pgIv1NCIF1zJ6s8LX3eKqECmulXXiViNhGqegmaY
Bm3fz4vVwhR7RLC3j0wMTMcDXnOR8EEt+NmlqSElQfY4ic5O3TCfmbRXMfIecPmq
L5gqF77KTGhchvCbmpKEXbBDylgPkCcRG8zorhSKEbIPTkfHW6UjWuytcNFeNWrT
iuZ1x+tsP0OUEUiawYKqcLsXd3/bOefIukLuTSN20gnZSgY+PwEK6v5+Faw5S8t3
X1b6OZucx6eFHOTxxO4ky2UE/15CRV2IYdHclMk0m8qRLqTGk9h29cYvUqO4GdsU
7nXno4jo+Vem1StUythqyyE91gk7CUq8A7fFLdwp/eX2Jg+BrenHth+kbeWc0MUd
LvGgrL6rmiGsFSdjoLmCVRX3qRQY1c1vI7vEYCMa+Po+EwJRSYrMtmpm6ZWBBK+Z
l+1pW/NSFa0QZaA5166P7fnVkFOPF9K/RV+bXIH8hflyRHcCJtAEMhEfz9XyJnpk
BdjmMx5iCcfis5UjaqLae6LaeNgqh7pEWOm/F8HC1tTrKUJoTdD/s05bZ4JmzULr
0mBnUfkgFB46yydY0r+WpH7714ONo1y1m4wb9SPzBnX/6bjp/L0/9ZiGfUPhLIld
NDhGssOpwFtCiBCrCvT3DqCzOfnWXWYap9R2g885DWk5gq0v2bEmunQvSfllG9V5
nDs2gyZGfpbQ/OREROh90kieKptfZxWt2kI147cCYOCIz63c6HDndvHJQagVcZUj
s4V09h6Tf/7jSibKwrQWWSGeOtkWmrdROcvGZbIAqtpxnAVKCO3IZi0cifa608ZE
1p815k2XoNqpOp6D1kUVICKR79Y2QH+klIbMBz0QusDsDfvPtYgBmmEgxEtE0tQC
pTUUCEQFvjJFCJMBSTkRTuejYiyUcQagPuRxAxgBXxWKMGIrIN1YvL5rqtLOZLIl
w8Ya7Qndo0Dkb1RHbBhseVFHivC3VuHtwPQsdBc3w/vXsshA4oQGE2nesvtHIF0H
T1dVePH/xtbyU2yrvOvvmdzsBYqPskWZI73xI6eNYXOuGpKmK/hJdzBKbeo2I9+a
6J171v7wls9AJfb4lzwMxYu+pVWhZBuFcDezf/+ypymNnLT0w1BoxuBg7eVdufk8
rlpxV6TOHSzkn+WCfXCXrUvkojeA0eihzh+Hzuz2iBUL6teCBCtwOu9BdOsdH/lx
3NmyfmioUIyuxA7K/f/O9Bs0DbP5GiOBW12GOwel3wSYY/HESIz9eDBALyVSK1M8
VwVQ02HJr2fdjV9Iw8ZqQZ3B8czj9YjuAUid+ZKf45w1YZrE33qaXBl31kLsy/c3
uRhZSWRtbytJz6twR2R7HaOmjodYsQ51huGhPF5MRTKeJU6tKoiTahx0kKu1/ehu
GEJsWW6wez4wxwGOGMmpa5BhDlHlV3CjW/Ce0xWFp9BVdhAQd8GJUGjMNXzF4Kt3
9r4pQqjaSmhGyzbVZoBKvNZIrVyzj1eSjjBqQvJOfGfNCVOcDe5oO6vkL9IhkIV7
x8+lYKCH0N2wS6LeJ9JlzRU9cVIA4Kum65MMvxJmJngBhNJ1qtc3JglIOgmlIaPa
PFx4t0h86Eyj3Dgg7qxOujEAwiwPL+k5yUsIIMbPJjAj1vp8vV59ZA6V69RDRtrl
Iq/Mbm6l3AycTVnuWYQJFje2hXKr9PkM0vOn2zxk00S95v+Kvm5N4cRu+NrSwVqx
oYM7EZMbhs1G/aeXZsndUb4WwX4DJAAAlJ3CDhFU0dEaZHIomBxplbUCqFksfL5Z
28YpYM5802QTpa8NQSaSrx1PQEc6dnGE/yD22RZBifzRTMOPypjGi8GqyQlSugca
Cvdrs9gOT3gzIoUSycD1vhHzfWaWtwXnAk1EUAhWxqRJX1/CCmA/mWW013oepONk
N2WA7pFnwcADfRXAvufIHeaD426vLH9yLi/e61F87U030q1UYa4GxXvSTJpZi+Kq
oOrnBa2LgTauLcnailRZbNCiECTKgT3Yvtj857tymOxf3WnpbJTJCytEXbtWSaRy
lL11gGouKWBfXWWJia+ZM+TN3yOaD0yZTjFyjnGEBCdb4P24cF9wCnKICbSSaMJg
Birn2CVDvcyO4qHUo4oz36MnqPldFbHY3fbskkQZrye2/WD8P/CFsFgIn7TIVLWp
ifmbWOv3djM89PSeF8JcNYL7gMfglg9v1r1CI7jyli5Ionpm2bok1IzsnmrCU/eX
puzjIwTqOeFP/ADlhUQhgQbQiIv/4YRz98Yfsiij0WHlZ2n9vNHRtJ1AtpWyyQ99
QjuGg5JMb5mA/LhTHPmKgVfpIlRenoUd7mwgN59omcq5wHj4p45XgKcOpPxRoFPX
kKAr9swIi9jAXh++iUuA6+SP/Byw/5+lMt4U8fsLknKwnc4LRw1YBdHiiLm0cSpv
73LvusJZpmPYBznwA4UhljOW3hLyH3tCDY4uqzXOvjEQdtdND927TdEJcG9z269o
moZLAlgn6zgWkRVFTLH1gboQGT0WqDzPvMXpGFuy78bLp+h6LddHyFAGkr6or6N8
ULwttOQjVFnw+eH+XiCMtIEoWe4PtkHHotW9aJaiaJ3cuH9i+0mokm78k8bOmVjx
DDu+L+BLFpgpo3WTwoGc1cvsy5iWNXi6NdJ99V1ME/oqUpGpiOeqsjryc7sg2JQg
E4G+gh6kq+F6nRkGXwyYA1gDtsWO5HrNX1Hy1emz67p49XdMEhv5ROPWFl2jthWR
pT7E8+jhF5SMRjO40J987vBFr6NUM6wqqmYFTBvNutIqW5o6uEAUgokC6ogVsf9o
AQJrjTkZsglj2o8pemNL4ZMcDGJs+QkoREaI9FL77af76aki5JikaQEpQpydrknf
ijpl2Tnf3EpOekmPwWboQJiY+CT8vXkJGWLfXWFu+kwbCWCU0sv+1Asa69a1FyUf
JmIEfg0W3FWvjjVSrI+FxWEfyKruRBtiKL+2Dic6sHqLqWlj9Bmb3nyU7ET5qi1h
RKe/rnhKJ5kAEgp9eioZM6m4+fklOHL6ZXQTHo+81vfpKCAoWA3yjdF7hUUO7EA0
hCp+pFqYoVU0xX4XLMOd7dBzbyAKU+oxJhMA4z1PMsNWgTjX8yEKvm5w9LvFDTIg
4+3VfdKnNR3mD7dTPr4/lUl1ZkwGZ/+1atH4PjzWiJsUYn2DIHsYUIFpIY/iF5qL
X6QyFT1VKHIXDdlvIn6ihAn1TCgZg0wWs2zBnuRSD/a4LFbiycT7Z9oTzFTZ4S8z
KEZNKojRT7Y6uVHMTsrtOyTfPPcLah/Hs0sfgje/0D6JhqIqsUTizb0ePCkkkEoG
n6XVCjN/MLR6iaYsexZJxY4MD3tfCfIvtnrXa63RmEGcEBjca++k0V0pqMXiMmrH
jDNusrE8sbsWx2zFO1WFk6MYRfdLrhmsja3mpokkUTrEeBxeaRM8px9uUlhnD7Nz
8ebTttNC/zTGAP0AarpGcml2aASuXoQIjZT3H06VI9k04J7zk3r+6HxkkVz2sgFf
9d1bijwyPU3rQM14gl2Z2bO5weXKdpHNt3r07JQnl0w9AKL+x790QHLVz4oT71Yt
IFacIqKmXQ8O1qHY65FG7rnshIOrFHtluKvvicCG+k6hIYF84ItWhzA6vy0n6sl+
PgTnpIVmAia+dh46ASnxoqdeGQgphfXAARsmKXWeagu3iLJSGYRT9X+Okt0ThnZ/
T4jV8PfjdFOLSikft08slwvicNygtak4e5AMYI88YLAxV30Qy553xnWdgZs5mnZ/
nYMVXfQOAjZyxp3GV7ryXs6HJh4cA7LWJIno42ZWUUVn4R+xXzRVaV8IosriS956
wgITIcNn8zDbXUG13tguCBM2N6Wpsy1ofl/nsnUho//p5NjdsGORC6QuJjvmLy7y
5gvPcLN1M5HlzBQx5qGEqBglRRwr6DXzx9T6dYfWdF3QTa46V5Z+/jLssOaw38VB
VP+5ubkjH3xV9/rWnN7moVzka+XpOWdGLADzXyfSCjvKsSop9M7C1loCPyGwfoNu
eBStAed7JXoQ0TV3q5NcPEe5EEYl0jyoRqGkLzSNjiNqef6743wUMmzib+KY4zN+
wHxp4Js7ShM5Ptm8DjtJD0a+2LfeKqOF0u1pmHy3QbWlPw7cPIuLXay4WpQ0x8lX
FXhJBU6eEjvMNYqMcOfUfgmpcuMl+aa4vhDmZZ4ZQJ0XXXs+RDBgQxdhDeAKYHRA
xAwHSV0GTQnFnGQoqf7zVCXCbiutqocJnCRl8FxuhC5W7Xa/ZX+PCZHfxxwCV4Oy
FZ3uRLmSQbuIR6iV4VHPxyhkWKwbO8Q1uQJgqjtUwiugfWEjgh2fO6glixWlNZHM
NG4YGifkPSo9mE9SdsqYApNBDHdM5Zo93HFfKkfUIhC4+6tSmcKmkNG4X47obvuR
l6Fc0KhLnHuYAqepEu8l7tAAhZNGSNGjXR9LCCyowLGkhTTAMuWOn12Bzv3eMiQ1
qyxXPvqA1OgcnwwEcrRWULF/HTBrlFuj6E8Jhc/8mMwYLIf2ZtEqUb9PSHOum3cS
Cz08+OfvMXQJwhKSxJBi38+dhIug2AvGUWiAS9knM83fkwQmUMSlPZKPv3W4Ri/n
dli+wabeCYslrtKK/R0L6tapduuEPQdzta4IT+ZAVzpkX1iNbKsjWzqmJ6HbejZ3
89/4ZAV9XllGFXB3KLqfKtJzina+BsWHj0sz9fuT9d137HEQbSqIAMiRCbweh0kr
Y5ddBT8keMA9y16Mh0tCZgPlaHR5uu8ZzoR0lceYfov5znpbU5AMDJRKY7R5mLX/
S2WMmkr/VgEoJ9shg1UaMw9DBsSKbmWSlz0RcNI+1w+7BX3z3EdNrD3NpE+mF80X
4/KhtbcM/Jn8lECQSuagfcWePKmDE3GBDGMMgi5B/T+U1csPDZe0W4wNibfsdRlc
i4sB4elwm8jsgUWLz8pUo7+NkOhlglC5ppKlFgUv3O4Uh9Wq801SSsMlQ9C/1jhy
VzMqm/GNly6QFp7XerX5AHEwzw/sEFtNsdqJkkNXS+STceuGRIZgdN77BRBr/X8M
KIBDyI2WSSeNKE/JJw3E5jCppTnas4sqknAxqyifQHR2QrKLPNnNEljWQwsLd7eh
EN1EKtPl/3+JqZ0JuK7xSLG7jyUyVcxXJHLxFQ8sEXkyuZBygp7C0ZKnaKzk1xuF
HqQr5uEeeWqUHSL8yPFEoGT1QQAyDXHd5ggz97xwH2wE39lz9cNvN6vvC8YzxnLe
MQ2wfyvfQU6wyOIAWO7OsrSJHnrJqWIOw0fpxHmfavELwXOd6xVxgc0RlhFEVMhe
X26wRW2SeFo0fbcadm4Fh13n1hWQAkEipNt6i9ITE9uHOvbCb7kmrzfpWq2kFPGX
STOZu6m7MBtlDxh+9XS6WeScBlWK+JhKMSok9PnHUwGpq9s6uxLP6ABIx89ju1km
cFg/lpvCfl6KjQueWdLAfwjMIGgqZfS25tdJOxxZIawZZ7HbIaFBummcp8TdHeTR
2un29UaFWmIVrM9bwE4Q49Ije2B/azI0NmUnDVx4FdN3wXPS+UQsHda87IqcoGRm
pFMeqegVgmASbM/YYGQhh6xcoZKFxBmTVBpA09hZmS0rXS6dt0kTOkPHdadFSpVu
QhebEB5p2UeyQvIm/ZQ7nDaBQoRARnLZBH+QhBC+/TSys+JEgEZCxCIiwOP/wuP4
64KwGjE/4XWyNqt9RSoVClDsluktwi+FRR3gP/uov/XBh3cZtJBEi7CNwr8l7glM
HU26bqSSHQc3SdLJi3TUP+q5XJePA9cwGEylkSjTzteA2Ft65VCkXLTlMuiUU5hZ
rDI6goHu43JBdpZkSHKRm8eOA/6+SFvJeLItPt8jbvgfqdgUZNTSP62OnvQUIQ7x
N0rlncfTOIyhNLFmEhy8mR3DoBdVDxIYmJpqAqyBHNlFVwgfXkPUkQUJi7Z490e8
irkWwasKIqXCNJK1zBKPc6Bp3aQZVAZUGYnREAOWF4ux/BkLxS/ax16YTyRevFFn
eP9U97qrUnfQO1jpQQQ/hDNbhF/8vXOy7J3YHdrIou8l6qie4tcQ6TtvJSm3+VH/
6fha2aQp/j3fKKeNJ+4JDXA2XtGd2Qw48AALQGLrOpfp1nplfhjdqzDCjAnX++LM
el3W5SGTmLJbvDGkebBIQdrej70BMrBwvr11w2Vs3z9wFJQ1mSlstQ8sh69JMZfn
E7L76pI2eeorx6U9IX+XcCmMlryxlSFDcLQOqy97t1fXoFevOAGQPx7BUfsbGYuD
Je3ElhavqS/qZTMw+UVBmlSCA/ynS7jzlz/I+5o5Ajmmu9rog85dYYBsLQjsFQCB
eitq7z5AjHrj/UfbBzTM7xyjtdSjsWoLOy3/hK61GycGW1DlplhbC9AfpATZErOW
p3u1IGNOzK6mwhbrETo6ENYs66m8x+EdZyCCV1HzieoWVKtYxKw/MEHjI9X8bKa2
W70n7Gfqh8qBmCzw5z1S25ShBmsYg3Ko15yzEt4OcScq2SxlXFMWbfTJsKdV41ZM
5p7Gg73U9aVe2yeeLyvYZ3fOxFt3bijm+XLeLh2ur6sGw6MGsvo5C641Uu1uGFt0
9YQ5Q2j9rrucAe5sxy+qL6hl0mJOIic32NzDFkRtI09Wf/unAws1iDjBFaBXQ14i
runUesf+thNP+d8YY8uvS/fSTHuX/7eE2JIjjFQ9aMQXMCqLnxloVqof2I8W+CYv
+mUZbhM/HRELcEGAtaqFJPGuLIwTjT/zea02hRmGCm3bs4uZqTw2WCkbvSYBXa98
EYc9W01nAc7BeJXh0+xRV/zb5Jizi29O44RVNQ/FI2JbHGTh0ECAaFY8ivq96T2n
ehZO0jepnKAerkxNCXmvO9qDW12V4U6eh3eIZEkltYApZyFkm2mcEMG9NJOPAXbK
dPymXCrhJS1Dp3p4qNHpt/cqQM+yQvI+I+fwpBP9T416bJY0nWR1Ws5jPUVfD1E2
0MmVskVPlCkC5UBBr4a/2iqsdIapoIt0fXHk1khV3GMLhHSypj6mPlmA1Y35tbl1
Plsp26aSLdETSE5+6mX0yGCZrBgUzmdm6cy8XK1jY5P17Cerstt+g2SbU+vkh1/T
FSqYDs24dPXeFqIGnG+SHUl+T4zpKOBA5V59fSNzyEt75IKyQGKSz5L7Kxvh7XUE
iwiGBxkH51x939lEPiYTd5gJai6ey3pPn1HrXr9SKV12D+NCr+GRqDHLhvI2EVgI
Rgn65VQle4Wk1FQr3NbRXT85UaFRG809SUrcW08it5GzvU+DeGTcswXsSjHKOrLv
RbM4dZiXve7PvVb89seg3qxt5s+5oET1LHHzGQbai6tXNu/GnlFJNmAiqNbC5Kj9
W+wZ3ERbmiEw5fYYd+wD2eJNVX54spP5f1gvBiCy2i1RGGZuA3ld8z6V71w4sF35
xCGgqy1P9stp8dIkLHDTj/byLUc2zi0fqgOxU7DuCPPhUHsErMm3MGDcSzA4ALlc
m49TMj4uBOOSEDAmPgyrAkWw+575OHnFelLviwwzqCZKYJYSWvLpAV+zqsjphGvq
JPzzK5n4Phv43A9mI/shYexepdJIyTNmKf0Lxbb7sVrwNjbcY+SGbmY45S89Kvn0
VHz/g4IfgnGU9UlObeLkK6adqjW0P9ZjjXFb21ez2HpCe87mbGvffioLcWxD4489
BOMEo3KKQTdz3dWRmroTZt+zDh4IWVdT30A6WfNcvYuYS9jK21/UlL00kEpT0a5W
EJKv2YHC8ZylIrbewVYwpyZUyuZ7CgwtaXfEinS/kSYlPimLHsB0WBbbVJfFEiQj
CcHe0mpWe5XjBBYs5YnM7PPeB5E0VGy1CvdkZDZOKIT0x6i1mD2ZzfJw3L3ku3fm
32nKG1KbE958ZE7zYKZwuNz3V2muYoQIAy/3grIqCUDWMVll8OdmYpu04VFA5x1P
xwbI3DloDzbVfFwgd2/VFcRPbY3JTyk0eWRkTZlJ8dj7PjqmEq39SL1b7o6CfdrH
QXaxRdXB6iH95B6d53wj99Z+4VXY3MNUCQVSp4r/FneV06glux+Z3sJPbnnHwNAA
0Zj+qe0fObPRn1TdHIsldkX0F4clgk+spKNbo02fIGbVp6Gvl0km6qNo1bqHSCzt
Yws1unTVpvh+Hcs3vcmRJ2WY3a38TMNXlejia3VGGW1PuMv3vMb7Z6/9nqItkhbB
HhWGFqmh9OCcA3S2E4nLTuCvx30e9aP7GLG1MwmaXZZtRr7VodEg33ztToTfjD/k
NtRJuaTu1ShwESOa+q5KgOTpzMHowOkViMLqKVmMYgiTSsozZU16ECaTd7Cqp/ub
Bfckp/UyN3oezKPjRsTjxvocFJP/foRfkiq676DPzP5DCAkiTagD7oXjfFLtQSNv
ZkXoIoV/CoitAVNvOedaDAHRAlgUkTFydSvuUfs5K960io28mulCCKnMmxyFntDJ
4T3qCR1ZIgaQCoV1yNeeAZRZlR0gIruao/0zDXK9BIQVUtjh1OJHt6xJJZKPo/x9
JaUjsOc00xA7OkgRbK47y2mlU1/B16qdYnu6rHxeGO7SbCavNVh00D457wh6cyUW
6LUxyBqPPS7qGiHpwBRL/WJ+00JsaN4E14UP94tRZsBOW7KVj81tmN5Ev7N3QTp/
6PuXT3aWUKwKYfdho8oFaikL7kHvN3SyCI4xs0Pkxjsrv2eR3lcQMLtmwfCf/Y61
MDdkbZMbwU5NykN1cF7BjVTKKlTPdIyp/a/ciB1pQa/qBYtszUO9jH91I2K9xCjQ
uVY9T689OslFXRS5ufKZuIg8L1hSuQTo7Nqq0iptfyJZOp47Rg/g6Tyrpg1xlhwp
GjGX+Dhp1jXamwXqg40oFmRSx3w/O9owvRFhU28usurpGJgFPfSlAdE4RFK30Lgd
0Xx4OqejL/+RHyOuEqukMFkEaxqYWaeKFj1uoPYSYyk1NfmheiDCREFyEtn412dA
JSzoqaeUakITeW+rcaY4keMDkC9yOrz0/aqA+IhGLRb6CjxW4PRZb1UNz0SUBUwm
0Jhc4dhMzS9dzHlB7dOCsoCqOecFs2GnpCFN7qKW/RudVRqWhXHACajnpVbtq4kv
UzADi2Cou38PcGkGZzGgvXPAzLd2HHB9kNM67cjhdEPJcJWeXHIoLGNSTGwM+JWS
UtpvRJa3rETRmgDaqWgrk7xLPoeFg5FnW6G5Ev8+nQDtfm7DbJ2wFqESZNx8NgBD
4Ju3p5LVdAqYum53vMxTK6FXctX93QJD5gh0fkxw12bGD4w4UH2AQhGdot3w2McH
lNHKwQ+TJ04X4aHkkXXmEdGqoYpdCoGwKMXY/cqQ4bzqvOW8h9vTSQ0coufv9As7
JNnDTvCpOak/DL0yMG66TOYBkNlbIxcePgbz64x7tkJp8IL1q40mdXMuBWKQSfHy
cb9udyX6u0WdKFNPk2rRD0DvFvteUEVhTUxxaWJPVrLVkMUfm6wywP3NM1znRUi2
7BJqGWzaqPH8UuQ02fhYIO6J3OdQhWXCuw/hXsiiG3WOXgSsOguWy9mccW1P7Kht
wa3kK5eC+u4E6a/+h2AcCPgs6u53+sxGWZxn6wHVGKuqLfOOGvVlN0zZhpb8wiyi
iRRxxGvpSIrIyyM9TFhrBbUkyHNJuUA1xpThBgeRA66B/4C7o2qWcdmU4fuAdAK4
NTPJ8QT//fz9jBXeAie/Uwic43kjqGyYF/xFRiSJnDscZKPouMSx+fzXPi0tJeUe
HN3LNmeiXnM6D9T2/GBpjLe+A5Ty7723+9XSBmUU2GWFnIyp+W+dnx70BMFW+DTl
ij76MbF5Ybjdt4N+CRl839UaKz5+UXGbWPn2mllZ91FmJ9u74OPoIql1xj/A9Lfl
ftcX8xRt81CzFncKzJlAcdZ0ogKZuRIu0OXOXPiVodwUlG64TFMLbmKhYwUKvK0F
Qg5ZaK+XWIcS6HFeQ91Fpm1blehtOH1oZulHuVEtK/x50ypkpIFVi+rPvhf2pAC1
FbeigmRs0Rab0C6uBVhH9cjfRQDW7x9+tlocDsrJW2qVI1R0wQgbf4eEpE3S0IW1
X40HFXbL6VxStTdeFnF/9jw5U6I0zNuTCRd4KN5GYDZ1bOVMYTIseljGYVi4z/8I
/gSWE9aCRY8GJyPTOx2HBhV2MA1AhyJd+9z62mkr6dcDE71uooosm+ZhN6yFMMfX
m+UmpdKTSl0v5XH5G8h+q31WuFvcXGro16L5Eh8OAjfXdMGGXZ+upY3u9IIUhQeF
Ta29SQBPCl/n2NbjTxcTCF+mPTMDM37nTnMVWplMQw9/ZRqk4Pc8jk0AHepNru0y
tGFteyIFjYsfdAdqtEuxK0AlXYUgGngt8YodRXrsdEdpGB/pbMfDUmwlQxBAe350
ZuE3jq/hA2VIqkqXaR5vmSzAjlRjvEGElq/8+p/ziqlFyM+vq/PAS+EVtB+dp1XW
h5dtnYEZ000OBsWBC5V1ny22n3nAwExkwmr7634HXcZTSLL88H1Zm2LM2WgWlvuZ
BrPLUuLdpJHeQpv+7SqiBVqeBczQfd8+Vzxv4DHvIPt9qomAnmJuxnfQDM3g8WtA
Cv3tL0rThdObbz7vs+nzD6wTDqI1gONXfIW4gsoBRdlwokaTyA2RZW6CHMxe19Bc
Igs8brbqDwIWw0/nQDzX9ISG9RufPjBNeM/tfvPQtAufqd/uaNwmTMju/HvRWbx9
wru9tT4V8bGQE06sXhJbMSXZ0h2Iz5z2ebQ9dfQts9hDLqxE6ZaE++NsasLULEqk
QrhilPR3K69coV3ntLPayRYe4Y2CiGv5HVQKty0TItqHfQTEZbfS6bqdmc1Cl6+s
n06aeEO3VRlv+a+fe9RhoPWDrNWd0zna7KPW5dRQnoMtqkOhVXoXpzeN74EuCuqU
djRy364xCvM/66Xdv1ybPVSkPGK6pYYrxO+9sl+IBfrSqV1kYLQG0IA5XrlMWb9I
jCTRbVncIVuCCygJ2tJzk79cqzg+n4FwIuNxYZSeWDVe0jQDCstT0+L3oQaCCpTX
K9SJVjAl88Q9FH5GB/8bqjNZ00E2tjgmakMn2d6vVFdHSYiNv0GZfy5CVAkCjSL0
yQweI8BEI5nr6hg5z+iWf5Sel5XsXPlQKlMzJP8Udrq04Kzc0o1J8fImSBleD6XT
On2aE6Jn5LlgdJ6+0bFQHIx9sfJFySWAzl7aEGACFYU98/OqJ2iA2zPourSwoklK
zLuQxSHL74vnGZOPi4y2nnIktjHkkXb+QbVEE5QfZG0VMW61ljuPneEbtYb1yq19
C+T02pD2t6Pg1gWhlf4ReJW4TSD00XQDwmkaawgkxrhhMNxpTYm3Kqp4OLI+X4jx
Z4qqf62D7A1kvNFGB9ivC1BAgX3QvdzgL8nIIyqIqVCzEnoVQXUG7QOe3yc5pwn0
/jqkK12/HY+igIycjkDN3xGgzOqMlGdZ/tE4alfqVtjNL+sa5+mFYATmM5u3M69e
sSJv6mVXBGXq4Lpjo85GOjpzEK/oZvh+R4dgBlwHT4/Mar9BAREHMDIVS6QRF4bV
WGxF2qjlUrn9R0ncuUKNKMrH28XkAcaB8QbPM9n7/rUh8Pl/TL7DPmRaFP4X48Ux
a2OY1nDfIEBCCPzM2p21j3stbiSdCW6X/lXhHh2d6QxOedN7gpKaOAlr59cy18Sk
PvuUfsadVbe0YK7kpuPGL7lOMaOw1ZwtaBl+t7yOQRZzQdeqR5AGxJdEGWlN1Px5
DGXrdZ4ckFne7TJRB/kwUh2sGVS6Vo+VKjztzgcoSCrnan+A9e5QLEJztBWJcYyt
u43KkV6b491q3FJwMpvIjcbAcAF1E07+yBIyeCDfHpNH4uDa5xZDRfAVgvwpsKEt
pcJgeAh+81MAoxrpzo9oxdr90CkIVyB1IZIgDITkX0MXLzokTHIxi3+d4dLZDQCP
YN7UQv3N26/QPKp514eahI0rPEnHVSBi6EmD6Uk3I6K3WJZzK0mWxOA/9RMRvVdw
HH5JNRiRe4q40keroRs0ixnTfc0LWvB25D0DyZd0u2FISUSAt+q2/0uxVukCWnPe
dD+rQHYlvuCpKYPfk4fe6C++tybFRHz9QsnlY9jtZQah9eiZ8Agd40oq2HKHPFS0
xEkzsFjvVT8Kw0OGR8kmdxoD6TgQtXjDN5UzAM2rWSKxTVwrXanXI7gVPm0/50zq
DIXOELaLSHXjkK/MeEF//Cq3VyjC9cwtmjEjmEzdbTY45+ASoXKnl6UE2ETN6j09
DOVBJCkh2efYmRG9izdtWNNSVu71Ho7Hspu4iXqoEYOsmYR1UYrDd28NOmaz4LoR
aVx2qw3CEdKxmy79j8XiSMdKO6e+eA2yo9hnAaoUDfUc1j+sFeRxl/itpSIujdJE
BU/jpKOcW/SI30DI70k6fWAeq+U5I16kdm1uA5Zf3L1NtG0cQtg3S69lbSZLtcz8
TNX2BZ9OPaAyeW7Rne5y+a3zRji3qhydAbBnJ6xYJymWvMu3iSVdA4f2GXIZrRQ5
zFLBz26Imu91NYRDtKX5uc06+f590hsfuU7b+qhRd1hhP7+JdSYnz7SCz/ITjjjI
E1cHobmkqpxOQrRid3IE4o1hLx/4kS5//49jRuuorhEZuUHANDrAkfw/msfzUDE2
NlFQpxPG/mEOG6xiza48tw1CFGM8/kQ0SqV35PgxuA3TChSyzif4/AsU623Ey5cb
Q4DyPMQ9rMIxW1nBGs8ExltXiRIOntq+OxstDyQICCgBQjuyfaocle730shdv1jJ
FqLWW2/geCUFieV6ySRlDMnMvcKRcIQ/X4QtGMqTaRVySsH0h5HT5nHLc56La1A7
3FUaHYEl4r9pQRRSD4RobO/XnAEkGlXZejQ4HsBWypR8kgOE3UjDr7g4HPmntlU9
6+5+M7nYo+wqHKgMeVwiUhNOoh9dSmssdTfWuATUWD6UkJTdwn+XFPvliCiuXhcB
vlm99r99hImoJFZmjHNBwh78728U8HviGpJMVXQF63u/v02UCGjdkFn9Shy9V4vO
lL1ZhStePEjO3Dwf1iV9daKydm+4Ku5C8YxW620achnV1kCQZ9vhjZpcqB/lTV5D
e3fLkHaG3WauRG29hhUg8QQABFI45Q0dvMOxl/X93+UJc0/zT1PaEcNyEJ/al0b+
Rq3U441ewRU5easYkRtk/ZgGifeEbC8DUYZ3Ml0ik8xfNdo5QRZmSE86EthqYp3C
RvZafIRxeTnMk589+74dOlG0QpyVcArTJaEGGZzkAFGpgKLAsd3W2gRWxz2sBKTz
tQ9jpMYtfSiHvNvnozyJcWSGly1TFVAPMtZ61zgONINsPo0eOpiiyTxqwT7ftrkk
futtnnmy0EpURYqSYx0IYeDQdQuq3soqSpNvkVBacR8doEjyjy80+aOvdzCj3DM5
7saXFxzEuLPlW7hDs9NqzvNfSLuK1oPSSL1RPSBqwRDyaRgFgQIZ7NMKNPysAdnD
KgWx2jMJ5UVpd1ARCnwNjeegePc2nsXHraUmRmu0KE++d9qhOiZhVfrgZ4bCnGE0
gNnRRnofbYGZ2sEYlQlD6Y6MnAW87CahI09s2vdX9yRVb69Wf1u8zU6M+Ng8G8gy
r3aViRFbnzVrGVBHb2OXznqwpvuIWKYgNVmKbDThYFPny8S83/2hPRmhXQfBJ7Ys
h1CjZ7FJMlUJhyC/MtM9BjP/bgkHee+YqQ6p/CjpBUEi1143Xd06R5esQwcjoaHn
8gJ7De5j8QGy3Lb1ABUv+cLfSj9hu5YV7TDHXYJJaAnbixNs1Drs1GoON2JBh28N
MOanVbe04vJw7K3jFpKKfRYl8iJlT7mpsD3ukRqOaEHjiHE3Jx6CBe72oKGKizsj
EucqoVs3Hp/mRDNu7RBfPSutMkWefSsWhJrawib8i4oBVlTqO498kCDl51IGNbrx
rujOZbdkuqgHdP6qdzoOWMAF9aFDF9TQ49i5Me8qV7wYvpt8QiyIVXZ9ixyESgN0
VwT2N6xevuXj4v2+UN1xeyigiRJII44VBBWZuTKU8VFFvgmFieKAHv3J1almOk5v
LnvLAIl14tDIDPGeoDgiEqVBqZSzNCeF4lRdpzRYSAqF4ZsEj670XgBmsJUxllww
wS+K8fcjXlMmnntBGpyC8AOvTE3JeaCKsQWbn1COVQL8fqAYzM3/mCxhYOe5SFLp
uU+UgIZDyIMhc3SjtyErA/5xvNiuKqnvV2dfzvUvAjbpKSxoy+BqfCwJpLhH7YBQ
c1y5YNr87bSa83g2G2lmxAtNd99BwNhKrCa1bR4TIAbVvRQcJZD9xuYy0DKrpfSr
/cBAUgvM70cliCUw62yqgDqXyYJ8lCv2POQ1orMH5bg0B6McEYZxWk1sfCa6dOPU
WbrhYK9MQhHMkvCtwi3PPEfs8F7sVuh1Xi7VzxSt85/mpgvH5RYINMya2sEKdQKl
evDuFd4ECgqUdhqhI5ySVLQBltXQZnHwE5ZCjTJmyDDQ2ymyM9u1JmpsSo8l+caA
S6JL6kwKAOhkQNzvMcHFDQuQTouA7sh66hQ+BvgfuIOTBR3fLR6r6CzpsvCKjEC3
wIWg1ypGaUdJsdvpdjLgD4xO+PpkyzaY0/XnHNumKCOJMGXPVaqrDu0BN73jumWY
ufpGAtSLSlVjY4ZPzYR/DkqMeymXoIe2+npaLa5aJUIEUDJMPqV3QJ/VdKrwEHI6
mSMNiudkk1fDnmNoUJalgosOZ4QZRtq2l9e/vlcBiiCD/uTqoAsqk10phXjvMPcE
+elUsI4UGGwun38EjTmK5e4KNXct274hbRO/hxrxY/GWE8xafGOr98aGfRpsJLso
Zjouf9SL7HpoF2HrtdZhzgqtCkl5RxKpdX5X0fesfbeVFNDt3ujwIfIZvh5Q+Flj
HB1LoHVuZHrT2YHqFHvYNQSGqcgQalFkYNk/zAEVgMuvkbn/S5Q3dc9RWXY7bWJt
FVXnumA8x8s1zroUtERS1BIJnV7JmCT8hwGN4gZ37QmGkcLc8Z42aUyP3Y6oKG03
gUyJBsywV8Cm+dJpNjLctVrBiH1SsGxU+ycTNG32fSBDvFGPVfEHNC2H7UmhJNxp
mg+v6w8nj61OhtzokZUrgysHN68Q0F8b6OUE4koAFeCu7vfUgAzb4YzhRnknGxes
f1BGSfTKpJJMwGURHbPXepyuiQD80EOhYKYsAMUKKgYZqn7VdJw3YqBv9bsPdf1O
1cdmS6ectmVuN/9w8Rv6PKPCqBsAK9gWyAcTI9tkk+yWMt0iSucYVznM+14qK+Ln
QpSwZ09T6/HWmjt05GcKFdG65kn5CBz2FAby0aR16vHHigPw5c9gq2aDwm8oS9e9
RJ39/i2m9WW6QS2D4WU7oaxQmuN8xzuiCsGXnOIaEwrDYXcAOKUzEf4APrNbkV2p
c8sfjhVhgjybKdHAFGUUGxSZiukLJ3xAJC5FnCgjkNvITToZdG9tD93yg5wxMs9D
gg50ZZ2+VDrr/hJUilkDcEi1mogLldAJRigdaMWqRW6H0ZaePUtpsbX/vwQP0hxL
aZxaPFF89KpZHefA2bpqNR0tDrEg+ERQ07L/sek3OyWeEvzeq6yu+MbS0TNAOJ2b
yML0TRdjH3g/DH2yXziuZTmOnEJK+MmxRfw2VrGEC4B/gP8+TNx45E15lFcp1v2P
V6n4+j+q61Ze+bAetMFJZCogYl9Ml7SCHoNXrrZSdlkvv9AdcgsX4Nx6KV+jLgPn
Fm4lxjuWI/Dj4scrgdF8i0fhIxD0hNJhLLzaOGv9ep9N+JhpGEBlhugOE3r0d6J4
MDZtwbykK2W3VOzyk4HPdOumy/DgX/82YQlAsp/Qk2gpweeTyqNv4+S4iP/HnDCs
QCgnVVmV8OBSDuXkLyvKhjsi+m00sZsVXwMDHfca6vzflPUNrVP2RCUcK/xZE6PJ
jB5BJzUC0Rs5MP15NujjXrDzxX/0MStM/Jz8EkJWIim3dPOakLrROwY9hwWP344P
qJEjwLCwgmiADU305xBgNyoiD34kNgK0gLqha97CfDzCnuTEbmodDH4kCMm08H77
1cHDVZDlexZlFnURy2/u5ubym45fHyCgDLRnBku7wu4pOpFvgcLiIVydXDhChNS2
rnQvyKJM0y1fjanA/bdADd6IKzk8qKm7QDw/29MrgOUK8yuYCpR4YRnAyaAg3hLO
xxI7dK8cY6RBmDhRUg/KauzABUYdDzwFfCVwUeongkes3xFX3LJq97TSM6ZqBnkc
h77XIrKiMjJmVsLX+z89erFzbgH1kt60l0o83AxiD0ySQ2RDIvJ7DzEX0uxD59hp
r6sOTG+3R9dGxVC0sZaZ2znfTr4/4bG9kP16h32kekvj6ee0dOdS/xXT+l4s4YwX
1upgn7gV9qfF08r/u615+s2m2jMh71L9R4IK2y67hUSr3XgB0i+xAgo8KIs9NHQ+
B0z+cB+ChmelVeNDtfNaStnnnSdt4sJmEdxzoYPOH2oGZy+C6AT2xHILNwLRPkTH
0IK5HBvfEEzld+0K5aVAeXC1axZqUCDbk2LeQkq477QOvFqMmmOPVqoDmBqfQ1rz
MuQJtSg2ZrvJVoQVaiSK5XKVMrDefSaa1+je+twT2xnKeGRLzjdudkqGRbnsKVYI
djIqG1WjBtyDaNZuCVjf1QHR+Q3dq28vN/m9snpR1X5P45VmIvGNQJ0UQVcrMwoo
0ETq3GcLgPXnIyztdEXZngzasTUeHalpSwq2T8INyCGmBqOhpg0T3cA1K4NlglTA
ffp6Q4mXQ9B8BB9VpNZr/+1a1VVwe9lye42vcOpBhJNppoBEIsX6hd5/MrBx8FOJ
5NZUf1PNWVtH00CFM0NGXKqDE5KFYKNqgvPAVL0qlOKivq9rt3TrwPHGKWIKGSUW
wlZ7MJe/YES1sImYw7Wmcubhk5DSkNgcIOtmhT2XGJbm7axNufEyOV7MCyIArFUY
k1siHTxjNCFO21uGmj6OFT8waSDY0sVL+NYy0yvlRwuA4EC3KBf+UhwFdfFi+ZpA
47I4XJHiXopVz/zywv12nGI/33iw6hkSUQRno/yfeHHkiyMnLMR7pStbWzUuD4vg
VUlwfS5iQQW3ABLMtO/xKlDnWaQUR46NIeQeGRBR3mTJhrTYgOjxqpM2pRtVOWxY
Kqkvghe0HN2Uijd5tyn2vHbJ0UqgC61NWX1UKKdirtE8x4rQmJaLmh3FWs/47K9a
wO99lECTJ++ASW9k8DhbHjuXDkQxSiU4rI8B7NBLS/xMrJfvzr9E+tnCPm6SWCpF
tdQ4EYEOO3PPcZEOSnRL9Q6XTThP4v5mP8+dd7L8hG3eKO1QAikgYbQb5Cw50IUY
unk2WF4QS1GQU6761n1c9q3QQuhYLuxEuqXugG0Me+IYoXZeOvQcZuJI6oowHCus
SbrzBn/gd6wBENy0/bCYJ4wnmZp8br0iYkjcpXZSy25tms9F/1fQdONpxKkqJGW+
Zi/ssDIJrr/T4E06RhPjH/ybzaY2t1K6B5ydDhpJk31D3Q9jUwwyNT9DAAiNnerI
ju0cI/9uaDWFLf0qcGChNsjIG+uelcz5VTcU2oAjYbg29KsM9U86xJV9oHVp6TzN
fbIBkKupg3jpKKi65wMeyxD6/vcQD2xZ/QG7TjBYpWpPHRpeMGzhyhuf21Iqziil
NeP/KeM45YjIy/wLHBesxLYyj0zoXZt3/qw8AkFfpdDH76IrRluXvTTvldOzb9F3
y7eJtF3GxDs1B/fZMx3XEruNpQZGtbDaYvQ0GSPz7HRS5JdXiTRqacaB7zRJvrOO
ub0ukKsE9QQFGE82xBaHLxYhsSYp+2dqn5mOMkCg5s3g8SDdfNKTUDIaqvNoLDgV
t/ZYRvolewb68e8m8wS+uxNVTJOT+hbabc+zdHmtgmxoYqIk56pVD+Y9VRe3b432
Jam0O49OvROIwhPu6Y4Jenf5GVnsw10H4V1F+gC+mjqNFQc5hBoOhq6MFA+oG91m
GqlyMq1qi8WkHOdi7OQWKx3N72vvJYhntmFoaiLDViDio2qK6+Ab6H4UvwPB78y3
3mxbSfwyVsPpzg80SF907VjMswQ2z+0ljo2fQsrYDxZPym+ygbzrfoQQImjTQNnW
MO5YssKT1hFhnDedrMZRON1YazSETF4r3W+eunFyrB0ZMi0nRtJqkakiuTy7YTjD
/miJ7i+Pn1YO82N2XobZ+Ep7I3JocnhsmE1DHKeTPw9JRaWsllcg0GIJvOJv9Bd/
ZSkuNRJr5HIjNCXLnw9oHzCgF+Dhl5Fr5crhXUnVTogK8gsFRUds7/eJoZEfFamU
7lOmGBeBI0Id9OBxd0dmlsbxu13foK1Ls9GbeA6RTk9ux5qlUkBPYuLjwggzngk2
tjfDJmRKEEK4WrPsK1d1pTl7Z1PJll9btFO0jBHaWTc3E1V6z/TuU0KemhmD5FUb
XiwX6aSrGxARhEAJaMngkxJv9QtMl/kcZ6KX5PACjQTwRf87zrcvSFeSNBW7zu3V
QN3NFgJdRfuIvvJ0m1Jf4J+aVyAkyCDQXqdjiAwGDP6mrc5Ikbs0I0aogChkfCA3
XhO5cF9okkZntbvYQ1S524zyrN9NasLRKLXfV5WnJQsCltndkPC3Ae9yhLqvJCRG
URzPtYGPmrfg3lJH97XsLXM2TVINe0ePdjKV45Bj38BErdU3KU0mDlvg772dfhTJ
4hmuc9w9akmxTnulCQCPGF4hH3C7wGAPF/A8MbaZwX+bpOPTeEUPIAl2dVHLxXex
WEtF9XhekaE68U1DnOXeKY60ZEJSpKhDmO8XGxLAqIX8i/aHD38EWiGEWfRIKDBb
2hZfsbsQkNGfu47LH8P4EAMIcIEmo5sfwqi/QsC1xBAHr1I7/RbJvmZumM6TFSDP
NbbKs0ktaRG1La/iSzk1GXcKYYB5gPFlRDvnagdrnAtRRiI654Kg+zcllyEkX/Sx
W8S53M5JIRxXb5mcU6oP+WTPujjS7ACjGLnzEJZQ5ZqcYt6RjMKWi1vno09pMnzc
JFy0MgXXFm62I3scLlnfuvGt4lwNU8NaTsb20LKQO3OksXk4amx1eg90uQX+tEmK
L8g/kxoIoN923+UtELBxAgBYlbDD9LN8qpfgvTXvfoeROJbEqJb6tHAWC16w2Ft1
FXxUlS1NsvLD2NuLXA1z0cHfGuR+k9SYTqbEgHGXhi8HHg27Q2iZPEUoakjqcNYK
nhCK8azMR4JI7K6ILRsJzVHL/XCnzSfYiG+v/t8CRjruJDyOR4f8BCsNMwhL/GY+
0qJ9hUxTqic+WfVrCxS+fBAO/ykYKE5aBh/ZvS/WDOzhLxh00T3u/cTw8WD7Vk9k
CoflHSbHG8rSW+LqcC76A4AMDAi+Gs8hT1tH5mEilk3WzMkT8LzRGXuqkbjbxbG7
ltyCzzUNnVjWtmVchCYw2gWOl+LQJelGWIOYLuInJAcVIcU1cp5u6ZxSmFuk3H1J
vDfm8mdQ5MmNRy9oGIlRHubq+DnWldJwU0C5AxNRJfd2deqsSSMRKguNaL0Ejn6i
n9Y83feR4FaClbYGMDuF69OpfdzEjb83nYF7J7/IDd1tfQmHy+hMS7JXzEvYo+Tz
tYb4M2C+UhrB3neLXFXHPkQ9EaFwZUyxposnJ1i2Fy1ZxJTbaLC3ZzY9NKZBRncW
V3BGrTrWrVVR6E8a45GYKNdUVs79RIk4NogDVSrTyDxCxkEy1Feh2HiMFbkEeIFJ
TTfc2yFXnpaAXemGRAFWOQHe99uEkQ3ux+NZwb8+THxpbqkw9GMjuB4Gp5pf1vhp
yRB0SE16Qf8VPsxwEvMkOGY/59E/1t/YOeUxmbL5z3jLwb39k53DzaUzB1LIUDfx
sfxRl199c/nA5VQCQQFhB9dGubAScvAv4xz+tSIulLVox2WY7XhOCQcNWxlnky/z
f9e10oHCGnYJ9YfGgkaJFLH/x8PnNvj3hD6Uv38Pzq13k/FD4bFMaWOM6bJAlsvH
0XEKSdAZUnUnWjvMxasQ/SxUeVv8/VhH8T7ABHbFdFTzHSVy5bUUYorerqtDH/k6
eICIvPKH30FF6T2HzDiX0Lqw5MnFKLcU8IKlN83q19Z17tLE3lXPCNnoNsumHVbF
YtvVm2Lb3ZdidV7hCm9D70vpxUZxLuRcxaphJPJ0TbVbaUy07TYY3SJWC2VZpq+A
QZn30wssAHPaZFZlnnleD8CxOw22fqQIxk1/HvalbrZ1lqFf6/Eco9ATsG7y10yr
lCfIixBgCJtjCXDUyb/cCNvjmzz9I7yKQ3lzG0XRsAAadHYTdqsh+pPXrDh45+bX
P2v0H4mCUSOmRx8wdfhhkuupUizooIdKeVv7UNqe7X9Gg+Fd0MylAar8Pgb2bfni
tkiEH6U4WqQu7VlpFx2Cgpg5zw8L+uL9ZjoSVEcBP6UTzrWbwjjSqXrUmMYpjiXG
N+yys10GLy/j6nVJIUU8Cgn/DYkaYmNiPNhZ8DXiAjL6ZdHSPUGj7eTOR5Pb0U1j
tcSIk6X0q/dRSZYyLdD4ZfgHXcleUng2ZugVKChk5R4m1BSAqnSWy4KinZhoihcu
yBVknKeDlJQwVoqSnGth5a3aZLX8q4nFvdVZejJSybp+3YiSg4Lwb93O4BTWeo1j
8WdWGsW4GRgtXXwPGij2EfHRpC0xPr4UvRe4vMet8Y5xQZz9WFLFtS27T50B+AJ6
q7eB78A2CBwk7EU8prkCfJct0qM3oPYSj9XOQQtqTdIKPGMlhFq34nn67hQ0sKb9
BqdrSwFE+v4a0W2sHIu2VDfT6BpTvYAGhYywd8gFXxs1uuNUv4GjBQSBk3MIgQKR
bohG5YhSKcJU/pFGDDhCYk3KESZs+35/8rpE331NXAu9UGvk0midUwhCPKWG2oJN
gQxFdOGHXOKxpyy2/+jTv7bwMr6MJOo62dpnUn35/K5azMXvy1FfSd1KXj4SaaWK
bt1A2GoOWtLRb0PhgXLCRV2vUI93TFTA6ZAxoUk9vKZ5YNGk6/ODHlYRFt8zTlQU
qqyg7s09lirlsGpVXtmKanoqPKX4hHk0q/GKm0EsYLRMmX89CQT0zYV1v/68rpVG
tc1BrCuzSmGeNrUVQ6+O645jkM2awxNVQlJ7TRe+oh3pFceP5erSTsByRJPkxZYV
iYJCIPxJk15fYAdx+bC9BgWmvP/EQsM8m4DHciunwLsOtpLWY32Mhhcl2+Sn+xiu
iCWOhMOve5Lw7a8RsPw463wDm6Ok8EuHUpDOHFw/7V8j8xBXLKH+bLy+B/waNnec
ZzEnOCrIBoguagic0KINWMZNRtL2bVKmS3KngqxFFOQxHUN0PgtiyhHswck8QI/d
fPtlhmXHJfxxUdWfMrb6gHjPAJiUGGIQOtLf2kNuUCZPzdFExb9zIh3Ug5Xh9HWN
tzQqB/kCUrDgYA0QC45Sw3k1mlWgxiwnj6fxAYuMiGf+FB5DCRZm0D9VyhhwEmap
tKXExedXjlSnXqtL0Sjbnfiaif494E7JRDKnzbz/A0fZ+/B2CggQczAhWNyhpUpu
L7Xuc82D319NiKQ6M6X0FEh9VEtFJWQK+AH0jhHi6CU1q3XHJmZtLrZgUw/vDay4
SabKudfjJthD3karUb/QkPBmcfeJMgGwURVcVaxys7BsGMFmb0q6rbXEfym69wro
4cQCglMiT7IWOIjOdhjFW/Sy+gacfsIZGaB4ph9R4gly75UMYoQmZGaMyK3N1Bex
GJOOM4FBKiz+fWZQLkUFoZnwhnFxEc2HdLTQmuWe2Wsg5XKcgHvoq3zMYGPE9+ZD
tDAXe5dBF1TgvczzuhaBnBv9k+4drR7HkSGFltHaqEuxsjGlsIjd8C5Vz1dGxE01
by/SVjwwvoTWeWmdhKk/RjbINr2z7leuzlGyjyeZTBs/pffq8mzk0fnoGxb0qZ49
fjjbJFGgsv0NQxVbmET+MIMaF9SQZljn3fuXHB0dvttchJTvKY/0kY7E+BbFBM4o
wMjYAM3s+uGQ2OaGUcPqBSbM9U7Bl0mMhHNal7cHUijQNmTuRYaRWCaACQI2IBEc
MrGphYMqtB0JfouLGgl045t+GRCeroLyBBWrcyTi9ScjebqIUxJzTbykimjZsW8A
e7NAbuQ7x7gqTqzP+9BtjgPhdTricMTt2sD2ASzZhPSUUeu69qp+xt49rXSODqHK
iJFLpI6Hvtjei4GOWZYGZtlbmLeQR+jIM9L+3hctvyI1C/SVtvRLIe2vsmsr03PY
HR9L00f1C48RwXlwmhPMBrNrgcPCyxYAyrendxjEbb21Z0eX4P27YXwpUvHKsf4X
OJlvrx+5atIXfJRvTaya/hBuWc17w22cpMPlDg8G8i3Vdya1VZrrsgjCAZHBbFi/
ek4oodWo4uc0lLEYujuImgmOrKzL+KQdN3ELk8YOx0TtOPUY2nT32kjMWGDWmhGv
tLPadV5PXMMgkOLIfwwCcRWbl4cP1i3xr3Hm68dLk8ft0SQKVq1qjyRCm/FZWH4c
MaBrPRXycOmd+9FXc4K3Zn8I884fDb/GPXvgyQAzUtpipwfn8zbwKGKKuCTGWjlT
vykUpzq6dC1x5WFyb6wklC3KxCtth6UGQ3YmLzzC33OaE31s4tKgHu8Z2by2emJy
+03zALNjtK/d1YWbvPKMcTjGvQyivG5fjX4pZBHIVneMpCIFLonDgLU1oEMS6q5j
3l8uZcm4gyZ7hCDhGA9Kd+74HaH1CFIh2aU3zN/QzN4DPCsZTYx19WW9dKdyfnka
P+4d+xAWt0CZzIAr3zvRcCb0ANDLo83zTHCjRrvC20WuoskwdoOc6QluGD9krtw8
UmdrzUVgfOBceM8fSFc8IfzCOcEZawdSJ8OGqMsjKbVzgsHT0E32c9dru13KV+5Z
Oe2iw88wyDeB/Qrv7fItn/dHVCB6jj585A50aQjChQCTD+c+o2hr+ItOsnsNr6v5
jIvLYcCyoNy+AifPsS5w1hBgC456EhRKjTsQ7OspvQAysXqwqCJ6cHHmGdhP7BR6
iII2suJT+shjgfO0N32pTg3q6wkMUTF0EBeXGAuerzzUH6J8/h+ZzMERakpWU5KW
vJaU9pq1dc11USlEQJaNMGtqnC2sZwwsaWfxn1Sirs9+WgwNrn9ZiIBLv6Mg24l+
RI36vzFLHDgHv+y8i1hCS8oxBJbLdh+EmRvRPvG6jE4Ugbz1tdvJ4FE8/QhxgpOg
esLd0UJXrAKN63gCxlAGgCP4mi6wZJVBki8zKyZCtmvkPpBdffZkvsIUb32y+VEg
AAfLl+qIVjQyBjWEDbOBjI1YqqtlvqiHgzjY+NoQeV/67RVxGcBV/o9OmuvfYvc6
FmeTzs6XCYA64FhJIjGGC9ziMjxzG2K5n7UnLfU3jkBON1dplOnf2JoksjXB0Yls
BPS/hXcBEZ/mDlBwsOxAT0/7t5BIjxR6IB8IE7XGoxwCr6NG372RLJgqCk6EwFJO
tjN067fbac9PH/wgNiyN+smayqb/b8d/6eXcMzGzm65E0uf6J5JUjj9LjXBvbami
hKLX+CYLCaxtZRGMHzE6pFvzp/7lZmHpCY3klyxBwKufhlA3AXB1YmdipNnCjA6j
NXxWcaSfObwNtnMTtg/WOtJiVcy1kCl5OANfK69TfVTQB4fZmJkNIRcgXEt1PLnn
3aEZWZ+sOlOBvTrNaP2OsO8YWt+dEnssXWZ7wlWl4bkTsPzeI3i6XTgH5+vtqyh4
LOtqiE2LZ/samwVc0pZlTiF0GB7D6/7AouZW50IuimWzjMbHf/T08Lq7fPjQyenx
GXXqgAym/VlPduGk0xuJSIQBNFTj5hQ3trEInGccFqCfIqUeNWQfZjjYr3CpQRYg
maw8is6eYPLpt02552X3Sgh4j1XfiHDa0wzJgH+e+RbyRrp8qnj2WBHbSIMrMC2C
BBdnFurQo0Q3CUhKIQRsmCcITUbllQmihJiKRJpMCd/XfpF+1lPyr1rZO2c+86Fn
tX0b2wxe8MI46QafKf7H8Xpw+QH4iL+BMmxgM64eSjxgB1HkCd70jG/3YlHTWmu0
/Zxf+e8WaK4GnUy1P4J543wnrjDlVCPcZjkHWMapDqO7G+C1x1FLf0LM+s+R53w6
6RUtUmS0iW3012OkM15AA/DGsJ9kQb2Xoz8ffkXhyMln7Sorwik8AnnecPutUltp
eCxuXoJoSw270ZVUWVJ3ownG9vX067FXaQ2LkhLiMP/eJOOY6cwy0o6uSOAbbxsI
FobH8VkZHYJ5qXj4mR/lQcceQOkbqsXOwap0o4DAiWHKjzXu8lqGisNSWfD00jzr
YtNYpNU0xRrzKXFyGbB2EAm5uaNUIe/HEjkG6gZKK/kXmFKf1VMfEd9uAwlyU5HO
C3I9aDktP6yTsZCIuKGBwqHYhepPlAG177IdaMV7MYLvNFYeF3UgAJ4iAd0IXylN
dt6kw8SVNxxsz8/0zdQCiaRY9CKAXMLAF1uDJFVf1U8mI9Irq4qssjD8HT7W2v91
3DK5AVRS/+oFOiYKH2arnepRdPA+57qUDAkuTMIaAgyGtkZpIsn2u+zNLm+L3YzD
jqytZxX0Am0NY9WMLeX2+F2a1gGkPtvlT0TReFiy6dzdkDSk44TrZUIbaCKf24LR
mc6M+76/0Q/af+ZQG6pzY317iisVF1+lqkfmfJjmwvz2mctQrupGmjguqouI2djj
HIFfGkDGRnYUIo3isz4xJ2H4DrKfO9WU/ngSNYqJD/RPkKBZCV+2uepMxF601gRc
drfsL7pmX9Ca4GMuw7fta34r9O+pe5jTx5U5Gjrwm0f+CnKbtGZ1nl+6VnXWQw6U
GJfLox0mkzsLW6UZAA/NGdcl8OXw1f3BV//Ukxge9zAUULPb/u6IZkeSNmCKSysI
ciWVVZtEwPO5mWyzmI59GKZHZhLr5A12oHwQ6VOceprR8cntnM7PgTrCCpKCj2H1
WqJ8pBFrXxwaomKVqcP+ldxY79RevWjl4f5nDtFKLyTBEKsHTWmytsx1fvKWGofd
HdD95LZtHMsxBgNkYsdgTOb9fh+eaWpRoQXOErvYG52GXh5VkzIa/3c+ZSRvEabu
DfzJ+g5JYIcBv5ViSkMxIJE/YD6Hpp4rkkS6zMzzK62OYYyFmHWHZmu9zOhQ4hkZ
lvWVhabbVICy8ukiTodaLKinEu4WaJjA9NC31XxgIeuRkoEu8fW42ZWXzpJstjiT
pi7VPkIX7ZNH+wGigNbORuyY2Ri7CIfZal/IYSfoeBd/K+NyQ9rmO1jQ6JpNosBx
SIQ+BhrP0BR5ql8mIY7d+bd1Emj53lUd/MH1+x6y0QzVRCayBhTe5mPJfmEuAtVn
GoIlc7J5IyTZ6ELVwhKcN7GWaKHubIEgVMljJJ2TJnoYEn0eHmpcwYTLvCNl/Wut
yGjO900O89AhBP43DNHUqgFiV74f82i15LCDzy7h+3ojoriSTxiLgDmVcqyEa212
1WsFJeAnZDfiOVlxZImFsaBiHgc2xnW2jQA33bkCGpl+wrZH0TkhVNuLsKLew/7K
C80bdddgPmFWoo7U8mC7lYX2i8xYqPAdLD34FnZBaXu2xl33FvQwgnx2WGUKAHd4
5MvUYo8tkvaxQ14Z5nzyu327Or9KdXiudCIIoD1P42Kd7Iz2/XJx1aSL82iMrefX
+mXDtxDhEQ38Wi/VuEZZhaDe5ycP3Gyfl02trQU9f0H3r/BbBQtTT8asATfzO0Js
m5rNpIVai/uyY1xm1sPYyiNGlN76wG5+C+PhUNiYp3girH5oL3mwxU3YwraaKYfi
nk8R8dt58f4JHohiBUmtHa+EMkXfmrQ9BmJ+PTFbos5x9UgfJpMHtNODtOwLXCRx
lG7Fg9/aTb7R/zQ7BuEx3FAG6uN8xI6sxvsrT/jdPK0xIRg6CTfW1GiDT7SIGz00
IpzP5Z8IB8EjzdryPgP1RC7a+mpTVigkLViz8UoQ/JFLHj7Y7h8oko8uosmQGZVS
gSt0rtaE9TlWBiWBNvMsvDpO/c3wbOD5O0Cbr2qe76dDG24Q5rM+r3ThAj5SVhyk
u86WkLkp9heVDaCdbR7g9mG9dY0eaOCfNxymL2BSSDLJYXQul/L/KTCcbqdYhSOJ
cbEF08g4+6b1BGPX3nm9lcfJdfjGBp+jmpgUzunJmSzw5wy15lx4/uyQ65bbqCzT
HCqMY6x38pfM7gWyzVPaQanAl+bKRiTxenfDCyFVb87Hfbf7qytiM7LOmrf0LNWu
TxKkOlJn8s4mpO4CpgqmUQpltSNBe0aqVGeGGvO+9uwQ6n+gLIcFh0rgKpGTNWdq
FTLsCPJmgQumcUzYWSRNRa9lv7h99Y4cqbQfBHt2i2UW+geIFGDgx/2ZhsQM9u9r
JtsqhZnckdfbbUzmu2KKZUZVabdEQclBGlmXZI0naqJBmpxcI2v8DgOkIrqblvmi
rEslMMnUjcIYXlG5jwP1aChI/wm3rkndieli6Kti/FQodBzQpd4cT9c5evXkC4pz
kId8C7TCcVAT7+i5Pkcua13SYBXHjh4VbWn26/OAC6P62858bHblOPG4Fb2CBK59
xqCULAxtkSjNcuSO39IiTxj11cg79/RkN+P1ahPSVOt19AEY+pPnI/b3THW4M4EN
YtgnUobQhhwRcDEeoFxBwBPVAWc2Iz9K6MuDePaSF2u8AD0iYEz9z24eZuDgEb6E
7Ea3VQwkAdkEzEdnSUiOH9L7DmHyP2C6A0f7VgHHrthHLAkRE6s37ZnKrnXh3aEY
wRoARWN5bVGg6MrWXZkV7TupZA6Ae3nAuyqlq3EZ8mTo4/PbnlT8W5KBj4qJmHae
Fv4O2HTBSimlNpmNBctFkvLfKAh4FKzp4r/IG6hPEoc0EDRcQ8xg7MIYus0os/Cs
WXbz8P7GHJb2fcrpUE7unCrhpHUJ5y6hrXMBoUtGxq3BMmVGtL3YBnHox+KixNDa
flN360+RXfENePLHTTFKI/pgQPDTtB6hkAwES9cQmS2ja9mxeX0dOxyhxcUuYVQi
iKEeded+OSYVh4a98UJpb7BdgIkSjhQlY9ti5OoQB7NAVj5+GScvNS3j/dSXOGZC
rR3QWTF2uf147xnzKiRcum5FSIkjgr8JUlJ7Fjx8PkpxmGADojGYmGWfLBtIBZnD
zIz2Q7+FjBLuyzlukFTlJhuwm+lUkbOhb3de/a4lwUz9+Fp7lC6wUfURegKuE7S2
dtaUUHJ34jCx0KvRdfvvl2kYhz//nFXvWEgeQ5Gk/5cGWHm9AONkRNx+fSIpx6Jd
ZQLXO+WihG/1xyZ7AxVS4+tew+mSLyQcnx9M3tzV4peyclwqPNijWfMRuBjVIKda
Nx5GkWTXkr61ZNNuD910D3Nmq+f70y59dhls/KIUMK6RYBJTEQrRwWKnT7q/veeJ
gc93E4R7u00LqwMyItVthJZeX6qILUuhjtwTZw0zfjic4UjzWtyh+vKTIfLKIsWe
2ILkSU3YovuHf+VlYeab3KSf/TTwx8ZVTE3AZ2Rl5wMI7q066Fo5y7jmVgYPuUzO
lbnqqX2SBjGPQJ5Qhvnzi2Q18vojhVuUyURbtSxgNwE/QoGgkgnvOr54oxItAtK4
wbaMHqzWy3VYx+NLBg6PrBdIaNf1oxrrTOrH9mCzv10gQeFnqlViACwxo88KrVeq
wN46yv5sOjrDfFvnok1pUGfugYDF9wrY/WVybYRz5bjfCyJJLIO3dOHXiDoRJ4Aw
/KBCgJiacVaUcmOmNhEnaYUyDGjEKk/RXZt5oTrDJEJnf7fUn5eJjw0HV02wCegs
nG6RGVwHzLKzeS7xS976MOUavFXfAKrWXMYX0Qp3gJrlGOnIdnDNwaP9bjpr0gxs
vFBL9DFvhttc+siAlKZgQsqkMGhq92OXueWCNqj1QFmZyauHaBxGI0jk44rrrYDZ
YuuI65XPRq7TMv5HaEtfWssMg9002GzLrDkcjORbzAKAhwc2xuzMWeqHvN4DMWd/
yJccioK6lg42B18VvEAEXUHaQ6RWxn5BM1z+ODL/DUnM+VtXwHVpGdr0dHcAT2cn
e6mq+N/7+8xZmMCw9w5exCeo7y8N6SOwnSvJM49y4ZxApYEpCPclj/ds8riMnG+L
yuA5I0HnpgzYN8elWBolfC/bANHqNetyvhh9tc1YIBJgWj65/+S2zLx7vJW6Hy7N
LmExzC5aMpqER9Afl/x5a9YgZ7/H98D5grd1nKk73FpXHKaLFAExb3Bj65beAjBj
qEQl0a/lHoQGItHAzS/7rlg4cW8ZlBuc/HmgSjbJ6wkKaZUdu2A+bt8h0GVRilKh
xmAWEDYWjsjoWAmgKE8G0lssjvaiHIJDQIYbOsfEqgYCz3FFrWZFmjj0P/P+RxEu
iMyxUZRJjMvSuMZFgw/BhYnG5Nf9Ks0c9zWWg3tBV/fyjSg2S+ByX4wm8UgZfEa5
BXTKPPLuIbwSESMghGQrFofi1YHRMUwUUx55UweYYXKedCBfe9HNfF/ew5FGBGvL
jnXpcip4KPC+5Qgd8Y8XrKU3vpglXRMZh+/lQ4C720YPs+7qHiooqQPw+H0Frp/q
rIBuIXbhJMc7vKIuW6TS+b/X1xX14qoQxc93l+10ZZRarVvwJwlVWxXjVAkhRFxK
eWfvgByXsqaK6EvuPdWaBhGf9yxAnOuwmHSIh6UTFTU7cZMSa9CIZhjs25xqs0FU
wN0aB7oYuMXuVQP+rSIa7a3VJi9Bo3KMijuaqkMXVoCMJ6mBVTF8F4lFbUXjXQSH
lteGjjB3T0z+dPTRrhz3VlPKZMklMe3g4uWu81tKOkIKoaDoUfiBYQuY6Dci9LHn
tMWBRwvIFWSqiLQXVUFX7LyQey7eyPFIj//71a5IBXXuYj7dTc7ctM9FX/i2Arwo
4nS00XK/ihYFUKHxxrypA79D2iO79BeWeRFvmD+6LHuUCZcieTOIIpXdd3DsuW76
TPEIu3jYn6rBbfHdVpuusuMRuJxrlHAdcATBiUniRJ3vgNZPmIhM1DAE1Jk0elGH
N+jteh6zRZm3ZEs4YfFC9thJ7kdCGz0nwpo5rngnQKVITtvGcURs8lQQe3Bi6Bsv
9ANSTMnE7ZutuP5QjDx8USLLKoyrWgA9sK8AJ1SQJTiupvb/whOH2X4khTMxuBAe
UdoP34rU8cDTHsDr84V7Rgl2GZuq/q2P13gKcwXoS2rH3OLKps8Sr0Lr4z/dhWfW
0xLV/XQR0d4V3tinFYVJkMkVOcFJq75kdP0WFFU7aWBLiyfq85EA2EDxLb/7jzqn
3u0Z8F6naAQKZE9ue0E3demm1DYPbH+OFruAO5xBxConmkOOYm8xQJKRFb4u8m3O
Zv7XEj70lHr6vhWg8SaRwBm8I4rUk0k4EUNFjmqQg1Uvy5Cn3Moj6FxlvB3dRlvu
I/19sr8hp/bW/v9q2KEAJSZKwm99ldGQvMdv0dAgCxjf+ohKiWbYHMROEcXdoG1n
DhhV7SZ1Uvr87iCaslKGJxnOMIVwox2Le9TWu3thKzY9vOaUCj2OuHA3pI3kpx6z
iPG8YbMLYXfPXxrayjELtdq8XLyPBbI9CYrtfxrMLtpXMLeGgXW6FmNzVPAG9EKC
9tUILz3/bQSIx/zv6WZrzEcfv6m3XFWLXUz9SFuMM2na/QFyMJ9BhEBhJs22k6dX
wqPUi6MoTvWsU4mgzFrx6kiENNUgxJ07/N7StDOVmJJqxYFWp72djYdKrBvwDuU/
4zOelBlNdeQxT2oADQauVmIdnCWeQfGAUE4TJ7IrySYHpijhYLQExc8BZpuC8LXI
wm6lPckHX5p0HLARLjBcYtS6G7BTSo9RU3nUHUdU4kFhKEXqJrFM8y/MG6AcfG0T
RACWQ8Ry5X5yypqwKGFwGrQ2qUYbhAX0ObydiY6g5RT0TrHs3jHKXF8oW2D3zu7Y
92dK+0mJnIZApTm3HKBZku8U9J+9fx75r7mpWsYcDHTvpiSpneSJgSXorcvurj3j
NQMgECqJvzQyFw25GJbHHRSlFpHbMtdzruMCExNNtmmkwmWUgBw50UeI79Y48whd
9jCX5gtVToFrwxUNwEKKe/j2UdW71peHfOuCYJlsUEiuxLIwYB5axbA6RZ2Ld3q/
P8IW1wlhvdNlKRjRKniNesPrSa0EIP+SKkqnf+xTV3iwC8t295ugAeAyzQWppNuR
sH0gZDRnCwXES7M+A7y4RAndTIa/UqlRqQzElve4wde8wa0XrN/PmR6NQR24XFvZ
Wsj+aKqTWW7kEB1DIqgEA5KkNj44ZZh1qw1DGON4fILxsDvkjZgGSAwvWb8W7c33
pezeRatyAVzI/fBAhWaUBM2zV++drfd4d8iFws+A4+Jl9eDIo4oKX9FV9UTZmlHK
erlrtmMAxQ17olrqgqXsPJ8pu5ilsqGWkBHHZpC6DTKWuvJfXMohykaHMH156+OB
9ajz48VqSRlHjd5Qo1rpgmragLVSjC81JMDjd4n9RB+Zp6Ifly5P/vOqnnnOKeSJ
jLE1jGung0B+st7Tpiap3GdcEvRqodm/BffapGVxVsEXJCQwiRcZD+VpzVL0LjHu
l+drhAI4o5bsxSzeVhlWluQt9GxO682id7gnAGpkjkVxcCi+y0bIYJwluk6ZULsN
seKMaE2ymohymw02eLUiQTkYDK2bG9SpQdPPQCy0DzRCofuznoW7bRgBrWJtqsxH
tyuyGvHshBuHQOANrGCUFSL4IVzMCl6WmcmntGwrKc2YaFYwRVCERewuY6YySDmS
zsKpIK3UZI4uNNYasImAuMck20FccL4qhhiZFZpa9LSgXtlZ8oWVlNSWbbDghyAu
W3zU6i8CUuVYPqUsQT+kVzBcXFuHfVmGrCDnUCkwJMZxDLnzh57Q6JHpNdtLV8Li
S5g8isebCfTvxcvt+Ww40ux2z3FGnpfXN4XmbKmYdCJuCrbq+BMkXG6ZQyed0PWT
z4SXu/LOTHabd/Q/WFh+7ySJRffJKXgmHiAKxzkOZGgdVRYUh2g9g5EWLSXjH83i
2NL/JrJbl22jror2me3EqnVxPBzvWzRlJhTVl5uuc//QJ5/fVPJkTLTzGNu83Hm7
LrImMj8Gpg9Rb7CmaOYVGYy44F15rxELXQHMWdF4LnTxu+nLvf+PHlzSlMb27ZXB
903VTwhpqgro97k0Rt2WL0L4DLwAWFddUOS7gsCSUm5sowyf4rD0ihDryVSRbLbQ
mEeGGOt3+Mnk9wnKvNWNkNlyT0dCon1bL8D0EEtsngxiU9xCVWP3LpYCDvGfbyyF
gt6/xBNtdfgR1eHK3nXW6KgIu3EaFxleOc9p37adr8b/WZ5GmMzBNHXl24UnOgfN
ruuAHXJDI4kRFpVWDmHPup1Rs/bbppKmrhNp66sKr3/1qtRThidJg7oYyQ8lSQ1G
MzxhJT+askA2wJ6VF9xBktGsyABaMqXXRcx2edOgn0rP+JynehxK8P7idY0yNVlh
2aXrMoF6+y2GtH9j4RDXNQ/DhYmLWlZoTqDd3f7sQS0DCYWTGH0tGNRoXbsNFazg
fWcSxg+9VAqOT0szsbBCG4U0tsck01j2b2P5eajfMYLslGHdXQuoIRyr0UizqDUE
Gwtrr73NCExQAayNjK0vC+Ib3WvVNjO83vRCMBHSR2fFYuHr5w5IcDJ63i6O03Ao
c2TCd9+cLN21FnY0kzHMF8EbPdd+BhmFZnL8+C/KNEwCNTeme7icOz/8spButJIi
0H0zQjxzU6PYlk2Gfw4P33UgOh3n/foqg4Ynv8TuGhszqKaRC7ra4bHIfDXQKANn
ZHGDwkHH5LSTpUwtxjDx5iu90Qiul/r/+VKSq4en+4J3WAJ7PweQQIBUmDlRjAQd
b3s63pWCoQURp7c+xw4ZtKpAIGJtN29Rqfq02VCBIWpUDviCQB31RGWztH81WJ37
lP7QdhHQQKlc1ziJ21ulMF4KR4ElUtKDpgfMBIK+NtmpTeWUUq+f+Avc4jHRXPHL
u5V/Bc6iy6VZJQOTWgqUryfY8fUVQZPnNzp/p174jNoEiuKak70w+r2EILrUt4f/
yduq0AKKIdUTTqqpSLjCowCS8IFdW/f02kcmiHcCRVBtLrNeO1MbcnnZCt5sixGp
57FfJvYAQBkdR8PEcyZIRi+zBQOSLX31E1dUUQom2b0XDxwROsbcs8M+/im+32NK
1LJ+VnVOM3KlUYRrKOcEYyBGBWbZ1Rg3W506jpDUUYVAPeMEDx79ijmP6nWRzWnZ
LySP0YXKNfHsf26ZuYOkKx973G1X9f1o+f/7CHFze6nip5Ef/GNBmkF8nfnnY5Zi
K5lQ6jQBmnYvZYCyxiadAyBDhRutiCdyTxZ5pCtE+Dc0Q2whHYhA6la/fckjXtUw
f1p51TVZ3cc/WDMxBqrUVLt0d88LHsRCMmL6W6Ij5X+xU0AgBYnihjsN7J2qxLmE
OM2SY70PIqlq2MakFXvfrFo/H2o+Pxqui0tRIjaMYcDa5MKIAXVfwr6+sfEWHc5y
rgpH5snKQC8DnoTEllMP3Nh1BX3oFuTeBTTcJQXv2LSqFU/ZiYZRWu4eQLRIEM1E
tJTAh8uBZLt36allz+cPfxZloDbk09A3HmEzc/0tIgUK1XK6j+sAtrCJtAj0wmcb
EpqPYgteSRiLiH218eUTvZja/AmN6BjUZ9RVVUHoAqxx1FUJo/f89pumQIXOG3ti
uJZFaQi1P8ryOkvKbfB6rgRJjaUM/0RHGGz++lE0gsTIIko18e1COu1bRK99/Nic
FgUzyYpSjh/zvz/ZTbJ/NSHCCYimYbUmTZY/lkWRxMj4ZTfTclXS3dOQ4f7ABUeZ
7num4tkwAG1xcfS0KUrtppY/iCbxhjeWwaKS0VR86mE+6qI1QS/PWe5qzPpJ+VD6
OIsQp5godWtag9qjupJ2WdRoNua3rcHYTB+fnKVCr5U3pf8P4f+Mm8zbqpvBM0T0
b1jOuF9SoZ36/p5dfJO4LO/oTXxymv/ciD4RHZiBhYhKD5D83r/Ks62OhLKMkpgR
XHIrkYwrXajho6nnQVTMRGCm0LhSpfABkqmbOtX/IZEXhTt3IM33z93HcWZfxiwP
qaal38lFHP5qfXZLmLt401acAJP61rS2y6lOxnvgRxTtujdXrQyySS1Ah4cBwsap
cGJJPIDEP0tgY7vhTFI+zHrNJzOoDW+GhcXbFeHRT/64jMLCZ4ddmx7Yy0OAGqNq
6glgJcwDiO39658pC7GyWlaXYrPE6i4wCllWuB+57TbayZq30OZOTcjCtdvhiXUH
7yMMjBpz1d760MuYbwP5/nwReIy5v2ZmTeIMgNUdvJZQb1CW2p+gQOVs37PbuCf2
p7DciGEOmJ2ClkRjcwzoM8HwSwyKFaLdroGLB8TTpXtmv9B4g0w5u+Hdyq1YlNaf
gRoBW8rcXEErdoUAaO6EE8wd+QOnabozHuVJp5MjzXCIlW12zr0zwKmqdfpB2r2r
j4KKWKbxDMvQ/krCnB6vU6Z/xrzrcJ+EXCehrHVtbsl3AVi4Jsf2ewEeeqOq2Rdo
IWJKdyQ9T2i3Bu7/N5OQRIvBWVy0wBluVouOdPqp6KEzbNAp2IfdBkjIejnQAO9l
ijwwOTJ51Htx9ev0iuiPbS1j54wTFHOakDjzkOhvBQcVGxwrHWJunxj3sZwYWN4i
k7xm9uS2bgQeW0sQqST2V2QL8WyJ4dN3/B2b+m09rmICUMc4IQUELAjfSZWwv0f0
h6VZOjehzKdRLzO6qBTkfWfyqRrNjfrLRsPCzLUPRn2MHfQaaY98PnAxdNzlGVAQ
cER8SAZU8DoJIanc6cCOPLbH1unHEIB6De7tJ9nHycj5AB1p6y6K6oRPamau5CGN
Llg1QhqIVuoVqC2CnECshhLPchNHXKDwlPfKrHPzVKThb5NFwGLLhhGFSeGZuIDE
TVptDcCvq0f/MVe7ZhEYbY1vW2rmwgoZYHqBF5am5CSA+VYUldeEBrIgmXpi5nfR
ZCx6dTPP8Jk+xfeQ5o1Cu0FnhScuGiLKif+GeyEA44WcR2U4a21D8V2GSEP665A5
jgQE6maP+7/vWqZsMk53dgCdlTAZU7RhJScUvf6F4QFQDSv7IDHMOrDb4knSAdWu
UYke1CyJtDaiDpRy2tXTGNQgSifFGEV20EkZ8Ja+EQlHnwjoP7Kwl8FdhuJbKj2W
sxrXqhFHtn3B8ALhed26On+UnmMEq82Y+kE2vGOenfXfvrbdmIN3W9jU02YkLleS
9ZX7si5B2LAcGp7tYYOz6OvyVAOwUm2rNs/7vhRFxQtPfBsVfP3cmFVP5EuICozK
GSZM6zoadHnoFrzdtBBx3AookZ3K+ndQbK/fSwkRWPxu4Misv8DTbFawJeJ9Usjc
ST25YnGd28QGAVgvDMcool+BQOFRKK2LHXXVKjc+ZEYLROwmaNzs/g88MsGPh23W
ia1CsrUgDOsCAJLkZRSO0luO6MoWnKtNwzBvgqWol+lgZ+8HB9kXiYghKVq7Bpuo
ZMG8bcapxLwV5MGMUExVpRmk+ENTsV8T0LURpyQptfNOT1ouBqIohVPKc+LEwyjU
zOxN6vMwRS2wv68DIM5dtgDPeJcHeDgekHgNMxeWhxceAMUXbaw5hoqJkLzbIr6t
IL04eusVa1S+cmcc3yjvRVNY3Jz7uUC5WXbeG5qsydwzjaWXAjfhz/tG0D88Li/V
x+CGVMWBweB72hrG5NBWJeCEWyoqvFdTdbaBf7xvRtPWIx/gSJolzrBqGFlG7HHF
AejKVgWkMuaCWL+8ZkMQ6JHJGUAm6cAtuiK19J+GsI/NuDwqoh3pje1b+rBL475q
8UCRWEAkFb2L0jV4Ibv/7Elt/XsLznXV5oPgOOlACrmi6ImF/qcIFna3h+3qRn7u
r1VLuArWeNsPrjGSY3p/7VpMY47v64H5JYEfa/8v5apGFtVGE4xPhQVegzLO8OHU
9r8M793VMcfbWEPuV/ujwOwFs0yfXtGw5cDed7ZwRC+uYFJAsmghSApF/D2LFCKz
Y9UBEdx3w1XEvtpA5c1s8drHYxKu6CshInZN6G9r58pWxxDMSMCEu9a2pNvh4CR1
OdGRI7/uTAwtXsncnJTw63zy+f0/l2bzPNR2tFHuJD1+UTEfAGmQxDfejoCvL+gj
bQjd1AOolKggyXwEwUGPTpCc1XPuc5mwSTDhNOCmaNHoCrpGcjwCz4cNhlU/oIly
aBDBvnmVBLq6Adnno0js7piuINdNBXWnXgS9y1R/c1+Cqk1Fq/WRLkT9vvTBBEUH
ezy2gyYX7RepXxblhresO5kk2TjKr1biz+CkDUw3CYK8VI0C77sFYPOzOg3lkpna
Q4VSgFGiwM93hG0cQklu4R8/CEDOsFOJx2SvOjNKSTWngn0s7XwnHVjedu32dfx6
+fzNlykdCp+oXboJBuYSj9Ni2TmcN6GpYpP8via08/2q4YDKoybBI7vmn2GzHCEw
iDWIL/DpbsicuGKXd3NUOPDi21H5m5AHchYwj+izR1X8bVikES5SGgPgdbv501cV
RpdZFe7gYhsH/fV9cYaFObRxyV+Ui7Puj36kuDVj+o061rn3cKAT2rfp2b/CIYo1
cJyWhfblzOza8rZciIqAudgqIhShsh5Y4T/hvW62gDXZrdYH5XvoWtO2P3FkfhxS
z2yuEXABSvNl1VCOgs6USOaSNsi2XbRHaabIrxUrEPZTgWIr7ocEHd+s+wSQsBWT
I5uzXijdHJ4WqVJMLw3koEQNhHCClhPyq0iBaSCbOhoR/QeX06o8lhtpa+GM1RzW
K2nTWa8KCX1kzVmCQH4MDyDyHVp5f1VCUKJul4/S5uJqu2C4kSSeh1qAKeX7WSuh
O6o3QEX2v12hi2L/7UVJFYtqlp0Aa/BZq65SPKTNo66bQOYb8zYIET3zBbWtfzQc
rkzRFdXXSUKzqOByCM9YNUxl+Dlst8jtSfbTUlwBJujR/j5nar/IxnvNqXMKNG1K
IvJYnQaGBNUXFsmmw22VS5qH5UX8oRo4lq47qMGjq7UvLt+WKs9nUnuGTJs8aT1y
ePy/PJ4eJQMrGMYQegBlqre52aNrNTD2LpW9stj8tL0RDY2qDz9Dz/FAL/bBRUFK
ICfi3F95C75o1cLNeRqDng9IzCFWgnR/L/zCN5YYCh1jfdQHtnG5XUZXsa37BhTz
E+6FjxUrrFfMWmqII5vUII9kt7SZl14u+YgaC096S6gmaE5tyaHxDMeKMlwVowy2
SLIxWjNY+m1NeUuJ1CVR1EfuYC/+4tj3Et9da3fw7KNYgCuAKZ6LXFTWKW9IsviA
R34oomHEuea0wm41qhAoKWbGmeh1oTQGKF8gkStWrYjcyyteZ/OQML3+6hWjnhwP
rE2p857Bowjo1ffrIKjLFh2CXmDTIm3Pfknlsh5ta2m/z3nIMXIYYFe+bKgrwpcX
YxbkhjDZYY0hQGBpmqojtq1iTC/DkEeVvK2U0IZmIeoX2Lk+CR1OKnN5SKta2P2I
tcWcjHnRCOIBcvxWE9cASLHF8wLHDBJ/Iu3jI0akaVUfdw7Nh9vxd1a1Qe8EfZ18
BtIawTMdFb0+VABDx2yiHFglFxXy5RAxiSZY+9SiUr2FvrHiwFbRw40FVjww5q1R
QuffFZVwOOI1ga1d/ZDbDQtatyG3VXx+PwB5mn8jj/YJLbhOTNf5aaq0i291YYpG
JMORyAGdsl/+h4ajyeEwd+NIFdQVd5nEVz8Gm+1KT+2cYw2i+xUS3sTwwOhNyMBc
wlPp243Ij6JZoZgOeb1l3V+Pz5tvMFzJgcedODjGJGoGXsGyCcpsQjFoQM+AmrAZ
lpZHvnmX+E51nZvn2y/Mb35Hb8ugHACOyd26rylKRKxFZ3uP6gCVRFtq/LPKickB
qdp30Xh4pCAYeouryGVI33kpcQAv5soFeUHr/Tr4IkK+b1hZAXwY5sJGkOnYpbTV
+Yqnr/OdSPEMa4OhUsZeD5qzsxQwhn5HRNUtoX1gsYijilBceDiaByYRF4HA0AD2
/tJ1Ub3QLGIZLYn7BWgyzr0mQ9u44fI+eD1DcM+3D/2fOnGZGy76ENNT8d97Dipd
zLU43LwVzl/yvuCn6nc2Lo4MJ5rU9X9UxH7ZZVksqxS8QhYFu8ALzsL9+HUhk0Sr
2ursol72Ih+0LguEGwIsHKiL1d7ejHIBNJPPug96cPg/tTa5gRAtkMP4molv6O+p
rlRWp3vYXgqktNwlxPqLs+TWifpSHryNiBUURd139H8G37+UebachBl636e0sPb4
KKbmyJrNoofKKq4Za3UykvqY6LIL8vTJkbWK7hyYpG4NnhHyMIdIlsJrjEvyDjhN
Fe9vBVbn+5A28Mqx3mOr+OcpWMze1UtAZO37ELSjWdQIi6aLPz36goMfYiES0npH
eSCscRRfUiUsmXZrJ4+H+MQ+LQ/cko8ON/pZ7x0fAhGCPMhl/rdrXzdlss5XZqxD
8BK7KJi52AOIFuMEUaUk9q46tQPLAE/KUG05l51I4T+sfKUaxA7LLQHxcBbATUbG
eZbpnsaeityPUfgjL2EV65BdEV/ZAwt0JTlARQfX/7QxCdgnHPV6eMhppSv5Vkwf
Zx/gQ1Pi6lNCotd7nKKxmdK1v2kBNdd9Aw34REcFz6CJSD0qQe72RRvukaqX7Wig
Mo21wWpK95FtWv1w6bU9u6PHpF3ce1uoDi8+1aLv+9t1AuZ8he29uFGHfrWUL7rG
+H7rm2cqSapVHaDiVvFoRxvYjRRzpdeGl42FXJ2P2thKd5YfbdCoFQcqc9cheKe+
BOFjoKxliEMgAHZmjm0Nn043vNy5J3Jr7nKsA2HXEl/YpVyECjOP5GpLUTSt5yb8
kGAZnMrP14j8pydkbHM1opu3HH4nvjzfFjOCXdSYH+W/ubt+126qlgtZeBQ4uEqC
8NDH9O1/2Hg3vI1Tg+ZwOlCORUd9x0ULWox7OG9a6gkjk/EBUMwRXuU1pUqJVJCD
2Do4VipXZXmonV7kj7+U5WrCDy7ehTsW4VyUPWm5ZrjZ5W564fjosoAqJW+efwf0
HCM0hrFD+fjeuKxnWwqAsWFpJdJkf2Awwc/sNaeTW7LZv5VG+PPUFTumpGMMegAj
oVOjnfJcnfvpYRkVDyxgKVwEgKSWOmS0BXIuk+ZQmA49+zycBA0k1YDqy5C840eg
E1z5LHeclMcz16BCfctUNHDFNnUraSKTCEKvGEoZTRTmA+VI7BYVI5nNPkvyQYS0
C6YCrzDhoJKDqUSF4FJiHCHxi1Ghm7uuT7A20dSJ3V2W31E9QNETcnFHsvlvgqEY
SoyPtsYtKVAz6RaVavgbgvoULXnsKKjHhy6JZRRMCvsSRTa2qreWtIcpNribptxC
tud+2rd42mOt4WduxYwnh+vxStlSun/pk1BpBpBOPPvyo3d4TZ2r9me14t+qNwd2
RZx67RysEB52lMdVNcGVyUE73OmxAHTG10fku4qv9x6yLBUMqlzIIq0MKRo+bKop
D/aAdZw96rEp0hiwOMDf58QnAE1didenjeD9mBQZ/2YS+JBc6S73d9fv188SZNiF
ho1aIaEc+NOwJ5QDTyPhAAHTJr8oBThdWnaV6GI1u3EgEaY4tV1H5ElzRBYIaBZz
CO5Rra4m18HPQ275UumP42dgxdzPocmYX2xFRCL4qj9/m2HW3A87gpLEEVWSwFDF
wEvK7kcEVysNtOq7wXHoeGHIl+4swghHmDyvcvhYhr66XAAZW4XFz4AuMrGHOjxt
YXEiyaGX6sdnAY1GNyMA3NFNjHGWco/WjkXpoOZVe6T/83+kFvLx6iTq+vVnjfdr
6YQp8Oz8tmKfX6o7uXuY1YRQzsmWr/Mn7WanXvk3fF4mxp57hb4RA+T4VPPfon+R
R7fcQSR9vVE4M2d2AGcPfCSj6dGKsmA2c0c7UAe1JB2BIps9DkSUuZ+QTGLTC2vn
T0bHr9XD17UnR3lI6YiJ2ykGhWsuK+cBlX5HjGv3LsLexlPhtsyKyBG/WjMlJgc6
kGOYCgGPlSV/hEgcc5ACiTvryy1eAnnY9i85yUC4RNjxFfKeX3sz/dGKH4CmooU6
M4WTec3pxiY++B6bX0awRxVplAk7vmKfPagYJem+y2cIPZYDxqpIzXQfygvWDIb7
6fPjjJ83jBFWGFTy0e2LeZWB6qh0Jke0EAxcmX8hRsJWEss2UvD3tWhiqa49dsJ6
1ZErx8lFkMVxw3hUB7jz5WHlP/wxqOZnU2yBQD0BtgovWyVAJLFVeoWP/hBbM1GY
odjgxzJP+Q+jPKc5An34GtjNcpcb0uuSAfqe0GzK25C1OmJ45hV4n8Uqyr368tLw
N41iGFBts745yS7RPyKQHIVhV39D1mFFDEJuh5ELEjlp/bYWWd1OWdBZ5yqj4U7D
qlfU0c0+6geP+VL79/CHC+eJNtm3Rqi1oklGB3fmq8H17O6/pBfi3EtveGFgnQk8
vZCPpgtYEP9M4OnzQR2XIeXk59JTu3woqwGM8zPq3SL/OdjGvlAvEOurP3uuirV1
epxhM2COG5kjbiGdfe37UZkjF9am4fPx7NIT6GDrFezDp9mcZt9Fp12tBCPDjJYJ
9eq1K6m8MmFPVgCft3xgbX8STmbgRwjSLJN1JnBwPqVeaEyXvX5537ZfvbchayeJ
XURAKbrtn7BxY+HAnpqFePiZh3aw7Ye4/0sRK/0dUwZ+XMT/IqqJkPPdvqj/0EAw
HmpreVK6RaT5uaNAP/tWZLc5AZEDpi3BiXEKU4Gaux9unFkpCfJQPS1yXKgNnRLU
QIo4AzhXiZBX8ai8QnYvNKnmiORh/v0NUmZzv6HNXJcM/38DHHvZO3HA67teCoC7
9GDfMdalDk+ldqRQhE3cOfJd3L+Yu9pEEzGxl7UU1eWZAXDDQiT9qAdk3GWmx+xV
BeOKzPLeyrrslyVSHUMVO/6SIa/6ufP6DeHS0/h0wPsXXjRBoc5V56v3XblU6GqK
MopuzmmKiXoVxv/WAdxFRChIoo5Rya8V31Xj8rM5AJYVaLOZgY2OKNqiopJyCUr8
nIAXs1W2hCn17mmVdG/2R7fFm4d1r138lwPIh310EyyNtPVTqPMpqLXJVyOxFaAd
vXeNtADEW+pl34YyYDIAL3XtDjk7odW6aUaueXGg00PUXRSovboxxu92P6Xr3SqR
V2cSSPa4rXV4KiSFD42pRaBUz75UDmw/EfkZyvuOMwzG9eaWd2okiWtNbBne+sxn
N2oBpy6asMdCDS3i5ic9L1Ay0R7XFFx4rMgFtZJS2r9rvMaSz+08uEeCZ5+ch6fD
M2gfMpleozmEVvOYWyHBFZjAeSNlo/i94csj8CSoFTmRUzKqKaiZvtUJriamEL47
8IgvQIJMaMleS8YtSP43fsqjiFcMgrxL6Qs6W+khnU/q5EswiUGAThbB0V1OWGxc
Z0WoI0iBLHVGGQ9X4Kl7WlBVtJ6RFBVb3vXb1A1oMNpeLTA3vOKXoLzOZ1QqmxoF
Tk+m9tx4P2Q8Q17unVdBQkydyQA87gIBQ3AmeREOk7WsKPcICdivmR9n5U5IufHo
czpgrjclYbzgg0jnNdyem76tC6XoUhe3OPe5RrcsXlpXovOEvIAA/JBS4ey439pb
6oGzgpjGFEbYulG39kwqq3q+bbLL9sNZGu/BXIrf+YeLMswulPsdQWPyj2nIovwM
8aDO4CYq4B0V4HdvGK4DPFOq5bDPAwN6rUUgkK5QXfN/ahHRrrfOwleeoHnwmpG1
AcE46Uk6u9IIYLrUeapQ5Q2+P/h1pApT4A+8USrNrX9TOjOFvFH9GMSTQzPSXMAT
rGvGc9q0TMak9ugV2A7gyVahcDCNX0QbUss5jMnuWfug+51n1DSV0jbTV4WuDuUt
N4JngcPsY7x/j7TbOiF4zLx/lREKe3tjudqzaBTwlD2hpTaD3QWcbtHrgNr7GZQR
FWzrk2QmHBjOokj2Ml+fbwTc93t94eC0kP9/AQyFEuRJNwWgA/Wsbwyn6YG1rnfn
420KFg292waos9fYhc5etGOaaDHFNDwlusc1by76Gu7xpCnfH5c95wwhSFCY71Ml
/xmBvB6DuLw0pqeixNx56VMTSekdr4A4j/pn4Dd/5HfN6ijAJH4YkVpMfTP/boIi
hdcYQLW9jmXbKv5A14Y1e0cp7Kf7+BWiKtNbBbXKdto41hdv8TvIVcozd+g1X5/M
lwLUViIEppSX4tciL9DHmP9AK3sJD80DtKIwI0uvEstKu8UDq6lOC5nkghIoKhvL
fVjqGXyxcdBuDO7DfFnGlDYSU6CjAnpQFxNDTvG5h7gzvLLkhTxboswMfjkYHZu2
h1oOF923URGYgqY1ojPX6iB5toE5+FfdDB0BK7EGPD5IJALuDzgaqSPoimBy+MQw
wB0DFFgd2vdUJAIMclwBbMdwAs1zfWFPfK8nQCYUazCBgq8lnX7y6Rn5E7iHRGUK
U9TUCQL/gTeRjHy2gOgtW5xQcap9owtWpSTzJ3En8SJDDQPF8SAPjct0uCJNkczN
crBzUuvO6FD26gLFY9CTPcM+2Au9bmgeD1Fil+Q49k7OZ7L8fa+xb4YtTb5BckAG
EGYd+XciikXoI22ei53+bOO7RW7+PMfXtpT5AovWXjsOtXEVdHYMd8o9Sm2sg7SC
tODsPCF7Capj1soFObpzP/li+qskB+y/GUq8Oxz06UjkCkm9f8CZP7hY2tIyPb3Z
yHWmDgMXGZjjbkTGIyPadSSedGt7oCTQLoG2uwJMRtIlaiXV8mXIoNBc2Ny8XE6H
cmXzGzyvSGZft6p/bR3wPdo1sW2l+IpBSjR6ZIExEG1dF+Zx+2HWyhQqwRrOirhk
fn3nXlQbr3PBTwg9pJUrIguprI7B/e/6yvvZhq6tnB1RHHVamRZFgqu908Rd05AQ
HJJ7Fq1onTWW48YyZJNYBuUBnhAL6Zwcwm9SSehcuCsn9CbNAuda5mTzhEywO03N
rkpTy0Q83mwaSPtK9aokLlFEhAIB0muBBGlu8fvNGCdDgI6Wq3QpxKUBh/Cvv6Jx
u31AOxjsgs47CPI0HPGg48tMIasNznISkyBkKHUBRVPTmYxu6yHrWGwB34JkyvOz
vMjZXVP1OQgYyWTjHJx5hYBMp9PfkMLSGzqYJoDrNzoFIDq0wMhHd7AACe86VsUs
izuF6U+B0EgOY7zCCpm4R2mgKBg6Z8y70hZhnYKoMaNp71bD8yeQYCvIlcnw/JEr
NsTAuEuexSyZcA+oVnz2Ovttrpq3IOCTSR9tO5R2gu+6LiTyU4BLqnH0mZRJzDtq
ssNVh/rVyrR+1VOKi6pfkQzAaZDJa2m1D0OBQ7z8c3lWBfSt5V4H/JcpmwFtLyqQ
TroPzi4lvCvpTY5rNrQkc6KWwCu//XCFKZfLlh/ETfJ9PN9JkaKWZvRE4xCmO54M
CZl15wKoxfn8/2RfM3oci+yvlxD40TU4mK5WV9fvL6ajNd1sjsBoG8lYdGq8ktT0
pBnNK7O5poW7/eTKaXCb6NwagF1fYsX4qwzLdNKeT5X78j5i4pylgBL1AoL2tJxw
Z6TTkvQwDvPFmymQ4fTcOhXfHIy+2rTbP5C4t1Wk3Lssu/fBNT/M5pw0W7vUTR5z
vOkunpXmo71Zty0ZraHoiMAEg9W3hE1BmaheZ11AO6ZUkECPyi3T8IIw2l+V9xdj
YNH5KbTh9Hu1IqzrnIImkY2VpCQUnQp+nkZMa8MBoZ7j2SbngRBveSY3KSvxXGoZ
HwacrQN13uw4/DyERl0Top+8m9IHZ/oHIgQaK2XMeOEnrLePCbNz03QuW+kLcNmo
tFhG7q9JuayaD2KmMjqBu4h8b46F7E1qH18Ab/LB40AgP4thzDKfjPss46MGeabP
zm2jUYf3mafYC6t5GVwQ+6s8exA9ZL3CNeqDO4Zmj/O+6Z8BkbAecZDG8mJZRnIA
2ZIp5VPUR3UVvX2GenJ1O74JOEISPEulEP6HK8TMZij/oWnzk27OUngkVLkt/82M
zy7/zNSEGPa15eOrfI6fOybQTr+jF21rm6XhmfTCqjWh611IotiE1sb8mVwDc8WL
/8E7CoVudc+ELboTP5k2XDotXOUNkYWJMdn/gD0z2BHoFQgbN2CZd2alusVRHdBb
mtjuoLT3l/mYTzXYIUTa8TTdemQITUztJjJGgacJn+ah9y9oMb1to1Iz5zvt6RVQ
S/77NgGIjZr+0ziOT3zi3ow3X70K0e6gswedO+dOTNQCqkR1mPT0LUXbBl+XpBlN
hATm43LEIzORviPq1moBs/KCt0V7DHBNIMju/RzhhMHzDdSB3dt849K/dRgC5sHB
wnJ57b3PpfJ6fRlM5a98JwB18Tv548R92aSP+VF9z3xdv4drUkb5F4MqtzQpZYTI
Y0VV5ynAlXA9Ff3atIwQF1qlDsWXYLw/foaL5nsSTqOU6TA84OIojgJnMLX/Ybfb
Uv1cd4q+Tufya7003h1jz1Mg3irI4g7Y9QffmMuP+WL0ZvOd2ltXVn9mBEFfBNbh
ucS1iBVtaN+tSDfX1xkXOCqgMB1WP4+nqTn7RkzktMJK9CEjVIIeYH7Yov8dmeP+
8Vo36yaWvb7LjGvJiD/lgXD+7OBhGfjlaynXWOdtfmhZbBHFT7jKKyGZQMIU4gy9
TuuTYWSNu0PIJF0Qa3iFR2PY/MBIBajSsDWE0+1G7/HqXNfSgXlBPoaAS5NuaYwr
7+6x/c3poVee7BFeC+s5WPuNIcjlBNmWjXomZd9+eKMrNtTAMPPFsiHPEUq+yE5z
0bkFyskvTKN+0nhaI7eB5rHK9o96VZFcURnQjqOYhjxwni+QBwscudjU7lzmdVyJ
DSfUGqabchq45DGL7wlvLS12VBliM8ONQt9QOxi8u5DKQ5nEb9ULcVnRGc8kn65x
WUUO6+6zTDeDsqEoOnj0HesuDJ0Qr/tU6XoKc9wuZIYjt2M74Cv8KkLiAru15muJ
en2w4mWIBJ2zNwYifhjOnLVT5ia2BX8kfXzkYfY9O7nSNQX2XZmPeEUYXpEL04Cg
IjU8eA4lJfrSGmMXI17/BuD0nQtbu/J07GUup9H9sBXzsxUR+Guqf7R/BQqVjmlG
yebgHZm0AzgG/n/UyT9SmB5mgsrC1Yvwmaf+w1E3m1bwQt/lS95uF+B1qzJNWQmL
7E1OpDmccrxrjFpZUh0MrscpK8SiIzfRbAAU3SzDOFqeGZcic1WNGf33He4vwjPF
R/rY1VFPz41eePwun6E7hn0yjZWdXcdh+w4BTKKZWYwcA0x/tdnLKxX9IQhnIhxc
YYvDaQ4RJU55XE4lArGiUpunSxp2sfQQENhLsjlzG5XN08QG2wLksvQ+nMkuWs12
HYQsjeY39y2CbIzaoGldXI8msD1iceJSsUjmZTyLMCtdl+PdDCCeXa9dFsi3HoRD
WbQHhn99J3oWg7OE9RVLer10dfq0NI8MtMFI9gESM5p9VNTpsVaIo/1rnU5EYw0S
xKDCzcne46iPt2w+2v0ygENQfoTrH8WBgEi1igYu+8FIpKtbd4NqKdFgAX/dSoxR
3xtbnk5LZts5IUbnBSLeaSVg+FdOtNz4Zaz/fbqWYFJDnOjYvARoyA5YCJv2v864
wQDJs5Ir5SnfT0+BW1mL35JI2dRi9vbq5ajVARZsEXzb+kgF50n3Kd7St4lZMhhn
o0gSp+PewygFH5FxCvzUDT47Py2GiG88BBqNMDKBpgtwJExOnXrJssAjStGf3CeX
LF9L3u5//IoWZCYiCDnuKwChjZeq/0KGtE9yqpqtROl/IBXSnhSTB2wapDupjBgC
A2KNoIytUbfzeenth8C3NksllTBC8RUBQCy15S23k/xEGw72JMwxtj9CYneXHVtV
PM2b28U5UgzOWu9V7s5jc0qILIRrttawj0VrZ/ORsTNZiQpWpmp/0E9YXBLv9ty/
fZ18vFnfR0l4fwjoLFkp3YJt5tBQLRHgu6PBza6jv+7rop8vuI5uazSEgUajrQr+
womzbuDN/aLvNadmO5rl7+6cG4P9z6PpnRnwsHntFc8t7LbgC1N0RCtRftONKOPD
f9Xo0xF4V9Q8VfMuZM6rFbdv/bJmYxFy46bSrJ7mMzCvEy4YBxE11ifO9X0cIFOZ
mJcGqq8D8xLXdHt+4UYFHOZfqBXelasK06RTF7hQdL9AW6r/vakk+QIuVQWYVbJ5
+lNAc+3iXPBA7TV28UkKRBQWpdOVi66w1KEK7+2KXjQ3vEcVbjwmoZ5K7C7pSCN6
9fe/WQQ/wBz6Rx3mHQSZr93DcA+AGWEgTagmMclG7At8kLPxHhpX7kagUfKRP7Tj
KPpQJ40Yk+fGycj+TUQD3kNN2pMx5rH17nrETSfkz4QEUrmMe2/h+BnSfkb/hSR/
DR2aBMT0kAgydWFejkBd5unBbL9T7CdVdOK7Ze/CUqkRBDtUDuKcYvAdzknsIosf
QLtrtHou1qSOfrLEaqWswEqCMJXUnGAsLoSbTQvcU9lEw6QjAowt2LeH0rTFekNW
eM91qmbPCAdzku+Vh0Id+c8cIhAKWTvhDBETHKS8DMHFS2OfQHoLoX7lwratFvWh
GovRn95xHjGwJqjQ32hvvKsHgyXtYNaSHXWEJ86pOSweVvQboLPOm3i8LOcZfQAX
H/KQEAp5S3LfVMo+xdSkscDyYT8GC7PSI/B/BhY1xUKBlUi3mn43417gL+wRO7LF
w6EMXWd80IAVhioJgqYspmqxFCu3PPEIB1rGa78u9sX9NQv6whpcb3WNk8sBgdpU
Jkrwy5REZxs8n3O+xT7gQ6CiHPO/wzK8sM090uSsz4bFRSJ9urSjNzR2wiGbfPaA
v3JbkVcyoF38FUrn0GtR0vnx3yKkh/2SEOSQJAbhzcHiLYg9j753zyEoFsZnJ+zn
IgdUkKdKFeKzl8JMnmX4LwBvWjyrcb/DRfzv1n90jKSxvneWso6VV7QUb0s/FhrX
cGTS7wDwOBmnUOtJMNW+HECsA8yBrlrBN/smPV2wZQdFLdGqWwDVE3RWXkIe0A1n
8HVvMvlATuBn1U3kpnYZoDagtxJPBhECB19jSQtPPhf7f2pR4tVJGZ3NN1UAU5B1
Uqdm2QFkX6ma8QiVqOuBjqvDQionseqSRqv7yEfmLk43jdh9lizP8na47+edDyTp
X1UAe4u3+IEGyTXbiv6g7FcFJB+hpGZJi7kbVf7Pbiv3LUVriU9chbYuqRjOXCFd
kO/lpAvcF3mw5W6v614Ie3AHIdlYMogULvXiiwGvb+ELerli8gFz/m8IPPAyO9oh
AWpkw/40z29Wz9cuPVDVMY9CAakwBpVLxZElHZ2C4sdt92CzhQCQj7hLZlpWlfei
k1vUz40WcQPmBx9jmfXs0YJWHjzISKMp7Gu6Yn3ud00HD8Of+fGDuZ6kfy0NeXHp
yAmsaiHKTG7FeuD3svwzRE8hquX/FW9yL4OtgSWuCgvnjxfr+ZO+/UI4KRRcUyKB
6Ga+Knf+virWsZilT1ESnwFIBHSe5WqIw6LnkXayWcC6yuN9IY2MOHrKKFFygdGX
Wn1JYDMtOsKhlZOUU00zjQH3v081X1r1UXsFAFQHSnHWAt8uYWsSiaZ877hxnI+t
k62TT5atwnaraROKw+2GjikJFlve29cnh5nFzq4AkcF8FcA0ITaq8akQNEPGbsc/
8cbSyst2rN7IfN6shJg5miDUFeKiotyxuSWw3nEfgJXNyD9KSo87ilg85LLXV7rx
weS7b1lQQfqEZFTref67L6iQJ5CO4tjIHsfJWnQG4T4uiwShSkS0B9c+WUs4kTny
CeYMaYeUajjZNM72ZKEz9CVFqXrmL3l3QzXbBnwl4uNwPYnVH911OPRvEvqje99i
Fl6NEk/D6Z+E9hSA9IKTMCx+o72+/k7btz/kO+k4zR3DBR/kS1GTVBx+Xpye6aEA
zQQTfL0Y2+BIU0Cda+ARlBTzGwD7KTbrEr6K8cXypdfP0/ulmU+6PtnRL8v0Xt4n
lYYqGzEJ0h+twlfFC696JJzkVGcgysdvm3vg50bE0ZVzdGxWMn7LY5LiZoNoW6hz
O06QQvUB5XySP0p8PZAcXW/TbLcQMuXkXG/F18lt3cQ+jf2Uz3Ggmg9Ih2w/lu+f
LNtsfq+7qJkpafMHym0XyCSxmmjmbGWfrHGCGg6AJO2qQRkySt1NfZaO0s5vu9gX
4JCzZCJeJSPeBJYP5U9rY1GszgL/Sl/nXK5m+pv8+nv3MHuK3ssk9kN7cFe9FhpZ
nR/ENsSaOyGGkRoEZ7wQTYetkatB+VON5ImMdR20mt5inUqsU7Xilw9vhmvcsXW9
ih9Oz3WeJBjSeAfbNQHsf/EoYP2b3GmGXUb0Qlryq6eZ30dOANtLMl7lFmXTADlU
liUDOzjnc+8+re4vzbfEgz0+NkDdGBBo3tPWjoCykCbyiGN6epJOVda5HL3b0keK
G2uZb72uizzc/qnQocpg9Ju2klvkFJeDeb4JjgPJ70wZuhAbbc369D3Oob4M93Ej
hAUArGuzh1/oAYfyZJX0wZpK5imnN7URdROCrUpkJsz5dpZ0dpAQmfWCvlPiEDFp
meG73d1IyfqgYajAL5vdoHRQelp0voCmWwtKib7X+alxHL8qbN2DqMazaG6aOTrC
+g+SXBzQFreMl2tJf8jVTgqQwcsi8ZUVHS5cdHRzfSGvUZ88y7X/WwSXVLSsvIQ+
RL3B4W3aEI6cBsZ2hz3I6MEh2/wyipiw3bJOsvUlBXbEDtKJcCB+kQ4S24eKyftW
RNZ/+J3nQsJOBWLFiyVORafqRIe1PqFRIxUrPwYK19aayppcXwCk1g9Zxm7Hb8nv
ofbFFYkrF2FeqngiJFYjaVaKHe1sRp1N0t144QVyXJMelJWqWKu6lIUzL2X/T+I8
B1qqR0oLZVZb2pdHME2kmATUGG5mYnIJfZcfLLnNBYnbhTvxOHRPxQWWTmwwG6nw
L70QrVQT60uFFElrBLQHCoCQiuR0ScPc8WxrWxNUP5SHfqDv82ppLMC8BQSFH2tH
NTVsh6FAdxFP2/PDCiMs6k++rKJChQhO4gjfjs1k3xxbW2TSRFv50QYrHMCEhozb
+Lu/YIWIQ4Gd+BTz3ksvI2ia0HpfDl38nDfr5D8yYM8JcjfcvoeIzktVhYce7VRP
6i94Q2CJrFwn6zRafKtZQ4RWqsZGJogkOqd6igK/expli/OmN4S3pgrg3m8lEkSW
p4d8LL1l2xCPqr4F6MIln1o/PR0AZ54iuHDtE2K9jq9MtNUqhBjuPapjeCqfOwmv
AzwsOjLySS56RucFc0fgD3Jt5faEDBmyz2zDPOQHVWkzJhfH71hF+ftcJJHbcRN4
R77AkHB/0qTntgBVN5rJMEosNVOoFYGkSe2hTfDsHPNLXGoLKp/yWKqngLxWv9z5
P4YLkZ7bEEIruNhEOFwJIfriwrvnVwcu7EkAdjcjtM2So3CWYfMkOx4R3vj9fxbx
BCLCfM2N24MV0K7SZkRYXIcmF6IfTcPKXDXa90W1EVYmUJq5ifNRyGRunnwzN678
4dIhObf+qqGD+vVpCgJGINp+SivvSrvIra4HO38Y8hx1m+9B2hPb3BAXnBARMvIS
hZNvXoIklk2d03GOlUTeb+rpO5UFH/0rVnZ+77TIqRADi3t0wsL+oVcY43K/6I/X
j4sYYTBOnXJ0Kz+mQXD1eM51nRpO1aL2yRzMfCaj1qiPvsyHWlo/H65s2wQhwFmw
rzOODsDTIHK0wMAAR30qVIZ/mx1nezitbozXjyZvZds/2arlj1IacobWMcnGnnUC
gYlsaoG2TLf+EAicLl3qly6ULOcb8ErrTuh2TVhvCiQTI/LsGMkOSEhcfqfjBRKz
PbTjuSjRjjjGYnNfI8zuos2ZGqSqjFbtfBdU6m44ovoZxZGQGDyiKD5fHR7dCfSm
1g+y6c93dGpq+D4CNSWdRmToA4m+LEH1ForaAXzCcwPfGEc6xXbz8fwNYV8nFZHe
54sNtdeUXqYXvCGME3mEOmLrdZ0ONsxpypKD24xbofI0Ug/zsFaA6yK5MHyhmamd
6BXvN+Sb22t1/GlYS9qhJkVwi4y1KACYfBpNMMX2gmS7IP9tqvZQSQKK/pnqw8Dc
UWbKHLKNhMiK6bPsBNAjL0dHT6UD7xTGaiT+JwKTJVkI6R9IaO3m0boVrAKFeekE
in3aWiW/Enhoszu0difb7QGHdO3BAVj0fudHmUL4Iks2H0V/z4t67ElI+n9FxzDI
2V5FeCo3P+a1u2XTaB3OMOhBY8WlG8MUAsy3kj4VrPw2xJAsRBHqCbEGOyT9nRH0
lr3/qqDDpyZceFUcGEWB4JF9LgG3835J/QmkZ0bKln0XE3c4T7oKNtAz1l5E5N5G
A6KO25tc/o5is6UQeSWRpWVVEFzKHHT/omST7x1Taen3arl/I5v1JtZ/G4ANrYFR
M74tLvtYBOek9KelP8SCVlu2ap5lzgc2pATR69jbYyDl2ZQLC9sJzJrmAkdeIMiX
9eNBntKvtl/6GoSnMDR88yJYlzSj6LPMmwYxFelNghMnnUxxlCzxS28WgREaHgjs
pcE/qetIGn7INmrnLzkvhETo7pGkZM2SClbiwUB4JZhmeikZF6e6MQG8E29aWOZV
aSZW3qG5ZNlQ3AN1tF18zhasUZaN3g6b1utKgP7bGNK79U/kp22wcgsHZjtn8I6e
hPjZZgg2ITwMhzc09OfbYNDNoWM28U9803dLJFRRonieudkhOKEAzNvyPJe2y5A0
3O1pEWIxZcCnw5EbK/3hLwo94PcZFgeBRXGjZTW9swxrXkxXHOBntxKdGfkxUqId
hm45Fpco1t6ZaGkT5o5Zgef4Pg5bDK0ms774xPJ5J5zWqfBWvBNkq6thaMjfo7AZ
aNP4hGowsbJaAYfqr8K1Z3maPHlwf8Tt3QIKD6lDAQMBAb6zElwUJZ6iRE0WSjJo
ljacYVOOuHvI3pW2LAJE3d82tFjjDmf0PkIOW/2m8hhPZ2MmbGnUzMot1Qal1zDP
G04IRHEjh90pYkBWW5yWSJ6m69r9wYQuD1Ow9izpmpUJamC2ScBsWEWbEm76R0Yq
qhIqj1GXu5KIpqQZAiqEFUvWq4VNKil7oWRxAVj0n44JcVK8kZ37LdTLW/wqSb62
JpVy/+ohPuLxWBdOIwqge0EBQKsNmWOs+ensvHAFuLSeMTJnR7r1usa2Ecj26cCi
PETVX9jOUEfrLO0HycsYL50tvp+esrq5IO6DCRQQweweZ/pqSmkt58TLMnzvudV9
N+R/dmtQHWnxNHR9ZS271IIrcLnUjzjTiUbn+sxEAUQO6H/1mg2/V9nYKG5ZlooF
omouYBtyF8xB7xX88f8Hw+z6f7IhwjGrvEKr2V3tkaQR3yZ025BUH6Mvb1uPz3PT
JXycGihPg3PSD8ftwZJ8YDy+vPbSRj4o5adEQTLtT/UVbJ2iE8IbhXxB4WKQsarU
o28UFGlAeEchFcV3hb/L/Sp565zIHpwS3seVTJhVUyIYQK0ICQeNfos/kPyFVsbw
NgZQudzxe0aNR98JeCOQHmId3JTOKd1BDJcchy94sjrm/jSSguFt5od3Y3VkkuO7
az8DtOCvmKZuwsxgmClq/hyEGXnGMcqU7MrZriHZVHRMNHq2QQZvNxa9cCEpAyXc
Sf0gb/H+yVDWcLfAkOSBbR2ZP7MRejlZJgacSRAgcCaHEavm4PPu/ObDFQRwaPqS
LwQSvjMa+dy0Bb6CJQ+7Cev1Hmf7OiB1YFgB559IZ+JdxlKj6Md0VOL9Qo1gK64b
sLOB+fWouam9FY5hzWRgtC8iFbxOoxYJQpAxsLULkk0ZLjbMD162G+dTK4QxNGTj
Dgr0GDdymhtygkS7VTLeuAFXNpcfbBmcLx1RujGV2Vu+QNFUMQ+ewLV/ZxP1xLSk
MI77G+V5hmf2D5PT9uJCZGE2E/OcXfHQEVZzGQ0bGhLcSC1N3CsR8V5Z0/v3Kc7/
U0zYnBojfzUHiNI2NgS9XMpvKWPTCrqPr45nT0I7TEuTVWdUIH+yDjcxyEiDij7g
3lLJONXvLg+XohIOODd3Ccy3U32gSstm/KjvnlFb788bdnV/LMGEOtuL+niOSMe8
xOJ7601cborto+0OkZO/uQI/X+u8sFPk8aRp1AgSgiTrYrhm0FrDhG8H34bKzq0b
2oshMe4BXZEsZMqc9K3T1QrPN3O4s4/oh65OYjERaZLSwvcIRu+cuRr8mIcDH+sO
Oos20z7GgT0k+HWZOVO/2nYIXlzzhScnlGXDAJtseTkX1DFWdoG75BTqdbRXi2+a
YxOxt1nZEVPTtncpwHIWAXpnFQwoyqauyIh49YGZhqOSQRif91xKvTWpXpoX+CBN
Q4PKReoMl8p8liYtxYBqPFKO3O78DWsvUMCBB1AzB7vTVSBb63JWp4EOTSrzFiVY
+IpW0DJE4nD8mAZghxdbt5eZB2uC4v2YmX47ZqeWKjIepeZggaqA2rIhDzAktPec
IUgJZ5wPYM4bICbVh+5HzjHA/FPyC2zOPLvBLXFtN1+4+Uxcxv9z9qpPz8hsoLgF
NcwCsYaFwbGT564zO7BMK7gbD+9DvxZj6VTCxakjJXtF1nosCSwXbwCyh2+yY8Xc
/apHzhB+J14uqkatYK/VVuYVAZcDkxhEUeJbpY35cf+JyMDuwLcOmpRHZiQiezjI
YnRjbxafL3hFKxxc93ilGOcaFiDNuWDe0yrDdMH0rmgzVpHw6QNtK2No248PrhXV
QWdOeBaNcFaJLayruDVxMYLU4Ifsl4cACbU/n+0gNLT34G9IC7yrOc8TFTBxCmX1
JzCB/AcGi//k9kL1wESllybkEMXFnL+5lOmgBQpCDtwUlVdFq6ysEWZmSOejtzcm
lO1MJiv6jPKvnmrx2aZqAmusTfZTGH51glq/HuVNEbgxy7YPu6H8O18rxwFuAUZY
BOTN+W4ZYjbFLxtEMQX3kPX/9YFbgHrs734w4+wMVUa0u5YfSPwJ9Qa1fZBUTGiR
4VHL5vBxafhfv0LhH1xMUi8crO0cLNVlxtneRwRrpiy3y/SE8VqiPqspxjuXAqCS
dsWMRMKl9kHO+VliS9frH7C9FkfQ8xKxDVmZccMwjjLvNQTVYmf4HA9r9fIqsdlI
dHOCxfXL6m+e/MSe276KCLBlE5lFGijm/y4cquA9GN0UMzEHSpd9O3Na7jGYfT3c
YFQByH+qM7Oacx754ZFtDOi4rBXMLnABVURtuvbWPT5dvyMTccut5VULxuMfZ385
T7CDAxkUUgH4EvHHyDR1sDP0akSPfjNVWQ1cU+ts7CpFvBYiNg9O/uNfp4n6McHh
Vqawem+1gN1wOIDVBzx50E2sp+bj0cZCH7GEsFP4mCZu2oaDEQne2XBEMjx4ajW1
jrpOFU5XhTOMjvr7vK8maUkvp6YU/kfDKbLNHo9cmZrS9asHkHWPdaw446AznsH4
0IUZiut4+uUMOh0Dv2EqEEmcQgQodaoAegyR0E7OoEqeUfz2qoIhbEmcE+1OnTu6
Zat4tCFBMnKW2xRHSW2mM1edk9ENvBYnMsQQnosstx8fTpCPI1rtPfPJSZIB6L6d
1gyjiQUVsGAZf1HvpZvWwZ93kL+LtR2u4MsG2sP6uJ4DiUUAlXrTQ8tySKzJ8DO9
6dnDXDIrd5Kqr+Rl3q4G6eY18UkTsNlzF63a/FZtUk/7nfNXBRLclhNcFClEpWAc
/41QCT6+Q3TT1JKTeEMOXs0W+Ehi/hPzDetvfBADGI+aMz9jWV/gydcLntYUC0Ax
NkCGMy1/AYRm2zJu1OCjVC+8myhvpQiwVARnA5TcqMYe9j6l4zglEHwZLgmSazt5
G84eMF4rvGHELJnudnKe/AfwkHkz/9zkfiufBzGIxh7H1iVvMlEVAdVbz8TAY74H
nIWz15GBkRAFvMs7HvbyGdvmUthuKsOUav4woDW9E6eOWE8sLeq/dra1emNxH07m
XkcrPBbccJC721ih6zTsxhLCxWi6tHxMdUN5oWh2oSnJh4blE1bUKmBIzn2yMlr3
s8k8WzKiyjlq3tVpKJ5xAIT9veGkFAA+adOul6RhuoXI04K+PySmZrogncSKJBPl
5fBKPafi0ZANNcNGjzQugMdcShsWzPIq9gPN9sLlvQr3/iikZFEs3awSJif7LVKm
i/eRw5w+6pT+3ovAT1icT4dUo+byMSPhEaTueJmVjPrPEfPQoQZq//XbcGPBErvZ
TYlihJfvx9phhUWCVxgYKpceAlOu2MkFKdV7NIXyGhGpMFsBlMYVf+AGVbHjkGcc
6ObWeiVT8U8YJObOv3HWGaf2hAFYj6ov7p/uvDvp0VwfCja84d4YlpPDAGqFxcjM
9MyisCbTjrXvyYIDKNNBN86IcuaC7DX6+nx4qk5YeABNhUegzrjihNfw836B/fa2
42YJcizPzChRueperOFDR6suphGK7zNvX3GBFO+y36+ZzXjBPCPo6U5PmVROFEGH
yCjI3+p3+bq/sqYEyVdTesW9QkFUBRdz4AP840TOp5nlR1hA1Q9/jb7C+ssXbKe6
LY46YAru/8nv9gc8vKuoHJehEE2bD7tXK0iKOGh6CeDk/1/RRO0sDJv+rBEqfLuH
2POn094+lDfSEI+RujL2iCICtojhq3VaQNPGFirrXo8T5HIXpR1+STsf4zoUnkZZ
WzXqplJkeSURtBrvh+NukyxN8sSCT9k6SCF2Jyy8/pJ7MNKJpOre8iGCXZBTmCZw
VIUga/hdPrmLoFcYSXN+2x/buOCF3hUgm6mJagY2Pm+qsv2t3nY4ML2DMFZFtzmb
S2Yjkg8ksaLiZCMo2m2EWZmBjvYxStSfsVGSKEbJvN+o8RShilDpRSHpQEZkeLXC
KCEsr4vwQukRwqH3c/NcL+810FdumDoO/7FK7gmwaoFy76kE3nP3kjy8fgvrivpH
JuoQ139/5hBmAnJpimCa/lNc/3cgZMabbC6SjLPNyY6/r8HjFfE96AJyuPgarszC
xrVwxyB7/Fbhz95txjk07TZM3O51s6u8sif+W+z7gSut69Hgj7BqwR27NW8iXoE1
vCCHuGVPTg7goMWcF1MRPztxpi6NhLvYP0FZ6fabXAri3ezDVCLx9p0h99hczEpp
D/wxpBphdqWeGe9l61FXPIkmtGxZmuZPkzYx1jbVLoG9+NGG3yMW+fQVOOqNVoKi
UtVr1/4D3SrPxgl2BPtVDmFUFqHJlDnmhVLKipj/y9nwPsPDnzAt51GQbv9Hsjm4
mEQW20Gdz2+HJFaR8T7sjVWAtlAHYgB9RtB2TTvDhiNdFkxv+3k8kvAA3SeIaqvi
Piv8L/vtWUINu+UsIgzUv+hgcGPEd3IEjLgrpAAV1BieN2/2MQxYKfoehh6VjoDm
nTrSYpIqkLegypZE1hW2UTgM0L0mrnRpH9q7flUuSv2d9ane4ih5pPsgL1ulmuET
6jlFE9bq/td6yeEYGptQtrcLlDmGMWyu2YnKkKYN2ICsfmL27amCCXJCrk11mpkI
NerO/Zp7ZsfZyEKUceOAWd3ItzOURvfnYRm8srIcYkU1tBJ6ynBIWlUJ8XA6icoK
eY4nTasYuHT4U1i403gf734SqbI4qW0Nd+nSRSelOl8140HBECQd468UIwbzKmTF
DR3ImQV0ZcRx2tueSpXLRI8onO9AwObH/OHSk2RuDubnvYhs+2zV7WvoWMBV0UbA
YFM0mtf+8zbio3XYlteEunikaJOh5+0nwYkLycvuaYXfGSP05Ctp79pUrbvwzbqZ
1R5JI5j5GuIjayH3op5h9XhpqBigQuL1Q5tly3vYlYB/5IOvvcy6pZCqaJymOaZL
qHK3qj2aLsDgZXAL54ybfqwjDQrElskdg9UWGghtGKADYJY/08W4mPtXmVruzKGJ
o9CkpDoT439kCx7w6XlVHjXqBb9egVhfHGrxCsRm9ggp1QDvEO2luKFU46StrSQq
00mNSjPQ2UqCc2RqBaK8fWpCPj5c3ur9lZ2hJR2+eER2xx1XmBNBp2VGREK8K6B3
9JXmF68l/fxhZPC3SVliZMr+vnRmIjPMzPWcg+h8xv2e7pDSyp4Jstqfzn1B6SKQ
26WEt6IHaELdqneNIw4Kd8oSOvx6Olt4vTrCmGOT9iPfKAAD0uGaXGvo5JllrRS2
p06loqHzFB37/fto09a4SaXEXRi0LfIxdCXbeGaMvBkouBtVwnWVNQCx7hL1knZ3
EhKstK/52x7LFQ0pih5QHSl7T+sJcAeonDxLVMl9U8xsshzDO26rZkdMWiGWde0w
JsS2T8vMKZ2wYCzHcbj9OiQQkrWrRMjLwYTKouo6tDpfw+74B4DY4uVXATI7Zq2F
y0CLKrPnUMO/uPA60GMLlAX+7sdqkwpX1XaX8sAzEzydGsaPbSAbBCKAkW7NEGcy
PC//7m57PYz7U9HRIcxa980+C2iYN7FMqUnyhflfHAxScXe1Iy9QbusYgheSbUDU
UTUDmqubHhl9DAztSRqLqccX43dwdTd8RqcO/5IVXdnIErGRA/Ja4pdpKjJsRuV+
U3zNI4VC6+HTOBpUTNmEnonXetVyEerTms3MVvMQUIigOqyJFjfs+Er+bqg5MLLx
xiFAcEFi2B9DIPATTPwadMWlV5Dl73/LfbJlhW+8rsJ40C2Xgip5fSaYhN93IiIP
YMeFkvsfq4fz/UM1NfgxajWS12xmwxDh1oWWVGmKV7TjDmat35MlaRJcsfDEUZ16
AYzNgKD7MsjcAmPh9gguOdbk5rfBuCcOPHucW7rLeWO9wo/1MujfPUD3s0+AIOaD
moJAB5D0sTxIlPXMLaaUXUyfsKr/aCdFL1LvF9DSqvaBaErVivm8rwTpzcWZUN56
IPu7pTJoHpWy6ueLwtRbX5G9MI+qfeDvndAG4C+fuM1ls8zKyg0yWxxFn0iD/B3s
TNJM6yJTpdqsK52m/Hqir/1FM+MkTQqjK/d8vcA+CM1VKFavgRVzePd0C+69/0Ry
FSQmy2lHsMcYXDmtJv3EELdV+HUjJ7XMbsnI/tTNW9z+UZxuqplQ8EBgGhifWfTa
0UysUUKlfU/v96sxZruZQAHcvBvT/DRR6CYgRfv2ijmnRm8bF0K2qD8FHUc8p/nR
wiaUOs4SNRw9nG77E12S4vqRVlULyQFAqYJElYDYbnEmE6bbGXbqtvwxQ/Uagzy6
arP8SZ/wA/38Bc4hCecQaIZYcz1BvusXT9nrGFqJRR7r41j/Te958nXMCzHV1jul
eQomf1M5uHSQ8N8o0boyW7zTATZwRheC5cQ+qcHhHfYbLzBs3OV4+CeiF8bCrvXS
tIAzV+ntZT7haQJ/ryRZ34I8DvwWstIugCHKhAykxRIJpM7CMlE3nr3RQvJohml9
+EClXnkR9Ng7Rsr0ckFLQNrn+T9UnoRlR2girj8mbhugvKt0lu9iFz6j1TGVF3RX
K3OYS/h/Wne7GKwuyihmtNdUyZkRzYBD2pVfNhXafqWY6cXlHLC2y8UhJVVcHpuI
c+xz0qpqnu9kmRGJxXKclSl+GSE96mguk94uO08QAEWx1VfwZP8/p07cjoo5z6dj
jkP+uUDIIDq5aCMRkHYjf0fE7fU9SSd6VH98bHj34+YKL281/6JgCq1MZ5FyE040
59YcUA5XqcILtCaaWZ7DNmls4iJsvtBKqZnPXLQrATu3yVDSIvMNH2yeoCY7kso6
wmKIGQNDjrviTJc10tfM662Lu8dHOiCcQUsltPleTsH1gCaae59PYkDhnPKsVxs3
8RqZrlGolSLLl1aLeQiwL6f9X5qWbTnG5/GPYCUWjWT8tHUR1BxYeNvpageMt5Qs
KSmBoIk74GrrWgukfG3DLj2RCjYdq73SyJ7AsSWDgO0iec6NA2Rq9oxfmJgAA55A
aGbPsBB+2oll/j51r1k6OqR8Q9RSegBYp9BFEEm4TH12UxPfuvOgNTS999WGElHe
SHjxCfUlWmT/8Iqdgt1t4e4EzjhQvaFLVubLvSeggfWrZa+kOkFASHd81CasjLyG
6bLzGhUI3JDipDDlTsmPv/lRAbv23ZBevnbr8k0fbee7leiRcC2wmq9jIIM5U44v
oFJYyhXr+BbuiWw1qHfDeBd7b84hWfBF5ApGNHpVF8vl3EBjxBwAKxKE2DQZJCrx
8sdR3t270qOJ2WvTkPbiZj4LmDjn/4HHG5p3zigrD0LGm+WfbN7zNIfOb5vv5aO3
IKQTLzVyjdPXx6majnOj4W5Ye8eFF7F0VAW8WW0dorv8yHES09RTOKiL9rllhAJ8
n5oE5HiUrrCyYx/9QnJdlzO+AWkKWKtZEsI13ssYO4kFB6YhdtwDLugepSLHKTvk
axVowIajYobQ0F1LY70Mo7FeEN+jMUPob1eXsFDQbeQFds6fnrv2kjiN3YorqCOK
VRR+jLRbOHYpU0brGOKEjo1CTmbNrXjOlUl9I1ZIeTx4Y4Hkn8Q14YtBpmOFv/Wa
MsqrUChIRhDdD4vmtiwABBNaIQbpz+nQkvFhsJ7Yzq5usx7pjd6ejdaA80NcMYdx
lWK/vagsetepv6Gb++uModn5R1SzHOGIbzNIFpUTkVwgo2EifqGKuo4pOsgyEI/8
hiS9VoE2pIrWZOJ2l2a2YAdXD1+PzChBuBB1SiuRtiC+yK+2qiZReuITDYR6tQyH
7Xqh5pnWv/9SgQawbmbBkOwL5Kykq9e3n+xNjP9yNW0a2sxL22peYXUsV/Q2Srp2
ibjfAWLmIZxQEDQKwpte29M9jcOam9NF94c53+jRUg0YYQ8T9YER5sYGx9jYjb0i
WVlcdZXbARW9yqOmanl2gA+IfvBqBp6oyDW3Kgs6LCPVPv79EqSumGKqstcPcXJX
TwUrbc9o4+U/+YerGLEwFbbCkyw1Mohiwgx+B4N9aF+/viSNdXfKlC6BdWGuSbQV
f/d6El3C4myrhnD8wb3LK/BgBjHZbqZaAhSXpzVF+geZ1eAA7PFJlVLSeRAJxnMZ
zs0fXBCuRucwW5pqPKo6HpwI0Y1r1qQfKiXQ5Eh2cCK7T/KNnQo2XMSE5kSLTa/v
dC4JGNj7b6cHmOmGM4Qfu2rwfwz95Q1pZPjEigIACOxvG3//iu1eaV3ZUN8TZmFD
v3UWXQ0OAB8hRQ/1YoFzkIQ22uAWSaHHNZA9NzTojpDUQm1rSm7QR1DMsxQU2tOF
+54IMDtRCf20viR/7/Lfbf97SNZJLnkdAKv9LFz9FXtkfKrNgknDrLojbb0NE0F0
R4N+oR+krENz9htiZpmiumYZYZytVIhtSPyxi6yy16Eht4ei5TeFo/JJhKNy8bT/
PIfy0/r+AIjkUcQ3AgZXPydXEcioeQOm6AsybAyKyu09LSZMqI9PQP5AgWsFflPv
CZmYl2vHefNyiTaEsZVEsnw8mrClrxm2RGaYvAJe1o/hByuKS+QnfS7Gzx3dna1w
IwIUQqJsZ/sJkOd4+nXalFSmA60/6TV1jYDlFFJOnSikBdppy4v+zhx9CV0LbJ+K
kZoR9jmRmog+Pmiv/r795mBlLSh9vT2KBIhqHbhSbSSEPmTV9n0ZKAj7T0VT6HKt
snFHorw47e/kx+jJr68GKgr/vDQD5B7ixIvAkxMDYld2HEMhPA4og5WkX1KGIKUa
dOMI/1+ui6ZjORv3uw6oDxVVmScmG7/fpoOtnpNOt4XlcYLsM1/TdHL+SXnK+kPj
lNI1GF+689TXWRt6S9h0lSkeU4AWeFVPPHs3sDn/5+pCGp0K9wZbImrYTMQPAUSB
q8w7+CVfQmwaUIOHCZO5eZCbbONtYekUdBCFoKTe2ST3BdUauX6irkysGwbjRV4R
lrGrN5CWsiLvuv/az1NQK41naYNyLm+kP6CpgyBEgNBIAl4hU8ZrFsgIFvZRZDvj
8JrAN0EabaDUbn9lpBuTC0flZrPf0IhUXq4tfzqcQ8KuDp+FMvDQ8rBwGRfKrBPn
VmKLUHQy8UFzGSy3a83DFZ4uSsshR34Gtb+Vg9UiAPFYUwZdgTZfUE6wEgm3Y8Zm
my4KIxTHk5ZEE86Tvzup96z9OrnTLDs/nOszJIPhrxntM20kJBFHX9XyCitgxpPg
6BEhBbBMqpAeULwtowh1hrJ+/eeCSASjxlbIjnz9h/Xp4G4HQpA9kl0AAyJWpqPN
leH19f02jPsE1LD0gvwZ/+sjfa5ZDepxhFVYC0rBz6qbCJAdfU50mzH1PtOr7UOc
BPkNS3PWJrk8DFqYxgZeEZPq5mHD+aZKSjmhCPiysu0+6l3A304WKEP1s+YvT1P8
5BSBShmoMpOqGyyFsoYNc/0c7q9I+neHfE1BaOhF3V3qzdkpT/PSwTIUOGODgVi4
/qpvMW2w2WeF5bOKGpbBhAKgRN9K4ltFzf0pthN6oW3LpzoXSfWJFPvyuTW2wY+I
pjv33v8QT6ulNyjrIVQkR8fibnLNda0Zbl+wQZ/lOrNluZwZMUyIkw6X9hAv3GB5
PfRO2CGVJyRa4uyEfWnQ8RTDk1VO2pknuAeTNHufz//Dwm98XIy+35k0gtYRWbDB
3SDlQ+l/j4u5sxZ18lEC6geBi1ekoe/cAUsrJ1kLDilTvqnvKcSd+v/Lm0kAkf/U
welJgc7ZaNQIZSSmZFUsLCRN924OyWG9ajyOxsOb21tSScz38vCQs8zGbhXF9DIM
9I66HPIGG0QiGZ3kQ89Jz80YNlkhYWLTZvK8QWcymz0L6A4TRFzavih3nuir7mU0
LW19qLYE8nvVTbYOZw5LJSb93XHm+QjIwnIompTiMEBqCxTCfJ955TeCggPlPd7n
HvsxOjK6D9Tib71SioMEjlhtRQWCoMX0BlV813XELEyY6KETsn6TcZZroRz6B/+9
FpkxOeauIFQ5g9wVcMV2rvjn7nnE3V+kPmKitEqiumKg7j5Yia0x+4DHTDFJ037v
2kEKEAdjjIe9UE8GTfpjN3tFthKxqUD2dTDiDgz1EO4k/v+6w4Bqi4Lnoe9ykLJ+
2KmdFPHUsK/h8aXqi2IAvJv+DKj3vaseuIxZvJEoAgMUTywuCb8wSuo8/cqRGY0W
oRjWcT9OknGf72wEi8MucS5WhylMQvzMtUwknku+vyvYuWJFEUry6ugWZf3QNRME
z+39TeWgSFBKrTMrDR67cbEWNQeTPGff5k59gkTbSQK93l9A5UrAk2ZrVEEcgO/x
5HhVGecQRksK7cBF/AhypvtEeZce4q2QHknsqhj2To9H5NtlVhM0bSBjnymrqdLX
8INzxl6xSEh+nl4N+bXpOqxsbkRN9T/NyCf9AVQHf2+fsWB+jSfO9/kvXOYmA5ye
BTdAf+WZm+X8kVvWO2Es57w/QlSUWWFpHkr/veHMZH9yfAbAGoIEGG0qA4hNsxhg
UI+epfvafI5P4DilIgLfXxBb1yQW0awqLsE7LOsAW60hLcuK8Mjq+DujmVtrC5mX
6mc5nMtmHQDJ4So67VzV8PpzUB2GiSfySjRrqXjUxWMGJx8hrTRp8gHfke6gfcew
/ia9CKPAF+ERlQoLJCzQZYRNNoLL5J5LBjMPhm2TzC06uW28hR2WbtuB+032yznE
r4PNzH1HXEOH5NCjrrF4z9LPqxUj2hvGQ5Mtyu1pX8S1O6+RXOMgLtbEAmRTlY42
cve4y4d1PmnaM90gtisaZzeL0wnRR4rXFbgAkkhZA5D9paJWkY7GE4x75C1RouU6
uQJwEqoT0aMTcu2wimdpzjLjVZ5NJ61qqaLTVjkW48lOGlQwu/A7BRUwjWgaSd/c
8ZLQ8emNGOpyLvv61U1a22saKuL3x+JiuqzZqfllgvo7DqXLNaLWVBf0ZegNOEZk
UzouFjc712OdAWg7hNVoKPgnRlsXfZdwreHhqF0T/NEQDiD24F67c9gBXktv9Uu+
4aYCuVD2yGbYu+ClaWXUA3HNaUDs3MAWr8MUD4Slo3N+4SFxjNwOZ4bBeg5hHFOu
Dt+W5zoI2alz6lMx2Mm4PUO7smt58HWn8wmFBG5JPCZMMfgtTNrPcKzyfe3HbpMG
5jqi7THaoCYLSDNu2zvPO9ehPNpbW2HyACKnriejEGWLKgOVbJdaqhjm47N4TxAu
r9TPCcVpAuQePC+l8hihOd8nxdNCimX0ire+OY4v74QnMbw/3fDeOqm9FC5sSLZk
k0s+C3JYYs97aysSo7ZUUUgtXyi+PfgGVe9IfNTTZ+OFtTUMKlEiXL8WSWhaeTXg
RKON7QfJ1I50o4Uq4Ky7yLVQp7xEYxIaGZBhxgaV7oePJBosCdD65gi14o2sfhfm
1ugB6cLH/2Og0NQE2XKlvGVg6frZmjQNa3APerjQ78T01r3R+1b2ORGS9V5xtHGi
4C+y6DcZhMqojjAVuFHc3sbPydowyfTAobc2TVdOQnMK/ajMA2kY5g8En7YW6Lta
HdOGSl/7kXTHp39069gUBDECl5pQPNezwfh1ce9OyHpngHPNsjZGQk3pFhHTA0//
XgSq+XXqIQQdwx9JxcJBgYpBdmP+yUGqNHtLXPHyyghfXCzvQXJ9plXyLTqZO6OH
O0mxEdpKDmuFZzzuHkYgq2tIjpXBDuLLEv0wWUoBuOo5U0onyp5adrDP4RDR6o2W
EW+mHNeWuGnjQN+jPa3Wg55uoCsEEM39lkh6ilLERjMirxsFbkR6ZvwTrBGi7/f4
goyc9bem2GR+G6q50Mq2GJKfvqWbizMJ4XgW/1YxhGBTVXuuPozeLYOM9kuf4qoV
pLb0h7x6yYpN/u8O0PeOGad655Hg4Zlmi89WMi8nu6GAlqiafEp3iumoaJ+qlJb6
Y1hC3wW6ygloMalyR4E8RTS6Tw0QIBjvuBG0XvdjCG5cj0HKPJwT8im0p/S41YjD
4HS+s2vLBz4fPnTImrnSr2FUIjEtq0ATEYYcXB8ZilmIULED2tTrC2GZ1rKyD1wz
SW00yWsZsR054mMi9YeNlM/f7X6ISYwctlWYXXgIx3UI4H2wk5RBweJK0hzxAWrg
s0dLSJ8kprf76RqQPb7LhFm7vMM2Vw2eNMicL4khOyu8CEPEUYdDTgze3E8brqJ1
b0/jOh1sDIcrdPgba/ovHvkWDQOWcrfv9jR58eknU4l5w3hKQcT9x3ZLqXzPXUhv
N2hvAZlxMwT1BQvV3IejGwVBlurYr2kjMbvuDuAvG7oY0ISAw0ABCCb3N3kAj84C
lTMr1bvhs7EQT4EmDtqs+MVFGno4NZUd0R2UtEwj0cyrpj6mj2C6oY795SEGX/zL
HOKXSmmK0h4lJWuWs2R5Dqx6e58mns10uoDqrga8bGcatU9Sp3hl5zj05DA4J6Gc
M42BVFNq9US9cAVxdM7aVCm9mYn3G15eHAlZS52GcRlQHu2yg5RJBBUkcXy6MfMM
65svoJuVtrt2K/YO6dznuMMzL8DHoTeYKMGKMXiob/8xWTYuYbZf406xxpZG6+qP
KqUlwTNefeg7BF8FsoqTVeMryoeToCKP3FXK5ss3XofiouQll6tg5Fu9t1PAgS01
KF+a2KZA0MyTfyS0HR+lwCIzBzNtAK89Om3bpW9ntAKA8uKGSnOf3E942mqo8uU0
w6Fbc/4xawmCKBGNpoNwongKDC5/DemSss5YHk0wZMktM7ApUXmGd4XeumnIZGXq
R579VSwxr9nqBf6pU3gZ+UCEGE6hdjrF1CllbkZuBTdf+eje6uPFACNyglHtW/Kn
qmcLoGsnv8p6vc5S8AsrDOeLg1+Xs37GdxdPHoGWTk9PED2cuEkBawUzwT3WtLms
KchYz+lgXLF5KAEfX6TOgBjWI+ke1MLSTcZdrMcICumPQkh/Q5ZzLpzJO7w0Fl9/
bPlecNZdm3sDUm724BVgbyZDaXh/D8KEHT1QddmVYAQbWjWntRw96CYWe+FP5xjY
3vK/WIf2AOKpJfwrJWznTtZpDY2crT1/pzZlSHChQUTm1MLOtodpD/iScTJljA8R
v9T3N/Yp0CQ+EbgoJuLTnSuIAnsz8vbm49A8MNYygt2sGwc8rUISoHQv0IoHyXcj
a8UbaN8/ykx4/7caeH8xXHOR5ejaXcMCL98I0zUQH17GPjWlmTSUdNNEMuUc1q4K
Sy8cY8IpNHvrMNcAEqlXW533djLsXReB/mtmGyB2Cu3T1do89F8WJY3wRIE5k5IU
xx8naFZUedtUuGy8Or5K4RxP+qkKUtZ+D1hLaZbHRfOF6f8ZY9qb0iqenMTmrTSv
L7ss7w7/o/5KKxH2BW/jGPchrhoFl+vb0HLNHTzhN299lZjBgiADt0t7LKCoZLWL
yE2t/Kuex/HwoMPCyCmslIISj0eixWAD4CmBK8DcX0cl0XW0ec+tnAHrU4SSRVdB
dBCSpjzqzfX+e0H+KmliYipDei9BHJ1b9+IKM83YbjHtwhsQyY0upNZMsjmXBvCp
HT4QCEHkH1s1nTyYWfJmjyPVVeNVfg+YHBbBhAOi+IHq1vbvOt8fQBz+x81HW1QF
UaLfWLP8QW3GecYpKmyU1pGyE9af15/8irdJwt5eNwW0tm1Pi/UJxVTK8TiL6k3w
zSQOmILo6d2do4hlmox48UZ09xK9VuR9EecvIQhCjF+s1qr5oeVKaof/a/3OuHXV
TZrMA7WanEKH6K6u90y+Vxh0QMJliz2TsMAwydA8Kbjo3gRwZtfrkhtQncXgwVwd
+Nw6Xe0P9GuAgoZnbN37Gra8/CfiD7yTYReE7WCbui8LdLC8x6IyX3dCKNuNZziq
vMOZ0DIYNZlK1fQRym72Ad50q+Vyz6sFY/Ubp5m6DTGgY6zpSPeXxXfpGFMFJpyT
EnUyf+7EQiBdq5CPNwu0yi5n6w2vHLHhyJ+wcfrzbnDOdBI//TJA9w+KmfIJc4al
Bmt14w0xvNW6/pQArTZKAUCoKW2jNXb6RrsL0MTpOj2I4pUvayshSkRXKLEWVLgy
RDKnhuImN/dGzFULW9lM3BbB9OUoLHhw9XUuAYAxNDLQ03puhUshgOo9WbYASVXz
2SVEYi7HNhLh/FXPL1hkCvYI+5M8niRrXih2W+bdE4U/9Rlcf93A0c5/m2Bw7py/
olh7GGyuw6HJO+bAZvPDHYzqqqbWjyO+TxGhHwWoMRorVztBpwCvxZZbKwXRj4Wk
1Y1BuZ0NGF/0buGb7HPkG2Smy5/vKRq55zU50IC/N2oF6lEkh39tQCwgka59TI0t
XqG3LYQ0cFin2Q5s1WYWwxHzYgqd4G+SFpmUFTI8hSF61yIeQ5ao2HB/PrIlkGt6
ss8vljSVnLKW6ADVb7lGNKvJbDftp6nAEu+RPSXrlu293tRqsXQUancb2HI0H9dt
9KfLF+t6Qn06ahppW2nyPHt9ieZKIpOHbIvREe8BSb0gB+t8mNWvb16a2bdKS9nl
Pi3mHPXoSs6FhDj80gS7ewdzn5LQsGzJkrXQDSFMvRj8tjuKS284OOfBJ/vlFwC6
MRs8iOYACbglyt7+NxYKbqD4gbqMnGkKnhtjf7dwf8cbxmUNmkByBhgLp9BDe95k
6BJXnlmy3hpbAkZidmLCAcWPl5Jau++AVGQkXGX4ANw3RpQFjZa9p6mEqjsW1iYd
5nuSdRh6bzYwcx5MfhLjLpmBQDQlXXzHQL3wbLVL25X+ZATWCzSeIlY0CFFna5eY
5OB4kyIASosfIO5hfoG/EZH6BaX/W2KTLHlGntfrykxDvPoPEXV1axX18RaD7k0U
OH6XNVPrYgfg7CY2saRk2n7O5dspRCw88RTEXH1Rb4Kpz6XixNA9FNgbxgHR1bgg
B/ViO/+neI4mhD/Fhq8/Rz5nAzMjeAepETj5McRh+5sXn+hI6k5jBDILnVHWP7RC
sB57wWMEFxq1rFNrsc33c93of5OGKZSMNTCbu2EoXU2t1O7n6SPDIabol50XaB/1
LSx3n3CTWAXMvB8dLuX/+ptekmPuCxXVhCIHeR7pemXiFFiI2yAUBQ34y9vyRWk2
yhgCc6kZwGXsYzG9XHEL2wzYjHgM4oZ2Q/7zxDQazI6FD+V2pQQPn263w2ZcgQag
odNv/3azqr28U/56MzdNZaw2h0fUV5cW7kp9OtAIq4MRzUmU2WcB+O3vadrNSgx5
6pWwlW028MFv1y2bNH4UtQKO6v43Q5TjTCOUJlfMfNishLzhlXUWwbw5YNHfLKxM
ZPQq+qorOWQlloJt3Nh9FB5sPXaM7cf1rXd6e0GB2h9jvihYWxtObjFZXYXo2EyN
31REfqbCgJ48A8byVkFvQK2CSPkIqXpQSiq55D2hQW71mc/HqeCyDhQGW64hkYtt
Oi6UqiV71AU/7WsOKaryyxTQqlhln6FG8tjBZDQfOs6bf/x7/JGO308SHVpTLOFG
58BCK0uF3Zr7hi1KUlKD8YceJ6btqxROuj0d7VR6n38uoa+HgAhGRFwJnEQploQl
Wdb9xVOD2sYapEXdAfXyrrZkpy0F6DTTBHgl2CR/WZz2RnXi9Moj41uQ9PmEggYg
6SPI/fEspoYlhfnSwzGGG0JKiumQYo+5CdnEjfqhbT9IqAhk9H3R1Gdp0nK9KQdh
bQ0WLgauGLSAip1S4JSMdEWsgfA403H4BE063cXcxyStmlhPPkU68Pp+Ehlwunwq
jh9heVdCD40lbx8qIG0KzfoUKt69DUnobyPEFZf3qgqcEtg+UN05VgVVeB+5UYWl
XGPCoNskOtJNOQ+++bWhs4Du8G52oYdUBvnvq6qd5VSyY6NojGNhDoGnZ7T/lodM
XjJD66O3gve7J3Im8CJZLBnfdkVqN50eFlGF8aE/jD5+yszIBL6l9KJxBdj4/mX0
jJO98U5N0nt4fX6xHD3nT1tOTz/ci8hIaM+5cjjra6lCrLI/fKKLaGMYO/tWAfCV
Hc8QdbChIKJem7XpPD1QiTsX1GagR0bG/0tN+lnXy03XcN/2f+zeLbLapMXV1BmF
pRTiFjCoIa9b8p0zDk8ABVh5qcha7noa15tzABeJoIRitzF6zI/7+cUiHga5oMJ+
k/cSiIM7XUsxcdLElIIYJvFAvxRm6N6ejp2fcFEENhzEU8spfUd5mULzi5QImLlV
/K8kDBCZEAK8PvDgLTF5AO1knjmfOMb+GUNoR+Z+qgPSM/MVSukIooTPAJqnxxbf
PAr+IDtzmsBEHkdRuBthIcc1PWguYWMRQQmLpa8e8YIVthhNOufrUuQMi54fpPhP
iwnekt1iLKz6MiGdHXy9iKmZG5Mb2e62ntJOWw7NWXylqCGe/bC/ti8hL0rz2GJw
QuyOITmv3pBa8IYGuBT/NzXylra81QUFjnZdxUcqSAuSoVXiIwaIHeIDA0w+vBb5
aNbDAvxjobQ9Izy2TrzbnRtcSmsuYLasykxfpb7xzOUZnCy8X/Cm4cbZ+28VLjs0
G1VyYFxKlPuBKXnEk78TCmMlQ6tH816s0LnihKBT5I/i+yvBsVanZ+4gMC/DQz4e
xCNltOc8aRibozD2k7vwXfaxkpQoFZUJ0aUv7BrIX3d1YNug1sF2ZTpfQiX/kGWv
25zZ3m9tYAhTUygucGIbFRccu5oOZOi1Qw6d+rNaUNploA7O4pnyK3Ft3d1QhoA9
CdOSAZ0vbDoAkei0SSYpb+Psgwk4wEVTpSK/nGqfrtHsqmZnSb/yAT0Nfe9h6nN4
puMC7+oKhvc9x+6QeY7HnMqR72oVDULLMAnwDPhyMDF4cwCz90ft/imfkCFnLY/O
78fJnR0jtNqzLhhF4LgnvJ6jlgGh5oFZMRENqwwIT9GvX5BmCSy2zFuKRhK0L/q0
1NkgKqFeza2RpNw4jicTVL1RHBM++FZ4MnRIM9TMt9gMYlfy/bxnsYkbzQhCG3id
IiPvF8hnWXMrYvIeVhA9vAiMKgJnOcxvIl/o5sLMweJqXqyh9v2DDiV7nGVflhRA
0vOGBMUcB+wjIO4MS2/uYcqmOToR9VDkITkArNspSAHX0esJCIW+7SKb/+qAS5sc
75twE9arBr9NQprJuYC9fPbxJT+SyvGZNMXKDkMWUBUuqfCvT0Bk67gGtr71k8dv
RzZD0lwenrZn5mtfeSXrJPGQ72zcn5ug9ntJ0KdcwjcFUyyqo4wVfP7fueklq3CY
+Qn8UZvkF1BHrmt3nJGvqicXBFJyTwsICdVX7/FFmnXF6dFx2LNHyNW2sAqXk9yM
Md2qFeUe4nkY/n97mQ+JUbsmd2RdVwJb3aTpkBOUFcWkfo8KA56WcgEyBiXS+Orh
eWXGmj2LiKK99rO+YUVRQbN4CsMRBmLtqkOh54hFimFTSNpbdWQq3hyUB6ubXjtk
CJax6HOi1Uv+i4KY4rq65HxsTzkXT1sfvxyVKl8/eBwun9+DLdnoSKPRwMRDo7Af
BT6x2/nFJBVOAk8IgEGDVfPtYf36ZHhlEnpkwqniWPGYzM3Rjs5BxGHCqINfwqY3
7KhaqfRWFxW8dNg66gW99kG5EifGmh+K+L9rddjtVakGg7wdlhPd+o6P2r/gMRDe
tgAbEWumaJN9UbbaJE9Z0Frd2XvU0wR7AWmwzRU1tSyuDKmNOaE2cZwJxsXf84EP
ZrJRlAZ41+IqadBeUDXv5FcrzYcgGuIf29P87FnmcsX4nBK213c6GGYrIHIdNwsK
O1C9TDrDFJXvJiD1F1Nl8JxrdmLbPNG2gFyBnR/yiz23StslhfFGaykmxZ4wnUKP
IXBpEhrxi7AHvNLTa4nMYQePJyaE0fSUE5Kxxdl67xiPRDBh00pqPlTVHjUqggND
usNh4iLFqOBPFnX6bh4E/9agnWWvHTUMq6xFYDYfDmofLaZ4w8jSvszPYXJ8a3H2
R3qxFRelK+wtSm/RrC8U7C45hLK1EPiREZBKfMcPomNC2y22nIP8GkFqsGnF2D2P
fXvw2C5+eDFZ4qVlS9i3gR1IVeSonvNjRVr8uAPBrV1vtT2PCKlg2Q9bzVkAe2KH
8Zwauwx4ug6mUfSA57jamKSrYiITuKRwTZd995JgWcWHy/D720EI5EnJ1pqrzWVS
Siw5r5R2twBsDTgU/vKPX28XYc0wb3gNVQ4waQNw3GK59HUACU0Mts2lDLtieeFP
ES4z2dVcPhH40dXalMo/uujTB2Of+cp21IUxSqqplDdfL1uVEPIjdFSlHI1geC50
HVx8wNE2HXQ6FDPp1q+Wso3LcpeCJgMUhYbmltmshkoEtEG6PSEiOP4s1vtk3UE3
LlNwdKaSjlYQRnmnn+HIxIL/9dStwJzVrNK7+y+1tf+HoD3Z9S5AZuT41oZkH/Qv
GU48L9kqljT2rYnWP7XvRPv9hD3jfR8sSr3hdH8G3ojyZ16QedIw1UgCmSMXUzr/
cCZrY/xeDJgrduvnWRmobe4Hs8Uk+PUjayv5kd/lNFlRAvwLXPwz4fVv7UHVVpYj
JtZIMh6ioYi4GhxNUTo03w0h9bk/IOl9O7blF3KExz/ZfIIsCf/yy02AnHgQMdBW
GroXce8BVZ7KkuvdBtoRq3bJL7TzHT14wzTk/rhjeWFFXrhb5I9Xs8uP2kcoLF0f
yoeptftsa2BUQIX3CsUExgUvbQvHFtAcaEYfbSdh2VGx5sOQyK//yRLskviR2nT2
xbEEGENgeVdXHQFC9VnnW17nN5y4ZooFj77Zb3NiTtF+CmUCyEfD5w/RmmglXjEp
eG0nC+VO/EoCPWIRBwyyobJE35U3zBfNawxuLuN5WSWCCRh0pOAamfc3Z4x7VU8I
rbOA8er+iCNRHHBYpjiIqqYL9JB2aEWbE40mcI5P5fmWlgp4h6cBwmBEEDpXvw2R
uEos5W9KTn7OXgw+iVLU/4xE75Mx/O2HDHbq3agzJGLIEMvx+5akHBpl+TX6KHmq
G7NoeJaD7+AWfCOB6xjUp22FnyfH548RdE3gV3NZIp2tJH00yWD5pLVUhgoK3a8u
cmqqphiJ2qsmHc94DPzTwAe5M6ExxsAurVPBoFoZiuHn7ef4iaoeRH7KXLjpj5Io
JO68+uUndE7i8+G2OVZhmrE67vl6X/OCKIZpR1zBqpMJ0NUEol+liW7j2ixfEVnC
MUQx/76N+Dlr7/EbEhNinGmlx6tcT/2OviqeoQqjz08FVSd4781Rx5PKRvYVgC+B
LQBe0Upxi/J+5HnA2ffrsUEa78dr+9TaTuMEapi5hyzBPJ2e0FEFv7GiOIlZq+dZ
aYD59ce2d/R0t0xSYKacuTMNaX2H3RdxYT/1vNmKIP9Nz2gRHRjj/vbXXYTNW/k8
yGqfnD9TkJnkevELJmQRUwG2nYoZYOaIZAfVYY4Z3t3Dtm/UsY8bQQ1nINlnn3dA
0f6cTS4BBZhTs/yRhBhAwvwTKjpSku1rbHBzrtCqHZKlpPfK8eNoGoqUcy/8bO+H
9AW6NmDR0r445s3UtIICabTfooJwpuvgd1Qf7xid2aLvMrVlIUrcsbkKuXCHbOCY
l6DATHQSIs8GKyliI+uLoZy2sBEAA98jZRSP1Ob9MIbPAIPnfQgcwuNgImIcMnzl
gtu0bS7+BvcQYafMKIKdDMk+DEWeIIYJxxSYUItNbwFFjz9Ci2rz9MFRZk9LQJl3
Dr+xhZwOHUXY5RFpxMV/dU4pIKm7TCwhK20jC3DcFrNscDVse3Wxm+cq4sil6nvM
JxstfMlx3JBf6RQCWifMgsVLuHJer6+k6tZRjRXijEC5pTIyP1NOqsfi9o23S2SM
F7B5unYOQ0+phSkIydgKljEScruiTsJj7eBzSI2zXNY7DoPCuphtzYFUT9S3LjfA
vMmIh4kY7IBsu81Z+VB9hQgsU9M/B4P1rmvDl5aOWbafiiA0kBfnFW4FbU6igpnN
YUhdfCMt6fccQYRd9vPaPQPShCjPSpGNz7SrhwzX9+E0ZZXtTyDrYNk4jBoj5YIz
36MzdtUJQtTMdMHrFZRLsF8lVjmaDAvKb7/JiX6IYK9Y/0Himb6PR9bw/pVl1lVP
5yMDXVoZaVnB8Su7acdhC2+pWSpLuYVwVcFxoMgGpyVgP+HFYn1wDkwnc9TE9nDa
sBPOV53E1FIA6OeQKSoN8IFzclXOB58CX5j8hMPF7o/P68NWMCBgeW7vQ24EDH2E
xwobLAQolme26mxKyoTSV1fCB+Ew1i4uzeaJzNltIKoEn1A0+GzlhBWC5BANtwLs
pbwLZGPc3EDVwZ6vdI6+3pqG029WoFaWA0/z9LjxxPUqEfQedeeIt3Smh49nm5nA
TMVg1AYqmwrJXEj226s8syRRsF8hqDARI0JilLwwiW1tOpkutp9aOv/xczxJFR+J
hp/9HFngXElIl3q6XUOygesD5fN/ztpxG6HUP56usjlAbJPD6xyO2TxqGwUaGoSf
qv2LHQMzxQYbSjMlCENzMPu3QEz2i6tF8ATdtJ0y864CkihbWjmvUPSFDic8/z/E
vqYzg+0cMHBfe4Qt6TsHKeBYBzpCcT0eWUwo/LRaZkMZq2eTEP9yXuwV6MR0dUJr
mcGC/Q7/OCTwTwmreslqwQSNtj6FEn2rxnYuZMNaW9kSvnnpEBLZJ9MsBotT0jMZ
8SrtnT5O7cdIOp1cZdl38ma/ixYEIj2RS7I+tp+7ATPgunF4ClHFrhXiWUl6djRf
/KO8n0FFHNJQZJBFJiG/LMpW9kLbWVnz+NNYofe4eHIqxnzI1YCejy/XjZ05tjRH
397M2jMZHe5ptqUNibioEZrM1EIo9Uk612sNAgKyyR/R36gKbJLWGbBIXp0j2kWW
h56HhSNj16L9JSem6zToG0lzeJEPiabKaKwrGRMiackQS1HEpbVhuR2t6QdtrW2d
1oB+hyW/+bCx6kh5tY2Pouje4mVk2a5PQXpkaepEdrth9mN9CFzesXQjKrecnzbQ
KzLNyJvrxIcGdsmznecW37G0z7imyEqRBkJHf9+AC5mHT2yXzla8ytPP+B9x65J3
/4GVCrQ5LFD40P2CKEDZprdOlWvw8wjRnKTp94XIKqrbjx1Qglm+Sk+a/PaBzBdt
3MpfA8+pt7iwGh3ZifwmL1y4v0v8kITd3QWrVSSR3JuFp2lpIgVn5bMJYG5SoFLJ
STRj0N3l06cR7JXLwNl+mjQYcU8xGND2UKD0i1SP1PtyIodLEivYZlerNCfnltBJ
S6vPXr5dLds7IHuIy+RsqVyCRtL5Y6eaqMAVNLMP1qHBcwQJp+Ub47/zOSg83E1Y
mGUFg3hMacll6MjUUqJj7GrwDtpg62B9OJbZqlw7j+osRTniIeziGNPnJvDbyFZL
9Iz6Pg2QhM1cUM40mQScmwGGfYF20KD1dJ7cAmIkw66qnYNLdnVN3OFEcP4qU2Te
9P6v1xNE3JrZR8wRMqHf2IS8cZfASd3rI0TG+174F6H5VcvBYVwFuWJOMckwD9FL
gXJ4Rzjrvmc30WoljkK66+F2B31Pf5WL9QPw4bStHlJ3EGRRQVzo4exsNoCsIDHc
rTZYLcJY4qsgfORKD8N82e2SDY9OT9kt/aIl/iPrOyDaSTkTp0buf54ICNcwChSJ
A3nViY4YMp4vXxGElneiygOy0FpmW45JBUBJKXccZ24ju08DEJqt+GQ2qmt2WQAs
wgSFl+04iWP9cAe/wcWtEglTXhkUUJx2+SYsV/ZdAzjaj9GyQWDi7dLhz9tpxNbq
Y1YB0QNIN+PoJBv5mFkzlEKID2o/OEgtgLgzbn4UUWbChfJGhcBNJ3zXDLbSqWd2
8egjPaAe0p5Ly3IKxWSWQ+h+eW5OlNzWki+ExnHshNUBDInPzb8/cFiMPVhwC9hD
TekTReu4bVy9Y46qewzGpj4uFAWzMqinqw1Q0v/zxRuhTZeCVIGJNIsIQrT9OKtP
6JTc+2zkqMGSxdJHu/IyhK0U4J7aZ3u5TULyxBM2RZSnkIMoIEuKy5UOWoord8Il
71WBYS4AUjBq7FsuSpHFJb6rM6C93798VYa2efUqm7SH6DKGYCC+aSWMLBKoerne
uTSGn++AKUafSXbiujeegp6ZctjKaqMgBdqtJflynjN50drkuyB+EjRilKkzDuZR
hwpZEJWjpQ8w7xQ1G961GQnRYLrzy/sQS52Fp8P03d9RFEGSotFelR7jW+KofGc1
ZBSWDQTJTRi1dC5vzMgcdjVwLccFrjE/tEOOS6uskmUAe157cC5oBGZ/j7ay8c2n
gjnWGKMw0PA5FN49hEdxozkWM/dO5VyXTkDWQaV76LXAGp+/bKj2ZiWNPcGNnTqZ
uQtgkVqtw4wkq88m42HIeVIqkDTkFJsISunX34qcFYY/F+Mv+R6tnnYaic4G8oi3
YbfmSYJ5Gy5o4CGN0xHgBvABOqEPR+DsRC7mwWcZuD7oRktkuws6AiZuvOfWdPMf
aNDRPLR/D9hm/N9ef+722G80J/Vcu3OFKwcVnD3+vsth3r38g5l8NxNvyQflZwTI
+y1k9hUYD9am1U3mrMBylglrTMz6gyIWQXL/451Oi4sGtquu+hZXE5nXDfvYvMT2
ZkMoN/Ld+TLtKYb/NkT2IdfULZvqVDlPJGwKHR8vCGh6fj3lnfp6aAHXfvhAAZY1
vCwQEaJod2jZwSnBVwghxJ6AdsQDevgsSQObkGbGaQQo9Q5gQdJuv+3RxygRlWL3
uVj9Q7sC9Na1CIM2P8/3YU9OMKoUFxqzizWzZFRJciVkREyYfpGW7Bd1aueCIPHl
bkJiVI7TDMFQo62p/ZO2xTPL7QETa8qtq46Dznp9U5404NMzbLKqpMraI4wD4/nY
/cqUN2QuTC7tlScNzgaB4u2DjUXfj8w7dPBrs3ei701GycGZTauDdBBn3+Rjs8oP
IuBptKrKM/NhowighKPWb6ABNYraQwRS8deX1uAMJ9Z7Dr6v63WpLkNHKiP+bFLH
xxLq9L8yRNezgJ/1NW7rcDmYVbdCcJvSWPXdOsw2bq5bQC61DQCbFVI8rbmpbSWN
facCpHJjFTnloXCr6xwhm7Si1xYkiJF+l7TsPoFO1KaKo9jHMmrOIW2mPXLZbIWn
weN+utgDkgA5WF9CdyAMcb8IO2Mdgb8vwY//vqxbc6KNllJ7tKSbSD/6cXTNrFvY
s001/wYENdVlm0HFatsC7Mobh2KVA/VT17jwUE5k89Q8NEFDXtsHT/kv2PC8098h
U3yQiitNfCa2NfdXFnKzuSUAL9kDk4QhVEK4WVbhxyPfH1YWkYrgs2n8zRiTDMNx
pazxvhXBwGE/h/35G2MiuD52cssy8OtFiZGxO8cfK3rNfBHd9XAm2/tl8WlP8VhE
6h1cvbsgaP7lVuzVzPWOuTPNxi6itGKByu3LWPp1whf24oR5oCjv+aufBMBKpdey
jy30lSNSzug6YMgAbePnxrAykjTUd/QSz+razY98E6rusL0QM15nQy1pWxXjQUIJ
0fqeMqXB5iSOGmRKkTgqOrq9xtsszGRccTuWWiqw7/NmmPIiEu772FLNc2+EClDc
A7OfIObPv6pfz/x1GVU6icz+QDv+8eJBeOOdK/faMm8RPgeCAfI9RuKdHl5XleHw
4cV8+9Gmev/mOa9EF+X5wio0IY/T22PGPGIKlRIu2tQM/PtPT6w4quTDANrLEODr
IRfFvbpfHc4P0XfbN70SygNnYCS4eFtpRKSRA2cdMzWhqmb8JHrwa9o5G4bzh0cr
m6uswBVJ7czXR84VTBWWP9tYpyX1XE3Zu5f2nKtGF7MTxyCx14bbNoPTjeubzASZ
rK4/JRq4nsRVe4F1QVtptSRL3PLy+0IW9MF2k70IrpoPZAIJsr3yNN66xGlmvZDF
4nTo6aSlRRSuzG9S5fdvz79LxXnqNuefvDE3LT+IGEjMKc4PaQ2g1soMhrhoMf6n
3/H3QXh6eMdsBhHKCeez2I/QEf3gOBM5uAQld0UuFt2XhiG86CJU42RcCEXS3umv
l5Dg0n6NVA/P3xmbAgGfjFxwD/G9kwMkO2u/CUZHL2Es0j4FborS863Wl/Ha8tF0
FLXMt4E8dRGq+In4L19slZIJ6Vk0olG2nLW2//RT4Bw2JI/6afMajq9i/ucXlxfN
by5pgSN8vqRCYkkhieyNuU8jx2wEJ9WmJLUL0hPVqCMTsK7KsYWAGr45AYupPS1t
GsauPPwPx0e7FrxoSb+TsdL1Aeabq7coUDDz+uHJCHX0Nlvr2qDcQ9QlCFIDKKMi
WnHRxQ6Xdf3Kfki1k9WM/8cyhJcXfEDTXvhb1jJvnfIgMsVnB34VrIIulslPwa+U
v7F0KZaoxNyyojNRk/bIUlwPFbJyEWNEgrlO+pkKjk/Nz5PXcYQaqqp7sp8SxELA
HPgjsHd0aNCTgcqIOttNLRZmnHgrcduDAKwQLmDF8JF92kLXXgYGcK9I6tC4n4CP
/iH/ZAAsHFI0Af6VaPEg6DL2GPF15ilz8vQE7BHTWMTKjG/IMAg1uKzrFWQg/pt+
5+n81fCQBQ1M0/LVm3qtPjaP4SNzaWTgjTGR6aSDT5D9yaauycIeZbIflwfTJrjz
hvVynnP4ELdnKLUhb5l5uznQDGzXD/An+qmOpod8xU0w3xzIIzC/cEhJGSM5c/ON
9SfWG0zmr3yNBrv+WiHasWAtVx9CDiJMEs0MLEYmyaPEtORwdKi7L/A5i40gii6b
tvE/4s3DuLkSvNSmhvJX0yUnLEICMuRj9e0RlDPXgcXSqxKdIq+3GsrJA/KikYdW
zEc5Bx+JT60gq08YkeHDn/AFksXCWE5vSsVAg+IqgtGc6CVoJp6h88By6yOax3i/
wpKuqHJX0oao9/8V1/EnSnizm1o8aQz9vb6rvbdTq8Ez++kb/Xtu6vGrg1oMG8+F
Et8e4ECgAd8W+e/B1kh2oP3xpya5endLb6Ta11XX2BkJFH5k+gv11qJi81FYG41M
7lu8DpUj2fR+Yve33G+k3k+bFAgmbKTK7byLE8Q43+m4j5h2ATPshjlGvfVq/yZh
39c+PwQqrjdHcMvQjrTDr+PViCi8Ghh810PxxBVPF8OlpWpkANY0eXTZmEXU07wZ
or7NwYywhV9yhWe8e744Tx9MYD9panVY4ZtQgmC3U1hojdw8mKsWZHWJV++U0Zey
Ih1OFe65y2Se5Iw3nCl+ldvZmVeOafT8SwPDocjRvmq22t2kuMYktctaGQ05/0Zb
fIjGG7CXZJ9W+d7E3DacBtXRuPXzUaZ84Wbm3eC9UQUkVWGPezfyzxxU3u6ypv11
323XAwxbzCoifHnMGR4XWqU8HMoT6l6scXGta0l5Wp2HjSQLqUNp2Z4GrmjmrXC7
k3tnHPSEXeu2fVikAREcaihUdtJf4F/m1+ZT+NnJM2fKepbgIesP+jO7SreqgDjz
CnTgrgD+x1z0S4XZYJ4p7U9yCADrxZVbZBn9oh5vvW4OprRAg86nJoT7VM1iLfN4
FVOnezqF1rdu9OtECoCdlSFA34bD8dXMJz93bL2RlbgMMurasLsClU8pBG5l8Ax6
ImMcR5vODKqO4NGmf7E6WyGBqdEs2GLTuNhWpSSE4MMS89hm/U8yo+bN3jG6Fnw5
GcdUEwyWlkc/srsaRrbpPgbmIVthPihEr+vUCDQGrRNv1wDdD6eVDvAgMGAcOYbt
Ai4W0dws+IP7cuUiO5va/z7F0czRiR2gTPrH8LfPa9ve58B7r/149+I48cFlARlF
u0qU2UjyHChJIuhtm5lrkF5HnegoZU7H9pRBPnmOOe0w6l2qPc/ofyFe/Jn00hla
wyLifI+6wiKkqy64/tqrTNdvSl/OQqSsaFuW+HLzHfs/yzFXJTi4VfCLpfWyAq/6
RFY24gxGl8xegn2Do0DabUjfTjXRnWvz1P4U3ISsjlOCtSQUmI03eSXd0YiEv7Fj
ql3zC1KqejRTFzm+8uYP3jf5eh6mQ59JkGdWpYIGlsbmOU/1EySHIY5PUMkWgC/P
CNZe5Sod1w0lIZjudJf0JtFolCZ8LkzPimYmhgQFiOKKzNBuTH9kdZGOFLSwRS+Z
vmlmUrBePMvB+l4gS3Tzskx+ZPzSp4y1M/1s1jspj6EgfM+RpKhML322bGxFJOEU
3iSKbgIPU4JwLjhkdGi/lzD6dvuSi+4GlzgsaR/flteZJL05Cah5XDkxFYcDIBpH
7ObqYt+8CgKjSIc6QdegPWEjA61maZTbC0FyEfOql+XG169WFgSQHE6JgZz00Jrc
XJF7+tZjH/Put5UBBZjW2RgNtgbsmyy/vuhppv2mYTh4RnJmI30cLEBhYfHYSPni
VHFkZiwcKhVJAkyS5kLxQ6kHnoLuQh6+4CSMSO9LZMDijazPRu545WWm0Zs79otJ
IWXbDu4jUIAn+BpuA1tkyxpeJrS9j0iC8iFx3s/oyk6PEmwMs3h1lW3ZsdTpKmd/
KDTghjwffCh215ofr7+onj7tBCrRrOWR+CjgFluGmu3TXIb48gyH01LLFgmm+Ped
qufWwhn7QMaYGgTRNOt4Fi78EpkAcfxWrf4OF8UJb0nZ7gu5+xGd2ZJbSGMu7/f4
NRIw5EbUWdR0Rjt+QQhou0tiq7oah4fCGTCLDScJNtH+iTDoGNKCY+i7bY6nsG8D
q47DnV6DN5tQMtFY4kdCcEG+mhL4XDnZ0dfLFtzi13Uo7hfXk1ALuSi66mScTHiu
QVRrbgoeV0TyS+GzC6R2VTWOoa+Fr0BYRr8m0299aSBicPcK8z1eQoNNBC6B3dGI
0uBy8IpLM01yZyrX1AmQbyV/teZHRc6Lt13/+wZaM0dXJzkk7PLEofFW1DCjN3n+
GV0ac4q6gwXix7rDUeSu4eX7LLbn8aQwbKLVOWcORe2WeftjFOsusDvbk2bgJSoL
NMGVLPU2TEq2DtX4b9AA6sOAbg1Ga29TpKMPduQDJ5ffouGUNW+kPIteyjC+HuUh
RzXUEN/d9wUEorY+NwFMkxkbvYVjLbStXSPs5Eex2eVz6Vt7OI/XeoobLOWs05pH
D6AWG18xngLectgI6Nqm6KXUWxOUGJMd3wdfHMRUgTJ2lGiFONsbT3iM79FJh36j
caZ9yuAbH60pn+p7pO3ifiFngxwSTqAGlq76nm15/3T0eEQjdabusT5ObX3DPr8M
R9T/ee0IV213jtCnwpEjH3qMzA98mi97BDcxGXy0VH8xeQ3TVcC45sYD86OEV8im
7L6Vd3pR2GGAs7dSQ9iR5MId/tuUOQrJBUxZ1Nim8UDGBbzWvAY6qADwY4Fp4xT8
RMYDY2MbPdJ91XeXzYCyYsNvJ2Bwy0uNsRUv//gbiG+5OkBwtMhvyA+Cw0+eEess
/ndjgFaXJWOgpmyXYz3PSqgM9mWboHFLIAy5X3NgyCQ6xAPu5piOGembwry55I4v
AQ+LvzTh2Mzqa1K3pDkZ7Wb2RIkeo2pzdtmaFntexoELU175vP9wwZmRVK81BkFR
DqrHCyAKG0tE+d11ZFPSVqvjRyQHquQfn8GivJaOrmPTWlk6hXZ0KlOX40Y1WCbT
B8B7Bc+o0Ql9BF+kYQlwyzKzM9Zyr3/K95zpdkzxmlxDUtlzgIT1KR/Pb4xDpV5U
EZzswpGFDB2nYN/BmHfgfkiWxa4x1elp33f/aMLkCSKQezonoJ/wBqUA1Y9WpLMV
zx7Ehp4SzFxIz0iWPHvb+3PX7Hzt/tWBTSu6BiEUmwJLwDjgCZ+ZH2dfPDV3mmoJ
8W1Li8WvA5ctS6N1bOk8eXWTX+4Rt6SHxXpl0/IlCifdr9kmvPaAqowWbviTNHup
75U46i0nrGEa2jvtgRyuBesqsbCLXPigPVhnDVMlPb15QDh2a3+2PUwRo+p5/62+
8VIHvJElcdgrjcCPyynIL/U+MuN1NXOBwGmwc1mI6gEnL5KQsyNRf7DdIrsN5hsB
USr86A2gPm8uTmNDvIYT7PQHGYOBhc2JzYKvHKNuNHGRuLKmsl6zsHGXF0gK9JPw
BGWBT875azX2ubPbP6KuTcHdrST+lEHDAnPOHh2dg2brhZqfi8Hn+WZTjFBjXy0t
pq29e4t8voWp33GIx9gDUNANOZEF/Y5L1LaW0Id6ZvU3gs4F7Uf7UdYPPtftdtpo
VTQj8CuDVk1/VsRHhayEMQiT1iQhPnjGnYIOzFI0L9u2mXSOyuvlphTZ8e0uk9wF
yd/Vd+H85xvNVEy6Bzk4nE+ipw7vlmCbSF1KV/T/BmqgCMNeGqYpoYGRK9tLj+t7
9T5xVpzLeG6Yosz3FtbexBiuv/1gSw6Y6a3SO+ZD63egbuCJzBC1TF2dvNg6ovPL
wUSsMSBi2jt4VoMFlKqUI6iZHgxhZlNvsFwgSnBGtAgi18Stky+7aKvM2Fw6zqxv
QGOl/p4+fRN6ubwl+tp2x4/da3uu1Mk/hFv91WpJi0He7fCePsou4v+JvEPw1o62
ny5HBRzGQ0u7sJnnGb9FWBUM/2im9WGBUcagx5/64RotWbUB7516Xncf20eywln4
+4RaKaUk1JylGf+f3/2nadn5RfQOhAAD3fMp1IfkhRGwmSxSXQN2FteqJLJ9F4ZZ
yaO3wARaTXkJ7W4cP/a8zrnOItJ+Lkw063OnM4hVIwWi73yJYMqo3d/l1/p8rMni
XF+deVPAkWKtCYZTlbuZdg7l4JjJLsvReCRubvjyhg0PDrQ7GhHNOBnTn7SDFpOt
Mwj7lcb0Lq3JEmrUOM9z1WKpSoOMffpCVAFdsD0+6N0gvfNVwuVSsCfoVqnjq7MS
DUxfP3DeOhJ+9FZgM2BzaCdotKUFHQYikQ882+CH1yJjrP5CEKfLQUSerVRW1Uon
xq1c/711fovWtutm50Lm8sXLbuRscMwjHYjuUGv4ahyzE1OPvLsufgB+m3fMOFnR
5ggbH5+QBOuVF22j7DDMD7LzgFxM+oSaEUImhfpf1uAyS64t75pDJ/AgaKCSkfI5
jbbHC+qADwAZZjGb0bfxm44+CeZFRbTOOxUL3PIpJhmJRxBy8B2xMTreKhwXfTUM
9DNUIpUoF5qre1gfA/aDY3LqEu6uQ7CWYPwKP3AVZ/9etUTZfEJqSiY9y5K6uHZ2
uqCYaXDJebocZy70RAqCXC8VkYRG4LyZDwqLHJBjUOZjrChKcTbWOcSqvwidejqb
i94O7w4qD+eq4ikPABRdH6fWt1PdLbnKmXkmjNMNQMwqGH4DQ8VXxfPQCAu0k63J
f+64e7gEjq11NRr+J4xY4MxCb+mzyVboDpTVdxUtj85IoMnLVL+uxVXvuXhPwBFf
cdEE7A9wHDP0qoWNjliyt+ErzVCHuxozLeCOYy5iTg2kar+7Dy4g9/88EfZ0eJU2
z7TizDG2C19oUs2JG5XGnyPKfhXfsLLgxWmUm5yn9IBgDqZTDlgsmDqM+4RakVeW
cIDriG93CRIq1iYA0kQF5/OqSyeNFV6uEJHdWFs7KpvLyH+o4Re76Me7Xmm17kT+
D8viGFWrgZUj8V7/igYrCCgMrHqvuJwK9zSwpiFguN9M519WsfxBwHJoF5zypqrm
bQIeIZ4h0o2d1eOhLWoKpbOXqASSzDPNcipncFZ8bG5r+ftLbPvHzMkc3xmTuG3R
BpuDR3dfh56Em2QeMOhG1mtPNYDd9luAGNNZYwPZdXl7kD1pVKCCL+K2WYha2fgt
TiSZ6CTJHnnH6xXmZu6KvAvYaRhOhtuRgORVqbIR0Tg0ezb5fbLgjYKH4OeCJAju
hQZGhy0lxjBDeHRj5TS94Ecq2rVoIBmo3uD4Z+258o0lA4+YKNCafd2ESkSVj+c8
xplkidg6OfhkFwkoh36+6lkDg+B2ViVU066B0C3+qq1AFV0/wx73TxWTQLvW6MZV
8crbRDunekWY0LMP13H+tIbPfFrC1GZnsKC7XzKEpcx2BDhxSfsWMBWCEVya/v4T
RkTaV4SY6PsfqnWls6qNZG7d3od1kdji5zGdVkUW1YSauJi9hL3JDERsjnYYBlNY
A/tp/XxeeDzhL07wlZsXm3TjdLASIl31QbGieF06skF7dOcO1QrQi+5XVw9jpVry
YMu59MkPBpF+sbUUsCHgw4Sb51NL8byXXRctCV+Bsn84uhCOAvEkeCQGBQGU24Ik
GHh2BX2p1RaVOBOmNzpptsWRc0WVEef8Mpyhj8E2qdDd84CtZnsIGHL5uE1PaKEe
d04EI32RxBoYy/RK/fejJu3jeXGJgDjsFxsX604m8KC3oPUnoyLFKZisHHI+l+jS
IdZsRvCRZx1F+k1Npd+EvJinxG4jhM9lV4GROExWxQQDNoJjc7uhOYHMxLgS6rhc
bVQrAsFegwCGmacq8+49tQjvTIpgaUQjctawekA6lwP2RMozpsh+/iW9VsejB48f
sio8vxmf+yXjP/yTtewFHDNUqiIDavu9I2nQ4mT7oPHMPlek+YgqceqDvVInO3M/
X15c4m9gOHzdTFIP0G8MJyEotUX2waxqDxa0Yg7OayAbuHUS8g0pYpjzATxoraQP
GP2zb2LjND938zyXvl/ebJNRgBXRP7PEcQqFaFJn2JkfeLYqiNLFbT2AKd9v27fv
JAwGe1TnI1hBVBdwPXA3m4wqzvVwEbke7oTGtnxQKdISP4+1UKohFjlY++498zgd
i7RxFhMHttuv7mo/HOJg8ysKBS7H1nAjI+UsZD+nJmsrCzEykdfS55Np4W4pupOD
mxHj9OZj/bec58YGoXYBL1vQw4ur3ZK2FvImLip0rPzV7EB4QCDxVkK873Yn34MP
9c+UYH+Y2WyOXeV8H7iHgIETmzIFjJrnWPZwtAG0ID968kC+Azhp/EPZgZ0N/9SV
qonxEVL6rz9xl7pyGZhi7j/aNBv12dQy/QhuyNkXIyiSx4oDLVQ4H6o/yUokCXxR
luWamth2T4XrFszi6yWJrJ/eL99TV2q2865ytIRtXU+2pxRZWbZ/9zGlkLQAvqjv
j176QdilGF7SCCvNDqh1B4ATYGjewdbjCnq+kvr6iqqGaCh4cSnGF3yUxgf5GuLj
v/Vlq0S6ct3sgP21UlYb2A7v4Cas1+Gp0kW7Wo0EGR52n2cxfWgonOV0ICPVG6K1
fH7GnPpgCnJO8k6OMFoA69QBCu/DIkvWJyl9j6/BI76A3sIMn9Vxdnud1VnhWvZW
2EsyUytEcQEuvTpLSummt2XHGghpzLZJyR5cqo+C2JFHgJ8NAVBinRdfqKDDaUYK
PWHFliRTZHKZ/hrhNwarwXfbwrYawXCFh9RJzKxtRDgSoSoZuORDZkfchVANkAJ3
d4Un0BsUYnhsjEpGI5Sx479+k+PXMNnc4VoQeAsf7UgzwND+ZTvadrB8THnh/GvZ
a60JSN1dfHZOjWxjMiCYvhj/yXt2CM2VMhmpkzKdwr4wJ1/HVHzLLd4F1+aPyc70
a0NL0M4MJDP1in4OzVBI9ZnWWjiDzFE+UUHCpXFfn2VMKdLI4F14It3DQbH2MnEn
1UnfiGSlbd2H+0+2j/aRMndkhjsAF8mhvCLU2Kka30Clp0QbhLSl4AHiKCU+PTF3
+jl7yU/oNJ9oQBdmCV81+lIkeQdRCNbxlmon02aPJMsZl0vSyiEvF2VUw+/0QRnP
RzSVfK0FzAaQ/djFZhnpbwkyxEz/wRmxApmzhlfEYi7hmRCaAAMD6kOxhceQaCQt
pv08rND3QNCEUnOz/yxwTzbGRAhVW1pjjkcfnwfP2rtUrRFQHveQXopDx2jCWY5D
2tMrC3KXi8BAvcET8+ax0SzG9c3HBA/k86JVxS7d4HAWme8mFpIyZwI3VXzvD9mA
kPMj3ZelOrJ7sGsxwkeRcVUr75ZlUS6KFlVfM7CY4hQExM3f9E1HXSfTfXyW+4Qn
X1ZZRqvZhnIHfti2qZsC66s+7mJ+VrB7Mre8hojpxmgUtjERS0RsApdnng3Kj23E
nUTUR5LqRZv54FQm73gcDd2/efNTW4B7vgoORjH9IT/bSf7GjEbWDHV/1O6aO1gd
FlI0tMd0/GsLGVXmAHymTKLx0SB1+zctr0PJrqp1Cbm+zAEmwH4UWvyDgbBndAJf
yFVxFtzUmQSj+dGsRfxpuF89hVKorijhbsvaucbb0Wg3yquZjQ2qVgK6tTxbWR8z
IWK6IdlRo+uOWKhofd36aVPvO6mt9z7yRRpNyuGMeHXbocfGyZ9jb9cxGPXgbDeZ
50mhSEW6Y9BhtQvOIReWt5c3zJO2IGn2pLphKUljC5+pKcexHX6PovNpyMHBjc89
ThgQsuWUTH2cH0AS3gC8/I1Lh5krmHhZUoGiqjB0Vdic7JLK37/qr/mHwCSTZUdH
7jvhc3EUBNQnns4ONNhgohAWdXiCkCz8aG2sY8VW6nGW85CGyUYbACsesT+oFuxw
eWfNcn+0EX6jphN8WHNRK3Ujw4jbImEAtvI09P6+OBNu1zMXlTA8+xVcV+IO5pWQ
Yov5NJ2kMaBcLZKFeTe7iwVNNrKdCEg02zsRSmhEmp1+VkP1+/+OGxAFiyMvQ708
S2eIxC6Y9Jx1mvwJnbdgl5foQW6RSjpQhEISwo1cG1HtTiGAg+ckgAv/2IDecqEm
rSjVh9r8HZImAZeOMM5svpxCvO5Vmt4rHk7ECaZos8hD5wD1PTf2OHjwjaPR7JER
a6+ztpWrMLl6xiug1jF5g6GaLnLEhV8WmLlpKksEiZ6pG1hgdwvSV50KhBfPK3SO
UU4AW1i1MsCnjao/naSQTf1tImVyOsvunxhGzgIUyQgIxfFqEvDxtInnB4+BB+lJ
cGRrL0QyJIW1i1xeEivVMTHLNbhFUQFuVIEHFRCoit8Y+zCG5If3NgwX9FMmlGTG
bWRP8BYKY68DUmmD5GEe5oWonRXvZYVBw+id6KnkyYpVb+fk86RTwb6CY9hFNI/W
MDlrVFk8FyI9oLDFgkxEA2SRwaofo2DDrshMNSGz4SG6OIR0bF6CM7Jm1VYcPo1z
sRaUu4XBgam3bc3RwD8GL9hhidJBwYTTt+0ySsSZ+rPmxPg+JwgYh+JzqgkqLXov
13oNYsp54nxV3EJ8nWJyFvrCYXqsBV0cw3rI7jnqLlTXmA8wCKhBJNI5yyJ+GSk9
nDkOT3L8tkvY7AxT2OSk4Hz8Jieh+XItkHbOXxfHJBs6zLPHg967lWIQDX0gHMbi
HXwBy6QsPTguP6SdWzobFqpylxUjDHC/CGnxMsT5PYD2XswX4bXB8zenwjdIBuyv
yOirR4GJ45brav6P8xfcPZ7lSJm3ALOzhntjXcnIdcwxH6qDmYY0n+mx1WPt9jPU
JcwL+a282rok20JCMcYWrLzgpw5Dk+i+8ceXHQnffnfqKz5zDu47sCEtL6mZAevd
vlo0v2VsK9kDM8Tt6PtWmt77THKQ1VPJYZXLP755JuVkbiznsHFCFVXkFWSPT5zH
YlzKvWrAcclKyYBlBH1qNMtA/uCKaEtNdDssYntPe+GmCVNLfyFDQwGJ33i/N15n
olr0Vyi7wP37r71bAuT1SSr/tptGwNvraz/DioaSnyWcZmXSc1B+nhTN/VXUL3J0
wXdBa8hwQTDlLHihiGjBYF6iepg7HD2huEuy//hhpDrXqrYoNbWuVRxOEF4EM4Bc
geFhgm0iRrO/8WbVdf0mwGOx0DkTuau/RWMu/RCqpYShFKvoU1ZHevXWqwuFnvRW
oFGnX+NAbH7cLn7+d1FrLfF8xKPd7G1WCRzpn7frSs+eZDEnFt0kcENTA2Lyl8oz
lwSoRYvGbFvikPQT11G94098hc0M9RfzTXItHyrUsEVbJOnlBi2EKuSncIZgR3VE
ahQ/2D7sGOxF5UYAR0scvSiYCBRLIdpTOd90KAGj4hlu2QXMbClE2ICeFLBUWrCm
i0kuJSR5sKeyqM5LORvnxQTkzUTVnmFVFO79PjYYTt7htVeOASSPyRbhIanEKiq/
tbc/3dQfacTQDoiaFsxvxa+rJg/9Aeqf4PkFk979ojNn9JEZBCJiwykvJorIspWL
TQV6XaCHGuDWQeKy6a3eeX7ximzDoodN/w6kDMsei1bdvAun3/5xz/yBf3KwW9D2
qJpMnpNfuTwFNT2rEAV7wQiHZ9Vxg2DRuJfTUkE2eDcuhuoRwflxlD+YtEUG3vST
Grjc43XAIJaaHW/P4F64guhi+l1cO5cdBYvFoy9oVNbezuHmp78aNRkUdR4VYalW
pUpMXOxI2CxjGy8fRMiQec83Zfu1xdBhnoR6etkH7coR5NqpESosx383Lj3Cs3/3
hF+SaZFCpJIQqJY+tLrdbMclo6dYMgc9LX3TGb8WiWFM98YNhrYqd+VyHDGtWr68
kY4xRIIGPN6vIsvcbqAKtPLsdNPMX8VMhM5C9WhHTemqWzRd+m01rFcCwZV2H9rb
iQlpf1v3SOeeV5vB6tp7QBw3S8hZ/CCUxzkt5kdxmyUIy0p6PsnX0Uc5wHOV6WIl
xUXzOM6tpw9DUiBAwexDsu/zhDkqGhlD1CBw+91Rti5brKly4tylOQXqsBoV/uTg
NKRLFl6Bliw66mQtPqkS4vljiy+QrsicAZy1lgCYgqfzLgAPdAVO0VNpgmM3MshU
DTK19xbgNRUVsnk/tMItdPCeWRsbbiFb8xLsx5erBlfPKh6nnYFM5QNttqMNPjAa
JZpRgPSOwOHIXMVwlsXnNhIyS8Vzg5xi16ITRq+dD1AAA57kv111sbECV4IIWHDF
IMIZb8iXeU5mGV+jLv1Ui0tiPhCMG1Gfz11H0Wrsa+mnvoAc+EwTo2+sbR41ImJX
frg4PJT3HzFAK56TXQuvomYD/4Yb47zUzOT2bT6gHyzaNUmR2aKLSpZJOMwsv7TS
aMyHeH02zf7q3Ojs346Gc+vybiDBOoQqTtO0HD5GJm/0nC8caLvPcKvIIEpIxSqN
NAq0R246avmxQnHH7cy3dPitj7MHt3SinbnhID/XMf2FaDQAf4FVw0C79nH08mTU
IcOQunkwHfnYjKivIggJGVILb2B9RPdVHiTvvH38YzyOiQv6vwWwDNDY8OleCxfd
YOM22KVhiLjKL5L0XXvJuaiEpZ2n2cWAgrGsH+6ytQy+6vESPOsa+8pRzFU9FVCf
xFaZvHtsWHiSIDaWA9KRS0DYZ3M0F0l/vwUiVKvnGJU9z5fWDHckf5K2PLxctfkV
soVZnhmhTn7BZ1cdC2AtDQdaz6vl+pKlEOrUYEfqxAXcSbz1tBNyhPdHy0K/Pob6
u4Ai8k0OpjoxLjKiyEO4IPgNrEbnmo2pxQyt5XukJ/JwNLjbp17EDXdQDeku1wsc
D3u+BZ8b9+ZENNFg8t+tKGpALtIDuhaCWD1YUNoRVVGcuDafMea8gviSeNVUeRln
lyH2NeyPdBwPfWC2RsjSxQdEhoUcZMVz7E0Y52is7iYNv1CfH/MPaK2GJi5iO8gw
+CifHpB4xhiFYtQQeWw+r92S2ebnZVBW5ecCl2F2DGZxPHEsSz7PbvmxP0BX0x9b
fPoSAAeRZGV5+1FOK64Ph18eosnQkk8Hch1rsdAzT5AlVwICfLCkxb+PobsC7Qfe
zWuOmt5BVKfDG4XmqP/33Hec1CyLSjHsOAaN7KMIXvsBFe5dQnZZF6NDOwiwoFHc
mLoOkrcbsKygAvc/QMRJNqzwR5l5CZZ6kNxXmI2uemkXLXYrZODTSCTuLIgzJQVF
ZSHEtWCrCBY4xQG9cOvinTODHhmVag/qQ7pgpV+KTmKkckWTdLyY8uWn3sVhWHIh
0QHqtpmcig79geK/BAH5QDlBv1N52KpxcvjOcX585TBlxgHfo5PjSeNE2Bu7DWyP
H6kZPZbcwca5cBgPe6cwU2TjW81mJS71rb/Ht90FIktmiw1ESdAXAuAKkcLcCisC
F3JBtBM1hHx2Yeo95/uMMF483dbYXjiz6R12A64D4e/8hlcIUvLCzf6BjGzgmi9o
/LwLdFvce5SVH9CTkriObH/Tt22+RXzTxZeJpKDJEeEzTkN4BBNtl2/Qrsxblcg0
zjc8AFrFzLUf7To9v/RuGkGzLJdKzfqJkVU+LLdr+/8D6gTQ+eeuWeHe2EXVUVNS
pUF1tHKsEL28bN+Q2UXTIDlj6RCv0CaR8Z87TOa4fEr6E4n3wsmrSjpbawCzGs2t
ooUinGgo7LGWfjZA+B3lTCrIbzCM4iz7w9vp/VmXoXcKQd/t5R0YZWNBPi7p1D33
Lv/ZLQXCr1buv2T4AsDSDztZmJ7tVXLq5UEK59KgbTI2hJc5sQIqWiuYghis1/cv
RgDJjFRMvSY9jNFtOqQBZa4HVqMvNB9qtyHAxysUbGSI5DWhC4WYjh8oj+1Wgg3X
GGOdDB5slsxgFUE3QgNoFLI53Nf6K60KenTvZ4mbkQg+5KLPmXOKaoVbJw5bxfDP
d4Pmu3Kqq7RjqtSUAShdTYyFEreR02HEY2vMLYugeBjoJeGHj2dVCIeptHK7uB4v
biTGV4D+mbbnkpniEuVKXBxHIdjVCubJ6iVFdfcPNeR3dfhNB3O7XC0Ds7Ezj9Cl
rX7FLufG9SLM6BzMebUpD7Q+54dJEJExbvw19CJmSd+Ecbl8G7PojKzkeqeA7wTu
F05RX6+sNJv5imO3WyKNj5800xftCRam9eq4kbKqaXMLgoB5SllMmPyV+ScKVId5
8O4CTZcXm+EjOo50qFDgzRadrIFpFZ5LF6T1Z+zH8uBIre979oxydpuyIDBCF7Ht
3bnUYCYgGcNo1TN+u2WvV1twBL7dql1XOmTP4J+AFkV9+3jF24ztr3Iy4Zz+5niS
p0ihc0ol4O8U3AHMm2DHPm1fFNaYffMEa9Ru/bMqqZV2YBNG29XmQQp6ypSQ1pzl
k8GxZpVdw8OLT3lgK1RF0FoXMxyH07G4Rsb64O2mCtJoepj2NNs1RMaZRmEYk9Q6
SVwvlYlJOnUHH9PAINOicSgJ/6qKaQU5YtV+rddviJhgrJGSVaBnFnrSicDslpBt
7pK49PUhDq3HSkri9xPRSUdZgLVQ20Y1XlEgH2QL3bVcuvq3fQ2pqkv7joyJK+1A
uFF4IRTTdTEw3PGBqzyzYV9YnvchDnBHxZ72z7OABbVZZToCXSdCLpMJRyisrSz6
MFRgESgGKVNzq+ClkJ53XXCtxhpEa5+snwhXZttW3Mo54ugYDNR3O18crjn+R7k+
H2nDeOf6EWcQ3YHVoVn39oHWCeSojljlgtShejViWPJGIKMRd2+5/Nlr9wTmYAIm
cf3TBSlqdk9woBKvUBbKPvoRqnahnhEYuk9ZpGQM6Dk4gJXNAS81TJN68A8xa1C1
aS3nmI4LYg11dgtPNwfYIGQmKZoFghSgxKfDQ3Tq5KiCaT+7dBmFCO/4nilYfIq3
QK4Brzir/1tSGhrpOLcOCskAq/o8nGCcQpVM7s7KCeQHX1pufXrPBbahD7XZXMxK
jkuvyVf++OmEc4mK3mnTwo8FPDBtkYrySPR8fwCym+ssOEyUxTdYEOxWjocvOYaj
C3KAtIHxUS0W4fxcXSIW4JdIqVZtwSqpYmeYvzEYBn3Pyd9YgacynrTPLDwfgDHP
uc71FYF2fzJDw7dYcuc55wPfeYuWvMglyrW6M8DQ1Osb7aare/OL9OoRs/biJMUk
HX2EV6rG47hHcFn5QDjL095cG4NfM8drw8/+mYSQIP3CkyYiCIP77IZ1PWqMFs5h
rw8CLGwODRR7013gHqlCIThBLrDrrFwQXnsSr/X2NPKwygRbX8KvwLKBfCcxtX9u
OHWg71a0TQ/dbBZYiuhH6Df51il9zJRKrIDF6tZb0+lbfjl1SPotoUKJaJ6XF++K
ry9ZzwVWUOVgDn5T/DudRc91jk18OttQWBAKuGgjqylHi0E4UZStD+ejxy+sFXXV
f+/5Z75k5WOGjYGvxqFIUG9kKAXLniiMKNSxbtbhKVi/jXA6d3qAouVEbvuc+xW+
2wuaRTpjkQyygDTPae5ZS9sL5SPc133jPYQjQHpF8xnSu9KMzrQOlykZYPLAxSXa
amBhfqEtppsd3lkloY6JC10khJ0rh6fMvM1A+ZFf1jR2IllCTfe/dxpv9XDfyNpC
am6RsA2D5od7jjaL1bkxkqwnZSRx4Vv3HXDTBxj555Xcg8+cZ4CXExixy8ucOw4H
60Huc22tdyObTDDC9Lhi5naiePvrs/O1ZBN43Io2QuvJka5dwjgklMR4OQ2xmHhu
/p5W0tZqDA0kp2ytjcMTyzllegKDhzHWZSpfR1Va2Yi2Fye0tYXZKpp8epxrUiJP
WsPNTAYFPszwU3MIStQGd5VF/r6FZOUTcvctprPsxerFgkkzn5PARN9H1hs+ABA6
4pM8oY+EMhD8CRKX9QU9ApmccSufnvN1/Doc2F/TAykvPd5P36albgWyvV4/nPBJ
AQYHllG+HROl5UBjfAAlZcJMtoRuuyBI+QgntNWMLnf4eO1YtJsbgAFQBJYTunjt
/o+HNFlYdtPdwbHF3cQROWUtIm31hINseYAyAfUQyYGVmsqM3VPbjUCUIQab36cs
meWeetKnl4HeXi37wNMKIY6UcndRN2T5dfmWweWBWm6429Uo4aLP/Ea6NS97KIXf
F0VyCyeysPFQ7BEQBwxD8CHo3nV3TQc8CqNuzucW2H3xGkUMMrZ4pqHr3mx+nnT4
wY7QYaUj8m9+MqaDGVjkF5G+EEtxU5HxZ1hRw1zTWcj/E+597fWQB/y8hOsOuegn
Tb2LFlfytD2N7P1/5xza4jg1Vb/Q1D9IcsSXWJjI5Gkv0l5fZygPhvZ//G32J8B5
Adjsq35v13G2OZGdgC1LpcNiZ/Q4P9QLKxzQuITqYivMQ+DVGJwFIbmbU4II9TAx
+XbkLFlD9EtBU5i94dzPD3sUFituLV544sOa/BXZz+dTPhofPVDvjxGDwvzr5mEh
sLcnlKPOsUjUOPswxm89RiEmWxdnz7/XmOAiJPDSsObrkHXjw7zWMka2oeZW++DI
pan8n65EiScwJm8KQ5IcGHOzj2QRkMqngfccWtAU2IkYnmnJSZ326Jp7IQmhZUlJ
DLAfS11qorQot+JC+rbN6S8/BYEathrT2XLRLb73lX7G2od/q7oRRA8nnAhdsDV5
4PX3wDCLzXiOp2vVTEbFe6ep+D6G7brwzEsmicQxcs/VX9R3K6SlVfiiH6fIuiHk
VP4wg4fzgNbx3cH8cRfljkV/WvoO4Likpei2HFraaSKO9cIKL7cTXbomGdcILgkM
KE/bpnkQpbh4EAWdLuQ6sZGwhCaHj1LWdGa/dJTJiZTUbv8Tq57k/bv/ATPe6/o7
/8BAZvK0r75cRV4rgiLCdnUwx1/BDgH38XSYiLmnd3SXD0tXucZDYGVxAC2R8iMN
mpISOq0ECHEUsy/v5R3iHbhjmNcpoqzw3LHx6PHRVqHl6lf7GJu5wBJJ19WKYpkZ
GwOWF/sfbmtyw4QOdXp67kITmoNG2RWsLpM3f/wlokUkKlHFHK2g86hrkpUUrrTy
u3fGd8IdtAcu1KUXQsZYpBA3JF1CMeZt3ebWghuijtAppMtSiG+U1g+MMgiqoZ0t
YM/LNN6SBOE3Mr0jEFUg+LTqOKxksw1xOKe8CImHWNiaBY7HwEm93ZDGsIqnzywe
IL/z448Cd0MtbIwIa0V2M6yu71ijhLpu011QwRcKVcyxsiybea8QnGPLOBEEqrIv
XeofKUEFYGv6swZriOuDKyYEWfTQhc0FzTWQADIzXcR50XOCvSmY5HdIMigxE0wy
KkQ8hQpVmBYVzgpyUW6BqogjVZnIxuD1uVfbIUyBVyMnvUD1xBFARLSKAnxTAuhb
9sXLXnL7lSkLjDrrsP8xTx9x8/O35Uhhk12+QdMCZrBSLDyREZPH0vJzP0Z/LkSF
kd04vSH5O5+74MZoJIYq5eN2/69agKe1kR60jSRUEWUzO8lupLLFxkAmv2g3RAJx
WclB/VgLTVkPEQwGvf2IJo06xQWawCriN02wc8JBf4q3jOMfEzb9utBRHCUPml4X
rie/JAQn/iGf24lFBC+qzEAOIjEODZED8B8yI3zyOwIXhpnxwj+UW5AeZDS6Bv0R
tqH4rklWHboQCWKFApLg42RRmYvFAdIUjQ6kN+iRi81ilw9CEgaz3xsQ0SpsiFxJ
Kgo0LIwSgsZRhYjn3gtKQNjgcznCuziWQgDgOPiD3PxI3VYY+ZJzUkISofHGIxlA
DsZs1mJHfkqtT+f38e+53dk3+AhZI4zK2M0n9JZ7lTW+NkqExKQ+sTfBA7CIP+Fc
+TBYKIWrdqj9idrmoXPK/zBgXjEa4/MBbUlQMvAJ1z4RYXi8Ckm1kUEBR2OkZ8Vz
6H99zl43deTVupOxy80J/nwNIjPploKHgL4gvJ0g5l1PFHd4b97Zqt5iB/XzkJb8
cK+Apv7cukKL+ETGlPwLPZuwgvXf84ZDpASlgKFtgnlq4PiGspDBY0IAG9cZH4P4
vhyuVAgPTmE7o8feK4X8pg5YdFmc3WFpspqGdR3BcKYv4fLq1HkcjnNVvaydwHXr
4vt84cUoj4zTF2ccuef8bYc+u1v9VCXc1mK8sCeYt7FJenWiBK7v2yPhMx17pCbE
13HvyFie6Ge/zKVsc4Dtye4QA3DkNcNPEfS93nMmMZNyeCoRmoZOHLpVI4lbAIUF
p9L5u46t1bVv+UD5gMwwKzQleq7h21TYwC5vKRAHRhFPJm5torfsnO9QyJHuFXDp
IUhxpGilcIuCJlL+GqJh1mc/F8JVu+UW6ymaKfFcobQE/Zlsjzu1/VtLE10DZUai
ukhYRvcZgE+aKTxd1aeeUkGaV9ekvmXM6wcUQQV/MJouqqPqQSnrMFNpXPpsFnOU
Y/fx69up6uOX+sxVLjnRxNPolymxQNuDT2bXMhSJN7kE7tZjYWfmcFHLe7iAorIG
GXrKHt3LeVGSAM/vfDhHCbtzSefTqI437jVOpu6BtelWCcQYdI3MP71RVxpwcC8T
ArkMYBZrYiTQZKpmF5fbJtpf0NR7b16tPCQChE/i5BZeZMG9vpq9+SUSFp3+WUum
xUr8J1qe16MIsmr5wCVS9E1sNQYEbA4/S3n/HqNyMTR2eYlEvP2epzZH1LUXlknD
PJc7GyB83w6N4+pV5/f3IORPMGovji62zDHiLVulF4Lc0Bou8OrMXCxMIbfawwxw
zoJfYdkf6lEFo09QUuPsvqtJrE4faqvYfIKh9lGJAQTTWV7ZGBDx5GuYWd5DzK4i
FPRGZl3tpjPAP/krzV6ulhblLBiNRvYpWi3sfE0698QdFG3qEy9vIq+xNfRfvH5d
E+Czu/YwgYPsPhyd/tOTkvGoehib0njwxSz4yW8K7mstSItBZqURcUcSAKudLrbr
SjHki0d2L7DEmtoNAFoIqy8acaVIO38KjRGZs9x8R+ED6XYggqqdfJ4lROOHtFa/
qg4yG5Du6kCuZCrBF2yCsleqJmT8dKHLbqjjSq6T5cTlhRDi6WTLEy/+YYSKtSG5
KK7nP/kWHOAQlXgsnWxOw1YMXDZotZ4AtitHEQnwGw/8reHAIMYS2V9bJ8FHEAk4
d4Z+TsmecTJ39Ebp/yaRuslIT6zVi3QxAfHAdbVhWS9PAX7m0M8vDkwz8VVm9Ygl
YCJQ9nwfEFrpEnZiAOPOLTuj1Ou/mMyXXThBeBokk95s9FZBfLiOA4xZjDVPK/zT
yDwEhECSVbVSjLLFBGiOTz9UMd5/x+UdUeMc5vqJgOzpIEtMRfXE+O45axeUw83D
IWp6PEw/afHH9QPZh9/5tuXFCwfB8AXJA5paYYN+UMhZZFNYHN3wXf2VZ/3WcC6M
e/OlS7tzN6UYUVnC18mVJYK9JyX0c3dyyRoKQdPxUp5zKmy8o4nE/tTgWYx0TeDB
85B4HHch8eHqEQwvg/Y77J4Is/mdaesk3EWqbAMluCb9OHOC3k/8JU7KswQvoxC6
4tdv/HWXGHzi7pbiVaqwLbs0+XjbbAyqWSQgQNEE1KoLqcbtAGvbrs8/JazRaGyh
X0g7egUca5uS21JIhU26GWv/I0TP+/87w76gYLFoXV0WDiHRBL+LgyuyLiIRzw4V
IPbFV3EcsqJPGvkAXYW2TlsLZLIHjdVyTRclr8SbWY0aL+wM6rsXKL1S6PavK0e4
wXjqxo14+tobgw+M0SR5hCJdkLWfy3tYDyxZ3At9rmPEHvYRn/f0QzIM2FN7ah4Z
KOKcGRcWnGaH0J9NY01X0vHAm21Jeq7RTPkEoLea+P6ftGjSkv4tAkrPo9136TjS
/pBzHv6PVTSeeypk28DLlc0JSqebRZM3iszH+RSumS3GJtZvE+l25OVryX/1cZda
CFH/xkk17OvY6y6cy8mnKeOMxBeG0d4tOyO9+DbBvlEI3ONPR3DRwA/pzuQ3QDsM
SsmFJ4LN30B/wFOnXskqn7iRfk/aMwb5+K6brIm3N/0ItQH7vMDBoAXNXytBEk8/
YfaNm61I1PRybtrw5noDF6fu+2N7/gj0rWa+zSMaH9BRD/BXP8R30ldACAxgvOGr
jalnxdl87N83sKZ3gSCB9xqdFI7bzua3NpzDTwhaWVJfgnZEBHQv9xSu900jL1P9
Ak4PczR39ybj3Z/ExBt42uU6HZWP+KahMSy3Sqt2vZ141AAYpVnQE5gK64SRQ30S
/bkCkUwvwli3d4WbYxySYj9Mht5PEANwaWnFPqY2URtAOQBzsW03lcLg7xcC48Ja
B0DYEhq92n1MX1XcW1AL5+HpAIWWkVq+1ksO5hvARuQht8++PjppbDD+gIYyJGmy
ag5OPzNbDU2mI1J+956VcQeXwFoZj9iLdj1fD5R4b5Zsjst355XhF4eOExsZ9l+Z
bNAAvvD3FtJZacNCrJWbW9SIEmWE3xjApdnNa3Cq4fsPVMljFQelIy8kqWpcteQD
S1h6squr46/1SaJy7HHz2E358YaXXwpOKQD/pCIgB6WHnvNj42HJsbTEHYbu9UK7
iSsxr1bx9QcvIhK5QvCgfiDiZG9Yw+LjvCUw472aVKWZfVb3b32q76N8O1BnWVSq
6pzwVUe1IXhgff6pHyWpK5fNYOGw9dbjR4kQurYpYB87emXYAFCBwWilCHUioypK
32SWlwVSXy8sBrCc3UOaIVSC4bcfY7yJfCEttnvhRcICy3EKe1eMJSh0p/JoPYoz
+BRpMn/wmPZ26S14qSozeY5/BTv4QZ0vkW73lClbKmCnl8fWsKRBKLnKV8gFC/Bh
lMgsV4whnBlra1MDIfDsWF3bPgjMFzhsv+asfcjJ1aC0H6KK1Vp2pqFwiEY1maXs
kKJZnvzFXSuRoAAzRZa6b86JmwigLpn946psSpXrYgC9EV5x/9SNfyxdrUOdZmRZ
cdBJl4I0QaYvT6vWQObMYHvF00QDZkMNFVMr9qyPoTf7B3acryyyfQq0AZOUAJi1
uERrA/MpNng7m6l+qrALbYPpSkzuFVsS7Ys6q6nIMWn/KG2hT8QNaszCUEsFiCEj
e90xQFPu41iFKIoQCFOzhX8ajcG4PQNFW5q4BF2RIWF2yDAfykfT+KB+pBzbBPa5
r/DpHkfoMqScfvC87LJLk2h9LyFnWq60hoQAg0ikVo2v9LbCxS3Iq6i6bxweDHnp
3SDT0nYlf9X9H+8vn/2FH/JE34IlHspmndbjI6NyN/qakJjjKvBJILyp8dVI8to7
4hoEEhxllCQ0SdG0ZeRkzEruKyW4ip3cLQuAQb9tpZHCYbx/7Bce2CUcmsruX8eF
oNUlI7dUQCB3/HthG2/aKbe0BGlsPWdt5wnB+DuHEBSWjsCMSWtGMAKiYKkJD4Rz
Wx3gRo274cbz+VE0Yifez+Mi6397Por1DLRyM8i3XW2STy/2ZshxttPA5hcJwItp
0yx+4BaKHOtlNfbdnwgJKvxfnsf3Ug3t8yELVL1mM+WMvFMDPChShra22UDlPwEg
SqiaEj1sC/rQXITAWj4txPdDviOLyaeHtGMaAQM6ja0bngYKKCm5PwwX/T02epgC
JHLtxsjOTr8H/wZj0zW5TdaVQ6Wg5qZyEHzvPawG3Zvd6asKVHp1d06X2YKlC9sC
mxGkNrU0K7A2kdjcxihbPaRECKHVF9iSbjoEOtRvW1Rv2kkb48zlu8muuFAUU/WE
t9eSTTddcvjiJ2FKEwunFQt5ATA0q7bAbl8kQ40G/bc21/7WqeVMO2OwytpYfXP4
TIs2mwsAxcZK+otgroJ4BpRU/j5kQkCDIndnZyoJ2CVgf7L+I7h/W9uGtCVza0U0
TXcV902zNYxF4q1kGTOypGSOprAnx02asWoi5wWoeGb+nE/HxtT7r7upqyvJVYWS
vSpPEgTHxw+NIckRIIUGplRfbQSiEUbPaN2wFxIUsHNqBnpwUKGp/QF+yYYLPLns
KbrcBwcYVaIDWB0GJcLIM4RlR1y/6OG77VSMLwQFnXNWOvDeDEm6OoPZ1OGFsBxQ
SdsBSK8ikHIFe+VnV15D0UMIwi/c8hOdiCb/FbTCWnBGN5qwhvskIknsmz5MVsJi
cPecp0/w4ZWLu57qeY7aRLGZbsxnEmJEsq1FVo4ahth6LRXrkDykA6V2vedFFr72
aTq+Hdm29MjQcFFjtngp5tFcZbT+AavDbNv5dLRtnrJYdLtGfU5YjW5WWhqbYhO0
AUepjCpGV3ldxDUkmXxLeA5nTe27n/fIokqjrnVJsqWGgh6nysgmVIYQwNKtj5r9
QIv93WHjudbzWKGmhMLpUBuS4CkAHULj7nAm5+//EsglSHVze72X7eGHxkXYAGYZ
FtPgJEudVS2nr/Y63QpSCjGTDDtK+nrqUy9DNVybDEnwu1P0tH4iu2myR7kSsoOC
MgUkr1WJWRX0hLXpxvnoFtgkG9KL9uqsYBpmP2GBuVkRb/2dMTltftPTh/tboGLB
T/IZRZ+goqKjnfj2Ahpv6ZgsHoHbS1Y1Bjh81u5ja2e7vXMOfTmOyq1PwJw6rMXu
REXhoZ3tvWijAgvQyoNkTMhdqgSO0stWyepBq9Wq357xQcGf8rdOse6P9ULuhj5e
HPFt5flbzicsdUDG4+WWmOMBf7R770PuSWkEncPZGCdnGjPrl2VIR/3KYuQNNiXc
sYt53qZ1ZyEMsEJH2zLiXpI6Y0d6VRW3QDvUIgHFsXx6CoR2FMGoiUQR/NXLNgsz
reyVMXyAr4U2NVJAKh4TV/yMLi9jUv3dqWj1gTREMQS5Rsh2uJ3qJzZ+2Hzr00+u
sKmYCb40kn448gPIJquM9w7ScLZE8hsJ1cm05Ja6be19GERtwWaE9VkVKmX6ZGPy
3/2V3TwyIPGbhilfTBwFHzbVQDBoJrsp4ZyEckiE9T7huiRhE7OV8E9I04GSSJew
EqitHgAvt3poQXEm+0Svzb8TZa/2XMYrxH/cq9VI9IQuhKqBKtrYlPx+UBKoN0K1
s5m6et5N0l8Cu05eSckYB0tHSxAhZT+vkFjlgTBn6vtQxDMjDRAsW/FaueROhTRd
0SeDVlZuZEQ49nOWRlxbsr+XXLkr62E+R/G+deLZZ2ZBaxv+NaxhoULPWYIvbxwM
D/vaOryjx0B5by+tRs6XBXKtUwkckBQjRLaYcUrQbFq+gLCHQr+E4QzD5zZOQ5Bf
IAPoF+HukRDWu0ngI3S/BdoUrsYD+OfyH02yZn789KZ/OW4ds4aEebAQrMVuLJtq
0yL8u86A8/y+kPEC6T9WHvOokadhfYXrlryikp1PIvefFelf1RBqiVB9+ylB4pbC
2nijVqNNnMEjbjm7WtRvIzelQpTKZs6hPNT9G0hUlL3dNjmnOrgpttfC0hLuzDm5
cDsXUND080+iLNoX6XUyrF236DsdefxtFIVkQ/2uL2RNqAdZEa8c6ImwCmKK9I3W
E+TMs8vUUArQfKeG4UNgQah3uIqtqBM7DYLrifM0muL5YVygne3x6uZ9+4/4Yjeo
UpTx8m+J11mBpLUDMuP7AZY7oXKemJ1AFXUaQuK11YV9ZGW2bgE5KUOy+qMF4oQl
NzaGs+L91+Dp4hU4hPy/rJS0xwtaWQ3U0JPYg/VSMiL0Hbm6XEHHmpHZkxF3HGHH
xFkbGRcXMYQPp3+2a2W1F/CasSdopBOdsR60MPMA1yZWtwOH+1ekNWOLpIycWrQM
eyKNCNAcH0uuQcgQLrK8V7KMivfm703y1mKItv/KK0SmfAJ7Xm6TgNkkrDCSnmvY
A/Z/OLnCvukkIrEmjP+RdYthL7XecyuntDyA+HRORkBVrhvKxmm9sihz/mpHnSIw
tPe86IL2QQDpsSyXsaBJBL5T2vs+iSWzbeRZPwF/xS0PLMA+yIxnRzsJG65aXn3Q
EfjQHmHrBGpnSOVkAvbVBTdtl4vKyqvY33mYhNdugEM83Q9Q0Js5CgxAAIefpKqt
XxM/iTjofbxoKLSxdz1ydf9fLMbL0kWvQT8vPxrSFP/kHW1TDevdgDWZ5uKhMy8A
TwuK5+6kaEzIKGN0irn0KSZeGFRz4PKS3B/MtmaxfiK8C90bcZEDukgrembiI1mV
7tGNh5u+UDqHgp9qEuq7DcEs7HdB959Mezd/Zk8Hr4xZdpl2BEMRslcsautvxoEd
uquykpe3yxvicxKHFKFW305C5S6iCZ26Ti3a0Y/eBtg/6B3oqTxDTKU3O3MtTkWp
10qvY8sHO1ieu+mglK4h7PN+ab016nng2V2F0ORGiwSpcNd2uc2RFw6d3RXLrBBG
PUpPrfkch4SLGxbxSWx8AGkvHgWHY7EYZbzBGLX9niOnXC4gSQfye0rdrs3vBetA
q3WdhGEWhT2EFP7HnIDrAnwgDt675sDk19fSTlj2F9b+43Hx9y8xCqTTOJmulFrK
uYNfUFuFkw7emN0hQPJlwebGxFxm6/5SQUBdIDXbeEf60pDolOn7ADQ0AAgXtthf
RMRJg6G+xb0cNUA/uy7LIQNsXipqggbD/q0G293QlqigieZg94IcsI3YnC26iKTU
lKheZKMokgBovAWEji9v0UhFo38r2o6WQLaYTUN3B69b6oVAPAyvw8uEc3g4Em4Y
VJSa3onp7PmQ2NpS4kPNe7+p3ncJ6aY+Pa9oBR4+pK17eIQQmFSiqaxpd//KVatt
Z0U7Tfq58zTk9v/YPuvFQWiC71O1H3q17gUNxnFzRPx99IrPxL6MCPOIpdq8asiG
EEoG2QB5P4jTmy/J9iBLsw0dIQhgURia1ZYbpx8E6trxWl8tfqorBqqLPZ7DEFmV
sswRGG8vO/qfd76oMxqZ2tiFWfGVNhlAfQaxrzAG++FtRQwISQaD1OlPucWWtakw
ky0YHbge1LoXK2MlkrUxXdE1fCbEghYVoooax5mf3SBS/r69k6pL47WsL6Xpr2aT
Z/klOgCxVrFHMRxsonlsBUZcbrqZ/hhLpK4tuzzvyzQw3Cnec12ri0izKixyA79L
aJRw0VfJJdtkXf7m3B8rmkkmu3n3aidHaEOq72qhCo29hGy4KAIrV0QhBnJis4Le
vtt8ct3346AaAVrPXZHLPK3S1pocuk4sr9YUOAl0FJ0Yw8/ucB0buqBzTPiAgdYy
8TjRL0WQxDyBCJ0QAYUrQ4vzjNHCj1fCfabE2bRAqs+W/EtD2AsCiMNQP5V5uW8g
ChKN5tNlbXE/I/99PiG46/eLGA2Bx1J91Xy5sGOEznBfaczyt0TlMvgVUYdN51OR
w0Z9LXrZe/yqRipr+qHAZ49LZwh3+FhR2MF10Bq2kj+ZRDuZMpH23BYrOo7G8H2L
RbS33kKXZ8p5tMADjHz6L7N1H6RGs7rXpy5cR++1NVCwYQWJQbDSIeYHWtHqtC0P
4Y8GsCd6lxbVSeLX+QdI3s3QUYGybpHjkvki2tB9NCgWHcfyoACFE2DSD7Cp7bZ8
lFVuz0P9YfkiN/kNYI6clv2XgS96W4wyJOhMQYGV/AF6FYUo5Rx/NUPU3+y0Thky
3E1zIwJzSfm6xttCm1rVt25VWWrMWGOtPBvm4pYJ2kGIColvTjc0lAxKVdvzOGOm
cc4fRCgXTJPNPr+PEanGNUvg1UkntYWAZvX8MZemC4ser1FLfzOGbOdbTTzKDupp
yc1EpAtg6ohXjWM8EFYe+aq6YlSlk6bIVBOblewzKd7U0CQ8UD+jSbRdYQhR2hzn
j0dhrs0m5LqnLEprlriCpoOquj8LHI5nOHZPvJeHjA/pJsSvksiU75kB8MKM1qFR
f3AjpkP3g/s3FiS8ugjlNWBLwnnyN2te5+qw4ay+8PKOKAZAtUUbusLGN7qlkJu6
OorzrinbDzfMoUCmWyVeBXwCutVYVlOIqs88RHkqcy6Zn3hcZtWZTl78WiiUR2ry
/hMoLuBXaercDqOSsfG3H2P2stOObw2YEWBWvVgyyau8aJ13Jyi2r1HnDfHKHX9X
6raKRxB0lecug2lcGWpf+QcLasIsnELAvZuzxkt0/hgo67Z26TknFlpPlSKD3FQN
/fDhORX+gu4TmTdp3dkHQfeT+OD2Al9lHMnF2VDJd94Jn1Pwx4bZ2mHY0mB73nYc
w3V34IK5Ah/Netxp/bNExs4IrYIFlfkI8U8Nf0SExLjxRWRP/b6fRa/vnzgGt5v2
CV1sl2ud0Hexon8mWrwsMGXg7e32MqEihKsHdqJP3qlV9uZxiAmkZ5hqbO9VgLeu
Tx/72QaT9/FUwtyJihd7WpIKxd2eKSPZ3uLfa1whVa5dk0qF2Q/wCF+nb0XDiIms
Q39q7ldcqcP5t77IJs7AnIOTsougacMdiBJJdLNAGMzaUpNGkUYY8/n/ipyF1MVm
ks808m0JiS1JLcvEtT47ejOnff39YGReTpCQo/g1kZeg8VAmvrUSxZSlVQl2yauy
ah/kYCtE0syo/5xfTW+HkiwYz7CfbipUUuz1pzTUIy7cAFBKL9glH5pbMxkrpudC
VmUfKTV9OBcR0l9cEYzSktbUIrda4bFGKsezq2/tEPe+I8qe9/xqZ+7pKHLZn5Rj
h9gD9k3u3hynegqFooT1z7TV6JIXqogyELBr4BS9Y5bLuQscGTKQFwCtA5BkZ7Ps
2HtlJWzrCpGyNf7J178SGhXhaoRRAKbpcljdk7m36Gb5fq9eSBKQQ4Q/SHgOtSPk
DSxiixDYQUmB/minTbwEEtpxCe6E43Iu4kX0Gqcck5d2Ng72jOAsbIiFHdsKw9hY
0uaaJwuFh8hDAqrH1IRuz290wx5sV4L28odUt6wswoycS1Frgb/feIL8J673RkN/
AXSuXe9qgtZ9OeFehRivDvsvsyfDy2P+whzcWNjXewMQwpvf1FOTuDLqTQBwCGqQ
e9MPECsViU5HopvMPQvRnKiw0p/0ToGOI9BweknTdq2UgEZZNFyTpOOnoahN0swa
3apk+hMnGDegF9UMHSN5o2qMuGBfTk9Bh8qzh8PbOyjBeIk4lMrbMKOqmpizOa+C
rGG/gRXZyhDOM8/1VtlnfNAIV5VL47JZQf1ZWnQTnUjbCoZMwTN8l/xls3/q8JHN
JyMehP+0lTAcynaJ3LvKBtIfPeT1KZsg50V7B9Q8px3cOxBwTb7Z8rCaDXHzbVkn
X4QtzykoEY2usfeMsGXROSuA9U5Pdl2rDehrSAEseN7fMwVg6z3xFUehUqgGPm2P
8s52ZKM58xbz5JOxEM8a+Wfj2yJGSALgYAtNrWfaHv+OCKWxb2h5PL7pacrETHOz
JVr+KyqqR+2hM/OMRXhmXcWdh2JvQ/gB+VRVTlkiVbp2+17IcbqBPdT7GCCYhmnG
1wVuetrZu5dIRFHuKcHsD+DDHMFvztQzZ+CQxigV6oRvX9yj+CK30GKpIZinZqN+
kJjDmMFC1DkrRoyWMGOdZOml8kcX8DPQWdoCLY8Wgjz63KD31lXIXTP2D8jb+w0G
4hk/2WDFQAUGkvGvz5NVIt/0UB8m984XT7P8SLyNIBqKS7CSyio5bM0cW0u9Y0cv
kU9wB/lzVYgnh1ZEA1269LLsfoBkjpyibSFjTNh33tHJ6Q6Kch1ZAL191T4hCWvQ
663uXRDvFyC+tdlGrJxknknf76J9gPvpoFM0lj0e+YO9dXAq5jB7mBpEnnrwlIv2
ofnN0aeggzf2eRolZQUL1LwrHeCPhOE3rSNKempW+RROyG/qBHHha7jl9fHyNaob
G3vO7LiL3uwlzzp980WAEJlKxkY7/p7uqFMzResWd4zdVfWwEmkOuWwGiuDpFso/
0ezZVUoIyfxn5I2m4A72o3Hx1xXOwcTCAz7fXIoS59FeahP2G65tvg6aO3J05yEX
baKNsvD929soBLbWonV9CLC3LLkLUguZ4MachGGXRpxPUfzvkaSxbaC92qdSIZ/G
g2l/z64zTCMBTabmjDs7AkGlwUO2MpuBHj1mPNMycoT2dymlm52pzitP/4HjjShE
ocJngt+WLw+p8yq2tMRR/s2WCdITkp8dcSkCHqpaSYZLF/pbtPKWAVt2AjT3AyWF
d+PIrSGcGhbY/ocKKk/ynBdsv9APQsFBTRGU5NaYc0Kr/2DyUXpo2gnWcqCZfgPC
3Q1kz23HbLmsrXAVis+Zr95OfNIDwJ0sDp7IQ2zJj1ycF4A5PUEn/llfVCgQPPHF
WeA30OwefZJXYuwFFieyXhoNJBg34IhXrh3Vt7R8MFfSlHuA2bj5Jz0GLuVhGp7K
AWYLBGlaBt3gJHgEiCcXiQhjT2OktELB6w7HAvczNDxHkdec5iNv15Jd/z960kgD
tggLg8+4z8rDIVHXX4MEGo6zcy2gRuJtbg6WhTNJp1CT1ch92Ky8d+ABnxWmVbvV
3lesuMHXEE4t0KG7r892FunqIOro1/5vI4ZjKUKqTmglqxzKNRFWJZzX1YsjDL7t
5k3IyCHk/zJU+0EsCTC+XF87FsN/XIkLGODYBucq/yh+bspOrqyJCaHV6H/YAHJL
gQ175MmXCi6KZo2lvn3VI2zQkLbFaG4/rv+NIa5nxZv4Uy1GezHZEB4zu+vqZET7
fBF8leoMlN1HxFfB7rU2DZSqjWvETyLC+S/Jh3LjwB6W3OhVWV4JQeim93x4W8TW
iZjTdxcJZfbAlcuJrNkUSUYjrO7Sq6nnRT8tZZyq2JT8eFV5W2IvtDdukK4IYKEL
8JU7aseOThE4/m880wr98+zsCFuPbEzhNGjyckzPe6FLuRr7urNv06bCeYTdEpBf
kvxVlFQPQSAs/Hdw3WMDX4yZACdGJTgpxz9xCpel6XWQhVQvR1SNA06B+UmWmyIM
QngVlw3lsv+2ma1nv6qT9EepndRZZHZ7Hekcn2q//JWE272XjuRy0cd6zDQWvofB
pVjzOCulcJ4b8x4ttRFiNBF9J/h5OLPGiCFV721bwx5/xmsKFOWWQ7oFLoMXpg3N
1L+JkL6EI52jXiBRzwDnwD7IXXPczjAUkEa3Dk3XEWZ1K07N5Xywuw0fcNHjEH9g
xAa0GShi5DEjRRB6Bf5mZp8+X1eG9k2qsImYDu6Cy6p9YBhHx5+Mg63vqkEZA974
w7ypElSb2kN3ZSdwaK9L+Hrg/6NYUdL8wgrQNWigmKCsBgRsQ8VHpbk91e60ayLq
YeS+P4qrx9iCgMan0+I0Og9WDUXluxNHDwY52agRGRvbHPdlFjszSt6ezcJtm2aZ
JWCeTWFvxOCqDaq4RTXpuY3OHGqBbzZ9E4NUJUGgqW68Zx2INEvtweBkHv2fkvHv
vkkIjWxgeg9PP3cl8e3lu9RCmb6ZYvm3pTJS7o4f8sCdvIBWgy+fqFY/cfQBd38S
w7djSIhoZ6zFOZP3gpR+vg+I8lzYSwR1tX4Z3B6SJTlvGMAWrlHmtPeVP5E7gkGL
a0Pbnren5Dhvg89WRm5rRTg2b/wQCa3isfhTyelDWwanS1EUukTZr4kQyjK1keGw
Jzha4I5XyDNIHuoL3IfWpVZI2pKYN5tSJRCpzUa2fs8klKX02bJ5VSmKgz2oG+HJ
ys8iT6Xw4l2Yz6c+HAmk+8pTxALk97Zgqv2nd2b0gVrhbS1KngL146JqU6v6ROWo
4l9+uPjIZuJp4A9RosV7AbfhJ2zdg/WNF0MxKqqyHh9xYTReeHnvC+FMqNXaZFqJ
nHlFqD0409qgIyMAdMOrvv5LwotosxaYovX1ur3tTIeI7B3BHy/rJf0KN754v97O
rCjo9Hq6JOWZ96Gw1HJ1YRIKHwVBtCCWzobTvkpjPMtzDAmn8N+7J8wuSux1shSw
HhNSZA3/CXtiMYk/TxuP6ASrzZCJKqxVIh9BCD4pipBWiVBaFyH9byvY6nVqC+iE
dTYCdKLbZ++vZMTDZKP9pTD4tzU8ZmhfYuf58+r+Xkhi691R8cSQdD1vZiNoR+35
QVkfX2/wdr8Ahy63JRJGCIXHE84g68PQiRCNCWCx7l6act2oyWgdOv63mD+JMGHC
mEj7M87aNf7+RdrZLfPTFAUZqlwkIAvVluV5944NUA+Qi10Hv/iVOj7ukm/DxO/W
iyjsIW7k6Ix8eUEnhQJ9jWCWDL6c0gjjTQIbdJ64bNu7Au3Mln3de1cGmgmsYboX
MpAU3JIliX9LTWGHHDijVF+Rwjej9SyZ8h8p4F8zQaUyC/zHW+kslN5fa/vDKZbf
Jm5r5XUoYk9uIJMfe7yfyB5rLCLHr1i6PQihjjutoQju/4F4QJr5LjalOmoXuiIz
iKg3RP9kvZJagFLtLhwBlM7pB8A4oNW0RT22gAovux3wfNyHYvqLzjpuzoqh6YH5
WpSqYzHPtvyrpEKddZcMdeNQnYrTuGgovgn4ycufUFqfzOqGobaVqZaxvGxwT3dN
l3QjSvpP5I+jwDIDPzGIqaI/JX27EMRJMPmM0idf0R5QFG7Rvz4S0L7sPDw48tx2
d8paIWclHJLFFKVO96q1VFaJUTacgDklCEsjsM59eYGQuoMKmL7n9w9NEyw21A1r
F3YKvT5COGw4aDw8ZmtayyHkRuRMkHX9ID/+sAI6iqjDOk3XeXLDPw4mmbiyuggM
aJoGppl2Dya4cmetB6dMEgNcCBfzdqMkjWBouO32AYXrN/2qiVqm2K9zymwyB1bd
/Dt4kAs5MBnqzalwQW9LG5ZbP6eo9PZmTvlzxqmC8hybsjgFuX/S4U4ZJD6ivKUG
C6Cqg2KRjDVLt6AicUd8slw+gTBh0+WG+5QpVuZOPvTlQzWXYYsytC7S01grQvzO
nJgMAopUtdQUXyin/rOxUYjA0i3p7ii9w4KK3UNszNdwQjlwbRJEI+KHICtgo8Uu
APrMunaY3KhBIsaytWg75W7zf+3+NXzcw0tVDMEx15/QNa6Yj3q3mvLNsVwHJ4bm
6sgq8F1M1uiRmQRd02YHd8r+u7Bss6S70wklTWOpVWowrx3UJm+GjguqxBJGMmbn
KqoHmipPTV13WNpaJxamYZPY/i0xi5Y6S4mNjKfJycoaDuRLFxudSeRo0DRhot+x
wO1N5nK8FBTDtVlgPI+YNcB2JpxZrSH09qTrzNMBpKo2xA0WMvgyQbsLjHRTgi8c
DWbbYC6U5yx/6G60uvX6cw5sh4jnWXxtffgGQbMDpwzgqxs2puuZH0tne46vFr9X
59nJ3mmSLtRVxf3KTjRaOm8BT8u889ZLJCycaPXjmZ2JAonctHT8kc7FZ14uyeor
rYCLHRV06OQ91JdlWPq/c1KqVyBXPhuawuhwc4O8WwAt1cRJyQOiaeEwYgk9H/A+
IC3LvvujxjHIHnGB5LFSLh1rg8tB8rRNnc7UK9c/E085cOiudtpItNT2XVvTyV7Y
UF6rmsoOQSxFYapmsb5kX1oJIlKJsOT/dGmOlYW0SYQmHyNQFYji+K7tOWaJ2fus
tsUxXGYhMAqgA8o/xT5tFt0nacrehkrZsCXiwmBI0eJGj19Jrpl+5vt0YnwanQ/s
QI2cTtygFX8OBJY2SgqWIsgplFXXsOmQdsjl8H50fiiqMibt60xLFCTyOpPuSQ4B
34ycT7+CQD+Y7LF0TkUmn8dNfsdrwIrU+ymHolY9101qWpxiCbPou80XBimQwcL5
SeQYXXJ/PW3NMSrO1HA147zCb0ugu3RFkqzxP78rzRFSzqF+vRHN2nkso/8G833k
E8uJYoLxV48MHG1tUbCqEzZwGcLrpUVJnEvL+S5s+oCD/ikf3nCbTX1VgF9cPPva
/q5r6UakPWW0hoV3EjLUmxkUEXoZDink0ANV+ba5976eEihA3w/ttMlr+Dpv2jqU
+mxY6bc72xtVBjNNm6Zqr3CUmfSi62SsZijGCaO4AU2ib0y2y1jfxlZ1K4a9APw+
DtTmPgvn2LVdxu1fNMViYLW7QgxUK8htT/+G9Eyi2DHiVC+X5KH1n+85fjVqsNNs
GdDIX43g+Ww5QVPWygVIMgWYomTM73vcboyIFRSux/9NrykiGEYdkZq90Z68gKuT
6Aem+D4uJUh/2rF/ijcuHFX4cwie1rAXZzYYvxco0/RlTGfTb+C5D2rLKaSmzRTZ
bRC8Fsv9d+FlAjzEPu9s66sLbYXxNjAV0Ea+1nsv1hC/Fkr5U6a8CxI/Wj819Hlw
j/SFgC8slQJuEeuTGdsZ0QvvNvaSnBn/RZqfbQ5cLGBI4xUtCXZ65oGjjQsMLEdG
+3NGr0YdEkIHPajEv5sV6Aw2Rd2gavujkbTmBJ/IIhzTamZp53D0os7TuJNdluZ3
2CZFowh/DWv0qAyMWkAoeNwg7Und5OuWifr0OjB8UDq66vxeWTbsU4M/XeBLp8JK
kZ+nsWE93U+fixK5gqsuURjtlc9EWDxI+GD0iXcRh+yAsviJCbdFH/Iu2WamV3Gc
DUKMVM+snKvSGO9MGbrLKxjz+AqCBVf2ZY6+pPumu6CH6STSCUM2hWrwwuUrF2jn
KskUmr/WnAtBpe1htu2nKA6GmJ5QLyTQ+Zw0h7hvVkY2CXGmAD5aba93tyzG8riU
6UY3vsAzr+vEqTfuzBV2kqbRQoVL6y/KYH3EVlyUiLWnbTwugejKxWF1d725jYmT
jsbmfP4XVT+HMGRsbDPH8tNcScMSMOkDeZyqiKv1P4Qd9qTxP/3r6lMVDXI6KUK+
ueQFrnj6/UfBxUcRClU6fWTmfSQd6ekJsP5OP001y+F4lRgo3pVcVyAQMShFHFwm
Jug7xMCVmWrNryr2gjVkWHP3I7Bf+9++bGGlVZ1YoHthGYwdenvMNpVtAascQuDn
B3A07y2hytqxnFE6T5LDw+70qNo2YEg1ovMWt5sJd87fbNJCb6mllYjjne8nKAe3
V+6ZokKX5Bkufjbv32/Ub63kAsLmymI3U32Nwc+2pIl8McFfdD/zzBwKg+xAvoml
3dwUj2W6sK63julze+tCDBzwch58RmecSKgqhchSUX7Fbr6irUWzU0Q/AxVaxtFj
PVS/3uI+B+s5/iU7JR4WCAAeTDaClwxf4Z/MarU0vAeO82pmp9TWkh/YbD1tKEg3
Sxgw7QbGnmPMSHerPHR7BzaV5hajnU9x+TvcAyTfZYFEk+mXpaDJ6lxcz2yFb8Qf
NxYoRRn97fn5u6QTBPxJ/AGszDHVW468KyM/vkgdEy9md+2ZAC+nZpXDRi3WWeD1
Ylln2QOxIjowHtb7JLEfM4mgTkkE44b4oTfi+weI8+2dBVj0C8RBoD4ystzG5E7o
c9K46R9S6n78GRdc413XtI47mqufo1VCo8EHQ21cnjPRidkEN0sDG/qNAGhCj2xa
GBRHwLTrBDmx1g6wR/hMb6aDaUFFZ7cvu0Uxv2nfOS7Ld19MgMOGssoCL8P68syo
+1niO03GyegsDrFf8aCBxDIHXapMOFSDPk9GRzoiFwMHkcXGwk/J+nwQ3cf6Ab/H
1hI2BOWO+CKCYInGl6VV0+mzXhzmNar8W1lLiZIoiQaZMFfTst095Yl72twWY46v
5NeEAYgMDdWUUQ4a7LDLqAuXxJa6y56kr9q1MXM7QolzCkdhmHLsp0OyCY5Uzlwf
cRrBQSEWmzeOtd75TPyWtxsfj/oybzbD4NQt4qRb6TxkX2z3rkMdHq7Z/E6BjRyU
5xjMxi+lpmscO4oFDkXA1BHpDc77Z92j4GlpN6p6oU0FzsIR7vYuuHPJbkba6tXx
KdI4BKkbAtki5MDuCEcoaht5xXY8cqMDLexIap/IsN2MOoq4Rxcon0AhhLUP+kpe
x7BWFwY47Pl541thbVDx3ZQvPY8Qu1jGvmf65TOUFQ6jznGL3aTLcXOBt6b5+xmV
LS3OYJ/vX0x+D5T1KBAa1HitiJ0W9cb5rqNuLfXmwohRRq1765CXcRtDrLeHXs35
m3FuRnOtM+w71SWxW7b7Vyn4isAQhtEaDlXZrqgt7bBBk4azntUIsrJBZHhqpLxI
47FSA2Jd1MlrDnfYvH1yJKsXULWg4ysqrRVnPVK1lZuTjcm9SbJBP3lgOLYEm1t6
GF9BChUSH3B4tSr8D0USpeHiIhhYXZw58R3CbidCBDD7OU+rcMZhkHCHYO959Sjg
QpGEc0auHjduRitovUk0xY+58Dd1jx2SdP6gSK6dIucQqf9iFWt1ZbCAgCwFXVXK
AS8mzraIawFsj4pqFr1wkEoiGSHP4QmikGfU1UIEZ4hhG3WMQ8po62Kw72LoKQy8
xvxmuEjXxHK5zAGi7iHetWXy180Mm02H01v5KSZFXuXYTfuVSzEWEt+DacnFX7AT
gWb5jRRAypE53amlB1OGq3moijcn37XFXLLTAeM2U6JXY3x+kwuwfPPduWfy0ZUG
Ns6cJR+VAj+z3pe8RGeC+P3vNUHhljnvypAjopIgp8Y+0nHq2gXju9QARUUBZILn
sOu9Y3Os7j21OE7JUWd1vrkHXgdYCedEHgTXujcjhE5VrINbltDyVn533IppXnaj
+RCVAUej0AsiOFVfD/2FlXIC0fuj3JfeyfzRAk0nKy6Ww5zhNJeN0qf6pUByPHtx
iTPF62LB5JiXFs86ODohRWCnz3Ngxhz2KjjoEfWxnZ3TRhWBm09bV9fgdbmS37YV
FjoD+DoymBGsZ+x566lNsxY8yBRXVuovrR1u1Vb32QVL6ld78ZiilDU8lPSFvX5s
/k0l/JFIoudL8kbk8KDHoPqkalcxJhd8xIj6k1e5SdDdGZ6fuq5tDShsKRKqDF58
aXMEthebn4U5FAkcplSbf2jRfJxa2lNENblx93yUl8yKKLX21Dllx/pPTEUeBKZU
IfOhhSWxj9deIoT2OhAzXxveVDZUmayQGTV6rG0p0T5eoM+NbdaXQb8/dOwJzrxq
0Py9J3WEWlM9tVxGbTpCSL15vI0qB1IoqNxoQqfGiCsincbDpcc15txAj7/VlYDA
fEwpAgriJz/WJKO4uLEETiJUff7ZWzeH+0omHHzUlEN27EBc3vOiLIAjorpB7AH1
MgALcHxQg7IpFdOeHalCcmNXzri9+6zl9qGuIExtV9tEdYOJiQly6qsTdvVzowBr
X8U2X/shY8Ib9coXtMQgaMv4wu+txiJV94v1EN4CUNPBfUjoGhU9ziIBkq+eHim8
2WdFLGoQp7Wq9xxE49Zxbjq3x94pfPu8AjvhHF0emxZNJaUcA19Os0Q/DEXsGipq
yLTmhu1nKbuICYQc5T2zLBhU9dXbGbBFKwR2jzRAIql1IkTv9ME+Y8WkTJ0wmRPX
1m7Fdcgw2ux+GcjL9mK1rlDOG2+xpi6hoYOXWYdGfn6tDYojmqYN39LOlNnBtpgu
ZTyfBPR2Rc/10M42R1usMrYbew1kxeOWr9F2VEqBuy8hColHwo3uKHB7IgrxsEI7
tpOE1h9J+yCyOWmbMKwdujqzhXHiaj8HdlLDR4aeO9oPDGMf44ybhiO1sHXMYUpu
Omcknvsf+uIz7hAI5PIxqn9qmYIJh57OG/5NFNUBgXpa9fdqjm9hnWVfKiwi+TS9
dqGhs2qELLEThym8C9AYRMsMiJrQxtLa8c/fHavuo4N2yBlnO6TEUbCaqqYAJ9tu
GzUPsA+2lGBh3owIZ6H9Gjd5pNqItNhrH2DFEWbelSl0f1OVxPZb/s6kqvzFQA66
R5caEFHs9GeET9EPJAWhvQ984L3knJZ5W5GlYTeaKKFFt7wr81eIyc2AzM5Ix1dk
nHkstkTg1qsaNJ0XAj2jlvdqMWxiTgrPumeCEk0hJwJH0euKklg2iMf+4IY75gM2
mwtMiL3Af4U+g9wtJCsy7/LZEDy4eSpSLVxaDEpTdWIi/VkEnR07xgAF2/olD/Y7
W6DohNlRhBuEt3ukGdloDJQ1kLUOUymzjY3eVMUFMtZ8gIhz4xruRWbIFLPpiXOs
Qmiwo+M1EAWrPfjxtFWZakOAGz+YRO01bcIKAA6bZsNoHS+o7AFjDIowNmpA/EpL
6xX9F25/9ACeaeEOHWZEgDdJsc6zR9EaznbsCMLDBSMoAm6JSRAdxOC4MPCH/Tmp
poYkrT2BviuzTzUFCnEfrqrBHy4BoAexmuNo/bCPdBfvzaGUWCh3kXSM9aM/ZHYe
vDL4pO0fZMoE1pgHU7PpUZMvkI0nWdm33FU+rToZS21ZAvMRypymLbtZQu0+JwNI
uPD1apovIXXlfMjuleUYB5Jt2YFw8A1oTJs1v1ZWMHy7vIB0EAgVuCnNX7go7Obd
kE77x9f1oTyhel2KQ0JdwUN44gh/aCdeIvJDFaWPIeQRNm7HH2SRUjAbd3VPgDZa
m7W2jwkO0BfN4UFX5eTwPFgfHeNRRUdknfiJy+HwlOHJwm/izQnwhQWXYlDxtfy2
WAOapk48GLxuxeDoZ8zdohPyX7FfA5jZrZP5l0KY6QnpHohIUKRZ3cldK6km76sX
yr7Zb5qGX64goz+TkbvytXIsGG8T3WLiZEDb+m01iQjYvOHK9js08rOWEghz8ikJ
xZgtRUCvfbsecUC9tuJHUinYlOrMO0CU5apErcCc1k70tYyNUXeDTXJthPaqsB/9
QKGOIbvLSyu1Qgz4hlmfLyerW968GoebRNFoWZyh5IjxKWFvBOzvAQk25HV2p7vd
V7zGnJ+lgdSr+hkrBWMoO+B6s6+VEHac9GY/DMhDXM/vStRJSnej6l1bhrn2mkzk
QBEfdB0nUl6MaYTeVS5DMGX+dOXiLrCHlpMEdVMylqPWEa/ELnH6qlPFNY/oaMm/
Y3iz65vg2CPSJYeZV1d2SljDerv5AOaAMdU5gBKm9TYU3AojZM7Qpuhsk4fgh6Yf
HfVpRLV11813biSmGyelaubdo0+UhXiycTLZ08P1gd0RxloyyAjPOZarMN6dIEpa
NiI2ASdVFbbiqRp1ssrVyln6Jfmi+xlJPUpnzkl4iAZ72x7EQUPWJPpFbFFyOo1m
KHec+BwDRKrPtr7JetRpXSgN2l1UsZYlvBnJGbTYmtWBO7mZbxehUEXnoSIs0g81
4rmRudcUfonWL9Ud0cay/70gl3bwMNIlqVXVfIIpmjL2iuOf+BwBY2JKyxTdJ275
f6dsS2EukD1qqtn+C6FJHmmgqSQHPNzWLwM77yR4ha1214tsKPWZSw9CXdHxZL3L
NQA8tIOlGeBrCNxGwbiMf3WvuOUE5aq6Mcvi8Sxgbz9Jft+qmVWi8KsytA1ims/Q
6DMa4UClQ+Ro67WarOQczItg5Vo7FXnvHVus4ezKn6HFukBB3iNahvZc5XoXnXRy
B/NrhmJd3A1JsOfmj4c8fTyzaOnwXHvhyNF9bvd0rCSBJjIeGhlgfUETd0oHW8qk
0VOKs8vJzR4kgHhBNHU53zW4/oromX+73wgOM7u3fl/VUR/NLHox7G1YVf/JV8r9
eU+mYF+QipD0paB2BioJy3wufFTrStqSZFPZMSy/ZxVUL4XnOT0fd0TswDwQ4LDb
/jT6MT8/2MmXpV3nsMM/FkElLBLDGl1QfSgdlLg6TDJFseZjJkUCyy4wT1hEu+PC
zHWKI8C3QCGyEGttSC3b3+A4R5vWdmlCXvlmbeI4FIfpDtE6UO1gS4Mll2ykNqxh
59tOtrpl36oye/1rQjHNg7RJwoJ3JcF1YqXuqgbtPHDXEKOfBfuGlRGxL6mxBOQR
ks/WbvDry+LZ+B/DVeNTel92lSEq6EJzPoi/zi2Uolr/dMgJf4aBqjLC5DjQQTPH
qH81pdBgkGL4DGnTYrdEg5jfLZGfy36LL2xQWiGicJAyiNTtGwHG0h1gX4Q3iU/E
M+CXxAR9igx75J7X3UEn7n2sm0N9x9QvdUZLM92ATxyzmxbGSVEBflW4vxLw48GV
yeXi/soMqZq2AXDr51CAha84fMiTLhzd3dyAUzfep25CsAE0qSEJTNQR5AUyGcD6
0GwA0RVALdvh3XEy0ud7qzMTCzZdEYb/zP/4Z70IV2j2XzYLP7MHnB9WHMlCr3Ur
d9pnuEENIfuzDUeN3Gqq20vnT9+/Ifm4ReMoM+w7puuCBXS566Y/XwMYR0RySstD
YoNm5Zf/z4QYooxD9B3HaHo6rt2mxVZBgAO0/fFWe5bXEK4YtCDmKBoB9GNY4ZZP
zTUGApnSWtbHuGmLs+kI+Z+h2lPzDF+MrSHYfdgQJKNrrCqTT1Aabb3XS+UvjpwZ
OfARkuW73RGtv9dbTw2c7OFbDuQWtV9NtktraCujIbH0RNvPGvBxpu2YUv8SdjP8
MbVA9R06kMaYfQXyZoIxsIbQaR6xOcZJZJ2o8nCqoB/PSu0XwOQBsdVtS30E6noh
jtBeEXnNevxuB2AjZWZwN11mQx6GVIzIv+Omgc+M/hgGZdBsHM4xANtrspwDXfyE
n25p9mVu4LtVrn65rl1RTgahYadGt0ZT7kcOKj+X2qlJp2Y6ASSJkxLNMhf/ydMx
+klJgt9bTmUK4uJSzRZHEZwYAwiM8PPO7qJrh3VKDLUBbZKtgL8iXRqyxaGCd43u
DUn/vWk/9vi9u0EDUk26i4nXYE3HfkYrcjgWPvSudOVD6fGj76UiiTiDo2g7Y545
0JHMEabWvFmHui7x3zKeVuV6dlnGgieZfuQ0gy5LR57VydIEjMJd2znoHCGFFTA8
PcZC/t12qUPvJD9fEUtbkVqN+orXiIjj2kxcgTg7DR00TEBskl0YLfocoW/dsL4X
DZf+9VlqeWZfJ/X3yCX+EgzvTjsOXaHZSAgGWySmMFA0F5DpxnkoZlB1rLq/BxJt
n+qBceSKr2mN2kaUNVeBzIxpxeA3IISKFiLu1Jj5pdiC966BjtypZlqyarH3/8yK
1nktWcF+fht6ahx8eFUzuoM0J/+a/McinHZsMBdLsP+gQuej8O3ILDFLAe4EmPJm
F8tmvsC/heOroLYJ4Ndm0HetatNm8xM7Kh5lDxPVC2579YvTC7r0lkrRdUQkOWLy
1BwHQ/dpjQAmnHigERUUzrWCeAYxxFHa/rm0MTFuWP8GQ+rpAXpYKhUQyytugtiC
nqRjSGKcOEUuRxwce+9pPmrCUcUsaD60l/8d649jJ1afJw29qJgv6Y65280sc1KC
LywWb18cK5a8RhxdLGnjo/YDQFehoU/gTw16BFzUO+w5jTDvGxpT/AqnizK5K5QR
F5Sr/On4QJB1zi46Kkc+jRPCyDQ7tdr+9LYSgtDh7lWuhy9GodrPgWHcHl5b6nog
VePoCH1eVkQKNs6PeDdLV+MHXjLGG6hJBNuBaIa/q3m4wbCRawPppqkRzfKWOeDS
o0CJAFH13EUmBPLGX37CDXnaQraQDkVF9J1ASAhm8j7VgqEqWvqdWRA1Ck0gWCnu
Y1YKcLnblzc5Bk7yr2j3p+ne51Yo3aAxNzjoqrr4OUgX0p3bYgoar0IRnfbGLlG1
Vx4uY9FAP/fSZ5ogx8+eQp0hJ2odhPOo0KDauHv+rqvVxam+PJ+mFX+nn14UW0Ow
FSKhx1zcG4YMJdCk84/cP6EvkRZQZREvJg5WHqapNSO/3RgqKDuaJ0vvztHExMzf
u8DP1Wdd/Wl3HxOkRjctU8lAt1dNYLEr056jt2N3UU36F629M31WE+KMruB74yOX
40l6G2C4c8Bjp7Zi7Dep+NbM5FIucWhab26Qq6pJ+MdG0qIda4ASbf/lcovemKfv
uzqWr7WA9tbKgZLsDcKKUiCoQlwcuvVlSVPJkcCsElZ5wm/Rt5A5Ok6eS7JTixLd
Zmr8VqtChLZ9RaX27RpoMic/Zw0PSFULW+i/zqaSsqktAb+WpXdyOp5BsF1vPQTm
+3Jeij7OoU2sKi6RDEASREc7SGf4DpHjyxuoGKdxE5jAq2pi8hP5gioZwNC8SXng
W2vhRO/6P5qsK5PQq9/RGhuvGoiA/OWyZlq52Vbci1QNdtUy8zHNOHGCr6SyRFXb
BPCD0iJciYrnpmctbBv0w1oVc1PaMrtjtD0ar0+DvAaCmpfZscGXwKWPCeNi5gD4
uEZcdPH+f2lQiq6PkKVExe+Y1Ii8brnmsqEmxZt2vwz0i4Kh9MA5R/El8xsq3627
77Sc4dQGEPh5fA2mtOddRE+c/hgIR0lIK0h1VsEleqqqJ3lBPr8C7FDQMLABp8Pc
AWk6h2At1lXUP5y1dWxwr+CWVY9Xga3SWAbOTNjzlPlMjzg/C3fg/kdHNz7RSvx7
GuJnxDkYnRwPlx0zgh9QmD86IT2EhWOQIJTtc6TEvrZPg1hswAt8B9TuRKEl4Z7A
XSEv0YaLq7IjXfLUqF2C/Bq7b7XExIwTuMQjqapIrSmyBdYGROlFSGzUoR0biyod
fC43kWoZkVa7PP9g2qU6h5BFt46fD+q4Ac6Dy9p/5WrsxMMH7LK+DziMAkLmBRjE
LIwPPYcEqUM3Lm3V1FDA9oMhP/YHp8GIPIJfwpDW7zuiPg+6aE9kX3ZeSov0MYni
Esvk2C1ee6XJnIWByjyrYi/6lwVBtoCZiWOveu56A9gOo/tKasJY4L1dimQpKtBE
99z5dZNfIqdD70F51h31EeHSAfmxj2tg6+mEHrYd0B+78T3wBows4b0CzDDwy8tV
dnYjtfHJMX+N7ygWXyaPhiU1TEmQnb4xSVxcAM0Cq++U8Uy3v9ALH06jj8JD4Ufi
fRbQVptXLyGdRuDiaJYIZd8XVlb4GhjZTOg07Kb9UmHt3x8y8jQD0FdI+wc11nYd
dJ7yoMVxkcfsDIfhKgRtUEU3Ywu9vjQR5yYPwXQPGCGlBS27cAU7pSayMr4GHKP6
FjQ8AFtjr31apc/sBaJg+Ek0n/C6R8NvR+ckqx1dkUClYIFQ30P/ePepfJlfu1rp
WHCmzkcBCnXOI7QjLqitvWhBMsJyI6jw6/PZwBPZvbl1PVCOAysprcEeWiDEl0kN
xXu3ArfK/DapeJK7EtVVMc6mxyAF+qxDg1uVUu2XjzhMRGRHgCA6aOBXv6wLl4LA
BNsATd5KGw+LdSE4hQ4Jp1bMhow2SsNU045wqe7fwia2OWFAHdENTJv1PQt/xCRR
zBictLwWq7vu3mGi3v786/LoX+dJ7a5of+mDRdVFRJx/2rFpLeocd5vQwOAZQDzB
0MtWjiAn+bhq7oZ2AFdmTTbKb4Pk4+zZ/EEGY2oYmIkR9bh1UpQbW1KdRqgHQB/N
r1jWqfoLtAWRg+qjkW8zqw9HZbrNUZRxaOG7jTpldf4W4joHbhONiqp+APduuaYF
tBJP6od6VqondzhUsL0z0C6iH9tFrY/2q7RnQmW2ZMSojmyrh/auNmDbSrOeuhVS
ZU+SEcillnahk8IHe+dw1ywDNUtEesx+m/4zJLYeb4WmhblnBELojfjvHNcLI0lj
tFOXDoXpCgAboRrs9+O4Ru2n5L4TOBBkKWY+Z75FA4RoPsOZWUc1pbUcrt35kc5w
MqvN61rUkBdpnEWnaRdQSTkZD/b0K2LfuQfpuCy6wrDxjW56ux1tiXGeDaAuRcl5
a7a4eyZfCDZlSw1D9wGn0fgc8QhEWEyyqV5JBOJiVNuPi1iOHgKLjxdyhGDxvskw
F1MNbI5YZRptzjJvtk6WUxIGd2TjNSZfkMSPgCCtr+zpa4vnLMGPP/0IFO9FUAa3
WKfdyzLL5BEBFFr8oadjpot5w+N1ou1v6J9Fn/5cLdzLLhnY6pdzti9KpVREEMUP
a/7+hx2OCfB6OtyTk6hOOtSykOD7Ct7x7ZnNo7Rogtor7nUB4oohFC77eLj2McOh
VZUNqIJgzKUQLg4pF9ttQnoBFBLMkfJzeZF3Slwx15g7y3UGjMoXDkKXYCt+NP53
z0VUiSBSJyePgfGRJ1MTf10+ESvzQyuzJmpLLTXSIfpbebfr1mQt/OIBMxaWBzek
d2HEAckwZae9JI3Ot/+WtXFxLD0e1lQz3ndpxmv/T1PNxeWPZ5t6hDFC9Uvp3dhB
PKXzAJ2hnfr5gkIbnP/yXavwmJLHD8sAHHFE431alfjyWiENXVR7PZ32lS+/s8HR
8269q1KHoeoxIOHW+p5S2ub68wJBe0QRCJgUPcprUBnlLHmnGs3hrpIChsYoaaIP
b7BC1HcEUaKw91P6XDPtJ6DzLEyJbGh4uxR8oLviEqLkEQX7/acFvTN0khtIEFJO
rVYuBG8JYPZiu5HZ2iTfUgHZwKtyQGt0xp94QCCGJ+g0fs5bnvwazhsRVqqJQpMI
aPZsMC6DFhR6k8R9GveUNX3R8iuIAngBBrTxoF+h6A/uk0lTP9CqaGgnhDp4YjX1
vm0pIa2L03vyQ2RyN7Xo1IKSWnA0GdC68rUtzDkmL3pUA16HRAftFb9w08Wg5HFz
KoFVsmrF9XnkAONBe5hv1HO+r7PyLhrTkQT4iRRzOGL4pB809SUp6Uf+AvbtgkDr
Gzz62Nz1xzCxlQe+XiqRS2CGa+JcNH+j16aEBBcgx13lng7OkbYdIoL7Imtmqlmp
/nxTvmAQNr+GStk4LeS2LssX3+vOweNrEWpELm4Ciubs05E3XXyar+bw3wk68ANX
VNf9oz64n9jxy+vsONNVSgeZtXiPkimdcyetImP/cqVwmFouR09uGzwE7NcjHeoZ
a35TlpX7U4BN16NkUXL3ZVKQUkW3MismGxsIo5jkLLMJvBlp4kuxVVxdSboEcZVI
bfy6tCLJ76jHQOoDAltE+6fERx1Q2eiioMmVaV8uY0feQ0gLs2oQK+2c2OseFXDw
IIvNvmeGipE3QRsvT9CHoZHX3R2RcJvgptm90WVRzwJm3pXQwm2nGVdFM9FtKoQK
YYCpXed3uEeBf0Z/4sugwtg+9mq9eev2j4HQiv9CHRQH/QaKq6vVZiB00ciUIjgG
aOYmCNqsoKMLTdN+WoEhoBvsi5CIz6SSj/d7YQDDySrx8PGhi7Jft3tvl784Wc6s
gJ2uSkFPbie68thWvM7+UcKFvFrtAa9oX46QL/qWqXkHuiGjL1dPVxlCW9aE/qvL
SyrWshMvpguTLR9rFVqXeraQS3TuDQDBq+UHeoVGMfqH0AOSq2d6/yyKSBBarNRM
vlzjkzWHeZ9EXtEroZHgigeyeEI0jh5LJMpX4OpV1ab/6/Yh36FB2PniF6cxL2iq
v0mpZishPEN3i5JJLObIUuPFsEo1SL/Mi4xfwZIvEDU0BFHc3vUNdVvx3e+qRcai
NZGIYMdQRZE7lmi0L24PQVDxZFmRl7fquVwLlaKejE/mRIN8e2aJuhf8Hq/KEhsL
pyAeyik0qMkzs4ut3mXHe2qt583qYDsWoZY2bHgKuR+UXDYdswu1PRPtQbQBb5WS
H8PZxmmlj8Bsk7wbAid6s4U82iAe4fjd1b6LdU3JnCK0xdH2TmUCeyWcDstbfLIb
w/bojbgcNEkhEIqWRLIirJcuM6wIgY2jQb7lgzAGQe5p/J8Qipi2cuybvxcsqNQs
Xm/uVGQnr4vjzXDf/bz/zXvpuvkhHfzefqdZfriKNvHa+JtRj19otNZUtnMuFr2w
1IOlXdJLrpV+0AuNfaGn+JA31EJ5nGuQ1t5LvE9OwTnJYoplJt0b9T4hMZPfHbkT
RbaGNKHEaX5TkzAuhoAMvZGfYOU/pD/HHp0ti/1PL0ZpgndpQXY4NTNBwKgEwlzj
HgWDeLCw5C5fy5M/sp3WLkEWnwymnPwU6+s8dnatxR50gIm+uq7H4QFOnZ5AC3uf
AMNtUoc93OfCv65lHuWilYr/BkVg4BNvQm4lSmGsQuDM2mDrJBHYzt1AYKzDUUD1
HVrvzl+CknZ/8z6uZ6QlyCummSZnDMCBkoN1RUmajI+CrCoVcK1FuPUFrjtRfZqB
ctTIFLTcVmSVjwp8jujmqEGpvDw/LQhMxK/lez6mfPXgTs4vIVMnuCXWm0nvTsHQ
HK0Q00dLcvTFFUdRdyzRjKxbVk5kcm20HjKugN/Zn6HtV3JD9SRW3ZtjMpxpIl3A
eobk22t3K3LWwUvJY+8DYjvtkwmTqUHFK6tzG6L+X+x4CzxROvBH6e9242GaUi3s
1gTzHS3C66aEBusCYv/eYDGcD/IuiP2uI/ekX9GiyfaMpsgYdzTX7v2VCUrA7NT+
H6VV9JHurP+hmEcvLA4qEfqyn9BYtGfObDL/2M77XM5k3w25U0LDxfsRKpDtRyNV
8dvus8Ft2npjZEYgP/1Bc/bRHxpb/gPkUuiiwrGVWJv8KiMXjpz1Uz7qYkWvChLd
3UBWALSUC+0+OPKHKqCqJgX4Vlcw5zjekhhlPPOt7zz8l7r/WlVfEabOiOnpbRs+
zxNSvEVFNgSrTtEX+/Hwpnndwn+pfMmNVBF1yLIzwJN9sZkZScvofQtbEDUaDuq2
PI6fr4wRrfYwbJBrOmhTSEk62i8Z6qpEZSR5ns5yyEp8fWO4umnJuWk9rFoXsjX4
ecOJ2PkQmFQU1eY6uTA09sEFhOSvzrhPjhcDq0oEzgAyAPAsuDwLBEuZaMd14sN1
s7zqI/kuEmvd0GXB1aO3b0BisFUm33bsRqip2tyhX8AJegke5uxKsveeANrxjJ9t
y6YBBRj21CamaLoB0jg1Xm+Syk84BIALBu39LptBQ3xeiWDe/Cuyl1+Il/LptWW7
cM5gxchmfEfsEz2jWTPjnu+pufo8RTGYnheDe/WQtOUp4izd7J8rG2Ik1BS7vD32
8PhIbAuQ0TWd/wyL2C0ybvR7MgwsrMLGHCFaL9Gob4ofs6OMhD321WT0x8AmRYlo
0l2Bn+5plsERgdJKXc7n/1hv/bv0KcFcAd1fApy9ESpi9Hgl1vEDTIpro0YGRIhh
W8S+F4S+GfjQi6N2ULs8WYQsY5uM5dU9NEy0vCXHALYaNGEp6TXlJvY1APRJLdIc
FOUEHjdXkzGUnVRHWO+0olu8RYiDrsB3nsRyVSMSoZaR7o2qEahGaef/jWWn5LLb
xCAODhTKEOZqSV94aVgDm/KmBWorTV/LTrADROrDIH61q6C5PcS3LFZPUtHR/uHu
jQOMQiJ3cT/7N9o20Gfn0Ql4RH/PNOPXjw2ogo/F4hnQXk2Oc/60V0j7B9Prelnq
gCm3y0ndi/PEUybbiAnc/43lW1JdsUOxlIqgJp0zKNFO6o4hV2poAkCYAtpabIgj
tg9oYNm8AY3G1iERlG3/5cJDKH27nsvo8RUjv3MJ9QYmg5l2h+a6MN7XIygNQLyy
DWIPA6k/OU+YjRyaWjHXmPeWF2IB+TYAYaBgZO9vioLGF+mh1nelXmKvJ7FsuwEh
t61hBUf+jnbFYikRh/d1oaQyXZdnEaCtBA4RW5MT+Hrybmpkgzy1cZc7Z1f8Fij3
mRIf72VMbEFrxK1ZaGuRSD+V+ah+gmPtcBv7uVfaVwFqDu2qR14lYbRMPQTNcAZh
d5G2qUv/J5W5ddadw1lkmlLDPNCOq9YIbABmhawxiHTHQQadaT91PKX8oL+ShU+W
kk24SxWZQnGll5G/jiZ1dLBGNNakh+DTKsi8Dwuv0ILnratAgif2rNx/8ftgODpZ
N2qRdujm4bByq/keA3mMNZbcaUHJNc/NRs5xkG+5L3ax6NsmVyi7BQBup2ysPWtM
s9SgWZMzTzT9FWK+l3PNBk0mICppW75xi4sPtcjpraAirs/woh2REydpmye3wf3L
ErDkJIGMvYyKAYh83z4vra19Eg15Fhpcov73tSE4dK4GlMA7yXOAMwykzEeS4xJz
DfBtEpcaOawIzxIH0SguCkjXf/MLP0UHqbXjvi9at9q4Yoi7PGMWspW1KBlK3X83
eXaTJQJvcXL5qDt5lRu47afjNyTy4HfHD0NnDFoR8oMx85stDGp0RgPXgem1Bjek
7U+4AlhoJOmdwASCgAZLz/zlAMfnXKOPUqsehc6vC8jNE5qQnl801fTlX2HiJsLf
zgCLkfcP5QPCHzcyMgxeZXmlO03yBNUuJF45x98eDMg25MPp4L6+h7lm/TYF3jgc
HZdb7VBtiEPDZXOzBZdJ8jLtxUOV70nsWNNRzuL7OzX/0b7saMEs3dgtidZIlPYx
0T3q+kEZxYfjqX2uUlvqVuBherUWxlQbnZ47VwHwIhkbF0oUY0XWQBGNYEKKHMXt
ICUVmSErZXRver1xtFtTSyTdh780aoCjBsNQtNksHrOCBoBwxXuYmXuMK3kU+hW0
Loz9p7jN9g9TdWwejE3bgJGk2uwJlT0BjBFyLpLiontnFHnTYGyPyeql9xF2NBWD
CvBoyeFC9/B/z9T7w5Ip1EmBg6bxuad2x0LRMirpBY5lmctL5SMZgjPnoDoX1RT8
bx8rn4iN7f9yCIE8sIykkdKnr6ztJ+Tu+AkQvxw0f7TtjhqsU5WV1Y3Tr9mw9D7T
7qYZFoJLKSTRirFK2IeMTdFPGqvCvFd9dmjibTKVewLgm8x/5Yp3aAcQgiYSZGm8
foHcLkQl15aRmxHfby6OesnYZRzG0oJwNHwl3vlWuBuaXxipiq7BEls8dNAcxn0W
+iwkEhP0Z1pbIzK4xnZI2rUp5EKWKhFTu46jfWDDFSRW5M/BHADL1Agb/UbCntvL
/T8uq87JeZ6qtY4tV3mrWpukXLw7LlelKUJ+/8Q6pRp19CPPBidBHRiwVGKt1LMv
PBzicgpXCSXItEdGWuF5NdZ/Cz9cM/PD2zRNcwULMq2UkiWhTEQ8vdtrZ3RTfJ0r
agZo8Rre8QDPheAkqESWl4SWMl2nuihRazmQBjhUbQEr9LdAhMylWolJ2ILGetGU
cawPlZYP4N6PR8haK1QNFUrGGJs2jCW6H8oIY6m9ilL2G49FrTRljLkVTvtdnSbm
v0I7VgWAts7/S/U6wtVPEBJI8gmLHzeREQjxU+RfZXuyCxpFj49QDwf3FpJzs7pA
Jv+IYB9gNpPeFd/FK3tRPDYX/M52ozM9pU2jnEMfTM/xPIBpIU1K1B7UZtK4J8IU
6n3KpcFUuYFNiXAD8DPyiknovyShS/phGug1qWir8gP6FdxzMoc6HacJSX74HRY7
eBqwlzLlAmbbFPh+BGPcW7ZFZUl82Crsk0WF8ZxGfTum6VbROJx6/JgFd3zBCJZQ
90chxzN9p3OBVR5Qiz3TAbvWK3xYtWe3O5IgpMnCOk9FMggnbQip/GI/jCxOc9VS
IhfhyPmGqzABsSVIhkKfrjewpjGBdtf/FhFeuplHhh5fKMJGUdnxUYN1rPa0a5yn
P4bgwnK9hVxDcZd1ScCJ0aff5HsB49dO2tAVW1yGdssMris5ThrryvU3gseNnZTf
X2iNQV9Qg5aBJXZoI+rl932YRJ6iCwviQozvvmb3lKOD7mVOk38hAQtNejdFi/Ty
2KPFhQUhmCmaBTAoOQXuFQZa0LPugY+UOtNZBBflDckFL+gXz8Q3JFPzUq30eBtp
Ge7670XTCw2H8E+JOQlQn6nTjpe0I6HfEw2yQVgkqQpMN2wh3JJ7O9pDxQ0gDsjF
ad6Iu/3yr3tki7MwrgiqZ7Vka6jm/rKv25+IJp5mDtTGDAo8mCzzUf2GfyxERtBd
ZX9HWV9yiopL4fFOwyn8+PMst2wUVdswqyrIlDgWkoDsH8WzUbeyFxIPPHu06ZFk
iYLpaPsKLtqcKbJtBVxEDPDNSZngsF5UrE9XfCT5KJuonppmXgFHtRSu517MxH4L
YXcSpevVFnZrg2D65j2kEcvu9VyaF9ski2izJf8avm/QQYzYZfqI8PFAMBo6vqnV
EQ87Hc5w/spU6C4OUvNAqiE4dVirB5g3RnraN+z30+tnG95XXc/EK//2+wVTxEVN
WSGmTCD92HjdbYgrraiXUKFXZ4zI4d9VcXnxI9ywdcylra7B07NPnX61epjx1dTR
nu7GBraC5eSQHoJwaoS6gQtT3B8SjmvHTq8B3bcqUE6K4+Sftdo8FJtcDyYTRUeF
iJVqfWkeKRNuQHM0EuFxdbfSBeGXyFMZgJcoZ7LMDD85AwN62UUtytYMGUtVapOU
zg2Y2UF6hgafefIkTZOGj1gS4Y5FKBcGjp7s0nfL7xCoINzbTP3tXryxNyiXORnS
fJpX3gG1MiAeL1tt5/vCdYi3II6S/i3VAXh/CMgd1OCQ7fuXGPUzggd9r+cZM2g7
Ptx89AdzikelZaD9YCPiSzlVqLiy9dZa83ZwhDO/AVP0mv+aRRrRJKMwrk79Nov7
1VCUtFt7Xu8uFaCamfhgQPhQmO2lbnNyYO4Q7zJ7aqxxT3HiL3BlS521j1KGdvih
TC13mo74x0l8OCitCSmh8NzzV7eWNerXxCcuEKsEHb+aSkxIQkjMTMLOZjDlbtbn
OCSav434mn+9c5CxGHnEza3AM6Bn8fzrGFHIMvFbndXnEOAZxaUt9WzbTdsJA2d2
P5VtAYw0YFUYcarWyuCZItWSC7b6ISXOQBMkq3B6id3tZTUErUbJ1VQKdw6fVW6O
YmqCeQ2MFO47uMmOjvKvFMtVVr15FqkQO09ijQZFT0c1EoHHrFhLagSoDy7cWT0S
dK9N2PZkoUo4EbHhbzSCJ/KiVTmyi+EnOqZ6qYNv4yKVzGYN7zxmImN+dQ2LRTnQ
Ju9kg/eDOMqJ31SF7KMZOeLML6Mb1serA2hifX8RqAjZOlZtpURjBPygkpGFo4wO
hON0WX6AJTsSs4iXHfT7T/HFyfftSqeLu0FaFpGEREN/h/f2EwXWdR8KpJXPyt4Z
2H4WuG0eprJFgOAi8E0kUXVCu35tKhDhv8qitJ5A7RbAf0ftK5Ic4FFOe4w51ERe
kYpu+UAIUbHbVAWrWGSjo4/4SU7dQLnkYfKgCU9ASdOnQLSRAmOjo1oal2ug1Hh3
4O582ZN6tOyj9jbyIa1oTwEsTs8zv0Xvz7oWECgJpOMt0XLtRPl2XgXFCbrELheN
JQx8e5F9ZlZFDbTUb0x8CaBPl8JvJik86kZ0seRs9Z/6WjClC1twErQrdEhxrBEg
43AHwBc09W5WZBDykMqfczEB/r8ys+jmMOgxJhN3gtEWQohIa60orUJpRQka2O07
UCV07ETkMIPj+KcJCN4kbxntbCFkE8LhRI0648xvkwOdrCBa9ESO6tbjOVwkWahp
ue2t8ShL3AF+LNUfPtjTTUQ5rtPzkrY51u6ybaSkT35qNEjJuNUPKGuF0IjoI4n6
E1XQ/TGJKVWEG53xXOhh69mqxHEkc02O/4nEYD2or4NiOKLm2cJ6rYcG1J3NR7uc
9ZQSm2X6wY+J6+BxrNMlziJsuxFtIHcLA5ezv0AoSXduyBTnfsPUNA6ncH/m8HlO
+6j0fcj3vnWzknJSGc53kifUwGZba3RLzvIu1eJehYaiBthdtJ95Oh3z8BNZqruQ
G16Z9Szx3MGYt+MGazY3lBGxG6CEx6IFPDTnS2h+S6HXoWd2W6IoSuMb0RDxWBhR
+RKbojzvrWxZJu1A8Sd4PmkDrV5aEP1R05VUGryDHuAkFDHBMrxyp44Ibs1MrZUC
reygKj4OHxLyuikiqsWQrimHdEN7NqLk93aZvKMQdJGnl79Kh4geYdRi9I6Ypvvz
gtc7iOhbyvRQQJoL+Tcp6dxm34OLi+oqQXh0CikMWv4S3jwR4zhvTBRh76OTZr2g
zW1fhEGGuxkIU19YFq/iM/P+FLBrBtC3i3u85ahyhVj+r+Q0GczuTlnwme06TY7E
e8Zv/iVzzn5Pm5huUsA4VRB9BMLs3iSpeI8EoWrC53Yncye9xwzDVgm8Vl5fUMFm
WHaDjVj9+NBYjav679ljwZVfftZ3GcuUllAlqiBQb+oYzV296j2L7Cl8msnyTJso
FWMe6qVC5DAVdCSUjANl84cmdnTlKklgWUcwHu/ctQ/qVIZ108+9qxlvuPLyt4nM
q/6f4NAyhwbT4hXKq7BBDHuw5/MGiepwxn62vmtwebrgLMZgQOtwaf48TLDmkWC3
smagpb3OAhNeHWiKuxL9losbujWaixp8Ii4srx8ikBamWXbIIReNGtBazoECht6a
E3pCoOyqrsDx+mYC7K2d0kTGM4EE+RHTeCAw1cB/JA1oDCGuW3cLaCLV32rKlkj3
k/+sGfTTYobni1ujQC0dWsCLOjnT4arQ9DCiaSRU5H5e0uj8fEctvfVRF4NyNiiT
ZW75RMZGHeiE+7Uqe4xHIUr5/S2SXaQMiBBquE95UG++O8vOegfsuQYxq/GDq2Sf
2toNHNzgq0gh24V3pW1blUK69PiY7bykYKWUOBHJK+8QRWzvJCRq/rCKyQp5ol8d
C+0eoLFItKB8L709p5FFZgwvzAUZQw0t6JAIxj6rYV8zi89sedx6CnqRL0GQOjqZ
cuhJr0Ht6tzMTQk6ubJ+cFFzlnYW03cPrgzP4xmdz3Kugz1oUDfby0rw7SxbxD27
BvWAz1m7mKpRazGWtAyvYWL34rwCJPTlrHESfAchXHg/qYmoiT7OM0zRqZ/rGqhh
JIT7IxKwcU9JIFC3f2t9Ij7kR7O/uIl+zj9cvEfUiaC1TShLKrbzp7NG8ArxIULD
FTICT4ivXDnOCvbB7ARV80RKWHBkWs9+5ifH4FmmyUplyHAd7gVY+iv3jnfn0lVv
uJQ9IF5rhTztxgHxPJ4Lp/V2U0Gz5F9XGp4LARxhweFx4Kpthnys5y8KZOGBjR9L
N5Qf/ugxWCshiAfRHkExhYcIwdPvIJUVnxRNgFt6Y4PYaKV8my7ssmjuTKgaX1pX
5wfNud3LglT1uG8ffU9AVsmGR/CvIpGoyZ0jvtFnoY7SNNK8HKeMS/a1RP4IRs9f
gKdJVYRCAf2t07X+ZUEdJn0OYgQ62d3sznzaxfRv1/x0sjvGhRgZqZIr0OnOO8n2
1izHmFNjlrHoJQX2rKJKeuluiI2HelCuF7q2j6uV69YMGfhBei0BNy7lOH+lWXEr
LicOuPU8FY12EpS6gbk7edsiDigqonRbPky+LSeib5B+0lDcTF3JAua6045PnJRu
3KhWKp4ae/QvXAEX0TDb7hTivQLdOk3caJ5bcQ1ljQMiR0IXQ0Rx1AvGAQSTdYFc
hFCb3maTnu1nVFl94bsHtnZnjCj9fcXDD7uS7UxvlkWBMs1Xr3PqzAZoTH8oOhB6
5APCXRnbI2SOEXDEtTp0SpMYQ3kx/UsZIT/RRjT8VW6U9PFWQKi1pJ0Bh3B7mUYO
d+Y1kFeIxSTTwAh+CevPvqNDETQAp1eQHj6Ocl8LXrgt2NLEsw3jkU9mYQROoDPA
I/lgj5UlZn4MyU12m9vUKci59q/SuW3ZmNkX9itjtNZeMKuex9fjMNd6MuMecNR5
wI2lvkJwsVGoUNPOaxOJKUT5AmncI4A3RHMAySpC05k1u7uXD3Z1idlc0NBmL8vl
Q8s0Ya1n9jbcYgQ5U5eNvpSz3CPGs3b1QYlw3ortzgqp0NMDbuDNfbGhoUN+Q4xk
jguUvpnE0VORiz3wlIVYSVY3b7V3mlL+9mGdmbi+mwGHwlFRuEJ0lKyCuwIYIiMk
Id+NjW7MjdxnNjYShE0AwRsu9g7JA7YpmMIP97eC/WnffY0tGrK5Coz3C+FqUPvD
t4s1vsMmrDWJCCqUH7lmzJtvU8oDreAYayaMauu2uNP0YvDGCFWf2GkPz7DLe6WW
dBqAx4ZbKGj6XmRvndysfFcbX9CTWj+nW3jC+y/MPaYK7+fkZKGyA9hi1M9JtGiK
xlOy2oF7qfRjFlz7enljciS0NGq6YDI6HEBuZN4sjwvtfL4XfSz9OZU6EpHqJ2xL
YABKbbLbcPgGygk7cMUUTQF63aRdQXMkS4C45eUYs5eyQyeY0q/IC4kRQZiqv0QC
aDIVYALGIUZ2iTkHvEgJd1viZQCWvM7o5uyHaiyjYQXBJIuDr23FXv2AhGLLIQ7c
ifh96pCTLz4kcczbXdqcZ5jwQrOjdI2nsMZbaIqNZxjZkohzgcxVOj4Dwewc+p2A
P0VqNil1mZn3u42XdJvKe5uZZuvYkIyxHGEei/YoEmiO9i5jNwkxOxyMJ1WPI40/
FRueLXc1P3UYcaYrwahJAVgsktcjNrNxAfL616hFV9NxXEXDhJl/UPyWpUsQ7Kc5
0BuCY8HaFHuvnOjL4YEr6JjNB0XfpLDHMrwF/EQp8VziLn7yIKFnYTeVbcK8bH92
eEgpE2EZhnKqIZnN7vA6ZflrV3SwDC2fuzRgP9QmG0f906xBcu3E3lFd9Pgbyq2O
EDM5RCjdxzQmvUnCEodGkUz52DbRsV00pM1N6tW917EpX9rxUmRh56GxBeGrGKZl
9me19C5/wQF3xUdJq6KvbEMQdfPRoKjjTsZZ/iPK9zojQtQJdQzZO2s4p3bw4sWL
AXbkvJ4nKvIdQwDnsgDfg2oag81eHPSSwTJfISXwDCUg3NQEI5EIFPsgko56JN1s
2GwotacNNTGo27W5KKvrMlsMkkUo/tsYD2LvJfjD8Ax8Kr/XPWh/zwGTvwBPUJiW
16VGU3DMY26FEOtS/shd/Zl/Am9hCKefRIKF2apEgWHwk4kNLMN3W6jSnq7+AaEr
BGPYtf+1t0GravEP6dCu6xb/m4OLNr6hnPF4Oq17tYtLMxvjSqhgJ06PD3oJX8yA
P3gDoIp/UwbqXiqb3mJL2IHLXJzPUq/HJUYvNO/wXhZ2CztcoqH0YxaFQvjcD4PX
tIGkXFlmgzDt8pQX56iKf+jqXil4eGTQL9Ta+U57PL/9l3ilhypX1laDBY97oNCc
ODNKojr6Q6gVhn2BOpJ1gnbvRN3FAM2foDPumgEAC8f3IdMJAstBb3Xb47U0FBCb
4Cxhik1o1cuXIJVU/0ihoaHYhBrJjlY8moNpeJRP2Rlye/Fn08dFbR+9Y2T/P9PG
zW1Qo6CF7b70QTOpYEloP/j1cKR/f8JUj5GfaRpq/CoVm7/RqW7ZcTxCzJ2Hmk65
DaVz3qBKLFmYX99Mw+cOX+0kPKbdoUsURfH2Sh9KNqjHjpAQF/+qSuZcAYw1W4RE
y/ccQ4BA1UM+KTZBUXT05BEy9K4XfgIVTkfq4dAKAwo6nDs9J5/YHj+7z7h4cFKP
v5kCkpfv+r32qDBN5fQVMwjragwre8+us9ccLKD83A3y4f/jULl1JqyfTbA53yZx
ur7czbZKWYTRaeCr/V/nhJxJPK07wqhDMH2jA8wW8VISGuIFhr3cgOfTKACkXmAv
/G9ABJ8DlHRx7MaDeWd0m0QNXqA8mW6tFgTQ0LQ5UbG0yBLz6giVM3kKwikUuJzh
9YXcUH4xR5b3hrz/fh06SVOAdDoEj60IeVG7MxER9+kWdeDvrH0qJmRqrzlBW/qY
FGjfZZ57WR/vznlrq71zVnyMIbslRDMeSqO9nr49QeXmpKteG9sSM3A/Ve5P4Fcf
kbzNwHbDlQmfNX3jnrWBDleDIN7a5oqrbip7Woj61hcky6zbLFR1EHe9cCPiG/rU
8edvumi55MJZS6i2s79gmqzSiOxtrgeYnakxXGMQv8ld87ut/21L3wtnD/+9/Rwb
AZ6XMZMnp4luqOChognAIKRJDbkfvyE/D1Bp8PWR0fHhRP4+c5jKlMkdSrxgZ4A6
7euAC3i+CZnNr2trM4BDXxM378nX5P0i/CbLdnOJuCMOz2gvjjf1E/wAVRzBqH47
U66wewCMGD3IB9n375JqYpvdbBZnhVOSfJ5VBwYQXMsTR2qQjfv01PgeKFkN2pue
AdR6cb9T6Kc0hX1LsfQPlGN6xswjuiMIX67h5Hye4uTqNcgU/YrUEaRIj/PofSnH
DQF4Ebxd+K/z9+ulgB5SB/Pw70z5O9MQIo2Z5SwZfq48SSdIinN0ssDrQ2TzgsIk
o5eX/z5YBTUALVsr1Vk4O1/AhEJErNEGw2ppgmUKChA88P6kPpTl28ErEkCIl4o/
Oy3FV1H22moaGiPSXXAkTGhmrBdpUJufJLdWXoVWionBNhJ6CQFublVbfq+MHmjn
h10yqPOuFzeYyWWPVhVBcfBr+6vWLo1SgA2uWRs0VdWXRDg9VGBYdlqppJRCTLjz
H7N9QsfCwqGI+8/EXYF57LnPM50HJgU/LsXTHH5pyfak+qeTkgxenJVjJmIy/whe
PzPBaOTXSSxUms4953Q7MLjxjfHbyRdAilJiand5FRGCCudySzxlZ3q8x+nv65aW
zPpBCChlMrbpRcS7h4aLvuaL8CUqNTVvpH5/Np29ww7A+37clFTeb4Xynrkg+IhI
T9DU6dtSVlnGAJyY2J67HotR6VFw+4P8xQpHmEFDJg0sMqkeuvlmYwjUSRNE/1dv
9V99APprXAnPxpsW/aCGiWU8RcQ7O5oYAtulxNMqWb6shXFZKqXOXW/xphoHSyLs
ZyaDenejSDNOOJRX1C9Jt3DPucfRpqiUHtzQo5QDe8alfgLAZfsRbCC1HpfO3CKJ
YtOsVkuDVt8uUljnlMxYw7tcRrSLqp7m6/1GFy2vl14QFgPp9itDmxDwZaNCNJ/b
eK6+8V6V8VGyRF/AoQgUGZr/H0NbGgqEizC7DGmUK1JAu1wLCgwxNbCCACyMKb4x
02ePz8xsS11p/81jLWZbglZYo5W/fJeetNgo5fb6YwHwXlnHIhVUjcYJZn78wNaB
H/P4mTw6AV2Uk876d8QkCBfa/y2Liq42cO+oXofo5DYqm8gTyqYYkalErVq5IVNr
8rdPVRsh9Jikym1/owwOAoRoQZJnJUIBgYySKKyDP20ix1Sdbm7GAKW6CK3lkbUt
ixx74ZOkbRHXqQgN9qdelJtJdL5uc0CMXggojpe/jMkcR7Mj9QE1pgfzE034t3wZ
jwowyYvbovGWgwG9lkaHSdIpDSHBLcM0vl/ZneJUV5os8I9onBmb9C73gWJ1yT1Q
+F8MF9EXS1rST2hmM5G5Qnxdhb2MJiei5iXTOJBwOR3S7vC/I4B7O9Ihjtbkcbly
tbIqq8RkBFUqNCOlc6LZSFzZKLY4NXyMlia31p3W65bRfJlqxaj3d6ME85HCl1cF
pgOexNfy98vdKC3eagc4Ogl6w6mP4xyDygoow0SIn+GGHcqZ4JqeKyJ81tKkhrgz
gZ3G0pgaYzX32wW5XWPQFoBwcXQmgru1gKLCw3iIm4r7W5ZcMZFoW9pk3vfZrMh8
J556w6x7GdjNew+4bhxP6dTtJwi71wd0lww1h0HDiZzTwxTJi0zf0094VfNAw0rU
xAdryHuCZn1dwpbijVjBe1/TOzpG8Gg7a6pF0ppgJ4uSjkftUgMMrSv9GWXApZS8
GAIxl3Ckch4/TTmp2RXJQ/eU0dL6C8G+wgfhFGqCpL05AXlLbbrgP4/UMAEjueHw
NdW7v6VhEKNQSfbcHQC11ns2yFyQBiEIqKyHpYaRvakW4+l9mkBafTdRXnoe9ndi
xGy8AEPyObj8WJsN8yjt0jqYiDZ419HQ53caMEYRYWn22eFrZ7452SlFNXube5w+
DI3skkmCllCiAi3Gz5O17ZWSFM5WWju7dvblGduIisWEwlRAE+GyRKn6EDOv3Ct9
2qi7ZnJjvDvyb4gO6NGmSp0LIl3vDyga20132zd/gPK2ZLMa9jTNydtcjn/33ztQ
l4m/wOUJv1ky79gmM7+nKqInZ8PoFTBYHjUK5gmobNJEhcZWLo/lrKyCFdvQ+Cv9
c02n/bKBz+p4I3oCOHKwOJnQZmnozvBMAy+uloe6YWn9EWPf8cnrSfwoYdTQy83W
wCxGlrUtf49qleNX1HAoZvzG098xTQnuNc/RwM8lVYUrMEWDioyC0udU/WCjjYNy
BdW+7CbwC8mR9FhQMlFyP2dzx4B83QXuEUwdOHyxrmPGd7WQ1MnvSd9vbNNifRCN
qO512Tf0fEypQMgGQPNxdtmnncNyN7/QBPAVJJ2mTHEXEYXjxAAdTnSvr4AKVsYn
l35kTqWKczxr3sndU3dNQzzcUmmcdkLW9HvyMBFS/pmYZlwSXAwWeacmLeHKqDSE
Od0qgX06BrPbckkpR/hqPG3teAGzvQeseDZgmKSTQ9uFZE3pjLWaLE/DH6U2jfRC
7+gfnJ3Am0EuRGPKAdpY4gHJv+Vxf8tiSDLWroyvEiky5YZWlWPYqM/ID5WhzQdS
VPjcIJKBGl7hVmIfup4Xz57LQ1L0Rp82TTefknGdTT8w3Dr19Go9S/ynymhVsnE8
WOI9DAKsg1fOqJsiN3K2kFoLOPVTSM7zqbDY1+6+41dkDE7RyhoYruE0d7hRsTi+
gDlRXR27vC80uxjqtKk/i1cN+BBdk4z5410pc8Q4fdToMkAaa0Z4UPlgiW7FfT58
843kzNsjq9smCTz/zbW3O3tKuu+hDNiC97+ziQOuh1W5JMHad7w3Pa7OYkxcySQ4
Ob92cFyYwV6FZ11xLt+I/3eIXJl1/fxSHLfyve/IzeFhJpnESBvnU6sadMNC9MSF
diMEctpipThWS3Bycm+eLcMpXK80HPl64RhhLQpZDgfoa7Dm2vux0iCLAnsAGZJy
QqtxuopRJAU2cn2k6merx/lw0cFoojuND7PTtRrK4d+pryoFIQ3C6dXQEnYTpgvo
+BM/JJghX3sSusTqWCBL2gO6jhWzN8TdjH0j2+xf4DsgJPXLQ57hCk+egbapzA2l
dFskfAvEWfCf6ViIulk/tVe+PMluaqhkz03VUz/eF2B1IP33QiXSYv5tGO1+ZMcF
kpTiO17FFcB/iajDmNQu+m2mIWp5xUs/Asfj18SvTCm1Ax76PI3nXFI0L4T4Vi4d
ZTUkzKcMQVAZQqvrsw9Jfsf8MOHBUflp3R6BKd+kvLzcMs7CtCNTH+wG+Lx4CLH4
w4KrmLhNEfVKVMIfH+iDh3fcTNvkUrJWa9pbbvkoPlqljTlVXaW62gg/aSQnaRGf
xJtVjMjkbmKJh4cLaSmSwM/PO5S99CTT+ggsM2HlxImNETdpzSsK2ixvubjx+zAb
w/16FSnfQ0ReEOmmbl5vOoGaAt12CIm9A9G0RJWUnB+uGIcLI7/77vpc/+t0wF60
2OxfEpMg3jlyd0SEla9esR7EZuWKFwTPb5gFixulP5r2rEE4L5qjR5nYcUYebSed
XT73ZjYY58K+qXoFmC4XeYYf/8/cosDnnE/zKYKTOqim031XCtjicLHvSr6kgJYV
U4BLeUM9z0btW0GZQaV6lAY02obAAt0W4Jd+ZHyR5Y1mctvT2ZhyzGROpGLz0VB0
+rh5whAnggVXnoqo0zzg7nzVsy6E503CJtls3dnyC9UNA6DVQnY8Crj5WpHO/rG6
/0G6wsU+71qAALoZjGvorC7XG/pqXD+1xpTgN33Tv5j4d5oIZ6E6Jno5q/OxIZXr
WqH2w3xh9qOQKhIveROBoOg+KgtpcQLnvJRkFFtrsYADE5YwPj8xxX4JVHx9ze0Q
pgMjXZM48O4HXwTQFRNoFn0hSRVtZTfUeUDAL8NCDtMyFyO2O70/T40jyjh5+0g7
QIX1Guuhx3/AJZmG5FBa1FGSoyNqPEAJD7/bkhs9q1nWPR7GtC28khQzFx+p/Fxv
MVwOchJicY/ylGP1aDYOcVAoVtoD42B3velWPuFQDrIm0sUbjeG6JovSXmzn+mPb
UcCoHH1vJ+V2yUAtASRzzbJVMd6Mv7fe6JXToKBF8Mpgozuk8HdyfmXonmVL/wBy
L8gNq3UXnUFmknowfL2mEOiJ5mcHgzjBKK/nEpX6fgJXTdFF3jHhcCL/pR9ENQNE
viC8Hgeg54TWdtQwLP/QPUIXsBYWzlUkta7wTk5CNn49zNZvIJqcKHpsU0Oku9+f
EdSzvtDUPn9Y9m4RbSI863l59zjPe7NqTDS7yFaU8UHpFCn07YE6ZOtgllZKpOzk
x4Xp42+X8N7N1Q/+4bzvdp2vRjFrUyJI/bnhIYJ79ENqsGfmyudFl8/qFJygYn1q
oC4vyowGRsCaxra5gxYIQvlzGrG0DBxwKoorQhTnBv98WDj330KSCFTB+n6GOlfJ
D4vM3tjY0gvq2ouQ2QUw3HKjrzq2nP7/cJG79ZBbKjX+AuVN2kNdTVKjPdRErBDl
yCvSvInIp3gCExVbQoIkdo6amqIBHmfoUjeS5bECZ0agEEW1sXBl5YCSUT7cXbj2
UfqCbvhPKOIULbeB8sZAzVYSGP4RR4mBsoX9S+8jvFIyJYLwpwxu7GPb3Zp6P5E4
CSaDSkoljKq5UEbvQvjsPCV342vBkJK4YHvA3nRjk48StY+FwEupnD2kyzXrsx7q
kutAi4++GrJ6OTkSv7+I8Kd4GlwVc+Bp4Kz1Vgkxm/ov06WJzOrrNx9c6Kqtk0XV
uT1jHw8cPIvIiNVunn17KZsXdj0VmGDd/dhlcoLSevI0ejZfeoFdjTEsjaVXVbi8
i1DI6Y8CLXo/u0axUBo/1tBI8Q40vhvSAz7amAc+rqe64sDVjNxZgCPZRRpCTh7+
vbcrQyrqtLhuFj9n/66bmEUT7YuBI8A5RlXkGUD80B8gr8HdGBneyc5OD25cA4l3
b+bt6UTUsMWZTfRkhQZWyt4hmQxAgR593INPPfMMrW7EA6B07GHMi2MVBMmKQLWU
c7YjLg0Jh2vNyCsvm4BMu3N+KAHGi19X8vwJtwUI2i3pPEtBXm2RCzeTlPQCBnMR
ath4huV+QQEUGFDBzRUvT0U5yqadkdJyHIn4cAQuBaXnrSGAk64lARHZTHVEHIly
LfnkRqlluTbH+/5C6VC+RHDSwjLDY2Om8RdV89ILxUita+t19i4KiQ4meOOJg6g0
Ubx1lokQK+bunlQmd8ALh2R77c9QS4LoNFTfUtP2vZ8MVeaEh8LofPie8QedQnQE
rlmOJ7Skf6E8vWUx6fQijNpgTy787SDkdlK9koLiltqUhSPrm7GNQ9chThqnIYDL
KQ6Di0P/MGOODylSZiVzL3QJnlHZvR8ZKQvSAVPKYDeftwvjn2fV2xm2o+1GmQww
V5+6t6l3AhGnD5/YjZfiCpXtZX3jyG4xlh2vZ2aDoyH8OaJrt9B22OBVsNF4kjae
XMkPUfeayingDx/ey0xti5vE5nXziThvHh90Xmpx9r/C8Hua/0GRX04AL4sducEx
PgDdxe6HCcfGaqtCeSeNDmhKZKZax6FyZs1VGKAntoqRONGGqbq9FlnbJz/ahz/k
zVxks0KvWHbz3L2J3d6+mSCxA7CDjzD8aDg+5DgZeb1KEKWG3Jvve/leiHMw3ARE
ztKulp22ZjRi+HATLvFMkFDddwZBVpI+KeZ7c0wkbSOFixHKKApkmXlatxuXGloV
E5TzCAUfm1TTOP7QWVEHhYW4TCIjaS6stmQWOE6EHH6LIQquXTNnOtpKdVq0Qhyz
oCDgWbb/r272SXLfQGPDgwnDjm0Td3vMbGep79VE46aZe+0eu5CySa/seGTYZEM0
tQ1OSICYhg66gBEC2NeqA7VVhdJCRmsO3Dqo8mbk2umS/hORDtGjSde4qpWSKhaR
4dgfmVRcij2ABVoe6X++BXzLKm2398vQkrcJkrQYKxS3X+wkZvJ7TURP876Po7bQ
Ogt6yK5yLdJ0b639ruq9EHQORcDPs/U/pCJdWR1haSWwk9ML3+V3xtsuB+tab1PV
rQ7yytnxo6paIJ8LbKgebRSmTu0AG9LpVb5XuTa9CbXO7D1XgFbuC0Nx2+Qag2qg
lVwFbs2M6KRjeqpzVg6nxb0D7NgmrGLrbmUSrAkm4fR9Gn0J+x7hOOinSj0iY+hr
TfYLx3kX9Qf8dkvaez8Yj9s/4FBFc72GG+lkXmQUCl+vBXjBLPVx+1uOIb92gZJV
hXnpX/fykBatBA7HcvDzJARXFIWzvHtmTlEmZ3KqzIYUaElV1kgx2ieE2MTX0T5R
uPBkSTtkoih3RzWsS6VagCmwVlHKbJjBYQazhQpSNiXr2fzbhK2ccMWwKtBDvOvl
ITG7OrQWRyookbkpxEST08MfXjnWxHQwWJHrx7hgq2nH0YwBqrwiLLOkRcYdBg0T
hUZDaCJBc3tayOO0vKP+/iuYZyo9B8BneQ9mZYxXRRN8MiR325dpKUKPLtA/1nlZ
epqeybkatOBo1m6BB1BFidIfcW4ovytubvfi3Qk9pz3tB6imkuLeTpPOZJmwaca7
R1aOVWaK8VLwQ+M7W05Z6jnBpyfRRYhjwgcz4ymhVTz9JRTIlJ5pAJZQP2OiIn45
JsxgwDt2JL3MNxkqIsMKieyeVgvpfQqcJJabIavAHXPRfWrLJj9P7bv7lNyGWIBl
FwkVWDuqeU8HqXwbv4AJy2dO6DXDFb8YZit8bkuMVuZ5bDCGcHmI0nn6KVuA5YwK
NaiL2MGuy2YU6WD/dfDDu7PXDv71lgZIyxkG1/BpgbXk7ONPv2STxXHIGBfAuyzz
8OlG8Dh76vF0+oiw3LropFJiY03C1Nj/z8iVR4OSZ4XZrIz3KhG8vnvJh87cQGeX
gM64NaBrXLMlWQL1Pq5v605S4sCFw98/BMNVYjt6feLftm0mSfTtpd1pnHmUszc8
ZBPz4Se+ZJ2GjSfMr0b4anORQfk2ThPBQZdIjtumEJ9EE1jplKzqV5SX1Uj63EdY
BloFfqM7jXMrd7wtD85dmPckXjN8HG0dDl7j80J3v8vIG+RwQ5rloW9vEsZEFmom
gV6D6HsglwqPvEafAP3ooMSVkxiJaRytWlpL0LVy7Rmm0XjeaOWcnfBh+f7mnkF7
DuEeTJYzGDksxaqINKeHAjuEMpRkrx7l871gxU020yucExwUQRSqhgvaoTNiU/p7
rZW2Wy0JgXBPK2XizbKwYBDq1AcNeomIIGyF+IXnGeaz/XkWGNDT2VPIwVkTWVcG
8tWYsHLfn/NXGGxch8bqZwFIAEEpTnJQFA3K98tCFIcq+82bBTWMBxxRb9pQCZYp
jFdxVcSuFpcwm//gUHUjf7QH5NW/+rrncV3ReWl9cknPWmfBAmXlVWn1nKQgR3NS
x2MWQdO/pqyw8NNcLA6qlmNAapjnBzbWGETxFM5bVguv9DeSaogada8N0GUNevEy
xLyf5ZagyarDUOyMuylOlQCbD58aJTGwmXVLJRtwk5WwFZlIbkIbH9naJgQMudiv
8fWop80vn2IR0aFX24RzJOS2X0saarOGNqEV/IWP7Fk6HuXi6/5ic9kIl2LbonhK
FGXexk9jkekFGcAZxINA7e5zXgYRo5sc1dp9PTPRwUwis/q3YpbYzHHLD8TQ/MzX
16Z8jNAP/PMN1lskIflS7gONsCVSCSfSRoid+nutGEY+p2BuHGwykNgNiIOSYpj6
jHbGiOpRgeAdXExKwupYycBplX1jtQW7F6eDk3DH88eanXh1WpPo+cna/GXuZfTR
UE3kXhRSA/JDbJg7D+qlL8jw+p06f0MJqCzRXXRtmArAc+pTBns1o1gU6dDxmSME
sfJLTyd8ST2VDdsCyRXRDuoWEWtonSaw5XNtM30/1twNnjFeObWHH57nvw5sFKf/
qsLdtAhOV3EF52JtHtkIm5CBbFzoSk3o+SFAoCBlObiIFGBBETTu1d4NFXJQePb1
SOWNCJsjdhNewMNHayTObERu+uMrG1lBjoXjE4tVPiqRy7rTxphHOtAkuzKXLofi
2tNqSzwaet4JYNCvj0Cb/ckiAActfGQdtZOg39xPWAH0lor3BHsJUcHZjwnkeBjc
TQZwslgvj4J+hlDN9NyljOFqMvY5ajEPxWd/WNdLTnIKN6iSLMaxm8qDNJBO3co6
k90ucutvJ0dugkmqn4Cc0JlU28krhGljMunjDvItIrC/d8v6HibUQeyXf2bDzCbd
+wVFkkOMumSdoxcDUU5uOLWpVt2LsxaTWADQNcTztJnxyFlQM2uzPko/BmjiF2Ex
ZQkaWOsZzh5KeSD1Vmgqy99Y1GVAn+LnFVQOyw/SAIQAFSpf4c7ms3gfl/7of/Cp
je+vNioW9dUnPZa24RpF2X1rWkgw9gkx9uQ40Ee4nMV8PBsWa6EuWpLNrxLYDk69
uzwaUA9Ct1XDl3mBAt3zhe3Pr2oM6F4n4Fz+kmrwdH8orU+cpYoZhDAApspDGP7K
GzbrYdsfuxM6O4Uax/4Hxt38NMGrJvCxo3ZE+28afsyvZH9N4MOYVo8DgGn5pz6j
0JXizWheCWdc0rAUutgQ5L7YSq8Z2d7J6LwOJlrFJgHJUfB5QqXCqdbLkA4E5QiS
1KzkmQmQ+kXW/t51IGXLbJj458g2ICVXHSExh2TctXA503IEreVO+u9DeAfpHTdo
+H9uh1ibwk4olwXmQLqKj0z9qMYaDLtbUQh2H5Ct55KqqYSXBN3q9smMbV4BC1BT
Beld69zVS4gVKC4MDkXJZrLuesOQ+ybeyUPmEddOEA1RwhiqbM1aFaT4+pMAI7pi
HxVxjuUDnuPba0KQxCQEbVO4hI58jpbK8vFNZZzIS56jvLrFKaQAxaqWIGynClW7
QR8bSr/JNjVJTC7Kr3i+aeDjAUmesByyxGpylD0Sd/ZQ9OU53tSU2i5fwGXGkGmH
CdP/nLYfg/CP8mQVVzhnvKM48e5/V1SWJ4WVFeoxx18gsXskFTQR/MEEnX1n05ZR
onYxeHGK8bNC22blOQBlQ3kmgMl5eDCEoxYK1dq4kjfVoKWJhYbH+GjH3MurUww8
TjfQER51I6OpwndnUL09vl+6LsT7HtLUxZb2RJJkEzuEcmueN47eMPAd4pSsFIwY
l9r7Bi5SFe7g8wlL0jX7XMwuM1+vfqJS6zMB6RGpp+CiMW+Mv6oei8DcMkvMpQxz
/m4E3Z3cPBzCIyrvnyhbubIf0+WTkmzZCg6Ikpuho9Ooaxw1F28KEbwo+RJWLj7C
Nl6cUIpxSo0mATeod1MvZTe3YG+PelSYjHzLOkhzkJcduCp3c7+gsKoYmCvWSAN3
hAVD/X/XI/ah9sxE1yCkQ48wLJf9J2w72f/4X5AWt995vsDVDzPbYKY97qQNvvx1
Zc9vejGtuZlU75ZEcXxYI4Li2156U8dV70s9kRBc8DhUCf+gCq6JbVvuXX7L886u
6zBTKD6Glczs0S3UOPk0BgLskmrgdXIbaiEov86bp/7QkkPLRJ7Mz1YvrM5jQS2m
zelfPMKb4Ac5oa0Zl8uiF7gDpNjqP91abSJcV7nkA5TOBwoSn8dmGN8k4mOtw76W
mWivk5p3NGCsCZ/vFhjZH4ai+pE8PXQfw0XHTrRoDViFb0N4mUFo2XEIH0ox8n5G
I18CewUxGLXZNl221P9Cmkww1lh3s35XgFqmwYH7l7j95NagxObI3efDYNnLzic6
wrq3t320fVurTXR0h9W1b2/c6nVLUJGh2atyNHCNmipvPY6kMiOfjACi9pxYMkDx
XC2oHrt6t+OSX+HoiBE5aX4+o7TPWuyomIG2Gd+M5ng8Ku8ofj+GMXEsv84AldS9
1Ym7/0WtbMGpkE1OwJLjadMKEZqAMJp8LHHamoI9y+9SG/Y+4pcTAHjJsGgzh1Tj
hVxtKzUvGPie66pxdQCD6iI5+4PVDBDlFi0kyKToozGlHhXlJWrvm2mV6PHWM6IN
fjY0El2jlQaLih4DpkjMocQxwfuRpaUj8s7U9y2f7LRIe6IlEJugvn7QHmSQmDKL
Pbc2ZscSNo6/waB24Sq/M7vEbxOv6SNVQ8Dl6GTR6ee0IvkrnZ7SCxeT07gownD2
06CRHtpsX6zt2suWHrS081RW9MOswe2F3MyI3bZykh+t2kfIPDyQLaImXpkLRo2k
5/rccZxzpzg2L2v8PXw+n2m/AJ2C6LkOXW3ws9ScSelTM75mTnborG/ZSZrvmNyf
uS7GpJsj21nzoSpbS0RWVoclhbGObkSS43q6bvfuVzpr48qcnSepmg+K+bNcIZct
B0qRjziSyqFLaqdxIb23Nb5p3g+liAmxlW6vwmwAPnaPeipX3FRp4irw+503sNqs
JNU1cxnvAyEN/z0cQA2SkBFSlIFwUBo6eR25Dq2IqV8EM4hVq4+Uf3KCFtzJ7qLQ
iM+egZJCgs5ZB14wgMPkj/q0eS/EjSfkllb0XJBz8HTPjnxZygT6ZFbrhNhFxJ7j
6mdYTDqZHLI2ynlrGl0Kcgq9OpR4JKAr1NSdpWRto65WjKAPz9505HDGnoRz5cup
dmJUStBzPtO4+w6wmWiSIr76WovaLVYNkA0ZihS5VcnieCtaKcBEEiKxko560UVx
OiGttW/eWH7TS8ucz07lnKbSxSfapYBvUaFis6hik2tWqRX47fvYU8wYkiCEp3mT
4f1QRJe+CFj2od7YNUKLjfrJ9a4E8SAaBjRl1HKKODJakJ0ouSMMVNe9g3h58lvG
0y/5cB4vjBvaiYlPPUcNEEgtnEXEPLJqCceNxc2pldo4dCjUdNUHKBr1lZvzlQCC
jvgrIs3Kaaz0/7dzvOetXHkRBDjudcz9hknNYPAyNlGn6B84PGqX78wlBBK1Fw2o
889qvCSvCCQEQByExUJTJw5SexHd2bD3aL5cdOWgY6+cx1eY7pJ0/xTO+KWL887p
/96nlFoo3gkbv23wQM7gwd2HtF9kqR3dUO6NAOr/kQ2OX+Dk08OAMPYAnH661unk
XU1Rw5ng1CByS/FilfH07c1BZCoNeojCMfTw43b8rarBW11Lq+aTdBJBmNCoiNcW
XZiQshEZ3hNdsgCZbrbIArGNj0vLwtQaEnoBUrE7maewuEskMfxA7VvRqbi0Cr4n
yxz4jtbeJyXGe/rwh+R1scY4X9VONefVn7dpnWTeu6QHyBUTgwV+uJdkUWo9Rfcy
U5JS9L28KkBNUoztuDPKH0E9jn3fNq6avoR7hqb2gu2Jum8dOqYuWviZNOKwoDtS
KF0oxkEj8rEoyKFh7oiG2tRVrxhB10SpHbEjFshb3AdeMrSZVLIIArKSlXWEMyyq
Ctvez3RsF04vPP8BnvEZB5QRVhspg3sb4/YUyW5j9i05Mnvxfsn9SLE7qtFGgxrq
JobdDtXIlYineF05bY08k4BByLfVUlZ7zuPnLT45en/LN4hEwqtvG8euwXFEgT9n
D/Cf62c5Dn6p/kpSaCFfeGca9gHqNXD1j8TFzs6BYnZKiytNdMlvNMJ3zMhaHO0Y
C5+p7SjQnijcKeh/2zv/gaUuYastsIObmSVmwklKOdgUxsFnGUD+EfLLCWcv1sVP
OoMh0A4GMwJsGpUD5b3FCOZXWWVB1cVW7QnxZUD4SnhC7NFxisCXrLZe07BeQ7lP
irpkEuPLxR6byLjy5Cqp+civ4G975dRURGNmmFehMgJYqc4x03fXLvCON4vDISLS
1gy+biU7vGZX/TPdB0ZyI5HnIILjsjDpyiKQ8An6zMAFxrhB3syojqC8nuDJR6nZ
xmU4Cd9zU9ZcfIoRhWbGLlZjScGltu+oFl2JdY9CIANeJTLNjdZ+8s6mwsXFbRes
i9BVcVCuepwe/D8d4TlzXqOAU/gAlL3w/m5JD+LVyPu6FkqRx2R9+jI/1HNNveoZ
9e29kbC09HaUxVdYOLqqNXzdP+o9ydd5OfRjTsTzvXUngz/vUFkyCUzviejuhHxq
zvSKeta5kH5Yk502VG5JqMw/nOMd8MQNHqhahEsuiDwRh9Y6MQt2MRUYIDMewzb5
Zt048Ed07aCl9MvJ8zqMNXc+S4BOXk1F0I54pU6MdeHwXlVMR6Pf75YhzHNONVam
f2a8RJmMGn8wa8SCoIJcgQSa17wjGG4rZ7beeww+iXyfc1GN308uJCifc1N0nmNM
iwIBgMVl+V2OqdZr4pCo3oCjh88NBnVg1BGnml1sYaZFJEflQPSxVusw56b3AJOg
Yy91+hsA3ZkX+konVq7evfOWF0662DCe7jCh1SPKCLzht4KI2Cwz6OxPkufYr8Ca
GU3iALNtLPfX3rS7HwK4egrXaJeTJAAcCkuJYLKa0BOJSvvMrt1JU5U3J27jQqsN
bBwljeMWFgQyXRrpztLcNWaSrmTbeW7aoDt3H+opHpyDpHi+tWREd8qJiFnoHMzZ
hr/hHMCFt0DPSkWBgxMy2N0xxM9ziBappaInNq6eBzNVaYIt0VylRdQV9J0/oTHu
I7/ZLUT3R/0e5I2DxybCS+6h+yzvK97HdlGuyi/1o1MArKeSwjMwrDAbCnjgWkMK
FHM+uHBHWTwo0yv/MKe8I/MAnInlr+kuZ/+tXa+0kfXjf0QLqStJNO1ChLr/b0UR
zWclVeAy++/4wPMtKE17Ia3vuR+QQSB6cjxlAqaNnvQKRWLn3xrZXJak4n0K1aLy
gjYQ4XrXdNZrxvZKEbN6wXrgIjD298MbdUCDetsEk8Khpjn2oLbWKOYOpETw3BRf
YY2UNEYN52aBcOd5fJlDEbd+CBvbWIp6fFtXiXLrK6Qt7podli+SoE9NlS1YgX4T
Yf/mYOe31vq3BR2Ll4i/zLujEasOdttp4hOkyXRaagZiiwanfcmvReJeZ8DUVtOG
RkrpKiupW180f6b800XNen6gVAvvGZRGcLTngu8nf2SoNrXjgRV6jaPJMw8Cq9g4
9LlgW5LY+bC9R2QTfsYPfGczvUzhSKkLV4ywwoUz3tlOoWMwpQKMrpe5PB4sV1V1
7UXmyOK2JROsu1vBT1wpGpzLbZP4lmqkYgxFfsreaNXxe5F7NEiXGaFVu6FhZf2M
Lhxy5CPzliinYNnbwhrkSkm1pN8egho33JXhE7ceoTs/CFeeolo8IjD9dEO8y/Zb
T3jRbW0rHlWSEmL0YqeGqLCcsib651wQHY7Iwy01pbM0tIFgA+vB13TNam+flaxb
ZLzWwT8ScxXRfemP4gR4Z0pIP1uVsc9ABSvGrSZxfzC+TSPArPk7t6tz6I9AuMqX
sIe4A5MOEGLV+nPE9p4dcHd8RmyNB0CdqoDh3Nv7xyeUL+GZD9SNcWW2ElWqaNk9
wZ14NnQCFr9tWI8YwYK+6HxACEUKXs0ENCvRigLsil/O7rbRevDamF0IWxhURPjP
2yJ46HD7OdG3/TJ7opmTrpt2UsN0RoO1Oge9452yyqxUJhHM/sSQIpeurcDi+TCX
blzHFEsd5IoL9viOsndlQZYAdWiadNdmdJrHqxbh4BSOfG4XwCuCy60EgZVCZ1x9
x4iNOMrIOzcPgRBP8k8k8W7xVF4j0ZB0fM8FTF5IsDWAW6zx96jOMT4o9e1jYu/X
9eg45yJPk6AMGVBj4txKahXCBBTeHePES/Ej7ZJL0p0hm9wIPIqHHSb1t5BNuS5+
JTxzwiYFpJNHjiqJHr5hidq8+h25gGryGvaEltUa3zdagAKsnAKtj2WIikpMeUhr
eveT85pcmDUAUCnStRCUq3bLMGliblKr1j/+XOy+731TkwxOsCQCkJBfbEWxu7K5
bNcIStYto6yOfSuTZbUFcL1PIfyIjdQwSqtWwM9TbITaqlyMRq1IeZZoUQdPt53r
viNqRssO/C4cgMOhL/SWtgxSVmkDuiOlHszDeBoHjc3S02RYhNg+ItdN8cKrwQm+
ACm6vHEJv9X/40Xz/BGOT0kYl27HvJwQbMaG+CuzgQf5+K61/VoYrMpXMtJ1ixgu
n77802IWQSHlmhut6d/ZgwXfhYLH5x1TN7DJRm5Q4MJ6aFl0qLtHf1cRaiLYgcnq
kWoYyFtcj3fo5Zad3PvjI6dGfaXpr7uEsAmIDv4cs+yov94ay0iw/SF6sJV8RQo3
K6gr1gbM6TCwZefxzwqZT0T5ySvvZm/jAIAmXrp+0UdJokoZMRWcJjeA2hsVazSe
G+AvXMZBvryPs4RBqFhPJOgQ0nL5uqms9tIjDD0U9nO/nb1zI0vzMXHmSDmtMR7K
qq+blePJMu9xo2djRd+r8ifVbWXG2GpQ0U273kqWX1G5+SbxR3kne2YDFsmsgEdt
Vc2yhpOzP8xFPfO47LWzezFyDFIGUCFkGMAj2aAAkZSizRSRojnKFLySQDEewVJa
GEr01mp+j4IiolT3lEJZEgraNfwN2AMT7jVccE/XHyN9RFAveT5tQapernAkMdcI
wyk31gdeEd+zu95e06kDlcqDo/JocmgWU0F/sUWaJcj707Dt+gCInuJEVNb0BpyW
ngbRjIW/Qx8pI/cjrbZH9QwqZDVWvQyZ5zfFyBD4R8wBMaS830ZSk7fWfmq17obh
IyJRxVWwK05HiRTyr7q/AjC9o2Q5+m22zTU5choYjVR0AsLb6bgoygv/T/xzJmxr
62FYzSbHvKTCwyh/KQvuBqDH7O++ZEiv+BHYgQ2t+Ft5/shuV1bcJCrOFWxuDuXO
TOHttGRQ7WqVkQW9wcmyG7jVG4HRrLcWZVg4kZ17deyExp4r0qxGGCJyixc4nB0d
jJltomWIr5zzCTn6aQsuI5N+tIZSTcv41SAqw3oOHOM5CAcapSVXiRIlvJ6mtH91
0erbXaMFekTNb/sidq6SHhY2JBSgOYh1XILtXiD59MhABXA0QZIxmt/BaDvV28GC
VqteykmkZmc3jLZv+teTspazpKYBpFG0qVhaXRrjYxMKOCnCaZu261oThdSz0Jzs
++qE393aLS0fsEqo6rGi6MGM+iLVvnuL6hyHDsmrStdFKcIYT1Q0DcVoJlQCkB+f
LXF0LRpB6RB/BWPqo7nLH0qMmgFnDQgfBxt7T12LJVx9tLyb5uFE3XLZdZMH6GLP
d7MyV+C2WKMKdOSvhaILhUqsaGuy0Ukn9jxsFWcspFmPFVtw9hQPvmJp4Gr4agnM
9HMJHPzUXVEPg4fmwJRCMoGRev7kXtJ4r8VRfv4QLmDXKeFVXJ5ACmZrVsqr1ChL
Fifm1NPEILr6vs7ZICdbl4Ee2cEisds63SGZywp2oKkjK1minsEBtVhysHq6Bon4
sdrV0QQ0wP07Aw6pDDcOzxDtezt0qmuiyd5VmW94tj+yW1rxoRXDn3nwyVHstzcA
inbIBK7kJgtH8Tj2B8A+gWrWN0fcM/fBwaFOG1/Li3OoZQfFW7S+FXtrHV6Fr7AA
O/tI3ArZAsloSEy3spvToM2DE07Td8DeINlw6DtnVfg0ILI1f65DlQjt2hk6SmM8
kgBBZPsDkQ6TR64e5IvsblHLlSj5i23PAq38RhPRi0BsW7fD8KnpwJVB5c+2w8uB
4cZpPsAr858vDs2pa2S640346kfP2QKciapmVvbgwh0moqVfBa8FFpURUk8qvHnW
+A/MgaDiIWKjIe8DXwmsfImKkmcY3Qynx+YX/+wfPaUuLrQvboZB4zrDEM0pfGvp
JgIu4V+8JWL5gtl9VNM+Xw8ZVr3APU37UGpvhQ8TLV0p8iWmV5y+ZpKd/ZyaVzef
leM5RsBt5RPDRPwKVHtl2n1OjI/UAuE3AAxAF7yR5jPzuZNmMpC45mUv9vnaPwi4
Vl1qPmIa4Len2yuFnh23W84RKmtwB0+29hHWmdAT7in16ttqGUr/BxgQIwBLxsPl
MLRE1a8VT1cB/Ag7ClWwGD8zdfQtKTBsZQNHgl5LMsPfmcbtiwwDugtHGytl+R6Q
qS/GjDH2YtBn01PDTIrzcMTwwEM/0rfYXgYTd/0D9COF4YLljkiS5WGlxg1N9bET
xvGqP53X/pO5KZk+YdeowZ0l5WHiNZXVbCC11Fd489WrGi94XylwjOmBRjHIWovs
85SZK45slxD+QrVATX8KMWzNm2fpW8W4IfwmLiaDIATmcEyk1SBsIFkCc86HMlcp
deb4tPIQ63yNBTFtKkbFwI1Sfbc1u0qLRNrcq0MOEySQUe++L92Qnr1Dx3/O32oT
J7V939eQRqniANbMOBlzuEp1bKA+vj5EMGhjQ+esJ5UNP4l10SCOis8+YZDQOucI
uan61Vbi+SEIW8EVp6R65BdVoo12nA2DOCbYl2oSOjm5vmYFL5jLAyBucQWcn2v0
3zqRM1hH7wC1xPExe5E0W13VAQc/nZmn/ibpdr4+2vxdGEhhB7jGhYFBVZGRKVof
Kl1VtFeH8k61Lfh4ZwMbhE7z9X9NukY8v3L2OY4BqyICsLUpxMn8SrliiINKSEad
cnBtr9hq3kf829RrWHmmXiy0zzrPupGi839hpcGBD9Bxn5UqNK5PRFWFVk9tTeDx
glVSVi4dNlHeP/2npVZAxGOD+039bLfwNkCOOOK3S+YgHDuNCjOWK/Ie3OHrceZJ
fieKnHNtUoMTAkgUUKHpcEUmlKZ0v1j6czTB5cHafuQ9C+OWIglCzoB9aReE80AF
/n+Il36J4kUSv1Gh3ljNennz0C84nKGVQnt/9C1JlazDhh9sn4dnE6AseLz8VxWw
LQjXt8a4VsmVcy7zdGCwo40l5+SxxTNaHDkfg5+r8/7Q4Alwo6i6ywuo5ibpVBkh
waTsk8m9tYIzlqkTBkmNW0Z1Hv8t4oJzS5x9zLnBZF5RssGjiRxrZctO23ytv4ZH
2hHuqNdon4Y9deGJNNokMb2mPngOAwI4Yq3OjH/0JvWGnmphE9pdfX+Ja2AuWl56
M18VHid7TOXR9NfeLHLe/Yz09Hm8Fkom2whDqP2ZufeKW18G4TQh0dnisyHgfTJm
AhnUd4EKyd4AIQMwxxBm3Hwrfg2dvTYI0SAM+khBfV29OXKylSBBG66Ie1xoyzBP
/ZHvv03uH28x3j/3BZZCfjYkhS9myx2V1kiuFQwkXV0j22IY0RmiiS6BnikhYUQn
Av5cPGqQ8TXJ98mSNgiefDBXJ422eeojWwFhXwE+03PaC3tk059UmpnVRkYIpRHA
5t9sFGq+i+neHA89zn15K+ctYFhjftXCKkET65UCpbha+jdsKX8nr9dWHXM7a1aQ
6UVgkuNS6AC4vTyAXh/eD/aWZRXwLGzMv5sqARwVG3eHI2JQx2Jxx+DxTumTRZCF
FGqx++7VXLGj6PPumDxpUGlAdETojF4GtfqhzDH1O6U1la8dCrjfHtzlsvI1GiMQ
Uu8E4LT5zhneCTEobvVoMfGnwuLjEatB5FsMxo1Dijby+ClIhvietuxuUwyweC/e
YQv8SUP7RxJ6FyL0L6xlVv9WxM0ywnc+lrUALgLiOSx7tFSUsjw4+EVFL5Pyq8sd
afOgBE0Anx9q1ADs8bv9dwoR1MQscNQoPhrF04s8c/H0C+NBUajgO94b5E2j1Hy1
1HdYQX1ToDWk07upRP2rAew3xqC/8mfAbRUbiwjUQrh5hXBifsB4u2qBafybj4oH
76ckZ+X71b5koqSLM9KyMnDT0gTwCvRvp4St35u/omMT0gi9jUEF2A2uj17oOj+b
biOpm92JrVngbQZPWFtToX7bE2ZAjxKOqgkvgSLXm7EmO2EPyhhgtc1Wm8R/CNyh
tE1IBwBGenHVN9SS6+D0yHG6y7FX+FvqZJwZashukIF2KK60/R6hMUQ4rNZGXpm5
2zakwvvxhE82/6ixHRlerc3hhEPy+Ra6YkLgcOJrSijvxtFLP1d0i38+xvsN1+xk
BlmO7MQ6nWQEoCWKY5DwIWtMu2sFgBvbh3JMNfPfb+XBjzJa6romNLKpewmkNLIn
5pr83uaEk+CTWDmOuPC3d+5rABzGQRMIn2x693n/FOfAwJI2Q05jGGMC5Ww3uczW
od7JmOXofgsH6H4esayMt/tAlgMJiJ3gvoydKh8eELgoToQNR/ceQe6r6UfEnA9L
D3i8hEMChTYvuOSGTDWXg+ItFuszMVebukW/muG8x38+exQ7IWA+Bd+rjhWTsLkW
Il+38mK2OVoclT+wDLHH7wd1lnM28ZwDLTYykhLG18E9XekJkxBViQ7njSwEmjjR
5uWPh9EJ688ijpoTD9gLewPBow2ROXTNblnNj/dhyK8FKLt+JqN9ZuVCXLNP2hH0
OmBoRWONZ+yayPqinF0gq7f5HLiaKE1D9xrkK0pwPTzW4h3Nq410Ii6u8HMHZaFL
sb9EV29CweA5bGo675q/92WKg45aX89Om4CqWICTvQcbZuASrRh0VMKqM/BVssW/
ZgxAQBNj4r5pkxESb4fFpNrtZBhxJip77kfTJMu3L3wa8AtkOsLSVnyLgB8Tnfy3
H23OG3N7H/Ie1QhRlCeje+me8plhBXiKs1wukFT0RM27W11EDvhpIG5T1KCWLaen
6oo6vajhH21JkIlxIPq6U+FCtGXhDdiQroZnIIF1XTVQYV9U0cvHLSzjNOgZKEuA
sNCu+SBfjereaP3Jzx8zyJRFNRW78PckmVjQfGL6ow191HvxX5wvUAl7Zi+O6z/I
yyWWc+olX7ChP/Q77J235fYCzWpwVzuoIfWuFaXeoJhbK4No0KbmFURugHhjM9Kn
XoKxKgDZ/Jywpbj8fS/45heHLbQhXMkswZE2qaxEO/GQsyjc8jfqLUaC2zywYYbq
VSBgyAEVrpnANJ6vQy60Yu49xc6XmAICi3kEfA7a7BP+uaN6ObdfM/wvFsJjsNEf
n3U58oP7y1nVagJC388gBE2xxFH4kjY0ZG98+EZMjNxji9VS3dlJaG4KWOtMF66Q
Zkt/ikJnb73bMFhF9cz5IOkoKZLOLzqcmmLdH7hZlr9oQ1kt7sBEiS93zIkRwLAQ
9HZgwuS/wktiRHkGxiX+4WUMMPgcNUx3pRTvXFZ//JuGnxa68PNehZQNr0klTRr2
5Hc+QTcElhud2vWBxgPKXnvyXUjJtweYJrOfF6GwLpwnqZnN7Yi1AOhKD1nRGW2u
eHhoIySeTRq9RAbYNLlXs9m45Dce+nzwF2YVP6FqUNjwySwFnmcWlavsoV+wcCFc
RjEnU24Fe3fi0Cb8uFeLaLG4p/FIGXSc/oXg1u4vVHlk1B229E/brnAkPNiZVTRG
RNEuMMGJfnLim5ilBQ8ixQ8M0X1U0lRt8yKsBIP4nngosG22r4jjXk6RUDxNzi+n
vaCJHYmt/vFdBqblLGdllg5seS5KbseIPqYfAA55ymQl7R/dCEWYmZY2vbFJiFt8
7m+22VFVuf5h67S3yF+OIhOf8SvDgYTpMuov5L9VTmqwtFIBrUyVLj3haeCQeABD
kh6rh8/fR+K03bH4ukZQvzgHyxuTBMLjATx8DX1Bzql3MWuE8vY85AZfLNjTW5lS
en2+AbDHYBo+C/pgJ9jA69COBk2a9CJscGzX8Mn7ztqJivFI2gT8xFtTKD9LMMRb
ooddBEV/2u3DgmRRjL0VQr+lOfv8HwCQTIBxRJ+YFtLE4+uO1agZggA+MLBdifAS
eHuTdavbz2iC9QxgvaSHrKxw2AVHfTLygPVvPaahHQ7L8dy0w1fqprb49SXFtNqA
dEDrIqJJtwHGYLV0KzYwCoAe1ETF60Flh0PyT1oJe5zqDgS/us96v21FTSoanQ1G
bYogYIY796YQPyOkrrIAaVhvQ17mH7GKjkkj2+qQqMcL5R2SKHvgDojhVlGTcWJw
6gM7Gm8ZF9hwLIRUc1palKHnrVpdwJCXWscXaSGcbLILKL57Aj3NpyvT+NicMCX9
k+uNEfKqElLA6MRj0Acl9mc5AsJceccT9+g7rJ3pXMHUxYImtC5xqzGgJxtvg7Oy
PA2D9U2T3ZCmthLlDlZ9BPh7zgcyhOivRythncqAcC1V3Dq7AbIvEN+1iO8gRggw
8Bv18K9rF7qxdYqutHSbA1UpjEDHMMb9V45pPF9LboC0xN33+73D5WGrS8OFF7Up
g/efv+sD4Qt2kFu0FIQavpL2Ueba11yZLEoZgmCEYKvr56RAio/1EP5Beqj+EqPc
e4ZxpftAFKaV6iBe0sVH94NgcIqIUYoA2sRniyLjzLLZUMI8Jq0Wa+SFGGANfClF
p3IFQWVnlSsiGNGpILCYpz/FRa/huvmZyCPqLoXRK17AF5luBpE9nd7caid8Wa6+
6KOjB6z1mwvgiLf4x0L8uFRDgWn5AZ2h0RNF2Y6P4dQS3h9relDRFWJoljGHxddk
HpCuyy+tzfEYwiFKhVmVMIXZsd+gDzyqnCfUEXwgooAggY5PRzpj6bb5zMu0RtFv
jIxR5ggdjVKMFpLpvKexqfhlD5xTuYnfnMpFJLyY+b+GmxL8QgIsqoJLlL1BfXxQ
GxvFQlGDjCs3j0L+fVzYNqm0ZxgUvyg/AiU4CYRUJDIVzS7fZ5twSjd5rc0G2/Zv
Ayqpvae1MwFQZ1mgP5nlStrwzciVf6UUd5hz/6MNRZWVBSCXbRCf8VshUr6Efd9i
+b4XFHoRtu2GYMYs74s632mD7wCE2AcLb4vcpA5s4zXnmiWgeg5W0F3Uve9/8Uf1
qBd1Z+PnKZ2gl3Dt9/9O1Jzo2q/g+xqCWYgp8msAgI+FFjeJas4fK8rRoy8TyNNJ
y11lllqMSuddv3sYeSE6ZGYjcp9VT5kxYH0t7n/O/Halw703h45hnw7PbbtzlokV
0Xz9cgdzH3CSqJM4zJS15fcjv3sN8SCsbygk9NtJrADQT+1pVKpfBkJMYhOTfrVY
PzkWVk1LGfUIATTqNdWmPpdJTWI+xIS8AxnkJtxaUhMr35hAUAT9qlgxTOFhF2tG
svBK9F3+IS0R5l2lBvt9qhOv4ucnAiB7vwim0epYrD+SPy8lCPECLTlyZu/dpQdV
cRyIk3vz776MxB1RukvqNYSDhboqefOOWQiyLpWU31dQEGitHhRBdUkAvHWb49hA
nahSyGO67SOAkrQigFe5I1/gabohLwHuyXn9yrRyOdbYjhEg5Y5mYpn8QnwgCC0D
wASzLNZaxyyJMvLm9xTRrW/gxgwRWF19uLQPG3Dej094LW7y1O0tUnytySnyLq28
M8bgmIXKeWIN5VZtKDYNRWgXMif5GfZcOZmPe6iYdACuM1HBLfQqw/S/rKc4ByFu
IhpzMp4FRfdxwuYnDotPP5Q2vmtMHKnD889Ki6zXDVrGkEsDWEQFhD/9YFgpi11n
4hl9ycIH8KWIaqS+zA9XSeoK8WDae7wY9i22TI7ekNPemSqN63toel6Av/vvZG2B
wYf+5Fm9lqtaZi2PGVZKVcXgeslrC+M1LkDo4iExrCKpX2hy3r9b0uAzCtPE7BKm
k9O1lMBrnpOZx26O3F0RaOPRz55yX6HTZgHXULLXXs58J8ByfMzb0OnytMI2UvBZ
p3iPBa7VuQg1R8Whhxt7crRrk8TcsHbv2CAx8vcZRcW48vrhPKwOuy8LPijWH76S
Zn8zdWzWut/Bu1yvgGGKZP/5QM5tQksnnPezfUpSJhED3qsJR+AzWpYCvrOyEmnI
BUwE4fke6sG1MecYf0ZmYMLzchdQe99sJ66vfJ4TdBSZs0PupKW773V5273OKZet
S3BsIKk6QK6xx7Qi/KHkjadvNNLL6C5XUIGkYV/DUbdMvK1tjMJ9fjf82ES5M2kX
70065ytM8Iy8AdUywby2mF5Mf6GbzcQMCB492/5/2dwMQfKInm5clBVt+VXt2A07
rOZTb8kWkzfprLr9ABdxGtiD3Yof3DzfbOKBzbZ/p88my4J5F2BKZsRDHWaZphRy
258EOluuAs48Y42lBnB0uK917m//t7PvVkuR7jNDpFKJkEIRNm+4wSX5r6gfMxXm
JyL7VoKJkoRkqokweUGEfwR06uGGPxTq7a4sWLaLVfkIqL5civm5s38oght19biF
+e2t9IPsdVO96AtU+Splaw4dpQXkSRuvc8ddYUwMVb5lttNdwgtlOIafZ2yEyUPn
msDBGG2ZCG7l5TjynBhzyPklP/4y7k20UdHP6p5gx9Nn3tX38wZ7qdBXRfdNaw5I
V2hlXlslZ/PgwrTbsyWMLJqVqKWW4jjn9kFYS35OywCx91E0EWfBXqntz7r9H/7V
LSSZDBfMei0Xc6GLXXwo8SfmY5GmIzwbpnwNBXAcIEaYgimEWFHy+2Q7NJIKlpmu
lndoZnnOIml03s5f6WhaeGiIMx5fLWCV8ZrvGeJbjJoI/FBAFAUm59EH9XnfyH6d
CeG5jAzzUpC7Yxz+DlBhecX3oUTl1FJGbdYupZsZmBLcijuH7ssldAcfuaIei2Go
B5X4RwEhjosJ1iTV07b4/PV2n4adZAS1crAgGesu68xrveZrnqP2yQCHnhLBAcCS
XZ6s8xU8TB1wSRBXxJRczGu32KveBo++lGy2Uo5e0P5Qx+NgQb4AhnKOzYqEFtx5
QvmuDFh1By6fQtGmrGcgga21FiCI/5P7bfdITJ5xf2J78jJ7wxh6R8hGnt3Xl00L
wiofpmtUvtuid+2G8Lg+yCEG9EB0Dd3Eb7dt9cHjAVbb2qlnQrcq2tWSnJNecst1
74HyvCTjZa04iXtzEnT49A2K8qSCtZya+OYYnyitzMRETdjaVDWvH350jqDRIidM
RrG9aLBdhPFMd1Y5MHhJJOpZD0ND8q2Ms58tsp7HZ4S80vHg/GeVPSVzxrD2z9D6
V/V6khFm944GTtSnDMUxzakFfD9urd/+Z7HiZHLx4pJ4DmTOyStztkjBhMJEFSDJ
3QZl+QSpGFq48O6xKWPtBflMnd0S4L9s4omT0kiFYivBl9sJZFvMcjyg+d9DMw0I
y0DVzDWa5hIZ1fezKpD2DRzOZddU3i2V/Td/M/u9Q9/jpOKg5Mz1bNp9dBCtxD9X
x43/B3cdaU8fCeGNmoKgvThns7qrnZiz/Hj4ycBWYiWg1LuSp9WtuU5GwcoGlHjS
Z+iAvVgopHoMboCYeL/qlyPUQfCrV0PEoGnGjB1TpyPrm0cOa5XhX/fgq0DlZ8od
PNHP3DjOV3ulu5swd5sCL4QcPkSbo7ZXWqwyvz46anFMuZO5DpfZTagy0t7dTkjK
uvxnDuh2AjhKHV3BsY4HYiFfRQb4DP+dSnlIdFcnSxrHB1WjyGxbdxFr5iGcHn7k
zTWZSslh1NanKmHpF3Ih0JsugdyvDRHDJLVwo5o/IeHNR0rwjjTU1SqDT7kh3owU
765/DfHry83nLIKaT1Y9qmQ0weZd2VuRvoHa0DCnYWSbo7VX9qIa4QsU8jSlii+J
SC5mQTOxz/u7L/cjXRpsBG8oE3hVI1tTRI1x3fQsbThRK9s6A1EkamvPlPpzPV1B
+Hiw0RAv5bl0+z1SEaYLQeZDAnurPN/wOH3eB5fl+Rg8AWejz35vJd+dORqPfka+
AbUQez2HcTtj+OeSopebDuzT/hoShSeFenh3PQnIdUVDXGXfo0l9QDb+dGAT9haE
M7wjr9SXH+6xfFsiYz9XtGRb1ePl+SKJ1CxlNHythvQMNgrbyBzTyKASfuCyHpbb
p79mUWGIjpzshho7I5QUzHNHN+79PHT9Dxjum66SbTKMg8nc4PmVdj2/S0dNmFdg
TXmXwaUAUbPzvnPZ5FwVI+ckmvoscApmcsYRuttwxIpx+3szWYr4TQn2SCSK/DFQ
AhVMQ9Z/QcMTSMOMRsioEW/oljPpbHURVec7cFQb4SrERMPEPOQtBxLOmg4EmVcB
dkw4fBS4Zuv/zumCr5d6aMnV0n97CXrxFeq5AzjuUmDYg98jfrPF6f/eQ6Y0tWZa
Kbm+VtExxQySCBj74sQVEieM2v7LN79YdUwxBWfjxHB+sZcGtJRrtquQGR9vdAJc
iKTfd+nTugC1qxIlpkJxgQaVEkRtUW1P3S8bgTDYtfnIjT+9hwJSRO92xcVc5BAh
X3Wh3YbQa8KHTovQwhIUwAWR+Zs2vsj5tdJSApgpvE25GuWqQsCoEpDLyxtcsfuM
boVRDmXIqSuTGlUsBlfT5imI5Co3PY5ZDjJu+Gw85m02mtvG9nAvxB04A0h5S80J
TBuA0TRgqXeGtXDCA4wnACz2PNMePysb9MPukDknSdltIltbsybpXhV+y5Tx5QmC
D66wyHaO90igLYehKJSgvGE5ZX+rLp54dsqhARt7HeK2mL9+JKiZ2Y486BydBomQ
4XQkzPN3r4Px1/bIy9JEmEhvC6gPBGjPT+yDUE5b2EURjDw7p/Ox8JbHmfFF83tz
S+hUBSFS38MZhUu8BGo+6itoXlYdY3qhCBOi+8/L2+Rt62l+1nR5QpXvlPpPfjw0
iGmTvudJMoPG3RV84f8NOTjiCk0VdO5IKykBszfmCr8pDRoBwJHtQwv1vMGbYy/p
kAGod34JRB0Q/4CovnbrbSmKeA/F0pB28RzHj7AcmlhL8g8L3tCOe6LtDpZmKtoH
GI1VjtIDYLBWwrRBeKmZiLk6hN5yPvAyo1CJJS1DB2zT/HY7SRk86QTJg/PThrlI
lg2Q7cNEFY0Zo6afFrusOoy4qfiKRpV0W0x/oY4xtP3RX4SgHF8MX8vFKBgeKNS4
atEk6u79OidDN6iARANQ7zDSG61lNprYqUu/NdjKtHJtkCycUFw4o834YpOT0L24
0PanE6PsqPnrFklfyAHV0fgWGUeD0/xtglZGyy2x6FdzF1RbVnGalmYblBtWq7xk
71jKoXbEtng6U8Ht2AjCbcsA7XiLBf6x21I+HOSEvazoTgG5lQE+Pr7RPtll39IJ
t452NxZbQnVpn8VgHXETqJqGPP2t8o0QZqT07Oz8tGGgwteccEsKXvANqLs3oXGo
96JyiDcrBs29jrVdEUSMMjtTM0azOPzDOre2wLI3dRA7l2dvPBBNiha8HADmyjTk
fbd2Hdx2kB8Q7X8GPrPXBh2GdXk+9nUwLLGSk+RCtWHsyKO8fAVS+s78L8NJknwD
yGqOKZucYCgq7YabjrXEcQmRJ58IMqoSA4R4buVJZYZ7bcTWsoPXtaoUbwL5WbYj
czWIa1Fw9JKVVJsGIm0PY4DwZaViawF7tpBW+DkthxyqaoIT6JsCL3ooB4fTo8p2
TkfWNV2RniyvUyCwtySM16TyUYuIQ1XDBJTSxHnGTIq6LUiKo8NFWrC+d35hDj3y
4GSW/pptzqrjcCQK8bBaBe6ZdCfCvSXEzdX9ijN9AuO8dJsmYlOgTMYN/5boSytp
BHvPh2ErwL+E2SPYP77ABaFylL0CE0OMpbGba62a3kQcS1KwbwphRbhzbYC1NkPO
1GeDon0EWlnlMIEAvi5c/meGO3e4vju0xCsKdfk1oo/r0klJt0Iz7PLIerY3s3Uu
y4ljVZ14O6ke8CFfW9O9XLDs53CoucRVO4ulonQWgMnwrVAMjqCFg5eIO4JCsNNU
Wp37JmxN6NefwCnV/3CE51LUut5275czewJ4Cujm4kIR+mNFOEqhDdWaCY5OlJd7
7YtllAyGNaVRRr8Sw7EQgq1SKQM8sZLR9bHrUwK7H3lFSs7Dcyy1oTlY8ruBrDdR
kqV9LjVIBUlzsiSXF09lbLie5kDn2zfFkeFZkJNOXrs0W4OfW7MeqZH7BwiKliCm
D6aD3aeq3AwpIURYcDv7iyTCscVPHQiBcpH2nxIyYtbmLD/0ZM894IuV1EpH3GSh
AwVV107LwfpgKab1MOMOOQSAH+oqGhwVOvbAEou+PFYNvB8ebz0gKsD9WoiboBj0
t5/pVVyEPlU2lr7TPmuob/Sn3myDIjeC2hr+WRkP68HH3twKRYz02/oB9HwSja5S
HYgdODQORMmUk7wDOd4QNM+3y9gn0oIZa8PMAFHiA6TWaAadiX2qdhJNGIS8dstb
7JaynqjrBCqOtdmEisIMpHefeJI2vbhDiNTJhvDzqnoQE6vg7d7tzMg+dU9k1YNs
6epEQznDhXdVdZJMEgssZ/p6eQoLxM8oOxNSjy6W2xDlKVXt3NbMj2mDSGRnpgtd
4/vHH+j4RJt2vR10YETJhBO5YY91+KssL9gAomn72qjSJAehEc3aEK2rxXpw3rjM
s0G3RvamsB6IiRiqvEkG8jtGd8N4e0dD3JTKhpnZDxC2m8WATEz1KMnGoQOLUUIO
Wkq9rWeEMNlEATqRVqwLlV+NGAfpc08CweVdx2bOvH8YDlPL7ZhP/q3qc7UKDqXT
pWioDmCx5fwi66lZYySEd5YQfJvYsme7tOmI0NEyaa7jhvTRbPISxjK7wnhpeLxQ
KpKIm4iHfTrcWyES0qurHkE1f4BWbEfdlJvt8izt9LeSssrHKdj97zk77BzqKd5y
Pl9jphvMD9TPIWzMf8bW8JF+3Blk1PmMiUfOEehJSSGmsMWMh/EUvvycJduOG75J
YxCi9ZRxUDLuRD/th6IsRdpzcko7c1NCuI4Q4ZwM9ouLA3NgvJ72bSdM5XjAjdPG
LcEwonotpneo2GChECdmYrOqITT7uB5PVXpljGAKgpvfaZrxUNh4giwZfWXMwc51
roScHPib2GwRLvmBUVrH4vBFFfzJnWK2T+j5nqCWjRdl2bi6bb74sOpRK5693AFu
STdzPJLB6Hpog2NJFKMyAo71jYNPPtKz2SEhVlsH9gIZGX3KlsbEGN75mBrUREpH
Rpi/bidIRYNVibVCcC62yDR+9KpW72P+jd5XYNeKdirqQNdhwDPcI0/BACmrBzLs
HvpXMHBuDLO5aoziMCvoh8CfwsWOKBfajXD0DLVP0FSPeJhNJZT5vRwntoPwLTGO
c1r4aCXwJ9slzVHI6Qnq7J4P6LWCbG809leG5kBoqfOFdy/xlnYe1DSKTjItZMPr
AMSk/uxtDyAITq9f30QfbGuQyWwAQLVeIXWuCMrmMDTrR5wGLeaCMBqgpQ47FDda
TFpKXNC/eG9Ym9Y7DaojNYgPyvEUcnhtYL5LoyEuj6l8i4qhVaJZ6ttbIdcMJYbz
iY/r33QLVTDi1l+cXvjw2P//QaT+X0N37NFWnGyZmty6F+BZZNGRzB0k0UHh68Xt
0iPaA5305DyfwAy4kwSPDB8odhRgpBtvhUowT6HSPLIz1WphaEESDjiDiENJzDKZ
DsHkMBz2R81R7qKSCbIJHNCzAfc/LmZHA3dZdK1gZg1mihHIoy9B9ANNIxDq0Mka
Ll84tHMiu4X7is7tFRf1ZKWjhmkJ2qx2oCq2feP9verj5drVHuhh3CcD4c0mxnU6
Yw7Me+uNnIsKnXuk13dfZdmuornkh0X3W7e4lpVaWq6PvwYDtW2Ha4zum/gAQlQq
WdwFUvzfbBf72T/sR+gByKp/9/fQPiGTJewqIFfXI3lwg/2LzJ0AZdf04cw8ddJH
Xz6JMeM/3MZ/qnWRe58yskSxTgHnu08q0YMJ5bVQkDSXYhBF3UCze/JUPlrNEWSo
xe+bQVcn4eJMtELOepA80tZtly/qf9jlfODqT1EoRwMgSQkt66ut/H3u2pGFw/qM
CK1Mq61EWS+Y83+DTi+aEgdOiZ7fiF+A5FPcobjLiUlAaXWyPIWTzxhbtzYLZ3FS
CeUiCJoB1Mnp2Ku7z1KbO73VrFu51GSSmDfWMtqbkfpj0BLBOrj3qIejdDZT7zpZ
i58Jra0iLLaTyO8wbQcrJ1BuNIATqpw7XpOq6IK/vZp5Wd0umTCfdWz2EKOUtpzP
6fHaTwWD5ISmI/LKZOmxJuqw5Bn4xAHxsDum+6TKqf30wXfMqegAF9sB9y61u07Q
Clkf8UGlEYNwFSxbLaIbk8CPhb7WjpBE7a7O9Wpm6tCDsrphEv4L8Qou1rPvwS/m
woQdMb5j0qEuk40b5rUzKg1xu5uczhZrgAq+2rCwQAuxdKvNKjg504qoQRSqWQSr
KxWz0wpgQLISf91OcZSkW1WIKoGent2CYoio9KxrA7uPZYIEjCHi9kzdDVcJ6nT9
7jYy2X+vkDLPgEU7bZox1O+i1fCaZd4W5Wuf0uszYxRzCSmQkwG6bNhZq1D2xlBT
DR9Muq7GZyop0+lpXmh1gest5hLiU9kusJrHEXUpluHadF4n3bSssRQv/+q3jHX5
TBoJ1LSPx5ahw6U/xjVT55fm3eV0HJihCCxBwJmCF/lJWITQ32/ovnFXpO6C00ui
F8oSi7XJkmEVhiwTFMwI58rfiFkuvWUbRb6oUf2c9ibZaMUCjx9A5bSmaYPr22fs
WJjErkDmuRsM/gAZnDzUe1h8G6KA2SAc2HWU8kX3nQCS+8LxN0uDgEtkyP6yok0s
1UvcNQii9szA8VUCCzp3My0HnwEdog6oYL7doXxVSshzFPBIy1z0XFXqA8HQ9Ft0
94oKIiyhQB+i9OoswxF0JPIBkSLmFJcSBKXYLAlS7tSpyzYcGcGH9s+BUPu2rFI9
2MljvikjbY6Xd45qW6ZDfw47D9Os6hyjsuHifNfExUNKfHQMqtTsbmzMPH4ikESE
hcUbOA5YtjmvQSqsexNYcRfLEQ1CkPyqX939tKj96qN5tfyhzQzteFrEPId62GbL
Eqas3OgW9Td9JbQSc4pgOX5euJa0LREtjg5RsQl9WZUclc3Q1nnurTJiG/ytnZBC
DLsbLCgzT2s4ep7Qr/uMtMNq7Sxf8yrVDwss1PZAUMu75AQY9qo0q9A9NoIlVZd4
pTAcA1fb8xgrgAa1kp5IJvDJsr918kxBePDHAeWNdPoLf13pCYYyRxO+pi3Ic5vO
N8NhJxQvElaOEga/j0sxiwmpJnIHAcsjXWGO94WnSlVv3X1A3A/NyuUKzGDXyYxK
3x185eiWFycJ3NYypsU+0WaffBlHOCvPheaDHuIWKiFQaaeNmsbOjywe6tduEHwH
FQ8+UcdE87WL6UsDellBvrYPwDGyJEPS5R5UFUbxbmwNTfHyofpt5tTvQKpjg06n
RWfO2rzhGw+Gq7OI9TbHBlrhyr1prpdv2KiDcz1TzxHY0ejY//z6Te+dJR4KfoMr
7ooLybIerg0sNM/x4YQNbNfQwMcz6oSPc+Wi/TgoZ3/FqA8fQOjJ/P1/HTN7+ahV
DMqyi31MO0jwNimwJb7lOjetWxFrbJcdFrKvTBh9XQZy9V1qskw5J5lRuroC7At+
d7wnPeHqAAC3YME2lMaWqdME/mOzC6xadtI/9IrnIvOYFBW0+oljaqq22yXgPGgC
bVBUKQWfQdrA3A3pykmUcm9OlqeEFic5GjWKemH04xfZM5idubBFQpRNK5mg5xRj
sxyPb+49JbYLhLi1ImAsVBABOXDYnO7+7bHb+p1EN4mZ+m0Vt+RSaJL65mFHfnnF
kpYmmRYlypC3clVapYp5gylkFnmMEq3qdU9ndduiNPeYvUZvN24v/ZXZfG6DZomb
Mrrqf7PhpVWBTYbjnoORuncM/6SfliJyOcON2zq7vlFG7HQpoG1wKqXmyj6gOddO
L9IOU49bUGSp5honpnJhvM5Cru3aXtJIDHwqq2V+z5t2Mm7dLKZjUHnASNFnfFQE
M49o3MiIyVj4skgIFMNdUD1P13NHGmIohm95xNgw1OgPPe8pqSkNreT6oXB3p6cx
9UGMP9pNBffElbjbObLQ8AlCvJxFjxmQ9uZVNe4i8ttZSlwaOPzpkwQIMG+WO5RW
11fMunUIZGiTI9AHuaLro79h4IHBn3xUVJwk2nLYTPxmYmtUDsLNAuRVDWCyVwrF
Y9Bo3DgmxyzaJm0FY7CVS4ATgYUGTun7mXG/5s2s8TuKNd8K3bCQZ3Y87qWHx+9p
/3pW7d+6CPjwfwYp0kw4teoF/00qiM7PSNJiM2hs9cLbXJbhVcQxaNcYc4d5YQo4
O+ck0dS1LYfrpuOHBe42+UBhJYBNxfo4oboWND514HPEmTOlNlH+j+SYyJ/p5UNj
DccvFy7UHApEmCccvxRYbk+kt1OKhiEfz6UcQYeAIFvrvaFGqNsjeLIJ85piCdWt
h97uypFEZSTJNJ6hQiqYxNr3/PvgX7sAzdQbgOfcKFhqCc3wPE7xsRB7BaAsjZRi
IxEz2hL/J60WXNZzMScdrnFZROCelVvSCyStHGYcIuBSUUvThEoMM1tcWMvDBnLN
otcsrdRkNN+AJcLNkDYYkNHNJOdN+ssKTyWbpFxlgS/Zl2L+G3jJmdED9/wpkrH6
7PGqyJt4AOxdMZyjCPhSiyeoO2ty1VmS0tSO98bAlBdmXhE21Tui40ZP6hR1C+CN
J9fkR1DrWfmAqtwHX5z12Rjn73jUt6dfmGOgLCy12HJq1vqsqOJBpmaW3/aXMQN/
Ow+OqPayj0hDKEDs9WKvwjp71n/HMcRG0SxWYFNzdZkkD6Mwd8QSRPO5pmgsIeW7
kHIEs+5dyhfSTUzW4RdF876Tn8PYUzfeU9WgZC7efPNs9t0psTzR/fkngE41lms+
7JIBikN72Mx77SjYuOePp4q475i78WevU6vVyoJPl4/IADpP/q5AeOaYIoGc4I6I
K9Jbn8zYvetfN5+3y+ZSiA7zokGNRqNzw27OChujn1RXBJWXCNGqc6cL1FzELUBE
OHVK+xDwjVEOAfnK8c1Jh0kMdkAawOM5mWfPAsU16QWGvllTMEQ1/Tj2ZomTWVmZ
qlfOHcFxs7gC7qXaah1dJNUs6WgEN/mqCO5ygIOH2dJLXSjs6ApuMrB84gFbii/j
LsAXJXQii+MEYR83oqVW64bnil8kzr1j8+/Du/KeS4+gx/acQi9FWZVbuvH0Qo2W
TkmiJ1oOnqIVPZzHhGLSH3HKTW44lIPPIyq+d1JTHx3G1+tSQwqnQgt5uP4DB/Au
XOPBCqWdz7HOtRMXDDs99p5SYBWRZqDr8sCCAmIwjcd4h0H6veFc3ZLXySZb3Dqx
7G3qo2qTeF4gFHkmcg8hyLtZ0GO8nhqeoQW0+Z/0WlX5QGGcQePx7A1+VJfsuHXH
MCzkE7NMvnTpWodp9dNureEyhXL5NAZzQsg9MQQuZeF1gASPNghG9MFLABG0o2QQ
v2MoM8daUK7kX6ZFcCdLLlORTS6gFM/TJp4shRiFg4imBex/QNO8V+vMNwOF/CG/
IOiEa3KlDqOBfZjFZXkpxFJGnpqZKlVRnaMKvFWridD9DIYtv7SxT6vQL+Wrb9tp
GcLuxZpzqzyZSypUCz6itaYmKuP0ALy06Z/NrWbbf6qFr0ftfC195EHTYmMif/z8
2s2NucdPg/wJX8HPM9W9RFOT5SlavSzPGDS4uBYcYitfgGsCbaeLY/7Qqo7DpQ4G
7jCC96gw5lB/wW6na46qqoVN6R55WyWLx9Qk9BIzjFT+FbL7WVQ17a/YtJxXH/Hp
wI9CxqbraYHEHRLrNN/z+UZIpd6enjpop+z2qV4UyazepTkdJXxq3WRup+rtTE3N
0wO+aHD8Iz0iIJEn9ffNYhHjzjA1wk4Tt/PStUMPguH6csnaswrCAPwfcU7iI4Dp
a940ek7IsyJt7dFS/FDffCl13ok6ouX591uvQTdjTECX9LrJJVC5HuCyHMTQNZwy
TyHh4VD5nqweJ1GzfJ4KvhyQhdG2u9JmiuDifbj74ukF86GGJCKus6LGbYn6ExdH
cgmMj7xUowkfr25PB803iPWYVOZ+NmZv7IC2v+57gP0JCbRAMcymEBV/PzAMmM4o
1NQ0mYMrAFENExoaZKFyo0RGghYdTCrQ3w83Lmb5xbhdxug2HoM8+5Xn9OdssX63
lrDY73EoLtmN7n+tka0/t8oBiNiSKctjAFTg8rPfeHDjINDnkb9hCI9y4K+yaDn3
j3DtP3Cl7i31nYBhNoV5yh0RW0NP2w4dHoSSjA7AOwHsdFDzNTJiyhjbd5rONPJ2
nLxuN3jz5UEhFLp2JtGJA77mouoKZRVOlAVYVAL3xQnxRoMWOoDqe5uRQvpuEnkb
9EBRGc73N7Ms9/SR3avQyX8wBhVVMI18N6WvnI01QO/oXuI3kIZTeyE0R6Pgj1MO
5PfLvhE4I95JrDwUQm9YKVcwcjuPrS93ajwsyB+dV4mndZ7tL5Lasknin8WwG/tT
jkBRm3Zn3nw/nRqYcox1/rjGQjsDCTkjuyzDaJ1TulYFlHrs5UUyH3Y5Whc7zLRz
TPxMzq1I2g+RBa7jzHgQxsiwqzO8ZAA1BrtlCAN59q96FN5dVk6i6er4cYJ/eW06
mfIq/bpZuFOda9U+Ft5rUemllHgG2MJBYa6cv36GFEMk23RbsqVg/U8abwSaRWBU
dmf5AwqN8ods9nqfjCUpAAX67WY2p9NCMbCZwBQMTVo2K9RwUU3B+o5YCl117Lrx
7/JWFv8KYnB/3ze0vY2hFtHbalHO5j+tGrkTMzU3BtpUPqTwoCKzniI/nkwFvcqt
rykGFfSaK4FTzfVgdSyC2dGPxzTVmOhb1uGhF08gfQjHo0ncgO9gTA1ZhD//DEUH
4oMq19Bqo7rjTe7wx7JdJyuyji4kPTK0X1pV7NOKNmjg6RS4nHeUosE8U+R7B3Qu
jagjRt+WjWbfGAEmeb3wVF035RbkTJFMJThRmud7mm9+3umfEZ2QS1cGoisZo2HJ
ZM8+AClgmbmDpbYPFlgoqV4cBTH9TOi0hm4TZxRtfT0FTe94Rjau7ZI/hmNqAYZ/
xJtW8BfCOAVDxRcw8fqaUvkXbzpCBqB87ALW0lzTTrq9vT6Wkvl6PziGafQ2Zk1l
ZnnCadm12S8hStZlIqb3iT2WLH1yDFjjoI44m+VhIqsTNmhYdcfk0/pFFyU5e1Vk
s5AtTLpdRpgjvAEOeSNKHHJNJjFtLYoGzCdppWiL1QlrbRXhphUs4D2qimgexMRs
KV4MTtGSG4YQsUWCWg7iRSCUy8qT8t8zBrjXIJiJPWBbYZHNhSToAPf1+WVEIb+P
OCEJEBML44jpMyxnps9stdwKs8zvdBRspL0fDWt5FJQRGwhwqAOilyjhDiQlm5YS
XlKOrZNOiwboE6d/OnsRi8aszT4iOUp1IDlmwPrfWz3IGe2w7wWW19k3iajEg2pR
YsOqHgx8a5FHlHeY5DgvFKWIIM1zThx3sqbc5VXtT6d8dEejSVntAdyqPeK57ASD
9b6ERwms7EYCNQP1gQhrLAByTaO8/Wi2l5BCjl4iPXYw+6YX42H7fg6y2tCAlQ6U
f+mXImh7UeR05OGaWtB/fEKqQLB9bI49RHOkmNEPtFhuwTQCRH9kxq/2TLvQcaNn
IMr7IMq5ULrFj2x+8S8i4C8fLSwkXOAhXx6cM8j3QwllwMrLxHh+UEADcYfaWnj5
tk+hZGoVG1JZSB0M78h6y4x3Hi1v1Yfi/lP80ABS8sZi2S890p8PoyO56GI3NwAh
HB/ynQQ6gu1/gLF0PoU91PHqCR04kjNJphE0JDMSX2A5NpVx5YGNzkSLKkP/VP/k
NbHqtr/bSriu4Q26pVACpHMltFmVwU5vxxMPXLViJZr69G62pP44JS/ZuR5LfoNf
hyxJ8d7jmsY56G1RwuEoGEGmtfSL2U2vM6KKJcOsOh7+xR1JHPo43IiAUlINKAWB
dpI2dehsFQIpcajV/F+DDVzQgGzmU5dEN2ruBXawbuaxtXyh8YD2Md3uGiqxMZwd
mMWYQRcGcY7PldGzhJ3UCze4+jB1VxSubpZ2CkoomSgKy+2kNsuXv0IUvGjPqqrE
ayHMU+YxBQLh17pQfc/6d8T3lmBz5V2W2Y0I38atXcT42gqnqeKetVxXEOUH8wsq
iX7A3qyZJPdFmQUmYQbrSmTGeid+omknBlA570piGjbY+3+5L91tzZtAFXCCIYM6
jx5QFXIVunYNd05SkmfPE8lEY6qqGAJfnTKucenVSqvPeB2SC4Jm4lS9F7TmWFLQ
t5r8lRNSEGN0X4qYNOuW53zspAMO1+8T50lpmXFyt3W4qBOIRGEqYs7Aa5SOuklz
H6ERpO2N8931Sw/dyEC/y+KQ0NXlFrGuq6sn/t8hRfk5LjiMOYE6XLT3yTC1/myJ
fIl19ycbiDW2X45+/t+ufZq5keWh+0wq4XEHED6I6l06x5P28gEu7WjF09HHc1O6
NF9Yx3R7Z2c46v9b1J5rtEtUOaY6Ao9pjQIgP6q/K63kCsgLNGJ+8eYdyxEO6Wdk
P+W5l21d5XtswPJOc1K6jmc2Ui2LV6zoBbDu2JrZruyWW1IER2HaMw8f2ofmn285
EiC0UuZNx2KDpGi5hDB0nGwq3UZYTGWxWsMkSeqvESZmDRH7hseWFJX/shqaPkUg
XyfTqaHoT0s0rGtdKRwiWvpKauug8A5hlp9Viu5UpcwVFdzeKF38hBzxmvquuNXO
uA62MAMrj2TA2L/SdDDK5cYwLXUc/8S37zyrKOPEgOtWAe6ngb6tD86UMFA3n3I8
8rBUZ+mdSbVkYGH34H+cCzQqj0jUVFiLHXN+TRTsp2qbOQ5vfmwqIFxg/rWiLJLz
LjIHFl2IZkWHb2Fvzf3hM0Ss4WnwOOMri1TuLQoldk+/dYGE8y97KwJ6ekMY3+Ao
svZpj7hztrdyp9Howp+Ex7N3wUG5ZsQiuetup7UXw5UJ+AWU/FVGfmWXHA0bA2oH
BMI+/nqk215DM/IHvO9vYUEJGHKJjmrq/r/AR/Hf+EPmzeyCSpbv+6l88MTAhDR8
mtkM84Xkj48FalHToxXCCDcs+JiAGjlpoiZiMOHIXyM9FefWc3ZScd4POhZYvk5N
fmJ0J9B5WdFMd2REFxactJMMjNjI4QhlfFsUTKU4TNfwbixb70khWgBYdcHNzywK
9sB2mmlQve3p6+Mbgd4giJhte1mbuMGPL4A81T+hoHK2qO5LDRkN3WSfn8gDPBL5
QVNp+F14jkhTuEpa47JWzJizgQJu/vYnUkcvp8TjLEku0a0xuo1MCNmhzYPg3V6T
cndtXebke8xEaXb56NAfYK2pAV3CYM3QtsIdbL5LUisg+cqWzdlhgF3JMsy5CFxH
IW/LrgZIMFT/linc5J3SqwM1cRelbXCuNTkps/cPXDkPP6n1fkBiP4x5Ywz/U1oV
kLyYk2/WSBhHeObozkuF8NoKaoXJbVnqhCne688FafWAkvuhkb1QGeuN+I15uaWw
wvGDP0cjmjUqQaj6WF6YLvf2pq1HE8dBvZPKigH1k35NqdItQvhBnNHDegGJCsMT
bI5LQR1NvtCvn6Y7mRTiCGlhAxj3Jse2hJpjsKIYLbLd9vFIVb38kXoZFSQOYqXt
xOXys7L/H3ccdhmd/ODMXRt7F19qYPbOzpRWs+jrdJSxIT5tmLE0xlXml852DvrQ
duAzDWWZ41aru40Oo81AgoF6HPH/kw0kBDZDjFucM/6Tf0oq4jUe+zOP1uVfY2PR
IsR0stU+E2HtUCqhlPvwUvqEDidZTB3RbLlmdc2jGG78eEwSZucsOUArZT/jOP+1
aPuKKldktwtMyqGVOJtTMVqf58uuNxIdx77TckYIUXuZHH0f0jZl19BKZOg640N3
5VUf2dU2TdkzbKlscqS8MizU8nsYb9VHRfd7WzIFZ/cfC4P+0mZbptWQqCWVqKTV
DI1QEfFCQxFQw8TKeymHhE7kPsoPNhzZ1+Pg7boo5YuIJttxk0P3+zagNtPf3WMM
8dFrcnulLpE42y3v1JvIxebq+iHIxYQ61Kq5/NtWaNP3C+hRHTzR2muB7YS4cEZw
oHIS4VnCP2AJolFQkj2bcfi12oxKCtnmAJhCiCJ5lj/xq4p+eF1bN2GDmLKUxmTo
ls1L7LVeDTMs5EyFhagCeZCDDWptOT+MyQGJjsHEnLiSyYvBICSO9wvvmQggcsLE
kJGZsVQ6gl2sJgYFuM1T7+T/6PtztnnLJ2vckLUprm8M39E0+D9apST1/kBeozr6
oElXCmzd7eY5lkj9Mx20kvd8vzxg7+kTCMpY2zzh1tavdD2Zuvef3wYGVrbz9hAY
u0g/ewW4dadBCddCB/+ssDQ+UdSUbDlBPyjE1fPSqCgYONbTUb1Ih1DTnch+ejsp
uEiuAgCzQSyALEqrhbR5elCzn7my5Mp/sMH3NR7uSXeoDKwkwAsT5mjwo7re/UJp
HVliKL99nx/slrk72pWWr/gLXtqmR2R1YwSg1W94MGKwvUTBBBk5nCSqjTCIWc8p
1EDljlYpBTdP28seuDw4JHbD7lAzq2M/bv2XpX5mDI+vm+UhovxPXxNSbykZ7cMw
rIyZjcXwz4pWL0C40Oz+YJ/pxyLCyo78fde/Q4+8cOmceAOzuyhjpj/6jhl+9DqA
XqhYheJu5TEYNXeTuhR4gP/iBFXA0YCS64yuyP3xYMwNbBQaaI/kwLSvvmF85kH8
netPVX7OlUjOor6I6mIsBu6o48VRDE7gZuBoNrgxSoWMfWKa77x8MS0cmTm3HygE
OzmQXalhdkE2QOgnxXqUdRULDtMss/kI+oEYOxlFgiwR5Z+fxWwRdE2O88ZT8mET
Fofr3J3AFN8ZRgLYhjtLVofjnnjO/ZR06j2rGEh+lGFpvuPe4yJe41lo1NZapAvj
5vvvcbvkMBgfJWjOrCzMjSByb16U3/EraJ5N5Tb38MJ8XUKjD7dnX0Jr32kKLkOk
jcfm/CwWNPsuUVw9mH9TR58HIu0lKvOQER3X0abINUKokIF0Giz6ujYBnxwglTYr
jwe0cZBAPRqzTZNJEgUY39J+Dov/oUHrDWJRUzqu8mOm8otJBV0UFXJlZ1gpOj+g
4kzVXXQp3wYQDxMUy54QsRSdoO3/bq7taAO2AwqKEO/D70gH6/mDK9LNEY9qrsRo
QPjmMBt4XPLFDG+GcRC8/5vwesvTD81AZfkVZVZGg++BI7mi147ac8yliRkXxme6
alnP5Nk4AwYYoi/enPofFIrkD8UkAugrnymegdEnHv3NGVPHowD/At9X23Ydj/Ji
LveqvjpBwjZUaZ9UZIGRlig4IpcBOwd4KsWoXqamJw3l4njfVaWEzjMFJXhsdJ6j
bXWTORU5m2QzbBBwjfoXoOzZ23pca2K/60/urGF5p8QuBfoSGqt0AtW5if38BkRC
13iwVoYOIh348bskMAFy63i6OwTyN3dvvDXc/bbgSZPWSakA5Hf2KhupQLNw32ot
YMIwovIgbaOUwZXFk8g2tDluvz/mrxPHCQONBVabygCFlatISfy7yh3DKXZoQL26
9rx3o1IRNkSE631Gt5IeF8JkZ2uEyLxGnZDylTtNzk5mA8GjPfWkbOwG+X0Mg6TX
1iecIJB7xskF5iFQJYSfQXiiCU8HrE4NK4aw4AUmsFRHx+oWjehJCVSQBHISEI7I
4tD+MmNbKdy9hHktI9J1wbMIofIfI6t5yhK2sZxSdF7EsG1BcMbpvSZjnAPN/xEG
tFwohktRHNdCFFYVXHqq0uZ/YG1fa32k1F4qSRGsDL4rB3WnKXWaYz1N7OkuRMq+
EluZjRGAUXrzXFbG8nq9IkBJUDeALI+z7Z+si7Y7yGm73izWHnY3K119tbipgb3m
adJhhJZGNIUirYZLD/CPgPGF4Niv2xa0SC/h6eQqrs9MzhFPM3TJjWUOuhzoHlQa
VVmiUmBdPKV02V2/hDSnBioMgiqWrx7PlaCa4yXqWpPWSzT4zxTheR/6V0pQI0xb
HTXpLe2HFBXFcgDCDXqc92IH0MkM8kbHA9OS03T10ipHO7aEPDis72CqkFIGb1PL
/iUbK6YKmR0B4KQrFy/4dKZgv5BhjvMZ5Qa0GbACc7YYHvDBkqfGaTKLN5tUgWkO
pIS3+oGIacGNcD6yeKK+uEfF8vxhoPvmgLEh3+81Mx0vyrKO6LFosXBEQJ2EmNXV
2/d377gyamgt4/QAuq9UYZPFW/CtMrTgyAlX4zRpLRW61TQYeJjeQMxDpYgrMIdw
ibkUiyN8qd5G04jN9QU6ITaX+0e4gYgRD1JULhbu9BcMTQ+dRs27mgpN17PhdN7I
9hW/Ax3/l0s+gJjosqxTiwdW+RCVzPwqO90/gmYqdQDXE5NtvpbOaf3S0YbYTlSu
T1AAqRgJ8RUHX2FM7yBDaKcSK0lpra1NbunDjHFK5v9errj2iLLNUK6BUT2WcmlJ
eLJrnYkq9sKA9sKaGbPxsT2TCYQuWUp12m3zHdR/HKwDzAtVNiC8fEt0s0IhYxJq
pagbuJDigXkXVrloCW8BmdYyKPk50S8W5YNV3Bn3mxQy4dCH0y3YYo6xE3NuCvfH
9TLHuXgJoQSpvHJ+ZGaWfvPOcc3EjfnfTbKZBjvbZweHD9Zge2KF2QHYTBM53KEw
Bsdw1btLXpC51UukCseNp1BDZotiDH+P4dWw39pHJwmIWrYtRcs1NMpfiqqNVm/8
bM9t77lOENK6OMZSKJt2gWQIMYFszmfB9ZXwPKs4jPLXrWTjkSVBcAoj+iDzcgKm
0se9txxeDbwgX+v8iz42FeEaYky/kxCf0rg2tIxC3CPuTuiTX+F6hWatmlL5vK0S
KOXzfbxfDGYE3BeWoMDx50iGWGPgfXRjoC1jqL2FYz/6dXEANpK/aE+WC1KEzAfc
2Go9JRTI+sw2KvVRgw3SLOBtBtgaBjsB6P5zQxrEElLMwGeY2o2DaS6g3h+6rIRH
37WvL8FrSMprrwFIbA9MxiFs3IVdPapUsuyzjaXdOsY0GlPjlgMGBRsHppk1z59l
Vipfb1XN9dYaUx18NyPSTbf/O7SciWtb6Anet3CsM2GiLu2UPrnX1pE9/FBooj5V
Jf1YoJ0RrSbPfyzDKSTpfYTe2ES7I95dEhNh/wGkDNgLIAFoRhcxbWPt0H9/fGVI
fEUSacQkjxjRnmiTjoQ5oB29SrsdAX8vYgwI7K3o5Vg+e44yiIO+YgHK5oi93TTo
KO+ummEPU9XIaiZuK1NVoHFUV6CHdjZEORFz1Na4WARr3jsasPgg/ujx5GO1/aYS
BAFmVV7qzDLZfvLpUwgYkrU4zgnG/Ov/oY935ctcbvEYTUdw6/pFqHgiOFvfCf4T
pa001YIPOVldJc1YkQi90v1iwu0veINPrIICAvt1JBdKMvDbyGdbe9V2KNskGZkx
drv0gsYtGt3Vv3L8o8GiJWgFtwo9uqGtI25CRfbamZYk3lmlmYhe1B8CIddR9IPK
RUVdFhtysZck5Hb0FYws5y5nbmxS7VehmQhow/o9BK4wHtJlaVI6U/I3pVYAqYHW
xLXuDZyZJ+BLZL07CYW3AMBuGxoq5jio4Tm3zFDhJv8zPr+VgoAyVk2pWoXZ3axM
P/tOslzQTNg8D9SFpHeh6lSL4A/qowBXbv+3oHOQQWdgSmAcPYEPWRbZ6RPPBakr
q28lsF1tS/indppM82pSK0ahWfEzme3hNURrnAVF7oAeefJjSENJYAzipWLRhrs0
DO3uaiqwyym5/EA+m9YQjf6tiK92Pch9diV8a4BTv9obhwx53vZe1yivwYe/izlT
XDcBPJFcsLgivbAYezCUsJus3lRD4mpxGH1E3Fr5zDl9DL/n+E4KFwCAt+po5dvT
bZzD5sbGSYxzzjv7M1MIapYF+fIlo0Z025cHB7UKaUQU00rONvaQDEPkF6X9dcQh
Az7758Tn2wflA74jbBVgMWl1z7n4KfPv4Uk/L3mlO3cIT+d8iH4h9P0xtVXVmrRx
8hDW8fTJ0oBtXC6Ixw1C2habsvQSaeYH+Y2znc0TrZnlEXZfn+DpvZUPDmojaj5H
r9NsM7ZJb9h77bAJe1/x5zvYc1kUcdbGb0ercNZgrwkGq6sy8VVovvINHzR6Xk4V
wpelKyxEadH0PD0TgPSTWFXNGQ2vnDEFvUwfKW4btfhm5q5CPskySb4h/0Rys2/r
8MJ+urGtZeudg1+PbH59XkTjxgLSynRZEm4ottoWgwEy5KhxlY+xuaN/ypgymAj3
bwv5e01Af8EMHXFlGw2KBsry8cCnVOcKZc2imMs16BK3IsilWSCTt55GOHzq4KMk
Y6MrExS1Cf6uQUn13ZVTd7KwegRTQY5zcqis7EZtsCLarnI4KyvRT2j6wgup1yku
x7cLTHAqByb7ft+G+t0DzItNRVt4GfsXVE5a31plR34vrkI2VvC+2yT2lmnvueUZ
x3x5tEpJ3AGrEmFPlp9XTCqdfpIe9HV2xk+UbGcXatAXMu7Tc5oicDacoP1E95xz
7uhUERlNUwx16AcMxvjJys8WSilok8yWkJatD9w3O4HhinQArbvt9DPJYXyEtUuC
Ah7rwKoUbp1t0ni1l5/iBoXKUqehb1cvX+3lIcwURRW33EwnRy2aaC3bCQrqX7La
lsDwkRxPiPCgKN20QkdsaKLzlNji+UTOT9yGV0jG9XkDOv6al6i334nluZEUz2/K
zXcnBZVSNuA74AJMSz2RWX+Ov8K0jUlsdqnYnTnInRmkEjHhr5n62IiFVOpkJvlz
AsGl+WTgK0hGHEemWn8E7VEjRfx3/fooVu2teBwJXnj5vO1kCaurF3VTmxVz60VV
NqN7ZJ1qm0N4Qb+wSBLN+pM9dc9VsWUm5xtlYke3PHPaB4XAiXPrJOpxMDlPZV+P
qP/KhnpSYwve2+lv++Lyo487vr0VINgc2E5pnndKkwCOIVK5pkQCZYIVnXhPWkzm
pLCSFpHh3nyKITbuBabYv0xgzeU+m6ur4Sgn6nA+yBY0SbMoKlQ1HK1weyjqWEVX
X0xmnS3udIFDm/nTHAehO4JYLOUikNlYd/jqaMIwXxaRneAT3h8/HFnTECiRpmKj
g+VPy/WyQI46OKgUrixSiIlbgs3hxl7yWFSxgWaeGGF5c21OHU8iLBl5GmjTVJge
eer1cVNR3CAYmvvqYYKQRdZAeOZMtUP4OtdhNFXAAoO1pMQcq7oVyIAgjz+sUL3i
kn3iMnHP901dTp2BlJ11LmyTGoCMM6YJtgf1PkrTXFlSEt5iNutlNi+FGExrX2+N
dGS7b4NK+wOJHKhB0tAIXmEtpGM3Q+iBcenBruE+D6d5WHshM1m95n5LMRNlbXdp
2bqL9I/lowgtWu4auzX9h+vEZbewgbbuKr/fFgX8o7Y4XIuB2W5RfQq6OHU3sRDI
D7TatG/ab8WsVCLZF73+I6hcW2vrWLP23s6+7cFFIxEQYxey+vlhnxMUpU8qjUEc
//D9FTe9WzgMbTZDhKx16aC4G2ZALXl+E+TUcOknNwKbegRsZECaLmOcaCLblPjx
VrsVE6bYVXGDqypNz85P0zHJzLOJL+ANwOX7oE8U8TTBtIMnnhMzlnqEkkz0Aihj
/JnETrXR7fGXYmoT5iM9+Sv4KafOUiMKUxP1zb91t/N1ij1QF8djtIfeCavc9NNM
Eyt0CRGGTg0HtnsAfB8XZcj/SqiaNsvkutZyxt032ZgmdX+653+LBu7C4vhX2G3e
j2rwFtRRXXC2dffSDZ991qfOwwLNRXZACTtouI5wJo92L7dxcpvEW7nmCdeGl2dW
mucDTeELnSeKFMxpIxm3qhFS9i6e+9Sbq0hTNjzX9bo18QBGo2ueqx50QTWuDDag
cPajppjGJeNzoUkXFdEJgWaBvgzQp4lqdOV1yC8uY5UGarSb4sWBL1aLgwte+QD7
ffvEQgwWS/dQs1E4+588Sskgxd4mePRo6bFZf5vIANnJ3Z1ajyf7/5XmjU6+v/d0
yAApnQoBS8IOqJ6HtogiP8naQfzAZQAFKG3C5jaqr/n6PZdth4Dn59GgRgAkTKIM
+PKIoBAf6PGdIc/DpbDvN+bYw7SF8BDBD7aHige5fXDRfIOGcNlS3Ef/OjMBfooa
hGnKxVc4vcjRKZ2T9SoZgnrN97kCBLkI2POEndBn9zw2V/FXt2IyISLRCh04exl1
JmoAMZEafTOt41buAhfOkyhS1pHiE4OcRkAm9qGbrDg4JrdJFDOFKb1ynWIGnH7X
mlYivPeGZ52dPEm50RX7PRXYbn9Ah7j/KWc9GIK7Sg5a2k4EzAwURhOE3ucjRIwp
5LU78ynsYfyR/Jlay1FNFnkQhytR/wgKGucwkycYE4Z5gDuhCHS41YBzz/5S3LXH
9iLbc+BewlSzaHz8amRsg/KW6Yf1mvJ/Sumit7XL0Tm5na1qJkDDEg/a+QD5FMaU
9rCZ440kqNHpaoePfE1ZAUC7BgJnq0IybnTVOSze77v9rWk6MT2WSW49zkelctoa
VKdw5za0DLmCpIeK9Yy2pUeu1YYO0vZSSP3bzogMKhsvmKAcPm2FMtvTKDtUmUlK
ZSSUaCRpnBbJ4JsCkwQtx2fNBwxAuCQPbwR6F2qwr9rcjmv0vSalztdcq9IN8z3L
kBmpEGvT52HSAvu374Twd1eXDfj1ZiXA5kf9jtAMKVTX54WZcOhvZsINExSJA0wM
hVfQhFDuZEQSnSJgVL2qJyetueFiTIL7VGCxQr+T7bSJ4lHrJEL2ziBpl3a25Jpa
V9O1ClhmcpNFHosQTG7GboJdFtoCf9iXSWV+d9P7FXUEdJsVVvtcEnU2L1tjovzn
L16IDLGmKu9sLrirnva08pcW37RBFa9Ecu12gdYheebgrjkCQPfp3Em9Gd6VHZVR
mVVGMIGIGfcmFuEDj1W6NJJHOknmtgMO5ar6sXjoesRi4g4pmXq2QZCNA9ArX9k0
syVUou8fLQFCg0LuEeQ6EIx3vqgJ5+PbSL+drb7ywAZrrxjunb1PIbD90516fniX
o9fkkosI6/EsRWHgJmnXf/c98uYIp3x8Ox1LX4MhhxRO5BuEMugAwooUczp8hCZC
CnfpyJmYIv4EC+v64Nt0zpM2DJwH6E0vaDGbWxM4HWBzW562jOL/1uuReiV1D7ao
BV3Ixd8z4NubyfCLbpouj1DSL/ArNq8mZgQLKQD5LpCTrdm9jK08MkFnDVYs5kpR
tpimD7mX0zjext0Eu3WMCjsbB7j0Y7UrgjALNzAU+fci+sNNJUo6LwMRABKkKBED
CBdX5JmMkBbrtAVR+IBUIofza1PFZWFB7b4KPs2eOw29BWqcbHyqvj0DVgcgZ4Lv
XigdG2ncEzVaKabkvSn351qRpalPy/6Ich0+PDI/B3Xt5ImhwJkb2egZXArBZJRQ
/JZ2X9hxvDEgtnKVzex0yh78dTI/C/nAPUcUwtMbKJbF0KRiZuG5rogMrWnHqh6Z
Ee1zx9vVrAXmEuRPDzOQWbsulaCDi/bb5/5OgqBNZIxzCcI9XoYY/OYcsbmzidUa
akWO1y1cUFt0QDNngyoV7+zDTvqUs7bxZGuNodLchSoueYJivVs/I7DaqyLU3prp
wgSIgS8up4julQiAAQZq3bITx+UAuX4U4x4Sy+JEzI6axIeISF32/zIOf6lIpl+c
hGDKc0KNEEqssPmA4+ShQ7VT1jJluwP0Nv0F05uAfFhnihiHlMNy8O0Mx+Miesvm
dbAFlUHrQcXVXJ3lMzJbD9GwjArFwORaogtWrBl00mlBchBHMa89FwQttmJ3xokr
jzg3TpcFjpLukDZxNUPKeNlTREh7VWPjMBhytKgKHXLcY+A60DOxQVAFfHYFOAbn
f4BmNRH10F6E5dzNB523D/y0hiRCFwnlpDfJ4oJcG84wEWNyBiKBUvM3+nx20yRF
w2cAMYREjK8rMEd9wkHtGDlYLf5kFr7YHyE0YU9R/Iv2ewHOu7yaZoGygEwp54MJ
FNg7nrufuAdqp9fhke/6HX8j6w8+0iSaxkMKlyBPW9DbuOcObKceWlkEwHG+0MQ6
MsIXwV2Ri7l5djoJnHQMKsUbiqIiIwCIqTD10sMiEn7lIhEQRZhEEQKktKd/c/Ca
5/FZF5Pk1OQpYjcOPwJALjRQ8S7D75KoHyV2xpasFfjgsJ5j7M/28ZbWKbZnscKf
8EugXHiLtddwmqVo47oVI+CQ6JpgnFXGOdApJY4NC8+CBQ8z8GnNey8McvT73Se6
fiSlDCkf7PeWiXO58mBlGDIO944diI7TaJKxSe9et+GZ6iunX/XVcV+L3VqDt2tY
aepFhuoLAPPubhTwhkToOKpuvGJAJAR7mMUUWqOxHEQu28NvhBFg2kKpPfeT6/Fo
aNwvd8zwav3iugtSNealuA7W3X/owxxMfa7yWIOwr22p5bW1f5HgZdt8wuNDrF2U
Z4rWrZLC4yYUSXp0gYx3mD1UrdyF2MGuxUiog/TUShEY3ASZTQWolkdFQ+D+gltA
k0sLhG2uQ5W7fPYy79G3lSXVupFTi5GPIJkte8HtSevwHh/AQdkZq5jNM4aMkH7k
JZFr+2azkO6WMeFkiZbTaDKIi7isUD4U7KcbRnXyBgTBPv4Zqtjj5FJNt7evpwYJ
Iie8F4D5MVKL6+wVrzVQiSEZ3KtojM5Vu2k2TK/+c537ouGL2L8sWSa6DPbNlRNd
ORib4HS5EcV5MRKE6k+kVj8GzZLaYYxlKLbz/8NLeflIFBOsYrjbvBrIpxvOpBox
ldaA7teQdTh+jEZray4iglGjvKE/wl/XxvHCyK97uKFcya5xAdSBZfYKtT/WJpwM
Dy2Ml0kPl4+t3/8J0IaucJeEyVo5rHRJqhH9s9LoD2GKAH2PdlHud4hGeJxXTVYB
+Vfn9eKP0m/rQj15L6sCnXX67ihFk83076ajLMRPPBv2eCuUb+1REM3h9VdgiBvV
pcene4DIkA0f32Ts+nO+0Sow9evxlXKKZLxsMxr+NGtIegcJLoWF7nkTs7Iilbx1
B9d9SUjGPKuYk1pTiB7zmvaGcSYE92NnsZVCT8WoVFSriTyhmHoIfLuPWMfvOCZQ
Q7lTP1bOz33JewCKk+jmiqf6hm3nGmVpAVowvwpLWUuCJooW8UCa5ATYDH5tPFEB
AVZpHFNwiJwt1aCV/7JwWWDJYKAQx5Q2J16nEBpCPdmHQ5Sqibu8gYX4dIVrtMaO
iLcaLWczZrf0wNAhhwzM6N99JN7fBFLA7A6ueEL8roHWDA7yhWImKrlmM3RPPTfR
xuV8IVoWAqzVLbTyA1tco+m3//hafFy1aDZ/FuJl0imNnpuGUCm+eHO3a5Z+wS4h
1fjq6EEEvpC2wc2O0zuwSAKTvIKQoKSZA4ex4oAwAHV3IrCfoV9bMciymWXNqk9u
oR3aM9KchvyNj9onGMHK6MrZMAd+njFNhYXhfE+QEP9MHOkVWN5TlrAR1VuS9w6L
MJ3tPZUSpvP39D1wt1rMmWhPzvNrCuZkDxkBwWhmoreXZXEgtpvad2Vu/URkeVVe
5VXreH+akSwPVO9mZONM+vLE4YKXiaWlPDK7bhOMyDflbLlKVt5Lq9G8PwPtG5vm
vI15QpAUdebyyM+azUCMrWJWZvCL3pgSifI0gS6jzzZHg4ayrKbylw3xl6BRUjV3
HA3RyAkNyob5/3J1D7AbVqntq2LGPhuIbDaHgYRynMAQUZPZF+0c6pZM6FVSUT2/
1FDo3Rwuy/LyCNc/se1JXxDIPY8N4d8cMNtAEJbQi7wmjJiYqZSr4/v/puxKBp3B
eiZvW+A8L/QAmWVcigBB66HbxI5MnCqjYCPWACzVMoVC/UXJbuMxiuoy+Qv7Dsfk
mxAnJhe2vGN93omJ39enEd+PSb/7H0BhCxZEhrKP351J7qU96ef3kyQZA6lUhhA8
EwnubCU54sy4XwsJXyzSsyiiwDzdcYHLGI4GqwdWy8OGHcOgG3AqGSqjp2rsv1dz
NFjk4tY/WA/EFMN4iK8nyJbT1ILkWxbIhltq47xVXvdLH+p46U7R3/VKuVJ2iS8n
XzEOMs6VDiSDvXawVwET35/hVLpOCBE2XaAjdgSgcrmSZ6wphNWqKdeUssxhX+8y
USjbLlVidVlEW9a258hkLpNw6qISg+K3xu6KKEIqLw3OqpgwOpk8z1QgBkeQgqix
X/CXZJ35YgLQ30N3ILABdUg9UJ08Xz2T22oE/qz6uaJNo3nRDo3w53HncATYTU32
2HX5cH0Rh4HhIwzBIXd0KhZ+mHZ275moLo+Po5hUiV+V6+evNAQJTxSNGVcQfnOf
VCn3mfumhN/K7/B4dx5fpkgQFhoxRAP3jbPfSJxn1+RjR6lUBauP3ggem4OSmXT2
6op8yXnepUFO5rjBuhtMTmBs/5kw5YvRdgN57y53J+hYdDru0O5Sovjuh4HCBQZh
+zYczUH6m971BKOphn4m3saVXe9lf3v8qPIQpKESvgnG7y5E4z7D/va0swY07QkG
jLzbk1W4Iuhmn4olEcXLYAG+3iWfY70avEjrPVQBR5ApcNyJL1sD8x9SOdMDykv1
KImxMDNuMYh7MzEmPGcySx7NTq+1OwjanbdkbmNftWZ2pIFPh9uKhM+mRDb3p5sl
f3oH9fLZ/H/t4wmo3OaRsI35mjwQmMVm1nbRMnH/qptXyKmwhi5uDshcMd4HphoV
z10mzAomOCRaB43BqpBftRexn9oU2bk5cer277PUH67qawuE9Z9cpuxxAzApkLr2
LqO5/JkAiAYG3GaUPdq9Krg9sh52WQ1EciWmc2R4Ha91m8LYumuL3ZeOdVljHHUT
rRDPDVwDCYuho6n7ipc8gv1cyGYn48UBvIw7+Jn6S2SV3xOSuN10JgzPWk1LvF+7
QLJkILXBvGf5MLUby5JY4nth0+t/MebGznbg70LAaCOtAGvHW/DK/8brBCHkD8uy
kMlAwKcbSMuqLKFNOCGyKaMBWIJIyf0AOTss4YLe74OoFPbWPIweY5maYzPdaHrk
mauFR2iFi+vfcyUnF/qdU4Kw8XCM4Yae7Ex3cu6CY6JbcYaijvtKadWiI6mtO5yp
DwdfUT/uY0xpYPM7UCMuZ1xmoXCrHNkvGco1kOmySdc9xXn4hLGf62fTSbmpEXTF
soQoPUZUrG7VHoWSeSs8Xqfj6dcW86rNxgHHL5LyaFq/ZPDTYDBOHDLoV+73Sd1a
3EzaKn8TZDDLabMl7uSP1CSfhKrii7QwbFDmTO1/MDqTq7GoU8hzIF11hW8qmqDf
bLUVkKfhp7Y5c2bvdcZqs0JfcBvVXmvpbzAj7LNNiN10IjuPyBoD2ZH3XqmIfics
hcKJkL5CHL8KOJNWWY5QcT10uF4LmLtAiX7HXbCzYVupGoxvAEaVpoAopUbAPt1+
HyJmOIbyz1dTuJwEEVvvNWpCIsyXtfAuiGtZWnEmvc9MwvCZ/LgJOEMEd5Tdc5gv
x62Yb6eYOjNF/Ml1u3cjM2trXLdRJVZBLn80usvd2Vu+G34puVmf01YTqoa3H2wM
RruwxwZ3KCwmvicexQzvnukFmAjKRK+aszaSKw9N1u/k6KvZnmVEO+JV1C2ELDiv
Vbn4cN5V5boRp6LdyQxNnhIo4vThiNlzqABqKwXJ293ipMJoIj6H7VFP60VZJ2An
U3QdbDkR28p7cUCUQEIuPrFZx/hUuqSzmuht5i1sMYJynuuoqUkaLSeSP5qGwvjg
BCFKp8bqPoN5VG6sgn8M4ew2vbs7Gt6xS0P9LCNVO5p0WT71RgoU7YLn7flDZsil
LRRCxJA70dCEJOTTkyyPX2SEU2bJCZnw8WsbeFZ/PLUF3b+6qk2+Tn+1k8XjbOV3
Kzjv3WEQWx7O9IMYQ4szgwQDuKnw9E/R5HhWYI8wqgzkdPyNDyUarBpczSaxDWpp
6meVfQxWsocruCm9+q3f8s2SjTvTrLHHMH2P42Kiq2Z1bVV/5OGJNZpRH/n8mJzG
iSbTyAwrPp0LOOyKPEYPVB/xqyJm3Y3M9XG/Rfbgv0VPCKCRNhfqYCC/ElnTDfYi
W795rweLfi3fM/qGb+JELekc8b8R6n9Q+7vKWQ6kwgCIYbgf/TwZcmS/8qduJGXd
Av22eQhUcIAqbl1kfJBxqQ3i+g/HmSGzGI9zdRRY6/FrRXE4nv1MTGSz1JL57S/k
64PgFIVCoFVhZ2ltuF+y0dEFIaXSocQMBVpla4PUN4uQZ5swkPeLx4FO7dTj7YvX
I55g+Y9gWdfQvAJABPeHdAzHsaOf1ZSnGhYHEYjvBvW3b8LSxhsvQ3pbqpGrwmZh
vYZh+63GpyuMx7z7Xm1PIXx9onipuU8gQdpzgXQ0PKkaTO4imYbKG0CKjco+3SRk
Vk3AI9r208A72WV3bmPPZeAFDp+EzWLbIu8OeWAuQul3iw/P2ex9jvX0lMM6LusN
GV0Ik37QhRVyK9jldDDb2597syzEHN+3Ni1EKRs4d3gKW9WrUbm6x2i50bUylUmh
bRgyLx6IcJSF+b/WshRkllMl84r5pz2lKpzzXHwVBtxJ3Ebarc99qN3kSodnGV/M
dkfdxs9gFKDeEoaebEl5FnI4MEZr73PfJb2eTB7CXafBQouzChlyI0EfgnTV+L+5
FcP3ARTD0v8K25prz3pHkL4nuyTNVIpUf2lCEITxiljs3ZrwPEBvjOf3pqNK1Ri/
fp571LJKs7eTZreEpsehLpr7ql+/F1SGu1B7BcjTSjTAVyoDnY4x1xbCkhbHK7qE
0fNwvJv/uXe5aibSEmZMXTWZxWfpoGwAzUf6atSRYynD86SVGIMm+qlDKya1gmZz
VCy/ern1uGr3CafpW5IL6M3uugENcOJClr0V8aDTagt0uoZAkiZ1ZsuAKSS4wES3
hUFsGDj3cuwScbEyQXSlFhUK+Lcto6W/iJWoRCCNzqxytGiHhPAWJriUSudeHtBb
8+ph4cMPksvPsY+fOYkBdsWY523Xun0gRr4TlGyxPBHHvf2qUckFOavaicAUVEya
xl4vCzCjBUQFkmK3sSCwQqziH2ksCG+IQocTWf/uAEBLVFM0TFG0kq+boG7Qy95o
JogyU3a3EYRl1ntcEOR3iwmoJwwwunhqsBdDNnK3V3xw3N41D887XU+TYL1F3sKS
/eJ+V+IEwr3kfvFTkwuFwaZ/1VSr3fkEP+KVztMUp5D2nS8bcWX+hOwSbSynJrAY
Ci7LfRVEf2OUvHc+daWNiuHhF/rMOe8XYZH70s5ND8fBpHEdfLK0TbcHsDOpvuo+
Z+QhPITAoXtI8wonoNptu28VDhIMYkscoDaiZJcjqPkg6JwwncgzZKHKadiTqNi1
y3NkdnTsGNzJnZ3zAAqaxrd305yJB3JNzro8smARLnjBw6ybPtjMa7I/aloNZxRU
nFnJr6paSKqP4NlWGw/U+/fMtHtY3Ya7VtdD7CzZqJNXDioA246z/MvDXzk1w0Jm
DQw0Yk+S5OfEuK1j/7ncozRtPNfkmCV0AvB8va/zIBwApawjLNnyfSNlGX6H6+VO
xMB72A0Nkpoeb7b2LdJFz7pkYXI8u39RAO5iwk/GUwBGm9xR1lMaIF4fRs5aWRHQ
ZVEbfAo7pfZtdkqYl94wMf2UOKx3KGVjplG9BMGjw/lFpWY7Vg2ajgef1TiK27zB
TmumaptCXQKXKWaFpmT/A4ma/0fdea1EvEKkEo67xj/ANpEh9V84+o6U4ebnJvsj
ziLgFkfXDza6QZsXHtz2iuszJH/cogmkXqgYOd5fpYdPYWsg79JxuY4Vq5mG9HfQ
4hB2+8aSY+Zgv8+gztUWYQ90R0DSkLW1jUiLflvHG6iwO5qIfjCGQfkmdHblyQuT
RF+xauqG/tahjcV0F67SKUIOjRHr2d1MBGs41Qo6QV18wlN43vnfubfy89k8DJkb
eVwCxkVnMR8mNQ3Yx6UFqEnmY3be1/lXcjOi5+nsh+ok06duWq+zQMXL7YMRXwCt
fgwCcVabiUoDPVy4WChEMnvh53YCyWhjrQDKCIkI+O2CJKFvIoPKWW/hzsp18YHb
NQCdybRsLtqDnWBLdk5DjGUepVmfRrXuz+YNrBFPW+enujxbf1vt3+PKN36YJzfD
b3PjFflcjpYYImb71v5yCRMGvvNVU3zm6PlmNOCIy5GWH0O8inyHuiypCiaB3amw
SuejC+w0jGUy6pjBA9eNk3Z/GPulNhNdUCkx/oLi+cCqi/gZEC0U8gOVw/VhGhlk
BDNhMVdln/fq6U8vHXg4inPFQhyZrIcdNi4A0v+Pu0f5AwuErQ8EWTNu+TxpwzBl
kGutgOUrtM0UCM+QAnTnM/JYaURS5iK8i7PSvgQ+o7SUuWfO8EaUtfP1sDiZtCm3
ytmK1p0QvTubruGWjogZgdfoB0LogdoHNM3sJ6IV1hDmP4kdYVoq0trckuDLQTbV
jIZCBodMJOh1StpG6zE7GLzUbCsJb78/Vk3shpgdQFbphTqbUvL0VAQJb0ZbOOTW
ht2dKyWfn93JvM//IESjE6s2NALFCpqeR1TtnvPc6Ssz2srpnj1i0k2pQWfT/s+a
s0vYGlamutW7INrChui53lOq1obeKCrfIyKjy5RldRHODqhh23sIJs9zKq+obBvv
ehpPPaJPBTcSqBy1T3x+75eYqQfC5R0F1OFSeN4LAv99V4eUC0x7pw3oHT6Y3Nsq
RyXI0mXf9FfRf7s5zrxU1r2hLdkPrtZ6I0THSjTaBqv0eyd5Ue+oYVrSSk1b5xQ1
HDS+EPTnnJ40ohrycIzvFUc/rROTA5cLn9WKyuozqsa6kXhIAUut1XwTnJ4cfi/o
qCXX/BrT0yxf8ic4WsUL/HCVX+mmXAY3iWXZl1UAX40S4MUqkFktj47OJh4dyfZV
kW1N0SNpddZCcW7XPZkD6W/W7OPhukJx5ddb61YDf7U5uGxqZdKzcksxe09iNgV1
UFiajsA85p/HHITRjRbQ4U6Q1s1ZA9MmDeJZkC57chOB2g4yYqj+HTG2TE6OrLyK
NNa+DHVj85RKex47xXD35To3P4S8IKKGGJkopH++B1HE3HPEPe7oG5t67gPLZypD
WjIg6M5fvCtYCMnGhEbXecrzWdrgCvgV9hefj/9Hgl7quEHFnLO/4WZBcL5AiVY+
IAOr+QX8f2KVeZzR5Vn4o5MHlEq3SVCH80LKVPbcY+n4rbeQ/3v+zO6wCM23O1WQ
9wnz8MveNn0LVACoVRFlKFsVWjUSAIv9fiULR+zxDbVWMlGSRNgYLKzgKA+mbqxC
wCSNj71KXkybtiws8JcGY4o+EQzIsb2yjaDup0/CW93l+PpWA8x8YHRV07oksW6V
DISVWIWjLRGWfvy72wOYo41lZA7I61nI403AlHyiUAIRbehIsxFfJ+V0puBDyFf2
ZsgtkSla7f7IqWC4Vaj6yKIBAIrjtoBd2jelrDKXe7at7XJUhw/oIQO4NbcHyWdE
09PXWYcOFmOrO8yJpuY1geZdKYIvPvbeiRdr+1AldGh8TVAWVCzXhsFkSnmbVWYr
Scy8sedOe1JS2Z+Hk+U4LdjYp1vNBMsU/u8a1lgERlwRw/SytoV7pVd3oZa9//Kv
fUPDAn3kO8R49alWwepe2ZuNDjLAdu8mYYXhaYVNmeEFRAiVlyN9R0B4ASLmOZdp
ts1jX02vFOtjhaMgUlWukmG9I7CX7dR1CTeFbhpDZMpH2UBFRTMTuiWn8Km2NW67
hFlvIQaYn0myhJ0h64knKcMj9A8diELgJyJASsz8FvhWaCV0t+tHn6QODSxwYFM9
II4dHJqxHo5FPFHBQY6297vSKiCr1VdqAarpP8xSya605ApMl8qTaCDA5Ch1S6U9
mxju2QylkWQ3eG3yU8wIqDoGlMo/BqS2db3l3XDSw8CvVw7K/zGHRNO8ZYyVCRLo
Tmb05y7Dokzng7PwD6yAEzRnNtZAeJZ0st0GNpvIXgTHQSc+ZXetf51oYB2nv4gA
PcIyclIMqi7HGzyoO4sFAjErzZc3FOCat4ptvxYV5V0OaXch7i+QRM+ZslLAT0el
lfWoiC2CVBtVatZwXZgvuhx2wRqbx16juXSXmCyJ47J1beUZPTz8AIGPxGVNb2FJ
1TXWc4pV8w6AJXEzrJGBR2tNcM4Tc8sgkbHcZ6vhGtWxGVeRlV2mW8RgLubkuzF7
IE8nv4rTTGNYxHUjQjnPBC5vlwLCUs/6dNc0wTgRH1431WSo57Wx4jrFHKhH7RYp
bQHn4eMrzUGFp0dYCs/DdMCbRMAcq3zIFjUB9wMwO0c5UHHibmG+BAA1y/sWAXHN
lpJagSqo+ETMJ+V8fThqM4NtNCAEdFDl5QBUxctuaRAd3B358Bx8wawXn5mavYF5
N5k6hn11cjb6IZLCAxCLOc5JUOxUIUttiX+7TW6083j7K8ZnzsFdg7WOvJrKuovA
3YbzUbFo9XALGp8j072TnVKK9aK5X3T97s/TQ9+r72BuTw5v32znvGIAWI+Ad38O
Fy+l5HAHyiN9Z1Ex4/rZkVk+llNcqL0VDgx8jB/5idBo+vrFi4iGzKnq6eW8HZfZ
BRcwrvr/mpVPu7nO4xVc7ltz3zgRPVPICfjFTOyJsbYfEaYAjKKbuwGcy6RscQGm
qsaHGQtkz8uKji/5zbes//vFxSBOCLNn7CdBGqSqA4kBR6XHrmrF4gpx5tXCD3OW
vGOufUpMe03926iaw2BNWOJrtevBv7GSSqHjqrxvDTij/lfxSAuWeG1FMgZhbfWo
Zu53fs/+Jf9OXocDZV5fiGvmJi0FDNbefKYRvDC8C4LoKCbX8Sj5bsXDbycgpA7x
370pK5AbREoZnBsMbVrlMpWOLCvoXUzkvx+dEtXz7BtFUFqmSFmh7vF9uWH91GIL
TfpEcii8ZBiis8LB0WQM0oRcIjFWBcldf+PEHpJuR2GIy9zMzhLzHeTzmiN//mqe
sItL18E1X1Tt2YHKjcVOAeCd3kQEzt6+iXHAlTMGnYCxlSLNDFLmL8ZkUKJlfkQC
G8Ze8FGwIOEQFx3CEGHSf28dCKdHz789V+OgsEa9b+c0y+sO0FN1wHYBzEVrKQ6v
Cz45N9L9lw+PYApj1cbzriGCWa0MkaLWNddKKD7Lk7vz7IGUtVzSHdHuK68o9MAK
j/Uqg+e1/CPWSeuDHBoY3ee4FT4jWIJM+7GrDVLOd7EB5dqsC+E51CzZUyLhNIi2
SSRiK8DDUqoeimq/M+hXHZ+amvohaCj4Z4DGvRyiHl3et6kd0K667WsgPy9C9aVW
RSyvkS3tPUWDAeSO4IgPQwarazjmNz9w3l1+OWrVgWoQLQ5sBwNtljg+Nns+CxJ9
7scjSSga9wDUFFxE43JY/H37os7KgUUKTf2RG3fkBQL8MU43UYEneWAI3KmM30TD
1NOf9sRa4036mMY99/1MSEr7pG7SbUSTfVR3RGGyIXIdgk+J9Wnyy+kRcEUNHTvP
V0isGQys91MAz6BqUcbgqeV8OtKvnqKZuyVWkVGxlEZSiNjQ4WQKtnoj+SDN7OuT
LK7a933tlHprAWJWA0PwqSmnY4ynIYol2HTBX9B7XsoMFYdWbDNrdFbWKUNuL29y
ZPuVZPIkuL01GCleZXqRN52zU4zaKoSRC2wP0hA3wxGHT2hUDCel4rzSENIkjb45
3EL82k8/JAd6iZkHfK4wPX8R56pVC2s5WKU7HghWH8LEQ1K654NgOZsyQeIRKdY6
TzrcrSs99B8cIC+9IieWFx+SvXCjDsqiWCU1TTlPOFqTtG/kf2yg3EsiniNp4byY
mA+BvAx3YcKgXrVYU6zD3cuLeyPuiuJCfwE3L7baDUZduzI9f5NWyiENm9AGJO63
uj+OSAlWQmH76gdJ8WL/NW8MiKLYOXkF+KXeOwA3IgKS8dneGZA0q0BbgrUyy9gs
b7O2G6E3Hw3nrzBvFAEGZkAG1tRskVgMYaBUC7PezzY5OJisUbmcqaNxvQTTIFXl
hQI+QhKwOEt3k9QuiG1kAj6upK/D8W7hr8cf+xz47xHTBDAgHSx7NzE6QOc7tWuj
hiEYuELkekVgoCZIlVV1V/RhjGDaZuqYzOJJ5Ast4HqATsn7gMrVf+d5FsLH8mQX
NAEdHsy92UkrAb6nb/uXFM2jO/GUeueZn62rEtyO7Lqu0VeL/nTeFrDXAYk/FK62
AEE332hAla9IX2twR8sGNXJjVzTXJi2EFiClEaGoFBVjoDTgnG9jIwb+vmJ6WCB2
A1HxTjgd61XgUWylZoNJmqOfsnxtgH4p6Cvq7btd46t99WLvMqjuqKOwUcW9jHpK
25vczR+sGGXDlVV9QEO+myfd9oChDZVazOwvEYaB8SS6lsWv72eB+bTZ+Zr2b1Rj
C5307NM7FlA0L1ulOwf+DSYtU2AnYCpbqOlNK+lo9wp92flVRGa+YIqBxegbYwWk
MW9WaiIPbPTlaKHNSqnE3cl4TnHvP80bxdMTaTr6uR5ynlcQ0Y0O9NsQDhdtXOCx
MqqelOkoMforI2A8l9DLYpUt6irZXyqiJX+9+7W7GjfG6616fbbG4NnHvuvsWtAz
mOox0ESznQ+jdy3RABRJqxV1lu+T+LWQECE8qsiEE2FcXEJMGv/0+3aZRSJ3HDJj
Lwc3/MZGCI0F1go9ZD3qSNsF8tigS7kXGby/gXAnlfAQtA7UTwDGQL0mJlpeGlFa
ruwTqfo9gkQXzQHzHZhvUdpDsqEgqTrOcXuM6dNzLLqjFJkGkw12mcHEqCxYuYSr
LsBIBdRRK2mFm45O/EI7/0gGfh+82dcfZFfLQshq2RG4TfcYGq4jaG+Z7+m7n+8h
K8ayzuSao9Ua62plsBoUEVr8/mhU2EKMC0/3jZ+2AKO+38mWCvTNEK8KeMExCRyT
Bpq4Rn2P6qlwHtsRn+9jMBFkOrXIF+nJXlKIRb5GQR2zUzuiyyhq9wqNC5wGBZ5m
SaE7Bwobi/8loh7lc6bH/zwEdJdFN4EbpynSBT8/2nMszEh1bPPTf/A/bNMefYqG
Mopefrab+FcofEHn/INVqYcbTN5NPmbjskE2SLNSGH2LaaXMCaK0e/Vh9h9/LQ6i
dkkh0OzGBwkB3VXD4E3oSYO2iFhI5cybJzd70b3DYULopxeoEQXlklFb7wQE7PZx
koKamGM4c5jxdEdf+/LBKLi3+jQ8U3ZJS5CznkEq2ayeOFuoSuvVHk9ylXv1dKRb
C40YbDJ2mtrJocju4RBwT0TZeEwsJ2PH/4MW+Bjr6bXigvgiCNpVMWySSNnhyg0l
ILb2hIfCHYa/7mMpV2SpuFNerKyMeJubrSKQyzFgzNS7tZEEEF6Fg9gex0adUVwm
k77fa7FGjjbkwTUI2/nVPMVjBgEdNi2bCkNgNO9rwDIvJus0AMwpfS09qlg9ciet
gGPyIZxziDK3yYdK1O3+fOZFzO0n40mmMPHuCGYy4xifYISgPqfXy2JSf8c6lC5k
bximKtAaZGB1rCMJnLJw4aLeSgHah3yOXuy6ucxzQcz6peEJ0ZYHIrMYoTQbitRu
bIOz+j0Dfq0rsEvPOlTfamb5rE+izccarITNbO4ZBBLs0WoU8+wmJdvnxlCUCFu3
1J8OCsY6LRbVHc2gmBwwFeE1Rkh2wcMcE/DQdNXaekBAAYC2AnqJJI4KzDTrE/1u
i2Jjcd2lXriElz4XS0FVGbJaxQUngt2f6FT0PcS2Cz+EVi6NAh5+1Do1w1whWNM/
Ub+3UJH44hfYQjQbRNazeykFaxspFFeU8FL7GGRjCT+vH5Bhkr5V4KSlIM9uNFVr
k1gBIDAkssP9Ps8/XHMVAghGegjl3K9N1FjaD0tTpcbDO5/0q4E9w1PYJtV2GYrI
ZH+ej8223UIgtQHQVNORhJ67qoXXPoj9ZWv5OUMTUNx4pePt2uBDjVPtmfzARlxu
OsFzVG7h0Apju48EZ2TBwbiuwHhADcNfA3XrAczmh3ReYMppvQhcIRL00hNSvV5K
MUxXUI/1UVwl1dC7e80bxtNKGDcL26tm8P9ynqNwvvRegKANnWCBERV5IkzSILc3
3u16jx4ymud5sXdhpXhoS0pElX9Ye2hbGCZxSGR+JPn/zcicyRsPfCQs8QVfcqD1
Qm3bs4G1VX+BwuxAWSfL+QrglZ8idTqlHA81eJIKpa30LJbZ1d+fSlG403Or+t/Q
budrHLcOSXRPMGxUR08yy6L5BwlyIT2QvlMd2UDEyZzPnujCSDc5BxeHoDNwunta
dQbdzgTjfhRHkSIIE8FxCzqxnFt+0bNe4hKdHZZ8EvIjfU9qTO5UazwhrtBDqAl5
ZvdMDhcHy1YbozX7SJ4fqS9tHtU8kLr71xHyKIgW+PFO7k0cbgE24dLZTgFQhhCR
B9aSscD7Z2DN9i4Ci7WHiWr1mhFmGo06/Ua0rTkNVWfXTWwapjtZ9dki5QzF8iNr
YZh8e2qE6uzXPuj/01sbJQPNSSGpNx54Z77bY3sERbiXXhplTb1aB5Q83skfg0Ow
u669mhSFTNtnFCI4jJfZlDklsP/3JC5ow+EhsmnGwcmbCcOXTeJHlDwvUxxFHGzc
Kme/5zxNwCuCrGuG7nplWeqNuaS9oqzBvhRg2MbjzAxtiIUDV9irlzBRjItAF6iu
d+S6j29WJx+igwoZfQjd3m4UQgRk48uV+mjrX6CLRA/FbQLbMLo5xnTBrc8IrMzf
PtWs+/GE9uIE/2sVbWlHM4pkSS276B/apHKL5IHzA01dwND4OANP/XgHhpDsJ2GA
dpZ7Swk5Zwu2jN4rnSBInGbb4MeEoYnuRGssP1x0jTxjryK0N7KcZGLnbkSqQIxD
zHkZ8rumDrl229Lfaq7W1KgRhHDi8XVlBIFXagGJji0n0hOKlcoOiwG6PpcDt6xX
ySlfpjjwCMhaB4yPI7nL9ONf++1esJOiYG6kaAI1c89qY6Nzy6LK9rhouh4Kn8fj
PAglQfYJM26wwOvJ8jkCXsfunWz4a/m6n6Buqos6TzGL8iU+k6On6jIzCITWlu2t
IducSmg0AzdIND2zz8IoHRr37YpFrjb8C7dMzxNdBt3LnyZwx/uYEPvxZx7lEpaA
YdoBETX8X+1AkLmnk+QrT37H4iVQcfmp+N92ljzPGrxGrXHq+QU1v2aT8f5YIYL9
brPovKnY7Sj6L3XF0/gRqL4m+3oKk22if8rZbSFQxIecNC4n/hCg4OWhKYAA18yA
htqPynlk+BBKYDhbLtHB8Xf883wTsUeMo8NZFDbVlfxpibninam4+KNGJ4kbO99M
Y831KgX5mo3cisrapDUSvAnFuT8HqG0b4/wEG9d5Lfp2l0NaD55M73Wd2TUnBqT9
tkT24FJyp4KHqGCtOsZoPZCOJFXREdG45jlTtpcgVR85OlS0kbIeQZwDbrKsjmNZ
Ymer7QY2MMMduRNvvb1GEYUReNx70Zk4peuYiF1mQk1nD7/zOxzSpK5ceDhVDpiB
iToFkmRpbOQi4GtnHHL5065iG4a26Rt/IHOJUuBzBCDFbZ+LtrMtGgJmZy5qWkbh
cA1cpevcc0sK7IKOa3vZKIuOETVUKpWHSC2UOarS3vCFn06eCJCMlSSyw9v6yyvt
0B9zOQqxqXh5xr9q0El6zdpNCP/iAVbJ2YKk2pRSnLx/ZY++IeQ1zdCbYcqvfuqt
ZWMYQNVvJwXsWc8iQX1xxzfGf9YH8bq1m+mHyDPqsnkx6GGMXXf51QiSqAgcD+m6
qmfuNfxViNkOyZgYo9VIpdfAXh3aFeSZ0uBRRglko6hCFvwaSvmmvXLRNz98hF2E
Ug0OjSBYvvx7cjUW0F5IimZh7T3QXLPDXKp5OWNL7Q9IMn1VTddrq2A+YKP1sdGC
+ST0sxckyYr84mfV86aFdc+JmOl3XbmXp8itJbGD3PhsHiPNPbNlI0LaTCRuPEZd
yvu8g7zVjlqtkLztp4gWsFDZtYyeRwet49nWP40t+HRG8MG245+cN6OUQF7PnTFO
FINRcIC7E1wL20lTr8FUF2e4ITpUF9iZEp3MRq50OeJOqfqzLLBotweyPHZXU+pm
bG+N6ihr5sENAsNZ5zhAPvastlW4tpMMpEzhgv2GQJma/QwZ0FfQ69GKRwNAuqBL
rhOoL58Uhs85K2SBCtFsiq6/Xyvh6mCyOBttRV9As/d0DNNpq/hEXm9gqT5fZYhh
M/70NrWmVojs2B2lUVJRsJFOU+wveH7xNd10sFRTpgPG9tXMllgwJ/fOyJR4T+2I
scdN/LUZHmjYIUZeh/9NZw+dqDiF/uc3iSzJf0krzjLzhOB8j/WpaqAIob+ydTIK
v+OfofGINUb/f6kZgxWlcFQA+RlXvpZ0ph9aV2cnbXTX38lSS4PL6JwODPUHPf9N
yo9tHH5k42rCaNsEWb/s8nb0b8PGNBekCekkqdpURw0NakiMOfQnRzmrsjSFm3tF
mgAtt/f92Ti8tpWxbq5y7SCXnAsGa3es6CkxOK0TKzXPhinaoKcf/VkOBgL/japw
Fv2ah0+arn17/JJ6QwaAb4GbciHgGsmxdkJrVPMIKUOSBTGLpZ3e2gKJGlgRtYoc
jDpgE1euSoI+8bdtA8U2Zy4n9VNkrUk5hMJaQx44p2OvcBs+XJD3DPL684wWtLpP
/qUvIcIB3U99w+oDQEkWzGswjMfrpEJif5THAkV32h4x74bmBFMPQVE43kiECNQy
N28e7NJXwT1fafIVtgRiZK84GW0GgvVgCGk/HgJSd2aeBuI6EfYt6SDnAoiqmwPl
bRO8hcl0h0TL1kRMfIFbVPuFfSecaTyDBO7vTUIBbCp8GyRcWWrP+/nF9RJJiDcf
JlTzY0aSXnN9Tzgkjo6U8qYzpWMKPoQ4vhgm+3YJ7MCrsFYqpKU1SNh+UZz0Bmyy
4vbtqwlyfzZHl1OpZXTfULA/TemsamZ4y5mOTVCW+p4n1dq4WvpMkxuNQasXMm0A
gP2D2l4pakL7eVdCCkMlQdVtLlKil1kXusc8f+hqBOeubKjOdiCB4Aot7ktbys43
DTqm1Q5q1MeUU2zBFynyLLEsZ8tWWaKlZ199cYE+MS0dPetNOxIchDeo9x+GEpG7
mf0X1KHGrfxvYdacYKJuj6QRltlIkdz5Bmwt8tes1De/8f0dOG4acoOVwJjIS+Dd
ZJ46XyAvtmPniay4t1u5mqZEgfKFWkpXLJb7SgPQ/nqSMRtfUOOBOq2MH7pIEXO0
8z3rQnkIkxD2pGFuZK0WO4xUhn1hedEH+JNcYYi4+Z/QSZuLFedqTK2/Pd+JKcjx
hDmo9MG7L9TesoHG2Qt0RnDxSyjEFN6rSIEaz/ffF3nxSmL7VvQY5NFJ3mgkqxHF
znJRzN7FOqx5q+U3GyPpFnxhBpxdq3oa4pIeF5G4ArQfrRnPT90eIZJDny07M0zf
0iP2VWI3xG9h8JaIzEY7cXSNqgobQHO3Rayrqrlj07NIqbUkWV4+UDzPzvgZcaJt
MaN2Lk3tvIuF+mgk1g3W7+CPH3aUl8rTOmvOipJj8E0K5oXqrlmcTEM4DmC+i4Xy
YrdapcQ6zwyAa/aREsfc7+vmRdhMsp1dYY3qts+yTRjPdJxb81cj3E6ApOHIFzb7
doKeNgv9uiUD4kxMclZpZHcYSo2KD4X167kNgLLwd1Cudh9K5jAFhVsHSs9pG3KY
lD4yuIRTU7aIEY3PLFKs5pu+sKctDkNaqj+eTx0r5iQEiD/lh8+4TqsllylvIpd3
Zo4fE6mHLRL5EAxfSXSt8rxzGw0JoBkEhjpxd/EIZZA0VJD4+MrzvVV1N8p3x0+J
8TjXYtb+F3I12LPokNUVOcAxKlTFe1XcUqZlK9V8zjuTyElhQ02kxdZcW1nFMaSR
cRf0t+0gpmKODW9GCZQUm9IrWrBzzISH/2/ZNvGTHyB9LZqLZngNgAYs0pvM5my+
5VfIec0eGD+PmsuVYcrRec+eA7EIMa3/DG+noTKOMYSZ49MzmJvpGGNREJlwWRRA
GcmpQvig7W1myPGsxvu7hDDZQu+RYjoifUHLTye01U3PPYZw0QlMQr5DwA6xU8Gc
WEMCmoGvYb1igRJZPudedGny9pFJv0chBgGmSBtdLoYEvn32ZAQ64HjbRypK8cUj
uhbNPL3zItVpMLIK8JkjXY/BwKR2PBEZ/obQ3/bJ8Ut9MdObamy83/Tb8CYby/CD
9G682zw7pCaUl46RDHDEylY4jU9xNkThf+GwPGu4RKDeOFwaMmoU38rAT+0TSluX
Tdms7Ht/BeQoBSZcMhGWeVzuibqLex/DCokIzkUeWvikTNmPcirtPsyV/su/ohrC
SjkhQtrohPb1RPVec/f4DuNRx+EdLMdN2y5INdRmUS8jb0k64/+B00HH93C1132z
KvuMXn2uGGLo8eac6c840ejM6cElOYqtf0NEa0xS1QQOTalJGCV7QgdMxvT7J/er
Xup0GHHxsdthx1RZ9Zltrh6A/gr+KBaW3vBhPZhoB3OSdKi0xJo+RfzHCD/AyPzC
90yOWTuBFamnNBiX0B8RfEoxjl00C/l0G8J0q4IYZbaPum2TFkhlF4TnT3MPt89s
vCGWiNmbvi+bisJP2gRm2PrK+ZI+nMErylE/GTMWKx+aV4N2fq90KE97jKFoZAPP
KOv8nID6LZaPnU6ujIN5+V2DOCK8aA+jfmIvTz+kk/8lJZMWWPr83HXv3eU6IRP1
/KdJCD2eLXN6u1gIKrP9aSymqk2CX+8eFvgYhdbTFJ7d9Zz+jXvB80hgImtCzaip
2SyxJDXHJJr6/a3F4P3+UsSPG9Kpn/ArAO8blyQn6MQROH6kpYzLqiNYy5UE/KJy
FHTjh4RTIPneFDfsa49s4prQCR35GkbPZTKk3jZiBApQvRGzH8BKP3MpwU/a0DzF
FJGJXthIjU1v2jsjbSkrwo2+P/1Zs0+6bbKwMDSiaeGRFv8YPRuliOEX/LtU+aBB
8SakLvyAiF3jZCLQ0os5ewNLRRHmDZUN5K4chCfuWqLPzE+Vcx0cnNO6FCTMOU48
+R1ORuvjOzyENwYWmPNOq+BZvK3UFRXR5IfDrWrptFfUqVckcB25e+8wXke9Po6z
eIlq75xBmNYyH8VnmKoRtAZ/nD2k7cbyeD0EgBi6al/JIR2F8N0fq0nU+6iwt36K
mEQzSMuaWSYcUa62/7oM2gKEVUkdDYsmF7XfRBRtRp8fzNhmllB4SfqCtaRaA0WZ
Fv3yp7glOdKtR30vFkXsmv8jOBrJHLSITNeqC5hWxsSKs06OGndeSAUpao1q5kDc
JfgtcQwsoGLIM6lipx33lXns3i1UTFQPOMqUWIpr+PUbq55prNDJpvAu+D7JmSQ2
B7yvFkLJNzAdSrMhifviF0bAHV636R3qa+goC1fHElmAUToSlwRMxX8/wM/sfo7u
mjIFDQO7kbbRWgShi0gTmDxI4FWzV/f2g1EUsaXlerB2P3aMYTvRtYWiLiOEaSva
QVkvSecWeaB/z4yew21tvkGKDyIU8LVUvP/fuzHfsb4jKeLG0TBM3JQKjsA9b8rl
LKUq/9aKnNkQfNXMVrsAkJ+uyP3P8R4JCiU2dY9SNy8epwyVeClZonG7ErcxSoSM
uS3KM2s/Lv4m/0H0WYti0LXUD2M9XXZajvV7/b2AgP5h/1dkkawLk0lS+g9pgK2S
AJv6pYzt2XC6fi0z6yyYcmnltpzWINNmawAFwOFbu6hHpUHpHlGiN6/1PX8PARJU
AgUlk8GbuDSRI4lPhwsBDCnz3JWQo/yMD+35KNXcyC6BYSNhPNO5bf+ZvMEVZi9r
A6qoFh7wabepFonCyW0MYvkw8mcVJb/0TKwd05PA0AXRpg88FFDUdLAaDsp3oVy7
ddzBJbRsrn1Ux70JclS52drKVCPovzfcktiiGN0nixnfzhS65R4AyPyXWaK6/maE
BQDPNqqV2io7j6BJOofsH+vHZhn4D/8iODaoyvPgMzvua9qJf2aD6DuCfbNkyCPU
i5b+Jzm0BZa62VoT4gS3kOzey7OwGmyi9YhRNRzMKkygPke1euY6uImMlwj+QEK9
TuxJtT/uZCSO4sl/Fe+MQhdFRUamkmAixez7Bz0L9+VmowkaiPjWxC68PMzs6pZn
x1T7c+l0nQNzsz5lX7K1IsIkQY7/ug5/LbLBdXDs6rLaTqxg86OZ01Tknh1g5DaZ
TlxvQh4ooiwVLzx1Ut+mFU1rtPwckBVJ/yrPSs7D43E+xqbIoSiQLiAXMIjgzk/u
Vtz+PSWmeg4qhYpbqrQZHZnsnHEseaLHTZt0FBdwgasmIFdY7z/KWlAUt/G0/bCG
pEux1bSYRKf19CExUPCgusmyAkXE4+4d4yF8PcPDSII+/3t0gAQGZ0IaG5Q3OUIB
hF7g/FzH2CdqwCzBFv8zT0lFt8bG3jReXoM0+N7zj+bpCnK7O1kCSNJWM8sEndlZ
HZ1umxBdicnpQVgCPHCtVHG7Yataneaooepfx5NHQSxImqexGCzujLZPDy6+HXgy
9BE0XLo2CXwcjoGekNXkcOJfKELliR4gKux7UY7AemdjtO7d/QJUrsbC+c0O8ioz
68VZNlt2ImDdZd+7O5x/sutp9BaR8vRxJ/050PwfRn0MO4zWBPJKmAcayHRTaJt0
zPOY+Q07bjOE23CltLdeBQ8D71zJ/qVr9Kj3xlVIDFC1YDBisuyos7ac0CDMFIm8
Ys1mL/0TT2qKRzvKoycFlvBMXkYREzgCMVNBUcwufKIlDzKyQHeyyZlrCNOjZ1Vv
7Ld2y+xPB2bx16kiKrVObvViEqkJOVloMS1b5dfhbaYlXqaNpFgxmKdiSZMAEDeF
yPg+CKwIgD0dzVk/RDMWA2D9jAqOcDv5iOaGh2g0cfOttxJoFZ7iDhV/wu5lpgK1
mr5HlPID4NBoZknXsTVzI+peCv1lUTOYthT4pNPWqHHd8x4Tx/sG9gMcI7rwV9JV
7Pfl7JoqnlfV3tUG2IWCJAaQrqbyWqGnCNWFImLY9l0v1y+h76cj1qseh6xE61oG
DlLHs2yZ5HJszwjRWmqIes4ra9xnGtSOacSe+Km+MrdpmNS92KXLe4Ui5kvNhgfc
Yw64VMtQQQxpqlNaE1YmzCUrNQy/5enCOfu8Bo1CcRFGcZSrXmQyy/lb21P/65hM
KOotEgbJq161aEY9k+q7ZMSIo/KYUuWE1176C20jL+PQINz5Pph8nKBHIaE6CKiQ
Y9VS99Im3utyUBxAfMKN5vVP46LVmlgr/b3ycaFKjAmZtPGxiHYgstEMqxV9cznk
qkr63G1qg04AQfKnXWI48YX4O7sPJeGkAl4tzHWXXlfT8zqKDas/cu2qFB+h1ZSE
0VNihaFmuvBAOy1oIjxwKyWLePMgZl21eZzGEpqZ2gA4leT43NZYlPsRhSjq8Kkm
o+mDNeQ+Q94xSt4/csBFV3IehXP6xv1GNXiw7yuJjthzD65jkVTZaPhIRCoYfYb+
hU04dTC3dW8MeYsuTRYSLhUX4QLc/cxfWnUnGxqRlmXWFrGhJ68h3VDlK5h3WxpS
Sbr1AKSyi77bOVIomdQII1iACPmT9W+WhfyBCeJUEgnKY6k4NipUB4HlkmuXEIum
HMk6F1/HcN6Sw/o+lr5Gk8d8A5sL6QJfBULlsR93g5oCoQDI6UtN3+943jgbr2PK
TjEgSf7BS0uNiTutCfvRaObAagPpd9K0sEW3yJJxrtNykomuRGPzK5XeFKC6srsQ
NyMXwC6O4YPPUtUe2wBanHfhGbsO+FtdCj+uT00meypT16NbN/9qaxqXY+plx/xX
fmyKdeAL5dYQXEq68UulbXCA10/iMtbn06k2N4aUl5jX/Jj6wkMJjjzjdbULGdAS
r40KzpsUoKBwD5F6H1nWWBNaOvvaVFaHNIVd3dP/2pE4MTRR7poUpwt+dQ60lQWD
lXtlvgZbdlUQmrXR3RehzxAWBTuXgH+m1AkLqVJuCU1ER0LI1ahVzIs4tOLKknYo
cmq656nd9Fr2YJREDr7lLcRudUbO/SJBmuYAVx2PcFCjd92U/8kIExsOxGb2wgN8
FUipdLjUKEfVaO3n7sk3PpjqGAh12MZtyWQmcHC7ZgzriKGC/UX9G6D0YkwE2BBU
5w5BWp2QxgAFpJVsJ12XB0FChj80+1qrBUgsyTiBr3ytLjA0NNAkZTWQm+l00zan
E4DTUi9cBh8XFF9snfbbU+UWewoQYpez3GECZppl+LEH/08PG8+hdoySbwIMwBcQ
wvc4ugKErUAF0MpyIUKblw2EtKQh7jR3I0HKscVgNT7Y2124QwknEJhyCNIHPXJx
06Xh16SM0wJNqI4Wbn5Q6x5JCn44aTmgHn7C3tY9G0r1O03/uVjJHZi0YJK4Sa/e
yQxCUaezlxzBd1m7+eMutVv5jn0VMtpvZkDjoN7De5gChL0zNNrnjr/+NNtJVRJd
oBIM/ezl8E6DZGilGM0WjcY8Q2HJYN9HZRy5uAJduNTgDU87vouqRYwm8/CtaMVJ
yGNwVD566xrUPcZxKbe0nhwKVGwtM3TaioI9pERaEABChMCnYaA1tUbXcPXmHEPQ
+/3TNt/6HWNqtIbwhaASvTSur70lOfvgUImz3twHDFa0bTTcNI2vzUHhHL8BmWGv
6v9DtYLeiQPPgUxOJvfW0TZ/ff500HDUd4nvspdkeAPWxmXTz3l8n8yKKDLSFhJN
Hk1RkdLwVoNJwXrxQR1OfqpjaXpZYCeB1vrcldFX1k8hrtOLgmU9pj9+7KKtxqL2
P+QI9b4Rzh3hDZVzStxsDb8xTgm7LDVJbPzJcD3pVZBdYVh2Smm0XCe8SyHR39oM
mylzzfTjVTUbEg5QfZ5SgAVpcKCwe7NCrnmyKRX0YD6xlBTdPr0mVBRYXhnaf2A3
2d3YuzAONkS4trfpxEiGBFcSX0YqtVONI4YXRwmcoE5av8loHs7hdqK8nTvkfJw5
d4IdTdqAUuEdpfLlT5/0NFlEYhkyNehwUERbal/9U/H2Fw0hnEVxqY51CGvkB+S1
V5Mx2TDS7/5JJr0d5iGHACzYLOG4fqh8ymjF0Br7AYWDXPPYcCEwBj37gB/R0lF+
JE5VpiECR3RejYZtk58e0kVkjcM0VUFnoAFUdr8lxW0i61yNBz68epuxRPzqcfMu
TqpJFcJP3FNtLcHpaXTXiOkiRiCHZyb+oQHsq0TdL3tY1uCGzoM9iaGaAJeIx9Um
BtIih7J8H7MhtdLqy1Vs2L/Hv3cTo5SJQvYplzBv6LnqM9fUEgeAmdjnXPpjWklg
SUwBosqvJf33CkasT7Pvb9pnSgLhvaRQ2mQ6LULQzCVhWay2MU70/BRoRRfMT8y8
4So0hBooMeZB3ph8cTKN6z011CtqRSO/tBDMdvr2c7uJGPo0x1LcKdGqd6dQpqWc
rsHQuUteDntrLRkzg1USuLdvs9MQDwtnNiEeanhd+ksZP/5j3/qZ8C0OR8/CgF+q
7Vaxh6T3l3NFcJCWpvBvcv40mKfp6J4m2PY7xjxyyf2L0wKgThErCZx7j9+iJFkM
txYhTM1S3+19XqhXR630UnJ8Cb4yYdOK6nwyWpXC8AEL7Bc6C/RWzY2JLdPnESk1
jHCRImA+jsKwr+KfOi0A18axmdsR88+TQFY8Z6KKPZJg6otH29VVL86Xve4Kxi0/
jIj6gkStslB7Vv2Dg+KM7rUwQea9EQLbSh0g6JNPPcRjM9T8RodHmP6cHoTrnnH+
y8NVPuikOVmcH5QZjLCW6Iq4r48qDMEMbZjJkxZUyIYBOxGdCjl0QYTgheQ6skWV
eR7L2OEFBMKB0vPp4JJGvEw5oXY9Pvuf5X+egtdS9w0ubBJiRFb0lCF8ONbc20MM
XBCEAxa070LdcikXQK5IveJsIT0Q06ib1s/yBmDebIIxfokK+2SvSj6Pm3loM886
pQdAsGMmGt8YIKCrG+Y1H2lTQxALjaBypnc8sVoO2lR/OBpF7a7fDv4oY0syM5Oi
+NXovy37T26SbqvZAH725UAfK7OknZDkhfl8eHq4eYs2zhy5OYsBD278UHgfvep9
uSy3NTvxJnvYJ/UA1zHA5RnCu/qD5+ilwGHbkZw0vOGaPylys94462tpLlWbsbiE
2REkk0hCGwapqI/EvoL4sEmOhmpiYbCmoI2CQ2TebPb5rD39us9lBrUKgXYgyaBC
CdTpwDGzSJ9TA+kB0erAtS7zKDw7yQFhrPc2eY8Nm6ngrNqNCtkmzhxx3uUDeYdy
QoH/gtICKC4lA0c4fwfJfhf93Szuzk1eSN34nXZ1yqApwsFQV4OUEWA4WfeLshD8
JT3qMZPAxZ/IbBHt5ny0a2VIAd1aJYEHdPT6IMyisCW7UtrCMbACEUdk+AG/5wgr
4dr7C0E4at8+uWmObjmEcWV3BH3mgBsBXI14/i8NiNgB37EK0rWoEnq1YghhbCDU
Ud4t/Z5gmKSoA9YHG6gNTpkXw0pKpaLJekhnrFeEOcV+uy0C3ZWOyHae9BB2DNYS
3LWndNKIGeOtMcenhFNR91vI62hgsbApBmkwEv8X8XmHP5q67KFeGM73/QM/PCqn
7BwfEfxyzxXLwToEfRbwAN7odaIfGlcRlLlrrG4ylZg3wmiHEIsYdGxROEV46Hd2
z1x0Qay+rPYRjZbX/ePywsEo+uplvS6F2zLPIPKbSDW+oETVJUfRhZRSZDgpqe0y
o0L4wdn9dYaxgAzqBy91+w+5k/mkKIJDotJQnJ75nbSo/G1g9cmvTqS5iZR4b+Uf
mLyrmq1GlfLTwW+DqOtnDM7jIU+1/u5ggxjXNRxy3hj+Kj4OynaauPqeywepLesR
v6jXYvz9Dk4KUwY+BP71XOc321vzd+vvAGdWi3sGtJbVdzImgJwUgGqI18sYRwrh
Hg3iDiX7XleOCWQRxEjYMSn8fwDsEQC85poP6T+ifW4XL8He/ssnF0PfaQNlaQiK
JMg3pihkl7diKR/gGo4R1NmY6P6RhmD82KuItxklEAqt9LGGVZnVbyy6PvoAVyI1
Zyn+TsL2xokncuYtwjVph9EuFzqUGKE4FfV06cYsKzUZiP/Lt2jPkQOS1SNRc4y0
cSH8oFhiYKKmn13CRNKPKDthDiLFxTgFJAP58n/mSBU3cFluxB3yFYVEdQfBlVY5
CXj3g2JOMo4b/WcJo1jBSjFr77oCrlxxMe7puciuekFQsBE3yGti60PYnZJdB6PY
O1BjTg5Q+/XpRWOxAMCwdpEujayzIrfHD+8xFli8JZq292QCa6ayRyyDj7Al9WHz
WGVsPD105nFUR7ojF/Uw7Js5875Lc/UofpIFkrSqksPsDTJyqjJgG51WVBl5BN2h
KF+Jux4iD99U/NheY0jOWEdCxz0YsTLb6EcWRIeNEUmkHUXwALznrYDy2FkTgMP5
YJIavoa4F2qJKucMK6LXUBxpKcozYdiEeuOhfRmb86CzFbas/K2zphRw/FB+M9sk
K13PyqJkbnQoOFedUuzI/6sGTrQQAIRolIeDe990NeoxiAokcOPs4Cgn728VC2i6
kpXDeCQGshVJpeN2IdL2Ppbbru/wvSIWJ2+ee+s+4n4EiTNXl51qlrs9eO0qr4NU
69bEHPvMhYxTcayOfOSUqfPJtDhg73MRd38HEdSsVOgZD6vddCsYC9qiH2BssQfq
pH/2u+E1CkgcSRvTm2qwmMtpBQQPAm69njkzgNbFI+zGeCHW+mWjrMD9Ur18x8u1
VMWUEzLD00/lAP1USnr8fI8DX4ft3zBCPMmQ/oQ3ecdp+S9ROyRuXsQeGrpG1DCk
hjxyIFrKO/ee8ZR61J8ECFuI02OLw3siIeZa66e/WkWAiXDGaPKeZwudVglUT7TJ
WCG7CK6X2xSSlT9B/OEWSocG0iRJHd2KZMa7GPv+nX61Xz8LiBK1HoITC30ov/mt
krWrTTcOZ9U5Vi7yCJGGH0e9i4NeRsR11p7a7E5iI8PJCokusPQOt2LUNrXmGj5t
oX7bSgtPhglT6eFfVKmWQzzv3f08dLHHRpZfjEUQzRH0UbJK7cp4Dsoehl3fwHUW
bn7Swo4ssN1xP2agPpzQRggCe7W/4EmucS24BrFkIa2BOzAkfKo4w7tA9OAWEr0r
oYK1nFo1PhDrMjuGsVuzeFaLTdQveRQMm42NIPtbXSm2YTg/nzi5BKj+8MMqy8OX
qmmRfy4hf9tD6sWiHiUE3mhBz/lREPBCxvugcvsMsg4VUCqiB2zWufletTo5wggG
Tg9t2V/Ut8iaj9BEcbOyF/cIcoE5NV37vOgLh1bkf3GXGqzrNvm29tFS0AQjP19r
8fQC/Um+WFONAaNe0Y889Z4lQO5/kRr9xRzzmhRAAi8t7fjvOhMwTfHWXDDgfBXs
cu1Xx7FWMYzlS1k/krKT/r6BcWXMm4pcjr2q5AjZKd56ykP0q3MHdQdAYt+/nVgq
AAYlvGXNwKuOl2n1pIj8V/HZxUsJhzQgaE/B3lJJw9BmXU9K2oLP+xK91aMNmGKZ
nB6JIIJZ7AOQMVTBjQMOJZpDILAOoiIoTJhnI1kqzc2QlUkaSYFz6uFlXrgRVufe
1G47NTxis5GonpjYXX2LOMmk017SZEX12LVgrNMsXGkKIlBbp/fxgipNDyyT6ykt
DBbe95Wki0gsrD9ky2dra7tLAsKTxxTnUdL7vC79T9D7LCCD2gK0r3rAGIIUVDF3
LdjR2Wj8DmEH80WbTWlxJKzz9sVBHwVKpQSFrRzaA/RfCSN4wqDIZZAWkAXByfCE
kwCBa8ZBx/oXe4nHUFnmTO0pcUjBxbDT7xQTl8LFj+9oleHUhQBIUtYvr1Oh1EiE
4zVfhUV5NCi4dgnUiwuG8Jh8xkcZejZ3bQm9Lf872lFK7fUQLTxKSXAf8pofTPZ8
420DnvD1Uj9jJfJ8xNT/dTYAdeULuA2EDd1RJ03imMGj99kMSM7+gEb5U94EGW5h
Ii0MGmvuQGYFfTRqLTO9Lmef+lAUDvS2NIA8Srh4Yy/cnFTy1EW0L+dzFsVVPEe3
qyqKnxHWQRPT81GL6dhR0/3bAXqAMjBZpglLKfmX0J5R345yvatUedDkTuuzBK3m
kIF8k+uOATUGoTO56RJ1ymCZEXLlwJ+j9aAHmbx8C6Qt8FhV+8WgpeSL0tn9xiWW
bQOBoql3SX/vKsyT4L0IjbvqvyBI5191mXYPxKAPyCqo6RN0Cw4r2T8mjXCfKg8C
EVNmrnHOoN9HXAJKGnqU0sk0KjU6mHxjVn2S/tvgbZan2dHMpY3K9QlsT4BAlpQn
I124gPs4zE4GWvV1tkNFLXV2aULVfa0M/tiBac1X4z7oPdb9pXdqgyAM5o+Oq8YW
nvUeU4lpTvePgB/44GU9ju5ANol1H6WvemB15SwuQEr21PbuABHKM3LIiNvtKM5j
kwl6i1rGMM6Z8Y8MgKWVxGhRqFQbSaY0qoRdnMSun4YvYaeARkP5ugtVO0MroFVc
FO/uBNTvmPk4lX2l2+LAZx50i5OlsKwR4/i34hLUo0maaW4AmVWBOO+igFTHrI2g
TOvV/rxisqGAllX30RCZyk81re7UIeycCTvkydVJ7YbrMguvnr+Q3ap3DS5h9H/l
Wf9Ly8xtssj1y6wrhGSKw0gnuCkcdOM3pBJK5vEWkbOJCGmwERDG6hvNu932iZTG
L/+dAGzb1P7gmoIyWWcRqWj8eFe8Yv0EOUj5KjFd+gWGbFh6fmyTywxFBJU0O3W0
CUR3ivwTbTuTS07ErgSl3Fx+qOnSqjyiI9m17JL17QnZKXmZ9tmWivDSWbZe9PFK
wAUJ5huvACXAh971m6e51WbOKAgMCiHvs7K77p59V5cy0JwIywXjcsJRH580Anuh
tX9pA8t9iapl03Xcg7t64U3kfmF6DPPDdveBQnFk4APZKDI1XC/MHiInLBEQmMXq
LNyOcmPFKjFCZhfwAXYdRAKO5lG1zWK2VI5Hwg1EH6f7gKUiNJ2te8jV+0IVAMCR
AnSPcDakcv5S0oq4mWGJuQW0RH9jpD8HYkhgU1ksOFVH6e1L5xSpvUkOPwJ5fA61
CNGZAevvgT3UxJ11YsdVwaZUjwkVBCBGQxihwgM1NjeEAb60NuSBIWt/cVMr+s1n
Q9Xb6Wsizi4iL7W0k9EI3Gsji4KaCgrjO6DVeyClEdKmNQjn0pSIAcFg955fi2oo
caFcRTs3OBP7HgARWpLRAH//0WdDmv+71CKKhWub58WBVOwpfaDOAPMKDdN6IJnM
eXZ7QjnAkftH+ZKPNnSinQ0IerNRH1yLTOrkbVM3jtHwf0eAIGabnuf2XM3R7Loa
c4S3LKA9ZxxQVbRWjxAFKSUDeOvrXl2sJe2RtihAYT8qgDS443AEJQK8BHmPzVcd
KjXR2labRWLZKov041FCxCBd56dSe0wvdJ+E0oD8xfavhD8TcqpliGnEZCGBInrS
7QLqJAGsjtOqaFcQgXUGL6onn4bgg5Jr9I/e58JKnfevQ777HS1zXsyf1DP3Nnjd
nGNISW/SM+t9SYUFXpXmHGIHctjf3qDxA+QlkDriX8hgHdo1zxcjLy4bNB+/81Wk
IqNPnWL08cWgd0szZxAGtdv+W6pMrGFvUgVZhdY0uYwN9WS8j8XmIMh0AA5zHv+z
1jNC+IbBTbvy4uWCU1eAB1281MAXNYjaI+RMpRayiUQUiIsB/q47xtrK0clgX3wa
aEEutLbYt3aYfIuLRdIuZQkI+rdfsA+IrnkTy5svPANksHo6PN6DkTdOUsc5JZHi
YK1CUwsa1tqu2+mcR7uM3agxWq/nmYrIES9FWuM7j3IcKZXqRXtcK3L77ZgAjLGQ
s0YFvY88AcbIy4nfPUV/qLOoUIulxTh0cKkQseHcMYPRJbNhkbRr5mV3VCrYiqWx
7JcE/M/xYvW4HzLKTszxLGq7kLjiIWkpPCwEgnvSpgxf3nVpUGLVqxVTF5q+rh6d
ReAiFiPp6Zmn5cL/gsVCgadcf5qp6ExCGByCZtq/kycN5ELjsPqx7IJ8WmDqT2Kp
gXi8oKMl7S5Mmcwt9Nqe9/+OgKF7ZdFbxVTZ0tSWwEPPHojtY9ie6NFi4lahB8G+
CU/DSOvRguQZU+1VwngglLGgjPfeHjpI7HauWR2IexHhwroV2H2oyz9bospWei9n
9++EIoWLKjnlKvFb2mCWV6tUIJcb2oCTaPOCL8nO3kOqrpbbUAqTsscu5JWnHzgG
2hwM39ATzGXQUJrCJJ0DnMkUkNtLbQxih6LHIJhoQdcJoRejTHXmjaJbTMLZHNw+
pR5GH2gsFwQs01KuKFitHjYQfYRRjUUTp3nBeK1gxPriCALt+CUT0MRGUxOXyJ/K
jeEPLLF9u4cVye6OkdZ4/lfe45lPJMPtmqqteke5xer5pUfe05wbzVkCPtZVC0I/
XFoi6FqFMbge3/tTGFFxOu4l6zAMxDieSRWhKP4Wy0Y2MUi3PvcHYEx7b1psuQw6
Z9qFiw5NZVN+6NtGhdFZC50Jv2WjLFNr6htj0WDPRNaX1fhmJzkYVtnJKZGZp3vs
OM8oBg789a0oGT1QWgE/d+woIcejy1S1kQ/o9QPbu+iaVaIkHnMfGYs0wWxdpPFB
l3t2kJ9vTEr1yRj4uMje9k37WEmc2QRxkXbVgZjVfvlA5fq86o8N6IYPtuy0NImF
FoRFOOnd3UAZgSIV1FIOEzHEwd8NaRNidt0qHyIJkcaSiUTUZlDxTDhjbTL2NJ9R
PENPV+rdF+mJEvTMVBGdKbS8HQQIPxLePUcVvc0LQM4jY7AQ0W1DIrkeE9XjJdyE
WJTyJbHgRALqeh6+/mTt+oabMr2CoQ2UBB6J44cVgc8b/eyXzts8DOzU+NVxj19w
NUxy4c8bRg926s/dB+rBFn2YVZqLeZ0SGEscfxa/secxDvuAOwE+82Rij0ygOyDb
d17OK3JYj8ERHx7pKUdpM1awynAtRqqly4Bq7ZILh5KuaUFj4moAmXlVoWPljeou
+EVzbqcfeDSDJ8iRCSn85ZckH8nGew2TyA4TqBe7Kva2+IfSqwU2Q0Z3S7vsP72v
A3PIbeRw8caU7axjIHiw4Mj9nj1th1MUjxvI6RquAmHTSQZSYdavS1dtqoSAy3qX
dizkVvt066tRiwFVNJdLNoQ/bqScAA4uKDsz4v0xxbXz0ZmGSNkNaqC8dTTtl3cW
C07Ev9T3jFSg8/1QXIY/Lw986cYTUe1WJ8A+jLk54bgIdxmHhBI/7EPCYRIihgV7
Z6OmXR7Kl9QVTI+nBi+3TrgM1tF0sX1rbxn3vjV59Bz7ScxwnbGFuKq+iLKremCC
+LfAznuQsjcARdQQ3+yIDevmBUd/aznlVXZDO3/2EWbTkqePhzmxK4+B+pAvekuw
zSH8ICQtq60/fcSNmLaSDw69CqC5IXBbWxD/Mds3Wu9ouhCEFGbO8C2WzBodWnhL
hq2O5kiHRl25/f5BGE8ErM3CAGUoV/0OejbRuDzLUV+T8r7vZDDHWAjPARSD3McN
jWcpvJqwumiUP/UJLMBuK+mGkoUqDg2SJbnVA2RSTZ+hPUWXan3gZBIGXB7zJUa5
cbXKvcxzPXRunoEX2sg2kw0zcKB7L4QIcPQUAWDzbFNeapq6awKn1WjDCWDYjWnp
oV+aw71E8yx7Z+jmqYKvHw0ifJ4fPhCj+CJPhoCMFEmBKE015TyMj6NX89eZZVL7
bjBZNxq2B/ldQx17WyKDNGOLXRmwvVqSD8NzC/ztb4/+I/0Wx8samdc5nJJKkQVj
eV6rddI22QGaovt5ultY2kxVKv6uQNW2a1rWIVAJ42EW4mDz0lQ5HKd1WiOiF67s
A/AkoOCUwW24xpKRuHUF8WK728Ec5p7LGHW8J1pO9dQJVs8w+WG+pyMJGy6KfoMv
YaJdT9cg/mURAsi590hhPfi7O4KtmG8HBpvUc13D6KvNXunWs2NezE3jq6IrB4En
7Roj9rnxjbIVDldbzo2yhGJKvlbqosuNpfMBckcHViSirSsMclNbLSpM74akRJul
UT4nz0oY18pzeK7xjZ5iVj+YfhWKZO1ii3WJnunDEMNj/JPVL0RGzrFanZN6lY9w
rTCkVfRwP55D5yrgCl8WOoXph8Gz1fY5LCzo67A1KrQPVuQGmTDCifPMRUrZIM/D
B1A2OxBjOPONNwgOSFR++ieMEnnVJE/mVHQ/Gz1C9EC+G1RFogEiY3Ys2Usvf5vY
wn40kQrikHHH0eOLDEgRoqpKNy5rRm+4xHXD7uJjMNs7zm5aJe2sTpbjoJ+hHCQY
S/xMV8DJ0QtlQP5HA1sBAcF6ChiW/9LeE9cS/se6BQFASaaqtHuqJlYZRDFnvFfd
AlfvQX+ALVnLjm3g7IYIdI5FNBDJRPakAhiXFPRcAAeWCUdTAUdnGq5QWWAIb7OO
QKVC9CVsFu+w6543q0xnz+yK6whzzkh540VIp4HDbVZPId6x1IbwTFKSIzFbDMKG
c2h/NZb0nBNK1xxtC+z7HzIfclaGSE995PMO3UwhKFKdYtAJJr/fYnfjbFZgHE4b
zshZuvajmgvHmoICEO0JD+EPZ0ruItABC7vl0MsdFIoWjy7U/5hmZeV3EBO6Ea+c
2OUAQ4Z+qoRZgVPFpiZxmKdUobQmtF+RlAPtfodrQcJSJdWddy3F0kac42koICnY
h+6w39GL+CToxA56c6uM83I+arr0Ywlft6ldDav4d1HGHFYVxNtbEV4ei84dBHzI
a2/C01L3a6fy1ASWXEl+CiUXDrr6lDrLJUk/9i2eWRbyGGt8zOln3IwA2TixEG0b
vcfIfKnVNDSBUJxNXLJRLojcmvU2A4wr4SKL7uM9znNRSwryvFYVefaHjp1Kiwt8
TqIWX2qlm/SSAX+1SM/lmgtI6tmqaHw+IXle5w+KeVKsdne5alNcfKZk9IQQdg4t
LL71PW/4NHpXXbYMi4A0kAbv227dqiYs3cHY1kBze/VWPM6Q7ctjBtHyKG5sZA71
9qTC1AUPqqjmxbAOd7CMhXFFCC5nTGNAqUe0B50pzALXXs6GhcjGUQN9fnR54EZH
vdIe7bJ7dbpXgwHy9afe6WCJFNLiLqIAiCP8se1Ixbm4U+xU0/q5TXl6PY0xRwEu
dzkUMF7khaxEwte8a1tzXF4tV2N34Zm2HbmBv6t201UrNDaKulYI8wQSuWtAPlBZ
hCuHhi9Q28NPokK7qko6pmUFBTXUNDekTzS8p69tnjFlIwNsnuyMrQ2F40GxNLOT
hp8C04vPmvGjBMYVNJS9TyhCKMTEZoefmbLOLxpssnnuIkKto0tR3lVhQT39m6VO
ui9FCJUrN2Ogzg6IR9IRuTmTVFkQE/qHiHqMxceOIA5oC43fuVAKlKvGwpkdxyL8
tbsrWmLVmxri6NpULCK36mYLeGw95Tmv8t4lCO72Li/5GnHhTy13VDhbZlGU0DsV
beK//mjMKPo3a8QprYo4qMG9MeooPlJU5CO2FKVjWtnqaXkyE/BX2GFvMa8V7SXX
a2zivY87PQifZPPYnehVD16NnPm+UXIyhGBkTJWrUDDV3Bu/qivJGjxBRUBBC90J
6USRjdR7PPv70mK4BZwHv4At4vW5nJJpGSXsyuweq8QyH9jMWsUKLxp/ARiCj0LF
0TYGeQnPr1yKHn4bMdEUvYJViSTHZz4/o7VU3E69FRDAHscsuVV0mGZ95tGtuAh/
6KUeQmL1VfVhOiz0u+91MRPX3aQFpwP/PSHkeH10SnoRKI2zCFpenhNBxFzVQTxC
WLsl4delxGckLqKL5DGGDHzN7YaHAcEDT3DeyDl5GggkLs2X4lJ7trYWonw8IVXW
yJhC+1NN7B3tx4ImdbpEduCIdgB2r33wDDeRjrevpkpMLd+lF6u2DFNJby7iQmkv
55d61EFWscbzc5bXtUc0nvt4FFWtyQ2YkaXg29yeDQPXxR3pkaXfio3qvZWaUuMk
49b0YOazeNJyejZEcsP095XcdOp9rGcDtCFQkjxfsHkTUXwxzL5zvxsrZIjp8yEr
I0d7KfKVZBzfsxOTqeqtWpFDmbPsSSE+p8a6k/5mIl7sV2omoT973OBi30yTk4+s
prEUn99tLCl2eyi9sk1kIXJavDhIbLaOPFCulT3tTQtAGakdLB+B7Yh/4sUwPrsc
/bYoSeEprkgjG9+QhMpc8rdiZGUJ2CBoNR4/7elYDWKmpMXRV+P4yRMZD2yMeVbo
bBeqmVs+e0OXTEHGPlLB1E0DVuCThgg0WxViD96PpJfyE/MZ4bjXJsdtWb+mt76o
5F0sZ/1YB2EM83LuOg6obB8BG3p4SynFBKYTjXtHqvqPMGFVr1B8DqXDbx4F+8rZ
qYXihGzCRzo146Pa5C362JVC3u7RspJDgupcBXq5/o4U+LaHaPM0BYyC5pzNJ9Q2
BPiMVf7vLT9abWN3J8jRwVirzN9meB6OG588FM5YaI8TqPk4wnL3e5n7WyvJZSmL
Rv8KZ5Nxv0WoIblI6ZJGecq6BGHdQ8h0xYGa2ze0HhBwerGKfPpsNAacx/BksJLr
eqpIx0fSkX8sBKc3B1v8Tldcyqtwd5q3BVdt8uzTX62RvCkYrpo84S3pHL+XFnoA
sEnhwJEx4vlb62KjKtcRPp1NnJwi0kg3buscfq2xVG78JdSIJIarBiH/1kzoKGjH
XhhFmwjalX9KVMu1Kt14YLl86YD62Ew8gdarRXzPeXh5Xr01m1kxP0HQ4m2d4UOy
xYKH1lYLZ9vkuj6GnckkuNNsYz/JSRBTX73wOjDlnINmoLnxKV5Bb0HPwQDEYdkZ
uEbIipYL4bB2T3Iyb9RHeUCClrX9RleQB86z95cEg7jEsRXHwBbuu1PoxY3x4ktz
1TY9kSWfSShT863NrlNyFA7U2obcjtSTCtTTDjc+KsDla36aRmD86Ilet/w+LWiE
NLC0rLdlMCWS9ILZbrP8t1WQhLCYCwQA4iVUrBoQ9A8ISU7WN0dz/MZjstr3qvxp
juAu+GUdWGJOIuDi87rTLorsBNh/yrO+ti7IqDzalJo9+WqkjGom/KThpk23oqU2
PmCapRxYZrPMAzmq/noA95oIzWeCXN46L+9sdLsES42/1KQU0fgL02q5pYr0IZaA
hV3H34sxL+fFpwJLdi0TMqPI42njo4xBt6N0e8fX1KlA+lns08rcaj978Coz1gSa
Pd1NsuVeYTVcVjFUVLxgXSdWHG8TY9b9oJCWr56LIBD5uRgdOC0PShgsm0i71gxZ
2pjdqSY4PX4fehOEcjZc3qxBs+f5Ryt66qgUldZFypn8SP73+s6Bl35+jfwgP3FQ
dduoLg3bXHei39Bj4WsqbILwT7O7QxqozeRD/NdEj+C9ShOvBGXj0Xzu6QpD4Jjl
RZ0sKhRDHnDJYlSSsgbXnzgfe//OhUXWuIlXXTxfXx1lkWRCSLtxNqBhi/VhJdpa
wvKHplt0yTvwlTnajZAZc7hG+FaJzf65NLB7ZlWw6IMg+04ecDCiyR8SVrkjeWqh
ge2UbLqZg/b9WKLiM8ZJdqWsFaqn2CDQLUetoKcwLUucXCPyV8Oh4g6dIde6/rRh
gRDPXMOoqk0Bks8t2iDsbhjxrMPJYNWEZEcieAgdY5zb9LPDoy/dOz4OennLS2n7
utxzoL4zINofkce4+hPZB2dBS23vtvb7cu6UwP2MtP3kSjoJeV658gxQ2bCVjmsW
pGY416IljOWmb85lnHr56n/SGnR/iGA5Vxn4GB8PXOrp8gWMxEdHS79bmjyp32tN
zkSZnxtMsfHb1ML0jSwG1VATHpE2S0Wh+5B73AENcUgL3WIdP/zXUOwBYSmLrBR+
vSw80YOlJv1R4EoPECjZB7rfxpiUcGq6T4sIiX0+deaWwnBTjWeN/n3DCBbIigky
OkHiiqKgFk36ytGkW6XMc8W5kyq1KAOTyeMDc3eOFXboX8Ubqh7iSTJIP2JthQ9z
jGyeY3R308efENuFOgOSCXSC3/qYOWJa76HYzI61+GZfg69lKxweL0VX3SGN4erw
wD54JSbwZBJwH3FZtQNIAYNNerN/0qe2Mi8gQ7mVdS10FLs2A4MJSwStd9ifCbJh
OSDeBQa7byNB6wiKh5t8Pp21GQaj4j3qMKhoyOTiFSD9KoBwY1z/jSa2rKOHbKRI
ZChr86soDzzGImV6mceljrQp40N3RxyRR4ocQnqR+h38rSkf6iKS4BOqQXk/cMiT
ga/va+mbSBVJfK5SlnXtXSfUu4h43sSD7CzibUB1un8AGLarxHdk3CvPwxz7g5zd
M7bkKDgNTyrpTfoQrWEZTJyxqefFEusWe0eGBVsjv74AaDmlSI94Hi1+smP9P6Mr
E5XIlT6i7mSv8iHlQ65HoG8kNXDFI+Iuzu8v5GzDuzQliP0FBJiTqd2yb36uP2j2
LnHrsGLF5u/9xs0b7EVycuX9R4mTsYsn9+DQ9mVejauapO4pQAWmY6vjtPRXK+Pf
YgE6EALGMWy+jDl37yuaCxMCOFuL/I1ZRzTt0YDQQDZ0XpAZudRgdXKKJCf5pS2q
Kr+fT8OAQAYF2zowNEoabP/hS+NyRWojhbJaJZjUaPUYQl0oL5gAJuNK/P1MZ9Ve
nxCq5CYsjSNi2QURLKEmQwu/Et13PHRUBEDFLp1CpUT4BdbNXTqI2JVNIhfZz3li
ABWSV8ZSpdcjqma5Qw2GcAB6iNMqMussvD5mjfCIhRAlnsmHLUJWLF81wr3rFwB+
Sc4zvOeDt3eOw9/wWBzOd1zbRADD9WguRT9iOHMnMv+rt40uNQEQaOS75xUhcObw
PWzo/nTvxSQu1Ee8azQ9oZ72Om9VEAIHZ5STyG2SqOVd/9DDeRxtvSTb6jGCGFtY
NNNoOPMa/6maaBYP6ksYk4Tyz4au3nopoGcZOm2xpxIK0TlkWzPeD36T85C57H5Q
FHvNRn55ql/MYuQXc5NIBWeV14/VWExbVNMnHydWll7DNlojHr3vn9o3OJxOUKUz
TvMdGb6oocl6EhV3qrCihwin5kALZofEvVTBhUfMHc8DxcP+4txoAYu8DAGtu6G2
8D6olrmik0zmpd2EpYSRjXDMOxos9UAzw7hRKWg3eGrUpixYaWWJuE1+R2k5IK3/
WcHeHATjKiWC7mN2CMB7rwaJrL3H8GoWinEd9d7eSPBex8qEWLr67JxOpiN8CO52
jiZC3OVH8HwZJPX5vsixuoxGwX7GbJpBbNBuxIBGj/syWLOxcaBS2PJBpt65SqM6
zHAB5BMiE2g16KHG9+d6wLt2WjdxPVQMxf333BjXBGRCxvkfK2xVZD0lpjj7I2mA
/xTQkkb6FLMnpDiL7XQBz9GRRlZ0oz9hEUjcq5rTkLcltU85SvXwqy8fKxHHyZcH
T0dMt7Z0BIi10BKMjunYdH+DHeQs9IJRhD3wcZ7aURbUcsjeB/rM7onlltoprDkV
9fTBPnXzLMatq9gmmRSsouMFENUvDIEoBhCN7u23BoFFuvhhjRpy4Y4MPXr4j8TR
Zt/ADYQAAhmloQWXHbI4hBmyXxFKdB3jkd0VZUOvFxcTAOVlo6+oSQ9A/NScnYmW
p8dhDlcBOnF5kSwLA0ny5dqHzBBQLYhQBFi46e+zVLwEsWfcLwxWJsG7pb2efnzM
ZTYf85FjhV16NusmUIOZqBc/B3LHY06GiwCn2yrNFC5qc77qyMRfGTLUUpOjmaHf
a6WN2MP2qEnc5gBU6hOM7jnZ6vRy/sNcwe/A0XXJpRu0H3XmzqDfq3ihykBo+F0s
JEKNH/uXTKnF5+cRbaAttbhK9vHzM5jfO2Mo0JGAE408o7ucwWknmK67vh87F7Vn
NsRQsmgQmX+Mpm5UfeSF5xXA0YljLAurlU7Uzt3smknbFS8YuywTaIHwlUNngb8r
jcxeF1xFOMSbZ0NctT9CjsmNZ4Jy4ek81u0ZXLp5CdHTXQxGg4HmJtqIL0WuO01t
8N64Ak6dpoFCpRvDO39v7ClfGJeqkWdhFyR1mZEwzTlKKOjjILuDcO8R8QTyRNAh
eYiF1BA9m8jMUE/RaEQvkmhZk3inKcePLXaFe+PEyLDE0Y3aQjJ9OlA1WChQWLEM
caq/kvdP+AXKmhETUSmssoo8X9g1RzDwYU0Km8q/SQztrKDZDlFQV1FtGxSRz2Wz
xzChz1rPAcVqIsU5Tn5tCaVjNrs3+6X3Ues9o64bGYy4bUqovoWmmwMt84UXCYSo
Hwr1Uw2nlRzMdLCZZA2YXRyXe2IlvXMOsg33sNsWSdizzmL7vqzwC7XNZO3SEbG6
gZpWgbuFrzf7o7RsGTVNmFB0vLTnzf6LK22CezP8pLReY2tJBRIgHINze5EjpOJ6
JkQIpelq+6np8k5ltlrtbvUNru1M3vCtQbl+cJhm6Ps/Tuqkjgs3E5RAN59Nc0Pz
GWdSFMKRRucE7AJAmVF2XR3QWCNqv70Nsji96wMAVoR8M72Ki6afwbutLS39fqow
37wxiD1Giz5gCKbGcixtfdD+s8SXfSo813sYXL2UScey8Swhck6qHbHwx68b2g+H
JHorZAvxpxxAY99Ev47JzR7OK7t90Vz+ZzQqD45+eko2LRVPgr6KyH0niVpx8tMS
8moy7OJQmZmt1E5QMLx/02fMNO4m6JQYfPAOG8b9jbvJHiiW8Z4xQPBU7NG2CYSL
+HakoUvZwc9Ph8W5n7od0YilBdXY1qKKe2p1zl89YJsUiJ2MI9cmbrF4dzedFvJu
fyVUfeXr6YZmgeODBmg3l+12lIcbsy/dynymFHQiZ3IEwAAa2tEKz3r5OxsvezOK
7PD/MB+AkDCzcD59Xds1Z5xMfg8tGPYFzAFIj/J0AUnVLQrhL5GPPELemqR+63sf
LeV85VDa+Isoyl+d7xz2PSQD0c6loZFwkBMok/FQZmGu209IDQwzP934vs+RTiJh
c6I+R3yWxyJ82pVPf3d6tJHg3byDIweh2TSzkfjOytTjDVlmbuwLBvjTeAP0yz1o
X2s8/P7+j9RJXPvbhamvT2ykE1zXl4UsaUmEtZAMjT0OC+6dkY2/PL9fY6pYYAGQ
KVlWmbwPZVPHYppDglp8ZqsLSfQJu1swxS0DLe4Mqz8x5xWKGzzvJMrj1O7jLbHP
Lm4kkCXjGWvrBfrRxn7mJdjnbUoZ0LVes9Ypt0vOiRLQgelsypQz4MX9t/mujz4F
BhAECcGianjduIpoD6jqII3EYADI5YrkeHlTCaiWeaQBcPjN+BhCEES6d/xKyl6T
cfsUdakmbzlH+Y9HgLsRepymXzwfxHFRsGUt4bH8xzVqxaR1lT/7tNRf09rRwhdc
TsRU7xZCpoopeEZOWg6Y2S9dD+xX85Lhkth8zxQeShyJp9vKRB8FCt51pgN2DPOY
4IoKxh3zMCugUTXARKkk0dQbkgWEaHkpzZWVNv5dT9MayQ0Fdvb4ShPZlZpdCsKE
fYftlMH5IYKlm2VVxplpV1kGpwttuPvYYYrhJCx6DBA8DkmPAbr9ScPIauKsmdkK
JZur/mu/8YaqpeuKa53rhA/7EfaaJI4wioDHM/UTqCGlzMlzeOzuqzoTjURbzl5y
H3Hup0DakFOlisFWEMmxbdohe8vZS/RQ2mUTJcRdFVrRj5oOLtUomeUSosOahCh6
08uNFCkweQZBR94XlECont+H0FqEAfWE+nQ/X89zWhDPbEvzban5l8LaYCFvJTFS
/xEiHKYehP+FjcYo4RgQdJ1yehDbA4aTUSvmCkEQtDFsz6ho39b/PsRh6nUt+7BT
kq9nfz54Dnx1H9aFA3NbM7kFvJYQ3tkXB0CNfAquI0irLDToAjh511VG1lCsDHXl
sRUMtcWE2oqmunF20ou+vt4cOlxHoerg8gUDbXJit1VShKLIjDYKsjaxENUfJvqh
n4A4Z8mbM23wCqp4Jc0Xqzvlgddsa4LszOasUc+JUdx+9jOc0wwTI6X0s9GtsHA7
2YF34iUbusEMzPPGceomiS6S/mZocWQTZqEwVJp4BaoZiKqgs7haeXvyw4ZSi9Ps
a48UdgDhnv+F5ig0cIq0z2jLbxDBChKD+cHrhN5uneRaGh27c9Cy3tDl+FyXZwpX
WzluAZAAuTOei1pMKyzh3BC0v7DUXhJltT5RH8O8XsUG9JI8e+9pba/C+SEPb6VP
NAA65TWpnBkfXXgAxrj8mO9KtRMl2P4I0DxcS/BwYMCTLt2Qtk+S3+lxu1AZ7ciR
wo4gv9WIoervdrV7c7qeyhvCav0d1eNnv6xqYb4wG011GY6bBrt+DcYETzdo4Bcc
j34pyjVNRHv65IXfn4PXCQZPJNBEoAVkbPencw3fpGmmU7/oogWl6EYGeh8/2BLQ
CNEKWGrWOWEGSQAn/oD08RUnirYbpPlq1zynzm85xvxJclld/3stwyDhXn5mA6NA
uHWkQNG0zlpVY3lOyDXpm5BOw80B+7ro5RT0qsmjUzQkkRZWEkZhpaN3D/41i+jX
No8M7CABBmrqh7t7ydtZWESothtVQKwyImh+54vBH/pIc9hvQ0EjLkDNN0RkySIi
czjch2NriKnvo5YjekoJ5Ifp3+4V9UGZhNdu67j13e/sHuMmeTBNPpd/KQZIZAZm
Nls7pK5qIs5FNaBe//9faXakJlAHA3oGGNnlc9Xw28pufm6Vif1JLnQiz49d+AFp
zUbePSvEmcBxrw4+dCpmitliTcefQZUBS5bNkignHyxIhM0Up/kIPlcs/Su62bTU
GUB58kQlPbGkoeH1z5IkwXASI8lsC8VfDDgFPvVuEt0oPIvTe57asivJEA5+4PbI
MUjj5mgO3aPfQqSwyskBdNzc71NhwGPr0dfgVr0vZNNcac9p60U/HW/YDfyZNkFm
IN3uRWYFPpmExP7iLviY42RUw9HetrUAfuiwIQ8gCzOROh3ucnsu30WgQqUf875u
m+ZMGX9t1CnfILCZxYlf9ngluEw0JjZ/wlQoY0kjvNxNl21sPTk8Y9jJV1WXQQqz
Zj1AzPM71/NMYz9rp12JOqvxYvd3f66gm7ByRYKKNCnUcIfzMZSFumSVYneMfjPY
PGx2n41t0KcblNcqWnSoTbmug3P3FFyl5SzoVN8G4c8vy/pQuOwHQjHM+4kYw1rz
t4zFWNSOzjM5sEHJ0GwXcTeENRzdIMWakNvmnDGsIGv8GNxjHzHc5q4EpmMo30bg
BrCWjd74KFNBforTr8L77i+5I1jVlOgDjbM7Rr8crvjKKbUVd1P3HhCAbuK0fnGW
2zWeDKzCYjUnwdInu+KobVmAy/kxrnZn5hjE19sGdtKrExN1FGwElbGvcmFLtcTz
XhjBPHek+sEKi9JQHudw4HO9yN059aW8vHgUobgkwusK/KDM0Jw5Jwfn3JKIN8Cy
bZyYTUbKKKn3WZfTl4rcsyPvT2wChLgwU2w6WtwKF6gnANmx+zHE38gWTrN6vw8S
5IiEmYb8COg9PYipYABCwErRdL0C4JfnKa0WJGpB0TWzEoB9+ULdLoioCXnRjx1B
Mt/vkVa0l4oin1z7ndG1u9yxRCDeG6BvMDS17xYPCwc3tkseo4AT2XxjJJ8o7pLT
syZK9xslfR+0AsX5ZHvKxwdWIZCw7iftQNvz4DGkFmicPF/7mmDACtevWDo20Oux
tyIYzs58wIGJa3itFZ8iyPJO7HwUWWwVv09mwaIjqRLTjJjwxphH194Rk1AeCW94
HmSrB8ZD+gBhep2tEPD6XHw68Xyh0tnFPLRVgUBIyoZjJ76nMOKJ+zapg7P71lv3
5qnzIwdDDW8w7ZR7t1LQU2vCgOTZ4vbA7ZWpVTQ2+UHmd20Gy1OjdAI4Vvg5CUcd
mBEEGyO0hP6asscGrqxGrfcQx7ui8uDXXx1Gi1ENHZuRcpcYwzi4FAzESl+oypXb
sprAu1XjLCHc0E2fJEE70ccUUvgF1GDR1w7WoPU87b7GlwJlo9JP7rF6Vd3JhVWH
4GkA7gjFVWE9sDc6pTlEIzkoJT2JQzcYUXPmEoB+Hdxup8VeimoPXJ4HsD3rSRhh
UqNmaHZOMAJAPt3KO/pChRi1vfHUj9M0w5ZO1hevsIvEldzXTyZIXRFHMrYzDkAQ
msQwyl4zewfZzX+vEguCYMzApGG/LVenMLszOxrC745Sw+Y8Eai+0WVo0pX7vwoj
gZjfbFNfLW+dUH8wmphC6EeC7CN3hYNwaX0vDMdAq1Jy1RXLqed3MCVmvictYVIw
gwaQoU4EnXDwFWsbGWhEZOwBpOcv/nnT0f5C+WiyqAs8kTbniqakEWNnAmvJcIMj
0o/jBRnD/bMgnj5NSv4vPO/aU8VWaubyoa7bH8aNUOXp/I2nQ9oA2lNmbot1tk1R
Db8e7AsW5kq4dd4eleDGlKpkYBdCMfp8hfVxfVkK+ruGlao5nDmQqHEk3y+Ho5R8
nOKyd/WXGIQw8XPtojOCRc1NZr9Rh9+3EQk0+mNiVv29Mfpza/t4eNsjZT7zq37/
46mfClV4lKTW0opdqIXZIAPmCaboxDQ6kSBiHG07ixjCZwU93XqkLxfprMEzI5iC
k7oZjDhMm5SW5InGIh/E/7gTImR9IAlrdwnRiMnrROfvmyPAIgONS1/as+AlsKkn
iVq1C3RdBbwfzCmUQNNPEnx38rCLcXkGf4NQCQdvYqvZ1IYycpBlNYzrW0i2R2Lr
bavmqIO6C/mRzxVBnpULFmCjMbiIFRxdzMMQBSHDolBNGB01Ja0UxNVBeRxoxTx1
VcViQRmnEDEI5Fh4/zxgf5uUbgqr0V3F+gaUh+9Yo7mqbJf5Vugd+nNz3DqyVDIu
rOM38xoNmQ4TomujgbmO2hVV4vFxZb6AOMM0LX9i7nxzj8iALRwhspMzEm6Sjrdv
kq9gdpLKqd0QHJl/nIETxR85pyh1Po2KnQK27bAU0FimrtosKU/drKiDVtcAx3WI
CvKRflWtfGj7MkHYupEQA2VRyroIkkz4ag1c0IT67BFgjdr2Agvi6fU2cGpIPCB0
R2oocqjQvAV9GssE4CSutv/rfbEOmhmIcZvh3P/EQmvE6MVZTcnbPiFIE+NfbvaV
j4p7osM2TQBFsWREB2OTjXrkeGdAxllZxsUgrZppB/7PGB8SeEx6B0H2GAXW/6pe
GJ7dPTKYP7ff/r7EJ1+EFj+Tk/jMWuk+wC4InLTeUu5WdLetXJMSfpiy2JWwsva9
yujFt8oSoe3iNTnfxqLDisR2C7og70sZ/vF9cKUUanI1rxjI3jeaMfDwTP3k7J+a
tFnlmi3Apqt+RjrPxyM10v+dvuH16WeG13PqFFBmgEdMjx1yeA/rdugWeWVgWqoO
Qvv6DpRJxtpsKif3Rd+dXmNFYbhwmqdvFREvYuZ0+RNeb1b55Z5qI3U3wZgPglmf
o8+TSDR0Rh8n1Rrh4VfpARfayYbYHbDr+DOxuBNyv4kg4l/1A7PEghpRYJ99IYJg
k5M18huSRyOjLMoZDGq9YhxuiBXOZmkqeSiQtyRYQfh/8uNh9SQLrlqf1QOW0d2n
0ol8wqZePOeI8Dj+imaf0u6wowKIECWhAFVVYkVp+ZZMRG8VFrlbeOKAcJfuSWug
EgDvOJFbuYcLKnCGUO4iu1PbW/YeLyHK0rgtRn2icubrVTi625rU+NCPOmFc4/3R
/D/Zl6C0uZP08dKujB3LeC63+my4LceJU+xHBfLVk4k+EYZTaMu1XPmrDSn7PL13
5sazyalm4i1g92xEsg5jjeoxMq2lnRArqY100viVDsO4JNHXCNXhnDTHOG12Jh87
hV2ElrxrgF0ax0JMsx7c8U2vCzjuIyg/DIKq7qTPtO09WqSYFmpIsN3Ms/9GWUCJ
21ARwPQhivSf5PhMAllCRjDF2e8AxoGW9tXzL8BxmwHNTRG9M51cq6yvTFQi9RV7
Va/ihLwXdQLxVeYEpdFY/b3zg111XOeyNIq9KQzIxHwvcLewI5f9/FYyheWk+a1E
Qv7FYckCHpkV8HO89VgV4lTcIfw7C/fIYUOtfWJTHjDFc5DxNsT2bs5Fm/xyRUW9
TJ5BztKVT6zzjbL8qEJa3y/gzAA6G8uCJzBrh9LQNUop8K6/WZHMMfITXgJtUFxh
nUjRwe478qFAENnbgeEgII7ZNC/NB59K+ePnQVavDfcjHx4DUYZ5wgewdV+XnxEa
8kSIaPliVXWKh/hLWo3fVkslzcQSmV3nIfmGpiGaiLxw8+qAlUxY8ZUs1QxfZyh4
3bHqEVXpROCrySTlr/wXv9nJzyAB9u3Yk910vZmaTsgNYs+5fkdn/3E/ElVtQviL
5ZxhfJMgt4cCkQF4fK44CrTrZ1miBcLVCK3e6o0jXaCdP9x0c8jYR2mxC+cIZE6A
sj6EK4intTvVkBb0NrC/IedkBSAmnlboWT9yZmN4rpQVIUR5CJnZNtRlwXErzHbj
AaADtX8sOjZ6oMv9AuhyZGqYdWsJFf4hHFZYzwrx4EpEhAQz6aUhaNz5CG2rS55j
S/YviYoJ+xMX86s5yGHsTmKf165pIl0GHOpnAbmsIEQ+G83PLo+4/ZO96A+PtQ1j
IFu60ZKQj6kjowQTzdRllKSrodBtaN2zlpqiVn9ctpuL27+PvT53kOpfhyt6anpU
ML6dB7BGtk/PNTw+b8i52U7EJ5GxddKdoXcPNVjWAAqLs/3+xOs0Bgrm+nCeYOG7
gx1OjxBzgrNbVuVCChnhyEtl7Tu3+nH2JMLxMBXJpQWSM5d7Xsg3YwTSq0HM4sXe
BPlXddwC6RpzM/2FPZpP5tauWTYz1fZagn4mkh5Q4zm7XwckBYnvmhjUvMgve/P7
iGMYuEaWOTO7qWMvhWS5W38bz3RYyQnM2cXou9UYoNFFM/HdwQ8s3+3S/O1Nec4J
zK60sUBCfOLw7CjulS26ojN+C2lWAgVDaZl9+Uq8cbB4jnPicf9QdL1bq0cGjG3g
uvHOGO/s/h4j1GUkryMRpi8zUf9vI7QZwwn/jEEnuC4ghYNmRDQ028h0vRRUS5jZ
39fTLQ2c12bj/P5n59dGemBm7AelGQQnNp4xrZhO5CMnXS9dLW95x9qs8IjbXm04
9p+aOvN/dGuBco6Ryv2JCU6NPkdbJCBMEVeI5XROEGLUz6Yj9c27hKUaLGx1DtYB
KUofMhY7D2VD6MTwQt2d8cHJ/+ejX295WJncuo41TtcvddjxYmyGPPsmrztL3Ktd
cLbbK8lMa8IEAqisuYRGrDytyfzfvR73noZWSZKpv2C3AD1j1SDBwfBTIkqYHMmf
DGCl4oabLvy5vU1ilYdrqBqHMcISaQrPv+4R1mMojrHuqaYiQtHypqwK6aVAkceA
aYXlB/xbUB49N+QX6cyh5/5KBmadEPWnGeY19+Cz9xz7XLJGtNhXLuEYfUiI8d1i
Q0fKUJMEzWDwwbxasPgum6KOCWb89AnLuIYDrLXnYHN8XE5H430w9lQn3eUSq0BF
Zk+g6Wq44toAtIilGQhJdBA8UbhXC7WZqXW4VaCGLT3p3me+jd20u5SbbgwS14bW
45nuaoF+UifVWweeIEVVVhviekWynwYSdUFDe1OYwcNvQl0RSa18trX9hs1PuBUE
26A3veb3tjSTzMyCr5muuGYlOSu3QEFDS5W0cNjH/AUmpj8AzAzm56g7l1kM7/CY
Ylt0WogWd9JPQiUF7kFKl+R8sSa7s+VL9Qq5q1yBz1tspsTMt+dgSWJ9ETJCPA+v
CoIYPLStFcz3mH2gueWi5UodKGglavb4R4Yg02gmIud+GPdQD7sMiK0l8ufGRETS
H7C55k7JJMraHsmSfAgBj83BVZwUSUi8NSFJcbLeUUPHdZ+NVJraCun4BUeO4r6f
Z70/J3BSkjiyCBEKDzytenxuX9Lm2l1ErEqteo4zElraVPbLN2N2uDIqmy8fu48L
mgayZ25t5fbI/HCTlu/EsMUPW/D8XRaTeqv982rff8RCGxnNv8qH5kapBy39ctQr
vJ7Epug6WuzOodIGDn1/3ZlTy1e4NeNN1sVWYNWslfo1VALlwfx9XZvXM3LlDuo8
386S0MCKRAsFDHr/vaIFnXKIoGAKNbKW6t8Y8GsajdNRfk12D6EQNCOaESaHacuM
SJ0FN/gG7gBh9c6n+DvHEqnX63MWB01NNcWU0/9zIdYdjnAEv37w4BCkJqCDLD1P
x/Cr8jmI1VnIrZzjvMBh+LAXvSMN5zJ9RFzhIlWjG09jumvxqa5LxmObCjj0iwji
enqdXI4NzWMRGC5LjQRi03WRpT75d5coRdgN5/ZZv+atOaeeSH61lykSliH7d/db
WWHcUfqwoiXP6keMoUngmDb617wEWwZdWpSlECAU5HVmWhFcNPiF9T38opH/7Zi2
7Dk4TObHT22nzk0UfxKfP7BRcHBscaQv5EoN/uYFcSuJUgs5vXRyh2gWX/RpV89L
XQfubYxBHutXFRMHd6i2+tjfc4Gb1jjBQ8/O+E5O8SYrBvQSBCresxqsEtL6f2nm
UI7aBjRpAfdYO78xYlJgwIZHKL0wV7HdB3G/iczaDEr2LyGToUBTGdag8qzdVqEJ
anPxEAvKb1yGKWILWNCKnINXkR8tj5o0/vzSgzvsIfvpDuEKv07U+6YmnRtDsQ+O
48XVehOhM+TBUIXYbF0ezZyq39gcAxuTgCecvWVQ8a1NmOs1FaNR3AlWMSqULKwq
CFuXy3IRNUOEfrzeeHF4Mf9tVHOA1cNSZ6RZ/vB+JuoYOGqlTVOLV2FUGN3H8QlM
aGIUJ4gYFugMSJvPPkftqd6+clMYja7ZqdObdrHHh5iusS88Vd5ipIAlYnkpIJOo
ngug6m9wljg5uqwmHAqIBHyTYhvW8WFY0zmOgccFk5chRxAaGMlwV66VBfH7QBgh
Fzz+mBuOVWvjyyReVn5LzpDkKi4spQpa4esHs3K0lBI4t7HT/t70AY5QCK3avOuo
BV3m4mayxsESmohOn9MKl017qVl7ecH+S3c/b1gSK4Wrbk/iUX+N+DxJ7HU4MoHv
WaU0cLNjqexBgs6QtRqzHAt8m1eh0ImhbFkC3hEm95+srLqstnHwOsZ/hwTt+52C
5uTcVsAxlzlm0878SYVHZCQB1kA5iIpcetbaHmynivzWDPF3QnJswFSxYNO8siGw
UrtxyVZat6sQksFTigNg+KUagBjqQZv+9OVzePGAi5uWRL9sEnkOs2uh4Bv9vp0V
W/TPiPCHTYyd/MT+a20LpRG/Mr0mAMckdE//0Yjbxz19mdyOyzt8ookLd1NgzVI6
eh22ntvBL3ZyeE/vkeRhByIJvR7LipsIBgyop4Zpsfgrwzi/VBT5SahxMACcQQ4/
Vqi2Ypl8GbcFaxLdxzZPnt5azcVGMZT+wtKiZ46qRpEXS2T31jXN+9MPsLV+JluP
KIvcr3kDZ6TFMM2fPiteiKmg97VaS1EhX6QYjLHP6VyTAbuxSvboWK5mCBQ87aKN
g82VPwcJT3wwZPEWaQg91tUDvzX3Dyi3yDo7D+9WOKky6hg/1pU9J/0kqjjtY4KK
pd0nqIyzolFZBicUIiNENdQ9/ir5sjA+pA3di7PqutG2QS9FzXVHIpwcroFqJ5J0
hbYc/1JkIz4Nnf//0PSJHP0pRpmE5EK6MKX3M6tHUVZFX+8IoyByPm/kFqqyxdmz
zbC8MeD/0qGKIG+HIalA5nwae/wmCxLCDTJus7kigaCXFwx7Y/qn8D32nAdaWKZZ
BKqwupmFEPEfBzACkH0G6OnniyU8j6IF/im0JuUBvP0hTBTtrlpg1FXw41facSEf
uTvQyUvuHtzxY99GC3RuvJscp+ar5TZcR9li85BK9vq/8+/NNTmFx07ZL+STXjqf
PoALUbbwE1I4x5cFpFjcHegOmhkc5e9Hw+BoNYxjGXdb8MVsYdeFati0/0uYeG/0
P/11LmQCM0OqHL6j6DzXnZS/BX1IhJJmja3a8cZB/LnDvj36/84yNLQo71hIP+2f
56k9w/RFpDW94/TeigwVWXZXIAUh9XwMGjzmQzRb41+eAZ0NjwktrBAx39GCKeP1
aL1v5maAWjhcKmKQRVckveVRKkMuEn1k6zzFiduMzb5KQux46TwgEdX5DsfiCcmQ
5YbP8jrNCupoYvrqyoL3WP1PACr+Dd1KcnKA6Bd55lwHCNx1AKhzqX+MZtfCoF3O
m8apUKWGpfTcbHoSBq2g3hP1cDka5UJ5tRMvSPRRlZJD5TIIoDEmgzbr8o4tXFSo
oGS5bdgnSLqhHsEapjFgxxwIhLgVGI6iXYMPGY/ttXHgmfn4rS4jtUmuOMXUAKnA
FkMNlUtV3vcuM7UASLFGTU97VFeHIjv4sB+xa0nSbhnlwgZztiJTxbvsVyfFhU1r
qX3fitAlATIcLXZgbzBSlV4drB9Jtf+d5FPJtTVTWV/UrUMqBFLBbN1HqD28msbe
dIVuAeLQvo/9LKEYKq6OqxGbXFExatBK+ELKtB0P6EL/CSSsSY9tnQgyHvTkI66s
x7UbTzy5omlMmhKfWwiIewqq+nNvU/eT1NNsQrzUziZAKpBepbv+jiLvnGzEqOPb
+9rWEuSRBICF6N93V4n7eO9eDVgg2VcAXiKQF2NdWmnN8psa5ieOmj6RhaRmYkGt
v4ri5csAtW3iUFf/w/GNluYzXhRkQlcy+BgTcB1fi0cjSUZO57EHOE7+9NZslYd+
Qnqa+YZS0VsX4nG/RGWpJWQ0JYaKnVozUC3z0ve7TO5bJ29qndeUlxjy/VZDPObS
ErD/m7HlWznXEoWF422A110ffPHAdrHCV84KbYTIpaNWnMsFA8iVJYsYt6jlwT8C
/EPNEdBgFCpQl4hNEOhj9tydHkQdfS8ZzMJCaqCLQ8qw8zhT7Wy6Mtmj3ffL2PR4
d7AGhxo3vM0Q114Kj0zgQvBAfqHaTV1nKVcpjnijphewuoLN2RHlyTNAdma/q7jl
QyJ+5bEOmDk1ofVjrtmOFqeog61O6qbOGH5t23sHGldvEcKXY3Ju6RTnVcqLWzGJ
SHAUb0yZTPTsrvWedcsDzOaMC0qysqLNNC/MYRcd4/296TFa5iiWykmzJqs6WEpC
g6+ovUBm/VtxAZLdh3LDFsllETSyU/SODKN8BH4c6KurqDFKGt5wEtYJZakG6NUn
d75YBLYVTrh6nPkyxVKW2jri0XKVbV8jW3DvfGEi+BKZKRDl3RNDijc13ZZUpBoo
6T/GsOUoMePtswrTt2xh0cBGb0CjmaQ4o9LqzwcxLEPX8SoxfbHZ34C3o+KU3hAe
GrMZB2yi//A2HnX8VMZJl3ztaYMNPwI4Errie6GuUdWMjFKIgxOc68FAE3lhwjC8
uNtXCNleEmEXcCoxoFidhlBTxHxBh6HQfl8fz8nZ0gqRaq4mIRUMwg5q9BHopYD3
UbRgf4xFvKAiY4lcpTTMltQTqkph/622HF7Moq13YlMEHOu/FnA+YHI379gZJkSB
h5ynbukmzVuQWNrHXthevKaBx+Wf2tiDPUivaRDy5CkOtmE8kqSOgwM+vQzTHGrl
69vsEWuwJynIr0AvsNdMxyr38LVoglR0l4jipoK5HNO/YYw7igNkVdth0nQgqeX5
AI8KZtkTxd8Mzhkn1Pt4/Bpgu//D9/jK1l7K+hfE+gGy0c7RAQ8HDHwJjWCwV+tp
ZMhtkSDaW+LG6qdCUIhuhwDpBFz74vvWPUXn/dYq/bzwhS1F7TwQB1fpHMZETM79
yXjI4BQAjXIJvw3634eB1R/jyNvzYW4JpprYhQh/3lCucQDCNK6Ua3A38Q6Y9a5h
cFWOOPhr64LGfWv0yvqZCOeYgj3NF1FJnDKZpffXNFmCkSuMm9IIIYoHIqnrn8sd
2iaK4hWxaMmihQtNCyV8fjjn1rQWQiiei1cDpKf8QmM/b/JWK3/4QIbcRTFd/7Jk
Xa82mSJjnPkTMkq/9jsO9orPPXNcqZVoElKIM8aUWPyA5gOq8HjuNOZDbCO5nqO5
fMqSb3BlS7biupyNKgiQsXIRnnr5lbBMNPTzfwm+KFYhEal9j7o4DMsKzafroQy+
bp3cjQc/uEvMOV17jOFvsiHkU7gYiI4gCUqwiAf0MCyshEfCXL7RQPlVmoSDeHUt
mha2bQGJFxH3DqO196XBUmUe/H2rKmwOj5yNTsjMafObYgGwT1WEZGNRqoK+FPWa
MMoPgvEpd9HoR4Hlt6vF9rSdxPzKAYyQaSc5pLD5Qz9uldynsCU/hDTd/QqPud2Y
Ril/so8x7/TyqNPLIO1T6Ov7BNnOnnxdFpmf6hZkZkDgF6CCZvJSb3JKKmx2P36R
OadtLESc/ML7BVEWzpKKoehzFxg+eUxJTlmwiXmznEAapnAlRNHMzkeTKFjGlNYe
v69cbUHYTccNV5M/UU1WzB5WuS6CMqqB1f+yjO+AhdFJRXtUHBJDwoCdhIkHMkPe
jZQWnIG1Dt8VPElr7H5RMnW4diUJHEq+Ahohy2+NfUa5PXIf45wmN4jnoX+/xjk9
UnU5J21z0XbxQsRn2eG9orlSwKDkQ8o+0q8dvVR704IkDrG1FoxsynR0vUtWGKqH
s54w+hfQUt+gOMewklF/DDpux7FAf7znbQVgAoXU6hLw9Xx6hmyc3mX9UQkSM7bv
MtdC8Hq43IfTVelXt3xVLCUO5UIzOMJgaS+BvhWI4+NYzT6isixbnWq3B8uDauD+
V8xaZsjP8JDMN1lWd15tTY6p50Gy+iWEuNtSlqm2MUbg/Fr+yXEbOIm+Z4Zk2nUG
DjtX5c+u4jpuvmNF0bF6yN+1UrNqIXBscm7fnDzuxN/ccIQHKxXgmGwZoeoBIXen
fjT07H5qid+dYZI0d5x3e/OjOQAXB+uDxXwND8SQgsmn9LrIBZ8tpogREePpg5hL
cjElQQablbETHhICUxYsbU4ERW5S854EqsEzMe5ac6F+Mfa7jyWQYjFxN5fQenEb
EG1Tgam6pViBRQZSXF8Wc/1npqObW0KvUuFEyyz/aKfd9/eV12IPQr/rRe12ZpIo
NHgyeQLJ98cE/A3gf/KrIUw7NANy+jmbiRJXvdqIpHfCmgLwL4AmrJuWsgG4Xbi9
y/JRE/xRThwrtWlM4A/5byCfAtv0mltoqZuIow4aavRFEC+tm6caV/lZqPshphqj
4UbH4gzvY+UFu2uK/2rVb/AoxygO3XH0lLLjAg9xL3DDYzEbMzkqhPwwAOX4PZPl
JzYqYdNtbxpQdfv9c4DQGGtGWl+eR3BZK3821Z0budzlkw4vXjeBgLKM1jgHC6cG
DBF6ds4l5mavvIVOCevel3jDcbLv1fPdZlN7bxagUd/LN0+f+0XZ8uTl+p56zRxa
FwXMOyJN0IcCAbB7iDcfwQDudxW/4rPkNCU5vYYXOxVVr22eoMMHcBTflc0WPPTM
xdayl1KHLyIoWvsuR5QJg31IJb4P1s2xkwf5+5EW4bCkD5rsiwYPCkek90zCdtYR
//QeWzKGTaVXOLERCuvW3KspzEKbLIkJvuQsW8b59zmTNJJ09wMZWwdU9o4SeIxW
Ajy4m+bmELV045Xk8f7wV2wU+wsgev+UWE9chohzzJgVaQzL+d3UZblLXuxBk1b8
sditPgnCE8ftPBB/++KDQIdqno0nC/8Z+U+07ElSjYBcVuNpxXUpeINMfrfXgorP
u4bflIoBFR5y0594HJGCa1dlU7czOlv+/ymIZjgELIZ4BSSEaEGXk5grThUMuG5d
MhvUN/9SqEKIq1DNyCXF+yrCIJN9DqclEC8asxHsHSKyha0xCnbexpqrH4DKPl14
O+N9mGO2zV6FnXlcXad1FAH8bAoMk/e24Y4xixZsHO13RfyP3EgvSxlkjwa8zyQw
AVs+zLVdnqSTzSawzcGIDuAa799LwN0CCX1b5jROqlFZEnYRwQR85m3ynLjMyVFJ
K+WQHhdDI5wrF4L0Dve20IgmnqYsU6dLWtXXPqsEsPwLTVun51amOqZk2sNgIq6s
Aj49Oy08takqm6B+7/s4Ii64fTdFIMl2L3nICZdXZyl1baDXVxxkH3sA4oX6sqky
tAYxn2cXjSoQHn4fKFISRy24T4Yr/8EfBawWhYah/dSIc41pUYtTbksIYwJyg65/
xZnd5Z/SiOVzTXio8r20gmBI/uOiSzTK4QgtohFkhhikIm7fgx4x7LpaYlmQj+2O
kcRchIBYiSf8Q66V5REPk0MortOLTuUDlf6r3+CjnX/5arQXQIEABC77bbxJz+nV
O/DRWlEriiSmt5V7OnhWj1HxoxBHmw52VQ7PkGGj1FbN576KPbChLV8U6qEO7pNW
X9qW5FzUOSPr4x99h71nTckooRgzdYrQSzzqVhx94/793faodk2UhJ+QRfczL8ns
UyeOG/0YSrQB9BbHG5p5ZaXCqpastwEwZ6Xkb1payFZrFUhQ+Bgrh/Tikm/clYMi
J8S25kmWUyKiGmVqKwtWmAzV9BiQ51wuY79Y7jlXow4HHPAHTn1nzOYrrfOnYJLK
P8cO7w8HgudfvBf/DAJzBQgaFQr8l3jIdBFT76lh9rdsjyGTxpWRaM43RIWA1VBC
vkrL48RM/C8UtnkLJkbT+lAKOr9nFdbx2VNNYX1jApLc+TBJMH6mlm//IXahkVHB
E6xMsuR43aXl8InkyV6hg2ZvoeKgaDCLR7KRhQyeINWXWu+ALdA/ZZ1csU1o15tm
MWLAPTwKF6Ay8CYKE2VsSJTn2JXN0UD5Kjwm89Y9lojjNg8ZDdO9jIgMaE7mxYOb
nvQ41+rhxoVA+AlpbI3fUS8IjNB/0Khhxh7e96HB6JopDB94FxsKv0788g8L32S7
WtahJQ7dkydyPoH2jXaS4qTOqAvthHYPjx67aMaP318EsxuyyFFclEiPV1gxr+qi
i/yGGLRreCYgD4UIRoPsMcbRiNPsj2MBmzv+3VPjewVDTz0FwE4MfVPzKRmlS0cb
qNRmNu7u/cqji426O+Cztx6WC8qHMoVc1S4/6/H4Lrq5zgbs3xo8zMvBUp1SCG86
XORyYKPJLnzSRKo9khKTttHvaO+Mf2eNxXQgriPK0KP+74MCjFt7eko/3dTqv6y0
vu3blyBsWM3M0UDfqcN/FT6S9aynYibhhKHM9P49pfDhNlnW10a+tf26oh1Fk6na
Wdf0Oo1uNEa+vdHYT7OXeYg9XvN0iTJSonyE3sNpLtNVI3sNgxq5BQ4x1RWS3qxC
ert1gH+2hqKQFxUKY6jTs2B0v4zaQOlnkVNzb1eEjijAXqFxSQtAF7aDrtAPtY7C
kWJVG8km9eAiEANLOiF9kWywxZUXJXUjMv5sU1MvoJ3skGSwi7cPWgpPvLh2a95V
iRDiwj7ih4f+QkkGkohQP+E7Zezd8ggM4hhyWpxXkbKIO5I8WHqgjib5bhJ467h/
o1pXzDfjikcjoey0BBQh/xH0k67pvXdGId5G9hKVGI5hgO9x+Lm1XqLP9dEtM9H3
ephMsv5nyIGlhZLHFjfCLtCjspQFMG8L1+apOd0VezqlzuiAjfcRdN11MZ0Kmayl
VFddDEamqpbagvDxH+Ssr1wIT7V9SvNakYU812I5HzneiCaO7Ytv8UbS2UOaEgcc
MdqHNaIugXf1k0apqnsTn+czDL8ySDApTDUkdaMDkGrrAs1wcYJxWBmcAZYlZzqK
ad6sj29hPb+2wm/22aB8PkYQlD23DkvIXr80PSbIYatWiXu5tqYEMggWO1dtRlOA
9g0qOkPrliADMfxAFz/vhgPXdgR3lNCGoE8Rfu+qUFEGblMxQlFs/GKbASteWD2U
wlVCm2iTJr9+5TbwWz7k/7XMRvzaqWYXz8y4++CUUQdnSkggiscU7bv9sRAyRCUX
0gIZgsz+yqjuRu3yuK6DOo+XQnNkQqMhVUNe9S86AlvHhgzN9TkzgRTbwxtsGf3j
/5eGtqb8tA3VaQfpAgDrDwkiNUBeMFbCt0A6xCoH+H2bLfSJWUWfek03x0zyfFNr
HP7PdYfvpuYrE5H73aosX07fks3Y8S0jlL//jTjuTld3QXAeYzx5MR8ZmH7dWJha
rp0XB8fGU+PnJ+wlet74Rs1MWqRXm8hVy6tiUCKXIriFJrM+lsjnjyQdj14chyX4
IxXUwbV7JDPQ7F0Q1dWke+DU0VMP63qBnLDw2Q6RbdBV6Q7/sO2W2KVxUynIkBBE
Rs1wstbYI9OlZ6NAOrv9tJtpi9S6Sl8nNnif2TnkE4GeWHocp+OfFwRsf4rEuWFa
scTELbfqubhqfQ3eyIBt0Y6UQJM+/lPtC5WJ4D/5E5gLXOu35zFrJDM74dsWjFe+
zNTrU/ibW1oZCAq4zjql3rXss2ZyWAjoUmBO+cjvkBJofOFCA0mpn8490tv7hkqO
IgjCdHraVoglqxFjNiM5xxnYJidTELf2Bds9ubTd+zNK1hGIxDbQjD4/a6C2pYAz
8OvGcZqIPnwK38w/UPwyu09zObm+IpAmr9a5QVoMikBdlXn+TAGVkli/PwJqQnEj
/eZl9q1hKM/Th/KjZU7kRky0HIhXWFVXcQ8Z1Rp5HSO9bXmBD+KK/tIqqLBE5SiC
WVN+US6aT3+GWiYatOCeVUI6NTb86JLtQ/S1liGa9CaBTM3z0WOURGRATpuPU5Po
yV/09QOeRQI+hVgGV0Gx3EeLF2lUQvBPot1aGyVRow8yUn6Bf8LQndiGbkPXdt4H
hAbMIeIN9wPOYSmaGAM+9s5KX0A7NiRHpRDSfJJDl3tmDK1syn94TDJIdxxNvw8E
lnx1qcfiTHxp/jdAUYN86io7iQjS1rDRICf1sSQhP7O7MFFVDZLDhbkIPy/kCoPB
CRTQX08oITLKYV+IEffDlUyOnVwKcoIxxj8LKqMOtcrh8bv9+l6rU1gebyj6SfwB
2O9hrmB7gUzYMbtWCbTQ1XT97+Oc3LudX0uboD91eHnRNrn2j6h6Px/idvShd8hH
z1VGs218512FonLGsVeNZhPSEWMbKvljTmnf22aC8DpB/JqQef222o8ZA1mIiwPF
9u9Q72nFbV7P7ZrqbWOOJBkXI4ng4jJ+shMzAfoTx5RTnlygVEqtIeSQjIgyBBGt
r9tuRjZDtjYnP3vcQ6cMz3h2HPCCjpzRk8DqXj9QZILWYBK2CKgAVZUyCnspwsLQ
nEH3p+JsV+lHz9u4xSZlF56JQQaKe8fL8/Q7OsVq2iw5/NeynjDyyPC8sZA++sUf
YdRCKe56UzJuFeEC3nIin0GD3gqU0J9E+I39cL8F0Ztjgbt1lgRewoTViS75hj6B
lt52cE7Kc8pFnKHYcHj/tL1JB8JN1fta0tWwZ8rtOK8daJgNMhbGo2+EtGQnFZSc
wt09xHtvzF1ktMzKr78mpIOiCoD3j8FZM38lWyZrBLldDCSjA8PciJYLEMP4773P
wU88O/qI+VU1mzqjw/crQrwQCKV6EEtEUCkJpJc6hAY9mDVbGbufkCfouOLYQVib
e67XWMH3kFDfEl7DoDchRrLCrR8u3hUndO27GAV6h2Msbc9rqM4BdCCF8RIGbcyq
0VA3M0a1kcKZubDooeArlfB5f2f+nArLPmDhi/TnEy2RrZIXRtcImCL35ejk8BCz
5S8h+DdbMuokJkzG9Iq0F0UXdN2s0DPtkLmQKQgwOT2K3mc9Y3QqLKVj1oBfuH+R
hWnh8CUHP5tuemvFuTC9ciYDVbstINWb5V7+3nAO+Q2y4AIhExmpiBaG3MzfgGGC
XHzYNb/GeesYP1IHvbuJji/HH5iUp/baqSyG7BJk8Cxxl5hoxrep373RSQbBxyPs
EzllBj39Kl/stUdUmyjxy2GOwQwsOQVUcB/Qkc175rwgCPMEc4qvQKtCFlc0hf+m
ARBfuAeJdMC4bEWiB7xLqzXbO1DGrwEvZKnEgMyuqJTsm7qig90gx3njVnTk6ffo
ypyirIwUmT1Qk7qaqaV4mvm+KXa9C/5EbAbzcqWKp4k/Wa6RqG3FlVSjGEFqaoR/
OH7WhRNOpJAH2XJ6yjHj/b/TE1zK5vta0AT1OS/v1JfsW7ODSgtUxy2HdD68CcoE
t/ZtIq3cUVi3TXT2CSrqj3gktfw0Y+XYh05IHtzFWVwRNAR0ZBxXTyWkNsfLRJVk
arqzW6Rc4beQU1192B4VzktTV/zrM5FjtuV147+qe2LCthrlLwEsrDBkSQcuRUUr
r0iKgZc0zSUER5eA35pxbYKa1vJuTrd32BiuWQBTM/Lwk2PpYHx5Cv00hpNHTNrC
HN3nVMyVoIVUvDWD3fLRJMwbcCswPLppnW14okumkSajVM+UZ41FzNNJDhJfdhvs
bnyFhsjqITv1GQEJySz5H4fZtbMpt8LvEZQPmuMrLD3ZLP45sTA9bW0aNrrzYQ0u
hPyhdLcYiECulgJnbE3vNb9E7giZffqTNYSrIFlRkweXmUvNkjNDLn+DmD3TbItD
A2AQdVVmiW1La/+rbXuxF9A6rg3VvmsojEtm2aQyIwhe/uvePxLcJh6ES08V1pru
Q9yt7eubB6r4NEoi+i82Ss5UgJ82/ETHtJNA8as08cTWtWCCPw9U+kN2s6ucWqKX
ptoiYDyME2wBZKm0piXvCPGgl7awsCI5oC2JssqAz+iapaNijxvTrYkZeGI9JhEh
y6EgqpIZSmQOWTU5M72uXAkiTExeuptRebhZRjXEXnaiUMnNn7d6Y4MmNy6RH1/x
NHQfdoyRPpGZOwwgLL9IlPnN2q6Z98E+0n+L2CXvWD8P/2qb2FdM62qGaH6b/4Xq
AWxfAuljSRUX0z1Wdaipo5S0WcCWQG4FfCdmnB6BPOVpdln9JhWrsKbdNhH9kxup
QHDetjT7/eHdM4v2r7Lc4mfdEQZz0iQR1x9fPzaoVfVYD+Q/Umb54AGffoJbYF4J
yO1VD5GHk3j2xhHEdUOzvvQkOYv1q0LlM1QxcbOSmPWpW842S+546ogaT/2R+xp2
UrmaYQevN95eUra555ZIeOR19AOUZLLXgqWM+grR5Cm6v7ymGg1txAMKTa8OlgFL
VV2B8ITUG0k8Yaw/YrbkZuxp5LbEx8hzFrEvjc8YB9Zj49lrZjdODOYAafzrMaRb
AL5RoG1baUZV6xUpvlMO0dvexflVdWYPh4wtRQ4lheMiBrpxZw+gRYdv4KzXanDQ
RrzExCqdrDpH2r5pq0Yip0NsvwAI1K9oZ1pY7T6VmkHj9v1TpRHvtieKxdG8vRWp
jRXXlv6pocOu3qnpMkz45TOBeZcpiDrsukNJE+7O/81kOXhYjMJzZiXW3wb4IuNO
YoN6/kGrs1Q2aikkafIizQ4EYJKxJPcX8bYrV6JViLhL1ut8eCSUvdX5gR8HssWB
TXrIVEfqLQkpEPhu9/JpjbXeGwIahiRFn3XcutxfIktJlo+SAdFiijM84VLkRFns
3ciYMbn3sPK0zAWkmDWbqMgOhlq+kyuWLgA0STIotFKARXNE4UFDB0xN3y+/Map+
kOCzfgZy7CmZm4DYno6757p6KQN3lPY/pAmdHiwDhjc+Ybf+Mi74I0za9HaBwDYI
5tOUEr7h1suFb475v7u9towpnTPmUPQAbaZ5VeHx+72sUCgD0NEeFdtpcznYxBTe
+KmwxtJCYTy4NE5l72eCsxNUgCpGsMG1mobLSnNjcqm36OK+AB+tAdLGIZD1d396
V3bet9il4JCXO/0b7/3rcmmx8IH4ZlduJ6IapspwwUBBWXpALfnF0bRcDdcpZbQI
JnC5j1OIq5f953bobcCCOlKg1bbW0XW1R5CxW7E8UAKVHnvkAzBmFqFC6+fZ+r/x
Wr/vEL8TmtWCnc4+sW0I0s3C+fDUqiaDAMSVWvf2IQ/0w7sqVeu9XWpM6Clzjzc+
puSXzCS+Zo+q+2MdoIHJYekOu++jRbEp/Oik+v/wHjeqDDnTdD6PQ1r/MqENwavT
zB7k4/5cCz5Ur3Ah3e/JDmScIO2j9laWwmCrWlcEQeKoQUdhkJI47wwOqhTz+bdt
HehwBHG8A0JuoxFWcqw96cFxRTOFlo4W94DuDBSPZa00A46oZx67HK0Ywb2uNVjl
76BI9dYz3NX/av6h/rTyBZZo0l0ransCmqlJ2QhKmCiNLG4mMZTTd9SLBQQkVduJ
nxlEPUQ+s45Ihs+j072m2UCig2GdDRY3YoScDBw0mCNBxyNEyzD9CepVQOTDC/DX
1N6Wl4r99XnTjjr+sRKB9b7spnahSzvQnioekduKl5GJhFCjWXS5H7rITMaIGbCk
f3kHoSvgoxPYZ8AUCNE1bc7CpjU2NGuaVPD+gsbndKq+XyotpNEVGI762rkCe8bn
GZ8gRIDU57PJjGSr1POqxGBKsvsGNp4I971C5IDybU619xvQMO3NssGX4dCfL757
5pXWDWhdy5zwPRq3TYJCvwiH4ScoiGcm2mUXCt8H9ZEZHWq8visjkhUstZnGzR1v
5GDmVLHVVndBze+/x52BzIVd8jBDy/eA8t1vAhf63XrMTl8js7V+zOJbsApCxXk4
rh42zNuQgfQ4yh3QApiPX087WA3hYN2JYGDWnGGMQKjcv014hgw8yIk4nMYeqDn6
nh7gzOGhfslw6esARlUR/OD/fmNVFwHBtZlaKnb29JIcNjCnW8qbFuqp6DLxwTQu
jPez/h1//T+slo4WDF/GAALU77RPO7l8JELSn6wpb57TwwIaC2eodhW1CBm0aqlj
HdaXXT5BhHT0V8pKYfEho2f13BHVxSrrke5boWxdVs1vzu5QhMjJOv4hEKF0Lyg5
6hXJ3t3psw1Y0zKz9kc6uNO7+FxA9bJ5symeD9qnlrhC4oIgovPGZTmnSaaNmPbQ
sKH+5pNEN0bs0dM3TLNl4jKN1IwMsxYbMGxYYoWcFyxM7cYMq2VE7NOjc5Ho8qED
dumoITeO9gaQgrKOWr2JvactfusoHeCHx7xUvvZoKWmAT6s153ouSRkF2T3B2Gew
NFc4326ZfaD8BCwuR1AkGF2cssZ2boH+hEr1huN3pWfV4DnxtqTDSDdbGPJLu6pf
fGHoPLVfic2hHKg9z1UjaRJT4s4bsY2i6rxtga63VsgaPVwA1u7m+YOSi4PaWdxF
AQwijzxCCObeq+2RsJVWENUeRLaK69uShgM1N8VisXEgdffBlbr07rVsr3wg0pcG
QAREZF9/1DJ2IzZWlfZRMweuiLvrWQIkl0yg1JQ+NQpL4HcH1ZgNu8IVuJzJ+00b
VmKELydRRggQh7XYRMj+bO36UsyfyaT+pzKY1I4Dv21nw+vHDTRAdpUzyyjq33Uo
JOrbLCIu8O+ehZ6eFMzI1mT4X7omWxLWBV82rUTdf+VPPraQmkbdehLh6TP3yGmH
MJqG7IMAgR/kVcmVtGQ3TAFwiek9aLIk4PqxOovoQrGFbJiCzmyuYCWX/uEgmnR7
B1kaW0J0Kc2l4O/FK8O7Qzv5FFi/mhZUUNAfXHNEOaSUVJxqPZ63ovHwdDihR8z3
kMd93Q/RgWABpz6u9RHegRBHIhafR9wsnpBTHKTttBVKJ7hUa5liNuQ/V3qR1cGV
03AEr3/cbAZVpSDWOa0gabV8bZZyP7n6OFSIuzfcCGfH3j/o8BWf0X5zcmPy2443
QhsQlRvpOADL8hNjopeQJQEExwoZk3tp/TIYJm6UdU1Dp2BmvPpOWa9/aEHphT+m
eWWTpbY3Qe+IZCOy4tRx2hItALdBjI3h5WL2F5MB0tSaP+ngs1Vo+mn8XDKKtR+3
wJY6pOPWY8pWXvKrq5+W1IU7qMQg6PzQwRBsi4JURGIYSU/OenmHHBz9K5aemPG9
2uHhzKNdUu4mqwrIPh3nf6uJiFSsNB9ZuXoeBkC+ZFnOXN4Ps48wPeQ9Pg3UucFx
8WOaW986zaU4CwDetXbOCh3Ml48DItyk3EJ2DJS38JdmMinBi4T952sm3F9E2nEW
KS9wJO2S6rxhjRnOIodGJMQ6MAEwpYcsEfV/Br4A08yoIjRh2rTQjrfE88WH1wk+
ZzXIHbcg53oCW1SoTUdV+mE/9eshL0wGcowX2FNnODgY64GB/b/ulVGkMk60GlqU
8KOKtTKQ0Sn5fnU1hahbn+iF0c7YH+PrapQ0fZf2eksznTcI3gkgGLRaUZpgEMdk
LEQRM6S0+64DkMs8QySXYgbHqVoW4iMGjHG7BfWLcP5fz+i2vo7k75VTTN+D3+kV
f1F5eeCuBH8SH1JOF5xlt8qe1vTHwq8HAZHRCC6tV2HSAQFmzM+4kXgQSA/vLixc
rjg1WQHJQBN1in+Jci1m6x9A34k2EbLn99P0w7mL+Z7r+uHvsCC3VBL+XxchoMCX
VCGSo5/ONyktJttj+ovuYsA77F9/gGQk+BLtQiQMDgivFhlpLA7mwVCp2gHTGSkE
mDbHi8rGUWBpkp0z03ZMhmD1NcL8LXC710d6Q87vNnjUal8wS9DYqaEVcSRk62wu
gCUPAZtouCZn7f4FHuxSUI5CbOaAG+bjhd4Z6uZA1DsnYsB2fhoiKPQ8cGY/buVw
/5+39iLy4Ef2oFNRBtMkvrmyLQoVP4EiVCdOtNwLGixOvqfavvTd+FAF7nEcKW4s
C2+FBKAcLfZ6QKoqpPnjBfp9OWcQaVhQgnnBhh3TxEk7Erk0S4dCJ3tKJSj55RVU
ijljJEcyAHI15hK1bDdBL+dO70+Xw1rB3a9+fWXlvPALFau+6qzBzoSUPbVhCUvu
76tBBHt6MLrfG7w2NXjzJUIGuClJzfqedHWzRMHW+9dXqeWoag0h/K2LdjMXlv3q
Bw6nWijvB06zIcYNQdK+tN0aE1hWaiz9OWOxXYFodVBVAvW8nsH1LX2+uZjXfB5c
mTUSxAKxPOjQp1TFEuYjZC8HEa/naCP4zaD8bCX4FDuZTHmRMoykyWijiU2zIhKl
U6qjO0pvyqMm97YL0BX+u1cZqqIVIv3oTren8GLAcYgZRxP3/IGOOHt1IJd/lcp/
02OiSrRPoqYK6gPZhTr1Nns1XYMwSkpdPh/j7l8/2Df2xqHCUBtI0UJpqC2cjiLJ
eghVJzYc/hQ/XIuAw/txrlBqFiYbEnJSU3hlRsWSyYtHX1e3ucKG/GK+jGbbQIw2
1FPtbKpVSm6FoEp8b4GQOTEPez6UG6sPPqIHyOOzcmVx5o7QcncIaFz7IT0a5WQY
F0Cl/6cUWQZwo87fNd2bSXRa+hds74e87zvN/ymCDnqzGBrAivVEBZ0N1D3fLRXu
l7EgiOHQAVdYJjKyhRuINPcGZeSdqZm1gJZkZ1xbAxfYsKqgQxpQDUuCxn7O+I6D
MN1bGHGZX2xjYeWSKjg9NzHOMcDCiCpDh6J2Bu2S3TXw1mYxQpgnl6ZpEi4dgOry
9MLkighOFCflYJxh1BpymsdCS9ebzfa7D1IoY9f0YC9HJutUb5CY3ultvUt0+wZz
TNARJGTOac3x0HZJu6OzMWK5dEdZ8b1UvF9O2z8tAcioKytxajkt9IKKsIH//5qn
G78bDLPOVmWVRiWG/iVvT/j3Xv8NcQcREDL3HupiTDoTTE8l1DVqkhJI14Wyg9Q2
W0EXPemtLeh2JjpfPXOiM5ufOPWQPi71F+GpTjoPIHoUPYB30rjGwDHJ7BoO9wtR
N1Vqb1FvCazjHJcwVB3i3n3vBun/f5jbJeoq9I4Ncj78Cj7avsT+p9czqV0q71te
86Ua4Uu7pR0yn/f/g3awJjkSP3cUKHxUbKQ8zFAVb4hUm16x12bnVb5mVNV2k8CY
L/GJtBJZ3cX/jhtE4ESQlVT9j6yifLkMFwU1Lay/fIgvu1mY63yz413Uic/c/BAk
R6DXSksBpoKQsQjAICAjn8JXTmEdd2X4omCxFL4qGswUlh7ElaF7g977zaHTskJ7
JUoUUXAY1agP4L6IwkEMV66ackpNeaJPBrxazM5hGK36M/Zm+rYsBAF4cl+WqIQC
U8PnQgZ68nr3sMRmSu2+zJPXdwDme9Lmo/9UJeUVQyN8H/5IDelzUO3V3/VSRYjt
0F6yVZ1C8cBwejUW93thu/ofK7xZFMt1g21GyIjecRoej5BaSoMbFOXKAmJWDiRB
N3ujBmTKezoHpRL8n98H9VthX5pZ7vNEY1HpGAi6ndA4bF2zo5FPnWL8o6K4d/bQ
pNgGus7qeGVGm5o/O19s2PEtMMx8SCcsY2FYWtwcli338/eF3s+IfFApHbn5OS2u
2lOU8f/FiQYVgpaNuv2wJEIZIPvRCLHr4TZAZMAGqltUvQXP24l8HHhu4tPSVTD+
ap0UBuw6jP43MZKNQKudDaX+HqJ/kkkIqbd0p9LDg/W6ZKg2NCH6dX/TUilBflqA
Cp7Febwe1n/DPx+ds5Q8BE2UaB5iWjqfo65yAFOWuDDWXleSMuqQsjI0Ek7DVbW1
byQxR7uwOQjibEO1gINE5O9yat5vnx59iPS1jIRt3k+dlTkfmXb5+8mnit1QEUNu
i37dPKjpctBWVRKRhugykQzoKwCsrVWDdW0m2mwwuiE1sOlOwgTWmilqb9bxcBJe
pP1ayv6udSCzquYiCJGlTKlxGLtJvKmuQNxC5V2Fp9Z0R/e6dCRLGRkXcYCRNCeg
S5eP1GDPJI4DXJnBMoHlQNL3uU2ZqIsghzexEEwEHYf7HEpPU2Ah9B3EZ41i60KB
GO9QU3vndFteZT/9+dtJp/m/8g52FrOxYs4BwxJqzWTRKu5FRm17JqJS8vqp63i9
G+QfRLznh9x9FXUPPDPd7LkZ5o5TM8HcqC3z+QVbWFXaT9F/mUCpN3zyY8FN2sc7
EgpSM3J4rrtQ5A4WxZrf4Jq6cdCwBbKU/QCNo2XSb5FMXbudgLqKUDmXsmSjknzI
LMIYX/pRFwoLWkX5oXlJkOc1D5DcwpO/sdXjuick1FWKGpQ4cCvaBeRoG/f2oQW4
wNm1hWL3OwEMSqFIHxNVZjNtMu1cHvGiR6Lz/ZfREYai5XhF0NU5tI3ME6Bo/Dl+
lf+QUEe2IpTpEudNXxEIltvTPln6ym7Gezeo0TrQq0HLSJ17JglAhbOxO3v44d2M
gs38jYCmjnk7nTFpKFJ3DTo//BQS/eSo489KioasNrOPqD8DPjw+O2CHCEFWvqj5
UEN93ySJh/YriVAigJ65TVeElCD/IbCyMi6XZqJp/qOB14dI7ZqXut/CkNV6Qo0Y
pNjLTXil7a6yDp2xnKZno3/MgL46U+OdB7XBiINHaSNDp3KrfOWvEGG4Sc+I+wb8
ADvszGiDfEflvFJbEZYjNerwiVvA7DjyuZtZIJbm+Uxi+v4dGTYjk7G92ZKKh9mI
CfGx0gfFRcWC9JemPRsxcK4Y2ePpT3+16SN7Do3UcBT3iPOVxpWjem1JJgKIZGSU
m00xIAtlhasCJOlTsQV8BTNyKoUpFnSKyb0b6gitGy8+f5nMWGqvQlc+YFmj8I2T
XKxo/jiG7StDIKKULwgYmn4itfW4hhQt9JkxJLvBLye8qWBpv2FfQbxpEZjH3nwx
2cnd+PP8nSB4n4ejdjP7zdpA/2ELdRNqzmXIFXf17PsyQKAU/T3S5k4OcOuquG7y
npafvlkvE4kOjql/T1awcVQ+RPVznydrcFqPTEQHJqxaUu6+49iRQJCmlqGUs0Iw
zjXQ0oyy3y7rp6xFuwWo5/ZMCkDL34XEdASA52NjFF8medPr5Zi6vY3IlMzVi/3P
1YCFXL4W4z8uFxMGaAyVctS6Fpq0p1ao1GfkNfwjky7WAV12k+SOTbEpXkkOMsQa
qTrmusNQIxS1MB+yXjAiZtkK18cz6Y7lqO1dI0kzBEKWiAu1Oun+67TQ6/SSy0l+
hX2ZIDkuQu2CTfIxqT5IFR4RFHt1VKFk27mmJz+V5/TwH0nTHamJZKZYXARW1iwC
ySBCx9uACIst5hZ9oEYfTcaa5X1i7bNIu4Qh9yaDUTKQXwChYXTpu3sPanrxNcOj
NDzkb2wmnbZQM1kRZHDKC9IH6Xn0k9R9nfLimbd2/rDwTCPHKMi5jOWKorTmwo6s
DVse0RPQSTgEOeqmT7uwv0ZI5L2WEK3Xy+jQpePgeZoZqTnqbS5v9ifQBL44S9Li
p0N5j7rmJc7VQ8nF6eKJGwSj66ViUTnnQ//1BrZaBiA+w6AHre/4vj4knTXF3dy+
ykAx99rSFsh7Gfrox6dAi4B3/gj6wd3vDVWSaqJzsEupaWdTpy2HnZCzuTZh+pM3
uEtS0LGt4iewmZhofqnonuXncZmCzgj8FuHSdWaY5XkbnETpQSsFQDNP76CUbuc/
BgT0BNJBsV3CxL5ca21+E7/OpNay0tztxClNmOXtTJDOwU3E9k/WaIGKrdKcj5XO
F3aeSLL/k3+0rYVjkFBNovFkLXB5rH8aTh0kO/ud58YljOvNi1MY0KENHYEB83cj
OI5Babtnb9wtcI9rK6xOAM9lhCD5Js+YbefYaf+9PydZJzeeRIOlahSoVt99lEHx
vfYovnAP6VVGRthEodyIKCD4ydNF8p4cJPAwiHiObvQR0OZUCkXlfRECsmGVCz1m
mlbiqxN9QtCdO7rW5/jSsRAbXTjgNoFWu9DWvp97k8GfSLrdxRnzwbWhJpHPF7d7
GDviYE1j301VZgtvat6YvPNODYPfrI+Hef8RgV10qB+QVa6aby1j25GkCoHXJDWi
mLEqP4Llpj89lFSK4/lJ0rtfv3mNhQUmhK8M5DplxSP+hDGUEUOiz6fB6tvPezRs
CuTJbrPni+IR3afwSOwXZtQxRHaeXY3UiEEv2A8Cy0gC1+oYdG5D7Y7osdy7ZCOY
shV+H11oKb6JjWISbLjQsoxo/+yKtwdUNU2VwCZTzRrnB9IpWAH8yigKrJFcP0zD
cfYpmTAGnU1o5nqq7Cai1Ptinf7L5ZS+vXH1fCbcce8a/D2tr+mxJUGKcACCSYFl
CcU4Xd2Cig9vfACw9j52X86oEDJiV2b2uCVUgNKClkevWgQll+85OLhw7VvdI++W
U4BqdHCJPCIVrB7VsRH1/ta0AoWrfPL4+HOThMrnsC4PszgiqjJnzn5MkL1YvbcS
8GCM45xOSDDKmdpruf0VDC05XqZgz20LesB/5gAtKBzYoR/DHF9iEriA5HSNm+oP
LHhSeTHepskLFevkDXJ/9re+lueFKYQFrFsDwAeF0GL8nYjO4PryZKp/VaeMev8c
/ESBTX/lZLh0L+B9h11Bckl87xvARFTBzQKuSKMh/iLz69gw31eqBXeSXRFpAKM+
gQdm+JyA377jlR2JjETDNk9WIBSheYGy/B62811tEztgghrQGjAnMEAyykaYXbwO
BJtxpHgYKj8Wt0P79YTCON/Z6Tn1LQEDpBpSkVrd2Qj3ty8f78wKMDz1Z5Eb+DCi
LG7IgrLxlI7Ek2BZeAVPBcX+DGSh0ClPbrF/TXiqzFnwq1GAFCMfYq8Ia4aDFKLR
R3zDyS1T/q4RdXP812dvmBNYdPWVeDal3ZyH0Bo1VwW5lJ2uGmUVfrB8H044SQL6
An6qjQziQ9JgwO6Tb3AJ1+C1v9t/BdZXF9EopEptfjF78Nhknyzv3rtk5dTfOEoI
/wfHnw2D0dqg/u2+X6sTecj1BFoZ6jF2IsekW2QbdyMO840QsjdxJZLzy5Phwa8T
peGhPnMroWYc+G0rv8x2W1WPc2TlFlefnJHRzvqBg/Ns1DZvr5QV/ovGhYdJqCgl
yHjzGNZkqkle7i9lAEasF66nDGwzBjwzKvzH37UtzNDfLN9hyKYJ4Y3/8QYxSm9y
wzHgMSX7PMmzX5Ja3osRBXXiEGGaVQ1CpmzsckuJ2t0MWW6bBxeiU5Xx2Po/b0+7
Bz5QCtjaOZni8wz+g2ErsP2T4mD7E1Jok193oQPMTUBUODUudIEnLdcJ98PHtdVF
5V7JBHbwAVXTPUMVOgz/B6bueSNYeNAY8qpecmCS1Mh+keRw2IfS5mViGW0x/9Lf
91mM0z4I1NgRdduCmy0ZrPUtI1PB4IwTELuqFvsQQ77mIBuDtV8ZFjlztoPvhi6t
9V5Ro1+Ed7tMu0881kEvKanTOWx2pdut8MXx5gfXqB++yGry44rSQbO32iHDW/zh
Dt+vQkamVTpybmg9nAhPksBOA9N4ueXBCoPxnyz7SfA9TIuYMqHUr+I6snXYyTTq
ZbX7551S5Fi/MHATeykf9ukKmrVM0no+5Uyt3UxRv8QcsJaP7gwFZqKNT8lggIfz
9zYSHoDQ47fWXzNOPJoQkehitYAJrv9ew35T1d3JFNVDQxju/tnzC6L0V5Tniw/R
agsW074LYR0atYA5oSSRjz3Pd/7MEAaEKorp5p8Pb6eGnqDMsFyB+nYcaeL3wWQF
6TjDS4+/xuqAmortVgq8Ecr+T/b+tClccyZWjJHsUNhXZXZHePW8Hv3jEWVyIqTb
xiZm6Rc4ULRWFZoTAiMKFz3mxrFRXix5l8QY2HriBuHlP+E8X8yYq/80l+M+yWEV
UYTeAt4Hst2QHkVdt2e4QdBbfE/+dKtq5BLakWix4DY7vs8s/+yx/kFbi6hOehR1
ouCBhuSENmLP4x38/UZ8AgSumtnLukaFKWCRZFAJctWxoUWffo7QRcJgDZjFQczH
RPJZ0N18tNuiIzu2DG2Xj0/kDms1jivn5+G+l2blZoTFmIvzzkml/KllFrD0vlSE
TnNcdgKJEYMIbnJ3bgg4XfbNMM5tAyA8GPcfoxeoSqf9QOQiXLAIH4fv0Q9yLROB
7AQgO2oMcz+1Cwkc5tqoFx1h1jxs+dIpB/I4Rc9m1DolgdtyfRsUCstLZREFFfDr
j0at/H49iaGNCW+bDGvlwglsv0gDBJYgpOcuRZMo4p0qRtkl8axbUU8Y3dSTbJnd
iIY44l2LAVReGOEdkd8srRSzTCg1obdBD6T65YMYZ02KDlqQv51jV9VQn18il2v4
VS+K3iyIgb5HVGrq/nCjG6b5q/FzTm769PTGpl6WZ5egeoPkmYL/e0skHpfh5YGA
QcC7X77IbmCC97ABpZ6v4KCmd6n8KZEQRY+CrkYaNGmKBGhU1dqWILFeuPfnEXca
Q+uFA9lqcoCx5qwq5++5w0U3v36zRS34OrfYPE6s7Xo9vSEBvR99OLywpmOPfwci
jrtGRsSh+jJOh7PMLgGDdA3VhCOGDKBceUa46NtjDoqCpSFySqyqW5whCX+8LoUB
huyN3r4sBTJCe86hV1kk9usoChBZGJc6Rho8O3RChggMHvCY+W2D6DTsKEQas+6h
283TN3BECcDwMEf4JILcRiSrGV0ZIdkGsU0lZQtCcZpowjcUG2DcuzbVGbI2MXue
2+GU5CimdWSGbZQ0HUlBc2LSl2n8SJWOQ/AUhXstZI+ngCBp16RVS65S2e0+pBvS
kGcXZz1i8sNPLjYHDYrR+R+DGa6NVerSWZvPpaeIbD/G8TDcK9BIl3NnhIoHXIPy
NQbV95amzlkt4Im58+g29sOp/TRdt8Is31TP7XhDyTF4H1P/Qcn242wQc7KtySmk
wmaHpXOsOC8s7jUUytF8nEVuLJa4+6JagYjKWG5u6DWb/TSWBfYd7Wv+5dPsH/40
b5pC01Jb1Mwuzan7edL14yKjBSscGSnmRJsp2+71ZQparXyAFeXqXqK1nQI7WkpX
63UeCnloEr+cr2dcBLeEWlWTi+0shyNmznFNBwWsPX7iihdKeNIGDClpYokCWxuJ
5boVcLWShcJz1seIewTW2kmmy10165GpudIoO9VdnqwzGwFrnid/iOWJZHVRvgQP
z++bzeag6zeXeXBmytfDAs9iaeVLagLZq7coZ6dKIsFygEP2tLN8A6A/5Mu0wrWm
H9ZVHURDe7J9SSkEwrny43Cit5/HWlcfw8w/iFu5ir3O5xwUaNV5WyqrpvJkvBJX
dm9E7XISUMV09cP7x/UJMy1TIfSwyi8Qpu4X0eJB7MpGxgEqEQpuorYO3NsCuyrX
13sIFe9zJZTRoJcScWdlGW52Q2nBUBxtpePiNIKgvXm+zRsX+SMm6R1/bXGjn6Ml
a73+igXQidhlev6rL5Bu8X3nHoVynx0V9VBZh2c4bXsPJZppbDAWwTYSeCRuHH96
PM0XivtRrFFMiT3Wf4jxqK6Wt4YAUwrFOzxyQbD2KKsWb+wh6GXZepItTZLCyh7g
83HoJtt9kHjIXSAhA8Shf4LZgCeGicIMOtM4vJt7jgOPR5MFY0swGV0WO+W2xYHl
Qn3P4tajQe5e8sPJSg1HmxRv/8rU8hqMZMG3FzBpi0U3vz5Glgyf8e7wgskuk5TJ
RPNiIGWXsvOjwGFiJTcbdLqYZR4cSCmvoaFMnvJpor2D+IStEgNx/t0nJ7dbnBCT
00vZNKEL9CSZafgF2FNXTlydN/DGLOdWuZ0pAmGir8lwJZ9MZtWKC+jh0kxWW/x5
5CrIunqqmYgi+0OZ4tDstMRHHEf+dzhky8X2dtLHR9/RTlydvMTMoDT3ihBLTjDg
cfmQiaItgZDSHuXQZwXy1ZeE/G22PzRi2lptj36dccQ5D3nVfCtBsxeL7y8aRN19
o52wzFG8JqmJ8nUPY5DIy2Lacfjvu/Qo0vW1TtB3rJHvLw2jkGxsNRYwJ1I5WIAy
NzmGXPLWB+Gra+J659Fxb1uIAw/6xfnz8f8f0iiZBVtgk2Ymr49fasdj8hDhfasc
sqAE93AJcDUmtQl5dfwRYTiutkzSKfDVmR+3SSmJCTEh8RH8+1jLaqpBKOLDjrHR
4oVXpKXeNqgXyGpL7/6QyTn5Xyi9z9TeYQ8m1izVqu+ZYNT3/wv3r3qgZOy+0+4p
ZHjKyrtglmtrsBEy9ryiJsZinMTuSHj2TqfIToHa1AFfBFZniYXDvgqjVfrDhmsm
3hNkaaAsd78C69QjCP8PcasPnGE3jgrth69BcG6LZQn4oc9MTkEU64C0w6h0qFaV
w9aCi5FGSJVUqwqdnPr6WxAghIjCy4Zl8wYkJyv377LtKbhvmF4oHD9kjDOf7RFJ
qAQUd1lrycOr+P1qw3Hm771xD5zQl5nBOi2/WxGZFDFMHEJkA337/2COkUFqzUKt
8NTBJNhwny5+xLreVAJdTnSogDd67ffPIegIQVzNYx+Qrx+8WjsO843NIgqTjyRQ
6/oSIb1XXJ42UgH8N7EzBV94SUBoAjqJN+AM1Z3Q5fwyDMDXjf4stQJkuzjqTpQi
QncW0jW4dx2R5AM/Lx3MpSj4pXYZxM+v0fUloHCC+Wh4SyfOIhYs2LDmtd0dh5uq
c2rZ/i3eHeEr/5YA1+EgMX/WkJre+k4QEyTup0Jbr37H9wd6HllilufGY5SglC2c
dDLjvZzcANpAiv0gcGHbdA/MgB4/agCppVO/TdN3otRdNVenkGnZ1SWc7uur+MHN
GamePRcWPBB09A7hYAnDYAK5LFagvwsGkX3gbdo3SB9jSAV81twa2xIQDd3K+VPt
E43dcWi1XWYFufeOqLv9eMCZ7A1hA4fLrhuKkic8de5HxyRcvtkGS2jvTV159xdc
5pVWodsZqVgguGUAMWvAv80k0TNVbXt/wVVmtINaM68HPTucRKbnqhtL6zK64yyC
8D7c6B9l9eD5OUSPsPtKhEQs/9xbHiV+StxfVkncZfe0lBwoqvZc61i3UTtVVe66
79TJv1TxDqmuACS5kI9HGrqM3aFMAMU5iEi6qjxaCa4ADIBrcorrDgAtj+cHcPkE
2FcufKtMmRETEF9lQYdoCC9b79IZgFQmfiTCZmAfoWTtoe+2FThcXH21EMmw5k8g
C9nyMVnXxqfew657+XTDXzOmn2j9g/wm/qbkyyhYIcJyT1FHB5hzTV+MQMn+m2jU
B4Gjr8t/OgdL0eS6mKVwLVMHFkPORn59slFGq2MjDZCi6nRG6poGEcImi3YtsGGk
iYHgd2SMOd5FlWeO2GNC95xkflPXyIoftd64giNraPQodgpKzAZIWIHTa9/kG/zA
Ub1s0kYYecXZMFUd5JchkqguofQz+PF+bjLgpnVcLYJsX8rzWnnnENrKoNx85/t8
506UOkjv+/P/URd/op33Iof42lEkJinh37wnGrdzQl8KOlupM/c6YUQYX20Dm10R
ZBaVTwaOW+0oRaM3GcpyvIsVKjliYfUXCYgedyBtGD8Y41D9GNeWv70c2hJy3qAH
f/NeNjvp7y9jbmwhuU2FLLIv5d77npXr8mPe0yMyvnyJ1tHNFVDHidn0gfjqRxpY
j5T4W15aF0ITk8eUQ7I0Twud9CAhpwLkzTYqUGK4zKOVwu8huOrWR+uLopMx8Qs1
WdfBMigPeFMJ9b22uGJayCtsEH2bewA6FX1KrHaICwGWUXYPZ392iHwn2Es6zmHW
2gh+ElK1zzgZvuEGUVWywdxTJpnP4E5jO6/T3MNiIotZFAIhO8azxKbBwJ9mgGQj
Qniq1SablMcsHtSNplsdOYVmSQFzq8if0C1EjwYIsk77St90geajh4GualMnxAxY
n9axQwlJptS4xpJgvF/OZagybNxSOhcAz1fMl7CEYCGi3h3pFHoxxOVhQjZBYHF0
Wkx05/HtlcZacs7hJeGEU8UlYguK+L2v6ddNmU2tNiV0T1sSF83+PhrKpNzCHAtR
8CXyozpsyUOHWPj3YUDBWqKMNPdNulbxQIcOFnQE7vnILyDjbOlxlelOjRTLDltO
Rsh+Nr+0zHqy2Ios95EulaRFD8Xs+QoItIBC2QfxPa3pgUbe7rOQRUvK9AM9VkbP
mviUKI56bNY3cTHhziUw8cA/3gzz2Q7jViySu5PX21OYn6NEAUitpC0sw7HNhekS
y+fUnjLBijifuykZSvJgfJMdGBkvIKkwgIm2UP0NzU3NLk7tFzTPE7H6idn0F2De
Jk6ES2cBK4JMrB24z3XTWJQWhLG3w/Gg8EfttPr4liDiSGW2gIhXqRC4incPNpm2
T1OXUWKt8B4r5xNGxd0yNne/VzzjNNSW84H/T9NP2Xc7NWl/SZ8BX3ExKcmMoUr5
Loe83V7AdHT4Fg2aYerPyBGomRlkWxYn9mnbELTTtxqMxJn7SaP//ZZnAznEtt24
LXdFXAElIKV+k1v4edp1UwDjnAiujE7rAQbWhWknevpJIjpHUfQg6mZbjbtd1dFc
NBa2enUT7M5MG+Ls+bDUkgXsrWgRgXnRBfm6fR7R7JmleYPgrwM1QdZLLmgGuJkx
tovfT4uP9N7v9f3dw3gtu1JRE+aSadspHQiPaEHs/tjZEuBpEo9A1BrVVLa6l/yW
FVEOznLSFwuZ4Bx85T4mTI4FmHN7aJC78vckjnX/aaqtftYgcDHWcbTgUghtVU8r
K4aUDRM10Hmy33VGvFmKj0v8o6SH01ZltkZRVdwoQe9MB/sjhwXu9Yf/RixTfXog
+D/vri9FG/Y8vHwMhAgry0LbFXeN+saOzbZqyPWDn4VTRRmwyxU4EISmwO5rymy6
J2Lj35tdVcMv6GHIHQO3CD6z2kJtU42mKxSSO2GJCy19/fZ7VvQ0A9M/F3p7TOpR
4PgI7Fg2Lt+bdDTRNUYmYGBgM27X03kQ+BAW8PZFgpN6zpe3thodYTAgp0ELGzLB
+6Dc7a0HVgVy0lB7AdTFGiMElmCgBMmxkKf7g8t9g8wWtBcWJjnK4r2FgCX/+HE0
7iANLsqAUbGg6l3qhnQcEytRw6WbSgdNikeSEdzFGow6rjdsQgJk6YNQmY1fUBY2
lrdQQ73TAT0p/WSFU21UGEYC34lfWzocgGJA9DBw1aOf38lkQ3t8wWxI8YJSG2BS
jZtOyB/vBb0EaMAJ+iI+D7+AHPPY4m5TIyR3Z/CQydBVv7T/JmsrlMuU1jTWdV7e
ysLlysByhtc4Lw9K1cDYSyAMLNqPJ69Oz5poChbgbO4rjFfKdeZFqp8rLZxmYEWQ
/dOdqBneObIOuJqiXF7znq2s81s1/Fz7ccJ3JMPRRQqvq1BSl+h8Y1zxl20oQQbQ
VPO7yunspLTC4W7YOtwYwmSH6qvfQDpXFSAdtz7K9itU6n81mOnYWeMMYpW44SGo
NO4u2iktcJTJ17mZIlV1PrYoBrbuwruvM0x2Jl0BZLzS9H1LhtdAeF4PyFzQLKeD
GjwtEBEUj7EAhbwT0PZVGPtnYUaPjmiZ9yy/a/u7rL9lnrH7O81xuiXIWDPCczC4
wGsBoyrip/sUT0BPCq/NEe93lTVaRmjF5nfxlCPyuzdRozl35gfUW7ZpeiSZdWuc
XWYQHNY+1GxIEx7bJkqbd5hAyAF5Y4q+cx1T0E11ZOtCBWzLE3S62jQJJcCQCXuX
nUfet5XcE+vyeqOFmCwOZkaW8xEnxla9j2C5r6ne20yQbtkNTMGNypowmu519G6w
Mwh1z7qqp4xrub2J+YQkwf8PDL/dHH1Xe74lDD5l5atzQK/P61kekoz8MdM+9nzG
EEXgozdQYS1Ery3vSh64l6Iok7N2vr55OMLZr7OvUVD2PnAUV/Amx55TZui3ZDtm
PJ6EaQWj1GalZ9Yts4V0p2gyHQr0p9yIAcNWGBUWHNZeyWoG6JJPoNgcudruK2j4
9A/KarHGjpZdMCBXUVdBIBG6xnOlZA6zHoQ5MWz76mzlQDt2EV4JybgS28QsjrmW
kdoV06906gqiNwHhmY8S1lZjs8iHF4y0hlW/1Hj5kgJYOS/oG1YtE/GIbpCFneb9
JS4WIHnwMpmxP4MvY50UGUPiXYzD3QlAbuzY4bai/Eauvkm+fWMkZnwybnD3/ekF
eIU9NvIqGyscTAQroHZzKC8x9ezZQLInoTm6z0uo9ofg5ybtP0qM7E73WF7Vxnku
Wn/pcazAq+EJKtEffr08GyjhEgjUNLZWxdolG69333lxOpn9As9/BZZfIcUz7x7a
6Bmtqag2dDW23/Oh7898NjMqDZ4hd2CUSxK07u4v60j5UcFnoG2UAr0M7gFtfmdp
uKtnLNp3IB5qJan5YXqgDhyXLh3nu+E/edhm/oqh2D5wxNkuXuVRQhFgtvXEeboi
T1Q3tBKU23U7qVMnb3s7Wdb72T41+bDMG+P/bdWs2W/4aR/SygvHrAxk5B5m6L9B
B/a7QLeOApD+Xz9MsFF+lYE3tukxSLf6+5NwhGC9nWhxuAvKEM9C6wqGv7PjaU5t
RWv++I21c2MvZV+A4LiqyuCPqAFGVuU4XUQxzqw5b6GsOJ7C0Q78k1hzOtqUnSCm
ke/LpQF8BQP9YI3Dkn6KP70bUrS8iYj71eA+ivHxHKBLX6qbB0R4EzWnl1bgeukD
ZYYIjCI7JvjxztoMFY621qLv6QOvF5R9nnp64uFzSAKCF5WVB2VOt8oRYhv51RB5
Wvw8b2uCLJTBXcKMBrzFewOn9gtBoNzOWcYKvld/R4XZxq8QAKew3r7CGV0ANPfh
weanl7/JJoYCxsZfOeC4OH7xSkZNM3OMZHKMUI7WALvj4ZgNIj86EdYponu10K2B
Dr63PUO0H+a5dPVFh+m13I0Jsvh1vG2HZqbe+rVxqDwStT0I9HcZbOPxq1Rqom5g
rIm7fyHp/EJL6wupfwXrP78jYFoKAVhNoB3RAfgm+rPLHm91LfD7Dknop21Bv2/+
2pI7gaUB/QOGfP4Sbi1h1qzRv3o6mF5+jnMZ/wtDohfOkPLvLRcOkbGdRaLEyRG7
RugbgVCUF2r8AHdsvOZcVwr2bmbNy5/oZkjr5e1etYPKfL/Y7EeLV8MwsrQ6/Z+/
NdB2TLTbe4MfBXTuqVYOQrj+tX3XbyZZ9fJq637zm0/Z39rkanVgY9nRVhHMq4CQ
gCWCFqqIWR/dDoPZRovrvKUKRudYQk6lmJPjeEio5haKoHzttpkjdeOMB4qzBxJf
VMi0+6b7v4PS/sVyLEwRvq+5dVlTo2qgLxJ7UzqdRnxusTbbbRld8Yoz0/qQ0AON
Gfois0lVJA0JZzS0VP2peU+A4RaXKLxPhySs89Gl/09f65K+J/mf+HvsIIA3qjMI
KcxAtoujsQpHsvlf77dxGcdnJZ/FhIQA9jpGsn5s6ddfsvli9jj47wa01DwCek9i
QoCIN6eVVsKTbSXQ6CyHxrHEt/WyqIAatnVtXEQpuV0OLPcgDpxxbPZI33R4e1LN
SXIs3zDQBIfzs1tUrU4ouGRwaf6dvLEC7BmBuIPxVxkHJzrAT1gDFPT1pNPDo479
90MB4kfSO9yJ4X8RoQzA7mhcJbSymMSluvKHdH7RFTTbN5IxGIEZMb5bfdq+oyVN
X/2MCMiA5Yg2fIPIyh3Pn5KAEsic4ybdMTU9WYESZSTrmjY5CBxG4NZe88pvcBcd
15w0gANteEWniwq8jllScif/VwrQhM/AyqlViskpd5d+F/GRHZwvgP7w1Aw1fFHW
lLetdyutih3pztw8AssUekqxM18GDUlTlQqVAQfKgd267CibvRJsxdZXmSYa/X1l
S13r8wEBmgkqMXuXqvDhdmOiRU/K/Jy8U9FihRwIU9gfjSlpdW9oIdmXIQc30Lvp
ATDtj5waG7lJXJL3uGOWizETI8c7/PI4IOo8/7jDLF7UY+eY2GTtxpn6hrVMDSpQ
U/+7SLVEWMuV6AcMv2/s7+JALyDCKLkHuOmJqGPTxP+8+1GfA+899EeuK2dWvD6p
MZdH7xBdTh1S668pNUfstFMI0y1MSGJxEkqalwfUv5LOuwuYUgPbZ94K+7nbjiNm
5lG4qrEWSX24UR2LUJKNHUU2snTauSTjc6o1I1Q3CfGwZABH2RTzHGoSwaFt9/Dh
zMNsfHfyWifAHzOr9nQkobV9Pso1Ia4p0nA6X2C+t/TzTgKd8lu9BlyDqsOEiI1I
u8cJBY7zV6ZOQNZHWL6PTTC8mPzwMaO5mXvQHB0Yxg3L4MovM9+xLPdcA+yrLlFP
K2Cb56tFhf3vNR35hsgD9VXMpwGHUpjZUvmONx45TgECAkRemvKIQ2qTHbUhCYsl
J6Qvei/AA+2YrZNxueaYJVkVbMsrDvXDvEU/GlAuPiGMJDr7JlB/s3S6NgoTl7xt
lpYgEwdNmOZrTAUml1eZrLS4ic1iQ6VWJLBvwfLZMUWdkByfexI+e1d2p1SAYhY6
RKSL/fWSgOx5sCuvqhqhsszTvFMtBmNVVWNNYb2WIFS5JAD7pHjzJ2FSfD63sDfp
9xmz6mO+qUsnkLM65j7v7w8YNomQwvJvEJkGAJd5mKA+dU6OOZtQRZjI8nOJ7DPd
RmS8HQLX1bRNyZ9BJjuJqaSK8xWOy0CZdrv0j5HI+p2/zt9L5zE1YBpZg9xntSvG
6wNEIAmRfg9uoFZlIDObiHVG3b34ICwf8iu50+2u9t6sRKoJdiDG3mwTp505oKwN
ThNQ6AlITEWBHcPcbV4Z6ACiGUiAEbpmh+vdIL8eSJGuASa5TYWBt8HgTj4ngVnX
M0DXhASyAYB48YO01w0tKSYMGtBLPjYh9bAfiik/kv0IZBPcBny41KZwlcpnEvDJ
yjM7Y31tbiIqrN1naHmL7xMwyz9ZIx6NxJtfUfr1buLwtoh8R3OijXm9H+2zgM1V
xZRiDFmyWxH6Wp5QbrNvM//aN8fXDG1SS5EKUNQPQYKTNgtcbAKfzGezCbzz6Ycp
HKRQ/SQKampNNwgMm1l4ZGCBvkZzb5OrhL4/pNcLVjuxTgjz4StinccEitk/g/hT
oxcmkCTAZW98tEpj/1Qeeev7sf/aKYDt09YDuHMFG7UQeGaVTCmPLo8hLW3Ol+IL
/T4cttstvfzKVFKIZGJc015h/L4tpFieAbbW0GNg6dwhQnZVcW1Lew4WWB8Ks7QW
cSJH8XpzLl8Y8DXdxChN1QF+w95cQStjBU9VaDJZpXXsB5lWe0EwszjyIVJ8OgWB
lGoKgLxldnlftZJrJ/bkY28d/QDcufI/iFxl0HoZruNm/ZvVzdOQN0iIXSyLFNe5
qMdlelBOmL4Tbdv6LWGATQN54/y7fii11KL5A3fBF6SzfroAr5FZNDnw6EjjIKSE
jTf4pIyoYtAf+hIWsU3PE80qHGcPFS7EGdyFhVcwCmicliP1qb2qrPEdGs8yRcX6
SI8VV8Kn+vfTP6poC4NtbNa+31dLMGDh8JPP6bDuYRIUw9RT68u7ENl3yTaM7qhe
ZZTmdKwIpXkaaPlHAlSVIIlzWoHf6FOcJwLmcKgiEvDlZzBBmOGmLuKsZ5Kcq4iO
4/lIUyrd1d/F6B+/3oxyF0caJ7kjFN0VPM3fjbjPro8f0tBTpcGWC8KIUeMb/zMb
ypphZl/kzSIW/7LSfUz2PIVjNwD/upjtk0OxHIlFUJZIAOjhcOMERYhA3U12B5Tq
hG0RcZthCi7rLxxrbZeIOrr53RN0bjf/FCe1ohoInkitPnKpuYNo3B20dmLMQywx
Hh6ywUGzAGGT0dqEhlp/ZYwK8k0WZjol+CPliA1K27Tl2yjiJ1PdicQ/dH2x+Ihg
6nZkoa49h+trm9k2fhbH2+XEZqZIGxG+wDBpCjN5zs8T3JeTmQdsF4mr5C+Jp69I
MO3iAjASHvBHMk/1tkICFgmJw1eX8diqWlLQRkGBEKB+O+3A7T8DZwlY6Hx4whGk
qdQZs9mNpRrdC/abcv9kUQc7FrMN+M759c5HNag9AoUljmK0TWyA8bjYW0NHTR5A
aX3HndPKVr/MAQq8Liy0tZHM+s0KKEZIk98lO/ne8m6AX2A82s6DzdtWLhrX1jqK
+BNA2OkZakrticxpjYHF4BRs8Un3oQ3Uvx7oRe5LMaOvRl+JoWGzQP79vOEhRJ0/
1PW/VJtdJzyn0wZv8fRzy3VfpcNQ1R7b/PRNPoisX9PstTztArhf45yvD6WKB1qO
UeVeoxC+Y4gKdUtyLBraid6hl5LcAx/hZOGALrFrw2l1zIPP/LBKJVtA9orkr50f
WjB1HchPNONAnjp8tF2YrP4I784g+czcf5UhjSBRFelYYk/zdrHYD0gHQf5eyFwT
6FDWGF0JzIbvhhwmn94qlk/FPpDNTg4IQ2v3TfAlLv4kqqNlvF3nsvV2ea/wkuRo
KrK6/gSJTY0LdH8sK1Aame9W9aJXA7Bna8DBC9687NCcHwWAM39DqKvijVPxcvax
SfKb2uzYw5oZo12uAJCY2V9vUCHGy+TpdQXHTYFOkQ6gU8skW3n6VdF+ZRuB3TIz
Wfz3yWqUGcePGep1GtYPgmpizylVBmLb+spLYZEb62RgdLYeENM1qcgDJL9NBrfA
1qkckG6m8Gf6j3Hcz+vRUjQd130Z3+IBpcCcy041zrHr0ZZZWGLfTmNzo8ETbdrz
mBj0MhWIFc1GOU+stPrsslG9dSVOXrS/V3JPe+Cw/32BH3ffHPCggZQ8an0+cO9Q
LEe+kZUBN29EiCePWk1LFmWrDWljjhHg9aa26NesFDSy+5ZKCTjkHHsCb2sIjpU7
Z5ld0YKt12Rx5PTkfcrfoCxW/AbyzVpes+L12NGDGsj05Brsa2/Hd3KsQuP9KXQ7
fEo8/pAc/yyVu8yuFwK4qNW2Hrl2p+ybPAfkF5SxeTmE0C+Yos71b1cuS1kuIgAI
rnoCmn3mTu2csPxbGfBzobPJBbAuFXv4hMb7HsN16Dqghg1syHm72yBKB2TkyKz7
FAcQS+U4ZAgm42FkQWljxfLcsGPXVKrTuBEssxityKnfHrf24ue7r1ukY47N5TlZ
o30FDNnlGDGxeWbSmwKA/+o+lI5gaB8+mj/acBn++pJK4bq8YqLYgwfNn1W4ns2Y
w3VOQgbmMTRp+AoUmViJa7KZpEBR3URhUy/f/qQQpJv556/4N8qsk+2Y3YExdfTW
Vg8nywNx+QO8N+KAkXM8XiHoV4ByCNJ5B+Rgiqp8odflWeA+MQn1AmAAaTHnpRun
d6kjEU9NNhuMU3TYR7kq61orpHg4KdzY60QX4dfrANsHN9nRtZ6ckuQh2hGnETOD
gbxfiY5Jd/hNLoc9HFQaXFfC273yPl0aNkILETRF0QiiZ9O5EExMdF4Q245b8MsR
PaMg/uRZtm1HizEahBGGKhFLWYNruu482q04hiGDR5wAQQEUT0lAqNLz3TIhzf3m
wRoCQf8XfLAB0kE7KCOuRdW1n2LhbO9VurKa1toG2XV/BqWnv7f72EbJsZQENzyT
Bu8Ive45DCfoYgF5WzYvH75YN5jrDotFWUJk3mVd3HkOqVGvX2Dzsg+bx+KmHz1P
u38f1R/JhOgYHejv8ohxaVDLWh8vIlMfYXjGKR/LoYTKmcZ7iGv8KQRygklizPnY
dSQYg4qAD39AN0gXog3qzz7CWwjRJLzEURt1hj3YC7MIvR6YB2mEVm5MUiYQ9NOd
i3ATHrpAAVeFLrYa05viBVvqHmHGadRM8jn37uxwme4i12kAtoXAeQbuRLpFdeD0
YLXb4sm5qPJ7rxIrHmsc4F8AQNtf6VvlMpAdDm9QOOAH+V6C6N9+g3YsapXP4Ljm
wkbXLqCY73r74CfV7+Ud3jrNAkG26ohOU205D+B/LbvoLD6qFxBsvi9tTLc287im
qE2ZHJZRmkj9KL+Hk8XQCyYh8a829xthIKzv1UFPCg2HrKXmrlAwrbYaf1dNzZ20
AiCc+XAMTGxs/V/Id6rbKrMGbNS1FNMPou73EX8/2uNUgU7ki7TyOBy/LZmEBTGA
hk/4DCIyj/0BYe9ceV76nz3Hx5H5QJHKyKXNLkx3gaXy8ViFwNVtjFkCdYqAPF4V
6jzbfBfqWQXubzUmPheVD7NfLWYqAh+eSJjWIRkxwSbHVdq6LGwu6Dowe49RCYGH
mzmGDjZA5HxQ4ACjSHnYP5LJlhdFnkNR0+RtBoYvYbrM3V9rf48tIbowW4u2ZkGl
XTcmWJekiOjJqYf0YaqIP2cuTqZoNbMzN9VsdrkldiYbb6UO1LLiWnQrzXoZhibl
lbAnEPrlERL2OzRrEdpRr+kgbhCySIQfHuFULgEhsx5itaQlQQfOdfaGQLmP5jqk
hUXLpsVrRgQxFsueoAmlTkFJFPY4B5sdxrtLA6Qep3bd6NXq21bvSlM6PhPvmWFd
+gBuCOhFwWOendjBw7py+IkJSDAsgSJLgy0K7sVRVuNdLXpSNE1mA2/zbNKwggiV
q/UL13MVbDz/7QZsGi/9nKINlkRZ095I4+J4AoyFAaPjKUWlIE4LnM6gcxjTVpKi
PyEKG2dAp9cHqSblhZqyVdWXNbjiRwlMd4AeiD6iTBoxqyaaEPWrE4goBiSPd1h5
0Ix7+vX9GocLg6X2Eko5cj3NJGzPvrlzsYSUyBv25wmvU0jsTge5HNyuZrHGzk5/
1iJrjKuAQBPuOL0cNp8cL+O37ivTFBxThkAeYN4tZ8ebrVoPAqy6Se9R32npVTWN
G9FTpyeW+In/fekYovR42Eu4c16pn2zRh7qG1TDNl6xsrswcEiWzE1J/7xhoE17o
mjx3dzmdno1m0KiTTLfQ9h9DCNLIwFnRQlN2PhPlVTzu1n6f4iNu2GBQKwHm4BV+
A6dxoku+9ByJVKNgFVNdimwvIPpxUqOjP0D/F4BYPY4naWrWnSZ15NGuKBqzEUZF
aZgr7WGMUZQ0WD+GCGVwL+KMhXXLn5QFH6t9gBjoA+xsAf0mdumuPLRgQ6/mi4DF
KBgsXpp4baf4uqlvxdZoOxk+qMN3XOIMVI9WndZNQt3NVyhB9tYNxZ78FTEaNsYa
uYGXJ//qmdFRwMm6l/Cls0N6CiZvJ+pguBcUeSVuvTd5zVXAwfmLJAgiAd64Yt+o
b7fOCO/Vyj55BmdVn9ibfjTU+f0oi3XxGTYBIX5iEuqQKB41uRkx9HFf5TdYtKJ1
H8ORdqTN7A4CXVF3TNvFiY8URHCfUQuSBY9kO4cY7lTWaUxq/d7z/tk+zatBgfjL
z7HIxVa5OZxHID+wGTvwq3zK8fePi6EbkkvtAQCvM/5wyaTp8tQJ5FUOQFObjUiU
EqtuRJFWZdypdtN8gxvXpK4YoEoCytiwHBg8m53LzMUm+8JOQ7OmvAO/+vynIJ7a
UvPexEpV4JHK04pajiGilfiWzLxq7aLQxrfmf6YGugdUIr61qObxlKPJSCfcVR1O
l9xr5U8lit95gBmykPWRlIzaZffHB9lHfQ35O4blXExeeQ+R+HlijH7Fm91B/9zm
5ij+NvE05dQ/Tlhitd0vPNsBzgEXcSZhuaAcgFWz9j6tYimkbZLFgTJJ1x2ZM0MN
W+CvOD5MQWyrKyUJ1mLVYOoD8AGdF+5wVldVs1Z02d/i+XgTvMCE3/QAadSdXuKs
+ucCsyPjeXyGIykZJcPwLRFPd2UiLo36prL4VcueTyM8Z1654V6MfjvojxW9OLGX
E0/oLmqkocifUOpadPMnE48EuYuvZ45+ZP0TohDL5ujDDspiVjqtmj3Yd4xCGJis
KF4izqOrmJWBcc+AEB0gFu2pNQNT3r9znrs8ETUK324l6I0N1DK1sjINxv2Hhhkm
HYyE5XzLec+UXCUaqE2dWHkwuHowbLvXMe3NEEryaesOnRZ+gmeI1TCVOV0UlPvm
mVrtryK1Z5XFSTDLPdQ05Na5zOq2QHjMfZcpYOlaxPBR6URMZK6KDFML7e/xCtIC
35jUsyZ4oS7tbV/BV6mPIfNZtPIhkIX/XQqWbaErnnKIPeFNQt8lEvIJvIT1lmP/
vLae3IMDo/x+0Q0Dn6QV2PdYtaLBpH3+7uiFbUYMLq3xo0VgwcTJE2TWN1sinfhy
NkVAT09jhmVoXtpWVmrSkmanqKVpurdzVC9Y4+TygCTsoZgKH75VT6y+4/VsL9If
ckFnrIPiVRfepdFyVVu18HIZn4RAYjM2fiHGSzkoXWSNWR5UVvRX2hqdp6rhHbse
A2O7TkuW+3qtMiWJvKxstC9jNFWuYJPIwGFI/5UebHz7akPRcLyuazEi8+/VQ7GM
QnaC381E967zlBLEkveZ9i2+51/TJCsKNAPuPl7qw0+MgsCCjNGmqtCST3xjYus+
Aj7O2LuYU93yA9i2NFWkHxvQzke2oOLhrQxfXwZvxc4Sc8safACF42Zkzk6NDpKi
/r0edwqXjefbomaYHb3VKw70qEnI1AppGZ1Vm6urRhZR4tWP1itUFqX/rMk0fFtm
+Fke3s2HTOHpxvMgL19OsLS1xGnC4XQ6/KKdxY9EARyXxZBUMeA8khhyjOEAaNLn
xZJTIL5l19H8d/IJQxO3Vt4efpzGtdNUGHT/8e84NocWnj34fQx5ah3yiS1IlBVB
UK33s/ph21leWf3ALlL65+IcvktIRfl/EBa7n6OQu+uO3V9n2H8002WqFe0yyDah
8HTfhOWhMvMEg+ii6d2P0A63PfefIPvjGwRLNIQK9EwKolZts8NArjuoQWX42Rkh
XraN6eHWh7xBau8wb3mWtvSHxKI60Xrsj55AlX1qHiTNKAUmLG7zJLHYy0+IW9wJ
aFdNsAZqS0JB8F7de9S2L1SMiwvj9H7/d0W5+TPuZfX0nndbm9RRL4dcsywiyBdR
i6i07YufDx/SIH27FAG6BVCaVBWiAHEV2c/SSFQ6hgGqmp8BNhmi8IEAw4M+MeWU
k+Z83FsZc+x8ISZd4z7WGz7LRW5LloUhhAbsINGRKwGBAX0zRB+HEvK4sp7d9JMn
omDIFOR5bC1z5d41FUoLAtUy8dpjfShff+hQNnQhdEzfn/TG2PYO/74MajM+T3Lg
ADv0+rHRsYmF9RvVZqclO5XubxXHeNqXIQhrMpxvXLKHx/sstCVvZxBZJ5X9Tdf9
05M2+zMAv2hdluI6r5GgASRCRkBJyCqcU+6giUnp2TealHUcfB2XuUPELFqJrUn0
cRZbgoVv4y3PCEueJ1LqgyggsEu539IhC9KZ2t44KqoG02w7SSaAmERvlWSivd/0
m8rDhBEVHcCW7L9QucMaACiAc8aaTif5i9GquwaYiS8+9gcP0vXb/wBSTlQ6yyIS
BG7npktYCcaXyxE/mO+cuWNrPg8hgHk+dq4o7s/aCK63g4rg2g5dyED9cDqsNF+U
k5WcbxKCPxKjMsOO9TndHaPle8FvQt3LA+Byv0JJ3pN2PijZ1rv4O2a7fv9IxRgA
LkLd9YfKaDQp504WYvsu/M9EFHzhaHaG0//kTZshqJ0Pp69fkU3gJ7crzCasEu+p
2JqMpDDLONxvPx20WS+9JslDJRJbJaI6HJ7VJ+viM2SqF5Y1+eSwrblkXQYI4TDa
apOCchUuPN8O/zVSzBqPKGxYkiHTq14RnC8r3jUqJNPgmAH/UgEqAlw4MuBdfXbV
cOyBudsI891vGyCRkIAr5bi3yYXWrjtZ9ejdfLW+hv5P007j3bjmW9AOSBpoPRuO
EyMlWyCchKsugDk9w31Kb3jU97zF63U7F1LWctJIjRmxIVMQ6aF5kcy+Q1NGKuq9
hB/YC4RpkHZun0hHoD5xw7qY7/mPmcGdi8II1mHIlpTZKJevs+vutI55AwUobrsi
90Qek+wtJYyG8TWEaSvCjRTuwdzP+yiaFJOEXZeeluYuOW56PhdXByv9Urfp0hfU
sLWPa4XZY9jQTWk4fwo8H++4M2j9uBczWTkPydkUduLQr9k5sViDXhS0xgNXYKve
yrvcOXLka4UMrpZt7oPlW8aMVuiUYr/ktfeqR7r1fJFKzowcnlqwp00RPffAXs3I
3pmhltcmDHaoh/sN3SoSifBMedpGCdExX13yIkPU4ULgxncYTmUkixFtNgMzw2V8
W9gEZWokuXxB63kth3Px9wAG2LOK1oy3iw0qMbrwUM6KsarjC0Y4jbA9krV5YDkd
oriP1+74PWODKkx2c9cUUAQhVeXajBqvm4myXpKi487XqyOr24Yt5bTWPGaRiNl3
/JkQk2G8vCQIV22oGECK1sF40+IIeg93rx3XumjlfuONm8rc3v1sriVmtBUzU1YT
HVF3HHBfId+waj6/uocKlwSp9GaOdbxK+CUZE3yL9GoevzCNSTh8NJzAhjOC83UQ
mRxzJQJE5QRwomkhzhyw5coiC3iOFaaofxY/7HF4wpw/R+phzywGZLYRYHZfRkL0
b/BRmDH/hJtulrc3U8vAkITwg/8eeG6cFtsEJDZYNh39PjCZBeVqGSYTTAGP+WCZ
Q1tNLa65CTIxKDYxBgeJsYP2BigyjYhn4hdAutcNG0eMlxcJb895KMJkakMGeiIJ
ZiaZnmrZiUm7yTWdTGXHiOq88ufaWM05lAdrkbIFBL9YBxKmsJgi1QGDl2MoEC7m
f6reK/zbKa1C/8nF/6umGb18JqI9wdLUsDU3CZVlncBcx+Qi3gwDrlWQmFIjilz0
PkuZ5eN32ViJT2NzsPlPfpnyXWX0P06AK4zFVIjwDF658BGRhE5o4yv3vNPJiqlA
fuS2eCdWx0nkfdnJ3ze+RZ3yr9L7tSEALrCuehUkKp5qx8epzx5LJcf7WVB3Bk0/
0xwpZ6qR2YaFtiHEelxTxQN9pRRNXkmdLrxQMTv2us+9xgzhQ0Nv1aKSuDIjzWr1
Xm/EUmjfCndYnxiNtvZ0qQ7Fk4tKblL4PyXaWVBUiuGVnQZmMojfjthUHoUqZt6g
rIT3dv2q1h9qmYPvWrcDcFI+0k3C5APGtMsOkyvNtHMHrh6lLZ2Ee3gk7I6cfz53
ISepQraiRxrYb08aJajQHteE2vzMyx6oa4e95iIhICQXw/F0cE1bpA4q5GsMbMDf
7OuEbem8XdmxejUKERRiLq46reGMqpZ5lmj3W9YEfGhSaRtb9MVzZfRICOUDuX+i
spYv8MxMKjhJ3ZCSX66HXmMHLxOQ/y3mpB7OyH5Kv9fqpwUISR1ujZ+RXA1h16qr
YugplYurPel11VbhBvxsnTvb7QYm1ryu5+4B2CQj09PR0kxjWjAyDcqSajAXeo2k
PkPL1hBP55McWWmUAOx2fzyq7XJxddFGt0hB3XAlguCmetV2gabwPY09oQttk41c
Ap/mXCjOL8IlHhjpOAgQXfvYa2p9WFDm8iwndk92aucuPGgeAOA45kJ0FcwzPXmF
2ovjxAP0ghV+spKWp1oQfIlcsxkwMfzkRMOY4/dfg9PvsVxNz7753+K//xaYOLr1
gzu3z2u7PeYJP6uA2v78ZZpA3wCie0Vde+JCq1qp/0dcdcVz4+6lCu/2rYpZkN29
UPQrJAqRwBXphiSDGiToYEET0DoOB316Af0T6giGAI10l7MY+j7XXRmJpUmRYxo7
DcJ3fpEH7FbGzkDRJ7kkfXFxFKnX+3H790641P8VhSIEFHvkEV3Qzc4WVGn1e5BX
vgknLCKI0F9MWYTjk9bVXTru0eHSrGhr6kaMBRex4HG95dtMq0hSzbguSJUy2c0a
2fUcs2OMl4+fKg6F5TvIUx0xWbx9wVqioU8/4EVBwJs95B1qwil9BNl93DPojviN
hSd9sLVYtWEF5BcmzWCtg+D+FyZ0Qa3W9rCNw6GPmMLYjDbi+p6GKUdO0v52iJQV
1+wRemKcxiqGf4z/4prDkh4JikFA7tQa6BRnYDF0IVlYon3ZG++Opf7Z0AFjh48A
+RgIVy7J49zXOOpz470HyN57Qe370IyYYHwZCdc+A01HUyzwmKi9QTKIqym7r38b
g9j7vOwKj24t63Bn9ud79NPE6PyiNCNnpEHpMokWA5bjowUl3W9l9nAk58PGIQwj
B4lDWPT/TM/CWKeXM5q9G1PegWBcJhSb7S/4NNCJTNvdnb/vZIx81u6edHAiB+ke
au0K85b3Ox6K8nOC4JPCmXg2PgbiCcZCTpCr334YZ/cAJBGTSaO2SQcQN2NUUpw7
G9V818oQKai6vcTVpTvBcUv25CpvNkTeT8vQCf9MkG1EbuC7POLGMnhHsVg5GMNJ
vvyPgunZQ8c73cEexo03oDZZGBXuH2ksICaCtYSnKqnRAPdwKIoIcSvxvsr5UP0f
43wb35E7xru+e0ttfMtx3aDz5mUIE2BHGpR6kvPUtn4IjC8kiSMY3wEH377s420E
hXl/gpLRu4EkgHMwYtjk6Utkocb+Fjuawb5l/srlmn1W2JSZyV92xWgUhRs8Cvj6
hrfjrDKzEHtaDl+ZGUO8Od183k6tEHIF/KGobMpbwJCoGRuAPKcq372ChmGgFFw7
s2FfRI3/paJz/1uSlWrOdtniNB7l8xN+oTEK6pwOo2wrEe1GYpjuuz3Kk9ab3FdZ
W6uBtfUCktSwRC4SOEjNsAuZxpJv/+T/7q4TTMGvFWSsMsrZzXQSIU4q9B27XaFS
utmMzRJV7Kwjg3QuqNunsyKXgFEV1s+fDDBTwQ/bT8LuU9FmIP0VsD3x3S6xrV8e
bqAa9SlCvYXZ6Nggg4eeJLuu9BDXF7IrxK/VzLTlKhFg8mC42mlBT0qrD4PLVCwN
d9U6zXrutQ8MIavTm++tLppM1PI2E6+VxFZ4oZ/aJdHa6R7s0N7mrAMqWI64sofI
11/sX0gvyuO99xRsfLVvRWjvXFfWmIUpkDns94CM5LjjpznScsf6xrC8qoIEQkw8
7Fg+BFJoy5tpPVZyrDqZkiMJpwf2qe2NSMeAZNjOvpTeGumZuo4M9WH5Pr+OTRM4
sMSjSZE4O4i4XKStOz6LXSvnH5WEsqIcMBXNzkUTA+DKWXdA3HLz0t9h44obpiQ/
zoVGUb1Px/6q9bZf+SH5QsBSpb+13Q3zxNzIQO1ZF0Wf8bTkLq2GvaW6nitTtQVe
OvQ21C+qT5FfqLfL3/Je7Od/FbDumtjRWvSkHMLEGnM2IzbmDlPY/ylEzLMhrQnO
d0201V32D9oZY9bV94r54Iq5mtVNFO8OfcokPyoJs8bOpODOZIp4+c4poeqwJkGy
VF8m75IWuqMDPiBuuyHxevy2Cn7Gz8mgzqhnLx6oXnAX05XOx2c4UUMFQogi5aEp
KHnGRXzGBkIfZNYDum9J2rkl/633eyXiS/Zri5KVq+kflnWRZpfMAm4j9x9i21lS
pr7PlJXIfRL6xcgrAuK4WI0luiLKHY1qDXrmQ0N3yqUOQlyDlDeD5a40OLVT8tAr
2zHV2Gvn+rmp+XwzcWkmF5H4BJJDaKcMRl/spbuuia/4/cQQMqD659S+4FX0mgBI
EuyYSkGrqMU2aPGMVoXwssnCA3NLPM7eipzkPq2D8qkPMYfG18bHlJX3oQkuncik
DHeagXRD1Y9K1pHqgSU5wTaTvcfmxmm1LBNrplJwf8zyEMa9zgdZvw5QsbaSAWe+
lIEtuaH2asaEoHEdybnLlfdc6EU53X9qQoc+c+Z2An8V2GQow8uZYa267wCBJ4NO
k6n5lckD/uK5wYreMCOJfmfyXvocDjTEihxnbfOLyU7CJXWpvtuaXTPH+S+90xie
2+ZTRlF9H/+GDsxIiqi4XRxfMwpxmznGXImY+BnLaayos6DUz+64U/BeG1lcV3EC
AuMs+hxWiChWp74pHhqhvEwj10qLtrrpOpm84uHzqhyMTN0NWe/OqEFVukSgdXxL
udODcg5/G1tNPn7guMbXkisFxE0hmak0orTHpdV/R6PfRGajuJ8hJk1QRbWud+DC
Qb7TwRXLHqVqZidjvYr5SpfVmc7K2LYjzqP8qxuS+aobPnUTKbcCwu/0YVLE4VDw
7aO6EQscGWM59mx4cBD4M55U93SLObJOVfenK2bfiCY1UQqe3Xy9dIIwxw9Wk9Cy
oi1WKdq0B/glVeLJs6r4risdyGDs9sUF2eR4tOnoa2uEj9/BDims6b3jqZOhR+tg
DpK0115IgsFG8MZhzq6pEe+AVw6Nl58bZgpSmoaTDCn9VUDpXJo7o0ZwNUPe9pcu
/IWSdp98NME4DcPfj1akUvYkqlGIOym9hguAlkD2V1bu191glAajKWcnDfBM6kV3
kxTnrk26KewVZqgaY6X6WrW/pEV4PqoKVMxfv5qeLQBfbyS+Gc7GumUEnhjCqbQK
leyzcJh09i+L2ouDwjtBISMEj1A5LCEQeFPeKtG11ISPJHBK1OYEKkzQCbj5ebPf
OPe8aHatiDeguPH3pkDjtb9OFZWLU70T1kWFbqgiWt4nFQRN8GTRSxsPTY3IvvLY
doYfbQs9vwAu4QIMXZMGNLN8/GNTAOwtSedIg0ETWt+TVVW/GkdRoL72WSIjKfm9
9t/GkQrxJInch0MBGsQLXWMKULQfn9paUxpcMzmBo6/6vGw8YOAHXax620H4ZZd0
9PW/YvO1yTD5myrJB1kAGCRZzWnwlb3/yOv7D1ZqzQimSx9vMYj1vfK8611K8eyi
dP4C3UePsIyNouQnJweaiKNtmxIcEg496YJpd61bb4Zfa9QmWAqkf6Z7Kkth6cE1
F64ZOB+l5KWRvkYuveSB6XAY/CXBOJaLf/v6sJr8mqCcc5GPJ3q1Cmz+Puz3sSVA
cPiVxkZYG32pLJC/voDm8EyqI2P8+BSgljXpS+hvEX0eymIlZUcdvbiJBLG76IXj
FZeHP9/sKhQQKACzO1uZXzZzobiVzsAmykS2x9LwkpI+GZNKfid0MKDYFX2soLXf
TbvxHX1WAZLsAkGvFTpkUg8j4PE7y+zpBmLOx4MlGAPzF67PIRBYSh4QAnZ0QCX0
OZQOHp5vhGLrWDJVj0EezF3GTR+jgA9KcTg4+r3hn1ZaEA4Du5i1H0O/VRkxEu8N
p/j2cqRznkh28N2GYVQguIJV1yeywZBDPWns0VWjsOl35PsGKcr3A82/Z+EvkBa0
Xh4dp4XSfQoX1GeHcdKI6Qg7+3y+HXuJpzfiUeZk4HtnWNtBh+W5gnbrEwWXo14Y
ZhXjzAso6vXQq3sTSJLj7dbaEhSwEW4I2XSu/o8nYVEGRtEMXo+XrV1C1WGoHmYv
KXL0+nSCJXk0JXYODMZApq9betGsMiAkOTXjqjARKpElW4iPNgp/es8ron8yXYpm
a4IfWzvqC9GPNRmGRKQ4BKC2hWAZNGHsZCec5kQaj7VEXxMyIMcwPRQAMuRkqSbA
KyppkG9wgrz9e9NcohGxXihlMQ+SVq1V6rCtj65uOnvcDfME1xCKLSsOwbNfRrbQ
6i6k/bma/XkdT4u+zsmtt8dvP6nz/xYwZ6cWXsh7+XCDYKQEhrolKw2lu/7OKxzN
CQ0yx34pigHDijQ7wW60eCd+EdguulH6Br9vD4yRJYkBvEAAFcMQA6/PkimBCl03
vY3nG2BypnTB0zzJxRiF3PULJxnbfy6kc2nGmx3eQCuatxdXuyAnfMaoXc8nkC4o
LxfxQKtBrytOKoMbyfDJPrhpB0q2FFKWxBhqEIvwrpBfO+6nkb0eb1z5X1Vgl35Y
1Jjd3P3NtGhRL7wjDi0r1k4Px/E3FT20vYDy3Gs2UBlA+AhoucXdt2NcdRYIrHI6
Z7XgQKrHU34odK0OzB5rA1AayQw2MENc3Xif564DR3KmLIwI1OkTEb9QWChDbu4z
77eXNu1mWK170u/tC2TjSKIGEPoYWt0+UbwQB+wfz83aU8ocWiYLyUwStGlPBeEm
pqlBkvXqIlu6PHz7BeJ1jQdbPHg8R+hnJDudPpe7expZ9rk/lhc4a4Ltoeolc+dc
fjbTPiqF5qb/syxpuAZoDouuRbBuLjCp/QWFNEa+b2zbMKPXeNPv92kcDFsrB5h/
IkOIJ0LFvvigWS0FB87IU4RB7XFFODX8C9h6VPvbNGJlY2DOETpv4yIQjIAtrH69
xBEN7acHcfm9q2zv/Enr9fa/i+cSwcaJbvqOQCgHqJX6Hjv6vKDM0kFnUvoGtQ4z
/BHUjN1Cp2seQ3MLYaigaNUpLyuPgakJlj1uB22JVame5hqB4FTSMr06DLIzJPzD
91EdivUivxQ0B/JGfGk5ip2YJ/waP791LzuUVhe1aAOWV3nQzp+pHe5gOdQPum3M
HbjcwYodpa0jTEC5K8RXdVihFHbyFlwKr68VdM+5Mal39bXSXtx6uKpy1BYKd6yw
JFsexboX4OQ2yD/XHle/mO3G7LAp7wgdXx/pa02VThVnhZsxqqhms6sb2LWMxufY
75MXSZkpS+8SO3rbLNSE0x1kqfR8m0DgVS/3RdPy63Bs+QTqL/if5hKMDm2T41yr
BK3McrwraHB42E/JDxLmroJ6BRjNq8FLML4om2sDWkNK0vhR1tG3l1hEMIaFnfK2
40CSk9/BDZC5IWxSgaTNT1IOxIiXLo7VPAblUjg7aK2eEY5jbirlVi2teXRCrsZT
01KP3T3k19GGoR0srNFFRqeWHNBxuVo/P8OIufrFFqgAVtUCpRtXiFfOVXiI6ZbO
Ovo/NTI868XFHpNhE0/rixLXYemh8KuYri59pF0HU76NKzuzw+RpLJsHTLoqCnN3
xsgy7Lwr4sTwJFIidp0Qxp8TMESxoHMQVnLFSb5MFVElprJUhCX2MNcxMZNYP7yz
MvE8bm69Qq65ZiMZezC/uWPpL+A6rVD2dAsJ2ed/7kwkAb+ZMu7QkXsJLe3g4u5Y
0GcbG8949ZNtq0pcxI34IUtmD3EBRsIwXslogHbAFEqquSXL1E3h/klSKvphme+a
kcVz8RIsAAhOKncUQ6+Iedr965BinYtJNwMRVP6xm1ombe0/n2HrccZAIBWyz/jH
Qbkmo3sXBDYvlGoND6kk+MVGHgo7Kpp21ILzv6AWyTLTRe8nnLQfiGtDB7IJ3raG
zdFNYOCTD/mnJWZGeSegfVd9+BqaoKlEk3XspT6JfiypvFkekHKWFs+Z+TTvXv/q
JwIv6vKiW7JxxnYhqJzPeTj0NBFtCk9hcaN1uBL23q3PpxfmquBd7PfnoUyfW2tu
0u66+QQtYG3nZj9DVDa4FP3oYW3UH6sPe68oQ3mXwz9/5JVa7J1+swXTsSxV8JaI
wyb17haflQh8z8Uz+MTjLpeQRO1+qkPklIrT4ky2veayausgzma/Y5RjomAoznjr
sFZcBHejhhGqKhCRaaeNBvURWwt5r9gBunShFwCFtrf8BREJyrFZ1na/x2CkU0Ds
uLbdfgTdTO8vpOr4RxQKMznCXovs7wSO29fjHmBJZyZRdZ52yF5TekB/SooFvlIN
z2b13pRNosgOYtktmWvxrlMjQz3dKl8rRdPcteoGuts3CpZxUE3P8UQFFfowu68Z
sKpdrjPxbE8lpgc59IxoiidMvEli1tT9XGYWnf8js4NtDhVBWqF4uXDqyaIYnJhN
1hrnKm9U6YWkmC3ac6dmwL4CUwK56WrRUEhYMBbtlH0Fek2tv088JywJC7DnY8dY
ssLWyBo3NgruT8Xe6XSo1Jn3+4xweR1Epsb3T2ch0OVJrSiJhksvAJSqBiS7jXoY
F4r/tzPgtFt1J1bIoAJ54H/M61OrBie5WKUEuXuC6G6049YvnHS2Lva283a27yOz
y36N5/ye+bQtGVVhYyGaXACevYHEwke6GJSWkIJee20XRnh4jDquhnMxLaLOMocu
pgZOqL6QQX+MxllOZ8KRIZWkKyO/ijEhsaZcvaJxCxw9BDe7Ve9aIp6Rqf5sklIr
XGjBeAtKrUFmbEfYQKTKCGY3fab0cAZsxWuiXQnQZG2yZCfRIKOoaM63tn9SQLvD
xi863sWTt9qRZXGPl2t5Vh8i8hrauXVCGgUVUyS/cZ8A03L7I1jPpOJ9Wbcl7CBV
87tvpY23HMdmPebFV+Ta0jwv/I3uAXZhQAffLwGsi2xGbbEnq8PCe9cHp+tCSUz0
uwOmZax3Gh9njjxKuAXeNKhYu4gBnZcofvNxQYvR/npsBpDWXzInekpROgYcURBr
YaGaNqwK5DjkQjE4rZHYPbiaixk7OA+Ik5QjgwNg51+Sxx/HNsHBYmi9gELDIO1N
jbCdzI3Dejl0mB79acSD7bDTd+5KW5rIk1bUVG3cqYClF+0YDs1SuhD+aLR3y5db
L7PZuJBO/ext8HE51tiMLCZF2zRApMe/W55rrzotTrL33olxAH2Q37RUSA0pFwJ9
TGR9E4PDHit92L0ueiLuFbsW94RrCWnKSav0Y3W/r17TuQlKI0YSy9HRVsJqdIBW
KmcLoi8GkPxmTTzAjyJYpZW3ihcpbO6kNWyI618Erdyq1eP7ryfd4caJ1aW8r2FI
D1Wc8kEESKQtakS24bxwq4faokIT9aOAPKaozqOyqpN8ZKLCoNjRSW4qDMaVih8o
/e51dCNuHENbkfaj4Pl3wnIFsA+UQanP5vcHB3dRF1RAq67ZCkgIaE9XpCO04gZH
w36eSq8/nF3nCH17h8khFsEUqQ4tDVfdzqH3gGfe3xqKb6yxSUW5pdCAIXgXjDGO
CFUb2kKve7mBIL9PiP2hBS2dMq+8kMYyJnOqvRebZf3vFPUybiFZrFC4ZSieug3Q
Kan2NJl0RMPmIkDGKXZbk5KYiv15gRvCElJjcgxvIr96/EwVF/ffwY/Gtz0dQ2IE
xUX/+j23ua5CJ9GMJ24n2gzxjpkl83EPQH8qnAiLFDU8+nm5uBba7emfPwsRkR08
yPPcuqqBzVxfTcGTNPafnVdi9kbFNX+Wa9cBGBnN+wHSb6AKfHNbLQ5FAKXI4FAD
JkGw27nnLwoq6HnW2u8SczbpPlJ9N4f1RaXAsnOcrbA+Dk/zfbm0WwtdRFDz5m9u
bBHfeSGEI37ipapTE7947rRorITfq13a2BET6Ix+EXwpJ5e9oqHNkGozZfn3672M
z2UMhBvtySMWQDcfEVLrUiSu810E24uoyewQHGdV7taS2qWcWlmTWNUIN6hyFZBg
y280BQZ0voYuenlIb8RTqkbRwkg/tRzefucPM/4zH70psa09OqV+JOeiV7w8/wZA
in9GucAGwDFuetHsgMo1XNHFHqqW2A53rKr9mzt4Zc6gQ3ifZLgbfIeLAWEVt+cR
KPMkIBFo2hQXWYcFpUeiSUp042x6D1IsoC6g8yrT1k/Jxo3bpgM/GEv9ij9aDvp7
qrfmIzqUnlj8ohrIMrhfvEBYqD1uw7tG7DM2cI/d7t7OkwCBGhgjDOxcTnSOjQJ8
SXvjktdfSqieAPYmzZcGBtW04dNsS9k3+Nmm9YrQkQMVbja1+K/ZqdnivUR9Te4g
4mlW1Z4OysqIZSIyy8mh11RrE6Z2y1sE6xliHyqGCK2wy0U7Or71pzfh5IgRYDrz
tzynL2PGIfDJd7zeNELi+HPcD8fOEVaBRMUFY6cWcg+D2PjAiiSdOGYNIcBOo9Zy
zrkBKbKpsqYTUjaLrJEAoLLc2U9lSuDfVvKn03sWmnCyGbzhJ4neYkDQ1j/9c/fn
sWTuB/NOvx0SPlkEHeIusuIl2vkM+k4Wil+qcWCVyWcTA4KQ4rWJbXxGuGmqRHC+
bJEAEk16M8J/qvzj2odA+4U65hI+rhDMFnfNAGnXwka4Jrz0YcpGQxn5f0/LDBoG
9FYLQ/q4HGW3oZfE2gakrksUauyKFbNwbZACCvlxxMsbdq1yLC/w7qgVag36lG+S
HKCyayhV7kSGIzBHlLsmE5wIU8mYSBgvFjKJCh7jn6K+BD0SvgW4jqGeRdrdUpGh
SmM2MvqEC9Z7Qoq9Km2PtgSf2Vf0R/a5dzC17C6xbHil58AtiN7G/m3wr4dY3bMQ
HjCBjnVxOMdjKZOhPfbP8Ws8iKr+tYV+LgH5NA1JHlJjoLN5BFMrxm4dS9tt2gv7
pvZERLOfaarx4ZKrEMV5JtOgjRDBc4vaE3odlJp8UfjszYJaNKxhx6llH5LYuo7q
r+mo4tXQDJGmFIbUbF9hvCQP9Q+iJTuuSYzx5+s7xTPelgdwW2JiU7815/fpAQrF
ORKwhk1plIeuz02FpnJmbxgU02k1ntjiS80RhQdEHySvdeqNT3yvbnSuz6eCR5EC
LTRTLY8VCcIklb7PfaP4vTypgDSDMAZFVTkTr0kBOMXSVkAbME5UjqZxOH9/YpOs
Adqyy0NZ+Y/HS+CgL5jDDcZXOvHI/IlHqwwKlFmps1XcyBwAiWBuIK6GAHXyMcFy
x5j6rLc14RwefYOuxihmy3XcOhje2AVQNm7V7YhaTB/mFna2xSIYFgQixWnPQzlx
927jqH9gkeH/msmEwTDH4m6Vp0MVevpn4zs+WgjWqnZ0XTXqdyxR6ymVubMuhK6X
x5a8mStp7T3KH8GWtL9En5ZslfsSqgx0Hldln+RMKBpclLGcx9PeO0iIPahVRAW3
0YAy//TKifgZVPhcJDyOPLiz8yIaVys1IvUyrOh7jRuKwSbuyV2hULuAsWw2dTP7
Jsuv3iDOm7GNa8by+5ocuHG0ezaKXyKGCXPqNlkDu507gU3cVrN/BkCQ3m5d1F98
b3brnd2jTp+rLp9mvij3KRLsKQccRGrp2aZacnN2TLZvMSpP1LIEW6u1dXrWvbko
5A/PaXzJWQ7jShk0c58is0WsMZe9oFRdIR1PusPSwDXRu46NM8mxHKyrzDu+uJJ3
tuJFTb+EJyWGkZ5uqFH3WGHMMC1Qf/IlOvALayiFjziX+7mf4FkumsHX+qWNHxFY
qAqI2TqvG9jF1hRZ4N3zQ4btcKAQmEijZ92C7B2OnJ2vRtLBw/W+Y6ygu0q3+sM1
PtmUA/NR1sUwT0tvozL/0ayaqZIxNIbXCSFNwU4MrESrzNp0dNeRkbRzfPzpll3u
/WrQ9Rbrd+TGb60WsIwQv0suyRy61X7/0ZY7J+HQ7/u35ycbnCUzRskHt03Sz/0+
sJw36ArYX76Dp6oIj7XJZ3TXnX6h8/hbxv/nd2u1hqZodXurfk4SXYjhAQ2hd350
YKZhNn+29OMdNxCA0/ARru0k3MZez++Qd4z82tZXLR4pWFQCsCGu5nnUtWbQUC06
KQkeMNep87KvtnvSBVQP0gvUTIBdEAQ+oxoa3ozqVyfl4ye9+SYucqd0bh3XEVu4
RBlaXLrGk88NPZXZj/2KryWYTHmJo/9b7E4SQfZAt+AtbbzF/XkCVSD9aRArG4Qq
eSX5fmmerC1AkRGgQADBLpB/8W7C2Gqg5VIe+hLLByag1v4VLhXcYUwKzPmAsAMk
xJW/fFD/A5oDVXQ5YguiEJ0YO4j/DwDhcV8KXKWVyBXh/JEJjbBlgdw5g3escvHP
AJLDPhs5V07+0UeQ/Dz7qPP6v9w83yoTiaDsFJNN30IkCR2YvQ6n/DD3BXD/Y+WM
MALpaXGy4V9/sv5ulA4x+6crzDcZhklBKxEWd810i705eeElybWvsg2brll5lixA
/l0Ur/lgHVwuM1t8n4i/k1piJIFinzYZQ65YoN4A/Q9OzmWfWA2siMFQHQpxHSE6
cCxEKejGToKfpy+vNJlNsCzOiPNluag96EJV4Iq4gOOGZfkozeE7aElrOkLMSILT
gWnfMKr5hmSm4Qb85X8Oe9r8pYZRnSyVQaVwuuU4pcAVdTlx4mZeYAHE3cJX6nBN
EgN0IU2iQ5CxBQlBg9y1ErtDUzGRkjnQV2tmYnVwv6YtB345Nrim+t9/26opCRZO
nGOPxvB697Cz2tz8rjVniCI2c7qbc0LyEPExbtllGgf29Rinpw/UeeMW1nfufvuz
lcXLbWMtf1FyPZXR0JT4hYxW9dci6pB3UdJUI7HGixSRd2e/SxlDHgudrleVFIE4
mI2eHKPiQZ5QIsJkY3skKJrJJdjjqwPZVS81HnO1I3U5D0CE1I3BTj65U+NcTPlu
te5q8d7pv8vTKF9GYZRilRYOSrnJPfseDSmZQcKHd04i4cvCwVi3SUX4P0FMCcOA
jn4Tl89xvtbP5Topy1R+Wf4h0tjOSD8HCPHkNsRpqLbNUhKzAY/NgcB2IMj+i/8a
nI4ygYRKkDV++BtvkgLI/DN9FQV4wFrTQhtLXrx6viLtCXWZQpPPBuYDW9lwRubh
VbaAxjPN94eEUEHQbpuW3eTKF/qM2jrcsYCZC2RFtP7bqQq2XhgEEWkyurt9w+bN
2NWELfrnjB8AO0Ey7+0FJYfUlL7jUfKRoVZejEQw3bRTEd1wTSUHVLaG8Eqb2FaK
JZ8/7PMF0awN7kjJXbURJAXqz5VsWvOa7ZQVWvPUjJ3dEUlXJboxf8Fpk3qhfGg0
1SJrnLakjeyr9JuMGxZkr7PbMHFpTf23QIFCZjDrWAamvFDku4F11qlbdCkEr0kP
xnQlqpLQDgAuWESCAwmSgeN9l9UzQs27RQU8MVzCY2an/mLkQpGiyQQBy9Sd5pq8
iadEw6MzyjQv+nEmpmlLKW2X7Uoztutrb2BM9ppdphc7vuZf/zjAWe1gLrYT4vSn
baY5wnPf+M9iS7hcNP2YRSBjGk+lTIAVF4mQqL6NtpOS6L/ls0/t2fa2fw67tF0l
+x6VJ0IkV4xnmKJ7TH9UX3Etomb1ICp1mLbqxy/b6rhGJ7g13wblb4yUUWQt4JX0
6cRpKbms5rRP5gFh/pcW6EAx48W2f3ID44OZW93QdjweJn4H1gvHCzWCLZ8i4cMu
6r4Mi/UMHNhz4FyZKqcWo86B6f+l0tSsCngUvrBORi15cC4fSaksna+P62GhWqr9
Ab81rJATzmO3+SFmGAdakpmlDG04+lzoSvQrn1hOIMUk6jbEhnnssFkGZXipLSsS
GiBaAN2I78oM8YtMSio7McsG1rh1A97n1GdsXHFbBZ0rErPrrKmWWgmBA0FQ9P/y
nr8ZJV1CfHNlv/mHkqUh8Wr6VmQd3//HJEWk5tLlx182QN0GB9Q6FGvqip08yrjq
ZF+OAJG10XrVHgxch+wXl/XY6ZXs8XwSvuY45kjkhemj2IMWOlGQ70tM9U8xrcTQ
2TfjICrFi1wbVQw/0KNk+jrslmRRt8/ag7KqjprejYdCezXeAN8I23byqzUEd9FO
uu83xB0VYQZMUa6ELQNpAuHf3j9iIPiUADbT0jX3bkce/7GZg2CvsiMySwCb5J3m
E68b3sAWGIB4ImSfEeFjYLF+lYvoIR241DrsAUSTV/lRNYJAN+QJK/1+9MOe5Moe
Gay60kSIzVoUinPI9aBJyO0ZR4aLUEAxFlqzBftbm3YJUF4+b+aym4mCeKVtUy3+
Lhi2xqMcgamG8p7uSWCI88Jd5w9Ut4QwLqUvHevcxn6Gac0AQVUyBiqtT4kiVyrZ
aH1IcuSQ9IGA4Yb0qi0PwKDDgxD8I9KLdAdB82u29nQMDWlZDMJlWsJWNjGgmxVo
4Z/UIOgxUFL0xmgyATl5IV9yYumUiOOLvfKM+ErORBrJNzGfXctLX5XcnLh31s7e
+iNruyYA8ovsBYCzpCnaomgyHBWuqDi3BMDd3mqdxuA3yS5Urv8zOdP/yPJ1WGs3
e71PPQjzSv5w0jDYN9ptshOSTJSrc765qmwVxDuKdrLAii4xdjkFc10+mcvckfNa
JKvMy/ahY9ngtSyH+5tpCWMcGSRgqVksskfy+m5OKzQjedV9jSdZTaT29gAC+f3m
WMibqt1fIGpwNmWeVkpPP/AXkw5KoKkv1Tybe4Kw7X/yDMXolT4cYCCJXZYU0Tnm
9w+uR9FtoeozjE0V20x9n/CqBtZ7obQSC/+LN4DlTQb0uFImdVBMVIaHNp1jpQNa
5MuVCWx0JBlmh8Y0g54YFoX7DDbUYNJW08ihibWQ9RlP/Q1TC3FIHH1ubpz2LCmY
JWi7VRef4yVkbWYzoY+PeEdO4OJAghWkbHh99RZ2ZPDJkrwcQRn2227QjunZ6MRJ
qHqu63+YY3cxZXpRrOiaPSfFasfEjDJSg/nDFK71fdFLCa/RExy8Ie75TZWtiA9W
8lEREjP4KL+lwc/VHkdRL58dqVrXXy5+m80kT+F/3II/NjS4wb2oupfcn68S6Pxt
JsH+wIg6c5KuJzvt7m8GV7gPCZtwUJDnMzskk0GLeP7FOulNYUCfzsnRUBVTS3/B
2R6SY6zkyx4Xfnca9ZhG3jEvRlhmtDwe++oTCCYKnatUs6uPQW/k9i2/OoQ0qQZT
HgmUOkPfkywnVRjk38hiI2uBe7l8fH56pBmyApZda7f5nvlS3K95G2ipbC4yTW+I
fBy/BGA0riQCZczGVVH/M21Vky6zyw+mWrTJlj1pEjvLVrqnP+kuM9rvz/3j1P39
dQfIjbL9NMqcMzdqWd7D9agW9bEuKK9gE5ZXVBSXsTATGA+JU2Pp9TYpGB03aOHs
Wu6PFwvL3OY1zjjl7IL7vZ6bF3Z4V6Vz3ObugKFFvCkC0+q/ckk5P7rmFuXzCpcn
WB6IY40V31A4TZ9sJjDlW8fwMisRTOKYo7b5tUj93tM+02/EBpj+ysMJmzGB99Xd
e5PONjywoocCKvlwOp95xQdDjieHr402w3z7Dah1RhCiuZ9d21h4tQQHu1PG6ljp
FYeMzh98KK15b64yMkTViAD7S2HgZp1Ma3BHNlaLPuFws3HHQzKpn9bUthNqLoaW
bV9pKdcZ+j6DhC/ioWThwLsGzmBr7ofU4tljybtHzZjfqb5VfCjExh1eOteB8HeY
koyvCeKtCAyl3rGMuWXb98yqgCg68bMiZ0CBfyhWvBAJdclLquXnIpvahn2XbOA/
kF06Yaf038mYTfU/6YFiLf+khc+7oEh5Nm5v+mKooInvAQF1vD3vJ8xIxbo8R/Ss
bM9OvyqOIpppCPcsWMpQm0cfL7kfIHf24B+0BYxmqIlSdpwOsj/qfjIIifPqn6r7
2ynOmWBKrZxGqO4jduYwN8qRv155Hzrb28cCYR+q6okjvElIJUWq2oqUGZLCFtTP
HCFKSAFMJOqkgLiOBbp9NqzOC5XBveZ13zgENoOTB77X/SBJDP5pGYfaoqVyIE2a
G7CQzkp70htE/Uof9nE2bJvGquIOZ2UfnIR6yWc6zRRsjrOu9jjOEHF5LNoakRNg
2Dflxc0PxgikpT8i0o5Q0s0zwKe3X6VMskiEvu9hqnY6HOmqiztG3UqvOBunRnXy
Y52nHzWH3Xy77VoBqIhazaTHIWdXibK7jXTLSpWxE8VfPCWgrkVmYXb60J0LKJ2X
tNAg+e0Cv2LlGpOtTLIlaKg1YGnZAQ/pC4q/kBmj5+1pQS4uc2QwJkmzqzhGOAev
iVrUx/at4JlTvdL6Kmbx8D5qP/W58EVgl9OcVNeeO6iB1FAvtF56/WNaXRALvWJW
aqrzGwkngpL5aGAUZslJIqhyiDOuMGCE+q4ECraqOVQ3IkxChgQUUm3mZu4ODGHO
Z1yIvnRZOdDltF7UFmJoxK+Pkc43zlFodvSRVDJcnQmkik9UAkdDUHBgdZLKRQbC
G42wtrHtx/NI3XoswhKJ/7N1Vbmy6zRz+tCkASCj7K3WrsATbPz5qPCAb0d0fi1a
I82+z9TcnwJ22P38WzEcolr7Pt4hSHc0nqFnGK6sdNuY95xuSholIq5sqMGYppoN
HpP0OWMy4+4ghBM71jZvU6Dhj6LnJrT/rurl72V4IaSuSgqk3YcDum6pwvg3Z97D
m9fIO5sCcd1uwGhDkOSesC+nvjYBuL9SN0OLOxnFky6Z11eZeagB/iB253gi2xMz
Flh3cv/+ayetWgph9eJ9w8ia2JUHsCNDwtEMC4GsMOS5rPw97sbOpIYpecKl7HrM
ANyry1hlCdr7k+C9xYlM8cLJdujEWc1OjN+yCRjM17w/yLWuqVOZAmSRaFFuBBnn
R+VntNC1X9aa/zqNIOY/ltn6cEIA8DiV3+1Td/S1ncXQw/syj5PM03Ids125MmDm
AdTJYDncEgywVA/SqbPdeGTv92kklsPNaYclk6ssRpZjna3G3yu4c6jhYjRvAQvo
ol0PuZjjRP9PYyHwMJibLfo3U6WEyjC1SBiHxkgXqBuf2SogxMA7VcQ+rAhOtrMG
2rXvuLqFu07ZFSG8ClFmG9UjnwMUqQy6sdY5tAd8DREFuvqJoZxD+sDiigYy56PG
VyAUkLkUVnGWpXoz+M2z3xuFGZ4Fu1/jg4xbOaD1RERK4UpwfNqRVf1gxqkw6xS3
HOj55XQKa0m5g3c2AHPVwkgTk3dnS9wRBX6zm2IGpmXOL8Kua6Pm/bRavoH/5JKm
LrlT1nBESdk1CP+e8Z65adX/Y7o6CpWIEUXm2CTKums5nV5OyzoejG7A3RDUtver
NdsmVOIiFaym0lPi1fmQYQJDVhIxBLjA+JJJ7Io43sMVbhYxr4zdJcKY8q5Tx3Gl
s/h7La5yWgbPJoV6JZocgYuMF2ZGBb13sJOMY1UrtEleZ6s7lQp/DxVGJICQCVnM
hGcF+3k+3TS3NMDBAkeOJ2LzMSBkBOrJdk5Hn7wRkfhQAIZVMEQJ65s2oAFaFqVw
TSwihDIpIaYs6hrmtIAbMg12it4aj9nAoyhEIfBWPq9JCxtqQZrTuUjjRdCGb8xr
dyGn75ntSgDBcSVv0HCDWt374AG9MWHkkx/oxl+Eu7LTtfOwYNdgRtd1teP79jDa
z+4qVpzTr+XlELb7s2GoO2M7DO0ZBlOIBZahSuwtvyLHZdS/o/zbjRAMhFm4t8lM
uZ/NfUk8+ZNd7DXqEdUDRZxHHY8eDeBPhl4yqsUfKzB0EA6+1YZF9Je47pkVQ5Bb
LArTEQT1uLxteMNxpJfBVdYC+M46z5dGTYhTxyCCBMfSuq4DZUQWTUOVblR0ytUJ
LV9wzMliyCnZWsfGA4ekJvkdItmT2V7cOHerc3SaIl+FTtZzs0EysXhaFfKGSzha
4o2ycI/s4ccQa1uMuS7JpsJF0O0gZ9RDbit48BwqPxeBbKNuE18SI9HqCPwl6UV8
UCbNt7WyMKcWo3K6wJdrq20AsufUjrcrF3I7eYQOvqgf/DZLYF7yA3hTHT2BL0mk
P/aPY4MZpSIrgHaZFSbkW7R+GNIsRoEy5HJduLPMAO+k8mFBTIz7eLfMUA0vuFbm
vn/fIXpOXc3SiVixzjunI/a6+8PZV8iD/rslQj2fUqhlMrlI2RHsNTgaJDr07czh
PxJcP1glV7NHMlb81gft9oV35GCezc0eGO/dmKpdKuG0c/jzJEQ2EIUmSLDVy9WL
q4yCnZiy6dWl/RBBrQ6Lf0M7SUJ6e8zRzrMlXTf4N6Vjka8iOF3wAIuecrJZsfM0
sPASpwpeekYlSgrzR+FpOHlgkVA/5tQSegBbxniD2Z5oBTDn0VE8+0mnNmzg+0ED
SJ+WM9aU0TCOW0aZLe2iMNnf2NxEEWqB3ofT98qObLP8vvOaMfXzATka6sRLxJdQ
OnEWEbjvZioSrTbsGxJ0rGgBess0LnKgQfFOMqyvcrTl4OldmDLNpcHWWa+CNJHQ
zmp/ufxLP2fKwwyPIqxZ7GiB3isDz/VtXUiXOUsNHzMosBGM/ylXc3F84Du1caOg
FJc7eIZESMi8LS6gPm0QLXVPsO00fLjuFF4WRTi7CtmeG8UF43GDJnmHMD7HETtH
6dPuDKxs6+QXXeO8IVfijRCct+R9UeuIivkE1h9xnkcjuB3I62JFUb42zler5jC3
RLbFnwpszxvL42IEd2SxyaY6b+LVEDX4rPItKCkqeiJtRAo+vzb2o674G+qV/3Vf
7daTjniDBJSGrzFq5JsLwYgM6pVyQjoOl7Yz5AoRvI8sDhC8G6KOIAthVMY1aqld
n8it0TVLO4f8hkfJeFn6e1S3yFewJqAgGjblHCeMT1zJCD0KKdz2jpNvBsg3KDmc
jxTMv+IoR6hM27MHPVB/O9TV3bpXEvtLisjUpbPAbHmcXIi3+rJaMitj7AeMMOVR
2rI3AlQyeGwd40xujOB5bB1AgaGY3ySE07ijwB/c1Z2droO6767CU5jKftrDFqr3
Zu+pE+yNRm5Hvji2yhKIPg3BRLsdKMB61HZVdMcOQtfK6JAkEzIDnk/D0AbiooUN
UU1rUCD3ja0NVL+jj8XRaeGO5EFw1gcEfsfVn81vwBhs47/pOLlP5fC+HCmfuu9u
zXn7A09yYAFniGoF5Q5ad7CuZCzZbxcxoAWtgdoaRv+l6GpcADTHdCMRtO9YgzTE
4O1QJuqdO59Tk45vqFXbqDPwDpQ0zDeVMUxQYpytfFafdbNAUxiJKCi/2KvH9p5F
2jjAgpum8iCFfo+lWsE1jtlT6fjoTx6G4SfObjyw1zsqmSIcEIYuV5XxOxNcqd3K
0YxOiE+UVkkUVBQkRq7XpYDqEfpFkBBo+b86kxH97RTr2vfPKJUbyFFxxM4SrJM0
CQNszLHceD+yIm7eP37h9X1IIf5TPgEA2ROuxRotUZmCwYNfeHay385R1vd39QCt
KOJiBt4H092Pq6LaLZuY5rlYmyEE6yDGQ/2BMELWHQYIvraIvl8cZQ6Fi4rtPN0S
kavxMeGSksy3S6vT8fEJB5D8u1n7/tp+pzj0S6V2d3ZkyeDQMLj8U27+jM1b3CDo
A2Ry0OO7S8KrAPSS6gTzfXgcEn/JiEsXHm6LJRCtnjMYUFL6Dza5PC+KW7pyu5ZU
F/s27BPMPtrWWRFzdMIEVMJogrR7WSXbTmd1NVvuzE8o09g7HiHwbiqAfIIM2+Cy
EHmj+VN74dedWfGZyjaqYq7JbvdAMIuuVerKkYGy5BKRd911OYTkU0d6LwIPejWQ
Gj4b6WjqB2iHxXA8kXL4KLLlulpNsqPIXH8HKuIrfl6xRz48+1FhsrTibnimhSW3
qxdg7cQfKbQ8DNww4D8ijub6xlijBuXMYUoRIhNoAkjf5Vd3cijRN6ncdcKpz3oV
lrFaEE4bxyfNSHXhGY6dj5LwtswBISGLUldMzM9Ul3bG10JmK8zfZf8zSO0YimCd
pQes9ySicviwfXM+fAKMeBAYYmN7DETJT+KAyFhDawv9giqJvFHnN+Cs/SUIyVfv
CB5LqE8a/IbCZuQJ3Hi8bybqbliKaDCWO3f2gPWkPuio/ZjG1rmU+h2xc2mUdc6Z
DMjpYJfJOQ3n+gZ1SfvUCqCg31T0J7yDp1k57mzNpvkoNz+AYfDlqEULqhQCLNXW
2l5+oy8dOMO+h5HfQAnXZ8enVN0mteCBZRoCv7/pcnP9regypzzUxAlBIIGWR90o
VaBHOjUsGkc2N5s8pn+31dt8IvT6fxUoorF1yZFX4pxS/gkEn3zukqBzQq6xusVG
iW4RQGzLF8uLxb0hSI+bNAeV9VABGdZbUqXN6uZ+MrF8niefpezk0fj70iQEf9vl
k9YO/tcPoIRRfSRhPC/+1uV4fwcgDHNYVmSX9mdm1e4EjH7skT+LFe17VcBcfBIA
HwLvIOTVOLFVh3PUJilx4A2Arzgbx7Paz5PLRLOg56nNDxKehl2qgO/BecJTy+od
keD+LujJIPn3pvB2dbxxOVEuCGxrfmQQA/rH0LKIk0zM0ne1xrqLJ8m7yOlVv+jy
+r/vM3zqwaD7r/JVUeZfE5mFEjwxxtlnryoMk8s7vC0unFLJ/uej+pd7t1I1PqmN
4OeOIwVAHD8nueb82xHS/+uInQ4ny+1Kq9s9xMCLxdBiLYPxV9sv2jI759J6igBm
OqWeqWOKGed0BDG9aDzABAAWPsMcWJi3F4wtaoYkPWQpxZ8Q+4lsCsZ6rPRPOLpG
Rd+mJwPLz+eLE1zSqUBicKoMjCR1LeSceoL8+xZVix74DWWAe0Yu3kuffoDGGDkb
l+7zpatdQPNfWRRXNRy8+0/Cq8DIAPsJEmvyRfxOySF7AH8TX94bRLXpJeT2fYhj
m1xKp050L/POBDERk13MJ1QQpgt+WebdQn4yQyeem5iZShqQFkRKco9D5mIJcgpP
R1j2JXSDxWOLnsGt2O3itzcS1f1/uE66XvPpFgkZZCV4VlBOF0hYtRwtKJKh4Szo
lOSfd2RQOrYiAv35jqadwE/GTaPxDYSJ3wlr/nrd+ozH4aOqdBPqVTWk28pMbLiX
Za9arLxc09Pc1px/cFilKFOzj2qNlyU/F3FblJDHPPZZcp70A2vl166H0fCl/dRU
MxJ8bDlcGY8i9NwJeKxH9S33TpjveQqM5NkLwUIrWZLkkXKVEWPf3BT3ZJvk9rjL
2bym8QCzhMHlTctgeQLD9odwzYAuV//HyYkIYeXDxhXcsjZmzxE1WA50v3SRFaJm
AZawChIlFnuMyaZ9Hg7+jPAZBJymYP9EMFwj1guvIFFaGYKZ7zHz0fgK6n4mj1mL
8HRZ92BLFEHysKGY1Xge1WFavQ5D+9MNgqXE3BWt0kTw/LSkoBM8h7smrl8R6qYi
UP2+vi0yheShc9VhamjFymFkBmX9jCpzbGLqvxVO1EfBUOd9BPYvbA5LTNrgflgW
0GgV0PXdQSaCdprUf/9G4foRdBvYEsC6AmynIRrsMneMOdWDvZjnMXwVGSPCnDwK
EAvb30YalgMMAlV6Wn0mS/gPISgMHx59wdUvDoCKc9AGwAznjDMkgGU37yE3Du2b
sMzc0CoNbeW/YkjjUw5t/38n09meSraJmS8dSqJqWqPltftKOi3Ag9ooqdjRBT1u
+VCbcb5/Fc7Kc4jJ6ux8aevKciL3nb2xohIScQbYXYXecl7gh66yNEimwCREhb2z
9bZSR+g0gwL5fveHx9/kFADZygsD4bsbpdhXjosQQrx+VG0J1puz4CAgrKVjsMv+
efJ8hAUSZold/BF25wnLndgvTFXE6Jv3pzHNZIz4bHnDMNiJ8eTU7fiCiKSeilqx
7VkzjXhPUU1plIouDcllVvu/2PH50BZkP5CGqiYreJtnPF2tkjU/1DzOMPeU0yAR
X8V4zTpkD/ykmRsFwEB5OFmugz81JvUcr4t2zrrrBvCoUXXF5ueG/FminwffejSU
4KXP7xTs3cr3zzV7JI2tAxTrUX2S9OwxzvpvIBptBeiWcFrt63WOUUitvI0mOr3b
88KnkbDFSkOMfL/uMT6BRtfn9+vIW8Knlq88OitcwjsqNzWLsRdCP6oK2FMzpjq6
b/rCAO18TktgfeZKqZnbi+05qlyo1Jp2/oCW/H9f9hHUQwOg7fvmS4EaV9291g8b
Qye5VGAfYJMC0Noyk4muR58TfQsRUU72e21H9xFFA6jRjyxcxwhGWvSVvxnthGe1
AyPGY5ESFjK/cFFs/Enuwp5+WrGccCsLjOvArWAiKZsxfv0chF/MiHt6U2nkVlxC
SPW/PF3xEDyITY2nKXW4ozRSP2GzHhCeZSPXJ1zEcPfk6q5GDfvzf+lS7UXsefl/
4TdpTdoyhO8dh3G/zSnObmSAtpjqGNXBr5FqTnRSF4I///ObFTZb8pYr2T/UF5zW
coSS9qC/PKyzQDwRrNEBt2PbIGnj7xFZQeuG03pVcoZYlzGHxIye14ugFErQEN8g
YNrvaXQjC/1cgGtncpAocDgcOA0FGaqojLlxQMvV/oN+WqNERRZYQ1kV9Rs/eXDD
N+ZDqY7Da7veLDDEr4InRNE1nZDK/wsc/qU4KAOQGZkC9HVzms+m49mK+IpEkHWR
aqYeNt/gtLsdMMApY50OILMFqlhKq6N7ZoaZ44OArzyQVdwEsxDU7uvazkqJCuI4
mUFFTqLlkXcEFLeYP3Cb8wJIIqvt/A4f1Jz7ezpDEGgstuCWIPsy3iORtScUo/2M
OUYHIP8W5oiz4yZo3egQq5zJxR1AfoelodtC3trKPe9RwSEaNZNanD5JzBI8cobs
zbOz/EiRwSLp0Ab4YK922/pNtYlLT4OZMCU2PE2eVhzPvyVD0ynjcPaII2aIxbpL
hghaSHR2eWOh9LceciukwUhlruwDSmjTPdvcioGD9s7Foj5Pb+Hu+5tnI93eA6KO
a6Y3NRmD8kJ7ekEe9Gat5R5Z/Tslmo8ON8t7bSL313wS72ppPaiHd7xvTn7n8FIR
IranFxWeiDRbKb/AWAf7B4Ous/TmNJA+iq8UKblGf904jGFodkHfJ64XtpJYO5bk
AztAI7Hk8iDU9fSPntshVG1mt+CopvVc9FHFJUpRme74wLQdRFGIOrZHON/eF3gg
r0Jk3i8ud5R79aCPSJJxTL+MvPbMHoD9fDugAeRoJuYIIU7PEbcEWCxgvHZVwY2A
qDjk+Mc04P0pHvieE3b7SbR4t1lsr0W1rzVTMNb3gcRf8vzDO3wEboa6MSrzEbWV
UrzuyGldILMM/UOUlYCUbA4Kqu17EIeiRxawFM+5susw+jxNBqEcTM9YKCVaXny/
3iFS2vG72wjV77oU4iKuKRNOK9GY+h29ov9d3klv1gCzQ9dPKFeUA8iZfn7Pllns
HycxE03Q66i00VYeU0iich5gDHq0z9IcyZpf/1mT9LPY9NvMXFVD5XaLKHUN0ifv
nX0N6p9eMC9VTV9O6Nv1NdTnXVdW21sRey8YmvovXwSuvv7qn7ie8YVgWxCi7feT
X6j0UkoeiGFtHoMRYm3pOdLSJAzXiYEab8FgIBvOZPkFw8/6hei4zIJ9thHwN89T
R9d3RSRyjPX890WhEfXcMVcVHxOewIPDjjlbIKoo0kXnPJ2SudrzNQuBV0lGQoh6
SMTCDsObeSKCnbvm9ReLBV9Oxf9UhacSChB/8d5veWrB0G5j9wvwppevVaaoOvdN
NL0RWFDlomqFDmYXNdnQYu6apCkOSs5x57lkItjnyHJfEH9QXyYZJGFLTW05sihO
Z17nxnL1zJs+x5QWFHnkd+9dFc996N2NEy4Ie4u/RMSBMmoG4Ga1VGalr/UTVVZX
+g65rXUR7tubXk2l5XnKT7fd9M7emFTAqyrK/NQLzeeEnvz+mt5h2wpTcoFtd/Rf
7+Kd5AHS0MXoY/EHrIXSP3AMOXJtWXo8TVNXXYrImNC/igPw9w84uZnwQgnMR6QV
dEew6T8Nh137qkcwT8AzHPiQ7vbIHG9I4uiWtBrlmzEqHtK/MeG3RkBKDNvzmYkW
PYyWTYoegawpRtwxLYqacT3l6m3AhLEkV6zFlTVXRF7jwu70GGCgIsbuODzbVFlE
Mw/2Hc95rLabNbkYSw7qFR3ud1gbVa9p6aqtITHb62Jbfqi8kySVRgjBgsgIiEK9
V5Q3UVihRNtiLni3D8cYFtRQkX8qtx6yqxjyJJCzOyE9B934BwpMIhPv70Mk6HBI
MB+jXaH7N3j3EMmSt+cLIHBkdNIh+yD11AfSsv1/pV+lpZ2qk0D/5aw5s5oLh2qx
G+Oq5ETiO8k2+mZUMixx5I5aznIxCGquR2F/+bGSlxsLM240sSvT6MLGq4ywaKm8
Pi1UaJxA1eIUs6b2APmhZq3Ac0S8m4IEPDrg3pSqJlnUZoRhRTwYxBo9JVgSd8Iy
6GjqK0lbU6fwWaX0SlrfhU0WbYvb+br8GEuFe0pcQk/SvH9R4yaEYa4aZvX92MSJ
j8HKpqhpcqh2rcS5H86pUF036XIe3otQseC8A6GYvrLZi3jm58NMJMF4xCifrgor
BUZ2vhwYQjiGxH41VXK8kG43Wqz4y0+S8oaaFSbYRMtXzRpT1hYoi4afGl9thcaC
gTkCpYkO35DrrrtBFKgrb+oVuiUbF6JTIeRkeNx4mguwv/bb2X04rqu6myG6njjh
evWFxHHfNVjYCLzAGpmlW0EzxTImm4n5ebd7lCzCVsAFkQ7livOYCJKsHfJz9ChJ
bN2TaWpKjhiVj9nBj9Cj1XlT1bG5fwjgL7bHBYKz8GG0+lmpjeykhZBaW9L0vJY5
SyyF5Qoaw7DPjqHogCMejUuNF6+9SmsQ7uvorfKXygrgqXg2LvacAdbws3LiK7uH
PgzjZoLpfGZe19+e3nUUOa6eATM06rT5AAwR9/eLB7eUNFAQJpySUsP61OXre6hI
lp1n9l2ZUDfCFP+q27aOHo0vVpmrbM7WQNgR4KWM6mDyRv7DOE3nyi7kbL3rLEIw
GnSdT5vZQ3BkAGocOyDW57NFJwlGAPE2mG8J+YWQ/6RCSyALSZtXrp1z/6+F59+T
qHUAqT/iL8jw1vJkjdbd5VN/iqi3Q1spkfyBIpYItL/wntVE/1qiyjwg5Jljmb3m
HIj8aoWXqSG0YubPPr2zoQa3Gefnd+orziXPPFMgw7A5xaGtCrC8ML7uykZ0hcRo
3SqO8Nnr2Rwffa5mffRa2kMXUG3qu71D2+6oOhKPId0Pp0ugCiRoGf3i3H91Xw/D
GnaCX3kkWXyTtZ8E17ocWQUjnLJ7mtR9SyburGS/6S3TMWaFy5LRNR94jO+j2oBX
HKOiOSa0iEClYQGLR5Ea5CyrkXv6V5/6VI/UTM2JPkQTLltIh3iUb0vC7V4ZlzEY
bD5s2c2Hfc5VZ7yEyuRi/fK5lh4DQNdwmhpP7kShOv+ch4TOVuD42NOnkiiogD2R
cjt/gMKpZwyj4xQsau4MjH5hwgPZne66+/fOZ8GMlDIvl17iXSaJN+I7zUWQW3mb
hyWCOb+N6OP703+5BMbgVeQmZC022DJxFQhO1c+XrJwr58+j62/+8+1HJC8DXEjT
DWoNhTlV+MudeZKpGyh+GhCko+1xH5GiW1MedmcApHRGffrUdOYWmz0HQ/ubzLbF
kitd4wWF5jlt1Mu4d6YRwJDiiMF6aRdK+3nQONwqW2h2c8qpB6bn3bz5W6WLgiVq
NC1nV8mLEaAKYckitVi104qBoqlW1Wu31VLT4F6mrLohzAZcy0mCibbG+bqRtSDZ
K9ews96tNsIFSGzzmusL5jWiD6pn/0TbKjrJUlwjJhVj+MwCuPm1OKyA0jc8sxXm
8IONMjAXc9Dfc9iDaSzUo8ovgVQLSaNCS2il1U+jRPi/gMw0/Ya5+gAUGt4lzYbt
3159eFeAqqIDydyobQlEtVcsKsBFg6Za479ze+dZi0TNlwVEUYPoPmNRdGjwmbqr
fcLckZeBIsMQZ5uSTAjZ+iUJiT5MeOh/C5wmXJuxRk1fboei2yy170Y+CNIOePBX
USOcjUKkwUgCd0mqwXRcUW/oSSkDCaqjowtvIJ9nTBTm9RYY24SZ0Im4y76TNCVn
21ZdBIpe/f+op2pFo044prdKFlCsOJk2+Z55FDC83P3CYlpPpJb2NlfN/UnWGHv2
Vks3q7Z/VB34D1jWVyCZVgI/xuYeUje7H3kSfDT7CqZkUWYBT99j0ct0Powbsiv8
00frsTAwQw9YIwruljrBp6s3FdCylDHKEBhI2+/Pj1/sAJunpjHxGCWgXOzKDkgt
O8z6UkvR6gfW+SRxqO9kloM6pSsTjA1IutcltUs200c+paa+GqqSAN3gADMHBdeq
U8OrpMsmqVHCSvLWaWlqPPYgpaTv9k236n/juZJ03Qv5QWrOZcVXVmfXTRcxwB+F
v+tD18+xgHshLuErwPHm2rTkwNsM9tK7SuVbHyheR3aDSDbCj9cA0gfCeUMrHwxP
COnu6EjuumUqenZ05ImfggI/WBKLqbPQQWjeJop9SGvcvn05Q6yXXr2YFD0fTN3V
1e093Crhqkj/+0l/NSkY5lZXqzFyhvDSVjqwEgm9egMvLl8KFtDLK+nk7dzJ5wke
rJ0Hpes0RVLwcTkqlOjP9v3NFzyv6gdOuuDNMCtOjlrmKtWqF0MTUhT1qmKEMxxA
Fi1uDXgAaHaTyKGLk3lAbwf6zgjruYVfB3vr+Dijy1RCoVh8Xtp1CyMol3uyHNUj
6EP+12jIrENd39Bl6XR+VsRphEbn9/tW+U+CFf0dHoh/LEkxao7rXhy8MgjglPfk
gs3V9vEVbQBVqzaeTL2X8yz1xAF1Pr1hQ9MoyYanZwLCVPlHYOUnct10ITM6gb0g
7qwP6w7KIOhlNARF9ijV738qt7JMTByEvVA0OJOsdTAbE0LWwN8j3LLgQgUcIK0R
Iit5QRozJAVFNFDFemkGi/zm/XpmwAdJLRofS19wZ9LsgGaiAT/YHSpihwqJb+aD
LjA3gqaqsPs1u5t+SGbS25mNOsqOOKjfu2cuW3VQzacZj6JF7g9n47EI1BE8pKK5
aRfFZalVY7Peq/gSFcWNPHRg3ew94KXdj9yj8sFSUZjFe3Czha1bAyAv8YXTTLl/
zI7Vl9VOwxHZ79a47pDDdbtqHBDAGSeyL5903mHfSmp40q3C0n8lZEkBDeU3Uc4C
nf8SeucdchWczV4eIPR6QV9M0mmthKfiS42o/cETvA6b0szP2dVjMu+8ignCszda
ydkehsWKWXWFtyPkT8l3SiSQ1+bswTVNhBHjhxn4sFQZOs4uXNK4wv2qMRWANveC
8NGgxQfoIMKG8TW4gJE6V6ZOmfTxzmVrOKc3iND5RasddcVdCclOg8/20w44ek8D
AL7bnrrel5lSCun6Spln0J42EVeLdvj0g1fbyyMUKSO/Hngp9jClv9diFolGhtbZ
G9ch6h09ePN/x6qkrm42HdEw82Ijb1ApsjhbpwkLUI3OxcISIxzAGPf7f+EJj5+h
l/naO+GnR9s7NCPB10JpdDLp7vPp0gC77vxUwdxytu5ht89ciQXmUAzPwZDc9PDz
nZttmtntX8Q2qKHCK8ATIPr0OxhUTuAUDMMO1Wij32Rlw5ixlNu4IyGS2aX7GDQj
9K+2S9V3Bz4IeDPhdaXh+lz54r8BhYN6I4+/zpxxbDZS2s9qbWFbKiEoU1hYLsHh
MeQEsF4pNgWi3QmC2u7tVqag2Ew5cMa9XeGSe1fL5Y+FjLbfFBw2mKKfNJ65c4Ci
0KntaewYkt1JjsvN9L66WjRLrEYHiTNKCw2Q65QthXb2N1cFR1phCwxzmwSQdTgw
PSUmpDMtYpNqLF1X4meokqRIT8CQ9ic6YrpUCQlVpJ57aLz8vVTUaKXPrkiPZQH8
35sT0QZTIKBB5NpiAunSHq9RdtIY9CYqVwgnKa4OliPI0i2RCasSB9TslLaGBL7E
Rln1F/1iIAEM1PdNQjxG/6vCyTKBFa6Gn6LAymul0pNnVbzWykzR60FpHx5e0z01
6OXyBHd99VSxA4T3x7hn8+4BlmwbRl4IgFLC6iJ+Gan2PiKvl6xcrhVzxm6gIYjt
j2aVwcjf6QuM/LhOGJYvMI/F3cC7Y7Xd7IOwEiqXHWJgnvgjNewJ4M5oLjDj8D6G
X5nT2Z2Rlfw5SfqFNvs/DHWODLXZlbh65/b05BMLyFjwc0BPXxlvA2uT5qCLOipJ
Z78bYb9FZG198SVTkgGYq42uXhLnpzTxUtW0IYw59hmtTVnPjjyValVik0/OI6sB
3aN5m/0bYm2byLj9KGTh8cinZWBSgl8UDEM629jwu915Y8TrAQ5r58wJijteG5VA
I95rHXjw0WRpa10rVM72VKCPHuf3UPb0D7tiorl81j+VplPwRymX2wz5tZUTosKj
nJP6T1xkAFBgre6NgowVUiKLs2Hepv3vlefZBWlf/bMypb6jwV1r7ev+SweiqpMx
1ca8jelsEyApXvbE4MsaFbp+9ySthb4x3oQsfJlYsAVo/eLk5RkwgUow3rVnQvOu
53xNiY/dXJVgH9BvobXwUZM+PpzsK+1MrxZ7zqnrOJAoGyuW43Qvsr7K1b9Ei9/E
FH2HH1FlDehF42IeGyF74zXa2b+3G+mS09MdAHikqfRta0Gb4zXNDMdjvPgu25gu
ukXwVjImj+hYm2SPCL7cw9enBAIAyeqX3FFNSywvYNohWH5PK1HcYeCWEmbikqy0
ohveMNpMlb7sPn0I4//kaLHOyhOcoH68Lir4FEz6xd0qCgMjC8wBRXCc1KK/4RWr
UI+ZHZ/W2di7dkB0XwL7IPxYnIfNDdS88eaUztHsrrMnOqiZs5pfFFGl5R2rNMMV
nKNcNOOB+JZdeL+ceYRkAaPpN8DCQJ6BqjhUjns+rfeiufoXs+AEOK8t024Vhw/v
VnYCxR0qNpd7UY7EvaKXue2CEuF4g0zN+1sIoU2nwaYraVJxVYenuhddvxnHxYAB
DyKKADd3Xl1B9Z99GGRHOvezyZD5ZjDAXldcknnn7J7mpx6QCYov/TBL0ilJHPx7
z6yMnVzEtLTNOis6viZGlmwmon3VeQy4/Kq0hggB6CPDJn5GoAkaLqWArogWG5sA
Kw02nDA1iuDSJivz9ksXfstOVbq4dzhcX8ilSutXYzutA/i9SFcnWTV4+xm+pLao
hlRazWSRGGxT0gbJ5nHEtGsUKw/nopf2+faxKoxPi8Gj75Jownmb9JqEfcIthOta
41eOLBgVc58V2z9hgE8hJ6e7FpNSndxsokxtk51yCz9WgpYszMXvPtDfmrgjFb7r
BtdwYf2gBe/5ViJ539mjlzYbemfyXbOWRNjJBsxQ2+7wtux/xR1MCw3KUwirckRR
YmMRYBjTwbeshyxDgu0pr8xoPRo77LCPcGLf6tFD9kIFrbspat7xeC2cwuI6ZC7l
V3jdrn+9H0HeKjHTPGFqrPMWRofnJzRDUKddp7zEA/e0L8c/vRcrINZJgS4rfr6s
JXW08f37KIkdNqr6u6yhDP4baGcdBXlwAiwdjsw7QZDVg6mLNf/GETUvBRK0w0S+
ELsP9RWVKWBXNL+a0qjzbzSxo15roZuZGV5SftemnEwceayul0v/E7Es1L1ZD+qY
xnGKCbH5uKX7oCckjB86J01W8+2iTtubXLp26/5RFmR8fSmZEkT6lIiAj1pYaDOm
R4/ZnFwZuFCTy/TBd+C7Q0m7TiZsCVdcE2DmbCvof8DYgAIlPYvdTpk7Pg8t1bme
xQoma4CV+xmOd+7iV8VFGrFqCrX4eZikeqU+L/Yfpnfrec2A5qvpCadmlhWCiQt2
8yeW5squy/T7zsKgHbxa++9B2YZq+SmUMLv1QzYuRPMMf46VFT1ySiTdK+YZd1xC
oOdAb8f+UoiAuv9E9W4AsFBWg3HbcYJ12+anETUJoEVCAGF++6KLPFUBe3zu9u/0
zYGnDVae/BodWYx+wHRRfL51rJcczS1/DES+nO3bfJtPHHzZce45i4gPKmfS6WG+
OLwNSTkuxDVUXIC+NiSuarquGgWKsw+7jyXh2Z+Uh27DE0sa0/a0Y9ORj1zza7gH
YdeM2Xti/bw+TqoodM7VlmWP2jIYU+cl2vbbLUNKrXLMh4YO/yuOIKSDPqruXk0M
eIC6IZLEvOli6xK5M8a7JIpmmWDM4HBEJ0dbphcApUoE0jIyQCjGMzvKYvftMIE8
xFY+qxfYEn3Z7EbDdDA0o0z1bcdRW3Lx2jJhgzNxbD8urSE2jE8/XE8qOFNl8gnF
TN96VjYxONDe4Kl0WZCt3W57XkMYKLp7iMnwrIUY5iFJUUIyK5tnT/Eei+2bYzvV
WipSPje1muhMwnZZHO8AONec9Ro261nJvdKj7AADAs1xJRAIsSDzGO7/VqU7eSvi
5DQGOZptAlPN5ElMrNx9E8WNEG847mnUlCpO22vFvOeReI7+j7EzbH1BHrhRBN4y
pLWTJBO/rqHj19FsEmptwIsRVEW//SnZOxg7YdRNOWLQa5yqNf/mefXsf4Lslw/1
vpEwGSQcxE4aTaGcUq49nwFzmoRLXL3NHWDhwyskEB/2PQb6t0FNH40ehnT6WP4h
GS0yj8W+ZFNL/UHSjA8CkQXrAtdr/0FJsh49iGcNLp+njGLwIdA6KhVo3kV7XfIv
3q/gQDNCKX4ox8D4CXUa/xRB1T8iflFoU6TL1wmZwMmbQ4pvbsatJQ7r+4wAZrEF
XXrhPYSMir/iX7+PE9WrR+Lyi+BJN1aTzC01nSCsGJGuZSdXpCkim58W2HHqwuB+
+08gZBvwirAkTutPCtd1CYkLZkOWKFozBjk/eC06OWolSTdn3evezPsZLe2Pz7dK
zI4LvPR9rYStOUqVeS7y1NeaNqyGV7Pu8TTQlLUPimo0GW31NsPNJjKbIglCcZhZ
vJrisEcMQ3Fu+/2+3iEyZM6ZQqsr5VhGsuDl/uDa5FAIpBXUR/BgKXlMbqP99xU8
CcXT/xtVmG9JyoWdXJVbjRdKN9cOtBxlyRJB2ilkop2NP81QFleVDM3cbrduj3lk
bdfMNG8CJzhdRdd+3NdhVmcZHb2itc2sPn9F0sMWFKhdvKev4EIAhQCJSH61pCs2
Qyysib4oyMxtwgbkubTVcWxfmZin8hpsclQj3FtH8zQccJWEc4VYwCVeefy3uB50
rweVDF9RVVLoyr3RhkTny8YigssrvjpBQHkrr8zo3E6QEml1ve5CpEWSeS+BqTPF
D9K7zDtOd1fnHgm3c58OODCUKgytGqSqaJPaOcxhey8P2ga+5NKVvBKUu3xrs3Yh
LvhzlPlijuv2M3XTKpwrn/o1APC8T5f6DrzxQM0PWfflshf8ej35gdnjEZ2s7m/B
B20TrGyDmg/yIKP5eg0L5l3Y/KrWwK3OVH+aAy1frNabDUfPOcXD3It41xELGNnp
yraHg7F6QFyuyx9LDz+9zVU4Ekbfp7zMKideZNFA8kPj3uA25RoXDgmP18F8KPQW
57dP0m5cnv4L7XOUzySHCfBsX24ndsQp4hy/CX6qXUSy++ZvdhnYJSJaq1m8W9Ax
2XZKaaoeWOD/fOB/JIoZwc1NDOJ/WYVhwqx3g248VwycEkEtPIgr4GRVcDVKw4/6
0REqrCshi2IvgdJkYancFgdQnvVnePQUdyQiE376oKuY8AVWKnovlqITz3sYDksj
1XY+QVUG7EH55NNvhnbQX6ydz0g5cxWN2f0hQekpi8GkIA1lh8ZYUwOwks0kYe+l
8A8cPh4gQIK6HHeSyMKFsw5CNslo96Z66nx27swdZa+m9V4BbSDokig66iOs2SSk
MLexnneRr5piGyqjhKmsATDfYrVKZNAPmekaiOZ1BSgKnfr4q0BQ9nwpPVkwXNDK
7GblIKHPHek56VDZInM0R66L+gNKVnPk8xXGPjCbLmqQBE/n6etmgqJUZPzrRNgb
+N/yNuMySXJqBUEw6tirCzu7mrMVokYdsXzq3Anb4bHEM9SFOL4SEq33LnjCheTn
FffQwCqzPURjs051fyGHWH8nsOi1PAOwYbsbM4Y/wQYD6Si7FM8iGq7BwFPeXiko
lJnf1Nrh2zWSG+TT3x123YyqDbJXsmjGLVY5Q6s+o4jaj3w2yBUN5VPCuSb+aSad
QgLpKYqHq7zO4kad7tx9X58L3sC5EKY72dkA1+uOJsmWqwaTH9Qazt0c/G4H9z3J
W7s2OQYGQetd5ivhWSgp1a2TE8KsB9FaMuFxHKJRAmYOIbHaTh0lqEpig2uTpvqI
VXPzgvGIeCFENFXccJEvioedP+JIiigrHChaarZUVmY8RZ7DPntLEPLtb+UbbtR5
jIwpIMnKyxbAZovQIhIhZaE5DlLuDJb7Nr1qfdtJ2l+nFLW39SNK4kqikJSMPyjZ
Ksv2peGGiZMUucS+XHkZtJmmzDTdqQ/DWeBXQ6bANQP+LLIM9sprzDcJ9dcDqDhE
UbnhMpccdb7ZFkKPcBwXjI6mQXjbkUUNjRyKVroBeOFB282kXZt6RNfjpWjt6/Mj
ykvW/2vH8MLX1Vep8BaddknREYEQ0tj/USdVRSTmTbgsWCIjvMpceypd4MWE/URQ
KkHghKjWzidI4/5YsUXzGeJ5mpdk5WUIIgLi5A5V6QUftc6EsqUnOqxAO+nnF7cQ
h9YSmRzJrMfvzWu7VyxLqmorxcGOt3JTpQ1AOrTMzmKvRC00KcfjSqYmPHl0dTIH
/6h6KKCEkD3X5WpZHj9J2G3QIM255fQtT35HvaZ8NYdk5ISbrShpkp14vGOWmzYz
Ure4mKtfWWxHqT/OJe5gqmFl79gkqjLRC30WAc38Dha+4On3nw24CaVL46JRQ848
aboKlxpGv23vC5vzN4D3NEPLAZEQt9D+7csvwEaN45eCsgsYxfNcC5Kg5YT++SV3
oTjmPDCdMtqAtlss7TL1ozYNHwzl/OhqQFkW5keNOjbFutAPVtOrGDQ2WX5YNe8T
8CO6aBKHxDIQTYjeEWs8ipgM04+yLkxiuE5y4D0DijvSdx83UlLvhjRt81L9z2ce
qv+U9G4/OTsOzI37ZM6TMjx3cjEpPSA3MIMpyJZyqLmgnPZso8vTT//dstdBoTde
AXl4E1LpWFUE0emciAY3yEhy9GOOWvmtITn47KYPunzJ/eTQKg55FxxCpjRM4Rbu
iODfEd/1ncFBr6ANa3QGU/uuZyV0wCgc9J+biqjNCkyBdtrOwqtMyJUwr+gx1Qn4
1RBZPA4ECbeD+mFoXM+EapVpurnHJhl7T9/9OVCQjUrmiozLTbzho3Bn2JCc9QCk
iW66Y8WTwhaMKLDWfYA1DZlSqkxFxa3HeM2YepfhJnlKH6OthQQKu8LqWzgDl7Za
nMPlq7/f0cHl7xmaN6hJB8p8NYYiNjUTbvxNgf/jqp/mlx8YRObyTCuSBqAqKOjs
yGovvgGJj4Y4ppkEtA9Ts7UmR+KhWYhGt1lE+igH88GunEHoR8Dd/ZldUVtYjEpW
eX0zi5l6dZKAm2mjLgwM5qAfrUgrA8g6Gf87VpDrN5nxGOMc1QcarAP0foL082+0
USQemC+IEG7ICQDbmh/qaDlmAi3Hs1Fz1BBakyLEgF16ojA3VuRCtGksyaxF54F8
Va5yo3xC4hX6BOVwhxBiDP9jEpzQvcdizf5RqtUhvOEm/xUyOeMj4AXfLsxffIY4
Z+mSuii75AtDIQn90LGijmo06sdhH+J017GaiQzAMXTYubBNA5YkAXSbM4wzYhav
oYH/Ntcj7o4kFoq/bPSbzmIO5NOsbfDU2alq1DAsrvRuO4mS2coeU6YED/pfknuA
XfuMVwGB/AWc8fr36CJXfKwuUHI7t3wwF2/E/cLQN/U9rQmcWXzVGl1+lpoNT0rg
sXI7yWzWy3A5V2TNBICiRrEAsjBwpMK1uUW+qtcRjVnw1E4bnnkYd+h/ogQxfb93
0oxbyp/tD9gl7oiP7I32wBNKe2jHH0PNnsOfs0+PLVVjt478JJt9DYpJBp0K7K6R
TAFq6r7eWLjBRA/zWDgXb54hWaJSNU3TRHPmyhCVJN9K9PqViiXNMqBnioFFZpco
VfZiMN29nZZjoyaahuxqdnTquWJrEKtBmnek2DDWdVDDBdxsrvJscuQNV+mZ1dcW
jczXYsO3reXL0yDZnPcqtxpUEQUcqhUKMEIZR9PGilbjBRZC3SRZNWRMMdQEpjUL
vNVx2pNYf7c8hYb/m749oBV1nPJEOfnTXuPb8H2B/8shLMxZYfvFZRS9PETtk3US
mDEQ7WaMRSdz/iFpBxDRvaEbX4pOfotzsSzFtInSoIVaJrxbYdbHqy41jSNg1TNK
g/VB/M05I/eu1bg1FHURTvWPCDCARG76nIULsZqcpf5/hgSpqe41vSxIAOsm+h9G
xwV9JrB9stUU7ChOpFQk1bLz4M1sm3I8iDe13HN02lWkXJ92MQbcVRFNz2x8KdDq
FGrGNUtwWqx7eiL9D7rtEaQEX9Mp++blCHIMFc8nlQq7RyVrgjGIf9cz1AlmXfc/
vD0ktvPevHWQNzKG5BlYw9EDq/inTWYx/xDh2Ie+QMJsUbe4iYyBPofV8bE93Q5p
zBsxQmmxH8CHREP4ZK/covrHQNwioLMBTl7mrf+FnYXjrnjhTwlU/8ZPy/gxFcmr
B24A4Gxta0yu8Yb4i/vqgU25Nmg2osk8vj9NULQYeEt2iXz2iSpIvSU/yeHZZZuz
uXDlxGOs1//7YbzodV3nCitdwvuD0hyRSQKhKpNEl0/itUKSCaWnFwcZMsIJY6x6
Sn8UhdizXWf9spNEg7jqoG40Xqkn2zqOUB6TFd0XG0Cw9F4OM47BMJZaD2i7c74W
6NbgBu1iIhvijXCCorH7T6QW1LUk8nWoM/QCmnSvxCs8g4Iucz1nCZvnB/Ba71re
4QvVspVYA4amqzacozmm7iTe0hipm6kbrxZpNcnE7TxmzA3Ct+/C4w9Pa4OO9BOj
zapDinGDMPD0uqqhv2N3qSE4WkahcruTB+NDzPtX0+7WeOsv3tOp+Lxzoa0Gp/H5
PqEpeqSJ40sD0fzEKHvl/ehKndOrAWOMbx1nzyxjC2u3C4enkvCO4meiIXk2niBH
SOjyHW8MG7Z4pZnzYmijYMkdGTis2LAPJFMe+8RAKeLDe4YaNFob9izbkzCiBZ5B
gP2+lhPU4SO1CigZzcaiogmRRzLV4JGoXEvBkujedHjp9BSFYg9t5njwp+nkIgHD
BHXY95HKb65/tvFJ0wDyzuB5eRUUXQ4XVbpKiLsvCPYTnqeMlfNHLr7m5rvDSQZJ
gcIpE318hjZzqkgWDCWajlONQJe/intvwTeP0OQN+3YyKasASG3/oqcDRi7FtXFm
F0324B1c+yHXBb7yVQXTMwEocWbQ9r6ACDK3ov1mbSNcjzNW7JQp4yCY6Bqn/PdK
LjzhgvoAS4t9VfQXD4fGYTvuwzYRMCf+4uvzULEJkERoWatIq6vukNk+ZVzP1wkP
RYPVyoO/UMaUaMvkjBVpSOO63ne1hjyKwhBOb2IuxUHhjjpaDotT/VojiYue3Ugq
32vridhstf3YzH8K+MsUKEsIjIGYuQ3U2o9YDiJv8hfEpJXIO1f5bhrvGg75xvmK
3kE/ERykSElbfZmFqOh/xgoRZXHoRCCsBnn9b+CuCkUjzfJjBFFIMsogS02hehjt
B1hln/y8PSKvIFxJ0TZlh2zZduk8C6RUavnrd9ijg15szCLxQbz3J3hwJg9EKCHy
7/dMaB7laZTL9xw0+Zxa/uiRBbrlIpwtCdOkaUekj1yAOQTlts4GkTmSjCKXBuD1
OU7cVstTXRUwdbUAT5Id6xtEOt6jnYUdt5MOw0i7xDXrp2Qv5nXX1856Dpo/2A9n
LaX37gDIqthhUEKckZlZYeyJaXpC2X0n7sxMFj4gC9QQuTH9Rh250arbP9XrzzJS
bcBD9UaN4ya/psw1g+bXDRPtutKKuaDVPzS3yFyJUWr4FBs88nJAngI4DXj4Abvq
rAX7kTlUC2VAuJPyvlUKqMM/4tvRgB/M+uHArVYCzx+Ush5z3qr4IrlaQrUzNuI3
AtKyqsi21OjuZsxRnFacp7VYuB22d2/r33xOue5vatu1ujChGO0UiCG1lC4DQ5IR
v9jSLH5KSFqk2XpOFMYTR3IpnsyLAKRh05k+EfQyOuFRzNC7ydP8jx5EUTTGMkZ5
Ix8MwYwMT0aHiyquI8TSuXBQZVQDcru3KJgOfoSw6LlJw1AJUpOMVSTW3RjIK9sV
wW/R8Y/9PtB5O0RzAKgQzlP7E1QnFXxjk0jkzC4qFsVFyfV7ucfYLnyQPuzauiaI
t0QPsg8QfaDYMoFo4A6hzzhCLybc17zEI2EAj4FrODMtKFn+MyjVsJtuFUSdsnzc
71KdfavpVZSabAwt6Gyt2M2qyUzjV/Fp9ewBM2CFoLAE4w7AJAUdGwzd5GQYpBM4
lIWyrEkoZ14g61kEYKzkGo1w66epBb/TJ7Lek6gPqL7UvvrcJkvIgfFPm2EjPGwf
1q7s0y/Z8mbsiKLPrItcsYqLZoxu9KaO5Jnwfpkebu/GR+lFZWhQyMxOxBiDlE3o
Q7eW/AxYVAgCgx96eMb7ZBFwsR8hMXiAqwWxxwMCXTTpSH3pfaNp5jx+sHe223dr
euMkNgme1UN7IvGx/ECtIkJDwDPEHF+HVU3Oa3whAPfrBlHk/vGGJnh94u6SsKpk
Gqg1/fwhooMTTZnotDTiPQz6yI5jpxvBFdmNgq6L/ZMJGmaehDzdl6bunD0JQ/kN
zAkdahZGAhpWWVJjdZ3KtNDuQkMMjX3+xXxBVUpeD14oIX2aK/M9AbkRA8cQl+80
yg2FJUIoQDyyFs0I3IWrXw6zm6erGBS3Cm+5lc1SJPGTT9d0vdgCyzWkzeqIPLm/
AuTwpuAZ2/7nlbYTfx8XvzuUSr1a6vK8VT+P5M2/1xDEgRYs0uMv3D7/bwdhbQfK
LvucrdsSvAq86PpLNh7E6DHq31/0UOPMEa2q3jK0QUV5FU8Ti+ifAK+hwqqqM0i4
yuicVeKETcZZHlMJ+dSaXb9D59rvQdUz7wqseKCr7ocq3BuxAVLAbhl5lkJhQPaa
xf1O1Wo791nGj+0FmIabmU9NTDP2NkKriU4SmRb+JC69lY6ZVfH/rhrg3a8t/68V
XQbosaqf2YMEdUU8J+0UKzCM87NhYQzU+whQCwqAXriJDmAENf5aNo/qdEUDO6IO
gGSX1C55CEAHMqDqJbjPt0fOiiU0xXBEl78WEGvCZamnIiUT01WSaCA9AEf+qXSa
Q56A+deEOmwdFYvuzqJFbXGH2OUhWdwNx8FbAoLog0GhIMC2PcwK/Yq3dAezUTJL
WMz0HWfJIoUinzUjeuitBPXkflGKIQhWkT4yjGZaHjOr9uNTTxlkKiW//HXVwFy7
hMTxy+kg/8w8A20eE7Gk1ku3r/e3AnmczJCYL3c7uyvucHKT7Orcr+pmbEnGwH6f
Clxcvm27mwI7sPNeC0JOeqmM54bEALLViMfTwlVaVMYXsP9SAvqZoZ1U5jBESPTj
fyAV8NACkeLbjgHO2NDTwT22CBQfQMlLGtbgF7gosLobqBL+YAcFmdU09odVAboG
RTD3Qth01wK0SsNLtLCq5G6qKuiGJZLernW7+fTKKGDsFlQWNWD4tbzKNJgDNLcP
frc1bsJiugmw0FV0NB+x9oaBKlQvE2VjwlnMvmTC2t0si/0Dkxe1XK3usk1Gux9i
bKioPx2gxneLMflmdIF0l2efrT3d0pQr+SYxRqrh9JmIww29F2jwvBk3LfOYpc+L
+DqLAL//9hn6SpT2eZAgy73BUoYQWGl6TRYbp9uWkMMNdJ6uGjjEo5HxVkaPQgvU
cjD8OduQbLswq9eF/HzGhCrr5qkXELbt4KXel8A0Zg+f6yyc4C170mUWSOJadnpX
UlNqAcFj8/jZ+eZFnbGeXQONbICHKlSUa3BhwDyriBUOhnbhbE208UurBBANuk8Y
vPAc9y36Aue3wUFG/k7uGeVcadAt9oFG0bSLu69r8L1tUPO3U1+29mxbaYAvp1wa
HDQYByJXdPe/BOIfhfI8R8Ww5HsXjp7YNqpG4RbXSjeipXXgpNcW/mAmsLi86r++
HJWS1qmSCdrioz2Sbg5XD2aA9e8lSQaDZG5UX+Kcb5U0x7gllVk1XzFxXdOfq4vO
frxzM/AyJ0MIivStgunJE6dFwdbRjeYu6N1Iv+rDdfJmPsjx8DMv4OSTPQqPq2+d
Dw78231mOvGsLn5puC40K/Ok3fnOW+3NbVpJsHe6oYtHt5Lg1AQ35A6GAeZpbuEw
dWKJSSeFYCnhlq7nBtO/XyK6+7CF8nacMjy+ZVy3+K/JQLmne4/tdJmWOEhn698/
FcbkC2pUYDp9eXm6WFo014fJSy/++9bLDHYgxOywETMEYK6DBxVIcDbNiATMkJOi
yNOTmJaaFfie7EqcKM06N4S3i2v1AsCPEo6l0vvzlOi0H8LyyUl7TBPIi2no7qdq
cZVNjLXEj7n2o1GgFrPlRlZvHRqIrOIFG25KIAibkwJvgBGYNoyzevZ7TEKrr7u5
GUmv00MS2J8VVSVVKPei16Oi81OKlhDk5wZEsLt9n+w2PXPgiReEeu4C/Q1tir4O
5bh0FndQsVuLV3ujWmJ3PGscGY3BF7jrnQXs+e6ExGi5EPDnm+Y0EN+dyvLLkBaG
7jixtbbHvmXFpT7xAiHVIz6w/DZLtm0xstkL7i6HDVbAsy2wrZFM1nub4kcXqywr
TuWkp9UgbVY9++6s8XWeWNpFLm4aIv/K80uMOTxIh5jvRTwZCIt8uD9ZpytEqIfi
50+q/EhO/Yel4PbQ1kzTVEjXx3szk/4wUTuXXsbWNjiVtIONhT37QJVnOFxDO6tB
hcUN7sNDo+sB9Iq+AdyQP32ARSxqiyRenaZw1ZX5cmd61kLkTpmfTXMCcTRs/SCT
bVdKr2v5ITMiJtPrcEaVLRs6kK96bBNNFMYDYFvzoV+gAUGL39tUsbfxquV3AA7A
GbrdphVeGjzg8RC2AQgxPcz/VzwPHVsWrvqbEamxtj/DrljE75T1lxPaoF41Q1LG
/6jOAy2jRnjw/2s5oEdZELbulKNQvSBoo/tauXPgPnxP51fl1UnwUGKH9XerBT5g
TA1en6DnE3XHiD3K6QiCuO4rjc2HpKxgI0XLWgVaT+UeD6DlkqNvxFGX9pEJrVdw
kYAci0vDQe2/w2Urgdh5XC1rCP7b/CWFWCk67Uo17YtgycPaRXS53vhVo7xeoefk
5g+aXy3O0T9IA1uLJI1OcA8briBMPmQTYPmO5rSTbUMbQOA1aIU/MaiwPU/cB3fs
S6cbyw+DdhYoUrCMza0I0U8iVerzcbXuUjCbIOJW/fmOcs2F/NjnTwB9yFdb4B4n
dKLeZMiBUF/2M9IeRPEaVxMNlbaEfl2eFZ9GlHuM41wQORaxqIA3+hvKVwk9GvAw
TKEzVdW3O4xzlv2n6rTft5DeXeGRUyGH8PAaFxdwoiCKEDOpcwH9V4ERuaqeDOuV
jCqNikq6Sq/E74ZMRSLFNuFPlGUS9gMY0Dgq4z3z3jH04mCWKTgzB9KGiOMENbte
jYsr1MlCHuG4eCaEMh1MFWR7Ow6QaqwQx0o3MGsgKW6xgS+2J7Jj7BViaKvkbOEL
uan5AgGBtZ7Ht6joiNV4WKMZ86jAk7v9/cHPaSym0FVnYutcV9Tpe35ag3/tobME
NA0rjuKso/uvlJh981l/co0IBgXAZw+/0wSqh3I/+D5WVWSWdh8DdEhlKPFQGmKA
ogLaFLlsoc7zVhBoOf7ziJTGMjJtQN/NAai4JdfzxnEkhAmhpnchlAm3cfuJfjlv
+p+xBm4DzaOJjPtBXrDFd8Bpo5Q4My6QAlWgil7aPpP2D69JvBrof7BFcV0k7Y+8
navXFpUAJ+u27PzmKH5ByHVDQbj1co4UVat9WsV+ZQHXVczrrBp6Q0wItLyDiXJI
fV5eTzGTkm5tQwntyfBWhgv4OyX+yvyiyd2twJTi3Hh6WAxy2xZfnHHkpssqwtF4
vPPuPV6uJjYQkdCBLBUO63AOCKgPKs1f7j+hjRpdy+jJw33avtK0BizjN+grQZPs
2C7RNlD1CANTG4mN0jz1wzV2N4G3uBlc/is02Njl0DSx4+W+R2/xbTaJJ+5PI/2d
vgeAnLe7quUcK+psg/1gptjIPsx76tXcYpGeu07L2F7u9CBVXaj5ZX8XZMXo/Tu+
TaAsinqkzRNuNuuuS+6/SJp1u4d14GEMvAeL9kTSmCTAViWDGY2lQ27anhZt6CKQ
qQqdh1b8O2l7oyeI4eRr8Y530egg9YQrq0J5FtpHeVXS4WEdd8mkPKygxcJfPBGp
awvA+CBUlgSVnEX77+3AcUD2QOmlVf8eSRQeIlxadvwghdA4Qlx1sJZP5WYxgJAq
lHLibqliBzMuVpID0ZQyeWL83bsJLMFar/usj/NnI1T+TX1c7MvvehDcFHZ5x2Ye
IA9S/4/OfuaprGTeAP19/6coQVIvZqbIArkLyLv5OaBTOUjCzh2tnLkqhwr14NXy
qLhsPTMpyqI+LJCF8ua6SFk409i6ZCTjJmIlFiOvotwYQ9DGh5oaXwhu9AIKFuyH
V/qt2DNIiXhKQhVQYl9dBg0OHrVS/ACU99Z65elyQAMyzgxo+wj6KP8a/cxfYVw0
JY1oBWOueNPcyGtN9S3CX4XP0ABRF+glYZgJI9zffUKTGaZTXsH+pSfN480F5AzS
Ourtndi01QmPk8gExrJ4LfIpq4EX5qxtqJeoxqQPDqGzYIQfYpV5io6jsgVcoeKp
LqNo3LCYD5kFtacF8edPwrjeEXJEfy+5AJKMB3ajKQ6ul9e/bH2P/tXXHWWPY2E6
OZNLrZE2m36IV3Aw6bYRC2uoOKJAlNLNzuL0FfkcTG0jMjEMfiHyw5Bws1o0SciC
BPfERpGZFiuVVAxjdztKqwbBsWzJpwWGxN753BgMC6RX+TFGnov+jMCBwEiNHP01
qIoeZ7FeSKSdd3LbWfgw1Ctcxqcfioqn/wH1RXEf8SCKYWaV6GsSBVVxDXZ0Jt5P
oo2OFKALjCmyyCe2TBOFzV9qOVz06nQTX3Us4h2OVzkODncnrX7lRCaGGnEHR4tu
DQEtPwd0vRMxZVoImmpV9HYnF55up4hwzofoZXUvvCSrPeMic2Pjpw4mZywsrSRR
nUOK1Ed+P0kO+gy9BAcUSgxcDA7SrQCh9YFZDj1u6VSbYvKva2GjBq0OfLpUJbcs
FwA7f/ahdE4Wrf19ZF310Rf/KfLNSIhJmLMT6G9T23BDvshxebFI7p1CXR7uT/xE
mJA1ok5gqu8X0Tx4WsPUStAgDx8F9NYIHEYT5hGVpKlf54W2czFblwVipjUcdXMr
QT6KG8MmsPZtQPgF263Ci6zpqzHCxgbYMhGIPY0wJ319R3dghxfc5vzE75LoeUxH
a7KpbiqqONW63Gx9XBn4f49o2bMrPNuzPk0zrmwekf+PNcYk6BC9GbemWxq5Vw2/
wyAz5xvmBtJwchpfdknfvd1TR/W8Godes+YOPK4u2aKHLfKPLjvP4GvyF9f+zZex
uP0bntl/jb8LTIJqa/9xkVYvxfhCvA5gddgoVnAl/zfSGR3ikKqHntVXVAv76iQk
gSjpG1mKE3PeLkLmP569kLrIDsYXD418hafkesha95jc85Iw2+oBSOBCSEJ0J4vX
tQ06EeCodtMlDrTSXURW0BuOwxkTufuVP+qhjo038WZXUvSBae55FRMtG0FnwU1B
HysByq0dremZvtcNsChE2oOeEpDLKeSj2Y7du1Jkask7CaFwLFb2ZW3tBpGm20ZB
nqiDhIOi6w6DNbuagP/9Y2hZIlTHMbDQwX3vuStC3wz17tEb38Rn8ABe96CW0vPX
gGjzwNCPY4AY0yocRsfP8jW3uyx5QQFLiKZR5czY3+RmQXbEiQPcSKsIiYnXhaj0
IAk6ZVNR6lcxkT/u+j4D3q7Vm5+mkZ/QnL5Nx8eW8w5xiBQA021e62344qdrhZbL
w8g9D4DOYi7QKuaz0uhZ70nAnMC32IBuLSygcWdS/7xCDhOTI+bDjWzJNg9+OsE6
fJtphw1R64jvdR7Q2UoVdPK80rpMBQ1spVaLdEa7GZtPaQA6SfpaP9mSmUxQneFv
Tfk2YAy8L8fL1Spxzqgs8+namii6WbQQOHyBsx94/CZ00vL9gXwbLqVmJ1jT5jNS
8HHQw9HI/xTyxLugvBoVQb9x4IJIlKxxyCFkmURA/DuOHKWt5MbQ8iOjiWURWqpq
yzQavGe+vQPDd2JMY3o7LWd17U7CPH4uXTZrxRNS/YaeDMswPod1D7EKKY2V6rDT
gGFFUACQqgNrtqPTA2u/jd0RtWdprqiMgrF12FbVjetyq4WTLTggMoFGdlg72h3i
tz9dZmaPpfHrUQK7cU3OYCn1lQiSNghR5ngmfNDZH3eCmjXFJog6imo6cacvFy5x
qBKJ/jsejWsBqEkEi0yePvu+xhhLGtGbVLoGgHZpTeLn+kmFmj9iQnscPs9DSgVv
j6zTBCvEdRHH00ncVov5obNMNNt2GAPy8+OE0mHXnH3JCrRm3fBO8xnJuJPFcMpc
ECpSigkEQZfx7peaTvfzAC7DkFE/GPG+AO7v5WG7P4IS+R9QwZ09BfLkrULQBynQ
9ECARfUJFaRrMstLWVEuQX6Pw2yCFONY/UWFqKpVw5EQl/eb+xYQFt1bt6H912NB
Kupdr2pgY1pJari3sHiAjohQw44sNsWGwbtjVMg62/sA+APsKvDlpWBier2GP4RH
SVZLuyOM3DGsKs86nZ+pK2QhI8Y41VAfnutcm7+DdJ5wBsP0b+KAVZbmup/X+EKj
AI+HmO9UE12rlX0Or1l8JBBv9SbrUB6E/tQtQeY6MOE7Jri0ba2unsPT0a+GohdV
gmwh0yd2n4BYKN68YB7fIg7SUYeeN9udt2XW8DdWnSGH2ahkg8R9dMEIxke/SaUh
a9rDUAvY4lpLHijcVvWU6f7RsRQDf1XtyboBS4MTDhP+tk+3l7UVz6oFbCt8hawp
4+htW/HJfj4oL+QFW9PEBwdXjlcsFaUnEvMcJLSaYYVUnEaMhIBGdFfbubgMFxR6
DzmKaWQzeqksnDLwEF3JL8XmpjrkIX6lwHg1mZ555AncxJnHU9jOWb3t9mJD+7pY
fTTW8VMtzoRWx+/us+I9+jaFcy+fGffO9hB/WQd7igFD684py/fMduX+UeZjHMLl
6+l1Ty2oRVC2+GcEqTYjVEAuYgNavhwKV2WH0BhAoWjnijmAwWIVJsLnKP9uhTMV
t5tXSv4GBppVYupzRmxbRhA4gKRE24K/reMgInt7uVdrSKT20uyIz1tVRpE0RQed
xRH/7LNDb34rf25VkDKs9KYuJfSm9zp7SMAKpyK9actTRiIbPICGprPAVVP/ymgG
rTh6NJUruv9IGvpAeCeTzxCtFflP+fD4/PMLvVjO/O+Czg7dUUy6xobO0UMDRp25
0d+FJTKYSZh8b2lf8GEd5iMJhTMqgc3lPh4gh8uaby++iqg51F+zG+9yGP+pxikD
+cIbTM4TFk/XTJ9NRoKLKFuKB/Dk9hsSesWQERenkpZu/4PGuS0W/uFfSe6p5FSf
60TXRMDxvmSQFkMhfCG7AttaWk3sQUaflZ3Tu2C+1kViV1Am/XZn+ciswdSNFw97
joWmpExyexUaYvQITilBN33klQHsfm9QJIYEvv0qbwUKw5kyTkITLMl0Gd8/VMcx
NRTRLyxnQ/v7u3gt/tClDHDfyu+yNgk/m6hps6muNJyHx8NIBEQZs0G8dWQ5/0+L
6dtUKU/f29qP2Rc6tqx6HeAa/Wu9rem93F39fji+u1EQqV04vyu+vWc5f5nXTpvk
2HTycWt9zDNSy9aRy52oamZdTtKCJ4VtogdvLoh8UHyvlLmRUbQMRQYc9rX38XdW
pn8BVzKHr1Q1dgruVpbHc8/hqDow9ixK53d61XMx92t4ok90ZkHdMyQl7uW2Hs37
mj03QjnAyQwR3IeJIf3IV/3hXROsWeR6gTdDFI4/tuMxYV6ozSleT/4/jbPhxYwf
2F6LK4wqLFMLSEFw/wGpxFhHvmdCfN5CaqMSKtlcTXvqtdLoZyZnZHT8VmBGenSx
aSWDyXUrgI1pudxLpcfV6LEy00VN5d/pbAc8lxHNPOmXZTIrtgeTvhqwvVc2DINR
7NyfqcNWWk7sEwCI4qQvJKaF99xwkfkV4ZHxHwPqIi691iiV7OP2/ASyPVNv1J3+
dKuzXKZDo9V8iY7VUusAFypqTIClzzMenxkxF+idzX5GrrVW+tGiSv1JVWJvKmEK
iluoLjVwFb7m6JBtUycGgPgx45oGuuGxyJsoivcetb0AwhMbWsuFnmZmsfJR2G6B
wQti2fgcnGeFk0xrOD9zKnZ5MIvnmtWGmsixkyJwz9Ec1umrQ3vBAdJh3ZENQqka
brg3XT1yiVjDgxnT2zX0xOinupVECYKnJNJe4S6EbmXbL0tUFoIjzq24ysgoFRko
uQuzqdNl8raMzjS4MNdifdMdZAnKPHKTFpTQTXGClQeDlHf4QMl9jVmfAmnBuce7
8bj0bp4rrgtEhStUwWWTeB4uU043JNUOUsnNtx2Qvu9myOQkAzRk4xb8LSNmTbKy
ZfPHzU7v+TBkyZcYxJ/M3Bnq7eK+Ip0eGoDqFI72G5E1SvqkdUqgHYTzEV8JQo9U
hkqFfopMoI3IDQSTWBYHGUgPMbcP38qWwJkK7NxyqXqk+mXrXgfYXPiSiJtT+T6P
4R1s3bZg/rHGkVFVHFR8macAiterG+lXS5rPusiTk+Onz9hDByBv8VF+4QbDrrOH
k4ilT/NyAhJwosgqmf6fSeBfVNmx+UNqRdMv5mqw9/G6xE5bZDrB2sSMdMUnAjvd
mk4ocU3LMW+ftf2CPW8z/B80/RsmsQtIm3BINgFyBl2hiK0VbxAbkla8B9zKaRi6
3tUS1fzox0cSLXbeu7teqxMKASfWe2EEfYVtmBZ7Z5xrtqjDoPaoJccShGYa93yH
WoayfTwQGC40A7OAlSu/5cufCpR0aV/eqzHXGtxztZJupFk5I7hBw7zFYUUZnHpP
0HeUGhDIBebsudc1XufwGI1gTq18nLfjqIztHD8AsEGGXWgJG5/bSkhRtcoaXhQJ
lVHr7eUREbpVMRLPgjXy41JmoEGqaQqiIdA3EklA+Qimdo8njeNhyZrVAzALXC0F
eP0rGU9EgP8DJ6dJc3g4FbiVWOpCv/bgIkPgeuIVAP6usQRPr6moLOevAIgJJ5ME
6+b8prwzPa8TzNKxzLe1rAh988rFsv5gyf1lPSS+IZJ37EyAM8KWTD4amygMih/p
VWlyExxFrN87H7BqcZ5BIOgC54D/ySx3RCzPvoHdSTZ1muVBwEfCBIShlUO0VJK4
LR61YkEo724n++RKQ7z6RojVMgQePcf1/Br4P4UO9KkjV7WOIV9U3e/dN9vqDyr0
P2jAMhMhgkgLFIel4T8eUYieyh+u8zHH5mlAMfDXSM1Uwig1i3y8BxyvDOyAx8pJ
K4fBOGFFdAZ92HM/84Xc8Y3g/znh43ZXKpDpwE3hvHAmenk1CnoD3kHmtmn+9qa7
5JG+msU+hTAAnlti0CVJjyAA0TvhPA/dxkc3wgj5VZgwuXWJh2Cve3Cta4XyT1sO
DLl+sH5BDLru7V3TlB11lM+4XlLQGNNUSpUTNYlwQQncYz0td3klhzoqKLr2o5OG
z441c5tyVoV/3/eofS0udlfch4KCZix8yeGeaSp2NzpZG2PFDr2SsffrZUge8W1x
K16VLwh1yK11ZgZKCdrryi0JyQjNTbYdlHwJK6+Kuer759YKk4jlDrUxFv+1YMhU
KU3VM67mM9mTqSniV74eWkN1DYy/qyDRlo7/D2IzBF+h/M9eYDNF6URjD9o+OgCD
NDu48uXGXWM7IuXn0iHu+pynl1R12MsUAP8ls0bBFLieZylQ83LIfoCpnFAQA7ba
0dbIKLpKbnWUmfL7G0Ho3D1nt62/OkXpWB0H/sESCIQCoBSpLEDz3WZLnpPIj+sE
5OUT9EUHflMWkaGTi0jiQo10u1nEx8uVH4c89dFimzOhWaOTFMEpczCrOWJ2I0Yd
SkB3ynaY3jmcoIGVxwCdXTKDbiCukbQRgsycQj+H6y27/EpsdaSeV4gUBv/G3vkQ
S+5b2WKgLpaCsyNHxw0UB1iLRYvqXMXPKwmekm2XvBOlpPC7Gju82ckqbAwXkEKO
Hax3pV0jgi6YDazq5Gx9LJzTCpoWfL0obicXT9xNAujkIHUvJiZbpvNKMZJAmHgq
K0w1kaKnHz8GhRTD0FpFjo4PCcgcWc86giQUhWQI4DoGJuiI8upzo5b9CS+9nVqn
AfbVKwHSbMMGkYsl+vVX21vdOVMNLr51qzGZRN5nQTiOclIrVnOAr+h8A9c31JLv
zjn1Qg3EiT6zEqh3lI5qRusQucs5NHkBaVfAkOZqrMlxodmy2Kt4ieWMr+LXHxkO
bvKHVM3p1oxE+UaUCXRkJR6DZWvawe4EbP4m0GtCWKAwc+gWbB3Q1rOXv1p3kpYa
E7/Xs+OK/j6pyUnalqbME2vrXs+8qvqRr81vlYp5z7Y7u2PByPzaBypgbeBD+TxZ
IME5qQZdpe8NPIZsnMShlwozLY9+X0USNSw/MdZGIrFa0mgboEgv+CQsYNYcKWJI
qOszDhX5qHV116/t1C78vQvhnTF3me3ehlyMMFq1lxyw0NlOxUuVc2dWmo8Drah4
jAdQ94XZWLKWnceAH4sAkcXUPXFb7tiCQSxcefkzB22ulBEitHPuIPgvSM03/TOL
WSjYlR2Vd6R65UfqPdwFeY+IPANrluKVH7Dqu0qnlMAHe1SaU8J75hBrT4UQfN1n
+rD+N2+b54GEYFWquLkOsJhOELHzaNcoXuAXrpmkv51k/62tNmwnnmcgpjbXl7PI
QmSP0DF5gcCqWZycEoK8CyCagwZd1E7zTFY0Qk70N3TGYpWqM4FSBCJ/4SFmMuwM
hdE/N6RRF0YHngTgZi8Ab5B0jB/o4hbtmCyIeGpr+BSMyROrBTpH8GQLlE6Ue8Ca
PX0+9od9JaYgnVt0A6uUiP02X9gkgglIOHaE7VW445QtFOIosxElELwp4V40ivkE
jE1k/iZd3DuBicTL+zzrE3vc1bgwfArQ7CiCk9gCbxXFUAHRXDoAhSSrr0uA1J3Q
WtBOVEJd8hBErLU5b5bABNl93ltyubYMjWF+LM+OKIHLkoLr0y2kx3hMfgh686cC
Wwm7EUl+Xm/VepbJKknaP5DvTOoO+lZLbxXf3jnHspxM2IFw8cO+sbM/agPzzV1U
904mFjbPux1RfPVbUEJp0nc/HaU9pSe1FvGf2N5xU1Ml6QtW9hE/7fgKHgRf2OtM
6LI+3vBXXZB0hopbxPrpXDFQa5lXH12zM4zG05Porke2zmT0D46vzBl79Ky0hIfU
oDpJ0Zwu/3v6iDJ9vg++7ke2MC2C2K3tCm+0GhmfTBFukALy0HQG15WjmoEVChXn
zLOsgOAbdQI1+GMjTd5JPI5SXft6UVlf4gPTUHTVnaFzEikJdNDkgS8MYACbDKzJ
eMC7s7fYOnh6xBaW06A48JO/FF5Ilc2TwpEdJzUlPJamOXeplawO2LV81ujsU3Eb
1Q4Euzq3snjdMQu4/2ykrNhVd9xA2q4LGKq0GR90tnA4WmknpCVE06HKE4U/dfkG
PmYKN4OTXRijX9zdwgy3klNz3NF+QvlDTQeX7Iu/ywIQVzJcdss4O8crLNSAtev4
CcfeuNe/4LfMSPZYZ7rWlgmFTWry9cp+T55IuWmcQ5cKYPQdAeiYcB8TDiftaFtL
Q7HcyxvHYQhxd+7hE4WxSFzhhsIb1vcwU8htN66xsWQj493j5yPaeh8Sxs65CGLb
GPuaDqs5nkO+Ku5GOuJyTyxo2+Ad6NSwHqjrOL+Y2Dq+2XYSqCrJ+Lf3/2m5lsuT
Tp3MHKHvfrITFQI/Tizhv/sOVzkEWiQmszjxlqrPhY3RD74Vzg30E5sb5IJ9/3CI
m7inV7vYGTnrCjgM5BPDgQjtvZz7nr7w4HIvj/bkCojL2CbeFp3ghaRN/1rb4/5P
PQBQkhtXrzIJXHy5Kf1fr3G5CsndOdOZYYFu/VpRvrISHkI8czHJ3qXldnJ6VIBc
SpetgTyA3Puy7TzRA+LNtu8bV0wtH8DetiUdUATTG++l9R6rkGqpzzO1SVNSDZBK
Mkf/PKSNkE1lAnQ9w/39S1I0nfcNAcyUGUazUwudbb3b8cSw3W6y+wtZWsON/cHo
29TWbNBfZwffnYI0027tC4ckPNn5xV0xcXHB47v8uFPQxnSfcSgcpavb99f06TgG
u84iId8E8NmvE0vgJUX4GMBtsIs62dXnVoNbWHq9wDi9qd4ynY414Nh6q9ZjkZnu
M1In+N9iyL90Ea52oINOnkdsiRGaiXzCh6UD498NLHZaZ2hwlSvffXJleVbvuueZ
9Ex5Rg2QAas98Bb1UtKYhkmUtEDGWw9ytOCs1bldQir5exZFpnLqi1wk8zxarmBO
bXVTGspFIOcSMRODShwoyVjmd2ZmrUbJYT8/h3ZrlpYGPEGJ2bnjG+ZEN4+mNf8z
DLbbKbXHE2aU32pq4B1JFW+wHPWrf2JT0pBmwrj9KRnnLYlOIMOaalcVN0sXprMk
beKEUbLabn/alCO/l0X9cSThgWGnp82ev1xfMvEZ5J6UU/Ur1Uy6JkA2Cc4k6qzJ
J1Lg8HXzCMRbGqQ39tzqSchUyEt8Ih9NY69134zcNnIasUs+AdR56UP3ikJjpjVR
rw8CIOizSJMExNS8+X0ei0fydcEMPSu4J8bYXXjXEmO/Fv4IuWl60QWKjti5l29D
UuSRD1WRmEpfubWDRkJJGV8G0qMGM0eUExIKI29rzMx1GZAxHGyzOt7WzHnZ6Ocs
IJOaBUD9hWAVtdszw0fWzaT9ScLk5IuowrSn3rAsvXZK+/E/PWn6SuGunCy27Rcf
ZprZ9bFgjz4Cgo1LoYyNlOckHJDp09BKvs1gI2GD+XEGjd6sHMjGdS3pNeN03v/S
0By2ypnGvdpqVKkzgahMO5RT1evjXJztjeJ+L7bUGhQ5YYL7iNqqi+wBqPd6pIpw
T+YUW6eW8DO9CGmWuI+CxBYmoe+gOozX+83ekJmnytjTJdtyYMpnI4IlmtdBs/0K
yz8XeggHs7jPpBNBir67UZTGbvGto3tCnmvadjYa2ZfXt67HhPO8oNYFzIqyKEZG
ISlDJfsN3wPHbYyJYrjjeakYr48cX3BbkxbxFSZYsxdpRbGByaBcocI/SYXttT6H
oQGFCGqX6BarGXah9B/If38THRRxfk7LRIn/PPMsreL2z5I8nwZ7FFRwz83nMtUf
OTPC4kjOgkNNgNfg57XbsM27sEBGS+wHFx8XxaDDo9fuHyBHQeTFxNOYNr92RTOd
7YDNQUXT2RUgSUw4cjLeZbjDrs+TH8UlZwO1acRcdYm4jdj6lX+IAhxQnU+80wbv
Z3mCXZOUz5EWHhIRzhyJ/ncEO9OupY2NwY3w4MpNgdxhrXEHKKdVzjh3F6gXeekH
1SeuLnB7ynpSiDQbG1JeMiI5A4Q5DZVaqn3sHb7BMKKiZAr3ZM2UQ8lUGw6PUGeJ
rTkcKMQewPr1HwsRHB/h8N+6ECIu85Zt+bmiiV965VZ4t7Xl3wo8hXDxDNhaQIm8
wPsVCa45MSO9LxkrNfKJkc/NlSsVN0jEHd2b6jfLQLm+p3ad52EIfbKTgrVZxCu+
OAvtplQWgDA8EPAO+PdoA93hxB7aCm7sps2LdVg8bl5cvPYDTFGQdQ5PoE9ukbti
b9+O1HKcGDPxINfNvNw6poJUv4ur41dQR051bxn+JKPNgjXHsMNB2M9jxcje94jM
zmMMqsiRanNR3hIVT/B3lTIafEzZSh30rwMehpUX9dk3qd97wbWZ7BHyOEW1d6+e
zLS1Ay6zzAYvv5vFvTfJ+31FiOF2E5HekBqfMH6uhRfsx02osB04UbpYgVET9MHb
HPt1X/IXlta2JW/WnaUKQwSFnoDmcZCH5GiIrs4HON+gDjB7lGN4lqQdshOeO5RL
8v2xLrEwPtEKilYvWJVSqH4Upz/ElN30PHtaaeLsOoM4AdD7uztUzwSYim/iv0ww
Ghmt7eSn0UgYeo7Y3jMfRvKekW19fVCe4oFrndhZ6LCMZb4w/mIH3q7WkL9Tj7UC
sMsyV+lUtul0hH1V7v37I0hAOoKOTZvY3RsQciU1rgVz2m5ka2Uy7ltHv8wEJXHo
Es6iztyRWjwxw3eGCLkcBysM2jx5UT3tOLwUtzFdrqfk8+99AmAwd+kaqKo27Uch
Adnz/i48eVP/HsgBzXBI0kbDxRkQFn3gRp00QoXlew6vbY4EXZrlTdtJoxPl6BtD
9AIoI5Z6wsz3ksCm2T4DgPotypWnwJDl7r/NDs8mgq8BzAtiIJm31hMIioPPMN1T
42LHeAQdnn3Mg0U5E5umfa2Z56uCk6f16JRWPxd4u5AVoeXCJxX+vLEbuZj5h9/E
uc2wFbtnpSeuNRKuCf9/OmRId9dWK0Z6JmtCLLl+AiiJaqGSbllUGE9ppQanIPVd
lF+imYM0iY7dWTWUXd2IdZ43We22206mxT0BYTkoGU/sHTDuFSK/+hQ2lZU12A6O
4vjeNS+SXkerlB5q6T4iygGpckkfSwbelAp01x0yDC1K6+KiD5JXBg2Aag0DX77a
iQ9r9MLcC4E3vj0IfgcuWuMR+d5quxFsAj0Ivk7I0UdHMeWprIVSsdDT6uQ/+cLw
I+e8ngTqHQDvijqsjD3/w30XtSxTVtpIhz1uvtRiqsR7eDXBRwB53nexrdfkZPfm
94mG2GG5uK6kMrc7X7VVRncqqVdOflbLpNVPG5W2g1uAH5QE5BzM3HDC9NsztU5z
b38bcj1nPQRcMfDBCB+r0plVNUX0bDo4kuuizlKrQGBOTrsWFFcqSLjd/Y1ZSsA/
7dHj+DIQe3d+EnbkrmAae9xA2epv+wkK5B3bQPMOlqxlpdh42ZkKCzqEgh7lg+Zs
rXCgbpjmU+uBYkNj2wJ66Rjsxl+/4ZA/gqNmM0RB1rHg1fvUP5yI0EdDsjVoDPEH
E7Qar3MDyH8at4rLRfCG/SMiz14RA9thnRToJroeP2wPxr0/iZsTXZl3Ckld0XSX
mmGkdGuss/++BlXufLjxGXrnpI6MUkPE9k8YFgnPfzUdE2TpBnPkG8agV9wLbPKH
xSZMQ86JFOqvVWmsYxJ9OSi7Lt1Ef+sCv1ks8nmOh2+HixXEENLjTUitBrokLEtR
lq6wAU59SuZ0bV60SJCvcs8SHLrJukVFsQUWr40syrwJnVh+W8JA2237PLHgIf6v
nWgS6sY4xPoEJhgC6bxsoGW3CQeosWTYbUfPnuy8txwNw66RoPDBPUwxVZPeVSUi
4pVfQK/sGkI2/Ou/NVDEfP0HeP04gMpzKaYqgW+6hpYeWNtFZMkv3eXCC/j5RDNw
bJTvuGFfox8WEE/EPVytQX+fBRAAZulvdpzrTErT/41w75ey0IIWEpnmakMSx7oK
TByjA9n4IB9U9n0nX4nb7rmz3cIw1Qw5j4BNOG1/y4SxoElL1TyH6WFFZDWsHkZa
NsK82Y4hjHUfGum+dUd1EdqnNQU5/iDOTVaxhm9kQ0GhensCc3R1oPZOjmDj+7Pb
Xx0F7M4LEWZ8zma6tR9rJg7OMIyhhLlZEB5eA8w2u0jx60gIMkNc2s0BjHyytagC
TpAAxQOl7HR5CwXd5vc8fMffh9TJpfSYiZKu6GIl9K0ycqpImHAjNMIM6dtQeYzH
y1xV0namhX9xZbGZs808jzjnpeamqiOmdUUxtH+7h0NZq1/MKBGIkMH+/NKW7NPC
lki8GBbn0mCmjxHpDFDXMufG7QV5uUNlvU9viWEmQ25FoYBKcC0qfBNdFITz88eQ
swSSCMoG2Q01H/j6jn14dpfTZ6tlZAbtxYmA8QYxER189zgozK88eyEIgVSf5Ckg
1AFOGVCu29dWuYuFRU4nd28oKwXb9/Y7Imbd0KIHxLAUs3j868WX5rzlw9p56kQG
Y1Avg9CMPJ5NWVsOUb88IN9wiEtN/1vSYCeURW3F/KRnY2Bj6y35LWnv8tZsySmo
TuWyKd21RcMgsVVDc/lFOM92LRJX3ofKqg0xZrkEpX0hUjle1MHp5knkhrhBWK6/
LW4s27m8HiJIVOd88DAF16k1sBkEiQ7r879+N2QwtNCskMAMgduh3D0XDZUdwWiw
4lXt1XWZPZABjTH64/0cp+cYIUZdW8/AOlSWopcEffggbx2wSKzXA+uGlJHhiRGH
uBelw7jwrLqUY1vI0s10GoSUouBvVGwpwPvuzRkaJKw3xGLoiZJFP/Kll/fPk/sf
M4X36Po+NtksY2rihDVvhc8bxF1VyL24oCQfV2GEyACE9qbYVCF9zWjtDFbIUxD8
OhfgmCdFpiZyJ+q5kWABCxgYLNbHuo5lf+O2P1lYA5kQFxB1ILWBf/eQXrMHSfhW
tL/wyOyu36QGzpbhir2gYd/lthKK5H9QgeFW1gfCkASY0Wam7FNeNl+u3+TXgJ0n
krtcuLY4jpjg2kIuQrdvpo7G4N2isEKaxM0+4mbVQMW1XVx52gxWHiRj+iV3Sc0n
e5cw8yy7e+dAyraODuAnMNnevkogi2wqsAd0xk440u6+5I1EDvZcV3BJ8M5ZgGJO
5Apm7GXSqcScrlA0DJUlqUpWcFAOtPi/Vn+6NilKoQtrQ29MHshkkhMWVMoQT0tA
cL6THeptpG6+fIoKS4ujElQ5bCRv6lI9a8oZlN0amRWd7uTkbfnibScbqzCYySxa
FqgBHopaEETgGZuxdYL4fqOp+IK7s4RvVq7dttW4AHFLbE6HULGjcyAg/9huSI/w
LJOq5/qxpFdBxRZuZMyO8RW/mMsKATYkthPtnJlIFp5ZUXHuLJRAzPgbkyhgQ2pT
Ok0oZN9rxjN2dbDCheceUh0cJhWvtnNn33mRPoM0vZSXXB8Gd0nz7ha5f4Jc/mD4
7waLydO2tiRh/6PiDSbP/XxHx0pbwyKBvKH/fgt4fjiBLgOXLxm8nBRgUMqALNYU
pLDjXl9bZIEqAuuMcj38U09JWFz/olxKp99KN3Vr1JUODrddEVXRGhzUpNFcMQ0t
4C5FofQAtGO7JzAQOa4fQdqsgLP85YXwXXBOrHZ2OkBO3cFe3pVk+//jlEuWAx2K
PX3cqfltI8gsHMpHY+NZ2Uo+VsqKsxgeWRRF56oGi4p571hJwSSgroZzTCTstqxW
YjWi+YEE18aW3nDEwHYxMWlTLOHO6t9Dn2OwpJE5wXoC9LVxeREYJTofme+Fm93z
FPYi8yZ6Qf+PP28bxMJR565ebDjJRzhQ0aP+CfVSOCdDN5/VBpTCD7SRIhGpQrr8
zjolxfP0zNgg6tte0dkRanO1RydZ2TktThbXce2sEi6VGwDlzyyrOncJyF0edN9P
tZQdpC4ap20IMpwSTZ5gXLc3d5L4ZaDEtt+MbJbPnyZSBsGCAAiwWwCVDvvt7rLH
+7CXaJt6yUJeB+ikc3M/VZ454ixCptQeZXBMP2Rp2ej+4IvuB8yCLfNMMuhrWMLz
0kyrnBVX4QxBaBvgovobRncI/pJGyq4dKI1pRKlIX1XSs5n3+J2LE2UhIK/LtD/x
HgfLznZODOrPEZKkVapxIomlObMSM2DN3l1BQnZg/eL3MNsvbFSVf24pzAl1NZNl
qQi7gIQO+ZxY0zXAZhppRj6Z1lhW8Jc02jEPWw3flzbX8c1G/ZWtJMIFba1FWYem
lNqpqESRZ1t0S4UqoeZrnCNRCeSa2d3vtj5afq7oiVnyzt0R0phQQzScFqU+AeJu
/4rmC8wjpSrV72RyYV0yb90dNTTT2JDi9KN/ZL+uNP2Lfp75Eopx7BK0YftKB70q
QCeE5E+pW7lX4JQtL0g8GqiSgT9kZVoci7xig761nRcIFC5zCVCLpOa1HB6faV7p
TiQW1vXwcJdOneFZYGa9Y4zx15yiOCi45oY3wMzA4pLQrQeOVeXIbkWMSFwsyZwQ
Y50snCev9OjWLvU0EDbw+KI7pOvBlqdjLQrWtuhnh0QDpE7SUkFN/cwXDWkAXVBi
DjsNFbfXFNVYjQDJuwgXv1B6P/yE9MPaRURfrD/VuB5Vg4OFLSVIN7zAkbBkWzrb
Sj6evDqI3mUU9LK825uI5IW9XPP7m2EgeUYKKqHwrkXuP86f+Wuz64nLJzFlmcTY
JmKSy0KpRwoYKN+G1tpFL1rHHbLmgwdWtmyigd0EczTh1NxFaJFUffKJ0H2MjG0H
Awz8aNC+IUVEFUMR6grWKEeJhiZcJ80eauA4bU1lHtxeqjnxkbeZEXlJE9JDaDgY
bRURTTIdM31t+epu9Eyy+lgsK7BNdJprgaS15KLs3/Spg7bwBqUXNLUcV8MjZLQl
7X6no8j6Vy2mbzQUgjY8zejK67E230TlnJA7KB2b3KpQmzNSyOmTwskJW2C/dgKK
7gvBzDodwd/8gnQSBoDHVwmJEhIFVZWfJi5uB8QGRDZUQbphOBq3Fsbb+TnZw5EV
2KOPsTOdDNi67NtIZelRXdA7vnikSgVoX5P2Dr/bB6SLYJvGCEFrVwbGZN4EPAzB
hwv0LvtP1/6ZvQvrBpiTIKN5bao37FrSkR8WULv0jqNn9JWV3tlIgNAUKnStD2Nq
d15gYjPkQmpdMFB/EssOSIgC0MJoJpC8mIm6q3nk5Uryak+LgZzs1RzzOX3gHy53
3O3jgC5BtCZ4ZoB+1+RLkUqgDtEYhajp3tbvHhk6n7M3k6jRk026ooOrPRrN7vSg
WBJljLlLkJaq2C59xwUmhfx18yFHe6RAPUie1e8Uvv5vJtvs4MpTQkP5HI9WP5cr
2dRiikEXng6l3TkQg4t+JeW3hj/vsacf6yjFlbitU6PduKoBiMiLQH0vXC2m972U
7IJ898CDzNBl+JiQS2Irw3m/Vq3Q51FCFBRzToaoz74mRYlAcoytDKlq89Ng9t/r
ZsDLE4JlZFxgLF96jJ7xWAOfdBm6Zm+phgI6srCxFw3tvMsR0WFKRfsWVxyKLM+k
A3Uj8TxLisRkigf3emf+z8FVq6OdjEd3iycZWMb9G29igo4FmMtDKFFZh2HK372k
z1osEm81e871i06nI9z25iNbgg3ztA11T25SrKRbGeeESYHon+v+XWnVZrPnva4y
IxeGcjwNiBz5ahERvOgw5rHPFhXZnNiPGqT8kdPaeE+tm/8Kk9CcryTPeMo8SYsw
5obxMiQSys8ovZ3u3xZHOoGi6f9lcihsMamKLms69ILivT80wZQ3BMtY6jqbQyw6
1ybgM9oIuqxRlefJJW/h2Ul48cD2EM8CfpsQ6Hv0hgTWpTZpfFdtJK6ZSFe+G1KX
HuVVfGNwxsMrsD+BsbPsafHEpNRiv/gF3U9ZLPQqos3U/WH/ZVLKDOYJup93gxio
IWoQac7XX+TO+buJm3VWYYRVuTFgBitF4jxdiC0zJlPfwno59dU7A4OOLqSIV+kD
2bv81WfLu2ZhpgVoIia8a4hhilK01LPJNwFLIAKS63T4cMVTjB7uzIeQ5q5R9fSW
dhMKGe6PAgZdnfcC00hugbCHEwb7TNzox/87vluhDUPFA7MymzAmjeYXDKVrogor
41Wa6lNbznlZeeYD7dHnY49BFtoTC+rVuDVt1tXEwmpZ7K+fHUomKl/pIrfQltVR
mvDLqV7UeraqjHgO2sctW5MOb9/58BQMFMqqP91H5nQ7D0mlETBNeFOF8E2dHOXm
NC3a+FWkzbjVyoaH9dYqCS2AII1BLb9pEyR2fDmWVSvD07cCT97UIXDuE2rXrs7x
NOwtjvMKRLHn96S7EIpvOLdkSr9SS/4vGD0wFdTfYaVRmCFAAKxZGb4k/ug8iY+A
umrPOgyN5vilancGNFcg59lw/4syTZo0tK7bTXa9Ss1MQs/D5yNq22c//Re6ZBEi
GgGyAiJcKOEIO41QHpjM3ccHyE+Yw9dHEbtxL00+NEfJJhOns59CYknd1bfMIHr1
/Z1aPnHYQxcz3EwSq8GtYZHNR4t87glC9LqtZyjyRPXsCQlUahdFPdFHkeRfoyyG
1ZjkmdGkDJ/VTPji1x3trbqFBdXf1REzUsV3tMTeEc+e0E8yb+2lTcbHrzJWnOVh
isnet+NFvkJEuMKyB4oP+mVfYH2+usKNbKzyijxY1tCYDrh2ZSA824vCClok7/Qk
SiL87Awba2Xgtbrq3nyxFYuRsuyuP6Hr3W+N/5SIJSQscDyypzKHu2YkRNEnPlb2
R3bf68PD/loGHJ3E/RuZ5CDIAil06KOFgN39ABFLCR7BEIq9ZeEjZquv5MSNPlrF
N9hKtUrUIYFhe2SdJ1Eq5kpFjcTrU2KS+87Xk6COI4NN5DJiih2nL+/35ePspm8M
mlGl70O4USjAuCJLqikgsI6gxsDGl0IKZhO/NGfskjYNIwfWXAQwTQE/I8eTgdMe
+l6e6v3H47WhESnBBIxhudZN9U9IAUGTZHzKB4LjL7UubSUHyDRipey1wDoooaOq
fO13VKUP+bjYVMBhyYHGVOp2dG1to7sja3VCpS/Y2PrhHZUlfzCJWyBThIA7v7yQ
4d6CPaFSIlzP6ypxxOzMrwoywAJOFvjkGRn0cZFQsV2ERnUm+1VX60Yy18ujw5y+
bH2JxwvTj+UL2aq9C9SlTM0u34da/cQeJAXZcQA2C2oasi7MYuJGUOxFnX68TD4d
oAYd3RmUHwZvMA8S/ATSbtChvQsoHEKvjYOAAugeC4BjK+U3o/LdS2fA9KNKOzrY
ioccYb+cjRqNcQoC7JxABQcP/deNYDGLbNQx3TSU6vTUPuydwAPibf/qg2y0EMEp
OEki48kHgY3qwF4PK6M7LcORrwqbdata76uz2FqWEPVyJ+ZqPLgDQb0ja3npyfhq
dISTgAfxIc3ZORcwrBBb2aZ2lCLBd+H4ROC/PtrzGEYMspGTfhOCWn3TE01SWi67
E1d/FLEa1pAFkzrvFGA7DomMvQ+ScuexlFrNLSQqeoaZ2ZWBr+rhdNollZczhUS+
x0kd1AydCzf+Q6zX8nkntxCM4cYwCTk4MbTpHJ4yDO49vPclAmFMPcCy3RshfIji
yBmY0AUUycMdkJNuMpIaYKH/dFl0vh/NyZa0Avniv/F1+ya0oMOt02HqjloRYC+C
Ja/h0gWdk3Yh7QNjgWZXYCjaHPWPdzPBm3D7N3k7ZeJPEokigV8ZoqF+XRpb9V2T
oyOi/y4SEvIYXZIW75mD5qPwjaArBFM9NQ9M4n8l8U3UDRBg8bAVB3NDg4cpjjS9
yPI7kryMfyhbCD2+UycL6L2FZGVe24fJ6yV44sxcX+gIVBoeuW4yvLbME8t0N7UZ
GD7zFunof23vjr2A3ImBx/U9oZAyHi7hR/BW6oJ6rIaMF/vbx7uPyu7r7iQiz12p
U7Os3kqLf1hXbuNG4x6ZB173LlN7NIRGaX2dvZWprFrtQoyNBYiBYAeu/GupcxXk
+qGIBKbc+cR6qbrg/qYNL6OcjCeziiDtKyHzhdf99Gy/V+50TZIZQO1QVgJEOYqO
1YapZ/ZHg/gH3M4vkbkwwZcGNHFHsHMaIySt2udSuY5GSlLRP0yLEgELK58AwhMq
YrWYJzKchKgBGiuPhQT6YWJvznzmgw/2OtQcgAN+VxBT2zRzmU3OnDddOqSwWR7c
1MZT3A/swfYhUuhdR/pcOTUepm/kJliwVzb2gJ9n+Y841DvjSiMawyN+O+0ZcE2o
qQzVwPEsuoP720KCu1PkgyY36h5hxK/xWYuUaV9Wq6tvkDXpGKHX6KzK7w18RTpP
TNb+D4+iyEeBfNMj5sld2ocfXMZgTmrw/IlerIUyFKDYX2Xx/kJNMzhVYfpvLoGy
6vFLs4lfuMNUKk2WdG9AyNQRgmNduLi181tZrB4yOE7qVM1Y64oazuXuuLH3iZeL
3AXl/3IaEBKgFyQ0MyYud03OUEoyTIjY7/L9c+lft5rsws06P7zK0SJ/4CV1ehL1
wK/laoF06si01P7rKSmlBpeGhhUr9wBZduVeTnyT22HQYzp2o+UYSFCNBKExFLpT
mMnm0ryLIWhWzFX3BWu5hWmdxmBMxyBihHEO0Brcf/cGXkRxDXm8/Z0gL8rfeJ8I
4iiyWt4UHrfpsYWTlrZqVxBsYP1FaCHYqvyEfoEHta1bkHvks5oYH4QUpHQnRNsb
FmCELA450OoD/eOIYLzeHRyNUj4BioBom1Z4luCDQ0oQ2+DNcMOYVON8PnjtUokl
yR64VDCvI8FStnsO5wSfdQtZlj20oJ52BxbULMaNh4HnCj90CvXWangP0lq7ZvOP
VjZEU14vEZSm6LE6lzqgKLtH34Q94N5TGVxeNqukgDXksqZU7Xdf+CYpmA4EmOGf
LQ/YRNl5iwog/OliJAtZkMGTmYgi6+VENcb+WBYhWFbdrALcNCnguum9u6sWkxHU
ynmbrMVxtY3Ljf273UJ6PQAxFgCKzpwGXCimz6x7/qPbduDKp77thp5X1CXp5kD/
odozAhU+qZ7Yn2j8omaKqCTVU9UnuU4rlnBL7MG7/UrSoRVN8VYY5OnGVSF/e03K
ZyCILYO1dEG0HTcOomSK7InjYh7BHntwLbYTDpnf0y2lhjWHKy7p/iKcwfWbFeGg
brCBXcFKAerGFNKW3fkAZ6C1BtlI4iSGflP3nDLcUEc8Zg7HMDG4roV2SmNA5L8X
V6xbP1XFoHX5Vum7BXAen/AMmyp5rVgy4bWAAAtedvS+WhrlIZK8eAM/N1dlI9nk
MSKeP+AdLX/JGaG1TDMbA+pr016aNqN9mXfvDFAaQAGrZqUqpdpnMO4ACuTbmsDJ
DZBWwp3D8OqiYvcy6MjdVZdGxwZFqBJIASi5gBBMaPWj0lnxWzzHdulxq1peKUYz
qEIkO9PhSbs/fytmS2zpusqiDh/QEcxuVWhBHOc98Xzh+JjQSgroE7F1sgk0Z2Y3
NUdPD5FMNi+GZ4imo1aSXWGvFQK3pg1DD69bw72ttHRptXpnzNPhAf6uB5GVHE6f
1fkZ79DYo3cFTqLSG7+AhkiOxkkQy8yig98iLixmOdrtguZ65bSLjFsXt51d4xvx
SR0rTQTOQvJlwln0cnRw3uMhGsCs6wY17oJvMmWfdGCuirryi+ld2JjKQ0OrEEWR
P3qNxCsWrMnhCAvj4OxPqs1Evvg3DD2kp4lxb2srOZs4Mlj6LUgSYtboLkenj1xh
cv7/pVS997Iykes23s7CsfU8wa5/rAltMbrPS8OejJH+wB+zX+Umcz/KFaR/B2ox
+GLPw3ScoC6Ys3QW+gzYTTwwtjzh7IYDp2voh99AoxvXoahetr18D2flc3nBg4Jj
6sW3qnntg5GBHIIZ1LQolvjhOxMFZ25KsOuHXlcMQN6M3dhJF4pLYG07tuedWUdS
MkCjtCzL4KSFLCmcip2B1r0euPVns5H+bPl/LuHerbAR5BspqKLUYldtsDLNtsIa
OerbrmlrbgX3iYH1vJVIt5f9qJOD6iCcNFREfYHWOeJDH7G8tnyHkkIfhKtJgYd9
Tp0g3vVnBP87k44ZYUOD12Woe2I6diR1DzF+K7W5VohlPikgDgf9ZNT4qQGqxppz
k58UYtZ/1mi+bdDyXq59pTK1SjUOVKwR+4wv/UAWN+Zi2CelTFdEOzQzlmNwuf7E
SRDMci7C1Uc0YV+PeEF2k5nVBvPGI5T+830I8bUozPlG1MAq+YqlJnDqxig6aGDn
vFpPEgSL2oOWfz3BSlcAOdeDAravEJU6JIK2xmHWtxL4UyHDhaWHTtfHp07OyNQu
5fOYojPx5gi3v6JhqsPi89WaB40MR0tju9blzF6NlW3OLTBJA3K+HINza9VIyA79
+Ym22EpPb3IOQn6fDjQd/3O5uT0VBai2QNPelwZlS679C2pGngiJ9QSuMhbw2Apj
yCjwJRxB8RbrYoZEU4SsikCV7AqFJaUOLGQbcOa9rC0t3CUK83n1/VxdZHN4Wbdf
FEB12vdT0xXvlG8PQdGVXIsG2QuXA7a2dWs6Kj0K0/VFEwaM+5eQEpUkmnAEI0/i
WVOxRnCXo69z0Gz7aTgWF2K9j2EE3J2uxalecgWPFXqfRBTMzOxU0CYdBB8Kf/ET
syr0cSJ5lwq9D4MY2dxpS5+cdhoYdkPiTuPUTS9GYTQt/urVY+b20/EKZdJexgRe
joyuqw+/adWZujtR6x3FWgXgMxj2XLXkonAzvGY1h5VO3EIk6ow7LDUVK177mdlZ
qzVgUWc16u2CWDXUC8rcMfHWQueRjs25+JMO2QX1T+39e+sRl7oqID+BBKA5GWTw
7n4W0Ya9LHxuuKTjIXF0GNWCZNGOKHQ69NFxfXztB89VbhuItCg77p/6uXB8s1EZ
mCCdr1Uphav+gLhgXFPieo7wuJ81Kn+kTTQZr0km0Hdm58+0Si2bCDI+ZSVGCtS/
NcCueOJAGm2zT8SN1wpZmKdoi7pIhzkRR3G5ajpF355Gk/xsq9A78oitjU9rTFAc
06zW2xq8Avh69YIhKzEhfa9LzIUixP9oKG9PE7smBZHZBgf6i75OB3f31hF/Hi76
xFPHpMKGtXkMEZUobLW/pFunm9cQx8qRvUVaWErpl0hYqKxpDk9OYydXxWaWjG2M
0n6zX52DSJNSGbGgIZVD5itUUYKAK3SPM3g1+/Gh6S15KpWKimKonaZcDysY2laD
bbZdX74Nw6ESHqewOKpbSG/RErXXYbfUztXd6lE+kgP14SVHQdomzSOHG+nlOxyo
lM7PCjN2zJoGX0SARbNJngQ1d6O8eJTuZY2bL7LjkbRG4uqQs92uGjWXOK/ZKyky
rkpsuSCVUO0LcMTfcHoEDgESidQjx+DsuaqOUjiRCK7BM7q3wnojScWsuUeIgSWw
zY1UeiOT3OqUvVM423QtXC2UbduoQygfpxG+ptVxIeC0drezcQdi/ejz0hYjjssx
wJu3O7+R7FVXe/9BZh6xhEVOMT+533llL6HWu5OpyPMO12Cbz3ZDYUFpuEw/CINU
IF5MsADyT/n1NrODORcZOpNeOEfiFcs4BTtrOgJ5NEbx/JZFcDrLnXyntxN3DcOu
Jc25DHhww7rQuoPUrwunwkRYVLUCJbFT5cBlPvTTNwWe+rf4fkAMMrnbwO18m/4x
To883mGMuIdBp98nPX8EcxZxZLFYBJaR5X9bqfUW4UzrXspwai8sGoyGPlDUpa0Q
MZ/NuiL2FwGNtmmRjkvPhXGEVbVQwU0Bk4cbVUbW2ny+SkHXuErU7UVLXNoptnlf
40P4CkAo7LYVuh7Ac5xETUziPPq1Js2oSSOg8wOXo6l9F4gLPw5k+Jg29TrRidkX
i597GIpGwRLtPERbV6HKeLCPId2gsFy3t1LCJf2rCBY1+TF5Qze39gZhHwN/v2JH
yGGTZeSyHsLSsSUr8lX1e6+U5gKwvueWMTzKt/suhtrHiXG0EBGY1iLlvnD4mS3W
iH2y3x4gETjwnuRTvPplwmV2EtEjg5Ki+M4a65ll8Q24qxbVSj51tA2uhzLDBF+J
2aRwSpj5Nr7VFV6u8D5sK7oVYFBJf4IacHkeJo5qy9D/gdjAGNN2ttGfnQG9y0jP
X5Pf887k3qGUbfb2DigLjrg/24Kni4RNH68zoPEdXTrBLT4GP4JI4S3AEpg9xQQm
j/HIjNZDEL212WM4cLQN4yCMNyAvk8aKiGR1h2FOO9CGG2hg4yC7WEPpzCJHw7cQ
zhIbjz9CTMHD5RLjUubaOd7fCCxglgfb5WE13sG9qyIyKr6YtWZHO3hdRFiBX/m+
0liNhOLet9D/HIlpjOp5FA9KBe/2hdc+HquEZ4TILwHBmoTQqNEm/GkGNpDI0zeZ
21GLuJE2aknv8q4jGabVJh7WSfFIrdvt+QVgLJLgcT8eSHgibc0wcFuh23H6oO7T
yQhjPmibzJ4G0o1X0s1ztWsbRnfqKaRnB82ijZNkKbWMTvMGNDKkQudl82YMgKn+
iMc7q5u51h/6QZXZjciUtBLkZBicjqjBTALJo0fh3neacjwfgbs15Af/zux+2Y2y
5cQv9UuqV5JqVE0hEiq3myoq9cG8hASQyRR4UUZzOxkQRH6bwa35sy70vKo6bKB9
aqpGRVRYc8ck5Zi7TsyLlwnQl+X9dbaOq31BYOQPmBVlCqaX61QElMFbwh89sC94
MWytbBRpXcxoYsNo7RcmTsCg4K7Wdl5OI2fNZ3Ht+YgRzxWJuQc5xZohJjfT3gS0
O2Mo9o8hNtHU8CeLzuRriqxhL4BT2FriVvFcst31Gvx+aB8TuJlJyVFQBWfMCnr6
Qcsdywb6JO47FPMF9ep5TgNwdraYGbFuJz3bFeb8j/Tuw7BOBNZYkoIPX4dtTHso
lknugwganBUZKTuVn+pync9TbPxASEgDfwzG7L9cS6P7VuJD4CmhJZlwYIiwXsi5
PdyKJQP7meOdV80qxfnS1yIVcC8g0LCG/EIoLchjs4/LyJePJeoOezJLze1mQhBb
/cDS77RTM8jbZBzqSnNRcx6bN/9VfXwnbAP3GueubOXJi3J7WIbjdjjutrPalilw
nKvU/iT4OfgGyihY51Kp4+EBCIedXgPvL1enA8IRmkl5qTTB5EykRB6KyKg+u/nX
Skcgd0t6pWrxMHHP1eTEiu3C11X03VhthcFOPPMeJyueWZnx9K2ko9lcQxpvVzyS
8diREynvmLymqFA7392FWs3sQTFDrqUWbj7gIyyodquhVv/x5w3T8brrTbESit7r
84E0ReKvigZJP7HFPvJK1OXPtW5VFitRP7Rp6OrQE1F83nUs/CTyUug68RXjSDo0
7iXn7Kw4KFolW43BxUd32ech2gRRRVQPo+FX1VxH7wi8KlJ6REkNhdzNk03ThCaD
CJ5DjYwOY8Zgx7U+DUY0jESBnF0DXQJUh1oTXvaepu8cQ28JDD1YIxOKLZTqdN5J
V5c7q9I/orUW2GhnW+7FTRqAfCE+GZ42Kb1QZ+4qPewkX8qrFSLXTT8Si2q368Hr
N1wK3PdrC2xAtLJ7Vw0yXWEzXYe9zMTFzSRvy78a1lpmMw+ObxSwGvOnzpng2H+m
s2l4DOzuaYmgO2pBcuZotiv39IopHAK7JzhbqE/wU7gh/DlQr0nXd6W4glQ6B0if
YTCFIqv8P0ONWQjBI5V3Qif/zCGb50VcEk47QgYT7ikj32VRITu2PTtutgFZkOSy
x2oV+IXp9fZmkGWWnb4Ox6mNfzRNuqmGmHKcIINB7lO+wpGhJl98N3eOQlGMDFVq
NOhG4V9OvKc2VjvvpWcT5meSC3xeBYLUoBFCyororlggggaL2wf+OJjnYf5MxD+Y
KPqx2U9Biky9xRjaccxmA+6gymMwfe7LQ/CMgfNhUH+puT5e2ZZQY96cVhGeXwiR
vQWJV/TxRPWYcdV0zapeSwJR6G9jn2U2mKc2vKWAVeGAQO0pVBmPotz1QDFdlCIB
yncq/6HzlSCkAsHFNR1HgAHIk/SNg08u4pyX9glg0RpbptkHmUNpoevPFnXW1ctb
iSFfl4Uo/IT+k1BoO/xEIlCqP4kBIYHaagu/DQoRE70fU2/NPat0I0xsd/54P8DX
oh3wKOAqiYBcbXTUGL1RXlqSn66l7xlHKGpMJbHgPBUMBtQrLGzPjwWpAvDAypxo
wzAFPlQsZsKe28WnIzU3U2lsQO3mJgB763IFFZPFCUs8aFnWSs8VS4l3NcE/2azn
co+CXaMsVYdgwLC60u67od4x+w6wZ/c2V7Hly6A3Wx89lNZcnM8RjgUWbiY5NzkK
lHfbpPhYxJ5GR3OA9gsrLyJBtL5fp+2kegx2s3JlPmX1F9OfUW6vq2qrJhKxe8XK
jrZqO0z/w4jg/iKSWBc9+GsL+aKYK8EQ2v4EgY4AVRFkksEoopH1mrJaqkX4wruH
JAHAV/4eg1E22WjDpebF/XbI0n1rNjtCGpcjl93SjEjJdavaVy59wDcBOKwLP6Kr
1cMZhEVToXiEP9d3DnNXh4zYFr5dBQ/863DsfKj5KOYF1aVWX4sAfg2d9svsgZOE
CVfW+CEsiwWTvnV1p6j+1LYX6YUWrL3wstmAT+7zAz6Rbwi7GS6lEordgsM7X6Vw
fD5r+OO+O6Aq4rEivYPm5BUMp+NOWJS538GP0qhg737S+uiSs0xy2iN4F7L+dWzU
6qoPnrqzbIwKWGnU8KjWp32p99Fsh1Xnk1bhItg1fTsKnjrY8DQ6zOxmcWXsPe91
FRGnrlu9OwkHD7BXx+/hprikXsnl0CX3sE/8Pa0SctAd3YwijbO766h3U83Eh+Fn
FFT3lyFd76OBhKXz4K3c41tGPTmPtPtHNEAfXxv0EqJ3aUgWKf9j+ImPzGHbP8AY
blrDDHUBprM9VChCgh1q3Poo9t/o/dfDNZzKC3x2Jlb7bm5BmRm3dojbrMoHQ5i1
Ioj53d4g9+IbWYedT+OtyHMskjjGP9CwYAm6ZAe3bIF3qXoFx8OG0eRR6ygVc6Kp
IsTzcP/z4iwobP8svQ/TID2OJBsbwM7sZQu/LxTDn9M64tpmX4Zqa0ZHFfsTfk0R
xsSs+NB+bXdMySnwEbwNssfJfc01Sk1ufiKE0KqHsWcb3cNKI8gp2b/sgD2D6XuW
SgcTxVgbd95whdOB+sXDDdd3Z5BwVrog9f3hFr+Jgj9GY4NGv38r1bYD7lkiV/Fe
LstBFtvyirHKe5IxEIyFt2IAKZMddTv0iqmRBdobgmo2DRjIla/G2Lk4LPln/ikj
zxYJMAKECZy65ADb5BKuFm6p8dSDv05bBOezwcj/ghkN4svNvsAK3ohToNvmLYjB
M9/gCFs6uHZuAgIECsi2pHgFSwXMWuuSkQFizdWNPLnRIjZIAznVTF67fc7os6dv
fw4kLO2yxJn3uLbOLixoXOaLRkz3BBGjzZ25B3wMSwOqWBcvQPyJ7DilknLMExnb
9Sk95gXPCcOE+XhJgDxp5YPofHXjlRVKA3IgHMut6bAuS+6o6HTVY3X/LaeSYym/
rqMSklr1HGXtknJjKGX8D17m9FatVILNn2umLT+EDHA7K9sFypZvQjs30DQrBc6H
phmx9Xc2AW0mvp0jcSUP/rCR9R9ino8zLjAmSBZQmft3QnbiuvNqVlfdYlROmXop
mN79cExdA2OUQeRbJMdeE8hVxqazlPLZGXB8wyGfnShNK9lymN6Ei68sfSTJ1/4c
b5D6GH8rLJuZATOr99rYSh0KjJkWucvamIED/1rHMsRLswRHC31YqFaf10d+KKCe
EcBLQ9iyN8plSjk4zfF8B6IhhyngIH5Dqj5y0G7oLcKN6dld5yC5foDFpoAoE5zi
XCusuBF1OMgz0VlBR5RLm27PUXyuSBe7u7PvX7cUMzPVzCA2x8x9ajPDQLh6ao+y
LhFicphb7xme1pLgiBQj5MTp7bKpq2K4t6pv87/qfiGHahmR/5Y0qXAsscLA6dYF
ICeP1lCQEvAgH+78WeDB5KoX3izU6a8BSrhcRcxdbKMMKDkQ+Cfal9dx1cDExwET
EJe2mdrcaBQEw9S/BXcXwD7a+UnloSvaBU6APtCuSVfCsLYIFtaQRCf987UG5G/p
o/KdxSOLzl09+nvECdh75EvzBqpWr0kZXQ99ojt3MwUAkkiMT/44baSDzrDBbxz5
8NS6mCCuhh5/bxf673gpuwY0vpyNGw6THKJY46A5s25IXB/WFlaFihPda7fSXW2Q
n767WSmgCn0TfBK2U/VomXjqfsqU7KaYr1grSdNY0ysvqy5QcNEpxQb/pJWmgFNW
bLgtcYdCBGr++ojIavD6KwLb7mjFAJCNnIdkQ7ajmhkilHyJ299AibumhelV5INW
laqUNcVaWMbXnODtHE5b/5+jDx2wcmRelZuPiuSnQh8i3u238RwbESY9yKBMuBSK
+oWB8XxCB09sTVmaTfcL+5g7UDxUXBgRtEatvdMV3R+0w1KUYw7aka9e637c2fSI
odNXMNJVyYpfWZtnKwIsWTPYgT34OyxAH+ss8PyLOTYC8f+kdwlBoKDD6QNEEnxw
hjiokyNuRiobHRaUjMa8r3qNPpSjyTlt9WThA2f3bcGz/UrtbCMhwR/2B2XjHqvp
WjHebrncmce78rHLUi3r/vJEepDs9lInk4Vgg7/oD+z7/DLJPjCHEKbNntDwHHEa
RFvSCSPXz0fw2/6Kv05spl6dONtKjehNky+J2QDrtu1uH0PnXBFzeN7xY1uEHQtK
s3OD3u/cB7/NBglTh35SIRgKMDihtK6T8snQWjVFUveoZfYS4XlPp/+AGUYFnuUF
+b5XAZV/IRWOjcnMmPaCW+Hnr36p9WVoHoZc6vytLB7FpazKeGGg4iic24vFVtTp
TgAcul7bY5F8ereB0rS3Q/S4CXNo2X9g08NGC/iXHkDUChP4Onc+RiMMnhyicZvQ
+gms1+Zt3Dh6CVLjI8ttnAsdf+vAFcGULMvTqb/5fZSVA3Jt4vphRkFgG+WUjyf7
nZxZW5ryjcqSiEQ0Q+yN12ry2//X4DzRDTB8O2WKBdHxs/aMsiP/T9UaLSpSnBjs
OB1qFpIweeA59LJVLqDcMir+zLkPdRDXO8Oe/7vvT1Mfvap+eCsbiTCWA3F7mSNG
S37EwSnlwo724D1utFEvSIV/OZlK++9u07ymV5mrTAT3k1BifSlZHqLJhCh4wOjB
VB1rS+0Mg3Q9ZGJ08QUDzGS48kzTtCuCfKwOxw2pRnPGTf19UT+494zVy0TWiCJy
r6LqwPTIIRV/8zHZ/xu4bnYpFV2Go0a1Yc87sxv0cGRiZjhoe9BentpNJ+2OfXLL
b4vNNrqYPnw+TBx/iW8iJ8FlCUpRV30Kd2evWCws5XfGDx9PMfa4kisXyOPAmVk+
Sbx6Yin1NgWBIxqnQjCgzwXrtF8/MtFKLHuhHCJxrBp1c/UlLqSCGcC96WPLI+wW
y8mePVbXGslE2/DMosJ2omv4vhEOvyamfKqhvDRbQJijoyefWaZ75qe8q/KBVWut
hCuvt/IlbtksPLScJcxRHKzYWJg/DbgzV+hbP86xlZJlyJFZUfr1ceXQ0OUu+XZ/
c4zLLMJvhdC8wqECRc6I6jdoRc45wnePshKH/B+9PeLQ2sDnctSEO8hjTKVVLFF3
esqDsmrG/g3bYCMJgq+dZIEWWK4d6BkN4iov1eUGDtvmINyDdza3abRMWVcKSR5y
d6Hslo3rYlEIJkTg1DkhVcpFIUUDlxRvuf0QmI+FlQl3+GF61BNvWHcFa1m2gyOJ
oMR0eJrifRXOpQaNibJMOiOy44XUgOMOOk/dp60T8bhIdHTQ/sL2cBy0nqp6/xuM
0o+K9u1q6MsDP7CeVKQoJiU4iStsXYkEux5y949r0V67RFZlatklkRjhWPu/m3iT
7ikU7kK8ueOiFV3tkJ6YpH/pxQ+dh6aFxNe0t+PDb+RczMbDldsZGGlBOBWBFRZ4
QJ7Ox7WYU/gUUU3di2KtsjXVs2d2TPyvSzmsLbx8ByG0/3b0tsp1me8LuNaHzmG1
QTStqYh7Gyy2e2s7OO/NCmC/BUHDpPAnXm7Xfxg/MhXsxnqhB2Lim97u4OsT9bKA
PDhC/bo7ybhQeNIBjePw6+h3q+LhEXOI6hKeBv1iYPmu/+2mI28AIecKq6Y6FNNt
13QdBraJ5v07PJNm77vSGeQJObuMqChogi5aYRkcYFFZ4XVLYlNu9KcQ/ufxoe2C
2G04yZPmzZa6KdwqOMMbHDQO9kv1k4qq0f+uY3y94i0brEWMuvft+PX4gEsnRo1y
34tWRyJe1U2RYkHwDADetCxkEj3NVLG3SDaIOco2HhmZKqp024r5El7hhNKLPkdx
IJDccZB2xZDf+seYWLc1LuyjYIUOy9xv46j8Oz0Q0R7BWfGWBnX8urwJ58tSDdxD
ASSmOL9ntWf81Nmv00QUbsmv7EwJVuzKVXfaiio2DFc+pLhVWYCrbNEXpvG20Jnb
F3qCDsxkNtdz7zAYhlZ880zLjVyBiymlQKCgOxuhAurNlNgSfuHoDtx9IBicm+GH
I0BhtoslotCw8JKvPjNFKKv0LsitTiahbebIBo6X+vaHHTX3WiVtje/SwgF+6tV/
ZaJMyaEotYAABts+/pMU906cQnWlwWFX/guUN4OsqoOh3cRcZIy2eE5uO+GhsuT4
Zdfsd9jieEpJmaB860qwX4QnVKzrUkn7zRla0YqSZv6sX+GuD6hsE0HiEy6KWwdr
Un1FKCr6V1/XwaKMe1NvP2ABUpCsrt9rzOmh0r8kIow+MfYbRfQ73GjDo3Np/hex
BTd2JzRqRYHi3qfwYGnG0S3Iu1EChGJWbGZMHpZSeLT+dVbj3IeFZC4OWJoYBMlk
CRpMfPC3xNExRD5IrDPJPysB2p0HejtSdhV6VoHHwv4HMSaiZ4JFr/MjxcvkXbG3
iOGosC63JGL86tEH6j1gqnbts6D3AqeOs+A1kxytnnNUSJPmj+kXaAuPn09MSgNw
q5aK6NUp6VE+jZPsS34yhyI4Yw11M5LQ0x3525PYjtX4Az1h+mLFrZcZgmbc7N0k
kxk/tkcoJuDcxa9pi4ehCKJbBmmGNQHIzAO38jFlX2VN3z9NfwILp77DXzczUNuD
aMZtDSMFJicnDqe1D5xshsOIoyY6ijM2CVIEvwyzI1YjUkKHkG01HlMduMFESmMd
mjBPezMDhD8/mxcvR1Yyr5+NjtJp0phC/lwwbQmdPITpAHUcjgGlhURtbnwZEu0l
NzOQ5YvxufnJoQlAqHspmRsnDpPEnWT3vIBxmE1JabjahH77+BxNjl3iIdzDM7yh
Fq7HQQxAIX7crYkijCUwD4Btb3WokXBa3GQhwEuvPOf0J903NZMyhtFpkq5Zvq7x
9WLTHhNSEq8Fti116hnUb0XyhbZmqH8DK0zJU92LVbm4/NNNeS5ecO0aTXj1SFE3
5s+VqMX29XIJMD829HQrffWaPVPt1+BB8s0ud+M/nHi8D4mzaSf3f8Y/iLO1F84L
yTLr5lkhj3Ht2R0uOgVBnOcokvSDGnxZ2EIzLQvIB6iUSpWY1/r6Ua0/3coxnaac
1BZMREfgIkY3npePKnV68ewYH6ZatcXVRjn72JfG+/BSxrGlmhxu6bAw+bYaIMIJ
y8vlhCwVPOgpsI/jAC9FTiQU46FJmOKour4AytLr/49wtfXs9UgBa6C6WiPZl4qM
fZwy61oPBDpJI/CRS9gQR8fiiEbPeSW6zdoOawDnw0jVCuww8E8kk/41BJ6vqkOY
MN2jNg6/S/w/7fJgfUECXM4DzUMAvwgYz2f7wylNQsgEwOw2+hE1HOsb8qcS0bwK
CWQ+23XB1PU4HDY8KqhplyppSOw7+CNTbt/zDxtkF5p/z9xiw7t09FTaXYaxEndo
Ne0K4iqGgrSjkQF9narwVfQ4d8XsGB/T9X7Wwl77ofMifUg/GkWeCJ2WiH8p/jeK
NyjWtEf9v4WprWhy+9WkBe7vpbaJ1bSSSkU2JaR64tOGvvRud6ofFz4J2pYOVJoS
AyYZ/y09kaZzWRVr86nRBa4C8L1yHmbQrXUbvXketXzlrRlOWKBZu/Jk1+8iUg3x
tYsQfeGMbq+gL80w54CkGE8jHBqzU9jBPqGK/EdOX87DmGeKHuZfNO+BD6QtNMn3
h0XW9BsDrRP2viAG3DONAir/X6oiD9SRbDhahbbwoXkFEYZeS0jEuT8uQ9iu3uoz
Le4v7sMhlsGbu/jz6BbHf4quShcmrmaOo+rDMElTuPwEo8iMXqarMA5aTjUKToBe
y+NruT6erpAIDsekvtmEFdVn63KOffCJyhAv9/WzOKnYUFRIYe39Tl/4OjcAdklQ
ya6k3MFKWqtfdzCLu/8Sn8slhLtyOaNkJpAZujE8936UrA6kWkanZ9aB5Elz+QMm
yu9W2xT51srQ6/E+3q98t6VV5p0XYM1tkQ9xLhgfsbvQDoABSlYBZ1+dHbI1yG2A
doHQyretvSP7ScyfmNJyJhboU6ZTQ73EMuNzoFYuj2jvawB8IIovehkDGQNJxWAN
S5jfpJjxaPfQHun9asQ9Eqk8cGN/W4uunFUnpOtTQ5ciREwlZjSwJf1J06RuF33/
KgBgNUH3zGz/6EtSobQsyQEUPQQ2+X5fFOD1DLne46zPbWCI00SEw8N8Y6aMiJ0/
mYsNItSfC5c/Cgn47Ra1lCchWRJD0T3x5wY2aW1hUxcr+QOdW5vBlDvd7IPAmRUw
1gpRKggVMBjh518KvED/R55LEMqYnZXDNdHyjqnnQ7SPmtN4b+ZCV+LJxpujLvme
80wVysrjjdUtLBoN+LlALa6rXcZ4NfWsQf2TpQ05u9NuSzx6HVRzvjZs8Ja4T4IM
khYMchrFsd/SU0xupS+I3J4AULhybGvf4qkYGXMQQqszmZsOPEk5dmP4yJbSFTV2
JYYfTE53uQLIFv5rBRDsKqu5dozyFRJ9MbFBEyiSMeTSfgJvTeHdqjzGLUphfkTt
kMeSkPAhqcmkgA2DACGvXJc9UVIARK+Wr3/QJFGtUWEHoEbAHoFH0GH/b3qr5ZNE
PELHdEblJuNxNQKBOb3Fs0j3SfyU+CUZJUergsCO5qzfXu9FMxtk/1/29WL80YVV
v4zXpPbB5DDZp+XFRv09dzcD5OE74wLViXzB+o9IxE0a5BBHHslpfmj+XcuZ6P4M
YFyt1p+/iASKiU9VCJxOxD0IfgUffnLs7qtKDEHi7n6c4Z2YlKXzSy0fFoeD75Ct
LGnLOl2gp/HvPFF5Mz86/3nezRn4YLeWyRluRnnkLNKOnQ6tlXZCkobC7i6mFXaA
pKmTfz+XuzjdgqWPRVjPqk+17TJr11yaIjCUyj2NmHLV6oZcYDMrJKjh1gBdorUc
JUwlEr5KVI93RtLaqwPrYmFtrzivk9FM27tPqCFAx/FNQl/gtUoGDpr3Aa5+cIOX
ET5uBqsQEBV/A2FAChn7x0sEk2iLTxLxhow0prppnu5AYfCXaAgCrokb1zSYZdWy
3UAkw9fiPVx38mUlu8olaIs8FMXu6ZSHSazD7L8K5igcTzsDBPmkdDYGZkGhUrf6
RxqzcL7b7jGvTEhjYB4H1z9C49Wvulxv1vZAtcTz5ilBRJq7n7B0GnLo7vcgmlki
ZZOb0QudMqYdN3U8QxPjqPM5InNuhk7NWpxWtB1z4v3og3U+tOok2e7I+3Zj4O2Q
C2bkdWWO+oq5tvgfnqV/TigZMvP40PnVl7zSt0Ynf2+BdbqwotGB6cQTksDOQtHq
paUxw+iI1JefZN4segXVlY9CWA23IuxCk2WafzBy9Y3RI5Ff3GdwFedJGRiBTcJj
rNHQLhrZHAux0enyBm1DhYSInNh4uA2RoAZeahMJ1pdAtYbYZ5zEIAspIah65x2C
z7P1UkybOwSQkpvUVrBxLY0mNCZ7MsQo13znEQcASUZaRHbZ4ebcCXF7YUNIchRi
Gz6G3H0aLIQORr7yD0lL8+a5s5nGG1mgK7Mn2thpmTl7ooGOvpVcpUXlkQo2qJ8N
ErAv30daAvuFtcDbFPvZKoYuP6Q2Y2e6j5Z2QQaU4Y+cDCwTxrODaPsWE2s2lDDm
HI2HcmaYtVoBCrjZLzS05uyujk/gEoGaYOgZHZ998cC8rynuBkmgQtGFFpyOeaaI
UGFamcdWCCcuSs6FhuL9aah6oFx3DpASsmlB+N5xJszpWJbOauO72rnh+12VUM8v
fwDUozenddm3Ufp8nvq66DCS0gAUgaNIlPhJFOqxTKRhuSDsfkoFp7ZiNbJ0RDnx
Jfe4VbdsX/RejeynLWwMECgjePgJ8aMGyFPfvfIrwtbLG39a6HT8SwKifcsCr/IJ
XkmXEAPNKMlLDlCbvz6FAl9P38zGYG2uYGBHEmWBA89igyhJxNlf7tB/bh4SAZYb
83lyzKZKRgwsEK80R80mjM3X0N77xnCkxQJKJFBkNRXN923dHCUCUtxxibhbkMEl
1413WCA0FPnm14WgLxUzs/QVwFpTznLkH8H887TxypEjJ1FETzVof9UXrs5tVJMy
ijmB90MkmWYZNUZuIixvRzfzq81bETMFpfeEgEks9LyXLSFvnHkGDbwk/tuEfmo2
CIWGm06EBRNvCngeG5N8yE6FNo0qHh8GgMirNPlBCtLfjneFR+m6CLvbT5FI9jQR
RiJNxmmI+EPtz+E0uBBUQERH/B0MWBAvXICo0Z+eXIbrQWLgQAHfs6Yn3ozXRSj1
855GIVVjg3hV5z4cWV7lGhqj6ycx5zUGk0GTB3TxyX2optxt+SFm7Iwdu+Ls3gva
uyc65qPLMgS1WrcusQE5xsIfOuxEtZR0wxYqmBg/D3N6xQWbbda5VxJxjnnkQb4U
Ld1cdm+ryXr3dK7+Pm/TcXjAdlvzfgYyQJAjNzaV/9+HfgVAEeJTmWp7NAkVlkk9
EwkJMBW6oHDpIGc34OBCc36yjqR9KrSuvKWyAK4xttxvl7W2CaD0mHclVCDXb+8x
DDMl81BcC+VBJ8doaukQbvo3zHyU1aad88BFrU6wu1O1C8OxyGssro+Gv6dwsf5M
F1uW2OuzIgk+ALeuVWyq0zyc4w3NQBNGE5TygsZqw8irxuvhPNvNaIO/AuO5EvMb
01E9Wc2xJGm0zT3fBEG/kA4mkT9xoJMeQMSUeBFzZdiFDU/60tf8T89olUaOsFkO
8h+ltR17b3A79gJfBWL9wkzwShTZ9TblKbF5X4p5L/830WKQVYVaFu32ywGhx9zC
Q/0xg+E+qHU8TN74NF2vN2XNPsMRNfjai0QB1yOW8a1bBE3vQixVPBZKJ5eBCyI0
OvPZJmJ4Qbb4K19BwHXL5DE5eiykFciNC+V6w9iD9SnY8UZPG7V66H2kTmFTRQjp
QY84HVhPEeGbKZ4K5HiNJ1RXpCoJ2yDnjlY8bcip1RqTqU1uHXI10D01FJzmOVNj
cWe0oQ6v9FyGAbf7JmsiIRD8IqSTCTwfk7Htw/uW74tjv+5wu88k04RGHhSGPRPW
gyCAatgaJVhuixHYj6Jjg18TXD7XxC+BFRJFqNgo3m7uOcyur2JH2AKOk610ePFp
Y4oxsRZmDy9S6SIHsxknGt8oo7bxqjip2ivxKRumb0tQTcV/aHs07MNqx1318X0D
lsPyak78NSgwCvIq1FmNkfWDe9NXU19LCL1y+P4eAldZEgNPdT6/9mcb8GH7UGMk
kRPR4qmmLkDhD/Mdo1uBVQRugcWIsZtiCqxYtew2Mi25j+jWNxOPR64j8UhrIEHv
HtXcuLSKeNni7ctkmQr9Me1yXbG7x6Q0I2yx1ef4/JzEJLD6Vsplv+tpuL4+FuYc
rXCOdPC8hQ0DCb/+c65tPmb4dH2puJcWyiEuGZ9vH2gaeqA8hl9C3+rGwahbdmX0
QOkbU70MEpF2bFYtsvxyB5nfXniNB3r3fgIZNpfw9Wy4loF/EvLIVgyyMavZ+zld
TiOusXSV8bMkWHjYnXgA8MtEmvLldB+F2khDGRWP+0FspKPhCcOcveahe6yJwRpn
O6iZ3ESlOoe+xDn0ntjNto1FK/1gKpCLe3sZfMXbkjmQzFyQpo9WzGUjlFms5KLY
RQ3RlwqC8wOEKPR2G30p5oblTSJ3stR+xtLqfQsqqkPF8PX1I08jJ0qEvYMAa6t4
rynWbW8L4GbEmLS2bDCUkN0TJRXe67FlwcASz6ErimmKA0GLrriNomAgoZ93P3qA
iTwyOho1xmJjBgHfxzKWAAKV+GZMy1KuS79A+ynFAUfbUnrjRSgOBrmSayKOQaUC
F9bRspwrQTfuhULIZjtDhbecoB7eGE67BCPzPQTRHoWZyu9L8roNtIgfeQQ1q/P7
HLpQMs95N6c6ulHORUgz2XxbGlEpKWacVZ86u8w/EGtygR7pzRkngyOHlUgCvcmX
pzPmgZVvgXTKllAiRBu/UmZ2DW2qpNrucdfLpcU6V4VSxMIvXeALQpL8fXNgAPlt
HKuxrjX9d6srcyWR1vxH4WnFdRrUVQXmyVJ46KJIICJR+KVMo2MPQwlj05D+d57I
PQSYGwYRPGTxseSdIVEsyo/rUWTsMcbDxKDcHQ9385RjQPWNdlfdu9DOZYtv9n/y
O2sUCZGSCmH8VPT7tj8OFk5aUK8KtZQ/EttZBtnN3cC14T53dSNxhbqegPPc6U7a
icZ4UoeGc43NIb4jJyfINGB5nK28eXuzHVL2sGZKvbsnGGQO5Kl1mHVShSPap5xB
tfWtFyI3a17As2oGWu54HpDAJXw5kkfhjhWRg8Fj7HEQNxKVrrD4WCUj1ifOrFE8
IuniDfHEKG2HLoqIGLIw/hRV0FMprIbispmbNoiC11rWsU6/2/g7XgqHUO8KMPKO
e0qb+DQzty1sUQeDMZAhHX2t2COFuDO575aKcJCzg+1apJzIKjmm6S3SU8i0b7PA
M+fZWypyyWABMyNzfSXG88Iru3LBoatdTq2+9i1GZ3Wp4P0NXD64Ga5VS8KmfwfT
05eqgE9d/1C2VEbQ32kWWPUkRqrm4Sjc5ZtVhHitg0to3RemIMiim+3qNeHV0/HB
P/LTMpS+PhoS9HzAe9zq7qkR8yva0Rz282IJqKjwHWF/KT8FmdC6Y1gJQPI4yjDt
41rhQ5Ts9pvAUnTMUvwm5occdMmhZK9EpchA86gGQLNZIPK/r81CoyZPuP7o5/0j
jTTYP0U2kXQ6mXm5v4ntJArTaDI/+KBPOLb6MEavl0f59l6d5LoQbVSVHcvAxKrd
M6qyWZRCqMsbCGZFBosod1S9yFLmKQlnaiv09f5LR6IqAWWvIWeBs7A8jWYN99Dp
QZAc2ykduB7ez6swYT/oG7rImOQw5HeMrxU1qSR8le4B8fBdIEsqg6T5/0RSAjWj
FfCJ2e7AwgsrTO+uxs9tbvCXPOFzPZUb3iytHQFe/HiDW+CCXDkNwzSNEj3CqvWE
l3fnBlNTsOGamWdKMXL/l4w1u4P3uOqw/KJ79ieZIJNdGvqKlO2dgilDTasHJ0VT
IyUJiOpP61YhntVsxEtSqurChfocTHRejm0PULx2yeMUJQ+jkVoyDG49g6EIsNN5
ZD+yQ/BO3Z7LN0tElHAWh/6A/zKuveDNKhoiQRh/G9F2uReZXLA8vcFlG8gdzROc
GRcUEWAWQZSidUkm2TqB1h7XLaz10Vi23dScYHup4e640YyRMS7OLJMJ4bN0OeH9
+gQuRj9Y9CWkyNSHaL6ovBhw0p2UlUoap0XKe6E9GOrj0jjpzxYJ7Jc1UolnnTyc
QUxIVl3qZoHVD1f1oZGJUi7eWK3OjjL2dCjazhog473O2e/hodTTGyVpN6k9idVa
lq8I+1ZQqB4vJvaf3vuTwXnbtKcrABKgtiZwavLkAxM8HZQWNLnrT5WoiKWBYEwI
LwVRCfr0ujN8l0EPpmq9CqtXzF1hFTwEwDw6QFrJPrJ/gK/uSwurk6PwsgJ1/XZE
4LVIuW1T03r/DoJIKA9uFxYzctjHsgfzPFVA9MENcjdKIHvFRC4g0GPFy+kr/+12
HJdmioCQbuEHUHVde5SfXztUwOP6DgdheYOskHTXfGueRg+9kil4+p9LBdrFbYHT
DFTDCx8KGi6L11lXV5XhE9Th72oKVXvm+PKCe9lbWIOamUI3FPYGGnKB1JEdvds8
g+CYNh+Vauu9Sb4k46bnuP3Vxcrp4QtPvbFiArvbuc2RtvEGInlGrRpeJpoRBjdM
svXLvZ70uuFXSIJ5KlCV9HC16xic0yORxmNfJwoIIhvtdn/MPIt6RPM2bR+dYWWu
rL+S6DoUSIymJqYm/yipdISPNYtGC4wkImCRKs57v2xAMAoEwQMVA1WQzePqq9Iu
tJyd+R5+l9aOLBBBN9JweIXyXQA2JcB657NUxygChfYw7otGUtiW284oy25SojIG
8NoxO/+TgE5nx8NsYOwy5UYpvgHEWurXzMG7tTGRfP0eSoc7BUbmpjlgeqWLg51f
OYPeTGgbbylt8fcKaLbANDVb0oYCwlGuQa2ZJKqRAWDr9mYk6UmzGqaFWHcr9/8Z
WCPrw1GSwtPxMsoPfiwO6+NZLQKruAz4TR8EnhSBvFgEyFuHBe1Z0/Zxg34TLR/J
mYl1GEOh1eQBv07kfzbwzLoGQXaxKAiH1P3UqHaXogmE/8D7ZQQ1b6gVEmIVT8/S
Ycrib75xLUKuj2JxtE/PoT7Vdq5y+Sq+vN+aLuFrbgiucL5TXrDcqRYw5rLWRwnt
2V+FsVfJwj7LL/VHxRo+ZPWKzRK+tZgENpwjFrI3U7+lEvGINzt6vrHRXu9obNZX
LenVG6yHMnFKKwYHKTTD2xw05Ngpl8MdIux1Pxzzvb6XwpPEoOUYYbPl8E3r/18Z
n9T0l2BkWuvQuHbeiXstOJB6wlAQhDlrWim28LjXxBgtN5OMk2C3TLtwmrTo7qQa
3ZepW20GGTb78OvahaeBIGN9UNfkPWW4Or8kEzgMcxPchyoAwHGdNjwBOJ5PkFr9
4CO4VR2CleZNzvJ2GjnfaxzODDlGtrDkWJJTppJEwTFVw4Hqi8Twz1Ya20LLqYbY
bqjTBDo1lpsgjimO0ew3i+94B99MefVq01hC925bIBsT0ohZXIeFnl+/JOpx/NKm
/hgvoA5/Wz1ufGorsv5L7WNYZ7SW/78JezPWXfiW5BWTzBZVpClNytJ31PI+Wx+Y
2U3mXwPzjqhEG+LcZ6geG8UK2jC0rX7dIAQy/PjqNaGtI2YRtX5P9if/mss0Njpj
r6gpm1lEzT7WiyLA14qnGP7nTirBf1ifYFjJivwdW/7x0VwCt+7CYG66V64XMkFC
FZqiMMw0krLyfFMqAMeAFhwBDcXlnwKCWrZCQJNfUQMMcjZ8NSaZAkiZyDQe6KD1
5Fz0pxEuiOev7ZJt9ufWeIqP1zRN5XemWdk+7DN8ae/hKG4WYr7RGkR7A6lq/Dol
irmrgt12vSFBnZE33du35oqrG2Si+JACi7BcCKBrTKtAhvBxzV8YBxZ7shBYnP75
OhJGfWS3JygjHSceAKsyjzZuBWzIImXQPCqbdWHToyhN7fcSuT4S7uQIB9fqVbD/
hLfCQn4O4Piwlvo70FZM9a9DzebKDZtlGybEeiSLGqEJF7vGve6IYGuLHBHrZCIT
r3C0+Ax5QWv6s9C0ALIgIzbaERWIFyB2fmP5ui5mbq1zqXiYYESxL8RTPnnpQSV6
BuxNrAWZ74i7a0mzl4zPnDcPj+Akgo+pGix266MRLpu0Vki963v54PZpWcFcIOuG
4jYTursH0qXMfVGiz8hpLxBFM34JnQjxgMi5Ue1DJi1tVLGI6T5MH3/Nr4OViXPm
3pKO/R8ijXKTO7YiVdFwL0STX1cPmDvyWNPnxoWQssdwVoZhQlJiS9W4WL2vQ6qZ
W/m37azLNsr1ab/GnfiIrYMs4w2hs1pZ7FKNjklifVKTJbzLNpjExz4i3tdVAerF
/ErAQrq2sdXyxnMY9HYa6o0GO6IEpvpsjXDg2k09KsGnXq8IAHobQcKpfF+LwDXx
5WqRXEn/dcWzjco75HrlRRkWLOhje+4tiEga2JGuRNnzQco3qb673xGkpLsOlR7f
snTOtk/8IaP93hFp3jMb7UCRw8STMCgwT5tZi7zuPjheQK/v1uN/XtLJrhiKsozk
muf8HLwxBupAxcR73JzEx7vP+VZPycxPRvqtxj+1IiaGhKmDPMMJULRpOW6O1X7Q
bXJr95UpMXqDd0NgC7u9qo3/idWAoo1N4A59EfjaZQp2x46ZXuzdc5E2vONjCskm
NvSjzBP4tITCUt3ybflmnJV2rtQsri5IBl2JzZVSMUxDwSeOYFpfU17kmQdJBMKp
6TJ6JdZVAlKqaL2oFdqePQGiRXjPSFqHKAKfIwmyCycJGt3SEbG2Y8pLou2jhj91
xGCRU3qXjbuUxGgH1+79U7WY+yODg+ZpK3rSKEO2TdgVFCriJodC0lR67jp+RQF2
cIhlwsE5dA6iBqzXvhUzmmX+5gfhTi4CLC944nH23iNLbzKuQISbKHEpnROEnrG2
fE7UmyOyBiLLMaMlRG5G7MHZs5f5BbhChJWflluIkvJVWVj6XG6IX8UXYYn2Cukp
Tl1xYMTjfwo4Qw+pF/Ahw2c/LhKMwc8ZUP1Yks/YLWjVVU2AbG/HYyjvGAq0mwUj
U3ejHSPnCGghsgEjHKWS/NCZHVZzKQVjOOzTBz4uPfEMvCJTH1PWDdqVjOCMPuL7
MAs7lxYI7W2NEATzALwW4xYdWDFdPcGDSIjzM14H3pMtKFaoGtchVTmMIVwpdUN0
dn4MTzaGV10NTUKzuG7IOra6sCrmcpAZuotA/s4nOKNA3oAzVjGNlT4n3ElOym/f
5l/8UcBkMXmFtqP3CGtcd33+lbA1cHZPK9ch9LRN9rOY6SuT4gqiC7ZsGZ2vZaw3
mauJmVqwVBuPUz4ucpSzPD/tvIBg4bq7/B48uLjZIryeGid0LgAhC4iAUapjqUoM
GQEHLKukqNNn9SSclBk4fs3VgA0W2LwFQZowHemaXBKrXfMtUacCIqZTrwVfbJPQ
MEtCROV1IbbPhDEGm+ccR6ERiqJJAXPlYXsetzi0BbHeEjnkQCu1Vh8uJbLWFmN4
thfQwrm/AoJa6lUD2zQV2JkpTgAXAmLTr4sSDlpCKIpJ9WL6biTAXYAhWSxqSSJA
H8A+s6QPbRDdC+eX2UwJzHNawtbnfbu4PedCR9ESSZnrDICZl6B4nzyByvdKXa0Q
KRhd+QnEggfmeepA5W8lmhgRrvuYJq4DA1q0wF53JS+wQu7le09GbJ1rP8+eB43v
1WVDhdhXd5EdfBk9q8RhFPsAoFjt11kED0UOrg04Qv8k1tLNioFfuzsp6xtluAQY
3JWL0ROICgTM8FeZ7i4SYczI2IaO0CDucGpSbMK5wYDBLdnsMDk+nMtCvmPeQTZU
eTIQLCqDUq0P7OATdmLnSb/7fG7umxN+vMj5WgW5znpEsjegWUUK5NqjRlTROTOn
yNRUQo33oWiB3GJCv2Ep6AFgcUdobdcamtBbDDsxCaSfBEgbMa84M27BQ2Uv3RBh
s8FL9DtJlQM9CuLHF7OexyQHsnzu33/rzCy6Dr3RlCy4ocsCrxa7gEeiTfj/5w1m
x5JuCyRZQPJ4s4yEpTszEePdVp/QyqrPSVT6BuXg44yH3FQbQWWPyVHnnqp53Jck
szYkPkMfzDFRduN0mKirekowm6WRJJkay+ptnzYh7cG7EyflIi7WR+/pNmFk/PQ2
4DOmKnv4IQRLgj1nt8dk9y5Osszqy0ICJjloEEPuOyQMyyep/AP6zmSQXGHeK6Sz
QSUWdR7/yqL2L4Km4WDmT+cvz/3Ajyey9MdlBsUP/MaW5Q2I1ZUzuU62eikkDKgD
TsAdTzo1r1tSHwqF5ICihpOurD6npvanmLkQaMWwKlGPNrEf+YfRcWG7ckqxL4zY
ol5pQyQTp5THGZ6GeT8BDqyo9VwBbvFlzsZEe+/f5UHdp3OAnBwDwMji61H958ud
jSTMzXH37ENbrtqHMHA8+osJID9leQCkcR1QyzwcvC+C5c95o+BZO9OXRosrU1uP
Fq66BnArSeZQRBjRtONPvmwidmbH1PnwewVu7IQwSxvQKsRQjju5eHwy8sXffIZ+
/Au8qEOMS6cQc1xBaRxmR/4g2KU4XkKHipJHzPwEHsD5w357Hpe6EsHZdyYvgelv
96MpqIz+WE7gvS4/Vv1n3dbK5HBFqG4cIjSHIwMCz8GWhWYbzFyw1KEWll7A6wfS
+H3FxI11zyPb1L1OFky3Y2xlRauO7CWO4s+0Rl07UI8CqyC2xOR86JoGECHLoJQs
9vJkVCYPCOp+T80YupFS6SMaPXdR6w/iryHAX+3LYFkpRuZQYfDASDbCewPhmTyO
FDXr+4qi93OjYpjL+f9wBxsxHHbdMRJlwH5AD9UXGqyrcs8u1Au98b1+Fbw49smK
MX2gW2At3y/MSeDUEyiwLX/c4aW8xZtPCxo91/vNodn44yFXaUNfbUVPzMO1zuUi
jNRfS/0yNwcNHDWe1UWEKuofm9bmxVNrU1gjkZv/Qm4QLo7UTAcmUiR/A44WVTTH
9Jbf6+3WICYMK4+CTZALCDoeNSz37Qo92TOpA+ZbwLiso3+mS5pC3PxxasPbCKxj
46V330AYN6ZCUvewOLfr6J53EH2WGT30kkY6QsGbyNJJJJiAXmP4AzLnCvIG8Q1M
Nbm9uHRyf0me/UAiSA4PI3Fp6WcqnOflSzP3e97w/LBs/i4o9nLiPd3Ibq/9Ai8z
E5mkF5WuRZnenI5AtZnGKRP9hUDWkMxaxvFKNh10TdRuSpX302ywlnroeYsa3h+s
M4B2ZDFAVfKnWkfEK/dj3zKLaRyNWbLRU4vuh8tvhcHYOCiEJrVbX4vNBzYd52Jr
h6hpMv3Cd89TLvCfhXBoJHUapV0O8QMZXEmNibCogfBZyjgPGpUGT0BJY8sQdean
2J2QN90JjyEhElxXZc3KKanE0evaQjNg6vBehiwqKVbCmH9bZWkM+1uwb3qqfWg4
2z9dTTpS7By1MYm10ziR9UiQUZP9ImS22Qam9/zxnqlBmPsLaVoMOTiC3EBs+74c
VZN3XyESq/XIa/lxtEEQkMOsw9RqS7Bej5195F4KN9czAVsTfu/dl1KPABxTY7jW
1FEbmrrQVqLGc/K/4WyrryvUo1QAPJUPFvVmlvM4fp0bvG01PgcQkTQPqSmM2jvZ
h6DbcGMZnN6xFrmSTvxxaqxhwrTHwZ/L0/LEd941/YEmOfAQ5wGtWSvfgjbP3uES
pQ7zJdfH9aQ2GXgdo+TYQ9BaKMpdfnXe0JZrI0AC82sDnJCmOD7KGx7GWlcXgJZo
Rx8Fpj/vO6QY9yJuWPixPxBCmzUWKaBMiqr0HHUY5K1lhwmDHEA+R+O6qxauHTzI
69LdeHyM4uhmyTYK0SXkBo/eOyFAnYQ1KKGiedjoDdlIfUwtDsY2OuuM6f2CMRdG
8/HSTZlWhNYt16ZpfgV89pbUIo/wjIKiQjAas3kmv7Elq8KMtoLvBWyNQuZCbr6X
WKhR+57puQWR9gXo41D9w7D/xwIfAToaxnobd5TENSspYlfZALB6gOVvX4X7yG2o
hE4OZdBO74PrNZhU2hvRplS5hOPNdFvsyiJ3rckcdx0MweahDQ6y5c9OPfi3/EEY
kFBLSH9s5pRN5od/WHAS1KW8EOh18HuWUEFeYLw9jonA0P/njaYYSVJReetnL+Xv
cHn2F45SMpENVhW1v/fSqV0NyBmSvY86sBZe1Cc7e6HdoyJnh70wQe+Ca9JE6h+b
62hnZQaFb2jWb0uUAUyHXzo4D3LsDsoSAq9EzVoV7+NIuMqk2CU7OKWrHq8xIXrp
93O/9rup+krUiPeycsmLanXg6ok7YYmqY9BACxVmVYl9+JHyhzk8nQcaNm/akP/K
mI+vjGYxHiF2HSlmz9pi/TySEhH4d3zA3tqEpGlkezv9jfLwNL1q5lci1J3qJzMO
sh6VusOuRchAbWjzYQZws1uenPzYugY56LpwJ8/rBqa2r004ggN3yqd1vBHaOWcO
Xe5k4DmPhcbiKY3lAgiA13+Me2aV/qyBFyYb3eNa25cdwP+scNDVbpUFr/U65ydY
2nl4/1K8VqfHzEiGECxGG+dh9XTe3cZCZOz93KyU2Fi5qLL2i3wJzBvjjV4EIIkA
58SS1aLCjfXPzr9cuN77i9UV242CD0vTGjQEp+n5vG+TY4Wu0P353D/cYcigzGyV
w4XoxahtmMV9p9S8RAt+sqHHCbhIVTFuX3XFHvy48qW84rGiIIGZ9MN3tN2ZBLe0
n+gz146qYkzkXoLszlGM2sKqs9oqP8M/a8dri36GX/y0HcV4QFUsut8oo6yp8Twf
7XlqWSIULPuIj7HqbOVx96i/uZImt6+Bb5e0bpBBw9h2gF4DHKPI4ipa52UuxZ2l
voNyk53jpxVRfOmvYjBTr91Hz2UQqgiFddmau+ZV2Lx41Ap54nq020vt/Nl9Ik4T
Scn8uM57zAC5ukRtigGcPIzlohXLHzZByDs9c7WNGhwJvOMRcTnFXbl9KlM07Och
sX41OIySJznBZacUbYuQMSum0vMXc/T0kQ/yGgKbW79KC7GHpSsaCfBZd9qYdAff
tNwd3F9UGryOgoIVQqXyKOvCSnU3+jlKYvpmS/RK63Nz8j4+MikfBTiCY8p8eVFS
UmvLRc8heaKyw8quZliJjyvN/2yH/44/8NnnctyyDiAvvdi76VBzbJ/D8V2nz04+
3pWkM0I8gByuCLZDeeLyuN9cAvnd9qZlknlF6Cd47ZcZCGSv/Tdl/Ca3J9rQUtJ4
Z8uKR+Wj/whkuuC3kuzzu89/fMmXD6JXKDWCEzHPt3owUY0+wGp+KOewmuGTVb8f
ZlRdZ8KApO/PrSSQa9DSevtzXVklDht2gK6MyWxuLpkTKpuEV2QGpxNdKT1Atg4D
1kKyD5iu/ET63cw7C7qcdmoWYiN1yLdITz0R9V30efJHGWhVcpHYP+deWfEIKI6N
3DwLLQ/KlJPdTRDMDbE6WPMsf6wGrTbFH+7ywCtFxnW6VvIB66mdFRC21g2oytdp
sviOPr8iQ91Uvz8mPBYKdw1dsYEkYygw/X5qu2Lb8PSVh9AQfrKJx5lXRPA/HFZv
mNKvojqvi1roW5anofYakWEJTEjKs5BDgt27XbxajYM05rV3b26i/RtbFQZbsWc8
wZtD7HOhlqPeJA7iTJ4EnoBVcjCMuYgtSX90d2XJrojWDYmMnQWq0J0J4LDP5Sy9
tgvoke2teGnYWcWFhPAjYdbQ66Q4vGQdJa88jWniTlO9Q4K3pAdE5CxyUlBtq5NG
yi0SOGXSJztqprWjxin3BcdAYECcWvtOWcHq9pUz5o47ktS0yQSkA8e7iJDHt6YD
uh0Z4XiwTyv6/okJStucXeNk5ZP+A6yz8HHpGJdZIbBEsFseyJxb+MRp3dOj0jWl
DCNtGBnaIYTE1C4qYGbG/xXJc+jA654CqPD2wqYd6xm3b3okv+Wts3mR/PBZdM+j
3/p+hxSTMxKOJOa7HK7JmLsLlgtJJMUixO6iG6WsOR13IGoXBfHFmdN3/ERfLCEC
wXvYgtX/MYq/RoARVbKZu6XDeV8UGoHoUwZ4bJaw1gT0xUrPruAF35cryjQzSBd9
GVsz7Bk3fVw1AoCuST4JsIBJc/spNc4rPuszcbYVillquoxsNjq/atIyfgAq6P7w
vEUt5kEmusFbLAbSnqmQeYqwJU43LRvdTyVvT2jcW4Wxi9QZutlFsyn6OOd9Jnbn
KjpCOTlPKZJkQ8iMLkSrvUtp2IJK4HkOOLJbIs+5wefeRu1Kfij7Y3PZkhGHeXGb
BPQF9AUoYndozxxbvmoNkWtQ5bCTH2YbtOmaHbJSDYZ549t1/KhJSiNrRNWIVxyG
gEhCEckf3v5HS6HX0OVAsTCwPwt8oh45svmCaCS6IcgTBuyoiV0N2k7KG6iAOe4D
IdJWS68KJk2mVVuNLWZxFx33lugYplKMiHF6OF54X0g6X6xzKJQDVFmYJGMlyEs6
4OfUeVfYzsQq3SlRs6WDSaUOc4nFQwC7+sO+XY7deglcw0Bhsz1dxPh5/JD+WLDs
DTZ1x0urMNA9jXRd0Hx/UOvSCCSTM1UXb5ZGr4iyy1NWrYtmM9guW5buykGZa4Tm
SqJfQyOn8u0o4N9Cos+Hld1Ww7zijH++0vVyPhIDsmiS2T2uI2HsXcnfFdMU542S
E+f/rTZZ5ct4McGzLY9kXtiP0CDtUNFBmQCcR93tpskg+7PLljXUgssXY/+06AHV
em70ueDor3+2wbOrKs3bxIKbgA6VGXQiRge4rJqFndB9L0PlIalwru9x1uzcrk57
enLdMp1CKuREn8j7gsBXPKa9crH/x0AWYDJjF2OMTfdOMlzpIiLPsa0IrwSoYpOc
UpI1x6xSm6Iev5DlPZrE/NW6EPXNs6MaJaDvUGWoME5zsrsD93d2RlCo9G9bsKLX
i1+kM2VASzhxL6uPNHWfDAHnGt1Z7RZAYa/nkVgDeY9g9naLQG97j89Tf+ydZ7nj
C2ZFPx1TqxT/JFLYKaAw678cTWMIapZ7FRz76+YeAwHK8VXpP0lNrLIphc06BY6n
5v4C48B4GmI+bMkDo3xgSaAr1IzV/57eDXUjTjVK4mZJUUfyt4F3G6Us/KqLumNw
PUWbUdhCJ05tUxZUExgKHQfAw1VDYovFYv6nBiyBmo0cB6BtGv3IV+5xQrvYGuQo
85CrqVNUhtJ4zyhzGOoasRbv0BCWy1DbKua3RiC9nH5P8JbZBoOM/ENo8vkdc30D
1QzlyB6mFbjyFiPJytPziZG+4lSHMxXLqu+t/waif/Qi8YulcNAO5ZLN4sV+dk5k
bx1wPniIzw8oCMuFa0AcdU1FCmLFko6umEswND7leTofwo2zP3yCFXakDhC1Rrkj
XlCxD59dTO+oNkTWSogd/iVpMGCykOQCm68XSj3V1fGZdbt6Ih/Yg0J1pcrKZgQe
Kf0k8Xuei7affMmSPbcOmyG1fEahs1Tzj8U55bfNWnV3V9wFOQ38Q9C8t0gZ/a5t
IDIaQHqBmLSJHriMDj0vWL4914h/a8HIiB/d+PWSBsDBS5og6mI3vlVp99ErH3u9
CIbtdSDiT1SjhC/0HXUWLSXcSVxcY5ltQVEWCr7J1dmYMpN6gztyCTBjd8LLO2ah
6E1GMc2L/QhQhX8ugPOKvB+FuxSiA4tMIIfQ0TYg+Zfk/TfRHJuXhH/KCo3knwR1
ck34sq336PtY+4L1qMZxUgnVV46UoMdaHi0asfImn6e2Sj+sWrz2rWb8yf9cOyle
v4GhBfwn03HrrQ4DvRSINCPW6eN0UzxPzZ9SNDiB5WDNuJL7PdMq6EKrmxMGgaL0
+57E9SQYn9PaGYtuUIsIaDI2kNfdIQxNz+PIK4aflkRBJFwhFHG4HwfxYdsYyz9x
3LsP1HtL9kLd9/AES3KRlvE0h3kpOTipw98/kd3liiNGyquO80EplVa4UFHf/6P0
RjfXV0XfKJcQVvn7KsEllkOkpvoirpmN2bxtbrg5Vn2M8j0gVr+h5l5o0y/N2hNM
wpxJlsGx79PuLNTiyfb7DuNZaqyEp8eBk+4GbxbY5xL3+lPfnM2dzVsCIUMg6Fss
Lnq5kHGJ0s2USaEwxW+8EGN2Q6a7TzRAEDzvEDU9jP8LCYAxR6vghDOZvr82ZhIo
7gkNZNXLFhPOD/cm6ZnGpALC/TY3IfPlzNSQXqU2pyy7Yw2dCcqk5c4No4y9XsQv
9fEiKZYCy3KIEn/syfnGR6sX8QbrwwKExK2szYMGLKHwfWCqXhDHgq8O1AwFOaHQ
yz2CIsHKZbIZqgEQP0RMprsYfRMY70bHm/okkmNm6cIvQeMinYO+etI02I8OKiby
oa+v8NLWhzkDfZSv6w1tbBdayloZRgJ5rOSRzIHNz/HNgGPvMqUYEXEkj1pkAzf4
BtlhZvTq7X1xPdzD2CwUbQM7vfvQLmPZkdPU8dtBLSJz0/HAiIvr+tExBKzGee4V
1W2oWjnYDjX3pD78AWo+jWkXC2jVuBbZ7i/FvSmFa3cVxlIp5PTOl34RZxQauSUi
5xT0MhH6eeW0MafGMyb4XsGBz7PkWnQOmLyJKjOP16EoHFPD5jGQHROMFi+cBLo5
ncUeAHGcMvm/UV9W5w/Hj1lyR2tPScVw90NAhmEJzb27DO3YRlE8hUUdfpePkAcN
aD/ABkcsP27J3HSQYtFhAx4jF/W/gnEYFeRIHaGomChwAU15o+bNBml085IkGgp/
xtRJJw5K45S9/7mDLxKk428iY/LWFChgI6oKidRCnzDfV5gdJOxEbBbnlCkThbmd
EfCOnqWGw8N7Xh2ff1EjyylFmF/awIMIm6N2/pxxOMIg5Rh92a6/GU1JW4ctRL+M
OlJIZC1qYJ0GhcR4ebTcOC6HvN2MKq0asSzvlkKHWYji9Wy8L5fOj7JC/BILBvXT
5WHPYjAn7E4ULJPoZ9xFBzJtvW9FbSXf+HBVSJym8mzLj2qcTfor4+qCUIkptw7+
Z76A2fEWjqWIu7Sqevpb9GcpTiZIs3XzlxPnH53T3b1K72F/XWdVC3UmOHQVJ/e0
hwjT2vpWLSOaXutRsLiXoKEMaq8CSxoIIjUj8oNZWpe5lcWPQjM3JeWAUb20DwsD
zIxmHzPI/kNQHwEkmWMEcSxkzWOKn6HdWAy6iPPtd57H6GcAHlbaKJXjLdDWavyr
+0+h4hEs5fFHNBGfrfIhIFDVz1J+g008jJxYNvz2YqLVPhvQmtgU4rNvXBBzxTzW
rqOXkfbDzyoQgiV7Niscs7EuCY62zuADwPgItAJ/QfZfpYZNVkkaWj6vpit6lgiM
FVfw55DXbCzS1JhXdFuqR2c4t2G62nBz2WyEVp5mnIQc591nNW8NzD2PQZzF6dHR
oRf0dWfADgih95bcg65v/skLf7bUM+lV31Vh2emCVcWHo/FxNU9ZkThkBElHiLVp
TXQQkr4ou/MLbfGAFL/CdAfdk9wK4PcuYylUgNstXlIyijiIe1DcpyKEqF29Lqi0
zLW5s1O6JYk2mm4wEK2dtHfwZ75D5C2l7dI6hNdvYEhYYK+lJqE93l8oFlbUMZMp
NgRCyki1SVJbcIwDTHNB5TxShdTA40X2JaEvzY26fVnrDSSUa+RKCA1TlJkKwVIQ
RFkcs/OTu9Q4xF4gu0iM5Twpjl2+XSKFxkMgfYTh8l7Egamq9WJyOEYRPdQjY7JK
7jNb2CVLW8syDUqNho2uwuDZv5KuZsGb5+7VrVwXBWaGnWNc5k4c+69fh7DFfzfF
UyfA/0RG8fhC0ooY4NO8y2MGnliseDIKYnIcT7kShWmFur/hPRrDoqSfrvNSjYcw
n7M4fPbNTKbCxeJb34A0GEj03zRZBCat6dLUUwQxMqeZ0d1/BvBFcPEOnXc0FQvZ
+MJRa7G8/2Uiyk/o1dDr1WwszVsuRlyl4ZlsoVsPm5SLtbaS2zRMgH8e2hGxzZJL
NIZLg/t8hsnGY9PvE/Lnb1qogtNwZV2l+Ff+6s9B8Dzp1d8529JaJqyZLt6AXLDp
9tBKvreOhYGHwHx62TlJI+E4HCIUi+KNswoRK9+9f8dkQyIbtzAgutLwc6jqcsay
2sYVWnTVnelssBWOqbDCBqnfzhOBgry9kqwWn1E/YqW38MwoulsQet5OiO5mEEhs
irBRittDE0laIPnZeTDJUpwwqqxjEWAOZKY2CrOFWnze7eFOzbxAZCs4K06sz9UU
dX5uF2lXONVQr9w6kiGomNpao0krlT1oRDEi9X5SjsvALL5M2yN9sxA54rPIzkD9
CslSSct8bSz2K9WmO8tbcAmNkWc6Vs9HrUMYlwJ32JvVl1s32GI/+Hj/WP3LhOZj
8tNiTDNIiUjRqEFchiJ1k834nHM04T3fUT6k1aYn1odehVcqCSwVHmZj3wm8SG8S
gVnOU+rAI8e1YDteEzC1Ffz8KtGoi5r/Sz+FqhHFE/6e9z+U11OTwlQ1U3dmT8+v
yn1IsGCaotiL5iMWHaSvQLeml4WwukxzFGhDkzyDza7FpTPjiqDE9zyklXUKf01N
dCos4JXP9jP6bf2sIOYB+UBU83krDLEt3Rm/xQ2yPWbdB2HVqz7loj/WP9vHXLPp
Ni6+XeCsr1wFhVIBpsG4KuLrR+2f3P08q27gIKvUO2/Ll3rDI3R/Qy3VwTnAEd89
tqqeiW4BGJVjfbc7KAUxVRP92jJ9ugGyx99r+VHQZ2MWh5Lq+p5F7cWomnIPw2uV
35yUMOTalmtOvngzjVI3OiZCRi1eQk1aMJYgSJPFkUM8otvpw3Y8dXFP3CY/SeKI
5IqkUsyRDI49THgv10UmyK2RF/CvLQr1mNQe2FIFunF+w0/BHTEQNC/qFSYNciLy
liMO3U/XXdCJEYpoICn+3tLmQHq/viVLv5mkqzzquuLMWYJTftTHwraEP+D+ul0B
vmRuOTIdoCo/7MU+S3cwd1uY7pw/mWyxB0xlEk2eB/yNG4RuexugsLzWJ+EBivg4
m38bYQJ+XBkbjcWjySNNODwNlWdcZ5Psv0mV0Rqz9MnS2vi6U4QCVOhhs83MDdkL
tKQkgeK0xHFKkIFNkmb46UcW9RHGK5gkzOOvjrvG5VoACR2MFnc+ecKv4ZJzTUVv
kyns3KyyYTy/8oq9jud5wnPYMPP9FuQ3HmaNQw0pD9nu8AhddqX0ad1kxciIMZiA
+Pj22Yw3y4CfqM7mLnrmXMgjlFN68q/J0XpfutYBczFGeY9RqfsWnfCbA454cwo7
PwKL56hymYUwn9dO/f/PEPznfOYtg3+2cGYeeQZTSPbJ9sWE/uSnF3PKW7ssL5pA
dOV2nX5Mn4mee57jkgXePn5hxTiDkUol2o7D+J0Qi68vtZcD1ls5Ouikb5+PKczB
OHKuQ4Xdfkl9e8hZJBXOqKgdMxRLFC3JNwVK5JHcllzn3Ub4ywTIEs8Yh2x0n3WX
HmUALvNDpCOkZJtXcE80qxPIYDwDhlRS6Zfr8fjJbmnS58Q5rPy8MmwOgXqIGxK9
Rij8eK4XsP61b3WVYLY+Ls++2yZSKFycoKowCt7Eez3MoPS4TQhXZfphXuFVGoUV
+lBti1XviRAO9WdYFh/fiVyrKeZoshu8/CbIK+iuRWvK+W9KVWXvUtY91Sw3qhf8
ALfoc//K/57WCIsC034me3PZ45VPlARyjVzhDZ8vG1vN8Jauo7kO75UuBj2Wrrcm
vtqOJOZ0SI7ZuCMP2ye5LTZXstAZfebHTwGaI733JqTiyNUH4iUbV/4j5lbPkH40
wEVD+MAfVrTEhuC4HGiSGDh7veAW/ZRwH38dq0TjVswSVmZ7TMQXdmk/adDPJAbk
e9VxRNhNNUhNqk55mK3qYJiRqKsB65L6ScmJpXCuOF/GOpW1jOOgznh/dFPsRFCV
yj7HjiEu5dHCZqhO9Y0l90EkKpYM+PYSiZe7m+x/+O9o0ssGN4YbcgK05CfI43eA
3jIkTVrEf46D+Gp2Xp9LJl0n03LTKpxweBO3Uy6Ow0AohbNu1OuiTALVnunsQjcU
P2vlctmg107e+O2G5kMDeObwUg1yWISgoZHn9/BlPeMeT/Sg23xXIX7AZxNTygkt
dodkes4up9MikG8kV9t8cRt1JFXjyM6FOSG1vxhAgRxSeMJjuPZymV3OwnD1SKue
QcnbpDBxtvoOKmAhEPhpQnEe3Yufk9OZXCRpwTsj2Fk+ypISgXDMe6NA6KQXIQMj
g+Vkj77apbBA9BhNL9M5wWFciw4bGSTP1R9TbSaGfiM7W6SmEjlWS+Qopu+E0ehC
xHM9x6X6hjNt0klGNWaN7FMHSH9/oX2x/1Duq835I2OGSotgC5m0LvhsPzQpbcu/
Xgje0atYOwkX/UYFY13DS4yJb8YvBbssRXvwu0D+spZEZMRrKQ1/VfTQS108Dloy
bJ/PjVxFd4+v053PQgUwwlDuf2+zhBI24XXBTuTVAOPI7HZ1qSxn0XWtoYF25jnH
nG/iNwpoc5DdPai36BKwJ2ghxxMThLjJvkzpfWsZEXZkAKkAxIa6TU4XwAKMXg28
qJrG5908APGJyStwqFH43JU2zN5i2YdmHsaRkiR48A9jl5wl4InfWhhVAmzqjJuH
4AcgA3cij8mC3dNkznzLXtYQGOWfZaep//5G8lBObUXVKOyvJII8bmSoN2eng8bN
tNMJm7U3L8QVvB04lSn6eViFYb5VARnEnx9EdNrNgzHwHTU8/dfBIbZljspBtpmq
KzJbjXFFr39ulNXE4I0ozNRvkNg4ye47Sb+LBT+iNpipNDbaDIvt5wVMF44nuCUA
FdFWvkB0dXKc0/d8mSn4ZaOdHYoHXMGasQeufyX0lw1ZYpCZAaa3HG8nWnfeoDxG
+2gRlpPzHk+/FO9+wjmzGuNTvbpk2Kkd5Ky9RUv/jZ2kgUIsC3++rVYQ4XPgF4Xy
2SSXICiZZUGsic615gTP4WDbtYk8t/oER+loJcIsm04I+wNpr8yApzA8qJ7F7O+v
6nCqiISuNjB2NEwwI+j9cGvh/Is/O5jOGkIhZB8UfBCdqBPUhi9dQ+HuPvTCBzdg
/ydnRqhPmybH/U5dVUVuCNGblE61MCj5fL3PTiHz9aHWtTTQ1nbXVAKqf++Nqbte
0YOYKIHZtHQnCk/TULDkazambgBietEcPJqfL8fXuNTEQJRI0R9ZqQzLOjQI6Xt3
QWWi6di+vFSFZ0e/zU8fE3tfUWSOmC0eNsOX6fC/KjLdWdbKQHCo4IiZ8+Jo8bvz
fBizqM1eTVAXtuadQlpF4P9vMcrC/XlfrWjFBj2jkrtF5zMlPblETjxmqhCgcfzE
UZBZOHkBeDhF6T+A7eYQnwGLV2j2kABgxp7vHehhPIHz2VviKQ+ilIIsialo4XQH
6dnkVkieO31ttUejC1q3nq/H0MOKXgETivKN8abFCTXVLCEQdLhmdBZGYsRtPM2s
MYAYCH/kR2QszaaZEtLI976ZrC7Ip42X03UYycAWeatvk8fndLb2ETtci0tBB1ed
AGbV3QqXvpaPte2PVgmKvVn6IoDKybH4QfGwNNSO6v+3XhtHlh1+OE7DDw7NHDos
6tpBxGdTgBysyuTCrDtCHfO5OIt8cdr88Ei8C1yh2+mwkWR4sdl61nOCyjWF67s9
aVb2lgfRx6toC3z2ycfnucTAYagtxmZ6L8fnnwwRL1ztushNcjldS80cK8Ki/PJ/
ICJA6YIdGNB883P8wTyxk1hGkkKRpHQ2uT00/XC29/AjlnQbXAuVH5nZ2ZuwDnC1
gFxmt19+lT9NY18gGo9+0yiqEuMRPw2aVBu/u3e4QqqvH/LFPTW1KmshPPbMqjtE
hstxccsYEdcIR5d5ARm51aha2PCYeQFYmdAGydfaZl0IyVGDVe+KWEQ0e24yfWqU
9nC7QqlxchLdUYlm8PXyj+IhSX445AZtF3clev82MAVuRsgaSRG+NSFdn36oM+D3
LsjMVK/HpUqaOMjK/ZMxV/sT9LJS66V6N8oMlhPY0/NPW9aGQF5hXDWZ+LAVfFws
bWyVCc1hu2Te9hnxXvoiXIZXaq8U76VEYr6KeFpMs45LHH2iuvFkepCdw0cyp3jt
S6J6o7SPTxfUhJOWDRkWUVO+bN/vV3alpXpI4aeIQuZVPmC8pyfTAbdhQ0ZqrRsQ
V9rOdxrWMgWvmVQ//D0iIHNBg6pnltZbjIWrZlpQlSRyj63+FBoQryY1E1YDrGwd
Q17+pKK73KFj6DKLfTPrZ1zozVqLMnRfL8xjWKk5b4RVU6XhxwvD4M2lUoMJGFB0
wVwll9ogtZJ+Kt/N8GHCJsPg0hGz3okmyYowhW25VX57G0+V4RbpAadkky0it+65
pRnI0Ugfnte6TYA0kE39X3P1fiD+t9PAkL1pCT+k6TTrJ8xOTXj1T+ShZ9KxctR2
ps9kzjZ0r2k4UOjEJu5/ZHSMjPw8XVFnV6RIFmA0uqvP9gXX/kLi1U6wAFkhgsGu
LhlFTwJKd8ivLip0Uvp+BC7qcYtGyGVa96HTijPvR/cjY5OW9+JMpmtioagrNjUy
Z0IZR5cx1AKmM6DYo1iOCtVjjMG5rX06w+FOYFLrdKmqhc9+Im7OA4OFrXjyDzGy
Q2YZCUotz/Rabljf4NXt7v7QTv8KSR9JJNCkqBbkV5ult01VIVdmeyDczyI8V6xN
pbJDayQ5ofu80CHlY79NZrPXJxJ4lPXu3edHluNTyfA9QpLFVnSTIqo2VFA4rS48
PA/NRLRHDmGCSJoMdih+GmRwqtBFcQGuhN1ht4tbi5TzhEj1i5R48FB0X+4KN2fH
0t8bM0Ow+j4ywwWIKBOlCJCvewMwWBSgJF1wgphKKmAog65ddGCpvs1X6k2zJLn2
ST/8oIi0TBusOl0qUIF/fmhTPgPe115gHj64chjEt6ks2iiziFkAcx4ItLDqdV4J
QNq/CLI8AKih4zDUZKxIYlBGJAF26+c/X6eQIg/CsUqRGRZyq+NUw6cSW4dmWAEl
x5yUicbWDO9KPB8qTN7sbNr0w57ENd+wpz35U8nUdVLHkCJDq7uJDn5XqQmKY6tt
eCB2wfDhPAPnmXMGF2l6omuHz/QRUca0Xg5vPrmUiyj2jCebq1jYVPHXDHVHZhNX
TK/w4ZH1OaGwOzo8BmI5jFrhWr1Igw1cvonPmVAwTZo0R9iyzmv2Gmsm4XdrFxbb
Sh/PYfb8xxGizWE+LTMfb3wUZR02gGSn+Api3rrP6a9//3EYQKvj3dJ2KTBGA9zH
SlK8Wo0bZKLwAgcA3rQ+jiq2Gf4ogpYZ95LgyTzsQVqYMSsNIkEZ0PPI2qdc6v28
XYgAHt4XQMBsbFGi1Z9Vc9zlGOgEyBJIbW0VqRt71+1QouzN1+iXLZzVKzQixnRJ
UUU6myWlxJZvYrN8JeW+ydFW8BQt3VfZioZ84i+5SbOLk8u/rtYbUq3aNc5dKaOw
6EzOqSSWYFPk4AANKR2+eNBL6ovF+mCX7wEjTIhSq15Tw6Ys32ybHYF5/6LFaoVw
82Hqig7dSAGg1CcyaMuOqGyhY5IO3f6HlM3O1mrdwpjEGU1KTjJR9YuhepNvAeQz
PfqH111iBGT8ASEShRujo4d0s3LmKCvYr6SRZ0TuruLKZOdyDaYN62KVhxjADbXP
0uhkVo2F2Kl8xV6oZNiKR89SnKo/oII9Uj+gMXshkJrhzBdSP8ge3iHktCLy/f7Y
+4XpFu8nJKu77DqACiYYSgjEuyQrYeYg8A9s4FxPdBx9mKY/Eb1MA4O84UsWM89e
KIafa/WZ3E8K16rfF1zCl4sWNt2/ixrNp4O6F6DlJQMQ6N6lIWKwrF0E8N40GPS9
xM9hDZhFC5slMHLuwXAC1EvDmIQ/fTD40YxBjNED2hOme8QvJUeJXOVIneyorCDY
DsYb0c3FesCW6OS5HjHpDxIEbex2POc7/E95kZtZht3u4xNPKKw6Afb69hdyfSfi
lekdufSXcmgfMFbshLEo8hOAUQtoD5ISvFEeVNPe1CXm/NyURMsNPgXpTRJG0PhZ
6x00SiJvO8+F6K5ZLUYKrGDYUrQVcEhloxOQiwKwuiMfc51T0M7kvDr4nGvSm3P+
5pJO1QfTNnCcNKrTwNZg+ZBPFBWLZZboBw6LSqsv1xc+jMb1ToKLQDCqmL/FqaQn
E/bp4rAIinbrUPVXJpLg0ySvd+o0NbY7Is7tUvRvawTYdHfYhv90iyw2H1q79ClT
aL2sUYjqdCULnz4v+1OPVEj2ipH3zv7sZivQKOHPT+qj4Q31A3e7xCoNZv6HeTXj
he+GBmIjQrx07BAalTzkQC9RkbI/U0dBUxdcMglGsX/BAms/Aso2euF9div7CvlK
4qrxZ4i/st6slpC1uVotULeqBWT0AKOeBn0tSsUeF8K7iKquOpqq6M7JPxNE8vF0
oroxhIvbFBLxxm93on0X3nj9OoceVVlhpHIOL9FTB8N2+5B3srZNn3sXQn4Z94hl
whJrBRUvCRzyyLCr2ymRpa+DNxTRl3GQAYgJ+zqO8agWqgfj6i16ppez3aA2rvf0
CEXORASJ2rmAEep3bwARwTv2YcWell0I6OPFiW/uEvusdI5spAD3FSSB+AUNO2R5
+gClX/qZFat5MjBVoQJzgTfNcX2r+8gFgqs6hzg+ZvWwsVSChtUjtFqViNWSvuA1
X3fR81sjM+9hLjKjHERnsjLCypsjqQxOAOy0/PXVvtkKOQ5muFvuUhrWoTie1DYS
clwOz7phGJRUC2AAbWoSHD2SpRac/aiNSbYKMFpjTOY6ZJgiJULKudgo79WZdsNb
skrymynTf5L7q3+Ts/NsZNMLQQvSQH7h68c4YD3C4k3dnOk9XYkpl7wvF+JjNT/8
VREhg4Hg+Cx3StNasCw4XsRw9LObAH4lChDIAgWkl3+MokAaoCpfyLqwmtvLgQSp
N3NXFjpypprg1a73MfFdyYM98//eEvjUNP/DWD9JZWFqzBcG7SBx1JMxcG2NbT6h
FPhJJCpd2Xl/upwOyrWarn8NQtchcTAERDoOm1Ku93XsXj5XZyGeY+n/mnadqcNh
mpNyKABRE+cxZEtKpYkinFqFDDBlRPJMKkXqRVydaZ3wZKRd0Aeij54dEuPCyLyO
lUBmvfbfVDCYIbpJlFELeC8gyEMxtFlFhxSX5DFOYlfmbMUFWQQ8a3MllJzGJzDe
o59g4yKYu4xU3aKIIoHkVcrqDaYspZVhQaQPf5sk6u8FoqhpuNbl2U/UJ3etFwUB
O0b/+k7DWF7u8/DYyJ/y+XYiL/FI1mImX2gZpM2oEWTgsVekpmTCWg1bxOIQHn13
vLEAphkeYCPQsx7zsen62ZuWGKWDNfiaNmzZ4rQxxe9yh+9pcHiPljz4tQGI+nFu
qSNB525vwoEnCMuOJ1R0pNoCgEYqWijF1kvkYcU0l0QsnuUnaB0pBwJk/jCeJiFE
X/NcKP6/xLhVVICSYo315vbO5WW+Cdw9eHWBw/HEoyGp9SVVwurrlo9vo2/qZkoH
H3ZR5G9CYlKV8VUifQPp3+ZtNZYXXwQE18aHaI+xkhNzTMTSCu0tAssHfRKcPPwk
E7Car4lXg3o1WOp9kIlifX0H91cZKvyqHM2NpurIywG36+GHgtGqdenwMSPHS/4J
aqKSH6YtNe8GFjFjtfuVB83o1My2vD52ACKZdWDayurVoim1Zt7spsQju5j3aham
c1kLCB0yf/v1B2AwO9e/xAs9LHyeutTk83R4zNPvN51zIxQdaoYDv5OWCaESONNl
WF3Err8gW4FTnF8qIYLsoPnt6p+ZVm2d5OFWnWhrBV9PKt3qP1/vYY3LIlWTaow1
IvGgLkNrPpNk4jgeXDEY+zdOumPhzgC61rGIx5ivq7/ZfjMCu/ZjoHltNI8FPya/
knF/w2jIUyo57Jkat7HLktvx8VMGhi2KEEIXG432zVD1Zd4u1yQ+kYq1WAfqba8b
fb7tUXQ46BMURmK9vI2VUR4pLruVdhzwUF0Dnu5itR38KIAAjQ5LlswyA2XcStOS
HThWptlapGkBltS4feQ78Oly6a/ltuBvGyVAVDjPMuZiuq3bS42U/QYNUstotju9
6KtgjLYmVwB17QzvJfHflTKieTLATkUZ8vp6JBWeaXVcWAIDt8T2TnW69CaBUKD4
QHULJSv1nTpWE/JEVDMMqU4gNf1NIt7MJ6rbTM4OrCsRCBFZ8e2cKyetqOA6s7Og
zxDWzgV7uBLHjiVhvdpgaoxXyyuh85zvPpQL/H7mlt+xr4IwH8ZQtck8SmBC7SnS
bjvcJxaVjTqoHRajktzzrGGMx1aCtHt192+Ll0f6DY3dMp3UhwBeEYCPIPvnbUq8
GqFNpDe+mH4E7+ubIM9eHUE3OeB3BHMFqSHQDn0OGNqTz7QAZzmJjycyZygTzyFV
UCJXXu89Ai6L4HKCIH3SBOSoY53tidCZjpM4joivqZ5T3mnDjR3TPFdiqmDzx6V8
YU31P4Vlj8zymwL3VBHMaNxyGJw1ZdM4gFm0TT7iWIb08nQn1ybxGipHxO12b9+q
4AAiPTitxBsX2f+mPzxP75xxmS25GGrc/Piy6cBEkx07ifhr1NjvAyPkCCkXYLNd
VInlfLDIJWOG3bgHZOfnrXUDcu8exqMa7tbmtMM2f2yTqrHkoEaKT4XHbhkNEv63
DOct6vF96nyTSO+Rwf3KRaljYtooA6Aiwb8oc9vFxl/1j9O5cVKuzanZ/KFmRSOt
QhK+Gscdw+yCQAwinKT9x79ZFnHD0bGKPnuxb1EajF/KJlzf0hrGPAFQDXxSB+Fs
+nMX1dINHeUOVdKjmGPQRX7tq7fOeO4VUt0PmFNIJ3lwru96mnyK24ONe6ZL5DH7
NgLZ9Ck1b5VCmIvGEhJ3Rw6zEkLScNx3svBVnCH16DumWbIOFkdR8a5PfX0GRfh2
mN3ECjIw78U2t8ltOW9LsPTVylyFgsTYsO3TSfDJ4+/ct9PkONvMSJ93J0W+oNvG
oebqdt1yW4DXRLQzKwNroLcPpi9V/g4lsj/b2R30iZX+Oy3jzXrMHF4lHwWKWvzr
iYkZnc1QdUPuh7RV9il9A3zEsG8FteaamPhwedODPyQd74N0wcd0RqTU4dD9TM9Y
x1nUbYouCa5UXNrW68qJt2GaSrw/1WFoq0cRWm/gABzq0hJQEFg+sbcoh00AOJm2
rfCl9Z7bD+sPc8kywVxPJQkPE5zbB4Wu8ggb07EhHNQU1s754nZHkVvpK0H0crCR
/TkGDqv/a7jsAln5f/N53rUlOeoX3SaujVBHqgvGfiJUaL6+J0DZEFRpt5G+ypDn
2gNymmWcnzIB3ZUfY6dyFVUO6qh+6tdCTXlfRh31M27cudQpyVLVfHBHXzG19Cf5
M2bh6F/e9D+DGZoeeWcwMLKKQzF9X8z2s6vMnUT6kA+onQEGILtgUTm00krHnFU4
F5hntcUOeYIi0vLvZQcWG5OwmChsEOL755qVnOXi/kKI46/HmdPdWfvgwY+kmBtk
gvr6b0SXYF9GK8Sa7YPKS5LtS5vxJB9t1s1UREbe8qMY88QnJIdD14vKxzk4jw3i
ICc7X2d+FBxHh1vAROmIxMTDEdm6jIjIMKU3V9IiLF5/1RZa9Yaxv/LQoffh+kug
XZwTzIdT/nRKkl/pwtMRKXEQUbC+yKGyt1it8oLTKMGSB85INDQ9LDVxxrus2wYN
sfivefgYySOVW9ZdPJ3o85IsBJIF5+RBzGwBZ1B9p8jtDbq0+pV29zWvYcCH/B/1
ZszEGReU3P8b6IrXDGhrbvhnnKeZebHHX+AoBcLQ1kxxQVRvPmoc0DdV7C2tueX1
tSScmJukaeqGdfgTujoOGBh57IQRy1Ukrp/0VcRt+DV22ehQu7uV9k1dilYzZ294
GQd/Js2na2wjMkaCIn3KV1xmRBhopsuNHq1JtRLIdUqvJYfMwF7QusKiLM0sh/Ol
qL7hrzmJssGs/eZ3cMGH6N76beNqGrrotznmpXqAdIlBDN0jawAT1+JIsk6WXHac
IEQU4T6eJtTi25EJrZjPm0hplZ7wSQ2cjEHfKuqzLvY27NvoFbyKF55iPOjBY+q/
MS+0Z5EkOxgYKvNmcJRoaD99wijFgPDG2rRrTsBxW9ZLmoYraH9agF0Kyx6LjSLa
/fWBSCWGRtwqDdDg1tv0SeNxvpPq0Wd1mx8XxUQ+ZnujRXsxnLRx/1S4E7em7iAi
zZfy5Pm5xW162keqY4hllfw/gYvp7aBy4KrnJpoixSxgvSEd6WtYb+jb+KDXTjTS
SC9a9tzuhls1LIa99GOglR1t1i7LnLcXT/YdwqA/21JOvYzrMX5NbsVzNSb95WXu
2sdR6eD6ZOgzmvnZ4LSSbjk6X+lpyGvfuR5Ng0sQygzTR0F7GmnQBPBuEU3iS5Q0
ScjhU1qz+jIPVobOAAmZpgSbizk6joFswpRaZcZvnETNUUkljywmrUnEaLfcrWzo
TFKV5EpBPuYPGy9gWiuJ+9Rsg2op9dC3c3VFf415CTgMOzQ2HkyjlnHD83IqNYSw
CpFsUkexGAF7aLzS9eiYNEXJWxFOqsvR/siw5Ut0N7TgIEBiaYzsTe0TovOk5LgC
fAiCsoeUg9D1KcAJoJltA9ZsF23ArOxpbdTMzn1J+ta+YGUGAR3gLekJigBvNWDV
37XFuesLD4XFHopLvQVylydpwwVtGGDhwp8Xfyzk4GluA+lZADKyxtPFYaLchP5h
mrH6PJndVxJKintUauZCcKUcEsdFqGN21qcQPOqg9P6gQJ6kDi9kPCuOIBJS0MUD
iJlCGDXyvD4TV0i7qD+L6s9zdNYnceydkoVnDhVqhTwZ0AiLdN3SkAdW2v0yAlBL
MyqII8tU4HROfJaz0yJe+8TOHUXuo3ok96906OLix+3BWvPUyxl56nr/WZqwm/kb
R3gYGKnja5JQaRC0QwmT5tYftuuWFCZA3SlN5LEHvuq/oU9g1fvaIMOqvlj25Eyh
FJp8WPgB2HYfEok728TnoDnchkKVBCCSUwKxrCPz4m6dlN0BN4ABZ8eFY2UkxXMO
MxvYzRC/Q3PBRzq5rA2RtKutO4uqhy5NU8zHF4Zr5KPE0UvSkvBK9nXGQ0DYzYNO
/KswIXrc/84hn4MIGJ8dcidC83lcRU7tvtqrAzt5v9ORw3PZtq1EhvuHABMJ+DtT
YuV0Bbw3CIhMSpAXxPi+BVGhNv55FBxyqTnj5/23rbfCbyu1K1ueMPag35ydSYj7
shwsp5Alh/sWgr3dTHsiF9DLpvwDHOOL1oFxOw7fL0Jh0VCoywUygGbajdPcGLVZ
Jr9EHJU6Q1ubEqbiWGc47HBdrIZGyAAyB6GNZv2gfEyArOPu+0Qfjx4tqPh79Twm
qSymfmg8HHDl1VqQ086u6eOqtkSPA81gRLJZ3CRA+fzJgyZ5d55poT3NYoYcTu3E
Nu4b8REtJfg6wR5YbElegUqXOnUQJJX+xA4PM6Bq6x9s9H+eD5SL198ALRfpJXLd
ecvTOtdt1JSEoZRKKwlU5D+polUEMxhA6T627ulGezZh0mYXGkarLk6OKLOU/Vyr
+ldSxV8QiQ33BWqyN7HSlZHb0TXzzwjCpIvLDMHXMqlQ02PdoHTUr9hp3yEFcQvs
hnrpVgrM+VuShTOb52Swcj7o8Z5NQhk5U54DDwXMBN8k6JPyl1Cifnn3UYespH5r
s49Zi2IbYOIh1xvD/V+zzLO/AyU5TmpPyFEROD9ka2ADkdd6GrLC3VFWfvMYKJrL
8Ltlywl7CwNSZ/yKaYbpo1UxUHWn01qvYAHFFHml3Br+lj8d/BWp3fy7Ua9RZJTZ
nUlEHq3Hivn9h9/4NauvgmzICzguMbEAOUvaOJ/dDcIvyDghVZPWpRbGq32XTA0R
IHASKcLcjX2TdkaBhCyCtn06tNNRPCz+lImT/0pQGB3Txh7vC+Z1kgUVMk0qfuSs
nAn6Q7JDa5iK3dYFouKOSYFWcfivEIEwhlDsrFkmArmAr+3mFP8DNNS6u/0b0CNe
yX79FGKJp7NPDJ+goKLucsJSpJhFCM5BD/myL6mkrWPlqjRfSGKVBXxp+YWj25id
Pj6LVeBbTlSTzrL1hAkTbHZ8MIurBzmUUgBXdTDmQKIzZeiTgvciThSwPZtVrnrB
N2TJOjyxIOHToGeDheNLAMnb9NHooSO47avhYdDBpbw8hvJpwZtxN83dHB2VcH1L
OtJ3iDMSEwfoj8mzW5QGoIvB6zmKIBetzrTmjZsh9a3N2L1zmHyxWdN4rzO89CWw
khGngLTIkKT9JeVyylJ2q3SK/N4gb/gXdBiPKgLIc8yAu5bLJWPqHmTSX0DoSsKs
ADVfXt5IeRgUNvTLTyUrj5r23E+TkR24OvQaJR4UVqxvRf8NNyY50L8E2UC7gDYa
tQelY/XJsY1P6rBVjeuq2i6EdT06N5u1GvucJRKb0ve1RxJ0k5LZfqiodzTeV6xj
n77YKDMGQ+78JWeZj54cg6UfkvBC6lnT3jkaircjyX8vx8LLz5fqagv50XXtgXbu
CUdUGLH4/dRaybcKJjj61wxoZ8c7InYBdY9QgjnhnB8ewWs3krk3OQYPbeynoY3v
8f4PBOphJKKVHz+cnHAHfrqAHvADUiEIbSrwBQaIPI8+rX7sA3gpb2gLz+RUttsr
VHduVKJsor53eiwXCmbwpN2znLRJX/60InWJgCs/6BfTST7Eb6IP7cnorSLu8ZjC
QSYWwKB/YZpwHlgEnmJT00j8IqQR20b/9pWtXCUdOb0x0WFvP1o3gkSnQlOPSqur
srGqFtqSxnYa3mkBI7Qk7pWPhcB9d00W1K45D1Fi2q24y0RKF5tVorkW0Mom0oO0
+m6LZiW/reidNWt1XOtEAbfMFwo3bfrJ3qJPMwvDAXXhSquzHfEbMTM1oA+qlxiC
9KGbxX1IGjCQeQJ1PP6O9agDo3QoGOjvO7FGHKovygNSteKLymZFk2IpmHZBiMwX
0MgNkfdMKVRLkWktMfp0vNXshVvnQAMjCyZygl77vLcYAqMYzzO98JY5U+3e7yvN
eA2WiPkBh7K9XmL4Mk7AydP95wAP9dw7gCKXFDvK8ZhzK9OxKRPPCxuMgKk51rM5
zoicKzm2eJeL1ZPoL267jPX8XCL2GJnDpQtMHljScimabKKYE5psi5BYul9ymCOY
hk8qCU7VlV6DgyGATTi3So/tTX+XeRCDL2J7NAcY7YLROakGZALFIpnyo8JWv807
cNLJuETmJpECjW/d04j7WcLl49rjvVEMiYAz5Uw/6tpyMSZbuPc8eCNZKfpfHeux
69i8PRaJUsU7NB3LfAt+pYxnEIYqmYC1ato9O66SXKeB1inyKUlG4ycfoSy6PpMi
OD5BK80Kww1x+MOe/9wu+3Up/Tv8gxiZqh8GYr04xMX1ld9ux/JtsFP/73qletr4
w6IVflIxc0Ip5bD69F9aRGa+jAF3O4JPNoeBbB3MssgrN3031FAL6TluGsAHVkS8
8yhwst4BD7dmWuJPaKuMF+CgC8tA8fIPOjju2ks/i1s6KIEjSBmesajOAqeu51xL
cnn7yCI06ihlf8uczGk9mLqi3N6qhXUGgaWeZQgo3F9dAi9qUMqpFrO4/GVOz/Rk
iaycOTIjNdDqI+1zP0sDt0c7jN+LpNeFeaxolC1rD9oaLFOK0QuhGjcYREFv07j/
iwQjwJOPvWxTq7qsajTbRKNn+1ivtdbxByCR8QkwHKj1wIjChH1ujg/3bTo497D3
gyxzj25NVm77x4KMYYZS5uOC8sfHJdWRFz6ckLHnSQM2kHmaApctC9HKour1xjX9
DnLI3/ssgwfcbq+0cRmG8NszAzacsWyvrfAJ8FbPkWT1EKmSFFXsB8r5aie14acy
4U/iKGe0rmE/lICQRLoQuX6ol/gzIeAx9ovKCXhNUCj6kiIaaJ7gJoH4mIJ+bYWp
VVTdn5AirXGEjMR6WQB8Z8+Q8QaBDKaeeZVMr3HqLXl7lZUDTcgdXDJzccZJp6hb
d/x24zFOdSYigww11I5Ys+3EvpjxmWSn/geAMhKjr8E0fQpfldHQcBNaA0IVbWco
wax4HSpE5JsG3tL2jgsTyYAEZWoC+kzRT3Q6qQldeBNBme7z1YY/SXNi/VuFY+aR
9cPbYXTdvCTaGYI4lDs9LzcqZvaRpvNPzGs8liNHsKW+Io3bk/eK7wQBxZoN6/c9
25bgOjWgy80PPcZq4HaVsSXNAvGZFvbKJ/Z8W2yreYLqFF5CioN6V9taVblQsstf
kbr/zOQVKOSyxwKuIE6Hmejf1G8cbiCPDQE9XeZMud9NntxnOhOTvbnn8BSDLnts
VyE/JqbIYNzhOM/ZHvwLHynd1KCFUZs7H076zIvwkgx0t2AHf7LMs8ikZHKdbc6J
+x4FTXNv8LnBDPfdPdo0j2FAUSba38/tjiySWAPWTAmxI5KGy0pZ5L1XGibxbGyB
JL6tIMkupvDRNxRDEhFHCen0NkBfbct/8/OJHBvkAssQMjM8TOnl9oisaOoQfA+Z
JISqm3XB4T/F1K87lW/uzpczlr24NxTCUT8tROy6LxAK3usO+CORIRDcndDGOL/V
D1sn/460g6CPibsABAhgFGVM+fOGMVRrhRLy9zFr4GGYJktUNBTuSMlkPYCZbJeo
Cwpeb8SWjEthzLs1xAfXztwl8kZcUwizH99+eFt6FCmlEhlwH8jBZxUzLXOXLSFJ
7XA8vqun8Xvf5ouSRX8oXmD5FhnpKrkvZgLSGBvKW+p1EaapzrCADyF0d3Aoh4aX
/hxY4K3dDdJL+2IAa5NulbjfVrZ5ZVvhbNYUHOw2mf5P/RrECH8uDCq8Zzru4zm1
6WK3OE6NNaKc1a+Udb7GsKAJoU8vg0c3ZrHq3+HusFlnv3+SI8PQHQKzzU6UcsUY
cgU+jOEpl89K7L9vKlzQNUWpoNajcygjsw2iLilZiDn5yxCFp9r3Ueu8ok0mKBuu
MuMi0DO0NYlBBT/wSwwFGD2Ue0zONiPR1cdtz/X7wBRIAI7KkHIvr0lQcEEmJj45
M05ankZbUnHe1TPeYUmkzSvCfbgFmSVCbNIS9cuPdE/s30m5LDFFZ72oy8ln8Zsp
msjS9SvTGCCh8cJsOafbuC1GwpnZ0UEEYBi0aglObM8oGoHXY/Ui5J+9GqjfD6kF
uUXN8CcLawYEJ5fuSaDhVtqgdzF6uMpQu2r1Xny0mT97XD9wFdt7PYst4Bdbj7tO
mxec+PRXvufoIr9lm3xparptC4KMvzQf6igFSb8Xpxu9B6c3qKOulr/GwfO2Xdqj
ISJiKc131KDRDZRljdhv7e9anWSzQxW/wEzQBtnoejEWPNWymD/9kwFjfSFU4Tz8
FzfYBwTen6AS7i0GNtC8bpDjAViWIPOeyhzq9ffzDRdKI0jUZ5Tb0btIxfBnGBR9
ZaTpY4+epYgn15PSuNpKsj3t7JnVqjGVUPtnzB3+AEyUeXs9WzKmqVzkCkGQa7s2
/cIjoGEx50y+/vz9E3TI4vHcJ65tCeAR+4goAhdDv0/N0Vt1Z19L/KbFkFFi2nQO
MOWE+8OmSUBF7L13vfly7P3BJv+gYCMw8GFoOmsidviAw51YooWQZ8T0nw229DiM
U3OSCG+rkJGxKYep1qYaXIL6CeWj0I8xegHKKb+oGhniUEUeFeMvMO/g1oN56/s3
WzCRIQ01abzv840MMo7SAqx7ArzurfiVU0jO/911s0wQvkz52aHFkq6mNryJGMCb
rUFRT7jYhJtOkY/nhE0w42xzdBPTQCQsoEdMzhNcwGtXRwRza1PXj0IfLAnkBJyX
4nHvbK56UkXtcDuMjdQ/4Dkxy8HGbUY0q29Sz8Mq59jQhfe3DAVnIdSi/6mkd7g0
5KbYkW/rRKfZtlzmCa4iXZeCU8PnQJ2fbunCP6RLVfAW66SlyVOnO2LwuyZgRWCl
r+Tk2bpy/vpf7/h6J7gYiX5sck+Yxf/8NoZtVOZVci6fxI5o0ByTRMpx+4EUisbP
glfe4agNWeXxyuA9VcldeLcy0wk1I29y6xOtCUnQAuq93YeXLuIrtzqzao6adwzV
pm6L9dpEacZIF+95pvo+qj37u6MhO52tihbibOYp7hbtZ4Wo5QySk0ia8mqK/ZPv
KgUKY3thyekFcVDz+Xx2pwBEpYumdYeMoB1re3uZl3ntcuJP+Ds9TjLYGuGfyvQt
AE88yt+UIkaP9vfeYMlkNWzFsp7Uq34KHQHBEVAbUIaLZmAfFJxYtjSESFzlDsVa
bY6B57T7mGJyi5aRDCkwOCaslBi8/oc4j98XfdmuUmv/chkIWyk30zPz/ILhC8gA
xE/wX6nXSB3kpAfK+yxmAszrA1LOteeMP3NFdFcncLh0tLwWgd/c2KMYWqW1KCPJ
OT0DUOhVi0kNmXdfZGM+xE85tnU+Acct/V13P0ABrxCr88prJHm7FRveb9Fox2CT
REQJIyHHZyqAMCahrPwv6m8KvVrdSfLCfTqCjbEhBm1tAOdQwBdieHx0toEm/Rah
MOc2thZcGW5s5eGEy6+T2GRbK2EbW3DrXFixmpyTZoGFpgEsT/YgiHLMcCfS/aRv
qDmM6+kGy5Eofl84OBswW+GuEhivT5Gg0m+wr4sPzRHNGilguyNGMe/ZEkdyrdtF
e6C7tKuyqMYOp/eTaW1pIoZQYZQkyTSyKMURcQ7r5EiGLgXoMahXmGa2GG8Q01Gq
itEnB2aFR/mmCYOKNAueevXgHMIkPtwB73iJfLPQfDCyBEG9c55gFso6i+ffM9/h
K+mFnl0a+vUocnsjvF3Ssj+giWnP+djMtuDAs0KY2tMQftvkIWUZYlhvoQJJG18r
m1cbcuTGUtT89hj9++L3ysVeFiAiUxpnX3W5EyQogCqMoBbKII6zOZPD20zqFDjQ
F16uf4buiT6B9jNTbvZ/GCH+djOE6PXbMCFf5V1Pw1jGLAPkg88WztOJ2qCiAzZO
W6/VbZz3JadNoTovmVvCH0CeedQOHTAhaMMFaIeFnNOVCPzws89GkA3eUTvRhI+X
iTehWcxccUQkv6OojrVUxEpiF2pbYNfCPu6uAiZ9YBaWWQoso9dTS757AlPQKwyL
HX1c8RAGOT/MVTJYq3q6wWGs4/2t9b3WcRzEJWuYQ23+BhNDrlmhDHd8q6xIYMSH
SobIsfyd9aFImCqKNkz6yRSSm8Ztb2XPp3WL9n0110dLFRzQvt+r7BqzqYHWAo7p
9xeIACR8E4ZmSERrCG+OEO1sibu3keTe+ZpAYkcY6OAbocHxOMRZWa1+8xnN99vK
8IdsBLrTpAisV/GlccA5l1e+CN2D8kQxaVEe+Ijj6lN9mCsVK0Y+i8XtIah6Gb0z
uFRuWeIGccYDr29MSp8WKQqvDu9JiqRQmSL82xHvMuzd0eMHq46XpzBTwzDKdYqc
vDOPka11w6/japmRi5YSniVrfbwnbPmKGi1+ZIAMnD8Z0TQqhvAQXB0zmCqUUMlV
ZWYwnQUSc5T5pUPX42MbhcwRAFQ8COWPrY6wv2cZSogpaNt53XMnBnQqPlAxTQbf
uQySyCLe9AkBKK2+hZs8eOr3LzZUu6bQa/E9OowBSy78LV1yvpIyZP8JeIBCLnSW
6uGn28DvV58sYfd/PrVrpG50kaziHth7cJCwrDgF0knQITutJ0dRHNWv7+fJr2ho
9f8IkUrG084nEN5r8gHtVhLX09OycTzxbsqDFn/A66t6FUMTWrCU5rG7TsQFrWlR
CygSKzz8XQ8aWNBaLkLDCJti9yA5QxTzFbCj9FsyELFWf+jA4ZTu3mmZy2vJjo0b
eBq987Jk3C7SYG4cHqrb7fJtbClMFi9VIIc1zYhgUX/x4enrN3Nh2wKTp0sI0i07
g2gO84JLrqvnth2OpflBXJsoEdKRbYdEPThlkvliQA3cL/gbMg/W9bpWngdxJYF9
lkEYju0usX2vijBqH+ixJ12jicCMIV4QmWcC7RvLhL/mff1pGNbqOuxfR+wPgtTV
2GTsHI4DlnIhc+AJ/OfugS4pK+hkJ6ExaTMP6NVWuPNvLo02bbwPWmpfXji0nRoA
VXXrSSwzGlDcY8dKM3v9muX/pnQnk5E+D5yN8Qukv1fGDtayrBQBwMCzy5CjnX6W
aobw8OBO6olqrTy2i4DVo8gJRSTV/bp/mJXPlh0aEttjX1DiQA2OGXaKOXkLIJMM
ZTJ1odcTEOX3hvX+937Jlw8qid6WgYMkKUI0Ih5DXaD/X/f7H45lHpmtNglZXulJ
SpLvuSWksZ4kOtvzEEq068MgEeMLJywx7NNNmnyIcGxTJ9VgAJDLy5HiUQi3smqh
2PLi+RnoKlBFbFwfFjEanAZMVvnHFMGMnJz6agbzkvcZ+GOiBaJMm/y31zKpusVT
mlz7uuYiIQ+Fbv3he/YhkOCbi0YHYQOHKBrFRZlSkbC0bi0N8ZveKtUe77cOO2h/
DLJ2IBLf+H9x+CuAhGGvCgmiD/QehUWZzuxqvxnf/r1ksdekJHbg7O+AoANDspYR
goEPqNGgY6qh7g2ekjH4VYsCl8tdIP8M8HLbTHDSaJtji5RVQkGUcnobRSj8P+wz
h+AEQLcKm6nC7OwYJfAougb+lvhx8+MOWvd6MgP7tnYvhxnpiGXEM3ZV7onX9SrI
QC+KRjgLbpoyQ6p1BRk65JRHrtuAjSE8VU2Zo5h/JBZUPnuB5Wl4JgXS1FjZeF8i
JIu03FeFJl/DAXbl2l2MeHWY5BjI/yaXiaA8+AzPYiIUxIwNTn7ZpuM8kmJQv1w/
GYio5610FA8q+RJufj0iYOUneVct63YcG7Utm8X11dvIzxwSFaIWNY92TSzvVIup
pcmqXt4M0nuamARScHu43ja8dP3HVVOWoYIbbmwC/FVAlPyCNYMu8QC/rHui6c5n
Q1UqelHzvdmCpEEk8QXJTyIMYM3fS71h1Vsxy82LxOrrqhTEPRvwWvXau8c421pU
5cRHsw5gHAxrtdMDnRE1BGuTo+cjWogYu2gbgIfvDPYUIsm9xq9LgpFzs7RNw4Lr
siC+m6OPwsK353gKT1ZfTqtVkCKt5CH3022F6DdYS/NWUsuslrCgmJ2EmqBciZsQ
mxu4Td8rwISVPamYzHRQctJM0HxRm3p8GHmp5WUaFNoXfu/4+1ykcvydI7Rm/MSq
Z2tXSQIg/Lvg1B6qZScl2+7NvZ2EF6akg/NzqxcmKPddKidkBbsUcRhm3TlfrgSc
h2QrR/YHSAiz0eJw8k1cYauZcYcOZ3IMOhYR6H9yvFd9tyMb6wZjB6AlN/xeuIfu
MKsQxbgui5s3JrDtJHeSFaZPlq5JTEtJiMFF70oXR570Q9W0SCZR0zxl66Um84Iv
sl6p4CO+nnWT829TAjrWZclDsGsW/AviqWwg+0wrDfcob2Ftln63nLbjAe6eGv5P
qfgeSnv6sO4/1WFa4MgXW8j5721kynMYuV12ygAh9ym5spDwUjl5NDdske+0Ongg
T9Lggu3mWa8ynvOBYRDPrZ1pnIE7ATDDFrY2NCSi5aIGDj4LEL/SExXQiHjz/N1w
50GADao3kxw1lQz9pfq6OsD14ZnAGH/diSfXYw3+VnDskczXNixo0p9h69HL7OzP
HwBnXTpsOmCnyHfrX5qFYdwsZAZeqWuKXq1gsjzYIJkGuvOVBE17DN16mJkQOaUN
Qo4lVMzOeklhx9QzHIvy+3R4tugquohphlpLp5CdVgzNfU+hr4e7yWZ9JmeycVqi
5CPbM54BjD/5pRetrN734ThXOkKunqVzOWbtP1GPbJAY903Twz64xJbLpCsOlpdx
19OI06dUhx+XP1Y7MpMkoYPFqdEX+/f+FGMYMQvAlEgeo5JbEe8libZPpgEprKs6
rvduOsycdGHABRH93sGhBEoE5dgbIfXuMChDTqt6jIQqfQuKr4MVC5OUSqiATpdN
kOTG+SG83BzbKemuTVpVwj88E+LqXj3CLbTLwppHswINvoW8Q6yPzg+PnK/nDqj4
/VMiPMYPdCF5YVL+o4L+Fhd8OFu6vktPbsWXAf88HtRM6uHVvRouGuMfvDCKlS0m
MPImgXumE5mFGveYDdmzXIY5NDgSKTwfvsIYD88U0FlXT5OhJQ4rB2coDMWAcbOh
XKQpVBc5klhUWCtYkymG+neaG5VP/8qIs9OmBZUmk1JXg9Zv15yUjwv5JJH4alms
u4PpCv5Fe3pT0Va8CHJaVgfkEjNHG2ENPeQW+3nBGJp+Gre8EbBq7/qm+/TGhJ+A
214bDUpVDsgrPPE3/KFbS0lc1c1Xo2NxrbzbvN/6pA5lCs5B+BEhfFpPGCT6gPJV
QnB8w6TbGIH25EkMmY4xSPQvpEBH0WBk1EjQJ9tvKWe6oY1KhloZze0D04wRJy6T
ruk9chRK2NyOwonpbwZoplFbdlQ12yVqpCGdktNWnNSQbsqTGO41nxmIV2UQ6Oj0
NBiwt6UWYSRKoTKSXHs9HxdYFIntpgM5NRbzi65ZiC6qo5mEECmCW/hxMbSVYrZD
3WfM/wLqDhdytHK/PWKbLO12+HPiQQKlC3w9ko1lfuM440OJgfRTLdb8V2dzEWDL
8JEMUf+mOFMYnVVr8D02cW7ML43/FKyABtq0pa+On5xY/hJHPzCWns0phK5EfQva
ElpOtZ9BbvZOcqz34x8dF+C5QaD+Ng5W1UdAR71IQw+GK8YtloO5OXK01GKNetsz
2as1dkBYpuKlt/TiPuO7aJ6zmhrYDCSt7RkOrzY8nptsvHJm9YU7rx5Xdgb6xIfG
26DrcykgGz7eAO2kDQjCgI0m8dX3Xmep1UgDFzNF6OmzOeN6k78u1ELLj2v+NOFL
7I4i5+RlQV+7x3ttR6g9JY+MGqJdiQzwFf/iAagWP4jvGBCMnDewQM5WKH5uIxLs
E+/pVfXGrEDWvGjBVKPtpJftwodINpw11pXRxn5bgAQmZg5BVMAqvUOVVKxPEAFz
qWZk74opohvfkRreGll74qs2ZeFHLw1lASvMUUMar6Vt0CIpvnxLwdBHD+EHicCw
p1ptYWmfXR7ekpMkuzd0hpaESB8eUt3xebdaAZx4Mrf30LaOSpDa6mj0E9KYUs8O
qFK5Ep6yJ/OBo1TpxQ1sGjgke7uF2E6V9t3RAV/FNSPs5z4Ki3XzVihoLUXu9Zrn
VsJBNS4JF9XF+OA18QIlUAS/DaR7PFM2VmmwVqk/UYU4eyMx70yjkDjpw5wEsmNG
JTKwCyNdX4D5kqRVN2819BZHyEpv/1gD38x22vvHE9QeV+da953gXSBvxmZHG3Jw
GzaWANiZLTPEfN8HACbLA/1YBGMKhEWNB4mnty6HDHFdX3JpACYl1/VwuFg9sOVb
s5br2iQTyE+oAIaXQDYjn318aHz/jiIEhd8G32d3HpV7BxMP6JwlwsvvLCBddKtD
Yk93K1C4TzdDIrKpCVtfZJsCY+p8YEKULqOiFu6phoDOGNvcXth858SodgTNRycf
RaCcQCplPTKq9mWdJ9N1eIQG0bpebgj/SvcK1AZNcKxJrAYvq/JVVyKQFdHKt+NY
vg4rJZLcbEDuiKIZgNugeOgGALJv4RolLtdF0ZaGENIFUQp0XF9HXQNMmPcKkAf3
plNoNg5UZjYVnzsJK7ZWIAitIOGLCgRd5ZBl4/0bQ531OgDZ0jkg0bTrNkp9Dhku
Dx5L1jrA8cX5i2CLoHNFfMKNIZRWeI/931REqwCAv7DIRRPelyj30YdSbzxSyYql
9CMW/k5H5wDSmdHatI5tcukbwEEoQ7YEUjA4oTuD7Rj9cUgcAje7UmLS9t6mpk+8
fEJuXug6ReAhQVKNbY6Va7YHvEiwzg88xdFlQvqIU13FaZiC2YrtjQ4otoFc+kT6
XJKiVbgBqCphTAlfuqHcO4OK+Z+g5Qz+hz/CcDSpfYSjldy1HSixPuKnMmLvxwkS
uFv5H0Mf4EpSoeojOQguXYmodXiiVK23r5bAvbrh902IofbsYi863M+o2FGT5as6
IJCWNlubk2wntpBt6zqUCOqq6IQT5ZlmETyOdNQ3fnOiTCjuSJZhO/zQktB4a7JC
tP2zMGSI676CkNIL7POezcjHDnuaeVZI6bMrxpfyQmn+WfaRHwFYiuowq4gYlM4X
jegPHM2+GHXuIw1/DLyt5KeDi2hJGDdHXvZo9OjStSt/0mm78hABt+YjFzDeyv+t
iPnPRWnHLu3Spg6h4T/zi138bwk5Kc/RujK2yLvdZxfmPyLdyJxzGthN6oUQAojP
mSlI9IZ3gSbv7q6++8lECtewOokYSbYn1pOWyRHGa6sq3wlggBdVEiy5YT9vxj51
98nWZ6PLhtuI+py+d8ubXiSqYEdR9i98tAvTryXbmoqnMfLvwpGZkUmu13PBlyoK
rZBkZxv/pPJX5G4KdMVLeAOBqC0rja/Vfd2hStwYnd2dDw2+IP8awRTVM3W2JeRn
E/Br8ZAjcv29iajqkiT7St7Y++BqB6octV2kF9C3onEwVLd4wlO1Kz/bj2bUvZQl
y50GCkaU78+3jXgnQF6+4pILWonZCNuz97I9NmmWxsDFPvyQqhWysa0ozrtxJGDo
ThGJ4c+5CgtkCYumGzz0wBbZsnkKczZw8Dcj3mj8Y1jLRL5d99LSxccDtJR5j/nL
QXbniqZcPAaRwULO8Wot7Pgs9kQRTm8aJCHecg56z5dL338dDv365EpHlKzX7R1f
1yhMqzYED4NYviwJM32A3caK7K7pyjq/J9ahrihR+FRts5iDrW5W6wsw2uVEVn7W
pRjrCArXWTGio+HqXNBl2CyPsWOxI8fN6TGrPHoR8geO/03ttRu/DZXKsPXn4Ioe
oz8EwyG38MXwjHVLP6XCgNgemmeSRLarmCxvn8jVM7CqYevSIBATAH1UYPVsrUUQ
rFMzCi/OeiOpRpsPRibjZys8RaItSVGMK6KelZnMs+0OODKfqBOsnUijGo0Xj/jB
6ATQLrqRNvpiYdlQieuXZmkYVYBxggwpDXkmQ5Wiuw3K2LbKHlCWfhdM85AuZze9
UQSJ7kNrdmmIJ6+ZijwHCNDxA+jOHXKq6RZajBG17pzDFu1BAt4RC1hMbVRRNob5
Bui4zCQmNIootFekfuUjsIRQPeJDSiku4zSig3ex6BymY1wZgEn8/N5ReW2Nvvsp
cDJ8ZB9m6Qgoy+dsDGRhPSrHYAJKB5ciaAbCChPC+ar41NrVIml7Od+q4D8PnYks
AeP0kEgkyLzGOgUX+L12qPbFmilxZghr7qAjSm8rkC1cXA2ycZ25KpvcE2e5YJnp
5YMaSNv5iyIU0d6j5NPVkNVKm4Y3ibpV+lg/lrELWSIalNqhxtJaUJl1IXtONR7P
e+0RZ4oqzKcEbUE9k7Y0m7KNL1vsZplaPXJFdfJ9B1uV1CUuznKQEfFOd+G2urhS
fV2ZWECW0bG/SzEXNr/IaJMQ6DQOepEU0jSOPwTUHUBnQc5+8b8xBsb/gSLYVD6S
e8EnIZzCycneIRxPBDT4YnX4ejnwNxiKewSVq3CcDoIdE5/Jycm1DQNSCgbLqyFc
eT74+noTio9qQwMdQmDr9yJJ4uz/cmYBEJLLM4ilHgjvYwYC1JxrhJ22P0U9Vifh
gWzO+lKvQ+6RDE0xMD4vnWpik3mjcm5mxuDp/4XA8gb20NvnSy7e8EeJ9Kj5R4jk
2X9d1fhoquShJ5ZaFZJBx9/UT8wvAJG0dZZ1deBeQlH2GJng1xB1DpJIQ+QfCcdq
CSX+v/mkoUi6l9Hl0KZBu88v7n4d64e0wF9TW0GtZqmUBoYB2zZypQ85tn1Pacna
Yv6DBhK6JStGfZrwd8iinJc6i82RxpTY0lGIpNwN98ImQ5kFwh6sfHj3Qza2/VsO
X3UT0px961XD2rjGkID1LGZyTAdatSvaCYaPqEI+rbltkEFRHeTZ+9Q9Dpu/cc1D
6bdjvEuFq0ZXAELY3OArKjQjR97yukY7e2ygxXMtyTqOGRkw7Jy2b96sZEYSe5d7
vhNKvtDpBETWnG3xJkXYhhymLQmWhM/IWmiPagcysDh1hEc80qck/Z7GacY8JlW/
XFmWZpk7YCPJ/Y193OAX/Bu7EVsoEnCuF9tTm0dJi9LFeKqnzPNHmwFStpfBEMPe
Qyp7Ml5pqwVAwd/kf0FVl/OGVaJR6JcO12Clx5/GLzZUPcsbPt+ZBBXr6Ih9ko13
U3wzkm3ZUDjhmHKbkABaNf7Pf2/vZnrpP/i+EvKqlx+7fVVBNX4CwEAqhyBfmTnE
zPLDlLOKDXi9hi2v3/umHHDV2C/FdXslpKkUr5hvyJdhDpKQwFBkqQpYWz6huCh1
K1Coud/sX1oM9IlLRZar8hIIBsrxQU/UGwQnzynRp/iu/Tq7HxYUcNKwY9ksDb3a
bRBFn03ZYeLC7Oi2trbfOC8f9Hn2J+Rrm4FFdVrIUvh7P5L7XhJZUZCbJ3S3+Abe
GBvL44Upn06wqmh/YsRwEhDo7hNbz2iKDDHR2u1Idq98VPX/tdltJXbna8h0cRFy
AGMWS3BV3nfERAiiVW5hXs/oJCDOmovHoIEup5uTFOU8cy7NQdpe47e+efJstV3H
+5ZypxnAhWM9TOFlXu4+waiyzzYiBnPtv7T6oSl3JMvRad2+QHEqSBtfdIN67BoH
RZP9h9WRmlFRawh6CTMugTSQM/LxcGKMyboA7nr9++U/wwaXSvFCN73Ppqqr2FCp
XTqUc81oWa2kciLY4kTyg8qsDTHEi89nFz1uSsxi9uG9k1R/Heg09i9ApcgzgLpy
R5wclixsxG6hQo0imzDJ4b6qYk1McuKvLX4adHxu3IbGMi2OibNTvRnBSDqjz3hm
zOWpQHsB85EHgeYh3LYQlRhFD96Q5dLACwSnsivPj7clIQP/hzklSC5eZ3Aeu/aZ
EiDV2zXoUwYldD00x8Crd2h+RMW/OWaFMSINyCxNONFrxDcxKFuMJmQEMp52ALCW
7kVWfcfVnjCrj6Et4FC+UwzLgLdkaQR8rO29xmjw80CGv435KYqrOh/laFDE1nEE
jgD0NoyG6eACsmeui6/3yQnjfkHHK3wIfrZFu1VHG7kKaqxQA/0qv+ZbsKJb+JVo
XWEhm1ajM/0t7IgeAzAbRtUgZYDnBHeu1I3JTJu5ru02zaSNt8/fsthiYv5Iwf+0
HXXIeT9Y++e8zluUnoBfie9KdElE8citmDzTi3BCDz1kOep5Bs3r6aWMH6f46HAm
K82BMYyqNvnpwAD6RBH1QGLe2GolR6qqaz5hTVuvA6CWszayRwHH12YONFGR4TUc
Nsz+tm3pcKY9c29/T5Skv4OBD6OyaRsRIgCsGFhqP1Bu9wkgK/VBzVpdW1CkiEC7
wY0YeG9aE/l9jRNLDBTU9q2AepgyStUQXZSKb05CgyHbcn4mEl/XBjEBAKPuqMZJ
+udZj95pl8ppqcY17/fK4Wa33nsueXG1zoFrhxk5InCIC5Ij1uaOLPP9bA5+EzSw
Z4PKNQ/MCKMcDPIwzXrx7gdutqnWKpF6eFxyH7BNMb8T9SpJS1b57G2o7LMUNkxV
G/agpToC8qkPnE2f0oQmpdu2CXxm3doXS8IJltu1woKNo1KKU9d1yvoplT1wIf3j
utr1WCSBPeoZqk2Wv4aUcZdR9qdLfhdPQIEhhRNvVyzhOHon5s/xHKAkQOusKde/
hTz9na9p4u0tbIWNLEJNvkv6AdMoQvvRLpIJgf07RHQxyFZxleeRbchmos9/OrMo
KMTZs6kUJse4Us25o/oC83+oWhjp++9T/gZ/PEbgd3gZufp74sb2bc4KPPaYYbjD
b32M04kEXIkseFsjjbF+j6qbonJkpXKGscShsHQqVkXlhhmPPKFNu3HK4KrjIYCl
psP9q5NkEZYrhaZkm6WKzDRMZ4Ct1EQJ2nRKw9f4+9epI/KEA3USkvHeMZn8nWSM
Sh4ncC6Bv3jqYELk1TK4LKWwAINszsuoeN4St2dfb993qBHtutO5MzvapDszcExP
44skGEtSSONaf41tMgEP8FsHLhpwaqzWqwW1cyp2C8AOxvUqXh00jcspIG+1gxwt
1JqpMYgSvMDZu/eOhawuopRaiZ51ifS3z0p+cfTHrdWBJnLl6iRx+A96+pCVrGll
ji9NsQKN8flAZkNXHInfywXgKphbZQjWcDH/V1o36L2rKYXUZm/gfwttDE+pwqNo
Wzj9AFfsOj3pL8DLQRKmqpNh6xjX8Ynz1jUp5hY0vcF0pPOe0GP/NBFzJi5smNRz
dwnNe83rxG4CIW/SpD6tzAztwsKoLC6dnQjpVPyVxr4j0g+w7hC5RzsfRH1hxyMw
W0njszJDcOXNCh952AQZVigW/OcBPJMMgm2piOMHMqjak0uttdUHZDieXhBlprXG
UyAfSqmSiw/398G/u8nLcnjtBcN6cDLv2h5sV14IFP5DlJT5RhtM5Wgnzr+w/R1G
fv5t3DSl3qJuiKU30IZuaqQAGGfW7s6KaEnV1fpA5eOO4zHwmDOfHReq17emEsS2
j/MY/cYObJYKVNDYzPTmYTKhCd1NgnSM/wd7btF89dGU4SkSDBovWC0y9AWe9TzI
2VmtOt5PGV3zgQtcJI54seGYx9nz8UEzDGOi9zKlC0j5KMme2Hp15h5kGmH7xeUV
ckRv4fsFwh0fknGOxR0DesbyKSGReM9d5dNwX04U5oXNjO3Uw+gr85e4E55KBAta
hVDrojEBeRZuts1EckTXzFCaMv5bIkBZ1ZtDvETvlBps1TFHtE8/ory82pssT+xP
ELL8iZviZVPUyC/dYlFTFankFGzanHijqW9yzHfgZw/4b9dxpQnIqsM+vPjmd+MU
U5sNQGWyI0Kv5iS9j/Ell0a0no/sRST9cvAQ540042t1wHJYL35w2vua5eXV38bV
CGsVDdoZCb0CGgrlK6jy0BqHvu621Vf6zKulJ0GkYz8QXI3UkYK/badSSOtygDC4
kD+a6WOzsuX91JbGa/DopYIDyk5N5isK9y16WidK2voIBJ584s5iG/reqb3RbnBQ
xochRMHCOc5HUbuwrMw+GsGwbO3NYbzkx/uBL/mxbgccg/RjwEetjqIzZBiNoCbF
ZxpZMWzduD6IOfH0s4JbpBw2n1ZXXjwgVSp+Bsd0Wa/Zpy5ZLS12VsZoF+ABg0X2
Iz0Qt6OB5zY0AGou/ukOugFnlJ3cFbJZRu/NQa0DQjUAqrojNHyP8R38VAWTgKs2
BrwyBrBdZ+hKQQsV4JtzZul0UNAcub4pPBoPmzOtCiE7YwL+UnYzzjEY6WzN16aL
sP3CIhhbmcDx4aNae00NnVKgaGfjhe008np5spxY4v1L0QyGKNmvVeEaNRALGDw0
3iVIGk9liH+edd0oBCwrwrWbzsOTnp05q6ayCoXHrB2tBQfgndTk5lkf60gCKvTL
njoglUWVUTbwMAT1fgYEYPMUJF5Kde8DTFn5CY+msQYVHJghgJmuCvlGiIOvWHS5
bSIcWRFM1wpIs5vIIbvUNdgHLULHyj3klaQgy/AyBxxI2Suw3BjsHNTBfNq0NvMv
nMSYSQp+kSKvTA7my1biAh7/gXIg2xdpNLUEQNsG5/lxWrt7DUWoVaPKJLXEGDQ6
CJ8UawuqtU06NO0K5cFgV9qCneiq3Kz4zfG8EiRuLjQGMqZ0zR36aGxZYAewy3GO
eWdu+umo8PyXyBdj1h/6HWCqJHHgwPyXbcoYMkhUkdQv4fZrI6H0nYJpO/PANoiT
QljDIXWoiAVUcpzRQw8O65+9z/Ip0ds1o21blSBWI6m/ugzUXgaBbeh9vDAiT8v7
ozraDbclTNlQdvgyMU2/4OH7Qi4XpFXWJkWr2q97at4YDVdZz63fnhexRoYIkE05
k5KM+/zAaehzEIYGfDL1kZw5bQXvzyjrLscdOU50JaiHAo0jPvwQN1J52N/lvcBf
HeotG0dZGGRLgkISjN0I48GNbv3+A615Z9A0YB3S6/nJVp78X7kC6tihANGQYXyy
GAyxBPf5DS9NIq7PO8py+yulVpCjVGwPOH5RZc0WBfAq49wHr+PySAKwOFaHmsSM
I5BFGVWnWDdPwd02r4gn3wVVOE0Bru/8d/MCpJo5oAEmONoDSp1iXNHMNLtl5FaX
pUOpc+xfzgqAsQF7kLwlspTrEH+fknlYhLf/rmcRrXkdSEfdfzloRkbQycYU3XTn
sY4DTD+feEhpqK15PAgPmIPYfKbK+6M8pdOwWllF1VqSyYOSPjsg1nHoHGwOxXIb
oRj3Yi/E2EC4F0PHZgvPLhB0qVGX06onbsC4OavgZf4r4rmAlBwOlXthQlLHaGFL
V7z2GOICpJJH40KV6XdVvLqdgVcrFrWUvXz6Vh7nPZoCUhiFhmu5w9KgkAgK9HAH
JLj1bpuizwH8w0PKolG9UAxZDTslR706zoqehZwmdNx+Mgc4JKnlgNSlj46jKnay
KI4VEqvpgN2WJaKw95ekHobejSsS7QDa62dEffzkA+VqIF8n3nAxej6jOYBYtvhx
yH0vVbeauUNH9tpecF26tyUh8hc/XpCGN3CbvAfeXLCpTOMupGpCEkuY/XOYiy4t
y3QjT4jWpHIOcUeA/2IJZCkeX4hgaDsLPUCW62Hw2ZSU2Xiw7iJm9JrALdA4Oy0A
8tEn5XBer/BJbI+bPiHl54jsJYLPkhkDQ1EKNW5ONn6Dc6ozxoMMruhw6HbdJiuP
YJXN9VMEBonuRtbeesJrvlajHo2lkZJ45d0yrojwzJDojD8RyglKnAXlibEs/4C1
vpKcwnyIkhoBpUUbL33V76n1+wf717ktyASSpF91fcUi7D0RF6aWdpYNfFlW1usf
JQtehA0iLjzNz2GvtkElkNtCXG7j/IKbvgEwNHE5U5vsitIM2sexGSesL8LZNjxd
RjcBZN+6B7YOHSgDX94FaGvgZnxvi2Klvk6Dx5ifgPEzAPmJpt2eoniIaiRZMX2Y
dYzPNyJ1qa/FeERy6k8+DQmDhbfJkhyDTof+IjsG5Cmb0FREwzKjWjmy4juBT6KV
/kaTz/QxqzMP88IATSQTUB/b3f4taNZWJ4ySYX6UvYAj3P5OOQkimbQnFigp172d
wpJ4n12iq3/AF60LjIf77MrUCb6Y7CX/EcfPv73k98EQ+1zwDqc1f/oPgMfmU+j/
frrsTZ7qQiIpfSn7hsQbxsRa4eBnZi+CS3W+4uPKkGQ1SIu5VEerVqsVzr9gJ0wT
jvrVXP8eQgMvoX+RL8uIDLTNSu9PQEOkBw3hqM6BA0l5me8DR4pKpnIrAPOqLAN4
HBelNalnZ2IKHA25M2yi6Io5nK1PZt35pWARox5FLyUIY/TRlTF4408lPUa6DlHl
qPw9J/zgF+Mj619fmY7DikmaqJIqaC16nAmM1dMvZoDvmUOhDoW2T/DedYycTSxs
fKcG7hEWReXriztKV1pIPx1sKdSBAaxC6krED/uMepBnGFFUq39ri48mYyf9hdzJ
4dr6xoGASHFTGrdTdS4FljzISRUFghBf2v7h3ETBJekoktdtGTMYCZGtAhgTUBNQ
rMuDSKSARPHCeIbCqbedTw654YWrVTWrMOKeedrKYAtNJcuTATB0ZOcFRPct35aj
hXY2CmwHNX55kLFE/QWlytNusJZnOnAWetMqOfyPTa5QWgWHp+uHVidselPHVLjW
1+Rqw7v6xsxV9J72p4JR6KNmKb4fDjnRWhfRzlAnwE5dXZ/J7/L0JTPxpVTsCj/I
DlfskpUa6k3TyqmDlpIy4RsglAnQxhd8LTKMwCP/7vqWsCDmQTbcYurc5tu+kZTq
kveR2jv4zSNygAjTkQ1vcQS4jjCDG92R8cu538bkg5JnZMCKtA8ltxxihPySf+ES
C0a2yneDBieJXRNyHuUbsBsfdTN5N8hFrtvAJyOzrhaqhwkNW3G0M9bZwaL25mph
jMKq9rN42G7ulI++MUkMYSusG24rnb15dbHa0d+ePMZeOKK4ExXwbN9VMgJO9Xr8
08G6iGcptngmP2sWzvqJS4V96IgfJO+t/oB9tgI8mb5Ks459Zw1osbGeSLjhaJLY
xdU0B48CMDfSmm4Rs681gXrj0VsJc6UYke4Gq1/eNubc4Bpok7eMId/TRXZ4HU2D
EGLo1oMSXeyH/PiCjfUa+Ws12nfmUYbbFkuPNyg++Aso67QFVFIAQ8QuX4TUENcv
AorPRqijK/ucdQWwKTFzLEMx70UTP3GmKc2bPL93ZZqFbKWXf9UzlODrPEVjyNm2
rZ51s1jlZGnhaM9VgJmoBcdzQI9g+/8gRTu7A4XhaBwsmdcYSpwItr51LVLFM7jk
cXSGntzSZ0OLfX1ud1+9vh+b19dl/CoQLFLMQRw+RvpHRPGahzDjl0NBj8jA7j1w
Ed2vMygBZyUXCMzGGJ1by8eemwO1ezUSmi9Xiu9m6UK2n3VIPefIqCXPdMpRn6Z4
tXFTRstYBVpjpQauwy8/RBgGj+1fN3utXdZrk7gTsmb2h811r8qMdBDX4/4zBuDp
4Hb0tftP9bBnMHE9dxFaYOc61Vu3LNFVeo1yY+X1j7Ppe5/Yno74rI2FLSIhE4l8
eBSrSCjDKCsDUJIjEimqkwC6izjjQL+M1QH1p0r1ukIaGtNS+FnbF6q4VyZ7JD2L
AxMi7Jrjjct2cG7c3kDDyjxSPi66hbEMlzJp04Ya7ZwKI/i1cPBf4g8URkp5n70C
9IckGWdfkxZD+LHhE4db1WEcRs+WMfBY9PHqdH3C2wqyQmgwpZIIxpvRnC9evNvE
Ma1zcr/qnag3IndeXb5rOjG2vPoGTzXaYh3HnmtcEHPjQOT2/unALUbfzuiZJibl
6ynhkGJhBDgVCm73F7AQWsg0vvdM2CRlUJJ+barJ2rPm+I+WZTM0c078pu1VGF/B
JERMl5qv0b8c4rs9FzqaTe7gpubh27Si3/2lESKCucI5tgJG0xUhLALmXRga4njf
sHhn65cF9j5157JYrUsZQZurbCKJT2mNUAWu8YUqhQq4syVEu9w0xzV6MPnFyPj2
8cCQbcdwyKyoB4vEIl8E+kaXei7lmHLboiASh8fMwSUOH/tej6d9V2HZcqTiqfiq
T2LwcqeloL+dq0jpOU2HM99V3bqWXP40VpEDiwSTYaPFjmak9EdzMgpm2C26p+dM
5BSK6vkMDgY2+sL/WbGPM5Ep6stEJ1efAhpeTHGrpPulgcnKXVlVGGCXKhrce++q
u9q51YqXOXjk/45nCymNx6wOwenXCIt63wIZbOACTFeuGz9XCoZ9HMdpdBpbGy3q
gkXbdbc6viDna4l9Kqmg0+42z2zvMWgVWBUuo/yeSlNjfzQRRqq0uqIGrelpk0sT
ucjvzjv1yy//OU74vqakmi7qk7JBY+2Tu8JSS6SpNPYfJu5l5QATvP0DxGgz0x47
0wutzQPkwi8rHs5USEugRcRQ3DUGLYuEprBIMBAzCqfqWbmGvAYMe+SJPtRC4yN3
zTBGMOC7fnPITWvneA79XRExrH8VmvdTinQH+c+A7XjzB4I/TP5Kti40ZoRljqFT
RH8k3Q3OJzQ9Ha3vL4zjIuMc5DUN6gjGDBQ0ldOFf/j3OC8bzDQv4YR2jc0b8UvA
oigH7L7JQ3xSEtWnZDmGxMp2wnFuU4qHD330YIn2wduaX7ofPx32YjQBfP4dwy5K
6OHy0X67hiScChi/Cufyw8DJYT3yNkuntUiMunQDYUnbNNXATtTcLt9Rz0vSKNd5
pnH2+8UH9Z1ywPYVAadMv4/m90oF7KjL11MQnauVzjVKR7hNxTluMxh+1mGCbV2p
ULXOblXCVCxfAPEIgg8ZYMQ2uu05L7FAGzx0LQA10ZdHaVxu9uwpVeXy1EZ3+qma
7aNHloRnZJeQM5nxXLgGjm/RL3541PceWuE9AGGl8RT4ChfAaTuZno61Vtfacbeb
HF3cqtqaKj/fM05lYYBS2e2NX+P5H4BIRO1I7b4HeLslwyykO+E+/9oJqqF/Cpzq
ql0yslbaKOH7xOwVaC7IKHvJcAVrOuvvwKjimAPW35DZ/j1lkX4XqYs3QVkZ8JMo
4AWAHZ2vl3yxcuN7wz0FJ5hpLWvA+SBrEMaYQX0EHBq5azUI89BAXiHzSOeOozL4
yYePxpowtp+Fj81XmqSvmAAuOXqBZOXd4Cp6FOOh1B0C6USmbMpA/LJE9h37Bdip
LPXNxVDC/HZquaEMG52MFYBFpSNZM+trChAuiTxKZthmuadFDrTXM18452RfSy8s
JE2xO/nKmaHbMs3uyeP83iBlpeDni5n2FJA0D4WKh4v2bsHHndmrAK4dFMBgtes5
9XXVYR2NP/qZV2gqu+I7o23cHPhTCLSkIAReqZGf56E2x7YhMTA2qm4mA8bWXXdg
Ns1klUAIRR/BMtTCo48yCCq9iRq3zRaOcmuW/1OCtPMZqcgF2/rv9Rt/nZ8BqY/l
rrbpUEpBsc+4lRgaemAtJA/pcYxOPQYH+Cw4qTaj6QFccJzBwKDE5oMxyj0ED7I2
CpQOuZCqG/sGCrX1boI/mela129/tmn0bJWmKmo335de0mr75lpGpdNNQswoxJFG
pTnBAkNvVsB0Zgh9aLOKx2nvcfi7VTdKvsyuGVFrRDLXmlEsR2H2UNuT6l/r3UAT
F16ooWBlDbWjFhSRYPh+l2TxDpF3vbKGH3mdkGsGK5uomTVtFKmM22IMJFZAx+J+
sRO2tVsUFKaigyzyaFzRXrGoggD3kIqn4sxS20vChDpRBrKOF+5hXGsdNcAsLgoo
yeMl7HWKoEe6/JjQwzDDACsnEFffWZk+pYRBmVdF4Qkb0DsTh5/71+p2bpGsS8UE
7Li2GSV63wdFXkRSrsrQic41Ny7gtyrwrjs4ECXnUtZZrqtwGohaayjkw+LfHjkk
FLbzt/gg9YlIBQnmUvDPnNjCKsRAWeIgWYMx5YU44FaOhrG1diN0tVjNVv1yNkfW
jtSBdsKKPThgS7X+y5aQ/VqdZ5gYe5vqHo3IfqrQhCw1tlj7IFuTT+zmP52j+LxK
gYh6yo+ClRwj4PBTqOMEoh/dKDF/eQCDk4D0p4/B6upbQd3mmkm4FhFBmysUkOLC
yf2S6/BjvzMIC7RYRszf1S0mNNmVZTzzc1Td5tRGELawOaUpbsDmWPJdXp9RoSv8
m0ERjSHOILGL/SQB4Yghv91nr5oq51JAob31a6WF+IpinSluQib3yYMGH1sSs8Bw
m2fLxJ1jcMROYqpJ6pWWjfVQxQfRv44vQCArOkoOA95b5wZ4XVWHpbD8TOwnP/St
7k7UfK6uBHipLmrHPXAMZMSojmCKU4ZHx1jYFpceTOOWoz38Q9wvSSbflkcSxyFY
EWkdEwCPxWvjjP7RyhPIPRfH9V8nG4+h2Wfnp9mCbjOjaRKaWBXzEEcE/R40w0CE
4mHkI0/OdTlgNinZuT/NwzKzd1+IJZE+F3lpX+H4/52LZODhs1BWsY+qBrWZXGpn
iCaocoyAuIIs04PRHLltglC/kF2UkvcenABfli2mlamNQJ3lpbkOXU8s0cgeRw7I
IUhIM/BHo0Wk1Fv7679u6PYfYBzpjS0sg3jzFgvzkKkFch+bbPyeANKQAnslrDTR
c5QwX2aHuTIIQwVyrFg0NajJxNFXkstowH5ThbldXMuL7BkCeUaJBIGSO7M3qspS
XmYTI7ad/mWHDAz7A8pP5wt4ztQ533nM1h5iRcTaOdjkQHM7KVowLxnxJhdzZiDC
NLrYHA4FrtlbYxYzBkcqhSJh5h7dSVaO7AQXZNnGt3tvedMOcYFod8GbWckOc+MO
d/qjcfUFpadBqgtuaWShUV2DmNR8pRZP+Hf8vHaYzZRGxoJyPL6svpNwjPxV38os
mmfdZmv1D6x6wkc3mEgkCg7sNsXHQFKkzI1BGiR6QwYqM/xqFhvxY7+sTM987Xbd
4C2roH3ILIE0q9humnDgToGcfUpHGX8LMgb3jjzBQ+Ecx6bhPIqpDD6Lt0iaPNN5
HrpeXWxG4MTAmKE7IUxj1a9QYGedtKfLy6in3xHEB1hnQ2LEn0CVuW740LlxZ6zW
W73q4oyxUoCSv1//kgJSt14foIceoI0SmI90erM3JIK4GOh2ODa9x4a/xJpBu6A9
ZLcsUs3RwzbFXcQyUNthynucTMHOwuRm1gkhsR7N3tGWN/U4rztJ+HbtWw01iLZf
hvxRxqr4/xDEEzX7yjItzxg6s+R5brjrdG8WjQI1d7r2iQsQvZyxjM59YKc1fID9
2ZJaGAsz2qwD++A2sUllK73CR3WObUzK+VMSG0U6g4G5dPSIzGTl4wVvzx6wzw7D
9PnHa85nchcNEfRuQCJDvSGGFTnGBFJaEtDylfhvKP12HPL4XxQO1GEhJCxmVWcg
UnSE+PhzEh3B873T5P240gKvbp2fYilDN/PZ7dqQ3dJNYts4/VEK/fNRls9wePzQ
fk1u7tD14zxpyWmJtyOH7op2GblkWhW9+Qh6g3HHvGzvaDvj3mw0heBf4d3MyZ0+
AMlNuj0Bv38uAiGJCvSkdBKRQoo5E6XUO1y1x1Ua1SJSwxN5gBkxhiri8NWgiyzg
8CRFxpDeMRcIoVt3Gr9IZ9JjZPyeImhrm52qucnVahTQ2vfDpg1TPvOnHoeBJFW8
rxzTAIR8eUI72mgOM7JURGf7KLbI1+zn9PXU3GXvIU4FlBRWwHCPaAzj2iN1z5Ry
M/RWwlD4kDWYHzEuooAN1gFzOa1XwnmtIEDECDm3BoNeq2RcHECT0OlZ1xfKuRYB
pAb3w61lG4ZbN1goYkgOr/A8hTMxcrn9F9X2NXtz11EsweXF+2gvPEtIwvVo5xS2
UZngWFj37rrKTneGSSlGDnzJGey+ml09wwShRP0nbmsxTFAifv1X1+tW8JeDdiE8
OD3CnADRNfrYiF4SyashnH8SmZ23p51c6LYaf/cko06vphFKdckZYnOYiSH+iuOW
VEYruKZVF67GT0Sz3N2Z8Xybab2l3J9A4Bew3MZCBBI7d9U7pYD+IH8IJmw1N2mb
Lk3Aqe2NrHHPpUlLYoC73l9Fl9XOeeoOuWwMWm0tOicQoB8Py05RowtYQCIu70zr
PfEdknT9n6bW9UMj2Ew3CW58/IJTr436dAXq2T7BDBY5oqOpgW6MXRB2pfiqLswM
uuPyilUnyWPmP8jRcMCcJAWiSlbhGIVjc/NH/xiTSWTU3NdPToUm3SV3hG3fHkDV
NeB4m9oL+zvKEQMoyjm+h1j3wtrVI1ycnD5BFZ1BEGcxtJqk9oCyjlwB3mCLkmuX
Sk8c9U8VQbuFlIMJQkh04sKtSAzYfheMc8jdU5v6uzCXHBDA+Brx3UthFT65RVjd
G/AxWMrJCGmowy69fBQ7vBmDLNfvLFnPa8/Xa5LWPAOaBdkQjnXoZwmR8Jj9oe2f
qSyzlEKmIZKydK9DUrIj90EIJY437nKqlUJuGpqLdifu32cZlE28DY61l2tSOssH
cAvmdRKKJvOdHCIzqRoMvVf4lAVg4V04/lP/aTqyLivqulNc2CfgfO+uQ5B+MBfU
vG2zKeHCYOzOZPt+28UubROP4CzZL0vPZKVeCdchixaC/3c8zWymwVEzcvLG79w8
kmoPgDI+ppeBtEWnzuED9whJNjOJNlr5IUnaJeZLiDlsAEXhx5Ob1VquGScWqaw+
+Rpe6SjpX5l8zFRrIorTs5wQfwdb/pfyKeSLxyCY1utFuDcezL6HNpqVDDwg6xtp
X7eQ7hSfI7v53Rl9vkCBPvapgGebzU8z5f77wOag+8hUtbN1V+4JcNs5dDu/dL5g
G4+v5ia4dQMy7AGMrcAzNcBMJ/w4babbLiY+sfYSpcAtQkpvFt9PJKQQEcSXbYDl
FMBzMiqP5ECgPnQZ7zUeIPyqDm4/omdRFTrbJ5jGAbPflgV/0uP1O20LzNxN0GcR
/xtzrVCb4w1wkkk25tTPz+sUicBnKxEdI/dIgV2nFZ2RPC99TCw2IZEU0in/Vksn
rm2sDOZ9jJUWn5s1ezq+x9I7bN3Bre5MzH6ZHkavi7BgWtNahcY+W0q5LX6pC6OJ
p9BJGsOSOxRckZAFNl3+LHJNY0fPxVq78VLhKMabT25nPBhIp/7TwzHnIMXhVzei
3V0s8AjM9YTgUed5VTK/LStvZB7D5jxRyCxEzGeKR8oh94U9AOM50yFogJUhzjhA
rbeXTMR+2q3fyk3lgLTvkoS1UQIuN5geRUxICkAfkBzO6l2+mhG+cuIt9+qPQ7o+
Rj5vwpLfGrmo45Exqc1hQphPP1A+6mdP7bVrj2LkZXcKq6nzHBg9EY1jECU613ui
qgtt+bcXYNaup0KcXlcQQoM2y4zXRtqIe/1tAdajk2awI6ixZ8C7zjThbkKVQYty
v3EFnQ2MyJ2jPZoCoq2FgGkHp29BQ3hJCVJRsNRrYiIR++Y+zb7iZTawv8rf7JrJ
SgPKG8IlPkJ8oySD+qgrHB1MB6zPDJfvNYYWd/Skyutz4rLvSUtavtT/YFaqZedo
nGsV5838vFP4GTCagShFvLY2EyDawISmGG+cZcqzWpk58L2pPIgczgdj8qlkhnen
2M2xOGhh/Jkh9hsQbRutP8X3A1IPscf8JAg+uxS5U+GjHGyXaEwlMCxhFlGlxbnk
YrbnHLE2pemxHynHee3VCUM9oPPNSUlHn4sq7EVhCNSANtT6GWVgzcPOiUAYXXbr
oPH48w/wuxLK2yrfeJ0dS9sBCmgRCYH3OaslvwwBoWccI6jvUuirSGGn+Pj2UMAU
xqAen8X+guEpkeLeN6VE95lqzY94yqSx9sO/9X0v3WDXjxp17lrr6M3wO7pran/n
IcKEGu9eSE3KZuq/4EMMjK53cRm1r33G8dpsoBy43QZlifQ8x6Ojxed6GXKmCN9U
UnXKtDC2CR4kiiuFHZrObcHuEICVy/chCik68qyR2Ks5Mx8fZJgPe6lDFzI9X2ge
loepqUzIAp+KtOZ26onGDn4r0Z0L2+YDTTYqrjaMBgAzjbCttGD3yXOVW8RMQYgF
Aj3u6eAayapA7lOH8dkAabkHwl3jG+vELtIc7Q34XQJ1P3zzpp35AjYj2YIH15hV
o9X3wJuhLpADTdNkaNeeyI1oq7P2YqV1lNoCZhELp7YMJh9T/BotILD7FqnZC/Bn
azapAfaueVIXGk1PMEUKSjTVJwfR6TEBDpKK4YadvN+M29IN9lBNOUE/fG/i5Hzf
oZsf0Zfwwq+aa65gHyoK9ImYjeuwSGsuQBF1OLUf6hB7j1u2ScJihGvkVC3oUdiK
/v4BdiWAVwJVyurcJtqen3Tm3yNVNGSkis8R0npFpr5hrUyLm6y56beb6/sKPZOp
0lNfEwlBE7fNRWL/JDcolDRaLNDGTiuDVOt5gSndUbXwvBee4cHXScTA+/qi/I7S
FMTWh65QceZZtc/u0OKTD/2OVsrTz+ILKev2BZEmXOzLhp90GLDtzjrwPt3QuxLv
0Ti6HX9iq6Mo4hyG3f2y7XvykuenGoM4DguSuYHh9WeNZUKlfM03HSHFmIOXgLWG
R9Vq7ZaQ83IrK+LHUpbV0x+3esN/WbhbctEd0yFIoekwZqLkUluqsnQLBHWx2a1b
UpiIG7a7vh+LWrn5JMyrw7Rv8gYhU4xtTJoUbJSofxR3IeRfGnxxNsUJts5cdQqu
fdZ25pbCyQLNSdeDi+h30uYvnSXpvqdhDYKpIgt8wXRK2YCPV+xmoavstannRnhQ
z1pKRIpDi96lM0466e07ba+cGAB0N4qYVgsP1iIlUG8edzUf4N/Pioep9ezJX+md
mG6SK4ZXH8l004nZGflgbb82ZyutAtYPd12vN5SjFcRAVCoF/ZPB6CsCZWMcpjMU
jDFITDrVlvtUBVr+UGoJ74XNCz8p5fJE+4UkPFyrPgIYqAJbbnJ4duH9I1DMOblN
6RANHhDvGVjH52fPZc3aCGD1dioeCHLJwp195Va9MuFwiRWMBCE8o7KykT+eiumm
C92yt5cDNgBzmFbaZqZIGlUZrPRIL96wrkWkMc/aC1Dlp2jq3RRhKkCvpXBTpv5W
1DS7saKcKKuj548DHB9EQ9nzX8EW55gjcBr93qctVBLKkVFQE+cIXT/9ywYnD4il
kbg/Nr63tSiZ5ybmjLe0Bm8xGFW9w/9JCxCHD9PkRfUzMrUb08EHB4pORjrhOAZQ
RTXbyjTUYdAVAY/O2QK+gSjfmzAGXNt5EZoh/ql2oNlnk8Sg0IsV7FZYtlUh7FD1
momPfG1UZyhrmUaejhhzohiZ1P7/pNQ6KwEPA+vpOzDVZrQ4nCqnBYA/9P9VDbao
pWnDybh8dI2iKE7NrvdvADzGWUVNvkeq7l1uGwMJerPq3bFsuB/rgV9BCa2dsHDv
ufNulXVmfywVEsMhySnkme2dXI4xlEEmxle3DRdVqEcyjvz4M3FmEMw0szakX+5P
cjCr2uuCYj34JzIX0N1JGD32NnzsevgNvOZ7hV/lgxxpegyYUGkoMCSzXvmf86zf
/vw1X2Kan+p/wft9ynBWFRr2HYwCHVZ7EDr9rlvUSkAfgTMx41Ii2vQRhpRX6qdO
mtyYvCo87hYNXFw4Rut+NgzMOA3LtQwv/v0GF88s8rS4Q8FKulhyJb7Rwg/RMcCR
g8nz37d4x2f2frYWVUMWmfCpLVOK0DIHzdfA3Sjf7PnMIuotHbPjtye3EKmaUcdr
t11/9WUW7NoPBbAxP9Hff7aV1QVuvfyTu28nq7tHoN4M1mmPXlXqZWh9MkpQNO/k
qE8zdbpOoqX2liU5ArGGiLt8yx86ZmJXYkOhFLYhQ5SFYU/xOtPA6mU9AV7S8qF1
Pabq/ihvuZijSRavSHaTzel+nyRWv4PAUFS2GXE7jt7A8JN+WhJCt0dvxRlp1hjF
YnolhPPX2RDnnoDzBp6WVXbfu6VLVuuB+FZvsoH75QwWCVtka/aonHqHxJBAySKL
Vs5qXSuPewbwT0qWR9H0iBSRf0aOXN7snV09kq/M4XxsJWdFZTcESweetQf4yalN
LKzo3p6aRtSH359upXPQI74tLAg9qasHvNAD1W47ROdfVQCTE0EyOerd3c4uZ5wA
oHgpC5xpEUBeChB+N6vD0zDbPFoLujIKMbASe3IrFUvuVlba1QjL1xV45bY9//ZW
/WiETcHEdDJYNch3LmpR3uXfXatBo6+37Bjdn6RziwMPlcBUkYsHIBSao9h9+cya
e6IDd9NjrafPIrBVUZr5YYglsRDQrvdrJuqhhg8jxGOJ6L50Lh6XrsuEGcPSmYCH
vDbS/64NmQ9nbb5bFFpeHepf3DF5NV84vwhoLlxvaVH839kuRU2pylYhYbDx5kdI
MXuuYfT3mfrxrgcrCej+rSNTTNCacp/wDqEcgZWZPFiqhuFUWs6NZSLK57/1xrSl
yNwHExqvIe1AhFVbdUFWKKye3nqtGfERy7UdkEZSIVsh3lTSTTQxMfYGPKr7L4GL
sphsmM0/zuGOw4enugvyuTItRumaJ1P+xSV8OgznKXCi5rZuFlqlSp/t0PVr1wy9
A0ofU3S1toiZSfYg+Q49tI00VnMk1BMTCLncXJuUR42DLTD2oRTXeUbtZ4U+7eiF
4GmKvEg4/UIBugihGYIterXF8z5pST+YRyHn0cj7KOpxE4Kxk45B5K19Sxzw5KVs
AuZoL69lunG54rpFDOIEXcZtWpSe3n3PzHjWaYvZ0bpx0Le1ant4j7TH0+nuQBk0
11dKYvi5h0xYHXU88Qi0SBbUffLfuOIoxfmgSFN/87diZZOO2JWVNtFKOjrsWer7
ztEQ0H1HMoyDAz3wGBMcaZaS1krclz0TTNJ2z37wgg0fswvrc7pxFaDBStAWlNfO
pWQL0B2jUVBnMLtSYnJqO+DXDUg6z+iUj3lF1H96YuUEv0U7dhnNS4dhE/9wE0Wf
eO9l7ENtSkKFTlHx+1ArTuMF0oH124ssLBoxCVMqUA0T66CV5Q4RUUC4BMf9kiXJ
2ItwEI40KI0Y6ESKe59OVkVQVbVlVxhn2iVoypzxM5fL72DvgdiB+V14rVktaxjP
mUoWgShjbW2rfDNus8ZH84EiYFmVtLfP5pKVwjYxzXUf4B2pTQrHckmrVikoKIbQ
AQ0WDP9JucYoJcBBsz9tiBH68YvKuRT9EMa3TFZ27gffQrCumvDz7kkZsBgRJd71
vvh7uCsU7rabNJ+zcp90JmcY8M0T2O+x77nxzZQxYa99yYcHhq870eG1om8KEN1H
rWRzEY7BTIvk+GpdRPh/EiyB3MNQjqobAZRLUQ/5iZuH9J1jHZn1X/Yv3sGBRY8E
uH9/ovOj/2DWdoj1cndddEtVyROuj2xMHptqdb33RqheNOvUZN9P6Cms6c9GIPtz
DvxL5td0+qlfkhbO91ex6NsRLFa1SDzdt64ve/nFy2f5jQPt6ikZOOy4UUAKTXSf
yGMstx5gzK0Pq9HUHH52jkE5h7fNvyzOLQeGwM3U3gTHqDhLmoQMUt7M40PPJHdK
Gy0GuZISitcBMBFpNLzfLoD1qblmmH+WEJgA2Y+HwYs6CGzhIXh4JZd8K+QI4gll
7sMztyRphAxoufM0oEIP+1SCKIsps7uK+K2zu+uxQXCrFJyWuZIiQDCmoZDJBH2N
OF5m3PjbqJmRoJGK+HQLi8Ezx5GVw/U1qYqwwHmBdjh8I+7aMV63NmEioegIR/tV
Xy8IhtdkTZGQKfNnr0wcbMpn6K9QkpIVi2pD6jT3ChplsngODyXQNZMbxpuWNS9Z
CE44a+2JxG+/l/jDQOxXVxl/Xkd9ztwUnzxbyN24sL6WHT7TyVXuvpCHQ4eFjMo6
5rPnQSP5o6gV15OnLP21EFgrYhNm7bwJIow9ed68BL//r2nK+cXPiQOXZ4tQ6qee
OpoCd0wSFKvv6ZDfrqyUYJdyAV0pSTOjopdnoC3NlZvJ3VFCQft0ahDyBc+FEHME
qPznVnuys5bHdlqrk3Nh7qZElkmn/+3AradSjutY+T0LaytGuYR9RpZ//LGEcxO9
MOxgUh1d3h0RuphjkQdQLK4TYS1i2d/VFRy3bpdeWEG1Mr+EBgV4Omu8bB7ZmHck
TDSm9X8BN+9IZ1MS9BcYzos2WOIeNco9Zr8enuVxmYOkKSf7GHb5k5b7CZSumrbQ
lSTSbOGAzE9rNXb9kvsVnGLxqVDWqcL4hZ/2n1cvyd/0Kryjru5W8OS0gvwS+aFA
Ye3cuEoXRgyvRONUSwpiR7zf1LZyRzxjUzCOZtWyZF/82Nr1CvBFIQODMiXU71ML
4mOtBxzWcOZajBeCPphcf7VECY2g31X7o44SVxeFt2OzdYH/T0IzAJhUB8MKTqst
ySav6iO7z3Z8oh9pchRtFkQoCatFnKr07eZS98N+8huipaJvDefvVcsptCrPZuK/
Jhy6nzWRbDG6LXndIPlVY54zTH4gXMi+Npcz7AVE7IRYBBiEIK6vswPE1yaH8HDT
QJeZRpymg4zbXuN2NWN/I5AFX5P1LhkACSyDNcw7pbuRbP8o97NefZ8V7p6OgBda
hzq9DMH9Qs9jA+Ib39hhCsy2ywlryZ+IV5oAXqa8EZWg5cXBm5G5gIcqLmEDcpvC
sFOY1i4d+08IIiaFKMQOKS9kYh/j7foiNfIi2lEUFsTylSX2sxyirex8pxkiPCz1
of30BKorOe4gA2X93Go/eU2LHG0xf4Lb6oXv0+aQcGNNxP4pRM14t9EOAmcQrhNr
pIDjUXH8iwDkqm8pxz96pcjfpvNzHgbwxeaB7wWxT929V5yKuCGtr0vcEyIEJ6/v
YHR0eklSl+MSNBTgoZ9dj1a6m8gUoJ+oefgsH7T2vUehV3e9jB07LVdbERUOUaKF
9O5KYwRGLfqjW/qCm8iMTz0iazz4UstV6WxLTCoFNtAgPdK3dU/xtBd6GhKJXOfS
ijD40p7A6wNNYwuEfriFnVppgLlUM4POmbzltDsJii/C5TXcm05RrOyMR/txBXgb
ny0R68qi7WxnWKPFgZPVK7MeeOp8HRM5A8No2sgyNU8YgbwgJXs9lWtNfnECghBn
YG3xUaVeiGij48QeCVl0/HqD6RM4ZznTFbSdwTxOqNzbrRCFwYkCpGsEnim/i6o9
E10wKmW6eeB82XM7qdO90BzAs7Xx5mtkUO643OQI27/wzPs6fmTs0PangrQ104KS
I21eFBnOJktSaGCN4Iy5o9q0Qc5RY1Umyf6WvzqHjeS4xuExyDe/gXj6h4G0dSEe
dk0qE9kodu5QGYKvwaYstBzj/x6NYLldVzI3Sbrp8GYRQ65iWVkd69uBXAD+c4+5
/vAZLTBKb/G8rVRQU6ASkoTP1OzSn9ituJvSZcXSgYh+ftDNs4qEZJP1oJFq6g9U
Jy0r6YqGu7ld6Jl0r0+t5RrMkad2L2hAq/wcdT2th38jMvXpSm3c9OEnFQZ3hgnC
M7ofACtT+BG8XLmI5IIYGEVPC4UvJynakh2eA0N6KhDfFyilinDxIzesneJvSS/3
b3sCZXOWJyaO2RFRrvq2PXuw9I9Dve/rp8Uj8I1ghyV3jERSCed2MSup+q0s3Fe4
U2U/WG+0C6+GRkS1QKsVuTxxdQqGOd6RDtrfGB8J5cBAtaMBko4l6++lu/gaG6Km
co/5Cpwg1lPdtTjcPOZsa2np0o4GPcHp0HTsXCBnuiL83UUUKF22G8R6Blc+VfNh
WZoiDtqBWpvRZp0F1Tp5s98P3+0ieHKp/W030U8jzRpUJcGB7Shkm9Wf4bH05Kro
trZnhXqCU9RHHDsWqg9Pzdkziv4UI7pX5r/SF7W+r+sXGeKAKpzQWw7/+7qWLfqQ
5Ux8RsrHlK0GgI7XVcbecTKl+VdGEkG6JROclVinzZpzZqt8wA1DTWyZkx40fnGb
hRDNC33zvOI42KW8Pqqq8AABvPEIDKNzTWJFa/wMgM5Tm6kXmEvxkHZ0XIiWJvAR
a0xxWEuxaGeD84w8Jv4Tm3EPwgfDDIOT+X4wmKeOX4BLPfuwsQ0UFsVetSF6COoh
KeKfSrBcyzWc1X5vyL468uR2qEmCQQFQCxrWiwWPUoArW7bxIiDi5QRrN82ymIvi
/ZKyQExvs+7KVl764eCNmaeEQHev005+KhRZBvEgdFEGYaLog2wfFu+ndbFUUXvn
yTB3HJmLIPNOEIexl23/unp8n1fJ0TcNVjUEQnV92eCxDj1O0jooF3/AWqXzEt1Q
8E+dIm94RPH08/2/TuuHdY+CHViUyhqAUhT1M287ANBdGuAJZP7tRIPn+c5Ytc2A
bn6SJghZom4hz7mktucqDIWtAa4ZtOaax+ApEahCg+7RbtUR3BfqK4/p5/hqDYQB
2Vmv1Ipeh/P/dVyFIw0+D8NeMdtlqoq5TpVfYOn8iueC0Bt/SnubwKc1aPb+3oAk
c24P0I2zEoBTo13LUhxIaeUZ09fAMxsXSgKxHXsm7LqQqGNACm8t7I6EfRHW/iCb
C1eL6RsPxHzWKXCQZgc0c9helTzW7PFFYjnKFt74DygYyCIaGV9WRIwZxgsetx3H
ZP+LhBRdFHxqMyJh/YOjv5XALayG5qfPz1s79B+5e8AhFpO+KHFWvp6GxRofhq8L
2X93N35vel6v1IJnp0hjbXyrCSGIpaPmx2d718XowGUOrTT3k48FXoPDlNW/Fp2R
LLmHhQEdhvdpKoGC5Uf6rtvcZtt7fnro428IS9+KoARKCUF71mzFbmxG4lNolM6p
bHbw8kZ74jyH56t5V9LRZNASCi+suxngzS8S1QUo7c6tJs6GHVPcisRT6bkoLd+N
hkys2cnXwI1EOmPg9vu2fJErdjzkRL0nVa5U0RJRvMz0Z9bYWd8n3oLav6DEVb1n
1beiCZCiwuc8SDtnVwNLzEqpQTySB8Dd/EYaA2m7jZGnZokES84bYt/lWlUhFT84
iACE8bfNmbX6VMqbKSIp3Kx9qkP3PdFWOPvWHNoc0PFjKTeBo3vCO3JjQTO/UGYW
jo7DAWdaHPGXOSS8Dj5rSE2ap6z89X+YvrOCauvMKwdztwyP4dr1pT6RM9Be20Wm
djPVsVwddr02jaJ3n2WKUFa7CIqPpBeEoXAw/0khEOskB5WAnc3CoQPZBAQ3fAOm
q8K7IEdK84q0sNsHsOu3KmpeMgo9dqSy87duU2Z0RtYjzUplXylP9C/nOQmGWGq2
emwC7HV9yhUOpa6INawGxcAgu803whJmPAluweAX6N05tSJJ93gJ7JMaIkwTDg0d
NQ4sKZnuKGUsaN3S3pFmnl0Fvxpd+wuxYy4wBXuYKlwJEC8cgEkCiu4jiK82m4yI
M1a/uuN15qnyuTw6mdOvHEzH4m9EPKuXuWxkOKkhvjfox6OfYczLQ1g7oPZn4zUR
3CcgIimRYH4zS2hVg5gIoLI1csNn5LeDhCSubWooPAw3zdxSKpgspC1zH8OARJHS
h5bq9nhh/CIpsfBPMh9SNTcMNzrhu3TGWSR9M76Ty0hyQZcEcAHevwmDvB0M6ZZw
oY5kWBgC1FiDY7z3hpUlQjNBy1DW+eERwxPM/Hz0ilPOe/oPSS+cIyTo1rZG26Lv
oDqDwCFi/J/OaonmnDEFGvAuBCRcwMV/GFcJlqu+MTxwo7LI2ROLGDigC9TE+nTx
vCZG5SLSGG29+q3OIuduyQsDCzxJryXD3qevrpqCce42i+YDV1C9Efmy/clYTCrF
TVhuTCf2Ixw+VI4JFRq06SyNkKg0ZHQjHKIHQUVRejj/dSfS0ljkugluhNIl+GV1
D1WG2jWAiPMx/WVrgTOGsZW4WxlqH8l1ZEPtXI6x6ijrJQmbdLxnc5vX2RAQccTh
axxYvbSxB42XnKbl4T0K16BS45Ip9n4GzqzCPsdHzq6SXNQgRcN2C/lyjtfkOBd0
Nf7g4nPZGV/UM9RLlnoxmi7HH2k3YyuzZly/PiB+OcNsbMlErkfR+bJVW3PlZ7Zn
uS2aySVxy3CyLA8Y4RR13tGLAf2tH7B5TdfIHCSXD2h1IlQsK1t7iIjFyWFailrb
8JZwGMreAONVM1WJl1CmAIl0Ox7tn8La/9c4s7lXY5bLdtfXT1/wdewbLjMhKxEv
h7yEJmwjTz/E3yf3Rz1uDlcYLPpVfX7ibYCbv50Opjiiz4viFXjmX7uWBkzWsvGD
kXNawyyeML6QNWa4yJ9FjwFiFFQGw+0vNtEdDnDxdkF+oG7kmHn/e1AVO2ul1233
kIS5mFkllcl7lAYUQLGLYjEuWpEVRwnrpDFt8NIMeOl9Hnu//p0L1QVYRT+SQdTJ
YsrerywWg5cpu9I1K9U2pONfkc7BB1hjs0Qgs410F8QSv7kPlgoijn7/IDvAy1w/
KI0rMTBB2oqXtQW4jGs2OMFmx30ovVTewe2LhgUjU+IpeBIghK62JcRjUS5kWZ+m
urbyFSwJSUSzTkP6OvDksgPboCf+OBQY4kM+EuvIXhSZtPR/3mLF0p6Sj9HmnvtO
swghmf1w3HGo1O590d5dLBGmLt6lTfh/fg22aeYDsxNpX4G15AtG9Ls/0551QxEN
EMCW73cpa31h2aYl+H9phVG2k1wZ676qktBeBF7rnqVGrqFo/FMSHo3iFLLHmlKW
HM/hzm2nrsENUQ7SCeo9fnZLVk0IyPoT72rCvj0CvB+lx3/A9KCa0ItYmi2mCyBH
CyhbeUyZlIL0TqKcLFhrxtX8iHg0NG+NfvplVA5Fgxgr6p6lRm+4tOTjVL46cFwQ
SzxCGfTCHcUP1UiMvUmyD4903NaFuhklje3zWn/7AZvOGeIa9JCwS99+ChHHm/mN
GUNjD20qGI5HHLMRaCOwqNkRPZ7AV37561w3tHWajGH0J+DpVGo1Ee7YD5eargmG
1UUutAx/ThlIFlTZM05Hq//OcxSYRt2Z8EKcNIkFqeP0Zm8breV7PIxDqaweO4i/
gZ1sLvGWTzGMoePJ5AA4MRdrKj+NNTZ5kSRdONO1dQNCQiNEub+jmWnk1m/kbUOV
esz0E153EmugPdm6GKo7uhIbC25rHYr4gkyEp1WJA4GsPTFRW2umni8XqSHAJiMB
tJk9CXR61RLXKRtnslbe6oTYPsR87684iTKM7Ttbv8RDEH5Fa78GmmeUyNS6Zmkx
rpt1djpFnpst2E+K5esd3bbPhT7jpWmGJgFIy80ebsuVR4p25Q3BDBannwR8RrXE
dE3PxkmIHbpp4+daRBIzW7Mz4ONQOdbLgYMFPaanu3KIz8gc58nc0ZLZv44u6n0+
sMRtT+QSqDuM9+vYNE6itq0lT03U/tUB83vSr8+y/lR2wciVGA3b2TV5v/bApL9M
TAbCe6ypZUxrYWbbFQpFAh+kfYUUTe2hnHTBeScYY7nJFPdWkD4Ls2xln3r9bceS
SrnUTYTK7gZvtXGdSKT7ITpCsqkgge2L3lZQH+PhRXnW6/ITm0c9cNB+k+Fzb6C7
9LsGDO62HyOfxRBDklRs16Dag0YXuuROU3g24IiaNBkOCL0BGlblND/angFF2ajw
bgZdO/ASyGw9aVZEJP8Iiovd3/F1GJlvIjgy7ke5rhyFqQ09Udy9uwaQJ1HhfTvW
zazxGEkyB5PV9ZyWk3cECvEdt8hf6lyej9nNCmBzrR6ar/3qphGXZBWGDM+v4k1k
H3hr2N32ozIz1t1wd7Rs/DzHcFLkgWEhv29OnIXRzY2WFwMW1pVELZLKmbeHcg4A
YJdddHzM+friaRUHTkgoAwQjyU6pe0wmjjG+ua+mVWKbMiA8MiJlEuFJ14tX/60F
jtMX+YmbieuK1rjGU9ZsrAcOzcpbAWVDz5EkloeFJkDNi+djrYhz1je/782Off+0
QMB21250KCtwp9Fo+V1EF6+9Gxf+6L+xroDj6Mjmg4Rq3efYdWtpfyPZNcBZV8H5
JJbxoHt6dVXbR7YduA58yULPY2x+5No9JOFdq/wPIjIP7PlR9ZOc/9v5i2nwlp5C
EBKkkWeC8TLsQ6wPd4rNGkchaAcpkyJpTHOnkvOyn79iucBCK9cw/J+yS4Mjsm71
BnqqTCMA5pnNZmO4jS0hRqLxMQjX8pIgQNBo0AFj/iQMugiyHGRd5ZH/XHaJ+Wzc
iukDQsx1LjYDrL7INL+1kHX8m+Gq1W0InwsepVQDAdxn3Ai8QHEqGFquwIPp9u3X
lVYtUBRNAl/hAooMrjfYUrP1YMVuCCPE22S/uw6qy3HyqhvsSlP2N2jD5q6I1kRm
Hv7uX3oJ1y2zORXyJlZkWgODDFOLoWkRSK2xwwgadlV+fbyKS29daX/INa2DtehG
NlAzA4HZozUUFDHGASM+OaDMWJDmfRhvjmgM6S1zwP9Q8idsmVsRFbxC+bD2XITe
m+kXbVyT4Jp8SBDTIHJNDCuGFVl1uwPweWf4w/JVT/Iov/C+/qZ1fr835+H7TcqR
JB6lmgnENIth5rwVD0YnCinpB4vsxbTeJqHbEh9tVZh7V2tjlOsZ9ewYYLYCFEqq
KawTh5fA0avGUhBNyLT5LrqwzmxwKNpxHQ6WXBhzkdyRAhoTQFA73TP/5cTW694Z
4xMhE7yAYe9RAxPE5RS1NUIr1K1cGkl/RBgpfCGl5PwcffOeLQmuWjEE5pmaVo3n
FYohiEJ5cElKCuGnmaJOZ23xXsSXz6944giYFmU8Lxf3Ks2fCFF4HvGmd+5+Nl3z
Awb8IfVovXf7Q1WtZZ+lshdAXvYptDo2ahejOiNrsk3NZ7SJtK1qrQK+5kqjlZFy
P12WrzNM7w2UfnjY62MIzSJc/aJyWiCCJwNT1q5JtQRoY3oa+ymg7MjypVRvSNVM
RZbt38W210c1Y21ElEGSi7cYj82e6cUnSFM9BZGYYJHVABlRZDXvsdXlIw5M/RrO
izVbcWOwl9FkSsvWvWob0R4WBpLRkn69gumzvjADhEG5/xMmn0Rv4FrLsocRCJfF
/Kz+HQnme0V1/kmLyjdXGT0jZ1qoGo4+DYuSP+o7BfNPpQFdLQ7IDZtZkGxk3ikM
5EUrtvPZpnVvVV6Gr77b5R5rfkgfz6/p45Jdc8LDExCMQhwqPWcOsR20PhS8ZTWX
w9VeMBKcmADRwzctgxx40e1rFhsbBQMK2BOr5yuOAqbxmtpVlsUJpUuBVfbnIpeY
+LZS9o4AgwC5NjytxJ/SOObFZ4/Y2Mx7DcSeycAbtUkz5dzQRPWDd6VZ/N+DP/1z
MzEzN36DvIul4nUtuuz03Z62FZ/hpw7FztMfTA0J5/uPxdtWkavcNK5rlRazUcST
hVo8wmNNHw9Gb6yKsrV5FsLfg78PoSAXjhWpOkhmAyv+bA/mPOGjQcsDQ//wjKbv
AYErF5N134HuIMoAK3gSJ+fdM8n698A/YTR/SRv9UW2Jn00vbjyvPCWqYiFdQ16T
45TMA0zR+wj3kpgJCxexudn2b62P+CVaIVGXFawGxc/6coYuPrpchESI72oBseWm
FizAI8XE/mkJZoir4YrQsM1LngHe181bly3SJd+xMHjDKouVVr5ffy0wD0mDd1+q
p704C8hfpq/yblM18EjZt+tBkSU5HwhXX31hio6HaObKhdtQr/gXHW1W9WYh+VHw
vGWVWPCnxo6b3xGPdRvjrx2pM6n5bCN/4zwv9SnSnthilMdY4IzsovIP3nSO5wdo
DWNRR3xXHQXInbRv3TzD2O/+B3dCNbBi1UAsDG6j8yAiT9kwQdg0AR6FfPqrPigW
JitKYVLcUcLM3xa0HVlG0e0My5xM1cXaPlDbXh/J0SCDZKd7nv+BID6qv8qHREGp
nBv9ujj0twvPhIcj7HVH06u/f0zq8/aCJc7rkcAI3jnitx36BNW5sJxsBLVsxvKw
D8JLxn2Qo7d34A49ykFzveSXiM9aFJaUu007lKqKI1eM2dHO+lckAg93O3P4HJrt
mfUBw2DQsvgegSvwFdV5rL5OO44q4oRKf1hn6CZd7Yxb9e0bTfes6ENbjDtAxtLb
1xsEc3wdsglyhTrqxuI5dgBbdrwciPI5Sn8m2vx4hsDpB3vUb8ka76+k7yzYCT1O
cadMuQhYqfUB9UKq/a/tBnwKJqIDVdWiVlYZSxwDM+3Hn5wP5CqxcX/0b4yECj8Y
y6yO42ph5/GQ0YbDJQMr0QlkanplI37zhexfiOra3hmNO9vvWq6Bp34Rhzdz+VAp
wIgd68DKC3fMrJ0mAhcbPB3alBOXEiFkCbviD3XhUzVx5PO7dzhUGNudH2O7+R4w
oN8aamhmhklBWOYZ4CLgE4VyJQ5C596SveAVisgX5gWHEzHxRw7todKpchCCT7bd
NISzppQ/sbmlOs/hbdaYNzMxcsmMo1XT+DwYLXow2/c/MhvdJscle70QmpxupDJM
YX0A1kmGCD/cJLa90V1e0EX59icunJM+f9+fZAJWIe/6eUDwrTIY4VF2uOxN/g1r
vG5I7r7sx+q2wFrx1/z45uGeIySWJ7+YnH9V27HjW9DuJDpZuyGMJK6chqHNnByN
V7BNX/eTBeC3WmawISK5GuT7Y9++dmlPJCf8+to5482kuNEDGzY9MRw989vB6GM0
C7BZSUhjXxZB1L8r1K5SlGVLeLdHAS5gUO8uxV9/ganpuFweBxG4cDYMkGMIlabT
6qYAqd1Ylcnt++vHyZ9kxjnkH9F0RoXO2qJvh5jZmG4vlT1Bp91QhiFo2k9pKogM
Smo2uXD+H+LVZf0gDLA5M83wFtTVSKJOjS8hy+wEPiWld+TVXdRlJhhVEE9aD7w2
9Zg1wVWSe/7hZ1PVBSzZ0HfyO8BMkManwNArrmLRsrQ9ZlyUCSte0UV6GkAMLdqA
6rXZLB+E8kevrp7KZer9dU13yskzsBNnLZczauPNJBSiACEA62/6ZmOwt2uuDXpe
u/OHzAUipLnMvg09UunxSe6+iBZ8R/POOplwS59S8RnONWKMYgDa4aEP73WUEp0a
Q46ipp5mi0W2cKRtAmmexjrtHx7oIv/rJNgZaoaekw2QmLshd0oA4mgGXWZzeoB8
60oIXXdVx7vYWxrVhgU+dcOVu0JFcg6kVrnga4rccOcTAb9zdqUfHUt3a6j96GEx
KbQ1Pi9Fau127xt4Ro/mucG+xxYGjLHIT2kmgrMAhhT9rXPuvR0Ab92Q0o/vPkb5
Auso1ivc2ZteOQf010aenRlHblSMGD/XMbI5c5QOpGfiGtxVfz3Vdh62yRvP9J+K
vJaMveFhGOO6EQeXM9L8hkhiOL4f/la6tgKrszJAkPw2E6T/Kt82UdWJXV2j6LGE
Ivt82C0oBe+xk82tGiK+HKPGHpc5+vWDppc95R7MA+NnGBWQyQ4UdhDV2SRqh4DM
Fb5zh1pIqULWAgvqXiEs8DXRg8RT97D9M6gZJaJycEkHD4IBqobiy+J70zNED/1m
2t6M52VPwKvETNCq/zKmEgSCqLSzZyT3XHImiiHNr4+PYSyoTPiyxco89cqYhXia
zjcx9YH9cy1pWmEetZs8zCGyk1GJsVT//KlBQO6ynURzTQ5HeObrg1Pf5s8tc1RO
ZFPTclT1c+1majhTOGe2piRhOqWxVV8fGw+2nC6yN0kfqs9YclpliIWfjH1UyKlo
9xNv8O3IF8S4bMyLtoqpzxXeuI2bWH9HDEGnEdDaERysjz/4ACqzOI65Hh3H4wh0
clUoh98jhgKHF5if1yI+6rT3ZGMav4yfkgr475ck6MIU83K0p/LOFUQo1xSQ49EU
3MG8UHpYqdS6zcopqyX7OZVHJRi0FUnNI2CX2Kxjg17OOQNbb7Vz/uFJnLBDF3bM
eFWr09AqcUhq2ntjPl4lH1uJ1qaePIdKCJWmqXXiEnYZbeRsam2E49y3jECdBYlG
N6OdJR9Bz91YcKM+ic+roQHSTUm85/EeeIHcc+vS8sJGirh78BalwDhn7rFEmP6A
NJ/IpqVI5mf8DjOl6E7prl8Q97UtLNiJWBHPDBg79Yv1aVq3bklZ/OQmdUVxAADm
42bxG0enRl18PCZTVYSCxvZyZ28tyNvDrFJ1+Qj0UjZylhhCOEn3IgkrgaqvLv+P
ecuZC9Bf98/m4E0OfDm5OahuBD63KQu0M1Lr8uQN4EpMU23Q5sMiGr/JnEVWn8Fu
jfGel7Kn0hSE3UlfgOdSC752kvB/iiCWb+Duo3Gx/r8ZX+27wPU1I7i17k/5DKSD
tMLQvIBffmYqe6/1Bc3iARrDWdrgEl9D5Kst7csySJ4cvRayvyuUnw+6l/rdnUbB
JfAZY2QikfSaL7GpygA1PreSuef+yhwmb7VshR07kX5xWwJYHv2M6MNtvisakUMz
QbNMar6KRjTcPqaUCuWZ7ON4rejaCDXyxxHaQL2ic9jliqzurgMRTPY2Ndx8ltq8
3dYkNgWJyvm6EUTclKer39m0ngyLYueWNEacULAWtLSSqDXfnnCQjLB6+DRAvRoi
+gfpHPEkxMeYbm7uUxmjTm3L2aoWhzMFOwx1aWCjolsTsQpBpIXO72CzrCECDhkI
J1bV03sqRwGNaWRpe+cl1nNuCp9Y2HMrJtLMNkm9woMfWrqocOuaKT1KwC7ESIMd
QSAvhL/ltS1965csqugRz5HPyADCjBmCsBKhUIOJiR5Q4xeXl6ayjHOG8svco6g4
ZRy0g3zgEiam7KrNTs3S1O2EwlnFUeNkSyNPwqOE+uETDOeUOcsCb+ngR1sAkQcB
7C1PcT3ICjkwbF0G2UXyG/ENv06E7tqCc3KuFFAIKqSRLjtXTtHhSpCyEDFGyT5u
Wij1mlSr2s4S0fB8WxtGdCxcEp6L1wrpYD53Qai/b3klnCFbw0wX5NNgzK/OKs5b
yq+au13V54eP7FsS/Il75TJ1kJQw3RGIg1gd/VtdrDNull2Nr6F6zR5cdOhLy4E6
Lz2Gjiy8FfGNH5H/SNY31V5G1Qi7YOj6CoNgZeNLjtE2L2mSme/Ve6QpFPZPPWlv
bqGWMVdERlLXkpgSQ9/Gnm0OtaL4zsfF+LRUrX3V7M6VKeouFlQ+jwXi7SRp43uc
kp0G5qbp3lNqNzp/CFKR11vovv1dqOa/88vFXnxFq7ITDBqNGqidRqPumI0TLkI9
SMeGa5Kwhu/19ewUiZB/6I/eiBs9G+278aW/AS93zCmcGvWsIOifXm9Bm86Up33d
Xf7CxpKL31VPjqPvPoTcq9mazLm4jW0k93Kx/wm63N7FnBwZPnZrr4Vxz68vXw2q
IJ//geFpC3T1VJbXApode9PZzWL1LE8xh6l4XJXCDI9cWo+F+Iqd3+tS7R6l05I5
KQUhX1HnLMtVHpcotRJe0JUUEI2//R/c3qF7SXBwPueDBIgja98ZmwqlKL1v183/
bB3evZMlzKtgWY6hwnY+em8fd2Y6SLfMqPcIgZNybkPbxRxuYqD6AokO0f6XO/y1
qk3EfRZUa6Ree5Pqn/Kb8JeD+nI7+FmFZxbOvLe0yGY+BVYWnBY6Fbznr+s0hbx/
MjxpJMgoAXpHF2CjeqtsjHDq0u2L0iPCG7U8OgSgnj9adjzXCrV9DvJfdz3C2ARf
u6ANeQ148utGUQaE37TLuSngH0neWbaK+hh0ITnp/EtiLWAmpfzCoB2mMjp0RFmi
F6DZyD8wq/1T9+GW64koI5Xa4bopX0bTDPpHa+aekPLo+wMjduLanjvySDigl1RV
t2KjXYH7U3U2ZRc2z7YcxxYG/sFM+0RBl5/edv0XRnR8N+pKoECjF1t+DPbyy2AH
rr55AZlO7yTvYo0ZO5budwqca77drG7KbFBQpizwhJGFcMy8Y10KLTORxzT8C3nt
TYlLGkuqeuC3PAru3KWpnlEgAk21ExH2eYXWcCv9Z3zQT1rTP+NCAM/Cub3Lcuf3
By+YaKMTWf876BYNCseUv0AronnM4810NrptCv+NfutmpKxK6iTX37R9xe9SCPbv
4pulDDtMbvKzfbTGh+QB7xXMe/hUGBpEk6Ozy/+uAGwvjJ0vApVL3aLE7Z2uoYF3
N/QLSd9KNtfeUKrSjSwDs6ZdYgofddxieaHLViphQiaLtZ6oRB3ygat8F9xOADfS
q9H3tpNaZn14P8lpfdZef2W6gHOXUuoNEdaDZXHwPIoA917PdBKEpR5B1A1lIhIm
TFfSzgzA4ORemO0UI+6Tn66JoSNVbqCsG7AH/1bUDH3esVYmvWbCVGWKlmi4kwAS
BjlGU12gPCPHolOokPuNV2AJONNKKYTX4Wn0X/hu0/iEurdBhOJSF6z0IXfxmMIX
XOZYLgdrFQGM95asPRJgSqD8eDzShK4GDSMvtvYNgybkn4stZLyK2QgOBA4ucDtp
SeQnv0jKLBs+vfEWrKo6kLixAg69dr0f6NedfLVZRm/ye2t5XFr2dObae3RJ4JCw
4lnoSOQC+jipYESq4Gna1bSCxEK+mF3nmyOfzaljwOBZOf6HZXOqnNxf7tpiXoSz
MACkMBs7ELuKCzxaC8QeiW2/DDVx6kNg6oSASuKJpK/kLmMnPODQfi3OytYJMlnF
MSsuFqBDIHrpGglggZYIRp+KNreQlCkKj97x+1ZrqNUiml8GyRWPZAXgVBNkGYVk
CiQ7MQP/5jHamYrzdmQpDbbZ2s2KVcx2LG3s5XsMkIrw2r7Fa5i8Yu43Rx4lEGg7
+nXHV3m1T2AgWPtQqiVabPoH4geGO+Tx2IDeSc8NodJpYKEjKOKxley8GR/KD3Vm
KzLDa7vFyxZKsoHWRXtPZ0/MjS1/Va7eZgVIFVdCVXymYD94inhxjcPS9H5evqEh
htQMMjlsvP3ENiCMdq0+5oEj/bDT3Eq/nwy4/nCA7RUkhUg6nQOJyznjp1ZumW0P
nD4PZDeZwbomyNKrzLEmqemow5M4t0Z5WLKx5NMnGhMLL5B3F/PUyZG639uEIVXG
OTTzQ3w09+2H+R8zl6wJ6qGLXeKZ15q3deH1ROVMzmD6nzQ0s3FXhMGYoFX1yxdr
UFOT93MllDv/ZZGQCMW1IQQkrFEEJQ7TvlvmGPfgbsmTymkd/fpSaXpHOXVv2qfI
556+rlN9aa/P5n3pa4enxms07uSZlBbw3JorWOgdW48WFttGTqgkY4NYty1fqZq6
ZdBvXiTrjXd34HoAuF0EKENkNBJM6RhNknFyku1yb3cpZfXsR28qjuyQiep96sIo
Eypqfm8CNeEwossD4/W3F1w988bW1Nke0wiasXRo2trCsyWQpPOoX4seXVb0VYlH
CWIlynkDSbNVo4cBb2bSCmz51i0udn9iQIiFnksIdVeWzH1MF+hRkYjLudKQvjY4
jgwLyMfVqvJCUiVBJESVowo1YHlRmiMBeKHe2XvDg8GJPIEmpd/rTTmKnoiJduz+
8HR+FMp7ccWkNaJBxHYFzTooO27FzEq/+qlyI5cFB4ev1i0197CQG1OlqzrrBgqN
dq0Y7NeQabIFrpkkmSFK+zjnESOMaa/o3wWTI3oSlpbX9HTpIf2fwpzTBp4LjCPI
9NUu8tZh5gLJ/jBsS4Ldd10h3xXeeTf0jhfQK/E0LQ6n+MLV/xTmDJ5buA3EO+Gg
JujyCA30QeU6VzQ5ct/VCZiPGYe8kVWjj9K02EtdmnOSbSZZF+9Zpb4Ekl1/dAAx
RAB0N9uIJOUXkjF+2gEV8W8MRB9usLuWpDR1I8BzTEeEktYfq4D4C0N55T2Ik5P2
s25w+/6GMvrQTlj4Gnq/k1CC2cX5V9p3HPgtMim8zbeG3UZr2zx9uXFQBLp3eCQ1
JwFQ7ud8/cIAL79j7mka4tsl4IxULtJ8plUWhBc8VgumQewJSLIgjcdSNBGdZHUr
i7vsmWsbR2yBiZ+9C2rCRiCz/cyGCvveGSX+5rkq98xv6mDaV6JgjYYim0QOI3q1
R1jlWcny12ysKbvshRbzrEKVomJfIGPnad634YcLI/7HkhvudWXn+6FwnJeqQOe+
1Cnz+xtiZnKdtcxXWD2trOulLICN2SSIYrJrKgV6A01bE68f2EfV9D22gz3FvC59
2fnvZWqcfdoKZOGKT98ck6dQipLOEgztjQkqPcUVYduavBXlkrKKH2+pf8aEL0Iz
rmB8YTLrKbxfgTbmNQDT7xVv36z5467kxadUpQyhVS1bohkTXlcdk3jr0scRUa6k
ctBwvrg47mMkYpVw8PRtfCTVsVdAQY4avKY9sCuF/w1C7piVfLhzmrPrTvforcqv
iG1hUrCUKcivOFR3QjWCzwgGCX5v51RmZAvKRO01zsl1TXnlM9GXVcIbUlRGhLTd
idh3+SU3UJrJiqq4Da4SgnpNkaxfF2/Lkk30xAPDH+q4xjgZnm2f8tSTFfBYroSb
/cHo8SuEEcccx2RJRQc3ukAT0xFpRvWi2Fa4p433FQYNE2XW+hIihJbkt0c7fBL/
nLm4iJ7dF1zT5QGu5jMKBaV4xHxBlV9zf2Fv3wh6I2C3mMbUI438AfBZwgSn4qLp
JSwo78lb+QGw6OOJzNwzXqA31L47QGmwjo5d3Kma7hB//SQLUoe1SUTE9s9y5tZy
9IXo2yz0Tf5EZyhaFzMIGQ57M07vArug8zov5XyQGVyY6h0qG2+r10lryIUs5pk7
JSA5RadCTGxqv+AVcgrfZOcMpyn0GllupYQf8r1K6G9qng6SFP78AIQ8ce8BR1ke
+0aT/lSD5U+jAMhhMopCgCmfo8/lp0kZSslgpr/YWibbqCU3n9pOF+4r+BINhG3/
r/GRA91SA5L7wDVid2si0vR5d3LcfyXp2dzxcifx/mIJ+hbcvWWNrCpIsMH6LA79
HLgLz9SMxVcAkBWNdrhhE/mXSi9q2DqOV9pDa0QBU25VDC+/RXZS7raZZ3Eo/mPU
jZaHx/Zi4LILjqZZqg18GsjA9KLbqSyyyjBIc5TRMvrWFF9Xg37AR+7YFzTn9gSl
QV9vw20JUBGHHOEQF1ACv9J04KXZwwC8M027xMLwzAZkhdRO4hUF8kjddng/8QHr
y/XnYqDhWRs/gjibIRndgwe4vMrK6UhayhLLzfvhkNeMSlh9Bg8zenmaLHsSONiF
uT+66pOZyYjc6+zXV6j1WPp6D+w4ue11yrb4S3jh+XekXpbUT9tDcEykaiouQdAt
YCgS3VSg8FawBCHwu5WKbYey8Iij27o6wrKynu++lJBWugIu4yTTNyHwHEkOme+i
tP1NhPlCaZ432lgkcqiOeF1mvjh3R+88Tuu+ZakUHRCwM6fPsw/73EQtemVMA6r+
OVYzK6H+wbwSOeea6PQKp/J+otQri2Imk/Opr1H3ZCU/D8+KRyIrdT72Tbfh3iG8
VEdfknyIjtHDjwMZ3PigM43aKs5A+USAkaXm6NTPV5erstBqhClP7+3f/mTg/rz4
FXnu7cL0F1fAFOLeOvdTlkChGEtM7OEGC29c+UwEGR0WckJYW0yWAj2mQ/xw/HX3
WWcFulZ2xrFLAvbUFx9d9BY5xaI+4MvCEKbYmFcTph5UaPqC9Svdr4Cl62VfkWZ0
FarF2/cJBW7BhUsF2T/iUytegUFA2HeTYjgOx75YVCm6PGAThPsxw2Ipe+bX5+tY
ZK529lbIygEGYor2+q/12z5IHwnemQEINu8Ru1UaIUknQClVj6NsTImoawewmPkC
hzY1GYgoz7AXuQl+vZmMQpvwQWXIf410MW39MoKTh1AslDLP0RGHPJNBF3n64lq+
a0ZOQzzKFA/m1H3vSXx9jofFqrFxGBff6iVckZaaNNBOb2f+PwpK+KtL9CMbcAp1
97/Z6+xL52fyWcCcisNiRU0kyVO3B2oto0bs0N5uK1oe6JvcxTKNOGFeiOBCeAA1
6d3io58FX5n5TDRyPCQnzA0PeJDNnAngAcomHnLkmCVX9JRohhwf7f6Cdj/lorrq
6cYTl9LQVBECMm1tTG4i0PXFJsYH8r4zeY9HVWb70Fu2n037Stk8jpw8KDByfbb1
GREVXmaXPPocag5QuYQgQiBx/Ubrf3t/xLF0XSS2dJ7aENKVjKQIUvrtmXCgit3u
zQxzKtKtvMJGRsjrv5+jk4Dq/nGeUqyraTV7DlwanCtKHeZK3NHXCGOXXfOpxd7G
DD5XloXuEGtPNYKJW4cG4y+7ynovn8yru6J3v1DmVbkam5HIQQzDQRzz0/9cpgnJ
ZUjUXxqwOpHcjX3kP0bY6G4Y+fTGeRJH4yicBYO4inNqY/6HTcMTmY5ZSh7tgiNW
ok5TZltet2z56VuEEqIe3yHaYsddD4RgRaTf6HPvP7DGOWM4S+ufDdZLTqhIMJsJ
TswzM+bi7+CSeCHuxzD3NgM8iV70o5MJqjQCCXuPeC5sQLIEQcU8FBWUCSxmGl7T
JeX7WpQrGmYyShl+B/59swo7Ot9L4A2hWyxYnXuyfydLmzFnqffV5/+Km3wjN2ql
GnBXnipcFYHO5bmmlYTHA3tUsRwvxYc6sGu2XIHqnidc2RY1lAt//i3yTSnRNvJX
ZRy45ZPCDqKTr+x5SpF6KznyMOHXVSpu4wVZhPa7CWBkFLBfjn991kO8d78MdhgK
FJ+3vCPdCRPX5MbaU6A2D3hCvOmkLrgBRL92WdO9mq+KN4Fp/IUWQwe7QHgv4qiA
4HRCH7aIv3IgERtgCkEIwHQNsuksSRfiWH3uMt18ifPMZge96PS5pl/uZZvIAgMo
YxAdAM1VoMFJUfV12C8M9CNLrD5HwZXNyOErsB23NGjvI75Kp0NW6hxgi6IiGbyx
FZDcmLfGitO1b+uxJI9n7nQUDaSQvRoIrnKlPZV0Np2U5fFYFqaCSfguWNbPrdSM
WHJqmOSTN4rf3I14+XKnuPhQhGl8LtS8P455Oe2Giaq5Jkj0/8cWj7jLXGK/QAPZ
bKN87jVQsgcl6rCMH1VQ1X4CvZPPQT+M2R1/Y7NL9P3rTLdq3/4EfNi/ZigOsEuF
bgZAHZEJaX/62vMaWjz3wLq3LQ2ccLG7QetXxCKR32zqY7wWHHC1e2v+mufHG+1X
sCdgwOynbdDAQo1hMcBK6eUDJkEi4KdKIWvkdFpyCv1stlFLuQiEvP186ftG3ETT
6oXC24LrCnvqMeKyiLC8/yEOYZbxcGqFX81qk4XC7Zjx8pskiY4cUdApOCRLAsn0
IbW+0iRg/POYh1p+1H4vvc2hMYbhlpT207v9+lz35eXqPN5FU9L16f8Q28cSWWH6
Ffbodxo6jMmm0jZK8GmPVMHSJeJBlTcAm1Pk3nNqdWKLp8nA9FXhVFTwkqhE+M0U
vRZuo6g4ygLtSSUfhyTg9xao5f+xjXJUqNABhByUjGkKwKW/Fk0Wi5YbmsXT9j7e
4AuP1Q4uVaVb43DMB+CqjpNA+3tzma9V34QZJWXLremdcLxufwOUwbzHgM9Xx06r
iG0Jik12IJyMQ7Aqm/ZfDEG7OVZcP1uBentxeO8vSxkU8WAJKON8wxKaKvFtvp57
KcIZx0ilB0mXNhzSm8uJY+1/YQgSc1y4SrHuEyuEe2sPi4aB8VCFs32sVyYkYZvW
I4nxVR05BBdVXQSflfCYYEREWx82Tau7059ChIMG5hiNvU5WPYgXGrCaq6dKjbYr
L0dL2Fn65jZYKfpQWSQ6go2Jc8Zp8KlCKzu+5pf4yLYjoi8/wIalyPy7ys8ACR/+
s6aa7PlKm/Tt70ZMoGw65+esb52QoQ1VfFbORJCwSQf6G3QhqSD9dk4tBcZq0tJG
JQYRiA0vpERVFDXe6yALVm2l/Q84Xn+QhLAuoawgIVvIOFDquR9DHHdnpn0xvIBC
1C3q2+QimzTY1RmQrh/05goRqt1UQ2YvcFO/3FJDjE04LVxipJoCWQu5DqCuOGWb
Drwoojqgnqqbu75Qg8GAEoyy5PEx2+5vI1558NX8YaToywmIKZBmRl55K3x/DmG+
1WCcP94slIDD0fcGOTV1ZvbUxEZoXs6ZGjvBO6g+4jM3NUvsHnF2jERK7vSGz4uF
7g2fr+owBJ4ruvj4v6g9FGUyLWaH0QYdGcom2kmTpO/lTJdLsr56V5EiicCX/Qw9
CguaGOeFR+OXtgQi4XCEWXqstiEwIwP8/9Pwfr3KQLO1834ZAw0u4MYTGRi7zrB8
AxnoocZAnuJupnqPdIbuG5XFqrztRvYv29sztiQYTot3/foEomDKzWNbR0wqIgnc
OyTkSVut1vu58rS1oictt4o9gApPSc1V4J70YXSxul52ZlzwMiT0MOf5heiZto3r
FlM22Dxo4mMSqbIkymaGxwq4aZO/WMyoa7mHgyOD2dkfuzcKzqPQoHB3buGhnVgd
zXnGHLcRnzOpn8Dsqz4FIDPHD4ZRJVAfz+lOEkKnqK2lNmc+WUzR2Bz0m87UfS14
2tzbGbz5Rv3DhOpn0uFk3ziyuDTZjqbsGwp9fuauJ+9Z64mAmHYRYdFNhtBi2n2k
Os604k4QClnB5uJ0GubZAfj2AXuMN+sRuzxAGX2ncNOlQ3JwJMH8Vy+Oug/NicOc
fHuGXcY9U3vVCs7kl2HK+fMImzdMDY1RdJaQr016FSj3Iihw7FCd1xXg4ehfKt5G
7haaCtTfO+Pa+YEEGohGq0Td1cZhN02aNHON3czCnAnUeockzrRK6BLU9sq52GCz
MZROP6MwIhzNcJMhDwpoNa4gdLLHo4kQCqQHEKvuY3cv/8cppeZidD01qmYTRmlZ
ftsmqNKByFYIdwR/y7wtCSh5ZHHDimUCt1xc1n96oTrp6rKaETpgZFNZqW3oe4I4
M7yN22vodg1i2jBzrnU+gb7f1CZo4uoapOcSw55d8itmQ4MPmmWmCr1qmk1V/8Tt
gapeDiEm4+wFUJZ2s1XwEReIRusgxUKcqo2IXzUjh31Q7F5loPxma+RHg0Q6SpTx
s/fj1bFteJ4IDjip63Ftv2n6j5bH9wMuWMe3YqVyxD8SbgGV7w3PRM5iiBkya0Vb
2HIi7wvSHcRU7h10HXFnKgssLGOcKDFpNT37d4TdNwNGv4Dmc2fQZcvhEJAICNVv
goXYZqz5ILBQfIzbgDvj21ajm2c1nJYjK+JpYLmggbtkHlUFJqntUhqcmxM+Jvsx
Bb4XWDSKydnakiN2NALB/3PterjHQqQx4BE9HRMpJqpgnqI+E99GszYi54XkNeb/
A7Ez9pVYKdgqzbUbS/Xtqot3p+Vf/ocbYcagqVexm9H5nZvqmq7blkism/JEUX+p
KMROW/4MtlFdoHKlpLDz188tx163/c0erpCybZWi9bb20Re6dsha39tEN95mP1oA
NWcHHdYYMRU5mBXXo4lJUrhKrZaIyaJW3O1UagW9MatkHj7DTdw+ZwEYpDklPu1t
ujK9rZqSpyg+149SNr8FQ+XthnFe4k+EUl08/uiubB65Wl9Hyfm09IYHSD5sHLcy
V7aFZXecSRisrAhwtkfdyLcD6nGwPJft9ESa/mpo4x6Wp+cUJ0ZAD9JTS71zNl7G
KEGPmUzfoarJYcrijeLqIRTEhHy37FAVt3KHG+V36dxSN/cLAYZP7ONJPZxK5neW
dmkqYU6mOXwgKND280fNRSEw6AbIEP5r8bky9dx/pBqkGz0tuzWMM7ZPfUItGraY
E+qqrSh93teOi99U+JrvsXKRA19QcdiVNBe3zLDnWePCWaxLVxes1M8aGn140JxS
KK4CdrB1twCulSr5J2Dh5V9lYnMmtyJpr35yx/KKswtdFcwsrGv4sOeBXZAJp7it
yqyIqFk24BhuzXLb/XbHcY/+FuXeKxyWcCU8Y0IWvDa7d/yIspp5GUWcESLI+qcg
17w5op15CXKYgFP+kRwiyvZHWxDBgXnFRZOmFswUnQJV6vMJErlopxhKfc8+0tlQ
bd51ZjLcDdvQqW19yJgjrQW57eb8weQREeQrLYORuomczwaHk1ORc+zs8+coxpg5
NSiICXWpIRRwtlTdG9SMbDgZvC6Odhkb+wj/RiO8lq0bT8M0e7KI58eXrjklE6fo
i/D0WrESiN2bY4VzD1tbcRdXfRzP2lkk51Lm1M4s8sJSUyHAgrxDgy5AiOpq5Dzl
RdThukbl3OaGgCUaXRw7t57R+yF3tlM9E+MYx/ZIoKh7GDP32qBPuiO6zKC7JWGO
CMMIK5vmSCyaDlJ9kEgsYImnBHiP5ubewf6xw95XqP1Af0Z0NeWBAzdfFm48se+f
NN5YPqlHKg97IJyEokUEKXxX5IzTJJoZbN0vqhPoGZLyqPu/X4WE+7FiODNfTYde
E6fRPI29j/+EU554sRXsnazucTZ7RuLtx5dL84PTjobjUspE0OE3U+gZeSfOUC4W
7HtfNw7SxIa2CVU98IgxO2SAkcESY3crvro7ZCCu+LQQT9xd22LC1S3XKKBR8pEv
S6wu6ZCS2zFdQzdn/MtYgKjKqB35iw4KGcEeAEbpnMPLbh7YXv+tzPZn0Tszzgg6
upU+TXqvXUMpbWkhUXx1XUtsodVZAZIEuscFMEcJNzZUMPjWZ4gvAtVZxTGoPbPe
xSTpRbr43+IHVawk4bfuPodWco1LEK0a9rh2nWsuAusyNjFkgXfFATTTp+UuJV8O
AfW6qvMwSoN1WgOYNybJMga3rRhnnDtUWqAAIP1VnfSC3mhs7jJurhW3tqn96Fhm
9fq8GaGWZkBw5sgJ94VZdDG2Appi07L53I038rh+uWr/hGB3etVO/Ys4Hqenuhil
OOBOb8WuVZE+9RK6LDHq2cxEk3SFI9ig69jxfJhKUPkAcWeumx0LjTvfUYJrSCSs
s1xq4802cQV9RkpDXmJx/pKF3/pzv2/6jLc/JW3lSXUrjJ0yLFCmTt1lSx4Cr5Vl
gF/P3Zn1F8Kfj9K4sjRImu3W7HJ2tg4z1iinMDHv4z++3aVPf5TJeIfftIsaK0yv
oNmEP/dXe9XOxhctBK2jLivKvIYPZ53UwwZyvYvDRga/9tAjsDzg97hdEowQn1xN
h+OWAXB/vTn6MK5xPXVOLhvBCCTmsdSDQnPW/2kELiZiR7h5SPlWGpI5WSRYJ80N
ALOfdlsvDdTDB93PF1TwbGRFHmKhcwclnjv9xIXoVpc16d5VES3LZybBC3vSF/sJ
K8mOWn57YjGO4xC5RNa9Zet7TgsmppqAa7/t6+u0UquUTbh3b0N3+4TrB/Htpuii
QC2Obuh8bOkMTaobdXFh0N9SCVnc6vjF/c/ORuEhAqXyPjwUpI1w6YKq094fZqX/
hpF7ZHkUVpPAWKOOgufWcvTpBZjujQoBucacJkmUPuiSyKZcccxjy+Vl8JsO3J8z
gBkB7AxjlMVAI3wKcYJIidFdhLsyPVj67ZhJZbaVdWxtWXOhLjHP0p15i+UkBKYe
szEHvjra+KtaKZrm4MMAFeAS6x+KDWYWTxu6tKi8mAVUWM5JpNCz11UDIMEr8hoY
J/wF/1mdzXw+Fyqlielz71iRUlxnlzFaW6aRqNJ2RsJr89njVz0W31fVxNchFZ7M
rPQrCiFSJCx3BqZrxOkrPcaYjuHT+FM6o82BKjNDyoD+zgQ5B8r5+W/xskHsAd+o
zj7vhgeisDrIGVtY2jLQ71zLPitMFmdaHxlrQLKepJEpmft9+Qrq9gjZxsNHclX6
xRFx4rWhaloQP+OFCcIchFLAVBslhX8arLgMXPfltMZ+c0l2iwolqN75xEFTG/+x
GFR1Yl96HTUTDg41etBHdLylNyMHgXvHp09M1FQ67BUc/yf1jmN/677S3WUdGOtK
WcoMnZNF8NUHhRjgM+Ldl/Jrf9dB2IWmJszBWHto7Ggnbr3U9f/lcOjX8H7A4Cq+
PWPrK/k80YHJq+wbMymynrCxj5hnuavd+8KZRmBeSS30Dspf1QWLatFqZLVeZYWb
BCl2GG5oo4xt7KcfqD9Y3Cms9jZ4oAsrFzYY3EgXBjkoRQwi0x9T4+jgKCS8usbo
DhU8whY+CAdB3lqOzBWkI77Da3t+xDj1mkHWWMNFxPs1aeiNLrV905Ucqo/rQVOn
E8yWFks/niqX60WJGVso3/+388JirMcxQTST2FshBpI5XWpZGpfAV4zoc/aatrK/
eZYHcSzy/GoKDlW46FOTHjNjA0qmsK/uvrq0oyOpXpFzbrWPC61G2Q+VuXiLKm4A
hfXo9WAB2RnBaCYRVPqQVVhOG7W8qg9wJyuJSDfH7eb5btM8yFY/l7m7ag9w+51+
KgDldc5g6ExRTyxwHCgxuYtC+U3oiayyecdFoud8UaSFAt/A5dLioVxA3jtk7EsK
Nv5u9K5MkwX9aNYvQrd4EBNpRGp4ksgrzzybiN73KXIGiif+EkCYHmQJwPF0kOJa
rs3ibdjtJJ7BlHwHDfBz3ZIWqGLSC7+PohYRV/i7VXVsUGGJwpT3T3yQCa8KQt7Q
LYaXAsCrpJ0rUI2vI0v80eofPe6gpRIFQwBN4ONa8phCYvIw3M6Rj/E9kiOJoy7V
HyQ4nQDfGK8X+ywqH/b2/VQBZywUnyiMt6Q62z/LtQKVC9vy8OO6FbmfmRlK/LgN
A2IPtpAgG8ODvBNjKKz8ZGTzeXrlxO6BspUZwSejHUhRjD2ilBjUcUHU2Ua9BdKS
uwuAo6E4aTHKPRF1X5jLeF5rKYUEkH20/l2F0Dk1iPUEabHXwMo6zqBDATALv0+y
4ZRWcSskG7TBjvjUsR/rnDJgjbl+3XYFTA6CbEQr2Ub26Kd1bOCEkhCDBh0DMBlB
PBWzrsUkDeslcfVj1Z6lnic2syjO5+H0nqKz0yFB+Nd+sg3r51p5oBSuRdSKhhtj
uv1oCV9tfkfG3G4SV2HnM4PgJDwsdO2edc/0Qtto52g3gVf+ZchfLSUMmX3ArryB
EToxu+YU6rPWz9Rnl6iVgprQnuM0ZXU9GP/8breJMx78cfaIS387p8ylxK019fb3
PIYmfsrb5y/kec9cg2MBSL41fhl/5UxEqGf8YGZBKXiIMWFJ/NltLSBABSW8+u6F
Xl4bVM0FniVldzkmsxDVNdQOn00a9w5129xX789j3L+QifmNx0UhD2EwIrS3xO0K
HF8aSJSDzT5tHON+EsP46LomD8jHvQIr3qfDTG+O9VIJb39ulLHRGUMJxJeWzSN1
REcc6r5XN7XnST4A3v3A6ocEGoGkZKF8FtTZEgvg7QcwGFlyOPZS37qbAcowJ1s/
1IJv7U4vEGvw739TrIDK5PyZXzICjgDItnTALg4wAbhodzcqCXDqZ7PyYdohRH7o
f1IYZx8z6pTU92h2xOeX4K8JGavgXVMpzWBVwIdJxqPU4sb5F2DYyYdsISA8kqa9
QVyKkrDzjD+MzfMX7gNP8Ob+qNRrK3ILQDmrF7H26W2S6X1FEbOCw3orBOAFuccA
GZKARejUaB1bqGnpfS2f3Wppc3O10phSx9tSBxF0LcxpPjqRlEElmpuv/6j1a/9z
yXMHjYJx+w9A7zEkXtNetRgy8AUUJm/NPqTgiXkxR4ml5noYChR/jEz1RAVXBW5v
vbU02sxWmrfW0R5k7GMWBMlxI2QNDU4wv8Yqe7v5xFXsMhW10yr2Xn7OKpJXRSUo
hp/XOaUgSbt/k68fvrWJioc6GNJPKmmEjr4wRujkFcbXbNsyYJhFYEChXUBg7ssW
r6hFNr5yIVDRH87vyvaroTh0IGRsBKtisZAz3kUjLz/FiJyr5FmZ2LWV0bQOUum8
Q6k+8qVZK1fA7mf7Gqfy/yH6Ll+BR/Kq6qt+GNLgorKBEz3P2xQvc9KgUOp0xbGh
fwlnWf0RSsFTvPLhsQ7y2j0BaV1qRvF17hPPFu1SZC0UdoD7mJ29BX/KCHiM6nXE
nGhyuhT/lOKmIJIloMk2u7Ueya1yvNPXz3oAaZggE7bQ6ZwTkqdNRZwk4XDmJyl3
xaq+KSW/t2Mv3g/TuRaFHRaGlx4Vdqcg8htg6OEzj0btc9BaPBncTS0k60anIYrc
1XEx6qNSeaz68kJZDPxsIDcmfMUBqo/7CY3y/2LrSbuYZSPFUUCXSs2gj1igFcUG
4iTWEbMpAf1b3izYOhmG5t7QHs5CnuX3CZSft9t1UHt2ggHc3pTkQXZHemLTTdRY
EcRo+7VOwXhcy15RL7Sm4W7D5UeTG6Hcp/+JsUp3YgBYcv32K8YiYOSoMnhTJOx9
VKYBh6jhuAxTnfuE/bHPiXOLq61FrWPrQP/DQU9LUF1X2j6hgPQPVs9xFO3B+cEf
fT24p9qfJbZVJIP4fqhIxQHwreykpAIuZUqdRENeDzq1q3wh1hBdJ909bUyTE9EN
XetmqtsbzwbeuL1mZ+HbdeQ5t3mRhTn7/Ftojp68IdOhyKM0/+BrSNsZMt9Zc5RO
OD9qlwNlfj/beWs1MoTQ8fg0ipf3ZBr7CS/e25kOmIrYfZaxbpOvgflGeCVnb+lx
/yzGGOTn47nGUk78+CELlUIF6JsXORT7j7FEbO2b6LW7gVpRDv/JcvW7lxCMFlIo
6fEc2h7gjNf9Mw0FIva9/gLiHcsf9/ayeR5v1i7uryKgW8eAuOpqN0YDCEu1z96s
426Bu5783cUC3fCfXLPZTqDsqSSXP1rsLzDIZl4t/o0oHp5l1HxWP/PNYDX6Ykb1
tALcY6tMt0OXAvchbTzvbqd/IcTa5j50giNv+097bQ4E3ynw8kfMJAw361RS/C60
rMslsvANzu9d8topR878C775QZrSYvGrBkm6dC4nx2lntwRNAX0fLMMzthNqLJgn
+hGeNvbVoEfhxhjAI1xpLOi1EXFxqIn4zVr4IuuDt5ZodBkrJcGDcfX9mu7u0tJ8
y8yLAjvllCeDbWvJ69zEfZUr9ZylgcoSZ0BA4+O7vDtVrmWwGnRg3iDH0Ok0uSG3
7gKtCiJHdkxGnJojvU52ecVjL92Z9XYcTlRULhpLdvakWV845CktZrJdB+YVf0Dh
npQhYeZ+FCz+m2U3uMgTLnD+x2q2NPHsql2ebOlCTqndpffadKauhQIpf7wvtoye
uE07WMfCkp79D2EqtTWXResOxYWmQFiP9J+DPPmFmdi0MGiZSMqIlv6T+ZNUQEO6
Xt4szd4pqT2upyvj71gpZZ/WqGb0LDntIfEX5+5CS1xQoOiZN1DgK/KwuPyqrag4
DiYJMkaHUXvSMdOdx/L0LqqJxr5wSDTOH/EdHzhog4l49X4MPeXOSICdELUaUCCb
z53MRFYomPMmJ2rsuxgUyD+ThNiJ9422cN0h48OSEhl7QuX59Y6ai4vQFf/htRl6
LbIEkl6rpGbhOpEBo6a0auKTGJQTVshXavxcGc3W7BmdN4QUxWm2P9SiXk7PlHGV
+KekRrkFeRRXNm0U+CV1I+mw5P/Flo/NHLRBo6cRxJEG21RWuWWbIZe9qWojdG6b
doXQi70NtP9M0yOcRfUCaf46g5G/q6jI+esBq4IDG9V1WCArx3kBi4rR4kM9RRRi
NlF7iXcUfWUb7X57wRKqgT/cCyftdPKD2KDotrMlKmc7hH02rDH5V4sYF6VduM2f
t8CS3+JrbU4JuclQTR9sXcSSxiYwAdAXNBOh8m2Jh1QcJs8wj2xsPGGlqQsA5JP7
b60qYPJxcr3rTO4gc9omlJjkXgD478tzjnunFV3SVNE3KcnWgiiMmUa/hfbqdrmr
K9iRabScOfkrdvvXfMbzpJSgxLBaAHEXSWVbRPVe1LJ5iVK4D3lhewvvwMcpQXqP
Ki7Yrgb+DMqNtLLvBrWj6UEPH8E21jv53Y8uudZHar0h8d3ObS1AHfQ9ipnYWcty
zwJiEVAEm5AJMmhPkQHi6zRYnJx9eDzs/QAZNnC+c+622UfCb3x0uyCGYHrhSDmm
juFU/XoKfg/3abURkoeKAPHkZW7rp7+R78PJMNzeFvcmxscOiFptjU+iL5hIndL5
anDDdx/iM2ysGZPW6t7LzLnVqIAGkr+ihDk3xLxbjx9TtpkbxRW+3GkXBtPYfXF5
i44mWkPK4LL/ZEXlrzqEEuCqt6Mg2sUJc2nfhnmvexeV7VDYx3XTRGZZM0JAX7E2
TcqmCEZziuzFoaH5xh2W9rNj0lIiHhL9kN/sUEQXdCXgv/LZVwLsjyQn3rtjMOZz
OCZVH6cxk1wokUqrzcU/4oZjL9YXVkpm5yHe6xZgKOB0fRlEThOhn44sfYPNV80m
6ETXNMopiaKzubAElMZvYGtHUXZAcxp+dXQjChbn/Cyh/viLqus61v1Wp92UMEqz
aYUrBmAdnjnOd4+d+UK+Do2Se8QHaKR5pHR2fgq2dWl6nQp4MM1poUxMfE3U2KEM
pY4PxUe4zVs4z3VdX/IyBnHr6RrsRC07sdoUAde2prpM8S1JbDbaO9QcGzfVsMn3
IJhc3RAeYLhOvCedb9ilZ7jwQDWlFnb3RC9iIo3yVFvWRqSBJ6LkxJxFjT2tcCuU
m/nmP0rfKgzpb7TJZfrGu4bfEKXWYZwXDop0QiX26EajfJVFq5DK3qPxwHVepruN
BLf0pwe2nVGv/f4jzyBJ+yDOq0CkpuTElXCmQT2DDntffuwP4+ejUmE8wHlWirfE
RgPDknZ+auKXF9HKCOrFi244hpnGAYINOopJbyz59iAiXbaDV9ePazMWRJpGSoi1
IlyUEYyE+us0hVWFlp9T020WzXHlkHhgrpy5TDC4W5A9nnH1OFeqlX00pa6YZe+y
I9C/TUZ0NRF79ZdtPP0qHoz2oa1us0vFgKWbwttSMUz1m4YR4jWewtlCnmsLtUPC
rxZROoMIWSHifrQwEDBwbQ2ghjSO1je8er3tGEOVgaMQyfBOQ/kQ46amz4rlNS4i
UTvdlwbw1mYhpay3M0T+qpJCUnP0aFIFDxIxEDnXy9Nj48ntbszhvSqw5IXgNrIk
qeqwxUfIECcgOTTGpPPu8OSATLulqLbCBMkdcNfxY9cH76fN1Sl5nfR6upekvWWp
/CVrkvpMTjbFOgQgMUrQ6A8PLogXaEftBqsS2IxKvIGC7uUNgz9KLbuDPDZMgcZf
42XzkneqvGseNGyfx3EXm9Q484Yg7E5Kf5dkrrRDJIYOKWH8xnP41w4Ex6pZT+VK
v+d3VI3/bLI731g2wPhqLLepxTa0whBRhrYJcl9BiD2kIPnmgtHb88Cok77pOIWB
14n0wux+hRPCWCCjNXIlTAkaUnh+agGtA3RABEWHzICGqT5bKq9ToCUlrsBzdRkI
vezI/NJYssz6rbajB95rxAxZPAiLwU28PKppdPJTL5BfmkcnL3W25tKwBSwxfF7v
HI/aPkcWzPQvpEygqjI9sqzI5596PO9puvgZc2YD7SBz2RZR8auGChVfuO03W8Oo
NvM8If1aQDJJQMoqfgi2wUQxKsSNdfieWTfZcumL2HjctrD+G0GZzkd/cxETF/gl
b1Bc/7dKKuLIYeF+g3sqcVX3OinyKDWRurnWHwNGuFh8WKxO42H/Ofgkem6t/sV0
fRQjKuSTdWjxfg/1da0rxBOAJC0qrmAEWL75UIejZWT7wwR4agmfUnTjNFa/OSPm
Ak0an6JESaJuFQxKnVvlQ3j35OiYGljDNHY+DOnn1gkb2f8YNul/Wh9q0GWxJOrv
dw4rSsZV8vuzTjUDq46WR/J9WotzADsW0l7Q2cdpDunBx3JIMroBNU9dclkISGuv
cWty6IywiIcLpMNaaoIfCzz3o1NnxEMJzHvXdwgTctzwmJC4fwdr1c5qa484GfDN
Pftki1njAyCWOTD2OKI385x1IOG+Xp5nLI7bO7WVfhHcfQbl9n4SRG/4NUE3cniz
sK9Zfrkt6DSPVjNHUBNdcH+dPxmh7quy/InEjzXdYpRU+iDhB5dcj0ycoynfF/ol
WYqhyzmvMRMYhOKHhDQiYYLKIWYahhlB4m0fDwFaSWzOlSGAjvU2V9yKJWsyox8B
5yidpJSHkkk9yA0XCq/KujNkQ9mi5agOxliPBw/fm8hDJ4Ov+eYfytof9i47UZJ6
gqgKM3h5jax84SVg3YMKV7V11V6zgFiSouxngivqw5COc4LW7DNSjMAV2FPhCc6I
xP/NFDkC8V3jxvDQw/xuoGDECIB9B7zbBCgpFP3PDycdFVTxTAfz0uKjxT9kgCkb
zRxqtRmmz0vOnTwN0V3diW6kci9hp++JgWCE7mkpTND6tYFoRRvQN3AMMJT23tJZ
Xs2C4nuZro59P2ze4x0p/17a90h1kgp2ppk6sydsTrmLZWneRCF5um/Fq4Chexm1
2QtVVQJj1VHkncihXxt5o2FDGA04xn1IfUdPK0Q4F5wIxrNn8hMPPbN0hSGz0ktR
z3r5LoEvC7l/PSxNZ3DTn7O9AHiprtizIxkaqO+kwVaRc2Gz1FOIE7Ii7vrfeAJL
l0ByA79gsE7FAx5cj/X12oEzl9hFd4sEbTxYMyjC96aQBvIcuDAvolFJfJccR1eT
gU/t0NUozVZ0i9nnab2uoUBD2U1I2kV3yPgxL6D+e4+odGp8FFy9cN6kLhap7Y9c
MRKJ2WpQEl7E20oogLPMFqN+w52SvB//yg6ian8oB/46z2G3T50Ygbxadsnn7eW9
qn+YO3BTErI48mLW/3m3t2TyECmh4eiusCSOUyyH0KTl3E8WvSokXpu9UD/c2iAz
lukMoWYXDCuZyUVJuVv9VaIGfp3aiA2Hhc1DjsZvjb+ZykEUdRi8TzZRZqggIc8x
lz3oDbs4eNrVddZje4Ab44TG4ue3a9IezRYmHUMjDvYF0nHZvFhrV3zyVY51IUKn
EXJ2kY+w81PppKS3lO7gA5x6hDchV5GYR5tobVDLmIzi873Q3n7kitqmMEExohJ2
6XJWAvj9wNyS0eesHjXxQf340Vo6KId18BgXOrudMYX4btKxAP9BbcdOQuqiP/BN
sAVLb2xPo8H2ZMhwkMeQ+GC6lUDnBqyLJdYoAAZsI45yJTEhOw81D4vMKUjnWezf
F2EUuAq4uL9cBepiM5vG83M9kYEPwcpSDXqebkckqOZvOCMvuwOQSFcPAda5PV7X
WrGi8+g3qBXmp0+bKaZlm85JbrOk97K9hFeWw7FA+O7naegchxI9cLGK8TAlJTUU
vlci4MZ7PUdGWXXiiAN5pcwVs4cN+jH+3XNQUVbmgmqDHzBsOoBk8wo4wcMyrujs
mvUOpPEf3u1i+QxaWafxSwhvefPPbrG3dhdER7nhr+/fMdHRwP7jdJKALMrDGtR5
ajY6M1ihcA6yOEXWQOMo7c6koX6OGAy/nF6UNZkGZPssKyGVNZ2lZQpH7bIVilcj
sLfqNqY1q+v7HVl2HM4vq6Dws/++kF4p6Fgtc6fKsOyN/n42lGQJmMN9MMjWnv4x
LYnUMpAovMTApBvIt6o8h66f9EmQ/12cJHI8mIPTlvnYn92eWwN7n7xkZfjCcPJa
X1inLD/gs9VKOPVlg+rz7FuNkmnk1ZzOrhNJvYZpe5hmS3jihOwHh5MWAaEAFEHu
7ubujazKKp2SYSoD/A+BRJ0FYI+MeTIgnJEi+0Le6CqhG1knJ8TK/S1x1gwzT5OP
Va/5Jnml5bXRoMmewXdXrrTFldZRpAxDqQgY38ONTLNfqw7yzYpE3ZNJ0YWwQybu
u7e/Ay6z1PBcvixoVhbn4s7NxPvIxHvUyYgSrNcsbcgtcnNt0T3yOZcQODZagnWy
5ZdbHkuSsnO9q+oYroG1ElR2/pgBiuYBOpIHoqz+vucRv+ukmQX9JL46goXl1ov/
Vr1QjdsgNRUdbzE2izKs6QqJrMtL4PW7JmmVpXTzUzwUeIn03F8clxeVNXaEV02I
bFDUEkQOfEJUUeUkPyXWmcAtplROIwgSZX3ddVoLsTV8vovH3/T5ngQiU+MZXurC
gFxyS90A8NH+2qqUi+EdY/Uf/B5b5tG+Q/dw7weJvCk6ajQ2OPNwu0iVw7DtblGt
jgpZeobDYMhPfD2Uw1UT4u9NCFLjSinWP5eq6ds2PONQLQdYeEP1TmMZ/+CnGH9K
M/w4SuAPMTrOXNLYZzfNo0yofLy4ReijUtxbFv97aw8J8Ma0X8YvAawYFtIsy3n1
GVK3IxJnzZ5d6xIAlmwDD6/rcEjRSFwc9xI+58l+dQuOUIgn6TrlxYdlSCrQiNQ4
B+quF81jEe/+cw0mxIsoaevUPqpTJBW3acDz5BTchx5U36WybcqIgjKqJXM2CC3f
rWz2lleAFc4hEV2bpUn+nen1K4r4omXeRt8wGtP2Ff7WTWnknfMVs5tTN8TUe+9m
Y8ufsuuaVGwrEXub1/SNho3OKlWBEstidpuaJKFKhy64CXORxkAvgwn927qfOdIj
SJ/KqYIYxmcAetv9vU7E/T2iW3W7kAEAMD4baV4BgdV+ctVnDxRGN+2eySQkgIsF
DEmDRPwuoJ7HJE4DnU6fj5kEOgRC9rD7cHHQlxzHGj31LK3aSyGa2vw4rjnhqJ5T
JE/LHGy0jiGWu9zrsv0hu7KCeecaNSOQqRU6klSCnVYEpYlFaf+FoYI9qzDiUmsj
NJAptIPqPy4QXUY9sz6p1I4/avC+OMRR2kWcQt0PTZw8+E8eb/psCG8ZqWPmgWNi
YgGB/jiKOvdqYw0Ulblua33nUPyDHz3jt2jStiD3EgPAw1+cEw6SSIXrrvAss3SM
8tVw9fwtmm2Ljwc+Zn11owdFsVdvfNyzunogiPqw/Ntcx25nXBEWKWK04JnQlHuL
y5BjCOu19gCxihZvny8Ten9uMuYRWESxxXU8pqrL1LYULG2mOweo/abY34/qhvpn
uMYJvGRLhQ2UZKHNk12yYVc1JJIw0WZAuElVW2KeMWpTnzTlo7O50yp0Fjhcty/C
flYpI8fD98x7UNqqLiaTTCz45yn4rtgPfW64vaHzw4q/AjL32CSN7kNWINtU2ZFm
8ziO33eMVBY5U9KFkeuQeYQbigA+hY/ixMdHPdMpoo4YVN25Ds4ztBcX8vRR0vOp
E0Mb/x+F8pvUBrAoZUhY8JYIbU0V/6LaevUEHHuV3q/jgW3BjWe53zKyFKGrJgz4
QuGddO5rlwH0AiS+8N2F1ayYDeF1HtsyDBEqdKqow8OYGE3gvJENtlSGAm/8pBB0
Owe0WWisgLyueW0mPXDNwigGRzstaVdplUeIlaX50NCpvhaBsbbIEyPW5RPr/ag8
jo6zBSksa3HGfCXKH7H2mp7yFy0aVYbQ3IxEbH9R2g/f9dCUExlymuKeXeT84bsv
HtkIjBwxi3CbLZb6wJpNFcurrN0/Oj6gpi25im9O+5AD1OkAaBWJZYpqcUzMgF/M
mlfx3qBADPoLB1T6YzG3ultBCahJGKN0L12IdUTihq+Q+zhRWPNDVuuG14/QyenT
2smFBkK/oADfeosdJEh6BWlbz7vDLw2W/+VtAEcWllw+Je2pkLZJs18JN85b39pA
NjiB0U80OWDE8W3HSXXI1ZgsRncw9wdqYbJhT4YKJ2KAWPWA8Y/gT/dfgTyQC2Br
Hcl8uY7EQ811EILqkHDIRxIUCq3qEMZLYBaKwQt/RiQTGx0ITIXZXFIdAB+a44kx
BLGGTk1fVlVbF7s6u48/X4X3v7AkBfWsjAT13TupvHJahJcM40LGwBfLwVg3sz+p
TWUazupUP3XaNtmRcVJZMHXJfjm88C7MhIsczL5Gv6KLEWVWZ6sjYmDteqOZqTAz
hLd/8/6ip6qmJIjK71RaYsTpYSlcsoU8do4cG9aGIMkD4mOuK9IUdbOKhBVnigu2
YGSQBcKjYSokBRDZYLZ09v7spD91QAeIVwQVeb/bydabdD2mDmdYL5XeHJfmV9QX
Ao7WYaHPC96bIF07oeNAR+Q61b9heFQwsGidYDOFZ+4RJGcQvtwfjuFSGbfOqKO5
pgq4id8hYJx9sWN6fM9W6/T5Ia+zbwT/rbDBCvMtcZG9v6lNit5pTwATpwG+b1AS
2efd131kw+BL4gmcSYxWL3O+sMS7A2jW00pIFvF8HzKXcMIKgME9spTRQoQKMWJH
RTmEk+QxvdVvqgJ7HrDNrX8BTqoDNbEkE0EdS298rAgViODtZ1zevR7BxXpPB4uW
Sol/KJ0VbHm03VQ31nUgDvmRc2JiruPl6OX6PyH7cHi1+BnM8S7KZSH7VmEZ4/er
6Fw19r95cw/1Ukmr3oJZ4Oh14oEGphRInQDOvjAaXlXlw+L4rMlpPPaeUy+b/SFa
Gd9ZCPoOTlG2JYxtMyi2D35fJymBvNc+mYbuArx3LVfXpkiuXwsijCuc8pkMr2tM
14CTRjdd33bKYZ9AuIsTbe2et3+Ek3PWOe902f61TMvXYeneF28k8zSM4ffRvTfS
VhrQgsxnUzZXfoBSV6s9Ozd3uCeBdAyh5lBuUit7IX72F5INRVyqrBmS4Me8vh3Z
aQDXPP8mSUvzhIjIgVjyEwlWuykjTtCwRyBy3VAo1HjURsRWXcG7NvVfd/xVu6Vw
+Aa3paZMuAbpLtevs/uybYB+2BGhiLdoZrw2dpgi6hbgTp7eZVOOyDvNNoo3o+0m
tPO1Abxs4SH8pUTJToiX4WUK4ePSFxGNaRCJXaDxBq8wLK+TWzQ8WGLGv1JoaUHY
J1IA9Lg1494blkY02UkHEsDLQXO920HwJsBwj3cuCLHqwD2Oq1+8Z4mWjHjhpIpp
djDY24LrpwurCEQi5u4LgdesAkXKuzDsN3y4/wTl/T4lf8mWJsuQLtm1r+0R1sqM
B1rTfVRDzGiAgoTqfYR8XnoXfnhgU8sZ7J9BGXSBjhIsBfjEToqTLND/6sNawmLn
z9uZRTRN9sbtMR9zn+mw+Nr4o77JadUnBSzzFSxna61zT259MeXpk1OdSiJZFR9M
9JiQk3jthgGunusfW3GQ+cEZDToC1OvCREGLm3hAiC1ghueUBv6uEZd96wji8Nti
bCZedSh6oCxgYdC9chO4ES9hCuJg4/EOhPH/uBZFKAa+IwFDiIT31/w7X6RUuZIM
30eVJQlz8/N2ILaCnbc/A+mHMmZQ24C9h6sfg0Rp41uUih73IARr23saeCoibGUZ
qpVBjDEAbwTdgP6WfKrsdibaUwYgImCySZQPq7nAsiKkzMc3WkpZnV+/hQ8ivkkC
hmEgOoytPxFFmP9RQFbQsCSxdLdW/4mZs7lRzUHKuj4lEK6wm4mKeSfHg5XNQgau
aLhx8mMTTUZ5dMa/Dey7PJLqtsflzIbhMca8+OkEnxtKuwztzPnybYbUwjCsfaQs
wtfSaUpgfZgFZrjKUKS/4INaNlSLoAIzGmiWsKv1QEAFfk0mPqdjANe3FiUtzkya
OTACl8Xf2PWJ+6l7KueY/IzCPjaoJ/NXZfVgk4Px2W+q3TAnV5g3TeNoQFfv+gvb
waIidI8fxY3NKl+q20863jhrCr8XQnVoE3f1r8Iiyg7pefc4Po0vaYBngEoVWbE0
76CSBRhLWwQAH8XOJUU5PUOczr4D2tGmm+HM7/SJDjFhQ3+S3McgyMCyd46Wxo29
KOVqlT3mKtUVaf6dFvWkmYbuzazyaNO8Csf5GRx/AwSDTQNxNzjVa9FULuBmKC68
oKbBNn1g6kBohbCQvf81l/Qg+tR/WPW08+XS38lgHthbEVd9LfJko/xjORkhx4Lb
jVqQLaOULUEO1WZXLcVKhCB3oEIgyQb5MdYYDy73MZX9IBW6hnRmWdtYWpN/oGRr
2Vm2ksQFA43I38PdcIOXY3wQ1KmOvYyPi5TKvrCnzHAZ+54mGPLZNHWBfEK60Xyw
ZSK2yYZV/1rEDOCGMKctFx3e6LKwTSNkmYLwIA/sNPt+66q/LRAaBr73Tw2F7WK4
MNRlAOAY+nqu0A5CVcX+3NHrxF89OTC09GDWsbdxCWgc9UEXyWJshvhaTccHj0j4
bd/XFv8n07pgcpKZGJaDdWsC2/pZFtqJa7AscV2+7cDn1zY4T9aKfZNtBlH6OSZh
5+j3n/EyFQ/eSLwjI/LvD5zgZD0t1rqWi/UaZ8XhQPiRZtNvRXZBPbAteid35buN
9sfAqCyTa8S35S72C5G4qnDxjg8Rhp9+HYfjbylWw2i3/23lYrV81KYEMbh9/Adi
/QE/SUUreAqqUx4qauRt2WNHecqf3EIIzfuskx90wHUavsT8IEdB5BRejL/cXwVm
phdO4DfMoYGiKjcQDw17zbgRj0lUJkTwjgAJET1AYFW2MFnljuN02nCwyx4gpshF
6Gql/Bx14uFaBapusZUQhue5ESrWNnS4CyV18FPTeJas+pqOpUpJ+UvKgVsVzxZL
HMF766VJYh08Zz6KUMgVR+iLAT4Gk9Vy1Bc8Wxh+T/jzqbYHTkkNY6uCRSQbRZHp
UY4yWSC+axWKX+jBeTDVOxep6m3Kwy9V6vDNKGahJuBR72A3BnFF8cR+B9kRJSKs
s84NmO8IDR/Ol71VgR4Wud/4zk6CurCpvp6BQFdJ+21P5xKfnD2ZvOI4AmSkcl8M
46LY03jQeyvxWR0JSlZH4XSLPKQxoydJ/qTfgA5+k2m48QkDwD9TfCFuP8o5gcon
Hlx1k8weOPO0lf2fx+lqe3ppsn4bwpng6zPL1BMcQqrLUy8/n/MQ0gXf0DfJpNVF
jKjDrkz5xW7mok0kthlLs3BbrbxX8NZZtTRwSvZaq/98mBaip1pNA8Wtj7J3pa/Z
gyMQ/06WyrW0uiCfl5SniFLm1RbH/ysk6xa63YLOkCz8VRKx4r41Aejt0vf8wRgH
vIZU8ZEkQkwVdWnHr0LZx+eqiyq2kAoJci8Bz+DLuIGA3jqOy+wnQO8mCleQxuO+
pdDb2FqQZ0ygxHBLsBzONOsD/6QzMWDSMXt9NKr1HLZoTiL0QKxWmayp07LVHUre
0qpVa0ux/rl//xxjJ2ArFywUTP4UIgY7O+F8rSY3B1w6Mb9EzYuSd1NhF0fWsBOi
dhsbDRe20JvGCztURtx1JFt+8H6QgbC17SE1JxPM9C1lOWGqKcKUYxOicNT1+1ts
CVAQie4SJc8UXymYjb0T2XiwLvwaPO1fTXN0VPNizpKQ6r85A33p5EvU8ZN0ZaiC
NALeFrskpW1O4JK04gTY1rGnHrvEBP329jjG++pPd5ZbtIdIXQW/Q7z52FTUkXlW
8RCQ19G3DA8zFd2wg0xbhT5CmJE4lucfkySI1+q0JFJV0KVxniCdArj9Wkj81zQ3
2l7x2Sa8jxkUiR9Vd3NUCa1yA7XQkgfx/uyK7cplyy8OuMERU9OoG5J5cCqdx7o7
KUTaA67LMeJ0n5TzRJXlU3s94LNmvQPDVDBRwhCwzfh8NTENVpTOckx6fPeliN+K
+oNth6KGtqRS7M4PPL/J0DZehIx8344WyszBTtx25MW3le0yZqJ01KL8CmYK3e0a
6RfJsWZhVyLH5oxRuYSdVCTV9p7PjoIZwT0MoNlkdvaujnt2cZYGyTUxgR+jpt2f
nTRQr5D+Oi4HNbYgVf5ZujlLKhNxmZkhxlLzhcxeZuFmTcAY+mia+ryovcUVViHp
5OeyiY2sgrt+JsqLAYN3QPcj01/5w9p4Qxk+MwrwE8pDud16sQsM6ib9jRGUGvzl
h+ClIjBJUwc9MRpgfG69ZvBdcvqlBf27VipndlGg72V0FUAR/xyHvkolXfEvaHI4
3CNr3gqMOGoliDeRd8NnxdbZkeMWN//z0z51l2zLUytsgD8OEvzCvl6U4tJkgGOZ
NjZ+6XTdNzXvSXE+OvEykMH1YQUR0L2GrxuZVxGTFVHTLTwfXLmOPfRY1B1Gx2WK
dBNjI/RNHA7r/bZAUTrJwnKvSsbznk3Bw9LnYWqHzrVHvR+7qieJfbiQLcty6/OF
BEXnyX4TJoKpXzjwrTe7R7nwpYu6xWKENeZ+xTOyr7s9V2a6SFdPU5d0XzNGfHE3
1elFtKX5/3PrVI0I28tVN2KUfrHnK0UrV/MT247jkJ8aWVqZNHKvB76csBt2MdXG
h0lC1xI0e8eZBEsOYmZlMxV8+UHXNKQr38cPUg+l6HonZq2XqzgGePZWiCSJhZl8
OzTGpl11VyJFWubqHSUs4pbGu9zaPHFb2ntSQF9FxEJH/0GyRX54NB6Nr/l+M/qm
iyK37zP4z80AsPEKQ05dc7a0vQ2h735m7rVkKGhPWLu1WpG3mLHsXFjUUZLs6PkD
HJOzvN7WZq05REpnBT4hz37tFKsVooIT677KmwtXnpQxsO1L5DmGNDD1YO3JX8kG
q0vi762py8rRWLVy3pGTUWbvM9MloL60LVX+K5sPpopFg9d7FB7MAhhx6X2Kdbsw
/egpXx/MmQYBq+PEfZZK+6C+hK5a63k0j7IisecIP0RourrzDSnNiLvY6UK5ZfBJ
KS9HjyBq4Hm7Db3xSYeXd7s9BrxbW7qNNdBqUtVToQOz12vE3LkaumQcuWXy+fOX
nVSNcTZQtAkg+LOJlFPhXhnTteVMNOF4+4xtPNpnVSY8aVJWOJnVRFnsylF2Bpbd
NSHaU1Ut22euLGD6NHkjLzevvJoa1zNCvxgTfr0BPG4iH1jrl5ThlWT/uXnJpOfM
Kn2xAPniwmycYXGXfw7ULW5OPsPz/Neyq4sYBrUaTdQRDv11/H72v311Oaxyz7qe
4IzotMUTXCPbS9wXhhcxMaU0ydpgmzaWa5/wZvERl/oQqOaDJ+FV0B793TF2P9dZ
o1IvqNGJMjuVaynYOcC0EP90e3rau4324VSkDZ68rNm1BHGhXmFPmkEJi/FSDT00
6p4cDaks/ep5aQ9pZTlGZK7DRVmEpM4XDec4Om/CqdiMVwUCx1bvjI/qwdIOcjWO
vy5b6Tefy7Bpx+BAdiyvDpYldDrhou9f3Ip3E3spvkbBJNA+5Ra3kb38qOFnIhBS
921bY12+ofvGV10sR9QdJ6y1ph02/Emyzh83m9e9E8KthsdL9DzVvh4+p1OQVRUI
h5i1X+JKemniGUZ6CDqaSaVe85Jo3JqT+GEIOBNnkb+YiwXm1CWD8FMMATK+ME7c
fpA5xkPwPvXP4ydAURoweradthQ7cTps7N9X4jPILas0eBdOguRloXtuOJSvRWBP
efGhyCTdGyiedU/vnTT9gr+9LFgcdPwmT08BGKFH70KB8il9cf6x2PilDOQwQyF7
rO1Yki5uhFtP9q+x7P7hn/TJpqMS8FDc0miDkKvJ8YpPEOoL8rttF0oGgrf3Q4lW
SKQQ1khlQDLxUJuRRXhTv7W2uBnOSHWcKTGXaaRriv4uQ8vkVGpe3CUp5/1dERkE
E5wBERdPGnQMC1OepelEKdzHGhi91AX/ClYM/iYUcCwWHSRxLG/RvAoYfwyuOS/v
JbQJUKb3fZpkSd6tUmxFty1zqAB2JkIdjURACAZx5/bwDUpaK2xW6pbKVOdP8X5P
CtlkMd+9g9RgY9STeNedQjaF0D4b609qi/eXWmV40s4BsAnkKg3FgumB7XBs6N5k
gnmE3tqX4pBUylj2r0MEBckmEo19AS0B/L2hwmTQ7EfhjjmL6wfHuA4wqcAYsje2
pncMJu67zp3dwGW3GN1b5as03VBhOiWV4f8rqhosEOslpoTK2CO4H2kkRAYXUgbB
oGWfU/w5/FzcVldNcFFRtmRk/xDFaExyqRH2NspSVqlcRYq1N3BVqN437h2THzaW
XEf6aI2jBBbBozyZOoku++tCWVqwTC91VU0PvL7otwLfbJEX9SAQSAU8JFRyxLxA
RxMxGGTyBc/rnR24JY4zRLcRol5W/LR+CvqmluPlgA8909Phf7TFSDXsXccp0e0m
tuobG140yfSj2eCTvhJP7Rfuno+n7q/TeiznlEgztX1GjJNhkNSKUCmFPAsi+HoO
4Xsl+Wx3ZqvYsPFRPSpLoWBnvkHl1UAuIb/hVDzOtPK4dITYe7XrLi6Av/uW/Zij
BJFdOrr5b/DEAmShFgLss5yw8GVpPPz44ejlmhgcLEY0sSUdSCoStGFd+doB4q+Z
u7OdfrEcWHCCo+1GQOlgy4WHvltBeg3JA0B5nzXJ11UCQvFqNQGfQRMWajNcMBy0
YzG+I1RNuYRXLZf+sRv57H99nltM0kqLOyiKHaf6pQPEenr5RwRFdF68qNQ2ZQB0
5e9wnesyiZIS6iXqyFIYCWTwditcbDVapG3L3Ukp3uPWLWstVIvTlAWKmIFmKo7U
JouY+ZR2Vzf8Ske0RSb3ZX+9EvFgEZZvv7KubW7ycfMc5sU1uFvSGbLip8SlYiuM
RA0wrGxzyoU8LPF9wEGCPwvba3MoGPKMAiGap0/3EXmAjzbfLBAKurNwRDZw50gQ
PfbVagaHxKmgJ6F4i9AZBeV+4KG31KxLxpObrbDMXp7Atgc6i9bUQX8E+oJH5b/t
l6r8tRV6AcroaQIMJyNoUrUHB2KF7dZVSce1BOsiwFf8i5p/5/4mQMGSjYvrldoj
5GrC/5M7kf20pss3dtKW5N7IgwI7L+lqbA8NPtAbwoZNO46tdncjakpAU2blgAcN
ySxhNk3a7YIyQz6BSuSlid+u2pRPOY/soeyaSLSMwQMgpVyFxyXavoFX/esBdQM0
0KqnGm+DVjB9GdO560ewdiQDTceLRb1qx1yueGpHauzm0m96NBjDzAci81qJNnvY
O4kkl3AzV+CFeP8/+PiDTv7H6vf8SH2Zt1EEb0ul9WLoAGiddV7OoYK56hVe2hzk
Pc6jw+2CpiGgpvgYQ012jQn6EnSySYCFBjbfOTbUVHjYxpU9xcJ3R7CI520DXIcc
0Yz+psbic1KFvMWxqTNbPR/becCIbnluiJhkB7tBD6c3kvIP5H/QveAZO+0UK70w
6PKy70fFvZaTtVyTZGKZXQBO3VxEX5LwZmwE1yuAedaziXyFK3IU+HUReYu871zg
D2iJYoTCnlE1uQ5JptjApD37IE0SqcFzAZgEdQBAj9aKWrJRoPronx0zx/AIwcSg
BB7SKz100uv0UnBvW+M0hAwXfjrEU98PmN1boKpJd4cmSQ3d8ve4+nwWJXGkFt7w
Fmz1qy0kXA1AQf79N4VbS+wXuLZlYmKnHfEkYFDUDT3ov9okOXxanxTiR3rnIBQK
2Qi0H5a0EiB6fGtc/JUi/ixEvBTD1oTXOB2cU2ud1FA8l9veusocXZ42KRdMDnTK
OVkVLZVV163I8zHK6f7yx1ewgqJGJ0XHIjieXtimFjclec3x61GFgxY+c6VHrWzi
nalFVwQ0vBjAwveRcnndDrpm9J46y5p2wa59iuPt5YeWwAUdA7q45z7W5AMhjhEN
8BpVgtR+ZmtvRXTrSTx/ndMWjtBK8o/lhVjwzgbYQU9dOqHzxc0TKeYQ7xC/uBlR
IuiaJTDxNvKVjsDdS6+4HeFXFAPPDlJvwxSNLyfNCV351OLFIwJdfpl9OB5rimQx
9BNZShldxd/ucLI04f5YZui2lczIns6rctRO5vD6MsHvsYhva+9HZhHHxeriBcSO
2OircZ6rS0FcOC7n+8qz6VMA7XedF7VWoBuJLKE3GIw4vA+QGr6heiVRgKlU/Fpc
ad5oDRNCMcIPDmw88WXwzfiOnowZMQJwOCtFuIP7bL8qQ2X02hMZO5NUuZ+pwyIl
2vkjyKA5LLcx/ngYxaijGndCuc7v97kSrrszoQHqFo5kGqMukdq0kFD8QyLNmgF+
LJ0NPVsVHM9iljNWr/ELxBdt/QwrJTngqhebp+KexRpY7OOaAjxuM/MIFOW3YQLf
gzpoNpsYmMd1bDx2yv2LyJh1iSY+Y+A6EJCTwoHGJYV/UHqSU2HF+dKis8E/N2l2
ZVTENHn5MT1UqDNo2RJf2c9A640k37Gu2suG6LAOupnFmS2yfxy9zdikno8UB/d4
Z8AQ9AzhHFF5UMss+fnTie6KtnJnF5XTefNbmXX0H6rh8VA9wtqS67Ya1Cjln5bw
/cZXoG9c6gnWM53ps0nIEqpgmgAW2slODEU1be6aJ3btUc7yRY6z74U8V7D6cB/5
of1aImCKVKjXQLRjNJZQZfJ5TLZyIjzpmSiBm12AxOiu5pS0UufTotVZRBFRAdQe
LrxgXC1WLisROsDRqsm04dgAZ7qnedmMlUukimnYS+MFBO7Fyv15HBNWdcVvfaR6
kg/8Qi3tGz2fCGA3LRe8H6D+5no12zAtlsTudZIoveMeazqkvht1PgS8RWZZidb+
HwIuFtFeazc8U55/2AIBl3xsw1eQQ+2uIWZ/uZtY2GSvr/1Rm9Q7gprtf2cl77yK
WBiDwT4Aa0qT2zkvIAMLq6/ObMU1SyXg8L3zRUBUoWlmCnOriPK8p56saw+o/PCt
bHtW6XUgJU08qWm1QSFNybIuUo0cDKWlWDWyGNBxC5SNWy7q+UbbpT4N3J1Av5RD
Xy7usLCEAoPr3JzqJQNIOyDw+DiwEnoXR4ccjbYhVpYnBMds71dJvFj1BGIXbvkc
yHaFlJXHSpPBkr23o0uIkHimIwqO8RhZDYi97GKF/WxuuPkbNaKCXeDhtTh4CtjC
NkSA0Q7a3fzzv7d67GOMAtpDEd8xrn3dwdzXrCgkepMZJbSmyqwncRtY/gB7uuIE
7xcd1+hXNMavo+gL8s/S59qTg6tBgbUFTEb50XHbuHuzoxV8mKXhfqRxHggNFncL
3Byd+AYj9EdpVJ/E4BdxzD1VV/EsvEUktZWeGJKqAewHnfY2uO4aADG8fMnV6081
1jajzRXCAuuQMxifpxJxfj/RIjRJMYZoZxtks80JnLat5ww2lCxd8zsFI7zR8Yx8
iylODEgJM+wI7VEM9h2xUjp5i8EGnj0mZGegx7gpPCcvFhWwSTbNAm1CTEJLBZSG
KLCtVws6L/g5rJqud3kkXsjzDF+suTXTGiV1FtcKUjZUCEOIAAfZTvyuHSefkzFw
kCG38w/61xcZO98mT1QQe1Z57S5Stk86tZXp14gXUklLtEoA7j/KugzvqxdGgVDU
KDk+/rdYVpdQM8sKIQemyuNrgQa8tCxm1l4SkKD6uyrxYmrYQ9H7TBsbh1fol2Uz
ecQiCNUZbZ5pTFz4jyXFS5C5N1QGk9UFgKSB9KOG9sp3Ol1RjSI3l7AGaUdSOB1F
+FQF1eQXwGi+P74xwRDKO4Rty9vuv/A+nd3Sa/cZluy1RJD5EqYeqdp3z6xgRLvH
ccIuzLTNFBiqks8k6WXwNzDpx8yA68rhoZsDwHb0jtUqHJokvPuXVTAN8XiogSgD
yCBfnpfHc3vShvawwIOMpiatUNGrCa5DZ4mSDmEA6uqkM++BraWef3Ca0FcVI7pG
mg1iRG0LEGGyHbW2qrx4gPsdRZ2u4NsPWaV/tUgvMZA9RZhPUH+Bh3cCqH1IvGc9
hKTadvZDpPSf7GwI70Oc0RXv4wibVbcITuLxXa2GPMwhbv+Rh8fbAnEniMBN4213
04MZLzSxmnKfiOONstvbmjZuuTOjZN8IfA26S8I6CFsz1wWaXOixaEA5/XM2Vva1
HgteaR48RxYLEFMgn1LJS72dlCb6wUDqgEpzC0rxG6u6vl/jRo5wPqL2JFYLskTh
sRUINnbd/rRkAijHmK6LvprhdZQ+o9m9Jgg8kBkd4dJyMOVNrR1kimK8KBMm3PAB
Z2OzgNDOFMGJVBYw6zsSwK35Tahy/B3uHwUZNWm0zfFwmU0gVOQDEz9xnW1vLRo5
s/lt3cli3brPfqVcqTWNsVFlbdmE4jxXikPQ/U+APuFN20bXHC6xcCgcwmn1dPMY
fDoKLFnvlsueaQI0+kxNdIxaRQMwMqVunFwVuCAF/LD9t5CexvnzE1DMWsIJ8Im6
WcFTLBZYhaZ0BsGghHluemuhHoNTYd25HVFTcBI55PE2+81WY5zP3A7PSAJujo8F
IpbzOmUL0Lan/d9vwY5Ly43xs0H0k/JLI+1VMo8Hr1IM29xqaKktf5Ym06m4TPtr
g5p/cGB23Ute0INkAgZy+0DrO+MzyHXAltY4H2zYAZgjD6PygH15ueBwmr6PKlSy
ChLwvhvZzxr38opDsM1eFs6wEDijE+ZZHUu1d3GZUZ5rQ6TIa+RFWJs0dfqxSreW
VVMuh3OcLjGCWdLdo3Q6NozKsxFiRlR/mWDNbPoAx5Epj/BSR7dHBFY3fNACenWJ
mgJxWMvmelF/00YV/Hvka4LNsYTFZhOPoz9V+PERIjSk3tJ+f1+DYSw+RqVtELuk
Lk7NaOnoME5ReFmt8TvrIMJXJiV9a7vK7iuOdVimz6jTqDkXwZ5B7hCldJmJ6+hU
XsmrDRtJ9X9jmpHK4SWZuY712SSAhKl3UJNdTCfSqJ6VLTBRhZJjbNAfru/m5+fM
sp3Dtxbq7fhTB8oNfumzH3xgDYOeuffMu3UsCu+AavbnojbvSAYvle6tuej8F/sj
hezjBFzMBBkxZpmi62ajq5Rxlffx8OyQZ1/74qJs25DXh3tyZCzdS0Kp1xoWrwZa
6IEfD62IS13w7ii/MImO/xXqX7VxBdhpTwAZ+CWMzlreTwKZHMXcA5xDWQ7CU3Sx
FEVWM5JLWgmC9FQsAahWBrqluHbtUQhXaSzoj1JdS+KmZjzT9Mcl4NGQALUQKP5a
/cSXXs89P88M8kOPXuUKd7eWT3ox78zxckdYIPPYN5uZ+Z1EI6fDr6dCOoaMSXZT
WZVaZ6UKtoFovNtJJk6/eXhGwugVCPnYQsi/+QpJYnBWFtcJcjxy7FWJT+h6byaV
v++gIklA3iI//f7FLWNbP6XajFIGrA9wRDeOGpAp1LFRzHQHSAXIOKYzofzKiypD
F/GFEdydHApk9ZKQi+i6fEz6kJVfqu/QJnN0PcAq11KmVjk9qVdfTXFeT3LKDiWj
+yCdwfjq4CnccL8GVaGbbMflnj3ml0IWMVssIG+90xH5vi27YHZ99gCXz0CFbqv6
ZfR4ov0NxxawXKui4bxU8w11KOQvg2ZFx/nqHq0qXzXfqjtWy9qmTwAfbnI5XREg
NDPhZH+D8cZfvwtasFVyL6vcXWEBW1zsDTclvpJR0d9+mb+mA62iaVUAI+e5QVaY
M1HHbB6+3xNhIV/GTMPQfZ3NEI3JizgwZzhcByIh3E+27kn0rfwZISCKic1YCpUv
VoR+O174Fpt8PEVsltV7VQb7HxCVLjwZ8kHP2MKlSCspkLvqDuc89OBqNvZFP7oV
UbgazOv5UXtAJr7eDD5GJI1OoJ19Jzajer84pIIFrAht3F8661n3HpaCSaIFKBaq
WAiOQrrElqBBd+0mC2UYb8FkI8awI0MtrLYQS0g/tLtbvlO49CrRv4sJCrIENz/6
lG0KTW8QdIX+P5NT5bfOvei3wIREc7XERF8xhbdyY8J9rXr3zQUytq+h1rXFGKtM
wQDeKQ4fx0z8b8CA9/CIbiaB/ANyPGI9KmmIR+bkSg7d3v3+fUNPDnHsQzys8oXe
Gf5wNRedRuNgMSu4VYZGUDD2ApQ7XhUtDX0qX6ML8zM2dgdgk+yf9y627V/ipNgG
17KVuBkI8cLo1y4M0rEo1KPQV4h+ub8HybPefcQ7gts+69nWyGXAKu1QkVkzapg6
UC0OwcwUFntF2vLYJO4gZ5XMUauH7NEIHadRp3iKs16rUecegLPLgfeyFj8I07zv
CewRDFSIyrQTqLNOpEZXSAPJAMihzo+I9REVfWPWVRGugSgVadcLKY0WcX/Mi7yC
Szv3GfIRfGk4uywgCKvzc3twh2wOJCS9oJ5toQbVJfT64iip35Gnf1yE9rqsaE92
ftdZoaBDREPpnzOSIUOqoPQYm0TUFa7mIMVRyafw/MXgkeGKSI6rh/M6DTgDC3A5
QMpKGQc00xKHgfN6nFlyhKbPjUgr7bhZ2gVWI8S4N8+9r3LLl3K1IDf+OPbEu7RO
HF1lk3Mc4nEwO7imF9sagn54bgK2aXdhhVBqQ3dVbr3OPq+FUiurFjdKZpLNr7hI
EG4+ITsPJLBRX3RwXWcfYL9oQU1OkYUBld79jFnvVtlMHQW2PTT/eY/5I5AGiivF
uR5zZr2WtC6aF/d+xaKUxLzQslxT4fvJiI4MBQB8C1qnM2AcqZs234GmXpyXjv7F
B+guYGQLh5jiin4mZnIVb4BEbCsOjJv+eMfDDXeb98Nqlu/Pfvimrt56BBOljClt
s0t71XaIkoxoLbLXws0LPjl8RuO+nZ81+ByzldyO4yEVK0bxX82meDXIGy+Tk7Nf
D7A2vehvb5GQVTgbqHSJpFkG1iugHLgVDtUekCNADDiMDr0bVCW6DIzcAAL4AzIe
qD3FFO/hFtZ8V522AfsNjjm0HmPgtkBIWlMLPagcuG/zbk6odEiHxCVj/+IETjpT
toBB2PgJsedcsAmlAZNfQxzEpBqCDNS0EuqvYUQfsFfUXXf/WcCbL/eBpCWMXBlx
YdCWMWTZz/sZopgcU9k9eovKn0y/x1IFp/FOndV1usRWPU0pyQewEMYu1lsqKwVm
ejdyi2+HAaqSGTflUFcEzD66j946DMZd1wcrrWthTgjnHN4RbwSoiLQfzse6bw7w
uBT14GskgDLWmLir9UIJFeG2s54s/OXNEyZRw6g5A/NhQxLsv8Q5FfvPhgMyLDx/
jsA72dHr4GeD0534nxW9oFyZU6acKMr/izyhU2z4KbQW8u8CbTfW6nhWXUIe32Er
tWo9Ekkzkk6Y5eEL13T5qcD+jEBcvIl/b71yG8PvRuumZNDERk3GmuPTid3gDq15
ROBkwVkiZbnSCVnJEb58enY3C/zo00TRvlavJ4LwEKNsT4jZUqUZy5JXjt4Ffw9K
EsU+g28qts/fVaEn+RCIFRQDH+h5sgXDY5C0suw/j0fxawVBLCVvb+xwBXeUj0h0
X4SCARS7GqEJrG9sWz/+SluJLM1ApWwqAsdedqHaBHzI1UcP4I9k5w1TP1rX+h+Q
3OOtBxZxu6wb1bGCn2EouKjl2q3tdyQrLJXiObAvDGRqq1JUr9zyl6MaN9QtcAT5
4fOl8qOctR0/6lUtIHcNpUxzp+Y7gF+GmzkEj+30T7jftybg3c6ociFBS6jSG2Al
Eyrd2IKZxlgUdyEvgCKeX6Gg7T6qo2AKrwPH+o3/oePGMnRpRzOPKqqPM1hoOHr6
IEcE7F9Ah4GuIgvEYBjIy9PH0uW9H04NUn4HHRGZJ2SmVeE53o4cfWa3DOZK9+8n
2u36T7LfOKwqgnFm9VT3caay7c1GtgYcM9BUI99YVjmJ2aVI7Bs5WjS/Kt5BSj0S
Ft3yiADOL1d4HRJ7DkmffD2NmGCHxZh6yG0k2lG8AeogP2JSmSjwrvVIKlmlxGgF
sALgIjT3V8G2yXFyMIlki4Wfr1NLT60knTsC/M6Sk1mV/LFGuOTlnOw+dSMBrR6b
gcPyGK2IUKIzFFQKlkOTIl4Jsy7ItleQIYMGDTkeF+q2lrAdZ4Ip5XlslFdmtpVC
7ZHgLSRmMsQFsXEpUfNvl1tnsB2Dv3MCf5bJWilMWN4VqUs9G8kHGxb4mgdiMNdl
qtQ9VoqHG5F1FwFhuCPuYigi0IC8W2HwGqf2vfDwYgu5Ll8BBACFGWBX3+BlxR5Q
D6KTMriZXNjVBcHu4mzy9OmZF3k4linHu0eKMwD7m33fCpyT+C/8Dr9F/1qavstL
mcvED7LboptttVVIi7kA1TACCGMnRxm2FzxhEt25R1BUDrbiYohMto8ETkQhbjjo
+ZMgOvW1nAQ2jfxiaZUF6AT148FetVvmeOz9QgZCNSEVzEiDksu8pFGnhSkOo7Ev
WkotjYle7tOec83bixtHqEH70+M6V9iLfU4B+UaIvpOpu1Fuaxk17MD44onGrFHN
38WxtesiZiObCmVNQ5+g5llwRsIj90+fYciqYbbQyfZXD49Xn7r/G+wjpXjUyF6s
lRfGUW+IUDYZfeVnHhaw3Y+30BD35+dZQeASQY1u+Es2+rrtn5nCDT4GsbG0loxj
72b1j1UWq+El3wFuZ2T0I167anJbhvPJBUPxexhLSQCLCpMYW1nUhDIckqXkYZ45
/oIBL7+ga72LA5ZT179uX4WEeQ2oPxPimINnX8fj0rv1ERpy86NbfPbqkG/FtlPV
pbl9anOh3ibFwHln5HWtTpk4VAEzNF9xIxLVlpYhvb1PiOI2JC9HgJRH7As3HylM
JUWq+kgpR6Txn1w3s4ocrytyr/EVlQ4hlp6bdTPvL88aBjU3ciacRWsnPCumxW4Y
iwObLggTArW78SAqOFIsMOcBuufFHvIMGjB6fw26iaNEQI3OtUsU/jz/KFOyR+D0
d0QitiYeYCo9fbFTG8Z4LeBHfq23wLuT6sw29ucMDyn+7g7XOatuc4MZHkJNz+da
BQ9CfS/8xRDI4BNFXueQgYIVstdHi1aUNMryXQfW6b2XZb8Gds9eEQqgNdikCqrU
t/IXlFGx03LGGA0R5B/0iuXdumsm7yPpWmhqQXxs05oAXblR7G8xlmuzI52TDnq5
3kwxaQtdBeHA7stCk6OKMtHmQa1oQ62Z0A50N4oyKaO/ZCw5czzyrYyfX/4zntLN
/EvKj8s3hhINIMEFVi+j4l5LqrOvba2u74J1Pf6V8jMbLJYYvuj1jozAf7WFITzP
5AfEzMs9JJ7+kAHqn3hMgKcnWjYcZpBiKw0xKTGFsQficRSGz0fMrynFH9cssuVz
MLkgfvKOZJQBdQjMCRCB2WghUwCIu+ux/yBlPu10uiVuwVOj9BfnCnbL04Oi0tln
ej8LoyKwM8f2Jdp0JtHEAU69OdBevsJkVgHCuEcew0NGnz2voTS+4i8bRzqzhIl9
fwlWZtv7jHC/k/Xqf2wXug+JkGdEGuwIsy6E6UN0yx26m9zb54GOcBchWRchOFU3
PY8XJktSFp8S9PK/XQKVKsQ7+v0pwIFYBHIirhlPF1d+uqAQq/4PemPFe0GREFdG
/hMINm1+jGrO+5WpJD0wrqIH1FqzuQEe9F/sV7wR3ms3iaO74znwBdJEpHayAAdy
f3QswFUQr0zBiAiJUVgv3z5oUkUjqiVG3XBqKqUfBn9Nrb1uXfvJSlOg9HiShZ7E
v/r7duWQ5pIrs1aQ3lxcHHcx3Hrlz4W6M7ESDwxtDyg0Or4qgNsATLIEDbQtKPsm
O65nVnRsx/Ya83v7Cvyvzqs8UtqnAsz0dHdBA3tGx4LwoPwnQbOCPj7ONhkEFLza
M9nw1ls9OBaxHk6+t9OuLMd6HPLHKErDYYt+qh0JlrtXw9DPcgf/51JuKfYhkB+4
DDE8TDbua4+9/lt3TZN1ebkbDXg2LeXQtM0MXXhmLPF2lQwK/wmvlVN+D0sJnAwc
1MfJtdVC0qDZmXpbJXa0HKrTK0XASTNMATeIl2IcnkHgDhFatNgqBdFL38UvhoDQ
YkycyvabTtkZNzDedRKvweYDxlmt1tLT+05vMYD1wkL0Zys0D9SdTu7TBcufGd/5
/ATJPVurb+4nna0aW3EKENkq1p/yBzY12tFk9d23hRiQf6+OOyhaNRVKZoQ6Z3hi
tDLTB+dkA1QgaqXfvx00kDEYk770uZ5/KTTxI3oE1Gx1sX17XZktt4PdbzsYk9Pz
E9H8AETVyRWfaokjBGiRxJSNoIvFczQnC8T49asqsLy6NrI+fBDIJSiVDS5fIIOe
JJcv7oyTTPheofgdyhzlaL8eqoBuGuHhEG7r/uQdt/LT8zVeUY5pGnw6OO4i3Dfa
p56uutB4ViCIfTGIlh3DiXEs1Ay8LnBhQS3T1s6AB8hBgUJ9L729O27pfs8CQBN5
/uyaEpjGi5cO6vH+ieY8TewiN0RbyHnQzhyvZZ1YSA3Fz4Sjz/nkbMrEzYj/Sfrn
9E/6CymMO4NIhNR3vjZ4VGzt5DUDcWYBOpQLVaPC+ZdHFexeyTWHLg1HuU7qvzA9
c7iSoHXCPwF/1E1JZklgMFlk8uaSIDIExyTRXOftg+D3kbNxhl5dClqKcr7CqzpL
ZvogcajxqGMswvdfry9GM8DiUbm0Wi1C+5W7Mig5N3GEz7ua8ULwiT0M90Acap3W
2acAyrS4JRiVK5ZO7E+sqGk8nhUGKyZ1+8pZn/LZEDp8aLfkdy5vst2gscC2l16a
qfWw6NForUndtzHYdi5h6QaLjJMttE+dR6AxeNxNoNHqtIdM8rNKD4YPyM43HiK0
kC03xtADNJe4G1kKDCf6pBVWjylHjC7ZqvzGTN1pP9CUm9Dvk07W5HTCBSMUljy+
wSHkSkOiWLCj9d+VWU2KzRFTYPRKhqcGqGb4IFhaqMJ8SCE130PJIjj+PhA+U7Wz
dvDGkZGSjMmdwynPiub6ZcRgwoQbVGIB9nCZtzoLofU81kxBi6bK/1AxuKtnx+Gw
XWNbv3LYYFM16skCKswo0wWnLGaiRzfNvou/EuL4bH9o/ruxSO2CLT8oqzUmNov9
z57Tll9bU/7AydMLKG26L0vXmKgHtmZS65F+r8foATmuiJMP8wvI8nURqnjhar6k
rO9AaxO8HOMgmePV3bgYXiPRubZuy6gJ5d/N/JW6WRa6Md0KAwP7KLwr6Jt0xccn
2G4n0JoevDT5ACQVL/GxQMhUx+TvsRxXtW0RIc03eofg1aBNdQ52vpNQKQ7Dhkje
CCiVtdfB/1Zz23zJu781wT2IZWF9YrRnujs18z44WD0caTvJCsVM34+HtYRJeFI9
tCQcyHPreCuTN5q7yTZcMK8Vnx53pgS4uIPh+2lLS8howo/DnxHMLFG6+pWinPDW
/jPwNZm6AjOREW/aNTs1TX0eEn2/xq7cNPf3SgYlpA3VpVqe+m4DM/cq2JPGlMF4
NDh8WHU4joC0U2GVfXsr2GAW8KY/crmV4ospHSpB0VoY1R5cAv+nS4BPiVtIA/Bn
o+TAnx7Sc+SlUcKts88DARI0em+vJwD/0jrNHGJf1W+FIJCzI6XdTf/mZHzvlv1Z
sJX6VHJgeKTtnW/sRmbHKK08gl0CCjKZvniiNgxAMpCin+cbT0uZkxVVG2tlSwMu
spO4xRRcdPDfzyFtvx8xp6YE51TtKRcPRHgawpFab+tAxoE3jB3k/1HRCpP3gm9h
ooraP5F/R74X+t8B+AqhrHv6a2TpRm0BPc193KAaGb/tSnwvd16HaFDRpcJUXhd+
HFIEIz6TEX7FexqrPiFt+h/o83a2F1IvzWbWTQUUKgSm7ibDeQF5C87jHrkM6/+6
8066ZbEb9HE/EHZ6tnN7KkYOEdQ3SIn9Nr0Xg+RILGH9gNTDYJF1o9ar6ibnA2oh
DIehe7zkC06n2ptrpzZKKmK8SwOyfyOR1DkqZ+wJhKpQfBs00rexfDaliJZtvYh6
90EQdi4h550WHt53WswR0xeaE5Ot2LtOpfojLOu+y9ZKmU7VyCOMPGRyhUX5KwwO
nvplHhMg0DmDv+zcdWEJ0oxS8BZzQiLWGsFsEYV7wSH9gWU4qjc3mhEkFYMzbpzS
isJ4rqk5qEWDOjxmmQPA/Nw4bDMQmDWZg//enpycUUcy49XTZYR8Eafc3Dmrr/EY
qrXci6hPYLN3D+2DfUUbbvYr2GoO7+cxhcE1wwH+ENMfVB4MPwzm1vWz3JlJmmwC
RVKf5+ShYg9IfoFZVELDYwUQdi1Hc3797jC3z0kQct+4XN/Qm0fX8HZLHV+7CCik
Q7CVws9Yk8lXFzZy26sZjs3EzlCkroQszavwfqSagQdI90FLUVMXIaPwvRZ6zmkV
o+ws+1S9A+RapY5uOVcJUfqdg2Wsxpl5GfpZUrkbgQuKdYWNvQNjmRHhMsT4RE8e
AYqTNLqML+AJWwvWi9uZ+apgZglNlCMVmEpZsy3XKc6POQo0oxiYN9IaUxQZ7H2o
6baQQluEqevEivF3SU94NZxqrMs8qr+8mIUQUgN7CiEkTYNisiG5ONgHVUCTBHzD
ktk8oFqAhhK3AqubmIRxPdSLx0atPH2QL0WVgh3FhFjsCIwJuQckK6OHV7KYziXQ
OPnXGidWkmC+gwtgHkJBNW9I/nObMIAGwqFnME7SuQfpLNfRyebUNZOOjL4/ejUM
TV40yf2/oqJ+NADS6f2NHW/4wJl/RdRrcVq8S8GE5h4T8BeKFHTAYkZ0pSz7ACBo
hHUR4eKCdfPsjcWiPu6YNfP7V+Y4jKE5x02ouO0rYwYPLvUJMHkjY1YZL7e3TvR5
AC6kvytwqBAJg7eUz/JoanVdPQEwFNRSoNV4A3sobIUFM7VrLG9FgWP6BgQ+B0rf
30nnlf94/TPRdaaJfn+de3gVthhkBkd8T/V4FF3C+nYjxbNo7JfVXzuJ87G5bl15
7ogZzfwpJrqp7rRkJpU4o4PeFqPNGgPGOM2BNddB5ROIBtRfaP+1LaFtD8wS+1H7
lTO1Jm1itE2L6jhJE8xi+r/nMoMUUDQtEjxJnqSRJZAy0jTpnzPEN1K0pIUAUTTx
ogv/1LUqTZ0L/czCS5y6a9G+dtWU/OF4bX0j9SiYcmAKSkV5JEJzLy6Nfc3UlC4m
wjiJjbZBSA5ApSxNN5rcUhl3UDIaWQmLQjpua5VDjfZGgiRlDcWdDV1qMN56LLhj
gh2OL805MXz8/ek+M1xY9WdhlJBOwewroypyCUiQVcHnbuFuVWkW09St8mMLkbAl
bZwkLU4sroHcKRvZHGCu/b6h1g7S4mlGb8+hoy5tWtGzqVg1cVj+HJmsbv3gNJtk
XeZh+gQDyomNvGpYBmeLnfT2srHhBwyRKAyb4WaSIN/Yvu58GNxEEkr1BenIQ5+w
uv5G6p2xKmzkUI4Eu718WR32FlyfERjbNS3plmTxhUqKCfCFSNJ6uLuE3YdbB+iO
cISR2VmQh3U5WwlL2gdWwxPgvU/zh+BgrpuxhzKqM/0l1q39m4kBoDTY6p7IjVXt
lC/8Z0vwe2URgaQXjTMtpfMQFn+72m66Pf8Im/gHmt0B91K1ONoEmtXtqfvFeJDg
couimP1IoNIj1ru0AQU67bJSEzMUtzVAw3YZpHXMKLDpsgUw9206jqUOs5iSovqH
sMhZbNE0A6P5yKXX3stqm74aB/QMgOjALymPAv9Sp+u8uZuy9YyPKz4r7JBG6pTm
GtX8G1/DsAA0ycOUCmuW4PSRdXdDb2dVjpuBrowIOdrecyQ5V/SKYxOG8M5KOU0x
0fL69FRomOOyjVAzmudjbYZclLr+5VTgWAaAgyj7Rf9qP0NWNszotGFKyZ4aT5f6
8gKCIsBAo59cHW7B8rSg4WtFDHY+GqzC2AZNopr2s5rOP1yNfD/ioV8+CnOfWIGA
184/f65TRTdOR0poFY/4Qk4dHh6lxlai0GCRzUqBuYTLeERs86eZ//eJyw6Kb/Wd
OYEXMyVGtMBsEHqxJFSGwdp8Gg58VhhtUpb0kNTl1up0yn+eB8vUCpi2RdS3zuSo
ulIbCdshZwpXBdhtsIq+/1XLnzMua8lHGUpZ0U2eR4ekfvWiVHhv9BcBpqXtNLHP
xJ31OYH/Gn88ljQ4LIce0U5jQ119GT/yIipAxOfV9DCCtJpvkLywJJBfffBAG0j9
mjK59WVujlIYxBTvhgRAMyJ5Bh+PhV2L5X9eQEiH3ozXR9PODH8cAFq+wz5H3LwF
u2+1ToFppvDZYzPn110Ck3xIFrM68aFvZrQDHdp7PF1E7twF1v4RscIHFjXgCX7T
ZDHlUpqveSkq7sgCLUXymH3A6nSuuxmxnJAoXKCaPRQFV7yZtWDDDwX5hR+QsBzr
TqevSj7a0WUAqa4xdVapv8GIRStBdrdx/lWCk8aNEt9ht/PHLnb7JIPeZQD9SWee
szvNVl9PC8XyLo+u2JZ2YUYMhnI0z++1F4KGFqZbxO5xDd+HEflF4ecrs22aq8J5
MTtbOVkPoRiMZO7lFdiLt7Qzfn8SpCwj0jtV2UY+k9brgatceVGpAMNqz1GJCNhl
EKizis233dA+d8TSaPiq22Fhlf+34UXASjg83kAf2hPuAu51u3lDEpvfvV9LFwHL
0Iy3y3eg3kExyYAkukfn/ZuLWlahH6kslOzhUqYUAFgbaYU0opsT6Eg6brewdOB1
NBRxCrpsLxAt1vIuYlWZVc5O+wkYR6txKdHA/yUPCCAcv3aqBkNLJ7TewSyOsUPi
YuIKn94Tp9I1pKnZnw9YpnETwS8gm+j5yBNRPfbatHxR4MO0BXE8s79vfQZs+t57
BDo54lghpXXjgNU6pVTiJRramMsYKGOzPkNP/6owu1LyKHH+5h9TJJJv/Ych9sZz
sPoZHdmiD7OprfsncmsgqhtjistFj36efOaeb2WS/oUfyZgoQlNvC82KwXCbwpfu
73X8jMic/9sbg0fsDAdQg1DPxtYCXcmPfxtla8XcgshW90X4+Oo/4rUfIbjNOoAr
SRmaimlEyhp22DIEOh7J1yF7KNkAJr/KWcuvuxUUb8YuF1/NoLI/0ZagbRSPU4Xo
tzwOg/arudEYM6ohy8x74PDTW5PBZXM3sY0gGsNXWupPlmULCIr0kBnzf0YCdCGA
Rodg6M4BjS8q6kygiMZ6NQIJAGFAsQkEXGc2FnW4zzwmzMwEkFcFfhKovi86nfY8
lIc0rnoicb8rdr36h6aUmcy1VIhYLZIuMVDFpXShIuFeepdHjSwEXYAX5/fsJQ+D
/q9isMerYe6856SgwE7/E8/Kjm4yqj9CXkGeeMYmWIn3qs1HNVmNtOcU0hOhDFrb
OZ3p2pO8MGUl7blble3BIbWjfh7fSSpTmC3w5RXNLaxTCy9DJBHpXPSe3wwb3c99
oEXcQj6+uzl0fU83KSjJw0w+4zPQZq2zwDKMM/W/zbfX9FYP4Oc/2ZVjnLCzBR5T
/4BbWHXN3y1fsDHASzRVepBH7AWiXyvh7Q4kUPZn+D4yWMPyMqWkNWocpZ4ggM/x
nyLrzqbLDVfyXctPxpXcZYVn3NMEzDdXvBv+QlFmw7jPfs96dlJtrMMm+yuE4cQ2
sdY7iMJtwL0h5ZNSuf/eUE96CyJ1BvyMc5atldEfKU2z4u+GIhnPOMicO78E3wsJ
BOTlnVOvg5+vDVPFSRssJFVnY6YznZ0b/bkiC71X0nou9+yV8B/FuAhOro/OnQJc
EQZYWz7vzc/lKSxA5blkqtRwcGlv1Qyko54JcZbP8p9ZQ5qJ91J684nOxC0d8SRj
sAkKr5CkqOOLMrbtFlvaC0kTL9jruKhaMSlWJ9aINJHXejJlEGvDuULfrGwE4lBO
0jqos93Hmv1K8MjzwTKKZvqB8yD3Esz1+pFtf2Wy/IHb+4IEjxBqV9dhAi4KTtuJ
8xrXuv6NAbTmEoBcIxTF/IxACDfu2pc7KhuQihpSlfVr2r+BG3tMTGqcZCfhvXkg
AwpWv8KuB6Y1ZegdHuu5FH7J19GffubeUQln0XafCa++Vqlt5TCbQh2cGC1PfpY+
qD5qA7BVgfQX5I3oGq01YowArbX38IJ9GBOWMPQEyOsA3iuvfrbIhDJkbiIij7Qs
VWms7hWkV+WXPOLNBid6yRrh3qkEMkeVEWg/Gqax4ux7lNqMniXbv5nJ3UvezOiT
qHV5mrLhIuMekwRtwUFSXXdYNrMX0M+JFsg6hj9Ud4k2E0qEAVIzbQSBi9x1nc5f
vJhPExPw8hHQYfD9vSuJV5uK+Le9aG98YIf59WxX4011au/ty3schnLllucjTOk5
iCmludj9VhheGoJklbHiPifch3qsTTnW52vERLccXldYL8H6njZOBBKCFuk8dr3s
G9LB9HwFqaIjgS5X5wtS78whcOAidAArVCJrdIGAxhv/aYoYY0beLxSnRpGBPvLl
p+LyQXLUGLH7iHwf8KmXbdwFeclUgZSgy78M4hToRinucidhW4ZRmTFL6qPK4Ocu
cCIfy8qXvMj9GYT6obhnRPLinSTL07ChOjUPaKHWwxFxDNie5WvXI7BekW0kmKCr
DqlI4P96tdP8gnC/cfgcn6s0OQ7nlEhOXhlsY2cNgTRpCcovnVeJ+IIbqJP1WTSR
VhHteA6eHUcNP/dlXUhaWrF6UGgpNGzAyjzFP+ECvS5hk0bpBXsK0bvdbv2kQOVi
sQt0D5NuhPfxHBMtgOCxSeQR2t5NgrXblj1L+RzQe9LhULwPKn4yM9BWiBOQS0Zp
ra8kgQg42AVPc6foJ/V9TGISdhjb9u1m9zOgCJn6CKAXr+9USvjYYPNWo2zwD492
9hwOOZeNyykITpjMpUjjSxvR5cHf8w7GBdJI3fI8Aj6vy5NrWpyEHb8sDEyWwsVm
NXvJUHvSP8naS35AugaDgXvZ18R3umuhFRTw8BL90jbPSK9mdx00vvmqhMQaRv2x
GbD8NC7hki5ZKBH8DjAXJRecj4XbONtxlhyb0Zbve7iDwmYhr4sXtzgclpFmecS6
09FYNnNWDQq6xPm8zOYw7lH/Du7O8ZeQCmJ/GTjI0OJioOZuOtVMNpIqDHv4o2dh
uG424clqTHYbjUfPk/YMZfXK6baLkdVX9yU3Q+FpNv+eZjr4doNbNl5KgoTwK7yv
iVev8veM4mQEj2qBbz9Zqodj9AWq8wFwOFHdeAfVCbUmMuIGRuQ7A77qP9Bi7QZU
ZXK6wNaf07QhAGElXh5nA504LanRw9l2TyavyAapDpBRUefU1edrL3VPptQ/dcBA
i11n280vgKQpuiC/3El7JvQXLsCHNj5ZlbTuwKBMQiGp8LimpbkhL3jXHfvlVgOt
JtWhhRu/TwyMSr+o3PVI+FD/BkLyGmRaq0v3kpljRXK0F+ptAcUqPWjG8DQWSnU9
TtAf1QKz0qFSlQqtnj1ztZ1BzxXUxb+YcRCuLG85M5ldFDpwfhZq+UXnfqZ1jEHR
3dIpKjBGw/NqpWk3P2AeZzBPxJlvw7lw1jlzQ/3bgo/ByJ+t/xZCb8vdNaZ3Y7zq
XMioVxe+1dmkocK9IBrcre6fjezQHQ+sFipZTz+FBc7I1oq1wQDFkTiHEOwScnBi
1qLQP679q43Wr60B0YpZtHyxOzTwEAwsvgkpuPqxWU2ot/KiXb/sOCv0CsbJ7irT
CUpJ3AEDsEV0JwcC7yvY1ZUEZBl9SIbrYrsUDvxxmtOOVqyisywNmv/FNsmSmIOg
DIFkmt9ZqpcS2VHbJ7UOEuhm5+OYM+o+XKXQaeSiTdjeVpoJ/pia3tgoVzElmeFD
i9Lx95irzVi50GMQ7SGKXlYJJeUkdoDs/Xx6aJax4fRakO87wI1xyyGpMrHzgDmw
B24GyUW2GJAsw0uZ2+fXiaE6XYstBxlmT1p1wo4PNYBHzH8DiynWrMkTaYd03oTJ
3RlwHENFE9B1YpXXFimdP7i/ED1fbOsTb3M20CGwHTAPL3U7Zg7LxI0z+ew2YfV7
CsXwn22Yqs/QqVjBnmj/E2jeazUJyx7kFmclQCuwO/llSjyoClSJecX/L7kEE5OB
I6icxpbNRjUsed6lwYcaDFFr9/IG9h77MFo49H5pCmQMbSUx51Gv+LOw+429wu3K
2OpnpzNCVSb6mrVqGVBCfRz3zDVrV0ligDbc92uTsbpy6tw8Tcpwz5itHy5AN2nN
hUZLmyBDBk/HCHAPFV6AYepsAJJ2ibaDu6+IeL4/O/2VurxuQfn5gDhRaB8bQBLF
dkT4jUwaFLcgoab2mN0QGqMSI6qnRiN4PXaa6ZzLeA6rcj1cjehxlNwrbueXH/01
3x6b3VfQ50CpPoTloUyu/S+tlwksKaX6mKA5SpLiLRUFCH1qYRQYG0r52kXPXvwi
h+Rf0PV2gi956BNaKiMK4JbH9nDXrLlACWx9oOmXvFg5l8GkG4gQP7taWGkXkyeA
h7FOAcziwI5np9tsneTx2dR3H8q7rD0inZvXb9rE2ruw3ENakWGlVmO42MdnX2j8
u/zBfd+UzXEHVUVgZ6RoueM3ofj5XLfxwbdaBh3xmUlS3zqgBjfxhKRznM/Ja3jJ
SxUlUbfHxpRtcUi1zKhn9y2pwQwOKxqLjSo9yKu25l+TVQOaC895CaV4PBOoNSz+
TdVKWodKQHWc8imAbfPWiKAYMLHcAc1q20tGN+udSgjAbJpEXXsAoiy5DvqGvtPz
82twxs1SR1kgixo5QByVGlUu7UdjyZDlaJOUEBS5eEYwSNVeT9eP0jqgrLJyj+GG
Pwkx8QDas1IE51mqjY+fWJHaXOIsaOBm97VFx0itrDA6+lRsG6zsT1dlcu50QeYY
E6wDMjumGMJTsTgZxz8RrqJH8JcS6YoVFoDAUw1L1xPJwNu1pjqOKnRlFYgYGox5
haJhprFUGcKbOhJtD/g7dFsj+Bb2xrfJJ4HoqSWU2mt8rc/WCYk9sbEkBn79ecwg
kT3s3cuc5wGZWx1qzPv4GZEsymq0bP5JH1GJocFJcg0DDvZfyS0KaGqusLiyzD03
Nlkl/yq114NA6RmOcxS9nZV0I8fTVnkL7fOZMxHdoCG1C3barBG4XiyQr7/lruib
i+DLSPgFHm+BZ3fTTK9pLmbKYoI3uGQWjHjSERwnYFwpUIyOhALd4Xb64JXgXqdv
Q5PE1zZGo/DmBLBePkuG8STMD91ITnao5xy/JBKnedkj+lwIzZ8BioNvzoQwnqTA
dU+Xaz7TTBgjByoyLc0SpKwvIimBAKq0/kvRnLRvSVAEkYTGRwt6HdpeivSBGxtm
SByltgFlfdtWvAzjnIQQvy7IQ+GUvAoswa7XHUqRKzxBGOgi7I/35uhWguJvkjUe
pInw3YZbVlvuT1HZ2SNDjnVmnBFlcn8IeBWLdSCFYIziU7dR6mjW10UplLARMyVZ
XKWCX0vz6/pgDwrCygplnT9jQwncPuLXntwo/gs9ARAqeD3vW0S9JG5P0g0BapH+
kdBY09oYQJLQxhvRpQbQ+f1+fT7I4gQDs86LZp9DOZXyqUSZyKdjvZ7XpcxnyaLt
P4MEWsNETSIlvaka62rbIntRviUJlmthe0zXDs6+foRK8cPN+LpsLW1uDbrx4dW+
fzRQ1mFeb3fbaadZ7YsdKowQXiGstsgc1wM/b7nFsokVzDTNAqp9iUzxo9lDvvim
zZL/KghiH1VkkUu0HbrWe0DHoKUArytH/qMofXPK7FkSarPmhz5VTeSgb6dUvluv
MWSJHr9VQNOnNZKqkaj8lkqksFovejSgvF4d/Zf7+aaVw2vyTgG6ZCYpMUBDBkBp
9bDZRoiSLXsHQTlsqf128OL4baBmAD7vpO0lKYtEdWKMjTRo5K71tAWmY8+X+ux7
xKa3kG8FMd0gAAnXplZwPajKM4T28m6YwAt4GBF7OqAgniu/MT5tMGZ5/Q971h8o
q0VnreyWZ+Z/D7Ikd25o74OL2k9GzbrRCp+Y9eszm1fh34Bs1Zy6n69rgkhZdOKR
rN3Z1Abk4JdDNey7M9YxCJF17yIKw9qx1E5PKmGsLZYLbcPRp61FUJYmuefpL+lC
7dE7Vd6ekCwqDB+Nk9+TdskZMGj8kSPt6zpWSoxD8tIZmdWwAeDkiTEQiO+qpq9k
dDITqkOrRrw6C9ST8BYDQzj6arVRMzVsLIueoam+vAhOzB5CLo0VtTy/KKs12iBs
BLs+6RlGyCdeywkuMSUkG1E3ZJeBBNZ17z1n6tGa53yDWCB0aDpxKgyj0v++xKI3
F1bORED4/ap/Hu7F1T6JmPK9OapPVWtYETnNElbZmaTN3uH/cpkzD7Z+gzVIg1et
c5/L8fiXSldm8XbX9Pj2wb7i0Ri4qFH7Kocvjmgx2V5+QyeQZk3Xc1juLBx4ME3Z
OIi9DN4VMRJki4yW+09z7Wp2ycK+nF252GWXrYp2mzU6uTruZuJqaxSKJIrGuVxk
usmtcO44eeRwMUAcct+Iv/MwbBQRIA+D0tqMPTjZCKTr5ze75pGM7BSmrAGXJYS9
MkKd/8xLZmPfXqaIk006ttJCJhvl7PEWzunmNYT74qChgft6OzaocONRLlOkrQCf
O6wjoprhA+OsVtiaaaYW1orpP+m3yHUOu6PxWJU4rCWsLBoHY1a+Ry2LFtBGxhuu
lJSE4iGGdXThmIRAPOywp/0usC13kGgsWhjY39YskYWbLIQsrv8SjCkxPjRzAVry
TTS7filbvc3xs430YBjRhu/CTyYoC2FzqwMDCAJs5j6tyu0yy+6+7OTPymTm19A4
rhc3d2587S1drH4wwfBnGyWaN34p8PTKnjYNNzBBQ5KY31kQP7861UWOj6bGG8CV
CareuEGziz//jHyJHLClg33S2d6qsZEnBpkdvlC4QGDj6dlSQU1zbzuox7xySmRI
x6MHl37eogSUzDisYrEFE42aSxSAsLK+kIjkmr91tgwK9IDh2NtKZSK+JLKkdjXG
vK/C5KS1EaE7rlJANT7rQscbXCLK4LxS+ccXBy9AR+nUpN4ARFqnzi7qzybXHFkr
o5xxmB3iqrywX6/VpVOfMTPndQg4FZnXNMqtx4GZ/m/chQeGDNQgJSP2s6AJuenU
KASGKFkCNPwzyORe8PjwDGZgDwinTsUESKJ8NzRBPOn6lx6pOSypoBiTFbR2iqwZ
BkyfU4bP6t4oNIkYwwuSdZOM32fsP+zuVekvMdWFo1YgZ8XzBCrZKrBdEk/0TG6F
ABDbvhc7ttZhdCxu47P7Yff3q2UmoZD3xlY73wJKLEbddGaitfXnv5CrL1yGdmim
fawsbGDmMPcFV9WBI2uQSU69P9skMY7bNDev/WP5euouZCPG8qdiEGmE9tp1oJgp
M2UuYe/Fr8+9faMOsnakbd2rQkOrCmIJiHzpV/lStFjwG5Cya50gggo0QspSPbOu
hXwbDermv1AshDNW87q4s4E/2aag3TcAylcDbm/wNlPYD2EWCwgcxsMBQHU03/x3
4OVljpYyDU3md8/M9X/q+0s9MkXrQmnJVqeAEq1Ut4UYHJZpm3f9JTQmnNosv71N
cE1PoAVKHkqIoHNBsoQ1a8XtSIRIfDwOme9F6xuSu03LKAbKck3jQBsRMmr6SMvE
x89toGsZB9/UfMIx/L8SY9N6DrFmMImm9cYrQTRzDoSZqXAkdh3jaZ1fSUUbf++l
dR3DdTINX9xkWp7nYxv6w4DqOb0AAWFKRvZg84GLPjktjx5jsa4VZGmDRTga85Jb
FbtUYZJspm2aZWb/ce5gVgECxdXDqYtGVamBjS7wbJ6Wo+SOkBXwcqLjwI+VfxkB
67Lh4NK5Jv2qWq1KfolPEl0VpJcbtMzXAyh4c1iANb3OD+oM1wxBXZR9ThfZYxuv
CPxb9hG2400ouOh09iEPzj5uV7/ZbHHUcdbKu6F92CbVnAcb7k7t77s3os2o2VQz
aHlWjy0ZAljJMzwnYy5Vbkx98ovFy3YcBAHyYYqJK1FNKXs5A0Al7u9hJl2LTFP+
cgHyPCFdg+1F20ZaUmqEcVBxIinnK2r37hSyySewL8chNnunFbrsp/drQEsoI8nW
gxYD83vCNYx9ki4hhVTy1WdJPsX3P5PGMsPeM16WMMIegrAtfSbszHkyKuXyNDgd
o7gI22wwTESENyLPcTd1VgWzWOZnJ6ZLKFXFfKNTebW8nAA0M0KkhkHTSF/K8nOq
h/qP5pjyZyvsHtMFYASeq9qZksBYfKURV5a/bTriYMm4nQB0hxwexzP5lu+Zk7Ih
M8c4CxfipCpvsIBHKiLsMh2hE7ff0DH4pvh+zQZZK1g37dEKU8aMsrOxY4ozYTPk
ihZ7sBOXxP/Kl9BuMhaP6lvBXeU5fck3+GPIFl12+AalqsZmuHgQz1hocLjiXE26
rifKhGa1ghLA0ecsR8f1KiX536p5qa9W0r0beFMuxXPmZaTv5j4EjYL9UUHv0lY0
XJPcmpSZO8RsiMxivyl0GeDbRmJW18al2d79yoFPdB4n5W/T4KjbyfB4J2Z41x8q
YcBgeRIkqSOhezzK0WFKumwNCbCmh2/vIpsWtkPu1ib6M6P0Q/VMxnxsYiQy1YSL
4Z8EqFakZSuJGNlkG/7p3p1v/8WBKy00TsI40CiwA/2YpsKVE+/SX3IHUe40+Gns
/2sHU+wrNSdoamhfYmz6/TShHWn0FyVBbF1cxWTq13n+mOhhiNTiknNwr2hqWKcS
dN6LGKi/7gGFy10ldEczpy/pzWwj+7fhZ7FMNo3uj3nLkbV6hGabfuAQcKuPx2il
Y/5v+riq/KOvOVtwq51ovM06Io1wMtsMPzz934nNSZ07dsGj9fnidyztzFYV/nZi
rAT/LE5fUySzaH/I4HU9TezFU+gOeGubxatdj7Qd8sT8+OKejBcHDb5SjoEaSBPN
7MqcqtMqhasb6NADuje6CAbMV6oAO7q3PkQTuWPV+/9HTP8XnWYpYMszph5be8gX
rJTWIJOG37mf3fvgovZaA+5vYurANi5F7SIXHKZMEhUTjbGvdVm9QJVPRbX6disJ
Iv5YQ7P8meElT5UPtKGRzWdR6D2jUnKE9KpFZl+MsdBlVwOskJLUjHe0pyEgW1Z8
aQOLP0HbHjTk83eUH9uydUFuy7Of/xtc5YAS2lKe0p0msCa2NtDsymn4mh5K8xQ2
dhZuSzFQAwiNi/BOEJn/AGPvMAIrOopWNdGpcRbL56QsduPt680hiMYsSxfqul3U
rSvHCyf0tVqVlFw2uIQesxIcBamMA9ghQzPM5Odp+EhwkPk5HKVnRfTa56y4xlt5
5cp/6RSzKXo6Vo5Z76DpkSJ+CRU3tS74RRpLf8WxShwC3C1AEXcuWsIkg6fEGd0w
tkZqEl185Vr3KN8o/5z7Ye1XnvHMKRdUabwYTPMMNQZkRTSfzsGsXT2Hy5Gf90e9
wU0/zFFydQCUg8vhbo07BQ7vdJdI/XHAtQKNR7cDuOU+XapHZYQDYl5GAFt2ve2C
Mv6whZ8Nx7oDHYyZQuzyjPE2n7C/yAgAx47YkME9c0a8rUPhYA8Y8qECvvWmLwJ9
b76eGPAlHoMk0JtujT2LHVE0H5OJXw9MgGlTh6+Rf5Ehvo9iJL+oNctyMAMptJzM
mL1vFRP7bxiGSL1uKOIIH4T+NFkRxjkKDo2gXVHldDYkBOJgrUdZjzmGf1RJ/Dvb
bin4RhJrCdSPb3R1EUo5qt+5xbMuPz6Xn/+LcT+Dcjr6mp2/ReP7P0lkA75cjliI
X7NkLmQBZbeplU4pHpIUUocMzek/jMIV9nddqUtJjMQLa+Qelp3Gnh957TIpE6co
b2TatwtGVF6Pu/i+ysK6M0LoQCpSbTUIs27jmZGe55IMVnDQFXEsF6DfVMjSI2S/
8ZDnCAMwHRBEyTgoBmJNY1tZX5ayi+xdYaJ4o4NoDUob3ZXtq5IiSteonQSo8lWU
OK4SiqlXF5+PeszgesY921k2AAbf70TKs04ygVac0bISVi2V2smuj0P6hfav9seA
JAX1aKbtXlR9o1hn0OuleNFH/Uz8v8kNJoWvYEpoisn11UYMbjD/bLdld3LyZYc5
yjfHAQOI5VwggaJhRAvOyzDio3YTwgVi7ruMYltulGHcydwJikGzB/UY5JJI1SAI
WPqU5B/nKfaZIuNL6Hk7oKMZc84n15psXazM+rLQfEJ/AmGUAqSoSBV1SGW2UEil
9nwfzYHQDVU7Kp0VeKHBQl4eHGn2ipQkMvH5DWiFyDJfgrlD1LSOrxvRt20NBb/N
j0a14aNH/yhkhwp8K911x/mSNeaxWIIQLM6XqcQVWM46xhVn6yPtKob5Ls92G6VU
DqD1DOmrcYeXU2Vh06OP1ntJHr7D+qoKGfD7IkEabrNT/qahJS44K5DY0dQvshZr
ctOsjbaWR6h9A6MTzVtu30qTeLcpXASusGScT97cx/6iU4/uBXTq4Uuu/GJuVKiu
ZywSUtmxeyud9fGL4YdbP4oCV8L8uCTUdT0oA+U4yyrQzribENXFGnsIz7M7Op8N
ft0sr//iofcHn/UpzSnNHFGDLoD/hWnIw64/kSz/ExCFz4n/Fe9bVGS8sByVGVrd
0rb0qf8dVIMO2uuOGhJpGbd7Z3JSkVWS6UnyYDTi9hFRjLqs3rqQNzIZGVYRhm8U
Nmk6lYuJ/ZamIASE4kt4qsMPXBjO+20rx+m65gq4nwGHz+bddB0vzxaQlCaxj58F
8n06nK/3W1Ho5kcvcPx6WYbiVh87P5Dm2sgIADO2gZ4xCuZvrPWp0pRVGNjNEcLY
35SEQV1/a29ZoITaQYPHZqHObPEylYVkLjKyLM9C4a9h/tIwEf0/wTJ3oOq/q1Wo
yRCh7DgQeoCMD+JLalIqmL7DFwxWtSRWIDu9ka9vvqMK4lhhesE1LPmuU/BK+SGr
e1ZVkDex8B9lgPmk7QzAma033cAbBntZZgi2Z2zuV8a8CaS9lzWrOvMQuq2s/w6q
Kmf4GOxd55k5fCWKd47aRHTuIGPnulZ3CK/0Hbib1tEyKlWo/VC7D2sFTfjYhi93
cv2o+uJCbqpHbnVpraDaYbCIxnbbppdhQDxhdsTbv6Y4M/+nFO3n3LUMxI9iK5JZ
+z4jCy7vOjDTtsj8mMlAbjEr2eOW52S/62xe6oEiVINE7iHTwCsg0MXFSN8oDwA0
YI/AGG+dzbODQ3GdNdYKzWPWJIy/cJ8ZU+owmwQ4cEZEgs2okV1AETBiv1ojiqWn
jGxwkbg6LLtJlUg1bi9KxE0lM40NxwwzNvQ6yzECJxPjpcWKY7Yo98yomCXUPg4g
JP3lgGDlDVbPYHtOclyh1jftUS+9Y8SU1m5LwfdB8XBbheZxAZZ4ltvPt7cyi7oj
DWwRDAiddWlSd1Ks/Fdj42egJwC7fG4uT7kLmBxgzzAUWrf/Ra91upvNoLCJtnbg
xpP8tsmoGm18O1ZbQMt9QFP352erz05Da9KtwVc4sIhQjnMO4jXEyJzOlS9G92cv
GqB9DdgAM0EO5dhHvg3G277AxPolukASXwzrP80KN/pNQE1vGNa8XKPhjDs0ensP
uqpEB6UsUaJnDFIAvx6X3Ax62xET2v0Jo2b7alQVXeEbXDa4SVpiEX/dsA7PLFq7
pZE6XRNxIdiY4+TAVVO4IUIbF6YZZRklD/LG7Tkr/GAwBKPJ5QlHrVmo221EsmBN
szGniUtGAWAnjKEHNnhZqkYjdYIkuWB7eF0xe6vTJcXQTKXDBm+x7jVkxM1966//
y4GlKDPOM8SsMdUonaCh9s6Yz0y+KKsPKAXEszfe/xSzcGMHTcB38XLqdCFg2eDv
ZsZNir9C22nSGya4lTn2vWTh23096LiKwydFBAyEMicxM564PysCuPnqaRv5ePe2
+amg9jnGbpNiq+Y2LzRCShyorhuF6LhClSw3A1DUhqolvkhGQ6tY/cijznGrnrU7
jnrQajUGyiCfor3svl7IrZMnL5KBdnzYoRnKc5fBgnkOme5jZcGTBEjptKs2ypez
Sx9wHaf5wkoDCsfD7+h7CEPCoqQfHvNlb36BK3ZA53UDkLPs1sq0JEDtDsW/gnh7
7m2Z3H/bR03qR+wxb8m8Na0Ow4oSo7p38syplE8fbanB5EQKPhhwL0wHDSNR2B2X
8T6D0l8uanovIIwIU8uFC05pqQMzu8TMuljVfxe14wEZRsd3Jcc6f39hE32GyS/D
NN4YAwZ/Yis89fVdQANagz7K/P34lPuz9V8CzLMwC9XDPZS/0xggANy5ETnaoCh1
lfhl/c8jVpfKBuhFrwMRmI90Zjg29WfZQsPCeIfkEttJav0FklFnxH8ypoAjfoXp
bIrF1kdb09WWUzv1zWXnLX5mo6j1DhxT3C+qwYvw8qZuTKalYQhXAHL0IJ+zuR7j
Qlj3116sVQfp3+yQZrG+dqxnDn/ZkQ1c4ll14TyDcSv4++DNRDC5TEkqsEzUBB2H
Uq+x6rxIkQwewq+9lm/qhmQ4k4IC7iHdWuVVO4fTl0KH0uJLh89airdEEoCGoyZJ
XlWquuaHC0IYCydkbzHEH/0kKaHcxrNrQdXyRbk80eWMvbl24pqMibQHCzv3O7K1
q+C6jKKXb821iICOFLhc78yJN1Kr0fAzKhtewVjILttRxGd0fpfeScSgDjuRIx1X
E4Cf/pYlwY1qMbrZ8+K0NVwtMfszfBJEBonC8r1HzDwhSnqIpNR1NWx4+iEst918
la/t8OJ0ZJpOw28UmkbM18xi2eGV/S/mS57iiDK4IWeeI34Eps4hu8tW4ULTFe6E
EkAVXhh6zTLDb6aGkegYKyOy5N4+eGK6otr2x0cuz/TEb7YJZu2CpgildtW0M+xL
mpF8FPxRiYL1gcYOc4N/mLc1UNmbwy2mwBPRgfkZM2zeq/snq8TX4ZT6pvuYPFYl
nqXH/PHWWwFegP4eNI0MvPHQ0GKBlni84wOjjdnxJp2kq2S6/I78phYkWD+int5D
40KNv6lQ+gyL9EJewtBovQjs+l10qBxWVFXn1klfebvJNgInXdfNyRq/sih6RDoT
D3/BAv5uqWYX0XqK11L01bU8rLuqu2xiQQcFZKwGTF+PxvFPIAqdbsJS1oE5u58b
LuK6Ew1tJ/lUh4wEjCTB24+puhdVb+SyqTka+tt7vbx8oZjVCMi5Q+zwcAq/r0DZ
JdaqYCWftIUq92e6ajx+FVFgcPc681Pj0pLB81F9yO1WXYsU5HBWVxQ4ETwZvqWL
IYS67LB6XzLBsp8HSvs4pr6e3cQ0fopKypJjg3Pt1QvDT1kk+a2yLzUz4XoLWAYo
GGLunHSo7JCJe68eU5GF/6wLrZaEF77RYYPbRB8sA84uLvIfMuy07f4y5is2exT0
3WgM2pWzwogiWVKfuGE/E+AN+V+pYsT2FtHvlhCIVqktQb8GdrOZgab499AWNwm/
07cMw+yW/jLPDcVyF8uoaJjE6alqs25/wIUaoINP+DaL9uqE18joY9IKM98FP6EZ
lulkQY0s+OIxEwVIFyoytVdreuNnu+s4nNrYSsJImnzn4tDmmw8RKqmg9wplzagc
LUfMuwcNuBYL5GfJNPFY1elZL/ZMUqRNoDja3xhk80eclg6d5HjcGBLBUy4h7qPU
boeSXd52DlqX/o9F5t8VoGIvlMxt7ep1cHFkwXFzyIGkV5nYBKqsJmwXz5I8Ut27
hk8ArMxiO/uCAQ9dGp8PiVALWl2JmczQdukDca+HUH9hzwOU3WA04/K6ACSFby7V
Nnf3DwzlqOqEXNXhkUTPHflZKmEmxt/fklztntP6JQIjKH/DgOjeUBzXdoGBoHPD
WEC+4dj2NuyI+bFt7BIoZDWzHjKQ0UNeg063BjjGtkwBZcwXxhVK/vEiSnDDo/Vy
NuAUSW8pnNGMJyc91FUqFg0dv0n/0H2K1kPe97gWsvCR/NcsoFV3IwZn8W4pw8iK
pLKaSLfjF5wqPiYLoq38XLJZkk7EozVubH6Vsi2XxnbsaikJCkXxtYLMn8SJOAhL
jyVv/fnQzh8T6OMnqqVpAN1mmyvJAJFutga9WvJcQ7FmU1NSW2/VBHhzQ+zoAaDC
lKgEJ5uUHqVtfpqBjNeabCfyD8NzAlV82SboPEhChUIj1kU/o3XvM5jsh2TxUizo
um+4KQdcDzKkZ9e4WiowrLCfqu9uJ561BbpONS9kjMQvXSTlpkGbFnFwEuibyvJZ
tkposyi2Nvf4Bn4SXy3gAl5UMfMlGIwHHqzpCMPb/ZMBOeYBi1kYk/RPaZnTA7qG
1ezqrRn7HKui64WEH8sQ5MzzPrjMcjm00JMxk8wpMprB1yrYwR9KPwM5l2ilJiY8
P+ESfFMlGb1NW0TnJKTM/jriNmZbxxz6H8KyX7LaJeVt/upMr9Ay8BIRgqyYEOUT
0F4/PrgJvn3FAvwA+t4B2XPKvyDNDfPsAP7S7E0F64lhL2ezOzScGHD14Bil7r+D
YS/Qi446UfjsGabjw+6xA7Qt6rA9+DhK5C6F4TotQeV+RkOr91oKvASqmuW/fm3/
FtEV+uOEDURQmb1K/fNBljhDJRBt9yVVmDUKugUa5MFwMVa6/z9DVINhr3+LJ8jP
i0VQzeXQupzTxiLdeCs6UJ+k7Nqe8l8F5eP5nLqGRNfg1pOF44MiRUhtIvDnR7vo
VN3DIPa0+b8TcUD1XgMhi524iR4fuC4tCJiARjMhHWrCBqvwxEKwf3UEtoyQXiLR
/+fVyYFSECyPP2RiLALTdctTrBf22zKbkIorJ/rl7HOhtFE9antFZsX1dZUIWYCj
ksL32rIkMXqCSBBGAd5PrUVTBNJTbee040xgB3lLdQ8zOhgYtbju/rbxnlk5CznC
YvTFTQ6CCeeGiHfDaKfzk7yeezgVvF4pt6gGaeCjNZf7GPrTDiZaZIzGjuzOYNGZ
mkR+xV2x0nHhsr0AFNACGAdlct0aivFwEq0KPJoQ3K1rmo6/IazU4kCWx0iCjtM0
LEAH0TriPwsUoq5HnrtYk9zuwxcZH1TSQitIyznNPsHYHSHepwRwgn+DXLYf0U7B
1HL6BzJjiw83b5/dlwqx6Y9Ve3v/zqJBj5OQcA2BKPVIcnYgTQUhgGGXIcTv2B/0
EBxqf4ftmdpMPgJsLjBBcljl9o+bhXyXvHeGQN5vJg2spwsUkdXfuBB7CGRGUuHy
s4HgTFuNkoYbB80rbllTYpHEpcTcILIzKHLaADEBwCcXXRfnHwJ2rgNzMVKeey8n
d5+kc08eADjICTIRorciX6iyMgnpAqDRRA+GBtv/gNi1kZ1bRdrEWYAdu1FXZps0
LhJ01D+Iu+QXqxnoV2jAkGQg9TadFbWuaOBnHbokswWAEPnhdC0dx/qpA84DMIam
IyUVvzcLq6Mvjbkpef4eAfP8BEWeg6Cw2RIK0TQUBqBOShY6UPVne3qj8hyVlltv
LbXqyd+i5lz8SuH15JK023hBUka9Ub2nS3wumjoZ5Ut5HOdoPv94TIc4go+2Y6gi
g13eloha0L2d7B1u4rOLgxBrmpWifLv18/H2/lf+iHCSOFZ+GdAsvIKxxuupUpNT
A7avN3K1qmtoVdsL/SXHBVDGC1FdimxF0mnkGC8QopkbxV6sYMD31i+7A2CG3eYF
A1FD7Ume1g4gGWbeC92H+rVu3Q3z0vG+IcyhHbcQ52qb/wnSZtpAGXdpmHTqrdKY
NjxotBiFi9hliPAxmlNVX7zSPseOxvEqCnxX8E4Ts8neD1M4PwNsNUkmI9E6rJYC
K9L4+Rd6LurApNhOYzKSzbCKvExQSga6SoDNsVLyXbtTqdy4sYWrKmOASxmLzfUK
LOMXVy5HjNj5xnnAJjMQCfmM8hElaeuH58QbLiTo7ADNCbEveUVT7vNMW+d9+Zdx
KDkw2TSGFryn6zTWwz+RdMx9gYH9YjbyGFt6aTKgPtB3dvoAPRuYXeqoNjCAoJBL
9L9w+MWE1QGyHzSPOWICODeNtPMdEpaf2FJ14ELW4fGQhU1KpgOc5j56YE94CS/s
cvOGXWMJhiY8tu0nVjl6HnDDmVm5kEbjjcRCW+Y8jlHouEt42Bg8Sx+JXGdmmP2j
ffPw/Ekg/sslPcVZt3iDQX39UyaAg2Opmku1vBceLhALBiLPknmgXfj23M1yOUkZ
AdK7aOUZngO+B2DJvNipEriZt7KD+VpYy3JfhcCVXl1xlrM+YPu7UgAHcLI0PQkm
e/qFiMHFsFr/WGILxJ+QCgeueo+4usOYLYemqHOcaTYJg2Z5AA+rupAwMqpORqNA
/si30HvH0pbgH3MMweq7Mfszb543IJh2CpKInS4Wk0DAf+IqmXjyCzxjMWRTagSL
VhnXGdyOmWwzhfIAxaJ9SNzw2GfmrJm0jXGLA1EJdxwZHGD3ccNi4GjX1GqQPEOM
LpKNN3Ax5MTxFCjhrNiuhY/fvgibvqJfiZZ+uHvosvvLaC1KuoPTAIE6mzR60j5i
hTpOWXvYI5udfJLQRWe6LAvs0RrQMZGWqBaIodHM9w2WPwt56e21SvyhbXm/bba+
KU21Qs5lbTK+WTJi61hWXbOMIagOspLj3ZSnPXQ9upc9vTBsmroH8ULEliKeHR6k
V8oad2FCaymwby68GpPMPHkb05Wos9mEjft76YNhNt5qdH/0A18AvCV44u1iY9jP
gh2/n6DAA83z1t/gF9prX+uvyohDZuimslDbNWvUCQXaAMV8fy5sXeSo31W5UfxJ
L35B0e/6kNRmElaM2rsfXoJtR7ajfNo7x3IUzOMEkPMaqH0ti9i4Ftc6yWPivfHl
2zjp2sIcw2y3LWbKEd9QggGJVne11fl7mA0cb5UShfXmVfYiVpCQwXVfEu5UIM8Q
Goqm19w1GgxA+eZcvi4h2R/aZ8+VVpQjWj+ZAUcvu44Vp8onLhFnxunX6tzTUYZM
52UvLPqUb/yOXpHUHgi6+Mwh3MeoAd2j1HSbE3QO2s4tqdWIJEOIzhOrWyhMYQNI
mJ16+peU2sPwUOlErpY+R6OtZRwHH5Y50KNtSl12jqZxn2RP4kCqxP4ZhgvKAhWN
e/GDSKCVuhsf0wz93FZRgeZPZLA9TlpxwEickSULxdIy4XlpR/MCaQQte31PY5jC
WujMXHs0TMVH2PIw+7ltM1FvwdczuasmgAJWNLMdUvQpP1LJv9gIMrWe+tMnh9i1
Zhhj7Dl2gaysdMHBMbblbRgrN+6+p2VSG5CPTUHVafUWhfVBdSpbB6CH+TO+TREO
ng7avgy4wfQdWOe3L2DRwmnFGY5JSotNqkv7WmPSafGIGwqx+4zZwR4m3lTFUw+5
lIQ/SHJWFW1SmBgRe0yVHIzPW1TqMY+460YQaTP0XCeCFBgg94cfnojp+JkU2wx5
VR7URkGKgxBimiY5EDjp2t3wsvNUQMi39ZLy7oBVqUtXm6rZgRM0HP9JVJGKzoP6
hu9svT+HS5s1ztvo6qMXVe7I/eVkgWiRYKOTR3Z1daeXpYeX/EU3NyYjoObMJ9Jh
aEhPqofUNndHyB2U8ow0MtPwIbSS1K14h+PfG5GLrNmTJDXlVSPspGguwO2NbDVd
x+tU4XloBk5Q7Po6WIppNNFRVJQm/H9oqPCmC9HDw8VY1eD9Uv7mNDGZ4tJBSoTa
zNUJHjpyDVeYZi6T3PMQ/1Sidik9FKxetafvyfyrzh1RPVlWDn/5qvdUzggs3NXU
zvg+WhlUhfj6bsebwOWVfjg7mseZjsUgzyv3DfWi2Eqqaiq+0gh2Tbhh3+vlToNB
z7yn406JQDURxYLqff81lCg5El8/DzK/WjMGR8u1BWhkjJZY9pVUCblXLaGVM5f+
BNnpGter1VU4iUMDPceY2YsgA541io9Ok2b8fX7PobK9z9AgobRt9kf5JTvXt82u
gEgFsp0CXLT/IgIaRgSCWyj1biVnGy+hPfZHfrRENqtMsVPimq3eVUg1huYO+D/+
gb8dvHuFVBC5V8yvps6+tZB9YVDzRQLzL+YsFsu7julUMO81u4GBXXbCjCSRL0O0
T0PU6AqCkie3MSWpc9XBEetYJls3KogpS52cyha60alV0j7hnv7/pXs5sT47gdfg
6YMPihsZvfHcsnBhlDpZ3/DIXGD4eISbfI8gyhXrl4W8AigW2ovO0ASi0vmty2S5
lmJhR8y+h43F2hIJvIr1vv5TagVimlNLHos+cPd7MxaJghkgP+HY2TuwW5Yi5WYs
50t/ioAgklZ5WHC/ss01iMW2FZLJ5tlPE3nBFu5XL+omiATAaxfxUSOSptE85Moo
HkU+u3gCsSX8o0l6fP1gpmd6uil+zKl38HK/YXSYzLqJWAJEG9reExm56gMeU9Gx
DsQPVgxxfFX/w5f3UKKTkArkSId0ge7yK80dxGJBe92c4RQx/7res5MRivAbHWYJ
2el4jpLnnSCpy+KG+3QDEZXNH5vXzF9oItrGVSEdIrRvbNxHkoDLKp9mhGX8rY8C
wR01ZvtU+63LhekeLKmEkL1lIDPDeXZPEcAGFKOAn0uMIDBf5C7K4YqbgUNS7DF/
hcSCe1pG1iQh/g2kvD6gLo/xoWyNQg6nGbmYkDhI9SRhZlIe7AhDWPbw9bEBhmO+
dM4v7kw17ZGSqaH9nx4o89TMiDKzLYsYK8wznYq/BZwhhfy9mGaA5TaefrCoVevW
DBqD6rbkc8+U3MWwolAKThTobl1kXPeKcaVwWEme6vE78+TON6w3LgSMCIC3XDNJ
ulAuKdlxOiC+E7GGw2kqwZM8UUo35Sn40dyM1bOqe5xgMbJE3wZ65xKUl7XdRw8e
z2JqIHAgIv8dQGYe+7/wJPanjZ1pmLrjYunQw4EvrOV2OzEv7TbZ/V1TwMDPIiUl
D0p+AVLV+09sb5wJsTlTUwRCp59wPI/RwIV+ZOiz8jpQQgG03S7MZ3HXq+3lI+xq
D/vg+kxkc6JtWm4XQUL8/GI7K9vbtSRg8PBIgnXRXcNFuM7d9Jzc1KhRmC8x/0p4
iWJ26SqgF0NyqsiVQxHN0Ng5bR562p53o3P0VApGHtMdqpyAGr5zQMHEdCXTMlfP
bi+2msBQbEEHH1bTRhYawxnQT3HKoKPfYNdKO7kGJLc1ztPvXzLwie8ChqZtusHT
bT/qEvN/fuef9CSQM7IHlK3yH1FntKz4yj6oL/dilN2DLuCls3H/kpt0UHZzvMfU
16WNkkC+92meS4y9Jwyi/C4J3LYuJ5h1Z7WhxHgBI+aOxFv7TUzqObzUlq/d1GW2
0cGcHvo3tuylWzlA7/U5iJWw67OtgzfFa3UhaXSPdTdooqpksNDNbEyX0FKYMcTl
e47NFc97xZ+ZH5hk+55mRhjM0jRRS8zRP4W81oD1sCZ4tR5p6TelayR4KYJ/edBv
uvlg9plNiVK9RfLTVCdMIE8g9MXDP5GZ0k/LlLrmv4goOVPFJmJyMqSIAsIci7r4
uS9TXGz95vyfP4ztOS87RoI9aC25EeWbk1aUOsx5hgPi88od9Qe7+MVt0Hf49ZAa
5c1fAxJuO7vnDyVb845wykD/zE0/0PuuX0/MGBtoRzU7vpoo2Q6QNPPCXLVhqXoR
7VEYGIV9zKs+gpztay/Zeq56JGE2T5mBxR+mUCmMX4zzcdy6gZDYD/F6u16wHYu+
wu9LZn096IsN5r6DsgBIzrDZ68/AKhRSHuZVGD3aDHqGh0sxnAVYPWAzstqkdUWy
eqf78JYANhtX0hUq+ZmeI2tray44wbdsbxFehg1hUaitnprTeCuDK0m8KQdYniM9
gP1UtyEZ9q2fdQ4pSMoZ/Q8YTV6M4WnQf0y1ZNn+y+2Tal3xkHhV7C3A/rOsANwr
dSXkZl5/Pa2dp/KD9wijyuTjp99mG3/8ij9t3O6sxBE0+fu5Bhn0dymHUyu0Xw5w
Ni8lfDCT9RQySy1+fYo5LNcHuYPHX2qQhYNTwEVjJj7aTNE10zZs1Pc8DqYxVHQv
N4FVsI8lM7hXUwFRFwI8yK76oSsEJfZmp+TsQ9MomRhwRED17U0OundTY3mRFser
1e7W2X2JEx4ZdLz+tLGZxAugEH4IGWXzlkTADXiGpSCzugpdiz0RLLQiH+VHU0gM
Ufhm2xeOWt1A9aWL8W8m5n2eR0UnkPCqy3epYS3yrxcy1l024Mo6fdAANFZfMd68
5+cNnkybfrN5jWIlLye7RFoW81DozSSwhrLYKGJgUfCW56lL5WhOHV5wXpuTWNOe
8fyCz8nNto+OY0fmF9hm453rZP++NwXDuztc0zQJ060Wx1FRgYl2uK1hU4rjA1lY
yRye/R+rvAQU8rLlrp3BCy/cF3D9CXXYAVUuqHEPKNYZUZduTikClpqwLUjHvOXS
SNOA0Hvktlk4k+2YGnI9ge7pnlrvZHC5pUv4Zp/Rfb2RWC4QHyHmCSfZKu0RBtGF
7jWy8E+w4oQUDzka+RzZATSo71Dg5zg3r4JEojCOImDSl3WJ0aZgQ+m7wZAw+mQR
8nyh9MFjpDqgReElgmU4gPOIl/HftlUZEhBlgRFc1Pxpmb903X7/1VNP7/+bgoFM
FJQgJdqNzyaCE1uKgUe4DEFZxTkNjo035l/nXErfgR/CKarXf8KEFPIh+T262eXx
HWDKR7UlIxuHPU6+LOUr+uibJJrgn+c+ZKxVV2TtIGAQWH6Lwk+8upgS/Ds3HZgM
NF4A1WKvmnWDdg3wm47AFlXkQjiwHVTwvqYmVfCfvy8JPSnPOrbsdtBscaMLk7ky
hhXa4HsMCs/oQWB66SAkGQRbQFy/Z/2FU7kfclsriu3UU7I1pG2sGBApADbtqFv7
ELcHKqKrjUWkOB4EBgsk4TIcQlQvlWMMox6UsW+FAQlNIm1SZ/J5QHo0lK4iJ5LM
KtuRlTIWUb2c6gW0nnyseYQrxk1MhBWUA5eFvngB4MG0aURhP6vxIfWnI8ylnWUd
NMLB23bFE7VuJVpJBHvNPKU1L+abAHCxnKLhPvQ/1YTgzO92KD4FGm+ZbN09PV/k
X8atlNhIcHPfRD8e2DKi6lOeqDlOw1EdUVDNccwTrjvcLDSM3UrWbKVHhph9TLso
MuL5wHqBDmnrLBJ6c4RtPtzPrFHJgbVsruZDoTPL1Hw15Etdu9sCA4HiylXU6vgt
K1OgYlzLY+mD81/098b1RKj/+6hmg9xG32CbbBmN+Zezn1WNYL6HG3dOB4E58ymc
INHSney2kZLF8RqehgBtRzcu28Gxbu5MhDo9/P4kwb0EG+FDArIx9tWGQu8wqLRh
aBhh87JDkYVHkhKZbu7LgxwHu90P1pgZPXlwExCcDfIaGgskVgKRbx7Za8BTMiYt
uxvXYAhxbQ5CKGfu5XGEwcmA2f0pyB0SjBSTIs6xg9c5I9eVRXEB97bJIbLA6ca1
9Gr6MKT4A38aBlNr7jg/Qygx8Hh68IpbiUkZv819Y2ZFRi3YpQ4a95ItOABPfq8B
GLrw5C8b/u8Qnr1Dc2zDiz442/UlIczQqQSlfRfhtY7Qow7hQo7/AxpFYE2F7YYC
5mR2GVds/nwWCbjVYEeclzSGpyPnuXftnbmeBuBj2QnGgUFuPoVcclVHrmw4xCsU
RVebeGy+8v6ktu9XZ91z3LYWp4sDqzrS0avykpiTVF5Ew3TSpYGTEbXul+kjEz7F
ctb3OuXJvklCDFZnBgPr7Xh1nrRrs7JnqWJTGgiMfKTNBOcw4X6E5w6bbqHMwWwJ
sWGmo9njISp0iSlCxhcwu8I1krX56xtFJ+AOULcA7VcV5J+HUlbT3Ym3OHjsOLzw
KLrMulzafUtRnE2s7Jei3xwRXkNnmNRHO8vwRKz59pNZT+rAPziJGfQ+Sl8aBmMH
/x4Zbk3P1fLkJbxOaAgQ5aioZ8whVOK5wqgVK2rxKveOMTE7eFbRcqqQSpOjNwdM
MVih6JPu0LtcoXyciu3gvea3raHQxxmq+9lSQjVxJ0Fd9cwK7m0ChHt/QTSfPPbI
Je0DyRhaHdr0Gbi7nORgs1G9i/b/hwdkAE98j7VaB5mpgrx0KIprdYDRuK64avSi
9xDlg8VDArZe8ANQOH6dczZ8iQoIdAWNbjYp+5V85IjhSwMrNEF7rSDSINc8S5xn
l7J+vuWB85yaGUj1jSWweEzaowVngNcnLl0tV6dJ1wI10azmVeyIp+k1OCTqQQAs
8WnJcb4pgwcy9bEHV1OwVhcPeWT2LBYKed8MUMO8WxH+g/kerE/d8x4TB9tZAQZl
znzeC6HWCfaHjIYeKLf/qAxi9yOHQaU2NbAXP9V7zmpwsrnn/Njy8MYH9h4qsq55
w9crVLnBSeiOpyDt4Y5ftuJsKFVScekIhncKkWsN/1TO7eVhk2hn3TMM+8598lQx
DxKuntFYpFiDNzcfdQUaUsH9uOpdqba40KQfGxf08cIFsarBSjFNa38KfY4hkIoK
ooqBBnnlY7iIQz4UDBq7fSDZaJnPO9HtXXsR8NtwjjaXRHMMt5//vdeqMvOINGX0
gQMfyVVd2j7iGJw7qSgpIvadXRrfs/OPQ00GBJBMrjxGGnWMe7lJhrOqtKEfgsGo
P7mDXu+AWMNzt8+RwmTWBKA7JnqyPf9+iM/Hf+oCHc5HJhNoUNCP0O4yUDz4NkPY
JkwrBh3Dr+BNqr5Jfg6/ob3Pasf1B6K8VIqss6Y6E+/uWzQjw9dYc/tvL8vZhW0n
lQRl6sn4oEP+ix/wJjlTlt0CEEfvUe10k5tQv6zLbD9ku3FGiefS5w8ouKUhIuy8
60Xkfcn8rFZ4oyqgVtJi7j69yh5QirisYjB/L95a98LXJ3+dYapGjI9JYcc7Jvzc
hTHxyJwNPxC7vC8hjdXb15xxk017omB9EHF1gmhgZzjU7b1RPDv7/1fxCcWx+WeD
rwoqyt1sWmV9xzaRjUvhLoyym/TynWZhIsbzi/XBil/tTnoGjpNtVQCVQBeUgCo3
DlwhcgfcFFD1RkhUVJG4DlrNBWGA9IkYUTyhVwxRe11hpESxAZaU7KrDMHcKDbEA
S1BFQJeDp8W9ewa+xu2l56dQnL+dAQsnG2y5bMQMwL1wkcfStE+nldmjwa+qctAT
jQBiaW5AzW76AN1a3E/sEvbg/Ezx7+4Yw9BG8oRMdoE6JXHajwy/JJo/tG4dU0rp
RfzgOLll6iTFGDiLlvir3y8UDzRUtV6dARRZCG3oI+92pbUIyR6qxATR8fQP9HaU
tMQ/nKtVEa3yHccz74bsnXdJMjZCVitYZ+g8BCBdJOXroydQgly69w0M2pYd6noE
DcMQjrbJ0RGLPV0QpXqAfttHhhQWeVT0jL3wdfaNp8VrSoznPOyxxN3S492n/LNC
522h9wVER8lMxyiwhMDADY4t3BV/45cuGnAH0qijy4eWNFMINbT8VYwzuzrf4D0h
KD++/6dDTMaMy2fHRXsz8h5r2+161EEuW381sRMG+ayhaTrRhPEXVREszlI825eM
mHQW+wZXZZUdANkotWmN5MyszAajMcXzbf6c91QOOOpinngwAnoo8MXc8gH/mZsV
KqnJGlO6tZHdl4pC3rQkOms76u4cN1hBwnU1LjSIRCpv01PIiY68v/vzDX+/x/e6
5cApEnk08FJ8J1vFcvMibyAEbQlHpuDYYNr7RRD48BDM92ooSnHD0OzGti//l1Nl
siWneCR/8iZFkgBHYj1yDcMeBgah9d+5QmT8jml06o5ZxQf+GG04JDv8Eq0lztoT
hbd/tObVBoV6lkHl9+hpQLmvVdWzRUli6e79cgEtzmkcGJ28bs0Ao6psnXlQnJ7a
R+SgvBrciy7yqAZ5BR2LTBh6/NJHTypfpi30siqbC4dAuw1BwR6hIKx87MQt0AzS
4P+Cr5yNeEXj1TS1HNNqluHR3Cc8/6dCPw82adSiCACr4SLK3v16ona2ECsFg0SU
0zgHHAjJXfX/3RWpgFD6mUYGker8dZdTNqfJzqm/a5WLNVuHOq4lFNZK88rOu/i2
frGqA6UnQ/Y5WkXtvGmM3kVY+UDVMi5eqHMaNFbDGgxkSoC4JSVV/pLqzLO7tdVj
PsEFrNiJ8Qdlui0lZkHv92C4R8Dbk+r00evH4PMx8kPrG5TV0IQrVb7OQzeJu1rb
xG9Vk8GyDviT0cYeTJCwwrnhmMdzbQZSq8fNS32ffC5i+2pwOH38kx3ddNneQX6G
LR+f0WgmdWARn1j+VxDKDLTRO8Eqy4w1jGxy/G79HO2WWjKL2P7rmPs/QIovdEpf
8GYi5tXy1Uzg8B9YzD4llydJaGZMoVAiH3Sw5DisI05frTQVYviUaJjBiZ0CGO5R
lj3NnaePvP0JWWL4a8dv0ri752GxhjeivPZT4lSlDN/ElS/AZy2b0QvopYmgh+Aq
xRMvwWaDtX45hexOFjIfAN26AlxAE6DllPN5oEN7q3JFq82hpT3AtMnLmenKJUkV
9mYMDwOAVB340+OKm8q9AUVcayr1YYvQYoVlmas3a2zN9CRynsawpPZ6U1GW5NVx
FCICNXDR08oJWa+yeaxqAoMXyNQ9KyJTy9srYYKVI+FmzkzCuK0XigvJ/gaEQDI5
zmfCUDi/itJ/uDcF65Rt58E+8flJm2Y84AzzWg8x3ree+lGVjsNDPQghCNH+9jXe
fe8BGgxTTrh9lFlwyoVdMfx5NvlvH8LEODVl9BquiXi49vSAViWHoH8e+eW7GN1S
ffobFpHuvpHQ47JeVtxo4lYhH00MntBtSBuRd/pWwBNSbGBf0HHFFK5keeKZDlNH
rYrkaCax8J0GUNMkYKakFg26WnCmji3IX1sjqYG9mp/z1yAOjkkS5ymvOR5vkz1j
01PbjCavBnOat8IgOX+Kx7UKKUAeEE6UtmNFtY1i/ix/rB2EfaTsqy9c9mB9Nc/H
WMHSDnPPt891W2PVPEEretGanVVSEx8wXvbVgUJrxOK14zvw75Vic5qe4DnYiA6y
2TAq1PloV77jd6pl54xj2bv5hhWs60g3B1oax4UbV6+/p7GzO9K6iS7ZvsvrKrng
Ei8q0OLsA1Go6yirLkfJoEWpSvgCrobqb56Bu371ZP1zRQTJfLEcV3rW3S6hRErI
r+r8dfsBqWPrElRMfxVadc718FVkom/E16O7MxGAZSFIMzlxFVAtfatFPAQ5jnVt
2h++I3T8wEe9UNfbXDSrr7quDVZHTcp4B+eDR4X37TSWcydYIUYisuXTVPNHTeLJ
mWRc/Ad+dYneCeFOJXGDt7DZ695lj9wZoPS5CdL7QfEKFM+15wP19GiMg/3Ezsut
xqptrmFA+ZpKH+xPZLI2IuwUpMWO3cnu154ORjiPC2YCYhCcMKDRwoIqP26A1X3G
H+a4tSCQGKuOCTWONpbwgxjVC2pRB6J0193lXNasI/c5euwjTGyhrhmPxBOrx1eg
A2XLKfWpeo5FCxovt43RUaTKG1xrvTiUH52vUZtO0337maKbSk83v5exp8ocQe24
qdOc52WHA2M9OAycLh1/+BswJW8bM5aKiMLTN1OoIB938LA3fCqtKrRlSN264zeg
gB8DSNUrAEGDOIRBXC5uHGuv1atnNVhLI8XLkoJ0o34gK9POim40jLXQo2LcLxKU
kGdSHpnmqxKW7p6Xli5tZedAo+Sf46CAkspktrlLIv0AeXL2jtQf3oXduehKBZpR
goVMbWx4oXRwK1INkfG60zFTceFXiWXGT2UaNVfj5q9WU+5dDNpzNYO4Rf81qPxb
XhQu8nvpKD48dWIVazy2IqeusP8aNwzBEMcQSqSWbltHW1vWABpP8+DQzLkfoF59
dr7ISLKhViLvc155RzfHgUxQUS07Z3Ab3QvlnwtnXrpvsRfnVWiXOtaDYtAjCR0h
Yr9KHIhb0TwDcWRVEWyzc/JDRqFRDSxnaWfFsRSitfyPLVnPUf+iQjSk5N40HWem
VGHAvt7+0nQveNzZ0V8nmJTvJrygoQKkDEfUEZraQ4+XohzwhYE/XL37MonJOe4v
7XJGmQvZuzO6XKXkWkiUuyV6iMayw7muRZx93UO9qNqrKR8oTVVNfM9S+PvSWROo
FIo3wsCDYEHnkjI8LhMvjlwNrucNpvjcr66ijw3pWNyWuSQGQmMhL1/4a+C/yBdm
DBRRUZcnS1Mk2B37R6uzoRZH8vYTT1PxEMSUr/qA1H10v/+kxVczxfB8pBwD1x/L
FlrpTAYJCqiEEK4xr0EHn0pR7vA4YW3rnRLrxVfTgg7MjO5TSMc99atTF1jJZE3+
r5XxacLkk+l/axsZqyyYYXgSKz7EIaiTVgfcOvStP8lVbOL5wj3ld/vZpdZ291ay
pQRoBEk8w+bB2XM34dCxrIihm2zURgG9xeuMyUoB626MzDcv8iH942Td2OuG1WBU
l2OK0GpLioaWfGe3aIeY/0AImx8fYkprboX5y69Oqnq7toERTozskAV/OFosL0KJ
uRnkOccQ3mvT7CEGmV3U6kh0dbXgm9gLRVUj6/dyWg/eeFDNeyKho9gEgtHiknHd
PBAPtwGtiecNopIwRf7dH70+IlFlxSkdHK3owNzHbx3CTzIxUcyN6NP1iX0lu+xS
s3AHOyzvd2CmGEgraLOEqVcj4kLvYlEVh1v+Gu1C7tp1kZfR4NiYngdeEbsNVZay
eses5Vn1pXqIdPEVUswBYTr4oOWt8TJmhyd1/Yte08cxqd2u8KszI/S/Vpn17W+D
Uc27yOXOmUgqPeG6zqItl+Eajc8cWqM8GjXD6va1pA9S2I94UEYLrb0hpFL2LfYi
n3Axs8+f3QtchH7dJnIPBzjfEaJbyh/GbOkGc9O493SCZpBrpK6dA9x7D55dWUN4
y2dbD1y1mYClmgWC9jdJT+QHuNWKtI5bZ7wU9fmvzDBjfUtR3I1F60Qva32NkeMt
cTtSdTzKMH7H1+tuCaRZYn3+OLyMPycGu3468GrAhl2hd7EwNS7U1kZ5SgnIXPjo
y9qYT61IDldv4D5MXpiwzFF6Ca2t1c6la258lbf7XRpCWbpy0uRuyR7NcJF+1cvR
P5PqcK0GTQdHM6E38xUrTgAGVmbc7nnhQa/MvIu02nuEzYd4zF6t1qk6aEU2j2t4
cFT1Zpn8VWBE4w9IfLmWdHDPCMlSePnxLLUMcb3w1ERpZ8FAw6YZP2gIfLpOOfjV
f2v8mBxJyAToFWWCXw2ehb9hjfEBpmzJ/f7p0wQ5zhq+195K8e+2T+8t4JvC96S2
bTXShoYgyuiU9Est5ge6c1xpIFm7ek7OjjI19dccbvi8+lxjhDQ5lLeBFmdAVhjB
9n3BLxtOvMoUsQPYbTOBEcOSwe3N+1gv/RebzChnIc2xZN5GscCCOMvMw7d2E5R7
dRBxia3nsRK+zgnLko9pZdmw5GC38I3nc7+OZwlM2BmVY7nNli/zSnRhwzqkZ2FC
VvrIoM9VI+o+G/G/oeZrW9is53x1pwaEk41639Jn3dOhhUnPfOw9tBsqbXVs8oNM
zYDqUZqYfnGZ0aXId8SngwzW7CIjiObOLrbSGVXfBKpQ1jV70UnPcl/qfQFxA9oq
EaXKrFThGv2HHCgkMwbOirMQO1DsAmb5ka6tv41mTvrZ0a6reFbwoQ/OHwflS64m
sc5El+NHDzydLhVz5/7GiSOzS1WDSsa/na2+ut+0KJp5nYYi2jKbAHjiKfN8nQ3b
L83i41V1yWcUVOfwSYmHUqZogfJA/1r1nFAeHUjm2rVKcPNoVJQgeqiIihhlmeLz
0taUr/lOtNB8G8J5VZlU50jzcLW1eh1j5kUQwyZQDMRZIUvoaGfS55kbXg+4QPSI
gzry7BoW5xutBVcTiz+xNrFnv44HuM2LU6jiyfU/sFwcToOow3QstGPhVwHTRayi
s4jI/m0vmpHeivnp8VlurpEJaDsG8aZfG9yMQrKZHTOjcrZqIArydqlpN5HSL0CK
+VUyBFYB15WUznh5FTnUSnxWEwWJ9B1Sk1X7fFBSTkics33/TX9pqEd9fCPnkm1x
RHtqQEk7fRFGvVqrFAzZ0t+qykyI2HJ09OCACMJnQSAFG0NozI4aAH0JpzalOsSw
bdNYMgjCPWZT54bEfKi3FFt+OIAHJ9SLJwdU2e9CsMg0BsMf6HXT8ZCFsgYbX169
fjRl9QTIkY3shsjgLXFKv576vb8KvNDOTq1xXITxZx35ud+mbFaPqZVJD1rBi04I
RtV1jkgPxySCGSteSbRoileWtXiwKV4MoQKiQtaxQkvRbUxxyv8Nzbv2djpenVwc
0NbpDWRUuiDZ48PgQJsgDwXk6bYsk6JgZHJnOIzR/hlcDIiCT6odJwVyTTAcUS5n
3zy+gezGQ4I+m49JY1KmuKrwF4f3TqcGtmS+YtoBpIYVstMhfVTPWnuneEsTiPw9
cKKWL9XEjglQGC9FUStyRB1LDc377+tjN4x8oGI43L9KL6c7wcobM2YjTwggkpHb
5nL1Zo1x0MW+EKJH4cRlW8PkeBTJ4Sd+IU966kxJB81AWFqmqI8fVDWffXkGCurr
kl9I3mHKYtSwZuGrqdC+sHpHZdBTtDvHWovnXLiEzoVTAfnwFzPK/9c8avqgXV+s
FzPd5zW+zP3+TAryfV/7h+ir0RWVUMFlt967Y1Z2wvA10nVpK+rLGYH2Ye6GOwLR
mucKs1/egG92QPEEEY/Jac92wo7IsvfKKkV4+Y6+RZoR7qHjn+5Q50CM+iXlCUgK
yR7K4ayTiY+N/H6MrZ7I0fstqjnsr20ecSGCQhcs+36qLKf8Xt5AcoOHV/+uYHXS
fBKmFQ2Ikph0xPQWaGJllF65ARag3ucLeTiOa8ff/OBky7VPLAp9Tf/pSZPl/MN0
Hq/gJeI1+2JDCRPFYPkgGnXdKJ1AV1q8KVAsgjXbeUA7ilOsLodMzh4JhIib5igK
9Ygzi7Qj9S7CWXuqO+7fhm0lRPDzr+WJKilrpqY9iy9qOvRR4AeBFL1y3Ex1xf4h
6w/uUzmGXHyrINGABYvz6G48LrsGA5PKWCF2V/fBVM3q+j/MtBtgUjCZrPpsnI6E
C0oYY19ecR8+dI3SmYXmuBwyUEkXBNSNbicNt9BFug6qGyvewKD8+dBjqQcGxV5O
R/O2sf6/k4D2vlNwkzzXjhZua2d6IvWuFfuhVwqIQYf8f2keQ0o0CG8yPr6O5/G/
eJe0DVfMDZl6t8ZXdwBokKUBWzqZzbDyVt5TrK6uG05LbPRJzXW6sOjq4DHfDv14
uGLX3OQB6x/clrjdRjQgy7QsT7t4HGlU5iCq3nJE/oRB4nvz4boXX4YtB3OFUfIg
Mh1MY4HPvpqXperpJZOOn8tmlxrbeC+pF2MOEeZ0iRDZfVTgTCoiwGqL0wsCvHY9
fYdhxPVSnNhMSFAdC5YpiXkSInLWDNALkb43G7JFRUY0ARFi/6Y65ICt2wJwhFKw
uoffjWYXU01oJ1lWknLyWdisj7VxE9yrmyu0ENfTz1WAl4//KaJUJuKVk7RHWQLl
mIADne7yk4XOBNQoOA3dl4izAm5XptLcRgE9Z/9lcztf+SPwPVMu2NLRyhehd8Zf
D95KDeBVWh+z1iE3WOK6UQd/rzgAekrVB0tuvHh6abxnr3ckH+D4mS+r9adNMJ8h
vU0WLkDQIaLbHPjFiLCAa6Ulhc0TCevBElWar8kITcx7EcW/h2CTWgJF3nshueJS
O2fVIwC0FJyQyHy/M1czs0unaUCBKJvO70XNYpra8HZNoueDB84of4fXPBu7lGqN
KXQzm68rKevL2c5OEmb7hfH1JNXYFW3FjvYbyi6VE6CWMVv4foFcqsbjX3wYaaB3
pBek/ajZXAUl6bDRK18UxjLelLYQhR75FKGbl27O5nZG6mvR/Z2/pGDqLuievI6F
yyGTOLvkt95+mnWPUISWQ0QuphlUDE2MkaqGlpGpKsA9LRx9VBIwk4o4jj2p2lqH
bJQNLx0yhGKzh6xurd2QzHavKmvy45YVG/fH694Vbi0o9BdwJnv61foRkuc3YHqj
skkrgzOnJ0sWhMTkBK8wXwv3tswffruWxDpPGgjUArSlST5SWmpJ00pv2IC7WArx
OiFX3+xJym5+TLDXyLNE6uxj9nFMFqbn6KfLCezs+MZ2h4laEVVGindtIJkFUda9
YRlf9kAKzEH0PD/yeOnokzP52HqKePtZJ+1lcewIRFE6hbBlZVP3fmMy4RyB1JPN
nDXdqI8FNjg9fmAFWKNlyF5Mtv0se/oO/wTkc+CluZ+ya3DanAXFXzCm6Snt7vO/
hMOCzTa5IRxUn+OV4ZS/q6qu/Q8lKJGwWjgK6CbQxcqpz4MZeFTSxSBjB2rX/Q6E
vefIC89XxKf94vhshEd+nNeJT2VpbFyjNHNqLICy9W8/9BwIS+mq+dmUeyVKDpk4
x2A4nYvgOFM08K27u+BPQ4WFGJfydFdLrvS34gSEdbt/rNHzSMBR79Ajkl5+XSxH
N//uH29SVy1YP1dGoYsiybHJcYmS5RSVmWBxhDJUeaVbFffhVjIL/S11QCbsiPVA
VpGLG1ZbvqRNfpdPtGkIlTXoqXEDXwI9yKesUVWj3/nZOIcRyGIif/+2Qlrx43Ol
8dWAvml+fjleyAClQns2VBLZA4GVnPjEvUjTH/b6yniVHZXqz4XZ67AZR8tnyjuI
mQvO0lk7wzskqh5j7dwt1UgxkGvo1j5aS9y6NUU6/GycSOD366TjjGTHtOOHIYUR
IWM/W50VgurRVsSKWxmZXPz7vuUxDza720o3zYDXrjxKK6HqD3Bz6rIWdIiN8uXR
y5JA1N67gBH6wIcort+n9fN3c1plqNBHoEbdLMM7/oIuI5oSIlSKU1YAaQYgp5+l
VHxhwdYS9CZyQfLZ/XM9sSbyG8B3Db6HoMC2Ef4uK2niPyxEr2MVIF5ckqEeswvk
AmUirK1eHESUe6hXDe9USunvGtH0tpbWJZEjxf9e3zGLlnR7UfOoA1NUSEaKXOCr
YnD7y/CtJEpzNYtmViK1fV5R4o50iRRenO9zOJb9XyauN8IoiphBGnbtTPg43/w1
4BG7FHfqU1lNk5t57DFuH15WFusAd8GZ5S9Disw4Aok6ns9sIFQzKP3So7O2GDeP
qei/n1Ykj9P+Ka/mbOrsI0mpUgjlh26KQaavXcDHRCBLuiNPejWSKRonTvD6+uxx
V+0eOIgH2cwjN588FmNILdco9yxv7sx3xZZHueRdNrGX/BL0Gq2SW/B9N+lDTPkx
fNOxJ3lRivpFUIY8SBPVvXUryvxfHemNocuRf7jucRiDOnEUb7IVz9RkH6fFGC/a
09PAkkMgPi3zkdkcKw5Cq4DjcOMn1Es7DabIGdHJ+35xxoVaiTUU7TVWMk1N1M9U
990fnMYDsQhrhMn25f8gEbzp3/TlCOvWHO5t0eyxqrRHIlIp7A8c6YEXFc1UrgQH
eRSdAaikP4xlb8/DKGm94kkAPT6GoEGo9MQ2Is0TEFOlxDv4xaz7qVkmXzdM2pKB
1Tgomh8KQQYb7A51Yo3xNTJGaG3jPq5UIQFfAVZKspqYUkHJ14o+VLKbz4e4nmZK
cKD6E26VKIie11cqPXrLb3EygwdfHMscM3Ew4/SK0Ym9+pEsf7Rk4KUhWzE9yHC1
qScIjks0d2AcBsHgw/nKMlymlzYBl2CXM53mZNxUeKw6DVWL61O+yd3+y6E1+hvB
7eJ4Mz6YcpMNB8CIU35l3N9GsA+r7XNTSeAfvFDYCVoCUpkYAzuCJKvmgYpjylP+
Pv/rZyQTCLEW2Y1R+QCaruiPdMudY5bMvN5zctrlD5TdeqrUWRfhhRI00um3ZGJv
1ZHJlABoqxk5F92/FjilPWckx+qzkgYwQjZIG3L0XRB+FIoDNbN7qwvQJQFoC6S8
qDU1KIkZkjW+CJuy/qjuuTzD3SzBPtaGA5A2s0t0jAY0xN81oAqdn11jeJd7XAjn
23MqDpk1cLEPKcx439sKKaoCvC3nWpmyGnBOCcWJhBPhMnMlPfc4oG/RYVMpOPOy
vgfhUdsakGmN9ja59U3PDNJQhusnND9p3eI2N8L/G1/KOl2l40TqxF9+hHabciWh
9EJcCtjGABkTf0ZMv5+Y3CG2fIiVPRIFANnMnams8U4iLxIaci3YETn1emnpmFnr
l2AC5VMaeXhVc+jGoq8h+bSt1+ravtV6FIvT4cOaFwnPZhJNN//4u8QfbUGNSxOY
5VqAo44n0rEEQw4xaVdNVk59xxI8Gxzy2ah1aF5EiCR4QI3u+RwGxdhReJ3JBOIi
mx6lzoV0UOj+OTG1Yc3bF8cgI5s1XVPsb4e3sZSQtnfUpL9R+X1HdzA70SKAdsch
hvRO9ddkzHhZT9ac0eLA6Hd3zHpEl5HMnuQJ1X5aoKHGIsj29ZD/Z26IjSCFaGjp
h55MTaQH7HhgBxNJP5cj3AjaGuYlRcJtqd0Yk2DMUdrUlDZB1VKiuFE0KHNcxo1i
numypiSebdQUerLyqcJisC0VVarQwwNwVrsC5+lpF6h3HX9Y+rKj7mb4thv3t4A7
r4ryfAJ+9q9XHJCoxkHoD0y6WBFsj+DsnrZopV5hUFkKlnRmfZQfH1CXP5ZuOD57
UPLbcG+HkbQd35ltaPInWJ8SLwug8zoHeAbMKjkY+WSu6EEMEZYFv5cXF1NEf3ky
EMh3DUzoGqNbu6eeMt95cd8xL9NfGg+QgepQCiPPx75WuK1ljCfBJgQa/2wrazMm
BZln39rn/bTNZ52V3o6bUvvgbQka+t8OZLgZyOjR0MQJHPeOorVkqbbj/rmLTA3s
to3VJlxu2nbn59cTHXEXcK0qsT2AG16tByEIqSFc0ds7pRciClEnwjpxBkmIzVuW
89kJIuhiFOC3duHE7xWvHJybR0EoDWXDv5fGVDsBi9wfBC1VIxWdxYxn7SbzFdtu
XTvVlEjtYyzLLUxCG1QzRcTTV7KvyP9jDsAMPz43ZJJYfNtlM1OOPCPNr4IblFxy
ICJrC8VBYmMss7nUTmrCRjLsWpr5f49zBm+EAk0scvff63xKR7MBQsX+vUjr8lOQ
yvCb+mZ8Y13eaQGbq3j2OQZgpzAu55D+LTGOsOav7kG7GXDhsNBzhxCIUDZEUx9J
WVOBniKqmNaNiDZCQBFnjKMU488dDMyYE/HRQpxTPPgHmYfpMgcG4KU/G4AeDj2B
mwYbMxj3FuBv1Hx6X9Ogn6w7unoogDgqWE1fJFAmboieh71ccsu0G19m9+V2Jzaq
RME3MKCtjWrlvbiGwXFq/rOrSR3JaTpn2UEoorgeSjUI3hK4A/yUnHtVpAcS2x3U
ayWw1PINIAIVwl1H4EJV90Hk5KRWrMTWatKTKv0tJxJfmMJtMO3OIBOzIaUFnsvD
AIQsLVS8INAsEJvUWnEIktbtjZWVl5q/MV7kLXv9zFEV49vf8dGujoUgHh53cUc7
DpkTgDco1Nlqv0ClZ1rV85Yiw0PGuSgVSJqYfzYzEPpRai6ZxTRdKp5XpSfKqCZA
+GgXxWpsREidV7K05DYrCOpVKU9Lt0ud8p+041LweE/5hS3zc/KSEjIxikCu5yCV
plO+QDsKDzw01+VLKt30QElVbIVXEFH4fsuZ/1YZJVVSIZdtWB/PS/Hx8eT8zWil
YSwNOSTP8BmHQjaXNqR6qw1TWxhpV6uz2UVuGshY4tYnFCKXwPdGagjqxWZb/GIX
eTXQa2+gPNArnps2ZrhrCLlk6jZScCcCVSJQm0pENZ3Dx4bcL5zBJif9fG/eJXG6
E66S9JJ2YDCaNmeZg2ZXcxdjYjwGDXLQolua7LfHKUD2XzfsxenK0GAHFjjpHfhw
tM0wh/Zm4cqMoyKNIlRml4WK7CT/iqnZn0Yk64LzTiExW8OgimLUXzn6MzGK7Ztg
otTjFNw2PhxcAVL8xcK3n3VplplCdTEFBtEmeEwrvIi0gs0VX5kNiCXkCzWRVV3v
8+AJ4sQtf0fgknIyJpWfHNA+ypDjyp4B2DXHhvmn7IbmBWmRZGnAZ5ABnjevNLqc
I49s3sxzjsPPY+RLSeQEC0U6+NkKTuDjJytt+OujdhkLyGd6uCrE5Po3uIO1oycL
hY9THEcK/9BqjYAs3FknIN70GUUn4LizJ2eI5Q83JJvQfyuGxyqZH/NbU8K+qJ1X
AOGYzVe5qN3KSIZxLXb9BN52xjrV9AxFPIZgQwa/MiYq/C9U1s8jXFYfQhVGKGLx
Bww8bIBLtqQxPmK2OJr36MGxtbzug8KBywEc2F8E9SXKsTbCx09S+DW728DWiq79
H8eC2YZHP7eZDq6fsTHXE+Jn0KVDW2d4WB2A3SltFIKEqp7jf7vwIJxIXOCVybO9
L1cABuA5bk2c89DUZyq+2kitoF7hnGOXRdREfPZBw1wNQULMeISm41lk3t0t3YzR
NKquaIEjLamNQJs8SJ1k2+YCGlQUTqALmbvzpriTCZQPuoF4kf/4Xyiuknq3lWJO
ahuq8jlyfunIg07G10lS+hWMSOZlKbFmOkrQUTkZJfKXBy34UYLm6cvpUYtZPlFi
ojYDuWUCn0T41cMjK4ndqJ8HAJfzwccLTwnrxx1l4kVXryNDrsod87qDHwvUexZm
dXqH/x3bR4FOw09f8OYKqFmaOxFgWo+l+SeCe/aPYA9kFkYKipKfF8gN84JwB5fu
NkJm1udhhA/9RRcsZZkujL2mkzhdi+0QkqKPVan4XcMCqG3vFXy5tcLvRerAy/lu
BxUaE6M9nNt40zqv0ukDsTYG3eQ8xfxiUVwvL0jpRh5/ESOWRxiWX3n4+vXcfRKp
2521J4PbkcfJOY5vecnOonnFENo4qKX1btEMg5HJ7s4KuUhBl3Cnlb2yNptXzAGV
XvXNLq3GpdHwlwTS/0ZY8JoesIFuvlCTJ/k7GYGxeXfRYH5M3Gtjk0IKXPV4z/cd
CB8cueU8HuZj6x0T70DQYtVSaMRadpcQr1ihnBk+ASBf5t5RxSBf53Fu1LlitrBz
OJyqJMKapRbMQdxLnTTztvURqjWioOHlT6p6e7J45LvI3+qhqjzKCX4LEpX0gjyZ
PpL1J3aZbZQ3ADS3wH4L8tTg3lWNaSu29zu5gEBKgnT+7OZ1Tx/CylyZ+mPjU9kC
aFYZUD2g20Nd6Z/E5qNvcb5mST/Twlmm/3+utaMqnMF1uIgjgxgPM4ZtjcHD9BVK
r89kgumgNxv8UNwtNsRBFLkBLXP8jy5LKjCb5Fkd/DDWTiIEkZo32FpzmgDx2nU7
UD7G9B2Is7JcI/Q80nHSgHzktr0Ob7dEXbJVv+xCp9IUZfmn1Km9Kj1yZzCbajRm
lkRHkoCXJwyDv7bIi1OtFBFDD0qpvQkxoP+cILD+rJ3vfSnwivtX/eRAWmit53G8
xe7z3FszMIBZdSoiIdgLFcFkx7A0IWL9/Pyt3oCvJNyKyZnuFnZXPTefMAGzg7SA
mizXJMuyuEJ5oXMDaKf9pE8MjYA/6K8z1rfwCyUCmoeZvGTEYDqJ+nmxkIBv61Ev
Sf2Ngkz6HvaKPXLkY1e9l2aCa+TeqtMYXmU6OcF9KJxmq8KIBbc/8BKSQHiqQDN1
fYKEXDZDj1473l0RpiiMKd7+5OA9a7OXhkC03htsGGnIjHcAno8i5h/vdGFiTc5l
iVcnkkEzkDFLdW5DVvf+mTsAhSic1yMFED/ewxkUZYDts8823x4jcuX8vh5PEXxT
eZypWL0ZR35dKVFMZnwGX1tOuFuP0qtzOPugi3rqVepr5SiUfo31bPPeaXWfL0AR
4RbvWFLfKiKwCQHkRWcznVBYglAguKSBCyUeI6qxhSQJRwJhW1+JL52KlFN/U7Pg
iWmWAWFZqrJooqf2VDwi41bOoWeuqS6BNCH8eet18Jhj1ZX1utAaoH/8aElgpDja
AgRF2YMLkL+zXsfngTB7CwNbc0L7v2arTPULMojjihqSZzqsLziCZ6hV1c3rjkO6
rIrs8xA+ixMuumSm1N3B8pykOINrkdL4wQUVrrpr5hfUohAye/onPO1ZDYmh3X/j
a2PNFNBHlSGnk2HovzBGGeGyDs4BfczCpD5SehVy8zYxUiVoGegkCLpEHVcTq0/N
idgGwB9IIjnBbpd450uOEAJXsz8bJubDhgTye6i49ckdRf8rYzpCT3u6J4ZZReVp
BHkJbL3jS0YgpDd/VQoY+3a3uV0tDlQntlbccnwZ+VCNsbpwAeI7QeWnNbicM12C
gXvIlG/ABMUausmHImPuLKWMuQ2HfQZYZq08TAwd4yL82ZbtA2gfdB1DtRwHz6iY
CXnxtBW8UvcOeSfQDx3VoVv932UPitMJgnLNQ6acYVVANDRhPVRbDgDY+P0IkncG
E8mSLfn1mcc+yvYmraV/oTuUy23koMSE+OLNs44TbcjcO1xQEBQILOV9nPjqjAgm
VkLaE1UUi8AItr7i+mJDoZRreCZhzv30bFO07vi9iXe758iIe+ui2pvM0cBaEQwp
75XKD4Wwgj2k2PnNY5bz3mzLkAVkJcs/bhyR3opYowOg1JzyZbO1NdA1FBRoXGKQ
IfBMY3fG9JAeWctJD5+dpNhxthyKGVupU1Hal6WjhTgNK31TbUhqIJkadf6mptiB
xV9EOSeJCYLD/aHXBcUMFma20RwgBNYSQtC9MbUBKe0tYHCTLYaKzTLgpV/bTIgB
DMOgtc5w5qwZ1udKYSE1B+4R4+6+O5BlVlMAbaw5J4ORqWEtVakylc138ng/iF0V
MGtGGM0U8XgUBfVWh4tKow7eFolY9y0HMcgpBrjAK0fPSRXdSZN+WGBiXVgswI6r
kVfazGMYpqjBVfAt4tiVKULebnmOpFW9kuPPaXIQckhmMCcugy9iANV88IYDdITk
Z/dT5fKH1liV7RRRkKKPuWkum25zwMa47bZcVwOGt9Mb6xUsrQ7aYziyqeGcbY2+
grmfT1l8FPsaKVCeHcMkHoOmV/6y0ptSHCTUjODkcFQbmQH3hVcZUqhmUN5iGz2D
1VuNgqSU87WnE1hPARnR3fBMrprWDKfW7iaj+S/g8fTFs21xNh+CE+pB9o4e3Kq2
UCSyv/EsFF6APc0Cq0u++RWw1BfZlsIH1YT399XEawBL/WgHJCa4FAYu2vHKFlRA
hXpOBVOnItpeZxF0YxRDdxMtw0KEPcfF1EaVmEy5+GsZKqfbYHTZdlPd4RMlv8eE
/tYwfp5n5A43ELPcj77eNI7QNaXhKbrnRQUq0PDe3XtShevAEW6/J6drj7lh8DsS
K7TNkA5EUx7dMRoj1d1HYrwyJahIzuvsTPCWMFTBgauTp+yb+C0du6LoxeDXgjGy
sQ82UtIVBFcQS3uoc6Cdut2ZIGdc0RIMgD+3ow9o2motbooikCLHtaPT0tKxA6UO
FpkOP3OIWDcdrxtZOiEyrQrmm6hGDhM+YJL6B3xsKsf0mQ9NDt95ARvxkZTgSOHR
bpzVWHnPLO+NSytWTzi82VRKTS2l1pxsM/3ppYvVejEMaSjiOxAm6HqFP0xGKxKF
UY8ahG/0BY9h8s7W+p3kO248Mu1xB3i2HnULXHO53jFdez9QTrWfwhKRWcRZMFVN
hnFtmnGlNy9EMOEh6jLbMouXFdvXz+fKBL9ydv+7NIBTGQOkkFThawt7ER+lbmmk
AAfwiLw/ycLQJxc6aft4m4cIXW/Ev8oWn2T0yRG1ww6lYsP+6TkpK1fAN8KKeA2f
myH5epLP0u/R37CPPIDCWcby5SsLN6Wb2mzgqlPRemLfX4PwHM0wgGI1M9BSp3u8
wmf/3ix09XjeNaY/s1EBCMrQHp9CqHQn448DevAsoITd+jyoopxAeHXWGIJJ/lxK
yYi0lAV5bLdd64nrWaTJfmNcU+U6CM6aBFW6UfJTrTIU3Vo/IqHrDfI3VdAskg9F
5+xF9o1+d8wKUUqLTi4eFqsvgUUetex5sgIGrk92yPvcIt82lYfgNKttBiWVHhoZ
h/FNiKcTzUrc8PHJYK+GxXnurqbFNPYl4EjTvmWQWrG4utfQSjmoGtwsqw4Mm6D9
KaJnKU6lXpsraD2SEnYSCLEvt4sUP8Onyx9oq6rAAjRfmovxw0PX0wx8TXL1Aa+l
U+431tubDLMAAXYCjBJ8nSLRGe2bwBCPg4mp/xFFoC1xKqJd5vXMNYVK3xm9jiak
RzfpY5qiTcFtOX/o8lo7EPHUOmQOy5En67Xi6dHPu2OwiikgC17bQdF8xFU1IUKP
6sN93KM4lYOozrnLioRlbwWwmK+q8OkZMYj6fMchpRmxherMASkrqa4ASppATTbB
SHHl4Oi/SPcjgzGbrkgBYc8TQHMKN/Seu812Y5jQjYTPLTpneALHFCKttePb0Qsg
FT/UqfeAZjLfhdpE+MNNfCv4jNES9XOgBuS5crAs6m11t203AkE6VSZYiNAYQRPo
Z2E534eaBI2gHD3sxfVuVhhSV73Y9IcfEOp56IQGKEm1FPC547I+g/PJicfpNGsN
/q6oJA9gJAJ9y/yhMhUvO4IneYLrVQhkXuLPNBNX4UL4XfxhUSd5zvndjSgnplx6
+aV3y6/knPh5WrUVJZehDJGIVdNg0lc3gNnnPHluEh3PZoPwqRD7HqzAB/t0q+Gu
flk7tqWu+6aKkj9hv2oKPz2b483sfGpWI49oB+rh0SjDiJUC/vZ2+W+POf302G3q
iLfDWwpfPrLoODyTFSSLJgi/W3q/b55WgeMfNSLnCp5vGqyLOqFZxbpB5PXHSOu/
Fcu83s1lJYJF1NI+YOnbbtzOoYS+Bo4XriTKEXcbfTxEKjkpmn86ByWshlUoI+8F
Tc5cLH2wNh6sVBIG+/RlGrYpghMVh4e5PbS6EuIVc4pR4jCKwDGz5aVepRUiGG4J
Qa9BHDqHtMrOkV5VXgJEpXF0soa8JXnKmvAKXQs/mr1y7OQtMGySAkcFs85eUrrL
Ns2Vq9VAQYWO7lcTBYvYInzMQKF1NN3+mmEpJX9zChAYapeB1D8IK0ThDTphhf4w
WR3pwY8odPCDStbzwNcJC0EbRAbgZeV9WrqGya0YkJYqCE+ZJDl1H5l2HlD/mFpc
J6A3bOVZ7kBmE9DCkddEenJNZm5lU8jHcHtsYoR3xbwFJz2C9dPDxjXGfmX6LcE5
O06zLJzaaFQZmJ9YrcpZb8dB4OnoPhFR4rGRfwFnaTakdKXqrwb+Q9fVqsbT7YOU
5UNS2myStPhtPMQs0jmYHd/jouiv68PxzzoYEqBB4wOEf0jYwjTQABRQQI3vQzZO
IH7mAXyUXbinjoJ+kGaY+c45TgCNH8DnSCc31MB+6bvvPeJi9hN9zWhzkyjE1E/z
VnASphAdx6YNOno8mOqzVHNer9t2LTQVgcQYSCaSl1DU0uBBXYWoDFQedOkPTT3B
usMPVHYcIiDsb0aGylybN/6yMJfJaA2tQTswnRIAsNxYgMCMi3AfEQ1a0ueZE/PJ
C3+yDUn9FBZpXBFeKbjY9E3P/HtYfJYpcs5wvFeP5jyv8K2YPldpbiIb3EfCJZiF
SZX1istrklH+JX5neMCdjl+0TA51m9vGnbPpXJ1jmq4IMpbAds/37XVUqQTgCNVG
n+T/d2eL9MEsAqnPBg8wIcWtY2k/k4aio/nZOw8ZPLuzVpPGaqziMIHorNIe5scl
6+tZQJ0/+FsdQBWkv8GDwDuu+1WtlnBSXTxJFSuQoD4bFFIYPcUhIixUwILwbgaV
NCNjMAukK2HPPPTDEP1CY8s3QpMy91T2k1cBl6+J5aTi/ySB4qMXinCLJYVftAiZ
7ZqMJIDPm04vxM2ZW3WxhR3sCRoD0VmXVB9rO5wwmewv9YGRtRIkIPa0gl84ENbk
9gh3dcXVShouQsIASCrQArZtpFjxurhSMGH4WkJsaX5EiAvWuXLx/rBBWUW3/TYB
iK/WwPa1DCqHeMlhcbeZryj4PT28EGHzjv26AzrWrYz9nsUstY/O9mgcZxtM2iza
iIJiH+8J2FUwRFxIEPU5RkNrhJN5E17Ct/6AMU3pBgGQyB8hhPfAY47JB9o8xKn/
o8oBPfWWEQqMJF3LORYro8Y3hL7A94sN+FAvsEqzux1fmCAQaX+LAQDI/hZM5rhr
NCTeS393hUY7dsrEnA1maIcBquVpAgJd7RZcpHsGWPv4+9GCj8cMIJ40D0KpNcZD
UgTSHJVv6EJTboJSJPoV0tFnUVBKpwQNxIL1K6Grl+4C0okJ2Gos3+HHf3aL2G3E
wGAOv6sn8sWIZ3SnSP9X7uj5SbMXdiph1UyqbEwz47op+hAQNVRQlCK9XkLB4FeW
W6wyp62TVtTnRI9s0jVvA5n0TcpoVnlu9b6Rd5bbHcwL7o082JPjny1k9mSPrhir
zB7hwHi/yvPWlUQk952ogQCdytTT1ao934nI3kJqFDwAS1I3u0zOrnEUNRWe4iIa
f7yrkOdXts5jjLb11zY38kiz9OjjgyM/gC5EV7zv5JKEYzqMKE17mToagJw73Pu0
iM5Tnqbm0Dmxi7O8XhBnEXrSqN+d33y+dQfaDC0Pelty7yWI+LemPt1HG9bTtuO/
XPMxVGO+OMPJlyJ55EGYZIZf/BWksz7Zcg0hPOfyTcK5ywgZvogHZbxHG1Ffzt56
uLxysq7/MhmYqVc13VTsLIFSu0zbh+dqhnYwTgV2PMO0taZPLeLNPJyWolM2Y5S9
sol6sRetiO42EEHIzpKY3pydODAj5tsaQtOahj0OMeFjgYs+UQ1kDIXTl+ktlA3e
iEcwjCFC3Qtzx0bed3X3j/i/H5DSKP3N/dlHQjpAOocRwzZDBS74mcQuMtETFmu4
g8umZifRIEtcX2k6d8RjD3VUAETu2f4CYSHD1mMZH3Qkq+dtmvGQ8DLoOTBZwq7Y
hJETO3rP+9REQLJPW2BJaW0CGWCsVZdQ+URSE2Pw8lK8wfaimKmfIMEcMq67S9qG
E5ut3K2W6vkwh3S1Uxphl4m55/8q4kHElcFT5h4G5S1MomBrIk8IndvvlSZo1Rdu
AIPUu59c+LTfoBZzgF4PpCmlASMjkZebYbGBXstngLbDJ6CSehwVtsBdOh8AAsTN
ZEnjr6BSdOgaI+KWCTpr/Z0wI/hCQDYGxPajc0cO/ZfozyQpLQzTOXyijiIObGLo
qQFTpNGksYOzPeAmowFdAWh5Xj7EMlSPQNPjN2OXWx5FUqJqhzK5Dg2VHJKxp992
fepe3HbdS85Uj2namDY5F/aBS7oxL2/9FrG2XpN8ZEkZTbxhpPdZD4ol/0HV/8Cv
JNDZqOlpApklrtHNxxlQ93i0xQQZfvZt4ap+oxrcAcwuHaZNhVz3ORWMlmNl7Jdi
1u+3OF8yeKMycqZnkxtLzjFLWirbf+7YXdIPbQGnYxPkn7b2xXJOlzgzrmfR8O5i
mKaWRGkeeYfqz2fGOgVh4G/JLJYjWc3qwyECYdMCHbigxeYqlDYA7LJH6VJ6/gcz
NOajeqdF19DXP2dmIImeR2xevOfzWMb4wlaI5qv2Z/sgyF3gnSLxoAm71a4DOEzb
7aXHouDTF/IlmoVhL1keb5q7d/udMDJUquXO4wKIET/8FZzHfSjmglGeIL4J7LXm
TZgvhvgUcwJD4MiUFQUvzlRaQMwW9w5r4mHwLuRhIniMy12PjyXMjDQ81xeR9upO
pDeNVLWe2XLSQSbJG2XeCsPVZXN8Czr5OGLZUfqP2/mVL5RR6ZGyogu60p0jwHS6
zxz88WUh+UusJWe7yJwMYUw27YU1Jtakj6EmaXGWGseIRV9wQ4uLC238KeRG+MH0
2ywPHVl6eFOfiuzWrbMzaQDjpwXGhh9pXJvsdLQTPFyql7aFvM+cawyNIuByOzDY
+Y6TcTuu/4yjuC3EJ4aWNbqJTJufTDMAOg/zrhLCF+tTzDQDYSdbWmEJ/27Gq2qv
omjp8zdPihrPEGgdUIT2D/jb4ttqBlJe33iLvsmkvOinx9mE+AClTuE9ij7+KzzB
dCw7WuAHjb7nUSUCp2c0IGT1Hxt/evn7zbytJfTVaFR+y/Zu2QuRPcENk9u6JLcv
Dudy793FrJ6OOd22HhbPK5t7f90V5iKdt5mDVj55ZedZkU0XAV9beScL/ZBDNqOF
VZKayGaWYCUvsipAaOxQoDVvjdcw/WZWWHgeAfRqaNf4jZZ6h+KB7RLUl4eE4x4q
xMJ9ZQsWgXSw/N0mmB9LbflEb/u8tN3dLPgu+Q7fnH10tQ7p5ZkdUSZhlRxZr3pc
+BswyI3WkcxKNWN54Rr/j1rgwcjxdZoQBa6a+I1xVzL+5WJ5fQh4u6uTs/zbj5bC
/neiCEXHPeUWFmPPTawwO0GVlzEy2jzU6F/m9FEgMGG9bpoNEqWEiGAizGv0/Ghe
hibcZkTk+XzVN9tb3au1lP2RO2v+eieZYkRBzjeFXsR1DD3yUBw+aOzHdMmynQA8
onf5yL4wN74acD4uCQp/H4gbyf1tL4PefDiMbKa9iF2xYWhGqdtY998QynId7Qma
FXdrXchgMuppQdFj0NO9qlETZ6mt+t3pkrbV0hPW8KB3qChdmDMIc2v81LVt07if
efuRnmaEo9znHgktDYf7oX9ECJuxjByJ649fuRqlZI/FklMOuiSLYJ+un1P/gqCf
CGmFfzDvhhw5yOKmhsuyuW/ceh1NKRZpgy/OaOHHZU6v3ds5/ER10eDYT+faAWKy
Uvgyd1QcJprq6P7OyThuyEKuVfgmJAh9ei81n2cxjP85nFwTVGTOXxweNuvmKcuJ
NuiFkWSdkhRxE4wZxulL96zu5RjLZp9ZdjBtQ2V78ZG1Y+3soltWFt5XGrnw51Vs
XbY1IzdzPmyo4niYoc3wiwINDPUOpsBsfTDUlNpL2Vb1b+J6x5nyaGdz0UHKyNNR
G0dhGDOQCbUVr8x/0UeHtt5zh3bqNcRYgq6RH3VpvC59c0SgoKo3SpRqXGm6J34Z
3c5fQeeh71BYsfSb7CwzhCKrtH/lwAAnsgOJNClVZQmbDZG7RDLMiG3B7N5kPt6x
AtUP+wma5tjLAaSl/EnuuZI9w6s9mbZvoLUZIi0Id/uEZxMZAI/ra0Tbo9/f7F+m
uivLazbl3tgoJPs5g/MSa1j6qF6Qo/tKS65z6Dyxg1IvsGRtEB3ySolDL2gpIJbC
nlTNz+leU0zuitccl5+Dke77byP6lv9LlrvH4KfdOjebaJlVh/s5LXIkm9S0VFoP
qys/TKT46+1JkdjxLrZGlbDYgFo4Pu86mXkPUSxkaOsZp6rPTNNC6vVLNnPzpj0J
Wb4cv3fOEuipFo3ZqTheA5ULy5Xle/5Xbn1MDqa/eaD/MIfVtyQrsMmm/ByHmztv
CNYYpgsQPXYTvn5E32YRjARjBxQ0wU3o0qL+l3aiStqbtKZx5PY0QPi986/sUaPy
lo8Isb9x6w2OaWe517XCsIpNpqdDbptr91FBDR3J1lT9or6kRQjtI9zQBk3LsWWt
f85MxTOgsIRcXw65YrjFJqM1mfB5faSODxD2vwSE/EKeo6rv8Sk+qcyep7cCEzbI
b7yPQVnijz1eHglK3nLf56q8Sno8dAPI63TpGptzWtEtHqgCNcqde0UP72ZeAe1y
1AB+wqJ1QaZ13cfGLYZ9Mnm5SRucFeAnezmvoJwe40GT+kgO/QhQwKePXfEHyfnN
vNGZYzbho5LRFhfAhp39Hh3yJzunEcjdsIrf6+yKQTsi/UFuWW5sjt0Syqs8LAvS
/kJNQO+2O1RUUkugeaHYE/wrKGjSELmsJS+5kQPJs2x2C8nqx3DXLhppPC4ynRCu
1PYzyfAfmc5dUHwmweYE2dkSY3DI0q5o0BZy6E8SSboB4dFTBgVSSW53K4FHGQLH
QYjicW0tuxAlM5EgMfXiZzCFa4VRuhTKxyPQJ6qxBOTyKdP3F5AZAujg1+Q5WUCc
U2btM8RlnOAHtK5s9FJiVi9xHXhgLPQ5pgPGOFtmXLjBNG1l8EMA0p16cVlxPu9d
0x+F9BdP1i5ov5VUA6RDzUYaJEqSFlgdoHR3kgoUkzzQK+Nzs9Pp1ikoKLPOU7ei
zIP9pQ09e1HN3Ig+VFAVFQTDZihCS0V2K4A34Zse34dmxhe2tmchKo8k+aukyFii
YIqcANfWkH5CVbAn2QQItj0WMZ80RjX8Ap9jNqM+zzqOlr1e9/rgyXeflv2t4KaE
tcA+6mNvcqqVOnbis9X4rc7bWjnJFaLyYWXXOT5qqkBVWlSuTY5iEtHiS3ZBPl6o
5rli/AtIY8Wz7+CV8/y6766NFQtCTK+usmFWZdd2X0ginugg76+STcLvIOuLKdKm
crmS4DSmU4Xj5RmZoTP4VVeS+iTAuHEva0ROwVoqWj0mg3xDwuR8miokxBOpM1Cn
XQvqqwyUiaJ3xamIuqb6kigrPmIKJfmchYIbekHnAAdT90JzuUQrjVCR1FLwNSRG
h6N+uQsG0RIuWUfodQhsvhVMWTMFcdCHZVTCLD60aY+tQLmBDXm+kOtyuJQ5/sQp
guVACfWMWKYdsZ1tdszplsSwgxyp+KgdQ7INTVCcICOj49p1zw2Z86zJCF7QOMxD
KrJZiw7G07NhrB9Bf7afjp+y5E0wQkjF0dwrcZ7vG+0sKUl/SzhffG0UJM9IZTtw
GM/xmE8eUtWrkLlf+qA+XvePz3fkM8gK2G+XCH0guuGFGqBAqsb8jo6zsDFZ16mR
4MRJXCVfCC4k+2VS/Cjmoum03aB9BntWhsEBQZIqK1qTMslMqKMhvcf0es8jAUIY
elpIstnD/oAGc/IBza7oMPCPWt0urJgcpayfCX7DlNWtEaTC4HeSo7wBltlKauoa
ViwL1TWQQRIZW9In+YsY7m6nqZTYMU3gC8s5SAV5PFYRZY7ByqTiDZnqGMMtECJ2
07MJDIy6PwDDz71HcOZA2xUSOMyRcdJ55c5T8HJOOB6slVZVpTatBHLBNAy6w60Y
5K+doXHxhRuoB7rZE7F2n36hSTR9rTGQyIvBBKopQ1xxgElAiCY0DitS729IxLY/
X/AFWh2jQMEg5nx1RGxbyfxnoqBG+zEPDXStsMXdZne2y0aAT8TgtZuzUCkJIRE4
2kOnx/icsOLXqdmtHLPu2V6WfsjTBVpHrSJSwCWEm8gg2I9q4fqL3eO2EjsApEKv
FcgfJT5EtKrGB96U/nANjCxO9JlUpg0PoNxAKn96AOaIXCMzDvs/DJeEaCGaOY7Q
sd0Gz9gtHAQkEu8972xdiGp4guWRc0PXSXhTMeI0LX++dye679CPphV1ev92DIPu
8Ixw9P1grb8WH9RtKOfR3yvWGTWzPbPcROPNX4KL7g0wQ08PHcY0eYCZ92EN0N0Z
a1x/o/H9QQyQMpkuQKb3FhMMo4sTkh7IShk6NV2CKuWV23A+HFngAgKI6+gNat38
/w7bbd3yyVHHKtKIn+soPwmPQMb11SMdS+6pIS5/lVXXRDjlLBoMSTPbFJam/8R1
UAMRv1+vgkyyiwou+jH6UcMPFiZ289Qhh9vdzD/W22rBIcFqeTrFZEuM4AukxHg5
fOygtIs+o/Sq/bM/PqNmQ1e9+2P/rcivbCU4ryf5G1ys8C/zo+ncOdahAMSiqSM8
5iU8gzBHBad4h+T7+wWXAok8wOii9qVMx6Z5BTjiS391OiZE68TAKNb2aB3EGep/
SdArjytO4YVyaN+wG585PLfJby6vbgz3AoehEzpa6bOf1BZd+c49P41C567Cx1EF
tOCl5khj+Jgv8JPtDgoBwSyxKkP540MxmXuJSaKL8+nJvYaCVUzpiODK4nJqrn4v
bFGGv6e9+v5wAR1xtuAst+ZW+RNwl62tMzdSRjsfAZbwL05pEs5fXOinjpx2fJPb
PLYotwzdcxpgAprZCGudGt/7kBnHzFp4I7wLMO/j4BtgGvFGWWEod8VXUQ96DapA
Lwurhw359xN0G7u0TrkzJn6yARWxWkF6BH1k0dHl597hlcYN15BK7cvSptEUg6Ek
19/LNy5LB4/LoaC191ndDegdJCTX3Ggt7DdtQyL/ZEYv94lpcFwP1M7G9MuGqIv1
XZGEOa3t5rs/61JbGsuToyxrt/IgxB0XmUORHLBvio22dAzTfsj+BCQK/ws4vM1W
GwKB/IuuybB99jh7XveCVVs6n6LlAYW99z19Gy8futzw5Yob7Cn8RX9PMML+X9bB
6P8fCYBMAdmRYdLq5kS/1S8Z5Jrzp+D05WTAzJcAf90hJtJSw/q7Qw7uEdJPAEZ0
uYde4l0CYTigPcNNTQacPe4ScNoFqNnFKG/k1SDMoaHNM+HpJG6auQAtDbfkkpxd
B4zSd5xkXtcyu3R3zclErk3ZDH7f6IQRYDMyCfjo8WLmpiWVEh3CccLhqt5869xw
L5G1wbHVkw1cE0L7MNjXEizTuvnR3pphKuqiOSnJmpP9Vt6Kr0fz6gmom5Hg4c0n
OkJ6DBbpblFP9+2OjjxNQlCpxAIbgAoac8hjHkT31d9sSzFoQ4cp0r0DQEtQTcjz
/G/1xAbw3lE8lM0a3ummyrueOZbWq74r93J0vkduL8ZdPqkb59XZXPDrjJbmfdyv
xFfvTQBASJiouQSazPjzPuTQsqRyH7kggXZHClnhx+uDJw4wMJQ++AgjU2AvLKpY
YhHz1qHJ+1brQLGuUAEmdegmJmjHBodaDbHtztBRGapxM2gnjM6ZLVNznb0VZJnR
3+/cvna3Y4olJMWG9wvmcJAEkzAxwf/Pstlkiq1JPJyt9JX8bOS9uu4RjT9jgzca
GZGqcHqfTojcDNfj15OaAcaddCcjUuVr3Frp54hXwW1B9ZT3INLlZvcVrlqAEhSK
VQ2eSSsh+gz3kMADpfChHN+SSffE+B8seGkJ1YjEtHUpQUxnbm1WVrYclLaAh7UM
2rDx8oTRZlMCsJeVm5G9IiQz0kY4tET1/1A7X6R4smp1WwRYOn3BJpiRjXDq3NAt
rtFgM9TDAPex5m9wk3jy9j14re9vwD0WPBTfxEV1PevNr9bjqSsfJ5YGAlGVhLBZ
77v7NwKaGL0oTCLep/6Ee3NYMWchNNVBM8C8CFvwXPm8WA0SYz0csRnYcREVoYlU
UF8/4VJml1lFF5wm1oL6tY+MhAsgg/fbb3ss++CogKAWAfOvHcL2GCQ5PCd+4PyC
3tVbCeqHvnVlizG+i7b5g8QzxXGyo+uEFtISpKrPSs0kZ6hgj7HDkQpF5RpDHJJo
0AiHVrAuNgd3TWvuFffZFzTgG0ST1ujFUUEwMam/cOzdfoP7OeDNAv4w5K17BrO7
ttieNa9NxBfbkKRiHdZ47Kjj6gveGUwVfK2WUvTPQzUhK6qpLNV8oLEiczsXsQKX
ifuYzOy8ZPrFA7M23IpXzykTQMwtQtKe6FzI+SBeDWfar0gMzwWq3mY0CBARvbkl
j4u3bPrw/ZClWVDUyXWorrcGdP/2PlV6n0PaNP0pNIPg8OPw3+Oz3A0+6fQmDmG5
13BWTsBY9kXrAIUo4/sUMZSSzw0B3vVrI1U/CmR9/yreklUBp+4fnVjaDuZ22hy0
3HTEUWhGTbrS5oZRtq/lYm4k/kGQPwcnQbKzECX6DXiH+vWDVHBs3Y4xSHfO4ik8
2r0eER8VV4x8ouea2/UW4J5XPg9tSA8iW+afLX7rAdnTYLWwvmMw3+6LmSxncSqg
gSollgjdG5nVsXAZ/lYaJ49j/EDJEwVMhlZdpNet4M6H00rMxsZvCgZRQfkNNS8N
WqyGFsSSLI6jwJWTgzHAxHzxMelt6tbHYTnrUIh2KnGGM8pmSgd6z8re7IgVVT82
iUySZTObLgrED2zOYpy+8r2CeZVZcvZ3G8E+/3brZrzNwKebnTPw3ipuGUaQXNWA
ZNwzOxgSItGkiMp64KXJg3bdZe1LQeLNwdpP6DsZaPvHoAp+g0UmvbVMi9AaVbly
bFpJvNokKy12zTcFpD/f8kJCJstJ3CLCQniK6OkS20AbY+xvO0P7PIelVSWIdRik
zRubIRz+pvvGayu556v7nM7jxO8zMbwf2/sVO5A17JqUfv52Pcz5ZBWIn4dIdWhI
raVHNTEu3vShwF0856ii0mKJNQNZPiqvGEFNJFQ2IzKxoVzmG35fRmObQuRCskaz
DNqWxQS3lDY8ng84U0KCB5L5IBT+3KCZbY24spPWCQ6ML+Ks1Su4cy1VPDX1kgg3
+0efwB42pOFLOlTiKIMpfCGITSzizMhYr/R1A+lMPj/+D8YwIKsMhBFwJkM5gYkP
wg1K5QcIVMQkuO3eMiDRE9LmVWlH8oW3lIGTPUhMq6WdJpvw3LKMHm11eMMdrKEo
e7B16b8P2brRU9rBo/KawoAhhWUO6niumm64kg6sBWZb90iL/tZecTiu9pLN3cfV
yrl4GMgnion3PHO/i6Ps785LRs29VYEUZTww72w1OHyWLpbu9cZYUv3/u5kkdh7a
EmUHGCuAm2YvgU/zzT0f/OQfyJosJmrXcK8MN6ucwhI8/tpGyLUWAdbzz61OlqX2
GzdYeE+yiKVTECbsFb9eoEYejVj1PiksfATwaTH+DnTrwcs1TZW1dBFgLRnVUDUo
ju+e6ZCEenMfnuB+FURq0jwT8o44nY75ophLzzU4KDSHd2VvIVC+C4AdNcftF+C4
2vXvIZw2qieOKaZhryD+OD1CaLQnbUARWCYxzUwxbs76SQrrO2hnwyWw6eDRLZ7n
DGdk0RH0RQXBBiI+LrcriTO8dpbLC6cfuFKcwBC3YGTf+3C8AanswZ3TfzGfxd69
TT3aXgjf8TmwlDxKe0I3WnM9GszzJ5vLT0BSEL+nQyMzqEbeaeL/SQjacDFD3d9g
ZRNXiqQ+zMkTx0HTnQAfaQIGll4n1VTXY3diFn8FS9ExoJlczIQvfqJawCDUypaI
T+RN4Xr1KuTzt97dzovL/WsMLOmLolXLB9wkOgUYhQmJnyR+kWnp9w2pBtLmNr98
WfV6HVfwqfOgFHyQm2vS4uD1jtlSUSaOhshIls2oxh38r1v950duMT68yWaAMpBw
UyhLYN8bxPriNQHXtZrYkrGHfqPfj497A2DRUIAObauzuYM017oADcESKqarVeCB
JA22UndtyvH9A0PHL6FIFw4BSrFeFgHL7ulNj4wTb60F8M6TSSN5NTX801yVUTRw
D0cLUnqRHerjcRWS4TG/YA4GJx6brxJKzpw+e61d1evft6QQLi3s8CvdsvBkcnhd
bgA95RqhZ/JGA77zpez08bVWEqOPIEJoFOOYo9/4lbozqp5cnIik+oOJhGsjEv3u
+ltgXgd8bCe0J1WbkZO5iihMYMWjhpm9G/t402hPAf+IaweDKw1ssczVtZAy+S0d
rIWABB4BynJc9FHA8nmUYed9PfpIUTbhm71LlgjOqhC9gavmSkaeFpFdB/XmeqqY
zC1J37INoRoTf2U4oFWktIfgqakhDemoGOwAmnbbDsFAp0oZLEzLULbUJe00E0IR
NJu1bbEGN9hsxjpr3pvqF7AcVz2CW8IUlO1uKQcTsO6qTCTQCXJzkvZX/IvMIDVl
Bk1riktLtOVQy5s/71M6nfW6+RJXL9VgHIOhPy1nA/IJS8neVcQvqn35VQk1p50y
p4HVDXFCd7JFV5S458Dmp8CDsGhPEeYT5v1ngFnADaxG0Tn4TymbnqCJOkz6EABr
+0VuXfW1KWX/qNDin72Mb+4JYdds0NMxvhW0otaGBp/mNvrfo9Nuhy4f+RBg4pz6
akiqDLl3RYmAbzgaAAWVPLWrTqjU+a6VTm+1ilZ8cDBc6Rur3BaVjPKjUWnyzdUM
wVVCdVn7Xmn3yfrAPABkC3+pP97hxDwKupS5FXElthutA3TuHoZ++lbo8eM8L9Di
CFVMiP8Htr83/FJKiLmVrqiB6BWiXmfQSq+SrDqK4lGq/CTjiGvwVtfB29ECrLrz
K1I+eYGNcH1UnkezBJEecXrXg4ot2FSaTUEpmt1dh8oRMPoNIjzY+g8jiUrwqbUe
t95Eo2iruWV8B8FgGVyae7baQOKOWWJ3OiFCVbZSEcpwO7Q/n/j6O/bN2pQod5r1
f//Ab7utJiqKrJLNnF/XwlGAB2XM37PwpZcGc8nmOEDTbqD2wWf38z3Upo+OL9wf
drAXtprq94XsdONg9d+uu/aAh8G21N3p7R2ADd8Vofc1O5ICtqwF4NsGCH7CZAot
E9tnd7+Lgf6D/qchGEP44JizvGnVyRBb4VR78UDa55z1QqhdVItRVffvxkrgDxvV
Xd82tSuBID+mVUuEp2c69xJ0VP5UjNP0ZAqlzhFWV5Qetj9erOVc+V0kE9bPt/kT
YkNyoHpIhfUnBl3CLbeaFgCOa7FlJVpfgMSmMxF0M3r+oqe6ZrlA9B70WHsCSo5v
LpAK54WnTqmF7LzbddsjJmMc8A5lABgP4wUN1r9+PoeGiv1zcQOyWmk+3zyaRdGa
U/muwj4M+TFUnlwj6YUWaULoHCtKdXtSCTC3RTEIkc5C35dRvwU4GvJHo/dZa8CQ
aA6q9tmbOhQ/lEKc7k1flInGyzJOOmC91o1a0UAHnDTw/LkA241ggLNKFM6MJCDT
4vzgCd4j7iRRyF4eTE+5cJQGfGIYAXqF4B9YOu5EZ9NRElai2jZeOUGt92HiCTRS
49dWagsZDompF6ZEwcd6qaIGXo91I1agb7TcSb/RNlqvuIsQPBTDoaIecLFKI452
trxaJ4YHp/1pr9MUKPD4Bi4YEnxnXESzGhjK2p7Bc00V1DLt9D+wNg8vf2wTCa7v
H1/i7+nQmdWVLNy8NQQnHfBePMc2zAoadu9ibGYRj3QQKM95MspPJAFwfYoiBS9D
QhYwtOKTJVWzMe28gjR4dYZ3gEGq7RbeB78jsvW5IHGBFi2l2QP7DcEPAeYDuwD+
u8Gym7OjGHgteSSp2oHwNKzqgEHJNdH76tqhmGJPlrZ9Ww1VxS1I1C/KopoCblb6
LViOFYOPQjZOaw0athsBxzKSmjtBXP2dRQkd4BuOcuzSskf22DORB9TGrdy2ACTO
YcbMiLu/BUsaXGOZSjN9qFsyw/LLIgjv/WeShu2qfBgSnFrwuG2zXQJEPD1oQusl
fkatO83d35EJy/uk7oTIluTdShOdhwsu2JyDfoqTSR9a7bYfb/3z09ueIRRXTuvl
Fo49L5+45io0mYQE86ziKW7vbmndnr0z57PlHEVJaJZSSYjM+P8rCe3Q4AYcWiZj
V9FOjmli0CwuYqYPCc/cFw6ZvjniklAapDi+gDHQz+S/nkU+ZnuPuSTcRx5G+Qt7
0eUp6Pw11KyBtywMYOimoD/J43peP8RoUEBlKCRZ0i1Y7+QuVZLgnu2BaHnzSJRm
jMj4t1MfX8LSJzAO/6cRigi5c1miycTIjLowXMHyLMv/wFcn6t4tLIjFH7C0hV9s
gybFbEMKVanAyYRdcoz777PiAPSYJM+y6mKKeJ7O0PDR488GUb6X9VsRunPV7mui
Ee5NRv8f1M64TWswAVttvVmG7NQnfd4ZRSlvy5i773NNFdUREzxVAihlVA/WJKDJ
oqmfMSK+ssqIs4tQeTGLd9ide2otKV+nPV/Z9vrQos56c867/GiY6H6BATBSR957
Yo8+yP9NaIiQk29PF1EeeqFhnvdvrF4324CDFIxwD6vccKUJJCCxkBCj9k5kR0Pq
BpimSEyG9obKx4g/WfiOrIihrJ9Qob12xXZj8S7c+/wzaqaS+V2l2DKk6RGgOkpa
b2n8dUMwZysEWaVLUP/onOKkwaDY4+z4QHmI5FdeJMCqrUj42hI4+Bg27LdA4F/U
VrgUUdL+uggW1RBU1oLPnG2WBUn8/P8ye1lBVszAj8HriGXUevbx2loZH19pnLdE
HqMh28wTiqGnmvVVOJRqAzE4T3Z3RiAW2FuHOBfMnBK6oG3dnQbrwwYXdQ3xp60D
f0JBzj75hh7C0Wx3H+NaeV7RqvVHdjvd6TgbWJLppW5GdzAsAITbrx6dikrU31YL
o5vNNJnIs4pghbUrU5xKSwl61DpTDqOdXDm73jKrIllHTaoq7ypUqV1ZcnsS6bGQ
sdsvTmQa9dS1mtfGqzdcgL7eM8JVcHIaTNQKToTuxe9ioqGqXK64W2LoG0sFRvat
i7mGGPdut6rzJp8ziX5i3ur2a82xg1//gfwpLaQE9KgohabDgT606yc91qGzc8nt
6GGC7TjO7/ZFf1NZFBHl2nUsBeDb4W+fdRZTffzs+G1g5ORT5MFXHGGuzMWaPDW9
jjbf2FGvrI7stUJ4+/hpaQTNlbunpicvMp9JknxtvYPYZuvL/uXC4QlkmmEAuojg
m3j/y+hufceS09Tg3ppedJkO7i3gr89PdG/bNdh2PDNTgnI3akextC7mjMiPV7wE
YRyPQ0+ic7BJzOySIva2jsVHjN4sXs0VOR17YRcA9uurhK/zXY0Mbj9IgE9LYInt
kVe8WqFTjq0c6eDuxiN0rnRMhTB4cw10CCLgHe93xMknabyeTjmecb0weLUEi8la
vShHFcIcd10zu5wngeYsqMjl9wp9np/AdSqPGvXxA+qNIZat1R25euBT4fj2oDRB
EGHrlHn+eYj1W/oeqZMzSRnvCIhlOMItkrU9RZ7RBLrdYr3pO1MIUZlJqyhr8zJ9
n+Z+cdofRH6cObLH3rxdQcNZOh8Q0E5YVhyTrlDxUV4GTv8gx5TTeoZW19Hz++um
lIRBk6ZrRynh8HkR3UnksSGZsazStkB5qTbONJD0Kfts4JbRFENh/zAdz2Xxt/RW
4v4DRmfxDeT564WZQdgjCqs+O0pWG51m9OTBXj+cptdP7oijoR0TYIWOowzIGttX
Oxz/FpYBVNBsUU94cOyM3jgxbsaw/kSKCXYAaQcr21cwRePLaIUtvGRbpxjVI8IV
WnneCEOPSbrCl6DNFJF+gJWeSqN2fE3wjwnx5K7a/vDNGfZHkCwz66oP/6QAj3sV
90GktAM9vgVZdPPMtZEBXab2TvRFSrVLpDWNYAB783GR7503gZ0n8Wb3vNvhqL+Q
1PZTS9KIMbKvLYwGl3yMp+t6ajZLNW84EZ5YVrUWb4LLnyNKwbmqdC4Ncrsusjar
YwcFxsTqo88zb6P74863q/nNHHdSstI2tIbfu9Hct3ml+wWCQyoXoS+bgh90NvB3
6qZc5kTsD04XBuGANa1/42lTj8Brkztj9szJjuOpLCSLn7UtOiSmLjLDDzbaK+QH
Wy7NO445NiyKo0i3YFPPJw6TYlcgsRTGQyB8BS2F82QwsOZu46WFNsEyXwGPD/Wj
zHWKgOhRJqgS5jIL2sX98C+acqPzRl4JEhDN0JP9n06z36YHXKPdxr5SNgap5jv8
p3WFBXL+qqAQtC7gMUxo14mlcybeHQh413Th1ABWKa191o4nyzxDqF1HAlpYwTnV
wnL2DnIc9NwYeI6XqmPeib67ePm7OfAqiG9PwBbNQLsIHtWx+rNp/dDXVH6Jwl7C
LR6EtNqHrXRjbUg4zze0rG61n4PShDhGUGkiDoF5KX+lqc9+ZW6+JmnDHRz+b0UU
J5kxe7INXWqtTz322ptOrGx6gjplRZIeAGmzMTkUoxWcghcwBVYXbFcUfKBm6GVk
r8iVJHsPBosepd8UqrygGMK7BmPAByAmhEscv/Mx+R7Bh1B8b8PC7ebDbFriQi5M
+AbZdMPMVm/y5Wult54UfzymuFLuzbl+kUwou551P1gH8Zg9mFk9RPSk9B9v4LW5
mTXV9sXqzc1dtbgChkhOmD+rY8u+zXLVIpN94UsKiAI0Mrj3P+KxOpbcFTuoBpzA
BCaryKg0ej0T8GnzVKMxPbbBab1pTSQfiQsXIupIE8o0RduljWlU1bOxIIyH8Ofx
X613uFeP680Xnr1Rhoi4zhdTRft5bPqcfpGuWoL8JST14CCGlAgfSkk595+K1kvC
VDmQgos0WimX+5Ulpql1VhScPXAYE3XTBtWkE/EPoYlu5Luh1xhdydE0u3EP54iU
Ha8kKndDmI5LpZCWNvycYwSDnw5T6W/XQ3MX6DmjAcH1ml8DFKPevDchhy7PSQzM
qWN0FOf35zmzcGtjS7AGnjlcLsoKEYn55B1LwzUKChwHyRfGu+vWPj1npo2+tnDN
Mh+bX7cAoO1q7ai2fPnMgUc7PEXyqyFqkT9qSA6QG11+Qs2P+hZxCTOnfBOCTJAQ
NbiB/CcFFVxb4tZEX6N/SvmgZbekbMouyIujT58kyVuxc6a1OH7UuBJQcQqvdMrN
/iYjZthDslu19uVj89tZZN87JpLfC53kgufI85RMHskbn35Ei3f6WhnIbrAGHMaM
D34b6SH2A6gsYPweN+HhyN1R4ky8L0OegyfgJnfMHLNBP4SGgfcga6wSEPRGQG0P
d+BbML4Mp8R+s0zO91h11G1oPJCUC75XvRSt1NsdwLZroxR8EOVi7xMRznqfiuAB
lY91GRA3hSwASoPOArGlKpdzfU1B0i/8COabBPsd0WCRThbNG8SZPQ3/JhFqEr7a
/ffGGtc7ImyJJefAdUs7sVPE8Bfq69kPoqgrt4KOi57dqZph3Q3XFe89Li8dn8h2
ISUYIdASMt5bEDVhyKPDvTP35He9jrdnF4aSKxJQNnYEahM/pgLJqJcLPgTbc6Bo
ZuDaaz3PwjOLJ6ZjI4f+MqxCip+vA7hpw/7WiJ1/DWeB3cxyPJlu4b2u9MOVpEln
tyWJEYkpODfrDz5/CTJ0lQ6WXhA4k/H1rvg6R4m1TqvkpJhBUVtdOPWbF+LZbKvA
qM8Aj8Sl4cUEXDHGAXwJ/9nLwBgGer8lC7V89dLQQ1/R+a1i6yqPInQxEetQUfym
k60uBKwID5daxpY8JA6Cf9zlY3Z6lJjYySg1M3TQ/nOElXTb+AkSkUN+7Ghwuqg5
6tgm8oFF2PunD1x8i9SaXZyPCkmNKRh1uYVrLrkBxH6Lac9ZxnDvDqFnqWZYJc7g
5nx2/kaFkUFmnuEjj2qmj927hQJ6ddHzuqBpvAbvrlj5cnPkBkBH6FUCTlJmR0/E
ASWJs9FZ1glxI/AZgaWZfEBKTiahslrX3PqLUEX7Vtm2wk88nO0GVoShLFFJTI/I
EMu6oAwu6AgyEpf58S3gnY2x/JU9subQcYVGZCBVmZDxpOpWmDMpBB2slSfAyX6I
R02zyx4Bgg8kuBH52/Na/hYnHAsd3+iYmF8kADkFc9VoSaeZK3a+/qwurajJoCrk
agWODTnKjw8rkRyqQfbTrbggxnio0fqs/RWFprbm8D0Q3K+hq4I5F71drSnRYj3H
SX3yfNoXmFZ3JO8RDD2ZUqbqd/meS44qhCEmGAWqan98EdOXMc9KzuZ+yx0dkkZs
sS9wFwcC/NsvMJ8hyGgARlzh9ZGQT9W3JkqIHCKDT2fP7CAx5ogwM+M6A7zFJ0cM
skse5ZOT9Nk0kChCjKnteAiuOvXAioWC14akFszDCEv1dmDRP1murFCnsHC+Xl/M
UKqAphp5ybMdESeGI1uJ3DDLEa+oYi08GdnU06Z36e6iZgy8JeQ7IYvz2FWmZYPz
IYuP+xsQnnz7muLuPfuN7bAbEKJkvI4HZU0lP+lkMs9/vZtEexAvh+/Gk8+1FpPs
7IxydMIDmBQbFuNn8mp/LUoBiS2aZRP4KuW0yI3f8vpk6RXEZgzFzrV1duCClAa7
cNEUKxVKniDOzWm61dKXuEjXaPzmofsOGvAvvAdAIGli9uoAdh8BiaqCkieEuqG1
qcZeF+jlkf6ZhMH3mouBFg7CT4p9T3B4cPW5JtuMQzdDOhYYhTmCcjOjLtGTG5nK
chTs8xH9WC3+mUI8sTxNS/zkbTe2sXRQAAgPpMTokuujaKqlmhoAgnZcxM29dn+e
TWiarMqJEwOS24JhJA8JwSd7OKTl8vjICd5gb2bLUsvDphzFpM91Zzc6uAHSJeys
EKWNP8oWsjvPAyLT/RImhdNshhi2ZYX20HRXmjHYmfpObNCy47CvGlmSlgwFlJKj
k8RnhteiAet3JY7zGtq657uYKmimqAoC1KldEdj4MxXVt8FPDL88AgWP+Ajtmhi5
T5sAVtOKmJguNIZR8NByCSXNhecdFLDWpBrXJe9l/UgmrA97BBAaHDA5O0DwJ8hg
j34Mjf6rSMi10bmv+iV07neXbvWbLusGpL1BvrBoEq5zZWV0t0tlc6A0ypfea70w
KDYgr0wbH4QPRgbfbqnPbPht1GXfGAijPclVwrCs0AELeH3G1ERyLe9kkT2bZeua
tmh5dZ7XXjYVV6kZUPb4G8T7ydECK7z+fTkRp43bQiXV1xaTNtBI+gM/WD05PWZo
s71TZ94hWVNVGsneFqh0LsLql1sOjSk++57IVdHGjbIdWtQBZYQPpMcxAwZG30H5
YumfaRqr29OavXDgiUbLE6z/dC1AafH0EL3mXdJMO2dkhzoIjw0RiOEv+DNp2i1A
nEOre7i58LFNEPxlyuKfc9/aXDCxLLi5mLmUDnjf+OkvhJR1YBarhmQtnwlsz/eG
h65QPsQNCcsZKEIrAindnSYEOmB686lCqU2uUgovd66m5EIIHFPrlkkpsjyb8GUR
U7a9YLA1XwVUgzdidHQ8rIPFmg4weAHh+sZOhDkz0z2KIhaqsk4Rp2ed1wUGi8fB
SV6pe0ArKVcsKiN4ieEAtEqhEu95JEj9ycjqaKMlhtwyBfm5Wss7MZDLtI4hvLyQ
jnjOnjrqo2mYMgN3ZS0IQT1z3xA2tUjEImhrYEuRfRy9zQIzp90IXFBKCwEH5UU2
juk45h/EFhgOXT65sgZ1+h7aHaF89J8shQO/7mrOizDHD3TasrfX8yiHXkx1bIjA
2xz4pO6KDtSPeVvVjay51c5Mt7HF6Me+k2bRkiLPKf8wOblCsFrMdtJwftYNb9P6
4RtHxjUikEWiPEJSH0ixE7j2QNSaW2+GijmsKfVc1eyAYZbk0F/aSiO5Kezpxxm0
iJCVV8I68xNhBWVUKfif2A2zzftN/fw+ZpqLPeL/QxvxAynR32Eni8pwxVLfrZWn
bElM5ztTzJAsD2JyHNO4OhHqIgFCAqPESJB/y/7wfTmcD93tAmUCpMbLjqC2VXJu
M0eJsSitVlNOcqsTf8KArYDMAEJIydS3F+lJj518tn22IKogvnHOdO49q89ite2I
xnkNiB2xrag1dw53KRzlVKaZUdjGm1pOP0jvs062O8BIJnAdY2fmMSxeXiws3c1b
KGIDE9LyB9mub5DHqhsAs8hOvij+tQ3M6y0eSwGRMsU/vT9uQA7d/KpsOGNoKcck
KhCVz4KcNbvhNQPyofzJEL/CVzkB5slMhCmU/lLqGpGoH9T+JnGGjGcNlMp1++B3
2yHzTIcCElXWlRcc8vuW2D53k76t/7RAB1l7aLFmkWz32lAnVGTL8LiDrqFIedP6
cULAzNYbiF/o3zf4rrwuRmVFthpJsASNYOe0rz45pKTI6+QaH9ebGO5ietp024kC
ZE6HJnnYFx7EUX7yh8DEsapX95D8GaffQoIrewt70q14qvaQsuPMkkoxzGjYB6Nt
5KgbEUq6vmQPQ6FkJVlbsAU8kvHUQxnAG0AxTVzuzR5Cxn7n+uAw/rlU3qwKZAHX
wTj1ghS4Z8cA4Z57tNblVAyNuMcjO1a6FX+59v2DXazN0+ayJCKNyrXYssYfRhvn
Cs5hfUngwtVZYO6y1zYsSocolvqns4wuHuaU7Se+F+7zyXrgqtTlqVJtp4U7Dq6e
zBlp1RcnYBqxok4kCldu7SDG1eQ9O3uJVZQ4zFfrXOmsVKWLiRD+cGDW393+mkky
+hlr357GsgJxrFNNcJGSq+fbiJC6r4Xu7PTGAnCwEcuL6ojHmm3TNMuw0ntYjk6p
G0DAlr+Qb7UnhRxPkGJ1osvX+hfYph7gZenaFQKxzokle3YDGqHL/DjdHODVWh/m
T3x/RfWYJgxaon2g7OQdL4iH7H24C3WiU4uqQ+CNgjkFvipYR6TIf9uCpbS0fXnY
TSHcERt1SK1ZjL1rpmyOrNRDTJpAnbhDr0EFO9C901IwBtbyciyTcfQ5bdrJc9sF
aUOW+bVDk65TcGhRfivbsqoBjJPoQkcrQ9Zo9gJxlLJgEA3AgvuU14Ou7yHbzOGS
fY2v7Hhe6vrRygT7t9l03wHK8CXLZL4axU3LQb1m1g+DjFyTPElqkFplP1Fx2owd
7yPGgKhhRiTnEs3vl9KFwyUhTbBNgVompW6T3gGaS0E999ftVmU7bmHExQmVmrU/
fc7ANZ0Wojqmo1FeeBugRHOMH5LoOyeyRE2HzMD2c1Oa0qtR/zZzCAqIaGoJcE41
fOXxby3EhGJMWk5Jvp6iSXoI0D8ZcdIjXJAWYIk5TKKhAZHGq2fQJjA2W1AOpZk6
fuRcIPjOJdh6rmlxepo+w+oPTu7Ezp/I75a63Aq/x61YAmKXC9uylB81XxCe9I3X
nE+3F5nQqOPAb+K2Ypt3NM4zpO3HQgsuQM5RYYO2XGD8ORQx11r6N4/sP4k4leH/
7vmB7Qdj+QIqSUqdbt7AbmnPGCAn2XSpgdffimKvAe5DmzIiiRpY20MZMaZcfFDs
P2T7fnPZql7q4OfXHm7LUanzM4iP+GSoofcjKt+OFvRKgOhEwpvMs6ZkKfXfjJfo
PP0V1ItD0s/F/GD/r4qKKY1cnnoDg6bAkCaNhgNvHklU1TUajPiWkLfFlsctV/s4
KlSupnL5Lw/6j0m902SetROUpNMxTdkQmgp9DSSpl1YH2Wb15N6MSbEh6tT2PcU4
2Opjs4cVhmd+/IIYNBqLE67yzximMA6npZJ3N9n6Ob+chgvgQBJAs+5lxrpMzhn9
8opQwtwWj7ZR90qh4TiCUZia1446Z26+PjBwU+JaV97q2o2tBw4RXhsYi7CmD5n7
Al4T5BVlSU8eHxLHkXvANXix243yf5ArdTdi2Y6AtPv0kdrgLffFizpe+j2SE3fv
7NxeGibhKZWn6n+dQkY55sEOcctFz7BjcJ5HZkylAKwnPqAVoh08CcUiVJGhPsnu
0F3IcvyKdnCETYEZSFnLjwiSfSVIp7fP1yrEzjIY/SQPsElxq+G7F+nc5Vcr4RFJ
5ZfJkWHZnJm2l5FPvSBylssZegEH1vVPRkt11ZrxVsYYOVp23zjHC2yvwAGWoqqF
bh3rPMO6Lnk1zTti0hxcg8sRXKljCS/hTFm+w+eref73zldRH1Wt5wyEHO6OpKrR
zs69z4YXd3SMciOZOoWCqS5SwOJwysiVRuhqZH3wUuhBMVg8b2331tRWwX+ADS65
ty1S9tUqU/ACDFC+A5COerB4FNGh+kNxRgvctXi83eiCw8FvlrXdv5N0xufl1bnQ
s8NH9M6rRFL8vS1t0BrH+nwBkYWxThinXjxLQx/xBZWIwhYsJy6ilw41N5z908fk
NqebIFBXwKzYWXOLkQeGbfVaHL77HTEa63oiE7WMbdMVazyrN1So065vmMvbCzMv
OmTuLT+c8yFIRyHfSjY+kgCZAbzozjBFxHaEqxFZkG6cilfzcvlNguU8bzHMGLIp
CDtoaSlyt0cWiCJ26KWZRc1Mrp6VeJ7XYNKy1mMN3rK1reYgFDByhtGaj/niI6VC
8wCNfPVT9NAHCLji6Zd5OwV3oWmYAJfjoOq6uqouSVhKhw3xIZF74kFN/empu1dt
E1a7HbmZoqcCWME6MPzHerO11jGM+xCiug/7bz91Jjgun0Py3L3s5hJB83h9pfRn
NmW5K710A5I3KPZanAbb7RuB8TqS4+LW1hupUA5Z28zSMibOPf8ywk/QepZVeyJ0
/gVl4HHZglZexTJuI3MAz5p0lPxqczlLSwq6WLR8DIvU7bkCk34IkM5eFlowD+PY
1EtkNYylokHIQFcgEDk2CTU3JaYVgL36Xdqh2TaIDOUoY++27HSDUSV3PJ13ZhPB
XXzSSh8p5IK8YEPQMlRmtX/Ilu4WJdg5jpaLAoXW4Lvx5AyQerQG6Y0H0y5QHdQP
iyRo0FsAw0RCETCigC2K1XAOYgbncbMk4pUIvz8gdIhhb0CKXRyBOwiatGNL47nt
JDmfOBL0Kl7aZ2u8Ymie0GPrTW1qImVqyS5CvWaCUwFWyx7qYMjr723Dg6UX9Ewv
LsNP4FZJW6EBrZr9Xk4hHKVfNjGXQvYu0ZgsLV30aGK+GXp66a08Nqydv0DzWACl
/sZHq4KZ+1/Y561m6414FPnnoYyF9bsgYkXV4DW/6tHQbr3TctQ0w0nYZ8V1GzRU
lpU00VCq54xcJxlI37FhU+KVRAQyppqlNaQql3fo4fbyUrDJWVldCpRqRMFQzt4e
NYcRtmXNr/rRo4LN3YcEdoV0y401TsKLgLdLVKRFuE4OrNxfO3tL+PZKWsRVkWxH
ZY9SMutMjln6Gsu7aJRm+pr8oPAdaQMtKYU153/lX7iwmmr3paR5z30/gm7pEeek
y1ZZGISw2O7ZssNd4SbtEZxyd3vB3ZIPBuZeNEVxHoAaeTKyFfdPwnKaL0n8ctfI
oJ2yA3lMDLa1lsXeIqv5k6BhrnVud5vO54NEVL9/ueLxjaoIdLeAgsdynRnGgjTh
c815N1gH+rwQY9Vamy3TFEeV9tsLtknlzAN89cUP/FDwX79UEkIIeQw8cYW0h98u
2k2f50GFbhcw1IjVzvI2JHh1QCY5Ao4ltleN/vlXyexUa16oKiXbJZufBxdhRN37
WBC2tWezmZg2rjwE1QvTZx9zPn1Kmt1uqW04HP/MDtLuxZ5dgG3hHYog2AG+EzaC
hFsKShYeMPF5J2gbrY9iFZpGvIKqQ+9vbrcIsKItfvvcdGQ0ljXx5lTPKjPiSzjX
Ft2g73PBgv188lba/J4nkljljxQT+Rpo2wR0IYu+QGO63llRF8jWLCGZdH4kHwak
fCIv4A9aDF4aShmn09nPgXrcaIftX6TSJnMvS3Yrpg9o4bPJAm1m3v7Jd97AnDoJ
sPH9qPftKyXUbXReHZGqNOVE4QxcxJeXZfToEc0LC00nlj7vs0Sx7YtKVBPQpV4A
cz60rAoxxD6OokolCx636un8j5dY5vHxc/fEaHEtGRSf6O07laSC7LiTf5N26aIO
pKqD8Rc2amTNFqt0xR/grC0k4lCP/DQ45IQA537i7xUvfQUt4NsKprtKakEd5wQi
ZMifUbmNLRX/PZMjOPGFBKYhcIPlE4LtKml4qmRLJtnJ2TGG2Rxi1vimzYnSC+lE
iClr3IlqN04c+XOtcA2wqXqexyV8T33dyKbfXVFOyYdqo57GZAk5oJJtCvDngqiD
dllFNbveS6TqgtU8L95VXyWeWiVQ6ufh9jvVomStRgzn5Hi/GfQPB+qFlcVSLIEZ
Jp/TcY5ji6sUmjeBpWeDL9p7UDfTrIpxvS0is9aFe0G+SjB1ikurYn1CEPlmz6R0
A5RW81YPh5vLrNYZqteVLm0pmiL5zRAaXKn7lMgOVGRTr3fLeggF/VXznR3nQu50
7AEp2iwcyqlrPdGv4KuoFHdLoYh3yfOQ0a39IKNa7fm7zcw7tZgktRLhLB4cWfXd
V86kN7QvlBdui9YwlFs3KM/+ZOhbssQNVsnjNdExTgEQ8Ve1v1apDOeAD3Hmv8Hz
eN6ik0Tf4elOgM4L4kwlNWYj/2bQdyZjTHMx8c6+Y0BI85x4Rl2wv8kEgUXTNTTq
KPhuIlyrsa0NIDgy/uSmIwWrCg3r5bk8BKemzzUfvwVTG8BmdxfQJoCUUsqkKaxe
/hZT37TABbrgf57aZ1XOrvurMFxAWhqhWkuTkU1OTZXc+hBL3sBHvvPyYFPMQrXb
m+hAEtnJHF2pVwyt7gLMkon5xPN0ZrEYsTMBz+4mIqWOiEHdRMyTiI6kwKPDTYFH
/nk3t0FrgsWWWiyhTrWMOc4KDiptkYND0mWM3ZtgqtPRo4+zRatHpmgUTlM8QmFL
FK+ekifxxt9Us43IKDtrJnIJebdAax4/UmArI+iuqe+QpLaQcj2icWoMOilY2aC1
rNXBU4Ts6HXqTdkvcjod0RaaNnTJn3OtzFhS1JkQulgWk2k6dU0ZeLwHcJowNMFo
Uq2HlQPAM27+ThJzsvlkbiWv9U9rLnh9cpXb5wbb21JeLj1pSe6cclmcBbuGnIJW
np4cSHKPPy8/BpS8uuYZsXoW7adrO25nPviqjKCzqzvgJlluJrGsNB6o0p/Q0t4m
3gsNaIFYq0TVkwQMdaVtMHv4lEzU/54CWcrCztlr/uV81s2Lep4/lOhOUJuOP5fp
E89esgRZwcpKX0KO/DwoCy7DxeNr7eAM+TlaFns2YpowqQeIrgc0aTBQ4UnaNW58
/kN8wixrL53GC2myP3SYZitC10V/vG2/cdT0JAV4zySUefz6PQErw/x7pWGMK6fY
04ahiBtCPhLZmIm9kjqquMluh8HR00nJJDeAyjWdSvc4CB4TjoGP73GOb+/JQVdm
WmeVa2vIfaD6Md/QZRd4Ge6PuXbNOgDHYGokvi4nOH6iiK7cdpoEnf6zHMgsci6w
bY3Thq2tm83OtuRCg+I+DBa/UxTTHvlN0i0gTx0L4j/UZ82yXRYsq+eHBTJYjEjC
oTHY/SCzfZFvHyBfyICi34yR7bFDGy6Ui4FSO0A17haVTUFebMgwFtlOy6zLmD6x
YfLuBgh8luc2yCOxMTAavZXUR+i278XtLPe9/RTfAhqPIkRb+9WKUEjZdfNQcs3v
zzSxUJHyk/VJhgQbTJMSNpbOePdre2ZQswH1bTaLwFcp8IiFfhmxuSJ7WHrvPlT6
hYcBT7oX88TcUnw6L757UZVvHk4dGf5BGFNRfjx1nC4yzDcmC8Tf4wZxnbfYKbaj
5OftEIar8keWDCLsC91wE00SK3LanEIbNv4842dpStn3scuDet2W6ekpE2zwpkKE
nPwsv8sJ4KX8oEu+BsxulnZluvM2HjKI3LtZ6DyxxkqY0i55kD4Rjnh0KUA/O+5H
mxdMIvFQg9zXTie/OoqPz7sYWn+iU31F3/mvvXf68rH2CgcMmA5HYljYxUDumSad
1IXPsOtuzIbhB6HMBWFF0EI5Ipgem9kjaOt1LiQHT024wwuHtxJjd6qxItiKH+pG
Q6T0Y7BA2dBhXFN3ReJpSHy9ZBv4/2TnOSkwKpwTOY99ki1M3AItY2Br/VBnijBj
OJ6O4bVlksgIvcbYi+d08El036QgYxy5kriPDbJSJ89DYb6sRtqT/t3wjTRl1p1g
DTbmvQO/o+LWWSAD26UGuHxQqr0ikePW313iIMy+HwPUJn7ssdg/OTg3pqJwVj7a
GYfeMGVUPlf2iSgEXaQ4bjd9MV4kt2GV49ryEJSGCAnoF1Ei59SmltULkKzjEwgA
tGnzjAGv4xI1KHw2W2JrY/u4y4Pjl5Sw201XxubgzY35S/nmBDuQ9T4+y49Ws5sS
TUkAFLE9vp2np9ceZntixKgRhbstDJRv+uHdCA2PJzx+UpTnBEjPpcDwx7ONtKIh
s0UVctwjVHr2ixLT2Rhb/uJMQzCeQxABqdGx/9BLdLqEoU87mnYdi7rx47nKMkK3
hMF254ejWlVTnvrIamzAv4j5lkf1AdyG/bjPvwmlVK2jQFG1hI66ev2e2Mfd26pp
sjvrQzc9WjmMzyj890YfgqC8yU9mX5XN0Ai8B6HMW0lW3TyNncfKx5QyK+XOjCf9
bgffoRXXl0McdC9YZjxGXECO3he/9wmhEwYtcjmnkaPWVHFbJS0JpVIdX17HtK0u
0DaUqyVkQLgexqK9bDuYcOEnpIpUpa9F2fQG/X7MYbXggD7zpcT9fLi9VK9vtF3B
EO1DNrGIJDeT8PkKxWjNb4Jg4quZ8j5PVxKmgBzFqV632fVyOcY8ylufTNjGQ3Vm
hxf56HJTkNkRRIRxBMSkcXJAO3YMcQIPGcNKpHdJhBTSP9u/ywZZ/N41pPaZftgg
MDw84pURXOXLkSciXMFhigQ1oMqh8/5cby7vCD69k9hckSy+XOjpmaoUBd7onk+x
mSx51Mdy+RGO79Pbh9ik+OfecMfEGa0J+iHM5N1Aebqyw5dT6oVw7j8hMhGjJSIQ
T1K7mQqv+4WyCJZuMtN6V5QrD8uqcBwj7Ep2ZfCZzvqRSZeXAPFlxWH7KXt3JWaF
6JgRzNrNZYWyLOmdindPWMS1ByxFSKMuAMzWeTzX19/ow7DR838tE6vpFiPNlYBB
SuY2y/+CgjTXgvQ/eQru25MDuWbCFE8rb2OewcAdV8iM+Fhmhii6rQ6AC0jRJHfR
EQfjUix6OcqwSIMAcnxZkaJGFjmGnanV175hPN2N+Xn+BJ/LuV+0Z7CkTtQiPZki
LEacC3O1ygBuY2OUBW3OTPxaq69FG2qd9ZfwFvayhbGKwODkMgSyrb0JqRGwXIfv
R4v96s83hfLDXDhQmouc5h2X49VmzthuH4J3tf5WLlj6tHLGqAoU9v7e0Wa9qwNX
7wMW/TXabCbV9P2EFHUXsgI5CDP4wlWoys+6bdE7G7JxGauJLAKmZelU0eu3mPZP
MUcPNBtz3R/6LNkpvRSlC9jwAjXhgd11omVi0N90qQH9Tik1A0/sDDYVbmllwRaz
ehFRmAY8E68CrmvgldYHTzctFEjODVqIrsT4NXbYfNN6y/SraW8+pVJwVEod68bc
oJ1jwf/IXD/2aQ1x7LtEV+itDU39Ggv9ZeWm3wpeL3iROH0QuqkkG482K6/2veI7
90TjUv3pYxBvJPpeIZp21vm46BoHkw443VdS7k1LiqkViKvF69cct38+ZbU7w+eg
UaJDKIba5DR7hvKnwWRXJNCz+RXrY7GZWdPApRm9UtK1RRHb3IVOqCxprpu7waud
3Zfyj2jDUsTI4NWL1McV/i94PZVCWWfh6JV+z+i4UQffNq0eRMw/YmVHxvAfrzl6
6waGx8J1k3BLK1UjAjDg9VkiOWAnlGCSPvgD8rfnlrTRR+nW1SeXm5nG0ZlS82C8
gjw5Z5KFpOsaaDWU0+aYatjZcEI+9c7SEWbYMjtU8psBorIOLuz1WdAn4hExL4vc
A0o0I7KN9GlM+pnj7BR6QsTsBN3C+RnI7u7nB4CMP99ThjuSqu4KKFdgbw+CsEwl
0TzE6DBPAQeskrhoEPW8vuVDQEYmsZaaEmlOs1ZBEh0NHqc5mow25Sp7b+4m0lig
OXSgEOK4WGhrDwDVpGWdDQBRXRPnVmWmm+cjjM1yl9I7r/+GwfAHEP3K0L2YMn/M
QuOFIGcnSH0qTkJITZW5H7d9c4P6rBzlPhB14/HN+4GrZvlZKErNq2g816PPme8g
eIu+5HtoR/BpEepQ+DiqfzSVirkwJKKEPm56D8Vyphyo3GubODdXrWukcsZQ8Axn
x0q3PJhX58YjEj7KK5V7CmKS1fWPCWO/p+j+oeZg9TQpuL1xzYvXelU8o47KpM1S
RIOhIhzDVxsRK/SbTk/Ox/AF5DdqrRPs2D3PBN/9F0pstSu3upPvC58PnAhpVoOi
0Xs/dRJHhxl3OzWPFX1LT1nUt50KuzC+XrHEbi7PyFSWsY403dYzucFkX/t4BSp0
kVzlRWrZp88SXyz37RLXVkV+JY90jGYkZVzpxpMLfvt9tz2DFnEJ+jqwK97lW6rh
v0wj3vdyEbTVTDO/7jXfb7iqrHEybdMUSZTMyZDvmq4JBTBtQdmHHovObpw4zaSU
90zAu/nOALIQSuJtlK0C6DPa6z0ypn8cds5M8+vttnOz2Tl9MFZ4yCtFA1pE5eD1
KxSn/3UtWPR8a+C1LIcmMiftiigyOcd9AyvNDHhjo3uhzUlTuHMLmHoTey/kKSRQ
kkKJWbhQhg2oR+6ZFuZBArQHdzcmatIVLJyhZMTopWNMuQNlEG2+CLGlKpIRw2Pr
yMvMYW/+SiOrH9CTP2q2+AMZcurNS76ChQuLYLANUi4qxrmvnoKwz6aflnz8yd7a
bzE6Ek09mVfG4QPsWIfwP36VW6iMrijhBNK4JWyHUhEh2ZZltDdeexNw24+YYbeM
JqlaROcHogjgvbsEO/+LHWpQr5dUObH5EWhOg9bwjvTi3NARba8u3Qz4utO9PzKo
fFm/5ds7qZiNcpx6ivszzfBYunx1zZZZ1rKmNyte0/oCnfZ68EcLCOEE6V6kJTjH
UEoGS0wkzHA9hiI9AaDl1uRkZchO/jiaVTa91LExh/WdunH7q+BIJGSn7+vRe1/V
l+CXukbI7J48XYK93nFd5rOdeSLoH8tG9P5YbFPYVPU52CZ8NT0sKEDTPVYudr8e
+rChQbwNAkkM6r+Rx0w9z0/PuKydW1FWlknOmr6zQb8=
`pragma protect end_protected
