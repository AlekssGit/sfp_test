// xcvr_pll.v

// Generated using ACDS version 21.4 67

`timescale 1 ps / 1 ps
module xcvr_pll (
		input  wire  pll_powerdown, // pll_powerdown.pll_powerdown
		input  wire  pll_refclk0,   //   pll_refclk0.clk
		output wire  tx_serial_clk, // tx_serial_clk.clk
		output wire  pll_locked,    //    pll_locked.pll_locked
		output wire  pll_cal_busy   //  pll_cal_busy.pll_cal_busy
	);

	xcvr_pll_altera_xcvr_atx_pll_a10_191_6oxhjba #(
		.enable_pll_reconfig                                              (0),
		.rcfg_jtag_enable                                                 (0),
		.rcfg_separate_avmm_busy                                          (0),
		.dbg_embedded_debug_enable                                        (0),
		.dbg_capability_reg_enable                                        (0),
		.dbg_user_identifier                                              (0),
		.dbg_stat_soft_logic_enable                                       (0),
		.dbg_ctrl_soft_logic_enable                                       (0),
		.rcfg_emb_strm_enable                                             (0),
		.rcfg_profile_cnt                                                 (2),
		.atx_pll_silicon_rev                                              ("20nm1"),
		.atx_pll_is_cascaded_pll                                          ("false"),
		.atx_pll_cgb_div                                                  (1),
		.atx_pll_pma_width                                                (64),
		.atx_pll_cp_compensation_enable                                   ("true"),
		.atx_pll_cp_current_setting                                       ("cp_current_setting26"),
		.atx_pll_cp_testmode                                              ("cp_normal"),
		.atx_pll_cp_lf_3rd_pole_freq                                      ("lf_3rd_pole_setting1"),
		.atx_pll_lf_cbig_size                                             ("lf_cbig_setting4"),
		.atx_pll_cp_lf_order                                              ("lf_3rd_order"),
		.atx_pll_lf_resistance                                            ("lf_setting1"),
		.atx_pll_lf_ripplecap                                             ("lf_ripple_cap_0"),
		.atx_pll_tank_sel                                                 ("lctank1"),
		.atx_pll_tank_band                                                ("lc_band4"),
		.atx_pll_tank_voltage_coarse                                      ("vreg_setting_coarse0"),
		.atx_pll_tank_voltage_fine                                        ("vreg_setting5"),
		.atx_pll_output_regulator_supply                                  ("vreg1v_setting0"),
		.atx_pll_overrange_voltage                                        ("over_setting0"),
		.atx_pll_underrange_voltage                                       ("under_setting4"),
		.atx_pll_fb_select                                                ("direct_fb"),
		.atx_pll_d2a_voltage                                              ("d2a_setting_4"),
		.atx_pll_dsm_mode                                                 ("dsm_mode_integer"),
		.atx_pll_dsm_out_sel                                              ("pll_dsm_disable"),
		.atx_pll_dsm_ecn_bypass                                           ("false"),
		.atx_pll_dsm_ecn_test_en                                          ("false"),
		.atx_pll_dsm_fractional_division                                  ("1"),
		.atx_pll_dsm_fractional_value_ready                               ("pll_k_ready"),
		.atx_pll_iqclk_mux_sel                                            ("iqtxrxclk0"),
		.atx_pll_vco_bypass_enable                                        ("false"),
		.atx_pll_l_counter                                                (8),
		.atx_pll_l_counter_enable                                         ("true"),
		.atx_pll_cascadeclk_test                                          ("cascadetest_off"),
		.atx_pll_hclk_divide                                              (1),
		.atx_pll_enable_hclk                                              ("hclk_disabled"),
		.atx_pll_m_counter                                                (40),
		.atx_pll_ref_clk_div                                              (1),
		.atx_pll_bw_sel                                                   ("medium"),
		.atx_pll_datarate                                                 ("2500000000 bps"),
		.atx_pll_device_variant                                           ("device1"),
		.atx_pll_initial_settings                                         ("true"),
		.atx_pll_lc_mode                                                  ("lccmu_normal"),
		.atx_pll_output_clock_frequency                                   ("1250000000 Hz"),
		.atx_pll_powerdown_mode                                           ("powerup"),
		.atx_pll_prot_mode                                                ("basic_tx"),
		.atx_pll_reference_clock_frequency                                ("125000000 Hz"),
		.atx_pll_side                                                     ("side_unknown"),
		.atx_pll_sup_mode                                                 ("user_mode"),
		.atx_pll_regulator_bypass                                         ("reg_enable"),
		.atx_pll_vco_freq                                                 ("10000000000 Hz"),
		.atx_pll_is_otn                                                   ("false"),
		.atx_pll_is_sdi                                                   ("false"),
		.atx_pll_primary_use                                              ("hssi_x1"),
		.atx_pll_fpll_refclk_selection                                    ("select_vco_output"),
		.atx_pll_lc_to_fpll_l_counter_scratch                             (1),
		.atx_pll_lc_to_fpll_l_counter                                     ("lcounter_setting0"),
		.atx_pll_pfd_delay_compensation                                   ("normal_delay"),
		.atx_pll_xcpvco_xchgpmplf_cp_current_boost                        ("normal_setting"),
		.atx_pll_pfd_pulse_width                                          ("pulse_width_setting0"),
		.hssi_pma_lc_refclk_select_mux_powerdown_mode                     ("powerup"),
		.hssi_pma_lc_refclk_select_mux_refclk_select                      ("ref_iqclk0"),
		.hssi_pma_lc_refclk_select_mux_silicon_rev                        ("20nm1"),
		.hssi_pma_lc_refclk_select_mux_inclk0_logical_to_physical_mapping ("ref_iqclk0"),
		.hssi_pma_lc_refclk_select_mux_inclk1_logical_to_physical_mapping ("power_down"),
		.hssi_pma_lc_refclk_select_mux_inclk2_logical_to_physical_mapping ("power_down"),
		.hssi_pma_lc_refclk_select_mux_inclk3_logical_to_physical_mapping ("power_down"),
		.hssi_pma_lc_refclk_select_mux_inclk4_logical_to_physical_mapping ("power_down"),
		.hssi_refclk_divider_silicon_rev                                  ("20nm1"),
		.hip_cal_en                                                       ("disable"),
		.calibration_en                                                   ("enable"),
		.enable_analog_resets                                             (0),
		.atx_pll_bonding_mode                                             ("cpri_bonding"),
		.enable_mcgb                                                      (0),
		.enable_mcgb_debug_ports_parameters                               (0),
		.hssi_pma_cgb_master_prot_mode                                    ("basic_tx"),
		.hssi_pma_cgb_master_silicon_rev                                  ("20nm1"),
		.hssi_pma_cgb_master_x1_div_m_sel                                 ("divbypass"),
		.hssi_pma_cgb_master_cgb_enable_iqtxrxclk                         ("disable_iqtxrxclk"),
		.hssi_pma_cgb_master_ser_mode                                     ("sixty_four_bit"),
		.hssi_pma_cgb_master_datarate                                     ("2500000000 bps"),
		.hssi_pma_cgb_master_cgb_power_down                               ("normal_cgb"),
		.hssi_pma_cgb_master_observe_cgb_clocks                           ("observe_nothing"),
		.hssi_pma_cgb_master_op_mode                                      ("enabled"),
		.hssi_pma_cgb_master_tx_ucontrol_reset_pcie                       ("pcscorehip_controls_mcgb"),
		.hssi_pma_cgb_master_vccdreg_output                               ("vccdreg_nominal"),
		.hssi_pma_cgb_master_input_select                                 ("lcpll_top"),
		.hssi_pma_cgb_master_input_select_gen3                            ("unused")
	) xcvr_pll (
		.pll_powerdown           (pll_powerdown),                        //   input,  width = 1, pll_powerdown.pll_powerdown
		.pll_refclk0             (pll_refclk0),                          //   input,  width = 1,   pll_refclk0.clk
		.tx_serial_clk           (tx_serial_clk),                        //  output,  width = 1, tx_serial_clk.clk
		.pll_locked              (pll_locked),                           //  output,  width = 1,    pll_locked.pll_locked
		.pll_cal_busy            (pll_cal_busy),                         //  output,  width = 1,  pll_cal_busy.pll_cal_busy
		.pll_refclk1             (1'b0),                                 // (terminated),                           
		.pll_refclk2             (1'b0),                                 // (terminated),                           
		.pll_refclk3             (1'b0),                                 // (terminated),                           
		.pll_refclk4             (1'b0),                                 // (terminated),                           
		.tx_serial_clk_gt        (),                                     // (terminated),                           
		.pll_pcie_clk            (),                                     // (terminated),                           
		.pll_cascade_clk         (),                                     // (terminated),                           
		.atx_to_fpll_cascade_clk (),                                     // (terminated),                           
		.reconfig_clk0           (1'b0),                                 // (terminated),                           
		.reconfig_reset0         (1'b0),                                 // (terminated),                           
		.reconfig_write0         (1'b0),                                 // (terminated),                           
		.reconfig_read0          (1'b0),                                 // (terminated),                           
		.reconfig_address0       (10'b0000000000),                       // (terminated),                           
		.reconfig_writedata0     (32'b00000000000000000000000000000000), // (terminated),                           
		.reconfig_readdata0      (),                                     // (terminated),                           
		.reconfig_waitrequest0   (),                                     // (terminated),                           
		.avmm_busy0              (),                                     // (terminated),                           
		.hip_cal_done            (),                                     // (terminated),                           
		.clklow                  (),                                     // (terminated),                           
		.fref                    (),                                     // (terminated),                           
		.overrange               (),                                     // (terminated),                           
		.underrange              (),                                     // (terminated),                           
		.mcgb_rst                (1'b0),                                 // (terminated),                           
		.mcgb_aux_clk0           (1'b0),                                 // (terminated),                           
		.mcgb_aux_clk1           (1'b0),                                 // (terminated),                           
		.mcgb_aux_clk2           (1'b0),                                 // (terminated),                           
		.tx_bonding_clocks       (),                                     // (terminated),                           
		.mcgb_serial_clk         (),                                     // (terminated),                           
		.pcie_sw                 (2'b00),                                // (terminated),                           
		.pcie_sw_done            (),                                     // (terminated),                           
		.reconfig_clk1           (1'b0),                                 // (terminated),                           
		.reconfig_reset1         (1'b0),                                 // (terminated),                           
		.reconfig_write1         (1'b0),                                 // (terminated),                           
		.reconfig_read1          (1'b0),                                 // (terminated),                           
		.reconfig_address1       (10'b0000000000),                       // (terminated),                           
		.reconfig_writedata1     (32'b00000000000000000000000000000000), // (terminated),                           
		.reconfig_readdata1      (),                                     // (terminated),                           
		.reconfig_waitrequest1   (),                                     // (terminated),                           
		.mcgb_cal_busy           (),                                     // (terminated),                           
		.mcgb_hip_cal_done       ()                                      // (terminated),                           
	);

endmodule
