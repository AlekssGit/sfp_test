// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
kRx6O3Sj9PsOvEI3KIVsfAYdwfVNmddMo2qfeS4T/Sto3teEtDjKY7j82fKcUoci
DTzVqAFTRmd8o21hSP6gCVjbXI0xDJV33QSBiWnhbnXJij/cmh4yx0UvbPbD89Mc
lBEuR6c6jNljPBhh7WseL+HdJwDG7hY11hZLr4dLQaaugtP7xx0ZYg==
//pragma protect end_key_block
//pragma protect digest_block
sdhHdCd/ro5gHg8Jxwqb8b34hyQ=
//pragma protect end_digest_block
//pragma protect data_block
tcdJYD/b0Ly2tIRR4n398vavwyYiu7LUqDJv477Qedhv05aZ0sGAvdRz6yzvCAT7
c8MFgTO3te34MfdBbdPYJr0C9CvcPfbR2M7toJD8cpZHgG6RggWP90takkc1VfbA
8IIoDGvGvsuFPUKjtjZTh3SK+DAQjrNPu4tHlCCBZ+fr4or9FW+lVrCrk+qzu5qH
qYH0R0R05aCDL7lwWIC0HUB3x6V0/0uOoqPh+vwTDvl74jFX3adV6Pex2T7aRVaT
c5m/i1cdbfThKNtp6/OE2MVRlItivwfSK//pBZ7azY9/sZhsDrCI6pvnj2tGHsHf
H9FwXL54q5Uu1DyayS1DpVHNdZr9w8WcBxeuCF3wEAiISGyrYaLRiLV8fj9r2GHS
wAYgySANc3w7neZr17uAYKUjwHtxHdga54oTzmYnitTsT12SFLvnmXMMFJgWEOB1
smviEb7r68KAl7sPJhwDSGkePOvsoT0tfcc5gpbW5RJ/ldPhcV7dM6/GfW3aiywn
p3ZFCmni86hkaCqR7qf8yvpF4gGjzb/Se6MlCHSN4OB66Wcz6juFTGmXkho5wevR
y29glcN7xrZqRe0TOQK017uAZIlfQLqlIly1J/v8dYT8Dw03N2Vko0/fgLMJzJuw
xS9fKrFgb8wd1F4C5fRpL8oE0nwlDn9WTNdaYhKg7VgtO7w6Icvh2Rv8cMW51cg6
CcRISVNPhKE6xw0GjUzSdi86H1a2ag/bmBQ0CHa/5383DN64cwPCWl8QDNoao5LU
oyTFC0un4BLYIbfQtU5VXPxwp2UfmRoj/RgzzdyIVWiPXrTaRe7Vi9Iobdt+y00q
e9fSjYzRNZZvS4Nu+5KbWvOTNAO+i1dYmKH1pFNkfR4T+60HKlupMlyLbdlFanCL
VFtASSgENxNr61+skrq9m3OZeUI3ajna2XdodIvYwDolE0mSt7I7PJI9HGAJQWB4
xUjuz1Kbydun3alSiyqA0Ot6ezhJeMSESY3Enjsn+L0Hx7x9g9qYpJPEOilMPnMm
63tBafc5ivCzADw3tccCKvKDwOZLRd1FMIMDONhDB+gTGCVxohAjKFKSsaEDuTnB
YxdDn6ucQyyOgrqtEEtEUrwlDEO0V218bhg8Ikkua8+1jCsVS5IrIFj+mLcOm/l6
s0hQFeHOQbQtJo1BucLUccwIb+yGggoIRiIy8/kc3FT0tg19qsVdD/40XVjhvK5t
ArTnSaMIyFCtfIrX4Zeq+KXwyRKie5Fugv+jUu242wh23LkoqguZ3eYbS8LuVtBB
c8H8Idz0RVP029sdQmXSwnDrEFvSybtJPQpBYYxk+bsnAhCoFhCS1xeHbnyODS9Y
tJlEveFdVGWaJTsVgjHbMesJVq4SwcnR2qmeWarx4VQWRsahwVJuvm21AWrmnnZl
z0k6y5vN6cp3ZAiNWrVVxRf0VTvKC7BwbTpmp5bq3+BJifT0NXO3BfC4bKvPVnr8
Utfvyk+9JUeIITEFrlUbRDUU5T6TdJcurTyGvsvojsFK2kg/6SbF7ZawGJWoF7+q
RG34vUe5ZfdOhT657w+KgleX4PTIPrEXQB9QsXwgNsFmXBEtUqGwRlLed9ZOGL2i
GxKqtcjEuK6cTT0V0HsO7GznT33CmPSEBUvOz54BqWqaqzJrTa6USEP/BxtXcm67
xhB4CSMct1FrlT+pobhvXg1JbJZJQexCpBSjjK97zcfEgd+A3axwsQTL55AAMy3E
+JvVOf512w5hIhVIYnHovRUG42cup/mBAKE+id++1RT8xw1d6P/TDlKHqEYDl2BB
VUX49TqlN/Q+NFPYopaeFNGhdZzehd/0HCFyIDvlWXcoTJNBDcYk9TT38V1wEamB
F6WarP0v+XYWi4XNcp21cEum/+eAuKjjYeyG7E1SHTy5EjchjkAzUVHYT22Yb/ix
+jw6lTSuLWMVilHPcH11dgWbawFn6WodC4HBgVUjLU+HUdP43SNPElKytj1bu61Y
UT1diz3usobI+1y5amfI6Jp5gQp58l0tAs69IfHkc/06jsz5K7ZWL9dAin6Qds19
xSxyBXMLhjg/K1Z+5tR4kEfJ5JkeWcegsvyiQYznSYtG6co/gkkc6kzH+sZNlq9A
jQjOOMfZpnt1NZjSknuTB9zUYbweymEkdBi9Zm6dVniXbUanuLQlETNKrBeW34JR
mqdziUjJSg3uLSWsTKAEwar4xNDbbRoJMgEG2oOn8PXcRMk9QNXA7tyuQlzu/DaM
AEtNQg4ut4uHC2yIA3JrAWu/dLzuregfkfLBQaK/jhXDcOhOUyTfoe/AP3xr5dUn
knkGj9WltPJc7idIsOcaykfiN/07liDop79uZk82KA7wlDpGH/7B2v+X+Mke615R
O/NLy0i8Iq5uE8DRevCpP8Zj+N7YlJh41JnmoM7ns2i8bz+n45CiYiVT0Ysbowxj
A8Np1G8ouYpCa1fOhowS5cy8YDfntSLKRA6rZaSYbj3v+SYnjFdCmxTz8aEh3aB7
8DnXs0jC/nCVxClE2sea9LIECABCAbht5O2LxFvE+0kyemNdKlmcNlN2tfq0J6ij
ALrQ56J4ZlnFfiv4RRBENo5/US1CD85tJ8gQXbcfY0PBnGQMmMp9QDWt3eRjN5hE
Y4OA2Wo3sbLNLtLCXohVNATDIQoEpoI9TC/b092eP0i8qM+5nom0Eid7HEL/wla2
TxPiDPDr0QDeBpXOpquiyvsT9d5IoZcldaza6Wem6VCig3cybJthuhcJLasMlbs4
BjnJ7QW4biEuu7t/avH7lTP9MLPOui8ZEQl03FgBICr1U1MISQQo6pGOoulgwtbt
Hl5ds8RONHa7IL6M/LK51W1MU+uqL4CoXUumeDtP5bhVjDgU9w26SDbVdUmtZFdC
Z34lRtw1i4EBlP8YVrDhFd5t9suUjY5gpzh1OAKwPSczVpQb4tf4Z9Qx+cJCv0u+
Gc9F4MEp3aRYWGu59gp02vCwhe2z8Oan4IMhwMPqoWknQ/GjyF583ihVQ6lDHFGk
0KyckzwgeoN7LM93KPSRd+Wurz+Z0WTC7o9tRgxfFe7R1tZ5NgNrAsWSF3yqBk0y
eMZzG+AuOu91dglTb9hOi/pu+lQy9b1gXmy8l2fVzgM7bZS/YGKGDAzU2Oj7h6Kr
M+0SaDo1sCq2oyMQtshTEhG6VQuQRVExWzCgL3rLcpwgspA1Sgv7VO/1Bj364xb8
zQAgvXpaKANltme4+dFNOqEcrGJoUpnOlNdQYGZ1SyI1yN00nRmjOd21uEsb7n8H
tnIoWjyWCs5Lw2V2DdbplBLveMyY0WDAVPnV7ts6FvBBbt6DqkS5WKYKyEe/tB/s
eeTi3JbQ3yJ+Q2y+4VzwHcXa35FQ8VvlPmeVOweWBGiWFG6nUc1xeSVUOAf0pZTP
4DtQji71s5uk2U7yVenM2sMKfZodKdpN2QIDGhmkNOpzw0nIRijSUBhBqysgQeig
Dcl3s+qcSg+qk9lytEnbq0P/fGITdNNTzKn53RbM7TxGt/f/9Yfydna/GXpniC6r
6PNAjhc1paI8vBP7nl/UZtLxPp6bEF+QuN7uwmQ/e44ZLUcuNm8q1I1hdePcPYtE
PfYpCb1FcsQsQzVeXeZqu07JII0WFSv/HA3fXRs5zmWpBtBIXD5JuMg8BNnkgQsz
tMCWE+LlR5xN0rrVMGhQ8kuItaov8gpRj/5PrfgmMlt9AQ7BD5Acnznycm3jvuem
EiE615MRrg6HsgMmeaRAjbATIQpFLhkB5wNw9NdwIoxAvyOVKjeID1OeyWKtryAp
fS9EbUXeXBmaGu9Zzl6ay0KSmDHVSGlNRlOKz+VIoccwyR3kO3EmVk+v0fFQg6WY
ySEIeKzZ4iYU/fLTGMQ/OSmwJs98+leW0sz8rCV7k8fIF85LmaP7JhTvgDwPm4Ew
mRbhtQNUREwJEl5gAbQ8Yb0l2FLUQIeYnabyjID2+yTnBast/Lby+Bs8xpJr3oFW
Pcjep/QmwZXtQ80VNFPXaGRoIzjnKn0HW1I4FMwkNDeeAXD/uVw8UrbG6xaVNEmz
Hm3bvyvowkMkFcIfYuMysXqJAu837AuYiazBpx7vs0nBhqKoYbCOh5zo3EaXPdzX
UdavW9qDtnBl1CG8Lqp5eEPGMU8DGkZptjzrrSttW6pOdaqssPYxMl8XRy4VnF5b
tl/YsRd8HfYudnlytiHrKWDfrGbhCoaRy15o1lXQmxyI5eCXF/yi3on+femiWPR0
yuQLjyNQ4n62VHbZQLOY1cpR4Bw+Rgva91a5SyGAWBkZhGbU8lPPGOj8f7xwpRFk
CngLgUrsqKVlRP2vCHQUfZURcwxZupVxvxLXZ1lx8EEQlD0VUKZxbV9vE7KuSPm1
OSdnLmFnBxH8YrG3peB6BL+0mN3TiUhBWe2tUnu4lztUp8AQ4cD0XvGp9xwFkMot
g7smcDMq2k2OomlOm9sJ4o9QBkCHiAdu9C8zsvCuklat6zs2GW7lcHMMFKpF1Rhn
M/BnOqCCVDwtRekNHpGAq+9WbMFVwB+HxMcP5ZmRW5FShhsIomBenNCKmHew1MlF
9Fx541FyH/G7MibN0zzFxW5u8d1U6wtZT/MbH9y+cNWoY5Yij6rMZTZDw798VYlL
Q4rWrDgoXFNlmd71Ue/FdbgvrzxzHWYbF5es2GcSfaGghyPvWEWO/K9N6wlvid4Z
D/OhDU0AUuI9YoWlxbMGDSa6E1HsD03Hk7avNvL2B6VXR2Ol0h6cceWGb5d0C2uD
5wzjfya4ubnZzCBFOrjHdY8yLzx2U3/nwxWl/KmhA5MSnztvEK/V+ol4d/7TATv/
JNLFtewo/3S1Sh2UhTPPdwZNrlsAxonfCn28IupoV9zZK8Mu1hMbCULXfT2BbDGK
U5CVCXbRu2urhin/5WjIn7qw3xsNur3CDMY6KIDlzucICq2A6bXJymiM5L6aB1kG
GuCAr/71Bn9LLIJv+63xwRDL1yRous5xM6fvwi56OpmWKK7m8AAEZlN5LUZZSuQq
ITgkoR5qt6UX6LEGrc3NSwvWVpLghJlTbUn9xd1Bcv0al7IRMb63VlGg+WY8g0gl
MHDcT5Kfyph+wewUIjM0G1pmtAa/tVmGY+we1uf8RQKGB6QSrroIUqcVJFnV3LdB
HhXtCy+YDo7jV6g5rS0KlpZ0EH/vOKjWBf1GiNAwurXsPybudl8lXvW5zFn5yaHE
45Z7Whm9Jeo+iJSn4BuDhWIRSoONfWKI/3RcunI6+6Y72Fhcd7xx3gJEcfAqHX4Y
0BqJ3q+J5wKMvbcvma1sdhtsgBlOqjDgGI3x+pTKvFpCBp+9wHLL1uXFFGdiajr6
3OleTZcyWF9RqeRvuzm0WztRdavko34qW15pXU2BgrlG8iM0dBYd8FE95V0lD0f9
z2V1ek4v7Ox9gZN+2zftNr4RV9aDza4pi6KShts8LN45PpeSj9jtGlOXxcPm99w0
7Fvq03fHjpv6qM9BVzcPqTlg4zkd4GpyDnGl2D0SEeU/G0vGHWnAJhtgZg0KbjLT
xrUVB1I7EHU4KV0Divj1xxMPMj0N3Y9N2vBnSK8GfpHq2LESYR8Saoq6SE/Ni9V2
iyrQaz42H5KPKnZ768HJ/UlfkHi5o9006A05EiOwxYU+to/qYncizqud7aDm5NlP
FvPiL1uimMJwFKmOxrMX9Qc6jYlRJ5HLwDEO0bjzocUiXCfWLf98QVWYoe4s8xf3
5nqSTWgg3uchenzHyKqEf1ii/I5Th4/l/wtyZe0R9HLFVhZ2B4FUt7DozZrsL/jx
VwqNhzPZwcSlnUfxYzz/kIxU4dI/L/javlHr+qcgoeCIUqMGwudFgNw+w+qbz5l2
+f5aKF5xIWoHOizygBi8OR0u10QgORraDXL+Wbj1aXQagRy7Hg9WlAcvZSGYslHA
Rn59N0CmSVfN3pVaTBoB/JxG9OrbdaI9PQGCFEUHa3NYyiQYFshQ+EZa7cSyK/wy
mida/dO3+5+ExhotaReEnBEoAM0bZSZTx7/D3ND5MTErM6YWQU+j1AOwA9z736vs
5RxaBvHZ8ULIZsWRx7s+exZUAXYM9BvjvMAdgFRKMDhWSZWfW81F3/9efvW99vZ3
ZjdlvUuhTawHjTM61idIZn3QS3ff1ZDJRNYktdC1BN2ttPcFRX6ryq8FP00WzSk0
k5Uyv7N/+F+vsSfwXhMqWfaB2oRThZmM67tbyRqE99I9p+qkLaMejCDdFxmtIZwx
0HOxZdJTuvK5in7wgQ2WBjYvzMZqypxFEYywB3GRKc2/lhu8f7c1eCgA4Zng5KcH
p1CjNSZ6KOshB3QB+Od7UPkID/eZRMpypE92m/MMKXvCYMsUDKMJZwjcZFM4zPpu
ZFEVrKI4wfJQLzNMUg1+Ulg02izjfNlW3Xyu/jnAusit4l9DkVQwJYTF4IaEJFFC
ogaj5GU+/byQJ8TZbhgVnYdS6c4+oizJAHUYDkBSktcFIbNokskjvSqAX+NCIh2D
noktF+3rG6RVa6A4MohjwZStEQE5iGq+649c7FZkZmAY8Rq6w7U16WocnOfqZCsB
ZO9GhD3Mo4oamjTGalFeSyZZ4naksfmA0KAP1UdpiB8XVku0oeC9sUMdIlwussbk
Ruc+bWgdY2LAsnDulFRFNI4C+n3iH49DWod8x6tWfGXpRsgPxomLRX6H6vXd5ETJ
hn8jicf1vLzak6Z5cRodPgePsqCNDutQX2UcX66WxRP8kWO8dM3eB5MuIxbwXS/C
thkj/+xq2Oy2WBm+eu8qAckVYMdfQAAZAzD5b9Jl2V+PwGTqXCbTxclxzIFTpU/z
3Fffd/WRes3OWjbWnjI7VgObjQHhx8mM882FS2pMZoi3U6ASqMZQEj4SFZGvKbyZ
oNwNTiV+s1i6Y4ub2IxzN+5O2ZorwcSRd39NQS0HoaYWhOz1YtTr+Njxia748bcW
3ZL8uWhb6ubqYTJdZJxmyNlwLbCiRkMje8j2057X4x7S2P8PxfN0OZGl7SFwLzTd
29BUiBbYKLL3AKGGg43R3QWUc7SHteE9TtXaBgrbTFPHPIiBDYy8uQhWShrNP1Bc
dAuZQZ6/rTQoQSOdiWqvmLwbTRV+1jGK3ncvq/cmUOItY3YCaaabRpDA0Pe8V72/

//pragma protect end_data_block
//pragma protect digest_block
plKHKibFWXmt+GBw8l2bB2R4S7o=
//pragma protect end_digest_block
//pragma protect end_protected
