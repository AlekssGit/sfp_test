// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3sjL1uWLKuRQsE851yVnaEmjdaAuvg29LqgdA15JWgAaw9ZIGHsau5U5OX+Vu5v0
vH677VR9m4lL9aq1JIbV2hL1jFtlZRHgquwg2kc429qlAyfgTgxEk6qPAe2n9SI4
lcnp0JZfPK144ESl5Muf+lv0ZwKty1bIfjtbwoHzuEjJ5UpydCGYwA==
//pragma protect end_key_block
//pragma protect digest_block
Y1Q3QiGLXPyzt8vrcwFEG/YyUnQ=
//pragma protect end_digest_block
//pragma protect data_block
eHlxyrYhGl22pHMphKJ0+5j8yJ8AXibd7gvjbYf5SAChM/6Mg4Lxe2NDX1dDnStb
/TEfF9huzqZ4sWR/EoLH24iOP9uLsh0Zmd3XSdWIsuTRY3EMcPA7SbdzSFxOI6A2
Lo2Lg39hrLxzt02L3P7XBC1o/0jyqWWFEfv5GQv93rJwOUA1KS6gwLa6S9OhKY0K
SInuy+yAd9D3mOFJQ4hZ/jRA1CuZYP5WYGzpqAtDVY6sTU+6qbY4eRndkfadDdaV
RxKoEQkfItCOaobVp+ZrpS0dxKbXKe24aLxG4LzrGtn+TfZ0c12vuudqdtZfyPzh
bYqkP4xRmkfv4fXm3y+FV6/p1RQQ+jVMpkMb4tOQSdrUpQnWM4DxbKp4uZfWV9u7
cAr+Z73jJbRpyJ5iFz4uOCCtjL4cldQl45P2wZdUmFGYiTHLLQ9bfUp/Ax/pHtdC
MVuE4OMg0SCuCivQlSWbSvNbZ4zj59YD9uhsOs1HBec6Bg8wyFrOSJjVmN6YlFKv
wOd1ZkcFHlvMIxW3QGsYBPArTCLLUFmHFTtge1NgSG8S0mZrHK6PB5K/PJB3C9Lm
1jrDFE6ErRH2FJk/owXnrhBBJnQzO7HEkmpZe7nnR2xXDlg7XUu/31YjEMKxGC4o
meRHXwk8QS27tkhQLge+gXFAclM02Feu7OCtaIc4bJYfgHlU2g8e4T/90ykxv4wb
mDMNUx4o/L3A8oKlxaB+LaUxlg5f/boOyrhrhnJb1KZJy8As1mOOEAVDnAUHJ2hL
f8J5O0YkUMVhEg1M3Vr2lUTRdVZmm/gkuSnwhqlV1xZbm1tX8MkfSys+mVZ5i1v4
OttXjVLqM7JtlR0FZy5GDKo5HGpZxjWC/Cb2B4HKXD9RuI8pA+BOskk8aeFYYEwo
fRnNKlMsjvCChhBdWd1p9lsbAuVrj0QStLCm1Ynp6jFc7ZG3Mo6GgiGv9fvfem6f
Q+LVQM9AORHcddNUYuaGjYq0+y9K8mg6cpSIyjVLe5wygM2fQH0Um+7+SqYq5NX5
Bc1WT0VIevhxbeOS/Z5wmzbGdJsj45IPVWUViKqt78+RaScFdrG6goxC3Qev0s25
Ksq3OKoz3JWb7lZpisFz0iTuA6RhIT3UFmguyowkByn8rVjyxdk9IM/V0o1qHjQt
VpC2jHQqFTugMQCbymGFOaLGthq+m/KsxwwBhDCrHHrNw6szxP/P2f4MPpAIkhvn
WGu79rtJGcet2F0R1j2iOxC2PwE+lb/6+TkjQNhkmjiwh95jUlon6FRSDu9pZ8I8
iWZVyZFaw1K+KXsnz1QIkIg9hXh+uzJ30F+d4Mr8wrJWapPQb18/fcnniWLOfl9q
aeP6J2292HmOSOEHFTJDU26mWPOKKl4WcIASoZVvH2nuEue47RVIb6v7rTNIkH+v
etBt0k3yiI7um/p3vkAMvQ1qfJNx7CdVX9ZwgjS6btfEBmDpqghDFEiJ+u51tiRZ
E+0sC24gueh4b+/I0xbgRJc01oVn/MA/LMuIHopsPkBZkLkjoapAOz8sziBDywJ9
o1WoJSgmaM88bLNyB86vWxJ9lVtqzC8YEjwDSKtiRf2SP6CD+7JtOXU0M4gOSFxz
oA5oas7d3koRwEfEUNGN1YV1pphF6MJdfitlUbwMKeRX43/MoWQe1hEYYw4YVW0L
pSoc1OmkYt2arfSvWupCWTbWc5y7Xm9e1c4pR3HJ9dKXM0SiHzKqAJWI9hVJED0m
rebdRIG49KNSNMP2EY8IefZF9eYklwjcxxIT+W9l1nnohmVPlQa7/JHPSE4VJNmN
+C5NuO75M/FeFQtCAjw2L59Sxjvz6f3H0wCRjNlXw31aHqn2A53hHhhv+hNkPrQS
ZZdWirujIl3QQwkO6Q2cq5CpxUv7wgjQCBxiJZHUdW6nyG8PHiZgzocVQodt5m1U
eMHb1IgHS+3xxYAD4FwPBFx+rOYstW68tUIeNKfjtrGsARC0hf7+vB7qgKV3ehmi
UZKNs7He2c74/chcB4PNZHkIOmZXglEnxSUcyEhMlGdCVmjMEVy4/l2YcogUxc/N
Pkx+pT9Pwzlz+IiK4ln8QlwSvze5Q70U3Wsz5X1cP+8L+PF8T0QBT0p5iQpiTz8c
hgvie1StKShF6PhjGmXLW5Jje3VQrSxcNdIZRqZngq7vS7FzNfH/s9OcsWytpNYn
FH839OFXpDHQSccfUFgjrO4281+GlhLzDaf01tpbmlmHHefzee0DoxkN+voIxfCB
7ow2IWwpbDhn1B0naL3kIznM2B37GZlvQ4Lj/RjiRNcVq/u+bMz3A2JzpftREBpw
21vWxV/egDMzcktUb4incukBqtCxGWafNVcuIpniM77YLpGtLLp47LmzzoF6dKjH
+CrkkNKreWu/VBuXRnkmrt3xyknLtUUxH6V49I1ILA3D3GHv/yYnMYnp91KR7T1t
yucYYbzC10duux9/Vtf4CS1G/FowmncRnbDBt/vE17JfGtySvfoIVRiIW75YqWCt
bmP1xFCp3+yK5k+m4d1IP4ox/NBEot8ABfQ7T90g5RhwIzh2nrMZ8ASaSxImYGlG
MTxx4XjOqTkcLwNB9f3UsO377cfDOuatzPcO3Nhyxb6kg/xuedM4bZ8DCTkYDRIZ
P4uhQuvFJMadcruEOW7pDrsX74qn7tK+fjrP6ni3JSTjr+Nm+9EEsJW1Yju56Wrx
Z0xb5rm9itUCtxyviuoAUCoth+3SugR5PJQFNCk6UsO2Nb3FF0py8WD+3EpITsbO
CJnozRx+NOMBfK2lO59R8CYYGpVOGjE5v93CxE82JQFyWsOFNVgfVEjatLBKyZ57
6rszP70vBzeuMGQiX8TawDbxzR8Z90fn8hH3jTkmujgFhev0FQsvGE6W1yLHpjgz
+f6VTt36HhcFnFdlPIr9YISvgZ8HXu/kA6jrkywlwa1isvUGW5d3kIBF85r0xXMp
7ffoxOqACZ70G26lTAZlVgcd6AafjCVvLQG16xtztJKxEcRcwY0lanr69E0VuKnN
FpAjddQJ2l3UNkBvZ/NjDJ8VUx8158krd6BBVj9PmqIjcvSLIabjRBIbzR8U9IUX
rDj6XVKIteLLHFyiREHgV0P1em7FbALuon7jaHrxIrQLNFScmZVQz68sv9OjOP1E
xsCS3JL8ZcaSr4qdKseWXy9SGB+J8eIfKQfuTGjizAkZWlXKd8q/5WiKUCEMeHS7
I0V5CeNbTXdSB+wGDSx1NyjP1WV9iXdev2GNal8Yakh/LuZbQ8DtCqcX/l90n/z3
WPZBBD1IQmQAHq0s8UT+SZf3xpbtjyM6Tmu+CHktB37DAP7bW3ZR2fh4PQYNLfWE
afSyg3G1KRiqyIy9/mklzcN0jIYpT9bmRDbNuNZQCjg6eONnDFSmeJBQp8L541nF
b1XwuV9+hNrlaBHxBQwNDJ2M2aPaHkOAP95WgEV7jrIMfUxnkesdHqfst2ehfLXo
+2FeNzvkh4GDIbwAs+K0nA4riwt2smde2XW/Ipk4SXjVSZjWahVpMXYzXd6Zy0ff
6lvMMB9EafgPXYRuY0QAg4IfP6uRrMauZ8g1m44w47O/0lPTXHfIfNfSbSKvVRin
Pa3NyWUyZmYJo3WTWkwfUtP2bKEGz9XtFl+YirwD1ed1Z50T2XchDDKsd0xkgwIk
6Pk4FVct4WWlazP6to+Pt/5HKue7PiCMsZONOKZSSNY6RGeuzzegAygbPsY9J+HH
BuwsO9dPugG4/BX6tGj1GWsgBHsLOXmoNkPHLDx52lAoiuay6DY1EmDWMEvOcF5q
PiDfairzs4uLHJNd0HVuo3M8gY0Ir/OL16Puf+KEgMobNxCUDsdSfSOEkBvV47Zo
7AoqknUPW5N+ris5Ms37a0daGtR0adyfpoVdimte1YoV2Cev1efIpTPQJBaht9eA
0yy0sn0jSYBd0v1DVtCM2fikBc7EhJ5FFRW1XWHj43EnwgxU5fuN+qSCCfAwWUvg
EB4+q5QlfC73oUxS/PFCmOtPDC7L2V+uuT2ufCcEKHg35s+kpfDRqxE63Xsx1kZa
pGaaEkAO61dX/UKhgO6RSHQFzYPNoL4HAPXOCH5x+Bm4k8BMmWMOkHCsbRXTpKlr
mMI77MahVNjjJbb2JEWSSrUkaIJ73IHIwaNl0od+vCh4kzvQox/jp+cfq65USdj9
5pUucgJnNvNJNkpp+6FVSHm5ZIe7zV9Jfefh+dGETIU7Z0LwifXFWHFtLH6xr2eq
oG+oYVz0pgyZGjdiNCBYb+Evn35t5m071RoRXBOYT2ywbAE/IjB3ocaDVg4ScPDp
u4T5QEezqc+5fGnFbpwIzP+9iN8SHC/2mRChLzoyPWVz/Fneg7X5Xret+tS/p++j
SL+h8Imi2nWos1DcrDdK/s2w5Sj1y43dRoDY9oUhGCdcpy6uriMIV8Wk6SO1KSAW
q0l02SXICygzYFL8y5+a+JgkToi1wH6Y9KtnmaQti/BGKZLpljjWbjl6LaQvkROl
bEJrx2qlS+KObboI1uGFCkbB/0MTgjIG1k1Nepq2JpPuir1kp/e/a659l6HacPbY
1xTDbzWE9QetCisJ9tFuG+LmVcDGYG3O2OfjRBxVj+r8t9yAwulbmKZQeoFFOxgy
5iZSr+WYKGbKNxq0duoadNN2Io7qHb4+y0Tg0O3JnSFTGyRNX+RF+sKU1SDw0gcm
jrgcf6Z6NDrHpehWSn4JdgcNC6cePLqc19QALmI6MqAA0CJeWNZuc6utVQY3c+e1
K2bzNjrvVyvKZOOFJQA1yS3j3jyPb/j1MKqLKdvuyWl5jz6daG0mbIoAyFkVVfI8
jk1xSWK21BTTwjhWPZyszoioxb9QJmob+pKwlQuDXVb6eFgTScpl4h0QuaCWUScQ
42pxWfzZUwmgggDFU2bQB7VIotc+M+QUVwD7ma3vwpWlNoelfAWaaRfBp3B9REfc
Zn3OI/DunOYUsP1X5RTR+yMCewIbn1G+8Bc5htXYlOFZPwUaVKLrCgaAeQNM5sDF
C44vZEZ8Eq9H/LpJmod04Ca8ozGhefFLKMrsgbuqvnPrPtiN7+FEuWEwKiTq/p5R
bC4Vwq/p6+5Nq1Bbcr1aNNpNk73Nya0bFEzYgrzVxghqXOGLhDxa8Jcsf5GwqDTz
si9yY0TjZ/iSI2e4loi1NGlXKOBqwLMUz3eJrJnR2wYzML/2eAK5EGKNbeC/A2PQ
DWtLu+BswoQA8B6zj53at+QnK4CM9eOuJ/VdWWswKE9qm7Yz4nM7zd8lmzKmSe6F
Rq8SM5eAZi0Ns/KiDXFnyTq9QrdcrEjgcQ7CXZybqS565/pEOtHiFrFpypx+y8Kn
xAcreeaRbIa2vh9gPZaxiTLiLLAn4pLLVgHc8rg5nwFhE/qjmFaapTMfbK5FZAlC
LaYrbJefi+btFPi7EpHTkYarY1r7k7Xy9ReT2+57cAbnR7ZrZJ/JwexerYo+9tly
xSwpC2W3EvBbCI8ThV+1Orwwuiee52LEka9VHu8kEhqMlfK2+rJMhRo11NWdQexN
yqznKMBJC0UO01PAazUbRc+J4KwU5leDt9drv1AbBUOgVaIroKZDWINvIvgUF6nc
jgYnpGcCFYf8kvKdFhUXwzZexfD8aZaYlzSnF/uo76MHsPTJ60GGTqEqdlg9zre0
V5198+KC5nCy8ILUgLxjmlTDQm+OzC2MHbIt0435RoCTutdAv65z4jnaoMP5kbQw
rVJucDw3WMYL+Xlgmu1sxU8Lr5V6f1lwRy0JBa38gw/zi2BwxbHLi/y4wOQU7EBI
zs5piDsy0JzIywMyXfG0JgPL9lPuEt8Cjo2ZR4MZzSPzekd/tTrwWwpDuyIoCiWu
G0V3v169SWpnKxIE8SQz/oMJw7kmraAtbuYCU9f02f8EEfSFnhLYU0GhWKjhUGN9
cwxo4+K0Tlqd62l9byctXKz9wGZe5dbVhyPT7QgrHl7tsMzrnOOctKj8DtKR+BaY
jZ0xnX+c9sV0f8JMWfuBeJoMEYuersa2NtvdG5/Wj/J4iQyopOs+5BBlowAF7MKC
r+YOjdK4J5f5Q7+n6SbLAyDR+6NiE35Y+PxHxF6OgJNNcS8ulGasm9cYmEObB7Ec
yiEh6m+0bKnxfnv0xiwt57bVNJ3lVP1qt4zJJBd29MX5spBC9eWaB5QD56FpjxR7
bs8RAy9gd5NbPpBLDJoNUVyMjPPN0u3SrktJ4tjIYvB3JguBXDFqAOaeRGXjd4uK
sc95SHuQkzOw5ZBkpr34O+Gh8WoeR8OZkBo5PgSfkBvkz82/ARscF6tJUdInap3L
sV91wNFxOuq+6gwE17x+EplLEHnDY3o2m05O51ge/IbrTVVwZNLGdw85QDicl0Wv
4T0B/lYTh9ZDvEdKp+maVTVTegZWs2iqodtKJC2b4JMrSRhiE3m3wScJxuADpaIz
wQbRx+20C5ijw5flDD7nfd9boZTb9rnfkMMj6a8J9JUhmY5xGDj3vbAfYyNTJmT5
ijWJn8u26ws9Gm3Vv5Yk1hO2jslRzw8dHgD/0Kj7x3/6FSSE8nHuR7eXRsrxV9X/
0zgp5UVEcRgyNI0pJpnAEKr+oWuOYG+XBGm8l8kvhkAuUlRHSkiB+mSpGBl0+SRi
aWHUfkz9fNP6i0LbTvk6uPb0ORPv6PxRk3JNJmCSf5S0JN1NyXIjnU/bpn+zjxjT
TvoOtV7tCmIwaU3aDTqf00228jjpBOKhW779HmQePoaEwYsvvE8VwgNqTNGNcelg
UEtYh//1l5J8yyQwE5KD/HbTYFOtLHh/AbvZ0kl3l/XEt+XO8WYjJi1X/1nK2ZsP
ovqAtWNXiBEZICvPz1cSlh3sXuxbpsuJZg2ZpnHmPH8W++WtWS+/FHqaqUWSYVEF
cD9kSNniatNeIyneypZXVKwrcDK8JJy9mUdUDt0zWyBsVxkpLqPTkXHvtSIImUOX
2ZnISpmehQMDUxuseLZHmBsxylOANOIYK8bKgR966Ws58axB9VqAG1c67D2VKWng
TYuIUvcxXMhnlV/CK8Z3tY5r+LAQtzUmH7wdgLQ10289yXblDeVQRo0XRiUy3x6P
6GLXerhthDw7TGvCSeA5I98xMBYsV5H/lmDOgi4lUTMyWLVX5xbtbqhis1RGm0tS
FZIbvbLpYk2T5ktV+87fyvTcbNtW8L0YiDHmiZSKFQwec6n/ozD0iOanFA8kc7Gn
nbsiOYawE/X6wgwKRJfCZGmer5YtyxbCBNoxM1Lf+00gA9Mx9Xz8VBhVihOw3eMg
8I/8LT+oeSsAICzqLg8Zbd+dqlzJokrGEs0KjHV0ndyqR12RcSthW4YCyQLllRWJ
+dYm1vKZ30OVW/sFNPUgvlEUt3nf21l5DxAeHQmCd0B6cpwQieSYCqd3htItv5ae
zEnR0OpynfeC1VGj6d8F3yeSZ3MpOOo6TA2131Oy1XE2IHTOBsc6x1k8Bs1fFz9d
n7KAeFs5msEf+8O4MWz1vegrh7GRDCWJd6ZC5v1lXAOnET+NqzeNF6DhimuajRdA
AIg7H51DKzrMewjrfZCtzg+FDDdoMrwxIduEfhowA3IkIoqJ6ap4NczKOwNI1dHP
0NvXhJsXjVpn7pCroxuLJWSpMuylGmkkqY7jZmtR+/HoxkPIECZhYX+RhVcPAf/a
3O4TQ36ZXXIE2oOTsKZnyKgOReIthQ3GNndPby1i+FUZseWfjMG5nZdrw5PiOrcJ
rR+brhwgGEvwN0HAUICz30QFGcL8duLuR/ihkyGPLyYCYHzMyNeaTNJWHVGXdhb9
It3/QVbF5wCQ4hCXJGPx8ICqeYeqGi8ENH6EUPGa3CSBeSHaRCEnXJrhUet8Dhhh
0gOWLtYQWSEg5jOj5OvAmirvOy6pGNgYX2gYroa8CPlr/SV3eZm5kgzqURfXBbKH
meMajHRo1A11kOqDC2oZt3kVFptTexDTj/wj7E0gWrE7zAA5A0x5ZSH1yYWS44Rb
vvRdEVbuuR2D1Cszj3UH8/F6678wSxYPNG6OTLeDuVAQ5IOfjPbpBQDTOBb3il0t
R5aqfoUPimGmVxA9gKvKN5PvkS4GG7Th2QoMBDgtPZd2p5Qf5nPsRiB33Px04qyj
bdVNOfmAIhEpDHLJJw/Jp+3d8uKtn2wV7UEr9N45jW3zrb18R5KvMX5iU4iV0gfK
qmG/UCBQhlpATmSrLCPoBlA35o+tsHASpmiwo/mPWxTmP5Bjn+NsBvR9TKlbOCmz
H2TlJNRoqJKUfQEunG+WUqh7fnq1NDty04lRSzB6aVefPzRvHpvmnjWRCUPgZG6o
Cy6ZN/sEfEAZ76KrawkHVEonzqqtAZtdqSQzufgL2eApYpz0yyTfmKgC9Tt9Ko47
kkltXpJw3SUEQfwP16K5nZyZWvkOZudaTwHYEYEyeNFSk5Luu779WIGv9vtINn5m
HJ2RE5XR0RqPsMazHcEhM8lwUkb4bORW/kthnz7HvLVjzcHOybmCmFPkMVeyZ1XM
4sOz4jON6ESyAb4a9oGPWsWV1naHd80NvT+j+xtQKBRLjfqki+XKQ6K9FYLRpmjx
ETlVlpcL6T7+2dOJdyZDzKlglnRftuzxNV/Vc7CAFY8qFIcqJQeo+4lJbydQsi9Z
iVUzPa+jQQ87KTKwIe9D5td+pV0SaHhPNTuQU9F+WurhAfS0tjvi4ho8x6z5X2Ar
4XicUjBeOSF0gg3RxjD4P3bOuVIbg7mVuws4T7tuY3UWVJtlEnLdL30rxeP85FBn
FbeKqU0KLF2JW65eouQP1myvjHTraUbQh4i9WuD2XAy2TGFMQmT4QWlTlWbGX9Um
eKcLqbMgBBeLuaOEbDsja9F/n0p9rEfIzFK7WLSV8W+65SiqeJMtA/4HOKinMuiO
XXQqpLio7FgttFqoa6CzzfFRlRFc7SHcMMZKKKQN7W49JOgNlXfPVxPV5XbtfktL
paqByxC0xRCBgO6I78uQMw7V1y2IF4IaCeRoYRhIogOykuWvM+Ya3YknlFKSFd2/
7l9liZ5Gplz0QCtsIAeHJztXGsM2nfxQD0DAuw1ZS7KEiymnveBg6ukRppoC7yFe
EX2rjE4aYUjQ6PPVwVPyhSXhtyvy4BK7ShmzTw/TrXPpM1N5i7d8majVIIrVumjf
DqyXKlgNCBfpgc7sn68m1QtfIF/chzVkdD0ik9nBVoPvIinjTZQm/tXxqawnbNfA
xbEt9Lvuf64JDkzqC7H4WCmBcolDNTgI7S5KXlK/8fXbT10xg8pKn4PU3fWv7GyF
LCSZZnqZgbeT1ILC+CUal7UOId9ZEMC1kY/nvLWAu0+vMDIYClB94LUcxfjgxRcN
5wsktor+xkOHSup944z8x1Z+gAxnuVh28MNejp6M/xHGYogAUu/MXyQTje73x6vt
e4VYI872Q7enziUg6N5zinQpD08ZUwMEc5PxrGPboA0uMrmaF4q3vCpYqXgKQ1mB
1HxQJJiaWxHhWLXOmKLEHA8S+IMXJaYFk3E3T936eyPIlDIT+DTh1cJctL2WiFgu
09EuS8XU+VKiEFjUq8Ng0Tqzig7DijBIgc0VsbDGODyat02bp6b23Fu+01Y4qiRe
bSPAhnrCtihWYuQUyyjmhecT2+E4dasYDmasv7CUMHaNOVa3OAI95YXkNxPpmbZ+
Kdebph1uIxYVVs69RIsMYeVTB8WaZdf8R7of60jMG4GE4Eb7WuYrsKjJOu0FP7Kb
G96TjfvYUNj51TTtJNg2Va3X9kQ4eMgFgG9+GIZ669GzWpwTUcE3swug0fRwNui5
weyaffloEPZpKAWXYcD6O2jys8qeWaoSNWoktPZCNvGme0QRppsKRowDprwWz2Hm
q+77fDGfpy3Fue1+1q37iOBi2etV0t9LuhURAARNxwgHWy4WKDfU1UuoUSEonKNp
OtKkWoDhzHhYGfG51IltT7FvSTmikf+zAihiucKCIQPwTUrasxwgPOITOOPH6kDh
YnvojVhbvctYkB7SUraD+XzEzPWT0YsTsmfHVaewdBncMgl4fb5rvePETzOD73AD
4WmcSbvy+bpLy9wMpcDbOBPu/b/osFseCNjdVEZrl9MilzR487D2fFT8WiRBdYQf
owLT27fQuk759Bk0jeyFB14cEJ8CFcTwrjXtcSRYlHyuDv8bj2k+/SKZUL7ZA4OV
sfd1D3qA6NJ1ayipOsP9cRhNFJPcewgoi112NksWxu7BTnbfUuNbRidL1rcoyWD7
sRajuhNNoaqBDS6G9w7qkHG73Qz7lTTcgfyId+rP75mW2aGxRyfVD5JZnrVPXmnT
Vd61mUDx1BjxGpXTeKS/uU0npu4fmdRejFwH88HV/HMooQaITQdSykrc9X8kMvpd
vcXmjmGhDSLWA7XaPTbq1g9B8r6PT3g9XQCyeKLx/Uz+tRDQ+RRkCqM2KymuQtwx
ibkKrehWjySXFZQrCc3p1LjA/LO+smZ9L2qAjkyd2lucZmH3TeYgRlhfa2r3labL
vWGN2qLFMaA64dOYi+ZCMHSlSrOiVdDXfrIfBy3e1cD3/70hkdWs2265gsxjqEas
FgtCqCjtRFnHOqxJK2apX5yL8fgRAF7X3ve1ynhvSCoSQmdxMOVID7aCWd+k2crQ
T0iL9KGadfZwbVKRioPtZTkPrNonyeVyXl1QuiRlYgrqiPu5PobGoT4OCv1/GaI2
9HuuaPSiZjoz5R+bcGF3sObhFAx/sb4Oww7mZL+zuoKq8lVq9K5zelNXTbV18WLe
27vThdD2LtJ7+efkxD8c7nJTvHIgbL2vmYTYFSop7pXySGEp03D1TGI3owiZUZuP
j7G0xrHTp+Cm4ttG//S3yyFFVtqWQPqYxXf18QDxByBJVOk4ictdGxpI+cLSsGBw
67XQyFeNkIeYZtgnDBt3Oi3CVehF9AtYp+y8iqfqnkiKMibdCBudhbpogOpQUyjI
dq3rpGcjoqzNbn4fCbctemAm/Xg+XWLW/soeYeFZO2ttQFmquZCYQW/+T/j2Ja5s
8EdJf6jevb+JcjeLI+VXjWduC3IBDawFOd/8pXoCqSzdK5K7sGCrgw6jtYCRnDEx
ZalPSKm9LMHJC98w8RdvyNfBjx+FEISjZcqYtdo9WSxb8HwRfvgVz4/AoUt3zqtn
sxRX/QmvSnFw8dQJgMbbixI/GiXpGPcTK9CMjl7A4INlev4usbd2LhdJPl4m1Nzk
jWQbSb+7fYsMcpmcsmWqwiZxIhT72Q5BNWnpv20EDDK/F4ujO3DRUJVk3BpO10AD
PzxQk61HLRxrDYkvAssqMmiuBDtkM+xiFZvWESszJqjM/kQOkw6e65BngWnllir7
6Th6Y7xtM7tAMzh/lrmzEpTrNCSG2wl2HVT83kILPKL+Xfr0tXQsM4QlhCaU/ORN
IATX1haeldplW6/QKbWmpnEJ7jNwXpkUaTihsi5zDzAkX46PkjO3uchxAqUV/ntm
dXyAFZpSPpgZ1zZ7ceLp20iX5tFKbrwI5gS/NrZJ1drOryjHC5Z+eu+M+Ct2htke
6OCc4liwn9B9SSN/uiLMw911QdBND0Xk6bow8AlsAWWNZOamsGQieS42mK6DoFhT
cTEzxO931x9wsSzQNJ4/WTlwRJReYYoVUU7VL47zWuJEmkB6nZja6iQdKK8E5/pZ
4TNVHFFiSbJROhp39UpFWNw1Jzk1ebPffaVYzgRmlS38XbOoqs8hUdXssSKhQ1Fr
7CdJV2/V4KfLiAVTegMxHLUzKniXBdT0WTFzDQoRCdMHBHkkw5OgUDR9dVHR1Dxh
Rgt5FJpbexBqxyVp2+JeWI1KVoU4iAfryF5cl35K36IXUbSvPOhAqhW2MLIozxg8
ltWJQMr2NZVEh+oHAWiuq6c3hhQtBhKMx/uTJrrQ4Od/qGIRm9z9W9HM7ODRqB9e
bXomhPuuaGBH4Xcd+ClpAVvFQVsO3pWDEnCsXbESfbA69WMJiXqHPN2LzFLgzVsz
NBLqH3rmVXLlVp76ARAICvbCYibXwvsXCaX0I0jZCtdbNeojUvTCuxttfGrRgw0F
hVeM/yVt+dXmt/z5uOWtuZzf11MRflCsQvmuv2p5zVPTdXd9UjmEOBpE2VqBwcFL
vziqV773NEtKGzCi2JKnEops8c+usBzBNnjFuHTmn07aPt30xkruGw4uzDM2RnMK
4nPokHraItK8G5ycO2CIOOxhx2ttAiUL6RdpFrY3OyUabQVh1wYXPu/xdjDWs4qF
DhnX9THO+ggI1zqvdg8eHXFV+Jx7ShA6ucUwJNGS83vstSjLSou5KzIi+hNLaHoM
3z2WfoXev1c8vwdWCOHk8FEiKYRUkhDCF1HHTamxzsNg2VyXOFhUd/D/GB1iy8HI
z90pJ1m8Ct5YSFazCEYBLAxHCfErPqv6877Gf5fuwkCDj/tJ885vCE1rHP2WDwD/
W1L+tZDLRLL51f1T/WZxuMrcTQld2RxE6KifSXqK3akK+mkEl+L4BWRkU7welx/P

//pragma protect end_data_block
//pragma protect digest_block
cRuOfT5LyQN3rcKBSYqJAp39AaQ=
//pragma protect end_digest_block
//pragma protect end_protected
