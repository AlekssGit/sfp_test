`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
iIKrOc383QkS2yZjz6yYkuGThRZPl6jGD1Q/VySWJFUZmLXtWMxGFx58z2yzTcal
NDabB2s8ead8pQhFiarNKhV1GRZsZsS+OvhkaNqhSKfROhOVS0K19l8H+++BLiqt
JrcJ90jQZxYnMBIVG/Sl4nb5SzpvxALzJwQdEOMyYpY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2992), data_block
LRfGTleZAgol3w7piDrl5XCI9VQcy8br/wSMcgIYig/DpB0ropJz2YImrIW+FQL3
n9FXSBsnZZg9LnfSA5dp1/sSaZN7W35VvYFXwXccc9/yZkTRGRwJdQ/iZvSZ9mJ3
zzV3MznlNvn0FvHXjAw6W70qU25LBOyt/b2JEsME3D8tOeuwhDLo4IXVLbsW+7mU
a9y9NcxjeiyT0QeBSXow7xbsgo2BFsWPov8xdzvgn6P245W2N9jrrOibRugf5Dh4
l60sn9NgJDmg7zVECRPT9e11DA755pfl2aOsBgHBLUgVeb/gs1XFjrqK5NOv3ciw
fK8QVaqz0d4JpZUJjhRqUrvvq7f5f04po/GbaFrf6nYgLLMERCHnX8W9pG35vvCC
ITYT98kIQ+k9V5aJmSne4GKR+JEGwBBAfBNzZUkqqH9Y5NuuP7L7sfOLC9Zm9IeC
ffa8wJhqvxOiWomXMFtzclVb8dhpuQXSuFtT8xq9DV9/2w8XhRZjlbhDv6v8gqkb
cZCoFnmvW9LWNgqX0WJHbJPUZ2eCbXEuAVTvHB0mY4FyNoWpJK4z8ZmGlapJjYil
1Q9KL8qlWo64ewd1QF3+75VZbardat7X812bvzeN8c6mRvz163IabkR0boYj4JS9
cnwLldB/+0LV0tSE1sQeXpPrXXshfY5o1uFW5kTlaiW9DmVIuwT1u1Vl0Bz5pgip
FkdbCuCTtoAZB9bHdqHkuuu+BtcHk5yjAXLRYMMDlrbZxvrEcHTd9iFXeO0n7vPD
s1Hum6LXNuC5eyVmoxzMRTY2G9CYqc9nylE4JkOmWFFMMefCdL7Nt5HrxWqCbXL5
qu8xyznhJmKbYstRAcPoge9vdAvlA5K4Mcb4LARd/UoLkfCGadvumPsxo3On79eA
R4U4SHdbaPZYLvz7kuTkYAwTUVSaMwS5hNu8Py9AwKknHzRFhyEOQUGYukjeIkah
VjZDtHmVc7e1CoJ59xlItRW1qoQeOS+O8ZVHjRPSIFIfiLZ9HXg3tBBqSL4qTB/Z
JteZOPmQGAmDofVRu9unNb90wAC7dEIuJIC+Eq47FBG2Y2y39Qwwf2uf0E3SHR4e
P/UQNd7RB5IBGUEbMfIr7Yiic626H7E5GfYa0X1embxITgIcy0HWvJoPJpGfep+g
dd2nlaH30rdAREczxnccVSMBAQ5Av1UzYxH7Rraf1RexjifWn8WBF/HjpZHEwQ1y
U17baOGMyUBLWcyyt4/lNiUSU7v3kJDmtU/0r8O9VYTcCSqAt+ijN8luAtvQ88uk
LfZ3Bzt2fZca2o5OlmGByYk1ra7hid8Sx39oxNburEseavqg7Z/Jf/DNWx/nygdi
FGFO9PHhMWFeZECI0o/rItGgvUNvHXtSmIcdAjSlEgHLzdnNf/zDYbzJX9TkuB8l
v9Is8xxSb4CGqoFO5VBtJk8IPMT92M37AtH5beFuyNQnJgMKRRyQUyjetH+UaY0T
U51GLMkXSnQRg+RjQLaSzmpIPUcqaQZKb0Em0n2oWYypiJ+3rxkeIjfXfNhPOjh9
Qd2DAnx9FDJ0qNHVne4hn/qadjMEmGTRpJt+LWWUFYm6SDHmDgH8Jgy2YOFm4x2e
6Wrn9y1fVg1PQmASe6oZNR60jcUYKNifVoi2d+R7FPp7oekLc3iCwUviRVzQmzIu
w3tCJb+FCudbf2xGOmKOSneXqQGRvF4eW9/7xA9Vl92mx1CdH0gNDRjqOEc9/8RS
DJB8eRs9rHlbtgmjGeuYWsIuUe7XUfeFIn551+luAPFy83YTxf+Ku5J9HsIlcc0k
Wm0JjlUHUBRLvFYqrQltsD2fuVwt07Z6oX2XUBLbxIX8BfyOkqEZyEBGc6dNQr6E
yTCbiVyk+h/X4ynvzpxc9hUIcQyY52vZQ/sK2JcYhP9gqQAhZt1XjOVwSpbuz/IG
8QQGuAePcuZjAdyVyku+ct0StONIO8pm25d6A7+sAtsZoocHGHTI68dUbK5Vzitw
T+efHAhFtrF+196TRuopAx1FPIVZdSkYsY4+i91zpA/rw+Q2fnGec00EZp+j/9RQ
vKLWfdiATg4RJ9rnwvS2/BzG3n2yxT5k9Q4Hi3u/E+ZtDw6bUGsiTBLmKshYuDyK
R+cuBTUSfpbBf0ENSX6BQRXw7NfF2mBsZf+TBDqyVNhQLsfTLiqrIaLjo+HQkJva
E3PsmJcHY2zYm/zFE0H54MXI71ln4HVxKmouD+Zo1ekTICrSFXp/Q6EHSxS9mGzc
votLc3MQj+betzran/luMY8MOiCZqIHhEC4PTXhG3H3EjqCXoj5i38uYUZ1iMegn
JxzO4vWK+GAsAezm4zs1CVbsyJv/xrHw1OQf08nNPNThy2KdzG3ENmLThpYiEq0Y
q4PRlHeOqEJS4G+TLXXmGCLueK3jFVMQ1waD61Br7ae1Zx82gi8ymqOHAxFXad0g
UARmLk3YZEVcGU6ly91b9TwpJTIpfHdPHml6l/KF/X9C5LtrwL7F5mmNhyf1tY2s
nxuRym9y1jOk0hIx15R14anEZ9Pzr7BqtY6N137NoqgGDsNdW53GUjnezvHi40Ut
cFa86ddRfO7xmdoOfJ/jVLG0uc7nhz23bJb3MwgQOJ/bJtH545EstkLRhLusAepE
xE5+qtj7IaFEYTSE+z5ymlcd57ONpzzkHXBWVdAacW7z1eVqL69Cyae05QU1Fe6/
8MP8QWEoc+wf22RtImJfFGMmFLS4DLJTU7xeHWzpZTBj67/Kr1v765YGN0NiFiYR
ekLT0yzfWCUZnI0R+CIMqWo7QsWtzXgdkJmFHFYLOt1AcP+2WJtWe8Lo4v8dNN9t
pzxcyjwWVYYtk2yJhOiXaJMkdM4URZTSsQfLrHVCCIfolAwOrau+ZkcbybdIuPfd
2RL407DoVSjqh8dgpHOQq2aLitLCpsQ61+Ss33LYqACJkQlyqeXDqXOlmW1OXrbY
I5EGVjuaPbDk/+Iu8qtpNSNNk1iQQO/ll5VuByxXu5inEHA1rm817JziUai6uQCI
DSMjSpfNPD7ZNLM5XzXvPV8eLCuHs6hWy4tHR/B308fSGQ8dqT8GRPKLH2eADwTa
fp5uZxwR36LrgYEc8X43pLoUq0cV1RKL9Im9A5jV1rFU3tk1Uc4Rm9uZWs1p0XSA
C3zp5Tfhg25icPFsPU/pDABEs52rGPUZwPhDNTAJYb5hVOBVzAHQV9C9ltKvt2L1
tctkBprQ4ejpYVwYxg5NEjAp1ljSNAOaFPPQPO000Jv4dsqSRAMYpJbYUaJhB7ue
5ZaDAQKcWJ/w61FBeU+gD4JlifJ1g2WtGjsijQ0fSGh23DYN1WWCLFsbUrPWmQeW
aJtMpepFlDhL7ORm90oRF8t5doYIuc4HRqwBJLak/KHjUQu+ArhB7RW8eZyrjETB
/Fs19kTpRWEy8nBYergguQaSbjllod8PWncp0SiQgB4bs0Q1hyjnwP/Ke76ARM9J
M+M5EQ7l3t+I8Ho9jHkK81VA7o1UAZIzr44nxNKSCz3BDLaIV+Uoyw51662CxGPW
5hwRIjEAJfrst/bY4ZqjJzodUeGmH+b1MQ3NqvM0pRiY5eDKqxfNEKtFxlkGhQVq
p3gNuYqxlgizTzZuntkPgsv0lFEsjyFgyVEJJL5saAuNNuZgRsTifJVw78seoDnx
TSxuInk/QMR61tS5zFX7nevoOdKgNC1vr5PFS/43sb8Z6ZGdQw+yizJqsruEEKdh
jC2z0yQCQmrGK62hXIRwzCr+9JPlqL9T6iLmaV/mT4vSp3rJKj0CRyBDzo7nXhO1
zD+LV2stf6Ktfbv/yj6+lSJa2QDXBUW5TsW+0NrmMIHZa0VeL750mE3VuF0H0/D/
MI+RtByb6jZntiwiFSyN06c51bFN3are5vfmoiw+MlZj0tbOU5xcA6B+lpM/eoMS
7XrChjcZt+giluoXQsF93++sfyiBXRkv9p80kVhsgtCmIivQYCd/bGlNPYnUjwqQ
nDtiHbhs0FX4ph2C90KxzQ==
`pragma protect end_protected
