`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
p1hjKaquAQQaPagphZRNCPUBO08icj9KdWwXFObDDV+/X8kpWQ2OmFbC/esKJU1i
7cV2cFJJ3Ci2nA0LwciL3Op3WgyKqoc5o9RAu/e2QWEi/T61frwkB/YN35dktM2D
MbxiTVUSzYF5ZMI8tunftTjVKBt3ypj82vocuukqxaI=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 9344), data_block
uJvcCeZwXJA0QlxzrcineVQfgKvtO2RE+wHDyx2FGVsFOqLwIQHUM3o/d9uIqGuL
vf1FZy4VXPJgv+EvmOAluPJfGLBCZEJFSNQgxQtIvD2p2QkY8yBRQKNT+7ACEIWw
B/Qhhf6AHRjEsopdueQ1+p//0F8rucT2FQ2uxknWVplpMUE6iWu8jA1whC59qvsY
zTFTSA1I1N0W5IYHdbTY0aoIb98c5F108JyJUM1t90GDsSpYDzap2++17bbXthmx
BaHtvyRSkyQNoUQdZm+Qf8oPhCpvgmHnuisTbPzWmbts87RmsTf3/dpD2qrrs1J1
ZxTjpRWpiTbKBMLXGWXgKWkyuNm8Wsu7n9KgBzjQAZH67meXgHJR4bblU6X9KcXa
a6e8YeG3UTkeBI/ygb9ZLRVIxkWbbG+oeiG/CPxWe/XFmoFBmYcpqz2o5hzlHwJh
vbCiIcaU/WP1cMotfomfoBILXmsQTaEeFrrfRzmsD7IzhUM4/5ntEKcaIhuDT9fo
xuVvJSoOZo/hGmkLVMCB543XhzcQDQWg8Wy41nBui+fUqIXn7w1YnX/PQZ4Bd9/B
d3f9XVROe10CbFyZFqcwF4eQ8+9LSpuNfixzyV9BDCZ6vcF25neXyOBsyN/EC8C4
xx+wDuqINBt4Y2c/j7ORuJJYvQqQxnJ/JiEUKPmmbVodzRqBqLMrXxorgmM1DRQZ
xDBGaNNt0cxW/c2C8i7tlYcI6Eo59aqtXkPCKsa1ldI9T3sZWgTilWAIxDjV6vUM
pR/vvbOHd8T6pC/0tQ8RPyCyAYgbM5llintJkS+ZoWXP+wYfaCdMhiI2ZEAbeO7I
pPp3/r4/D4laWx84jwJ19t0uCWLVtCJuXkfsDmAaY+p+VRHW0EOwPHbwYecudDKq
BV1B/yWW1liB2UbDke2ivSb7/zxZjB2U7n7NAWSJtfnYh9+OVPxbZJni2xeLrZ0T
0dZtn4mqhylzEbDaWx9zWV8Ea+XY4layM49+SAkI3z0h32p4WGcERygLK+eYfyyc
IcSHGBKNJCYnGivYHbfrEH05vJZ5XcameRRfsybK1ZV3JXL09WS8Pn2/RnTNJYr7
/j5duyYjDprZQT0a/KTJghXZXe/5+8S5hrZmWrtZMVe/jVNh8kyxQtE3gRtwqEXa
1FGyYtEdhM56zpy7+qgY6RCOtUjvXKwaf58jNUC0Gk2mWu/GaMpztEq9ZZZDPXnY
ijkArfdGxoWZGzA+4WxIfuf02t/GyZoGpX/3pbVE2OM63P1KY6ea2x60H8/t88ZQ
gH83Ft8h2tKAeuj5YAWz8+mIl4fH5tU6NrGhLPYrt8fqryrskCddPMnfpe7xhnMJ
3CHXdBz8/RcioxhUL9/3caZOCh/uXLB4kAvXEdKXO5bjLvQLuZZNYHzF0YZfpkt0
cHLOZkaFw8HHgobEc/6eshfQ957WVX9WxPPz8Q+LbdmEukcxepPLlhj+NqgemRp+
jIAPMdtR7V5ntXuPIrz/uXcBWC1MIycUSkYLixMUmH6lpQ3ER3Voz+T1vW/GZtJR
i9m2cO08fRGFOtEEf5zqbr7DKee4DzmMMSk/EHnJiDLmrqXGlq8Soih1QTKcTXM4
/rFdeySR2RTSb2d3c0Vr6EQ6uTVnP4kO+TIhCTIE+isUlfRit7WbkaAjUs4oOuZj
73EBqJW20Qx4dpcj0Z+rHzqUhzzi1ooGDpMKWl1FF8sZgNX0w6UguebQ5D+Mgt/P
xTL+CzdwVajT6FY925WO34WYt2QuvFW8tjAIYMvdptfT3AxGCEdvp/1zQqFFZJ1l
0MD0zxJMG4BbvIIr9EKI0EMN46HsI0e67LLs10V4mIZnnxnIWUTvXZxk2bfaPK9p
PFFSkHrFGxMlcnU+sHRYQjs3HDZ1UT9PuupamJNNiriBUb/tmSldFELcx+QMJIv1
9JgIG3KV1tqce2AZn+0I8MbIcY/vTN7qoMN8ZeRIsZ0cGqwRaXPs9yUT3dGqujsM
ahlsWSW+nG3hyeiabUjzSSnTp94Da3m9DXVkdfRs8KEhYwNO07ALUQs7Yo+M3fEg
ySGnQ/Lx/VNkrqjz/7NgrdkuyFPj8ytK3a5Mcvmhi7ZaY4XVlYoaFOvS+8CAq1bv
gY6FePHnDRl7g1w9jTX53UnXiv2SKrlVxwHkDU3IuT/86QDoN3EPL6mUuZixOXNq
mT3HFThtpagiI8phmN3dG6SlSPI7uVtYxPvtamzXmKSLQR8TtKfUIXu1F2J64qzD
dLNcsNs7m7LlFvPBSCleuzbB3n9+FWgfQsYHwZR5XBcLzkyAVEMZW10cxuwo7F1n
Yq8oaGVAzS27JHQY9FL6cyXnzdPsd06EFqfAqHpX2RNYNW3c5nJ/9NLBbcBHfz8Q
sdR/Spj5vtRq/XHnPWu8yEDkZwsEoVJ6Hj6+Vwd7HvCCh8Q0s5xXHbIJylGsu3N4
4EgYyUas6Jj67jC7y9TvTiT56KHT0Jj9jB7qH+MqPy2JXPOIIWTzo7kq8zRKXzut
60R5S55YevF/ApJsD96x+a2HXtqpmeRH2XLYM7W/YzqhQezIqCeQXxwh0uAntXW7
LTelmdWk4Fe8Hk3iX/LG5lZfVs/UC8Zuq9SxUnxhNV7rZpgOC9FGRbXIWBnKlio3
SE7mHE5W87Mad2FXqUeyT6g/oA8t3JNlHZHuIa9xjxW3ATZbBpAlzG/44otapAi1
Y2Kgv8sQp8Sl3/BwNJEorQVoUdnSDkRjgDEaCZc1xF0svgYTufifVsK5wGBCwdzK
tnqdv6DSZtjaLn3RJvDAOKxZ14Op11ez3I88RXr5tsuMv4M1H+y66utucwQjD2C3
BpM8TV0RrSYiV94inZmtYjGpZWN+E5sTf4EH8hzEKh0SPICkNbUxRhr7AFNFYJO1
kucov/czDJmbzWiKfzVgX6I9f097tGW7AjZKtLoeSIMSTl8Mm8vSubZc8kV7oyNs
tZC7xVMXUGUUFK3KLjesvDGKe8yd5l9Ze+zS4sjDkOCqKs+rWzSwzL00F4X9REus
T/1F/mZQBw23Lyf6tu0gRt9PUREWhZLDwceDHwzXzwhi9Tuton2FJRt5R1vu5rWI
zwwuME59ukswRu1DE+6T+mXk3XMDTCGjzZZtZIPwv2NrmqXReIKSaIPwTaEsnMt5
TVeBfk7cew1s2BXKC32IyyD88r03pyXLDQf/pBvzguqjFvLEKZweoQ7YGUTgyigp
rZ1lkr12jNoz/BPayQYtMTtRLyNye64Csqg+vsQF9YAa2fbScZL2DfkpF2CXda0U
HuJRYDE/K/2+pOTVePw/+9w6oyO42AUUyFvTP3kfFP+NtmhwDPaqTwW67bGbXCHa
M+EnWn2jjamqKHchA4sqGdfrC3K5e07xqnJTnZOHr2r4k2mNXLSzvBNFFSPlqIR6
sBm8J35k/jrfjMwJfeo31fFwLEC+i/nxoRuV78F4NAnvNNng/5TRL9tJItRjZTbY
kXlhx6RkdQ+mYCzMAP3J8QcLuzP7tTR0WJKOV19mwyYGaZjjzEQBTSKocDj42nG3
QYojCoXmulb6tN7zbU1NjE1a0xvN+CyOI8n14nXQVHOIabMs768tY8SFHbUZYqbK
S66kSzm32xjLlg5R3UGmoHbbF+rTL7k+IrWwsFLEsvx1yzPycKkk+NC1FuvIwnrF
qEv4yGAG0IvrfywYcQhAqsHa/E5BeK8FROS5cQd5SqifkaiWrTM+y6L3/ghfZFxO
iMdLPdRAVGxvebxgvKh2XZl1qvrn3uG64Hs6+yXHeY+ZBRWpjlj8V6/DCL/6te8q
uZsLSGYmrue3WGOxM7AHoHeTGgI49yX1YcY9RAYtifRXVnvlno+oEZ4f9lwOv72X
3/5ZQITPAvcEmfpIldoVjhE/OzpquhZ5y5JqtDZOoUjV/s257Xl4mAb+PyUketW8
tzkGzGy6QJMvBfcTpe8X6y7X+/QzPxcDcbJfO7OQ0uPaf06bjgdOsoG6mKno9ZJO
JNGLfx4YkL30qET7J2Fj9Khns20RjO1CkKbZteEJvKLjQKuN5Y5Dt00P11IKbp0C
b7vh9Lq+smCqhFo1hvI90VMjHY9uDVT09/N79iujaC2lo0p9hEL4c606xGPvz1bR
QPqY+GDZGpdv/OMSOZ7/bnv87S/yEtfHxgXpjUU4PhzUlTCTtxL9MgT7n9koPo7E
P18DsY5atKBJ9zNWJAJZsVOncXn5JpOjPJk2i+nrcBpmbzKPOXKq9uC7UrKPJrQB
zNvFz5j2BjORG0z+7APP2gzk5tabt/ogH1A7otTRzhYKjQimI9yV3cx+mLeyggkA
H5/l04lNzsesV5Cyy8y6GdCAfpSsr2Ms8tTqa3cAFJgtxTKpyYXy8ELkUjlo13/E
YM6HIz2v7HhHKMjEVH0MY4514bELFFyM0ZaamDA7UpUHCxqvQwvE7GWVvU3bLj1U
UJEnd+Y0Eh/8y5PPZrzt3R8LOt8H73TN7qBIYj4Y5bofCpFy2hq2Fuvsdnmmv8bo
Q1M0iJEca5vmArniZkbHA057QwYH2I5UXWyGKvGLMdpfzPKsUiz22Y+sTgSaQTRs
Yrj3k7/zd0mIrrYgm3FB8U08fjULleFGsj/gNfI9gOdLkZHoazyxXGPXmy08RyiY
rSbIcIbHyfPrigK5T0iUqTaA4KJRj4/0hYAcLxs5RTOeY6cXiCp5k3G4ikD+xeoM
rNwkT8URR2M8vPn/Hw4pbHNN1kPmubilrzmsrzIep8ISDEvX97HA8Sx0lmvQ5xOj
w1ws1ZmsKUwTcHPIptp0pW/UzLbEvu8kXNQe180mTSDlOXyjHweOLXFJZlaYFNrJ
KTsFdcpKpEgikN1f2tC8UaRn4lppWOZABw9PCFnSyYbiYq3oFolvbEvcPRrgP824
U4Uy+mzG5YKGZy9HpVXss8ndoCJ94u6J80cAR2ds31vVannq/kw123ajmE9pUMUl
EnEI0CbcdynMiyyr57bLmGA8HOJTOjbK7IL+nYQH6A8YwO8hdu/03YGNitOiSk9e
eqOYcy8ljD/qFIw9iowdwmg1hRiAJjf6CI2po1NQaw6rGw5EEZdtws00xgP/WnAZ
dlXuGDYVX+wlo/KupvnEkDFE10X21pO+nY43pQu0ZFr+VsQpaGNhijPhkVtDjcZg
uYru4CA9/oq8+tfI7Q/fhelFVOdskQdi+ENxF5mJdSondjuAlQcf7gmN9DoCVjfT
ub/mkWn9aF2vLavWVn6UocK9VL/+x8M9Br3SowmeQ7O0/iLJ4aP0kPik2pZt8zUT
L+NpMD34rAstQWVRMxT7oTV+R6YNLlLSHpScEX18T+gOVXl1P7IPBGHlC0ejdOVA
Wow+YgH4V2/eUUfD3EUDQoE+QIAdMPhf1QKU4PeXcAXpLucwJUzqFFwzkOmFBkBl
dOlj4XV+qqeitTJH5KFl1mq4TfMA4TLbhNDK0bQaABBaeOqTIurZbiKaI4t4WG60
jKUSzzOJyDbNQ/C/+82ZsjkqyXqqWq3lY8uvvSngWbBIOwBFBPtpIKdV4koiZVAU
5L1S2rzLrosT4LoOuew5J6LKDmmyWfWwNwygNsGKuXqhmmoM+IHVSs80Dkfs2wUW
21G2yylZxqZTX3dqpGdQ13aw/tqXG55ysxTUDSDoGmCm0ds8NvFcPjFEeIjx3LTo
cfPbS5tiAyMFLGUs4Lijcrrubo1+hB/eNzzieGsLOvhjZTipzg6vk2HPjcNDxmxf
kbx7Q7o7mmIb+qoprRZR61pS0GAlZdf3m05vgUGbeRkgHQGowXPevvBFSe4ScdC/
tEBvgo3Qg/bPI8/HPZCmRQhRtg/uqeFvpMTKVpPTCPBnph9fmJWptmy5ayQjexxr
XdzrBSs/57PixQpBxFFjp1bwMxf2SW/LEmVUMBKcTGCu9rvF57BQY/WSGEuuoM7p
WHYUPHGDFc0sokDg6uWaclz5g0Yz4VD8qH4IFIO+ykx3BDoYT90mdpRl9Dl0AZjy
FbR1y9xQRXDX+2ftvJt5rJqjokd7eQbsWCct2KUdp+QubcqDTilS6xy7Y6n+6iwB
vUoLbYQmo4D3+KPhA5oO0YuAaWVqDUQ8GsFODLLOzA+qPeY7PnqaBGqXI8tnb/PS
KtvdGZVFPNUX3apxDusYuTUckELKuh5ee/FMyTLvJ5XvWycJO4BA8wgFCkvvx3UG
VzG/EqEwYAfJOvGcD3JRDTlCgB6O6BY2TGECaocyFMZkrIhFMcyj6zifKabfZbDI
0UUtOIBnRwBYaxTU/orABoCQNsatOHBOy0FU3jdH0MoQaSFCbwQDWtqqZJEhm708
nqQKKY+8na3a2LARKy+WZIt1l//tcun6fDbm/QsW8auLOJ+BhVcHxOJd5vSs8jg4
TPn6s9QJTv2S8Dd6cYFFqtezaphVYn2qukItlMcefSQl8BSCK1UlGSjzzNObGizh
obi/ynoZGHJUx0bVfvehJCi6VxOWyotEXOqRZFqImOt/R4193Ajq73qJRhp/wq5N
5TS/xDKpyUe+wuspj0QwJoOhZolpLHuG96jSUNcGAdAq8QEIIq5IdEBO5sKMt9Ia
buYYpsIwyaEHVDYjb2wBisTi/3qrg9RkvnuOMtlLoZqAiw7lNqWbw+WJG0p73kt3
BD5NX/hnA5BBu8HrjqfUpVO/rVebw1nyK1LZNR8ESM8ZWZqAJkHtSRUk8iU8zpbD
RC6X6RXZ9hvuV5qfNdggiemsyMIISn+WsoZFb2B/0Mu1fmVuZuwW0/eyL1RTn5dX
fM93PyH8CWnCCI7TOBs1ZjfQ+vEa1XQIV3GJD23n/uYVCU1+vYMUPb3OZ01JpXvK
jpM6hsf5oaUkvCwf/s0bvLyOsUF2pEpVu4OSYoncbLMICg65yHsARDxtuthJ6ZEy
5Ghlby0IuQ+8T747VXPMzQDrI7RKINFk5B9usZpo25h8UKUAWJPB3K0/r3Nmg8Sg
DIQEYzHsXYixM7nbzYNy7evaZ3TF3d04DofoGG6o78jLsBaI5WvaHm3a+Z45YoEZ
OoEbe7xOet6WMOxeU13A4oclbdaO/Z7PX2aiRcUSh4bd3YEgpPAKV0NS/T2GBhbS
GBx3GS36JmSEiFXNfemAp2/u16F/XruoMxOiWq6/Nxe+bimooxpAH/lp4jtrkI8d
XqUyJsrw2rg6fEMZq9NVEXskrmw7eTih7uiU22EHWgnhBJER/xGhEWjiIT24xkty
rNTYe5Li0VM7Zc6E2ULTeeTU+gTkBaGyKu1kKJk9d9ScHscZxJ8CoRzyG4gf6EWw
npp5yASpQoX3G8gs8keFWOe7/fZdZHiFZn0eEdETVJKtaVAeThNEh9gBOQ/9932Q
iKP5qXbxNXJuqP2YMiUVLri3n/xJ9x35KzdOsl2ZXDC2SQTvun4A+F77oNF+BNyl
jH/7JZDiDyBhFWNMsCCQeQTN9tUGAPEyMYTH6iCngYGBlPD26CDas42UHGRvHRBW
rYJNIwAjV1ImpJBCOs8tdZ6xDIwkQKAr7f+jDGaVg8Yr2m4tIdUkBJrpK2XR6y2T
ozlAJvMkgvS2DTqqX32SrrauUFUP53WzzaAfb38FCkw9tuhPwHE/jHe5EPaIa3TY
4HpJQXtPfzaJVmT5STZ9fy9y93AEM4RicNhckkGplVwSC+SIQISJ7XM4D/7GT47i
of9bipk+c9jFyLs0Dgy+7o9N2OUcKEraG+/Ik+EkQthSXSWhbGfzueHXb6Iv/zq7
+3WvnHOl+zr/5bXjfh3LdHvhO0kjg2Dnx63Gjx9HC6tZBQVuGMeUiBz9gO1sqSQk
HUJ5ZG8FQmr22Qt8y3kBslDVHy4tP9yH5kOHTY7A93+dIsAi4cAW3xYC1N2mf+N+
WvJyfA11cQLrNXOXiUKyaZSFpMJmXvCqfkSBWXCDYAXmdqjq55qIK44eezHp/7bz
wy3SsgX8kxG9ZWH/mvZvEsO0XiqP+p8iBypgMf00uD4EiYvk+HxAGqf6Y3382l1l
Df2m9COCv+Z9AEt8QK6oWKwa0OL3ZgYP4OnroIO/t2k2hVrHUq7al3RWApX9Dt6H
aTb+YTNTAp4tEoNUeJcmv12w5gyUyeBmPgdUaMp3gEjuUBLZLQ7CdBQqfizgAP15
bqQz1uvD7MjdLuFbQNTXo9w6gXwzY33yU0oq589m2k4l7j+EvLCQAS7VPVOoiNID
J9vFu2kK6VTnAbeBqfHInRpWnS6xUNwtxynRMMLnI8b0Q/mXAsbKXWS75TPcPagh
nuL3xQ5fWXvdcJCxJk0kSTQ3K4H5R7Qjp48IidTEBDuaYaiV16N66kYCys4eawX6
KVDCfLAHliSjMjtzQqIT/6A2dPTTgfLg9WOqJfKzH0ITAW24R0usnpup42OHVEwR
k98TxZERskI3K/Sja+voItMw4Uak8MPhszddx3qaSgu/kGAcbbA/Vjeitfcmwb40
lBsDCqE2U6A+Z/KK8GxXlTtKNLW52siH0wV/cN60JWcHwOhSt9bLGZZtwSnyJgfm
f3QmTnJMngd9vC0qHaDaK9R1oeOZhOoHFzVPm5xut3wdpa7cSQMmqYcuPvECoJQg
I7jycAhfKw+FAIEFIAnF3alCrjwb4Y68HJIA2OedxepT2stKw7hhZHDqu9F16hFI
MNEljThOGUoju24yNITUG/soGLBV3RAcJwAv/08JtUGZQmcowxQjDDmc+E2iM0B8
j/Dwq+zRqJdXHHZRnJtpplnB10Jld8qYGyoxoQXlKMCHENofAR/YrKyZmLqzYEBg
9xIRzZYh143jmSoidswBS8LawlasakbVTlBxg6skM69uuBYCTNZ1Ry8JOi3G2Ruj
6DULhcmXIDAkz2ACiIx43e6K/qHeCBowCO60lAQjUByiGQb2RytElVMb3r7Hvj7w
6pQSsF8RDpxVK0IyFYuZ6gS5foJ5t0hcfR5vUDTmw2FICVAVm32o8zSzR835ROkP
Q+fU1AJa+u0rlOqRvsNcFigHiuFC+CKuDX8LgfVVpddQT2q0FZGMVSg4wx+JW08R
XKknrnSuc8h2o/yu6wudplL04IyUH52mGmhAZlZ9lVRb7qjdqwi0djl2o8UCAZSk
hO3drP/IEv/23U/JzEpMOIk1/Loq7n1i2ct6d3chU9EZGXBZsNmNNiTHglMNBIrO
FypaCU3St4Gdih2f6S7m6PXyt2YL9BBM+lU0lEkAlGUcofk9rRLVsMzDLJOEpwY2
lOTTzjSlULs1umfWzPSUCJu8AqKSwQ0RqxGjRxISLa7BfUXxFJzwZBFvOaOtcCxM
QCCCwmrIsRXBfp9Q9oizQ2YwHL7YhenmC9zflVGXQuf++jkwzYLPlo+YqLNVDSFh
rxsiC2RWQCmPrePs8n7EsuQaQU+eqPOmoO9qZuFV27h+KlyWYAr+8O8PPcu5t6GL
qUKBdbxwz6pLa10LlmHrXHYexLzZ9ncqR8LJlR3WjMaX+y4s87IfJzOzOaveYoPe
YNraR7Cso+JrLNQZiNp7xNw3y0vEw9m9wvKdYo+4io02wjhNZ6vw/OLfrZxTi+Ea
Sdp7iLM14Sq8A1kX7ahTXDzM2oLe6gnjd/KsAR8WWchOPtszn/JPE3vd48WvPG7/
MGT/mIs8qtIx0jVXypMf5deDC9vQCITmOoHkcJ47yT1u2crR1QRCqolj9s5rzNkF
vYIxSZVKNVy3NM4PsvE+5+63qVZmZjpU+b0Fne6AHI127YxpHoYXhiG+QNiOP+sa
QQ3glqUxU9h8i4ohmmaiu2aZZBZHztAR5QvM0OaYYCh/3EUt+KGQB7SVp79VYoOZ
UmELrSgbLn7B+QkN8a3hlo0mrt0f6nFHVNMvlUXJXFQeJJeOSbrQU7WBzyDv3Dl+
17KbHj87TAgfMNJPQWtwG0Owqqv9EgKptcROpRwUt21MoGysjogNJfBrlHs2u3CU
PfJCh38lDTuTqNIGwRn2FqiNSIOjwiKd2pZ0Ahu57k7Js9JoJ3/PNcGwe8C0Od+M
jaPQQryzS6TwfPrTrEaMrJAHCy9dXFOyn8oq1zSYx6Cnt/zBBaJ5YgsqtqidC2E2
YU0mWhsRDvNe1TKUZnk8do2I3DGSVYB6qr3PORVjVAxPV1CdRK8ppmWFjv99CX3g
NXsWHYpEso/CZ84voqpE7qoQhYJ4GYrRgOzjV1Ot6UpNgdTrjcZ1lw5tVXz4gHY7
p8N3BrTTljUPP5veymgaOeNfUkujDqXsBORbTjN1ChsucgzQnFibEbXEfI4lCBFt
U7VmqqjKH1GCdX6iyZWX8vhpmE2OD8skiXx/ZW1EFl1xEUdsTR07Npy8biEzYcRL
8OY5J9k9YGhdSIauATeDDKTU71Lo58FVO+f9pBCd9k61aN7Efm7LJgkjzuijeqLA
C5Vraj2Q/WnIS0Q2L+3AFEdm36rHEZHz8rzaydairaCBPPfFDygQ5IxJv1O7Oof9
ZDedQVE1jweMJF76kjFPPwKfqmhvVQC8I3eIMKER9c93sl3JhoR5Hmf8fSuHdmqC
AL7+MpKle2juHZu50hX1FU9W8zsU5i4BipDsv0J5VK4pEygvKGTkHHbc0JdU30+g
s3Ix4gwqMmHM3Xgu7rjTKWAg/acaV5wLClYzkc4ojf8RvuRDtpL2pj3dgiuffAhQ
bd+f+D9tGmUc2UBAzebd3x+ehaD7YWjbsIeItbgGx0oBitA64gJHd7Y/qTDAqWkc
ZL3rriGyZvduM+tDRmtYrWgzE0edLH020WpS1AcmvuIkOFAk0PGdzYz0njQIkeub
IFYrFH+rRFOZIYo4AUFtfQfqzXdeR3deAt+zcE4NTU0hO7LtA6trUshnNpSMCri7
iu63op/BEke4Qa1HiZGueuKe4LrElV+1nc6DvrSw5RjdbVdvEwrS9KUkrj+83/bg
bYrWHFjOmztXb69H3SVymm8WxnMCCDQYvTfPMau3GnQgMeKnx2HOnypWjPTd65l5
v5xNGO5C/RckuaFxkXtg7TIu1GySrtpJNpcWJ8LRTb/TLGtZCtVpMIaJPjNbwKch
rJ8JMInasyfBKepipp+TvjIhtpaxFWZ3IwWgDeX/JksaurAZVRDO4SxV0iH6duaM
80lDNwrK8/cJ1Kf+MIIVYXPZrYQFlcXBRd8B15h2wKHd9i4S6fF4UrcE+Oyz0J6v
fTncFz1CE7OOm6DjDRkhODZLd5llccN/JJXkCiJoYxNRatkS8QhhiRC81yctRIX1
pJpCJg8XmEY9XXZy2YjbL1aXdKhb1QcLt+pTnJpVxMPzv3woNN2wMT/erZBfxrSe
ffse3PGwyr8YbMEPoh3OcwJ3GpyEdNHe/wj4QhOiv6GF4nWZSluPZOmJxwMvLsjU
y3uiaTCtYFl3mqut7x+CuKeJGnb003Gah8p0zh2OojfGNJRjESuEQu+oTJ/fcdcd
I25Uxz8OWa575udvBSSPMi8NT2Hedy2E60B6NhfIJDNlO+1thUNXIv8knDo8LlPt
f9+VABbORxDkbv0PCYRfZfWP1fF9H1grTjNIBspdS9dvLRURCyrG7D1LGUEH7ZLk
JqolAAbNa5CME1UvSWCOFxpcFTe0dc3lhRdAoUSX5zVAG03SBl8l0xg57Qb0i+P5
VX29pSRQ3bpp34aoXu8cHtQVlBRbKe33QTHbBLlCuYCML51CNUWGCrV4ODJ1O/Gg
nZWsxu2puA+lTuDLGjfo7KB0SnG5pWOaTiLCNuHSF5mUYF4z6qqkfBwkyRYjpC3v
DoGzbW2wprc8yYscfFiR1lI4HADM2XuPKJmIDJZDUkkcBGtqlmRDCC5c1qLrXUmu
pe0c5w4pzAV+mNR+HD8gNUWKlFdMoWYW87PfUr0VHUPu5JPNK7IiQSZ0fD1GkxSg
NSA3XNOSuWp4E0TE00+i4qxJgJaPY2Pb01g5GkEuvw0Z3aZogJ0+4zMVNyc7dKaA
CA7N2r4Th6WZ3PbdNxkq0msZC0HbPFvNQb+nBDv/ZR3QOMWQ/QvS0gBGbHYkTOmg
bsq3miNlJtEY9q5FD0slstBQBC/xDzvfFTjcyLotfRQkxb8bFnglNsabhHhEHvBK
W2xw4gB8itzTwB4HWTN7yd3mrkhSpll7B7nZ8HXLSGRpSH5Uj66M4MeIjgfNHtRa
y8ENNTIPvn43XqIjcCf+6dwDg93r4wHoR7PIqKrshJDLv+eSIij3uZw2tfgLGrsw
K20KR0yg1CCNKkGtP5y199FEs1BNJu1Xw5T5AXps/rIOUjHsNdHx6X61lFKsp0Wk
uU48mXbp10nMHQs+u+NZY5+WcCYv+1kyb1DgSKTVCxidK3KzTEGbMaPnpHff71wl
irEFG1bWhXqxHzabu5QYlCpVXB5o3cf/L/F5XeG511eH/f1jJ0mH30euWwmTBtaN
23crB1HS+DAbHp9E1WoIer1Nlu962iL/BXs2xC8qDPmB6emjdHIw8XufNmkgygy+
m4mtsa5Y4E1BlFVj5jGzgoTSgm0PFXekUdPKRaXssev3UFqH6I3MR2lAFCsj3iC9
kbvsR43mDQsom5tTN+riiHmhYe+GRH0V6imzT8Btijs=
`pragma protect end_protected
