`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
YL4kKKJDUhI4hPdxG8Q2yg4alWVfq00MSZuGpm/R3yL1x80u/A2PkX6nHMMa7ae+
mwRIXVlTeWNWv1GCi11SrpW7+CPhcai6oqsyZEY8k9wPrmzxVCKdxwm5hRXts/8b
2BA2MaHl4lyFXZG/ZIvWcsp8zFtjgKxjgdJsNXReO1M=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6208), data_block
+jupAORsxvaLgiidsOYl1sr/9dLa9IEJNk2io7itCUpFEaMQ6BKDlMwnIFrnP/hB
YCIolrtn9ptKMBlsIPp8yMBOyjI2ZWCCKXzM7ekei6co1cqFhDzun1yrID5KzmBm
AoTGPNdg2t+XjEm1JHoFpA087mLBsOUafJ7LHkRgsa9If9GRlQSVeDIexFBiKgof
0Xu3ibyiY3pgshwHXBrTB9rR9418Luu6OPxALmQB5KcOA1bDl5oY0NHbVnf/seHH
/092WA/wa8FrTFGLf50r+VbZJASItf9Ku/9Xac9UA5GaHkbs1ZAejRoF8d7gzRc3
qFfLvPqhVXeIPzXvju5mNndMV9PquKY4FmTeL1aSBDLrx4GjrioO5sWQJ4r+jCbV
SIurAcJYRF0KG4vUHBRLff9jfW8jYGAO1CVgSx1z4Os1LAkZPk0Px5RqItbSA3c1
vAoU9B9C1520OqbhyYGd9qRm7a25Ii6CAcvIrOGe6fupT6sGMB7xe9canLPGEMdX
S4KWnN4kJEf5J2sIbx2KAaDRckVohGHsiOlnrZpIVvovvD/cpibTyKMlftfVuVeN
mY87JCoipXQBSe8cTPQ/O6jIT2ZhAEQoVdzyodsnAiwNYUjrmh2MN9KTWCdFlBHl
h+33jGZvYAnLdt2EhGpkQ2XiaPH/yjdj0S/xyXcb0nh5NZnHM9V5V/JBrnxmsikC
F8y21+V8o+KIU6aOUyG5ZH+HX1yhF5IYYumchA8cm704A/wFt7xG4EJ1O7foJy0n
w3R6NIR1DRS01bZX/CnZsl5W3OY4FwUxZJnMPEg/4NbSmxkqlojLqFk1F0gM2VlN
bXeWkMevIs9MDuBgjZT4i8SZ9pP30hZ8URAD+lhQTUbejrktnTo64o1L4hVwl/eh
H7cizRBOqgKJq8ftRoP7DIY3vObwYrsCADOnNIepxCoWDs6pKt1Y4CiXDnJxPJgD
AMq/LNqrVwnlWQr5QpSMaM/DJdUprw8kkJQhneHlIxLiN66MAzl2jz2g5R1Q+IIJ
wk9bmV6ENpBbuZIepBy7JwHlu4JG/C9aDZHZTKM+XFjLYQkS5xao3cHgUvw/vNnQ
a2LcRksdUqPBJLShICpOx+6FY4DTCn8b26ouAJyVHMbPJUgLoFPgMQsuLA1mGtu2
rFXUlmwd+FXtn4//qVMY4TSXB0UwX3QzqOoNksz6VTQKk2p+I9qQdL2F5SCS7IGP
+Ushwkf/qoWdfr9Z9UaDnoZq0qSAuocRn4pv2TUxaguiIfLVxQ+Z5ccjD+raU/vT
RgvmuFgYzluyKcNfbS/lQAuLEVaAnYkkLK8G7fiJLheOzpc3H8MyytOLe5+zi68y
fhKCUUytuHxtQ3WuozVF6DjD9AvOZhaFcR0oSk1MIbtShK00xGqK6d5p8cXAXpO9
PT8lyslJUGnBBhvPAxWC7hIQcpZ/RBHDkCgnhhZP91mvGsBU+6kLo9CoVyeUNgCP
cjaCNSCEhT0r/Kvgp+91USGVefapw/khsNSSyQQ9zPYESXX7jpLyfIYTMjd7Qfl1
Uv1XoqtMXFQbbn80Fy5z2lr3wHsnVwelHLGRDNpmJUPFkF+JUaMcnXj0w1PXhZLU
EcNJ5RyadFKBMQ9ENbbXMFgnfAAAL+CvX7XHB131Jde6YK8fyEQYkmIzrpa1WQtM
WCFi1kser3LN/tD5O1fRsZaGAJ6AKEhaXWvaWM5ByiA/0Qdy7e2PGgcWimwqvLGe
EuiZas/8xMJtkMtfck3FrXwQ6qe1Uj6ba0aEpxKR3fH2NponY6c9LvD9rD9R3iMS
40/UVTXGzEuECQfO6cu9tNgOsQNQcSZnN9nhyiOpn4tVoO0kq3l4FcG1ueYvCzxs
W3a8MPgW6HaQ4qyleeX62Wxd6aqtiDz1gSvhG7BFJKKQnqicY+0Yt9lCrVd/mfnV
XZ8fxs8st5WH1G7/KGt9aPpihaFX7gH0a1KafDrbMcVzFv+383BF8A4yOwN8FC1R
SNn/a7QplKdP0sqNFHxvyy8vznog3JDPQBNwvj3ZMkYJTXvFJGrrKpteM6oDv2fb
3lXaYnYLJbeUHWqZEfBgPmq0VYhJPaw8DIqQZLn6boOXcdA14Lrt+a1y/1ztSqwB
5RT8noy3rV1uDJyu8GEMivjB0xi/dkenjqpa97qFXcR+yQqWxCCVysuIlvQUYh0r
WOA5kixK5ucoh6R2lkSFrXQnyaqupOSeQQK+0Tbun9LX6uyUbTAWD9ixrkufAluz
R8y9Ec9it9osLj+B7cg0yGgl3fqCX9/C5lAcmL827YNK0JV+GTESi2g66IPXIx44
HlsUGy/WbeTdXf0Dmd/Pqmd5oGfPEgQ7/VkyzOVyFgs2IM92nKQ2b6+OdhvyZemz
pVPh17q+henA0sIHoM9v9FZXiFIyeOXwnZCeMooS3h/2MxAvEPETsqIKOl5fkq1r
mDCmZNuE3mdtOGkmlxkglsj+flIfbge6qgTwvuWqMSSKgYsPPhvjzinIUXxqEa7D
oPA/J2BNLAqpS8AlrYymljyCg9M045Ojdtl7gaTT50XZ+yi44RRbey/bmnTzgTwq
6Joo86AzsOfQ68sfHalYU4uZy6iMLGJXrl/vVNsnHsZD9c08io2iDa4cy6HiEDuV
Rm9B+anuZqcC/L/YjsAt/Ycx8G4oBdJOTItbAzkZnfEb7xjwu4OWj/su1IZO10Rf
USs5lqfGQdERTkn3kiaBilUQrr7ntI1W46rPjOixwL+vq2ERXYN7zmyqxR2WOHM3
bs5DQyLKZR7BnaXT6JgM7od2gjjq1uqePn2DvNETRZeA0lAEfaqggyG9Ifd/4ZCx
3/IZgI1/jbnJe70LeKkfZLf8GVsyDZgUdIWpITzxwAuuUs98JBQEZmzqfpssvECQ
R3xyvAgzmkjm4IdNf0zjetGwMJp/67Y6M61epB70KCXSKdpu9WTdgkJ3uv7Y5577
RfFXL6fYonwwkWh1N6Q9Rgv/1Q4/zfYPHHC2ErXb+s4IM0uPUDBGqU4FrBRE7x43
4CdNP6HDXFm8bo1/z3viLDWFL0JziZdFGsf/f6Qdf0oeuEpyWH1NOxnCbI7TFWqg
YbEXx9aHPDU/d/PwWP5S2rz7vjhb6VhC2Fh83/MJ8ETp+0moGXMUSeuIlz0dDhDj
L+e6OtdR/3rwNQ0kX1wl/sbSnrkZtv0xuMgr9G4B6OmUuCeducsuLPsPQSvLUIm5
M3CelzhcnknAq79omfG9ycx/UtISf1qGE+uv7CdkxLtyKzpeHxGI1kOmfQsXR1Bm
fatJOzk5AOP8OmRRgTV2fLOdMfKgAmdRMsg91+appHSMwuMHOzSTWK4VMHuhcUtd
EbLcVYkylO5WrtFLIaeUNBWHer7gd9Ca/2G81eCRJXtjdgx3bikqUMzS/0y8yk0A
snBqLeJREhF0jiymNqkgr08VMIIIWXvBzs3bKCBvhHAVv/VcWuSGWe9D7yPFjzQk
7LZuGm5M8soYHypkcwP/nGLtJUN8AQxWKfm/CfFwoafzQ84BULcXLIV6ytSHcDW2
rpNWF2j5eEV3ee0yLrpN8otWnDiCEJpDA/YOXyMIvpm60/3WJXvApSJp3Qlmu/I2
F4RD1SCWSnfz05mYTAh4wTlnESgwkL0kB+1hKXGcy5UJ9bGCBbtKRbGB2NUpbNLX
hv13ZSkRionu5oSCN81uTuP5uH0eiYhxkidw1mR/Kykdqt9OJACaW7ooGJlBaTu5
wlF5okIrw+zilhorKy+grNGwNIUUcDqc98HcCzQc/7GnJPtf1+guaZ6/UEyrhNwJ
9/FWRcDaZAoQfLxJLHKFv9D9zjjqomrMzzgEPB6yTIQNhd0IUAWFjHU7Dgn8slVJ
+Pu4KarmzBqVYPSm11QPCXG7WdmhCNaw9Lcr4wvC9LeOyA4YfmL2HSfYxTy+QVEu
Rc1MJz6SxMKgAllrfsTZ1RZ+NWeGwiU/MqViDiKoEPI7SAoo5bDzp/fIwpTd+TOn
MC9yHpGR1HSnyHA8j2ZCIX9C0bp4eB6TOlFgS1c0FS444yp+TUD50SgH/JQDF6IT
6FMBIBJT8UVz9UrG4Rm384HW1/oYR2MRUmwfBY3GTaM4YqhuqmYlU+qeGLNERECj
g4Zui0Gp0w1fJw7Vju+0FEFueaVEO94DlK9WGoj4gnF4QrBB7x7wpw8YB30y5rS/
9arbp88kr2LFl97MqpQ5yRDbqiu9SPg+67AaiS/nhgD5BYhMFSoNGVShXe4sbX0h
AXjPhJTWLgCjmztF9kbfBbWPs0EurIxCWrbWdl7yNJC29U6PRY4G0JMngcVMFKfe
gNVS2TbwmSWodLFdB+ZiTnHWNJU9N3R6dw9poY9bBco7ROMMz5gipsLI4ms9yMRU
gDS0DcwljWYXunK/sQJ+n7faLijpX70PCcnpY9t7ZKrS75vbvglJkEUKEMuOtM4d
FG9uPDLFMzViZJcxMYaAINBTRhfYO9SjGvWbDNxrbPJN+LneeGvfJ1QGSh+ljn0Z
ylTYpCNbuBDTntiiLHUQgfAnPTAj4UwA15xr/suD5gFJFMKiv65f1Mls8stmLwbT
GZxT4S6mESEoMMvWXaXxPA/qDLuXNqnlAH5wg/DOMm+2CR3QAcJUeZuVS8Kr2wcl
UcmbeSAAAUC9JKanogTbmjS4wbE0N4yEVQQxq6txskOXWZYnTKVD6GHBi69BPd8x
yLqQELG64k8cfgNr3l8zUfcceRIevs1UWWeWr7ufoeRy3zN4HkyptY2vuq2Idwgb
r+vIAomNk3Qc3kRtZnTVjU5ox8vLG42QUsXpVtCg1/XzSXCrhq5mrQ50Ka1eYC3h
WuiMTVQ/ynfvj9rTrv3ENTS9eG+XxGc8Pe9MhKhOM1URrRX3+x7mzQ53f0buAfKn
MbDC4Ii4nB/s+IGFllj+YxNQqEwVwa5YcgFGGWha6IHAeYo5fuVwqm70FaOIVSkY
yoHP9jzlCLRHM/clGMATo8yMi2sbzz2f1HnsHJQvaLz5Ovv7M5EpPrIYwyy1nmCG
zYlkb4lPhZSyeO1GrkVvLWLgvnFpiYEj3pSXHudPKredtRcWKeAazesodWBC5gQJ
bp5493L4I0jiCHZWbY99ytqsez6bqoqy8PAbaTHey3/y4YzTLf+l4RB+BKciJa8g
irDEzd8wTP+xqo+KZt8pP+4bVGwisbjgDRGxporjgDq/wd4HMBet5tqFyxAUuZn8
SUWLM0I3+0UknpwZfvbKgEVogDMP2Lb/zpVCauxP+5YeFiHh4+44o3ljddr8JCuJ
QfvRSoGwvhQyxiYYu8uz3t1arhorlXRIvc9Mw0On+iaGKf4yoQXLCbQbguMPomDC
ZCZJY1NHaXRTPwl56Rl8m45f//yqY3LbjRjFjrNjKcv1xiOzb9kZ1vhUdOKzFL2I
5NIQGICE0p9+IIf/oOQEv3unHf+ZsQ7ldHuH6pdNEz0IXxITKGRGP9wnUh6Q85vc
VR4teHUAunxlUyPYaMWSCN4Xsd6a/nqI0P9fOoXcswc1WAdClpQ8/bQK/SXa4IDm
9rdEGbcwq4zySUBGOOi/pjEiYK1Mn9hCKhgNThDJMtcpnr4injp2Z1tiL5uyskik
msDERcu0ja3W8OsEE0ik6iByGqIfeRK7fY2D6eikw7QqnXRVBRkrkxMq5QZVZRx4
hUnzQwMigts+/2kLDJAwQkC5yrsvWQn9Wqp8z5i7mJLkCFeuPGccQX13OGkOfNE9
CGDCc2/nslL5Y1FWJ5o4MyQ21yJsMfl6mTuo+Mc2QDaBncqhzn7hHI1hGk09IyQL
OQ4CLMHaROg2SWWOA5t0Bd78glyI3JjslXNFEQArZCBRGAqychDVagvdTJfqU4ui
A6i1lLYzJoe8jUYylsPQHo7JN3ZeFm2FLOwBoiBtQUNFNcpFIdxJ073NJhx/kkp2
/dQLXUX9/H6Mv4R6C+4gb6lmYBdulBUv0+DT+b2s9YirHG7mPYDHtIqlbJqm7T56
VKxEWFhhX0nPW/wUrAmkNI0apTb5ixbEXXVs1SsdNw1nTQe4QN+kifEQxP5gyUGl
E/jEA450D9rsEC/YDBJ2eDhGARkoozTpx6VbHVbpm092zj7DDR1awr9PcGwYkaor
hRfQv/BeXSWdq7s5h3e5qDWYH7axpHJjg3yJJ/WcJIm0XSAhOejuNCZ37NGoaSh3
c9zhT+idw20I7JQrFiWvtKpufiXkRV3mYpI/TukL//9ZKLwXcPqJmb89h1GMLdV0
UdtpiC1KCz4O5who4sJ4cO4k6p90qGFUj8HQom8miscHRyD56e/zYgnlV9NNdqcj
j97j8nvbPfpOpebHWDAEoRjqgTIA0GYwXZeOChbhGXAzMA35/CI7kjP4jS2IUvE4
icyeKOsMpEMs5cit0hJr+zCstDGZi2xVDGt9r7nSsjKQNvSekfYBZICV9geUcZAe
hBIyirThHm9NxroCMiqLcnAaqXzDqJ7AiBj4YTBbNDTpfuan8TnWkyaPB/WQNpFC
HHkERyP/aY8looku1I9uAbgL40zph8FCwcucPaDuLEaE1FiXm6WRjNCUET7jVV47
UcMNe8SnmM8jMSzaMqn7+j9vVRsBolvcw65LQCXmvMRgSwFq9NW0M7pjaiwNk+1k
xPod0PwujIxpfxOozwGmDbD1hTGVWDUJYmgT4gKeX9CdrHw0vDtPTc77clA9T0lF
a6uygW4j4R2Ra1ebqjwxZkYpx6W/m9/lkftVu9FPSwqI6PRCFwIpk9nIu8JinmlV
uKKZgco0dKNU0kkJVhH9KS8EUp34/waUKlSuMO0TMQSDIq5OZB14la8a35u5TnoI
Tl+Gmsr/ZoRrIc5CB32pP3WqpFUCgXC3xafB9H497u7Rf2l+zhcNKwPcQA6JjpEO
bq/FMYnoqbSQPG1WGArPgCt7lXPX6Apt/nF2UazD6/ahc5V/2H5bKe8eyU7v90Dh
9DtJxF/UxJ+GwMapsrEnx0cdZEdLBbRuU7VwO57gNgbmT7PkQpryvz4al4Yc9JKX
xtFahVeogkkv2DMvRxqNIlAlGugpNsV6UQR1dtvJPRrmjvPcvRcAlsdMH58pNByR
gXs2ADnT8EdG2xpi4asNPYJM0UO2A24twCR6wVmWYtl1JDfs+gQJ5o0IoBAbKYmp
GTRY9S/Ut0VUqM3r+r0Qd5VgmAtRbSDob+i++YdEM9QH+EMTQ5v0YEjzNq6v8VoV
k49zaCL07lZozv+VDo8rZ9k2CIktOs1IggLmWfcYqXfgrP/VV8jCi7I7eQxR+P+q
j7KEiAbrgcenwkovWnitaS+AqhqoWWdr23MLAkOpRKTipk0088bgEERPFYUaN37h
af4KxVPKC4bFtG8P23Wnqt6sdT4eRXZ9J9+nAx6AnJE7Gq6F+543kNmmQ+8cpI9j
bLBXlbhZd+HtZ0k09/4z2gYUoTika3c4BtGm4EazDA8ft+UQhRxaD0III+7Y+4x2
3Gc4ZONi/UcG6lHRqlJzHszz3RpSmCSI3OgCW8hyfGqz/ZoXcT5QeBLG+AkE1Hbl
d5TniEuqJDGUOBAj+lhrYNdoXKS666WLef5htehBAXzwt9+4pUBvZ2VMiGCovUq9
P81O7uf0Tu6e7pR1E87FaZ3PhsXrC5boeNq0FUyp4Tr6VNCEUi2t7FMfjZIdEcKM
o3gEzEE3yIm0O/GYTZZ885dF0HuhVghENcdta3+r+rAebwiOsPt4rarDrsyhtGmH
4FGNmAi8F0Z4dD/Rg0iTT4ydBjUr7dQk3T7nhSqENt66qT4T3WN/uIgkgsyYnpme
GLKvuZtULF2QkUzAiz2F7vkj8NlXHqNAgjYzUPq1HaIdT/Zq4+8BiefBNOZs0vOf
CiEVdvR11uvZKWoPloKSbicwA2oOuaJPXBcHidMmIyycvfQt5dkgR4OWtay7b/aJ
Z19+QpKbAC+f3Fo3j3GvGTm56cKrxQLKV1CsrX//aAB/5sc8Q3r3pkt2MPZIGBV+
WK76YlGGzXVtgO70/Srf1TYBGKWCwxTrwU6c17hquMzhzdpoa+1pTc3Rc0EuNLmq
aXhhZ6+8ZnzP+ctWY8m2HxshDy2EHfZp2Yx4yHyf1mWNkh8r84EKj08ub1xUr599
JlJSkegt1KXSw0ulgBduA5Up3pYl72iFiYuFenN5MO3Cdl9rHKXEps8hLP3SHRXL
nmbOqi5Krs3h5SjiKXRRDxLdGPE7KqJrJjmItB0vugrJVL7SxnWEZ/Kmg/toA/qn
O0ciZpKrx0APFE1bzS6aqBxw0g1oXKBbin0fbIcsTLYDFe/nvKPU+ViVafg/tgzH
dLgjvHpURpzpkyXTTKxopA==
`pragma protect end_protected
